
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixcEcmHoldOtb ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire fclk;
wire uclk;
`_2_ wire holdEcm;
`_2_ wire [63:0] ecmTs;
`_2_ wire [63:0] ecmTsP;
`_2_ wire [255:0] ctrlR;
`_2_ wire [255:0] ctrlW;
`_2_ wire ctrlEv;
`_2_ wire ctrlEvP;
`_2_ wire newCtrl;
`_2_ wire [7:0] cmdC;
`_2_ wire [7:0] cmdCnt;
`_2_ wire [7:0] cmdCntP;
`_2_ wire [63:0] cRet;
`_2_ wire newCmd;
`_2_ wire busyOn;
`_2_ wire [7:0] busyCnt;
wire [0:0] _zyL831_meState0;
supply1 n370;
supply0 n532;
Q_BUF U0 ( .A(ctrlR[136]), .Z(ctrlEv));
Q_BUF U1 ( .A(cmdC[0]), .Z(holdEcm));
Q_BUF U2 ( .A(ecmTs[63]), .Z(ctrlW[127]));
Q_BUF U3 ( .A(ecmTs[62]), .Z(ctrlW[126]));
Q_BUF U4 ( .A(ecmTs[61]), .Z(ctrlW[125]));
Q_BUF U5 ( .A(ecmTs[60]), .Z(ctrlW[124]));
Q_BUF U6 ( .A(ecmTs[59]), .Z(ctrlW[123]));
Q_BUF U7 ( .A(ecmTs[58]), .Z(ctrlW[122]));
Q_BUF U8 ( .A(ecmTs[57]), .Z(ctrlW[121]));
Q_BUF U9 ( .A(ecmTs[56]), .Z(ctrlW[120]));
Q_BUF U10 ( .A(ecmTs[55]), .Z(ctrlW[119]));
Q_BUF U11 ( .A(ecmTs[54]), .Z(ctrlW[118]));
Q_BUF U12 ( .A(ecmTs[53]), .Z(ctrlW[117]));
Q_BUF U13 ( .A(ecmTs[52]), .Z(ctrlW[116]));
Q_BUF U14 ( .A(ecmTs[51]), .Z(ctrlW[115]));
Q_BUF U15 ( .A(ecmTs[50]), .Z(ctrlW[114]));
Q_BUF U16 ( .A(ecmTs[49]), .Z(ctrlW[113]));
Q_BUF U17 ( .A(ecmTs[48]), .Z(ctrlW[112]));
Q_BUF U18 ( .A(ecmTs[47]), .Z(ctrlW[111]));
Q_BUF U19 ( .A(ecmTs[46]), .Z(ctrlW[110]));
Q_BUF U20 ( .A(ecmTs[45]), .Z(ctrlW[109]));
Q_BUF U21 ( .A(ecmTs[44]), .Z(ctrlW[108]));
Q_BUF U22 ( .A(ecmTs[43]), .Z(ctrlW[107]));
Q_BUF U23 ( .A(ecmTs[42]), .Z(ctrlW[106]));
Q_BUF U24 ( .A(ecmTs[41]), .Z(ctrlW[105]));
Q_BUF U25 ( .A(ecmTs[40]), .Z(ctrlW[104]));
Q_BUF U26 ( .A(ecmTs[39]), .Z(ctrlW[103]));
Q_BUF U27 ( .A(ecmTs[38]), .Z(ctrlW[102]));
Q_BUF U28 ( .A(ecmTs[37]), .Z(ctrlW[101]));
Q_BUF U29 ( .A(ecmTs[36]), .Z(ctrlW[100]));
Q_BUF U30 ( .A(ecmTs[35]), .Z(ctrlW[99]));
Q_BUF U31 ( .A(ecmTs[34]), .Z(ctrlW[98]));
Q_BUF U32 ( .A(ecmTs[33]), .Z(ctrlW[97]));
Q_BUF U33 ( .A(ecmTs[32]), .Z(ctrlW[96]));
Q_BUF U34 ( .A(ecmTs[31]), .Z(ctrlW[95]));
Q_BUF U35 ( .A(ecmTs[30]), .Z(ctrlW[94]));
Q_BUF U36 ( .A(ecmTs[29]), .Z(ctrlW[93]));
Q_BUF U37 ( .A(ecmTs[28]), .Z(ctrlW[92]));
Q_BUF U38 ( .A(ecmTs[27]), .Z(ctrlW[91]));
Q_BUF U39 ( .A(ecmTs[26]), .Z(ctrlW[90]));
Q_BUF U40 ( .A(ecmTs[25]), .Z(ctrlW[89]));
Q_BUF U41 ( .A(ecmTs[24]), .Z(ctrlW[88]));
Q_BUF U42 ( .A(ecmTs[23]), .Z(ctrlW[87]));
Q_BUF U43 ( .A(ecmTs[22]), .Z(ctrlW[86]));
Q_BUF U44 ( .A(ecmTs[21]), .Z(ctrlW[85]));
Q_BUF U45 ( .A(ecmTs[20]), .Z(ctrlW[84]));
Q_BUF U46 ( .A(ecmTs[19]), .Z(ctrlW[83]));
Q_BUF U47 ( .A(ecmTs[18]), .Z(ctrlW[82]));
Q_BUF U48 ( .A(ecmTs[17]), .Z(ctrlW[81]));
Q_BUF U49 ( .A(ecmTs[16]), .Z(ctrlW[80]));
Q_BUF U50 ( .A(ecmTs[15]), .Z(ctrlW[79]));
Q_BUF U51 ( .A(ecmTs[14]), .Z(ctrlW[78]));
Q_BUF U52 ( .A(ecmTs[13]), .Z(ctrlW[77]));
Q_BUF U53 ( .A(ecmTs[12]), .Z(ctrlW[76]));
Q_BUF U54 ( .A(ecmTs[11]), .Z(ctrlW[75]));
Q_BUF U55 ( .A(ecmTs[10]), .Z(ctrlW[74]));
Q_BUF U56 ( .A(ecmTs[9]), .Z(ctrlW[73]));
Q_BUF U57 ( .A(ecmTs[8]), .Z(ctrlW[72]));
Q_BUF U58 ( .A(ecmTs[7]), .Z(ctrlW[71]));
Q_BUF U59 ( .A(ecmTs[6]), .Z(ctrlW[70]));
Q_BUF U60 ( .A(ecmTs[5]), .Z(ctrlW[69]));
Q_BUF U61 ( .A(ecmTs[4]), .Z(ctrlW[68]));
Q_BUF U62 ( .A(ecmTs[3]), .Z(ctrlW[67]));
Q_BUF U63 ( .A(ecmTs[2]), .Z(ctrlW[66]));
Q_BUF U64 ( .A(ecmTs[1]), .Z(ctrlW[65]));
Q_BUF U65 ( .A(ecmTs[0]), .Z(ctrlW[64]));
Q_ASSIGN U66 ( .B(xcva_top.xc_top.simTime[63]), .A(ctrlW[191]));
Q_ASSIGN U67 ( .B(xcva_top.xc_top.simTime[62]), .A(ctrlW[190]));
Q_ASSIGN U68 ( .B(xcva_top.xc_top.simTime[61]), .A(ctrlW[189]));
Q_ASSIGN U69 ( .B(xcva_top.xc_top.simTime[60]), .A(ctrlW[188]));
Q_ASSIGN U70 ( .B(xcva_top.xc_top.simTime[59]), .A(ctrlW[187]));
Q_ASSIGN U71 ( .B(xcva_top.xc_top.simTime[58]), .A(ctrlW[186]));
Q_ASSIGN U72 ( .B(xcva_top.xc_top.simTime[57]), .A(ctrlW[185]));
Q_ASSIGN U73 ( .B(xcva_top.xc_top.simTime[56]), .A(ctrlW[184]));
Q_ASSIGN U74 ( .B(xcva_top.xc_top.simTime[55]), .A(ctrlW[183]));
Q_ASSIGN U75 ( .B(xcva_top.xc_top.simTime[54]), .A(ctrlW[182]));
Q_ASSIGN U76 ( .B(xcva_top.xc_top.simTime[53]), .A(ctrlW[181]));
Q_ASSIGN U77 ( .B(xcva_top.xc_top.simTime[52]), .A(ctrlW[180]));
Q_ASSIGN U78 ( .B(xcva_top.xc_top.simTime[51]), .A(ctrlW[179]));
Q_ASSIGN U79 ( .B(xcva_top.xc_top.simTime[50]), .A(ctrlW[178]));
Q_ASSIGN U80 ( .B(xcva_top.xc_top.simTime[49]), .A(ctrlW[177]));
Q_ASSIGN U81 ( .B(xcva_top.xc_top.simTime[48]), .A(ctrlW[176]));
Q_ASSIGN U82 ( .B(xcva_top.xc_top.simTime[47]), .A(ctrlW[175]));
Q_ASSIGN U83 ( .B(xcva_top.xc_top.simTime[46]), .A(ctrlW[174]));
Q_ASSIGN U84 ( .B(xcva_top.xc_top.simTime[45]), .A(ctrlW[173]));
Q_ASSIGN U85 ( .B(xcva_top.xc_top.simTime[44]), .A(ctrlW[172]));
Q_ASSIGN U86 ( .B(xcva_top.xc_top.simTime[43]), .A(ctrlW[171]));
Q_ASSIGN U87 ( .B(xcva_top.xc_top.simTime[42]), .A(ctrlW[170]));
Q_ASSIGN U88 ( .B(xcva_top.xc_top.simTime[41]), .A(ctrlW[169]));
Q_ASSIGN U89 ( .B(xcva_top.xc_top.simTime[40]), .A(ctrlW[168]));
Q_ASSIGN U90 ( .B(xcva_top.xc_top.simTime[39]), .A(ctrlW[167]));
Q_ASSIGN U91 ( .B(xcva_top.xc_top.simTime[38]), .A(ctrlW[166]));
Q_ASSIGN U92 ( .B(xcva_top.xc_top.simTime[37]), .A(ctrlW[165]));
Q_ASSIGN U93 ( .B(xcva_top.xc_top.simTime[36]), .A(ctrlW[164]));
Q_ASSIGN U94 ( .B(xcva_top.xc_top.simTime[35]), .A(ctrlW[163]));
Q_ASSIGN U95 ( .B(xcva_top.xc_top.simTime[34]), .A(ctrlW[162]));
Q_ASSIGN U96 ( .B(xcva_top.xc_top.simTime[33]), .A(ctrlW[161]));
Q_ASSIGN U97 ( .B(xcva_top.xc_top.simTime[32]), .A(ctrlW[160]));
Q_ASSIGN U98 ( .B(xcva_top.xc_top.simTime[31]), .A(ctrlW[159]));
Q_ASSIGN U99 ( .B(xcva_top.xc_top.simTime[30]), .A(ctrlW[158]));
Q_ASSIGN U100 ( .B(xcva_top.xc_top.simTime[29]), .A(ctrlW[157]));
Q_ASSIGN U101 ( .B(xcva_top.xc_top.simTime[28]), .A(ctrlW[156]));
Q_ASSIGN U102 ( .B(xcva_top.xc_top.simTime[27]), .A(ctrlW[155]));
Q_ASSIGN U103 ( .B(xcva_top.xc_top.simTime[26]), .A(ctrlW[154]));
Q_ASSIGN U104 ( .B(xcva_top.xc_top.simTime[25]), .A(ctrlW[153]));
Q_ASSIGN U105 ( .B(xcva_top.xc_top.simTime[24]), .A(ctrlW[152]));
Q_ASSIGN U106 ( .B(xcva_top.xc_top.simTime[23]), .A(ctrlW[151]));
Q_ASSIGN U107 ( .B(xcva_top.xc_top.simTime[22]), .A(ctrlW[150]));
Q_ASSIGN U108 ( .B(xcva_top.xc_top.simTime[21]), .A(ctrlW[149]));
Q_ASSIGN U109 ( .B(xcva_top.xc_top.simTime[20]), .A(ctrlW[148]));
Q_ASSIGN U110 ( .B(xcva_top.xc_top.simTime[19]), .A(ctrlW[147]));
Q_ASSIGN U111 ( .B(xcva_top.xc_top.simTime[18]), .A(ctrlW[146]));
Q_ASSIGN U112 ( .B(xcva_top.xc_top.simTime[17]), .A(ctrlW[145]));
Q_ASSIGN U113 ( .B(xcva_top.xc_top.simTime[16]), .A(ctrlW[144]));
Q_ASSIGN U114 ( .B(xcva_top.xc_top.simTime[15]), .A(ctrlW[143]));
Q_ASSIGN U115 ( .B(xcva_top.xc_top.simTime[14]), .A(ctrlW[142]));
Q_ASSIGN U116 ( .B(xcva_top.xc_top.simTime[13]), .A(ctrlW[141]));
Q_ASSIGN U117 ( .B(xcva_top.xc_top.simTime[12]), .A(ctrlW[140]));
Q_ASSIGN U118 ( .B(xcva_top.xc_top.simTime[11]), .A(ctrlW[139]));
Q_ASSIGN U119 ( .B(xcva_top.xc_top.simTime[10]), .A(ctrlW[138]));
Q_ASSIGN U120 ( .B(xcva_top.xc_top.simTime[9]), .A(ctrlW[137]));
Q_ASSIGN U121 ( .B(xcva_top.xc_top.simTime[8]), .A(ctrlW[136]));
Q_ASSIGN U122 ( .B(xcva_top.xc_top.simTime[7]), .A(ctrlW[135]));
Q_ASSIGN U123 ( .B(xcva_top.xc_top.simTime[6]), .A(ctrlW[134]));
Q_ASSIGN U124 ( .B(xcva_top.xc_top.simTime[5]), .A(ctrlW[133]));
Q_ASSIGN U125 ( .B(xcva_top.xc_top.simTime[4]), .A(ctrlW[132]));
Q_ASSIGN U126 ( .B(xcva_top.xc_top.simTime[3]), .A(ctrlW[131]));
Q_ASSIGN U127 ( .B(xcva_top.xc_top.simTime[2]), .A(ctrlW[130]));
Q_ASSIGN U128 ( .B(xcva_top.xc_top.simTime[1]), .A(ctrlW[129]));
Q_ASSIGN U129 ( .B(xcva_top.xc_top.simTime[0]), .A(ctrlW[128]));
Q_ASSIGN U130 ( .B(cRet[63]), .A(ctrlW[63]));
Q_ASSIGN U131 ( .B(cRet[62]), .A(ctrlW[62]));
Q_ASSIGN U132 ( .B(cRet[61]), .A(ctrlW[61]));
Q_ASSIGN U133 ( .B(cRet[60]), .A(ctrlW[60]));
Q_ASSIGN U134 ( .B(cRet[59]), .A(ctrlW[59]));
Q_ASSIGN U135 ( .B(cRet[58]), .A(ctrlW[58]));
Q_ASSIGN U136 ( .B(cRet[57]), .A(ctrlW[57]));
Q_ASSIGN U137 ( .B(cRet[56]), .A(ctrlW[56]));
Q_ASSIGN U138 ( .B(cRet[55]), .A(ctrlW[55]));
Q_ASSIGN U139 ( .B(cRet[54]), .A(ctrlW[54]));
Q_ASSIGN U140 ( .B(cRet[53]), .A(ctrlW[53]));
Q_ASSIGN U141 ( .B(cRet[52]), .A(ctrlW[52]));
Q_ASSIGN U142 ( .B(cRet[51]), .A(ctrlW[51]));
Q_ASSIGN U143 ( .B(cRet[50]), .A(ctrlW[50]));
Q_ASSIGN U144 ( .B(cRet[49]), .A(ctrlW[49]));
Q_ASSIGN U145 ( .B(cRet[48]), .A(ctrlW[48]));
Q_ASSIGN U146 ( .B(cRet[47]), .A(ctrlW[47]));
Q_ASSIGN U147 ( .B(cRet[46]), .A(ctrlW[46]));
Q_ASSIGN U148 ( .B(cRet[45]), .A(ctrlW[45]));
Q_ASSIGN U149 ( .B(cRet[44]), .A(ctrlW[44]));
Q_ASSIGN U150 ( .B(cRet[43]), .A(ctrlW[43]));
Q_ASSIGN U151 ( .B(cRet[42]), .A(ctrlW[42]));
Q_ASSIGN U152 ( .B(cRet[41]), .A(ctrlW[41]));
Q_ASSIGN U153 ( .B(cRet[40]), .A(ctrlW[40]));
Q_ASSIGN U154 ( .B(cRet[39]), .A(ctrlW[39]));
Q_ASSIGN U155 ( .B(cRet[38]), .A(ctrlW[38]));
Q_ASSIGN U156 ( .B(cRet[37]), .A(ctrlW[37]));
Q_ASSIGN U157 ( .B(cRet[36]), .A(ctrlW[36]));
Q_ASSIGN U158 ( .B(cRet[35]), .A(ctrlW[35]));
Q_ASSIGN U159 ( .B(cRet[34]), .A(ctrlW[34]));
Q_ASSIGN U160 ( .B(cRet[33]), .A(ctrlW[33]));
Q_ASSIGN U161 ( .B(cRet[32]), .A(ctrlW[32]));
Q_ASSIGN U162 ( .B(cRet[31]), .A(ctrlW[31]));
Q_ASSIGN U163 ( .B(cRet[30]), .A(ctrlW[30]));
Q_ASSIGN U164 ( .B(cRet[29]), .A(ctrlW[29]));
Q_ASSIGN U165 ( .B(cRet[28]), .A(ctrlW[28]));
Q_ASSIGN U166 ( .B(cRet[27]), .A(ctrlW[27]));
Q_ASSIGN U167 ( .B(cRet[26]), .A(ctrlW[26]));
Q_ASSIGN U168 ( .B(cRet[25]), .A(ctrlW[25]));
Q_ASSIGN U169 ( .B(cRet[24]), .A(ctrlW[24]));
Q_ASSIGN U170 ( .B(cRet[23]), .A(ctrlW[23]));
Q_ASSIGN U171 ( .B(cRet[22]), .A(ctrlW[22]));
Q_ASSIGN U172 ( .B(cRet[21]), .A(ctrlW[21]));
Q_ASSIGN U173 ( .B(cRet[20]), .A(ctrlW[20]));
Q_ASSIGN U174 ( .B(cRet[19]), .A(ctrlW[19]));
Q_ASSIGN U175 ( .B(cRet[18]), .A(ctrlW[18]));
Q_ASSIGN U176 ( .B(cRet[17]), .A(ctrlW[17]));
Q_ASSIGN U177 ( .B(cRet[16]), .A(ctrlW[16]));
Q_BUF U178 ( .A(cRet[15]), .Z(ctrlW[15]));
Q_BUF U179 ( .A(cRet[14]), .Z(ctrlW[14]));
Q_BUF U180 ( .A(cRet[13]), .Z(ctrlW[13]));
Q_BUF U181 ( .A(cRet[12]), .Z(ctrlW[12]));
Q_BUF U182 ( .A(cRet[11]), .Z(ctrlW[11]));
Q_BUF U183 ( .A(cRet[10]), .Z(ctrlW[10]));
Q_BUF U184 ( .A(cRet[9]), .Z(ctrlW[9]));
Q_BUF U185 ( .A(cRet[8]), .Z(ctrlW[8]));
Q_ASSIGN U186 ( .B(cRet[7]), .A(ctrlW[7]));
Q_ASSIGN U187 ( .B(cRet[6]), .A(ctrlW[6]));
Q_ASSIGN U188 ( .B(cRet[5]), .A(ctrlW[5]));
Q_ASSIGN U189 ( .B(cRet[4]), .A(ctrlW[4]));
Q_ASSIGN U190 ( .B(cRet[3]), .A(ctrlW[3]));
Q_BUF U191 ( .A(cRet[2]), .Z(ctrlW[2]));
Q_BUF U192 ( .A(cRet[1]), .Z(ctrlW[1]));
Q_BUF U193 ( .A(cRet[0]), .Z(ctrlW[0]));
Q_AN02 U194 ( .A0(n531), .A1(xcva_top.xc_top.ecmOnD), .Z(n791));
ixc_uClkGen ukg ( uclk);
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_BUFZP U197 ( .OE(holdEcm), .A(n370), .Z(xcva_top.xc_top.holdEcmTb));
Q_BUFZP U198 ( .OE(busyOn), .A(n370), .Z(xcva_top.xc_top.ecmHoldBusy));
Q_FDP0 \ctrlR_REG[0] ( .CK(uclk), .D(n533), .Q(ctrlR[0]), .QN( ));
Q_FDP0 \ctrlR_REG[1] ( .CK(uclk), .D(n534), .Q(ctrlR[1]), .QN( ));
Q_FDP0 \ctrlR_REG[2] ( .CK(uclk), .D(n535), .Q(ctrlR[2]), .QN( ));
Q_FDP0 \ctrlR_REG[3] ( .CK(uclk), .D(n536), .Q(ctrlR[3]), .QN( ));
Q_FDP0 \ctrlR_REG[4] ( .CK(uclk), .D(n537), .Q(ctrlR[4]), .QN( ));
Q_FDP0 \ctrlR_REG[5] ( .CK(uclk), .D(n538), .Q(ctrlR[5]), .QN( ));
Q_FDP0 \ctrlR_REG[6] ( .CK(uclk), .D(n539), .Q(ctrlR[6]), .QN( ));
Q_FDP0 \ctrlR_REG[7] ( .CK(uclk), .D(n540), .Q(ctrlR[7]), .QN( ));
Q_FDP0 \ctrlR_REG[8] ( .CK(uclk), .D(n541), .Q(ctrlR[8]), .QN( ));
Q_FDP0 \ctrlR_REG[9] ( .CK(uclk), .D(n542), .Q(ctrlR[9]), .QN( ));
Q_FDP0 \ctrlR_REG[10] ( .CK(uclk), .D(n543), .Q(ctrlR[10]), .QN( ));
Q_FDP0 \ctrlR_REG[11] ( .CK(uclk), .D(n544), .Q(ctrlR[11]), .QN( ));
Q_FDP0 \ctrlR_REG[12] ( .CK(uclk), .D(n545), .Q(ctrlR[12]), .QN( ));
Q_FDP0 \ctrlR_REG[13] ( .CK(uclk), .D(n546), .Q(ctrlR[13]), .QN( ));
Q_FDP0 \ctrlR_REG[14] ( .CK(uclk), .D(n547), .Q(ctrlR[14]), .QN( ));
Q_FDP0 \ctrlR_REG[15] ( .CK(uclk), .D(n548), .Q(ctrlR[15]), .QN( ));
Q_FDP0 \ctrlR_REG[16] ( .CK(uclk), .D(n549), .Q(ctrlR[16]), .QN( ));
Q_FDP0 \ctrlR_REG[17] ( .CK(uclk), .D(n550), .Q(ctrlR[17]), .QN( ));
Q_FDP0 \ctrlR_REG[18] ( .CK(uclk), .D(n551), .Q(ctrlR[18]), .QN( ));
Q_FDP0 \ctrlR_REG[19] ( .CK(uclk), .D(n552), .Q(ctrlR[19]), .QN( ));
Q_FDP0 \ctrlR_REG[20] ( .CK(uclk), .D(n553), .Q(ctrlR[20]), .QN( ));
Q_FDP0 \ctrlR_REG[21] ( .CK(uclk), .D(n554), .Q(ctrlR[21]), .QN( ));
Q_FDP0 \ctrlR_REG[22] ( .CK(uclk), .D(n555), .Q(ctrlR[22]), .QN( ));
Q_FDP0 \ctrlR_REG[23] ( .CK(uclk), .D(n556), .Q(ctrlR[23]), .QN( ));
Q_FDP0 \ctrlR_REG[24] ( .CK(uclk), .D(n557), .Q(ctrlR[24]), .QN( ));
Q_FDP0 \ctrlR_REG[25] ( .CK(uclk), .D(n558), .Q(ctrlR[25]), .QN( ));
Q_FDP0 \ctrlR_REG[26] ( .CK(uclk), .D(n559), .Q(ctrlR[26]), .QN( ));
Q_FDP0 \ctrlR_REG[27] ( .CK(uclk), .D(n560), .Q(ctrlR[27]), .QN( ));
Q_FDP0 \ctrlR_REG[28] ( .CK(uclk), .D(n561), .Q(ctrlR[28]), .QN( ));
Q_FDP0 \ctrlR_REG[29] ( .CK(uclk), .D(n562), .Q(ctrlR[29]), .QN( ));
Q_FDP0 \ctrlR_REG[30] ( .CK(uclk), .D(n563), .Q(ctrlR[30]), .QN( ));
Q_FDP0 \ctrlR_REG[31] ( .CK(uclk), .D(n564), .Q(ctrlR[31]), .QN( ));
Q_FDP0 \ctrlR_REG[32] ( .CK(uclk), .D(n565), .Q(ctrlR[32]), .QN( ));
Q_FDP0 \ctrlR_REG[33] ( .CK(uclk), .D(n566), .Q(ctrlR[33]), .QN( ));
Q_FDP0 \ctrlR_REG[34] ( .CK(uclk), .D(n567), .Q(ctrlR[34]), .QN( ));
Q_FDP0 \ctrlR_REG[35] ( .CK(uclk), .D(n568), .Q(ctrlR[35]), .QN( ));
Q_FDP0 \ctrlR_REG[36] ( .CK(uclk), .D(n569), .Q(ctrlR[36]), .QN( ));
Q_FDP0 \ctrlR_REG[37] ( .CK(uclk), .D(n570), .Q(ctrlR[37]), .QN( ));
Q_FDP0 \ctrlR_REG[38] ( .CK(uclk), .D(n571), .Q(ctrlR[38]), .QN( ));
Q_FDP0 \ctrlR_REG[39] ( .CK(uclk), .D(n572), .Q(ctrlR[39]), .QN( ));
Q_FDP0 \ctrlR_REG[40] ( .CK(uclk), .D(n573), .Q(ctrlR[40]), .QN( ));
Q_FDP0 \ctrlR_REG[41] ( .CK(uclk), .D(n574), .Q(ctrlR[41]), .QN( ));
Q_FDP0 \ctrlR_REG[42] ( .CK(uclk), .D(n575), .Q(ctrlR[42]), .QN( ));
Q_FDP0 \ctrlR_REG[43] ( .CK(uclk), .D(n576), .Q(ctrlR[43]), .QN( ));
Q_FDP0 \ctrlR_REG[44] ( .CK(uclk), .D(n577), .Q(ctrlR[44]), .QN( ));
Q_FDP0 \ctrlR_REG[45] ( .CK(uclk), .D(n578), .Q(ctrlR[45]), .QN( ));
Q_FDP0 \ctrlR_REG[46] ( .CK(uclk), .D(n579), .Q(ctrlR[46]), .QN( ));
Q_FDP0 \ctrlR_REG[47] ( .CK(uclk), .D(n580), .Q(ctrlR[47]), .QN( ));
Q_FDP0 \ctrlR_REG[48] ( .CK(uclk), .D(n581), .Q(ctrlR[48]), .QN( ));
Q_FDP0 \ctrlR_REG[49] ( .CK(uclk), .D(n582), .Q(ctrlR[49]), .QN( ));
Q_FDP0 \ctrlR_REG[50] ( .CK(uclk), .D(n583), .Q(ctrlR[50]), .QN( ));
Q_FDP0 \ctrlR_REG[51] ( .CK(uclk), .D(n584), .Q(ctrlR[51]), .QN( ));
Q_FDP0 \ctrlR_REG[52] ( .CK(uclk), .D(n585), .Q(ctrlR[52]), .QN( ));
Q_FDP0 \ctrlR_REG[53] ( .CK(uclk), .D(n586), .Q(ctrlR[53]), .QN( ));
Q_FDP0 \ctrlR_REG[54] ( .CK(uclk), .D(n587), .Q(ctrlR[54]), .QN( ));
Q_FDP0 \ctrlR_REG[55] ( .CK(uclk), .D(n588), .Q(ctrlR[55]), .QN( ));
Q_FDP0 \ctrlR_REG[56] ( .CK(uclk), .D(n589), .Q(ctrlR[56]), .QN( ));
Q_FDP0 \ctrlR_REG[57] ( .CK(uclk), .D(n590), .Q(ctrlR[57]), .QN( ));
Q_FDP0 \ctrlR_REG[58] ( .CK(uclk), .D(n591), .Q(ctrlR[58]), .QN( ));
Q_FDP0 \ctrlR_REG[59] ( .CK(uclk), .D(n592), .Q(ctrlR[59]), .QN( ));
Q_FDP0 \ctrlR_REG[60] ( .CK(uclk), .D(n593), .Q(ctrlR[60]), .QN( ));
Q_FDP0 \ctrlR_REG[61] ( .CK(uclk), .D(n594), .Q(ctrlR[61]), .QN( ));
Q_FDP0 \ctrlR_REG[62] ( .CK(uclk), .D(n595), .Q(ctrlR[62]), .QN( ));
Q_FDP0 \ctrlR_REG[63] ( .CK(uclk), .D(n596), .Q(ctrlR[63]), .QN( ));
Q_FDP0 \ctrlR_REG[64] ( .CK(uclk), .D(n597), .Q(ctrlR[64]), .QN( ));
Q_FDP0 \ctrlR_REG[65] ( .CK(uclk), .D(n598), .Q(ctrlR[65]), .QN( ));
Q_FDP0 \ctrlR_REG[66] ( .CK(uclk), .D(n599), .Q(ctrlR[66]), .QN( ));
Q_FDP0 \ctrlR_REG[67] ( .CK(uclk), .D(n600), .Q(ctrlR[67]), .QN( ));
Q_FDP0 \ctrlR_REG[68] ( .CK(uclk), .D(n601), .Q(ctrlR[68]), .QN( ));
Q_FDP0 \ctrlR_REG[69] ( .CK(uclk), .D(n602), .Q(ctrlR[69]), .QN( ));
Q_FDP0 \ctrlR_REG[70] ( .CK(uclk), .D(n603), .Q(ctrlR[70]), .QN( ));
Q_FDP0 \ctrlR_REG[71] ( .CK(uclk), .D(n604), .Q(ctrlR[71]), .QN( ));
Q_FDP0 \ctrlR_REG[72] ( .CK(uclk), .D(n605), .Q(ctrlR[72]), .QN( ));
Q_FDP0 \ctrlR_REG[73] ( .CK(uclk), .D(n606), .Q(ctrlR[73]), .QN( ));
Q_FDP0 \ctrlR_REG[74] ( .CK(uclk), .D(n607), .Q(ctrlR[74]), .QN( ));
Q_FDP0 \ctrlR_REG[75] ( .CK(uclk), .D(n608), .Q(ctrlR[75]), .QN( ));
Q_FDP0 \ctrlR_REG[76] ( .CK(uclk), .D(n609), .Q(ctrlR[76]), .QN( ));
Q_FDP0 \ctrlR_REG[77] ( .CK(uclk), .D(n610), .Q(ctrlR[77]), .QN( ));
Q_FDP0 \ctrlR_REG[78] ( .CK(uclk), .D(n611), .Q(ctrlR[78]), .QN( ));
Q_FDP0 \ctrlR_REG[79] ( .CK(uclk), .D(n612), .Q(ctrlR[79]), .QN( ));
Q_FDP0 \ctrlR_REG[80] ( .CK(uclk), .D(n613), .Q(ctrlR[80]), .QN( ));
Q_FDP0 \ctrlR_REG[81] ( .CK(uclk), .D(n614), .Q(ctrlR[81]), .QN( ));
Q_FDP0 \ctrlR_REG[82] ( .CK(uclk), .D(n615), .Q(ctrlR[82]), .QN( ));
Q_FDP0 \ctrlR_REG[83] ( .CK(uclk), .D(n616), .Q(ctrlR[83]), .QN( ));
Q_FDP0 \ctrlR_REG[84] ( .CK(uclk), .D(n617), .Q(ctrlR[84]), .QN( ));
Q_FDP0 \ctrlR_REG[85] ( .CK(uclk), .D(n618), .Q(ctrlR[85]), .QN( ));
Q_FDP0 \ctrlR_REG[86] ( .CK(uclk), .D(n619), .Q(ctrlR[86]), .QN( ));
Q_FDP0 \ctrlR_REG[87] ( .CK(uclk), .D(n620), .Q(ctrlR[87]), .QN( ));
Q_FDP0 \ctrlR_REG[88] ( .CK(uclk), .D(n621), .Q(ctrlR[88]), .QN( ));
Q_FDP0 \ctrlR_REG[89] ( .CK(uclk), .D(n622), .Q(ctrlR[89]), .QN( ));
Q_FDP0 \ctrlR_REG[90] ( .CK(uclk), .D(n623), .Q(ctrlR[90]), .QN( ));
Q_FDP0 \ctrlR_REG[91] ( .CK(uclk), .D(n624), .Q(ctrlR[91]), .QN( ));
Q_FDP0 \ctrlR_REG[92] ( .CK(uclk), .D(n625), .Q(ctrlR[92]), .QN( ));
Q_FDP0 \ctrlR_REG[93] ( .CK(uclk), .D(n626), .Q(ctrlR[93]), .QN( ));
Q_FDP0 \ctrlR_REG[94] ( .CK(uclk), .D(n627), .Q(ctrlR[94]), .QN( ));
Q_FDP0 \ctrlR_REG[95] ( .CK(uclk), .D(n628), .Q(ctrlR[95]), .QN( ));
Q_FDP0 \ctrlR_REG[96] ( .CK(uclk), .D(n629), .Q(ctrlR[96]), .QN( ));
Q_FDP0 \ctrlR_REG[97] ( .CK(uclk), .D(n630), .Q(ctrlR[97]), .QN( ));
Q_FDP0 \ctrlR_REG[98] ( .CK(uclk), .D(n631), .Q(ctrlR[98]), .QN( ));
Q_FDP0 \ctrlR_REG[99] ( .CK(uclk), .D(n632), .Q(ctrlR[99]), .QN( ));
Q_FDP0 \ctrlR_REG[100] ( .CK(uclk), .D(n633), .Q(ctrlR[100]), .QN( ));
Q_FDP0 \ctrlR_REG[101] ( .CK(uclk), .D(n634), .Q(ctrlR[101]), .QN( ));
Q_FDP0 \ctrlR_REG[102] ( .CK(uclk), .D(n635), .Q(ctrlR[102]), .QN( ));
Q_FDP0 \ctrlR_REG[103] ( .CK(uclk), .D(n636), .Q(ctrlR[103]), .QN( ));
Q_FDP0 \ctrlR_REG[104] ( .CK(uclk), .D(n637), .Q(ctrlR[104]), .QN( ));
Q_FDP0 \ctrlR_REG[105] ( .CK(uclk), .D(n638), .Q(ctrlR[105]), .QN( ));
Q_FDP0 \ctrlR_REG[106] ( .CK(uclk), .D(n639), .Q(ctrlR[106]), .QN( ));
Q_FDP0 \ctrlR_REG[107] ( .CK(uclk), .D(n640), .Q(ctrlR[107]), .QN( ));
Q_FDP0 \ctrlR_REG[108] ( .CK(uclk), .D(n641), .Q(ctrlR[108]), .QN( ));
Q_FDP0 \ctrlR_REG[109] ( .CK(uclk), .D(n642), .Q(ctrlR[109]), .QN( ));
Q_FDP0 \ctrlR_REG[110] ( .CK(uclk), .D(n643), .Q(ctrlR[110]), .QN( ));
Q_FDP0 \ctrlR_REG[111] ( .CK(uclk), .D(n644), .Q(ctrlR[111]), .QN( ));
Q_FDP0 \ctrlR_REG[112] ( .CK(uclk), .D(n645), .Q(ctrlR[112]), .QN( ));
Q_FDP0 \ctrlR_REG[113] ( .CK(uclk), .D(n646), .Q(ctrlR[113]), .QN( ));
Q_FDP0 \ctrlR_REG[114] ( .CK(uclk), .D(n647), .Q(ctrlR[114]), .QN( ));
Q_FDP0 \ctrlR_REG[115] ( .CK(uclk), .D(n648), .Q(ctrlR[115]), .QN( ));
Q_FDP0 \ctrlR_REG[116] ( .CK(uclk), .D(n649), .Q(ctrlR[116]), .QN( ));
Q_FDP0 \ctrlR_REG[117] ( .CK(uclk), .D(n650), .Q(ctrlR[117]), .QN( ));
Q_FDP0 \ctrlR_REG[118] ( .CK(uclk), .D(n651), .Q(ctrlR[118]), .QN( ));
Q_FDP0 \ctrlR_REG[119] ( .CK(uclk), .D(n652), .Q(ctrlR[119]), .QN( ));
Q_FDP0 \ctrlR_REG[120] ( .CK(uclk), .D(n653), .Q(ctrlR[120]), .QN( ));
Q_FDP0 \ctrlR_REG[121] ( .CK(uclk), .D(n654), .Q(ctrlR[121]), .QN( ));
Q_FDP0 \ctrlR_REG[122] ( .CK(uclk), .D(n655), .Q(ctrlR[122]), .QN( ));
Q_FDP0 \ctrlR_REG[123] ( .CK(uclk), .D(n656), .Q(ctrlR[123]), .QN( ));
Q_FDP0 \ctrlR_REG[124] ( .CK(uclk), .D(n657), .Q(ctrlR[124]), .QN( ));
Q_FDP0 \ctrlR_REG[125] ( .CK(uclk), .D(n658), .Q(ctrlR[125]), .QN( ));
Q_FDP0 \ctrlR_REG[126] ( .CK(uclk), .D(n659), .Q(ctrlR[126]), .QN( ));
Q_FDP0 \ctrlR_REG[127] ( .CK(uclk), .D(n660), .Q(ctrlR[127]), .QN( ));
Q_FDP0 \ctrlR_REG[128] ( .CK(uclk), .D(n661), .Q(ctrlR[128]), .QN( ));
Q_FDP0 \ctrlR_REG[129] ( .CK(uclk), .D(n662), .Q(ctrlR[129]), .QN( ));
Q_FDP0 \ctrlR_REG[130] ( .CK(uclk), .D(n663), .Q(ctrlR[130]), .QN( ));
Q_FDP0 \ctrlR_REG[131] ( .CK(uclk), .D(n664), .Q(ctrlR[131]), .QN( ));
Q_FDP0 \ctrlR_REG[132] ( .CK(uclk), .D(n665), .Q(ctrlR[132]), .QN( ));
Q_FDP0 \ctrlR_REG[133] ( .CK(uclk), .D(n666), .Q(ctrlR[133]), .QN( ));
Q_FDP0 \ctrlR_REG[134] ( .CK(uclk), .D(n667), .Q(ctrlR[134]), .QN( ));
Q_FDP0 \ctrlR_REG[135] ( .CK(uclk), .D(n668), .Q(ctrlR[135]), .QN( ));
Q_FDP0 \ctrlR_REG[136] ( .CK(uclk), .D(n669), .Q(ctrlR[136]), .QN( ));
Q_FDP0 \ctrlR_REG[137] ( .CK(uclk), .D(n670), .Q(ctrlR[137]), .QN( ));
Q_FDP0 \ctrlR_REG[138] ( .CK(uclk), .D(n671), .Q(ctrlR[138]), .QN( ));
Q_FDP0 \ctrlR_REG[139] ( .CK(uclk), .D(n672), .Q(ctrlR[139]), .QN( ));
Q_FDP0 \ctrlR_REG[140] ( .CK(uclk), .D(n673), .Q(ctrlR[140]), .QN( ));
Q_FDP0 \ctrlR_REG[141] ( .CK(uclk), .D(n674), .Q(ctrlR[141]), .QN( ));
Q_FDP0 \ctrlR_REG[142] ( .CK(uclk), .D(n675), .Q(ctrlR[142]), .QN( ));
Q_FDP0 \ctrlR_REG[143] ( .CK(uclk), .D(n676), .Q(ctrlR[143]), .QN( ));
Q_FDP0 \ctrlR_REG[144] ( .CK(uclk), .D(n677), .Q(ctrlR[144]), .QN( ));
Q_FDP0 \ctrlR_REG[145] ( .CK(uclk), .D(n678), .Q(ctrlR[145]), .QN( ));
Q_FDP0 \ctrlR_REG[146] ( .CK(uclk), .D(n679), .Q(ctrlR[146]), .QN( ));
Q_FDP0 \ctrlR_REG[147] ( .CK(uclk), .D(n680), .Q(ctrlR[147]), .QN( ));
Q_FDP0 \ctrlR_REG[148] ( .CK(uclk), .D(n681), .Q(ctrlR[148]), .QN( ));
Q_FDP0 \ctrlR_REG[149] ( .CK(uclk), .D(n682), .Q(ctrlR[149]), .QN( ));
Q_FDP0 \ctrlR_REG[150] ( .CK(uclk), .D(n683), .Q(ctrlR[150]), .QN( ));
Q_FDP0 \ctrlR_REG[151] ( .CK(uclk), .D(n684), .Q(ctrlR[151]), .QN( ));
Q_FDP0 \ctrlR_REG[152] ( .CK(uclk), .D(n685), .Q(ctrlR[152]), .QN( ));
Q_FDP0 \ctrlR_REG[153] ( .CK(uclk), .D(n686), .Q(ctrlR[153]), .QN( ));
Q_FDP0 \ctrlR_REG[154] ( .CK(uclk), .D(n687), .Q(ctrlR[154]), .QN( ));
Q_FDP0 \ctrlR_REG[155] ( .CK(uclk), .D(n688), .Q(ctrlR[155]), .QN( ));
Q_FDP0 \ctrlR_REG[156] ( .CK(uclk), .D(n689), .Q(ctrlR[156]), .QN( ));
Q_FDP0 \ctrlR_REG[157] ( .CK(uclk), .D(n690), .Q(ctrlR[157]), .QN( ));
Q_FDP0 \ctrlR_REG[158] ( .CK(uclk), .D(n691), .Q(ctrlR[158]), .QN( ));
Q_FDP0 \ctrlR_REG[159] ( .CK(uclk), .D(n692), .Q(ctrlR[159]), .QN( ));
Q_FDP0 \ctrlR_REG[160] ( .CK(uclk), .D(n693), .Q(ctrlR[160]), .QN( ));
Q_FDP0 \ctrlR_REG[161] ( .CK(uclk), .D(n694), .Q(ctrlR[161]), .QN( ));
Q_FDP0 \ctrlR_REG[162] ( .CK(uclk), .D(n695), .Q(ctrlR[162]), .QN( ));
Q_FDP0 \ctrlR_REG[163] ( .CK(uclk), .D(n696), .Q(ctrlR[163]), .QN( ));
Q_FDP0 \ctrlR_REG[164] ( .CK(uclk), .D(n697), .Q(ctrlR[164]), .QN( ));
Q_FDP0 \ctrlR_REG[165] ( .CK(uclk), .D(n698), .Q(ctrlR[165]), .QN( ));
Q_FDP0 \ctrlR_REG[166] ( .CK(uclk), .D(n699), .Q(ctrlR[166]), .QN( ));
Q_FDP0 \ctrlR_REG[167] ( .CK(uclk), .D(n700), .Q(ctrlR[167]), .QN( ));
Q_FDP0 \ctrlR_REG[168] ( .CK(uclk), .D(n701), .Q(ctrlR[168]), .QN( ));
Q_FDP0 \ctrlR_REG[169] ( .CK(uclk), .D(n702), .Q(ctrlR[169]), .QN( ));
Q_FDP0 \ctrlR_REG[170] ( .CK(uclk), .D(n703), .Q(ctrlR[170]), .QN( ));
Q_FDP0 \ctrlR_REG[171] ( .CK(uclk), .D(n704), .Q(ctrlR[171]), .QN( ));
Q_FDP0 \ctrlR_REG[172] ( .CK(uclk), .D(n705), .Q(ctrlR[172]), .QN( ));
Q_FDP0 \ctrlR_REG[173] ( .CK(uclk), .D(n706), .Q(ctrlR[173]), .QN( ));
Q_FDP0 \ctrlR_REG[174] ( .CK(uclk), .D(n707), .Q(ctrlR[174]), .QN( ));
Q_FDP0 \ctrlR_REG[175] ( .CK(uclk), .D(n708), .Q(ctrlR[175]), .QN( ));
Q_FDP0 \ctrlR_REG[176] ( .CK(uclk), .D(n709), .Q(ctrlR[176]), .QN( ));
Q_FDP0 \ctrlR_REG[177] ( .CK(uclk), .D(n710), .Q(ctrlR[177]), .QN( ));
Q_FDP0 \ctrlR_REG[178] ( .CK(uclk), .D(n711), .Q(ctrlR[178]), .QN( ));
Q_FDP0 \ctrlR_REG[179] ( .CK(uclk), .D(n712), .Q(ctrlR[179]), .QN( ));
Q_FDP0 \ctrlR_REG[180] ( .CK(uclk), .D(n713), .Q(ctrlR[180]), .QN( ));
Q_FDP0 \ctrlR_REG[181] ( .CK(uclk), .D(n714), .Q(ctrlR[181]), .QN( ));
Q_FDP0 \ctrlR_REG[182] ( .CK(uclk), .D(n715), .Q(ctrlR[182]), .QN( ));
Q_FDP0 \ctrlR_REG[183] ( .CK(uclk), .D(n716), .Q(ctrlR[183]), .QN( ));
Q_FDP0 \ctrlR_REG[184] ( .CK(uclk), .D(n717), .Q(ctrlR[184]), .QN( ));
Q_FDP0 \ctrlR_REG[185] ( .CK(uclk), .D(n718), .Q(ctrlR[185]), .QN( ));
Q_FDP0 \ctrlR_REG[186] ( .CK(uclk), .D(n719), .Q(ctrlR[186]), .QN( ));
Q_FDP0 \ctrlR_REG[187] ( .CK(uclk), .D(n720), .Q(ctrlR[187]), .QN( ));
Q_FDP0 \ctrlR_REG[188] ( .CK(uclk), .D(n721), .Q(ctrlR[188]), .QN( ));
Q_FDP0 \ctrlR_REG[189] ( .CK(uclk), .D(n722), .Q(ctrlR[189]), .QN( ));
Q_FDP0 \ctrlR_REG[190] ( .CK(uclk), .D(n723), .Q(ctrlR[190]), .QN( ));
Q_FDP0 \ctrlR_REG[191] ( .CK(uclk), .D(n724), .Q(ctrlR[191]), .QN( ));
Q_FDP0 \ctrlR_REG[192] ( .CK(uclk), .D(n725), .Q(ctrlR[192]), .QN( ));
Q_FDP0 \ctrlR_REG[193] ( .CK(uclk), .D(n726), .Q(ctrlR[193]), .QN( ));
Q_FDP0 \ctrlR_REG[194] ( .CK(uclk), .D(n727), .Q(ctrlR[194]), .QN( ));
Q_FDP0 \ctrlR_REG[195] ( .CK(uclk), .D(n728), .Q(ctrlR[195]), .QN( ));
Q_FDP0 \ctrlR_REG[196] ( .CK(uclk), .D(n729), .Q(ctrlR[196]), .QN( ));
Q_FDP0 \ctrlR_REG[197] ( .CK(uclk), .D(n730), .Q(ctrlR[197]), .QN( ));
Q_FDP0 \ctrlR_REG[198] ( .CK(uclk), .D(n731), .Q(ctrlR[198]), .QN( ));
Q_FDP0 \ctrlR_REG[199] ( .CK(uclk), .D(n732), .Q(ctrlR[199]), .QN( ));
Q_FDP0 \ctrlR_REG[200] ( .CK(uclk), .D(n733), .Q(ctrlR[200]), .QN( ));
Q_FDP0 \ctrlR_REG[201] ( .CK(uclk), .D(n734), .Q(ctrlR[201]), .QN( ));
Q_FDP0 \ctrlR_REG[202] ( .CK(uclk), .D(n735), .Q(ctrlR[202]), .QN( ));
Q_FDP0 \ctrlR_REG[203] ( .CK(uclk), .D(n736), .Q(ctrlR[203]), .QN( ));
Q_FDP0 \ctrlR_REG[204] ( .CK(uclk), .D(n737), .Q(ctrlR[204]), .QN( ));
Q_FDP0 \ctrlR_REG[205] ( .CK(uclk), .D(n738), .Q(ctrlR[205]), .QN( ));
Q_FDP0 \ctrlR_REG[206] ( .CK(uclk), .D(n739), .Q(ctrlR[206]), .QN( ));
Q_FDP0 \ctrlR_REG[207] ( .CK(uclk), .D(n740), .Q(ctrlR[207]), .QN( ));
Q_FDP0 \ctrlR_REG[208] ( .CK(uclk), .D(n741), .Q(ctrlR[208]), .QN( ));
Q_FDP0 \ctrlR_REG[209] ( .CK(uclk), .D(n742), .Q(ctrlR[209]), .QN( ));
Q_FDP0 \ctrlR_REG[210] ( .CK(uclk), .D(n743), .Q(ctrlR[210]), .QN( ));
Q_FDP0 \ctrlR_REG[211] ( .CK(uclk), .D(n744), .Q(ctrlR[211]), .QN( ));
Q_FDP0 \ctrlR_REG[212] ( .CK(uclk), .D(n745), .Q(ctrlR[212]), .QN( ));
Q_FDP0 \ctrlR_REG[213] ( .CK(uclk), .D(n746), .Q(ctrlR[213]), .QN( ));
Q_FDP0 \ctrlR_REG[214] ( .CK(uclk), .D(n747), .Q(ctrlR[214]), .QN( ));
Q_FDP0 \ctrlR_REG[215] ( .CK(uclk), .D(n748), .Q(ctrlR[215]), .QN( ));
Q_FDP0 \ctrlR_REG[216] ( .CK(uclk), .D(n749), .Q(ctrlR[216]), .QN( ));
Q_FDP0 \ctrlR_REG[217] ( .CK(uclk), .D(n750), .Q(ctrlR[217]), .QN( ));
Q_FDP0 \ctrlR_REG[218] ( .CK(uclk), .D(n751), .Q(ctrlR[218]), .QN( ));
Q_FDP0 \ctrlR_REG[219] ( .CK(uclk), .D(n752), .Q(ctrlR[219]), .QN( ));
Q_FDP0 \ctrlR_REG[220] ( .CK(uclk), .D(n753), .Q(ctrlR[220]), .QN( ));
Q_FDP0 \ctrlR_REG[221] ( .CK(uclk), .D(n754), .Q(ctrlR[221]), .QN( ));
Q_FDP0 \ctrlR_REG[222] ( .CK(uclk), .D(n755), .Q(ctrlR[222]), .QN( ));
Q_FDP0 \ctrlR_REG[223] ( .CK(uclk), .D(n756), .Q(ctrlR[223]), .QN( ));
Q_FDP0 \ctrlR_REG[224] ( .CK(uclk), .D(n757), .Q(ctrlR[224]), .QN( ));
Q_FDP0 \ctrlR_REG[225] ( .CK(uclk), .D(n758), .Q(ctrlR[225]), .QN( ));
Q_FDP0 \ctrlR_REG[226] ( .CK(uclk), .D(n759), .Q(ctrlR[226]), .QN( ));
Q_FDP0 \ctrlR_REG[227] ( .CK(uclk), .D(n760), .Q(ctrlR[227]), .QN( ));
Q_FDP0 \ctrlR_REG[228] ( .CK(uclk), .D(n761), .Q(ctrlR[228]), .QN( ));
Q_FDP0 \ctrlR_REG[229] ( .CK(uclk), .D(n762), .Q(ctrlR[229]), .QN( ));
Q_FDP0 \ctrlR_REG[230] ( .CK(uclk), .D(n763), .Q(ctrlR[230]), .QN( ));
Q_FDP0 \ctrlR_REG[231] ( .CK(uclk), .D(n764), .Q(ctrlR[231]), .QN( ));
Q_FDP0 \ctrlR_REG[232] ( .CK(uclk), .D(n765), .Q(ctrlR[232]), .QN( ));
Q_FDP0 \ctrlR_REG[233] ( .CK(uclk), .D(n766), .Q(ctrlR[233]), .QN( ));
Q_FDP0 \ctrlR_REG[234] ( .CK(uclk), .D(n767), .Q(ctrlR[234]), .QN( ));
Q_FDP0 \ctrlR_REG[235] ( .CK(uclk), .D(n768), .Q(ctrlR[235]), .QN( ));
Q_FDP0 \ctrlR_REG[236] ( .CK(uclk), .D(n769), .Q(ctrlR[236]), .QN( ));
Q_FDP0 \ctrlR_REG[237] ( .CK(uclk), .D(n770), .Q(ctrlR[237]), .QN( ));
Q_FDP0 \ctrlR_REG[238] ( .CK(uclk), .D(n771), .Q(ctrlR[238]), .QN( ));
Q_FDP0 \ctrlR_REG[239] ( .CK(uclk), .D(n772), .Q(ctrlR[239]), .QN( ));
Q_FDP0 \ctrlR_REG[240] ( .CK(uclk), .D(n773), .Q(ctrlR[240]), .QN( ));
Q_FDP0 \ctrlR_REG[241] ( .CK(uclk), .D(n774), .Q(ctrlR[241]), .QN( ));
Q_FDP0 \ctrlR_REG[242] ( .CK(uclk), .D(n775), .Q(ctrlR[242]), .QN( ));
Q_FDP0 \ctrlR_REG[243] ( .CK(uclk), .D(n776), .Q(ctrlR[243]), .QN( ));
Q_FDP0 \ctrlR_REG[244] ( .CK(uclk), .D(n777), .Q(ctrlR[244]), .QN( ));
Q_FDP0 \ctrlR_REG[245] ( .CK(uclk), .D(n778), .Q(ctrlR[245]), .QN( ));
Q_FDP0 \ctrlR_REG[246] ( .CK(uclk), .D(n779), .Q(ctrlR[246]), .QN( ));
Q_FDP0 \ctrlR_REG[247] ( .CK(uclk), .D(n780), .Q(ctrlR[247]), .QN( ));
Q_FDP0 \ctrlR_REG[248] ( .CK(uclk), .D(n781), .Q(ctrlR[248]), .QN( ));
Q_FDP0 \ctrlR_REG[249] ( .CK(uclk), .D(n782), .Q(ctrlR[249]), .QN( ));
Q_FDP0 \ctrlR_REG[250] ( .CK(uclk), .D(n783), .Q(ctrlR[250]), .QN( ));
Q_FDP0 \ctrlR_REG[251] ( .CK(uclk), .D(n784), .Q(ctrlR[251]), .QN( ));
Q_FDP0 \ctrlR_REG[252] ( .CK(uclk), .D(n785), .Q(ctrlR[252]), .QN( ));
Q_FDP0 \ctrlR_REG[253] ( .CK(uclk), .D(n786), .Q(ctrlR[253]), .QN( ));
Q_FDP0 \ctrlR_REG[254] ( .CK(uclk), .D(n787), .Q(ctrlR[254]), .QN( ));
Q_FDP0 \ctrlR_REG[255] ( .CK(uclk), .D(n788), .Q(ctrlR[255]), .QN( ));
Q_MX02 U455 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[62]), .A1(n530), .Z(ecmTs[62]));
Q_MX02 U456 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[61]), .A1(n528), .Z(ecmTs[61]));
Q_MX02 U457 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[60]), .A1(n526), .Z(ecmTs[60]));
Q_MX02 U458 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[59]), .A1(n524), .Z(ecmTs[59]));
Q_MX02 U459 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[58]), .A1(n522), .Z(ecmTs[58]));
Q_MX02 U460 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[57]), .A1(n520), .Z(ecmTs[57]));
Q_MX02 U461 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[56]), .A1(n518), .Z(ecmTs[56]));
Q_MX02 U462 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[55]), .A1(n516), .Z(ecmTs[55]));
Q_MX02 U463 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[54]), .A1(n514), .Z(ecmTs[54]));
Q_MX02 U464 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[53]), .A1(n512), .Z(ecmTs[53]));
Q_MX02 U465 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[52]), .A1(n510), .Z(ecmTs[52]));
Q_MX02 U466 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[51]), .A1(n508), .Z(ecmTs[51]));
Q_MX02 U467 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[50]), .A1(n506), .Z(ecmTs[50]));
Q_MX02 U468 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[49]), .A1(n504), .Z(ecmTs[49]));
Q_MX02 U469 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[48]), .A1(n502), .Z(ecmTs[48]));
Q_MX02 U470 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[47]), .A1(n500), .Z(ecmTs[47]));
Q_MX02 U471 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[46]), .A1(n498), .Z(ecmTs[46]));
Q_MX02 U472 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[45]), .A1(n496), .Z(ecmTs[45]));
Q_MX02 U473 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[44]), .A1(n494), .Z(ecmTs[44]));
Q_MX02 U474 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[43]), .A1(n492), .Z(ecmTs[43]));
Q_MX02 U475 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[42]), .A1(n490), .Z(ecmTs[42]));
Q_MX02 U476 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[41]), .A1(n488), .Z(ecmTs[41]));
Q_MX02 U477 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[40]), .A1(n486), .Z(ecmTs[40]));
Q_MX02 U478 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[39]), .A1(n484), .Z(ecmTs[39]));
Q_MX02 U479 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[38]), .A1(n482), .Z(ecmTs[38]));
Q_MX02 U480 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[37]), .A1(n480), .Z(ecmTs[37]));
Q_MX02 U481 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[36]), .A1(n478), .Z(ecmTs[36]));
Q_MX02 U482 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[35]), .A1(n476), .Z(ecmTs[35]));
Q_MX02 U483 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[34]), .A1(n474), .Z(ecmTs[34]));
Q_MX02 U484 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[33]), .A1(n472), .Z(ecmTs[33]));
Q_MX02 U485 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[32]), .A1(n470), .Z(ecmTs[32]));
Q_MX02 U486 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[31]), .A1(n468), .Z(ecmTs[31]));
Q_MX02 U487 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[30]), .A1(n466), .Z(ecmTs[30]));
Q_MX02 U488 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[29]), .A1(n464), .Z(ecmTs[29]));
Q_MX02 U489 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[28]), .A1(n462), .Z(ecmTs[28]));
Q_MX02 U490 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[27]), .A1(n460), .Z(ecmTs[27]));
Q_MX02 U491 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[26]), .A1(n458), .Z(ecmTs[26]));
Q_MX02 U492 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[25]), .A1(n456), .Z(ecmTs[25]));
Q_MX02 U493 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[24]), .A1(n454), .Z(ecmTs[24]));
Q_MX02 U494 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[23]), .A1(n452), .Z(ecmTs[23]));
Q_MX02 U495 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[22]), .A1(n450), .Z(ecmTs[22]));
Q_MX02 U496 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[21]), .A1(n448), .Z(ecmTs[21]));
Q_MX02 U497 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[20]), .A1(n446), .Z(ecmTs[20]));
Q_MX02 U498 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[19]), .A1(n444), .Z(ecmTs[19]));
Q_MX02 U499 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[18]), .A1(n442), .Z(ecmTs[18]));
Q_MX02 U500 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[17]), .A1(n440), .Z(ecmTs[17]));
Q_MX02 U501 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[16]), .A1(n438), .Z(ecmTs[16]));
Q_MX02 U502 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[15]), .A1(n436), .Z(ecmTs[15]));
Q_MX02 U503 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[14]), .A1(n434), .Z(ecmTs[14]));
Q_MX02 U504 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[13]), .A1(n432), .Z(ecmTs[13]));
Q_MX02 U505 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[12]), .A1(n430), .Z(ecmTs[12]));
Q_MX02 U506 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[11]), .A1(n428), .Z(ecmTs[11]));
Q_MX02 U507 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[10]), .A1(n426), .Z(ecmTs[10]));
Q_MX02 U508 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[9]), .A1(n424), .Z(ecmTs[9]));
Q_MX02 U509 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[8]), .A1(n422), .Z(ecmTs[8]));
Q_MX02 U510 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[7]), .A1(n420), .Z(ecmTs[7]));
Q_MX02 U511 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[6]), .A1(n418), .Z(ecmTs[6]));
Q_MX02 U512 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[5]), .A1(n416), .Z(ecmTs[5]));
Q_MX02 U513 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[4]), .A1(n414), .Z(ecmTs[4]));
Q_MX02 U514 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[3]), .A1(n412), .Z(ecmTs[3]));
Q_MX02 U515 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[2]), .A1(n410), .Z(ecmTs[2]));
Q_MX02 U516 ( .S(xcva_top.xc_top.ecmOnD), .A0(ecmTsP[1]), .A1(n408), .Z(ecmTs[1]));
Q_XOR2 U517 ( .A0(xcva_top.xc_top.ecmOnD), .A1(ecmTsP[0]), .Z(ecmTs[0]));
Q_XOR2 U518 ( .A0(ecmTsP[63]), .A1(n791), .Z(ecmTs[63]));
Q_AD01HF U519 ( .A0(ecmTsP[62]), .B0(n529), .S(n530), .CO(n531));
Q_AD01HF U520 ( .A0(ecmTsP[61]), .B0(n527), .S(n528), .CO(n529));
Q_AD01HF U521 ( .A0(ecmTsP[60]), .B0(n525), .S(n526), .CO(n527));
Q_AD01HF U522 ( .A0(ecmTsP[59]), .B0(n523), .S(n524), .CO(n525));
Q_AD01HF U523 ( .A0(ecmTsP[58]), .B0(n521), .S(n522), .CO(n523));
Q_AD01HF U524 ( .A0(ecmTsP[57]), .B0(n519), .S(n520), .CO(n521));
Q_AD01HF U525 ( .A0(ecmTsP[56]), .B0(n517), .S(n518), .CO(n519));
Q_AD01HF U526 ( .A0(ecmTsP[55]), .B0(n515), .S(n516), .CO(n517));
Q_AD01HF U527 ( .A0(ecmTsP[54]), .B0(n513), .S(n514), .CO(n515));
Q_AD01HF U528 ( .A0(ecmTsP[53]), .B0(n511), .S(n512), .CO(n513));
Q_AD01HF U529 ( .A0(ecmTsP[52]), .B0(n509), .S(n510), .CO(n511));
Q_AD01HF U530 ( .A0(ecmTsP[51]), .B0(n507), .S(n508), .CO(n509));
Q_AD01HF U531 ( .A0(ecmTsP[50]), .B0(n505), .S(n506), .CO(n507));
Q_AD01HF U532 ( .A0(ecmTsP[49]), .B0(n503), .S(n504), .CO(n505));
Q_AD01HF U533 ( .A0(ecmTsP[48]), .B0(n501), .S(n502), .CO(n503));
Q_AD01HF U534 ( .A0(ecmTsP[47]), .B0(n499), .S(n500), .CO(n501));
Q_AD01HF U535 ( .A0(ecmTsP[46]), .B0(n497), .S(n498), .CO(n499));
Q_AD01HF U536 ( .A0(ecmTsP[45]), .B0(n495), .S(n496), .CO(n497));
Q_AD01HF U537 ( .A0(ecmTsP[44]), .B0(n493), .S(n494), .CO(n495));
Q_AD01HF U538 ( .A0(ecmTsP[43]), .B0(n491), .S(n492), .CO(n493));
Q_AD01HF U539 ( .A0(ecmTsP[42]), .B0(n489), .S(n490), .CO(n491));
Q_AD01HF U540 ( .A0(ecmTsP[41]), .B0(n487), .S(n488), .CO(n489));
Q_AD01HF U541 ( .A0(ecmTsP[40]), .B0(n485), .S(n486), .CO(n487));
Q_AD01HF U542 ( .A0(ecmTsP[39]), .B0(n483), .S(n484), .CO(n485));
Q_AD01HF U543 ( .A0(ecmTsP[38]), .B0(n481), .S(n482), .CO(n483));
Q_AD01HF U544 ( .A0(ecmTsP[37]), .B0(n479), .S(n480), .CO(n481));
Q_AD01HF U545 ( .A0(ecmTsP[36]), .B0(n477), .S(n478), .CO(n479));
Q_AD01HF U546 ( .A0(ecmTsP[35]), .B0(n475), .S(n476), .CO(n477));
Q_AD01HF U547 ( .A0(ecmTsP[34]), .B0(n473), .S(n474), .CO(n475));
Q_AD01HF U548 ( .A0(ecmTsP[33]), .B0(n471), .S(n472), .CO(n473));
Q_AD01HF U549 ( .A0(ecmTsP[32]), .B0(n469), .S(n470), .CO(n471));
Q_AD01HF U550 ( .A0(ecmTsP[31]), .B0(n467), .S(n468), .CO(n469));
Q_AD01HF U551 ( .A0(ecmTsP[30]), .B0(n465), .S(n466), .CO(n467));
Q_AD01HF U552 ( .A0(ecmTsP[29]), .B0(n463), .S(n464), .CO(n465));
Q_AD01HF U553 ( .A0(ecmTsP[28]), .B0(n461), .S(n462), .CO(n463));
Q_AD01HF U554 ( .A0(ecmTsP[27]), .B0(n459), .S(n460), .CO(n461));
Q_AD01HF U555 ( .A0(ecmTsP[26]), .B0(n457), .S(n458), .CO(n459));
Q_AD01HF U556 ( .A0(ecmTsP[25]), .B0(n455), .S(n456), .CO(n457));
Q_AD01HF U557 ( .A0(ecmTsP[24]), .B0(n453), .S(n454), .CO(n455));
Q_AD01HF U558 ( .A0(ecmTsP[23]), .B0(n451), .S(n452), .CO(n453));
Q_AD01HF U559 ( .A0(ecmTsP[22]), .B0(n449), .S(n450), .CO(n451));
Q_AD01HF U560 ( .A0(ecmTsP[21]), .B0(n447), .S(n448), .CO(n449));
Q_AD01HF U561 ( .A0(ecmTsP[20]), .B0(n445), .S(n446), .CO(n447));
Q_AD01HF U562 ( .A0(ecmTsP[19]), .B0(n443), .S(n444), .CO(n445));
Q_AD01HF U563 ( .A0(ecmTsP[18]), .B0(n441), .S(n442), .CO(n443));
Q_AD01HF U564 ( .A0(ecmTsP[17]), .B0(n439), .S(n440), .CO(n441));
Q_AD01HF U565 ( .A0(ecmTsP[16]), .B0(n437), .S(n438), .CO(n439));
Q_AD01HF U566 ( .A0(ecmTsP[15]), .B0(n435), .S(n436), .CO(n437));
Q_AD01HF U567 ( .A0(ecmTsP[14]), .B0(n433), .S(n434), .CO(n435));
Q_AD01HF U568 ( .A0(ecmTsP[13]), .B0(n431), .S(n432), .CO(n433));
Q_AD01HF U569 ( .A0(ecmTsP[12]), .B0(n429), .S(n430), .CO(n431));
Q_AD01HF U570 ( .A0(ecmTsP[11]), .B0(n427), .S(n428), .CO(n429));
Q_AD01HF U571 ( .A0(ecmTsP[10]), .B0(n425), .S(n426), .CO(n427));
Q_AD01HF U572 ( .A0(ecmTsP[9]), .B0(n423), .S(n424), .CO(n425));
Q_AD01HF U573 ( .A0(ecmTsP[8]), .B0(n421), .S(n422), .CO(n423));
Q_AD01HF U574 ( .A0(ecmTsP[7]), .B0(n419), .S(n420), .CO(n421));
Q_AD01HF U575 ( .A0(ecmTsP[6]), .B0(n417), .S(n418), .CO(n419));
Q_AD01HF U576 ( .A0(ecmTsP[5]), .B0(n415), .S(n416), .CO(n417));
Q_AD01HF U577 ( .A0(ecmTsP[4]), .B0(n413), .S(n414), .CO(n415));
Q_AD01HF U578 ( .A0(ecmTsP[3]), .B0(n411), .S(n412), .CO(n413));
Q_AD01HF U579 ( .A0(ecmTsP[2]), .B0(n409), .S(n410), .CO(n411));
Q_AD01HF U580 ( .A0(ecmTsP[1]), .B0(ecmTsP[0]), .S(n408), .CO(n409));
Q_OR03 U581 ( .A0(n406), .A1(n407), .A2(newCtrl), .Z(busyOn));
Q_OR03 U582 ( .A0(busyCnt[1]), .A1(busyCnt[0]), .A2(n405), .Z(n407));
Q_OR03 U583 ( .A0(busyCnt[4]), .A1(busyCnt[3]), .A2(busyCnt[2]), .Z(n406));
Q_OR03 U584 ( .A0(busyCnt[7]), .A1(busyCnt[6]), .A2(busyCnt[5]), .Z(n405));
Q_XOR2 U585 ( .A0(ctrlEv), .A1(ctrlEvP), .Z(newCtrl));
Q_INV U586 ( .A(n404), .Z(newCmd));
Q_AN02 U587 ( .A0(n402), .A1(n403), .Z(n404));
Q_AN03 U588 ( .A0(n394), .A1(n393), .A2(n401), .Z(n403));
Q_AN03 U589 ( .A0(n397), .A1(n396), .A2(n395), .Z(n402));
Q_AN03 U590 ( .A0(n400), .A1(n399), .A2(n398), .Z(n401));
Q_XNR2 U591 ( .A0(cmdCnt[7]), .A1(cmdCntP[7]), .Z(n400));
Q_XNR2 U592 ( .A0(cmdCnt[6]), .A1(cmdCntP[6]), .Z(n399));
Q_XNR2 U593 ( .A0(cmdCnt[5]), .A1(cmdCntP[5]), .Z(n398));
Q_XNR2 U594 ( .A0(cmdCnt[4]), .A1(cmdCntP[4]), .Z(n397));
Q_XNR2 U595 ( .A0(cmdCnt[3]), .A1(cmdCntP[3]), .Z(n396));
Q_XNR2 U596 ( .A0(cmdCnt[2]), .A1(cmdCntP[2]), .Z(n395));
Q_XNR2 U597 ( .A0(cmdCnt[1]), .A1(cmdCntP[1]), .Z(n394));
Q_XNR2 U598 ( .A0(cmdCnt[0]), .A1(cmdCntP[0]), .Z(n393));
Q_FDP0UA U599 ( .D(ctrlEv), .QTFCLK( ), .Q(ctrlEvP));
Q_FDP0UA U600 ( .D(ctrlW[64]), .QTFCLK( ), .Q(ecmTsP[0]));
Q_FDP0UA U601 ( .D(ctrlW[65]), .QTFCLK( ), .Q(ecmTsP[1]));
Q_FDP0UA U602 ( .D(ctrlW[66]), .QTFCLK( ), .Q(ecmTsP[2]));
Q_FDP0UA U603 ( .D(ctrlW[67]), .QTFCLK( ), .Q(ecmTsP[3]));
Q_FDP0UA U604 ( .D(ctrlW[68]), .QTFCLK( ), .Q(ecmTsP[4]));
Q_FDP0UA U605 ( .D(ctrlW[69]), .QTFCLK( ), .Q(ecmTsP[5]));
Q_FDP0UA U606 ( .D(ctrlW[70]), .QTFCLK( ), .Q(ecmTsP[6]));
Q_FDP0UA U607 ( .D(ctrlW[71]), .QTFCLK( ), .Q(ecmTsP[7]));
Q_FDP0UA U608 ( .D(ctrlW[72]), .QTFCLK( ), .Q(ecmTsP[8]));
Q_FDP0UA U609 ( .D(ctrlW[73]), .QTFCLK( ), .Q(ecmTsP[9]));
Q_FDP0UA U610 ( .D(ctrlW[74]), .QTFCLK( ), .Q(ecmTsP[10]));
Q_FDP0UA U611 ( .D(ctrlW[75]), .QTFCLK( ), .Q(ecmTsP[11]));
Q_FDP0UA U612 ( .D(ctrlW[76]), .QTFCLK( ), .Q(ecmTsP[12]));
Q_FDP0UA U613 ( .D(ctrlW[77]), .QTFCLK( ), .Q(ecmTsP[13]));
Q_FDP0UA U614 ( .D(ctrlW[78]), .QTFCLK( ), .Q(ecmTsP[14]));
Q_FDP0UA U615 ( .D(ctrlW[79]), .QTFCLK( ), .Q(ecmTsP[15]));
Q_FDP0UA U616 ( .D(ctrlW[80]), .QTFCLK( ), .Q(ecmTsP[16]));
Q_FDP0UA U617 ( .D(ctrlW[81]), .QTFCLK( ), .Q(ecmTsP[17]));
Q_FDP0UA U618 ( .D(ctrlW[82]), .QTFCLK( ), .Q(ecmTsP[18]));
Q_FDP0UA U619 ( .D(ctrlW[83]), .QTFCLK( ), .Q(ecmTsP[19]));
Q_FDP0UA U620 ( .D(ctrlW[84]), .QTFCLK( ), .Q(ecmTsP[20]));
Q_FDP0UA U621 ( .D(ctrlW[85]), .QTFCLK( ), .Q(ecmTsP[21]));
Q_FDP0UA U622 ( .D(ctrlW[86]), .QTFCLK( ), .Q(ecmTsP[22]));
Q_FDP0UA U623 ( .D(ctrlW[87]), .QTFCLK( ), .Q(ecmTsP[23]));
Q_FDP0UA U624 ( .D(ctrlW[88]), .QTFCLK( ), .Q(ecmTsP[24]));
Q_FDP0UA U625 ( .D(ctrlW[89]), .QTFCLK( ), .Q(ecmTsP[25]));
Q_FDP0UA U626 ( .D(ctrlW[90]), .QTFCLK( ), .Q(ecmTsP[26]));
Q_FDP0UA U627 ( .D(ctrlW[91]), .QTFCLK( ), .Q(ecmTsP[27]));
Q_FDP0UA U628 ( .D(ctrlW[92]), .QTFCLK( ), .Q(ecmTsP[28]));
Q_FDP0UA U629 ( .D(ctrlW[93]), .QTFCLK( ), .Q(ecmTsP[29]));
Q_FDP0UA U630 ( .D(ctrlW[94]), .QTFCLK( ), .Q(ecmTsP[30]));
Q_FDP0UA U631 ( .D(ctrlW[95]), .QTFCLK( ), .Q(ecmTsP[31]));
Q_FDP0UA U632 ( .D(ctrlW[96]), .QTFCLK( ), .Q(ecmTsP[32]));
Q_FDP0UA U633 ( .D(ctrlW[97]), .QTFCLK( ), .Q(ecmTsP[33]));
Q_FDP0UA U634 ( .D(ctrlW[98]), .QTFCLK( ), .Q(ecmTsP[34]));
Q_FDP0UA U635 ( .D(ctrlW[99]), .QTFCLK( ), .Q(ecmTsP[35]));
Q_FDP0UA U636 ( .D(ctrlW[100]), .QTFCLK( ), .Q(ecmTsP[36]));
Q_FDP0UA U637 ( .D(ctrlW[101]), .QTFCLK( ), .Q(ecmTsP[37]));
Q_FDP0UA U638 ( .D(ctrlW[102]), .QTFCLK( ), .Q(ecmTsP[38]));
Q_FDP0UA U639 ( .D(ctrlW[103]), .QTFCLK( ), .Q(ecmTsP[39]));
Q_FDP0UA U640 ( .D(ctrlW[104]), .QTFCLK( ), .Q(ecmTsP[40]));
Q_FDP0UA U641 ( .D(ctrlW[105]), .QTFCLK( ), .Q(ecmTsP[41]));
Q_FDP0UA U642 ( .D(ctrlW[106]), .QTFCLK( ), .Q(ecmTsP[42]));
Q_FDP0UA U643 ( .D(ctrlW[107]), .QTFCLK( ), .Q(ecmTsP[43]));
Q_FDP0UA U644 ( .D(ctrlW[108]), .QTFCLK( ), .Q(ecmTsP[44]));
Q_FDP0UA U645 ( .D(ctrlW[109]), .QTFCLK( ), .Q(ecmTsP[45]));
Q_FDP0UA U646 ( .D(ctrlW[110]), .QTFCLK( ), .Q(ecmTsP[46]));
Q_FDP0UA U647 ( .D(ctrlW[111]), .QTFCLK( ), .Q(ecmTsP[47]));
Q_FDP0UA U648 ( .D(ctrlW[112]), .QTFCLK( ), .Q(ecmTsP[48]));
Q_FDP0UA U649 ( .D(ctrlW[113]), .QTFCLK( ), .Q(ecmTsP[49]));
Q_FDP0UA U650 ( .D(ctrlW[114]), .QTFCLK( ), .Q(ecmTsP[50]));
Q_FDP0UA U651 ( .D(ctrlW[115]), .QTFCLK( ), .Q(ecmTsP[51]));
Q_FDP0UA U652 ( .D(ctrlW[116]), .QTFCLK( ), .Q(ecmTsP[52]));
Q_FDP0UA U653 ( .D(ctrlW[117]), .QTFCLK( ), .Q(ecmTsP[53]));
Q_FDP0UA U654 ( .D(ctrlW[118]), .QTFCLK( ), .Q(ecmTsP[54]));
Q_FDP0UA U655 ( .D(ctrlW[119]), .QTFCLK( ), .Q(ecmTsP[55]));
Q_FDP0UA U656 ( .D(ctrlW[120]), .QTFCLK( ), .Q(ecmTsP[56]));
Q_FDP0UA U657 ( .D(ctrlW[121]), .QTFCLK( ), .Q(ecmTsP[57]));
Q_FDP0UA U658 ( .D(ctrlW[122]), .QTFCLK( ), .Q(ecmTsP[58]));
Q_FDP0UA U659 ( .D(ctrlW[123]), .QTFCLK( ), .Q(ecmTsP[59]));
Q_FDP0UA U660 ( .D(ctrlW[124]), .QTFCLK( ), .Q(ecmTsP[60]));
Q_FDP0UA U661 ( .D(ctrlW[125]), .QTFCLK( ), .Q(ecmTsP[61]));
Q_FDP0UA U662 ( .D(ctrlW[126]), .QTFCLK( ), .Q(ecmTsP[62]));
Q_FDP0UA U663 ( .D(ctrlW[127]), .QTFCLK( ), .Q(ecmTsP[63]));
Q_FDP0UA U664 ( .D(newCtrl), .QTFCLK( ), .Q(busyCnt[0]));
Q_FDP0UA U665 ( .D(busyCnt[0]), .QTFCLK( ), .Q(busyCnt[1]));
Q_FDP0UA U666 ( .D(busyCnt[1]), .QTFCLK( ), .Q(busyCnt[2]));
Q_FDP0UA U667 ( .D(busyCnt[2]), .QTFCLK( ), .Q(busyCnt[3]));
Q_FDP0UA U668 ( .D(busyCnt[3]), .QTFCLK( ), .Q(busyCnt[4]));
Q_FDP0UA U669 ( .D(busyCnt[4]), .QTFCLK( ), .Q(busyCnt[5]));
Q_FDP0UA U670 ( .D(busyCnt[5]), .QTFCLK( ), .Q(busyCnt[6]));
Q_FDP0UA U671 ( .D(busyCnt[6]), .QTFCLK( ), .Q(busyCnt[7]));
Q_FDP0UA U672 ( .D(n391), .QTFCLK( ), .Q(cmdCntP[7]));
Q_MX02 U673 ( .S(n372), .A0(cmdCntP[7]), .A1(cmdCnt[7]), .Z(n391));
Q_FDP0UA U674 ( .D(n390), .QTFCLK( ), .Q(cmdCntP[6]));
Q_MX02 U675 ( .S(n372), .A0(cmdCntP[6]), .A1(cmdCnt[6]), .Z(n390));
Q_FDP0UA U676 ( .D(n389), .QTFCLK( ), .Q(cmdCntP[5]));
Q_MX02 U677 ( .S(n372), .A0(cmdCntP[5]), .A1(cmdCnt[5]), .Z(n389));
Q_FDP0UA U678 ( .D(n388), .QTFCLK( ), .Q(cmdCntP[4]));
Q_MX02 U679 ( .S(n372), .A0(cmdCntP[4]), .A1(cmdCnt[4]), .Z(n388));
Q_FDP0UA U680 ( .D(n387), .QTFCLK( ), .Q(cmdCntP[3]));
Q_MX02 U681 ( .S(n372), .A0(cmdCntP[3]), .A1(cmdCnt[3]), .Z(n387));
Q_FDP0UA U682 ( .D(n386), .QTFCLK( ), .Q(cmdCntP[2]));
Q_MX02 U683 ( .S(n372), .A0(cmdCntP[2]), .A1(cmdCnt[2]), .Z(n386));
Q_FDP0UA U684 ( .D(n385), .QTFCLK( ), .Q(cmdCntP[1]));
Q_MX02 U685 ( .S(n372), .A0(cmdCntP[1]), .A1(cmdCnt[1]), .Z(n385));
Q_FDP0UA U686 ( .D(n384), .QTFCLK( ), .Q(cmdCntP[0]));
Q_MX02 U687 ( .S(n372), .A0(cmdCntP[0]), .A1(cmdCnt[0]), .Z(n384));
Q_FDP0UA U688 ( .D(n383), .QTFCLK( ), .Q(cRet[15]));
Q_MX02 U689 ( .S(n372), .A0(ctrlW[15]), .A1(cmdCnt[7]), .Z(n383));
Q_FDP0UA U690 ( .D(n382), .QTFCLK( ), .Q(cRet[14]));
Q_MX02 U691 ( .S(n372), .A0(ctrlW[14]), .A1(cmdCnt[6]), .Z(n382));
Q_FDP0UA U692 ( .D(n381), .QTFCLK( ), .Q(cRet[13]));
Q_MX02 U693 ( .S(n372), .A0(ctrlW[13]), .A1(cmdCnt[5]), .Z(n381));
Q_FDP0UA U694 ( .D(n380), .QTFCLK( ), .Q(cRet[12]));
Q_MX02 U695 ( .S(n372), .A0(ctrlW[12]), .A1(cmdCnt[4]), .Z(n380));
Q_FDP0UA U696 ( .D(n379), .QTFCLK( ), .Q(cRet[11]));
Q_MX02 U697 ( .S(n372), .A0(ctrlW[11]), .A1(cmdCnt[3]), .Z(n379));
Q_FDP0UA U698 ( .D(n378), .QTFCLK( ), .Q(cRet[10]));
Q_MX02 U699 ( .S(n372), .A0(ctrlW[10]), .A1(cmdCnt[2]), .Z(n378));
Q_FDP0UA U700 ( .D(n377), .QTFCLK( ), .Q(cRet[9]));
Q_MX02 U701 ( .S(n372), .A0(ctrlW[9]), .A1(cmdCnt[1]), .Z(n377));
Q_FDP0UA U702 ( .D(n376), .QTFCLK( ), .Q(cRet[8]));
Q_MX02 U703 ( .S(n372), .A0(ctrlW[8]), .A1(cmdCnt[0]), .Z(n376));
Q_ND03 U704 ( .A0(holdEcm), .A1(xcva_top.xc_top.ptxStop), .A2(xcva_top.xc_top.evalOnC), .Z(n371));
Q_INV U705 ( .A(n373), .Z(n375));
Q_FDP0UA U706 ( .D(n375), .QTFCLK( ), .Q(_zyL831_meState0[0]));
Q_AO21 U707 ( .A0(n374), .A1(n404), .B0(n372), .Z(n373));
Q_INV U708 ( .A(_zyL831_meState0[0]), .Z(n374));
Q_AN02 U709 ( .A0(_zyL831_meState0[0]), .A1(n371), .Z(n372));
Q_FDP0UA U710 ( .D(ctrlR[128]), .QTFCLK( ), .Q(cmdC[0]));
Q_FDP0UA U711 ( .D(ctrlR[129]), .QTFCLK( ), .Q(cmdC[1]));
Q_FDP0UA U712 ( .D(ctrlR[130]), .QTFCLK( ), .Q(cmdC[2]));
Q_FDP0UA U713 ( .D(ctrlR[131]), .QTFCLK( ), .Q(cmdC[3]));
Q_FDP0UA U714 ( .D(ctrlR[132]), .QTFCLK( ), .Q(cmdC[4]));
Q_FDP0UA U715 ( .D(ctrlR[133]), .QTFCLK( ), .Q(cmdC[5]));
Q_FDP0UA U716 ( .D(ctrlR[134]), .QTFCLK( ), .Q(cmdC[6]));
Q_FDP0UA U717 ( .D(ctrlR[135]), .QTFCLK( ), .Q(cmdC[7]));
Q_FDP0UA U718 ( .D(ctrlEv), .QTFCLK( ), .Q(cmdCnt[0]));
Q_FDP0UA U719 ( .D(ctrlR[137]), .QTFCLK( ), .Q(cmdCnt[1]));
Q_FDP0UA U720 ( .D(ctrlR[138]), .QTFCLK( ), .Q(cmdCnt[2]));
Q_FDP0UA U721 ( .D(ctrlR[139]), .QTFCLK( ), .Q(cmdCnt[3]));
Q_FDP0UA U722 ( .D(ctrlR[140]), .QTFCLK( ), .Q(cmdCnt[4]));
Q_FDP0UA U723 ( .D(ctrlR[141]), .QTFCLK( ), .Q(cmdCnt[5]));
Q_FDP0UA U724 ( .D(ctrlR[142]), .QTFCLK( ), .Q(cmdCnt[6]));
Q_FDP0UA U725 ( .D(ctrlR[143]), .QTFCLK( ), .Q(cmdCnt[7]));
Q_FDP0UA U726 ( .D(xcva_top.xc_top.ptxStop), .QTFCLK( ), .Q(cRet[2]));
Q_FDP0UA U727 ( .D(n370), .QTFCLK( ), .Q(cRet[1]));
Q_FDP0UA U728 ( .D(n370), .QTFCLK( ), .Q(cRet[0]));
Q_FDP0 U729 ( .CK(uclk), .D(n368), .Q(n369), .QN(n368));
Q_FDP0B U730 ( .D(n369), .QTFCLK( ), .Q(n367));
Q_XOR2 U731 ( .A0(n369), .A1(n367), .Z(n366));
// pragma CVAINTPROP NET n369 _2_state_ 1
// pragma CVAINTPROP INSTANCE U731 NOBREAKS 1
Q_FDP0 U732 ( .CK(uclk), .D(ctrlW[0]), .Q(n365), .QN( ));
Q_FDP0 U733 ( .CK(uclk), .D(ctrlW[1]), .Q(n364), .QN( ));
Q_FDP0 U734 ( .CK(uclk), .D(ctrlW[2]), .Q(n363), .QN( ));
Q_FDP0 U735 ( .CK(uclk), .D(ctrlW[3]), .Q(n362), .QN( ));
Q_FDP0 U736 ( .CK(uclk), .D(ctrlW[4]), .Q(n361), .QN( ));
Q_FDP0 U737 ( .CK(uclk), .D(ctrlW[5]), .Q(n360), .QN( ));
Q_FDP0 U738 ( .CK(uclk), .D(ctrlW[6]), .Q(n359), .QN( ));
Q_FDP0 U739 ( .CK(uclk), .D(ctrlW[7]), .Q(n358), .QN( ));
Q_FDP0 U740 ( .CK(uclk), .D(ctrlW[8]), .Q(n357), .QN( ));
Q_FDP0 U741 ( .CK(uclk), .D(ctrlW[9]), .Q(n356), .QN( ));
Q_FDP0 U742 ( .CK(uclk), .D(ctrlW[10]), .Q(n355), .QN( ));
Q_FDP0 U743 ( .CK(uclk), .D(ctrlW[11]), .Q(n354), .QN( ));
Q_FDP0 U744 ( .CK(uclk), .D(ctrlW[12]), .Q(n353), .QN( ));
Q_FDP0 U745 ( .CK(uclk), .D(ctrlW[13]), .Q(n352), .QN( ));
Q_FDP0 U746 ( .CK(uclk), .D(ctrlW[14]), .Q(n351), .QN( ));
Q_FDP0 U747 ( .CK(uclk), .D(ctrlW[15]), .Q(n350), .QN( ));
Q_FDP0 U748 ( .CK(uclk), .D(ctrlW[16]), .Q(n349), .QN( ));
Q_FDP0 U749 ( .CK(uclk), .D(ctrlW[17]), .Q(n348), .QN( ));
Q_FDP0 U750 ( .CK(uclk), .D(ctrlW[18]), .Q(n347), .QN( ));
Q_FDP0 U751 ( .CK(uclk), .D(ctrlW[19]), .Q(n346), .QN( ));
Q_FDP0 U752 ( .CK(uclk), .D(ctrlW[20]), .Q(n345), .QN( ));
Q_FDP0 U753 ( .CK(uclk), .D(ctrlW[21]), .Q(n344), .QN( ));
Q_FDP0 U754 ( .CK(uclk), .D(ctrlW[22]), .Q(n343), .QN( ));
Q_FDP0 U755 ( .CK(uclk), .D(ctrlW[23]), .Q(n342), .QN( ));
Q_FDP0 U756 ( .CK(uclk), .D(ctrlW[24]), .Q(n341), .QN( ));
Q_FDP0 U757 ( .CK(uclk), .D(ctrlW[25]), .Q(n340), .QN( ));
Q_FDP0 U758 ( .CK(uclk), .D(ctrlW[26]), .Q(n339), .QN( ));
Q_FDP0 U759 ( .CK(uclk), .D(ctrlW[27]), .Q(n338), .QN( ));
Q_FDP0 U760 ( .CK(uclk), .D(ctrlW[28]), .Q(n337), .QN( ));
Q_FDP0 U761 ( .CK(uclk), .D(ctrlW[29]), .Q(n336), .QN( ));
Q_FDP0 U762 ( .CK(uclk), .D(ctrlW[30]), .Q(n335), .QN( ));
Q_FDP0 U763 ( .CK(uclk), .D(ctrlW[31]), .Q(n334), .QN( ));
Q_FDP0 U764 ( .CK(uclk), .D(ctrlW[32]), .Q(n333), .QN( ));
Q_FDP0 U765 ( .CK(uclk), .D(ctrlW[33]), .Q(n332), .QN( ));
Q_FDP0 U766 ( .CK(uclk), .D(ctrlW[34]), .Q(n331), .QN( ));
Q_FDP0 U767 ( .CK(uclk), .D(ctrlW[35]), .Q(n330), .QN( ));
Q_FDP0 U768 ( .CK(uclk), .D(ctrlW[36]), .Q(n329), .QN( ));
Q_FDP0 U769 ( .CK(uclk), .D(ctrlW[37]), .Q(n328), .QN( ));
Q_FDP0 U770 ( .CK(uclk), .D(ctrlW[38]), .Q(n327), .QN( ));
Q_FDP0 U771 ( .CK(uclk), .D(ctrlW[39]), .Q(n326), .QN( ));
Q_FDP0 U772 ( .CK(uclk), .D(ctrlW[40]), .Q(n325), .QN( ));
Q_FDP0 U773 ( .CK(uclk), .D(ctrlW[41]), .Q(n324), .QN( ));
Q_FDP0 U774 ( .CK(uclk), .D(ctrlW[42]), .Q(n323), .QN( ));
Q_FDP0 U775 ( .CK(uclk), .D(ctrlW[43]), .Q(n322), .QN( ));
Q_FDP0 U776 ( .CK(uclk), .D(ctrlW[44]), .Q(n321), .QN( ));
Q_FDP0 U777 ( .CK(uclk), .D(ctrlW[45]), .Q(n320), .QN( ));
Q_FDP0 U778 ( .CK(uclk), .D(ctrlW[46]), .Q(n319), .QN( ));
Q_FDP0 U779 ( .CK(uclk), .D(ctrlW[47]), .Q(n318), .QN( ));
Q_FDP0 U780 ( .CK(uclk), .D(ctrlW[48]), .Q(n317), .QN( ));
Q_FDP0 U781 ( .CK(uclk), .D(ctrlW[49]), .Q(n316), .QN( ));
Q_FDP0 U782 ( .CK(uclk), .D(ctrlW[50]), .Q(n315), .QN( ));
Q_FDP0 U783 ( .CK(uclk), .D(ctrlW[51]), .Q(n314), .QN( ));
Q_FDP0 U784 ( .CK(uclk), .D(ctrlW[52]), .Q(n313), .QN( ));
Q_FDP0 U785 ( .CK(uclk), .D(ctrlW[53]), .Q(n312), .QN( ));
Q_FDP0 U786 ( .CK(uclk), .D(ctrlW[54]), .Q(n311), .QN( ));
Q_FDP0 U787 ( .CK(uclk), .D(ctrlW[55]), .Q(n310), .QN( ));
Q_FDP0 U788 ( .CK(uclk), .D(ctrlW[56]), .Q(n309), .QN( ));
Q_FDP0 U789 ( .CK(uclk), .D(ctrlW[57]), .Q(n308), .QN( ));
Q_FDP0 U790 ( .CK(uclk), .D(ctrlW[58]), .Q(n307), .QN( ));
Q_FDP0 U791 ( .CK(uclk), .D(ctrlW[59]), .Q(n306), .QN( ));
Q_FDP0 U792 ( .CK(uclk), .D(ctrlW[60]), .Q(n305), .QN( ));
Q_FDP0 U793 ( .CK(uclk), .D(ctrlW[61]), .Q(n304), .QN( ));
Q_FDP0 U794 ( .CK(uclk), .D(ctrlW[62]), .Q(n303), .QN( ));
Q_FDP0 U795 ( .CK(uclk), .D(ctrlW[63]), .Q(n302), .QN( ));
Q_FDP0 U796 ( .CK(uclk), .D(ctrlW[64]), .Q(n301), .QN( ));
Q_FDP0 U797 ( .CK(uclk), .D(ctrlW[65]), .Q(n300), .QN( ));
Q_FDP0 U798 ( .CK(uclk), .D(ctrlW[66]), .Q(n299), .QN( ));
Q_FDP0 U799 ( .CK(uclk), .D(ctrlW[67]), .Q(n298), .QN( ));
Q_FDP0 U800 ( .CK(uclk), .D(ctrlW[68]), .Q(n297), .QN( ));
Q_FDP0 U801 ( .CK(uclk), .D(ctrlW[69]), .Q(n296), .QN( ));
Q_FDP0 U802 ( .CK(uclk), .D(ctrlW[70]), .Q(n295), .QN( ));
Q_FDP0 U803 ( .CK(uclk), .D(ctrlW[71]), .Q(n294), .QN( ));
Q_FDP0 U804 ( .CK(uclk), .D(ctrlW[72]), .Q(n293), .QN( ));
Q_FDP0 U805 ( .CK(uclk), .D(ctrlW[73]), .Q(n292), .QN( ));
Q_FDP0 U806 ( .CK(uclk), .D(ctrlW[74]), .Q(n291), .QN( ));
Q_FDP0 U807 ( .CK(uclk), .D(ctrlW[75]), .Q(n290), .QN( ));
Q_FDP0 U808 ( .CK(uclk), .D(ctrlW[76]), .Q(n289), .QN( ));
Q_FDP0 U809 ( .CK(uclk), .D(ctrlW[77]), .Q(n288), .QN( ));
Q_FDP0 U810 ( .CK(uclk), .D(ctrlW[78]), .Q(n287), .QN( ));
Q_FDP0 U811 ( .CK(uclk), .D(ctrlW[79]), .Q(n286), .QN( ));
Q_FDP0 U812 ( .CK(uclk), .D(ctrlW[80]), .Q(n285), .QN( ));
Q_FDP0 U813 ( .CK(uclk), .D(ctrlW[81]), .Q(n284), .QN( ));
Q_FDP0 U814 ( .CK(uclk), .D(ctrlW[82]), .Q(n283), .QN( ));
Q_FDP0 U815 ( .CK(uclk), .D(ctrlW[83]), .Q(n282), .QN( ));
Q_FDP0 U816 ( .CK(uclk), .D(ctrlW[84]), .Q(n281), .QN( ));
Q_FDP0 U817 ( .CK(uclk), .D(ctrlW[85]), .Q(n280), .QN( ));
Q_FDP0 U818 ( .CK(uclk), .D(ctrlW[86]), .Q(n279), .QN( ));
Q_FDP0 U819 ( .CK(uclk), .D(ctrlW[87]), .Q(n278), .QN( ));
Q_FDP0 U820 ( .CK(uclk), .D(ctrlW[88]), .Q(n277), .QN( ));
Q_FDP0 U821 ( .CK(uclk), .D(ctrlW[89]), .Q(n276), .QN( ));
Q_FDP0 U822 ( .CK(uclk), .D(ctrlW[90]), .Q(n275), .QN( ));
Q_FDP0 U823 ( .CK(uclk), .D(ctrlW[91]), .Q(n274), .QN( ));
Q_FDP0 U824 ( .CK(uclk), .D(ctrlW[92]), .Q(n273), .QN( ));
Q_FDP0 U825 ( .CK(uclk), .D(ctrlW[93]), .Q(n272), .QN( ));
Q_FDP0 U826 ( .CK(uclk), .D(ctrlW[94]), .Q(n271), .QN( ));
Q_FDP0 U827 ( .CK(uclk), .D(ctrlW[95]), .Q(n270), .QN( ));
Q_FDP0 U828 ( .CK(uclk), .D(ctrlW[96]), .Q(n269), .QN( ));
Q_FDP0 U829 ( .CK(uclk), .D(ctrlW[97]), .Q(n268), .QN( ));
Q_FDP0 U830 ( .CK(uclk), .D(ctrlW[98]), .Q(n267), .QN( ));
Q_FDP0 U831 ( .CK(uclk), .D(ctrlW[99]), .Q(n266), .QN( ));
Q_FDP0 U832 ( .CK(uclk), .D(ctrlW[100]), .Q(n265), .QN( ));
Q_FDP0 U833 ( .CK(uclk), .D(ctrlW[101]), .Q(n264), .QN( ));
Q_FDP0 U834 ( .CK(uclk), .D(ctrlW[102]), .Q(n263), .QN( ));
Q_FDP0 U835 ( .CK(uclk), .D(ctrlW[103]), .Q(n262), .QN( ));
Q_FDP0 U836 ( .CK(uclk), .D(ctrlW[104]), .Q(n261), .QN( ));
Q_FDP0 U837 ( .CK(uclk), .D(ctrlW[105]), .Q(n260), .QN( ));
Q_FDP0 U838 ( .CK(uclk), .D(ctrlW[106]), .Q(n259), .QN( ));
Q_FDP0 U839 ( .CK(uclk), .D(ctrlW[107]), .Q(n258), .QN( ));
Q_FDP0 U840 ( .CK(uclk), .D(ctrlW[108]), .Q(n257), .QN( ));
Q_FDP0 U841 ( .CK(uclk), .D(ctrlW[109]), .Q(n256), .QN( ));
Q_FDP0 U842 ( .CK(uclk), .D(ctrlW[110]), .Q(n255), .QN( ));
Q_FDP0 U843 ( .CK(uclk), .D(ctrlW[111]), .Q(n254), .QN( ));
Q_FDP0 U844 ( .CK(uclk), .D(ctrlW[112]), .Q(n253), .QN( ));
Q_FDP0 U845 ( .CK(uclk), .D(ctrlW[113]), .Q(n252), .QN( ));
Q_FDP0 U846 ( .CK(uclk), .D(ctrlW[114]), .Q(n251), .QN( ));
Q_FDP0 U847 ( .CK(uclk), .D(ctrlW[115]), .Q(n250), .QN( ));
Q_FDP0 U848 ( .CK(uclk), .D(ctrlW[116]), .Q(n249), .QN( ));
Q_FDP0 U849 ( .CK(uclk), .D(ctrlW[117]), .Q(n248), .QN( ));
Q_FDP0 U850 ( .CK(uclk), .D(ctrlW[118]), .Q(n247), .QN( ));
Q_FDP0 U851 ( .CK(uclk), .D(ctrlW[119]), .Q(n246), .QN( ));
Q_FDP0 U852 ( .CK(uclk), .D(ctrlW[120]), .Q(n245), .QN( ));
Q_FDP0 U853 ( .CK(uclk), .D(ctrlW[121]), .Q(n244), .QN( ));
Q_FDP0 U854 ( .CK(uclk), .D(ctrlW[122]), .Q(n243), .QN( ));
Q_FDP0 U855 ( .CK(uclk), .D(ctrlW[123]), .Q(n242), .QN( ));
Q_FDP0 U856 ( .CK(uclk), .D(ctrlW[124]), .Q(n241), .QN( ));
Q_FDP0 U857 ( .CK(uclk), .D(ctrlW[125]), .Q(n240), .QN( ));
Q_FDP0 U858 ( .CK(uclk), .D(ctrlW[126]), .Q(n239), .QN( ));
Q_FDP0 U859 ( .CK(uclk), .D(ctrlW[127]), .Q(n238), .QN( ));
Q_FDP0 U860 ( .CK(uclk), .D(ctrlW[128]), .Q(n237), .QN( ));
Q_FDP0 U861 ( .CK(uclk), .D(ctrlW[129]), .Q(n236), .QN( ));
Q_FDP0 U862 ( .CK(uclk), .D(ctrlW[130]), .Q(n235), .QN( ));
Q_FDP0 U863 ( .CK(uclk), .D(ctrlW[131]), .Q(n234), .QN( ));
Q_FDP0 U864 ( .CK(uclk), .D(ctrlW[132]), .Q(n233), .QN( ));
Q_FDP0 U865 ( .CK(uclk), .D(ctrlW[133]), .Q(n232), .QN( ));
Q_FDP0 U866 ( .CK(uclk), .D(ctrlW[134]), .Q(n231), .QN( ));
Q_FDP0 U867 ( .CK(uclk), .D(ctrlW[135]), .Q(n230), .QN( ));
Q_FDP0 U868 ( .CK(uclk), .D(ctrlW[136]), .Q(n229), .QN( ));
Q_FDP0 U869 ( .CK(uclk), .D(ctrlW[137]), .Q(n228), .QN( ));
Q_FDP0 U870 ( .CK(uclk), .D(ctrlW[138]), .Q(n227), .QN( ));
Q_FDP0 U871 ( .CK(uclk), .D(ctrlW[139]), .Q(n226), .QN( ));
Q_FDP0 U872 ( .CK(uclk), .D(ctrlW[140]), .Q(n225), .QN( ));
Q_FDP0 U873 ( .CK(uclk), .D(ctrlW[141]), .Q(n224), .QN( ));
Q_FDP0 U874 ( .CK(uclk), .D(ctrlW[142]), .Q(n223), .QN( ));
Q_FDP0 U875 ( .CK(uclk), .D(ctrlW[143]), .Q(n222), .QN( ));
Q_FDP0 U876 ( .CK(uclk), .D(ctrlW[144]), .Q(n221), .QN( ));
Q_FDP0 U877 ( .CK(uclk), .D(ctrlW[145]), .Q(n220), .QN( ));
Q_FDP0 U878 ( .CK(uclk), .D(ctrlW[146]), .Q(n219), .QN( ));
Q_FDP0 U879 ( .CK(uclk), .D(ctrlW[147]), .Q(n218), .QN( ));
Q_FDP0 U880 ( .CK(uclk), .D(ctrlW[148]), .Q(n217), .QN( ));
Q_FDP0 U881 ( .CK(uclk), .D(ctrlW[149]), .Q(n216), .QN( ));
Q_FDP0 U882 ( .CK(uclk), .D(ctrlW[150]), .Q(n215), .QN( ));
Q_FDP0 U883 ( .CK(uclk), .D(ctrlW[151]), .Q(n214), .QN( ));
Q_FDP0 U884 ( .CK(uclk), .D(ctrlW[152]), .Q(n213), .QN( ));
Q_FDP0 U885 ( .CK(uclk), .D(ctrlW[153]), .Q(n212), .QN( ));
Q_FDP0 U886 ( .CK(uclk), .D(ctrlW[154]), .Q(n211), .QN( ));
Q_FDP0 U887 ( .CK(uclk), .D(ctrlW[155]), .Q(n210), .QN( ));
Q_FDP0 U888 ( .CK(uclk), .D(ctrlW[156]), .Q(n209), .QN( ));
Q_FDP0 U889 ( .CK(uclk), .D(ctrlW[157]), .Q(n208), .QN( ));
Q_FDP0 U890 ( .CK(uclk), .D(ctrlW[158]), .Q(n207), .QN( ));
Q_FDP0 U891 ( .CK(uclk), .D(ctrlW[159]), .Q(n206), .QN( ));
Q_FDP0 U892 ( .CK(uclk), .D(ctrlW[160]), .Q(n205), .QN( ));
Q_FDP0 U893 ( .CK(uclk), .D(ctrlW[161]), .Q(n204), .QN( ));
Q_FDP0 U894 ( .CK(uclk), .D(ctrlW[162]), .Q(n203), .QN( ));
Q_FDP0 U895 ( .CK(uclk), .D(ctrlW[163]), .Q(n202), .QN( ));
Q_FDP0 U896 ( .CK(uclk), .D(ctrlW[164]), .Q(n201), .QN( ));
Q_FDP0 U897 ( .CK(uclk), .D(ctrlW[165]), .Q(n200), .QN( ));
Q_FDP0 U898 ( .CK(uclk), .D(ctrlW[166]), .Q(n199), .QN( ));
Q_FDP0 U899 ( .CK(uclk), .D(ctrlW[167]), .Q(n198), .QN( ));
Q_FDP0 U900 ( .CK(uclk), .D(ctrlW[168]), .Q(n197), .QN( ));
Q_FDP0 U901 ( .CK(uclk), .D(ctrlW[169]), .Q(n196), .QN( ));
Q_FDP0 U902 ( .CK(uclk), .D(ctrlW[170]), .Q(n195), .QN( ));
Q_FDP0 U903 ( .CK(uclk), .D(ctrlW[171]), .Q(n194), .QN( ));
Q_FDP0 U904 ( .CK(uclk), .D(ctrlW[172]), .Q(n193), .QN( ));
Q_FDP0 U905 ( .CK(uclk), .D(ctrlW[173]), .Q(n192), .QN( ));
Q_FDP0 U906 ( .CK(uclk), .D(ctrlW[174]), .Q(n191), .QN( ));
Q_FDP0 U907 ( .CK(uclk), .D(ctrlW[175]), .Q(n190), .QN( ));
Q_FDP0 U908 ( .CK(uclk), .D(ctrlW[176]), .Q(n189), .QN( ));
Q_FDP0 U909 ( .CK(uclk), .D(ctrlW[177]), .Q(n188), .QN( ));
Q_FDP0 U910 ( .CK(uclk), .D(ctrlW[178]), .Q(n187), .QN( ));
Q_FDP0 U911 ( .CK(uclk), .D(ctrlW[179]), .Q(n186), .QN( ));
Q_FDP0 U912 ( .CK(uclk), .D(ctrlW[180]), .Q(n185), .QN( ));
Q_FDP0 U913 ( .CK(uclk), .D(ctrlW[181]), .Q(n184), .QN( ));
Q_FDP0 U914 ( .CK(uclk), .D(ctrlW[182]), .Q(n183), .QN( ));
Q_FDP0 U915 ( .CK(uclk), .D(ctrlW[183]), .Q(n182), .QN( ));
Q_FDP0 U916 ( .CK(uclk), .D(ctrlW[184]), .Q(n181), .QN( ));
Q_FDP0 U917 ( .CK(uclk), .D(ctrlW[185]), .Q(n180), .QN( ));
Q_FDP0 U918 ( .CK(uclk), .D(ctrlW[186]), .Q(n179), .QN( ));
Q_FDP0 U919 ( .CK(uclk), .D(ctrlW[187]), .Q(n178), .QN( ));
Q_FDP0 U920 ( .CK(uclk), .D(ctrlW[188]), .Q(n177), .QN( ));
Q_FDP0 U921 ( .CK(uclk), .D(ctrlW[189]), .Q(n176), .QN( ));
Q_FDP0 U922 ( .CK(uclk), .D(ctrlW[190]), .Q(n175), .QN( ));
Q_FDP0 U923 ( .CK(uclk), .D(ctrlW[191]), .Q(n174), .QN( ));
Q_FDP0 U924 ( .CK(uclk), .D(ctrlW[192]), .Q(n173), .QN( ));
Q_FDP0 U925 ( .CK(uclk), .D(ctrlW[193]), .Q(n172), .QN( ));
Q_FDP0 U926 ( .CK(uclk), .D(ctrlW[194]), .Q(n171), .QN( ));
Q_FDP0 U927 ( .CK(uclk), .D(ctrlW[195]), .Q(n170), .QN( ));
Q_FDP0 U928 ( .CK(uclk), .D(ctrlW[196]), .Q(n169), .QN( ));
Q_FDP0 U929 ( .CK(uclk), .D(ctrlW[197]), .Q(n168), .QN( ));
Q_FDP0 U930 ( .CK(uclk), .D(ctrlW[198]), .Q(n167), .QN( ));
Q_FDP0 U931 ( .CK(uclk), .D(ctrlW[199]), .Q(n166), .QN( ));
Q_FDP0 U932 ( .CK(uclk), .D(ctrlW[200]), .Q(n165), .QN( ));
Q_FDP0 U933 ( .CK(uclk), .D(ctrlW[201]), .Q(n164), .QN( ));
Q_FDP0 U934 ( .CK(uclk), .D(ctrlW[202]), .Q(n163), .QN( ));
Q_FDP0 U935 ( .CK(uclk), .D(ctrlW[203]), .Q(n162), .QN( ));
Q_FDP0 U936 ( .CK(uclk), .D(ctrlW[204]), .Q(n161), .QN( ));
Q_FDP0 U937 ( .CK(uclk), .D(ctrlW[205]), .Q(n160), .QN( ));
Q_FDP0 U938 ( .CK(uclk), .D(ctrlW[206]), .Q(n159), .QN( ));
Q_FDP0 U939 ( .CK(uclk), .D(ctrlW[207]), .Q(n158), .QN( ));
Q_FDP0 U940 ( .CK(uclk), .D(ctrlW[208]), .Q(n157), .QN( ));
Q_FDP0 U941 ( .CK(uclk), .D(ctrlW[209]), .Q(n156), .QN( ));
Q_FDP0 U942 ( .CK(uclk), .D(ctrlW[210]), .Q(n155), .QN( ));
Q_FDP0 U943 ( .CK(uclk), .D(ctrlW[211]), .Q(n154), .QN( ));
Q_FDP0 U944 ( .CK(uclk), .D(ctrlW[212]), .Q(n153), .QN( ));
Q_FDP0 U945 ( .CK(uclk), .D(ctrlW[213]), .Q(n152), .QN( ));
Q_FDP0 U946 ( .CK(uclk), .D(ctrlW[214]), .Q(n151), .QN( ));
Q_FDP0 U947 ( .CK(uclk), .D(ctrlW[215]), .Q(n150), .QN( ));
Q_FDP0 U948 ( .CK(uclk), .D(ctrlW[216]), .Q(n149), .QN( ));
Q_FDP0 U949 ( .CK(uclk), .D(ctrlW[217]), .Q(n148), .QN( ));
Q_FDP0 U950 ( .CK(uclk), .D(ctrlW[218]), .Q(n147), .QN( ));
Q_FDP0 U951 ( .CK(uclk), .D(ctrlW[219]), .Q(n146), .QN( ));
Q_FDP0 U952 ( .CK(uclk), .D(ctrlW[220]), .Q(n145), .QN( ));
Q_FDP0 U953 ( .CK(uclk), .D(ctrlW[221]), .Q(n144), .QN( ));
Q_FDP0 U954 ( .CK(uclk), .D(ctrlW[222]), .Q(n143), .QN( ));
Q_FDP0 U955 ( .CK(uclk), .D(ctrlW[223]), .Q(n142), .QN( ));
Q_FDP0 U956 ( .CK(uclk), .D(ctrlW[224]), .Q(n141), .QN( ));
Q_FDP0 U957 ( .CK(uclk), .D(ctrlW[225]), .Q(n140), .QN( ));
Q_FDP0 U958 ( .CK(uclk), .D(ctrlW[226]), .Q(n139), .QN( ));
Q_FDP0 U959 ( .CK(uclk), .D(ctrlW[227]), .Q(n138), .QN( ));
Q_FDP0 U960 ( .CK(uclk), .D(ctrlW[228]), .Q(n137), .QN( ));
Q_FDP0 U961 ( .CK(uclk), .D(ctrlW[229]), .Q(n136), .QN( ));
Q_FDP0 U962 ( .CK(uclk), .D(ctrlW[230]), .Q(n135), .QN( ));
Q_FDP0 U963 ( .CK(uclk), .D(ctrlW[231]), .Q(n134), .QN( ));
Q_FDP0 U964 ( .CK(uclk), .D(ctrlW[232]), .Q(n133), .QN( ));
Q_FDP0 U965 ( .CK(uclk), .D(ctrlW[233]), .Q(n132), .QN( ));
Q_FDP0 U966 ( .CK(uclk), .D(ctrlW[234]), .Q(n131), .QN( ));
Q_FDP0 U967 ( .CK(uclk), .D(ctrlW[235]), .Q(n130), .QN( ));
Q_FDP0 U968 ( .CK(uclk), .D(ctrlW[236]), .Q(n129), .QN( ));
Q_FDP0 U969 ( .CK(uclk), .D(ctrlW[237]), .Q(n128), .QN( ));
Q_FDP0 U970 ( .CK(uclk), .D(ctrlW[238]), .Q(n127), .QN( ));
Q_FDP0 U971 ( .CK(uclk), .D(ctrlW[239]), .Q(n126), .QN( ));
Q_FDP0 U972 ( .CK(uclk), .D(ctrlW[240]), .Q(n125), .QN( ));
Q_FDP0 U973 ( .CK(uclk), .D(ctrlW[241]), .Q(n124), .QN( ));
Q_FDP0 U974 ( .CK(uclk), .D(ctrlW[242]), .Q(n123), .QN( ));
Q_FDP0 U975 ( .CK(uclk), .D(ctrlW[243]), .Q(n122), .QN( ));
Q_FDP0 U976 ( .CK(uclk), .D(ctrlW[244]), .Q(n121), .QN( ));
Q_FDP0 U977 ( .CK(uclk), .D(ctrlW[245]), .Q(n120), .QN( ));
Q_FDP0 U978 ( .CK(uclk), .D(ctrlW[246]), .Q(n119), .QN( ));
Q_FDP0 U979 ( .CK(uclk), .D(ctrlW[247]), .Q(n118), .QN( ));
Q_FDP0 U980 ( .CK(uclk), .D(ctrlW[248]), .Q(n117), .QN( ));
Q_FDP0 U981 ( .CK(uclk), .D(ctrlW[249]), .Q(n116), .QN( ));
Q_FDP0 U982 ( .CK(uclk), .D(ctrlW[250]), .Q(n115), .QN( ));
Q_FDP0 U983 ( .CK(uclk), .D(ctrlW[251]), .Q(n114), .QN( ));
Q_FDP0 U984 ( .CK(uclk), .D(ctrlW[252]), .Q(n113), .QN( ));
Q_FDP0 U985 ( .CK(uclk), .D(ctrlW[253]), .Q(n112), .QN( ));
Q_FDP0 U986 ( .CK(uclk), .D(ctrlW[254]), .Q(n111), .QN( ));
Q_FDP0 U987 ( .CK(uclk), .D(ctrlW[255]), .Q(n110), .QN( ));
`ifdef CBV

reg [255:0] ctrl [0:3];
initial begin: U988
  integer i;
  for (i=0; i<=3; i=i+1) ctrl[i] =
`ifdef CBV_MEM_INIT1
  {256{1'b1}};
`else
  256'b0;
`endif
end
reg [255:0] n792;
assign {n788, n787, n786, n785, n784, n783, n782,
n781, n780, n779, n778, n777, n776, n775, n774,
n773, n772, n771, n770, n769, n768, n767, n766,
n765, n764, n763, n762, n761, n760, n759, n758,
n757, n756, n755, n754, n753, n752, n751, n750,
n749, n748, n747, n746, n745, n744, n743, n742,
n741, n740, n739, n738, n737, n736, n735, n734,
n733, n732, n731, n730, n729, n728, n727, n726,
n725, n724, n723, n722, n721, n720, n719, n718,
n717, n716, n715, n714, n713, n712, n711, n710,
n709, n708, n707, n706, n705, n704, n703, n702,
n701, n700, n699, n698, n697, n696, n695, n694,
n693, n692, n691, n690, n689, n688, n687, n686,
n685, n684, n683, n682, n681, n680, n679, n678,
n677, n676, n675, n674, n673, n672, n671, n670,
n669, n668, n667, n666, n665, n664, n663, n662,
n661, n660, n659, n658, n657, n656, n655, n654,
n653, n652, n651, n650, n649, n648, n647, n646,
n645, n644, n643, n642, n641, n640, n639, n638,
n637, n636, n635, n634, n633, n632, n631, n630,
n629, n628, n627, n626, n625, n624, n623, n622,
n621, n620, n619, n618, n617, n616, n615, n614,
n613, n612, n611, n610, n609, n608, n607, n606,
n605, n604, n603, n602, n601, n600, n599, n598,
n597, n596, n595, n594, n593, n592, n591, n590,
n589, n588, n587, n586, n585, n584, n583, n582,
n581, n580, n579, n578, n577, n576, n575, n574,
n573, n572, n571, n570, n569, n568, n567, n566,
n565, n564, n563, n562, n561, n560, n559, n558,
n557, n556, n555, n554, n553, n552, n551, n550,
n549, n548, n547, n546, n545, n544, n543, n542,
n541, n540, n539, n538, n537, n536, n535, n534,
n533} = n792; 
always @(n532 or n110 or n111 or n112 or n113
 or n114 or n115 or n116 or n117 or n118 or n119 or n120 or n121
 or n122 or n123 or n124 or n125 or n126 or n127 or n128 or n129
 or n130 or n131 or n132 or n133 or n134 or n135 or n136 or n137
 or n138 or n139 or n140 or n141 or n142 or n143 or n144 or n145
 or n146 or n147 or n148 or n149 or n150 or n151 or n152 or n153
 or n154 or n155 or n156 or n157 or n158 or n159 or n160 or n161
 or n162 or n163 or n164 or n165 or n166 or n167 or n168 or n169
 or n170 or n171 or n172 or n173 or n174 or n175 or n176 or n177
 or n178 or n179 or n180 or n181 or n182 or n183 or n184 or n185
 or n186 or n187 or n188 or n189 or n190 or n191 or n192 or n193
 or n194 or n195 or n196 or n197 or n198 or n199 or n200 or n201
 or n202 or n203 or n204 or n205 or n206 or n207 or n208 or n209
 or n210 or n211 or n212 or n213 or n214 or n215 or n216 or n217
 or n218 or n219 or n220 or n221 or n222 or n223 or n224 or n225
 or n226 or n227 or n228 or n229 or n230 or n231 or n232 or n233
 or n234 or n235 or n236 or n237 or n238 or n239 or n240 or n241
 or n242 or n243 or n244 or n245 or n246 or n247 or n248 or n249
 or n250 or n251 or n252 or n253 or n254 or n255 or n256 or n257
 or n258 or n259 or n260 or n261 or n262 or n263 or n264 or n265
 or n266 or n267 or n268 or n269 or n270 or n271 or n272 or n273
 or n274 or n275 or n276 or n277 or n278 or n279 or n280 or n281
 or n282 or n283 or n284 or n285 or n286 or n287 or n288 or n289
 or n290 or n291 or n292 or n293 or n294 or n295 or n296 or n297
 or n298 or n299 or n300 or n301 or n302 or n303 or n304 or n305
 or n306 or n307 or n308 or n309 or n310 or n311 or n312 or n313
 or n314 or n315 or n316 or n317 or n318 or n319 or n320 or n321
 or n322 or n323 or n324 or n325 or n326 or n327 or n328 or n329
 or n330 or n331 or n332 or n333 or n334 or n335 or n336 or n337
 or n338 or n339 or n340 or n341 or n342 or n343 or n344 or n345
 or n346 or n347 or n348 or n349 or n350 or n351 or n352 or n353
 or n354 or n355 or n356 or n357 or n358 or n359 or n360 or n361
 or n362 or n363 or n364 or n365 or n366 or n370)
#0 begin
if (n366)
ctrl[{n532, n532}] =
{n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177, n178,
 n179, n180, n181, n182, n183, n184, n185, n186,
 n187, n188, n189, n190, n191, n192, n193, n194,
 n195, n196, n197, n198, n199, n200, n201, n202,
 n203, n204, n205, n206, n207, n208, n209, n210,
 n211, n212, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365};
n792 = ctrl[{n532, n370}];
end
`else

MPW4X256 ctrl ( .A1(n532), .A0(n532), .DI255(n110), .DI254(n111), .DI253(n112), .DI252(n113),
 .DI251(n114), .DI250(n115), .DI249(n116), .DI248(n117), .DI247(n118), .DI246(n119), .DI245(n120), .DI244(n121),
 .DI243(n122), .DI242(n123), .DI241(n124), .DI240(n125), .DI239(n126), .DI238(n127), .DI237(n128), .DI236(n129),
 .DI235(n130), .DI234(n131), .DI233(n132), .DI232(n133), .DI231(n134), .DI230(n135), .DI229(n136), .DI228(n137),
 .DI227(n138), .DI226(n139), .DI225(n140), .DI224(n141), .DI223(n142), .DI222(n143), .DI221(n144), .DI220(n145),
 .DI219(n146), .DI218(n147), .DI217(n148), .DI216(n149), .DI215(n150), .DI214(n151), .DI213(n152), .DI212(n153),
 .DI211(n154), .DI210(n155), .DI209(n156), .DI208(n157), .DI207(n158), .DI206(n159), .DI205(n160), .DI204(n161),
 .DI203(n162), .DI202(n163), .DI201(n164), .DI200(n165), .DI199(n166), .DI198(n167), .DI197(n168), .DI196(n169),
 .DI195(n170), .DI194(n171), .DI193(n172), .DI192(n173), .DI191(n174), .DI190(n175), .DI189(n176), .DI188(n177),
 .DI187(n178), .DI186(n179), .DI185(n180), .DI184(n181), .DI183(n182), .DI182(n183), .DI181(n184), .DI180(n185),
 .DI179(n186), .DI178(n187), .DI177(n188), .DI176(n189), .DI175(n190), .DI174(n191), .DI173(n192), .DI172(n193),
 .DI171(n194), .DI170(n195), .DI169(n196), .DI168(n197), .DI167(n198), .DI166(n199), .DI165(n200), .DI164(n201),
 .DI163(n202), .DI162(n203), .DI161(n204), .DI160(n205), .DI159(n206), .DI158(n207), .DI157(n208), .DI156(n209),
 .DI155(n210), .DI154(n211), .DI153(n212), .DI152(n213), .DI151(n214), .DI150(n215), .DI149(n216), .DI148(n217),
 .DI147(n218), .DI146(n219), .DI145(n220), .DI144(n221), .DI143(n222), .DI142(n223), .DI141(n224), .DI140(n225),
 .DI139(n226), .DI138(n227), .DI137(n228), .DI136(n229), .DI135(n230), .DI134(n231), .DI133(n232), .DI132(n233),
 .DI131(n234), .DI130(n235), .DI129(n236), .DI128(n237), .DI127(n238), .DI126(n239), .DI125(n240), .DI124(n241),
 .DI123(n242), .DI122(n243), .DI121(n244), .DI120(n245), .DI119(n246), .DI118(n247), .DI117(n248), .DI116(n249),
 .DI115(n250), .DI114(n251), .DI113(n252), .DI112(n253), .DI111(n254), .DI110(n255), .DI109(n256), .DI108(n257),
 .DI107(n258), .DI106(n259), .DI105(n260), .DI104(n261), .DI103(n262), .DI102(n263), .DI101(n264), .DI100(n265),
 .DI99(n266), .DI98(n267), .DI97(n268), .DI96(n269), .DI95(n270), .DI94(n271), .DI93(n272), .DI92(n273),
 .DI91(n274), .DI90(n275), .DI89(n276), .DI88(n277), .DI87(n278), .DI86(n279), .DI85(n280), .DI84(n281),
 .DI83(n282), .DI82(n283), .DI81(n284), .DI80(n285), .DI79(n286), .DI78(n287), .DI77(n288), .DI76(n289),
 .DI75(n290), .DI74(n291), .DI73(n292), .DI72(n293), .DI71(n294), .DI70(n295), .DI69(n296), .DI68(n297),
 .DI67(n298), .DI66(n299), .DI65(n300), .DI64(n301), .DI63(n302), .DI62(n303), .DI61(n304), .DI60(n305),
 .DI59(n306), .DI58(n307), .DI57(n308), .DI56(n309), .DI55(n310), .DI54(n311), .DI53(n312), .DI52(n313),
 .DI51(n314), .DI50(n315), .DI49(n316), .DI48(n317), .DI47(n318), .DI46(n319), .DI45(n320), .DI44(n321),
 .DI43(n322), .DI42(n323), .DI41(n324), .DI40(n325), .DI39(n326), .DI38(n327), .DI37(n328), .DI36(n329),
 .DI35(n330), .DI34(n331), .DI33(n332), .DI32(n333), .DI31(n334), .DI30(n335), .DI29(n336), .DI28(n337),
 .DI27(n338), .DI26(n339), .DI25(n340), .DI24(n341), .DI23(n342), .DI22(n343), .DI21(n344), .DI20(n345),
 .DI19(n346), .DI18(n347), .DI17(n348), .DI16(n349), .DI15(n350), .DI14(n351), .DI13(n352), .DI12(n353),
 .DI11(n354), .DI10(n355), .DI9(n356), .DI8(n357), .DI7(n358), .DI6(n359), .DI5(n360), .DI4(n361),
 .DI3(n362), .DI2(n363), .DI1(n364), .DI0(n365), .WE(n366), .SYNC_IN(n532), .SYNC_OUT(n792));
// pragma CVASTRPROP INSTANCE "ctrl" HDL_MEMORY_DECL "1 255 0 0 3"
MPR4X256 U989 ( .A1(n532), .A0(n370), .SYNC_IN(n792), .DO255(n788), .DO254(n787), .DO253(n786),
 .DO252(n785), .DO251(n784), .DO250(n783), .DO249(n782), .DO248(n781), .DO247(n780), .DO246(n779), .DO245(n778),
 .DO244(n777), .DO243(n776), .DO242(n775), .DO241(n774), .DO240(n773), .DO239(n772), .DO238(n771), .DO237(n770),
 .DO236(n769), .DO235(n768), .DO234(n767), .DO233(n766), .DO232(n765), .DO231(n764), .DO230(n763), .DO229(n762),
 .DO228(n761), .DO227(n760), .DO226(n759), .DO225(n758), .DO224(n757), .DO223(n756), .DO222(n755), .DO221(n754),
 .DO220(n753), .DO219(n752), .DO218(n751), .DO217(n750), .DO216(n749), .DO215(n748), .DO214(n747), .DO213(n746),
 .DO212(n745), .DO211(n744), .DO210(n743), .DO209(n742), .DO208(n741), .DO207(n740), .DO206(n739), .DO205(n738),
 .DO204(n737), .DO203(n736), .DO202(n735), .DO201(n734), .DO200(n733), .DO199(n732), .DO198(n731), .DO197(n730),
 .DO196(n729), .DO195(n728), .DO194(n727), .DO193(n726), .DO192(n725), .DO191(n724), .DO190(n723), .DO189(n722),
 .DO188(n721), .DO187(n720), .DO186(n719), .DO185(n718), .DO184(n717), .DO183(n716), .DO182(n715), .DO181(n714),
 .DO180(n713), .DO179(n712), .DO178(n711), .DO177(n710), .DO176(n709), .DO175(n708), .DO174(n707), .DO173(n706),
 .DO172(n705), .DO171(n704), .DO170(n703), .DO169(n702), .DO168(n701), .DO167(n700), .DO166(n699), .DO165(n698),
 .DO164(n697), .DO163(n696), .DO162(n695), .DO161(n694), .DO160(n693), .DO159(n692), .DO158(n691), .DO157(n690),
 .DO156(n689), .DO155(n688), .DO154(n687), .DO153(n686), .DO152(n685), .DO151(n684), .DO150(n683), .DO149(n682),
 .DO148(n681), .DO147(n680), .DO146(n679), .DO145(n678), .DO144(n677), .DO143(n676), .DO142(n675), .DO141(n674),
 .DO140(n673), .DO139(n672), .DO138(n671), .DO137(n670), .DO136(n669), .DO135(n668), .DO134(n667), .DO133(n666),
 .DO132(n665), .DO131(n664), .DO130(n663), .DO129(n662), .DO128(n661), .DO127(n660), .DO126(n659), .DO125(n658),
 .DO124(n657), .DO123(n656), .DO122(n655), .DO121(n654), .DO120(n653), .DO119(n652), .DO118(n651), .DO117(n650),
 .DO116(n649), .DO115(n648), .DO114(n647), .DO113(n646), .DO112(n645), .DO111(n644), .DO110(n643), .DO109(n642),
 .DO108(n641), .DO107(n640), .DO106(n639), .DO105(n638), .DO104(n637), .DO103(n636), .DO102(n635), .DO101(n634),
 .DO100(n633), .DO99(n632), .DO98(n631), .DO97(n630), .DO96(n629), .DO95(n628), .DO94(n627), .DO93(n626),
 .DO92(n625), .DO91(n624), .DO90(n623), .DO89(n622), .DO88(n621), .DO87(n620), .DO86(n619), .DO85(n618),
 .DO84(n617), .DO83(n616), .DO82(n615), .DO81(n614), .DO80(n613), .DO79(n612), .DO78(n611), .DO77(n610),
 .DO76(n609), .DO75(n608), .DO74(n607), .DO73(n606), .DO72(n605), .DO71(n604), .DO70(n603), .DO69(n602),
 .DO68(n601), .DO67(n600), .DO66(n599), .DO65(n598), .DO64(n597), .DO63(n596), .DO62(n595), .DO61(n594),
 .DO60(n593), .DO59(n592), .DO58(n591), .DO57(n590), .DO56(n589), .DO55(n588), .DO54(n587), .DO53(n586),
 .DO52(n585), .DO51(n584), .DO50(n583), .DO49(n582), .DO48(n581), .DO47(n580), .DO46(n579), .DO45(n578),
 .DO44(n577), .DO43(n576), .DO42(n575), .DO41(n574), .DO40(n573), .DO39(n572), .DO38(n571), .DO37(n570),
 .DO36(n569), .DO35(n568), .DO34(n567), .DO33(n566), .DO32(n565), .DO31(n564), .DO30(n563), .DO29(n562),
 .DO28(n561), .DO27(n560), .DO26(n559), .DO25(n558), .DO24(n557), .DO23(n556), .DO22(n555), .DO21(n554),
 .DO20(n553), .DO19(n552), .DO18(n551), .DO17(n550), .DO16(n549), .DO15(n548), .DO14(n547), .DO13(n546),
 .DO12(n545), .DO11(n544), .DO10(n543), .DO9(n542), .DO8(n541), .DO7(n540), .DO6(n539), .DO5(n538),
 .DO4(n537), .DO3(n536), .DO2(n535), .DO1(n534), .DO0(n533), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "ctrl 1 255 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW4X256_MPR4X256
`else
module MPW4X256( A1, A0, DI255, DI254, DI253, DI252, DI251,
 DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227,
 DI226, DI225, DI224, DI223, DI222, DI221, DI220, DI219,
 DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211,
 DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187,
 DI186, DI185, DI184, DI183, DI182, DI181, DI180, DI179,
 DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171,
 DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147,
 DI146, DI145, DI144, DI143, DI142, DI141, DI140, DI139,
 DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131,
 DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107,
 DI106, DI105, DI104, DI103, DI102, DI101, DI100, DI99,
 DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91,
 DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67,
 DI66, DI65, DI64, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A1, A0, DI255, DI254, DI253, DI252, DI251, DI250,
 DI249, DI248, DI247, DI246, DI245, DI244, DI243, DI242, DI241, DI240,
 DI239, DI238, DI237, DI236, DI235, DI234, DI233, DI232, DI231, DI230,
 DI229, DI228, DI227, DI226, DI225, DI224, DI223, DI222, DI221, DI220,
 DI219, DI218, DI217, DI216, DI215, DI214, DI213, DI212, DI211, DI210,
 DI209, DI208, DI207, DI206, DI205, DI204, DI203, DI202, DI201, DI200,
 DI199, DI198, DI197, DI196, DI195, DI194, DI193, DI192, DI191, DI190,
 DI189, DI188, DI187, DI186, DI185, DI184, DI183, DI182, DI181, DI180,
 DI179, DI178, DI177, DI176, DI175, DI174, DI173, DI172, DI171, DI170,
 DI169, DI168, DI167, DI166, DI165, DI164, DI163, DI162, DI161, DI160,
 DI159, DI158, DI157, DI156, DI155, DI154, DI153, DI152, DI151, DI150,
 DI149, DI148, DI147, DI146, DI145, DI144, DI143, DI142, DI141, DI140,
 DI139, DI138, DI137, DI136, DI135, DI134, DI133, DI132, DI131, DI130,
 DI129, DI128, DI127, DI126, DI125, DI124, DI123, DI122, DI121, DI120,
 DI119, DI118, DI117, DI116, DI115, DI114, DI113, DI112, DI111, DI110,
 DI109, DI108, DI107, DI106, DI105, DI104, DI103, DI102, DI101, DI100,
 DI99, DI98, DI97, DI96, DI95, DI94, DI93, DI92, DI91, DI90,
 DI89, DI88, DI87, DI86, DI85, DI84, DI83, DI82, DI81, DI80,
 DI79, DI78, DI77, DI76, DI75, DI74, DI73, DI72, DI71, DI70,
 DI69, DI68, DI67, DI66, DI65, DI64, DI63, DI62, DI61, DI60,
 DI59, DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20,
 DI19, DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X256_
`else
module MPR4X256( A1, A0, SYNC_IN, DO255, DO254, DO253, DO252,
 DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236,
 DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220,
 DO219, DO218, DO217, DO216, DO215, DO214, DO213, DO212,
 DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196,
 DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180,
 DO179, DO178, DO177, DO176, DO175, DO174, DO173, DO172,
 DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156,
 DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140,
 DO139, DO138, DO137, DO136, DO135, DO134, DO133, DO132,
 DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116,
 DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100,
 DO99, DO98, DO97, DO96, DO95, DO94, DO93, DO92,
 DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76,
 DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60,
 DO59, DO58, DO57, DO56, DO55, DO54, DO53, DO52,
 DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12,
 DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO255, DO254, DO253, DO252, DO251, DO250, DO249, DO248,
 DO247, DO246, DO245, DO244, DO243, DO242, DO241, DO240, DO239, DO238,
 DO237, DO236, DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220, DO219, DO218,
 DO217, DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209, DO208,
 DO207, DO206, DO205, DO204, DO203, DO202, DO201, DO200, DO199, DO198,
 DO197, DO196, DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180, DO179, DO178,
 DO177, DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169, DO168,
 DO167, DO166, DO165, DO164, DO163, DO162, DO161, DO160, DO159, DO158,
 DO157, DO156, DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140, DO139, DO138,
 DO137, DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129, DO128,
 DO127, DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119, DO118,
 DO117, DO116, DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99, DO98,
 DO97, DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89, DO88,
 DO87, DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79, DO78,
 DO77, DO76, DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59, DO58,
 DO57, DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48,
 DO47, DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18,
 DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8,
 DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X256_
`endif
`define MPW4X256_MPR4X256
`endif
`endif
