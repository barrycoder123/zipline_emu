
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_kdf_merger ( kdf_cmdfifo_ack, sha_tag_stall, 
	merger_keyfifo_ack, kdf_keybuilder_data, kdf_keybuilder_valid, clk, 
	rst_n, cmdfifo_kdf_valid, .cmdfifo_kdf_cmd( {
	\cmdfifo_kdf_cmd.kdf_dek_iter [0], \cmdfifo_kdf_cmd.combo_mode [0], 
	\cmdfifo_kdf_cmd.dek_key_op [0], \cmdfifo_kdf_cmd.dak_key_op [0]} ), 
	sha_tag_data, sha_tag_valid, sha_tag_last, keyfifo_merger_data, 
	keyfifo_merger_valid, keybuilder_kdf_stall);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output kdf_cmdfifo_ack;
output sha_tag_stall;
output merger_keyfifo_ack;
output [63:0] kdf_keybuilder_data;
output kdf_keybuilder_valid;
input clk;
input rst_n;
input cmdfifo_kdf_valid;
input [0:0] \cmdfifo_kdf_cmd.kdf_dek_iter ;
input [0:0] \cmdfifo_kdf_cmd.combo_mode ;
input [0:0] \cmdfifo_kdf_cmd.dek_key_op ;
input [0:0] \cmdfifo_kdf_cmd.dak_key_op ;
wire [3:0] cmdfifo_kdf_cmd;
input [127:0] sha_tag_data;
input sha_tag_valid;
input sha_tag_last;
input [127:0] keyfifo_merger_data;
input keyfifo_merger_valid;
input keybuilder_kdf_stall;
wire fifo_in_stall;
wire [127:0] fifo_out;
wire fifo_out_vld;
wire _zy_simnet_kdf_cmdfifo_ack_0_w$;
wire _zy_simnet_sha_tag_stall_1_w$;
wire _zy_simnet_merger_keyfifo_ack_2_w$;
wire [0:63] _zy_simnet_kdf_keybuilder_data_3_w$;
wire _zy_simnet_kdf_keybuilder_valid_4_w$;
wire _zy_simnet_dio_5;
wire _zy_simnet_dio_6;
wire [0:127] _zy_simnet_fifo_in_7_w$;
wire _zy_simnet_fifo_in_vld_8_w$;
wire _zy_simnet_fifo_out_ack_9_w$;
wire _zy_simnet_cio_10;
wire [127:0] fifo_in;
wire fifo_in_vld;
wire fifo_out_ack;
wire [2:0] in_counter;
wire out_counter;
supply0 n1;
tran (cmdfifo_kdf_cmd[3], \cmdfifo_kdf_cmd.kdf_dek_iter [0]);
tran (cmdfifo_kdf_cmd[2], \cmdfifo_kdf_cmd.combo_mode [0]);
tran (cmdfifo_kdf_cmd[1], \cmdfifo_kdf_cmd.dek_key_op [0]);
tran (cmdfifo_kdf_cmd[0], \cmdfifo_kdf_cmd.dak_key_op [0]);
Q_BUF U0 ( .A(n1), .Z(_zy_simnet_cio_10));
Q_INV U1 ( .A(keybuilder_kdf_stall), .Z(n2));
Q_AN02 U2 ( .A0(n2), .A1(fifo_out_vld), .Z(kdf_keybuilder_valid));
Q_AN02 U3 ( .A0(kdf_keybuilder_valid), .A1(n3), .Z(kdf_keybuilder_data[63]));
Q_AN02 U4 ( .A0(kdf_keybuilder_valid), .A1(n4), .Z(kdf_keybuilder_data[62]));
Q_AN02 U5 ( .A0(kdf_keybuilder_valid), .A1(n5), .Z(kdf_keybuilder_data[61]));
Q_AN02 U6 ( .A0(kdf_keybuilder_valid), .A1(n6), .Z(kdf_keybuilder_data[60]));
Q_AN02 U7 ( .A0(kdf_keybuilder_valid), .A1(n7), .Z(kdf_keybuilder_data[59]));
Q_AN02 U8 ( .A0(kdf_keybuilder_valid), .A1(n8), .Z(kdf_keybuilder_data[58]));
Q_AN02 U9 ( .A0(kdf_keybuilder_valid), .A1(n9), .Z(kdf_keybuilder_data[57]));
Q_AN02 U10 ( .A0(kdf_keybuilder_valid), .A1(n10), .Z(kdf_keybuilder_data[56]));
Q_AN02 U11 ( .A0(kdf_keybuilder_valid), .A1(n11), .Z(kdf_keybuilder_data[55]));
Q_AN02 U12 ( .A0(kdf_keybuilder_valid), .A1(n12), .Z(kdf_keybuilder_data[54]));
Q_AN02 U13 ( .A0(kdf_keybuilder_valid), .A1(n13), .Z(kdf_keybuilder_data[53]));
Q_AN02 U14 ( .A0(kdf_keybuilder_valid), .A1(n14), .Z(kdf_keybuilder_data[52]));
Q_AN02 U15 ( .A0(kdf_keybuilder_valid), .A1(n15), .Z(kdf_keybuilder_data[51]));
Q_AN02 U16 ( .A0(kdf_keybuilder_valid), .A1(n16), .Z(kdf_keybuilder_data[50]));
Q_AN02 U17 ( .A0(kdf_keybuilder_valid), .A1(n17), .Z(kdf_keybuilder_data[49]));
Q_AN02 U18 ( .A0(kdf_keybuilder_valid), .A1(n18), .Z(kdf_keybuilder_data[48]));
Q_AN02 U19 ( .A0(kdf_keybuilder_valid), .A1(n19), .Z(kdf_keybuilder_data[47]));
Q_AN02 U20 ( .A0(kdf_keybuilder_valid), .A1(n20), .Z(kdf_keybuilder_data[46]));
Q_AN02 U21 ( .A0(kdf_keybuilder_valid), .A1(n21), .Z(kdf_keybuilder_data[45]));
Q_AN02 U22 ( .A0(kdf_keybuilder_valid), .A1(n22), .Z(kdf_keybuilder_data[44]));
Q_AN02 U23 ( .A0(kdf_keybuilder_valid), .A1(n23), .Z(kdf_keybuilder_data[43]));
Q_AN02 U24 ( .A0(kdf_keybuilder_valid), .A1(n24), .Z(kdf_keybuilder_data[42]));
Q_AN02 U25 ( .A0(kdf_keybuilder_valid), .A1(n25), .Z(kdf_keybuilder_data[41]));
Q_AN02 U26 ( .A0(kdf_keybuilder_valid), .A1(n26), .Z(kdf_keybuilder_data[40]));
Q_AN02 U27 ( .A0(kdf_keybuilder_valid), .A1(n27), .Z(kdf_keybuilder_data[39]));
Q_AN02 U28 ( .A0(kdf_keybuilder_valid), .A1(n28), .Z(kdf_keybuilder_data[38]));
Q_AN02 U29 ( .A0(kdf_keybuilder_valid), .A1(n29), .Z(kdf_keybuilder_data[37]));
Q_AN02 U30 ( .A0(kdf_keybuilder_valid), .A1(n30), .Z(kdf_keybuilder_data[36]));
Q_AN02 U31 ( .A0(kdf_keybuilder_valid), .A1(n31), .Z(kdf_keybuilder_data[35]));
Q_AN02 U32 ( .A0(kdf_keybuilder_valid), .A1(n32), .Z(kdf_keybuilder_data[34]));
Q_AN02 U33 ( .A0(kdf_keybuilder_valid), .A1(n33), .Z(kdf_keybuilder_data[33]));
Q_AN02 U34 ( .A0(kdf_keybuilder_valid), .A1(n34), .Z(kdf_keybuilder_data[32]));
Q_AN02 U35 ( .A0(kdf_keybuilder_valid), .A1(n35), .Z(kdf_keybuilder_data[31]));
Q_AN02 U36 ( .A0(kdf_keybuilder_valid), .A1(n36), .Z(kdf_keybuilder_data[30]));
Q_AN02 U37 ( .A0(kdf_keybuilder_valid), .A1(n37), .Z(kdf_keybuilder_data[29]));
Q_AN02 U38 ( .A0(kdf_keybuilder_valid), .A1(n38), .Z(kdf_keybuilder_data[28]));
Q_AN02 U39 ( .A0(kdf_keybuilder_valid), .A1(n39), .Z(kdf_keybuilder_data[27]));
Q_AN02 U40 ( .A0(kdf_keybuilder_valid), .A1(n40), .Z(kdf_keybuilder_data[26]));
Q_AN02 U41 ( .A0(kdf_keybuilder_valid), .A1(n41), .Z(kdf_keybuilder_data[25]));
Q_AN02 U42 ( .A0(kdf_keybuilder_valid), .A1(n42), .Z(kdf_keybuilder_data[24]));
Q_AN02 U43 ( .A0(kdf_keybuilder_valid), .A1(n43), .Z(kdf_keybuilder_data[23]));
Q_AN02 U44 ( .A0(kdf_keybuilder_valid), .A1(n44), .Z(kdf_keybuilder_data[22]));
Q_AN02 U45 ( .A0(kdf_keybuilder_valid), .A1(n45), .Z(kdf_keybuilder_data[21]));
Q_AN02 U46 ( .A0(kdf_keybuilder_valid), .A1(n46), .Z(kdf_keybuilder_data[20]));
Q_AN02 U47 ( .A0(kdf_keybuilder_valid), .A1(n47), .Z(kdf_keybuilder_data[19]));
Q_AN02 U48 ( .A0(kdf_keybuilder_valid), .A1(n48), .Z(kdf_keybuilder_data[18]));
Q_AN02 U49 ( .A0(kdf_keybuilder_valid), .A1(n49), .Z(kdf_keybuilder_data[17]));
Q_AN02 U50 ( .A0(kdf_keybuilder_valid), .A1(n50), .Z(kdf_keybuilder_data[16]));
Q_AN02 U51 ( .A0(kdf_keybuilder_valid), .A1(n51), .Z(kdf_keybuilder_data[15]));
Q_AN02 U52 ( .A0(kdf_keybuilder_valid), .A1(n52), .Z(kdf_keybuilder_data[14]));
Q_AN02 U53 ( .A0(kdf_keybuilder_valid), .A1(n53), .Z(kdf_keybuilder_data[13]));
Q_AN02 U54 ( .A0(kdf_keybuilder_valid), .A1(n54), .Z(kdf_keybuilder_data[12]));
Q_AN02 U55 ( .A0(kdf_keybuilder_valid), .A1(n55), .Z(kdf_keybuilder_data[11]));
Q_AN02 U56 ( .A0(kdf_keybuilder_valid), .A1(n56), .Z(kdf_keybuilder_data[10]));
Q_AN02 U57 ( .A0(kdf_keybuilder_valid), .A1(n57), .Z(kdf_keybuilder_data[9]));
Q_AN02 U58 ( .A0(kdf_keybuilder_valid), .A1(n58), .Z(kdf_keybuilder_data[8]));
Q_AN02 U59 ( .A0(kdf_keybuilder_valid), .A1(n59), .Z(kdf_keybuilder_data[7]));
Q_AN02 U60 ( .A0(kdf_keybuilder_valid), .A1(n60), .Z(kdf_keybuilder_data[6]));
Q_AN02 U61 ( .A0(kdf_keybuilder_valid), .A1(n61), .Z(kdf_keybuilder_data[5]));
Q_AN02 U62 ( .A0(kdf_keybuilder_valid), .A1(n62), .Z(kdf_keybuilder_data[4]));
Q_AN02 U63 ( .A0(kdf_keybuilder_valid), .A1(n63), .Z(kdf_keybuilder_data[3]));
Q_AN02 U64 ( .A0(kdf_keybuilder_valid), .A1(n64), .Z(kdf_keybuilder_data[2]));
Q_AN02 U65 ( .A0(kdf_keybuilder_valid), .A1(n65), .Z(kdf_keybuilder_data[1]));
Q_AN02 U66 ( .A0(kdf_keybuilder_valid), .A1(n66), .Z(kdf_keybuilder_data[0]));
Q_AN02 U67 ( .A0(kdf_keybuilder_valid), .A1(out_counter), .Z(fifo_out_ack));
Q_MX02 U68 ( .S(out_counter), .A0(fifo_out[127]), .A1(fifo_out[63]), .Z(n3));
Q_MX02 U69 ( .S(out_counter), .A0(fifo_out[126]), .A1(fifo_out[62]), .Z(n4));
Q_MX02 U70 ( .S(out_counter), .A0(fifo_out[125]), .A1(fifo_out[61]), .Z(n5));
Q_MX02 U71 ( .S(out_counter), .A0(fifo_out[124]), .A1(fifo_out[60]), .Z(n6));
Q_MX02 U72 ( .S(out_counter), .A0(fifo_out[123]), .A1(fifo_out[59]), .Z(n7));
Q_MX02 U73 ( .S(out_counter), .A0(fifo_out[122]), .A1(fifo_out[58]), .Z(n8));
Q_MX02 U74 ( .S(out_counter), .A0(fifo_out[121]), .A1(fifo_out[57]), .Z(n9));
Q_MX02 U75 ( .S(out_counter), .A0(fifo_out[120]), .A1(fifo_out[56]), .Z(n10));
Q_MX02 U76 ( .S(out_counter), .A0(fifo_out[119]), .A1(fifo_out[55]), .Z(n11));
Q_MX02 U77 ( .S(out_counter), .A0(fifo_out[118]), .A1(fifo_out[54]), .Z(n12));
Q_MX02 U78 ( .S(out_counter), .A0(fifo_out[117]), .A1(fifo_out[53]), .Z(n13));
Q_MX02 U79 ( .S(out_counter), .A0(fifo_out[116]), .A1(fifo_out[52]), .Z(n14));
Q_MX02 U80 ( .S(out_counter), .A0(fifo_out[115]), .A1(fifo_out[51]), .Z(n15));
Q_MX02 U81 ( .S(out_counter), .A0(fifo_out[114]), .A1(fifo_out[50]), .Z(n16));
Q_MX02 U82 ( .S(out_counter), .A0(fifo_out[113]), .A1(fifo_out[49]), .Z(n17));
Q_MX02 U83 ( .S(out_counter), .A0(fifo_out[112]), .A1(fifo_out[48]), .Z(n18));
Q_MX02 U84 ( .S(out_counter), .A0(fifo_out[111]), .A1(fifo_out[47]), .Z(n19));
Q_MX02 U85 ( .S(out_counter), .A0(fifo_out[110]), .A1(fifo_out[46]), .Z(n20));
Q_MX02 U86 ( .S(out_counter), .A0(fifo_out[109]), .A1(fifo_out[45]), .Z(n21));
Q_MX02 U87 ( .S(out_counter), .A0(fifo_out[108]), .A1(fifo_out[44]), .Z(n22));
Q_MX02 U88 ( .S(out_counter), .A0(fifo_out[107]), .A1(fifo_out[43]), .Z(n23));
Q_MX02 U89 ( .S(out_counter), .A0(fifo_out[106]), .A1(fifo_out[42]), .Z(n24));
Q_MX02 U90 ( .S(out_counter), .A0(fifo_out[105]), .A1(fifo_out[41]), .Z(n25));
Q_MX02 U91 ( .S(out_counter), .A0(fifo_out[104]), .A1(fifo_out[40]), .Z(n26));
Q_MX02 U92 ( .S(out_counter), .A0(fifo_out[103]), .A1(fifo_out[39]), .Z(n27));
Q_MX02 U93 ( .S(out_counter), .A0(fifo_out[102]), .A1(fifo_out[38]), .Z(n28));
Q_MX02 U94 ( .S(out_counter), .A0(fifo_out[101]), .A1(fifo_out[37]), .Z(n29));
Q_MX02 U95 ( .S(out_counter), .A0(fifo_out[100]), .A1(fifo_out[36]), .Z(n30));
Q_MX02 U96 ( .S(out_counter), .A0(fifo_out[99]), .A1(fifo_out[35]), .Z(n31));
Q_MX02 U97 ( .S(out_counter), .A0(fifo_out[98]), .A1(fifo_out[34]), .Z(n32));
Q_MX02 U98 ( .S(out_counter), .A0(fifo_out[97]), .A1(fifo_out[33]), .Z(n33));
Q_MX02 U99 ( .S(out_counter), .A0(fifo_out[96]), .A1(fifo_out[32]), .Z(n34));
Q_MX02 U100 ( .S(out_counter), .A0(fifo_out[95]), .A1(fifo_out[31]), .Z(n35));
Q_MX02 U101 ( .S(out_counter), .A0(fifo_out[94]), .A1(fifo_out[30]), .Z(n36));
Q_MX02 U102 ( .S(out_counter), .A0(fifo_out[93]), .A1(fifo_out[29]), .Z(n37));
Q_MX02 U103 ( .S(out_counter), .A0(fifo_out[92]), .A1(fifo_out[28]), .Z(n38));
Q_MX02 U104 ( .S(out_counter), .A0(fifo_out[91]), .A1(fifo_out[27]), .Z(n39));
Q_MX02 U105 ( .S(out_counter), .A0(fifo_out[90]), .A1(fifo_out[26]), .Z(n40));
Q_MX02 U106 ( .S(out_counter), .A0(fifo_out[89]), .A1(fifo_out[25]), .Z(n41));
Q_MX02 U107 ( .S(out_counter), .A0(fifo_out[88]), .A1(fifo_out[24]), .Z(n42));
Q_MX02 U108 ( .S(out_counter), .A0(fifo_out[87]), .A1(fifo_out[23]), .Z(n43));
Q_MX02 U109 ( .S(out_counter), .A0(fifo_out[86]), .A1(fifo_out[22]), .Z(n44));
Q_MX02 U110 ( .S(out_counter), .A0(fifo_out[85]), .A1(fifo_out[21]), .Z(n45));
Q_MX02 U111 ( .S(out_counter), .A0(fifo_out[84]), .A1(fifo_out[20]), .Z(n46));
Q_MX02 U112 ( .S(out_counter), .A0(fifo_out[83]), .A1(fifo_out[19]), .Z(n47));
Q_MX02 U113 ( .S(out_counter), .A0(fifo_out[82]), .A1(fifo_out[18]), .Z(n48));
Q_MX02 U114 ( .S(out_counter), .A0(fifo_out[81]), .A1(fifo_out[17]), .Z(n49));
Q_MX02 U115 ( .S(out_counter), .A0(fifo_out[80]), .A1(fifo_out[16]), .Z(n50));
Q_MX02 U116 ( .S(out_counter), .A0(fifo_out[79]), .A1(fifo_out[15]), .Z(n51));
Q_MX02 U117 ( .S(out_counter), .A0(fifo_out[78]), .A1(fifo_out[14]), .Z(n52));
Q_MX02 U118 ( .S(out_counter), .A0(fifo_out[77]), .A1(fifo_out[13]), .Z(n53));
Q_MX02 U119 ( .S(out_counter), .A0(fifo_out[76]), .A1(fifo_out[12]), .Z(n54));
Q_MX02 U120 ( .S(out_counter), .A0(fifo_out[75]), .A1(fifo_out[11]), .Z(n55));
Q_MX02 U121 ( .S(out_counter), .A0(fifo_out[74]), .A1(fifo_out[10]), .Z(n56));
Q_MX02 U122 ( .S(out_counter), .A0(fifo_out[73]), .A1(fifo_out[9]), .Z(n57));
Q_MX02 U123 ( .S(out_counter), .A0(fifo_out[72]), .A1(fifo_out[8]), .Z(n58));
Q_MX02 U124 ( .S(out_counter), .A0(fifo_out[71]), .A1(fifo_out[7]), .Z(n59));
Q_MX02 U125 ( .S(out_counter), .A0(fifo_out[70]), .A1(fifo_out[6]), .Z(n60));
Q_MX02 U126 ( .S(out_counter), .A0(fifo_out[69]), .A1(fifo_out[5]), .Z(n61));
Q_MX02 U127 ( .S(out_counter), .A0(fifo_out[68]), .A1(fifo_out[4]), .Z(n62));
Q_MX02 U128 ( .S(out_counter), .A0(fifo_out[67]), .A1(fifo_out[3]), .Z(n63));
Q_MX02 U129 ( .S(out_counter), .A0(fifo_out[66]), .A1(fifo_out[2]), .Z(n64));
Q_MX02 U130 ( .S(out_counter), .A0(fifo_out[65]), .A1(fifo_out[1]), .Z(n65));
Q_MX02 U131 ( .S(out_counter), .A0(fifo_out[64]), .A1(fifo_out[0]), .Z(n66));
Q_AN02 U132 ( .A0(n2), .A1(kdf_keybuilder_valid), .Z(n67));
Q_OR02 U133 ( .A0(in_counter[1]), .A1(cmdfifo_kdf_cmd[3]), .Z(n88));
Q_AN02 U134 ( .A0(n88), .A1(cmdfifo_kdf_cmd[2]), .Z(n82));
Q_AO21 U135 ( .A0(n88), .A1(cmdfifo_kdf_cmd[1]), .B0(n82), .Z(n73));
Q_OA21 U136 ( .A0(cmdfifo_kdf_cmd[0]), .A1(cmdfifo_kdf_cmd[2]), .B0(n89), .Z(n74));
Q_AO21 U137 ( .A0(n73), .A1(n87), .B0(n74), .Z(n72));
Q_AN02 U138 ( .A0(in_counter[2]), .A1(n76), .Z(n89));
Q_AN02 U139 ( .A0(cmdfifo_kdf_valid), .A1(n72), .Z(n69));
Q_NR02 U140 ( .A0(in_counter[2]), .A1(cmdfifo_kdf_cmd[1]), .Z(n83));
Q_AO21 U141 ( .A0(n88), .A1(n83), .B0(n84), .Z(n80));
Q_INV U142 ( .A(cmdfifo_kdf_cmd[0]), .Z(n75));
Q_AN02 U143 ( .A0(n89), .A1(n75), .Z(n84));
Q_NR02 U144 ( .A0(in_counter[2]), .A1(in_counter[1]), .Z(n78));
Q_INV U145 ( .A(cmdfifo_kdf_cmd[3]), .Z(n77));
Q_AN02 U146 ( .A0(n78), .A1(n77), .Z(n81));
Q_INV U147 ( .A(cmdfifo_kdf_cmd[2]), .Z(n79));
Q_AO21 U148 ( .A0(n80), .A1(n79), .B0(n81), .Z(n92));
Q_INV U149 ( .A(fifo_in_stall), .Z(n93));
Q_AN03 U150 ( .A0(cmdfifo_kdf_valid), .A1(n93), .A2(n92), .Z(n68));
Q_OA21 U151 ( .A0(n93), .A1(n82), .B0(n83), .Z(n86));
Q_OA21 U152 ( .A0(n93), .A1(cmdfifo_kdf_cmd[2]), .B0(n84), .Z(n85));
Q_OA21 U153 ( .A0(n86), .A1(n85), .B0(cmdfifo_kdf_valid), .Z(n70));
Q_AN03 U154 ( .A0(n87), .A1(cmdfifo_kdf_cmd[1]), .A2(n88), .Z(n90));
Q_AO21 U155 ( .A0(n89), .A1(cmdfifo_kdf_cmd[0]), .B0(n90), .Z(n91));
Q_AN02 U156 ( .A0(cmdfifo_kdf_valid), .A1(n91), .Z(n71));
Q_AN03 U157 ( .A0(n93), .A1(n92), .A2(keyfifo_merger_valid), .Z(n226));
Q_OR02 U158 ( .A0(n94), .A1(fifo_in_stall), .Z(sha_tag_stall));
Q_INV U159 ( .A(n69), .Z(n94));
Q_MX02 U160 ( .S(n68), .A0(n95), .A1(keyfifo_merger_valid), .Z(merger_keyfifo_ack));
Q_AN02 U161 ( .A0(n69), .A1(sha_tag_valid), .Z(n95));
Q_MX02 U162 ( .S(n70), .A0(n96), .A1(keyfifo_merger_data[127]), .Z(fifo_in[127]));
Q_AN02 U163 ( .A0(n71), .A1(sha_tag_data[127]), .Z(n96));
Q_MX02 U164 ( .S(n70), .A0(n97), .A1(keyfifo_merger_data[126]), .Z(fifo_in[126]));
Q_AN02 U165 ( .A0(n71), .A1(sha_tag_data[126]), .Z(n97));
Q_MX02 U166 ( .S(n70), .A0(n98), .A1(keyfifo_merger_data[125]), .Z(fifo_in[125]));
Q_AN02 U167 ( .A0(n71), .A1(sha_tag_data[125]), .Z(n98));
Q_MX02 U168 ( .S(n70), .A0(n99), .A1(keyfifo_merger_data[124]), .Z(fifo_in[124]));
Q_AN02 U169 ( .A0(n71), .A1(sha_tag_data[124]), .Z(n99));
Q_MX02 U170 ( .S(n70), .A0(n100), .A1(keyfifo_merger_data[123]), .Z(fifo_in[123]));
Q_AN02 U171 ( .A0(n71), .A1(sha_tag_data[123]), .Z(n100));
Q_MX02 U172 ( .S(n70), .A0(n101), .A1(keyfifo_merger_data[122]), .Z(fifo_in[122]));
Q_AN02 U173 ( .A0(n71), .A1(sha_tag_data[122]), .Z(n101));
Q_MX02 U174 ( .S(n70), .A0(n102), .A1(keyfifo_merger_data[121]), .Z(fifo_in[121]));
Q_AN02 U175 ( .A0(n71), .A1(sha_tag_data[121]), .Z(n102));
Q_MX02 U176 ( .S(n70), .A0(n103), .A1(keyfifo_merger_data[120]), .Z(fifo_in[120]));
Q_AN02 U177 ( .A0(n71), .A1(sha_tag_data[120]), .Z(n103));
Q_MX02 U178 ( .S(n70), .A0(n104), .A1(keyfifo_merger_data[119]), .Z(fifo_in[119]));
Q_AN02 U179 ( .A0(n71), .A1(sha_tag_data[119]), .Z(n104));
Q_MX02 U180 ( .S(n70), .A0(n105), .A1(keyfifo_merger_data[118]), .Z(fifo_in[118]));
Q_AN02 U181 ( .A0(n71), .A1(sha_tag_data[118]), .Z(n105));
Q_MX02 U182 ( .S(n70), .A0(n106), .A1(keyfifo_merger_data[117]), .Z(fifo_in[117]));
Q_AN02 U183 ( .A0(n71), .A1(sha_tag_data[117]), .Z(n106));
Q_MX02 U184 ( .S(n70), .A0(n107), .A1(keyfifo_merger_data[116]), .Z(fifo_in[116]));
Q_AN02 U185 ( .A0(n71), .A1(sha_tag_data[116]), .Z(n107));
Q_MX02 U186 ( .S(n70), .A0(n108), .A1(keyfifo_merger_data[115]), .Z(fifo_in[115]));
Q_AN02 U187 ( .A0(n71), .A1(sha_tag_data[115]), .Z(n108));
Q_MX02 U188 ( .S(n70), .A0(n109), .A1(keyfifo_merger_data[114]), .Z(fifo_in[114]));
Q_AN02 U189 ( .A0(n71), .A1(sha_tag_data[114]), .Z(n109));
Q_MX02 U190 ( .S(n70), .A0(n110), .A1(keyfifo_merger_data[113]), .Z(fifo_in[113]));
Q_AN02 U191 ( .A0(n71), .A1(sha_tag_data[113]), .Z(n110));
Q_MX02 U192 ( .S(n70), .A0(n111), .A1(keyfifo_merger_data[112]), .Z(fifo_in[112]));
Q_AN02 U193 ( .A0(n71), .A1(sha_tag_data[112]), .Z(n111));
Q_MX02 U194 ( .S(n70), .A0(n112), .A1(keyfifo_merger_data[111]), .Z(fifo_in[111]));
Q_AN02 U195 ( .A0(n71), .A1(sha_tag_data[111]), .Z(n112));
Q_MX02 U196 ( .S(n70), .A0(n113), .A1(keyfifo_merger_data[110]), .Z(fifo_in[110]));
Q_AN02 U197 ( .A0(n71), .A1(sha_tag_data[110]), .Z(n113));
Q_MX02 U198 ( .S(n70), .A0(n114), .A1(keyfifo_merger_data[109]), .Z(fifo_in[109]));
Q_AN02 U199 ( .A0(n71), .A1(sha_tag_data[109]), .Z(n114));
Q_MX02 U200 ( .S(n70), .A0(n115), .A1(keyfifo_merger_data[108]), .Z(fifo_in[108]));
Q_AN02 U201 ( .A0(n71), .A1(sha_tag_data[108]), .Z(n115));
Q_MX02 U202 ( .S(n70), .A0(n116), .A1(keyfifo_merger_data[107]), .Z(fifo_in[107]));
Q_AN02 U203 ( .A0(n71), .A1(sha_tag_data[107]), .Z(n116));
Q_MX02 U204 ( .S(n70), .A0(n117), .A1(keyfifo_merger_data[106]), .Z(fifo_in[106]));
Q_AN02 U205 ( .A0(n71), .A1(sha_tag_data[106]), .Z(n117));
Q_MX02 U206 ( .S(n70), .A0(n118), .A1(keyfifo_merger_data[105]), .Z(fifo_in[105]));
Q_AN02 U207 ( .A0(n71), .A1(sha_tag_data[105]), .Z(n118));
Q_MX02 U208 ( .S(n70), .A0(n119), .A1(keyfifo_merger_data[104]), .Z(fifo_in[104]));
Q_AN02 U209 ( .A0(n71), .A1(sha_tag_data[104]), .Z(n119));
Q_MX02 U210 ( .S(n70), .A0(n120), .A1(keyfifo_merger_data[103]), .Z(fifo_in[103]));
Q_AN02 U211 ( .A0(n71), .A1(sha_tag_data[103]), .Z(n120));
Q_MX02 U212 ( .S(n70), .A0(n121), .A1(keyfifo_merger_data[102]), .Z(fifo_in[102]));
Q_AN02 U213 ( .A0(n71), .A1(sha_tag_data[102]), .Z(n121));
Q_MX02 U214 ( .S(n70), .A0(n122), .A1(keyfifo_merger_data[101]), .Z(fifo_in[101]));
Q_AN02 U215 ( .A0(n71), .A1(sha_tag_data[101]), .Z(n122));
Q_MX02 U216 ( .S(n70), .A0(n123), .A1(keyfifo_merger_data[100]), .Z(fifo_in[100]));
Q_AN02 U217 ( .A0(n71), .A1(sha_tag_data[100]), .Z(n123));
Q_MX02 U218 ( .S(n70), .A0(n124), .A1(keyfifo_merger_data[99]), .Z(fifo_in[99]));
Q_AN02 U219 ( .A0(n71), .A1(sha_tag_data[99]), .Z(n124));
Q_MX02 U220 ( .S(n70), .A0(n125), .A1(keyfifo_merger_data[98]), .Z(fifo_in[98]));
Q_AN02 U221 ( .A0(n71), .A1(sha_tag_data[98]), .Z(n125));
Q_MX02 U222 ( .S(n70), .A0(n126), .A1(keyfifo_merger_data[97]), .Z(fifo_in[97]));
Q_AN02 U223 ( .A0(n71), .A1(sha_tag_data[97]), .Z(n126));
Q_MX02 U224 ( .S(n70), .A0(n127), .A1(keyfifo_merger_data[96]), .Z(fifo_in[96]));
Q_AN02 U225 ( .A0(n71), .A1(sha_tag_data[96]), .Z(n127));
Q_MX02 U226 ( .S(n70), .A0(n128), .A1(keyfifo_merger_data[95]), .Z(fifo_in[95]));
Q_AN02 U227 ( .A0(n71), .A1(sha_tag_data[95]), .Z(n128));
Q_MX02 U228 ( .S(n70), .A0(n129), .A1(keyfifo_merger_data[94]), .Z(fifo_in[94]));
Q_AN02 U229 ( .A0(n71), .A1(sha_tag_data[94]), .Z(n129));
Q_MX02 U230 ( .S(n70), .A0(n130), .A1(keyfifo_merger_data[93]), .Z(fifo_in[93]));
Q_AN02 U231 ( .A0(n71), .A1(sha_tag_data[93]), .Z(n130));
Q_MX02 U232 ( .S(n70), .A0(n131), .A1(keyfifo_merger_data[92]), .Z(fifo_in[92]));
Q_AN02 U233 ( .A0(n71), .A1(sha_tag_data[92]), .Z(n131));
Q_MX02 U234 ( .S(n70), .A0(n132), .A1(keyfifo_merger_data[91]), .Z(fifo_in[91]));
Q_AN02 U235 ( .A0(n71), .A1(sha_tag_data[91]), .Z(n132));
Q_MX02 U236 ( .S(n70), .A0(n133), .A1(keyfifo_merger_data[90]), .Z(fifo_in[90]));
Q_AN02 U237 ( .A0(n71), .A1(sha_tag_data[90]), .Z(n133));
Q_MX02 U238 ( .S(n70), .A0(n134), .A1(keyfifo_merger_data[89]), .Z(fifo_in[89]));
Q_AN02 U239 ( .A0(n71), .A1(sha_tag_data[89]), .Z(n134));
Q_MX02 U240 ( .S(n70), .A0(n135), .A1(keyfifo_merger_data[88]), .Z(fifo_in[88]));
Q_AN02 U241 ( .A0(n71), .A1(sha_tag_data[88]), .Z(n135));
Q_MX02 U242 ( .S(n70), .A0(n136), .A1(keyfifo_merger_data[87]), .Z(fifo_in[87]));
Q_AN02 U243 ( .A0(n71), .A1(sha_tag_data[87]), .Z(n136));
Q_MX02 U244 ( .S(n70), .A0(n137), .A1(keyfifo_merger_data[86]), .Z(fifo_in[86]));
Q_AN02 U245 ( .A0(n71), .A1(sha_tag_data[86]), .Z(n137));
Q_MX02 U246 ( .S(n70), .A0(n138), .A1(keyfifo_merger_data[85]), .Z(fifo_in[85]));
Q_AN02 U247 ( .A0(n71), .A1(sha_tag_data[85]), .Z(n138));
Q_MX02 U248 ( .S(n70), .A0(n139), .A1(keyfifo_merger_data[84]), .Z(fifo_in[84]));
Q_AN02 U249 ( .A0(n71), .A1(sha_tag_data[84]), .Z(n139));
Q_MX02 U250 ( .S(n70), .A0(n140), .A1(keyfifo_merger_data[83]), .Z(fifo_in[83]));
Q_AN02 U251 ( .A0(n71), .A1(sha_tag_data[83]), .Z(n140));
Q_MX02 U252 ( .S(n70), .A0(n141), .A1(keyfifo_merger_data[82]), .Z(fifo_in[82]));
Q_AN02 U253 ( .A0(n71), .A1(sha_tag_data[82]), .Z(n141));
Q_MX02 U254 ( .S(n70), .A0(n142), .A1(keyfifo_merger_data[81]), .Z(fifo_in[81]));
Q_AN02 U255 ( .A0(n71), .A1(sha_tag_data[81]), .Z(n142));
Q_MX02 U256 ( .S(n70), .A0(n143), .A1(keyfifo_merger_data[80]), .Z(fifo_in[80]));
Q_AN02 U257 ( .A0(n71), .A1(sha_tag_data[80]), .Z(n143));
Q_MX02 U258 ( .S(n70), .A0(n144), .A1(keyfifo_merger_data[79]), .Z(fifo_in[79]));
Q_AN02 U259 ( .A0(n71), .A1(sha_tag_data[79]), .Z(n144));
Q_MX02 U260 ( .S(n70), .A0(n145), .A1(keyfifo_merger_data[78]), .Z(fifo_in[78]));
Q_AN02 U261 ( .A0(n71), .A1(sha_tag_data[78]), .Z(n145));
Q_MX02 U262 ( .S(n70), .A0(n146), .A1(keyfifo_merger_data[77]), .Z(fifo_in[77]));
Q_AN02 U263 ( .A0(n71), .A1(sha_tag_data[77]), .Z(n146));
Q_MX02 U264 ( .S(n70), .A0(n147), .A1(keyfifo_merger_data[76]), .Z(fifo_in[76]));
Q_AN02 U265 ( .A0(n71), .A1(sha_tag_data[76]), .Z(n147));
Q_MX02 U266 ( .S(n70), .A0(n148), .A1(keyfifo_merger_data[75]), .Z(fifo_in[75]));
Q_AN02 U267 ( .A0(n71), .A1(sha_tag_data[75]), .Z(n148));
Q_MX02 U268 ( .S(n70), .A0(n149), .A1(keyfifo_merger_data[74]), .Z(fifo_in[74]));
Q_AN02 U269 ( .A0(n71), .A1(sha_tag_data[74]), .Z(n149));
Q_MX02 U270 ( .S(n70), .A0(n150), .A1(keyfifo_merger_data[73]), .Z(fifo_in[73]));
Q_AN02 U271 ( .A0(n71), .A1(sha_tag_data[73]), .Z(n150));
Q_MX02 U272 ( .S(n70), .A0(n151), .A1(keyfifo_merger_data[72]), .Z(fifo_in[72]));
Q_AN02 U273 ( .A0(n71), .A1(sha_tag_data[72]), .Z(n151));
Q_MX02 U274 ( .S(n70), .A0(n152), .A1(keyfifo_merger_data[71]), .Z(fifo_in[71]));
Q_AN02 U275 ( .A0(n71), .A1(sha_tag_data[71]), .Z(n152));
Q_MX02 U276 ( .S(n70), .A0(n153), .A1(keyfifo_merger_data[70]), .Z(fifo_in[70]));
Q_AN02 U277 ( .A0(n71), .A1(sha_tag_data[70]), .Z(n153));
Q_MX02 U278 ( .S(n70), .A0(n154), .A1(keyfifo_merger_data[69]), .Z(fifo_in[69]));
Q_AN02 U279 ( .A0(n71), .A1(sha_tag_data[69]), .Z(n154));
Q_MX02 U280 ( .S(n70), .A0(n155), .A1(keyfifo_merger_data[68]), .Z(fifo_in[68]));
Q_AN02 U281 ( .A0(n71), .A1(sha_tag_data[68]), .Z(n155));
Q_MX02 U282 ( .S(n70), .A0(n156), .A1(keyfifo_merger_data[67]), .Z(fifo_in[67]));
Q_AN02 U283 ( .A0(n71), .A1(sha_tag_data[67]), .Z(n156));
Q_MX02 U284 ( .S(n70), .A0(n157), .A1(keyfifo_merger_data[66]), .Z(fifo_in[66]));
Q_AN02 U285 ( .A0(n71), .A1(sha_tag_data[66]), .Z(n157));
Q_MX02 U286 ( .S(n70), .A0(n158), .A1(keyfifo_merger_data[65]), .Z(fifo_in[65]));
Q_AN02 U287 ( .A0(n71), .A1(sha_tag_data[65]), .Z(n158));
Q_MX02 U288 ( .S(n70), .A0(n159), .A1(keyfifo_merger_data[64]), .Z(fifo_in[64]));
Q_AN02 U289 ( .A0(n71), .A1(sha_tag_data[64]), .Z(n159));
Q_MX02 U290 ( .S(n70), .A0(n160), .A1(keyfifo_merger_data[63]), .Z(fifo_in[63]));
Q_AN02 U291 ( .A0(n71), .A1(sha_tag_data[63]), .Z(n160));
Q_MX02 U292 ( .S(n70), .A0(n161), .A1(keyfifo_merger_data[62]), .Z(fifo_in[62]));
Q_AN02 U293 ( .A0(n71), .A1(sha_tag_data[62]), .Z(n161));
Q_MX02 U294 ( .S(n70), .A0(n162), .A1(keyfifo_merger_data[61]), .Z(fifo_in[61]));
Q_AN02 U295 ( .A0(n71), .A1(sha_tag_data[61]), .Z(n162));
Q_MX02 U296 ( .S(n70), .A0(n163), .A1(keyfifo_merger_data[60]), .Z(fifo_in[60]));
Q_AN02 U297 ( .A0(n71), .A1(sha_tag_data[60]), .Z(n163));
Q_MX02 U298 ( .S(n70), .A0(n164), .A1(keyfifo_merger_data[59]), .Z(fifo_in[59]));
Q_AN02 U299 ( .A0(n71), .A1(sha_tag_data[59]), .Z(n164));
Q_MX02 U300 ( .S(n70), .A0(n165), .A1(keyfifo_merger_data[58]), .Z(fifo_in[58]));
Q_AN02 U301 ( .A0(n71), .A1(sha_tag_data[58]), .Z(n165));
Q_MX02 U302 ( .S(n70), .A0(n166), .A1(keyfifo_merger_data[57]), .Z(fifo_in[57]));
Q_AN02 U303 ( .A0(n71), .A1(sha_tag_data[57]), .Z(n166));
Q_MX02 U304 ( .S(n70), .A0(n167), .A1(keyfifo_merger_data[56]), .Z(fifo_in[56]));
Q_AN02 U305 ( .A0(n71), .A1(sha_tag_data[56]), .Z(n167));
Q_MX02 U306 ( .S(n70), .A0(n168), .A1(keyfifo_merger_data[55]), .Z(fifo_in[55]));
Q_AN02 U307 ( .A0(n71), .A1(sha_tag_data[55]), .Z(n168));
Q_MX02 U308 ( .S(n70), .A0(n169), .A1(keyfifo_merger_data[54]), .Z(fifo_in[54]));
Q_AN02 U309 ( .A0(n71), .A1(sha_tag_data[54]), .Z(n169));
Q_MX02 U310 ( .S(n70), .A0(n170), .A1(keyfifo_merger_data[53]), .Z(fifo_in[53]));
Q_AN02 U311 ( .A0(n71), .A1(sha_tag_data[53]), .Z(n170));
Q_MX02 U312 ( .S(n70), .A0(n171), .A1(keyfifo_merger_data[52]), .Z(fifo_in[52]));
Q_AN02 U313 ( .A0(n71), .A1(sha_tag_data[52]), .Z(n171));
Q_MX02 U314 ( .S(n70), .A0(n172), .A1(keyfifo_merger_data[51]), .Z(fifo_in[51]));
Q_AN02 U315 ( .A0(n71), .A1(sha_tag_data[51]), .Z(n172));
Q_MX02 U316 ( .S(n70), .A0(n173), .A1(keyfifo_merger_data[50]), .Z(fifo_in[50]));
Q_AN02 U317 ( .A0(n71), .A1(sha_tag_data[50]), .Z(n173));
Q_MX02 U318 ( .S(n70), .A0(n174), .A1(keyfifo_merger_data[49]), .Z(fifo_in[49]));
Q_AN02 U319 ( .A0(n71), .A1(sha_tag_data[49]), .Z(n174));
Q_MX02 U320 ( .S(n70), .A0(n175), .A1(keyfifo_merger_data[48]), .Z(fifo_in[48]));
Q_AN02 U321 ( .A0(n71), .A1(sha_tag_data[48]), .Z(n175));
Q_MX02 U322 ( .S(n70), .A0(n176), .A1(keyfifo_merger_data[47]), .Z(fifo_in[47]));
Q_AN02 U323 ( .A0(n71), .A1(sha_tag_data[47]), .Z(n176));
Q_MX02 U324 ( .S(n70), .A0(n177), .A1(keyfifo_merger_data[46]), .Z(fifo_in[46]));
Q_AN02 U325 ( .A0(n71), .A1(sha_tag_data[46]), .Z(n177));
Q_MX02 U326 ( .S(n70), .A0(n178), .A1(keyfifo_merger_data[45]), .Z(fifo_in[45]));
Q_AN02 U327 ( .A0(n71), .A1(sha_tag_data[45]), .Z(n178));
Q_MX02 U328 ( .S(n70), .A0(n179), .A1(keyfifo_merger_data[44]), .Z(fifo_in[44]));
Q_AN02 U329 ( .A0(n71), .A1(sha_tag_data[44]), .Z(n179));
Q_MX02 U330 ( .S(n70), .A0(n180), .A1(keyfifo_merger_data[43]), .Z(fifo_in[43]));
Q_AN02 U331 ( .A0(n71), .A1(sha_tag_data[43]), .Z(n180));
Q_MX02 U332 ( .S(n70), .A0(n181), .A1(keyfifo_merger_data[42]), .Z(fifo_in[42]));
Q_AN02 U333 ( .A0(n71), .A1(sha_tag_data[42]), .Z(n181));
Q_MX02 U334 ( .S(n70), .A0(n182), .A1(keyfifo_merger_data[41]), .Z(fifo_in[41]));
Q_AN02 U335 ( .A0(n71), .A1(sha_tag_data[41]), .Z(n182));
Q_MX02 U336 ( .S(n70), .A0(n183), .A1(keyfifo_merger_data[40]), .Z(fifo_in[40]));
Q_AN02 U337 ( .A0(n71), .A1(sha_tag_data[40]), .Z(n183));
Q_MX02 U338 ( .S(n70), .A0(n184), .A1(keyfifo_merger_data[39]), .Z(fifo_in[39]));
Q_AN02 U339 ( .A0(n71), .A1(sha_tag_data[39]), .Z(n184));
Q_MX02 U340 ( .S(n70), .A0(n185), .A1(keyfifo_merger_data[38]), .Z(fifo_in[38]));
Q_AN02 U341 ( .A0(n71), .A1(sha_tag_data[38]), .Z(n185));
Q_MX02 U342 ( .S(n70), .A0(n186), .A1(keyfifo_merger_data[37]), .Z(fifo_in[37]));
Q_AN02 U343 ( .A0(n71), .A1(sha_tag_data[37]), .Z(n186));
Q_MX02 U344 ( .S(n70), .A0(n187), .A1(keyfifo_merger_data[36]), .Z(fifo_in[36]));
Q_AN02 U345 ( .A0(n71), .A1(sha_tag_data[36]), .Z(n187));
Q_MX02 U346 ( .S(n70), .A0(n188), .A1(keyfifo_merger_data[35]), .Z(fifo_in[35]));
Q_AN02 U347 ( .A0(n71), .A1(sha_tag_data[35]), .Z(n188));
Q_MX02 U348 ( .S(n70), .A0(n189), .A1(keyfifo_merger_data[34]), .Z(fifo_in[34]));
Q_AN02 U349 ( .A0(n71), .A1(sha_tag_data[34]), .Z(n189));
Q_MX02 U350 ( .S(n70), .A0(n190), .A1(keyfifo_merger_data[33]), .Z(fifo_in[33]));
Q_AN02 U351 ( .A0(n71), .A1(sha_tag_data[33]), .Z(n190));
Q_MX02 U352 ( .S(n70), .A0(n191), .A1(keyfifo_merger_data[32]), .Z(fifo_in[32]));
Q_AN02 U353 ( .A0(n71), .A1(sha_tag_data[32]), .Z(n191));
Q_MX02 U354 ( .S(n70), .A0(n192), .A1(keyfifo_merger_data[31]), .Z(fifo_in[31]));
Q_AN02 U355 ( .A0(n71), .A1(sha_tag_data[31]), .Z(n192));
Q_MX02 U356 ( .S(n70), .A0(n193), .A1(keyfifo_merger_data[30]), .Z(fifo_in[30]));
Q_AN02 U357 ( .A0(n71), .A1(sha_tag_data[30]), .Z(n193));
Q_MX02 U358 ( .S(n70), .A0(n194), .A1(keyfifo_merger_data[29]), .Z(fifo_in[29]));
Q_AN02 U359 ( .A0(n71), .A1(sha_tag_data[29]), .Z(n194));
Q_MX02 U360 ( .S(n70), .A0(n195), .A1(keyfifo_merger_data[28]), .Z(fifo_in[28]));
Q_AN02 U361 ( .A0(n71), .A1(sha_tag_data[28]), .Z(n195));
Q_MX02 U362 ( .S(n70), .A0(n196), .A1(keyfifo_merger_data[27]), .Z(fifo_in[27]));
Q_AN02 U363 ( .A0(n71), .A1(sha_tag_data[27]), .Z(n196));
Q_MX02 U364 ( .S(n70), .A0(n197), .A1(keyfifo_merger_data[26]), .Z(fifo_in[26]));
Q_AN02 U365 ( .A0(n71), .A1(sha_tag_data[26]), .Z(n197));
Q_MX02 U366 ( .S(n70), .A0(n198), .A1(keyfifo_merger_data[25]), .Z(fifo_in[25]));
Q_AN02 U367 ( .A0(n71), .A1(sha_tag_data[25]), .Z(n198));
Q_MX02 U368 ( .S(n70), .A0(n199), .A1(keyfifo_merger_data[24]), .Z(fifo_in[24]));
Q_AN02 U369 ( .A0(n71), .A1(sha_tag_data[24]), .Z(n199));
Q_MX02 U370 ( .S(n70), .A0(n200), .A1(keyfifo_merger_data[23]), .Z(fifo_in[23]));
Q_AN02 U371 ( .A0(n71), .A1(sha_tag_data[23]), .Z(n200));
Q_MX02 U372 ( .S(n70), .A0(n201), .A1(keyfifo_merger_data[22]), .Z(fifo_in[22]));
Q_AN02 U373 ( .A0(n71), .A1(sha_tag_data[22]), .Z(n201));
Q_MX02 U374 ( .S(n70), .A0(n202), .A1(keyfifo_merger_data[21]), .Z(fifo_in[21]));
Q_AN02 U375 ( .A0(n71), .A1(sha_tag_data[21]), .Z(n202));
Q_MX02 U376 ( .S(n70), .A0(n203), .A1(keyfifo_merger_data[20]), .Z(fifo_in[20]));
Q_AN02 U377 ( .A0(n71), .A1(sha_tag_data[20]), .Z(n203));
Q_MX02 U378 ( .S(n70), .A0(n204), .A1(keyfifo_merger_data[19]), .Z(fifo_in[19]));
Q_AN02 U379 ( .A0(n71), .A1(sha_tag_data[19]), .Z(n204));
Q_MX02 U380 ( .S(n70), .A0(n205), .A1(keyfifo_merger_data[18]), .Z(fifo_in[18]));
Q_AN02 U381 ( .A0(n71), .A1(sha_tag_data[18]), .Z(n205));
Q_MX02 U382 ( .S(n70), .A0(n206), .A1(keyfifo_merger_data[17]), .Z(fifo_in[17]));
Q_AN02 U383 ( .A0(n71), .A1(sha_tag_data[17]), .Z(n206));
Q_MX02 U384 ( .S(n70), .A0(n207), .A1(keyfifo_merger_data[16]), .Z(fifo_in[16]));
Q_AN02 U385 ( .A0(n71), .A1(sha_tag_data[16]), .Z(n207));
Q_MX02 U386 ( .S(n70), .A0(n208), .A1(keyfifo_merger_data[15]), .Z(fifo_in[15]));
Q_AN02 U387 ( .A0(n71), .A1(sha_tag_data[15]), .Z(n208));
Q_MX02 U388 ( .S(n70), .A0(n209), .A1(keyfifo_merger_data[14]), .Z(fifo_in[14]));
Q_AN02 U389 ( .A0(n71), .A1(sha_tag_data[14]), .Z(n209));
Q_MX02 U390 ( .S(n70), .A0(n210), .A1(keyfifo_merger_data[13]), .Z(fifo_in[13]));
Q_AN02 U391 ( .A0(n71), .A1(sha_tag_data[13]), .Z(n210));
Q_MX02 U392 ( .S(n70), .A0(n211), .A1(keyfifo_merger_data[12]), .Z(fifo_in[12]));
Q_AN02 U393 ( .A0(n71), .A1(sha_tag_data[12]), .Z(n211));
Q_MX02 U394 ( .S(n70), .A0(n212), .A1(keyfifo_merger_data[11]), .Z(fifo_in[11]));
Q_AN02 U395 ( .A0(n71), .A1(sha_tag_data[11]), .Z(n212));
Q_MX02 U396 ( .S(n70), .A0(n213), .A1(keyfifo_merger_data[10]), .Z(fifo_in[10]));
Q_AN02 U397 ( .A0(n71), .A1(sha_tag_data[10]), .Z(n213));
Q_MX02 U398 ( .S(n70), .A0(n214), .A1(keyfifo_merger_data[9]), .Z(fifo_in[9]));
Q_AN02 U399 ( .A0(n71), .A1(sha_tag_data[9]), .Z(n214));
Q_MX02 U400 ( .S(n70), .A0(n215), .A1(keyfifo_merger_data[8]), .Z(fifo_in[8]));
Q_AN02 U401 ( .A0(n71), .A1(sha_tag_data[8]), .Z(n215));
Q_MX02 U402 ( .S(n70), .A0(n216), .A1(keyfifo_merger_data[7]), .Z(fifo_in[7]));
Q_AN02 U403 ( .A0(n71), .A1(sha_tag_data[7]), .Z(n216));
Q_MX02 U404 ( .S(n70), .A0(n217), .A1(keyfifo_merger_data[6]), .Z(fifo_in[6]));
Q_AN02 U405 ( .A0(n71), .A1(sha_tag_data[6]), .Z(n217));
Q_MX02 U406 ( .S(n70), .A0(n218), .A1(keyfifo_merger_data[5]), .Z(fifo_in[5]));
Q_AN02 U407 ( .A0(n71), .A1(sha_tag_data[5]), .Z(n218));
Q_MX02 U408 ( .S(n70), .A0(n219), .A1(keyfifo_merger_data[4]), .Z(fifo_in[4]));
Q_AN02 U409 ( .A0(n71), .A1(sha_tag_data[4]), .Z(n219));
Q_MX02 U410 ( .S(n70), .A0(n220), .A1(keyfifo_merger_data[3]), .Z(fifo_in[3]));
Q_AN02 U411 ( .A0(n71), .A1(sha_tag_data[3]), .Z(n220));
Q_MX02 U412 ( .S(n70), .A0(n221), .A1(keyfifo_merger_data[2]), .Z(fifo_in[2]));
Q_AN02 U413 ( .A0(n71), .A1(sha_tag_data[2]), .Z(n221));
Q_MX02 U414 ( .S(n70), .A0(n222), .A1(keyfifo_merger_data[1]), .Z(fifo_in[1]));
Q_AN02 U415 ( .A0(n71), .A1(sha_tag_data[1]), .Z(n222));
Q_MX02 U416 ( .S(n70), .A0(n223), .A1(keyfifo_merger_data[0]), .Z(fifo_in[0]));
Q_AN02 U417 ( .A0(n71), .A1(sha_tag_data[0]), .Z(n223));
Q_AN02 U418 ( .A0(cmdfifo_kdf_valid), .A1(n225), .Z(fifo_in_vld));
Q_AN03 U419 ( .A0(n224), .A1(n225), .A2(cmdfifo_kdf_valid), .Z(kdf_cmdfifo_ack));
Q_AN03 U420 ( .A0(in_counter[0]), .A1(n76), .A2(in_counter[2]), .Z(n224));
Q_MX02 U421 ( .S(n72), .A0(n226), .A1(sha_tag_valid), .Z(n225));
Q_ND03 U422 ( .A0(n76), .A1(in_counter[0]), .A2(in_counter[2]), .Z(n227));
Q_AN02 U423 ( .A0(n227), .A1(n230), .Z(n228));
Q_AN02 U424 ( .A0(n227), .A1(n232), .Z(n229));
Q_XOR2 U425 ( .A0(in_counter[2]), .A1(n231), .Z(n230));
Q_AD01HF U426 ( .A0(in_counter[1]), .B0(in_counter[0]), .S(n232), .CO(n231));
ixc_assign _zz_strnp_0 ( _zy_simnet_kdf_cmdfifo_ack_0_w$, kdf_cmdfifo_ack);
ixc_assign _zz_strnp_1 ( _zy_simnet_sha_tag_stall_1_w$, sha_tag_stall);
ixc_assign _zz_strnp_2 ( _zy_simnet_merger_keyfifo_ack_2_w$, 
	merger_keyfifo_ack);
ixc_assign_64 _zz_strnp_3 ( _zy_simnet_kdf_keybuilder_data_3_w$[0:63], 
	kdf_keybuilder_data[63:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_kdf_keybuilder_valid_4_w$, 
	kdf_keybuilder_valid);
ixc_assign_128 _zz_strnp_5 ( _zy_simnet_fifo_in_7_w$[0:127], fifo_in[127:0]);
ixc_assign _zz_strnp_6 ( _zy_simnet_fifo_in_vld_8_w$, fifo_in_vld);
ixc_assign _zz_strnp_7 ( _zy_simnet_fifo_out_ack_9_w$, fifo_out_ack);
cr_kme_fifo_xcm51 downsizer_fifo ( .fifo_in_stall( fifo_in_stall), 
	.fifo_out( fifo_out[127:0]), .fifo_out_valid( fifo_out_vld), 
	.fifo_overflow( _zy_simnet_dio_5), .fifo_underflow( 
	_zy_simnet_dio_6), .clk( clk), .rst_n( rst_n), .fifo_in( 
	_zy_simnet_fifo_in_7_w$[0:127]), .fifo_in_valid( 
	_zy_simnet_fifo_in_vld_8_w$), .fifo_out_ack( 
	_zy_simnet_fifo_out_ack_9_w$), .fifo_in_stall_override( 
	_zy_simnet_cio_10));
Q_FDP4EP \in_counter_REG[2] ( .CK(clk), .CE(merger_keyfifo_ack), .R(n233), .D(n228), .Q(in_counter[2]));
Q_INV U437 ( .A(rst_n), .Z(n233));
Q_INV U438 ( .A(in_counter[2]), .Z(n87));
Q_FDP4EP \in_counter_REG[1] ( .CK(clk), .CE(merger_keyfifo_ack), .R(n233), .D(n229), .Q(in_counter[1]));
Q_INV U440 ( .A(in_counter[1]), .Z(n76));
Q_INV U441 ( .A(in_counter[0]), .Z(n234));
Q_FDP4EP \in_counter_REG[0] ( .CK(clk), .CE(merger_keyfifo_ack), .R(n233), .D(n234), .Q(in_counter[0]));
Q_INV U443 ( .A(out_counter), .Z(n235));
Q_FDP4EP out_counter_REG  ( .CK(clk), .CE(n67), .R(n233), .D(n235), .Q(out_counter));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\cmdfifo_kdf_cmd.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\cmdfifo_kdf_cmd.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\cmdfifo_kdf_cmd.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\cmdfifo_kdf_cmd.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "4"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "cmdfifo_kdf_cmd 4 \cmdfifo_kdf_cmd.kdf_dek_iter  \cmdfifo_kdf_cmd.combo_mode  \cmdfifo_kdf_cmd.dek_key_op  \cmdfifo_kdf_cmd.dak_key_op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "1"
endmodule
