
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module axi_channel_reg_slice ( ready_src, valid_dst, payload_dst, aclk, aresetn, 
	valid_src, payload_src, ready_dst);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output ready_src;
output valid_dst;
output [81:0] payload_dst;
input aclk;
input aresetn;
input valid_src;
input [81:0] payload_src;
input ready_dst;
wire \full.c_wptr ;
wire [10:0] \full.c_rptr ;
wire \full.c_full ;
wire \full.c_empty ;
wire \full.r_wptr ;
wire [10:0] \full.r_rptr ;
wire \full.r_full ;
wire \full.r_empty ;
wire \full.r_enable ;
supply1 n97;
supply0 n99;
Q_MX02 U0 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][7] ), .A1(\full.r_payload[1][7] ), .Z(n1));
Q_MX02 U1 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][6] ), .A1(\full.r_payload[1][6] ), .Z(n2));
Q_MX02 U2 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][5] ), .A1(\full.r_payload[1][5] ), .Z(n3));
Q_MX02 U3 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][4] ), .A1(\full.r_payload[1][4] ), .Z(n4));
Q_MX02 U4 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][3] ), .A1(\full.r_payload[1][3] ), .Z(n5));
Q_MX02 U5 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][2] ), .A1(\full.r_payload[1][2] ), .Z(n6));
Q_MX02 U6 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][1] ), .A1(\full.r_payload[1][1] ), .Z(n7));
Q_MX02 U7 ( .S(\full.r_rptr [0]), .A0(\full.r_payload[0][0] ), .A1(\full.r_payload[1][0] ), .Z(n8));
Q_MX02 U8 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][15] ), .A1(\full.r_payload[1][15] ), .Z(n9));
Q_MX02 U9 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][14] ), .A1(\full.r_payload[1][14] ), .Z(n10));
Q_MX02 U10 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][13] ), .A1(\full.r_payload[1][13] ), .Z(n11));
Q_MX02 U11 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][12] ), .A1(\full.r_payload[1][12] ), .Z(n12));
Q_MX02 U12 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][11] ), .A1(\full.r_payload[1][11] ), .Z(n13));
Q_MX02 U13 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][10] ), .A1(\full.r_payload[1][10] ), .Z(n14));
Q_MX02 U14 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][9] ), .A1(\full.r_payload[1][9] ), .Z(n15));
Q_MX02 U15 ( .S(\full.r_rptr [1]), .A0(\full.r_payload[0][8] ), .A1(\full.r_payload[1][8] ), .Z(n16));
Q_MX02 U16 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][23] ), .A1(\full.r_payload[1][23] ), .Z(n17));
Q_MX02 U17 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][22] ), .A1(\full.r_payload[1][22] ), .Z(n18));
Q_MX02 U18 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][21] ), .A1(\full.r_payload[1][21] ), .Z(n19));
Q_MX02 U19 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][20] ), .A1(\full.r_payload[1][20] ), .Z(n20));
Q_MX02 U20 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][19] ), .A1(\full.r_payload[1][19] ), .Z(n21));
Q_MX02 U21 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][18] ), .A1(\full.r_payload[1][18] ), .Z(n22));
Q_MX02 U22 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][17] ), .A1(\full.r_payload[1][17] ), .Z(n23));
Q_MX02 U23 ( .S(\full.r_rptr [2]), .A0(\full.r_payload[0][16] ), .A1(\full.r_payload[1][16] ), .Z(n24));
Q_MX02 U24 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][31] ), .A1(\full.r_payload[1][31] ), .Z(n25));
Q_MX02 U25 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][30] ), .A1(\full.r_payload[1][30] ), .Z(n26));
Q_MX02 U26 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][29] ), .A1(\full.r_payload[1][29] ), .Z(n27));
Q_MX02 U27 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][28] ), .A1(\full.r_payload[1][28] ), .Z(n28));
Q_MX02 U28 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][27] ), .A1(\full.r_payload[1][27] ), .Z(n29));
Q_MX02 U29 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][26] ), .A1(\full.r_payload[1][26] ), .Z(n30));
Q_MX02 U30 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][25] ), .A1(\full.r_payload[1][25] ), .Z(n31));
Q_MX02 U31 ( .S(\full.r_rptr [3]), .A0(\full.r_payload[0][24] ), .A1(\full.r_payload[1][24] ), .Z(n32));
Q_MX02 U32 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][39] ), .A1(\full.r_payload[1][39] ), .Z(n33));
Q_MX02 U33 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][38] ), .A1(\full.r_payload[1][38] ), .Z(n34));
Q_MX02 U34 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][37] ), .A1(\full.r_payload[1][37] ), .Z(n35));
Q_MX02 U35 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][36] ), .A1(\full.r_payload[1][36] ), .Z(n36));
Q_MX02 U36 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][35] ), .A1(\full.r_payload[1][35] ), .Z(n37));
Q_MX02 U37 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][34] ), .A1(\full.r_payload[1][34] ), .Z(n38));
Q_MX02 U38 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][33] ), .A1(\full.r_payload[1][33] ), .Z(n39));
Q_MX02 U39 ( .S(\full.r_rptr [4]), .A0(\full.r_payload[0][32] ), .A1(\full.r_payload[1][32] ), .Z(n40));
Q_MX02 U40 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][47] ), .A1(\full.r_payload[1][47] ), .Z(n41));
Q_MX02 U41 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][46] ), .A1(\full.r_payload[1][46] ), .Z(n42));
Q_MX02 U42 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][45] ), .A1(\full.r_payload[1][45] ), .Z(n43));
Q_MX02 U43 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][44] ), .A1(\full.r_payload[1][44] ), .Z(n44));
Q_MX02 U44 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][43] ), .A1(\full.r_payload[1][43] ), .Z(n45));
Q_MX02 U45 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][42] ), .A1(\full.r_payload[1][42] ), .Z(n46));
Q_MX02 U46 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][41] ), .A1(\full.r_payload[1][41] ), .Z(n47));
Q_MX02 U47 ( .S(\full.r_rptr [5]), .A0(\full.r_payload[0][40] ), .A1(\full.r_payload[1][40] ), .Z(n48));
Q_MX02 U48 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][55] ), .A1(\full.r_payload[1][55] ), .Z(n49));
Q_MX02 U49 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][54] ), .A1(\full.r_payload[1][54] ), .Z(n50));
Q_MX02 U50 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][53] ), .A1(\full.r_payload[1][53] ), .Z(n51));
Q_MX02 U51 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][52] ), .A1(\full.r_payload[1][52] ), .Z(n52));
Q_MX02 U52 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][51] ), .A1(\full.r_payload[1][51] ), .Z(n53));
Q_MX02 U53 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][50] ), .A1(\full.r_payload[1][50] ), .Z(n54));
Q_MX02 U54 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][49] ), .A1(\full.r_payload[1][49] ), .Z(n55));
Q_MX02 U55 ( .S(\full.r_rptr [6]), .A0(\full.r_payload[0][48] ), .A1(\full.r_payload[1][48] ), .Z(n56));
Q_MX02 U56 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][63] ), .A1(\full.r_payload[1][63] ), .Z(n57));
Q_MX02 U57 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][62] ), .A1(\full.r_payload[1][62] ), .Z(n58));
Q_MX02 U58 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][61] ), .A1(\full.r_payload[1][61] ), .Z(n59));
Q_MX02 U59 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][60] ), .A1(\full.r_payload[1][60] ), .Z(n60));
Q_MX02 U60 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][59] ), .A1(\full.r_payload[1][59] ), .Z(n61));
Q_MX02 U61 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][58] ), .A1(\full.r_payload[1][58] ), .Z(n62));
Q_MX02 U62 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][57] ), .A1(\full.r_payload[1][57] ), .Z(n63));
Q_MX02 U63 ( .S(\full.r_rptr [7]), .A0(\full.r_payload[0][56] ), .A1(\full.r_payload[1][56] ), .Z(n64));
Q_MX02 U64 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][71] ), .A1(\full.r_payload[1][71] ), .Z(n65));
Q_MX02 U65 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][70] ), .A1(\full.r_payload[1][70] ), .Z(n66));
Q_MX02 U66 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][69] ), .A1(\full.r_payload[1][69] ), .Z(n67));
Q_MX02 U67 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][68] ), .A1(\full.r_payload[1][68] ), .Z(n68));
Q_MX02 U68 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][67] ), .A1(\full.r_payload[1][67] ), .Z(n69));
Q_MX02 U69 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][66] ), .A1(\full.r_payload[1][66] ), .Z(n70));
Q_MX02 U70 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][65] ), .A1(\full.r_payload[1][65] ), .Z(n71));
Q_MX02 U71 ( .S(\full.r_rptr [8]), .A0(\full.r_payload[0][64] ), .A1(\full.r_payload[1][64] ), .Z(n72));
Q_MX02 U72 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][79] ), .A1(\full.r_payload[1][79] ), .Z(n73));
Q_MX02 U73 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][78] ), .A1(\full.r_payload[1][78] ), .Z(n74));
Q_MX02 U74 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][77] ), .A1(\full.r_payload[1][77] ), .Z(n75));
Q_MX02 U75 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][76] ), .A1(\full.r_payload[1][76] ), .Z(n76));
Q_MX02 U76 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][75] ), .A1(\full.r_payload[1][75] ), .Z(n77));
Q_MX02 U77 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][74] ), .A1(\full.r_payload[1][74] ), .Z(n78));
Q_MX02 U78 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][73] ), .A1(\full.r_payload[1][73] ), .Z(n79));
Q_MX02 U79 ( .S(\full.r_rptr [9]), .A0(\full.r_payload[0][72] ), .A1(\full.r_payload[1][72] ), .Z(n80));
Q_MX02 U80 ( .S(\full.r_rptr [10]), .A0(\full.r_payload[0][81] ), .A1(\full.r_payload[1][81] ), .Z(n81));
Q_MX02 U81 ( .S(\full.r_rptr [10]), .A0(\full.r_payload[0][80] ), .A1(\full.r_payload[1][80] ), .Z(n82));
Q_AN02 U82 ( .A0(n84), .A1(n98), .Z(n83));
Q_INV U83 ( .A(n85), .Z(n84));
Q_AN02 U84 ( .A0(\full.r_wptr ), .A1(n98), .Z(n85));
ixc_assign_8 \full.genblk1_0_.genblk1._zz_strnp_0 ( payload_dst[7:0], { n1, 
	n2, n3, n4, n5, n6, n7, n8});
ixc_assign_8 \full.genblk1_1_.genblk1._zz_strnp_1 ( payload_dst[15:8], { n9, 
	n10, n11, n12, n13, n14, n15, n16});
ixc_assign_8 \full.genblk1_2_.genblk1._zz_strnp_2 ( payload_dst[23:16], { n17, 
	n18, n19, n20, n21, n22, n23, n24});
ixc_assign_8 \full.genblk1_3_.genblk1._zz_strnp_3 ( payload_dst[31:24], { n25, 
	n26, n27, n28, n29, n30, n31, n32});
ixc_assign_8 \full.genblk1_4_.genblk1._zz_strnp_4 ( payload_dst[39:32], { n33, 
	n34, n35, n36, n37, n38, n39, n40});
ixc_assign_8 \full.genblk1_5_.genblk1._zz_strnp_5 ( payload_dst[47:40], { n41, 
	n42, n43, n44, n45, n46, n47, n48});
ixc_assign_8 \full.genblk1_6_.genblk1._zz_strnp_6 ( payload_dst[55:48], { n49, 
	n50, n51, n52, n53, n54, n55, n56});
ixc_assign_8 \full.genblk1_7_.genblk1._zz_strnp_7 ( payload_dst[63:56], { n57, 
	n58, n59, n60, n61, n62, n63, n64});
ixc_assign_8 \full.genblk1_8_.genblk1._zz_strnp_8 ( payload_dst[71:64], { n65, 
	n66, n67, n68, n69, n70, n71, n72});
ixc_assign_8 \full.genblk1_9_.genblk1._zz_strnp_9 ( payload_dst[79:72], { n73, 
	n74, n75, n76, n77, n78, n79, n80});
ixc_assign_2 \full.genblk1_10_.genblk1._zz_strnp_10 ( payload_dst[81:80], { 
	n81, n82});
Q_AN03 U96 ( .A0(ready_src), .A1(n86), .A2(valid_src), .Z(n90));
Q_AN02 U97 ( .A0(valid_dst), .A1(ready_dst), .Z(n96));
Q_AO21 U98 ( .A0(n96), .A1(\full.r_full ), .B0(n90), .Z(n87));
Q_INV U99 ( .A(ready_src), .Z(n91));
Q_OR03 U100 ( .A0(n91), .A1(n86), .A2(n92), .Z(n93));
Q_INV U101 ( .A(valid_src), .Z(n92));
Q_AO21 U102 ( .A0(n93), .A1(n96), .B0(n88), .Z(n94));
Q_INV U103 ( .A(n93), .Z(n88));
Q_INV U104 ( .A(n98), .Z(n89));
Q_AO21 U105 ( .A0(n96), .A1(n95), .B0(\full.r_empty ), .Z(n86));
Q_XOR2 U106 ( .A0(n98), .A1(\full.r_wptr ), .Z(\full.c_wptr ));
Q_XOR2 U107 ( .A0(n87), .A1(\full.r_rptr [10]), .Z(\full.c_rptr [10]));
Q_XOR2 U108 ( .A0(n87), .A1(\full.r_rptr [9]), .Z(\full.c_rptr [9]));
Q_XOR2 U109 ( .A0(n87), .A1(\full.r_rptr [8]), .Z(\full.c_rptr [8]));
Q_XOR2 U110 ( .A0(n87), .A1(\full.r_rptr [7]), .Z(\full.c_rptr [7]));
Q_XOR2 U111 ( .A0(n87), .A1(\full.r_rptr [6]), .Z(\full.c_rptr [6]));
Q_XOR2 U112 ( .A0(n87), .A1(\full.r_rptr [5]), .Z(\full.c_rptr [5]));
Q_XOR2 U113 ( .A0(n87), .A1(\full.r_rptr [4]), .Z(\full.c_rptr [4]));
Q_XOR2 U114 ( .A0(n87), .A1(\full.r_rptr [3]), .Z(\full.c_rptr [3]));
Q_XOR2 U115 ( .A0(n87), .A1(\full.r_rptr [2]), .Z(\full.c_rptr [2]));
Q_XOR2 U116 ( .A0(n87), .A1(\full.r_rptr [1]), .Z(\full.c_rptr [1]));
Q_XOR2 U117 ( .A0(n87), .A1(\full.r_rptr [0]), .Z(\full.c_rptr [0]));
Q_MX02 U118 ( .S(n94), .A0(\full.r_full ), .A1(n88), .Z(\full.c_full ));
Q_AN02 U119 ( .A0(n89), .A1(n86), .Z(\full.c_empty ));
Q_FDP1 \full.r_enable_REG ( .CK(aclk), .R(aresetn), .D(n97), .Q(\full.r_enable ), .QN( ));
Q_FDP1 \full.r_full_REG ( .CK(aclk), .R(aresetn), .D(\full.c_full ), .Q(\full.r_full ), .QN(n95));
Q_FDP2 \full.r_empty_REG ( .CK(aclk), .S(aresetn), .D(\full.c_empty ), .Q(\full.r_empty ), .QN(valid_dst));
Q_FDP2 \full.r_rptr_REG[10] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [10]), .Q(\full.r_rptr [10]), .QN( ));
Q_FDP2 \full.r_rptr_REG[9] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [9]), .Q(\full.r_rptr [9]), .QN( ));
Q_FDP2 \full.r_rptr_REG[8] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [8]), .Q(\full.r_rptr [8]), .QN( ));
Q_FDP2 \full.r_rptr_REG[7] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [7]), .Q(\full.r_rptr [7]), .QN( ));
Q_FDP2 \full.r_rptr_REG[6] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [6]), .Q(\full.r_rptr [6]), .QN( ));
Q_FDP2 \full.r_rptr_REG[5] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [5]), .Q(\full.r_rptr [5]), .QN( ));
Q_FDP2 \full.r_rptr_REG[4] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [4]), .Q(\full.r_rptr [4]), .QN( ));
Q_FDP2 \full.r_rptr_REG[3] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [3]), .Q(\full.r_rptr [3]), .QN( ));
Q_FDP2 \full.r_rptr_REG[2] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [2]), .Q(\full.r_rptr [2]), .QN( ));
Q_FDP2 \full.r_rptr_REG[1] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [1]), .Q(\full.r_rptr [1]), .QN( ));
Q_FDP2 \full.r_rptr_REG[0] ( .CK(aclk), .S(aresetn), .D(\full.c_rptr [0]), .Q(\full.r_rptr [0]), .QN( ));
Q_FDP1 \full.r_wptr_REG ( .CK(aclk), .R(aresetn), .D(\full.c_wptr ), .Q(\full.r_wptr ), .QN( ));
Q_AN02 U135 ( .A0(valid_src), .A1(ready_src), .Z(n98));
Q_AN02 U136 ( .A0(\full.r_enable ), .A1(n95), .Z(ready_src));
Q_FDP4EP \full.r_payload_REG[0][0] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[0]), .Q(\full.r_payload[0][0] ));
Q_FDP4EP \full.r_payload_REG[0][1] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[1]), .Q(\full.r_payload[0][1] ));
Q_FDP4EP \full.r_payload_REG[0][2] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[2]), .Q(\full.r_payload[0][2] ));
Q_FDP4EP \full.r_payload_REG[0][3] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[3]), .Q(\full.r_payload[0][3] ));
Q_FDP4EP \full.r_payload_REG[0][4] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[4]), .Q(\full.r_payload[0][4] ));
Q_FDP4EP \full.r_payload_REG[0][5] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[5]), .Q(\full.r_payload[0][5] ));
Q_FDP4EP \full.r_payload_REG[0][6] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[6]), .Q(\full.r_payload[0][6] ));
Q_FDP4EP \full.r_payload_REG[0][7] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[7]), .Q(\full.r_payload[0][7] ));
Q_FDP4EP \full.r_payload_REG[0][8] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[8]), .Q(\full.r_payload[0][8] ));
Q_FDP4EP \full.r_payload_REG[0][9] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[9]), .Q(\full.r_payload[0][9] ));
Q_FDP4EP \full.r_payload_REG[0][10] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[10]), .Q(\full.r_payload[0][10] ));
Q_FDP4EP \full.r_payload_REG[0][11] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[11]), .Q(\full.r_payload[0][11] ));
Q_FDP4EP \full.r_payload_REG[0][12] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[12]), .Q(\full.r_payload[0][12] ));
Q_FDP4EP \full.r_payload_REG[0][13] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[13]), .Q(\full.r_payload[0][13] ));
Q_FDP4EP \full.r_payload_REG[0][14] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[14]), .Q(\full.r_payload[0][14] ));
Q_FDP4EP \full.r_payload_REG[0][15] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[15]), .Q(\full.r_payload[0][15] ));
Q_FDP4EP \full.r_payload_REG[0][16] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[16]), .Q(\full.r_payload[0][16] ));
Q_FDP4EP \full.r_payload_REG[0][17] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[17]), .Q(\full.r_payload[0][17] ));
Q_FDP4EP \full.r_payload_REG[0][18] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[18]), .Q(\full.r_payload[0][18] ));
Q_FDP4EP \full.r_payload_REG[0][19] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[19]), .Q(\full.r_payload[0][19] ));
Q_FDP4EP \full.r_payload_REG[0][20] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[20]), .Q(\full.r_payload[0][20] ));
Q_FDP4EP \full.r_payload_REG[0][21] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[21]), .Q(\full.r_payload[0][21] ));
Q_FDP4EP \full.r_payload_REG[0][22] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[22]), .Q(\full.r_payload[0][22] ));
Q_FDP4EP \full.r_payload_REG[0][23] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[23]), .Q(\full.r_payload[0][23] ));
Q_FDP4EP \full.r_payload_REG[0][24] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[24]), .Q(\full.r_payload[0][24] ));
Q_FDP4EP \full.r_payload_REG[0][25] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[25]), .Q(\full.r_payload[0][25] ));
Q_FDP4EP \full.r_payload_REG[0][26] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[26]), .Q(\full.r_payload[0][26] ));
Q_FDP4EP \full.r_payload_REG[0][27] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[27]), .Q(\full.r_payload[0][27] ));
Q_FDP4EP \full.r_payload_REG[0][28] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[28]), .Q(\full.r_payload[0][28] ));
Q_FDP4EP \full.r_payload_REG[0][29] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[29]), .Q(\full.r_payload[0][29] ));
Q_FDP4EP \full.r_payload_REG[0][30] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[30]), .Q(\full.r_payload[0][30] ));
Q_FDP4EP \full.r_payload_REG[0][31] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[31]), .Q(\full.r_payload[0][31] ));
Q_FDP4EP \full.r_payload_REG[0][32] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[32]), .Q(\full.r_payload[0][32] ));
Q_FDP4EP \full.r_payload_REG[0][33] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[33]), .Q(\full.r_payload[0][33] ));
Q_FDP4EP \full.r_payload_REG[0][34] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[34]), .Q(\full.r_payload[0][34] ));
Q_FDP4EP \full.r_payload_REG[0][35] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[35]), .Q(\full.r_payload[0][35] ));
Q_FDP4EP \full.r_payload_REG[0][36] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[36]), .Q(\full.r_payload[0][36] ));
Q_FDP4EP \full.r_payload_REG[0][37] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[37]), .Q(\full.r_payload[0][37] ));
Q_FDP4EP \full.r_payload_REG[0][38] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[38]), .Q(\full.r_payload[0][38] ));
Q_FDP4EP \full.r_payload_REG[0][39] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[39]), .Q(\full.r_payload[0][39] ));
Q_FDP4EP \full.r_payload_REG[0][40] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[40]), .Q(\full.r_payload[0][40] ));
Q_FDP4EP \full.r_payload_REG[0][41] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[41]), .Q(\full.r_payload[0][41] ));
Q_FDP4EP \full.r_payload_REG[0][42] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[42]), .Q(\full.r_payload[0][42] ));
Q_FDP4EP \full.r_payload_REG[0][43] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[43]), .Q(\full.r_payload[0][43] ));
Q_FDP4EP \full.r_payload_REG[0][44] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[44]), .Q(\full.r_payload[0][44] ));
Q_FDP4EP \full.r_payload_REG[0][45] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[45]), .Q(\full.r_payload[0][45] ));
Q_FDP4EP \full.r_payload_REG[0][46] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[46]), .Q(\full.r_payload[0][46] ));
Q_FDP4EP \full.r_payload_REG[0][47] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[47]), .Q(\full.r_payload[0][47] ));
Q_FDP4EP \full.r_payload_REG[0][48] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[48]), .Q(\full.r_payload[0][48] ));
Q_FDP4EP \full.r_payload_REG[0][49] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[49]), .Q(\full.r_payload[0][49] ));
Q_FDP4EP \full.r_payload_REG[0][50] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[50]), .Q(\full.r_payload[0][50] ));
Q_FDP4EP \full.r_payload_REG[0][51] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[51]), .Q(\full.r_payload[0][51] ));
Q_FDP4EP \full.r_payload_REG[0][52] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[52]), .Q(\full.r_payload[0][52] ));
Q_FDP4EP \full.r_payload_REG[0][53] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[53]), .Q(\full.r_payload[0][53] ));
Q_FDP4EP \full.r_payload_REG[0][54] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[54]), .Q(\full.r_payload[0][54] ));
Q_FDP4EP \full.r_payload_REG[0][55] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[55]), .Q(\full.r_payload[0][55] ));
Q_FDP4EP \full.r_payload_REG[0][56] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[56]), .Q(\full.r_payload[0][56] ));
Q_FDP4EP \full.r_payload_REG[0][57] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[57]), .Q(\full.r_payload[0][57] ));
Q_FDP4EP \full.r_payload_REG[0][58] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[58]), .Q(\full.r_payload[0][58] ));
Q_FDP4EP \full.r_payload_REG[0][59] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[59]), .Q(\full.r_payload[0][59] ));
Q_FDP4EP \full.r_payload_REG[0][60] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[60]), .Q(\full.r_payload[0][60] ));
Q_FDP4EP \full.r_payload_REG[0][61] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[61]), .Q(\full.r_payload[0][61] ));
Q_FDP4EP \full.r_payload_REG[0][62] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[62]), .Q(\full.r_payload[0][62] ));
Q_FDP4EP \full.r_payload_REG[0][63] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[63]), .Q(\full.r_payload[0][63] ));
Q_FDP4EP \full.r_payload_REG[0][64] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[64]), .Q(\full.r_payload[0][64] ));
Q_FDP4EP \full.r_payload_REG[0][65] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[65]), .Q(\full.r_payload[0][65] ));
Q_FDP4EP \full.r_payload_REG[0][66] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[66]), .Q(\full.r_payload[0][66] ));
Q_FDP4EP \full.r_payload_REG[0][67] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[67]), .Q(\full.r_payload[0][67] ));
Q_FDP4EP \full.r_payload_REG[0][68] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[68]), .Q(\full.r_payload[0][68] ));
Q_FDP4EP \full.r_payload_REG[0][69] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[69]), .Q(\full.r_payload[0][69] ));
Q_FDP4EP \full.r_payload_REG[0][70] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[70]), .Q(\full.r_payload[0][70] ));
Q_FDP4EP \full.r_payload_REG[0][71] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[71]), .Q(\full.r_payload[0][71] ));
Q_FDP4EP \full.r_payload_REG[0][72] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[72]), .Q(\full.r_payload[0][72] ));
Q_FDP4EP \full.r_payload_REG[0][73] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[73]), .Q(\full.r_payload[0][73] ));
Q_FDP4EP \full.r_payload_REG[0][74] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[74]), .Q(\full.r_payload[0][74] ));
Q_FDP4EP \full.r_payload_REG[0][75] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[75]), .Q(\full.r_payload[0][75] ));
Q_FDP4EP \full.r_payload_REG[0][76] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[76]), .Q(\full.r_payload[0][76] ));
Q_FDP4EP \full.r_payload_REG[0][77] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[77]), .Q(\full.r_payload[0][77] ));
Q_FDP4EP \full.r_payload_REG[0][78] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[78]), .Q(\full.r_payload[0][78] ));
Q_FDP4EP \full.r_payload_REG[0][79] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[79]), .Q(\full.r_payload[0][79] ));
Q_FDP4EP \full.r_payload_REG[0][80] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[80]), .Q(\full.r_payload[0][80] ));
Q_FDP4EP \full.r_payload_REG[0][81] ( .CK(aclk), .CE(n83), .R(n99), .D(payload_src[81]), .Q(\full.r_payload[0][81] ));
Q_FDP4EP \full.r_payload_REG[1][0] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[0]), .Q(\full.r_payload[1][0] ));
Q_FDP4EP \full.r_payload_REG[1][1] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[1]), .Q(\full.r_payload[1][1] ));
Q_FDP4EP \full.r_payload_REG[1][2] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[2]), .Q(\full.r_payload[1][2] ));
Q_FDP4EP \full.r_payload_REG[1][3] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[3]), .Q(\full.r_payload[1][3] ));
Q_FDP4EP \full.r_payload_REG[1][4] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[4]), .Q(\full.r_payload[1][4] ));
Q_FDP4EP \full.r_payload_REG[1][5] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[5]), .Q(\full.r_payload[1][5] ));
Q_FDP4EP \full.r_payload_REG[1][6] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[6]), .Q(\full.r_payload[1][6] ));
Q_FDP4EP \full.r_payload_REG[1][7] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[7]), .Q(\full.r_payload[1][7] ));
Q_FDP4EP \full.r_payload_REG[1][8] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[8]), .Q(\full.r_payload[1][8] ));
Q_FDP4EP \full.r_payload_REG[1][9] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[9]), .Q(\full.r_payload[1][9] ));
Q_FDP4EP \full.r_payload_REG[1][10] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[10]), .Q(\full.r_payload[1][10] ));
Q_FDP4EP \full.r_payload_REG[1][11] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[11]), .Q(\full.r_payload[1][11] ));
Q_FDP4EP \full.r_payload_REG[1][12] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[12]), .Q(\full.r_payload[1][12] ));
Q_FDP4EP \full.r_payload_REG[1][13] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[13]), .Q(\full.r_payload[1][13] ));
Q_FDP4EP \full.r_payload_REG[1][14] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[14]), .Q(\full.r_payload[1][14] ));
Q_FDP4EP \full.r_payload_REG[1][15] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[15]), .Q(\full.r_payload[1][15] ));
Q_FDP4EP \full.r_payload_REG[1][16] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[16]), .Q(\full.r_payload[1][16] ));
Q_FDP4EP \full.r_payload_REG[1][17] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[17]), .Q(\full.r_payload[1][17] ));
Q_FDP4EP \full.r_payload_REG[1][18] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[18]), .Q(\full.r_payload[1][18] ));
Q_FDP4EP \full.r_payload_REG[1][19] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[19]), .Q(\full.r_payload[1][19] ));
Q_FDP4EP \full.r_payload_REG[1][20] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[20]), .Q(\full.r_payload[1][20] ));
Q_FDP4EP \full.r_payload_REG[1][21] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[21]), .Q(\full.r_payload[1][21] ));
Q_FDP4EP \full.r_payload_REG[1][22] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[22]), .Q(\full.r_payload[1][22] ));
Q_FDP4EP \full.r_payload_REG[1][23] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[23]), .Q(\full.r_payload[1][23] ));
Q_FDP4EP \full.r_payload_REG[1][24] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[24]), .Q(\full.r_payload[1][24] ));
Q_FDP4EP \full.r_payload_REG[1][25] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[25]), .Q(\full.r_payload[1][25] ));
Q_FDP4EP \full.r_payload_REG[1][26] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[26]), .Q(\full.r_payload[1][26] ));
Q_FDP4EP \full.r_payload_REG[1][27] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[27]), .Q(\full.r_payload[1][27] ));
Q_FDP4EP \full.r_payload_REG[1][28] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[28]), .Q(\full.r_payload[1][28] ));
Q_FDP4EP \full.r_payload_REG[1][29] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[29]), .Q(\full.r_payload[1][29] ));
Q_FDP4EP \full.r_payload_REG[1][30] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[30]), .Q(\full.r_payload[1][30] ));
Q_FDP4EP \full.r_payload_REG[1][31] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[31]), .Q(\full.r_payload[1][31] ));
Q_FDP4EP \full.r_payload_REG[1][32] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[32]), .Q(\full.r_payload[1][32] ));
Q_FDP4EP \full.r_payload_REG[1][33] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[33]), .Q(\full.r_payload[1][33] ));
Q_FDP4EP \full.r_payload_REG[1][34] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[34]), .Q(\full.r_payload[1][34] ));
Q_FDP4EP \full.r_payload_REG[1][35] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[35]), .Q(\full.r_payload[1][35] ));
Q_FDP4EP \full.r_payload_REG[1][36] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[36]), .Q(\full.r_payload[1][36] ));
Q_FDP4EP \full.r_payload_REG[1][37] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[37]), .Q(\full.r_payload[1][37] ));
Q_FDP4EP \full.r_payload_REG[1][38] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[38]), .Q(\full.r_payload[1][38] ));
Q_FDP4EP \full.r_payload_REG[1][39] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[39]), .Q(\full.r_payload[1][39] ));
Q_FDP4EP \full.r_payload_REG[1][40] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[40]), .Q(\full.r_payload[1][40] ));
Q_FDP4EP \full.r_payload_REG[1][41] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[41]), .Q(\full.r_payload[1][41] ));
Q_FDP4EP \full.r_payload_REG[1][42] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[42]), .Q(\full.r_payload[1][42] ));
Q_FDP4EP \full.r_payload_REG[1][43] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[43]), .Q(\full.r_payload[1][43] ));
Q_FDP4EP \full.r_payload_REG[1][44] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[44]), .Q(\full.r_payload[1][44] ));
Q_FDP4EP \full.r_payload_REG[1][45] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[45]), .Q(\full.r_payload[1][45] ));
Q_FDP4EP \full.r_payload_REG[1][46] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[46]), .Q(\full.r_payload[1][46] ));
Q_FDP4EP \full.r_payload_REG[1][47] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[47]), .Q(\full.r_payload[1][47] ));
Q_FDP4EP \full.r_payload_REG[1][48] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[48]), .Q(\full.r_payload[1][48] ));
Q_FDP4EP \full.r_payload_REG[1][49] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[49]), .Q(\full.r_payload[1][49] ));
Q_FDP4EP \full.r_payload_REG[1][50] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[50]), .Q(\full.r_payload[1][50] ));
Q_FDP4EP \full.r_payload_REG[1][51] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[51]), .Q(\full.r_payload[1][51] ));
Q_FDP4EP \full.r_payload_REG[1][52] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[52]), .Q(\full.r_payload[1][52] ));
Q_FDP4EP \full.r_payload_REG[1][53] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[53]), .Q(\full.r_payload[1][53] ));
Q_FDP4EP \full.r_payload_REG[1][54] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[54]), .Q(\full.r_payload[1][54] ));
Q_FDP4EP \full.r_payload_REG[1][55] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[55]), .Q(\full.r_payload[1][55] ));
Q_FDP4EP \full.r_payload_REG[1][56] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[56]), .Q(\full.r_payload[1][56] ));
Q_FDP4EP \full.r_payload_REG[1][57] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[57]), .Q(\full.r_payload[1][57] ));
Q_FDP4EP \full.r_payload_REG[1][58] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[58]), .Q(\full.r_payload[1][58] ));
Q_FDP4EP \full.r_payload_REG[1][59] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[59]), .Q(\full.r_payload[1][59] ));
Q_FDP4EP \full.r_payload_REG[1][60] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[60]), .Q(\full.r_payload[1][60] ));
Q_FDP4EP \full.r_payload_REG[1][61] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[61]), .Q(\full.r_payload[1][61] ));
Q_FDP4EP \full.r_payload_REG[1][62] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[62]), .Q(\full.r_payload[1][62] ));
Q_FDP4EP \full.r_payload_REG[1][63] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[63]), .Q(\full.r_payload[1][63] ));
Q_FDP4EP \full.r_payload_REG[1][64] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[64]), .Q(\full.r_payload[1][64] ));
Q_FDP4EP \full.r_payload_REG[1][65] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[65]), .Q(\full.r_payload[1][65] ));
Q_FDP4EP \full.r_payload_REG[1][66] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[66]), .Q(\full.r_payload[1][66] ));
Q_FDP4EP \full.r_payload_REG[1][67] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[67]), .Q(\full.r_payload[1][67] ));
Q_FDP4EP \full.r_payload_REG[1][68] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[68]), .Q(\full.r_payload[1][68] ));
Q_FDP4EP \full.r_payload_REG[1][69] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[69]), .Q(\full.r_payload[1][69] ));
Q_FDP4EP \full.r_payload_REG[1][70] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[70]), .Q(\full.r_payload[1][70] ));
Q_FDP4EP \full.r_payload_REG[1][71] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[71]), .Q(\full.r_payload[1][71] ));
Q_FDP4EP \full.r_payload_REG[1][72] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[72]), .Q(\full.r_payload[1][72] ));
Q_FDP4EP \full.r_payload_REG[1][73] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[73]), .Q(\full.r_payload[1][73] ));
Q_FDP4EP \full.r_payload_REG[1][74] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[74]), .Q(\full.r_payload[1][74] ));
Q_FDP4EP \full.r_payload_REG[1][75] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[75]), .Q(\full.r_payload[1][75] ));
Q_FDP4EP \full.r_payload_REG[1][76] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[76]), .Q(\full.r_payload[1][76] ));
Q_FDP4EP \full.r_payload_REG[1][77] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[77]), .Q(\full.r_payload[1][77] ));
Q_FDP4EP \full.r_payload_REG[1][78] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[78]), .Q(\full.r_payload[1][78] ));
Q_FDP4EP \full.r_payload_REG[1][79] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[79]), .Q(\full.r_payload[1][79] ));
Q_FDP4EP \full.r_payload_REG[1][80] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[80]), .Q(\full.r_payload[1][80] ));
Q_FDP4EP \full.r_payload_REG[1][81] ( .CK(aclk), .CE(n85), .R(n99), .D(payload_src[81]), .Q(\full.r_payload[1][81] ));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "\full.r_payload  1 81 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_2 "1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 genblk1 0 10 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 full  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[10].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[10]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[9].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[9]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[8].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[8]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[7].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[7]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[6].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[6]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[5].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[5]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[4].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[4]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[3].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[2].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[1].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[0].genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full.genblk1[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "full"
endmodule
