
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_tlvp2_rsm ( pt_ob_rd, usr_ob_full, usr_ob_afull, tlvp_ob_empty, 
	tlvp_ob_aempty, .tlvp_ob( {\tlvp_ob.tvalid , \tlvp_ob.tlast , 
	\tlvp_ob.tid [0], \tlvp_ob.tstrb [7], \tlvp_ob.tstrb [6], 
	\tlvp_ob.tstrb [5], \tlvp_ob.tstrb [4], \tlvp_ob.tstrb [3], 
	\tlvp_ob.tstrb [2], \tlvp_ob.tstrb [1], \tlvp_ob.tstrb [0], 
	\tlvp_ob.tuser [7], \tlvp_ob.tuser [6], \tlvp_ob.tuser [5], 
	\tlvp_ob.tuser [4], \tlvp_ob.tuser [3], \tlvp_ob.tuser [2], 
	\tlvp_ob.tuser [1], \tlvp_ob.tuser [0], \tlvp_ob.tdata [63], 
	\tlvp_ob.tdata [62], \tlvp_ob.tdata [61], \tlvp_ob.tdata [60], 
	\tlvp_ob.tdata [59], \tlvp_ob.tdata [58], \tlvp_ob.tdata [57], 
	\tlvp_ob.tdata [56], \tlvp_ob.tdata [55], \tlvp_ob.tdata [54], 
	\tlvp_ob.tdata [53], \tlvp_ob.tdata [52], \tlvp_ob.tdata [51], 
	\tlvp_ob.tdata [50], \tlvp_ob.tdata [49], \tlvp_ob.tdata [48], 
	\tlvp_ob.tdata [47], \tlvp_ob.tdata [46], \tlvp_ob.tdata [45], 
	\tlvp_ob.tdata [44], \tlvp_ob.tdata [43], \tlvp_ob.tdata [42], 
	\tlvp_ob.tdata [41], \tlvp_ob.tdata [40], \tlvp_ob.tdata [39], 
	\tlvp_ob.tdata [38], \tlvp_ob.tdata [37], \tlvp_ob.tdata [36], 
	\tlvp_ob.tdata [35], \tlvp_ob.tdata [34], \tlvp_ob.tdata [33], 
	\tlvp_ob.tdata [32], \tlvp_ob.tdata [31], \tlvp_ob.tdata [30], 
	\tlvp_ob.tdata [29], \tlvp_ob.tdata [28], \tlvp_ob.tdata [27], 
	\tlvp_ob.tdata [26], \tlvp_ob.tdata [25], \tlvp_ob.tdata [24], 
	\tlvp_ob.tdata [23], \tlvp_ob.tdata [22], \tlvp_ob.tdata [21], 
	\tlvp_ob.tdata [20], \tlvp_ob.tdata [19], \tlvp_ob.tdata [18], 
	\tlvp_ob.tdata [17], \tlvp_ob.tdata [16], \tlvp_ob.tdata [15], 
	\tlvp_ob.tdata [14], \tlvp_ob.tdata [13], \tlvp_ob.tdata [12], 
	\tlvp_ob.tdata [11], \tlvp_ob.tdata [10], \tlvp_ob.tdata [9], 
	\tlvp_ob.tdata [8], \tlvp_ob.tdata [7], \tlvp_ob.tdata [6], 
	\tlvp_ob.tdata [5], \tlvp_ob.tdata [4], \tlvp_ob.tdata [3], 
	\tlvp_ob.tdata [2], \tlvp_ob.tdata [1], \tlvp_ob.tdata [0]} ), 
	tlvp_rsm_bimc_odat, tlvp_rsm_bimc_osync, 
	tlvp_ob_ro_uncorrectable_ecc_error, 
	usr_ob_ro_uncorrectable_ecc_error, clk, rst_n, pt_ob_empty, 
	pt_ob_aempty, .pt_ob_tlv( {\pt_ob_tlv.insert , 
	\pt_ob_tlv.ordern [12], \pt_ob_tlv.ordern [11], 
	\pt_ob_tlv.ordern [10], \pt_ob_tlv.ordern [9], \pt_ob_tlv.ordern [8], 
	\pt_ob_tlv.ordern [7], \pt_ob_tlv.ordern [6], \pt_ob_tlv.ordern [5], 
	\pt_ob_tlv.ordern [4], \pt_ob_tlv.ordern [3], \pt_ob_tlv.ordern [2], 
	\pt_ob_tlv.ordern [1], \pt_ob_tlv.ordern [0], \pt_ob_tlv.typen [7], 
	\pt_ob_tlv.typen [6], \pt_ob_tlv.typen [5], \pt_ob_tlv.typen [4], 
	\pt_ob_tlv.typen [3], \pt_ob_tlv.typen [2], \pt_ob_tlv.typen [1], 
	\pt_ob_tlv.typen [0], \pt_ob_tlv.sot , \pt_ob_tlv.eot , 
	\pt_ob_tlv.tlast , \pt_ob_tlv.tid [0], \pt_ob_tlv.tstrb [7], 
	\pt_ob_tlv.tstrb [6], \pt_ob_tlv.tstrb [5], \pt_ob_tlv.tstrb [4], 
	\pt_ob_tlv.tstrb [3], \pt_ob_tlv.tstrb [2], \pt_ob_tlv.tstrb [1], 
	\pt_ob_tlv.tstrb [0], \pt_ob_tlv.tuser [7], \pt_ob_tlv.tuser [6], 
	\pt_ob_tlv.tuser [5], \pt_ob_tlv.tuser [4], \pt_ob_tlv.tuser [3], 
	\pt_ob_tlv.tuser [2], \pt_ob_tlv.tuser [1], \pt_ob_tlv.tuser [0], 
	\pt_ob_tlv.tdata [63], \pt_ob_tlv.tdata [62], \pt_ob_tlv.tdata [61], 
	\pt_ob_tlv.tdata [60], \pt_ob_tlv.tdata [59], \pt_ob_tlv.tdata [58], 
	\pt_ob_tlv.tdata [57], \pt_ob_tlv.tdata [56], \pt_ob_tlv.tdata [55], 
	\pt_ob_tlv.tdata [54], \pt_ob_tlv.tdata [53], \pt_ob_tlv.tdata [52], 
	\pt_ob_tlv.tdata [51], \pt_ob_tlv.tdata [50], \pt_ob_tlv.tdata [49], 
	\pt_ob_tlv.tdata [48], \pt_ob_tlv.tdata [47], \pt_ob_tlv.tdata [46], 
	\pt_ob_tlv.tdata [45], \pt_ob_tlv.tdata [44], \pt_ob_tlv.tdata [43], 
	\pt_ob_tlv.tdata [42], \pt_ob_tlv.tdata [41], \pt_ob_tlv.tdata [40], 
	\pt_ob_tlv.tdata [39], \pt_ob_tlv.tdata [38], \pt_ob_tlv.tdata [37], 
	\pt_ob_tlv.tdata [36], \pt_ob_tlv.tdata [35], \pt_ob_tlv.tdata [34], 
	\pt_ob_tlv.tdata [33], \pt_ob_tlv.tdata [32], \pt_ob_tlv.tdata [31], 
	\pt_ob_tlv.tdata [30], \pt_ob_tlv.tdata [29], \pt_ob_tlv.tdata [28], 
	\pt_ob_tlv.tdata [27], \pt_ob_tlv.tdata [26], \pt_ob_tlv.tdata [25], 
	\pt_ob_tlv.tdata [24], \pt_ob_tlv.tdata [23], \pt_ob_tlv.tdata [22], 
	\pt_ob_tlv.tdata [21], \pt_ob_tlv.tdata [20], \pt_ob_tlv.tdata [19], 
	\pt_ob_tlv.tdata [18], \pt_ob_tlv.tdata [17], \pt_ob_tlv.tdata [16], 
	\pt_ob_tlv.tdata [15], \pt_ob_tlv.tdata [14], \pt_ob_tlv.tdata [13], 
	\pt_ob_tlv.tdata [12], \pt_ob_tlv.tdata [11], \pt_ob_tlv.tdata [10], 
	\pt_ob_tlv.tdata [9], \pt_ob_tlv.tdata [8], \pt_ob_tlv.tdata [7], 
	\pt_ob_tlv.tdata [6], \pt_ob_tlv.tdata [5], \pt_ob_tlv.tdata [4], 
	\pt_ob_tlv.tdata [3], \pt_ob_tlv.tdata [2], \pt_ob_tlv.tdata [1], 
	\pt_ob_tlv.tdata [0]} ), usr_ob_wr, .usr_ob_tlv( {
	\usr_ob_tlv.insert , \usr_ob_tlv.ordern [12], 
	\usr_ob_tlv.ordern [11], \usr_ob_tlv.ordern [10], 
	\usr_ob_tlv.ordern [9], \usr_ob_tlv.ordern [8], 
	\usr_ob_tlv.ordern [7], \usr_ob_tlv.ordern [6], 
	\usr_ob_tlv.ordern [5], \usr_ob_tlv.ordern [4], 
	\usr_ob_tlv.ordern [3], \usr_ob_tlv.ordern [2], 
	\usr_ob_tlv.ordern [1], \usr_ob_tlv.ordern [0], 
	\usr_ob_tlv.typen [7], \usr_ob_tlv.typen [6], \usr_ob_tlv.typen [5], 
	\usr_ob_tlv.typen [4], \usr_ob_tlv.typen [3], \usr_ob_tlv.typen [2], 
	\usr_ob_tlv.typen [1], \usr_ob_tlv.typen [0], \usr_ob_tlv.sot , 
	\usr_ob_tlv.eot , \usr_ob_tlv.tlast , \usr_ob_tlv.tid [0], 
	\usr_ob_tlv.tstrb [7], \usr_ob_tlv.tstrb [6], \usr_ob_tlv.tstrb [5], 
	\usr_ob_tlv.tstrb [4], \usr_ob_tlv.tstrb [3], \usr_ob_tlv.tstrb [2], 
	\usr_ob_tlv.tstrb [1], \usr_ob_tlv.tstrb [0], \usr_ob_tlv.tuser [7], 
	\usr_ob_tlv.tuser [6], \usr_ob_tlv.tuser [5], \usr_ob_tlv.tuser [4], 
	\usr_ob_tlv.tuser [3], \usr_ob_tlv.tuser [2], \usr_ob_tlv.tuser [1], 
	\usr_ob_tlv.tuser [0], \usr_ob_tlv.tdata [63], 
	\usr_ob_tlv.tdata [62], \usr_ob_tlv.tdata [61], 
	\usr_ob_tlv.tdata [60], \usr_ob_tlv.tdata [59], 
	\usr_ob_tlv.tdata [58], \usr_ob_tlv.tdata [57], 
	\usr_ob_tlv.tdata [56], \usr_ob_tlv.tdata [55], 
	\usr_ob_tlv.tdata [54], \usr_ob_tlv.tdata [53], 
	\usr_ob_tlv.tdata [52], \usr_ob_tlv.tdata [51], 
	\usr_ob_tlv.tdata [50], \usr_ob_tlv.tdata [49], 
	\usr_ob_tlv.tdata [48], \usr_ob_tlv.tdata [47], 
	\usr_ob_tlv.tdata [46], \usr_ob_tlv.tdata [45], 
	\usr_ob_tlv.tdata [44], \usr_ob_tlv.tdata [43], 
	\usr_ob_tlv.tdata [42], \usr_ob_tlv.tdata [41], 
	\usr_ob_tlv.tdata [40], \usr_ob_tlv.tdata [39], 
	\usr_ob_tlv.tdata [38], \usr_ob_tlv.tdata [37], 
	\usr_ob_tlv.tdata [36], \usr_ob_tlv.tdata [35], 
	\usr_ob_tlv.tdata [34], \usr_ob_tlv.tdata [33], 
	\usr_ob_tlv.tdata [32], \usr_ob_tlv.tdata [31], 
	\usr_ob_tlv.tdata [30], \usr_ob_tlv.tdata [29], 
	\usr_ob_tlv.tdata [28], \usr_ob_tlv.tdata [27], 
	\usr_ob_tlv.tdata [26], \usr_ob_tlv.tdata [25], 
	\usr_ob_tlv.tdata [24], \usr_ob_tlv.tdata [23], 
	\usr_ob_tlv.tdata [22], \usr_ob_tlv.tdata [21], 
	\usr_ob_tlv.tdata [20], \usr_ob_tlv.tdata [19], 
	\usr_ob_tlv.tdata [18], \usr_ob_tlv.tdata [17], 
	\usr_ob_tlv.tdata [16], \usr_ob_tlv.tdata [15], 
	\usr_ob_tlv.tdata [14], \usr_ob_tlv.tdata [13], 
	\usr_ob_tlv.tdata [12], \usr_ob_tlv.tdata [11], 
	\usr_ob_tlv.tdata [10], \usr_ob_tlv.tdata [9], \usr_ob_tlv.tdata [8], 
	\usr_ob_tlv.tdata [7], \usr_ob_tlv.tdata [6], \usr_ob_tlv.tdata [5], 
	\usr_ob_tlv.tdata [4], \usr_ob_tlv.tdata [3], \usr_ob_tlv.tdata [2], 
	\usr_ob_tlv.tdata [1], \usr_ob_tlv.tdata [0]} ), tlvp_ob_rd, 
	tlvp_rsm_bimc_idat, tlvp_rsm_bimc_isync, bimc_rst_n);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output pt_ob_rd;
output usr_ob_full;
output usr_ob_afull;
output tlvp_ob_empty;
output tlvp_ob_aempty;
output \tlvp_ob.tvalid ;
output \tlvp_ob.tlast ;
output [0:0] \tlvp_ob.tid ;
output [7:0] \tlvp_ob.tstrb ;
output [7:0] \tlvp_ob.tuser ;
output [63:0] \tlvp_ob.tdata ;
wire [82:0] tlvp_ob;
output tlvp_rsm_bimc_odat;
output tlvp_rsm_bimc_osync;
output tlvp_ob_ro_uncorrectable_ecc_error;
output usr_ob_ro_uncorrectable_ecc_error;
input clk;
input rst_n;
input pt_ob_empty;
input pt_ob_aempty;
input \pt_ob_tlv.insert ;
input [12:0] \pt_ob_tlv.ordern ;
input [7:0] \pt_ob_tlv.typen ;
input \pt_ob_tlv.sot ;
input \pt_ob_tlv.eot ;
input \pt_ob_tlv.tlast ;
input [0:0] \pt_ob_tlv.tid ;
input [7:0] \pt_ob_tlv.tstrb ;
input [7:0] \pt_ob_tlv.tuser ;
input [63:0] \pt_ob_tlv.tdata ;
wire [105:0] pt_ob_tlv;
input usr_ob_wr;
input \usr_ob_tlv.insert ;
input [12:0] \usr_ob_tlv.ordern ;
input [7:0] \usr_ob_tlv.typen ;
input \usr_ob_tlv.sot ;
input \usr_ob_tlv.eot ;
input \usr_ob_tlv.tlast ;
input [0:0] \usr_ob_tlv.tid ;
input [7:0] \usr_ob_tlv.tstrb ;
input [7:0] \usr_ob_tlv.tuser ;
input [63:0] \usr_ob_tlv.tdata ;
wire [105:0] usr_ob_tlv;
input tlvp_ob_rd;
input tlvp_rsm_bimc_idat;
input tlvp_rsm_bimc_isync;
input bimc_rst_n;
wire _zy_simnet_pt_ob_rd_0_w$;
wire _zy_simnet_usr_ob_full_1_w$;
wire _zy_simnet_usr_ob_afull_2_w$;
wire _zy_simnet_tlvp_ob_empty_3_w$;
wire _zy_simnet_tlvp_ob_aempty_4_w$;
wire [0:82] _zy_simnet_tlvp_ob_5_w$;
wire _zy_simnet_tlvp_rsm_bimc_odat_6_w$;
wire _zy_simnet_tlvp_rsm_bimc_osync_7_w$;
wire _zy_simnet_tlvp_ob_ro_uncorrectable_ecc_error_8_w$;
wire _zy_simnet_usr_ob_ro_uncorrectable_ecc_error_9_w$;
wire _zy_simnet_pt_ob_rd_10_w$;
wire _zy_simnet_tlvp_rsm_usr_ob_ren_11_w$;
wire _zy_simnet_tlvp_rsm_ob_wen_12_w$;
wire [0:82] _zy_simnet_tlvp_rsm_ob_wdata_13_w$;
wire [0:105] _zy_simnet_tlvp_rsm_usr_ob_rdata_14_w$;
wire _zy_simnet_usr_ob_empty_15_w$;
wire _zy_simnet_usr_ob_aempty_16_w$;
wire _zy_simnet_tlvp_ob_full_17_w$;
wire _zy_simnet_tlvp_ob_afull_18_w$;
wire _zy_simnet_tlvp_ob_full_19_w$;
wire _zy_simnet_tlvp_ob_afull_20_w$;
wire [0:82] _zy_simnet_tlvp_ob_21_w$;
wire _zy_simnet_tlvp_ob_empty_22_w$;
wire _zy_simnet_tlvp_ob_aempty_23_w$;
wire _zy_simnet_tlvp_rsm_bimc_odat_24_w$;
wire _zy_simnet_tlvp_rsm_bimc_osync_25_w$;
wire _zy_simnet_tlvp_ob_ro_uncorrectable_ecc_error_26_w$;
wire [0:82] _zy_simnet_tlvp_rsm_ob_wdata_27_w$;
wire _zy_simnet_tlvp_rsm_ob_wen_28_w$;
wire _zy_simnet_usr_ob_bimc_odat_29_w$;
wire _zy_simnet_usr_ob_bimc_osync_30_w$;
wire _zy_simnet_usr_ob_full_31_w$;
wire _zy_simnet_usr_ob_afull_32_w$;
wire [0:105] _zy_simnet_tlvp_rsm_usr_ob_rdata_33_w$;
wire _zy_simnet_usr_ob_empty_34_w$;
wire _zy_simnet_usr_ob_aempty_35_w$;
wire _zy_simnet_usr_ob_bimc_odat_36_w$;
wire _zy_simnet_usr_ob_bimc_osync_37_w$;
wire _zy_simnet_usr_ob_ro_uncorrectable_ecc_error_38_w$;
wire _zy_simnet_tlvp_rsm_usr_ob_ren_39_w$;
wire [105:0] tlvp_rsm_usr_ob_rdata;
wire [82:0] tlvp_rsm_ob_wdata;
wire tlvp_ob_afull;
wire tlvp_ob_full;
wire tlvp_rsm_ob_wen;
wire tlvp_rsm_usr_ob_ren;
wire usr_ob_aempty;
wire usr_ob_bimc_odat;
wire usr_ob_bimc_osync;
wire usr_ob_empty;
wire \tlvp_rsm_usr_ob_rdata.insert ;
wire [12:0] \tlvp_rsm_usr_ob_rdata.ordern ;
wire [7:0] \tlvp_rsm_usr_ob_rdata.typen ;
wire \tlvp_rsm_usr_ob_rdata.sot ;
wire \tlvp_rsm_usr_ob_rdata.eot ;
wire \tlvp_rsm_usr_ob_rdata.tlast ;
wire [0:0] \tlvp_rsm_usr_ob_rdata.tid ;
wire [7:0] \tlvp_rsm_usr_ob_rdata.tstrb ;
wire [7:0] \tlvp_rsm_usr_ob_rdata.tuser ;
wire [63:0] \tlvp_rsm_usr_ob_rdata.tdata ;
wire \tlvp_rsm_ob_wdata.tvalid ;
wire \tlvp_rsm_ob_wdata.tlast ;
wire [0:0] \tlvp_rsm_ob_wdata.tid ;
wire [7:0] \tlvp_rsm_ob_wdata.tstrb ;
wire [7:0] \tlvp_rsm_ob_wdata.tuser ;
wire [63:0] \tlvp_rsm_ob_wdata.tdata ;
tran (tlvp_ob[82], \tlvp_ob.tvalid );
tran (tlvp_ob[81], \tlvp_ob.tlast );
tran (tlvp_ob[80], \tlvp_ob.tid [0]);
tran (tlvp_ob[79], \tlvp_ob.tstrb [7]);
tran (tlvp_ob[78], \tlvp_ob.tstrb [6]);
tran (tlvp_ob[77], \tlvp_ob.tstrb [5]);
tran (tlvp_ob[76], \tlvp_ob.tstrb [4]);
tran (tlvp_ob[75], \tlvp_ob.tstrb [3]);
tran (tlvp_ob[74], \tlvp_ob.tstrb [2]);
tran (tlvp_ob[73], \tlvp_ob.tstrb [1]);
tran (tlvp_ob[72], \tlvp_ob.tstrb [0]);
tran (tlvp_ob[71], \tlvp_ob.tuser [7]);
tran (tlvp_ob[70], \tlvp_ob.tuser [6]);
tran (tlvp_ob[69], \tlvp_ob.tuser [5]);
tran (tlvp_ob[68], \tlvp_ob.tuser [4]);
tran (tlvp_ob[67], \tlvp_ob.tuser [3]);
tran (tlvp_ob[66], \tlvp_ob.tuser [2]);
tran (tlvp_ob[65], \tlvp_ob.tuser [1]);
tran (tlvp_ob[64], \tlvp_ob.tuser [0]);
tran (tlvp_ob[63], \tlvp_ob.tdata [63]);
tran (tlvp_ob[62], \tlvp_ob.tdata [62]);
tran (tlvp_ob[61], \tlvp_ob.tdata [61]);
tran (tlvp_ob[60], \tlvp_ob.tdata [60]);
tran (tlvp_ob[59], \tlvp_ob.tdata [59]);
tran (tlvp_ob[58], \tlvp_ob.tdata [58]);
tran (tlvp_ob[57], \tlvp_ob.tdata [57]);
tran (tlvp_ob[56], \tlvp_ob.tdata [56]);
tran (tlvp_ob[55], \tlvp_ob.tdata [55]);
tran (tlvp_ob[54], \tlvp_ob.tdata [54]);
tran (tlvp_ob[53], \tlvp_ob.tdata [53]);
tran (tlvp_ob[52], \tlvp_ob.tdata [52]);
tran (tlvp_ob[51], \tlvp_ob.tdata [51]);
tran (tlvp_ob[50], \tlvp_ob.tdata [50]);
tran (tlvp_ob[49], \tlvp_ob.tdata [49]);
tran (tlvp_ob[48], \tlvp_ob.tdata [48]);
tran (tlvp_ob[47], \tlvp_ob.tdata [47]);
tran (tlvp_ob[46], \tlvp_ob.tdata [46]);
tran (tlvp_ob[45], \tlvp_ob.tdata [45]);
tran (tlvp_ob[44], \tlvp_ob.tdata [44]);
tran (tlvp_ob[43], \tlvp_ob.tdata [43]);
tran (tlvp_ob[42], \tlvp_ob.tdata [42]);
tran (tlvp_ob[41], \tlvp_ob.tdata [41]);
tran (tlvp_ob[40], \tlvp_ob.tdata [40]);
tran (tlvp_ob[39], \tlvp_ob.tdata [39]);
tran (tlvp_ob[38], \tlvp_ob.tdata [38]);
tran (tlvp_ob[37], \tlvp_ob.tdata [37]);
tran (tlvp_ob[36], \tlvp_ob.tdata [36]);
tran (tlvp_ob[35], \tlvp_ob.tdata [35]);
tran (tlvp_ob[34], \tlvp_ob.tdata [34]);
tran (tlvp_ob[33], \tlvp_ob.tdata [33]);
tran (tlvp_ob[32], \tlvp_ob.tdata [32]);
tran (tlvp_ob[31], \tlvp_ob.tdata [31]);
tran (tlvp_ob[30], \tlvp_ob.tdata [30]);
tran (tlvp_ob[29], \tlvp_ob.tdata [29]);
tran (tlvp_ob[28], \tlvp_ob.tdata [28]);
tran (tlvp_ob[27], \tlvp_ob.tdata [27]);
tran (tlvp_ob[26], \tlvp_ob.tdata [26]);
tran (tlvp_ob[25], \tlvp_ob.tdata [25]);
tran (tlvp_ob[24], \tlvp_ob.tdata [24]);
tran (tlvp_ob[23], \tlvp_ob.tdata [23]);
tran (tlvp_ob[22], \tlvp_ob.tdata [22]);
tran (tlvp_ob[21], \tlvp_ob.tdata [21]);
tran (tlvp_ob[20], \tlvp_ob.tdata [20]);
tran (tlvp_ob[19], \tlvp_ob.tdata [19]);
tran (tlvp_ob[18], \tlvp_ob.tdata [18]);
tran (tlvp_ob[17], \tlvp_ob.tdata [17]);
tran (tlvp_ob[16], \tlvp_ob.tdata [16]);
tran (tlvp_ob[15], \tlvp_ob.tdata [15]);
tran (tlvp_ob[14], \tlvp_ob.tdata [14]);
tran (tlvp_ob[13], \tlvp_ob.tdata [13]);
tran (tlvp_ob[12], \tlvp_ob.tdata [12]);
tran (tlvp_ob[11], \tlvp_ob.tdata [11]);
tran (tlvp_ob[10], \tlvp_ob.tdata [10]);
tran (tlvp_ob[9], \tlvp_ob.tdata [9]);
tran (tlvp_ob[8], \tlvp_ob.tdata [8]);
tran (tlvp_ob[7], \tlvp_ob.tdata [7]);
tran (tlvp_ob[6], \tlvp_ob.tdata [6]);
tran (tlvp_ob[5], \tlvp_ob.tdata [5]);
tran (tlvp_ob[4], \tlvp_ob.tdata [4]);
tran (tlvp_ob[3], \tlvp_ob.tdata [3]);
tran (tlvp_ob[2], \tlvp_ob.tdata [2]);
tran (tlvp_ob[1], \tlvp_ob.tdata [1]);
tran (tlvp_ob[0], \tlvp_ob.tdata [0]);
tran (pt_ob_tlv[105], \pt_ob_tlv.insert );
tran (pt_ob_tlv[104], \pt_ob_tlv.ordern [12]);
tran (pt_ob_tlv[103], \pt_ob_tlv.ordern [11]);
tran (pt_ob_tlv[102], \pt_ob_tlv.ordern [10]);
tran (pt_ob_tlv[101], \pt_ob_tlv.ordern [9]);
tran (pt_ob_tlv[100], \pt_ob_tlv.ordern [8]);
tran (pt_ob_tlv[99], \pt_ob_tlv.ordern [7]);
tran (pt_ob_tlv[98], \pt_ob_tlv.ordern [6]);
tran (pt_ob_tlv[97], \pt_ob_tlv.ordern [5]);
tran (pt_ob_tlv[96], \pt_ob_tlv.ordern [4]);
tran (pt_ob_tlv[95], \pt_ob_tlv.ordern [3]);
tran (pt_ob_tlv[94], \pt_ob_tlv.ordern [2]);
tran (pt_ob_tlv[93], \pt_ob_tlv.ordern [1]);
tran (pt_ob_tlv[92], \pt_ob_tlv.ordern [0]);
tran (pt_ob_tlv[91], \pt_ob_tlv.typen [7]);
tran (pt_ob_tlv[90], \pt_ob_tlv.typen [6]);
tran (pt_ob_tlv[89], \pt_ob_tlv.typen [5]);
tran (pt_ob_tlv[88], \pt_ob_tlv.typen [4]);
tran (pt_ob_tlv[87], \pt_ob_tlv.typen [3]);
tran (pt_ob_tlv[86], \pt_ob_tlv.typen [2]);
tran (pt_ob_tlv[85], \pt_ob_tlv.typen [1]);
tran (pt_ob_tlv[84], \pt_ob_tlv.typen [0]);
tran (pt_ob_tlv[83], \pt_ob_tlv.sot );
tran (pt_ob_tlv[82], \pt_ob_tlv.eot );
tran (pt_ob_tlv[81], \pt_ob_tlv.tlast );
tran (pt_ob_tlv[80], \pt_ob_tlv.tid [0]);
tran (pt_ob_tlv[79], \pt_ob_tlv.tstrb [7]);
tran (pt_ob_tlv[78], \pt_ob_tlv.tstrb [6]);
tran (pt_ob_tlv[77], \pt_ob_tlv.tstrb [5]);
tran (pt_ob_tlv[76], \pt_ob_tlv.tstrb [4]);
tran (pt_ob_tlv[75], \pt_ob_tlv.tstrb [3]);
tran (pt_ob_tlv[74], \pt_ob_tlv.tstrb [2]);
tran (pt_ob_tlv[73], \pt_ob_tlv.tstrb [1]);
tran (pt_ob_tlv[72], \pt_ob_tlv.tstrb [0]);
tran (pt_ob_tlv[71], \pt_ob_tlv.tuser [7]);
tran (pt_ob_tlv[70], \pt_ob_tlv.tuser [6]);
tran (pt_ob_tlv[69], \pt_ob_tlv.tuser [5]);
tran (pt_ob_tlv[68], \pt_ob_tlv.tuser [4]);
tran (pt_ob_tlv[67], \pt_ob_tlv.tuser [3]);
tran (pt_ob_tlv[66], \pt_ob_tlv.tuser [2]);
tran (pt_ob_tlv[65], \pt_ob_tlv.tuser [1]);
tran (pt_ob_tlv[64], \pt_ob_tlv.tuser [0]);
tran (pt_ob_tlv[63], \pt_ob_tlv.tdata [63]);
tran (pt_ob_tlv[62], \pt_ob_tlv.tdata [62]);
tran (pt_ob_tlv[61], \pt_ob_tlv.tdata [61]);
tran (pt_ob_tlv[60], \pt_ob_tlv.tdata [60]);
tran (pt_ob_tlv[59], \pt_ob_tlv.tdata [59]);
tran (pt_ob_tlv[58], \pt_ob_tlv.tdata [58]);
tran (pt_ob_tlv[57], \pt_ob_tlv.tdata [57]);
tran (pt_ob_tlv[56], \pt_ob_tlv.tdata [56]);
tran (pt_ob_tlv[55], \pt_ob_tlv.tdata [55]);
tran (pt_ob_tlv[54], \pt_ob_tlv.tdata [54]);
tran (pt_ob_tlv[53], \pt_ob_tlv.tdata [53]);
tran (pt_ob_tlv[52], \pt_ob_tlv.tdata [52]);
tran (pt_ob_tlv[51], \pt_ob_tlv.tdata [51]);
tran (pt_ob_tlv[50], \pt_ob_tlv.tdata [50]);
tran (pt_ob_tlv[49], \pt_ob_tlv.tdata [49]);
tran (pt_ob_tlv[48], \pt_ob_tlv.tdata [48]);
tran (pt_ob_tlv[47], \pt_ob_tlv.tdata [47]);
tran (pt_ob_tlv[46], \pt_ob_tlv.tdata [46]);
tran (pt_ob_tlv[45], \pt_ob_tlv.tdata [45]);
tran (pt_ob_tlv[44], \pt_ob_tlv.tdata [44]);
tran (pt_ob_tlv[43], \pt_ob_tlv.tdata [43]);
tran (pt_ob_tlv[42], \pt_ob_tlv.tdata [42]);
tran (pt_ob_tlv[41], \pt_ob_tlv.tdata [41]);
tran (pt_ob_tlv[40], \pt_ob_tlv.tdata [40]);
tran (pt_ob_tlv[39], \pt_ob_tlv.tdata [39]);
tran (pt_ob_tlv[38], \pt_ob_tlv.tdata [38]);
tran (pt_ob_tlv[37], \pt_ob_tlv.tdata [37]);
tran (pt_ob_tlv[36], \pt_ob_tlv.tdata [36]);
tran (pt_ob_tlv[35], \pt_ob_tlv.tdata [35]);
tran (pt_ob_tlv[34], \pt_ob_tlv.tdata [34]);
tran (pt_ob_tlv[33], \pt_ob_tlv.tdata [33]);
tran (pt_ob_tlv[32], \pt_ob_tlv.tdata [32]);
tran (pt_ob_tlv[31], \pt_ob_tlv.tdata [31]);
tran (pt_ob_tlv[30], \pt_ob_tlv.tdata [30]);
tran (pt_ob_tlv[29], \pt_ob_tlv.tdata [29]);
tran (pt_ob_tlv[28], \pt_ob_tlv.tdata [28]);
tran (pt_ob_tlv[27], \pt_ob_tlv.tdata [27]);
tran (pt_ob_tlv[26], \pt_ob_tlv.tdata [26]);
tran (pt_ob_tlv[25], \pt_ob_tlv.tdata [25]);
tran (pt_ob_tlv[24], \pt_ob_tlv.tdata [24]);
tran (pt_ob_tlv[23], \pt_ob_tlv.tdata [23]);
tran (pt_ob_tlv[22], \pt_ob_tlv.tdata [22]);
tran (pt_ob_tlv[21], \pt_ob_tlv.tdata [21]);
tran (pt_ob_tlv[20], \pt_ob_tlv.tdata [20]);
tran (pt_ob_tlv[19], \pt_ob_tlv.tdata [19]);
tran (pt_ob_tlv[18], \pt_ob_tlv.tdata [18]);
tran (pt_ob_tlv[17], \pt_ob_tlv.tdata [17]);
tran (pt_ob_tlv[16], \pt_ob_tlv.tdata [16]);
tran (pt_ob_tlv[15], \pt_ob_tlv.tdata [15]);
tran (pt_ob_tlv[14], \pt_ob_tlv.tdata [14]);
tran (pt_ob_tlv[13], \pt_ob_tlv.tdata [13]);
tran (pt_ob_tlv[12], \pt_ob_tlv.tdata [12]);
tran (pt_ob_tlv[11], \pt_ob_tlv.tdata [11]);
tran (pt_ob_tlv[10], \pt_ob_tlv.tdata [10]);
tran (pt_ob_tlv[9], \pt_ob_tlv.tdata [9]);
tran (pt_ob_tlv[8], \pt_ob_tlv.tdata [8]);
tran (pt_ob_tlv[7], \pt_ob_tlv.tdata [7]);
tran (pt_ob_tlv[6], \pt_ob_tlv.tdata [6]);
tran (pt_ob_tlv[5], \pt_ob_tlv.tdata [5]);
tran (pt_ob_tlv[4], \pt_ob_tlv.tdata [4]);
tran (pt_ob_tlv[3], \pt_ob_tlv.tdata [3]);
tran (pt_ob_tlv[2], \pt_ob_tlv.tdata [2]);
tran (pt_ob_tlv[1], \pt_ob_tlv.tdata [1]);
tran (pt_ob_tlv[0], \pt_ob_tlv.tdata [0]);
tran (usr_ob_tlv[105], \usr_ob_tlv.insert );
tran (usr_ob_tlv[104], \usr_ob_tlv.ordern [12]);
tran (usr_ob_tlv[103], \usr_ob_tlv.ordern [11]);
tran (usr_ob_tlv[102], \usr_ob_tlv.ordern [10]);
tran (usr_ob_tlv[101], \usr_ob_tlv.ordern [9]);
tran (usr_ob_tlv[100], \usr_ob_tlv.ordern [8]);
tran (usr_ob_tlv[99], \usr_ob_tlv.ordern [7]);
tran (usr_ob_tlv[98], \usr_ob_tlv.ordern [6]);
tran (usr_ob_tlv[97], \usr_ob_tlv.ordern [5]);
tran (usr_ob_tlv[96], \usr_ob_tlv.ordern [4]);
tran (usr_ob_tlv[95], \usr_ob_tlv.ordern [3]);
tran (usr_ob_tlv[94], \usr_ob_tlv.ordern [2]);
tran (usr_ob_tlv[93], \usr_ob_tlv.ordern [1]);
tran (usr_ob_tlv[92], \usr_ob_tlv.ordern [0]);
tran (usr_ob_tlv[91], \usr_ob_tlv.typen [7]);
tran (usr_ob_tlv[90], \usr_ob_tlv.typen [6]);
tran (usr_ob_tlv[89], \usr_ob_tlv.typen [5]);
tran (usr_ob_tlv[88], \usr_ob_tlv.typen [4]);
tran (usr_ob_tlv[87], \usr_ob_tlv.typen [3]);
tran (usr_ob_tlv[86], \usr_ob_tlv.typen [2]);
tran (usr_ob_tlv[85], \usr_ob_tlv.typen [1]);
tran (usr_ob_tlv[84], \usr_ob_tlv.typen [0]);
tran (usr_ob_tlv[83], \usr_ob_tlv.sot );
tran (usr_ob_tlv[82], \usr_ob_tlv.eot );
tran (usr_ob_tlv[81], \usr_ob_tlv.tlast );
tran (usr_ob_tlv[80], \usr_ob_tlv.tid [0]);
tran (usr_ob_tlv[79], \usr_ob_tlv.tstrb [7]);
tran (usr_ob_tlv[78], \usr_ob_tlv.tstrb [6]);
tran (usr_ob_tlv[77], \usr_ob_tlv.tstrb [5]);
tran (usr_ob_tlv[76], \usr_ob_tlv.tstrb [4]);
tran (usr_ob_tlv[75], \usr_ob_tlv.tstrb [3]);
tran (usr_ob_tlv[74], \usr_ob_tlv.tstrb [2]);
tran (usr_ob_tlv[73], \usr_ob_tlv.tstrb [1]);
tran (usr_ob_tlv[72], \usr_ob_tlv.tstrb [0]);
tran (usr_ob_tlv[71], \usr_ob_tlv.tuser [7]);
tran (usr_ob_tlv[70], \usr_ob_tlv.tuser [6]);
tran (usr_ob_tlv[69], \usr_ob_tlv.tuser [5]);
tran (usr_ob_tlv[68], \usr_ob_tlv.tuser [4]);
tran (usr_ob_tlv[67], \usr_ob_tlv.tuser [3]);
tran (usr_ob_tlv[66], \usr_ob_tlv.tuser [2]);
tran (usr_ob_tlv[65], \usr_ob_tlv.tuser [1]);
tran (usr_ob_tlv[64], \usr_ob_tlv.tuser [0]);
tran (usr_ob_tlv[63], \usr_ob_tlv.tdata [63]);
tran (usr_ob_tlv[62], \usr_ob_tlv.tdata [62]);
tran (usr_ob_tlv[61], \usr_ob_tlv.tdata [61]);
tran (usr_ob_tlv[60], \usr_ob_tlv.tdata [60]);
tran (usr_ob_tlv[59], \usr_ob_tlv.tdata [59]);
tran (usr_ob_tlv[58], \usr_ob_tlv.tdata [58]);
tran (usr_ob_tlv[57], \usr_ob_tlv.tdata [57]);
tran (usr_ob_tlv[56], \usr_ob_tlv.tdata [56]);
tran (usr_ob_tlv[55], \usr_ob_tlv.tdata [55]);
tran (usr_ob_tlv[54], \usr_ob_tlv.tdata [54]);
tran (usr_ob_tlv[53], \usr_ob_tlv.tdata [53]);
tran (usr_ob_tlv[52], \usr_ob_tlv.tdata [52]);
tran (usr_ob_tlv[51], \usr_ob_tlv.tdata [51]);
tran (usr_ob_tlv[50], \usr_ob_tlv.tdata [50]);
tran (usr_ob_tlv[49], \usr_ob_tlv.tdata [49]);
tran (usr_ob_tlv[48], \usr_ob_tlv.tdata [48]);
tran (usr_ob_tlv[47], \usr_ob_tlv.tdata [47]);
tran (usr_ob_tlv[46], \usr_ob_tlv.tdata [46]);
tran (usr_ob_tlv[45], \usr_ob_tlv.tdata [45]);
tran (usr_ob_tlv[44], \usr_ob_tlv.tdata [44]);
tran (usr_ob_tlv[43], \usr_ob_tlv.tdata [43]);
tran (usr_ob_tlv[42], \usr_ob_tlv.tdata [42]);
tran (usr_ob_tlv[41], \usr_ob_tlv.tdata [41]);
tran (usr_ob_tlv[40], \usr_ob_tlv.tdata [40]);
tran (usr_ob_tlv[39], \usr_ob_tlv.tdata [39]);
tran (usr_ob_tlv[38], \usr_ob_tlv.tdata [38]);
tran (usr_ob_tlv[37], \usr_ob_tlv.tdata [37]);
tran (usr_ob_tlv[36], \usr_ob_tlv.tdata [36]);
tran (usr_ob_tlv[35], \usr_ob_tlv.tdata [35]);
tran (usr_ob_tlv[34], \usr_ob_tlv.tdata [34]);
tran (usr_ob_tlv[33], \usr_ob_tlv.tdata [33]);
tran (usr_ob_tlv[32], \usr_ob_tlv.tdata [32]);
tran (usr_ob_tlv[31], \usr_ob_tlv.tdata [31]);
tran (usr_ob_tlv[30], \usr_ob_tlv.tdata [30]);
tran (usr_ob_tlv[29], \usr_ob_tlv.tdata [29]);
tran (usr_ob_tlv[28], \usr_ob_tlv.tdata [28]);
tran (usr_ob_tlv[27], \usr_ob_tlv.tdata [27]);
tran (usr_ob_tlv[26], \usr_ob_tlv.tdata [26]);
tran (usr_ob_tlv[25], \usr_ob_tlv.tdata [25]);
tran (usr_ob_tlv[24], \usr_ob_tlv.tdata [24]);
tran (usr_ob_tlv[23], \usr_ob_tlv.tdata [23]);
tran (usr_ob_tlv[22], \usr_ob_tlv.tdata [22]);
tran (usr_ob_tlv[21], \usr_ob_tlv.tdata [21]);
tran (usr_ob_tlv[20], \usr_ob_tlv.tdata [20]);
tran (usr_ob_tlv[19], \usr_ob_tlv.tdata [19]);
tran (usr_ob_tlv[18], \usr_ob_tlv.tdata [18]);
tran (usr_ob_tlv[17], \usr_ob_tlv.tdata [17]);
tran (usr_ob_tlv[16], \usr_ob_tlv.tdata [16]);
tran (usr_ob_tlv[15], \usr_ob_tlv.tdata [15]);
tran (usr_ob_tlv[14], \usr_ob_tlv.tdata [14]);
tran (usr_ob_tlv[13], \usr_ob_tlv.tdata [13]);
tran (usr_ob_tlv[12], \usr_ob_tlv.tdata [12]);
tran (usr_ob_tlv[11], \usr_ob_tlv.tdata [11]);
tran (usr_ob_tlv[10], \usr_ob_tlv.tdata [10]);
tran (usr_ob_tlv[9], \usr_ob_tlv.tdata [9]);
tran (usr_ob_tlv[8], \usr_ob_tlv.tdata [8]);
tran (usr_ob_tlv[7], \usr_ob_tlv.tdata [7]);
tran (usr_ob_tlv[6], \usr_ob_tlv.tdata [6]);
tran (usr_ob_tlv[5], \usr_ob_tlv.tdata [5]);
tran (usr_ob_tlv[4], \usr_ob_tlv.tdata [4]);
tran (usr_ob_tlv[3], \usr_ob_tlv.tdata [3]);
tran (usr_ob_tlv[2], \usr_ob_tlv.tdata [2]);
tran (usr_ob_tlv[1], \usr_ob_tlv.tdata [1]);
tran (usr_ob_tlv[0], \usr_ob_tlv.tdata [0]);
tran (tlvp_rsm_ob_wdata[82], \tlvp_rsm_ob_wdata.tvalid );
tran (tlvp_rsm_ob_wdata[81], \tlvp_rsm_ob_wdata.tlast );
tran (tlvp_rsm_ob_wdata[80], \tlvp_rsm_ob_wdata.tid [0]);
tran (tlvp_rsm_ob_wdata[79], \tlvp_rsm_ob_wdata.tstrb [7]);
tran (tlvp_rsm_ob_wdata[78], \tlvp_rsm_ob_wdata.tstrb [6]);
tran (tlvp_rsm_ob_wdata[77], \tlvp_rsm_ob_wdata.tstrb [5]);
tran (tlvp_rsm_ob_wdata[76], \tlvp_rsm_ob_wdata.tstrb [4]);
tran (tlvp_rsm_ob_wdata[75], \tlvp_rsm_ob_wdata.tstrb [3]);
tran (tlvp_rsm_ob_wdata[74], \tlvp_rsm_ob_wdata.tstrb [2]);
tran (tlvp_rsm_ob_wdata[73], \tlvp_rsm_ob_wdata.tstrb [1]);
tran (tlvp_rsm_ob_wdata[72], \tlvp_rsm_ob_wdata.tstrb [0]);
tran (tlvp_rsm_ob_wdata[71], \tlvp_rsm_ob_wdata.tuser [7]);
tran (tlvp_rsm_ob_wdata[70], \tlvp_rsm_ob_wdata.tuser [6]);
tran (tlvp_rsm_ob_wdata[69], \tlvp_rsm_ob_wdata.tuser [5]);
tran (tlvp_rsm_ob_wdata[68], \tlvp_rsm_ob_wdata.tuser [4]);
tran (tlvp_rsm_ob_wdata[67], \tlvp_rsm_ob_wdata.tuser [3]);
tran (tlvp_rsm_ob_wdata[66], \tlvp_rsm_ob_wdata.tuser [2]);
tran (tlvp_rsm_ob_wdata[65], \tlvp_rsm_ob_wdata.tuser [1]);
tran (tlvp_rsm_ob_wdata[64], \tlvp_rsm_ob_wdata.tuser [0]);
tran (tlvp_rsm_ob_wdata[63], \tlvp_rsm_ob_wdata.tdata [63]);
tran (tlvp_rsm_ob_wdata[62], \tlvp_rsm_ob_wdata.tdata [62]);
tran (tlvp_rsm_ob_wdata[61], \tlvp_rsm_ob_wdata.tdata [61]);
tran (tlvp_rsm_ob_wdata[60], \tlvp_rsm_ob_wdata.tdata [60]);
tran (tlvp_rsm_ob_wdata[59], \tlvp_rsm_ob_wdata.tdata [59]);
tran (tlvp_rsm_ob_wdata[58], \tlvp_rsm_ob_wdata.tdata [58]);
tran (tlvp_rsm_ob_wdata[57], \tlvp_rsm_ob_wdata.tdata [57]);
tran (tlvp_rsm_ob_wdata[56], \tlvp_rsm_ob_wdata.tdata [56]);
tran (tlvp_rsm_ob_wdata[55], \tlvp_rsm_ob_wdata.tdata [55]);
tran (tlvp_rsm_ob_wdata[54], \tlvp_rsm_ob_wdata.tdata [54]);
tran (tlvp_rsm_ob_wdata[53], \tlvp_rsm_ob_wdata.tdata [53]);
tran (tlvp_rsm_ob_wdata[52], \tlvp_rsm_ob_wdata.tdata [52]);
tran (tlvp_rsm_ob_wdata[51], \tlvp_rsm_ob_wdata.tdata [51]);
tran (tlvp_rsm_ob_wdata[50], \tlvp_rsm_ob_wdata.tdata [50]);
tran (tlvp_rsm_ob_wdata[49], \tlvp_rsm_ob_wdata.tdata [49]);
tran (tlvp_rsm_ob_wdata[48], \tlvp_rsm_ob_wdata.tdata [48]);
tran (tlvp_rsm_ob_wdata[47], \tlvp_rsm_ob_wdata.tdata [47]);
tran (tlvp_rsm_ob_wdata[46], \tlvp_rsm_ob_wdata.tdata [46]);
tran (tlvp_rsm_ob_wdata[45], \tlvp_rsm_ob_wdata.tdata [45]);
tran (tlvp_rsm_ob_wdata[44], \tlvp_rsm_ob_wdata.tdata [44]);
tran (tlvp_rsm_ob_wdata[43], \tlvp_rsm_ob_wdata.tdata [43]);
tran (tlvp_rsm_ob_wdata[42], \tlvp_rsm_ob_wdata.tdata [42]);
tran (tlvp_rsm_ob_wdata[41], \tlvp_rsm_ob_wdata.tdata [41]);
tran (tlvp_rsm_ob_wdata[40], \tlvp_rsm_ob_wdata.tdata [40]);
tran (tlvp_rsm_ob_wdata[39], \tlvp_rsm_ob_wdata.tdata [39]);
tran (tlvp_rsm_ob_wdata[38], \tlvp_rsm_ob_wdata.tdata [38]);
tran (tlvp_rsm_ob_wdata[37], \tlvp_rsm_ob_wdata.tdata [37]);
tran (tlvp_rsm_ob_wdata[36], \tlvp_rsm_ob_wdata.tdata [36]);
tran (tlvp_rsm_ob_wdata[35], \tlvp_rsm_ob_wdata.tdata [35]);
tran (tlvp_rsm_ob_wdata[34], \tlvp_rsm_ob_wdata.tdata [34]);
tran (tlvp_rsm_ob_wdata[33], \tlvp_rsm_ob_wdata.tdata [33]);
tran (tlvp_rsm_ob_wdata[32], \tlvp_rsm_ob_wdata.tdata [32]);
tran (tlvp_rsm_ob_wdata[31], \tlvp_rsm_ob_wdata.tdata [31]);
tran (tlvp_rsm_ob_wdata[30], \tlvp_rsm_ob_wdata.tdata [30]);
tran (tlvp_rsm_ob_wdata[29], \tlvp_rsm_ob_wdata.tdata [29]);
tran (tlvp_rsm_ob_wdata[28], \tlvp_rsm_ob_wdata.tdata [28]);
tran (tlvp_rsm_ob_wdata[27], \tlvp_rsm_ob_wdata.tdata [27]);
tran (tlvp_rsm_ob_wdata[26], \tlvp_rsm_ob_wdata.tdata [26]);
tran (tlvp_rsm_ob_wdata[25], \tlvp_rsm_ob_wdata.tdata [25]);
tran (tlvp_rsm_ob_wdata[24], \tlvp_rsm_ob_wdata.tdata [24]);
tran (tlvp_rsm_ob_wdata[23], \tlvp_rsm_ob_wdata.tdata [23]);
tran (tlvp_rsm_ob_wdata[22], \tlvp_rsm_ob_wdata.tdata [22]);
tran (tlvp_rsm_ob_wdata[21], \tlvp_rsm_ob_wdata.tdata [21]);
tran (tlvp_rsm_ob_wdata[20], \tlvp_rsm_ob_wdata.tdata [20]);
tran (tlvp_rsm_ob_wdata[19], \tlvp_rsm_ob_wdata.tdata [19]);
tran (tlvp_rsm_ob_wdata[18], \tlvp_rsm_ob_wdata.tdata [18]);
tran (tlvp_rsm_ob_wdata[17], \tlvp_rsm_ob_wdata.tdata [17]);
tran (tlvp_rsm_ob_wdata[16], \tlvp_rsm_ob_wdata.tdata [16]);
tran (tlvp_rsm_ob_wdata[15], \tlvp_rsm_ob_wdata.tdata [15]);
tran (tlvp_rsm_ob_wdata[14], \tlvp_rsm_ob_wdata.tdata [14]);
tran (tlvp_rsm_ob_wdata[13], \tlvp_rsm_ob_wdata.tdata [13]);
tran (tlvp_rsm_ob_wdata[12], \tlvp_rsm_ob_wdata.tdata [12]);
tran (tlvp_rsm_ob_wdata[11], \tlvp_rsm_ob_wdata.tdata [11]);
tran (tlvp_rsm_ob_wdata[10], \tlvp_rsm_ob_wdata.tdata [10]);
tran (tlvp_rsm_ob_wdata[9], \tlvp_rsm_ob_wdata.tdata [9]);
tran (tlvp_rsm_ob_wdata[8], \tlvp_rsm_ob_wdata.tdata [8]);
tran (tlvp_rsm_ob_wdata[7], \tlvp_rsm_ob_wdata.tdata [7]);
tran (tlvp_rsm_ob_wdata[6], \tlvp_rsm_ob_wdata.tdata [6]);
tran (tlvp_rsm_ob_wdata[5], \tlvp_rsm_ob_wdata.tdata [5]);
tran (tlvp_rsm_ob_wdata[4], \tlvp_rsm_ob_wdata.tdata [4]);
tran (tlvp_rsm_ob_wdata[3], \tlvp_rsm_ob_wdata.tdata [3]);
tran (tlvp_rsm_ob_wdata[2], \tlvp_rsm_ob_wdata.tdata [2]);
tran (tlvp_rsm_ob_wdata[1], \tlvp_rsm_ob_wdata.tdata [1]);
tran (tlvp_rsm_ob_wdata[0], \tlvp_rsm_ob_wdata.tdata [0]);
tran (tlvp_rsm_usr_ob_rdata[105], \tlvp_rsm_usr_ob_rdata.insert );
tran (tlvp_rsm_usr_ob_rdata[104], \tlvp_rsm_usr_ob_rdata.ordern [12]);
tran (tlvp_rsm_usr_ob_rdata[103], \tlvp_rsm_usr_ob_rdata.ordern [11]);
tran (tlvp_rsm_usr_ob_rdata[102], \tlvp_rsm_usr_ob_rdata.ordern [10]);
tran (tlvp_rsm_usr_ob_rdata[101], \tlvp_rsm_usr_ob_rdata.ordern [9]);
tran (tlvp_rsm_usr_ob_rdata[100], \tlvp_rsm_usr_ob_rdata.ordern [8]);
tran (tlvp_rsm_usr_ob_rdata[99], \tlvp_rsm_usr_ob_rdata.ordern [7]);
tran (tlvp_rsm_usr_ob_rdata[98], \tlvp_rsm_usr_ob_rdata.ordern [6]);
tran (tlvp_rsm_usr_ob_rdata[97], \tlvp_rsm_usr_ob_rdata.ordern [5]);
tran (tlvp_rsm_usr_ob_rdata[96], \tlvp_rsm_usr_ob_rdata.ordern [4]);
tran (tlvp_rsm_usr_ob_rdata[95], \tlvp_rsm_usr_ob_rdata.ordern [3]);
tran (tlvp_rsm_usr_ob_rdata[94], \tlvp_rsm_usr_ob_rdata.ordern [2]);
tran (tlvp_rsm_usr_ob_rdata[93], \tlvp_rsm_usr_ob_rdata.ordern [1]);
tran (tlvp_rsm_usr_ob_rdata[92], \tlvp_rsm_usr_ob_rdata.ordern [0]);
tran (tlvp_rsm_usr_ob_rdata[91], \tlvp_rsm_usr_ob_rdata.typen [7]);
tran (tlvp_rsm_usr_ob_rdata[90], \tlvp_rsm_usr_ob_rdata.typen [6]);
tran (tlvp_rsm_usr_ob_rdata[89], \tlvp_rsm_usr_ob_rdata.typen [5]);
tran (tlvp_rsm_usr_ob_rdata[88], \tlvp_rsm_usr_ob_rdata.typen [4]);
tran (tlvp_rsm_usr_ob_rdata[87], \tlvp_rsm_usr_ob_rdata.typen [3]);
tran (tlvp_rsm_usr_ob_rdata[86], \tlvp_rsm_usr_ob_rdata.typen [2]);
tran (tlvp_rsm_usr_ob_rdata[85], \tlvp_rsm_usr_ob_rdata.typen [1]);
tran (tlvp_rsm_usr_ob_rdata[84], \tlvp_rsm_usr_ob_rdata.typen [0]);
tran (tlvp_rsm_usr_ob_rdata[83], \tlvp_rsm_usr_ob_rdata.sot );
tran (tlvp_rsm_usr_ob_rdata[82], \tlvp_rsm_usr_ob_rdata.eot );
tran (tlvp_rsm_usr_ob_rdata[81], \tlvp_rsm_usr_ob_rdata.tlast );
tran (tlvp_rsm_usr_ob_rdata[80], \tlvp_rsm_usr_ob_rdata.tid [0]);
tran (tlvp_rsm_usr_ob_rdata[79], \tlvp_rsm_usr_ob_rdata.tstrb [7]);
tran (tlvp_rsm_usr_ob_rdata[78], \tlvp_rsm_usr_ob_rdata.tstrb [6]);
tran (tlvp_rsm_usr_ob_rdata[77], \tlvp_rsm_usr_ob_rdata.tstrb [5]);
tran (tlvp_rsm_usr_ob_rdata[76], \tlvp_rsm_usr_ob_rdata.tstrb [4]);
tran (tlvp_rsm_usr_ob_rdata[75], \tlvp_rsm_usr_ob_rdata.tstrb [3]);
tran (tlvp_rsm_usr_ob_rdata[74], \tlvp_rsm_usr_ob_rdata.tstrb [2]);
tran (tlvp_rsm_usr_ob_rdata[73], \tlvp_rsm_usr_ob_rdata.tstrb [1]);
tran (tlvp_rsm_usr_ob_rdata[72], \tlvp_rsm_usr_ob_rdata.tstrb [0]);
tran (tlvp_rsm_usr_ob_rdata[71], \tlvp_rsm_usr_ob_rdata.tuser [7]);
tran (tlvp_rsm_usr_ob_rdata[70], \tlvp_rsm_usr_ob_rdata.tuser [6]);
tran (tlvp_rsm_usr_ob_rdata[69], \tlvp_rsm_usr_ob_rdata.tuser [5]);
tran (tlvp_rsm_usr_ob_rdata[68], \tlvp_rsm_usr_ob_rdata.tuser [4]);
tran (tlvp_rsm_usr_ob_rdata[67], \tlvp_rsm_usr_ob_rdata.tuser [3]);
tran (tlvp_rsm_usr_ob_rdata[66], \tlvp_rsm_usr_ob_rdata.tuser [2]);
tran (tlvp_rsm_usr_ob_rdata[65], \tlvp_rsm_usr_ob_rdata.tuser [1]);
tran (tlvp_rsm_usr_ob_rdata[64], \tlvp_rsm_usr_ob_rdata.tuser [0]);
tran (tlvp_rsm_usr_ob_rdata[63], \tlvp_rsm_usr_ob_rdata.tdata [63]);
tran (tlvp_rsm_usr_ob_rdata[62], \tlvp_rsm_usr_ob_rdata.tdata [62]);
tran (tlvp_rsm_usr_ob_rdata[61], \tlvp_rsm_usr_ob_rdata.tdata [61]);
tran (tlvp_rsm_usr_ob_rdata[60], \tlvp_rsm_usr_ob_rdata.tdata [60]);
tran (tlvp_rsm_usr_ob_rdata[59], \tlvp_rsm_usr_ob_rdata.tdata [59]);
tran (tlvp_rsm_usr_ob_rdata[58], \tlvp_rsm_usr_ob_rdata.tdata [58]);
tran (tlvp_rsm_usr_ob_rdata[57], \tlvp_rsm_usr_ob_rdata.tdata [57]);
tran (tlvp_rsm_usr_ob_rdata[56], \tlvp_rsm_usr_ob_rdata.tdata [56]);
tran (tlvp_rsm_usr_ob_rdata[55], \tlvp_rsm_usr_ob_rdata.tdata [55]);
tran (tlvp_rsm_usr_ob_rdata[54], \tlvp_rsm_usr_ob_rdata.tdata [54]);
tran (tlvp_rsm_usr_ob_rdata[53], \tlvp_rsm_usr_ob_rdata.tdata [53]);
tran (tlvp_rsm_usr_ob_rdata[52], \tlvp_rsm_usr_ob_rdata.tdata [52]);
tran (tlvp_rsm_usr_ob_rdata[51], \tlvp_rsm_usr_ob_rdata.tdata [51]);
tran (tlvp_rsm_usr_ob_rdata[50], \tlvp_rsm_usr_ob_rdata.tdata [50]);
tran (tlvp_rsm_usr_ob_rdata[49], \tlvp_rsm_usr_ob_rdata.tdata [49]);
tran (tlvp_rsm_usr_ob_rdata[48], \tlvp_rsm_usr_ob_rdata.tdata [48]);
tran (tlvp_rsm_usr_ob_rdata[47], \tlvp_rsm_usr_ob_rdata.tdata [47]);
tran (tlvp_rsm_usr_ob_rdata[46], \tlvp_rsm_usr_ob_rdata.tdata [46]);
tran (tlvp_rsm_usr_ob_rdata[45], \tlvp_rsm_usr_ob_rdata.tdata [45]);
tran (tlvp_rsm_usr_ob_rdata[44], \tlvp_rsm_usr_ob_rdata.tdata [44]);
tran (tlvp_rsm_usr_ob_rdata[43], \tlvp_rsm_usr_ob_rdata.tdata [43]);
tran (tlvp_rsm_usr_ob_rdata[42], \tlvp_rsm_usr_ob_rdata.tdata [42]);
tran (tlvp_rsm_usr_ob_rdata[41], \tlvp_rsm_usr_ob_rdata.tdata [41]);
tran (tlvp_rsm_usr_ob_rdata[40], \tlvp_rsm_usr_ob_rdata.tdata [40]);
tran (tlvp_rsm_usr_ob_rdata[39], \tlvp_rsm_usr_ob_rdata.tdata [39]);
tran (tlvp_rsm_usr_ob_rdata[38], \tlvp_rsm_usr_ob_rdata.tdata [38]);
tran (tlvp_rsm_usr_ob_rdata[37], \tlvp_rsm_usr_ob_rdata.tdata [37]);
tran (tlvp_rsm_usr_ob_rdata[36], \tlvp_rsm_usr_ob_rdata.tdata [36]);
tran (tlvp_rsm_usr_ob_rdata[35], \tlvp_rsm_usr_ob_rdata.tdata [35]);
tran (tlvp_rsm_usr_ob_rdata[34], \tlvp_rsm_usr_ob_rdata.tdata [34]);
tran (tlvp_rsm_usr_ob_rdata[33], \tlvp_rsm_usr_ob_rdata.tdata [33]);
tran (tlvp_rsm_usr_ob_rdata[32], \tlvp_rsm_usr_ob_rdata.tdata [32]);
tran (tlvp_rsm_usr_ob_rdata[31], \tlvp_rsm_usr_ob_rdata.tdata [31]);
tran (tlvp_rsm_usr_ob_rdata[30], \tlvp_rsm_usr_ob_rdata.tdata [30]);
tran (tlvp_rsm_usr_ob_rdata[29], \tlvp_rsm_usr_ob_rdata.tdata [29]);
tran (tlvp_rsm_usr_ob_rdata[28], \tlvp_rsm_usr_ob_rdata.tdata [28]);
tran (tlvp_rsm_usr_ob_rdata[27], \tlvp_rsm_usr_ob_rdata.tdata [27]);
tran (tlvp_rsm_usr_ob_rdata[26], \tlvp_rsm_usr_ob_rdata.tdata [26]);
tran (tlvp_rsm_usr_ob_rdata[25], \tlvp_rsm_usr_ob_rdata.tdata [25]);
tran (tlvp_rsm_usr_ob_rdata[24], \tlvp_rsm_usr_ob_rdata.tdata [24]);
tran (tlvp_rsm_usr_ob_rdata[23], \tlvp_rsm_usr_ob_rdata.tdata [23]);
tran (tlvp_rsm_usr_ob_rdata[22], \tlvp_rsm_usr_ob_rdata.tdata [22]);
tran (tlvp_rsm_usr_ob_rdata[21], \tlvp_rsm_usr_ob_rdata.tdata [21]);
tran (tlvp_rsm_usr_ob_rdata[20], \tlvp_rsm_usr_ob_rdata.tdata [20]);
tran (tlvp_rsm_usr_ob_rdata[19], \tlvp_rsm_usr_ob_rdata.tdata [19]);
tran (tlvp_rsm_usr_ob_rdata[18], \tlvp_rsm_usr_ob_rdata.tdata [18]);
tran (tlvp_rsm_usr_ob_rdata[17], \tlvp_rsm_usr_ob_rdata.tdata [17]);
tran (tlvp_rsm_usr_ob_rdata[16], \tlvp_rsm_usr_ob_rdata.tdata [16]);
tran (tlvp_rsm_usr_ob_rdata[15], \tlvp_rsm_usr_ob_rdata.tdata [15]);
tran (tlvp_rsm_usr_ob_rdata[14], \tlvp_rsm_usr_ob_rdata.tdata [14]);
tran (tlvp_rsm_usr_ob_rdata[13], \tlvp_rsm_usr_ob_rdata.tdata [13]);
tran (tlvp_rsm_usr_ob_rdata[12], \tlvp_rsm_usr_ob_rdata.tdata [12]);
tran (tlvp_rsm_usr_ob_rdata[11], \tlvp_rsm_usr_ob_rdata.tdata [11]);
tran (tlvp_rsm_usr_ob_rdata[10], \tlvp_rsm_usr_ob_rdata.tdata [10]);
tran (tlvp_rsm_usr_ob_rdata[9], \tlvp_rsm_usr_ob_rdata.tdata [9]);
tran (tlvp_rsm_usr_ob_rdata[8], \tlvp_rsm_usr_ob_rdata.tdata [8]);
tran (tlvp_rsm_usr_ob_rdata[7], \tlvp_rsm_usr_ob_rdata.tdata [7]);
tran (tlvp_rsm_usr_ob_rdata[6], \tlvp_rsm_usr_ob_rdata.tdata [6]);
tran (tlvp_rsm_usr_ob_rdata[5], \tlvp_rsm_usr_ob_rdata.tdata [5]);
tran (tlvp_rsm_usr_ob_rdata[4], \tlvp_rsm_usr_ob_rdata.tdata [4]);
tran (tlvp_rsm_usr_ob_rdata[3], \tlvp_rsm_usr_ob_rdata.tdata [3]);
tran (tlvp_rsm_usr_ob_rdata[2], \tlvp_rsm_usr_ob_rdata.tdata [2]);
tran (tlvp_rsm_usr_ob_rdata[1], \tlvp_rsm_usr_ob_rdata.tdata [1]);
tran (tlvp_rsm_usr_ob_rdata[0], \tlvp_rsm_usr_ob_rdata.tdata [0]);
ixc_assign _zz_strnp_0 ( _zy_simnet_pt_ob_rd_0_w$, pt_ob_rd);
ixc_assign _zz_strnp_1 ( _zy_simnet_usr_ob_full_1_w$, usr_ob_full);
ixc_assign _zz_strnp_2 ( _zy_simnet_usr_ob_afull_2_w$, usr_ob_afull);
ixc_assign _zz_strnp_3 ( _zy_simnet_tlvp_ob_empty_3_w$, tlvp_ob_empty);
ixc_assign _zz_strnp_4 ( _zy_simnet_tlvp_ob_aempty_4_w$, tlvp_ob_aempty);
ixc_assign_83 _zz_strnp_5 ( _zy_simnet_tlvp_ob_5_w$[0:82], tlvp_ob[82:0]);
ixc_assign _zz_strnp_6 ( _zy_simnet_tlvp_rsm_bimc_odat_6_w$, 
	tlvp_rsm_bimc_odat);
ixc_assign _zz_strnp_7 ( _zy_simnet_tlvp_rsm_bimc_osync_7_w$, 
	tlvp_rsm_bimc_osync);
ixc_assign _zz_strnp_8 ( _zy_simnet_tlvp_ob_ro_uncorrectable_ecc_error_8_w$, 
	tlvp_ob_ro_uncorrectable_ecc_error);
ixc_assign _zz_strnp_9 ( _zy_simnet_usr_ob_ro_uncorrectable_ecc_error_9_w$, 
	usr_ob_ro_uncorrectable_ecc_error);
ixc_assign _zz_strnp_10 ( pt_ob_rd, _zy_simnet_pt_ob_rd_10_w$);
ixc_assign _zz_strnp_11 ( tlvp_rsm_usr_ob_ren, 
	_zy_simnet_tlvp_rsm_usr_ob_ren_11_w$);
ixc_assign _zz_strnp_12 ( tlvp_rsm_ob_wen, _zy_simnet_tlvp_rsm_ob_wen_12_w$);
ixc_assign_83 _zz_strnp_13 ( tlvp_rsm_ob_wdata[82:0], 
	_zy_simnet_tlvp_rsm_ob_wdata_13_w$[0:82]);
ixc_assign_106 _zz_strnp_14 ( _zy_simnet_tlvp_rsm_usr_ob_rdata_14_w$[0:105], 
	tlvp_rsm_usr_ob_rdata[105:0]);
ixc_assign _zz_strnp_15 ( _zy_simnet_usr_ob_empty_15_w$, usr_ob_empty);
ixc_assign _zz_strnp_16 ( _zy_simnet_usr_ob_aempty_16_w$, usr_ob_aempty);
ixc_assign _zz_strnp_17 ( _zy_simnet_tlvp_ob_full_17_w$, tlvp_ob_full);
ixc_assign _zz_strnp_18 ( _zy_simnet_tlvp_ob_afull_18_w$, tlvp_ob_afull);
ixc_assign _zz_strnp_19 ( tlvp_ob_full, _zy_simnet_tlvp_ob_full_19_w$);
ixc_assign _zz_strnp_20 ( tlvp_ob_afull, _zy_simnet_tlvp_ob_afull_20_w$);
ixc_assign_83 _zz_strnp_21 ( tlvp_ob[82:0], _zy_simnet_tlvp_ob_21_w$[0:82]);
ixc_assign _zz_strnp_22 ( tlvp_ob_empty, _zy_simnet_tlvp_ob_empty_22_w$);
ixc_assign _zz_strnp_23 ( tlvp_ob_aempty, _zy_simnet_tlvp_ob_aempty_23_w$);
ixc_assign _zz_strnp_24 ( tlvp_rsm_bimc_odat, 
	_zy_simnet_tlvp_rsm_bimc_odat_24_w$);
ixc_assign _zz_strnp_25 ( tlvp_rsm_bimc_osync, 
	_zy_simnet_tlvp_rsm_bimc_osync_25_w$);
ixc_assign _zz_strnp_26 ( tlvp_ob_ro_uncorrectable_ecc_error, 
	_zy_simnet_tlvp_ob_ro_uncorrectable_ecc_error_26_w$);
ixc_assign_83 _zz_strnp_27 ( _zy_simnet_tlvp_rsm_ob_wdata_27_w$[0:82], 
	tlvp_rsm_ob_wdata[82:0]);
ixc_assign _zz_strnp_28 ( _zy_simnet_tlvp_rsm_ob_wen_28_w$, tlvp_rsm_ob_wen);
ixc_assign _zz_strnp_29 ( _zy_simnet_usr_ob_bimc_odat_29_w$, usr_ob_bimc_odat);
ixc_assign _zz_strnp_30 ( _zy_simnet_usr_ob_bimc_osync_30_w$, 
	usr_ob_bimc_osync);
ixc_assign _zz_strnp_31 ( usr_ob_full, _zy_simnet_usr_ob_full_31_w$);
ixc_assign _zz_strnp_32 ( usr_ob_afull, _zy_simnet_usr_ob_afull_32_w$);
ixc_assign_106 _zz_strnp_33 ( tlvp_rsm_usr_ob_rdata[105:0], 
	_zy_simnet_tlvp_rsm_usr_ob_rdata_33_w$[0:105]);
ixc_assign _zz_strnp_34 ( usr_ob_empty, _zy_simnet_usr_ob_empty_34_w$);
ixc_assign _zz_strnp_35 ( usr_ob_aempty, _zy_simnet_usr_ob_aempty_35_w$);
ixc_assign _zz_strnp_36 ( usr_ob_bimc_odat, _zy_simnet_usr_ob_bimc_odat_36_w$);
ixc_assign _zz_strnp_37 ( usr_ob_bimc_osync, 
	_zy_simnet_usr_ob_bimc_osync_37_w$);
ixc_assign _zz_strnp_38 ( usr_ob_ro_uncorrectable_ecc_error, 
	_zy_simnet_usr_ob_ro_uncorrectable_ecc_error_38_w$);
ixc_assign _zz_strnp_39 ( _zy_simnet_tlvp_rsm_usr_ob_ren_39_w$, 
	tlvp_rsm_usr_ob_ren);
cr_tlvp2_rsm_core u_cr_tlvp2_rsm_core ( .pt_ob_rd( _zy_simnet_pt_ob_rd_10_w$), 
	.tlvp_rsm_usr_ob_ren( _zy_simnet_tlvp_rsm_usr_ob_ren_11_w$), 
	.tlvp_rsm_ob_wen( _zy_simnet_tlvp_rsm_ob_wen_12_w$), 
	.tlvp_rsm_ob_wdata( _zy_simnet_tlvp_rsm_ob_wdata_13_w$[0:82]), .clk( 
	clk), .rst_n( rst_n), .pt_ob_empty( pt_ob_empty), .pt_ob_aempty( 
	pt_ob_aempty), .pt_ob_tlv( pt_ob_tlv[105:0]), 
	.tlvp_rsm_usr_ob_rdata( _zy_simnet_tlvp_rsm_usr_ob_rdata_14_w$[0:105]), 
	.usr_ob_empty( _zy_simnet_usr_ob_empty_15_w$), .usr_ob_aempty( 
	_zy_simnet_usr_ob_aempty_16_w$), .tlvp_ob_full( 
	_zy_simnet_tlvp_ob_full_17_w$), .tlvp_ob_afull( 
	_zy_simnet_tlvp_ob_afull_18_w$));
cr_fifo_wrap2_xcm9 u_cr_fifo_wrap2_tob ( .full( 
	_zy_simnet_tlvp_ob_full_19_w$), .afull( 
	_zy_simnet_tlvp_ob_afull_20_w$), .rdata( 
	_zy_simnet_tlvp_ob_21_w$[0:82]), .empty( 
	_zy_simnet_tlvp_ob_empty_22_w$), .aempty( 
	_zy_simnet_tlvp_ob_aempty_23_w$), .bimc_odat( 
	_zy_simnet_tlvp_rsm_bimc_odat_24_w$), .bimc_osync( 
	_zy_simnet_tlvp_rsm_bimc_osync_25_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_tlvp_ob_ro_uncorrectable_ecc_error_26_w$), .clk( clk), 
	.rst_n( rst_n), .wdata( _zy_simnet_tlvp_rsm_ob_wdata_27_w$[0:82]), 
	.wen( _zy_simnet_tlvp_rsm_ob_wen_28_w$), .ren( tlvp_ob_rd), 
	.bimc_idat( _zy_simnet_usr_ob_bimc_odat_29_w$), .bimc_isync( 
	_zy_simnet_usr_ob_bimc_osync_30_w$), .bimc_rst_n( bimc_rst_n));
cr_fifo_wrap2_xcm8 u_cr_fifo_wrap2_uobf ( .full( 
	_zy_simnet_usr_ob_full_31_w$), .afull( 
	_zy_simnet_usr_ob_afull_32_w$), .rdata( 
	_zy_simnet_tlvp_rsm_usr_ob_rdata_33_w$[0:105]), .empty( 
	_zy_simnet_usr_ob_empty_34_w$), .aempty( 
	_zy_simnet_usr_ob_aempty_35_w$), .bimc_odat( 
	_zy_simnet_usr_ob_bimc_odat_36_w$), .bimc_osync( 
	_zy_simnet_usr_ob_bimc_osync_37_w$), .ro_uncorrectable_ecc_error( 
	_zy_simnet_usr_ob_ro_uncorrectable_ecc_error_38_w$), .clk( clk), 
	.rst_n( rst_n), .wdata( usr_ob_tlv[105:0]), .wen( usr_ob_wr), 
	.ren( _zy_simnet_tlvp_rsm_usr_ob_ren_39_w$), .bimc_idat( 
	tlvp_rsm_bimc_idat), .bimc_isync( tlvp_rsm_bimc_isync), 
	.bimc_rst_n( bimc_rst_n));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\tlvp_ob.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\tlvp_ob.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\tlvp_ob.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\tlvp_ob.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\pt_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\pt_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\pt_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\pt_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\pt_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\pt_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\usr_ob_tlv.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\usr_ob_tlv.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\usr_ob_tlv.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\usr_ob_tlv.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\usr_ob_tlv.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\usr_ob_tlv.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\tlvp_rsm_usr_ob_rdata.ordern  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\tlvp_rsm_usr_ob_rdata.typen  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\tlvp_rsm_usr_ob_rdata.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\tlvp_rsm_usr_ob_rdata.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\tlvp_rsm_usr_ob_rdata.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\tlvp_rsm_usr_ob_rdata.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\tlvp_rsm_ob_wdata.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\tlvp_rsm_ob_wdata.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\tlvp_rsm_ob_wdata.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\tlvp_rsm_ob_wdata.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "26"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "tlvp_ob 6 \tlvp_ob.tvalid  \tlvp_ob.tlast  \tlvp_ob.tid  \tlvp_ob.tstrb  \tlvp_ob.tuser  \tlvp_ob.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "pt_ob_tlv 10 \pt_ob_tlv.insert  \pt_ob_tlv.ordern  \pt_ob_tlv.typen  \pt_ob_tlv.sot  \pt_ob_tlv.eot  \pt_ob_tlv.tlast  \pt_ob_tlv.tid  \pt_ob_tlv.tstrb  \pt_ob_tlv.tuser  \pt_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "usr_ob_tlv 10 \usr_ob_tlv.insert  \usr_ob_tlv.ordern  \usr_ob_tlv.typen  \usr_ob_tlv.sot  \usr_ob_tlv.eot  \usr_ob_tlv.tlast  \usr_ob_tlv.tid  \usr_ob_tlv.tstrb  \usr_ob_tlv.tuser  \usr_ob_tlv.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "tlvp_rsm_usr_ob_rdata 10 \tlvp_rsm_usr_ob_rdata.insert  \tlvp_rsm_usr_ob_rdata.ordern  \tlvp_rsm_usr_ob_rdata.typen  \tlvp_rsm_usr_ob_rdata.sot  \tlvp_rsm_usr_ob_rdata.eot  \tlvp_rsm_usr_ob_rdata.tlast  \tlvp_rsm_usr_ob_rdata.tid  \tlvp_rsm_usr_ob_rdata.tstrb  \tlvp_rsm_usr_ob_rdata.tuser  \tlvp_rsm_usr_ob_rdata.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "tlvp_rsm_ob_wdata 6 \tlvp_rsm_ob_wdata.tvalid  \tlvp_rsm_ob_wdata.tlast  \tlvp_rsm_ob_wdata.tid  \tlvp_rsm_ob_wdata.tstrb  \tlvp_rsm_ob_wdata.tuser  \tlvp_rsm_ob_wdata.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "5"
endmodule
