
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_gfifo_port_64_0_0 ( tkout, tkin, ireq, cbid, len, idata, CGFtsReq, 
	CGFcbid, CGFlen, CGFidata, CGFfull, CLBreq, CLBrd, CLBwr, CLBfull, 
	Rtkin);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output tkout;
input tkin;
input ireq;
input [19:0] cbid;
input [11:0] len;
input [63:0] idata;
output CGFtsReq;
output [19:0] CGFcbid;
output [11:0] CGFlen;
output [511:0] CGFidata;
input CGFfull;
output CLBreq;
input [3:0] CLBrd;
input [3:0] CLBwr;
input CLBfull;
input Rtkin;
wire fclk;
wire enq;
wire CLBreqWhileFull;
`_2_ wire en;
`_2_ wire ack;
`_2_ wire [63:0] odata;
`_2_ wire oreq;
`_2_ wire [19:0] ocbid;
`_2_ wire [19:0] xcbid;
`_2_ wire [11:0] olen;
`_2_ wire [11:0] xlen;
`_2_ wire [0:0] sel;
`_2_ wire [63:0] xdata;
wire [31:0] i;
`_2_ wire ireqR;
supply1 n5;
Q_ASSIGN U0 ( .B(len[0]), .A(xlen[0]));
Q_ASSIGN U1 ( .B(len[0]), .A(olen[0]));
Q_ASSIGN U2 ( .B(len[1]), .A(xlen[1]));
Q_ASSIGN U3 ( .B(len[1]), .A(olen[1]));
Q_ASSIGN U4 ( .B(len[2]), .A(xlen[2]));
Q_ASSIGN U5 ( .B(len[2]), .A(olen[2]));
Q_ASSIGN U6 ( .B(len[3]), .A(xlen[3]));
Q_ASSIGN U7 ( .B(len[3]), .A(olen[3]));
Q_ASSIGN U8 ( .B(len[4]), .A(xlen[4]));
Q_ASSIGN U9 ( .B(len[4]), .A(olen[4]));
Q_ASSIGN U10 ( .B(len[5]), .A(xlen[5]));
Q_ASSIGN U11 ( .B(len[5]), .A(olen[5]));
Q_ASSIGN U12 ( .B(len[6]), .A(xlen[6]));
Q_ASSIGN U13 ( .B(len[6]), .A(olen[6]));
Q_ASSIGN U14 ( .B(len[7]), .A(xlen[7]));
Q_ASSIGN U15 ( .B(len[7]), .A(olen[7]));
Q_ASSIGN U16 ( .B(len[8]), .A(xlen[8]));
Q_ASSIGN U17 ( .B(len[8]), .A(olen[8]));
Q_ASSIGN U18 ( .B(len[9]), .A(xlen[9]));
Q_ASSIGN U19 ( .B(len[9]), .A(olen[9]));
Q_ASSIGN U20 ( .B(len[10]), .A(xlen[10]));
Q_ASSIGN U21 ( .B(len[10]), .A(olen[10]));
Q_ASSIGN U22 ( .B(len[11]), .A(xlen[11]));
Q_ASSIGN U23 ( .B(len[11]), .A(olen[11]));
Q_ASSIGN U24 ( .B(cbid[0]), .A(xcbid[0]));
Q_ASSIGN U25 ( .B(cbid[0]), .A(ocbid[0]));
Q_ASSIGN U26 ( .B(cbid[1]), .A(xcbid[1]));
Q_ASSIGN U27 ( .B(cbid[1]), .A(ocbid[1]));
Q_ASSIGN U28 ( .B(cbid[2]), .A(xcbid[2]));
Q_ASSIGN U29 ( .B(cbid[2]), .A(ocbid[2]));
Q_ASSIGN U30 ( .B(cbid[3]), .A(xcbid[3]));
Q_ASSIGN U31 ( .B(cbid[3]), .A(ocbid[3]));
Q_ASSIGN U32 ( .B(cbid[4]), .A(xcbid[4]));
Q_ASSIGN U33 ( .B(cbid[4]), .A(ocbid[4]));
Q_ASSIGN U34 ( .B(cbid[5]), .A(xcbid[5]));
Q_ASSIGN U35 ( .B(cbid[5]), .A(ocbid[5]));
Q_ASSIGN U36 ( .B(cbid[6]), .A(xcbid[6]));
Q_ASSIGN U37 ( .B(cbid[6]), .A(ocbid[6]));
Q_ASSIGN U38 ( .B(cbid[7]), .A(xcbid[7]));
Q_ASSIGN U39 ( .B(cbid[7]), .A(ocbid[7]));
Q_ASSIGN U40 ( .B(cbid[8]), .A(xcbid[8]));
Q_ASSIGN U41 ( .B(cbid[8]), .A(ocbid[8]));
Q_ASSIGN U42 ( .B(cbid[9]), .A(xcbid[9]));
Q_ASSIGN U43 ( .B(cbid[9]), .A(ocbid[9]));
Q_ASSIGN U44 ( .B(cbid[10]), .A(xcbid[10]));
Q_ASSIGN U45 ( .B(cbid[10]), .A(ocbid[10]));
Q_ASSIGN U46 ( .B(cbid[11]), .A(xcbid[11]));
Q_ASSIGN U47 ( .B(cbid[11]), .A(ocbid[11]));
Q_ASSIGN U48 ( .B(cbid[12]), .A(xcbid[12]));
Q_ASSIGN U49 ( .B(cbid[12]), .A(ocbid[12]));
Q_ASSIGN U50 ( .B(cbid[13]), .A(xcbid[13]));
Q_ASSIGN U51 ( .B(cbid[13]), .A(ocbid[13]));
Q_ASSIGN U52 ( .B(cbid[14]), .A(xcbid[14]));
Q_ASSIGN U53 ( .B(cbid[14]), .A(ocbid[14]));
Q_ASSIGN U54 ( .B(cbid[15]), .A(xcbid[15]));
Q_ASSIGN U55 ( .B(cbid[15]), .A(ocbid[15]));
Q_ASSIGN U56 ( .B(cbid[16]), .A(xcbid[16]));
Q_ASSIGN U57 ( .B(cbid[16]), .A(ocbid[16]));
Q_ASSIGN U58 ( .B(cbid[17]), .A(xcbid[17]));
Q_ASSIGN U59 ( .B(cbid[17]), .A(ocbid[17]));
Q_ASSIGN U60 ( .B(cbid[18]), .A(xcbid[18]));
Q_ASSIGN U61 ( .B(cbid[18]), .A(ocbid[18]));
Q_ASSIGN U62 ( .B(cbid[19]), .A(xcbid[19]));
Q_ASSIGN U63 ( .B(cbid[19]), .A(ocbid[19]));
Q_BUF U64 ( .A(odata[0]), .Z(xdata[0]));
Q_BUF U65 ( .A(odata[1]), .Z(xdata[1]));
Q_BUF U66 ( .A(odata[2]), .Z(xdata[2]));
Q_BUF U67 ( .A(odata[3]), .Z(xdata[3]));
Q_BUF U68 ( .A(odata[4]), .Z(xdata[4]));
Q_BUF U69 ( .A(odata[5]), .Z(xdata[5]));
Q_BUF U70 ( .A(odata[6]), .Z(xdata[6]));
Q_BUF U71 ( .A(odata[7]), .Z(xdata[7]));
Q_BUF U72 ( .A(odata[8]), .Z(xdata[8]));
Q_BUF U73 ( .A(odata[9]), .Z(xdata[9]));
Q_BUF U74 ( .A(odata[10]), .Z(xdata[10]));
Q_BUF U75 ( .A(odata[11]), .Z(xdata[11]));
Q_BUF U76 ( .A(odata[12]), .Z(xdata[12]));
Q_BUF U77 ( .A(odata[13]), .Z(xdata[13]));
Q_BUF U78 ( .A(odata[14]), .Z(xdata[14]));
Q_BUF U79 ( .A(odata[15]), .Z(xdata[15]));
Q_BUF U80 ( .A(odata[16]), .Z(xdata[16]));
Q_BUF U81 ( .A(odata[17]), .Z(xdata[17]));
Q_BUF U82 ( .A(odata[18]), .Z(xdata[18]));
Q_BUF U83 ( .A(odata[19]), .Z(xdata[19]));
Q_BUF U84 ( .A(odata[20]), .Z(xdata[20]));
Q_BUF U85 ( .A(odata[21]), .Z(xdata[21]));
Q_BUF U86 ( .A(odata[22]), .Z(xdata[22]));
Q_BUF U87 ( .A(odata[23]), .Z(xdata[23]));
Q_BUF U88 ( .A(odata[24]), .Z(xdata[24]));
Q_BUF U89 ( .A(odata[25]), .Z(xdata[25]));
Q_BUF U90 ( .A(odata[26]), .Z(xdata[26]));
Q_BUF U91 ( .A(odata[27]), .Z(xdata[27]));
Q_BUF U92 ( .A(odata[28]), .Z(xdata[28]));
Q_BUF U93 ( .A(odata[29]), .Z(xdata[29]));
Q_BUF U94 ( .A(odata[30]), .Z(xdata[30]));
Q_BUF U95 ( .A(odata[31]), .Z(xdata[31]));
Q_BUF U96 ( .A(odata[32]), .Z(xdata[32]));
Q_BUF U97 ( .A(odata[33]), .Z(xdata[33]));
Q_BUF U98 ( .A(odata[34]), .Z(xdata[34]));
Q_BUF U99 ( .A(odata[35]), .Z(xdata[35]));
Q_BUF U100 ( .A(odata[36]), .Z(xdata[36]));
Q_BUF U101 ( .A(odata[37]), .Z(xdata[37]));
Q_BUF U102 ( .A(odata[38]), .Z(xdata[38]));
Q_BUF U103 ( .A(odata[39]), .Z(xdata[39]));
Q_BUF U104 ( .A(odata[40]), .Z(xdata[40]));
Q_BUF U105 ( .A(odata[41]), .Z(xdata[41]));
Q_BUF U106 ( .A(odata[42]), .Z(xdata[42]));
Q_BUF U107 ( .A(odata[43]), .Z(xdata[43]));
Q_BUF U108 ( .A(odata[44]), .Z(xdata[44]));
Q_BUF U109 ( .A(odata[45]), .Z(xdata[45]));
Q_BUF U110 ( .A(odata[46]), .Z(xdata[46]));
Q_BUF U111 ( .A(odata[47]), .Z(xdata[47]));
Q_BUF U112 ( .A(odata[48]), .Z(xdata[48]));
Q_BUF U113 ( .A(odata[49]), .Z(xdata[49]));
Q_BUF U114 ( .A(odata[50]), .Z(xdata[50]));
Q_BUF U115 ( .A(odata[51]), .Z(xdata[51]));
Q_BUF U116 ( .A(odata[52]), .Z(xdata[52]));
Q_BUF U117 ( .A(odata[53]), .Z(xdata[53]));
Q_BUF U118 ( .A(odata[54]), .Z(xdata[54]));
Q_BUF U119 ( .A(odata[55]), .Z(xdata[55]));
Q_BUF U120 ( .A(odata[56]), .Z(xdata[56]));
Q_BUF U121 ( .A(odata[57]), .Z(xdata[57]));
Q_BUF U122 ( .A(odata[58]), .Z(xdata[58]));
Q_BUF U123 ( .A(odata[59]), .Z(xdata[59]));
Q_BUF U124 ( .A(odata[60]), .Z(xdata[60]));
Q_BUF U125 ( .A(odata[61]), .Z(xdata[61]));
Q_BUF U126 ( .A(odata[62]), .Z(xdata[62]));
Q_BUF U127 ( .A(odata[63]), .Z(xdata[63]));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_EV_WOR_START qi ( .A(CLBreqWhileFull));
Q_INV U130 ( .A(n4), .Z(tkout));
Q_XNR2 U131 ( .A0(oreq), .A1(ack), .Z(n4));
Q_CCLKCHK cchk ( .sig(ireq));
Q_AN02 U133 ( .A0(enq), .A1(CLBfull), .Z(CLBreqWhileFull));
Q_AN02 U134 ( .A0(n2), .A1(n3), .Z(enq));
Q_INV U135 ( .A(xc_top.GFLock2), .Z(n3));
Q_XOR2 U136 ( .A0(ireq), .A1(ireqR), .Z(n2));
Q_BUFZP U137 ( .OE(CLBreqWhileFull), .A(n5), .Z(xc_top.GFLBfull));
Q_BUFZP U138 ( .OE(en), .A(cbid[0]), .Z(CGFcbid[0]));
Q_BUFZP U139 ( .OE(en), .A(cbid[1]), .Z(CGFcbid[1]));
Q_BUFZP U140 ( .OE(en), .A(cbid[2]), .Z(CGFcbid[2]));
Q_BUFZP U141 ( .OE(en), .A(cbid[3]), .Z(CGFcbid[3]));
Q_BUFZP U142 ( .OE(en), .A(cbid[4]), .Z(CGFcbid[4]));
Q_BUFZP U143 ( .OE(en), .A(cbid[5]), .Z(CGFcbid[5]));
Q_BUFZP U144 ( .OE(en), .A(cbid[6]), .Z(CGFcbid[6]));
Q_BUFZP U145 ( .OE(en), .A(cbid[7]), .Z(CGFcbid[7]));
Q_BUFZP U146 ( .OE(en), .A(cbid[8]), .Z(CGFcbid[8]));
Q_BUFZP U147 ( .OE(en), .A(cbid[9]), .Z(CGFcbid[9]));
Q_BUFZP U148 ( .OE(en), .A(cbid[10]), .Z(CGFcbid[10]));
Q_BUFZP U149 ( .OE(en), .A(cbid[11]), .Z(CGFcbid[11]));
Q_BUFZP U150 ( .OE(en), .A(cbid[12]), .Z(CGFcbid[12]));
Q_BUFZP U151 ( .OE(en), .A(cbid[13]), .Z(CGFcbid[13]));
Q_BUFZP U152 ( .OE(en), .A(cbid[14]), .Z(CGFcbid[14]));
Q_BUFZP U153 ( .OE(en), .A(cbid[15]), .Z(CGFcbid[15]));
Q_BUFZP U154 ( .OE(en), .A(cbid[16]), .Z(CGFcbid[16]));
Q_BUFZP U155 ( .OE(en), .A(cbid[17]), .Z(CGFcbid[17]));
Q_BUFZP U156 ( .OE(en), .A(cbid[18]), .Z(CGFcbid[18]));
Q_BUFZP U157 ( .OE(en), .A(cbid[19]), .Z(CGFcbid[19]));
Q_BUFZP U158 ( .OE(en), .A(len[0]), .Z(CGFlen[0]));
Q_BUFZP U159 ( .OE(en), .A(len[1]), .Z(CGFlen[1]));
Q_BUFZP U160 ( .OE(en), .A(len[2]), .Z(CGFlen[2]));
Q_BUFZP U161 ( .OE(en), .A(len[3]), .Z(CGFlen[3]));
Q_BUFZP U162 ( .OE(en), .A(len[4]), .Z(CGFlen[4]));
Q_BUFZP U163 ( .OE(en), .A(len[5]), .Z(CGFlen[5]));
Q_BUFZP U164 ( .OE(en), .A(len[6]), .Z(CGFlen[6]));
Q_BUFZP U165 ( .OE(en), .A(len[7]), .Z(CGFlen[7]));
Q_BUFZP U166 ( .OE(en), .A(len[8]), .Z(CGFlen[8]));
Q_BUFZP U167 ( .OE(en), .A(len[9]), .Z(CGFlen[9]));
Q_BUFZP U168 ( .OE(en), .A(len[10]), .Z(CGFlen[10]));
Q_BUFZP U169 ( .OE(en), .A(len[11]), .Z(CGFlen[11]));
Q_BUFZP U170 ( .OE(en), .A(xdata[0]), .Z(CGFidata[0]));
Q_BUFZP U171 ( .OE(en), .A(xdata[1]), .Z(CGFidata[1]));
Q_BUFZP U172 ( .OE(en), .A(xdata[2]), .Z(CGFidata[2]));
Q_BUFZP U173 ( .OE(en), .A(xdata[3]), .Z(CGFidata[3]));
Q_BUFZP U174 ( .OE(en), .A(xdata[4]), .Z(CGFidata[4]));
Q_BUFZP U175 ( .OE(en), .A(xdata[5]), .Z(CGFidata[5]));
Q_BUFZP U176 ( .OE(en), .A(xdata[6]), .Z(CGFidata[6]));
Q_BUFZP U177 ( .OE(en), .A(xdata[7]), .Z(CGFidata[7]));
Q_BUFZP U178 ( .OE(en), .A(xdata[8]), .Z(CGFidata[8]));
Q_BUFZP U179 ( .OE(en), .A(xdata[9]), .Z(CGFidata[9]));
Q_BUFZP U180 ( .OE(en), .A(xdata[10]), .Z(CGFidata[10]));
Q_BUFZP U181 ( .OE(en), .A(xdata[11]), .Z(CGFidata[11]));
Q_BUFZP U182 ( .OE(en), .A(xdata[12]), .Z(CGFidata[12]));
Q_BUFZP U183 ( .OE(en), .A(xdata[13]), .Z(CGFidata[13]));
Q_BUFZP U184 ( .OE(en), .A(xdata[14]), .Z(CGFidata[14]));
Q_BUFZP U185 ( .OE(en), .A(xdata[15]), .Z(CGFidata[15]));
Q_BUFZP U186 ( .OE(en), .A(xdata[16]), .Z(CGFidata[16]));
Q_BUFZP U187 ( .OE(en), .A(xdata[17]), .Z(CGFidata[17]));
Q_BUFZP U188 ( .OE(en), .A(xdata[18]), .Z(CGFidata[18]));
Q_BUFZP U189 ( .OE(en), .A(xdata[19]), .Z(CGFidata[19]));
Q_BUFZP U190 ( .OE(en), .A(xdata[20]), .Z(CGFidata[20]));
Q_BUFZP U191 ( .OE(en), .A(xdata[21]), .Z(CGFidata[21]));
Q_BUFZP U192 ( .OE(en), .A(xdata[22]), .Z(CGFidata[22]));
Q_BUFZP U193 ( .OE(en), .A(xdata[23]), .Z(CGFidata[23]));
Q_BUFZP U194 ( .OE(en), .A(xdata[24]), .Z(CGFidata[24]));
Q_BUFZP U195 ( .OE(en), .A(xdata[25]), .Z(CGFidata[25]));
Q_BUFZP U196 ( .OE(en), .A(xdata[26]), .Z(CGFidata[26]));
Q_BUFZP U197 ( .OE(en), .A(xdata[27]), .Z(CGFidata[27]));
Q_BUFZP U198 ( .OE(en), .A(xdata[28]), .Z(CGFidata[28]));
Q_BUFZP U199 ( .OE(en), .A(xdata[29]), .Z(CGFidata[29]));
Q_BUFZP U200 ( .OE(en), .A(xdata[30]), .Z(CGFidata[30]));
Q_BUFZP U201 ( .OE(en), .A(xdata[31]), .Z(CGFidata[31]));
Q_BUFZP U202 ( .OE(en), .A(xdata[32]), .Z(CGFidata[32]));
Q_BUFZP U203 ( .OE(en), .A(xdata[33]), .Z(CGFidata[33]));
Q_BUFZP U204 ( .OE(en), .A(xdata[34]), .Z(CGFidata[34]));
Q_BUFZP U205 ( .OE(en), .A(xdata[35]), .Z(CGFidata[35]));
Q_BUFZP U206 ( .OE(en), .A(xdata[36]), .Z(CGFidata[36]));
Q_BUFZP U207 ( .OE(en), .A(xdata[37]), .Z(CGFidata[37]));
Q_BUFZP U208 ( .OE(en), .A(xdata[38]), .Z(CGFidata[38]));
Q_BUFZP U209 ( .OE(en), .A(xdata[39]), .Z(CGFidata[39]));
Q_BUFZP U210 ( .OE(en), .A(xdata[40]), .Z(CGFidata[40]));
Q_BUFZP U211 ( .OE(en), .A(xdata[41]), .Z(CGFidata[41]));
Q_BUFZP U212 ( .OE(en), .A(xdata[42]), .Z(CGFidata[42]));
Q_BUFZP U213 ( .OE(en), .A(xdata[43]), .Z(CGFidata[43]));
Q_BUFZP U214 ( .OE(en), .A(xdata[44]), .Z(CGFidata[44]));
Q_BUFZP U215 ( .OE(en), .A(xdata[45]), .Z(CGFidata[45]));
Q_BUFZP U216 ( .OE(en), .A(xdata[46]), .Z(CGFidata[46]));
Q_BUFZP U217 ( .OE(en), .A(xdata[47]), .Z(CGFidata[47]));
Q_BUFZP U218 ( .OE(en), .A(xdata[48]), .Z(CGFidata[48]));
Q_BUFZP U219 ( .OE(en), .A(xdata[49]), .Z(CGFidata[49]));
Q_BUFZP U220 ( .OE(en), .A(xdata[50]), .Z(CGFidata[50]));
Q_BUFZP U221 ( .OE(en), .A(xdata[51]), .Z(CGFidata[51]));
Q_BUFZP U222 ( .OE(en), .A(xdata[52]), .Z(CGFidata[52]));
Q_BUFZP U223 ( .OE(en), .A(xdata[53]), .Z(CGFidata[53]));
Q_BUFZP U224 ( .OE(en), .A(xdata[54]), .Z(CGFidata[54]));
Q_BUFZP U225 ( .OE(en), .A(xdata[55]), .Z(CGFidata[55]));
Q_BUFZP U226 ( .OE(en), .A(xdata[56]), .Z(CGFidata[56]));
Q_BUFZP U227 ( .OE(en), .A(xdata[57]), .Z(CGFidata[57]));
Q_BUFZP U228 ( .OE(en), .A(xdata[58]), .Z(CGFidata[58]));
Q_BUFZP U229 ( .OE(en), .A(xdata[59]), .Z(CGFidata[59]));
Q_BUFZP U230 ( .OE(en), .A(xdata[60]), .Z(CGFidata[60]));
Q_BUFZP U231 ( .OE(en), .A(xdata[61]), .Z(CGFidata[61]));
Q_BUFZP U232 ( .OE(en), .A(xdata[62]), .Z(CGFidata[62]));
Q_BUFZP U233 ( .OE(en), .A(xdata[63]), .Z(CGFidata[63]));
Q_BUFZP U234 ( .OE(enq), .A(n5), .Z(CLBreq));
Q_INV U235 ( .A(CLBwr[2]), .Z(n6));
ixc_bind \genblk3.b5 ( CLBfull, IXC_GFIFO.O.O.LBfull);
ixc_bind_4 \genblk3.b4 ( CLBwr[3:0], IXC_GFIFO.O.O.LBwr[3:0]);
ixc_bind_4 \genblk3.b3 ( CLBrd[3:0], IXC_GFIFO.O.O.LBrd[3:0]);
ixc_bind \genblk3.b2 ( CLBreq, IXC_GFIFO.O.O.LBreq);
ixc_bind \genblk3.b1 ( CGFfull, IXC_GFIFO.O.O.GFfull);
ixc_bind \genblk3.b0 ( CGFtsReq, IXC_GFIFO.O.O.GFtsReq);
Q_MX02 U242 ( .S(xc_top.GFLock2), .A0(oreq), .A1(ireq), .Z(n8));
Q_FDP0UA U243 ( .D(n9), .QTFCLK( ), .Q(ack));
Q_MX02 U244 ( .S(n14), .A0(ack), .A1(n8), .Z(n9));
Q_FDP0UA U245 ( .D(n10), .QTFCLK( ), .Q(en));
Q_NR02 U246 ( .A0(xc_top.GFLock2), .A1(n11), .Z(n10));
Q_OR02 U247 ( .A0(xc_top.GFLock2), .A1(n12), .Z(n14));
Q_INV U248 ( .A(n11), .Z(n12));
Q_OR03 U249 ( .A0(n4), .A1(tkin), .A2(n13), .Z(n11));
Q_OR02 U250 ( .A0(Rtkin), .A1(CGFfull), .Z(n13));
Q_MX02 U251 ( .S(CLBfull), .A0(ireq), .A1(ireqR), .Z(n15));
Q_FDP0UA U252 ( .D(n15), .QTFCLK( ), .Q(ireqR));
Q_AN02 U253 ( .A0(CLBwr[0]), .A1(n6), .Z(n16));
Q_AN02 U254 ( .A0(CLBwr[1]), .A1(n6), .Z(n17));
Q_INV U255 ( .A(n16), .Z(n18));
Q_INV U256 ( .A(n17), .Z(n19));
Q_NR02 U257 ( .A0(n17), .A1(n16), .Z(n20));
Q_AN02 U258 ( .A0(n19), .A1(n16), .Z(n21));
Q_AN02 U259 ( .A0(n17), .A1(n18), .Z(n22));
Q_AN02 U260 ( .A0(n17), .A1(n16), .Z(n23));
Q_AN02 U261 ( .A0(n20), .A1(n6), .Z(n24));
Q_LDP0 \_zzLB_REG[0][0] ( .G(n24), .D(idata[0]), .Q(\_zzLB[0][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][1] ( .G(n24), .D(idata[1]), .Q(\_zzLB[0][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][2] ( .G(n24), .D(idata[2]), .Q(\_zzLB[0][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][3] ( .G(n24), .D(idata[3]), .Q(\_zzLB[0][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][4] ( .G(n24), .D(idata[4]), .Q(\_zzLB[0][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][5] ( .G(n24), .D(idata[5]), .Q(\_zzLB[0][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][6] ( .G(n24), .D(idata[6]), .Q(\_zzLB[0][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][7] ( .G(n24), .D(idata[7]), .Q(\_zzLB[0][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][8] ( .G(n24), .D(idata[8]), .Q(\_zzLB[0][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][9] ( .G(n24), .D(idata[9]), .Q(\_zzLB[0][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][10] ( .G(n24), .D(idata[10]), .Q(\_zzLB[0][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][11] ( .G(n24), .D(idata[11]), .Q(\_zzLB[0][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][12] ( .G(n24), .D(idata[12]), .Q(\_zzLB[0][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][13] ( .G(n24), .D(idata[13]), .Q(\_zzLB[0][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][14] ( .G(n24), .D(idata[14]), .Q(\_zzLB[0][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][15] ( .G(n24), .D(idata[15]), .Q(\_zzLB[0][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][16] ( .G(n24), .D(idata[16]), .Q(\_zzLB[0][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][17] ( .G(n24), .D(idata[17]), .Q(\_zzLB[0][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][18] ( .G(n24), .D(idata[18]), .Q(\_zzLB[0][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][19] ( .G(n24), .D(idata[19]), .Q(\_zzLB[0][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][20] ( .G(n24), .D(idata[20]), .Q(\_zzLB[0][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][21] ( .G(n24), .D(idata[21]), .Q(\_zzLB[0][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][22] ( .G(n24), .D(idata[22]), .Q(\_zzLB[0][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][23] ( .G(n24), .D(idata[23]), .Q(\_zzLB[0][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][24] ( .G(n24), .D(idata[24]), .Q(\_zzLB[0][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][25] ( .G(n24), .D(idata[25]), .Q(\_zzLB[0][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][26] ( .G(n24), .D(idata[26]), .Q(\_zzLB[0][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][27] ( .G(n24), .D(idata[27]), .Q(\_zzLB[0][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][28] ( .G(n24), .D(idata[28]), .Q(\_zzLB[0][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][29] ( .G(n24), .D(idata[29]), .Q(\_zzLB[0][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][30] ( .G(n24), .D(idata[30]), .Q(\_zzLB[0][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][31] ( .G(n24), .D(idata[31]), .Q(\_zzLB[0][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][32] ( .G(n24), .D(idata[32]), .Q(\_zzLB[0][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][33] ( .G(n24), .D(idata[33]), .Q(\_zzLB[0][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][34] ( .G(n24), .D(idata[34]), .Q(\_zzLB[0][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][35] ( .G(n24), .D(idata[35]), .Q(\_zzLB[0][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][36] ( .G(n24), .D(idata[36]), .Q(\_zzLB[0][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][37] ( .G(n24), .D(idata[37]), .Q(\_zzLB[0][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][38] ( .G(n24), .D(idata[38]), .Q(\_zzLB[0][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][39] ( .G(n24), .D(idata[39]), .Q(\_zzLB[0][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][40] ( .G(n24), .D(idata[40]), .Q(\_zzLB[0][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][41] ( .G(n24), .D(idata[41]), .Q(\_zzLB[0][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][42] ( .G(n24), .D(idata[42]), .Q(\_zzLB[0][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][43] ( .G(n24), .D(idata[43]), .Q(\_zzLB[0][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][44] ( .G(n24), .D(idata[44]), .Q(\_zzLB[0][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][45] ( .G(n24), .D(idata[45]), .Q(\_zzLB[0][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][46] ( .G(n24), .D(idata[46]), .Q(\_zzLB[0][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][47] ( .G(n24), .D(idata[47]), .Q(\_zzLB[0][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][48] ( .G(n24), .D(idata[48]), .Q(\_zzLB[0][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][49] ( .G(n24), .D(idata[49]), .Q(\_zzLB[0][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][50] ( .G(n24), .D(idata[50]), .Q(\_zzLB[0][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][51] ( .G(n24), .D(idata[51]), .Q(\_zzLB[0][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][52] ( .G(n24), .D(idata[52]), .Q(\_zzLB[0][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][53] ( .G(n24), .D(idata[53]), .Q(\_zzLB[0][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][54] ( .G(n24), .D(idata[54]), .Q(\_zzLB[0][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][55] ( .G(n24), .D(idata[55]), .Q(\_zzLB[0][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][56] ( .G(n24), .D(idata[56]), .Q(\_zzLB[0][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][57] ( .G(n24), .D(idata[57]), .Q(\_zzLB[0][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][58] ( .G(n24), .D(idata[58]), .Q(\_zzLB[0][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][59] ( .G(n24), .D(idata[59]), .Q(\_zzLB[0][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][60] ( .G(n24), .D(idata[60]), .Q(\_zzLB[0][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][61] ( .G(n24), .D(idata[61]), .Q(\_zzLB[0][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][62] ( .G(n24), .D(idata[62]), .Q(\_zzLB[0][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][63] ( .G(n24), .D(idata[63]), .Q(\_zzLB[0][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][64] ( .G(n24), .D(ireq), .Q(\_zzLB[0][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][0] ( .G(n21), .D(idata[0]), .Q(\_zzLB[1][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][1] ( .G(n21), .D(idata[1]), .Q(\_zzLB[1][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][2] ( .G(n21), .D(idata[2]), .Q(\_zzLB[1][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][3] ( .G(n21), .D(idata[3]), .Q(\_zzLB[1][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][4] ( .G(n21), .D(idata[4]), .Q(\_zzLB[1][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][5] ( .G(n21), .D(idata[5]), .Q(\_zzLB[1][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][6] ( .G(n21), .D(idata[6]), .Q(\_zzLB[1][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][7] ( .G(n21), .D(idata[7]), .Q(\_zzLB[1][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][8] ( .G(n21), .D(idata[8]), .Q(\_zzLB[1][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][9] ( .G(n21), .D(idata[9]), .Q(\_zzLB[1][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][10] ( .G(n21), .D(idata[10]), .Q(\_zzLB[1][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][11] ( .G(n21), .D(idata[11]), .Q(\_zzLB[1][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][12] ( .G(n21), .D(idata[12]), .Q(\_zzLB[1][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][13] ( .G(n21), .D(idata[13]), .Q(\_zzLB[1][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][14] ( .G(n21), .D(idata[14]), .Q(\_zzLB[1][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][15] ( .G(n21), .D(idata[15]), .Q(\_zzLB[1][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][16] ( .G(n21), .D(idata[16]), .Q(\_zzLB[1][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][17] ( .G(n21), .D(idata[17]), .Q(\_zzLB[1][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][18] ( .G(n21), .D(idata[18]), .Q(\_zzLB[1][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][19] ( .G(n21), .D(idata[19]), .Q(\_zzLB[1][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][20] ( .G(n21), .D(idata[20]), .Q(\_zzLB[1][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][21] ( .G(n21), .D(idata[21]), .Q(\_zzLB[1][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][22] ( .G(n21), .D(idata[22]), .Q(\_zzLB[1][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][23] ( .G(n21), .D(idata[23]), .Q(\_zzLB[1][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][24] ( .G(n21), .D(idata[24]), .Q(\_zzLB[1][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][25] ( .G(n21), .D(idata[25]), .Q(\_zzLB[1][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][26] ( .G(n21), .D(idata[26]), .Q(\_zzLB[1][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][27] ( .G(n21), .D(idata[27]), .Q(\_zzLB[1][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][28] ( .G(n21), .D(idata[28]), .Q(\_zzLB[1][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][29] ( .G(n21), .D(idata[29]), .Q(\_zzLB[1][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][30] ( .G(n21), .D(idata[30]), .Q(\_zzLB[1][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][31] ( .G(n21), .D(idata[31]), .Q(\_zzLB[1][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][32] ( .G(n21), .D(idata[32]), .Q(\_zzLB[1][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][33] ( .G(n21), .D(idata[33]), .Q(\_zzLB[1][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][34] ( .G(n21), .D(idata[34]), .Q(\_zzLB[1][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][35] ( .G(n21), .D(idata[35]), .Q(\_zzLB[1][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][36] ( .G(n21), .D(idata[36]), .Q(\_zzLB[1][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][37] ( .G(n21), .D(idata[37]), .Q(\_zzLB[1][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][38] ( .G(n21), .D(idata[38]), .Q(\_zzLB[1][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][39] ( .G(n21), .D(idata[39]), .Q(\_zzLB[1][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][40] ( .G(n21), .D(idata[40]), .Q(\_zzLB[1][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][41] ( .G(n21), .D(idata[41]), .Q(\_zzLB[1][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][42] ( .G(n21), .D(idata[42]), .Q(\_zzLB[1][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][43] ( .G(n21), .D(idata[43]), .Q(\_zzLB[1][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][44] ( .G(n21), .D(idata[44]), .Q(\_zzLB[1][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][45] ( .G(n21), .D(idata[45]), .Q(\_zzLB[1][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][46] ( .G(n21), .D(idata[46]), .Q(\_zzLB[1][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][47] ( .G(n21), .D(idata[47]), .Q(\_zzLB[1][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][48] ( .G(n21), .D(idata[48]), .Q(\_zzLB[1][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][49] ( .G(n21), .D(idata[49]), .Q(\_zzLB[1][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][50] ( .G(n21), .D(idata[50]), .Q(\_zzLB[1][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][51] ( .G(n21), .D(idata[51]), .Q(\_zzLB[1][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][52] ( .G(n21), .D(idata[52]), .Q(\_zzLB[1][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][53] ( .G(n21), .D(idata[53]), .Q(\_zzLB[1][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][54] ( .G(n21), .D(idata[54]), .Q(\_zzLB[1][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][55] ( .G(n21), .D(idata[55]), .Q(\_zzLB[1][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][56] ( .G(n21), .D(idata[56]), .Q(\_zzLB[1][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][57] ( .G(n21), .D(idata[57]), .Q(\_zzLB[1][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][58] ( .G(n21), .D(idata[58]), .Q(\_zzLB[1][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][59] ( .G(n21), .D(idata[59]), .Q(\_zzLB[1][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][60] ( .G(n21), .D(idata[60]), .Q(\_zzLB[1][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][61] ( .G(n21), .D(idata[61]), .Q(\_zzLB[1][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][62] ( .G(n21), .D(idata[62]), .Q(\_zzLB[1][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][63] ( .G(n21), .D(idata[63]), .Q(\_zzLB[1][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][64] ( .G(n21), .D(ireq), .Q(\_zzLB[1][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][0] ( .G(n22), .D(idata[0]), .Q(\_zzLB[2][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][1] ( .G(n22), .D(idata[1]), .Q(\_zzLB[2][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][2] ( .G(n22), .D(idata[2]), .Q(\_zzLB[2][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][3] ( .G(n22), .D(idata[3]), .Q(\_zzLB[2][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][4] ( .G(n22), .D(idata[4]), .Q(\_zzLB[2][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][5] ( .G(n22), .D(idata[5]), .Q(\_zzLB[2][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][6] ( .G(n22), .D(idata[6]), .Q(\_zzLB[2][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][7] ( .G(n22), .D(idata[7]), .Q(\_zzLB[2][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][8] ( .G(n22), .D(idata[8]), .Q(\_zzLB[2][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][9] ( .G(n22), .D(idata[9]), .Q(\_zzLB[2][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][10] ( .G(n22), .D(idata[10]), .Q(\_zzLB[2][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][11] ( .G(n22), .D(idata[11]), .Q(\_zzLB[2][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][12] ( .G(n22), .D(idata[12]), .Q(\_zzLB[2][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][13] ( .G(n22), .D(idata[13]), .Q(\_zzLB[2][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][14] ( .G(n22), .D(idata[14]), .Q(\_zzLB[2][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][15] ( .G(n22), .D(idata[15]), .Q(\_zzLB[2][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][16] ( .G(n22), .D(idata[16]), .Q(\_zzLB[2][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][17] ( .G(n22), .D(idata[17]), .Q(\_zzLB[2][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][18] ( .G(n22), .D(idata[18]), .Q(\_zzLB[2][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][19] ( .G(n22), .D(idata[19]), .Q(\_zzLB[2][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][20] ( .G(n22), .D(idata[20]), .Q(\_zzLB[2][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][21] ( .G(n22), .D(idata[21]), .Q(\_zzLB[2][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][22] ( .G(n22), .D(idata[22]), .Q(\_zzLB[2][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][23] ( .G(n22), .D(idata[23]), .Q(\_zzLB[2][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][24] ( .G(n22), .D(idata[24]), .Q(\_zzLB[2][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][25] ( .G(n22), .D(idata[25]), .Q(\_zzLB[2][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][26] ( .G(n22), .D(idata[26]), .Q(\_zzLB[2][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][27] ( .G(n22), .D(idata[27]), .Q(\_zzLB[2][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][28] ( .G(n22), .D(idata[28]), .Q(\_zzLB[2][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][29] ( .G(n22), .D(idata[29]), .Q(\_zzLB[2][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][30] ( .G(n22), .D(idata[30]), .Q(\_zzLB[2][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][31] ( .G(n22), .D(idata[31]), .Q(\_zzLB[2][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][32] ( .G(n22), .D(idata[32]), .Q(\_zzLB[2][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][33] ( .G(n22), .D(idata[33]), .Q(\_zzLB[2][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][34] ( .G(n22), .D(idata[34]), .Q(\_zzLB[2][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][35] ( .G(n22), .D(idata[35]), .Q(\_zzLB[2][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][36] ( .G(n22), .D(idata[36]), .Q(\_zzLB[2][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][37] ( .G(n22), .D(idata[37]), .Q(\_zzLB[2][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][38] ( .G(n22), .D(idata[38]), .Q(\_zzLB[2][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][39] ( .G(n22), .D(idata[39]), .Q(\_zzLB[2][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][40] ( .G(n22), .D(idata[40]), .Q(\_zzLB[2][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][41] ( .G(n22), .D(idata[41]), .Q(\_zzLB[2][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][42] ( .G(n22), .D(idata[42]), .Q(\_zzLB[2][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][43] ( .G(n22), .D(idata[43]), .Q(\_zzLB[2][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][44] ( .G(n22), .D(idata[44]), .Q(\_zzLB[2][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][45] ( .G(n22), .D(idata[45]), .Q(\_zzLB[2][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][46] ( .G(n22), .D(idata[46]), .Q(\_zzLB[2][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][47] ( .G(n22), .D(idata[47]), .Q(\_zzLB[2][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][48] ( .G(n22), .D(idata[48]), .Q(\_zzLB[2][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][49] ( .G(n22), .D(idata[49]), .Q(\_zzLB[2][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][50] ( .G(n22), .D(idata[50]), .Q(\_zzLB[2][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][51] ( .G(n22), .D(idata[51]), .Q(\_zzLB[2][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][52] ( .G(n22), .D(idata[52]), .Q(\_zzLB[2][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][53] ( .G(n22), .D(idata[53]), .Q(\_zzLB[2][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][54] ( .G(n22), .D(idata[54]), .Q(\_zzLB[2][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][55] ( .G(n22), .D(idata[55]), .Q(\_zzLB[2][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][56] ( .G(n22), .D(idata[56]), .Q(\_zzLB[2][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][57] ( .G(n22), .D(idata[57]), .Q(\_zzLB[2][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][58] ( .G(n22), .D(idata[58]), .Q(\_zzLB[2][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][59] ( .G(n22), .D(idata[59]), .Q(\_zzLB[2][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][60] ( .G(n22), .D(idata[60]), .Q(\_zzLB[2][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][61] ( .G(n22), .D(idata[61]), .Q(\_zzLB[2][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][62] ( .G(n22), .D(idata[62]), .Q(\_zzLB[2][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][63] ( .G(n22), .D(idata[63]), .Q(\_zzLB[2][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][64] ( .G(n22), .D(ireq), .Q(\_zzLB[2][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][0] ( .G(n23), .D(idata[0]), .Q(\_zzLB[3][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][1] ( .G(n23), .D(idata[1]), .Q(\_zzLB[3][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][2] ( .G(n23), .D(idata[2]), .Q(\_zzLB[3][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][3] ( .G(n23), .D(idata[3]), .Q(\_zzLB[3][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][4] ( .G(n23), .D(idata[4]), .Q(\_zzLB[3][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][5] ( .G(n23), .D(idata[5]), .Q(\_zzLB[3][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][6] ( .G(n23), .D(idata[6]), .Q(\_zzLB[3][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][7] ( .G(n23), .D(idata[7]), .Q(\_zzLB[3][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][8] ( .G(n23), .D(idata[8]), .Q(\_zzLB[3][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][9] ( .G(n23), .D(idata[9]), .Q(\_zzLB[3][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][10] ( .G(n23), .D(idata[10]), .Q(\_zzLB[3][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][11] ( .G(n23), .D(idata[11]), .Q(\_zzLB[3][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][12] ( .G(n23), .D(idata[12]), .Q(\_zzLB[3][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][13] ( .G(n23), .D(idata[13]), .Q(\_zzLB[3][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][14] ( .G(n23), .D(idata[14]), .Q(\_zzLB[3][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][15] ( .G(n23), .D(idata[15]), .Q(\_zzLB[3][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][16] ( .G(n23), .D(idata[16]), .Q(\_zzLB[3][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][17] ( .G(n23), .D(idata[17]), .Q(\_zzLB[3][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][18] ( .G(n23), .D(idata[18]), .Q(\_zzLB[3][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][19] ( .G(n23), .D(idata[19]), .Q(\_zzLB[3][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][20] ( .G(n23), .D(idata[20]), .Q(\_zzLB[3][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][21] ( .G(n23), .D(idata[21]), .Q(\_zzLB[3][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][22] ( .G(n23), .D(idata[22]), .Q(\_zzLB[3][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][23] ( .G(n23), .D(idata[23]), .Q(\_zzLB[3][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][24] ( .G(n23), .D(idata[24]), .Q(\_zzLB[3][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][25] ( .G(n23), .D(idata[25]), .Q(\_zzLB[3][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][26] ( .G(n23), .D(idata[26]), .Q(\_zzLB[3][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][27] ( .G(n23), .D(idata[27]), .Q(\_zzLB[3][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][28] ( .G(n23), .D(idata[28]), .Q(\_zzLB[3][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][29] ( .G(n23), .D(idata[29]), .Q(\_zzLB[3][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][30] ( .G(n23), .D(idata[30]), .Q(\_zzLB[3][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][31] ( .G(n23), .D(idata[31]), .Q(\_zzLB[3][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][32] ( .G(n23), .D(idata[32]), .Q(\_zzLB[3][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][33] ( .G(n23), .D(idata[33]), .Q(\_zzLB[3][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][34] ( .G(n23), .D(idata[34]), .Q(\_zzLB[3][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][35] ( .G(n23), .D(idata[35]), .Q(\_zzLB[3][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][36] ( .G(n23), .D(idata[36]), .Q(\_zzLB[3][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][37] ( .G(n23), .D(idata[37]), .Q(\_zzLB[3][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][38] ( .G(n23), .D(idata[38]), .Q(\_zzLB[3][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][39] ( .G(n23), .D(idata[39]), .Q(\_zzLB[3][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][40] ( .G(n23), .D(idata[40]), .Q(\_zzLB[3][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][41] ( .G(n23), .D(idata[41]), .Q(\_zzLB[3][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][42] ( .G(n23), .D(idata[42]), .Q(\_zzLB[3][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][43] ( .G(n23), .D(idata[43]), .Q(\_zzLB[3][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][44] ( .G(n23), .D(idata[44]), .Q(\_zzLB[3][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][45] ( .G(n23), .D(idata[45]), .Q(\_zzLB[3][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][46] ( .G(n23), .D(idata[46]), .Q(\_zzLB[3][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][47] ( .G(n23), .D(idata[47]), .Q(\_zzLB[3][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][48] ( .G(n23), .D(idata[48]), .Q(\_zzLB[3][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][49] ( .G(n23), .D(idata[49]), .Q(\_zzLB[3][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][50] ( .G(n23), .D(idata[50]), .Q(\_zzLB[3][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][51] ( .G(n23), .D(idata[51]), .Q(\_zzLB[3][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][52] ( .G(n23), .D(idata[52]), .Q(\_zzLB[3][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][53] ( .G(n23), .D(idata[53]), .Q(\_zzLB[3][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][54] ( .G(n23), .D(idata[54]), .Q(\_zzLB[3][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][55] ( .G(n23), .D(idata[55]), .Q(\_zzLB[3][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][56] ( .G(n23), .D(idata[56]), .Q(\_zzLB[3][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][57] ( .G(n23), .D(idata[57]), .Q(\_zzLB[3][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][58] ( .G(n23), .D(idata[58]), .Q(\_zzLB[3][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][59] ( .G(n23), .D(idata[59]), .Q(\_zzLB[3][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][60] ( .G(n23), .D(idata[60]), .Q(\_zzLB[3][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][61] ( .G(n23), .D(idata[61]), .Q(\_zzLB[3][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][62] ( .G(n23), .D(idata[62]), .Q(\_zzLB[3][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][63] ( .G(n23), .D(idata[63]), .Q(\_zzLB[3][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][64] ( .G(n23), .D(ireq), .Q(\_zzLB[3][64] ), .QN( ));
Q_MX04 U522 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][0] ), .A1(\_zzLB[1][0] ), .A2(\_zzLB[2][0] ), .A3(\_zzLB[3][0] ), .Z(odata[0]));
Q_MX04 U523 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][1] ), .A1(\_zzLB[1][1] ), .A2(\_zzLB[2][1] ), .A3(\_zzLB[3][1] ), .Z(odata[1]));
Q_MX04 U524 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][2] ), .A1(\_zzLB[1][2] ), .A2(\_zzLB[2][2] ), .A3(\_zzLB[3][2] ), .Z(odata[2]));
Q_MX04 U525 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][3] ), .A1(\_zzLB[1][3] ), .A2(\_zzLB[2][3] ), .A3(\_zzLB[3][3] ), .Z(odata[3]));
Q_MX04 U526 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][4] ), .A1(\_zzLB[1][4] ), .A2(\_zzLB[2][4] ), .A3(\_zzLB[3][4] ), .Z(odata[4]));
Q_MX04 U527 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][5] ), .A1(\_zzLB[1][5] ), .A2(\_zzLB[2][5] ), .A3(\_zzLB[3][5] ), .Z(odata[5]));
Q_MX04 U528 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][6] ), .A1(\_zzLB[1][6] ), .A2(\_zzLB[2][6] ), .A3(\_zzLB[3][6] ), .Z(odata[6]));
Q_MX04 U529 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][7] ), .A1(\_zzLB[1][7] ), .A2(\_zzLB[2][7] ), .A3(\_zzLB[3][7] ), .Z(odata[7]));
Q_MX04 U530 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][8] ), .A1(\_zzLB[1][8] ), .A2(\_zzLB[2][8] ), .A3(\_zzLB[3][8] ), .Z(odata[8]));
Q_MX04 U531 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][9] ), .A1(\_zzLB[1][9] ), .A2(\_zzLB[2][9] ), .A3(\_zzLB[3][9] ), .Z(odata[9]));
Q_MX04 U532 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][10] ), .A1(\_zzLB[1][10] ), .A2(\_zzLB[2][10] ), .A3(\_zzLB[3][10] ), .Z(odata[10]));
Q_MX04 U533 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][11] ), .A1(\_zzLB[1][11] ), .A2(\_zzLB[2][11] ), .A3(\_zzLB[3][11] ), .Z(odata[11]));
Q_MX04 U534 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][12] ), .A1(\_zzLB[1][12] ), .A2(\_zzLB[2][12] ), .A3(\_zzLB[3][12] ), .Z(odata[12]));
Q_MX04 U535 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][13] ), .A1(\_zzLB[1][13] ), .A2(\_zzLB[2][13] ), .A3(\_zzLB[3][13] ), .Z(odata[13]));
Q_MX04 U536 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][14] ), .A1(\_zzLB[1][14] ), .A2(\_zzLB[2][14] ), .A3(\_zzLB[3][14] ), .Z(odata[14]));
Q_MX04 U537 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][15] ), .A1(\_zzLB[1][15] ), .A2(\_zzLB[2][15] ), .A3(\_zzLB[3][15] ), .Z(odata[15]));
Q_MX04 U538 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][16] ), .A1(\_zzLB[1][16] ), .A2(\_zzLB[2][16] ), .A3(\_zzLB[3][16] ), .Z(odata[16]));
Q_MX04 U539 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][17] ), .A1(\_zzLB[1][17] ), .A2(\_zzLB[2][17] ), .A3(\_zzLB[3][17] ), .Z(odata[17]));
Q_MX04 U540 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][18] ), .A1(\_zzLB[1][18] ), .A2(\_zzLB[2][18] ), .A3(\_zzLB[3][18] ), .Z(odata[18]));
Q_MX04 U541 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][19] ), .A1(\_zzLB[1][19] ), .A2(\_zzLB[2][19] ), .A3(\_zzLB[3][19] ), .Z(odata[19]));
Q_MX04 U542 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][20] ), .A1(\_zzLB[1][20] ), .A2(\_zzLB[2][20] ), .A3(\_zzLB[3][20] ), .Z(odata[20]));
Q_MX04 U543 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][21] ), .A1(\_zzLB[1][21] ), .A2(\_zzLB[2][21] ), .A3(\_zzLB[3][21] ), .Z(odata[21]));
Q_MX04 U544 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][22] ), .A1(\_zzLB[1][22] ), .A2(\_zzLB[2][22] ), .A3(\_zzLB[3][22] ), .Z(odata[22]));
Q_MX04 U545 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][23] ), .A1(\_zzLB[1][23] ), .A2(\_zzLB[2][23] ), .A3(\_zzLB[3][23] ), .Z(odata[23]));
Q_MX04 U546 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][24] ), .A1(\_zzLB[1][24] ), .A2(\_zzLB[2][24] ), .A3(\_zzLB[3][24] ), .Z(odata[24]));
Q_MX04 U547 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][25] ), .A1(\_zzLB[1][25] ), .A2(\_zzLB[2][25] ), .A3(\_zzLB[3][25] ), .Z(odata[25]));
Q_MX04 U548 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][26] ), .A1(\_zzLB[1][26] ), .A2(\_zzLB[2][26] ), .A3(\_zzLB[3][26] ), .Z(odata[26]));
Q_MX04 U549 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][27] ), .A1(\_zzLB[1][27] ), .A2(\_zzLB[2][27] ), .A3(\_zzLB[3][27] ), .Z(odata[27]));
Q_MX04 U550 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][28] ), .A1(\_zzLB[1][28] ), .A2(\_zzLB[2][28] ), .A3(\_zzLB[3][28] ), .Z(odata[28]));
Q_MX04 U551 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][29] ), .A1(\_zzLB[1][29] ), .A2(\_zzLB[2][29] ), .A3(\_zzLB[3][29] ), .Z(odata[29]));
Q_MX04 U552 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][30] ), .A1(\_zzLB[1][30] ), .A2(\_zzLB[2][30] ), .A3(\_zzLB[3][30] ), .Z(odata[30]));
Q_MX04 U553 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][31] ), .A1(\_zzLB[1][31] ), .A2(\_zzLB[2][31] ), .A3(\_zzLB[3][31] ), .Z(odata[31]));
Q_MX04 U554 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][32] ), .A1(\_zzLB[1][32] ), .A2(\_zzLB[2][32] ), .A3(\_zzLB[3][32] ), .Z(odata[32]));
Q_MX04 U555 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][33] ), .A1(\_zzLB[1][33] ), .A2(\_zzLB[2][33] ), .A3(\_zzLB[3][33] ), .Z(odata[33]));
Q_MX04 U556 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][34] ), .A1(\_zzLB[1][34] ), .A2(\_zzLB[2][34] ), .A3(\_zzLB[3][34] ), .Z(odata[34]));
Q_MX04 U557 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][35] ), .A1(\_zzLB[1][35] ), .A2(\_zzLB[2][35] ), .A3(\_zzLB[3][35] ), .Z(odata[35]));
Q_MX04 U558 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][36] ), .A1(\_zzLB[1][36] ), .A2(\_zzLB[2][36] ), .A3(\_zzLB[3][36] ), .Z(odata[36]));
Q_MX04 U559 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][37] ), .A1(\_zzLB[1][37] ), .A2(\_zzLB[2][37] ), .A3(\_zzLB[3][37] ), .Z(odata[37]));
Q_MX04 U560 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][38] ), .A1(\_zzLB[1][38] ), .A2(\_zzLB[2][38] ), .A3(\_zzLB[3][38] ), .Z(odata[38]));
Q_MX04 U561 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][39] ), .A1(\_zzLB[1][39] ), .A2(\_zzLB[2][39] ), .A3(\_zzLB[3][39] ), .Z(odata[39]));
Q_MX04 U562 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][40] ), .A1(\_zzLB[1][40] ), .A2(\_zzLB[2][40] ), .A3(\_zzLB[3][40] ), .Z(odata[40]));
Q_MX04 U563 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][41] ), .A1(\_zzLB[1][41] ), .A2(\_zzLB[2][41] ), .A3(\_zzLB[3][41] ), .Z(odata[41]));
Q_MX04 U564 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][42] ), .A1(\_zzLB[1][42] ), .A2(\_zzLB[2][42] ), .A3(\_zzLB[3][42] ), .Z(odata[42]));
Q_MX04 U565 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][43] ), .A1(\_zzLB[1][43] ), .A2(\_zzLB[2][43] ), .A3(\_zzLB[3][43] ), .Z(odata[43]));
Q_MX04 U566 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][44] ), .A1(\_zzLB[1][44] ), .A2(\_zzLB[2][44] ), .A3(\_zzLB[3][44] ), .Z(odata[44]));
Q_MX04 U567 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][45] ), .A1(\_zzLB[1][45] ), .A2(\_zzLB[2][45] ), .A3(\_zzLB[3][45] ), .Z(odata[45]));
Q_MX04 U568 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][46] ), .A1(\_zzLB[1][46] ), .A2(\_zzLB[2][46] ), .A3(\_zzLB[3][46] ), .Z(odata[46]));
Q_MX04 U569 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][47] ), .A1(\_zzLB[1][47] ), .A2(\_zzLB[2][47] ), .A3(\_zzLB[3][47] ), .Z(odata[47]));
Q_MX04 U570 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][48] ), .A1(\_zzLB[1][48] ), .A2(\_zzLB[2][48] ), .A3(\_zzLB[3][48] ), .Z(odata[48]));
Q_MX04 U571 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][49] ), .A1(\_zzLB[1][49] ), .A2(\_zzLB[2][49] ), .A3(\_zzLB[3][49] ), .Z(odata[49]));
Q_MX04 U572 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][50] ), .A1(\_zzLB[1][50] ), .A2(\_zzLB[2][50] ), .A3(\_zzLB[3][50] ), .Z(odata[50]));
Q_MX04 U573 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][51] ), .A1(\_zzLB[1][51] ), .A2(\_zzLB[2][51] ), .A3(\_zzLB[3][51] ), .Z(odata[51]));
Q_MX04 U574 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][52] ), .A1(\_zzLB[1][52] ), .A2(\_zzLB[2][52] ), .A3(\_zzLB[3][52] ), .Z(odata[52]));
Q_MX04 U575 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][53] ), .A1(\_zzLB[1][53] ), .A2(\_zzLB[2][53] ), .A3(\_zzLB[3][53] ), .Z(odata[53]));
Q_MX04 U576 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][54] ), .A1(\_zzLB[1][54] ), .A2(\_zzLB[2][54] ), .A3(\_zzLB[3][54] ), .Z(odata[54]));
Q_MX04 U577 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][55] ), .A1(\_zzLB[1][55] ), .A2(\_zzLB[2][55] ), .A3(\_zzLB[3][55] ), .Z(odata[55]));
Q_MX04 U578 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][56] ), .A1(\_zzLB[1][56] ), .A2(\_zzLB[2][56] ), .A3(\_zzLB[3][56] ), .Z(odata[56]));
Q_MX04 U579 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][57] ), .A1(\_zzLB[1][57] ), .A2(\_zzLB[2][57] ), .A3(\_zzLB[3][57] ), .Z(odata[57]));
Q_MX04 U580 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][58] ), .A1(\_zzLB[1][58] ), .A2(\_zzLB[2][58] ), .A3(\_zzLB[3][58] ), .Z(odata[58]));
Q_MX04 U581 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][59] ), .A1(\_zzLB[1][59] ), .A2(\_zzLB[2][59] ), .A3(\_zzLB[3][59] ), .Z(odata[59]));
Q_MX04 U582 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][60] ), .A1(\_zzLB[1][60] ), .A2(\_zzLB[2][60] ), .A3(\_zzLB[3][60] ), .Z(odata[60]));
Q_MX04 U583 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][61] ), .A1(\_zzLB[1][61] ), .A2(\_zzLB[2][61] ), .A3(\_zzLB[3][61] ), .Z(odata[61]));
Q_MX04 U584 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][62] ), .A1(\_zzLB[1][62] ), .A2(\_zzLB[2][62] ), .A3(\_zzLB[3][62] ), .Z(odata[62]));
Q_MX04 U585 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][63] ), .A1(\_zzLB[1][63] ), .A2(\_zzLB[2][63] ), .A3(\_zzLB[3][63] ), .Z(odata[63]));
Q_MX04 U586 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][64] ), .A1(\_zzLB[1][64] ), .A2(\_zzLB[2][64] ), .A3(\_zzLB[3][64] ), .Z(oreq));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zzLB 1 64 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_gfifo_port"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
