
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module ixc_assign_2176 ( L, R);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [2175:0] L;
input [2175:0] R;
Q_ASSIGN U0 ( .B(R[0]), .A(L[0]));
Q_ASSIGN U1 ( .B(R[1]), .A(L[1]));
Q_ASSIGN U2 ( .B(R[2]), .A(L[2]));
Q_ASSIGN U3 ( .B(R[3]), .A(L[3]));
Q_ASSIGN U4 ( .B(R[4]), .A(L[4]));
Q_ASSIGN U5 ( .B(R[5]), .A(L[5]));
Q_ASSIGN U6 ( .B(R[6]), .A(L[6]));
Q_ASSIGN U7 ( .B(R[7]), .A(L[7]));
Q_ASSIGN U8 ( .B(R[8]), .A(L[8]));
Q_ASSIGN U9 ( .B(R[9]), .A(L[9]));
Q_ASSIGN U10 ( .B(R[10]), .A(L[10]));
Q_ASSIGN U11 ( .B(R[11]), .A(L[11]));
Q_ASSIGN U12 ( .B(R[12]), .A(L[12]));
Q_ASSIGN U13 ( .B(R[13]), .A(L[13]));
Q_ASSIGN U14 ( .B(R[14]), .A(L[14]));
Q_ASSIGN U15 ( .B(R[15]), .A(L[15]));
Q_ASSIGN U16 ( .B(R[16]), .A(L[16]));
Q_ASSIGN U17 ( .B(R[17]), .A(L[17]));
Q_ASSIGN U18 ( .B(R[18]), .A(L[18]));
Q_ASSIGN U19 ( .B(R[19]), .A(L[19]));
Q_ASSIGN U20 ( .B(R[20]), .A(L[20]));
Q_ASSIGN U21 ( .B(R[21]), .A(L[21]));
Q_ASSIGN U22 ( .B(R[22]), .A(L[22]));
Q_ASSIGN U23 ( .B(R[23]), .A(L[23]));
Q_ASSIGN U24 ( .B(R[24]), .A(L[24]));
Q_ASSIGN U25 ( .B(R[25]), .A(L[25]));
Q_ASSIGN U26 ( .B(R[26]), .A(L[26]));
Q_ASSIGN U27 ( .B(R[27]), .A(L[27]));
Q_ASSIGN U28 ( .B(R[28]), .A(L[28]));
Q_ASSIGN U29 ( .B(R[29]), .A(L[29]));
Q_ASSIGN U30 ( .B(R[30]), .A(L[30]));
Q_ASSIGN U31 ( .B(R[31]), .A(L[31]));
Q_ASSIGN U32 ( .B(R[32]), .A(L[32]));
Q_ASSIGN U33 ( .B(R[33]), .A(L[33]));
Q_ASSIGN U34 ( .B(R[34]), .A(L[34]));
Q_ASSIGN U35 ( .B(R[35]), .A(L[35]));
Q_ASSIGN U36 ( .B(R[36]), .A(L[36]));
Q_ASSIGN U37 ( .B(R[37]), .A(L[37]));
Q_ASSIGN U38 ( .B(R[38]), .A(L[38]));
Q_ASSIGN U39 ( .B(R[39]), .A(L[39]));
Q_ASSIGN U40 ( .B(R[40]), .A(L[40]));
Q_ASSIGN U41 ( .B(R[41]), .A(L[41]));
Q_ASSIGN U42 ( .B(R[42]), .A(L[42]));
Q_ASSIGN U43 ( .B(R[43]), .A(L[43]));
Q_ASSIGN U44 ( .B(R[44]), .A(L[44]));
Q_ASSIGN U45 ( .B(R[45]), .A(L[45]));
Q_ASSIGN U46 ( .B(R[46]), .A(L[46]));
Q_ASSIGN U47 ( .B(R[47]), .A(L[47]));
Q_ASSIGN U48 ( .B(R[48]), .A(L[48]));
Q_ASSIGN U49 ( .B(R[49]), .A(L[49]));
Q_ASSIGN U50 ( .B(R[50]), .A(L[50]));
Q_ASSIGN U51 ( .B(R[51]), .A(L[51]));
Q_ASSIGN U52 ( .B(R[52]), .A(L[52]));
Q_ASSIGN U53 ( .B(R[53]), .A(L[53]));
Q_ASSIGN U54 ( .B(R[54]), .A(L[54]));
Q_ASSIGN U55 ( .B(R[55]), .A(L[55]));
Q_ASSIGN U56 ( .B(R[56]), .A(L[56]));
Q_ASSIGN U57 ( .B(R[57]), .A(L[57]));
Q_ASSIGN U58 ( .B(R[58]), .A(L[58]));
Q_ASSIGN U59 ( .B(R[59]), .A(L[59]));
Q_ASSIGN U60 ( .B(R[60]), .A(L[60]));
Q_ASSIGN U61 ( .B(R[61]), .A(L[61]));
Q_ASSIGN U62 ( .B(R[62]), .A(L[62]));
Q_ASSIGN U63 ( .B(R[63]), .A(L[63]));
Q_ASSIGN U64 ( .B(R[64]), .A(L[64]));
Q_ASSIGN U65 ( .B(R[65]), .A(L[65]));
Q_ASSIGN U66 ( .B(R[66]), .A(L[66]));
Q_ASSIGN U67 ( .B(R[67]), .A(L[67]));
Q_ASSIGN U68 ( .B(R[68]), .A(L[68]));
Q_ASSIGN U69 ( .B(R[69]), .A(L[69]));
Q_ASSIGN U70 ( .B(R[70]), .A(L[70]));
Q_ASSIGN U71 ( .B(R[71]), .A(L[71]));
Q_ASSIGN U72 ( .B(R[72]), .A(L[72]));
Q_ASSIGN U73 ( .B(R[73]), .A(L[73]));
Q_ASSIGN U74 ( .B(R[74]), .A(L[74]));
Q_ASSIGN U75 ( .B(R[75]), .A(L[75]));
Q_ASSIGN U76 ( .B(R[76]), .A(L[76]));
Q_ASSIGN U77 ( .B(R[77]), .A(L[77]));
Q_ASSIGN U78 ( .B(R[78]), .A(L[78]));
Q_ASSIGN U79 ( .B(R[79]), .A(L[79]));
Q_ASSIGN U80 ( .B(R[80]), .A(L[80]));
Q_ASSIGN U81 ( .B(R[81]), .A(L[81]));
Q_ASSIGN U82 ( .B(R[82]), .A(L[82]));
Q_ASSIGN U83 ( .B(R[83]), .A(L[83]));
Q_ASSIGN U84 ( .B(R[84]), .A(L[84]));
Q_ASSIGN U85 ( .B(R[85]), .A(L[85]));
Q_ASSIGN U86 ( .B(R[86]), .A(L[86]));
Q_ASSIGN U87 ( .B(R[87]), .A(L[87]));
Q_ASSIGN U88 ( .B(R[88]), .A(L[88]));
Q_ASSIGN U89 ( .B(R[89]), .A(L[89]));
Q_ASSIGN U90 ( .B(R[90]), .A(L[90]));
Q_ASSIGN U91 ( .B(R[91]), .A(L[91]));
Q_ASSIGN U92 ( .B(R[92]), .A(L[92]));
Q_ASSIGN U93 ( .B(R[93]), .A(L[93]));
Q_ASSIGN U94 ( .B(R[94]), .A(L[94]));
Q_ASSIGN U95 ( .B(R[95]), .A(L[95]));
Q_ASSIGN U96 ( .B(R[96]), .A(L[96]));
Q_ASSIGN U97 ( .B(R[97]), .A(L[97]));
Q_ASSIGN U98 ( .B(R[98]), .A(L[98]));
Q_ASSIGN U99 ( .B(R[99]), .A(L[99]));
Q_ASSIGN U100 ( .B(R[100]), .A(L[100]));
Q_ASSIGN U101 ( .B(R[101]), .A(L[101]));
Q_ASSIGN U102 ( .B(R[102]), .A(L[102]));
Q_ASSIGN U103 ( .B(R[103]), .A(L[103]));
Q_ASSIGN U104 ( .B(R[104]), .A(L[104]));
Q_ASSIGN U105 ( .B(R[105]), .A(L[105]));
Q_ASSIGN U106 ( .B(R[106]), .A(L[106]));
Q_ASSIGN U107 ( .B(R[107]), .A(L[107]));
Q_ASSIGN U108 ( .B(R[108]), .A(L[108]));
Q_ASSIGN U109 ( .B(R[109]), .A(L[109]));
Q_ASSIGN U110 ( .B(R[110]), .A(L[110]));
Q_ASSIGN U111 ( .B(R[111]), .A(L[111]));
Q_ASSIGN U112 ( .B(R[112]), .A(L[112]));
Q_ASSIGN U113 ( .B(R[113]), .A(L[113]));
Q_ASSIGN U114 ( .B(R[114]), .A(L[114]));
Q_ASSIGN U115 ( .B(R[115]), .A(L[115]));
Q_ASSIGN U116 ( .B(R[116]), .A(L[116]));
Q_ASSIGN U117 ( .B(R[117]), .A(L[117]));
Q_ASSIGN U118 ( .B(R[118]), .A(L[118]));
Q_ASSIGN U119 ( .B(R[119]), .A(L[119]));
Q_ASSIGN U120 ( .B(R[120]), .A(L[120]));
Q_ASSIGN U121 ( .B(R[121]), .A(L[121]));
Q_ASSIGN U122 ( .B(R[122]), .A(L[122]));
Q_ASSIGN U123 ( .B(R[123]), .A(L[123]));
Q_ASSIGN U124 ( .B(R[124]), .A(L[124]));
Q_ASSIGN U125 ( .B(R[125]), .A(L[125]));
Q_ASSIGN U126 ( .B(R[126]), .A(L[126]));
Q_ASSIGN U127 ( .B(R[127]), .A(L[127]));
Q_ASSIGN U128 ( .B(R[128]), .A(L[128]));
Q_ASSIGN U129 ( .B(R[129]), .A(L[129]));
Q_ASSIGN U130 ( .B(R[130]), .A(L[130]));
Q_ASSIGN U131 ( .B(R[131]), .A(L[131]));
Q_ASSIGN U132 ( .B(R[132]), .A(L[132]));
Q_ASSIGN U133 ( .B(R[133]), .A(L[133]));
Q_ASSIGN U134 ( .B(R[134]), .A(L[134]));
Q_ASSIGN U135 ( .B(R[135]), .A(L[135]));
Q_ASSIGN U136 ( .B(R[136]), .A(L[136]));
Q_ASSIGN U137 ( .B(R[137]), .A(L[137]));
Q_ASSIGN U138 ( .B(R[138]), .A(L[138]));
Q_ASSIGN U139 ( .B(R[139]), .A(L[139]));
Q_ASSIGN U140 ( .B(R[140]), .A(L[140]));
Q_ASSIGN U141 ( .B(R[141]), .A(L[141]));
Q_ASSIGN U142 ( .B(R[142]), .A(L[142]));
Q_ASSIGN U143 ( .B(R[143]), .A(L[143]));
Q_ASSIGN U144 ( .B(R[144]), .A(L[144]));
Q_ASSIGN U145 ( .B(R[145]), .A(L[145]));
Q_ASSIGN U146 ( .B(R[146]), .A(L[146]));
Q_ASSIGN U147 ( .B(R[147]), .A(L[147]));
Q_ASSIGN U148 ( .B(R[148]), .A(L[148]));
Q_ASSIGN U149 ( .B(R[149]), .A(L[149]));
Q_ASSIGN U150 ( .B(R[150]), .A(L[150]));
Q_ASSIGN U151 ( .B(R[151]), .A(L[151]));
Q_ASSIGN U152 ( .B(R[152]), .A(L[152]));
Q_ASSIGN U153 ( .B(R[153]), .A(L[153]));
Q_ASSIGN U154 ( .B(R[154]), .A(L[154]));
Q_ASSIGN U155 ( .B(R[155]), .A(L[155]));
Q_ASSIGN U156 ( .B(R[156]), .A(L[156]));
Q_ASSIGN U157 ( .B(R[157]), .A(L[157]));
Q_ASSIGN U158 ( .B(R[158]), .A(L[158]));
Q_ASSIGN U159 ( .B(R[159]), .A(L[159]));
Q_ASSIGN U160 ( .B(R[160]), .A(L[160]));
Q_ASSIGN U161 ( .B(R[161]), .A(L[161]));
Q_ASSIGN U162 ( .B(R[162]), .A(L[162]));
Q_ASSIGN U163 ( .B(R[163]), .A(L[163]));
Q_ASSIGN U164 ( .B(R[164]), .A(L[164]));
Q_ASSIGN U165 ( .B(R[165]), .A(L[165]));
Q_ASSIGN U166 ( .B(R[166]), .A(L[166]));
Q_ASSIGN U167 ( .B(R[167]), .A(L[167]));
Q_ASSIGN U168 ( .B(R[168]), .A(L[168]));
Q_ASSIGN U169 ( .B(R[169]), .A(L[169]));
Q_ASSIGN U170 ( .B(R[170]), .A(L[170]));
Q_ASSIGN U171 ( .B(R[171]), .A(L[171]));
Q_ASSIGN U172 ( .B(R[172]), .A(L[172]));
Q_ASSIGN U173 ( .B(R[173]), .A(L[173]));
Q_ASSIGN U174 ( .B(R[174]), .A(L[174]));
Q_ASSIGN U175 ( .B(R[175]), .A(L[175]));
Q_ASSIGN U176 ( .B(R[176]), .A(L[176]));
Q_ASSIGN U177 ( .B(R[177]), .A(L[177]));
Q_ASSIGN U178 ( .B(R[178]), .A(L[178]));
Q_ASSIGN U179 ( .B(R[179]), .A(L[179]));
Q_ASSIGN U180 ( .B(R[180]), .A(L[180]));
Q_ASSIGN U181 ( .B(R[181]), .A(L[181]));
Q_ASSIGN U182 ( .B(R[182]), .A(L[182]));
Q_ASSIGN U183 ( .B(R[183]), .A(L[183]));
Q_ASSIGN U184 ( .B(R[184]), .A(L[184]));
Q_ASSIGN U185 ( .B(R[185]), .A(L[185]));
Q_ASSIGN U186 ( .B(R[186]), .A(L[186]));
Q_ASSIGN U187 ( .B(R[187]), .A(L[187]));
Q_ASSIGN U188 ( .B(R[188]), .A(L[188]));
Q_ASSIGN U189 ( .B(R[189]), .A(L[189]));
Q_ASSIGN U190 ( .B(R[190]), .A(L[190]));
Q_ASSIGN U191 ( .B(R[191]), .A(L[191]));
Q_ASSIGN U192 ( .B(R[192]), .A(L[192]));
Q_ASSIGN U193 ( .B(R[193]), .A(L[193]));
Q_ASSIGN U194 ( .B(R[194]), .A(L[194]));
Q_ASSIGN U195 ( .B(R[195]), .A(L[195]));
Q_ASSIGN U196 ( .B(R[196]), .A(L[196]));
Q_ASSIGN U197 ( .B(R[197]), .A(L[197]));
Q_ASSIGN U198 ( .B(R[198]), .A(L[198]));
Q_ASSIGN U199 ( .B(R[199]), .A(L[199]));
Q_ASSIGN U200 ( .B(R[200]), .A(L[200]));
Q_ASSIGN U201 ( .B(R[201]), .A(L[201]));
Q_ASSIGN U202 ( .B(R[202]), .A(L[202]));
Q_ASSIGN U203 ( .B(R[203]), .A(L[203]));
Q_ASSIGN U204 ( .B(R[204]), .A(L[204]));
Q_ASSIGN U205 ( .B(R[205]), .A(L[205]));
Q_ASSIGN U206 ( .B(R[206]), .A(L[206]));
Q_ASSIGN U207 ( .B(R[207]), .A(L[207]));
Q_ASSIGN U208 ( .B(R[208]), .A(L[208]));
Q_ASSIGN U209 ( .B(R[209]), .A(L[209]));
Q_ASSIGN U210 ( .B(R[210]), .A(L[210]));
Q_ASSIGN U211 ( .B(R[211]), .A(L[211]));
Q_ASSIGN U212 ( .B(R[212]), .A(L[212]));
Q_ASSIGN U213 ( .B(R[213]), .A(L[213]));
Q_ASSIGN U214 ( .B(R[214]), .A(L[214]));
Q_ASSIGN U215 ( .B(R[215]), .A(L[215]));
Q_ASSIGN U216 ( .B(R[216]), .A(L[216]));
Q_ASSIGN U217 ( .B(R[217]), .A(L[217]));
Q_ASSIGN U218 ( .B(R[218]), .A(L[218]));
Q_ASSIGN U219 ( .B(R[219]), .A(L[219]));
Q_ASSIGN U220 ( .B(R[220]), .A(L[220]));
Q_ASSIGN U221 ( .B(R[221]), .A(L[221]));
Q_ASSIGN U222 ( .B(R[222]), .A(L[222]));
Q_ASSIGN U223 ( .B(R[223]), .A(L[223]));
Q_ASSIGN U224 ( .B(R[224]), .A(L[224]));
Q_ASSIGN U225 ( .B(R[225]), .A(L[225]));
Q_ASSIGN U226 ( .B(R[226]), .A(L[226]));
Q_ASSIGN U227 ( .B(R[227]), .A(L[227]));
Q_ASSIGN U228 ( .B(R[228]), .A(L[228]));
Q_ASSIGN U229 ( .B(R[229]), .A(L[229]));
Q_ASSIGN U230 ( .B(R[230]), .A(L[230]));
Q_ASSIGN U231 ( .B(R[231]), .A(L[231]));
Q_ASSIGN U232 ( .B(R[232]), .A(L[232]));
Q_ASSIGN U233 ( .B(R[233]), .A(L[233]));
Q_ASSIGN U234 ( .B(R[234]), .A(L[234]));
Q_ASSIGN U235 ( .B(R[235]), .A(L[235]));
Q_ASSIGN U236 ( .B(R[236]), .A(L[236]));
Q_ASSIGN U237 ( .B(R[237]), .A(L[237]));
Q_ASSIGN U238 ( .B(R[238]), .A(L[238]));
Q_ASSIGN U239 ( .B(R[239]), .A(L[239]));
Q_ASSIGN U240 ( .B(R[240]), .A(L[240]));
Q_ASSIGN U241 ( .B(R[241]), .A(L[241]));
Q_ASSIGN U242 ( .B(R[242]), .A(L[242]));
Q_ASSIGN U243 ( .B(R[243]), .A(L[243]));
Q_ASSIGN U244 ( .B(R[244]), .A(L[244]));
Q_ASSIGN U245 ( .B(R[245]), .A(L[245]));
Q_ASSIGN U246 ( .B(R[246]), .A(L[246]));
Q_ASSIGN U247 ( .B(R[247]), .A(L[247]));
Q_ASSIGN U248 ( .B(R[248]), .A(L[248]));
Q_ASSIGN U249 ( .B(R[249]), .A(L[249]));
Q_ASSIGN U250 ( .B(R[250]), .A(L[250]));
Q_ASSIGN U251 ( .B(R[251]), .A(L[251]));
Q_ASSIGN U252 ( .B(R[252]), .A(L[252]));
Q_ASSIGN U253 ( .B(R[253]), .A(L[253]));
Q_ASSIGN U254 ( .B(R[254]), .A(L[254]));
Q_ASSIGN U255 ( .B(R[255]), .A(L[255]));
Q_ASSIGN U256 ( .B(R[256]), .A(L[256]));
Q_ASSIGN U257 ( .B(R[257]), .A(L[257]));
Q_ASSIGN U258 ( .B(R[258]), .A(L[258]));
Q_ASSIGN U259 ( .B(R[259]), .A(L[259]));
Q_ASSIGN U260 ( .B(R[260]), .A(L[260]));
Q_ASSIGN U261 ( .B(R[261]), .A(L[261]));
Q_ASSIGN U262 ( .B(R[262]), .A(L[262]));
Q_ASSIGN U263 ( .B(R[263]), .A(L[263]));
Q_ASSIGN U264 ( .B(R[264]), .A(L[264]));
Q_ASSIGN U265 ( .B(R[265]), .A(L[265]));
Q_ASSIGN U266 ( .B(R[266]), .A(L[266]));
Q_ASSIGN U267 ( .B(R[267]), .A(L[267]));
Q_ASSIGN U268 ( .B(R[268]), .A(L[268]));
Q_ASSIGN U269 ( .B(R[269]), .A(L[269]));
Q_ASSIGN U270 ( .B(R[270]), .A(L[270]));
Q_ASSIGN U271 ( .B(R[271]), .A(L[271]));
Q_ASSIGN U272 ( .B(R[272]), .A(L[272]));
Q_ASSIGN U273 ( .B(R[273]), .A(L[273]));
Q_ASSIGN U274 ( .B(R[274]), .A(L[274]));
Q_ASSIGN U275 ( .B(R[275]), .A(L[275]));
Q_ASSIGN U276 ( .B(R[276]), .A(L[276]));
Q_ASSIGN U277 ( .B(R[277]), .A(L[277]));
Q_ASSIGN U278 ( .B(R[278]), .A(L[278]));
Q_ASSIGN U279 ( .B(R[279]), .A(L[279]));
Q_ASSIGN U280 ( .B(R[280]), .A(L[280]));
Q_ASSIGN U281 ( .B(R[281]), .A(L[281]));
Q_ASSIGN U282 ( .B(R[282]), .A(L[282]));
Q_ASSIGN U283 ( .B(R[283]), .A(L[283]));
Q_ASSIGN U284 ( .B(R[284]), .A(L[284]));
Q_ASSIGN U285 ( .B(R[285]), .A(L[285]));
Q_ASSIGN U286 ( .B(R[286]), .A(L[286]));
Q_ASSIGN U287 ( .B(R[287]), .A(L[287]));
Q_ASSIGN U288 ( .B(R[288]), .A(L[288]));
Q_ASSIGN U289 ( .B(R[289]), .A(L[289]));
Q_ASSIGN U290 ( .B(R[290]), .A(L[290]));
Q_ASSIGN U291 ( .B(R[291]), .A(L[291]));
Q_ASSIGN U292 ( .B(R[292]), .A(L[292]));
Q_ASSIGN U293 ( .B(R[293]), .A(L[293]));
Q_ASSIGN U294 ( .B(R[294]), .A(L[294]));
Q_ASSIGN U295 ( .B(R[295]), .A(L[295]));
Q_ASSIGN U296 ( .B(R[296]), .A(L[296]));
Q_ASSIGN U297 ( .B(R[297]), .A(L[297]));
Q_ASSIGN U298 ( .B(R[298]), .A(L[298]));
Q_ASSIGN U299 ( .B(R[299]), .A(L[299]));
Q_ASSIGN U300 ( .B(R[300]), .A(L[300]));
Q_ASSIGN U301 ( .B(R[301]), .A(L[301]));
Q_ASSIGN U302 ( .B(R[302]), .A(L[302]));
Q_ASSIGN U303 ( .B(R[303]), .A(L[303]));
Q_ASSIGN U304 ( .B(R[304]), .A(L[304]));
Q_ASSIGN U305 ( .B(R[305]), .A(L[305]));
Q_ASSIGN U306 ( .B(R[306]), .A(L[306]));
Q_ASSIGN U307 ( .B(R[307]), .A(L[307]));
Q_ASSIGN U308 ( .B(R[308]), .A(L[308]));
Q_ASSIGN U309 ( .B(R[309]), .A(L[309]));
Q_ASSIGN U310 ( .B(R[310]), .A(L[310]));
Q_ASSIGN U311 ( .B(R[311]), .A(L[311]));
Q_ASSIGN U312 ( .B(R[312]), .A(L[312]));
Q_ASSIGN U313 ( .B(R[313]), .A(L[313]));
Q_ASSIGN U314 ( .B(R[314]), .A(L[314]));
Q_ASSIGN U315 ( .B(R[315]), .A(L[315]));
Q_ASSIGN U316 ( .B(R[316]), .A(L[316]));
Q_ASSIGN U317 ( .B(R[317]), .A(L[317]));
Q_ASSIGN U318 ( .B(R[318]), .A(L[318]));
Q_ASSIGN U319 ( .B(R[319]), .A(L[319]));
Q_ASSIGN U320 ( .B(R[320]), .A(L[320]));
Q_ASSIGN U321 ( .B(R[321]), .A(L[321]));
Q_ASSIGN U322 ( .B(R[322]), .A(L[322]));
Q_ASSIGN U323 ( .B(R[323]), .A(L[323]));
Q_ASSIGN U324 ( .B(R[324]), .A(L[324]));
Q_ASSIGN U325 ( .B(R[325]), .A(L[325]));
Q_ASSIGN U326 ( .B(R[326]), .A(L[326]));
Q_ASSIGN U327 ( .B(R[327]), .A(L[327]));
Q_ASSIGN U328 ( .B(R[328]), .A(L[328]));
Q_ASSIGN U329 ( .B(R[329]), .A(L[329]));
Q_ASSIGN U330 ( .B(R[330]), .A(L[330]));
Q_ASSIGN U331 ( .B(R[331]), .A(L[331]));
Q_ASSIGN U332 ( .B(R[332]), .A(L[332]));
Q_ASSIGN U333 ( .B(R[333]), .A(L[333]));
Q_ASSIGN U334 ( .B(R[334]), .A(L[334]));
Q_ASSIGN U335 ( .B(R[335]), .A(L[335]));
Q_ASSIGN U336 ( .B(R[336]), .A(L[336]));
Q_ASSIGN U337 ( .B(R[337]), .A(L[337]));
Q_ASSIGN U338 ( .B(R[338]), .A(L[338]));
Q_ASSIGN U339 ( .B(R[339]), .A(L[339]));
Q_ASSIGN U340 ( .B(R[340]), .A(L[340]));
Q_ASSIGN U341 ( .B(R[341]), .A(L[341]));
Q_ASSIGN U342 ( .B(R[342]), .A(L[342]));
Q_ASSIGN U343 ( .B(R[343]), .A(L[343]));
Q_ASSIGN U344 ( .B(R[344]), .A(L[344]));
Q_ASSIGN U345 ( .B(R[345]), .A(L[345]));
Q_ASSIGN U346 ( .B(R[346]), .A(L[346]));
Q_ASSIGN U347 ( .B(R[347]), .A(L[347]));
Q_ASSIGN U348 ( .B(R[348]), .A(L[348]));
Q_ASSIGN U349 ( .B(R[349]), .A(L[349]));
Q_ASSIGN U350 ( .B(R[350]), .A(L[350]));
Q_ASSIGN U351 ( .B(R[351]), .A(L[351]));
Q_ASSIGN U352 ( .B(R[352]), .A(L[352]));
Q_ASSIGN U353 ( .B(R[353]), .A(L[353]));
Q_ASSIGN U354 ( .B(R[354]), .A(L[354]));
Q_ASSIGN U355 ( .B(R[355]), .A(L[355]));
Q_ASSIGN U356 ( .B(R[356]), .A(L[356]));
Q_ASSIGN U357 ( .B(R[357]), .A(L[357]));
Q_ASSIGN U358 ( .B(R[358]), .A(L[358]));
Q_ASSIGN U359 ( .B(R[359]), .A(L[359]));
Q_ASSIGN U360 ( .B(R[360]), .A(L[360]));
Q_ASSIGN U361 ( .B(R[361]), .A(L[361]));
Q_ASSIGN U362 ( .B(R[362]), .A(L[362]));
Q_ASSIGN U363 ( .B(R[363]), .A(L[363]));
Q_ASSIGN U364 ( .B(R[364]), .A(L[364]));
Q_ASSIGN U365 ( .B(R[365]), .A(L[365]));
Q_ASSIGN U366 ( .B(R[366]), .A(L[366]));
Q_ASSIGN U367 ( .B(R[367]), .A(L[367]));
Q_ASSIGN U368 ( .B(R[368]), .A(L[368]));
Q_ASSIGN U369 ( .B(R[369]), .A(L[369]));
Q_ASSIGN U370 ( .B(R[370]), .A(L[370]));
Q_ASSIGN U371 ( .B(R[371]), .A(L[371]));
Q_ASSIGN U372 ( .B(R[372]), .A(L[372]));
Q_ASSIGN U373 ( .B(R[373]), .A(L[373]));
Q_ASSIGN U374 ( .B(R[374]), .A(L[374]));
Q_ASSIGN U375 ( .B(R[375]), .A(L[375]));
Q_ASSIGN U376 ( .B(R[376]), .A(L[376]));
Q_ASSIGN U377 ( .B(R[377]), .A(L[377]));
Q_ASSIGN U378 ( .B(R[378]), .A(L[378]));
Q_ASSIGN U379 ( .B(R[379]), .A(L[379]));
Q_ASSIGN U380 ( .B(R[380]), .A(L[380]));
Q_ASSIGN U381 ( .B(R[381]), .A(L[381]));
Q_ASSIGN U382 ( .B(R[382]), .A(L[382]));
Q_ASSIGN U383 ( .B(R[383]), .A(L[383]));
Q_ASSIGN U384 ( .B(R[384]), .A(L[384]));
Q_ASSIGN U385 ( .B(R[385]), .A(L[385]));
Q_ASSIGN U386 ( .B(R[386]), .A(L[386]));
Q_ASSIGN U387 ( .B(R[387]), .A(L[387]));
Q_ASSIGN U388 ( .B(R[388]), .A(L[388]));
Q_ASSIGN U389 ( .B(R[389]), .A(L[389]));
Q_ASSIGN U390 ( .B(R[390]), .A(L[390]));
Q_ASSIGN U391 ( .B(R[391]), .A(L[391]));
Q_ASSIGN U392 ( .B(R[392]), .A(L[392]));
Q_ASSIGN U393 ( .B(R[393]), .A(L[393]));
Q_ASSIGN U394 ( .B(R[394]), .A(L[394]));
Q_ASSIGN U395 ( .B(R[395]), .A(L[395]));
Q_ASSIGN U396 ( .B(R[396]), .A(L[396]));
Q_ASSIGN U397 ( .B(R[397]), .A(L[397]));
Q_ASSIGN U398 ( .B(R[398]), .A(L[398]));
Q_ASSIGN U399 ( .B(R[399]), .A(L[399]));
Q_ASSIGN U400 ( .B(R[400]), .A(L[400]));
Q_ASSIGN U401 ( .B(R[401]), .A(L[401]));
Q_ASSIGN U402 ( .B(R[402]), .A(L[402]));
Q_ASSIGN U403 ( .B(R[403]), .A(L[403]));
Q_ASSIGN U404 ( .B(R[404]), .A(L[404]));
Q_ASSIGN U405 ( .B(R[405]), .A(L[405]));
Q_ASSIGN U406 ( .B(R[406]), .A(L[406]));
Q_ASSIGN U407 ( .B(R[407]), .A(L[407]));
Q_ASSIGN U408 ( .B(R[408]), .A(L[408]));
Q_ASSIGN U409 ( .B(R[409]), .A(L[409]));
Q_ASSIGN U410 ( .B(R[410]), .A(L[410]));
Q_ASSIGN U411 ( .B(R[411]), .A(L[411]));
Q_ASSIGN U412 ( .B(R[412]), .A(L[412]));
Q_ASSIGN U413 ( .B(R[413]), .A(L[413]));
Q_ASSIGN U414 ( .B(R[414]), .A(L[414]));
Q_ASSIGN U415 ( .B(R[415]), .A(L[415]));
Q_ASSIGN U416 ( .B(R[416]), .A(L[416]));
Q_ASSIGN U417 ( .B(R[417]), .A(L[417]));
Q_ASSIGN U418 ( .B(R[418]), .A(L[418]));
Q_ASSIGN U419 ( .B(R[419]), .A(L[419]));
Q_ASSIGN U420 ( .B(R[420]), .A(L[420]));
Q_ASSIGN U421 ( .B(R[421]), .A(L[421]));
Q_ASSIGN U422 ( .B(R[422]), .A(L[422]));
Q_ASSIGN U423 ( .B(R[423]), .A(L[423]));
Q_ASSIGN U424 ( .B(R[424]), .A(L[424]));
Q_ASSIGN U425 ( .B(R[425]), .A(L[425]));
Q_ASSIGN U426 ( .B(R[426]), .A(L[426]));
Q_ASSIGN U427 ( .B(R[427]), .A(L[427]));
Q_ASSIGN U428 ( .B(R[428]), .A(L[428]));
Q_ASSIGN U429 ( .B(R[429]), .A(L[429]));
Q_ASSIGN U430 ( .B(R[430]), .A(L[430]));
Q_ASSIGN U431 ( .B(R[431]), .A(L[431]));
Q_ASSIGN U432 ( .B(R[432]), .A(L[432]));
Q_ASSIGN U433 ( .B(R[433]), .A(L[433]));
Q_ASSIGN U434 ( .B(R[434]), .A(L[434]));
Q_ASSIGN U435 ( .B(R[435]), .A(L[435]));
Q_ASSIGN U436 ( .B(R[436]), .A(L[436]));
Q_ASSIGN U437 ( .B(R[437]), .A(L[437]));
Q_ASSIGN U438 ( .B(R[438]), .A(L[438]));
Q_ASSIGN U439 ( .B(R[439]), .A(L[439]));
Q_ASSIGN U440 ( .B(R[440]), .A(L[440]));
Q_ASSIGN U441 ( .B(R[441]), .A(L[441]));
Q_ASSIGN U442 ( .B(R[442]), .A(L[442]));
Q_ASSIGN U443 ( .B(R[443]), .A(L[443]));
Q_ASSIGN U444 ( .B(R[444]), .A(L[444]));
Q_ASSIGN U445 ( .B(R[445]), .A(L[445]));
Q_ASSIGN U446 ( .B(R[446]), .A(L[446]));
Q_ASSIGN U447 ( .B(R[447]), .A(L[447]));
Q_ASSIGN U448 ( .B(R[448]), .A(L[448]));
Q_ASSIGN U449 ( .B(R[449]), .A(L[449]));
Q_ASSIGN U450 ( .B(R[450]), .A(L[450]));
Q_ASSIGN U451 ( .B(R[451]), .A(L[451]));
Q_ASSIGN U452 ( .B(R[452]), .A(L[452]));
Q_ASSIGN U453 ( .B(R[453]), .A(L[453]));
Q_ASSIGN U454 ( .B(R[454]), .A(L[454]));
Q_ASSIGN U455 ( .B(R[455]), .A(L[455]));
Q_ASSIGN U456 ( .B(R[456]), .A(L[456]));
Q_ASSIGN U457 ( .B(R[457]), .A(L[457]));
Q_ASSIGN U458 ( .B(R[458]), .A(L[458]));
Q_ASSIGN U459 ( .B(R[459]), .A(L[459]));
Q_ASSIGN U460 ( .B(R[460]), .A(L[460]));
Q_ASSIGN U461 ( .B(R[461]), .A(L[461]));
Q_ASSIGN U462 ( .B(R[462]), .A(L[462]));
Q_ASSIGN U463 ( .B(R[463]), .A(L[463]));
Q_ASSIGN U464 ( .B(R[464]), .A(L[464]));
Q_ASSIGN U465 ( .B(R[465]), .A(L[465]));
Q_ASSIGN U466 ( .B(R[466]), .A(L[466]));
Q_ASSIGN U467 ( .B(R[467]), .A(L[467]));
Q_ASSIGN U468 ( .B(R[468]), .A(L[468]));
Q_ASSIGN U469 ( .B(R[469]), .A(L[469]));
Q_ASSIGN U470 ( .B(R[470]), .A(L[470]));
Q_ASSIGN U471 ( .B(R[471]), .A(L[471]));
Q_ASSIGN U472 ( .B(R[472]), .A(L[472]));
Q_ASSIGN U473 ( .B(R[473]), .A(L[473]));
Q_ASSIGN U474 ( .B(R[474]), .A(L[474]));
Q_ASSIGN U475 ( .B(R[475]), .A(L[475]));
Q_ASSIGN U476 ( .B(R[476]), .A(L[476]));
Q_ASSIGN U477 ( .B(R[477]), .A(L[477]));
Q_ASSIGN U478 ( .B(R[478]), .A(L[478]));
Q_ASSIGN U479 ( .B(R[479]), .A(L[479]));
Q_ASSIGN U480 ( .B(R[480]), .A(L[480]));
Q_ASSIGN U481 ( .B(R[481]), .A(L[481]));
Q_ASSIGN U482 ( .B(R[482]), .A(L[482]));
Q_ASSIGN U483 ( .B(R[483]), .A(L[483]));
Q_ASSIGN U484 ( .B(R[484]), .A(L[484]));
Q_ASSIGN U485 ( .B(R[485]), .A(L[485]));
Q_ASSIGN U486 ( .B(R[486]), .A(L[486]));
Q_ASSIGN U487 ( .B(R[487]), .A(L[487]));
Q_ASSIGN U488 ( .B(R[488]), .A(L[488]));
Q_ASSIGN U489 ( .B(R[489]), .A(L[489]));
Q_ASSIGN U490 ( .B(R[490]), .A(L[490]));
Q_ASSIGN U491 ( .B(R[491]), .A(L[491]));
Q_ASSIGN U492 ( .B(R[492]), .A(L[492]));
Q_ASSIGN U493 ( .B(R[493]), .A(L[493]));
Q_ASSIGN U494 ( .B(R[494]), .A(L[494]));
Q_ASSIGN U495 ( .B(R[495]), .A(L[495]));
Q_ASSIGN U496 ( .B(R[496]), .A(L[496]));
Q_ASSIGN U497 ( .B(R[497]), .A(L[497]));
Q_ASSIGN U498 ( .B(R[498]), .A(L[498]));
Q_ASSIGN U499 ( .B(R[499]), .A(L[499]));
Q_ASSIGN U500 ( .B(R[500]), .A(L[500]));
Q_ASSIGN U501 ( .B(R[501]), .A(L[501]));
Q_ASSIGN U502 ( .B(R[502]), .A(L[502]));
Q_ASSIGN U503 ( .B(R[503]), .A(L[503]));
Q_ASSIGN U504 ( .B(R[504]), .A(L[504]));
Q_ASSIGN U505 ( .B(R[505]), .A(L[505]));
Q_ASSIGN U506 ( .B(R[506]), .A(L[506]));
Q_ASSIGN U507 ( .B(R[507]), .A(L[507]));
Q_ASSIGN U508 ( .B(R[508]), .A(L[508]));
Q_ASSIGN U509 ( .B(R[509]), .A(L[509]));
Q_ASSIGN U510 ( .B(R[510]), .A(L[510]));
Q_ASSIGN U511 ( .B(R[511]), .A(L[511]));
Q_ASSIGN U512 ( .B(R[512]), .A(L[512]));
Q_ASSIGN U513 ( .B(R[513]), .A(L[513]));
Q_ASSIGN U514 ( .B(R[514]), .A(L[514]));
Q_ASSIGN U515 ( .B(R[515]), .A(L[515]));
Q_ASSIGN U516 ( .B(R[516]), .A(L[516]));
Q_ASSIGN U517 ( .B(R[517]), .A(L[517]));
Q_ASSIGN U518 ( .B(R[518]), .A(L[518]));
Q_ASSIGN U519 ( .B(R[519]), .A(L[519]));
Q_ASSIGN U520 ( .B(R[520]), .A(L[520]));
Q_ASSIGN U521 ( .B(R[521]), .A(L[521]));
Q_ASSIGN U522 ( .B(R[522]), .A(L[522]));
Q_ASSIGN U523 ( .B(R[523]), .A(L[523]));
Q_ASSIGN U524 ( .B(R[524]), .A(L[524]));
Q_ASSIGN U525 ( .B(R[525]), .A(L[525]));
Q_ASSIGN U526 ( .B(R[526]), .A(L[526]));
Q_ASSIGN U527 ( .B(R[527]), .A(L[527]));
Q_ASSIGN U528 ( .B(R[528]), .A(L[528]));
Q_ASSIGN U529 ( .B(R[529]), .A(L[529]));
Q_ASSIGN U530 ( .B(R[530]), .A(L[530]));
Q_ASSIGN U531 ( .B(R[531]), .A(L[531]));
Q_ASSIGN U532 ( .B(R[532]), .A(L[532]));
Q_ASSIGN U533 ( .B(R[533]), .A(L[533]));
Q_ASSIGN U534 ( .B(R[534]), .A(L[534]));
Q_ASSIGN U535 ( .B(R[535]), .A(L[535]));
Q_ASSIGN U536 ( .B(R[536]), .A(L[536]));
Q_ASSIGN U537 ( .B(R[537]), .A(L[537]));
Q_ASSIGN U538 ( .B(R[538]), .A(L[538]));
Q_ASSIGN U539 ( .B(R[539]), .A(L[539]));
Q_ASSIGN U540 ( .B(R[540]), .A(L[540]));
Q_ASSIGN U541 ( .B(R[541]), .A(L[541]));
Q_ASSIGN U542 ( .B(R[542]), .A(L[542]));
Q_ASSIGN U543 ( .B(R[543]), .A(L[543]));
Q_ASSIGN U544 ( .B(R[544]), .A(L[544]));
Q_ASSIGN U545 ( .B(R[545]), .A(L[545]));
Q_ASSIGN U546 ( .B(R[546]), .A(L[546]));
Q_ASSIGN U547 ( .B(R[547]), .A(L[547]));
Q_ASSIGN U548 ( .B(R[548]), .A(L[548]));
Q_ASSIGN U549 ( .B(R[549]), .A(L[549]));
Q_ASSIGN U550 ( .B(R[550]), .A(L[550]));
Q_ASSIGN U551 ( .B(R[551]), .A(L[551]));
Q_ASSIGN U552 ( .B(R[552]), .A(L[552]));
Q_ASSIGN U553 ( .B(R[553]), .A(L[553]));
Q_ASSIGN U554 ( .B(R[554]), .A(L[554]));
Q_ASSIGN U555 ( .B(R[555]), .A(L[555]));
Q_ASSIGN U556 ( .B(R[556]), .A(L[556]));
Q_ASSIGN U557 ( .B(R[557]), .A(L[557]));
Q_ASSIGN U558 ( .B(R[558]), .A(L[558]));
Q_ASSIGN U559 ( .B(R[559]), .A(L[559]));
Q_ASSIGN U560 ( .B(R[560]), .A(L[560]));
Q_ASSIGN U561 ( .B(R[561]), .A(L[561]));
Q_ASSIGN U562 ( .B(R[562]), .A(L[562]));
Q_ASSIGN U563 ( .B(R[563]), .A(L[563]));
Q_ASSIGN U564 ( .B(R[564]), .A(L[564]));
Q_ASSIGN U565 ( .B(R[565]), .A(L[565]));
Q_ASSIGN U566 ( .B(R[566]), .A(L[566]));
Q_ASSIGN U567 ( .B(R[567]), .A(L[567]));
Q_ASSIGN U568 ( .B(R[568]), .A(L[568]));
Q_ASSIGN U569 ( .B(R[569]), .A(L[569]));
Q_ASSIGN U570 ( .B(R[570]), .A(L[570]));
Q_ASSIGN U571 ( .B(R[571]), .A(L[571]));
Q_ASSIGN U572 ( .B(R[572]), .A(L[572]));
Q_ASSIGN U573 ( .B(R[573]), .A(L[573]));
Q_ASSIGN U574 ( .B(R[574]), .A(L[574]));
Q_ASSIGN U575 ( .B(R[575]), .A(L[575]));
Q_ASSIGN U576 ( .B(R[576]), .A(L[576]));
Q_ASSIGN U577 ( .B(R[577]), .A(L[577]));
Q_ASSIGN U578 ( .B(R[578]), .A(L[578]));
Q_ASSIGN U579 ( .B(R[579]), .A(L[579]));
Q_ASSIGN U580 ( .B(R[580]), .A(L[580]));
Q_ASSIGN U581 ( .B(R[581]), .A(L[581]));
Q_ASSIGN U582 ( .B(R[582]), .A(L[582]));
Q_ASSIGN U583 ( .B(R[583]), .A(L[583]));
Q_ASSIGN U584 ( .B(R[584]), .A(L[584]));
Q_ASSIGN U585 ( .B(R[585]), .A(L[585]));
Q_ASSIGN U586 ( .B(R[586]), .A(L[586]));
Q_ASSIGN U587 ( .B(R[587]), .A(L[587]));
Q_ASSIGN U588 ( .B(R[588]), .A(L[588]));
Q_ASSIGN U589 ( .B(R[589]), .A(L[589]));
Q_ASSIGN U590 ( .B(R[590]), .A(L[590]));
Q_ASSIGN U591 ( .B(R[591]), .A(L[591]));
Q_ASSIGN U592 ( .B(R[592]), .A(L[592]));
Q_ASSIGN U593 ( .B(R[593]), .A(L[593]));
Q_ASSIGN U594 ( .B(R[594]), .A(L[594]));
Q_ASSIGN U595 ( .B(R[595]), .A(L[595]));
Q_ASSIGN U596 ( .B(R[596]), .A(L[596]));
Q_ASSIGN U597 ( .B(R[597]), .A(L[597]));
Q_ASSIGN U598 ( .B(R[598]), .A(L[598]));
Q_ASSIGN U599 ( .B(R[599]), .A(L[599]));
Q_ASSIGN U600 ( .B(R[600]), .A(L[600]));
Q_ASSIGN U601 ( .B(R[601]), .A(L[601]));
Q_ASSIGN U602 ( .B(R[602]), .A(L[602]));
Q_ASSIGN U603 ( .B(R[603]), .A(L[603]));
Q_ASSIGN U604 ( .B(R[604]), .A(L[604]));
Q_ASSIGN U605 ( .B(R[605]), .A(L[605]));
Q_ASSIGN U606 ( .B(R[606]), .A(L[606]));
Q_ASSIGN U607 ( .B(R[607]), .A(L[607]));
Q_ASSIGN U608 ( .B(R[608]), .A(L[608]));
Q_ASSIGN U609 ( .B(R[609]), .A(L[609]));
Q_ASSIGN U610 ( .B(R[610]), .A(L[610]));
Q_ASSIGN U611 ( .B(R[611]), .A(L[611]));
Q_ASSIGN U612 ( .B(R[612]), .A(L[612]));
Q_ASSIGN U613 ( .B(R[613]), .A(L[613]));
Q_ASSIGN U614 ( .B(R[614]), .A(L[614]));
Q_ASSIGN U615 ( .B(R[615]), .A(L[615]));
Q_ASSIGN U616 ( .B(R[616]), .A(L[616]));
Q_ASSIGN U617 ( .B(R[617]), .A(L[617]));
Q_ASSIGN U618 ( .B(R[618]), .A(L[618]));
Q_ASSIGN U619 ( .B(R[619]), .A(L[619]));
Q_ASSIGN U620 ( .B(R[620]), .A(L[620]));
Q_ASSIGN U621 ( .B(R[621]), .A(L[621]));
Q_ASSIGN U622 ( .B(R[622]), .A(L[622]));
Q_ASSIGN U623 ( .B(R[623]), .A(L[623]));
Q_ASSIGN U624 ( .B(R[624]), .A(L[624]));
Q_ASSIGN U625 ( .B(R[625]), .A(L[625]));
Q_ASSIGN U626 ( .B(R[626]), .A(L[626]));
Q_ASSIGN U627 ( .B(R[627]), .A(L[627]));
Q_ASSIGN U628 ( .B(R[628]), .A(L[628]));
Q_ASSIGN U629 ( .B(R[629]), .A(L[629]));
Q_ASSIGN U630 ( .B(R[630]), .A(L[630]));
Q_ASSIGN U631 ( .B(R[631]), .A(L[631]));
Q_ASSIGN U632 ( .B(R[632]), .A(L[632]));
Q_ASSIGN U633 ( .B(R[633]), .A(L[633]));
Q_ASSIGN U634 ( .B(R[634]), .A(L[634]));
Q_ASSIGN U635 ( .B(R[635]), .A(L[635]));
Q_ASSIGN U636 ( .B(R[636]), .A(L[636]));
Q_ASSIGN U637 ( .B(R[637]), .A(L[637]));
Q_ASSIGN U638 ( .B(R[638]), .A(L[638]));
Q_ASSIGN U639 ( .B(R[639]), .A(L[639]));
Q_ASSIGN U640 ( .B(R[640]), .A(L[640]));
Q_ASSIGN U641 ( .B(R[641]), .A(L[641]));
Q_ASSIGN U642 ( .B(R[642]), .A(L[642]));
Q_ASSIGN U643 ( .B(R[643]), .A(L[643]));
Q_ASSIGN U644 ( .B(R[644]), .A(L[644]));
Q_ASSIGN U645 ( .B(R[645]), .A(L[645]));
Q_ASSIGN U646 ( .B(R[646]), .A(L[646]));
Q_ASSIGN U647 ( .B(R[647]), .A(L[647]));
Q_ASSIGN U648 ( .B(R[648]), .A(L[648]));
Q_ASSIGN U649 ( .B(R[649]), .A(L[649]));
Q_ASSIGN U650 ( .B(R[650]), .A(L[650]));
Q_ASSIGN U651 ( .B(R[651]), .A(L[651]));
Q_ASSIGN U652 ( .B(R[652]), .A(L[652]));
Q_ASSIGN U653 ( .B(R[653]), .A(L[653]));
Q_ASSIGN U654 ( .B(R[654]), .A(L[654]));
Q_ASSIGN U655 ( .B(R[655]), .A(L[655]));
Q_ASSIGN U656 ( .B(R[656]), .A(L[656]));
Q_ASSIGN U657 ( .B(R[657]), .A(L[657]));
Q_ASSIGN U658 ( .B(R[658]), .A(L[658]));
Q_ASSIGN U659 ( .B(R[659]), .A(L[659]));
Q_ASSIGN U660 ( .B(R[660]), .A(L[660]));
Q_ASSIGN U661 ( .B(R[661]), .A(L[661]));
Q_ASSIGN U662 ( .B(R[662]), .A(L[662]));
Q_ASSIGN U663 ( .B(R[663]), .A(L[663]));
Q_ASSIGN U664 ( .B(R[664]), .A(L[664]));
Q_ASSIGN U665 ( .B(R[665]), .A(L[665]));
Q_ASSIGN U666 ( .B(R[666]), .A(L[666]));
Q_ASSIGN U667 ( .B(R[667]), .A(L[667]));
Q_ASSIGN U668 ( .B(R[668]), .A(L[668]));
Q_ASSIGN U669 ( .B(R[669]), .A(L[669]));
Q_ASSIGN U670 ( .B(R[670]), .A(L[670]));
Q_ASSIGN U671 ( .B(R[671]), .A(L[671]));
Q_ASSIGN U672 ( .B(R[672]), .A(L[672]));
Q_ASSIGN U673 ( .B(R[673]), .A(L[673]));
Q_ASSIGN U674 ( .B(R[674]), .A(L[674]));
Q_ASSIGN U675 ( .B(R[675]), .A(L[675]));
Q_ASSIGN U676 ( .B(R[676]), .A(L[676]));
Q_ASSIGN U677 ( .B(R[677]), .A(L[677]));
Q_ASSIGN U678 ( .B(R[678]), .A(L[678]));
Q_ASSIGN U679 ( .B(R[679]), .A(L[679]));
Q_ASSIGN U680 ( .B(R[680]), .A(L[680]));
Q_ASSIGN U681 ( .B(R[681]), .A(L[681]));
Q_ASSIGN U682 ( .B(R[682]), .A(L[682]));
Q_ASSIGN U683 ( .B(R[683]), .A(L[683]));
Q_ASSIGN U684 ( .B(R[684]), .A(L[684]));
Q_ASSIGN U685 ( .B(R[685]), .A(L[685]));
Q_ASSIGN U686 ( .B(R[686]), .A(L[686]));
Q_ASSIGN U687 ( .B(R[687]), .A(L[687]));
Q_ASSIGN U688 ( .B(R[688]), .A(L[688]));
Q_ASSIGN U689 ( .B(R[689]), .A(L[689]));
Q_ASSIGN U690 ( .B(R[690]), .A(L[690]));
Q_ASSIGN U691 ( .B(R[691]), .A(L[691]));
Q_ASSIGN U692 ( .B(R[692]), .A(L[692]));
Q_ASSIGN U693 ( .B(R[693]), .A(L[693]));
Q_ASSIGN U694 ( .B(R[694]), .A(L[694]));
Q_ASSIGN U695 ( .B(R[695]), .A(L[695]));
Q_ASSIGN U696 ( .B(R[696]), .A(L[696]));
Q_ASSIGN U697 ( .B(R[697]), .A(L[697]));
Q_ASSIGN U698 ( .B(R[698]), .A(L[698]));
Q_ASSIGN U699 ( .B(R[699]), .A(L[699]));
Q_ASSIGN U700 ( .B(R[700]), .A(L[700]));
Q_ASSIGN U701 ( .B(R[701]), .A(L[701]));
Q_ASSIGN U702 ( .B(R[702]), .A(L[702]));
Q_ASSIGN U703 ( .B(R[703]), .A(L[703]));
Q_ASSIGN U704 ( .B(R[704]), .A(L[704]));
Q_ASSIGN U705 ( .B(R[705]), .A(L[705]));
Q_ASSIGN U706 ( .B(R[706]), .A(L[706]));
Q_ASSIGN U707 ( .B(R[707]), .A(L[707]));
Q_ASSIGN U708 ( .B(R[708]), .A(L[708]));
Q_ASSIGN U709 ( .B(R[709]), .A(L[709]));
Q_ASSIGN U710 ( .B(R[710]), .A(L[710]));
Q_ASSIGN U711 ( .B(R[711]), .A(L[711]));
Q_ASSIGN U712 ( .B(R[712]), .A(L[712]));
Q_ASSIGN U713 ( .B(R[713]), .A(L[713]));
Q_ASSIGN U714 ( .B(R[714]), .A(L[714]));
Q_ASSIGN U715 ( .B(R[715]), .A(L[715]));
Q_ASSIGN U716 ( .B(R[716]), .A(L[716]));
Q_ASSIGN U717 ( .B(R[717]), .A(L[717]));
Q_ASSIGN U718 ( .B(R[718]), .A(L[718]));
Q_ASSIGN U719 ( .B(R[719]), .A(L[719]));
Q_ASSIGN U720 ( .B(R[720]), .A(L[720]));
Q_ASSIGN U721 ( .B(R[721]), .A(L[721]));
Q_ASSIGN U722 ( .B(R[722]), .A(L[722]));
Q_ASSIGN U723 ( .B(R[723]), .A(L[723]));
Q_ASSIGN U724 ( .B(R[724]), .A(L[724]));
Q_ASSIGN U725 ( .B(R[725]), .A(L[725]));
Q_ASSIGN U726 ( .B(R[726]), .A(L[726]));
Q_ASSIGN U727 ( .B(R[727]), .A(L[727]));
Q_ASSIGN U728 ( .B(R[728]), .A(L[728]));
Q_ASSIGN U729 ( .B(R[729]), .A(L[729]));
Q_ASSIGN U730 ( .B(R[730]), .A(L[730]));
Q_ASSIGN U731 ( .B(R[731]), .A(L[731]));
Q_ASSIGN U732 ( .B(R[732]), .A(L[732]));
Q_ASSIGN U733 ( .B(R[733]), .A(L[733]));
Q_ASSIGN U734 ( .B(R[734]), .A(L[734]));
Q_ASSIGN U735 ( .B(R[735]), .A(L[735]));
Q_ASSIGN U736 ( .B(R[736]), .A(L[736]));
Q_ASSIGN U737 ( .B(R[737]), .A(L[737]));
Q_ASSIGN U738 ( .B(R[738]), .A(L[738]));
Q_ASSIGN U739 ( .B(R[739]), .A(L[739]));
Q_ASSIGN U740 ( .B(R[740]), .A(L[740]));
Q_ASSIGN U741 ( .B(R[741]), .A(L[741]));
Q_ASSIGN U742 ( .B(R[742]), .A(L[742]));
Q_ASSIGN U743 ( .B(R[743]), .A(L[743]));
Q_ASSIGN U744 ( .B(R[744]), .A(L[744]));
Q_ASSIGN U745 ( .B(R[745]), .A(L[745]));
Q_ASSIGN U746 ( .B(R[746]), .A(L[746]));
Q_ASSIGN U747 ( .B(R[747]), .A(L[747]));
Q_ASSIGN U748 ( .B(R[748]), .A(L[748]));
Q_ASSIGN U749 ( .B(R[749]), .A(L[749]));
Q_ASSIGN U750 ( .B(R[750]), .A(L[750]));
Q_ASSIGN U751 ( .B(R[751]), .A(L[751]));
Q_ASSIGN U752 ( .B(R[752]), .A(L[752]));
Q_ASSIGN U753 ( .B(R[753]), .A(L[753]));
Q_ASSIGN U754 ( .B(R[754]), .A(L[754]));
Q_ASSIGN U755 ( .B(R[755]), .A(L[755]));
Q_ASSIGN U756 ( .B(R[756]), .A(L[756]));
Q_ASSIGN U757 ( .B(R[757]), .A(L[757]));
Q_ASSIGN U758 ( .B(R[758]), .A(L[758]));
Q_ASSIGN U759 ( .B(R[759]), .A(L[759]));
Q_ASSIGN U760 ( .B(R[760]), .A(L[760]));
Q_ASSIGN U761 ( .B(R[761]), .A(L[761]));
Q_ASSIGN U762 ( .B(R[762]), .A(L[762]));
Q_ASSIGN U763 ( .B(R[763]), .A(L[763]));
Q_ASSIGN U764 ( .B(R[764]), .A(L[764]));
Q_ASSIGN U765 ( .B(R[765]), .A(L[765]));
Q_ASSIGN U766 ( .B(R[766]), .A(L[766]));
Q_ASSIGN U767 ( .B(R[767]), .A(L[767]));
Q_ASSIGN U768 ( .B(R[768]), .A(L[768]));
Q_ASSIGN U769 ( .B(R[769]), .A(L[769]));
Q_ASSIGN U770 ( .B(R[770]), .A(L[770]));
Q_ASSIGN U771 ( .B(R[771]), .A(L[771]));
Q_ASSIGN U772 ( .B(R[772]), .A(L[772]));
Q_ASSIGN U773 ( .B(R[773]), .A(L[773]));
Q_ASSIGN U774 ( .B(R[774]), .A(L[774]));
Q_ASSIGN U775 ( .B(R[775]), .A(L[775]));
Q_ASSIGN U776 ( .B(R[776]), .A(L[776]));
Q_ASSIGN U777 ( .B(R[777]), .A(L[777]));
Q_ASSIGN U778 ( .B(R[778]), .A(L[778]));
Q_ASSIGN U779 ( .B(R[779]), .A(L[779]));
Q_ASSIGN U780 ( .B(R[780]), .A(L[780]));
Q_ASSIGN U781 ( .B(R[781]), .A(L[781]));
Q_ASSIGN U782 ( .B(R[782]), .A(L[782]));
Q_ASSIGN U783 ( .B(R[783]), .A(L[783]));
Q_ASSIGN U784 ( .B(R[784]), .A(L[784]));
Q_ASSIGN U785 ( .B(R[785]), .A(L[785]));
Q_ASSIGN U786 ( .B(R[786]), .A(L[786]));
Q_ASSIGN U787 ( .B(R[787]), .A(L[787]));
Q_ASSIGN U788 ( .B(R[788]), .A(L[788]));
Q_ASSIGN U789 ( .B(R[789]), .A(L[789]));
Q_ASSIGN U790 ( .B(R[790]), .A(L[790]));
Q_ASSIGN U791 ( .B(R[791]), .A(L[791]));
Q_ASSIGN U792 ( .B(R[792]), .A(L[792]));
Q_ASSIGN U793 ( .B(R[793]), .A(L[793]));
Q_ASSIGN U794 ( .B(R[794]), .A(L[794]));
Q_ASSIGN U795 ( .B(R[795]), .A(L[795]));
Q_ASSIGN U796 ( .B(R[796]), .A(L[796]));
Q_ASSIGN U797 ( .B(R[797]), .A(L[797]));
Q_ASSIGN U798 ( .B(R[798]), .A(L[798]));
Q_ASSIGN U799 ( .B(R[799]), .A(L[799]));
Q_ASSIGN U800 ( .B(R[800]), .A(L[800]));
Q_ASSIGN U801 ( .B(R[801]), .A(L[801]));
Q_ASSIGN U802 ( .B(R[802]), .A(L[802]));
Q_ASSIGN U803 ( .B(R[803]), .A(L[803]));
Q_ASSIGN U804 ( .B(R[804]), .A(L[804]));
Q_ASSIGN U805 ( .B(R[805]), .A(L[805]));
Q_ASSIGN U806 ( .B(R[806]), .A(L[806]));
Q_ASSIGN U807 ( .B(R[807]), .A(L[807]));
Q_ASSIGN U808 ( .B(R[808]), .A(L[808]));
Q_ASSIGN U809 ( .B(R[809]), .A(L[809]));
Q_ASSIGN U810 ( .B(R[810]), .A(L[810]));
Q_ASSIGN U811 ( .B(R[811]), .A(L[811]));
Q_ASSIGN U812 ( .B(R[812]), .A(L[812]));
Q_ASSIGN U813 ( .B(R[813]), .A(L[813]));
Q_ASSIGN U814 ( .B(R[814]), .A(L[814]));
Q_ASSIGN U815 ( .B(R[815]), .A(L[815]));
Q_ASSIGN U816 ( .B(R[816]), .A(L[816]));
Q_ASSIGN U817 ( .B(R[817]), .A(L[817]));
Q_ASSIGN U818 ( .B(R[818]), .A(L[818]));
Q_ASSIGN U819 ( .B(R[819]), .A(L[819]));
Q_ASSIGN U820 ( .B(R[820]), .A(L[820]));
Q_ASSIGN U821 ( .B(R[821]), .A(L[821]));
Q_ASSIGN U822 ( .B(R[822]), .A(L[822]));
Q_ASSIGN U823 ( .B(R[823]), .A(L[823]));
Q_ASSIGN U824 ( .B(R[824]), .A(L[824]));
Q_ASSIGN U825 ( .B(R[825]), .A(L[825]));
Q_ASSIGN U826 ( .B(R[826]), .A(L[826]));
Q_ASSIGN U827 ( .B(R[827]), .A(L[827]));
Q_ASSIGN U828 ( .B(R[828]), .A(L[828]));
Q_ASSIGN U829 ( .B(R[829]), .A(L[829]));
Q_ASSIGN U830 ( .B(R[830]), .A(L[830]));
Q_ASSIGN U831 ( .B(R[831]), .A(L[831]));
Q_ASSIGN U832 ( .B(R[832]), .A(L[832]));
Q_ASSIGN U833 ( .B(R[833]), .A(L[833]));
Q_ASSIGN U834 ( .B(R[834]), .A(L[834]));
Q_ASSIGN U835 ( .B(R[835]), .A(L[835]));
Q_ASSIGN U836 ( .B(R[836]), .A(L[836]));
Q_ASSIGN U837 ( .B(R[837]), .A(L[837]));
Q_ASSIGN U838 ( .B(R[838]), .A(L[838]));
Q_ASSIGN U839 ( .B(R[839]), .A(L[839]));
Q_ASSIGN U840 ( .B(R[840]), .A(L[840]));
Q_ASSIGN U841 ( .B(R[841]), .A(L[841]));
Q_ASSIGN U842 ( .B(R[842]), .A(L[842]));
Q_ASSIGN U843 ( .B(R[843]), .A(L[843]));
Q_ASSIGN U844 ( .B(R[844]), .A(L[844]));
Q_ASSIGN U845 ( .B(R[845]), .A(L[845]));
Q_ASSIGN U846 ( .B(R[846]), .A(L[846]));
Q_ASSIGN U847 ( .B(R[847]), .A(L[847]));
Q_ASSIGN U848 ( .B(R[848]), .A(L[848]));
Q_ASSIGN U849 ( .B(R[849]), .A(L[849]));
Q_ASSIGN U850 ( .B(R[850]), .A(L[850]));
Q_ASSIGN U851 ( .B(R[851]), .A(L[851]));
Q_ASSIGN U852 ( .B(R[852]), .A(L[852]));
Q_ASSIGN U853 ( .B(R[853]), .A(L[853]));
Q_ASSIGN U854 ( .B(R[854]), .A(L[854]));
Q_ASSIGN U855 ( .B(R[855]), .A(L[855]));
Q_ASSIGN U856 ( .B(R[856]), .A(L[856]));
Q_ASSIGN U857 ( .B(R[857]), .A(L[857]));
Q_ASSIGN U858 ( .B(R[858]), .A(L[858]));
Q_ASSIGN U859 ( .B(R[859]), .A(L[859]));
Q_ASSIGN U860 ( .B(R[860]), .A(L[860]));
Q_ASSIGN U861 ( .B(R[861]), .A(L[861]));
Q_ASSIGN U862 ( .B(R[862]), .A(L[862]));
Q_ASSIGN U863 ( .B(R[863]), .A(L[863]));
Q_ASSIGN U864 ( .B(R[864]), .A(L[864]));
Q_ASSIGN U865 ( .B(R[865]), .A(L[865]));
Q_ASSIGN U866 ( .B(R[866]), .A(L[866]));
Q_ASSIGN U867 ( .B(R[867]), .A(L[867]));
Q_ASSIGN U868 ( .B(R[868]), .A(L[868]));
Q_ASSIGN U869 ( .B(R[869]), .A(L[869]));
Q_ASSIGN U870 ( .B(R[870]), .A(L[870]));
Q_ASSIGN U871 ( .B(R[871]), .A(L[871]));
Q_ASSIGN U872 ( .B(R[872]), .A(L[872]));
Q_ASSIGN U873 ( .B(R[873]), .A(L[873]));
Q_ASSIGN U874 ( .B(R[874]), .A(L[874]));
Q_ASSIGN U875 ( .B(R[875]), .A(L[875]));
Q_ASSIGN U876 ( .B(R[876]), .A(L[876]));
Q_ASSIGN U877 ( .B(R[877]), .A(L[877]));
Q_ASSIGN U878 ( .B(R[878]), .A(L[878]));
Q_ASSIGN U879 ( .B(R[879]), .A(L[879]));
Q_ASSIGN U880 ( .B(R[880]), .A(L[880]));
Q_ASSIGN U881 ( .B(R[881]), .A(L[881]));
Q_ASSIGN U882 ( .B(R[882]), .A(L[882]));
Q_ASSIGN U883 ( .B(R[883]), .A(L[883]));
Q_ASSIGN U884 ( .B(R[884]), .A(L[884]));
Q_ASSIGN U885 ( .B(R[885]), .A(L[885]));
Q_ASSIGN U886 ( .B(R[886]), .A(L[886]));
Q_ASSIGN U887 ( .B(R[887]), .A(L[887]));
Q_ASSIGN U888 ( .B(R[888]), .A(L[888]));
Q_ASSIGN U889 ( .B(R[889]), .A(L[889]));
Q_ASSIGN U890 ( .B(R[890]), .A(L[890]));
Q_ASSIGN U891 ( .B(R[891]), .A(L[891]));
Q_ASSIGN U892 ( .B(R[892]), .A(L[892]));
Q_ASSIGN U893 ( .B(R[893]), .A(L[893]));
Q_ASSIGN U894 ( .B(R[894]), .A(L[894]));
Q_ASSIGN U895 ( .B(R[895]), .A(L[895]));
Q_ASSIGN U896 ( .B(R[896]), .A(L[896]));
Q_ASSIGN U897 ( .B(R[897]), .A(L[897]));
Q_ASSIGN U898 ( .B(R[898]), .A(L[898]));
Q_ASSIGN U899 ( .B(R[899]), .A(L[899]));
Q_ASSIGN U900 ( .B(R[900]), .A(L[900]));
Q_ASSIGN U901 ( .B(R[901]), .A(L[901]));
Q_ASSIGN U902 ( .B(R[902]), .A(L[902]));
Q_ASSIGN U903 ( .B(R[903]), .A(L[903]));
Q_ASSIGN U904 ( .B(R[904]), .A(L[904]));
Q_ASSIGN U905 ( .B(R[905]), .A(L[905]));
Q_ASSIGN U906 ( .B(R[906]), .A(L[906]));
Q_ASSIGN U907 ( .B(R[907]), .A(L[907]));
Q_ASSIGN U908 ( .B(R[908]), .A(L[908]));
Q_ASSIGN U909 ( .B(R[909]), .A(L[909]));
Q_ASSIGN U910 ( .B(R[910]), .A(L[910]));
Q_ASSIGN U911 ( .B(R[911]), .A(L[911]));
Q_ASSIGN U912 ( .B(R[912]), .A(L[912]));
Q_ASSIGN U913 ( .B(R[913]), .A(L[913]));
Q_ASSIGN U914 ( .B(R[914]), .A(L[914]));
Q_ASSIGN U915 ( .B(R[915]), .A(L[915]));
Q_ASSIGN U916 ( .B(R[916]), .A(L[916]));
Q_ASSIGN U917 ( .B(R[917]), .A(L[917]));
Q_ASSIGN U918 ( .B(R[918]), .A(L[918]));
Q_ASSIGN U919 ( .B(R[919]), .A(L[919]));
Q_ASSIGN U920 ( .B(R[920]), .A(L[920]));
Q_ASSIGN U921 ( .B(R[921]), .A(L[921]));
Q_ASSIGN U922 ( .B(R[922]), .A(L[922]));
Q_ASSIGN U923 ( .B(R[923]), .A(L[923]));
Q_ASSIGN U924 ( .B(R[924]), .A(L[924]));
Q_ASSIGN U925 ( .B(R[925]), .A(L[925]));
Q_ASSIGN U926 ( .B(R[926]), .A(L[926]));
Q_ASSIGN U927 ( .B(R[927]), .A(L[927]));
Q_ASSIGN U928 ( .B(R[928]), .A(L[928]));
Q_ASSIGN U929 ( .B(R[929]), .A(L[929]));
Q_ASSIGN U930 ( .B(R[930]), .A(L[930]));
Q_ASSIGN U931 ( .B(R[931]), .A(L[931]));
Q_ASSIGN U932 ( .B(R[932]), .A(L[932]));
Q_ASSIGN U933 ( .B(R[933]), .A(L[933]));
Q_ASSIGN U934 ( .B(R[934]), .A(L[934]));
Q_ASSIGN U935 ( .B(R[935]), .A(L[935]));
Q_ASSIGN U936 ( .B(R[936]), .A(L[936]));
Q_ASSIGN U937 ( .B(R[937]), .A(L[937]));
Q_ASSIGN U938 ( .B(R[938]), .A(L[938]));
Q_ASSIGN U939 ( .B(R[939]), .A(L[939]));
Q_ASSIGN U940 ( .B(R[940]), .A(L[940]));
Q_ASSIGN U941 ( .B(R[941]), .A(L[941]));
Q_ASSIGN U942 ( .B(R[942]), .A(L[942]));
Q_ASSIGN U943 ( .B(R[943]), .A(L[943]));
Q_ASSIGN U944 ( .B(R[944]), .A(L[944]));
Q_ASSIGN U945 ( .B(R[945]), .A(L[945]));
Q_ASSIGN U946 ( .B(R[946]), .A(L[946]));
Q_ASSIGN U947 ( .B(R[947]), .A(L[947]));
Q_ASSIGN U948 ( .B(R[948]), .A(L[948]));
Q_ASSIGN U949 ( .B(R[949]), .A(L[949]));
Q_ASSIGN U950 ( .B(R[950]), .A(L[950]));
Q_ASSIGN U951 ( .B(R[951]), .A(L[951]));
Q_ASSIGN U952 ( .B(R[952]), .A(L[952]));
Q_ASSIGN U953 ( .B(R[953]), .A(L[953]));
Q_ASSIGN U954 ( .B(R[954]), .A(L[954]));
Q_ASSIGN U955 ( .B(R[955]), .A(L[955]));
Q_ASSIGN U956 ( .B(R[956]), .A(L[956]));
Q_ASSIGN U957 ( .B(R[957]), .A(L[957]));
Q_ASSIGN U958 ( .B(R[958]), .A(L[958]));
Q_ASSIGN U959 ( .B(R[959]), .A(L[959]));
Q_ASSIGN U960 ( .B(R[960]), .A(L[960]));
Q_ASSIGN U961 ( .B(R[961]), .A(L[961]));
Q_ASSIGN U962 ( .B(R[962]), .A(L[962]));
Q_ASSIGN U963 ( .B(R[963]), .A(L[963]));
Q_ASSIGN U964 ( .B(R[964]), .A(L[964]));
Q_ASSIGN U965 ( .B(R[965]), .A(L[965]));
Q_ASSIGN U966 ( .B(R[966]), .A(L[966]));
Q_ASSIGN U967 ( .B(R[967]), .A(L[967]));
Q_ASSIGN U968 ( .B(R[968]), .A(L[968]));
Q_ASSIGN U969 ( .B(R[969]), .A(L[969]));
Q_ASSIGN U970 ( .B(R[970]), .A(L[970]));
Q_ASSIGN U971 ( .B(R[971]), .A(L[971]));
Q_ASSIGN U972 ( .B(R[972]), .A(L[972]));
Q_ASSIGN U973 ( .B(R[973]), .A(L[973]));
Q_ASSIGN U974 ( .B(R[974]), .A(L[974]));
Q_ASSIGN U975 ( .B(R[975]), .A(L[975]));
Q_ASSIGN U976 ( .B(R[976]), .A(L[976]));
Q_ASSIGN U977 ( .B(R[977]), .A(L[977]));
Q_ASSIGN U978 ( .B(R[978]), .A(L[978]));
Q_ASSIGN U979 ( .B(R[979]), .A(L[979]));
Q_ASSIGN U980 ( .B(R[980]), .A(L[980]));
Q_ASSIGN U981 ( .B(R[981]), .A(L[981]));
Q_ASSIGN U982 ( .B(R[982]), .A(L[982]));
Q_ASSIGN U983 ( .B(R[983]), .A(L[983]));
Q_ASSIGN U984 ( .B(R[984]), .A(L[984]));
Q_ASSIGN U985 ( .B(R[985]), .A(L[985]));
Q_ASSIGN U986 ( .B(R[986]), .A(L[986]));
Q_ASSIGN U987 ( .B(R[987]), .A(L[987]));
Q_ASSIGN U988 ( .B(R[988]), .A(L[988]));
Q_ASSIGN U989 ( .B(R[989]), .A(L[989]));
Q_ASSIGN U990 ( .B(R[990]), .A(L[990]));
Q_ASSIGN U991 ( .B(R[991]), .A(L[991]));
Q_ASSIGN U992 ( .B(R[992]), .A(L[992]));
Q_ASSIGN U993 ( .B(R[993]), .A(L[993]));
Q_ASSIGN U994 ( .B(R[994]), .A(L[994]));
Q_ASSIGN U995 ( .B(R[995]), .A(L[995]));
Q_ASSIGN U996 ( .B(R[996]), .A(L[996]));
Q_ASSIGN U997 ( .B(R[997]), .A(L[997]));
Q_ASSIGN U998 ( .B(R[998]), .A(L[998]));
Q_ASSIGN U999 ( .B(R[999]), .A(L[999]));
Q_ASSIGN U1000 ( .B(R[1000]), .A(L[1000]));
Q_ASSIGN U1001 ( .B(R[1001]), .A(L[1001]));
Q_ASSIGN U1002 ( .B(R[1002]), .A(L[1002]));
Q_ASSIGN U1003 ( .B(R[1003]), .A(L[1003]));
Q_ASSIGN U1004 ( .B(R[1004]), .A(L[1004]));
Q_ASSIGN U1005 ( .B(R[1005]), .A(L[1005]));
Q_ASSIGN U1006 ( .B(R[1006]), .A(L[1006]));
Q_ASSIGN U1007 ( .B(R[1007]), .A(L[1007]));
Q_ASSIGN U1008 ( .B(R[1008]), .A(L[1008]));
Q_ASSIGN U1009 ( .B(R[1009]), .A(L[1009]));
Q_ASSIGN U1010 ( .B(R[1010]), .A(L[1010]));
Q_ASSIGN U1011 ( .B(R[1011]), .A(L[1011]));
Q_ASSIGN U1012 ( .B(R[1012]), .A(L[1012]));
Q_ASSIGN U1013 ( .B(R[1013]), .A(L[1013]));
Q_ASSIGN U1014 ( .B(R[1014]), .A(L[1014]));
Q_ASSIGN U1015 ( .B(R[1015]), .A(L[1015]));
Q_ASSIGN U1016 ( .B(R[1016]), .A(L[1016]));
Q_ASSIGN U1017 ( .B(R[1017]), .A(L[1017]));
Q_ASSIGN U1018 ( .B(R[1018]), .A(L[1018]));
Q_ASSIGN U1019 ( .B(R[1019]), .A(L[1019]));
Q_ASSIGN U1020 ( .B(R[1020]), .A(L[1020]));
Q_ASSIGN U1021 ( .B(R[1021]), .A(L[1021]));
Q_ASSIGN U1022 ( .B(R[1022]), .A(L[1022]));
Q_ASSIGN U1023 ( .B(R[1023]), .A(L[1023]));
Q_ASSIGN U1024 ( .B(R[1024]), .A(L[1024]));
Q_ASSIGN U1025 ( .B(R[1025]), .A(L[1025]));
Q_ASSIGN U1026 ( .B(R[1026]), .A(L[1026]));
Q_ASSIGN U1027 ( .B(R[1027]), .A(L[1027]));
Q_ASSIGN U1028 ( .B(R[1028]), .A(L[1028]));
Q_ASSIGN U1029 ( .B(R[1029]), .A(L[1029]));
Q_ASSIGN U1030 ( .B(R[1030]), .A(L[1030]));
Q_ASSIGN U1031 ( .B(R[1031]), .A(L[1031]));
Q_ASSIGN U1032 ( .B(R[1032]), .A(L[1032]));
Q_ASSIGN U1033 ( .B(R[1033]), .A(L[1033]));
Q_ASSIGN U1034 ( .B(R[1034]), .A(L[1034]));
Q_ASSIGN U1035 ( .B(R[1035]), .A(L[1035]));
Q_ASSIGN U1036 ( .B(R[1036]), .A(L[1036]));
Q_ASSIGN U1037 ( .B(R[1037]), .A(L[1037]));
Q_ASSIGN U1038 ( .B(R[1038]), .A(L[1038]));
Q_ASSIGN U1039 ( .B(R[1039]), .A(L[1039]));
Q_ASSIGN U1040 ( .B(R[1040]), .A(L[1040]));
Q_ASSIGN U1041 ( .B(R[1041]), .A(L[1041]));
Q_ASSIGN U1042 ( .B(R[1042]), .A(L[1042]));
Q_ASSIGN U1043 ( .B(R[1043]), .A(L[1043]));
Q_ASSIGN U1044 ( .B(R[1044]), .A(L[1044]));
Q_ASSIGN U1045 ( .B(R[1045]), .A(L[1045]));
Q_ASSIGN U1046 ( .B(R[1046]), .A(L[1046]));
Q_ASSIGN U1047 ( .B(R[1047]), .A(L[1047]));
Q_ASSIGN U1048 ( .B(R[1048]), .A(L[1048]));
Q_ASSIGN U1049 ( .B(R[1049]), .A(L[1049]));
Q_ASSIGN U1050 ( .B(R[1050]), .A(L[1050]));
Q_ASSIGN U1051 ( .B(R[1051]), .A(L[1051]));
Q_ASSIGN U1052 ( .B(R[1052]), .A(L[1052]));
Q_ASSIGN U1053 ( .B(R[1053]), .A(L[1053]));
Q_ASSIGN U1054 ( .B(R[1054]), .A(L[1054]));
Q_ASSIGN U1055 ( .B(R[1055]), .A(L[1055]));
Q_ASSIGN U1056 ( .B(R[1056]), .A(L[1056]));
Q_ASSIGN U1057 ( .B(R[1057]), .A(L[1057]));
Q_ASSIGN U1058 ( .B(R[1058]), .A(L[1058]));
Q_ASSIGN U1059 ( .B(R[1059]), .A(L[1059]));
Q_ASSIGN U1060 ( .B(R[1060]), .A(L[1060]));
Q_ASSIGN U1061 ( .B(R[1061]), .A(L[1061]));
Q_ASSIGN U1062 ( .B(R[1062]), .A(L[1062]));
Q_ASSIGN U1063 ( .B(R[1063]), .A(L[1063]));
Q_ASSIGN U1064 ( .B(R[1064]), .A(L[1064]));
Q_ASSIGN U1065 ( .B(R[1065]), .A(L[1065]));
Q_ASSIGN U1066 ( .B(R[1066]), .A(L[1066]));
Q_ASSIGN U1067 ( .B(R[1067]), .A(L[1067]));
Q_ASSIGN U1068 ( .B(R[1068]), .A(L[1068]));
Q_ASSIGN U1069 ( .B(R[1069]), .A(L[1069]));
Q_ASSIGN U1070 ( .B(R[1070]), .A(L[1070]));
Q_ASSIGN U1071 ( .B(R[1071]), .A(L[1071]));
Q_ASSIGN U1072 ( .B(R[1072]), .A(L[1072]));
Q_ASSIGN U1073 ( .B(R[1073]), .A(L[1073]));
Q_ASSIGN U1074 ( .B(R[1074]), .A(L[1074]));
Q_ASSIGN U1075 ( .B(R[1075]), .A(L[1075]));
Q_ASSIGN U1076 ( .B(R[1076]), .A(L[1076]));
Q_ASSIGN U1077 ( .B(R[1077]), .A(L[1077]));
Q_ASSIGN U1078 ( .B(R[1078]), .A(L[1078]));
Q_ASSIGN U1079 ( .B(R[1079]), .A(L[1079]));
Q_ASSIGN U1080 ( .B(R[1080]), .A(L[1080]));
Q_ASSIGN U1081 ( .B(R[1081]), .A(L[1081]));
Q_ASSIGN U1082 ( .B(R[1082]), .A(L[1082]));
Q_ASSIGN U1083 ( .B(R[1083]), .A(L[1083]));
Q_ASSIGN U1084 ( .B(R[1084]), .A(L[1084]));
Q_ASSIGN U1085 ( .B(R[1085]), .A(L[1085]));
Q_ASSIGN U1086 ( .B(R[1086]), .A(L[1086]));
Q_ASSIGN U1087 ( .B(R[1087]), .A(L[1087]));
Q_ASSIGN U1088 ( .B(R[1088]), .A(L[1088]));
Q_ASSIGN U1089 ( .B(R[1089]), .A(L[1089]));
Q_ASSIGN U1090 ( .B(R[1090]), .A(L[1090]));
Q_ASSIGN U1091 ( .B(R[1091]), .A(L[1091]));
Q_ASSIGN U1092 ( .B(R[1092]), .A(L[1092]));
Q_ASSIGN U1093 ( .B(R[1093]), .A(L[1093]));
Q_ASSIGN U1094 ( .B(R[1094]), .A(L[1094]));
Q_ASSIGN U1095 ( .B(R[1095]), .A(L[1095]));
Q_ASSIGN U1096 ( .B(R[1096]), .A(L[1096]));
Q_ASSIGN U1097 ( .B(R[1097]), .A(L[1097]));
Q_ASSIGN U1098 ( .B(R[1098]), .A(L[1098]));
Q_ASSIGN U1099 ( .B(R[1099]), .A(L[1099]));
Q_ASSIGN U1100 ( .B(R[1100]), .A(L[1100]));
Q_ASSIGN U1101 ( .B(R[1101]), .A(L[1101]));
Q_ASSIGN U1102 ( .B(R[1102]), .A(L[1102]));
Q_ASSIGN U1103 ( .B(R[1103]), .A(L[1103]));
Q_ASSIGN U1104 ( .B(R[1104]), .A(L[1104]));
Q_ASSIGN U1105 ( .B(R[1105]), .A(L[1105]));
Q_ASSIGN U1106 ( .B(R[1106]), .A(L[1106]));
Q_ASSIGN U1107 ( .B(R[1107]), .A(L[1107]));
Q_ASSIGN U1108 ( .B(R[1108]), .A(L[1108]));
Q_ASSIGN U1109 ( .B(R[1109]), .A(L[1109]));
Q_ASSIGN U1110 ( .B(R[1110]), .A(L[1110]));
Q_ASSIGN U1111 ( .B(R[1111]), .A(L[1111]));
Q_ASSIGN U1112 ( .B(R[1112]), .A(L[1112]));
Q_ASSIGN U1113 ( .B(R[1113]), .A(L[1113]));
Q_ASSIGN U1114 ( .B(R[1114]), .A(L[1114]));
Q_ASSIGN U1115 ( .B(R[1115]), .A(L[1115]));
Q_ASSIGN U1116 ( .B(R[1116]), .A(L[1116]));
Q_ASSIGN U1117 ( .B(R[1117]), .A(L[1117]));
Q_ASSIGN U1118 ( .B(R[1118]), .A(L[1118]));
Q_ASSIGN U1119 ( .B(R[1119]), .A(L[1119]));
Q_ASSIGN U1120 ( .B(R[1120]), .A(L[1120]));
Q_ASSIGN U1121 ( .B(R[1121]), .A(L[1121]));
Q_ASSIGN U1122 ( .B(R[1122]), .A(L[1122]));
Q_ASSIGN U1123 ( .B(R[1123]), .A(L[1123]));
Q_ASSIGN U1124 ( .B(R[1124]), .A(L[1124]));
Q_ASSIGN U1125 ( .B(R[1125]), .A(L[1125]));
Q_ASSIGN U1126 ( .B(R[1126]), .A(L[1126]));
Q_ASSIGN U1127 ( .B(R[1127]), .A(L[1127]));
Q_ASSIGN U1128 ( .B(R[1128]), .A(L[1128]));
Q_ASSIGN U1129 ( .B(R[1129]), .A(L[1129]));
Q_ASSIGN U1130 ( .B(R[1130]), .A(L[1130]));
Q_ASSIGN U1131 ( .B(R[1131]), .A(L[1131]));
Q_ASSIGN U1132 ( .B(R[1132]), .A(L[1132]));
Q_ASSIGN U1133 ( .B(R[1133]), .A(L[1133]));
Q_ASSIGN U1134 ( .B(R[1134]), .A(L[1134]));
Q_ASSIGN U1135 ( .B(R[1135]), .A(L[1135]));
Q_ASSIGN U1136 ( .B(R[1136]), .A(L[1136]));
Q_ASSIGN U1137 ( .B(R[1137]), .A(L[1137]));
Q_ASSIGN U1138 ( .B(R[1138]), .A(L[1138]));
Q_ASSIGN U1139 ( .B(R[1139]), .A(L[1139]));
Q_ASSIGN U1140 ( .B(R[1140]), .A(L[1140]));
Q_ASSIGN U1141 ( .B(R[1141]), .A(L[1141]));
Q_ASSIGN U1142 ( .B(R[1142]), .A(L[1142]));
Q_ASSIGN U1143 ( .B(R[1143]), .A(L[1143]));
Q_ASSIGN U1144 ( .B(R[1144]), .A(L[1144]));
Q_ASSIGN U1145 ( .B(R[1145]), .A(L[1145]));
Q_ASSIGN U1146 ( .B(R[1146]), .A(L[1146]));
Q_ASSIGN U1147 ( .B(R[1147]), .A(L[1147]));
Q_ASSIGN U1148 ( .B(R[1148]), .A(L[1148]));
Q_ASSIGN U1149 ( .B(R[1149]), .A(L[1149]));
Q_ASSIGN U1150 ( .B(R[1150]), .A(L[1150]));
Q_ASSIGN U1151 ( .B(R[1151]), .A(L[1151]));
Q_ASSIGN U1152 ( .B(R[1152]), .A(L[1152]));
Q_ASSIGN U1153 ( .B(R[1153]), .A(L[1153]));
Q_ASSIGN U1154 ( .B(R[1154]), .A(L[1154]));
Q_ASSIGN U1155 ( .B(R[1155]), .A(L[1155]));
Q_ASSIGN U1156 ( .B(R[1156]), .A(L[1156]));
Q_ASSIGN U1157 ( .B(R[1157]), .A(L[1157]));
Q_ASSIGN U1158 ( .B(R[1158]), .A(L[1158]));
Q_ASSIGN U1159 ( .B(R[1159]), .A(L[1159]));
Q_ASSIGN U1160 ( .B(R[1160]), .A(L[1160]));
Q_ASSIGN U1161 ( .B(R[1161]), .A(L[1161]));
Q_ASSIGN U1162 ( .B(R[1162]), .A(L[1162]));
Q_ASSIGN U1163 ( .B(R[1163]), .A(L[1163]));
Q_ASSIGN U1164 ( .B(R[1164]), .A(L[1164]));
Q_ASSIGN U1165 ( .B(R[1165]), .A(L[1165]));
Q_ASSIGN U1166 ( .B(R[1166]), .A(L[1166]));
Q_ASSIGN U1167 ( .B(R[1167]), .A(L[1167]));
Q_ASSIGN U1168 ( .B(R[1168]), .A(L[1168]));
Q_ASSIGN U1169 ( .B(R[1169]), .A(L[1169]));
Q_ASSIGN U1170 ( .B(R[1170]), .A(L[1170]));
Q_ASSIGN U1171 ( .B(R[1171]), .A(L[1171]));
Q_ASSIGN U1172 ( .B(R[1172]), .A(L[1172]));
Q_ASSIGN U1173 ( .B(R[1173]), .A(L[1173]));
Q_ASSIGN U1174 ( .B(R[1174]), .A(L[1174]));
Q_ASSIGN U1175 ( .B(R[1175]), .A(L[1175]));
Q_ASSIGN U1176 ( .B(R[1176]), .A(L[1176]));
Q_ASSIGN U1177 ( .B(R[1177]), .A(L[1177]));
Q_ASSIGN U1178 ( .B(R[1178]), .A(L[1178]));
Q_ASSIGN U1179 ( .B(R[1179]), .A(L[1179]));
Q_ASSIGN U1180 ( .B(R[1180]), .A(L[1180]));
Q_ASSIGN U1181 ( .B(R[1181]), .A(L[1181]));
Q_ASSIGN U1182 ( .B(R[1182]), .A(L[1182]));
Q_ASSIGN U1183 ( .B(R[1183]), .A(L[1183]));
Q_ASSIGN U1184 ( .B(R[1184]), .A(L[1184]));
Q_ASSIGN U1185 ( .B(R[1185]), .A(L[1185]));
Q_ASSIGN U1186 ( .B(R[1186]), .A(L[1186]));
Q_ASSIGN U1187 ( .B(R[1187]), .A(L[1187]));
Q_ASSIGN U1188 ( .B(R[1188]), .A(L[1188]));
Q_ASSIGN U1189 ( .B(R[1189]), .A(L[1189]));
Q_ASSIGN U1190 ( .B(R[1190]), .A(L[1190]));
Q_ASSIGN U1191 ( .B(R[1191]), .A(L[1191]));
Q_ASSIGN U1192 ( .B(R[1192]), .A(L[1192]));
Q_ASSIGN U1193 ( .B(R[1193]), .A(L[1193]));
Q_ASSIGN U1194 ( .B(R[1194]), .A(L[1194]));
Q_ASSIGN U1195 ( .B(R[1195]), .A(L[1195]));
Q_ASSIGN U1196 ( .B(R[1196]), .A(L[1196]));
Q_ASSIGN U1197 ( .B(R[1197]), .A(L[1197]));
Q_ASSIGN U1198 ( .B(R[1198]), .A(L[1198]));
Q_ASSIGN U1199 ( .B(R[1199]), .A(L[1199]));
Q_ASSIGN U1200 ( .B(R[1200]), .A(L[1200]));
Q_ASSIGN U1201 ( .B(R[1201]), .A(L[1201]));
Q_ASSIGN U1202 ( .B(R[1202]), .A(L[1202]));
Q_ASSIGN U1203 ( .B(R[1203]), .A(L[1203]));
Q_ASSIGN U1204 ( .B(R[1204]), .A(L[1204]));
Q_ASSIGN U1205 ( .B(R[1205]), .A(L[1205]));
Q_ASSIGN U1206 ( .B(R[1206]), .A(L[1206]));
Q_ASSIGN U1207 ( .B(R[1207]), .A(L[1207]));
Q_ASSIGN U1208 ( .B(R[1208]), .A(L[1208]));
Q_ASSIGN U1209 ( .B(R[1209]), .A(L[1209]));
Q_ASSIGN U1210 ( .B(R[1210]), .A(L[1210]));
Q_ASSIGN U1211 ( .B(R[1211]), .A(L[1211]));
Q_ASSIGN U1212 ( .B(R[1212]), .A(L[1212]));
Q_ASSIGN U1213 ( .B(R[1213]), .A(L[1213]));
Q_ASSIGN U1214 ( .B(R[1214]), .A(L[1214]));
Q_ASSIGN U1215 ( .B(R[1215]), .A(L[1215]));
Q_ASSIGN U1216 ( .B(R[1216]), .A(L[1216]));
Q_ASSIGN U1217 ( .B(R[1217]), .A(L[1217]));
Q_ASSIGN U1218 ( .B(R[1218]), .A(L[1218]));
Q_ASSIGN U1219 ( .B(R[1219]), .A(L[1219]));
Q_ASSIGN U1220 ( .B(R[1220]), .A(L[1220]));
Q_ASSIGN U1221 ( .B(R[1221]), .A(L[1221]));
Q_ASSIGN U1222 ( .B(R[1222]), .A(L[1222]));
Q_ASSIGN U1223 ( .B(R[1223]), .A(L[1223]));
Q_ASSIGN U1224 ( .B(R[1224]), .A(L[1224]));
Q_ASSIGN U1225 ( .B(R[1225]), .A(L[1225]));
Q_ASSIGN U1226 ( .B(R[1226]), .A(L[1226]));
Q_ASSIGN U1227 ( .B(R[1227]), .A(L[1227]));
Q_ASSIGN U1228 ( .B(R[1228]), .A(L[1228]));
Q_ASSIGN U1229 ( .B(R[1229]), .A(L[1229]));
Q_ASSIGN U1230 ( .B(R[1230]), .A(L[1230]));
Q_ASSIGN U1231 ( .B(R[1231]), .A(L[1231]));
Q_ASSIGN U1232 ( .B(R[1232]), .A(L[1232]));
Q_ASSIGN U1233 ( .B(R[1233]), .A(L[1233]));
Q_ASSIGN U1234 ( .B(R[1234]), .A(L[1234]));
Q_ASSIGN U1235 ( .B(R[1235]), .A(L[1235]));
Q_ASSIGN U1236 ( .B(R[1236]), .A(L[1236]));
Q_ASSIGN U1237 ( .B(R[1237]), .A(L[1237]));
Q_ASSIGN U1238 ( .B(R[1238]), .A(L[1238]));
Q_ASSIGN U1239 ( .B(R[1239]), .A(L[1239]));
Q_ASSIGN U1240 ( .B(R[1240]), .A(L[1240]));
Q_ASSIGN U1241 ( .B(R[1241]), .A(L[1241]));
Q_ASSIGN U1242 ( .B(R[1242]), .A(L[1242]));
Q_ASSIGN U1243 ( .B(R[1243]), .A(L[1243]));
Q_ASSIGN U1244 ( .B(R[1244]), .A(L[1244]));
Q_ASSIGN U1245 ( .B(R[1245]), .A(L[1245]));
Q_ASSIGN U1246 ( .B(R[1246]), .A(L[1246]));
Q_ASSIGN U1247 ( .B(R[1247]), .A(L[1247]));
Q_ASSIGN U1248 ( .B(R[1248]), .A(L[1248]));
Q_ASSIGN U1249 ( .B(R[1249]), .A(L[1249]));
Q_ASSIGN U1250 ( .B(R[1250]), .A(L[1250]));
Q_ASSIGN U1251 ( .B(R[1251]), .A(L[1251]));
Q_ASSIGN U1252 ( .B(R[1252]), .A(L[1252]));
Q_ASSIGN U1253 ( .B(R[1253]), .A(L[1253]));
Q_ASSIGN U1254 ( .B(R[1254]), .A(L[1254]));
Q_ASSIGN U1255 ( .B(R[1255]), .A(L[1255]));
Q_ASSIGN U1256 ( .B(R[1256]), .A(L[1256]));
Q_ASSIGN U1257 ( .B(R[1257]), .A(L[1257]));
Q_ASSIGN U1258 ( .B(R[1258]), .A(L[1258]));
Q_ASSIGN U1259 ( .B(R[1259]), .A(L[1259]));
Q_ASSIGN U1260 ( .B(R[1260]), .A(L[1260]));
Q_ASSIGN U1261 ( .B(R[1261]), .A(L[1261]));
Q_ASSIGN U1262 ( .B(R[1262]), .A(L[1262]));
Q_ASSIGN U1263 ( .B(R[1263]), .A(L[1263]));
Q_ASSIGN U1264 ( .B(R[1264]), .A(L[1264]));
Q_ASSIGN U1265 ( .B(R[1265]), .A(L[1265]));
Q_ASSIGN U1266 ( .B(R[1266]), .A(L[1266]));
Q_ASSIGN U1267 ( .B(R[1267]), .A(L[1267]));
Q_ASSIGN U1268 ( .B(R[1268]), .A(L[1268]));
Q_ASSIGN U1269 ( .B(R[1269]), .A(L[1269]));
Q_ASSIGN U1270 ( .B(R[1270]), .A(L[1270]));
Q_ASSIGN U1271 ( .B(R[1271]), .A(L[1271]));
Q_ASSIGN U1272 ( .B(R[1272]), .A(L[1272]));
Q_ASSIGN U1273 ( .B(R[1273]), .A(L[1273]));
Q_ASSIGN U1274 ( .B(R[1274]), .A(L[1274]));
Q_ASSIGN U1275 ( .B(R[1275]), .A(L[1275]));
Q_ASSIGN U1276 ( .B(R[1276]), .A(L[1276]));
Q_ASSIGN U1277 ( .B(R[1277]), .A(L[1277]));
Q_ASSIGN U1278 ( .B(R[1278]), .A(L[1278]));
Q_ASSIGN U1279 ( .B(R[1279]), .A(L[1279]));
Q_ASSIGN U1280 ( .B(R[1280]), .A(L[1280]));
Q_ASSIGN U1281 ( .B(R[1281]), .A(L[1281]));
Q_ASSIGN U1282 ( .B(R[1282]), .A(L[1282]));
Q_ASSIGN U1283 ( .B(R[1283]), .A(L[1283]));
Q_ASSIGN U1284 ( .B(R[1284]), .A(L[1284]));
Q_ASSIGN U1285 ( .B(R[1285]), .A(L[1285]));
Q_ASSIGN U1286 ( .B(R[1286]), .A(L[1286]));
Q_ASSIGN U1287 ( .B(R[1287]), .A(L[1287]));
Q_ASSIGN U1288 ( .B(R[1288]), .A(L[1288]));
Q_ASSIGN U1289 ( .B(R[1289]), .A(L[1289]));
Q_ASSIGN U1290 ( .B(R[1290]), .A(L[1290]));
Q_ASSIGN U1291 ( .B(R[1291]), .A(L[1291]));
Q_ASSIGN U1292 ( .B(R[1292]), .A(L[1292]));
Q_ASSIGN U1293 ( .B(R[1293]), .A(L[1293]));
Q_ASSIGN U1294 ( .B(R[1294]), .A(L[1294]));
Q_ASSIGN U1295 ( .B(R[1295]), .A(L[1295]));
Q_ASSIGN U1296 ( .B(R[1296]), .A(L[1296]));
Q_ASSIGN U1297 ( .B(R[1297]), .A(L[1297]));
Q_ASSIGN U1298 ( .B(R[1298]), .A(L[1298]));
Q_ASSIGN U1299 ( .B(R[1299]), .A(L[1299]));
Q_ASSIGN U1300 ( .B(R[1300]), .A(L[1300]));
Q_ASSIGN U1301 ( .B(R[1301]), .A(L[1301]));
Q_ASSIGN U1302 ( .B(R[1302]), .A(L[1302]));
Q_ASSIGN U1303 ( .B(R[1303]), .A(L[1303]));
Q_ASSIGN U1304 ( .B(R[1304]), .A(L[1304]));
Q_ASSIGN U1305 ( .B(R[1305]), .A(L[1305]));
Q_ASSIGN U1306 ( .B(R[1306]), .A(L[1306]));
Q_ASSIGN U1307 ( .B(R[1307]), .A(L[1307]));
Q_ASSIGN U1308 ( .B(R[1308]), .A(L[1308]));
Q_ASSIGN U1309 ( .B(R[1309]), .A(L[1309]));
Q_ASSIGN U1310 ( .B(R[1310]), .A(L[1310]));
Q_ASSIGN U1311 ( .B(R[1311]), .A(L[1311]));
Q_ASSIGN U1312 ( .B(R[1312]), .A(L[1312]));
Q_ASSIGN U1313 ( .B(R[1313]), .A(L[1313]));
Q_ASSIGN U1314 ( .B(R[1314]), .A(L[1314]));
Q_ASSIGN U1315 ( .B(R[1315]), .A(L[1315]));
Q_ASSIGN U1316 ( .B(R[1316]), .A(L[1316]));
Q_ASSIGN U1317 ( .B(R[1317]), .A(L[1317]));
Q_ASSIGN U1318 ( .B(R[1318]), .A(L[1318]));
Q_ASSIGN U1319 ( .B(R[1319]), .A(L[1319]));
Q_ASSIGN U1320 ( .B(R[1320]), .A(L[1320]));
Q_ASSIGN U1321 ( .B(R[1321]), .A(L[1321]));
Q_ASSIGN U1322 ( .B(R[1322]), .A(L[1322]));
Q_ASSIGN U1323 ( .B(R[1323]), .A(L[1323]));
Q_ASSIGN U1324 ( .B(R[1324]), .A(L[1324]));
Q_ASSIGN U1325 ( .B(R[1325]), .A(L[1325]));
Q_ASSIGN U1326 ( .B(R[1326]), .A(L[1326]));
Q_ASSIGN U1327 ( .B(R[1327]), .A(L[1327]));
Q_ASSIGN U1328 ( .B(R[1328]), .A(L[1328]));
Q_ASSIGN U1329 ( .B(R[1329]), .A(L[1329]));
Q_ASSIGN U1330 ( .B(R[1330]), .A(L[1330]));
Q_ASSIGN U1331 ( .B(R[1331]), .A(L[1331]));
Q_ASSIGN U1332 ( .B(R[1332]), .A(L[1332]));
Q_ASSIGN U1333 ( .B(R[1333]), .A(L[1333]));
Q_ASSIGN U1334 ( .B(R[1334]), .A(L[1334]));
Q_ASSIGN U1335 ( .B(R[1335]), .A(L[1335]));
Q_ASSIGN U1336 ( .B(R[1336]), .A(L[1336]));
Q_ASSIGN U1337 ( .B(R[1337]), .A(L[1337]));
Q_ASSIGN U1338 ( .B(R[1338]), .A(L[1338]));
Q_ASSIGN U1339 ( .B(R[1339]), .A(L[1339]));
Q_ASSIGN U1340 ( .B(R[1340]), .A(L[1340]));
Q_ASSIGN U1341 ( .B(R[1341]), .A(L[1341]));
Q_ASSIGN U1342 ( .B(R[1342]), .A(L[1342]));
Q_ASSIGN U1343 ( .B(R[1343]), .A(L[1343]));
Q_ASSIGN U1344 ( .B(R[1344]), .A(L[1344]));
Q_ASSIGN U1345 ( .B(R[1345]), .A(L[1345]));
Q_ASSIGN U1346 ( .B(R[1346]), .A(L[1346]));
Q_ASSIGN U1347 ( .B(R[1347]), .A(L[1347]));
Q_ASSIGN U1348 ( .B(R[1348]), .A(L[1348]));
Q_ASSIGN U1349 ( .B(R[1349]), .A(L[1349]));
Q_ASSIGN U1350 ( .B(R[1350]), .A(L[1350]));
Q_ASSIGN U1351 ( .B(R[1351]), .A(L[1351]));
Q_ASSIGN U1352 ( .B(R[1352]), .A(L[1352]));
Q_ASSIGN U1353 ( .B(R[1353]), .A(L[1353]));
Q_ASSIGN U1354 ( .B(R[1354]), .A(L[1354]));
Q_ASSIGN U1355 ( .B(R[1355]), .A(L[1355]));
Q_ASSIGN U1356 ( .B(R[1356]), .A(L[1356]));
Q_ASSIGN U1357 ( .B(R[1357]), .A(L[1357]));
Q_ASSIGN U1358 ( .B(R[1358]), .A(L[1358]));
Q_ASSIGN U1359 ( .B(R[1359]), .A(L[1359]));
Q_ASSIGN U1360 ( .B(R[1360]), .A(L[1360]));
Q_ASSIGN U1361 ( .B(R[1361]), .A(L[1361]));
Q_ASSIGN U1362 ( .B(R[1362]), .A(L[1362]));
Q_ASSIGN U1363 ( .B(R[1363]), .A(L[1363]));
Q_ASSIGN U1364 ( .B(R[1364]), .A(L[1364]));
Q_ASSIGN U1365 ( .B(R[1365]), .A(L[1365]));
Q_ASSIGN U1366 ( .B(R[1366]), .A(L[1366]));
Q_ASSIGN U1367 ( .B(R[1367]), .A(L[1367]));
Q_ASSIGN U1368 ( .B(R[1368]), .A(L[1368]));
Q_ASSIGN U1369 ( .B(R[1369]), .A(L[1369]));
Q_ASSIGN U1370 ( .B(R[1370]), .A(L[1370]));
Q_ASSIGN U1371 ( .B(R[1371]), .A(L[1371]));
Q_ASSIGN U1372 ( .B(R[1372]), .A(L[1372]));
Q_ASSIGN U1373 ( .B(R[1373]), .A(L[1373]));
Q_ASSIGN U1374 ( .B(R[1374]), .A(L[1374]));
Q_ASSIGN U1375 ( .B(R[1375]), .A(L[1375]));
Q_ASSIGN U1376 ( .B(R[1376]), .A(L[1376]));
Q_ASSIGN U1377 ( .B(R[1377]), .A(L[1377]));
Q_ASSIGN U1378 ( .B(R[1378]), .A(L[1378]));
Q_ASSIGN U1379 ( .B(R[1379]), .A(L[1379]));
Q_ASSIGN U1380 ( .B(R[1380]), .A(L[1380]));
Q_ASSIGN U1381 ( .B(R[1381]), .A(L[1381]));
Q_ASSIGN U1382 ( .B(R[1382]), .A(L[1382]));
Q_ASSIGN U1383 ( .B(R[1383]), .A(L[1383]));
Q_ASSIGN U1384 ( .B(R[1384]), .A(L[1384]));
Q_ASSIGN U1385 ( .B(R[1385]), .A(L[1385]));
Q_ASSIGN U1386 ( .B(R[1386]), .A(L[1386]));
Q_ASSIGN U1387 ( .B(R[1387]), .A(L[1387]));
Q_ASSIGN U1388 ( .B(R[1388]), .A(L[1388]));
Q_ASSIGN U1389 ( .B(R[1389]), .A(L[1389]));
Q_ASSIGN U1390 ( .B(R[1390]), .A(L[1390]));
Q_ASSIGN U1391 ( .B(R[1391]), .A(L[1391]));
Q_ASSIGN U1392 ( .B(R[1392]), .A(L[1392]));
Q_ASSIGN U1393 ( .B(R[1393]), .A(L[1393]));
Q_ASSIGN U1394 ( .B(R[1394]), .A(L[1394]));
Q_ASSIGN U1395 ( .B(R[1395]), .A(L[1395]));
Q_ASSIGN U1396 ( .B(R[1396]), .A(L[1396]));
Q_ASSIGN U1397 ( .B(R[1397]), .A(L[1397]));
Q_ASSIGN U1398 ( .B(R[1398]), .A(L[1398]));
Q_ASSIGN U1399 ( .B(R[1399]), .A(L[1399]));
Q_ASSIGN U1400 ( .B(R[1400]), .A(L[1400]));
Q_ASSIGN U1401 ( .B(R[1401]), .A(L[1401]));
Q_ASSIGN U1402 ( .B(R[1402]), .A(L[1402]));
Q_ASSIGN U1403 ( .B(R[1403]), .A(L[1403]));
Q_ASSIGN U1404 ( .B(R[1404]), .A(L[1404]));
Q_ASSIGN U1405 ( .B(R[1405]), .A(L[1405]));
Q_ASSIGN U1406 ( .B(R[1406]), .A(L[1406]));
Q_ASSIGN U1407 ( .B(R[1407]), .A(L[1407]));
Q_ASSIGN U1408 ( .B(R[1408]), .A(L[1408]));
Q_ASSIGN U1409 ( .B(R[1409]), .A(L[1409]));
Q_ASSIGN U1410 ( .B(R[1410]), .A(L[1410]));
Q_ASSIGN U1411 ( .B(R[1411]), .A(L[1411]));
Q_ASSIGN U1412 ( .B(R[1412]), .A(L[1412]));
Q_ASSIGN U1413 ( .B(R[1413]), .A(L[1413]));
Q_ASSIGN U1414 ( .B(R[1414]), .A(L[1414]));
Q_ASSIGN U1415 ( .B(R[1415]), .A(L[1415]));
Q_ASSIGN U1416 ( .B(R[1416]), .A(L[1416]));
Q_ASSIGN U1417 ( .B(R[1417]), .A(L[1417]));
Q_ASSIGN U1418 ( .B(R[1418]), .A(L[1418]));
Q_ASSIGN U1419 ( .B(R[1419]), .A(L[1419]));
Q_ASSIGN U1420 ( .B(R[1420]), .A(L[1420]));
Q_ASSIGN U1421 ( .B(R[1421]), .A(L[1421]));
Q_ASSIGN U1422 ( .B(R[1422]), .A(L[1422]));
Q_ASSIGN U1423 ( .B(R[1423]), .A(L[1423]));
Q_ASSIGN U1424 ( .B(R[1424]), .A(L[1424]));
Q_ASSIGN U1425 ( .B(R[1425]), .A(L[1425]));
Q_ASSIGN U1426 ( .B(R[1426]), .A(L[1426]));
Q_ASSIGN U1427 ( .B(R[1427]), .A(L[1427]));
Q_ASSIGN U1428 ( .B(R[1428]), .A(L[1428]));
Q_ASSIGN U1429 ( .B(R[1429]), .A(L[1429]));
Q_ASSIGN U1430 ( .B(R[1430]), .A(L[1430]));
Q_ASSIGN U1431 ( .B(R[1431]), .A(L[1431]));
Q_ASSIGN U1432 ( .B(R[1432]), .A(L[1432]));
Q_ASSIGN U1433 ( .B(R[1433]), .A(L[1433]));
Q_ASSIGN U1434 ( .B(R[1434]), .A(L[1434]));
Q_ASSIGN U1435 ( .B(R[1435]), .A(L[1435]));
Q_ASSIGN U1436 ( .B(R[1436]), .A(L[1436]));
Q_ASSIGN U1437 ( .B(R[1437]), .A(L[1437]));
Q_ASSIGN U1438 ( .B(R[1438]), .A(L[1438]));
Q_ASSIGN U1439 ( .B(R[1439]), .A(L[1439]));
Q_ASSIGN U1440 ( .B(R[1440]), .A(L[1440]));
Q_ASSIGN U1441 ( .B(R[1441]), .A(L[1441]));
Q_ASSIGN U1442 ( .B(R[1442]), .A(L[1442]));
Q_ASSIGN U1443 ( .B(R[1443]), .A(L[1443]));
Q_ASSIGN U1444 ( .B(R[1444]), .A(L[1444]));
Q_ASSIGN U1445 ( .B(R[1445]), .A(L[1445]));
Q_ASSIGN U1446 ( .B(R[1446]), .A(L[1446]));
Q_ASSIGN U1447 ( .B(R[1447]), .A(L[1447]));
Q_ASSIGN U1448 ( .B(R[1448]), .A(L[1448]));
Q_ASSIGN U1449 ( .B(R[1449]), .A(L[1449]));
Q_ASSIGN U1450 ( .B(R[1450]), .A(L[1450]));
Q_ASSIGN U1451 ( .B(R[1451]), .A(L[1451]));
Q_ASSIGN U1452 ( .B(R[1452]), .A(L[1452]));
Q_ASSIGN U1453 ( .B(R[1453]), .A(L[1453]));
Q_ASSIGN U1454 ( .B(R[1454]), .A(L[1454]));
Q_ASSIGN U1455 ( .B(R[1455]), .A(L[1455]));
Q_ASSIGN U1456 ( .B(R[1456]), .A(L[1456]));
Q_ASSIGN U1457 ( .B(R[1457]), .A(L[1457]));
Q_ASSIGN U1458 ( .B(R[1458]), .A(L[1458]));
Q_ASSIGN U1459 ( .B(R[1459]), .A(L[1459]));
Q_ASSIGN U1460 ( .B(R[1460]), .A(L[1460]));
Q_ASSIGN U1461 ( .B(R[1461]), .A(L[1461]));
Q_ASSIGN U1462 ( .B(R[1462]), .A(L[1462]));
Q_ASSIGN U1463 ( .B(R[1463]), .A(L[1463]));
Q_ASSIGN U1464 ( .B(R[1464]), .A(L[1464]));
Q_ASSIGN U1465 ( .B(R[1465]), .A(L[1465]));
Q_ASSIGN U1466 ( .B(R[1466]), .A(L[1466]));
Q_ASSIGN U1467 ( .B(R[1467]), .A(L[1467]));
Q_ASSIGN U1468 ( .B(R[1468]), .A(L[1468]));
Q_ASSIGN U1469 ( .B(R[1469]), .A(L[1469]));
Q_ASSIGN U1470 ( .B(R[1470]), .A(L[1470]));
Q_ASSIGN U1471 ( .B(R[1471]), .A(L[1471]));
Q_ASSIGN U1472 ( .B(R[1472]), .A(L[1472]));
Q_ASSIGN U1473 ( .B(R[1473]), .A(L[1473]));
Q_ASSIGN U1474 ( .B(R[1474]), .A(L[1474]));
Q_ASSIGN U1475 ( .B(R[1475]), .A(L[1475]));
Q_ASSIGN U1476 ( .B(R[1476]), .A(L[1476]));
Q_ASSIGN U1477 ( .B(R[1477]), .A(L[1477]));
Q_ASSIGN U1478 ( .B(R[1478]), .A(L[1478]));
Q_ASSIGN U1479 ( .B(R[1479]), .A(L[1479]));
Q_ASSIGN U1480 ( .B(R[1480]), .A(L[1480]));
Q_ASSIGN U1481 ( .B(R[1481]), .A(L[1481]));
Q_ASSIGN U1482 ( .B(R[1482]), .A(L[1482]));
Q_ASSIGN U1483 ( .B(R[1483]), .A(L[1483]));
Q_ASSIGN U1484 ( .B(R[1484]), .A(L[1484]));
Q_ASSIGN U1485 ( .B(R[1485]), .A(L[1485]));
Q_ASSIGN U1486 ( .B(R[1486]), .A(L[1486]));
Q_ASSIGN U1487 ( .B(R[1487]), .A(L[1487]));
Q_ASSIGN U1488 ( .B(R[1488]), .A(L[1488]));
Q_ASSIGN U1489 ( .B(R[1489]), .A(L[1489]));
Q_ASSIGN U1490 ( .B(R[1490]), .A(L[1490]));
Q_ASSIGN U1491 ( .B(R[1491]), .A(L[1491]));
Q_ASSIGN U1492 ( .B(R[1492]), .A(L[1492]));
Q_ASSIGN U1493 ( .B(R[1493]), .A(L[1493]));
Q_ASSIGN U1494 ( .B(R[1494]), .A(L[1494]));
Q_ASSIGN U1495 ( .B(R[1495]), .A(L[1495]));
Q_ASSIGN U1496 ( .B(R[1496]), .A(L[1496]));
Q_ASSIGN U1497 ( .B(R[1497]), .A(L[1497]));
Q_ASSIGN U1498 ( .B(R[1498]), .A(L[1498]));
Q_ASSIGN U1499 ( .B(R[1499]), .A(L[1499]));
Q_ASSIGN U1500 ( .B(R[1500]), .A(L[1500]));
Q_ASSIGN U1501 ( .B(R[1501]), .A(L[1501]));
Q_ASSIGN U1502 ( .B(R[1502]), .A(L[1502]));
Q_ASSIGN U1503 ( .B(R[1503]), .A(L[1503]));
Q_ASSIGN U1504 ( .B(R[1504]), .A(L[1504]));
Q_ASSIGN U1505 ( .B(R[1505]), .A(L[1505]));
Q_ASSIGN U1506 ( .B(R[1506]), .A(L[1506]));
Q_ASSIGN U1507 ( .B(R[1507]), .A(L[1507]));
Q_ASSIGN U1508 ( .B(R[1508]), .A(L[1508]));
Q_ASSIGN U1509 ( .B(R[1509]), .A(L[1509]));
Q_ASSIGN U1510 ( .B(R[1510]), .A(L[1510]));
Q_ASSIGN U1511 ( .B(R[1511]), .A(L[1511]));
Q_ASSIGN U1512 ( .B(R[1512]), .A(L[1512]));
Q_ASSIGN U1513 ( .B(R[1513]), .A(L[1513]));
Q_ASSIGN U1514 ( .B(R[1514]), .A(L[1514]));
Q_ASSIGN U1515 ( .B(R[1515]), .A(L[1515]));
Q_ASSIGN U1516 ( .B(R[1516]), .A(L[1516]));
Q_ASSIGN U1517 ( .B(R[1517]), .A(L[1517]));
Q_ASSIGN U1518 ( .B(R[1518]), .A(L[1518]));
Q_ASSIGN U1519 ( .B(R[1519]), .A(L[1519]));
Q_ASSIGN U1520 ( .B(R[1520]), .A(L[1520]));
Q_ASSIGN U1521 ( .B(R[1521]), .A(L[1521]));
Q_ASSIGN U1522 ( .B(R[1522]), .A(L[1522]));
Q_ASSIGN U1523 ( .B(R[1523]), .A(L[1523]));
Q_ASSIGN U1524 ( .B(R[1524]), .A(L[1524]));
Q_ASSIGN U1525 ( .B(R[1525]), .A(L[1525]));
Q_ASSIGN U1526 ( .B(R[1526]), .A(L[1526]));
Q_ASSIGN U1527 ( .B(R[1527]), .A(L[1527]));
Q_ASSIGN U1528 ( .B(R[1528]), .A(L[1528]));
Q_ASSIGN U1529 ( .B(R[1529]), .A(L[1529]));
Q_ASSIGN U1530 ( .B(R[1530]), .A(L[1530]));
Q_ASSIGN U1531 ( .B(R[1531]), .A(L[1531]));
Q_ASSIGN U1532 ( .B(R[1532]), .A(L[1532]));
Q_ASSIGN U1533 ( .B(R[1533]), .A(L[1533]));
Q_ASSIGN U1534 ( .B(R[1534]), .A(L[1534]));
Q_ASSIGN U1535 ( .B(R[1535]), .A(L[1535]));
Q_ASSIGN U1536 ( .B(R[1536]), .A(L[1536]));
Q_ASSIGN U1537 ( .B(R[1537]), .A(L[1537]));
Q_ASSIGN U1538 ( .B(R[1538]), .A(L[1538]));
Q_ASSIGN U1539 ( .B(R[1539]), .A(L[1539]));
Q_ASSIGN U1540 ( .B(R[1540]), .A(L[1540]));
Q_ASSIGN U1541 ( .B(R[1541]), .A(L[1541]));
Q_ASSIGN U1542 ( .B(R[1542]), .A(L[1542]));
Q_ASSIGN U1543 ( .B(R[1543]), .A(L[1543]));
Q_ASSIGN U1544 ( .B(R[1544]), .A(L[1544]));
Q_ASSIGN U1545 ( .B(R[1545]), .A(L[1545]));
Q_ASSIGN U1546 ( .B(R[1546]), .A(L[1546]));
Q_ASSIGN U1547 ( .B(R[1547]), .A(L[1547]));
Q_ASSIGN U1548 ( .B(R[1548]), .A(L[1548]));
Q_ASSIGN U1549 ( .B(R[1549]), .A(L[1549]));
Q_ASSIGN U1550 ( .B(R[1550]), .A(L[1550]));
Q_ASSIGN U1551 ( .B(R[1551]), .A(L[1551]));
Q_ASSIGN U1552 ( .B(R[1552]), .A(L[1552]));
Q_ASSIGN U1553 ( .B(R[1553]), .A(L[1553]));
Q_ASSIGN U1554 ( .B(R[1554]), .A(L[1554]));
Q_ASSIGN U1555 ( .B(R[1555]), .A(L[1555]));
Q_ASSIGN U1556 ( .B(R[1556]), .A(L[1556]));
Q_ASSIGN U1557 ( .B(R[1557]), .A(L[1557]));
Q_ASSIGN U1558 ( .B(R[1558]), .A(L[1558]));
Q_ASSIGN U1559 ( .B(R[1559]), .A(L[1559]));
Q_ASSIGN U1560 ( .B(R[1560]), .A(L[1560]));
Q_ASSIGN U1561 ( .B(R[1561]), .A(L[1561]));
Q_ASSIGN U1562 ( .B(R[1562]), .A(L[1562]));
Q_ASSIGN U1563 ( .B(R[1563]), .A(L[1563]));
Q_ASSIGN U1564 ( .B(R[1564]), .A(L[1564]));
Q_ASSIGN U1565 ( .B(R[1565]), .A(L[1565]));
Q_ASSIGN U1566 ( .B(R[1566]), .A(L[1566]));
Q_ASSIGN U1567 ( .B(R[1567]), .A(L[1567]));
Q_ASSIGN U1568 ( .B(R[1568]), .A(L[1568]));
Q_ASSIGN U1569 ( .B(R[1569]), .A(L[1569]));
Q_ASSIGN U1570 ( .B(R[1570]), .A(L[1570]));
Q_ASSIGN U1571 ( .B(R[1571]), .A(L[1571]));
Q_ASSIGN U1572 ( .B(R[1572]), .A(L[1572]));
Q_ASSIGN U1573 ( .B(R[1573]), .A(L[1573]));
Q_ASSIGN U1574 ( .B(R[1574]), .A(L[1574]));
Q_ASSIGN U1575 ( .B(R[1575]), .A(L[1575]));
Q_ASSIGN U1576 ( .B(R[1576]), .A(L[1576]));
Q_ASSIGN U1577 ( .B(R[1577]), .A(L[1577]));
Q_ASSIGN U1578 ( .B(R[1578]), .A(L[1578]));
Q_ASSIGN U1579 ( .B(R[1579]), .A(L[1579]));
Q_ASSIGN U1580 ( .B(R[1580]), .A(L[1580]));
Q_ASSIGN U1581 ( .B(R[1581]), .A(L[1581]));
Q_ASSIGN U1582 ( .B(R[1582]), .A(L[1582]));
Q_ASSIGN U1583 ( .B(R[1583]), .A(L[1583]));
Q_ASSIGN U1584 ( .B(R[1584]), .A(L[1584]));
Q_ASSIGN U1585 ( .B(R[1585]), .A(L[1585]));
Q_ASSIGN U1586 ( .B(R[1586]), .A(L[1586]));
Q_ASSIGN U1587 ( .B(R[1587]), .A(L[1587]));
Q_ASSIGN U1588 ( .B(R[1588]), .A(L[1588]));
Q_ASSIGN U1589 ( .B(R[1589]), .A(L[1589]));
Q_ASSIGN U1590 ( .B(R[1590]), .A(L[1590]));
Q_ASSIGN U1591 ( .B(R[1591]), .A(L[1591]));
Q_ASSIGN U1592 ( .B(R[1592]), .A(L[1592]));
Q_ASSIGN U1593 ( .B(R[1593]), .A(L[1593]));
Q_ASSIGN U1594 ( .B(R[1594]), .A(L[1594]));
Q_ASSIGN U1595 ( .B(R[1595]), .A(L[1595]));
Q_ASSIGN U1596 ( .B(R[1596]), .A(L[1596]));
Q_ASSIGN U1597 ( .B(R[1597]), .A(L[1597]));
Q_ASSIGN U1598 ( .B(R[1598]), .A(L[1598]));
Q_ASSIGN U1599 ( .B(R[1599]), .A(L[1599]));
Q_ASSIGN U1600 ( .B(R[1600]), .A(L[1600]));
Q_ASSIGN U1601 ( .B(R[1601]), .A(L[1601]));
Q_ASSIGN U1602 ( .B(R[1602]), .A(L[1602]));
Q_ASSIGN U1603 ( .B(R[1603]), .A(L[1603]));
Q_ASSIGN U1604 ( .B(R[1604]), .A(L[1604]));
Q_ASSIGN U1605 ( .B(R[1605]), .A(L[1605]));
Q_ASSIGN U1606 ( .B(R[1606]), .A(L[1606]));
Q_ASSIGN U1607 ( .B(R[1607]), .A(L[1607]));
Q_ASSIGN U1608 ( .B(R[1608]), .A(L[1608]));
Q_ASSIGN U1609 ( .B(R[1609]), .A(L[1609]));
Q_ASSIGN U1610 ( .B(R[1610]), .A(L[1610]));
Q_ASSIGN U1611 ( .B(R[1611]), .A(L[1611]));
Q_ASSIGN U1612 ( .B(R[1612]), .A(L[1612]));
Q_ASSIGN U1613 ( .B(R[1613]), .A(L[1613]));
Q_ASSIGN U1614 ( .B(R[1614]), .A(L[1614]));
Q_ASSIGN U1615 ( .B(R[1615]), .A(L[1615]));
Q_ASSIGN U1616 ( .B(R[1616]), .A(L[1616]));
Q_ASSIGN U1617 ( .B(R[1617]), .A(L[1617]));
Q_ASSIGN U1618 ( .B(R[1618]), .A(L[1618]));
Q_ASSIGN U1619 ( .B(R[1619]), .A(L[1619]));
Q_ASSIGN U1620 ( .B(R[1620]), .A(L[1620]));
Q_ASSIGN U1621 ( .B(R[1621]), .A(L[1621]));
Q_ASSIGN U1622 ( .B(R[1622]), .A(L[1622]));
Q_ASSIGN U1623 ( .B(R[1623]), .A(L[1623]));
Q_ASSIGN U1624 ( .B(R[1624]), .A(L[1624]));
Q_ASSIGN U1625 ( .B(R[1625]), .A(L[1625]));
Q_ASSIGN U1626 ( .B(R[1626]), .A(L[1626]));
Q_ASSIGN U1627 ( .B(R[1627]), .A(L[1627]));
Q_ASSIGN U1628 ( .B(R[1628]), .A(L[1628]));
Q_ASSIGN U1629 ( .B(R[1629]), .A(L[1629]));
Q_ASSIGN U1630 ( .B(R[1630]), .A(L[1630]));
Q_ASSIGN U1631 ( .B(R[1631]), .A(L[1631]));
Q_ASSIGN U1632 ( .B(R[1632]), .A(L[1632]));
Q_ASSIGN U1633 ( .B(R[1633]), .A(L[1633]));
Q_ASSIGN U1634 ( .B(R[1634]), .A(L[1634]));
Q_ASSIGN U1635 ( .B(R[1635]), .A(L[1635]));
Q_ASSIGN U1636 ( .B(R[1636]), .A(L[1636]));
Q_ASSIGN U1637 ( .B(R[1637]), .A(L[1637]));
Q_ASSIGN U1638 ( .B(R[1638]), .A(L[1638]));
Q_ASSIGN U1639 ( .B(R[1639]), .A(L[1639]));
Q_ASSIGN U1640 ( .B(R[1640]), .A(L[1640]));
Q_ASSIGN U1641 ( .B(R[1641]), .A(L[1641]));
Q_ASSIGN U1642 ( .B(R[1642]), .A(L[1642]));
Q_ASSIGN U1643 ( .B(R[1643]), .A(L[1643]));
Q_ASSIGN U1644 ( .B(R[1644]), .A(L[1644]));
Q_ASSIGN U1645 ( .B(R[1645]), .A(L[1645]));
Q_ASSIGN U1646 ( .B(R[1646]), .A(L[1646]));
Q_ASSIGN U1647 ( .B(R[1647]), .A(L[1647]));
Q_ASSIGN U1648 ( .B(R[1648]), .A(L[1648]));
Q_ASSIGN U1649 ( .B(R[1649]), .A(L[1649]));
Q_ASSIGN U1650 ( .B(R[1650]), .A(L[1650]));
Q_ASSIGN U1651 ( .B(R[1651]), .A(L[1651]));
Q_ASSIGN U1652 ( .B(R[1652]), .A(L[1652]));
Q_ASSIGN U1653 ( .B(R[1653]), .A(L[1653]));
Q_ASSIGN U1654 ( .B(R[1654]), .A(L[1654]));
Q_ASSIGN U1655 ( .B(R[1655]), .A(L[1655]));
Q_ASSIGN U1656 ( .B(R[1656]), .A(L[1656]));
Q_ASSIGN U1657 ( .B(R[1657]), .A(L[1657]));
Q_ASSIGN U1658 ( .B(R[1658]), .A(L[1658]));
Q_ASSIGN U1659 ( .B(R[1659]), .A(L[1659]));
Q_ASSIGN U1660 ( .B(R[1660]), .A(L[1660]));
Q_ASSIGN U1661 ( .B(R[1661]), .A(L[1661]));
Q_ASSIGN U1662 ( .B(R[1662]), .A(L[1662]));
Q_ASSIGN U1663 ( .B(R[1663]), .A(L[1663]));
Q_ASSIGN U1664 ( .B(R[1664]), .A(L[1664]));
Q_ASSIGN U1665 ( .B(R[1665]), .A(L[1665]));
Q_ASSIGN U1666 ( .B(R[1666]), .A(L[1666]));
Q_ASSIGN U1667 ( .B(R[1667]), .A(L[1667]));
Q_ASSIGN U1668 ( .B(R[1668]), .A(L[1668]));
Q_ASSIGN U1669 ( .B(R[1669]), .A(L[1669]));
Q_ASSIGN U1670 ( .B(R[1670]), .A(L[1670]));
Q_ASSIGN U1671 ( .B(R[1671]), .A(L[1671]));
Q_ASSIGN U1672 ( .B(R[1672]), .A(L[1672]));
Q_ASSIGN U1673 ( .B(R[1673]), .A(L[1673]));
Q_ASSIGN U1674 ( .B(R[1674]), .A(L[1674]));
Q_ASSIGN U1675 ( .B(R[1675]), .A(L[1675]));
Q_ASSIGN U1676 ( .B(R[1676]), .A(L[1676]));
Q_ASSIGN U1677 ( .B(R[1677]), .A(L[1677]));
Q_ASSIGN U1678 ( .B(R[1678]), .A(L[1678]));
Q_ASSIGN U1679 ( .B(R[1679]), .A(L[1679]));
Q_ASSIGN U1680 ( .B(R[1680]), .A(L[1680]));
Q_ASSIGN U1681 ( .B(R[1681]), .A(L[1681]));
Q_ASSIGN U1682 ( .B(R[1682]), .A(L[1682]));
Q_ASSIGN U1683 ( .B(R[1683]), .A(L[1683]));
Q_ASSIGN U1684 ( .B(R[1684]), .A(L[1684]));
Q_ASSIGN U1685 ( .B(R[1685]), .A(L[1685]));
Q_ASSIGN U1686 ( .B(R[1686]), .A(L[1686]));
Q_ASSIGN U1687 ( .B(R[1687]), .A(L[1687]));
Q_ASSIGN U1688 ( .B(R[1688]), .A(L[1688]));
Q_ASSIGN U1689 ( .B(R[1689]), .A(L[1689]));
Q_ASSIGN U1690 ( .B(R[1690]), .A(L[1690]));
Q_ASSIGN U1691 ( .B(R[1691]), .A(L[1691]));
Q_ASSIGN U1692 ( .B(R[1692]), .A(L[1692]));
Q_ASSIGN U1693 ( .B(R[1693]), .A(L[1693]));
Q_ASSIGN U1694 ( .B(R[1694]), .A(L[1694]));
Q_ASSIGN U1695 ( .B(R[1695]), .A(L[1695]));
Q_ASSIGN U1696 ( .B(R[1696]), .A(L[1696]));
Q_ASSIGN U1697 ( .B(R[1697]), .A(L[1697]));
Q_ASSIGN U1698 ( .B(R[1698]), .A(L[1698]));
Q_ASSIGN U1699 ( .B(R[1699]), .A(L[1699]));
Q_ASSIGN U1700 ( .B(R[1700]), .A(L[1700]));
Q_ASSIGN U1701 ( .B(R[1701]), .A(L[1701]));
Q_ASSIGN U1702 ( .B(R[1702]), .A(L[1702]));
Q_ASSIGN U1703 ( .B(R[1703]), .A(L[1703]));
Q_ASSIGN U1704 ( .B(R[1704]), .A(L[1704]));
Q_ASSIGN U1705 ( .B(R[1705]), .A(L[1705]));
Q_ASSIGN U1706 ( .B(R[1706]), .A(L[1706]));
Q_ASSIGN U1707 ( .B(R[1707]), .A(L[1707]));
Q_ASSIGN U1708 ( .B(R[1708]), .A(L[1708]));
Q_ASSIGN U1709 ( .B(R[1709]), .A(L[1709]));
Q_ASSIGN U1710 ( .B(R[1710]), .A(L[1710]));
Q_ASSIGN U1711 ( .B(R[1711]), .A(L[1711]));
Q_ASSIGN U1712 ( .B(R[1712]), .A(L[1712]));
Q_ASSIGN U1713 ( .B(R[1713]), .A(L[1713]));
Q_ASSIGN U1714 ( .B(R[1714]), .A(L[1714]));
Q_ASSIGN U1715 ( .B(R[1715]), .A(L[1715]));
Q_ASSIGN U1716 ( .B(R[1716]), .A(L[1716]));
Q_ASSIGN U1717 ( .B(R[1717]), .A(L[1717]));
Q_ASSIGN U1718 ( .B(R[1718]), .A(L[1718]));
Q_ASSIGN U1719 ( .B(R[1719]), .A(L[1719]));
Q_ASSIGN U1720 ( .B(R[1720]), .A(L[1720]));
Q_ASSIGN U1721 ( .B(R[1721]), .A(L[1721]));
Q_ASSIGN U1722 ( .B(R[1722]), .A(L[1722]));
Q_ASSIGN U1723 ( .B(R[1723]), .A(L[1723]));
Q_ASSIGN U1724 ( .B(R[1724]), .A(L[1724]));
Q_ASSIGN U1725 ( .B(R[1725]), .A(L[1725]));
Q_ASSIGN U1726 ( .B(R[1726]), .A(L[1726]));
Q_ASSIGN U1727 ( .B(R[1727]), .A(L[1727]));
Q_ASSIGN U1728 ( .B(R[1728]), .A(L[1728]));
Q_ASSIGN U1729 ( .B(R[1729]), .A(L[1729]));
Q_ASSIGN U1730 ( .B(R[1730]), .A(L[1730]));
Q_ASSIGN U1731 ( .B(R[1731]), .A(L[1731]));
Q_ASSIGN U1732 ( .B(R[1732]), .A(L[1732]));
Q_ASSIGN U1733 ( .B(R[1733]), .A(L[1733]));
Q_ASSIGN U1734 ( .B(R[1734]), .A(L[1734]));
Q_ASSIGN U1735 ( .B(R[1735]), .A(L[1735]));
Q_ASSIGN U1736 ( .B(R[1736]), .A(L[1736]));
Q_ASSIGN U1737 ( .B(R[1737]), .A(L[1737]));
Q_ASSIGN U1738 ( .B(R[1738]), .A(L[1738]));
Q_ASSIGN U1739 ( .B(R[1739]), .A(L[1739]));
Q_ASSIGN U1740 ( .B(R[1740]), .A(L[1740]));
Q_ASSIGN U1741 ( .B(R[1741]), .A(L[1741]));
Q_ASSIGN U1742 ( .B(R[1742]), .A(L[1742]));
Q_ASSIGN U1743 ( .B(R[1743]), .A(L[1743]));
Q_ASSIGN U1744 ( .B(R[1744]), .A(L[1744]));
Q_ASSIGN U1745 ( .B(R[1745]), .A(L[1745]));
Q_ASSIGN U1746 ( .B(R[1746]), .A(L[1746]));
Q_ASSIGN U1747 ( .B(R[1747]), .A(L[1747]));
Q_ASSIGN U1748 ( .B(R[1748]), .A(L[1748]));
Q_ASSIGN U1749 ( .B(R[1749]), .A(L[1749]));
Q_ASSIGN U1750 ( .B(R[1750]), .A(L[1750]));
Q_ASSIGN U1751 ( .B(R[1751]), .A(L[1751]));
Q_ASSIGN U1752 ( .B(R[1752]), .A(L[1752]));
Q_ASSIGN U1753 ( .B(R[1753]), .A(L[1753]));
Q_ASSIGN U1754 ( .B(R[1754]), .A(L[1754]));
Q_ASSIGN U1755 ( .B(R[1755]), .A(L[1755]));
Q_ASSIGN U1756 ( .B(R[1756]), .A(L[1756]));
Q_ASSIGN U1757 ( .B(R[1757]), .A(L[1757]));
Q_ASSIGN U1758 ( .B(R[1758]), .A(L[1758]));
Q_ASSIGN U1759 ( .B(R[1759]), .A(L[1759]));
Q_ASSIGN U1760 ( .B(R[1760]), .A(L[1760]));
Q_ASSIGN U1761 ( .B(R[1761]), .A(L[1761]));
Q_ASSIGN U1762 ( .B(R[1762]), .A(L[1762]));
Q_ASSIGN U1763 ( .B(R[1763]), .A(L[1763]));
Q_ASSIGN U1764 ( .B(R[1764]), .A(L[1764]));
Q_ASSIGN U1765 ( .B(R[1765]), .A(L[1765]));
Q_ASSIGN U1766 ( .B(R[1766]), .A(L[1766]));
Q_ASSIGN U1767 ( .B(R[1767]), .A(L[1767]));
Q_ASSIGN U1768 ( .B(R[1768]), .A(L[1768]));
Q_ASSIGN U1769 ( .B(R[1769]), .A(L[1769]));
Q_ASSIGN U1770 ( .B(R[1770]), .A(L[1770]));
Q_ASSIGN U1771 ( .B(R[1771]), .A(L[1771]));
Q_ASSIGN U1772 ( .B(R[1772]), .A(L[1772]));
Q_ASSIGN U1773 ( .B(R[1773]), .A(L[1773]));
Q_ASSIGN U1774 ( .B(R[1774]), .A(L[1774]));
Q_ASSIGN U1775 ( .B(R[1775]), .A(L[1775]));
Q_ASSIGN U1776 ( .B(R[1776]), .A(L[1776]));
Q_ASSIGN U1777 ( .B(R[1777]), .A(L[1777]));
Q_ASSIGN U1778 ( .B(R[1778]), .A(L[1778]));
Q_ASSIGN U1779 ( .B(R[1779]), .A(L[1779]));
Q_ASSIGN U1780 ( .B(R[1780]), .A(L[1780]));
Q_ASSIGN U1781 ( .B(R[1781]), .A(L[1781]));
Q_ASSIGN U1782 ( .B(R[1782]), .A(L[1782]));
Q_ASSIGN U1783 ( .B(R[1783]), .A(L[1783]));
Q_ASSIGN U1784 ( .B(R[1784]), .A(L[1784]));
Q_ASSIGN U1785 ( .B(R[1785]), .A(L[1785]));
Q_ASSIGN U1786 ( .B(R[1786]), .A(L[1786]));
Q_ASSIGN U1787 ( .B(R[1787]), .A(L[1787]));
Q_ASSIGN U1788 ( .B(R[1788]), .A(L[1788]));
Q_ASSIGN U1789 ( .B(R[1789]), .A(L[1789]));
Q_ASSIGN U1790 ( .B(R[1790]), .A(L[1790]));
Q_ASSIGN U1791 ( .B(R[1791]), .A(L[1791]));
Q_ASSIGN U1792 ( .B(R[1792]), .A(L[1792]));
Q_ASSIGN U1793 ( .B(R[1793]), .A(L[1793]));
Q_ASSIGN U1794 ( .B(R[1794]), .A(L[1794]));
Q_ASSIGN U1795 ( .B(R[1795]), .A(L[1795]));
Q_ASSIGN U1796 ( .B(R[1796]), .A(L[1796]));
Q_ASSIGN U1797 ( .B(R[1797]), .A(L[1797]));
Q_ASSIGN U1798 ( .B(R[1798]), .A(L[1798]));
Q_ASSIGN U1799 ( .B(R[1799]), .A(L[1799]));
Q_ASSIGN U1800 ( .B(R[1800]), .A(L[1800]));
Q_ASSIGN U1801 ( .B(R[1801]), .A(L[1801]));
Q_ASSIGN U1802 ( .B(R[1802]), .A(L[1802]));
Q_ASSIGN U1803 ( .B(R[1803]), .A(L[1803]));
Q_ASSIGN U1804 ( .B(R[1804]), .A(L[1804]));
Q_ASSIGN U1805 ( .B(R[1805]), .A(L[1805]));
Q_ASSIGN U1806 ( .B(R[1806]), .A(L[1806]));
Q_ASSIGN U1807 ( .B(R[1807]), .A(L[1807]));
Q_ASSIGN U1808 ( .B(R[1808]), .A(L[1808]));
Q_ASSIGN U1809 ( .B(R[1809]), .A(L[1809]));
Q_ASSIGN U1810 ( .B(R[1810]), .A(L[1810]));
Q_ASSIGN U1811 ( .B(R[1811]), .A(L[1811]));
Q_ASSIGN U1812 ( .B(R[1812]), .A(L[1812]));
Q_ASSIGN U1813 ( .B(R[1813]), .A(L[1813]));
Q_ASSIGN U1814 ( .B(R[1814]), .A(L[1814]));
Q_ASSIGN U1815 ( .B(R[1815]), .A(L[1815]));
Q_ASSIGN U1816 ( .B(R[1816]), .A(L[1816]));
Q_ASSIGN U1817 ( .B(R[1817]), .A(L[1817]));
Q_ASSIGN U1818 ( .B(R[1818]), .A(L[1818]));
Q_ASSIGN U1819 ( .B(R[1819]), .A(L[1819]));
Q_ASSIGN U1820 ( .B(R[1820]), .A(L[1820]));
Q_ASSIGN U1821 ( .B(R[1821]), .A(L[1821]));
Q_ASSIGN U1822 ( .B(R[1822]), .A(L[1822]));
Q_ASSIGN U1823 ( .B(R[1823]), .A(L[1823]));
Q_ASSIGN U1824 ( .B(R[1824]), .A(L[1824]));
Q_ASSIGN U1825 ( .B(R[1825]), .A(L[1825]));
Q_ASSIGN U1826 ( .B(R[1826]), .A(L[1826]));
Q_ASSIGN U1827 ( .B(R[1827]), .A(L[1827]));
Q_ASSIGN U1828 ( .B(R[1828]), .A(L[1828]));
Q_ASSIGN U1829 ( .B(R[1829]), .A(L[1829]));
Q_ASSIGN U1830 ( .B(R[1830]), .A(L[1830]));
Q_ASSIGN U1831 ( .B(R[1831]), .A(L[1831]));
Q_ASSIGN U1832 ( .B(R[1832]), .A(L[1832]));
Q_ASSIGN U1833 ( .B(R[1833]), .A(L[1833]));
Q_ASSIGN U1834 ( .B(R[1834]), .A(L[1834]));
Q_ASSIGN U1835 ( .B(R[1835]), .A(L[1835]));
Q_ASSIGN U1836 ( .B(R[1836]), .A(L[1836]));
Q_ASSIGN U1837 ( .B(R[1837]), .A(L[1837]));
Q_ASSIGN U1838 ( .B(R[1838]), .A(L[1838]));
Q_ASSIGN U1839 ( .B(R[1839]), .A(L[1839]));
Q_ASSIGN U1840 ( .B(R[1840]), .A(L[1840]));
Q_ASSIGN U1841 ( .B(R[1841]), .A(L[1841]));
Q_ASSIGN U1842 ( .B(R[1842]), .A(L[1842]));
Q_ASSIGN U1843 ( .B(R[1843]), .A(L[1843]));
Q_ASSIGN U1844 ( .B(R[1844]), .A(L[1844]));
Q_ASSIGN U1845 ( .B(R[1845]), .A(L[1845]));
Q_ASSIGN U1846 ( .B(R[1846]), .A(L[1846]));
Q_ASSIGN U1847 ( .B(R[1847]), .A(L[1847]));
Q_ASSIGN U1848 ( .B(R[1848]), .A(L[1848]));
Q_ASSIGN U1849 ( .B(R[1849]), .A(L[1849]));
Q_ASSIGN U1850 ( .B(R[1850]), .A(L[1850]));
Q_ASSIGN U1851 ( .B(R[1851]), .A(L[1851]));
Q_ASSIGN U1852 ( .B(R[1852]), .A(L[1852]));
Q_ASSIGN U1853 ( .B(R[1853]), .A(L[1853]));
Q_ASSIGN U1854 ( .B(R[1854]), .A(L[1854]));
Q_ASSIGN U1855 ( .B(R[1855]), .A(L[1855]));
Q_ASSIGN U1856 ( .B(R[1856]), .A(L[1856]));
Q_ASSIGN U1857 ( .B(R[1857]), .A(L[1857]));
Q_ASSIGN U1858 ( .B(R[1858]), .A(L[1858]));
Q_ASSIGN U1859 ( .B(R[1859]), .A(L[1859]));
Q_ASSIGN U1860 ( .B(R[1860]), .A(L[1860]));
Q_ASSIGN U1861 ( .B(R[1861]), .A(L[1861]));
Q_ASSIGN U1862 ( .B(R[1862]), .A(L[1862]));
Q_ASSIGN U1863 ( .B(R[1863]), .A(L[1863]));
Q_ASSIGN U1864 ( .B(R[1864]), .A(L[1864]));
Q_ASSIGN U1865 ( .B(R[1865]), .A(L[1865]));
Q_ASSIGN U1866 ( .B(R[1866]), .A(L[1866]));
Q_ASSIGN U1867 ( .B(R[1867]), .A(L[1867]));
Q_ASSIGN U1868 ( .B(R[1868]), .A(L[1868]));
Q_ASSIGN U1869 ( .B(R[1869]), .A(L[1869]));
Q_ASSIGN U1870 ( .B(R[1870]), .A(L[1870]));
Q_ASSIGN U1871 ( .B(R[1871]), .A(L[1871]));
Q_ASSIGN U1872 ( .B(R[1872]), .A(L[1872]));
Q_ASSIGN U1873 ( .B(R[1873]), .A(L[1873]));
Q_ASSIGN U1874 ( .B(R[1874]), .A(L[1874]));
Q_ASSIGN U1875 ( .B(R[1875]), .A(L[1875]));
Q_ASSIGN U1876 ( .B(R[1876]), .A(L[1876]));
Q_ASSIGN U1877 ( .B(R[1877]), .A(L[1877]));
Q_ASSIGN U1878 ( .B(R[1878]), .A(L[1878]));
Q_ASSIGN U1879 ( .B(R[1879]), .A(L[1879]));
Q_ASSIGN U1880 ( .B(R[1880]), .A(L[1880]));
Q_ASSIGN U1881 ( .B(R[1881]), .A(L[1881]));
Q_ASSIGN U1882 ( .B(R[1882]), .A(L[1882]));
Q_ASSIGN U1883 ( .B(R[1883]), .A(L[1883]));
Q_ASSIGN U1884 ( .B(R[1884]), .A(L[1884]));
Q_ASSIGN U1885 ( .B(R[1885]), .A(L[1885]));
Q_ASSIGN U1886 ( .B(R[1886]), .A(L[1886]));
Q_ASSIGN U1887 ( .B(R[1887]), .A(L[1887]));
Q_ASSIGN U1888 ( .B(R[1888]), .A(L[1888]));
Q_ASSIGN U1889 ( .B(R[1889]), .A(L[1889]));
Q_ASSIGN U1890 ( .B(R[1890]), .A(L[1890]));
Q_ASSIGN U1891 ( .B(R[1891]), .A(L[1891]));
Q_ASSIGN U1892 ( .B(R[1892]), .A(L[1892]));
Q_ASSIGN U1893 ( .B(R[1893]), .A(L[1893]));
Q_ASSIGN U1894 ( .B(R[1894]), .A(L[1894]));
Q_ASSIGN U1895 ( .B(R[1895]), .A(L[1895]));
Q_ASSIGN U1896 ( .B(R[1896]), .A(L[1896]));
Q_ASSIGN U1897 ( .B(R[1897]), .A(L[1897]));
Q_ASSIGN U1898 ( .B(R[1898]), .A(L[1898]));
Q_ASSIGN U1899 ( .B(R[1899]), .A(L[1899]));
Q_ASSIGN U1900 ( .B(R[1900]), .A(L[1900]));
Q_ASSIGN U1901 ( .B(R[1901]), .A(L[1901]));
Q_ASSIGN U1902 ( .B(R[1902]), .A(L[1902]));
Q_ASSIGN U1903 ( .B(R[1903]), .A(L[1903]));
Q_ASSIGN U1904 ( .B(R[1904]), .A(L[1904]));
Q_ASSIGN U1905 ( .B(R[1905]), .A(L[1905]));
Q_ASSIGN U1906 ( .B(R[1906]), .A(L[1906]));
Q_ASSIGN U1907 ( .B(R[1907]), .A(L[1907]));
Q_ASSIGN U1908 ( .B(R[1908]), .A(L[1908]));
Q_ASSIGN U1909 ( .B(R[1909]), .A(L[1909]));
Q_ASSIGN U1910 ( .B(R[1910]), .A(L[1910]));
Q_ASSIGN U1911 ( .B(R[1911]), .A(L[1911]));
Q_ASSIGN U1912 ( .B(R[1912]), .A(L[1912]));
Q_ASSIGN U1913 ( .B(R[1913]), .A(L[1913]));
Q_ASSIGN U1914 ( .B(R[1914]), .A(L[1914]));
Q_ASSIGN U1915 ( .B(R[1915]), .A(L[1915]));
Q_ASSIGN U1916 ( .B(R[1916]), .A(L[1916]));
Q_ASSIGN U1917 ( .B(R[1917]), .A(L[1917]));
Q_ASSIGN U1918 ( .B(R[1918]), .A(L[1918]));
Q_ASSIGN U1919 ( .B(R[1919]), .A(L[1919]));
Q_ASSIGN U1920 ( .B(R[1920]), .A(L[1920]));
Q_ASSIGN U1921 ( .B(R[1921]), .A(L[1921]));
Q_ASSIGN U1922 ( .B(R[1922]), .A(L[1922]));
Q_ASSIGN U1923 ( .B(R[1923]), .A(L[1923]));
Q_ASSIGN U1924 ( .B(R[1924]), .A(L[1924]));
Q_ASSIGN U1925 ( .B(R[1925]), .A(L[1925]));
Q_ASSIGN U1926 ( .B(R[1926]), .A(L[1926]));
Q_ASSIGN U1927 ( .B(R[1927]), .A(L[1927]));
Q_ASSIGN U1928 ( .B(R[1928]), .A(L[1928]));
Q_ASSIGN U1929 ( .B(R[1929]), .A(L[1929]));
Q_ASSIGN U1930 ( .B(R[1930]), .A(L[1930]));
Q_ASSIGN U1931 ( .B(R[1931]), .A(L[1931]));
Q_ASSIGN U1932 ( .B(R[1932]), .A(L[1932]));
Q_ASSIGN U1933 ( .B(R[1933]), .A(L[1933]));
Q_ASSIGN U1934 ( .B(R[1934]), .A(L[1934]));
Q_ASSIGN U1935 ( .B(R[1935]), .A(L[1935]));
Q_ASSIGN U1936 ( .B(R[1936]), .A(L[1936]));
Q_ASSIGN U1937 ( .B(R[1937]), .A(L[1937]));
Q_ASSIGN U1938 ( .B(R[1938]), .A(L[1938]));
Q_ASSIGN U1939 ( .B(R[1939]), .A(L[1939]));
Q_ASSIGN U1940 ( .B(R[1940]), .A(L[1940]));
Q_ASSIGN U1941 ( .B(R[1941]), .A(L[1941]));
Q_ASSIGN U1942 ( .B(R[1942]), .A(L[1942]));
Q_ASSIGN U1943 ( .B(R[1943]), .A(L[1943]));
Q_ASSIGN U1944 ( .B(R[1944]), .A(L[1944]));
Q_ASSIGN U1945 ( .B(R[1945]), .A(L[1945]));
Q_ASSIGN U1946 ( .B(R[1946]), .A(L[1946]));
Q_ASSIGN U1947 ( .B(R[1947]), .A(L[1947]));
Q_ASSIGN U1948 ( .B(R[1948]), .A(L[1948]));
Q_ASSIGN U1949 ( .B(R[1949]), .A(L[1949]));
Q_ASSIGN U1950 ( .B(R[1950]), .A(L[1950]));
Q_ASSIGN U1951 ( .B(R[1951]), .A(L[1951]));
Q_ASSIGN U1952 ( .B(R[1952]), .A(L[1952]));
Q_ASSIGN U1953 ( .B(R[1953]), .A(L[1953]));
Q_ASSIGN U1954 ( .B(R[1954]), .A(L[1954]));
Q_ASSIGN U1955 ( .B(R[1955]), .A(L[1955]));
Q_ASSIGN U1956 ( .B(R[1956]), .A(L[1956]));
Q_ASSIGN U1957 ( .B(R[1957]), .A(L[1957]));
Q_ASSIGN U1958 ( .B(R[1958]), .A(L[1958]));
Q_ASSIGN U1959 ( .B(R[1959]), .A(L[1959]));
Q_ASSIGN U1960 ( .B(R[1960]), .A(L[1960]));
Q_ASSIGN U1961 ( .B(R[1961]), .A(L[1961]));
Q_ASSIGN U1962 ( .B(R[1962]), .A(L[1962]));
Q_ASSIGN U1963 ( .B(R[1963]), .A(L[1963]));
Q_ASSIGN U1964 ( .B(R[1964]), .A(L[1964]));
Q_ASSIGN U1965 ( .B(R[1965]), .A(L[1965]));
Q_ASSIGN U1966 ( .B(R[1966]), .A(L[1966]));
Q_ASSIGN U1967 ( .B(R[1967]), .A(L[1967]));
Q_ASSIGN U1968 ( .B(R[1968]), .A(L[1968]));
Q_ASSIGN U1969 ( .B(R[1969]), .A(L[1969]));
Q_ASSIGN U1970 ( .B(R[1970]), .A(L[1970]));
Q_ASSIGN U1971 ( .B(R[1971]), .A(L[1971]));
Q_ASSIGN U1972 ( .B(R[1972]), .A(L[1972]));
Q_ASSIGN U1973 ( .B(R[1973]), .A(L[1973]));
Q_ASSIGN U1974 ( .B(R[1974]), .A(L[1974]));
Q_ASSIGN U1975 ( .B(R[1975]), .A(L[1975]));
Q_ASSIGN U1976 ( .B(R[1976]), .A(L[1976]));
Q_ASSIGN U1977 ( .B(R[1977]), .A(L[1977]));
Q_ASSIGN U1978 ( .B(R[1978]), .A(L[1978]));
Q_ASSIGN U1979 ( .B(R[1979]), .A(L[1979]));
Q_ASSIGN U1980 ( .B(R[1980]), .A(L[1980]));
Q_ASSIGN U1981 ( .B(R[1981]), .A(L[1981]));
Q_ASSIGN U1982 ( .B(R[1982]), .A(L[1982]));
Q_ASSIGN U1983 ( .B(R[1983]), .A(L[1983]));
Q_ASSIGN U1984 ( .B(R[1984]), .A(L[1984]));
Q_ASSIGN U1985 ( .B(R[1985]), .A(L[1985]));
Q_ASSIGN U1986 ( .B(R[1986]), .A(L[1986]));
Q_ASSIGN U1987 ( .B(R[1987]), .A(L[1987]));
Q_ASSIGN U1988 ( .B(R[1988]), .A(L[1988]));
Q_ASSIGN U1989 ( .B(R[1989]), .A(L[1989]));
Q_ASSIGN U1990 ( .B(R[1990]), .A(L[1990]));
Q_ASSIGN U1991 ( .B(R[1991]), .A(L[1991]));
Q_ASSIGN U1992 ( .B(R[1992]), .A(L[1992]));
Q_ASSIGN U1993 ( .B(R[1993]), .A(L[1993]));
Q_ASSIGN U1994 ( .B(R[1994]), .A(L[1994]));
Q_ASSIGN U1995 ( .B(R[1995]), .A(L[1995]));
Q_ASSIGN U1996 ( .B(R[1996]), .A(L[1996]));
Q_ASSIGN U1997 ( .B(R[1997]), .A(L[1997]));
Q_ASSIGN U1998 ( .B(R[1998]), .A(L[1998]));
Q_ASSIGN U1999 ( .B(R[1999]), .A(L[1999]));
Q_ASSIGN U2000 ( .B(R[2000]), .A(L[2000]));
Q_ASSIGN U2001 ( .B(R[2001]), .A(L[2001]));
Q_ASSIGN U2002 ( .B(R[2002]), .A(L[2002]));
Q_ASSIGN U2003 ( .B(R[2003]), .A(L[2003]));
Q_ASSIGN U2004 ( .B(R[2004]), .A(L[2004]));
Q_ASSIGN U2005 ( .B(R[2005]), .A(L[2005]));
Q_ASSIGN U2006 ( .B(R[2006]), .A(L[2006]));
Q_ASSIGN U2007 ( .B(R[2007]), .A(L[2007]));
Q_ASSIGN U2008 ( .B(R[2008]), .A(L[2008]));
Q_ASSIGN U2009 ( .B(R[2009]), .A(L[2009]));
Q_ASSIGN U2010 ( .B(R[2010]), .A(L[2010]));
Q_ASSIGN U2011 ( .B(R[2011]), .A(L[2011]));
Q_ASSIGN U2012 ( .B(R[2012]), .A(L[2012]));
Q_ASSIGN U2013 ( .B(R[2013]), .A(L[2013]));
Q_ASSIGN U2014 ( .B(R[2014]), .A(L[2014]));
Q_ASSIGN U2015 ( .B(R[2015]), .A(L[2015]));
Q_ASSIGN U2016 ( .B(R[2016]), .A(L[2016]));
Q_ASSIGN U2017 ( .B(R[2017]), .A(L[2017]));
Q_ASSIGN U2018 ( .B(R[2018]), .A(L[2018]));
Q_ASSIGN U2019 ( .B(R[2019]), .A(L[2019]));
Q_ASSIGN U2020 ( .B(R[2020]), .A(L[2020]));
Q_ASSIGN U2021 ( .B(R[2021]), .A(L[2021]));
Q_ASSIGN U2022 ( .B(R[2022]), .A(L[2022]));
Q_ASSIGN U2023 ( .B(R[2023]), .A(L[2023]));
Q_ASSIGN U2024 ( .B(R[2024]), .A(L[2024]));
Q_ASSIGN U2025 ( .B(R[2025]), .A(L[2025]));
Q_ASSIGN U2026 ( .B(R[2026]), .A(L[2026]));
Q_ASSIGN U2027 ( .B(R[2027]), .A(L[2027]));
Q_ASSIGN U2028 ( .B(R[2028]), .A(L[2028]));
Q_ASSIGN U2029 ( .B(R[2029]), .A(L[2029]));
Q_ASSIGN U2030 ( .B(R[2030]), .A(L[2030]));
Q_ASSIGN U2031 ( .B(R[2031]), .A(L[2031]));
Q_ASSIGN U2032 ( .B(R[2032]), .A(L[2032]));
Q_ASSIGN U2033 ( .B(R[2033]), .A(L[2033]));
Q_ASSIGN U2034 ( .B(R[2034]), .A(L[2034]));
Q_ASSIGN U2035 ( .B(R[2035]), .A(L[2035]));
Q_ASSIGN U2036 ( .B(R[2036]), .A(L[2036]));
Q_ASSIGN U2037 ( .B(R[2037]), .A(L[2037]));
Q_ASSIGN U2038 ( .B(R[2038]), .A(L[2038]));
Q_ASSIGN U2039 ( .B(R[2039]), .A(L[2039]));
Q_ASSIGN U2040 ( .B(R[2040]), .A(L[2040]));
Q_ASSIGN U2041 ( .B(R[2041]), .A(L[2041]));
Q_ASSIGN U2042 ( .B(R[2042]), .A(L[2042]));
Q_ASSIGN U2043 ( .B(R[2043]), .A(L[2043]));
Q_ASSIGN U2044 ( .B(R[2044]), .A(L[2044]));
Q_ASSIGN U2045 ( .B(R[2045]), .A(L[2045]));
Q_ASSIGN U2046 ( .B(R[2046]), .A(L[2046]));
Q_ASSIGN U2047 ( .B(R[2047]), .A(L[2047]));
Q_ASSIGN U2048 ( .B(R[2048]), .A(L[2048]));
Q_ASSIGN U2049 ( .B(R[2049]), .A(L[2049]));
Q_ASSIGN U2050 ( .B(R[2050]), .A(L[2050]));
Q_ASSIGN U2051 ( .B(R[2051]), .A(L[2051]));
Q_ASSIGN U2052 ( .B(R[2052]), .A(L[2052]));
Q_ASSIGN U2053 ( .B(R[2053]), .A(L[2053]));
Q_ASSIGN U2054 ( .B(R[2054]), .A(L[2054]));
Q_ASSIGN U2055 ( .B(R[2055]), .A(L[2055]));
Q_ASSIGN U2056 ( .B(R[2056]), .A(L[2056]));
Q_ASSIGN U2057 ( .B(R[2057]), .A(L[2057]));
Q_ASSIGN U2058 ( .B(R[2058]), .A(L[2058]));
Q_ASSIGN U2059 ( .B(R[2059]), .A(L[2059]));
Q_ASSIGN U2060 ( .B(R[2060]), .A(L[2060]));
Q_ASSIGN U2061 ( .B(R[2061]), .A(L[2061]));
Q_ASSIGN U2062 ( .B(R[2062]), .A(L[2062]));
Q_ASSIGN U2063 ( .B(R[2063]), .A(L[2063]));
Q_ASSIGN U2064 ( .B(R[2064]), .A(L[2064]));
Q_ASSIGN U2065 ( .B(R[2065]), .A(L[2065]));
Q_ASSIGN U2066 ( .B(R[2066]), .A(L[2066]));
Q_ASSIGN U2067 ( .B(R[2067]), .A(L[2067]));
Q_ASSIGN U2068 ( .B(R[2068]), .A(L[2068]));
Q_ASSIGN U2069 ( .B(R[2069]), .A(L[2069]));
Q_ASSIGN U2070 ( .B(R[2070]), .A(L[2070]));
Q_ASSIGN U2071 ( .B(R[2071]), .A(L[2071]));
Q_ASSIGN U2072 ( .B(R[2072]), .A(L[2072]));
Q_ASSIGN U2073 ( .B(R[2073]), .A(L[2073]));
Q_ASSIGN U2074 ( .B(R[2074]), .A(L[2074]));
Q_ASSIGN U2075 ( .B(R[2075]), .A(L[2075]));
Q_ASSIGN U2076 ( .B(R[2076]), .A(L[2076]));
Q_ASSIGN U2077 ( .B(R[2077]), .A(L[2077]));
Q_ASSIGN U2078 ( .B(R[2078]), .A(L[2078]));
Q_ASSIGN U2079 ( .B(R[2079]), .A(L[2079]));
Q_ASSIGN U2080 ( .B(R[2080]), .A(L[2080]));
Q_ASSIGN U2081 ( .B(R[2081]), .A(L[2081]));
Q_ASSIGN U2082 ( .B(R[2082]), .A(L[2082]));
Q_ASSIGN U2083 ( .B(R[2083]), .A(L[2083]));
Q_ASSIGN U2084 ( .B(R[2084]), .A(L[2084]));
Q_ASSIGN U2085 ( .B(R[2085]), .A(L[2085]));
Q_ASSIGN U2086 ( .B(R[2086]), .A(L[2086]));
Q_ASSIGN U2087 ( .B(R[2087]), .A(L[2087]));
Q_ASSIGN U2088 ( .B(R[2088]), .A(L[2088]));
Q_ASSIGN U2089 ( .B(R[2089]), .A(L[2089]));
Q_ASSIGN U2090 ( .B(R[2090]), .A(L[2090]));
Q_ASSIGN U2091 ( .B(R[2091]), .A(L[2091]));
Q_ASSIGN U2092 ( .B(R[2092]), .A(L[2092]));
Q_ASSIGN U2093 ( .B(R[2093]), .A(L[2093]));
Q_ASSIGN U2094 ( .B(R[2094]), .A(L[2094]));
Q_ASSIGN U2095 ( .B(R[2095]), .A(L[2095]));
Q_ASSIGN U2096 ( .B(R[2096]), .A(L[2096]));
Q_ASSIGN U2097 ( .B(R[2097]), .A(L[2097]));
Q_ASSIGN U2098 ( .B(R[2098]), .A(L[2098]));
Q_ASSIGN U2099 ( .B(R[2099]), .A(L[2099]));
Q_ASSIGN U2100 ( .B(R[2100]), .A(L[2100]));
Q_ASSIGN U2101 ( .B(R[2101]), .A(L[2101]));
Q_ASSIGN U2102 ( .B(R[2102]), .A(L[2102]));
Q_ASSIGN U2103 ( .B(R[2103]), .A(L[2103]));
Q_ASSIGN U2104 ( .B(R[2104]), .A(L[2104]));
Q_ASSIGN U2105 ( .B(R[2105]), .A(L[2105]));
Q_ASSIGN U2106 ( .B(R[2106]), .A(L[2106]));
Q_ASSIGN U2107 ( .B(R[2107]), .A(L[2107]));
Q_ASSIGN U2108 ( .B(R[2108]), .A(L[2108]));
Q_ASSIGN U2109 ( .B(R[2109]), .A(L[2109]));
Q_ASSIGN U2110 ( .B(R[2110]), .A(L[2110]));
Q_ASSIGN U2111 ( .B(R[2111]), .A(L[2111]));
Q_ASSIGN U2112 ( .B(R[2112]), .A(L[2112]));
Q_ASSIGN U2113 ( .B(R[2113]), .A(L[2113]));
Q_ASSIGN U2114 ( .B(R[2114]), .A(L[2114]));
Q_ASSIGN U2115 ( .B(R[2115]), .A(L[2115]));
Q_ASSIGN U2116 ( .B(R[2116]), .A(L[2116]));
Q_ASSIGN U2117 ( .B(R[2117]), .A(L[2117]));
Q_ASSIGN U2118 ( .B(R[2118]), .A(L[2118]));
Q_ASSIGN U2119 ( .B(R[2119]), .A(L[2119]));
Q_ASSIGN U2120 ( .B(R[2120]), .A(L[2120]));
Q_ASSIGN U2121 ( .B(R[2121]), .A(L[2121]));
Q_ASSIGN U2122 ( .B(R[2122]), .A(L[2122]));
Q_ASSIGN U2123 ( .B(R[2123]), .A(L[2123]));
Q_ASSIGN U2124 ( .B(R[2124]), .A(L[2124]));
Q_ASSIGN U2125 ( .B(R[2125]), .A(L[2125]));
Q_ASSIGN U2126 ( .B(R[2126]), .A(L[2126]));
Q_ASSIGN U2127 ( .B(R[2127]), .A(L[2127]));
Q_ASSIGN U2128 ( .B(R[2128]), .A(L[2128]));
Q_ASSIGN U2129 ( .B(R[2129]), .A(L[2129]));
Q_ASSIGN U2130 ( .B(R[2130]), .A(L[2130]));
Q_ASSIGN U2131 ( .B(R[2131]), .A(L[2131]));
Q_ASSIGN U2132 ( .B(R[2132]), .A(L[2132]));
Q_ASSIGN U2133 ( .B(R[2133]), .A(L[2133]));
Q_ASSIGN U2134 ( .B(R[2134]), .A(L[2134]));
Q_ASSIGN U2135 ( .B(R[2135]), .A(L[2135]));
Q_ASSIGN U2136 ( .B(R[2136]), .A(L[2136]));
Q_ASSIGN U2137 ( .B(R[2137]), .A(L[2137]));
Q_ASSIGN U2138 ( .B(R[2138]), .A(L[2138]));
Q_ASSIGN U2139 ( .B(R[2139]), .A(L[2139]));
Q_ASSIGN U2140 ( .B(R[2140]), .A(L[2140]));
Q_ASSIGN U2141 ( .B(R[2141]), .A(L[2141]));
Q_ASSIGN U2142 ( .B(R[2142]), .A(L[2142]));
Q_ASSIGN U2143 ( .B(R[2143]), .A(L[2143]));
Q_ASSIGN U2144 ( .B(R[2144]), .A(L[2144]));
Q_ASSIGN U2145 ( .B(R[2145]), .A(L[2145]));
Q_ASSIGN U2146 ( .B(R[2146]), .A(L[2146]));
Q_ASSIGN U2147 ( .B(R[2147]), .A(L[2147]));
Q_ASSIGN U2148 ( .B(R[2148]), .A(L[2148]));
Q_ASSIGN U2149 ( .B(R[2149]), .A(L[2149]));
Q_ASSIGN U2150 ( .B(R[2150]), .A(L[2150]));
Q_ASSIGN U2151 ( .B(R[2151]), .A(L[2151]));
Q_ASSIGN U2152 ( .B(R[2152]), .A(L[2152]));
Q_ASSIGN U2153 ( .B(R[2153]), .A(L[2153]));
Q_ASSIGN U2154 ( .B(R[2154]), .A(L[2154]));
Q_ASSIGN U2155 ( .B(R[2155]), .A(L[2155]));
Q_ASSIGN U2156 ( .B(R[2156]), .A(L[2156]));
Q_ASSIGN U2157 ( .B(R[2157]), .A(L[2157]));
Q_ASSIGN U2158 ( .B(R[2158]), .A(L[2158]));
Q_ASSIGN U2159 ( .B(R[2159]), .A(L[2159]));
Q_ASSIGN U2160 ( .B(R[2160]), .A(L[2160]));
Q_ASSIGN U2161 ( .B(R[2161]), .A(L[2161]));
Q_ASSIGN U2162 ( .B(R[2162]), .A(L[2162]));
Q_ASSIGN U2163 ( .B(R[2163]), .A(L[2163]));
Q_ASSIGN U2164 ( .B(R[2164]), .A(L[2164]));
Q_ASSIGN U2165 ( .B(R[2165]), .A(L[2165]));
Q_ASSIGN U2166 ( .B(R[2166]), .A(L[2166]));
Q_ASSIGN U2167 ( .B(R[2167]), .A(L[2167]));
Q_ASSIGN U2168 ( .B(R[2168]), .A(L[2168]));
Q_ASSIGN U2169 ( .B(R[2169]), .A(L[2169]));
Q_ASSIGN U2170 ( .B(R[2170]), .A(L[2170]));
Q_ASSIGN U2171 ( .B(R[2171]), .A(L[2171]));
Q_ASSIGN U2172 ( .B(R[2172]), .A(L[2172]));
Q_ASSIGN U2173 ( .B(R[2173]), .A(L[2173]));
Q_ASSIGN U2174 ( .B(R[2174]), .A(L[2174]));
Q_ASSIGN U2175 ( .B(R[2175]), .A(L[2175]));
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_assign"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
endmodule
