
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_kdf_keyfilter ( keyfilter_cmdfifo_ack, 
	keyfilter_upsizer_stall, hash_key_in, hash_key_in_valid, clk, rst_n, 
	cmdfifo_keyfilter_valid, .cmdfifo_keyfilter_cmd( {
	\cmdfifo_keyfilter_cmd.combo_mode [0]} ), upsizer_keyfilter_data, 
	upsizer_keyfilter_valid, upsizer_keyfilter_eof, hash_key_in_stall);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output keyfilter_cmdfifo_ack;
output keyfilter_upsizer_stall;
output [255:0] hash_key_in;
output hash_key_in_valid;
input clk;
input rst_n;
input cmdfifo_keyfilter_valid;
input [0:0] \cmdfifo_keyfilter_cmd.combo_mode ;
wire [0:0] cmdfifo_keyfilter_cmd;
input [255:0] upsizer_keyfilter_data;
input upsizer_keyfilter_valid;
input upsizer_keyfilter_eof;
input hash_key_in_stall;
wire _zy_simnet_keyfilter_cmdfifo_ack_0_w$;
wire _zy_simnet_keyfilter_upsizer_stall_1_w$;
wire [0:255] _zy_simnet_hash_key_in_2_w$;
wire _zy_simnet_hash_key_in_valid_3_w$;
wire [1:0] counter;
tran (cmdfifo_keyfilter_cmd[0], \cmdfifo_keyfilter_cmd.combo_mode [0]);
ixc_assign _zz_strnp_3 ( _zy_simnet_hash_key_in_valid_3_w$, hash_key_in_valid);
ixc_assign_256 _zz_strnp_2 ( _zy_simnet_hash_key_in_2_w$[0:255], 
	hash_key_in[255:0]);
ixc_assign _zz_strnp_1 ( _zy_simnet_keyfilter_upsizer_stall_1_w$, 
	keyfilter_upsizer_stall);
ixc_assign _zz_strnp_0 ( _zy_simnet_keyfilter_cmdfifo_ack_0_w$, 
	keyfilter_cmdfifo_ack);
Q_AN02 U4 ( .A0(n5), .A1(upsizer_keyfilter_valid), .Z(hash_key_in_valid));
Q_AN02 U5 ( .A0(n5), .A1(upsizer_keyfilter_data[0]), .Z(hash_key_in[0]));
Q_AN02 U6 ( .A0(n5), .A1(upsizer_keyfilter_data[1]), .Z(hash_key_in[1]));
Q_AN02 U7 ( .A0(n5), .A1(upsizer_keyfilter_data[2]), .Z(hash_key_in[2]));
Q_AN02 U8 ( .A0(n5), .A1(upsizer_keyfilter_data[3]), .Z(hash_key_in[3]));
Q_AN02 U9 ( .A0(n5), .A1(upsizer_keyfilter_data[4]), .Z(hash_key_in[4]));
Q_AN02 U10 ( .A0(n5), .A1(upsizer_keyfilter_data[5]), .Z(hash_key_in[5]));
Q_AN02 U11 ( .A0(n5), .A1(upsizer_keyfilter_data[6]), .Z(hash_key_in[6]));
Q_AN02 U12 ( .A0(n5), .A1(upsizer_keyfilter_data[7]), .Z(hash_key_in[7]));
Q_AN02 U13 ( .A0(n5), .A1(upsizer_keyfilter_data[8]), .Z(hash_key_in[8]));
Q_AN02 U14 ( .A0(n5), .A1(upsizer_keyfilter_data[9]), .Z(hash_key_in[9]));
Q_AN02 U15 ( .A0(n5), .A1(upsizer_keyfilter_data[10]), .Z(hash_key_in[10]));
Q_AN02 U16 ( .A0(n5), .A1(upsizer_keyfilter_data[11]), .Z(hash_key_in[11]));
Q_AN02 U17 ( .A0(n5), .A1(upsizer_keyfilter_data[12]), .Z(hash_key_in[12]));
Q_AN02 U18 ( .A0(n5), .A1(upsizer_keyfilter_data[13]), .Z(hash_key_in[13]));
Q_AN02 U19 ( .A0(n5), .A1(upsizer_keyfilter_data[14]), .Z(hash_key_in[14]));
Q_AN02 U20 ( .A0(n5), .A1(upsizer_keyfilter_data[15]), .Z(hash_key_in[15]));
Q_AN02 U21 ( .A0(n5), .A1(upsizer_keyfilter_data[16]), .Z(hash_key_in[16]));
Q_AN02 U22 ( .A0(n5), .A1(upsizer_keyfilter_data[17]), .Z(hash_key_in[17]));
Q_AN02 U23 ( .A0(n5), .A1(upsizer_keyfilter_data[18]), .Z(hash_key_in[18]));
Q_AN02 U24 ( .A0(n5), .A1(upsizer_keyfilter_data[19]), .Z(hash_key_in[19]));
Q_AN02 U25 ( .A0(n5), .A1(upsizer_keyfilter_data[20]), .Z(hash_key_in[20]));
Q_AN02 U26 ( .A0(n5), .A1(upsizer_keyfilter_data[21]), .Z(hash_key_in[21]));
Q_AN02 U27 ( .A0(n5), .A1(upsizer_keyfilter_data[22]), .Z(hash_key_in[22]));
Q_AN02 U28 ( .A0(n5), .A1(upsizer_keyfilter_data[23]), .Z(hash_key_in[23]));
Q_AN02 U29 ( .A0(n5), .A1(upsizer_keyfilter_data[24]), .Z(hash_key_in[24]));
Q_AN02 U30 ( .A0(n5), .A1(upsizer_keyfilter_data[25]), .Z(hash_key_in[25]));
Q_AN02 U31 ( .A0(n5), .A1(upsizer_keyfilter_data[26]), .Z(hash_key_in[26]));
Q_AN02 U32 ( .A0(n5), .A1(upsizer_keyfilter_data[27]), .Z(hash_key_in[27]));
Q_AN02 U33 ( .A0(n5), .A1(upsizer_keyfilter_data[28]), .Z(hash_key_in[28]));
Q_AN02 U34 ( .A0(n5), .A1(upsizer_keyfilter_data[29]), .Z(hash_key_in[29]));
Q_AN02 U35 ( .A0(n5), .A1(upsizer_keyfilter_data[30]), .Z(hash_key_in[30]));
Q_AN02 U36 ( .A0(n5), .A1(upsizer_keyfilter_data[31]), .Z(hash_key_in[31]));
Q_AN02 U37 ( .A0(n5), .A1(upsizer_keyfilter_data[32]), .Z(hash_key_in[32]));
Q_AN02 U38 ( .A0(n5), .A1(upsizer_keyfilter_data[33]), .Z(hash_key_in[33]));
Q_AN02 U39 ( .A0(n5), .A1(upsizer_keyfilter_data[34]), .Z(hash_key_in[34]));
Q_AN02 U40 ( .A0(n5), .A1(upsizer_keyfilter_data[35]), .Z(hash_key_in[35]));
Q_AN02 U41 ( .A0(n5), .A1(upsizer_keyfilter_data[36]), .Z(hash_key_in[36]));
Q_AN02 U42 ( .A0(n5), .A1(upsizer_keyfilter_data[37]), .Z(hash_key_in[37]));
Q_AN02 U43 ( .A0(n5), .A1(upsizer_keyfilter_data[38]), .Z(hash_key_in[38]));
Q_AN02 U44 ( .A0(n5), .A1(upsizer_keyfilter_data[39]), .Z(hash_key_in[39]));
Q_AN02 U45 ( .A0(n5), .A1(upsizer_keyfilter_data[40]), .Z(hash_key_in[40]));
Q_AN02 U46 ( .A0(n5), .A1(upsizer_keyfilter_data[41]), .Z(hash_key_in[41]));
Q_AN02 U47 ( .A0(n5), .A1(upsizer_keyfilter_data[42]), .Z(hash_key_in[42]));
Q_AN02 U48 ( .A0(n5), .A1(upsizer_keyfilter_data[43]), .Z(hash_key_in[43]));
Q_AN02 U49 ( .A0(n5), .A1(upsizer_keyfilter_data[44]), .Z(hash_key_in[44]));
Q_AN02 U50 ( .A0(n5), .A1(upsizer_keyfilter_data[45]), .Z(hash_key_in[45]));
Q_AN02 U51 ( .A0(n5), .A1(upsizer_keyfilter_data[46]), .Z(hash_key_in[46]));
Q_AN02 U52 ( .A0(n5), .A1(upsizer_keyfilter_data[47]), .Z(hash_key_in[47]));
Q_AN02 U53 ( .A0(n5), .A1(upsizer_keyfilter_data[48]), .Z(hash_key_in[48]));
Q_AN02 U54 ( .A0(n5), .A1(upsizer_keyfilter_data[49]), .Z(hash_key_in[49]));
Q_AN02 U55 ( .A0(n5), .A1(upsizer_keyfilter_data[50]), .Z(hash_key_in[50]));
Q_AN02 U56 ( .A0(n5), .A1(upsizer_keyfilter_data[51]), .Z(hash_key_in[51]));
Q_AN02 U57 ( .A0(n5), .A1(upsizer_keyfilter_data[52]), .Z(hash_key_in[52]));
Q_AN02 U58 ( .A0(n5), .A1(upsizer_keyfilter_data[53]), .Z(hash_key_in[53]));
Q_AN02 U59 ( .A0(n5), .A1(upsizer_keyfilter_data[54]), .Z(hash_key_in[54]));
Q_AN02 U60 ( .A0(n5), .A1(upsizer_keyfilter_data[55]), .Z(hash_key_in[55]));
Q_AN02 U61 ( .A0(n5), .A1(upsizer_keyfilter_data[56]), .Z(hash_key_in[56]));
Q_AN02 U62 ( .A0(n5), .A1(upsizer_keyfilter_data[57]), .Z(hash_key_in[57]));
Q_AN02 U63 ( .A0(n5), .A1(upsizer_keyfilter_data[58]), .Z(hash_key_in[58]));
Q_AN02 U64 ( .A0(n5), .A1(upsizer_keyfilter_data[59]), .Z(hash_key_in[59]));
Q_AN02 U65 ( .A0(n5), .A1(upsizer_keyfilter_data[60]), .Z(hash_key_in[60]));
Q_AN02 U66 ( .A0(n5), .A1(upsizer_keyfilter_data[61]), .Z(hash_key_in[61]));
Q_AN02 U67 ( .A0(n5), .A1(upsizer_keyfilter_data[62]), .Z(hash_key_in[62]));
Q_AN02 U68 ( .A0(n5), .A1(upsizer_keyfilter_data[63]), .Z(hash_key_in[63]));
Q_AN02 U69 ( .A0(n5), .A1(upsizer_keyfilter_data[64]), .Z(hash_key_in[64]));
Q_AN02 U70 ( .A0(n5), .A1(upsizer_keyfilter_data[65]), .Z(hash_key_in[65]));
Q_AN02 U71 ( .A0(n5), .A1(upsizer_keyfilter_data[66]), .Z(hash_key_in[66]));
Q_AN02 U72 ( .A0(n5), .A1(upsizer_keyfilter_data[67]), .Z(hash_key_in[67]));
Q_AN02 U73 ( .A0(n5), .A1(upsizer_keyfilter_data[68]), .Z(hash_key_in[68]));
Q_AN02 U74 ( .A0(n5), .A1(upsizer_keyfilter_data[69]), .Z(hash_key_in[69]));
Q_AN02 U75 ( .A0(n5), .A1(upsizer_keyfilter_data[70]), .Z(hash_key_in[70]));
Q_AN02 U76 ( .A0(n5), .A1(upsizer_keyfilter_data[71]), .Z(hash_key_in[71]));
Q_AN02 U77 ( .A0(n5), .A1(upsizer_keyfilter_data[72]), .Z(hash_key_in[72]));
Q_AN02 U78 ( .A0(n5), .A1(upsizer_keyfilter_data[73]), .Z(hash_key_in[73]));
Q_AN02 U79 ( .A0(n5), .A1(upsizer_keyfilter_data[74]), .Z(hash_key_in[74]));
Q_AN02 U80 ( .A0(n5), .A1(upsizer_keyfilter_data[75]), .Z(hash_key_in[75]));
Q_AN02 U81 ( .A0(n5), .A1(upsizer_keyfilter_data[76]), .Z(hash_key_in[76]));
Q_AN02 U82 ( .A0(n5), .A1(upsizer_keyfilter_data[77]), .Z(hash_key_in[77]));
Q_AN02 U83 ( .A0(n5), .A1(upsizer_keyfilter_data[78]), .Z(hash_key_in[78]));
Q_AN02 U84 ( .A0(n5), .A1(upsizer_keyfilter_data[79]), .Z(hash_key_in[79]));
Q_AN02 U85 ( .A0(n5), .A1(upsizer_keyfilter_data[80]), .Z(hash_key_in[80]));
Q_AN02 U86 ( .A0(n5), .A1(upsizer_keyfilter_data[81]), .Z(hash_key_in[81]));
Q_AN02 U87 ( .A0(n5), .A1(upsizer_keyfilter_data[82]), .Z(hash_key_in[82]));
Q_AN02 U88 ( .A0(n5), .A1(upsizer_keyfilter_data[83]), .Z(hash_key_in[83]));
Q_AN02 U89 ( .A0(n5), .A1(upsizer_keyfilter_data[84]), .Z(hash_key_in[84]));
Q_AN02 U90 ( .A0(n5), .A1(upsizer_keyfilter_data[85]), .Z(hash_key_in[85]));
Q_AN02 U91 ( .A0(n5), .A1(upsizer_keyfilter_data[86]), .Z(hash_key_in[86]));
Q_AN02 U92 ( .A0(n5), .A1(upsizer_keyfilter_data[87]), .Z(hash_key_in[87]));
Q_AN02 U93 ( .A0(n5), .A1(upsizer_keyfilter_data[88]), .Z(hash_key_in[88]));
Q_AN02 U94 ( .A0(n5), .A1(upsizer_keyfilter_data[89]), .Z(hash_key_in[89]));
Q_AN02 U95 ( .A0(n5), .A1(upsizer_keyfilter_data[90]), .Z(hash_key_in[90]));
Q_AN02 U96 ( .A0(n5), .A1(upsizer_keyfilter_data[91]), .Z(hash_key_in[91]));
Q_AN02 U97 ( .A0(n5), .A1(upsizer_keyfilter_data[92]), .Z(hash_key_in[92]));
Q_AN02 U98 ( .A0(n5), .A1(upsizer_keyfilter_data[93]), .Z(hash_key_in[93]));
Q_AN02 U99 ( .A0(n5), .A1(upsizer_keyfilter_data[94]), .Z(hash_key_in[94]));
Q_AN02 U100 ( .A0(n5), .A1(upsizer_keyfilter_data[95]), .Z(hash_key_in[95]));
Q_AN02 U101 ( .A0(n5), .A1(upsizer_keyfilter_data[96]), .Z(hash_key_in[96]));
Q_AN02 U102 ( .A0(n5), .A1(upsizer_keyfilter_data[97]), .Z(hash_key_in[97]));
Q_AN02 U103 ( .A0(n5), .A1(upsizer_keyfilter_data[98]), .Z(hash_key_in[98]));
Q_AN02 U104 ( .A0(n5), .A1(upsizer_keyfilter_data[99]), .Z(hash_key_in[99]));
Q_AN02 U105 ( .A0(n5), .A1(upsizer_keyfilter_data[100]), .Z(hash_key_in[100]));
Q_AN02 U106 ( .A0(n5), .A1(upsizer_keyfilter_data[101]), .Z(hash_key_in[101]));
Q_AN02 U107 ( .A0(n5), .A1(upsizer_keyfilter_data[102]), .Z(hash_key_in[102]));
Q_AN02 U108 ( .A0(n5), .A1(upsizer_keyfilter_data[103]), .Z(hash_key_in[103]));
Q_AN02 U109 ( .A0(n5), .A1(upsizer_keyfilter_data[104]), .Z(hash_key_in[104]));
Q_AN02 U110 ( .A0(n5), .A1(upsizer_keyfilter_data[105]), .Z(hash_key_in[105]));
Q_AN02 U111 ( .A0(n5), .A1(upsizer_keyfilter_data[106]), .Z(hash_key_in[106]));
Q_AN02 U112 ( .A0(n5), .A1(upsizer_keyfilter_data[107]), .Z(hash_key_in[107]));
Q_AN02 U113 ( .A0(n5), .A1(upsizer_keyfilter_data[108]), .Z(hash_key_in[108]));
Q_AN02 U114 ( .A0(n5), .A1(upsizer_keyfilter_data[109]), .Z(hash_key_in[109]));
Q_AN02 U115 ( .A0(n5), .A1(upsizer_keyfilter_data[110]), .Z(hash_key_in[110]));
Q_AN02 U116 ( .A0(n5), .A1(upsizer_keyfilter_data[111]), .Z(hash_key_in[111]));
Q_AN02 U117 ( .A0(n5), .A1(upsizer_keyfilter_data[112]), .Z(hash_key_in[112]));
Q_AN02 U118 ( .A0(n5), .A1(upsizer_keyfilter_data[113]), .Z(hash_key_in[113]));
Q_AN02 U119 ( .A0(n5), .A1(upsizer_keyfilter_data[114]), .Z(hash_key_in[114]));
Q_AN02 U120 ( .A0(n5), .A1(upsizer_keyfilter_data[115]), .Z(hash_key_in[115]));
Q_AN02 U121 ( .A0(n5), .A1(upsizer_keyfilter_data[116]), .Z(hash_key_in[116]));
Q_AN02 U122 ( .A0(n5), .A1(upsizer_keyfilter_data[117]), .Z(hash_key_in[117]));
Q_AN02 U123 ( .A0(n5), .A1(upsizer_keyfilter_data[118]), .Z(hash_key_in[118]));
Q_AN02 U124 ( .A0(n5), .A1(upsizer_keyfilter_data[119]), .Z(hash_key_in[119]));
Q_AN02 U125 ( .A0(n5), .A1(upsizer_keyfilter_data[120]), .Z(hash_key_in[120]));
Q_AN02 U126 ( .A0(n5), .A1(upsizer_keyfilter_data[121]), .Z(hash_key_in[121]));
Q_AN02 U127 ( .A0(n5), .A1(upsizer_keyfilter_data[122]), .Z(hash_key_in[122]));
Q_AN02 U128 ( .A0(n5), .A1(upsizer_keyfilter_data[123]), .Z(hash_key_in[123]));
Q_AN02 U129 ( .A0(n5), .A1(upsizer_keyfilter_data[124]), .Z(hash_key_in[124]));
Q_AN02 U130 ( .A0(n5), .A1(upsizer_keyfilter_data[125]), .Z(hash_key_in[125]));
Q_AN02 U131 ( .A0(n5), .A1(upsizer_keyfilter_data[126]), .Z(hash_key_in[126]));
Q_AN02 U132 ( .A0(n5), .A1(upsizer_keyfilter_data[127]), .Z(hash_key_in[127]));
Q_AN02 U133 ( .A0(n5), .A1(upsizer_keyfilter_data[128]), .Z(hash_key_in[128]));
Q_AN02 U134 ( .A0(n5), .A1(upsizer_keyfilter_data[129]), .Z(hash_key_in[129]));
Q_AN02 U135 ( .A0(n5), .A1(upsizer_keyfilter_data[130]), .Z(hash_key_in[130]));
Q_AN02 U136 ( .A0(n5), .A1(upsizer_keyfilter_data[131]), .Z(hash_key_in[131]));
Q_AN02 U137 ( .A0(n5), .A1(upsizer_keyfilter_data[132]), .Z(hash_key_in[132]));
Q_AN02 U138 ( .A0(n5), .A1(upsizer_keyfilter_data[133]), .Z(hash_key_in[133]));
Q_AN02 U139 ( .A0(n5), .A1(upsizer_keyfilter_data[134]), .Z(hash_key_in[134]));
Q_AN02 U140 ( .A0(n5), .A1(upsizer_keyfilter_data[135]), .Z(hash_key_in[135]));
Q_AN02 U141 ( .A0(n5), .A1(upsizer_keyfilter_data[136]), .Z(hash_key_in[136]));
Q_AN02 U142 ( .A0(n5), .A1(upsizer_keyfilter_data[137]), .Z(hash_key_in[137]));
Q_AN02 U143 ( .A0(n5), .A1(upsizer_keyfilter_data[138]), .Z(hash_key_in[138]));
Q_AN02 U144 ( .A0(n5), .A1(upsizer_keyfilter_data[139]), .Z(hash_key_in[139]));
Q_AN02 U145 ( .A0(n5), .A1(upsizer_keyfilter_data[140]), .Z(hash_key_in[140]));
Q_AN02 U146 ( .A0(n5), .A1(upsizer_keyfilter_data[141]), .Z(hash_key_in[141]));
Q_AN02 U147 ( .A0(n5), .A1(upsizer_keyfilter_data[142]), .Z(hash_key_in[142]));
Q_AN02 U148 ( .A0(n5), .A1(upsizer_keyfilter_data[143]), .Z(hash_key_in[143]));
Q_AN02 U149 ( .A0(n5), .A1(upsizer_keyfilter_data[144]), .Z(hash_key_in[144]));
Q_AN02 U150 ( .A0(n5), .A1(upsizer_keyfilter_data[145]), .Z(hash_key_in[145]));
Q_AN02 U151 ( .A0(n5), .A1(upsizer_keyfilter_data[146]), .Z(hash_key_in[146]));
Q_AN02 U152 ( .A0(n5), .A1(upsizer_keyfilter_data[147]), .Z(hash_key_in[147]));
Q_AN02 U153 ( .A0(n5), .A1(upsizer_keyfilter_data[148]), .Z(hash_key_in[148]));
Q_AN02 U154 ( .A0(n5), .A1(upsizer_keyfilter_data[149]), .Z(hash_key_in[149]));
Q_AN02 U155 ( .A0(n5), .A1(upsizer_keyfilter_data[150]), .Z(hash_key_in[150]));
Q_AN02 U156 ( .A0(n5), .A1(upsizer_keyfilter_data[151]), .Z(hash_key_in[151]));
Q_AN02 U157 ( .A0(n5), .A1(upsizer_keyfilter_data[152]), .Z(hash_key_in[152]));
Q_AN02 U158 ( .A0(n5), .A1(upsizer_keyfilter_data[153]), .Z(hash_key_in[153]));
Q_AN02 U159 ( .A0(n5), .A1(upsizer_keyfilter_data[154]), .Z(hash_key_in[154]));
Q_AN02 U160 ( .A0(n5), .A1(upsizer_keyfilter_data[155]), .Z(hash_key_in[155]));
Q_AN02 U161 ( .A0(n5), .A1(upsizer_keyfilter_data[156]), .Z(hash_key_in[156]));
Q_AN02 U162 ( .A0(n5), .A1(upsizer_keyfilter_data[157]), .Z(hash_key_in[157]));
Q_AN02 U163 ( .A0(n5), .A1(upsizer_keyfilter_data[158]), .Z(hash_key_in[158]));
Q_AN02 U164 ( .A0(n5), .A1(upsizer_keyfilter_data[159]), .Z(hash_key_in[159]));
Q_AN02 U165 ( .A0(n5), .A1(upsizer_keyfilter_data[160]), .Z(hash_key_in[160]));
Q_AN02 U166 ( .A0(n5), .A1(upsizer_keyfilter_data[161]), .Z(hash_key_in[161]));
Q_AN02 U167 ( .A0(n5), .A1(upsizer_keyfilter_data[162]), .Z(hash_key_in[162]));
Q_AN02 U168 ( .A0(n5), .A1(upsizer_keyfilter_data[163]), .Z(hash_key_in[163]));
Q_AN02 U169 ( .A0(n5), .A1(upsizer_keyfilter_data[164]), .Z(hash_key_in[164]));
Q_AN02 U170 ( .A0(n5), .A1(upsizer_keyfilter_data[165]), .Z(hash_key_in[165]));
Q_AN02 U171 ( .A0(n5), .A1(upsizer_keyfilter_data[166]), .Z(hash_key_in[166]));
Q_AN02 U172 ( .A0(n5), .A1(upsizer_keyfilter_data[167]), .Z(hash_key_in[167]));
Q_AN02 U173 ( .A0(n5), .A1(upsizer_keyfilter_data[168]), .Z(hash_key_in[168]));
Q_AN02 U174 ( .A0(n5), .A1(upsizer_keyfilter_data[169]), .Z(hash_key_in[169]));
Q_AN02 U175 ( .A0(n5), .A1(upsizer_keyfilter_data[170]), .Z(hash_key_in[170]));
Q_AN02 U176 ( .A0(n5), .A1(upsizer_keyfilter_data[171]), .Z(hash_key_in[171]));
Q_AN02 U177 ( .A0(n5), .A1(upsizer_keyfilter_data[172]), .Z(hash_key_in[172]));
Q_AN02 U178 ( .A0(n5), .A1(upsizer_keyfilter_data[173]), .Z(hash_key_in[173]));
Q_AN02 U179 ( .A0(n5), .A1(upsizer_keyfilter_data[174]), .Z(hash_key_in[174]));
Q_AN02 U180 ( .A0(n5), .A1(upsizer_keyfilter_data[175]), .Z(hash_key_in[175]));
Q_AN02 U181 ( .A0(n5), .A1(upsizer_keyfilter_data[176]), .Z(hash_key_in[176]));
Q_AN02 U182 ( .A0(n5), .A1(upsizer_keyfilter_data[177]), .Z(hash_key_in[177]));
Q_AN02 U183 ( .A0(n5), .A1(upsizer_keyfilter_data[178]), .Z(hash_key_in[178]));
Q_AN02 U184 ( .A0(n5), .A1(upsizer_keyfilter_data[179]), .Z(hash_key_in[179]));
Q_AN02 U185 ( .A0(n5), .A1(upsizer_keyfilter_data[180]), .Z(hash_key_in[180]));
Q_AN02 U186 ( .A0(n5), .A1(upsizer_keyfilter_data[181]), .Z(hash_key_in[181]));
Q_AN02 U187 ( .A0(n5), .A1(upsizer_keyfilter_data[182]), .Z(hash_key_in[182]));
Q_AN02 U188 ( .A0(n5), .A1(upsizer_keyfilter_data[183]), .Z(hash_key_in[183]));
Q_AN02 U189 ( .A0(n5), .A1(upsizer_keyfilter_data[184]), .Z(hash_key_in[184]));
Q_AN02 U190 ( .A0(n5), .A1(upsizer_keyfilter_data[185]), .Z(hash_key_in[185]));
Q_AN02 U191 ( .A0(n5), .A1(upsizer_keyfilter_data[186]), .Z(hash_key_in[186]));
Q_AN02 U192 ( .A0(n5), .A1(upsizer_keyfilter_data[187]), .Z(hash_key_in[187]));
Q_AN02 U193 ( .A0(n5), .A1(upsizer_keyfilter_data[188]), .Z(hash_key_in[188]));
Q_AN02 U194 ( .A0(n5), .A1(upsizer_keyfilter_data[189]), .Z(hash_key_in[189]));
Q_AN02 U195 ( .A0(n5), .A1(upsizer_keyfilter_data[190]), .Z(hash_key_in[190]));
Q_AN02 U196 ( .A0(n5), .A1(upsizer_keyfilter_data[191]), .Z(hash_key_in[191]));
Q_AN02 U197 ( .A0(n5), .A1(upsizer_keyfilter_data[192]), .Z(hash_key_in[192]));
Q_AN02 U198 ( .A0(n5), .A1(upsizer_keyfilter_data[193]), .Z(hash_key_in[193]));
Q_AN02 U199 ( .A0(n5), .A1(upsizer_keyfilter_data[194]), .Z(hash_key_in[194]));
Q_AN02 U200 ( .A0(n5), .A1(upsizer_keyfilter_data[195]), .Z(hash_key_in[195]));
Q_AN02 U201 ( .A0(n5), .A1(upsizer_keyfilter_data[196]), .Z(hash_key_in[196]));
Q_AN02 U202 ( .A0(n5), .A1(upsizer_keyfilter_data[197]), .Z(hash_key_in[197]));
Q_AN02 U203 ( .A0(n5), .A1(upsizer_keyfilter_data[198]), .Z(hash_key_in[198]));
Q_AN02 U204 ( .A0(n5), .A1(upsizer_keyfilter_data[199]), .Z(hash_key_in[199]));
Q_AN02 U205 ( .A0(n5), .A1(upsizer_keyfilter_data[200]), .Z(hash_key_in[200]));
Q_AN02 U206 ( .A0(n5), .A1(upsizer_keyfilter_data[201]), .Z(hash_key_in[201]));
Q_AN02 U207 ( .A0(n5), .A1(upsizer_keyfilter_data[202]), .Z(hash_key_in[202]));
Q_AN02 U208 ( .A0(n5), .A1(upsizer_keyfilter_data[203]), .Z(hash_key_in[203]));
Q_AN02 U209 ( .A0(n5), .A1(upsizer_keyfilter_data[204]), .Z(hash_key_in[204]));
Q_AN02 U210 ( .A0(n5), .A1(upsizer_keyfilter_data[205]), .Z(hash_key_in[205]));
Q_AN02 U211 ( .A0(n5), .A1(upsizer_keyfilter_data[206]), .Z(hash_key_in[206]));
Q_AN02 U212 ( .A0(n5), .A1(upsizer_keyfilter_data[207]), .Z(hash_key_in[207]));
Q_AN02 U213 ( .A0(n5), .A1(upsizer_keyfilter_data[208]), .Z(hash_key_in[208]));
Q_AN02 U214 ( .A0(n5), .A1(upsizer_keyfilter_data[209]), .Z(hash_key_in[209]));
Q_AN02 U215 ( .A0(n5), .A1(upsizer_keyfilter_data[210]), .Z(hash_key_in[210]));
Q_AN02 U216 ( .A0(n5), .A1(upsizer_keyfilter_data[211]), .Z(hash_key_in[211]));
Q_AN02 U217 ( .A0(n5), .A1(upsizer_keyfilter_data[212]), .Z(hash_key_in[212]));
Q_AN02 U218 ( .A0(n5), .A1(upsizer_keyfilter_data[213]), .Z(hash_key_in[213]));
Q_AN02 U219 ( .A0(n5), .A1(upsizer_keyfilter_data[214]), .Z(hash_key_in[214]));
Q_AN02 U220 ( .A0(n5), .A1(upsizer_keyfilter_data[215]), .Z(hash_key_in[215]));
Q_AN02 U221 ( .A0(n5), .A1(upsizer_keyfilter_data[216]), .Z(hash_key_in[216]));
Q_AN02 U222 ( .A0(n5), .A1(upsizer_keyfilter_data[217]), .Z(hash_key_in[217]));
Q_AN02 U223 ( .A0(n5), .A1(upsizer_keyfilter_data[218]), .Z(hash_key_in[218]));
Q_AN02 U224 ( .A0(n5), .A1(upsizer_keyfilter_data[219]), .Z(hash_key_in[219]));
Q_AN02 U225 ( .A0(n5), .A1(upsizer_keyfilter_data[220]), .Z(hash_key_in[220]));
Q_AN02 U226 ( .A0(n5), .A1(upsizer_keyfilter_data[221]), .Z(hash_key_in[221]));
Q_AN02 U227 ( .A0(n5), .A1(upsizer_keyfilter_data[222]), .Z(hash_key_in[222]));
Q_AN02 U228 ( .A0(n5), .A1(upsizer_keyfilter_data[223]), .Z(hash_key_in[223]));
Q_AN02 U229 ( .A0(n5), .A1(upsizer_keyfilter_data[224]), .Z(hash_key_in[224]));
Q_AN02 U230 ( .A0(n5), .A1(upsizer_keyfilter_data[225]), .Z(hash_key_in[225]));
Q_AN02 U231 ( .A0(n5), .A1(upsizer_keyfilter_data[226]), .Z(hash_key_in[226]));
Q_AN02 U232 ( .A0(n5), .A1(upsizer_keyfilter_data[227]), .Z(hash_key_in[227]));
Q_AN02 U233 ( .A0(n5), .A1(upsizer_keyfilter_data[228]), .Z(hash_key_in[228]));
Q_AN02 U234 ( .A0(n5), .A1(upsizer_keyfilter_data[229]), .Z(hash_key_in[229]));
Q_AN02 U235 ( .A0(n5), .A1(upsizer_keyfilter_data[230]), .Z(hash_key_in[230]));
Q_AN02 U236 ( .A0(n5), .A1(upsizer_keyfilter_data[231]), .Z(hash_key_in[231]));
Q_AN02 U237 ( .A0(n5), .A1(upsizer_keyfilter_data[232]), .Z(hash_key_in[232]));
Q_AN02 U238 ( .A0(n5), .A1(upsizer_keyfilter_data[233]), .Z(hash_key_in[233]));
Q_AN02 U239 ( .A0(n5), .A1(upsizer_keyfilter_data[234]), .Z(hash_key_in[234]));
Q_AN02 U240 ( .A0(n5), .A1(upsizer_keyfilter_data[235]), .Z(hash_key_in[235]));
Q_AN02 U241 ( .A0(n5), .A1(upsizer_keyfilter_data[236]), .Z(hash_key_in[236]));
Q_AN02 U242 ( .A0(n5), .A1(upsizer_keyfilter_data[237]), .Z(hash_key_in[237]));
Q_AN02 U243 ( .A0(n5), .A1(upsizer_keyfilter_data[238]), .Z(hash_key_in[238]));
Q_AN02 U244 ( .A0(n5), .A1(upsizer_keyfilter_data[239]), .Z(hash_key_in[239]));
Q_AN02 U245 ( .A0(n5), .A1(upsizer_keyfilter_data[240]), .Z(hash_key_in[240]));
Q_AN02 U246 ( .A0(n5), .A1(upsizer_keyfilter_data[241]), .Z(hash_key_in[241]));
Q_AN02 U247 ( .A0(n5), .A1(upsizer_keyfilter_data[242]), .Z(hash_key_in[242]));
Q_AN02 U248 ( .A0(n5), .A1(upsizer_keyfilter_data[243]), .Z(hash_key_in[243]));
Q_AN02 U249 ( .A0(n5), .A1(upsizer_keyfilter_data[244]), .Z(hash_key_in[244]));
Q_AN02 U250 ( .A0(n5), .A1(upsizer_keyfilter_data[245]), .Z(hash_key_in[245]));
Q_AN02 U251 ( .A0(n5), .A1(upsizer_keyfilter_data[246]), .Z(hash_key_in[246]));
Q_AN02 U252 ( .A0(n5), .A1(upsizer_keyfilter_data[247]), .Z(hash_key_in[247]));
Q_AN02 U253 ( .A0(n5), .A1(upsizer_keyfilter_data[248]), .Z(hash_key_in[248]));
Q_AN02 U254 ( .A0(n5), .A1(upsizer_keyfilter_data[249]), .Z(hash_key_in[249]));
Q_AN02 U255 ( .A0(n5), .A1(upsizer_keyfilter_data[250]), .Z(hash_key_in[250]));
Q_AN02 U256 ( .A0(n5), .A1(upsizer_keyfilter_data[251]), .Z(hash_key_in[251]));
Q_AN02 U257 ( .A0(n5), .A1(upsizer_keyfilter_data[252]), .Z(hash_key_in[252]));
Q_AN02 U258 ( .A0(n5), .A1(upsizer_keyfilter_data[253]), .Z(hash_key_in[253]));
Q_AN02 U259 ( .A0(n5), .A1(upsizer_keyfilter_data[254]), .Z(hash_key_in[254]));
Q_AN02 U260 ( .A0(n5), .A1(upsizer_keyfilter_data[255]), .Z(hash_key_in[255]));
Q_AN02 U261 ( .A0(n5), .A1(hash_key_in_stall), .Z(keyfilter_upsizer_stall));
Q_AN02 U262 ( .A0(n6), .A1(upsizer_keyfilter_valid), .Z(keyfilter_cmdfifo_ack));
Q_AN02 U263 ( .A0(n6), .A1(n2), .Z(n1));
Q_INV U264 ( .A(cmdfifo_keyfilter_cmd[0]), .Z(n2));
Q_AO21 U265 ( .A0(n3), .A1(counter[0]), .B0(n1), .Z(n5));
Q_AN02 U266 ( .A0(counter[1]), .A1(n4), .Z(n6));
Q_XOR2 U267 ( .A0(counter[1]), .A1(counter[0]), .Z(n7));
Q_NR02 U268 ( .A0(n6), .A1(counter[0]), .Z(n8));
Q_AN02 U269 ( .A0(n10), .A1(n7), .Z(n9));
Q_INV U270 ( .A(n6), .Z(n10));
Q_FDP4EP \counter_REG[0] ( .CK(clk), .CE(upsizer_keyfilter_valid), .R(n11), .D(n8), .Q(counter[0]));
Q_INV U272 ( .A(rst_n), .Z(n11));
Q_INV U273 ( .A(counter[0]), .Z(n4));
Q_FDP4EP \counter_REG[1] ( .CK(clk), .CE(upsizer_keyfilter_valid), .R(n11), .D(n9), .Q(counter[1]));
Q_INV U275 ( .A(counter[1]), .Z(n3));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\cmdfifo_keyfilter_cmd.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "cmdfifo_keyfilter_cmd 1 \cmdfifo_keyfilter_cmd.combo_mode "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "1"
endmodule
