// xc_work/v/23.sv
// /home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v:20
// NOTE: This file corresponds to a module in the Hardware/DUT partition.
`timescale 1ns/1ns
module cr_kme_tlv_parser(stitcher_rd,parser_kimreader_valid,parser_kimreader_data,tlv_parser_idle,tlv_parser_int_tlv_start_pulse,clk,rst_n,disable_debug_cmd_q,always_validate_kim_ref,stitcher_out,
stitcher_empty,kimreader_parser_ack);
// pkg external : PKG - cr_kme_regfilePKG : DTYPE  
// pragma multiple_driver_resolution
typedef enum logic [1:0] {ENET=0,IPV4=1,IPV6=2,MPLS=3} pkt_hdr_e;
typedef enum logic [3:0] {CMD_SIMPLE=0,COMPND_4K=5,COMPND_8K=6,COMPND_RSV=15} cmd_compound_cmd_frm_size_e;
typedef enum logic [0:0] {GUID_NOT_PRESENT=0,GUID_PRESENT=1} cmd_guid_present_e;
typedef enum logic [0:0] {CRC_NOT_PRESENT=0,CRC_PRESENT=1} cmd_frmd_crc_in_e;
typedef enum logic [6:0] {CCEIP_FRMD_USER_NULL=11,CCEIP_FRMD_USER_PI16=12,CCEIP_FRMD_USER_PI64=13,CCEIP_FRMD_USER_VM=14,CCEIP_TYPE_IN_RSV=127} cceip_cmd_frmd_in_type_e;
typedef enum logic [6:0] {CDDIP_FRMD_INT_APP=15,CDDIP_FRMD_INT_SIP=16,CDDIP_FRMD_INT_LIP=17,CDDIP_FRMD_INT_VM=18,CDDIP_FRMD_INT_VM_SHORT=22,CDDIP_TYPE_IN_RSV=127} cddip_cmd_frmd_in_type_e;
typedef enum logic [6:0] {CCEIP_FRMD_INT_APP=15,CCEIP_FRMD_INT_SIP=16,CCEIP_FRMD_INT_LIP=17,CCEIP_FRMD_INT_VM=18,CCEIP_FRMD_INT_VM_SHORT=22,CCEIP_TYPE_OUT_RSV=127} cceip_cmd_frmd_out_type_e;
typedef enum logic [6:0] {CDDIP_FRMD_USER_NULL=11,CDDIP_FRMD_USER_PI16=12,CDDIP_FRMD_USER_PI64=13,CDDIP_FRMD_USER_VM=14,CDDIP_TYPE_OUT_RSV=127} cddip_cmd_frmd_out_type_e;
typedef enum logic [0:0] {NOT_GEN=0,GEN=1} cmd_frmd_out_crc_e;
typedef enum logic [1:0] {FRMD_T10_DIX=0,FRMD_CRC64=1,FRMD_CRC64E=2,FRMD_CRC_RSV=3} cmd_frmd_out_crc_type_e;
typedef enum logic [1:0] {NO_CRC=0,CRC_8B_CRC64=1,CRC_8B_CRC64E=2,MD_TYPE_RSV=3} cmd_md_type_e;
typedef enum logic [1:0] {CRC_GEN_VERIFY=0,CRC_RSV1=1,CRC_RSV2=2,CRC_RSV3=3} cmd_md_op_e;
typedef enum logic [0:0] {FRMD_MAC_NOP=0,FRMD_MAC_CAL=1} cmd_frmd_raw_mac_sel_e;
typedef enum logic [0:0] {CHU_NORMAL=0,CHU_APPEND=1} cmd_chu_append_e;
typedef enum logic [3:0] {NONE=0,ZLIB=1,GZIP=2,XP9=3,XP10=4,CHU4K=5,CHU8K=6,RSV_MODE=15} cmd_comp_mode_e;
typedef enum logic [3:0] {WIN_32B=0,WIN_4K=1,WIN_8K=2,WIN_16K=3,WIN_32K=4,WIN_64K=5,RSV_WIN=15} cmd_lz77_win_size_e;
typedef enum logic [1:0] {NO_MATCH=0,CHAR_1=1,CHAR_2=2,RSV_DLY=3} cmd_lz77_dly_match_win_e;
typedef enum logic [0:0] {CHAR_3=0,CHAR_4=1} cmd_lz77_min_match_len_e;
typedef enum logic [1:0] {LEN_LZ77_WIN=0,LEN_256B=1,MIN_MTCH_14=2,LEN_64B=3} cmd_lz77_max_symb_len_e;
typedef enum logic [1:0] {NO_PREFIX=0,USER_PREFIX=1,PREDEF_PREFIX=2,PREDET_HUFF=3} cmd_xp10_prefix_mode_e;
typedef enum logic [0:0] {CRC32=0,CRC64=1} cmd_xp10_crc_mode_e;
typedef enum logic [1:0] {FRM=0,FRM_LESS_16=1,INF=2,RSV_THRSH=3} cmd_chu_comp_thrsh_e;
typedef enum logic [0:0] {NO_CIPHER=0,CIPHER=1} cmd_cipher_mode_e;
typedef enum logic [3:0] {AUTH_NULL=0,SHA2=1,HMAC_SHA2=2,AUTH_RSVD=15} cmd_auth_op_e;
typedef enum logic [3:0] {CPH_NULL=0,AES_GCM=1,AES_XTS_XEX=2,AES_GMAC=3,CPH_RSVD=15} cmd_cipher_op_e;
typedef enum logic [1:0] {IV_NONE=0,IV_AUX_CMD=1,IV_KEYS=2,IV_AUX_FRMD=3} cmd_iv_src_e;
typedef enum logic [1:0] {IV_SRC=0,IV_RND=1,IV_INC=2,IV_RSV=3} cmd_iv_op_e;
typedef enum logic [0:0] {NO_PAD=0,PAD_16B=1} cmd_cipher_pad_e;
typedef enum logic [0:0] {DGST_256=0,DGST_64=1} cmd_digest_size_e;
typedef enum logic [0:0] {SIMPLE=0,COMPOUND=1} rqe_frame_type_e;
typedef enum logic [0:0] {TRACE_OFF=0,TRACE_ON=1} rqe_trace_e;
typedef enum logic [3:0] {RQE_SIMPLE=0,RQE_COMPOUND_4K=5,RQE_COMPOUND_8K=6,RQE_RSV_FRAME_SIZE=15} rqe_frame_size_e;
typedef enum logic [1:0] {PARSEABLE=0,RAW=1,XP10CFH4K=2,XP10CFH8K=3} frmd_coding_e;
typedef enum logic [1:0] {DIGEST_64b=0,DIGEST_128b=1,DIGEST_256b=2,DIGEST_0b=3} frmd_mac_size_e;
typedef enum logic [7:0] {RQE=0,CMD=1,KEY=2,PHD=3,PFD=4,DATA_UNK=5,FTR=6,LZ77=7,STAT=8,CQE=9,
GUID=10,FRMD_USER_NULL=11,FRMD_USER_PI16=12,FRMD_USER_PI64=13,FRMD_USER_VM=14,FRMD_INT_APP=15,FRMD_INT_SIP=16,FRMD_INT_LIP=17,FRMD_INT_VM=18,DATA=19,
CR_IV=20,AUX_CMD=21,FRMD_INT_VM_SHORT=22,AUX_CMD_IV=23,AUX_CMD_GUID=24,AUX_CMD_GUID_IV=25,SCH=26,RSV_TLV=255} tlv_types_e;
typedef enum logic [1:0] {REP=0,PASS=1,MODIFY=2,DELETE=3} tlv_parse_action_e;
typedef enum logic [0:0] {USER=0,TLVP=1} tlvp_corrupt_e;
typedef enum logic [0:0] {DATAPATH_CORRUPT=0,FUNCTIONAL_ERROR=1} cmd_type_e;
typedef enum logic [1:0] {SINGLE_ERR=0,CONTINUOUS_ERROR=1,STOP=2,EOT=3} cmd_mode_e;
typedef enum logic [5:0] {NO_AUX_KEY=0,AUX_KEY_ONLY=1,DEK256=2,DEK512=3,DAK=4,DEK256_DAK=5,DEK512_DAK=6,ENC_DEK256=7,ENC_DEK512=8,ENC_DAK=9,
ENC_DEK256_DAK=10,ENC_DEK512_DAK=11,ENC_DEK256_DAK_COMB=12,ENC_DEK512_DAK_COMB=13,KEY_TYPE_RSV=63} aux_key_type_e;
typedef enum logic [0:0] {NOOP=0,KDF=1} aux_key_op_e;
typedef enum logic [1:0] {KDF_MODE_GUID=0,KDF_MODE_RGUID=1,KDF_MODE_COMB_GUID=2,KDF_MODE_COMB_RGUID=3} aux_kdf_mode_e;
typedef enum logic [9:0] {CKMIC_IV_MISMATCH_FRAME=0,CKMIC_ENGINE_ID_MISMATCH_FRAME=1,CKMIC_SEQ_ID_MISMATCH_FRAME=2,CKMIC_HMAC_SHA256_TAG_FAIL_FRAME=3,CKMIC_SHA256_TAG_FAIL_FRAME=4,CKMIC_GMAC_TAG_FAIL_FRAME=5,CKMIC_GCM_TAG_FAIL_FRAME=6,CKMIC_AUTH_NOP_FRAME=7,CKMIC_AUTH_HMAC_SHA256_FRAME=8,CKMIC_AUTH_SHA256_FRAME=9,
CKMIC_AUTH_AES_GMAC_FRAME=10,CKMIC_CIPH_NOP_FRAME=11,CKMIC_CIPH_AES_XEX_FRAME=12,CKMIC_CIPH_AES_XTS_FRAME=13,CKMIC_CIPH_AES_GCM_FRAME=14,CRCG0_RAW_CHSUM_GOOD_TOTAL=64,CRCG0_RAW_CHSUM_ERROR_TOTAL=65,CRCG0_CRC64E_CHSUM_GOOD_TOTAL=66,CRCG0_CRC64E_CHSUM_ERROR_TOTAL=67,CRCG0_ENC_CHSUM_GOOD_TOTAL=68,
CRCG0_ENC_CHSUM_ERROR_TOTAL=69,CRCG0_NVME_CHSUM_GOOD_TOTAL=70,CRCG0_NVME_CHSUM_ERROR_TOTAL=71,CRCGC0_RAW_CHSUM_GOOD_TOTAL=72,CRCGC0_RAW_CHSUM_ERROR_TOTAL=73,CRCGC0_CRC64E_CHSUM_GOOD_TOTAL=74,CRCGC0_CRC64E_CHSUM_ERROR_TOTAL=75,CRCGC0_ENC_CHSUM_GOOD_TOTAL=76,CRCGC0_ENC_CHSUM_ERROR_TOTAL=77,CRCGC0_NVME_CHSUM_GOOD_TOTAL=78,
CRCGC0_NVME_CHSUM_ERROR_TOTAL=79,CRCC1_RAW_CHSUM_GOOD_TOTAL=80,CRCC1_RAW_CHSUM_ERROR_TOTAL=81,CRCC1_CRC64E_CHSUM_GOOD_TOTAL=82,CRCC1_CRC64E_CHSUM_ERROR_TOTAL=83,CRCC1_ENC_CHSUM_GOOD_TOTAL=84,CRCC1_ENC_CHSUM_ERROR_TOTAL=85,CRCC1_NVME_CHSUM_GOOD_TOTAL=86,CRCC1_NVME_CHSUM_ERROR_TOTAL=87,CRCC0_RAW_CHSUM_GOOD_TOTAL=88,
CRCC0_RAW_CHSUM_ERROR_TOTAL=89,CRCC0_CRC64E_CHSUM_GOOD_TOTAL=90,CRCC0_CRC64E_CHSUM_ERROR_TOTAL=91,CRCC0_ENC_CHSUM_GOOD_TOTAL=92,CRCC0_ENC_CHSUM_ERROR_TOTAL=93,CRCC0_NVME_CHSUM_GOOD_TOTAL=94,CRCC0_NVME_CHSUM_ERROR_TOTAL=95,CG_ENGINE_ERROR_COMMAND=96,CG_SELECT_ENGINE_ERROR_COMMAND=97,CG_SYSTEM_ERROR_COMMAND=98,
CG_CQE_OUTPUT_COMMAND=99,HUFD_FE_XP9_FRM_TOTAL=320,HUFD_FE_XP9_BLK_TOTAL=321,HUFD_FE_XP9_RAW_FRM_TOTAL=322,HUFD_FE_XP10_FRM_TOTAL=323,HUFD_FE_XP10_FRM_PFX_TOTAL=324,HUFD_FE_XP10_FRM_PDH_TOTAL=325,HUFD_FE_XP10_BLK_TOTAL=326,HUFD_FE_XP10_RAW_BLK_TOTAL=327,HUFD_FE_GZIP_FRM_TOTAL=328,
HUFD_FE_GZIP_BLK_TOTAL=329,HUFD_FE_GZIP_RAW_BLK_TOTAL=330,HUFD_FE_ZLIB_FRM_TOTAL=331,HUFD_FE_ZLIB_BLK_TOTAL=332,HUFD_FE_ZLIB_RAW_BLK_TOTAL=333,HUFD_FE_CHU4K_TOTAL=334,HUFD_FE_CHU8K_TOTAL=335,HUFD_FE_CHU4K_RAW_TOTAL=336,HUFD_FE_CHU8K_RAW_TOTAL=337,HUFD_FE_PFX_CRC_ERR_TOTAL=338,
HUFD_FE_PHD_CRC_ERR_TOTAL=339,HUFD_FE_XP9_CRC_ERR_TOTAL=340,HUFD_HTF_XP9_SIMPLE_SHORT_BLK_TOTAL=341,HUFD_HTF_XP9_RETRO_SHORT_BLK_TOTAL=342,HUFD_HTF_XP9_SIMPLE_LONG_BLK_TOTAL=343,HUFD_HTF_XP9_RETRO_LONG_BLK_TOTAL=344,HUFD_HTF_XP10_SIMPLE_SHORT_BLK_TOTAL=345,HUFD_HTF_XP10_RETRO_SHORT_BLK_TOTAL=346,HUFD_HTF_XP10_PREDEF_SHORT_BLK_TOTAL=347,HUFD_HTF_XP10_SIMPLE_LONG_BLK_TOTAL=348,
HUFD_HTF_XP10_RETRO_LONG_BLK_TOTAL=349,HUFD_HTF_XP10_PREDEF_LONG_BLK_TOTAL=350,HUFD_HTF_CHU4K_SIMPLE_SHORT_BLK_TOTAL=351,HUFD_HTF_CHU4K_RETRO_SHORT_BLK_TOTAL=352,HUFD_HTF_CHU4K_PREDEF_SHORT_BLK_TOTAL=353,HUFD_HTF_CHU4K_SIMPLE_LONG_BLK_TOTAL=354,HUFD_HTF_CHU4K_RETRO_LONG_BLK_TOTAL=355,HUFD_HTF_CHU4K_PREDEF_LONG_BLK_TOTAL=356,HUFD_HTF_CHU8K_SIMPLE_SHORT_BLK_TOTAL=357,HUFD_HTF_CHU8K_RETRO_SHORT_BLK_TOTAL=358,
HUFD_HTF_CHU8K_PREDEF_SHORT_BLK_TOTAL=359,HUFD_HTF_CHU8K_SIMPLE_LONG_BLK_TOTAL=360,HUFD_HTF_CHU8K_RETRO_LONG_BLK_TOTAL=361,HUFD_HTF_CHU8K_PREDEF_LONG_BLK_TOTAL=362,HUFD_HTF_DEFLATE_DYNAMIC_BLK_TOTAL=363,HUFD_HTF_DEFLATE_FIXED_BLK_TOTAL=364,HUFD_MTF_0_TOTAL=365,HUFD_MTF_1_TOTAL=366,HUFD_MTF_2_TOTAL=367,HUFD_MTF_3_TOTAL=368,
HUFD_FE_FHP_STALL_TOTAL=369,HUFD_FE_LFA_STALL_TOTAL=370,HUFD_HTF_PREDEF_STALL_TOTAL=371,HUFD_HTF_HDR_DATA_STALL_TOTAL=372,HUFD_HTF_HDR_INFO_STALL_TOTAL=373,HUFD_SDD_INPUT_STALL_TOTAL=374,HUFD_SDD_BUF_FULL_STALL_TOTAL=375,LZ77D_PTR_LEN_256_TOTAL=384,LZ77D_PTR_LEN_128_TOTAL=385,LZ77D_PTR_LEN_64_TOTAL=386,
LZ77D_PTR_LEN_32_TOTAL=387,LZ77D_PTR_LEN_11_TOTAL=388,LZ77D_PTR_LEN_10_TOTAL=389,LZ77D_PTR_LEN_9_TOTAL=390,LZ77D_PTR_LEN_8_TOTAL=391,LZ77D_PTR_LEN_7_TOTAL=392,LZ77D_PTR_LEN_6_TOTAL=393,LZ77D_PTR_LEN_5_TOTAL=394,LZ77D_PTR_LEN_4_TOTAL=395,LZ77D_PTR_LEN_3_TOTAL=396,
LZ77D_LANE_1_LITERALS_TOTAL=397,LZ77D_LANE_2_LITERALS_TOTAL=398,LZ77D_LANE_3_LITERALS_TOTAL=399,LZ77D_LANE_4_LITERALS_TOTAL=400,LZ77D_PTRS_TOTAL=401,LZ77D_FRM_IN_TOTAL=402,LZ77D_FRM_OUT_TOTAL=403,LZ77D_STALL_TOTAL=404,DECRYPT_IV_MISMATCH_FRAME=448,DECRYPT_ENGINE_ID_MISMATCH_FRAME=449,
DECRYPT_SEQ_ID_MISMATCH_FRAME=450,DECRYPT_HMAC_SHA256_TAG_FAIL_FRAME=451,DECRYPT_SHA256_TAG_FAIL_FRAME=452,DECRYPT_GMAC_TAG_FAIL_FRAME=453,DECRYPT_GCM_TAG_FAIL_FRAME=454,DECRYPT_AUTH_NOP_FRAME=455,DECRYPT_AUTH_HMAC_SHA256_FRAME=456,DECRYPT_AUTH_SHA256_FRAME=457,DECRYPT_AUTH_AES_GMAC_FRAME=458,DECRYPT_CIPH_NOP_FRAME=459,
DECRYPT_CIPH_AES_XEX_FRAME=460,DECRYPT_CIPH_AES_XTS_FRAME=461,DECRYPT_CIPH_AES_GCM_FRAME=462,OSF_DATA_INPUT_STALL_TOTAL=512,OSF_CG_INPUT_STALL_TOTAL=513,OSF_OUTPUT_BACKPRESSURE_TOTAL=514,OSF_OUTPUT_STALL_TOTAL=515,ENCRYPT_IV_MISMATCH_FRAME=576,ENCRYPT_ENGINE_ID_MISMATCH_FRAME=577,ENCRYPT_SEQ_ID_MISMATCH_FRAME=578,
ENCRYPT_HMAC_SHA256_TAG_FAIL_FRAME=579,ENCRYPT_SHA256_TAG_FAIL_FRAME=580,ENCRYPT_GMAC_TAG_FAIL_FRAME=581,ENCRYPT_GCM_TAG_FAIL_FRAME=582,ENCRYPT_AUTH_NOP_FRAME=583,ENCRYPT_AUTH_HMAC_SHA256_FRAME=584,ENCRYPT_AUTH_SHA256_FRAME=585,ENCRYPT_AUTH_AES_GMAC_FRAME=586,ENCRYPT_CIPH_NOP_FRAME=587,ENCRYPT_CIPH_AES_XEX_FRAME=588,
ENCRYPT_CIPH_AES_XTS_FRAME=589,ENCRYPT_CIPH_AES_GCM_FRAME=590,SHORT_MAP_ERR_TOTAL=640,LONG_MAP_ERR_TOTAL=641,XP9_BLK_COMP_TOTAL=642,XP9_FRM_RAW_TOTAL=643,XP9_FRM_TOTAL=644,XP9_BLK_SHORT_SIM_TOTAL=645,XP9_BLK_LONG_SIM_TOTAL=646,XP9_BLK_SHORT_RET_TOTAL=647,
XP9_BLK_LONG_RET_TOTAL=648,XP10_BLK_COMP_TOTAL=649,XP10_BLK_RAW_TOTAL=650,XP10_BLK_SHORT_SIM_TOTAL=651,XP10_BLK_LONG_SIM_TOTAL=652,XP10_BLK_SHORT_RET_TOTAL=653,XP10_BLK_LONG_RET_TOTAL=654,XP10_BLK_SHORT_PRE_TOTAL=655,XP10_BLK_LONG_PRE_TOTAL=656,XP10_FRM_TOTAL=657,
CHU8_FRM_RAW_TOTAL=658,CHU8_FRM_COMP_TOTAL=659,CHU8_FRM_SHORT_SIM_TOTAL=660,CHU8_FRM_LONG_SIM_TOTAL=661,CHU8_FRM_SHORT_RET_TOTAL=662,CHU8_FRM_LONG_RET_TOTAL=663,CHU8_FRM_SHORT_PRE_TOTAL=664,CHU8_FRM_LONG_PRE_TOTAL=665,CHU8_CMD_TOTAL=666,CHU4_FRM_RAW_TOTAL=667,
CHU4_FRM_COMP_TOTAL=668,CHU4_FRM_SHORT_SIM_TOTAL=669,CHU4_FRM_LONG_SIM_TOTAL=670,CHU4_FRM_SHORT_RET_TOTAL=671,CHU4_FRM_LONG_RET_TOTAL=672,CHU4_FRM_SHORT_PRE_TOTAL=673,CHU4_FRM_LONG_PRE_TOTAL=674,CHU4_CMD_TOTAL=675,DF_BLK_COMP_TOTAL=676,DF_BLK_RAW_TOTAL=677,
DF_BLK_SHORT_SIM_TOTAL=678,DF_BLK_LONG_SIM_TOTAL=679,DF_BLK_SHORT_RET_TOTAL=680,DF_BLK_LONG_RET_TOTAL=681,DF_FRM_TOTAL=682,PASS_THRU_FRM_TOTAL=683,BYTE_0_TOTAL=684,BYTE_1_TOTAL=685,BYTE_2_TOTAL=686,BYTE_3_TOTAL=687,
BYTE_4_TOTAL=688,BYTE_5_TOTAL=689,BYTE_6_TOTAL=690,BYTE_7_TOTAL=691,ENCRYPT_STALL_TOTAL=692,LZ77_STALL_TOTAL=693,LZ77C_eof_FRAME=704,LZ77C_bypass_FRAME=705,LZ77C_mtf_3_TOTAL=706,LZ77C_mtf_2_TOTAL=707,
LZ77C_mtf_1_TOTAL=708,LZ77C_mtf_0_TOTAL=709,LZ77C_run_256_nup_TOTAL=710,LZ77C_run_128_255_TOTAL=711,LZ77C_run_64_127_TOTAL=712,LZ77C_run_32_63_TOTAL=713,LZ77C_run_11_31_TOTAL=714,LZ77C_run_10_TOTAL=715,LZ77C_run_9_TOTAL=716,LZ77C_run_8_TOTAL=717,
LZ77C_run_7_TOTAL=718,LZ77C_run_6_TOTAL=719,LZ77C_run_5_TOTAL=720,LZ77C_run_4_TOTAL=721,LZ77C_run_3_TOTAL=722,LZ77C_mtf_TOTAL=723,LZ77C_ptr_TOTAL=724,LZ77C_four_lit_TOTAL=725,LZ77C_three_lit_TOTAL=726,LZ77C_two_lit_TOTAL=727,
LZ77C_one_lit_TOTAL=728,LZ77C_throttled_FRAME=729,PREFIX_NUM_0_TOTAL=832,PREFIX_NUM_1_TOTAL=833,PREFIX_NUM_2_TOTAL=834,PREFIX_NUM_3_TOTAL=835,PREFIX_NUM_4_TOTAL=836,PREFIX_NUM_5_TOTAL=837,PREFIX_NUM_6_TOTAL=838,PREFIX_NUM_7_TOTAL=839,
PREFIX_NUM_8_TOTAL=840,PREFIX_NUM_9_TOTAL=841,PREFIX_NUM_10_TOTAL=842,PREFIX_NUM_11_TOTAL=843,PREFIX_NUM_12_TOTAL=844,PREFIX_NUM_13_TOTAL=845,PREFIX_NUM_14_TOTAL=846,PREFIX_NUM_15_TOTAL=847,PREFIX_NUM_16_TOTAL=848,PREFIX_NUM_17_TOTAL=849,
PREFIX_NUM_18_TOTAL=850,PREFIX_NUM_19_TOTAL=851,PREFIX_NUM_20_TOTAL=852,PREFIX_NUM_21_TOTAL=853,PREFIX_NUM_22_TOTAL=854,PREFIX_NUM_23_TOTAL=855,PREFIX_NUM_24_TOTAL=856,PREFIX_NUM_25_TOTAL=857,PREFIX_NUM_26_TOTAL=858,PREFIX_NUM_27_TOTAL=859,
PREFIX_NUM_28_TOTAL=860,PREFIX_NUM_29_TOTAL=861,PREFIX_NUM_30_TOTAL=862,PREFIX_NUM_31_TOTAL=863,PREFIX_NUM_32_TOTAL=864,PREFIX_NUM_33_TOTAL=865,PREFIX_NUM_34_TOTAL=866,PREFIX_NUM_35_TOTAL=867,PREFIX_NUM_36_TOTAL=868,PREFIX_NUM_37_TOTAL=869,
PREFIX_NUM_38_TOTAL=870,PREFIX_NUM_39_TOTAL=871,PREFIX_NUM_40_TOTAL=872,PREFIX_NUM_41_TOTAL=873,PREFIX_NUM_42_TOTAL=874,PREFIX_NUM_43_TOTAL=875,PREFIX_NUM_44_TOTAL=876,PREFIX_NUM_45_TOTAL=877,PREFIX_NUM_46_TOTAL=878,PREFIX_NUM_47_TOTAL=879,
PREFIX_NUM_48_TOTAL=880,PREFIX_NUM_49_TOTAL=881,PREFIX_NUM_50_TOTAL=882,PREFIX_NUM_51_TOTAL=883,PREFIX_NUM_52_TOTAL=884,PREFIX_NUM_53_TOTAL=885,PREFIX_NUM_54_TOTAL=886,PREFIX_NUM_55_TOTAL=887,PREFIX_NUM_56_TOTAL=888,PREFIX_NUM_57_TOTAL=889,
PREFIX_NUM_58_TOTAL=890,PREFIX_NUM_59_TOTAL=891,PREFIX_NUM_60_TOTAL=892,PREFIX_NUM_61_TOTAL=893,PREFIX_NUM_62_TOTAL=894,PREFIX_NUM_63_TOTAL=895,ISF_INPUT_COMMANDS=896,ISF_INPUT_FRAMES=897,ISF_INPUT_STALL_TOTAL=898,ISF_INPUT_SYSTEM_STALL_TOTAL=899,
ISF_OUTPUT_BACKPRESSURE_TOTAL=900,ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_0=901,ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_1=902,ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_2=903,ISF_AUX_CMD_COMPRESS_CTL_MATCH_COMMAND_3=904,HUF_COMP_LZ77D_PTR_LEN_256_TOTAL=960,HUF_COMP_LZ77D_PTR_LEN_128_TOTAL=961,HUF_COMP_LZ77D_PTR_LEN_64_TOTAL=962,HUF_COMP_LZ77D_PTR_LEN_32_TOTAL=963,HUF_COMP_LZ77D_PTR_LEN_11_TOTAL=964,
HUF_COMP_LZ77D_PTR_LEN_10_TOTAL=965,HUF_COMP_LZ77D_PTR_LEN_9_TOTAL=966,HUF_COMP_LZ77D_PTR_LEN_8_TOTAL=967,HUF_COMP_LZ77D_PTR_LEN_7_TOTAL=968,HUF_COMP_LZ77D_PTR_LEN_6_TOTAL=969,HUF_COMP_LZ77D_PTR_LEN_5_TOTAL=970,HUF_COMP_LZ77D_PTR_LEN_4_TOTAL=971,HUF_COMP_LZ77D_PTR_LEN_3_TOTAL=972,HUF_COMP_LZ77D_LANE_4_LITERALS_TOTAL=973,HUF_COMP_LZ77D_LANE_3_LITERALS_TOTAL=974,
HUF_COMP_LZ77D_LANE_2_LITERALS_TOTAL=975,HUF_COMP_LZ77D_LANE_1_LITERALS_TOTAL=976,HUF_COMP_LZ77D_PTRS_TOTAL=977,HUF_COMP_LZ77D_FRM_IN_TOTAL=978,HUF_COMP_LZ77D_FRM_OUT_TOTAL=979,HUF_COMP_LZ77D_STALL_STB_TOTAL=980,CCEIP_STATS_RESERVED=1023} cceip_stats_e;
typedef enum logic [7:0] {NO_ERRORS=0,CRCCG_CRC_ERROR=50,CRCC0_CRC_ERROR=51,CRCC1_CRC_ERROR=52,CRCG0_CRC_ERROR=53,CRCGC0_CRC_ERROR=54,CRCDG0_CRC_ERROR=55,CRCDC0_CRC_ERROR=56,PREFIX_PC_OVERRUN_ERROR=150,PREFIX_NUM_WR_ERROR=151,
PREFIX_ILLEGAL_OPCODE=152,PREFIX_REC_US_SW_EN_ERROR=153,PREFIX_ATTACH_PHD_CRC_ERROR=155,PREFIX_ATTACH_PFD_CRC_ERROR=156,LZ77_COMP_PREFIX_CRC_ERROR=64,LZ77_COMP_INVALID_COMP_ALG=65,LZ77_COMP_INVALID_WIN_SIZE=66,LZ77_COMP_INVALID_MIN_LEN=67,LZ77_COMP_INVALID_NUM_MTF=68,LZ77_COMP_INVALID_MAX_LEN=69,
LZ77_COMP_INVALID_DMW_SIZE=70,LZ77_COMP_LZ_ERROR=71,HE_MEM_ECC=80,HE_PDH_CRC=81,HE_PFX_CRC=82,HE_SYM_MAP_ERR=83,CRYPTO_ENC_DRNG_HEALTH_FAIL=108,CRYPTO_ENC_AAD_LEN_ERROR=107,CRYPTO_ENC_XTS_LEN_ERROR=106,CRYPTO_ENC_MAL_CMD=105,
CRYPTO_ENC_KEY_TLV_CRC_ERROR=104,CRYPTO_ENC_INVALID_ENGINE_ID=103,CRYPTO_ENC_INVALID_SEQNUM=102,CRYPTO_ENC_IV_MISSING=101,CRYPTO_ENC_SEED_EXPIRED=100,CRYPTO_DEC_AAD_LEN_ERROR=118,CRYPTO_DEC_XTS_LEN_ERROR=117,CRYPTO_DEC_MAL_CMD=116,CRYPTO_DEC_KEY_TLV_CRC_ERROR=115,CRYPTO_DEC_INVALID_ENGINE_ID=114,
CRYPTO_DEC_INVALID_SEQNUM=113,CRYPTO_DEC_IV_MISSING=112,CRYPTO_DEC_TAG_MISCOMPARE=110,CRYPTO_INT_KEY_TLV_CRC_ERROR=123,CRYPTO_INT_INVALID_ENGINE_ID=122,CRYPTO_INT_INVALID_SEQNUM=121,CRYPTO_INT_TAG_MISCOMPARE=120,KME_DAK_INV_KIM=130,KME_DAK_PF_VF_VAL_ERR=131,KME_DEK_INV_KIM=132,
KME_DEK_PF_VF_VAL_ERR=133,KME_SEED_EXPIRED=134,KME_DEK_GCM_TAG_FAIL=135,KME_DAK_GCM_TAG_FAIL=136,KME_ECC_FAIL=137,KME_UNSUPPORTED_KEY_TYPE=138,KME_DEK_ILLEGAL_KEK_USAGE=139,KME_DAK_ILLEGAL_KEK_USAGE=140,KME_DRNG_HEALTH_FAIL=141,HD_MEM_ECC=1,
HD_FHP_PFX_CRC=2,HD_FHP_PFX_DATA_ABSENT=3,HD_FHP_PHD_CRC=4,HD_FHP_BAD_FORMAT=5,HD_BHP_INVALID_WSIZE=6,HD_BHP_BLK_CRC=7,HD_BHP_HDR_INVALID=8,HD_BHP_XP9_HDR_SEQ=9,HD_BHP_XP10_XTRA_FLAG_PRSNT=10,HD_BHP_ZLIB_FDICT_PRSNT=11,
HD_BHP_GZ_CM_NOT_DEFLATE=12,HD_BHP_ZLIB_CINFO_RANGE=13,HD_BHP_ZLIB_FCHECK=14,HD_BHP_DFLATE_LEN_CHECK=15,HD_LFA_REWIND_FAIL=16,HD_LFA_PREMATURE_EOF=17,HD_LFA_LATE_EOF=18,HD_LFA_MISSING_EOF=19,HD_HTF_XP9_RESERVED_SYMBOL_TABLE_ENCODING=20,HD_HTF_XP10_RESERVED_SYMBOL_TABLE_ENCODING=21,
HD_HTF_XP10_PREDEF_SYMBOL_TABLE_ENCODING=22,HD_HTF_XP9_ILLEGAL_NONZERO_BL=23,HD_HTF_RLE_OVERRUN=24,HD_HTF_BAD_HUFFMAN_CODE=25,HD_HTF_ILLEGAL_SMALL_HUFFTREE=26,HD_HTF_ILLEGAL_HUFFTREE=27,HD_HTF_HDR_UNDERRUN=28,HD_BHP_STBL_SIZE_ERR=29,HD_SDD_INVALID_SYMBOL=32,HD_SDD_END_MISMATCH=33,
HD_SDD_MISSING_EOB_SYM=34,HD_MTF_XP9_MTF3_AFTER_BACKREF=35,HD_MTF_XP10_MISSING_MTF=36,HD_BHP_ILLEGAL_MTF_SZ=37,HD_LZ_HBIF_SOFT_OFLOW=38,HD_BE_FRM_CRC=39,HD_BE_OLIMIT=40,HD_BE_SZ_MISMATCH=41,CG_UNDEF_FRMD_OUT=170,ISF_PREFIX_ERR=180,TLVP_BIP2_ERROR=255} zipline_error_e;
typedef struct packed {
 logic tvalid;
 logic tlast;
 logic [0:0] tid ;
 logic [7:0] tstrb ;
 logic [7:0] tuser ;
 logic [63:0] tdata ;
} axi4s_dp_bus_t;
typedef struct packed {
 logic tready;
} axi4s_dp_rdy_t;
typedef struct packed {
 logic [19:0] addr ;
 logic wr_strb;
 logic [31:0] wr_data ;
 logic rd_strb;
} rbus_in_t;
typedef struct packed {
 logic [31:0] rd_data ;
 logic ack;
 logic err_ack;
} rbus_out_t;
typedef struct packed {
 logic [19:0] addr ;
 logic wr_strb;
 logic [31:0] wr_data ;
 logic rd_strb;
 logic [31:0] rd_data ;
 logic ack;
 logic err_ack;
} rbus_ring_t;
typedef struct packed {
 logic [15:0] addr ;
 logic wr_strb;
 logic [31:0] wr_data ;
 logic rd_strb;
 logic [31:0] rd_data ;
 logic ack;
 logic err_ack;
} kme_rbus_ring_t;
typedef struct packed {
 logic eob;
 logic [7:0] bytes_vld ;
 logic [22:0] im_meta ;
} im_desc_t;
typedef struct packed {
 logic [63:0] data ;
} im_data_t;
typedef struct packed {
 im_data_t data;
 im_desc_t desc;
} im_din_t;
typedef struct packed {
 logic bank_hi;
 logic bank_lo;
} im_available_t;
typedef struct packed {
 logic bank_hi;
 logic bank_lo;
} im_consumed_t;
typedef struct packed {
 logic valid;
 logic [7:0] seq_num ;
} frame_latency_if_bus_t;
typedef struct packed {
 logic valid;
 logic [15:0] rqe_sched_handle ;
 logic last;
 logic [10:0] tlv_frame_num ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [23:0] bytes_in ;
 logic [23:0] bytes_out ;
 logic [23:0] basis ;
} sched_update_if_bus_t;
typedef struct packed {
 logic insert;
 logic [12:0] ordern ;
 tlv_types_e typen;
 logic sot;
 logic eot;
 logic tlast;
 logic [0:0] tid ;
 logic [7:0] tstrb ;
 logic [7:0] tuser ;
 logic [63:0] tdata ;
} tlvp_if_bus_t;
typedef struct packed {
 logic [3:0] framing ;
 logic [7:0] data0 ;
 logic [7:0] data1 ;
 logic [7:0] data2 ;
 logic [7:0] data3 ;
 logic backref;
 logic backref_type;
 logic [1:0] backref_lane ;
 logic [7:0] offset_msb ;
 logic [15:0] length ;
} lz_symbol_bus_t;
typedef struct packed {
 logic [1:0] tlv_bip2 ;
 logic [18:0] resv0 ;
 logic [10:0] tlv_frame_num ;
 logic [3:0] resv1 ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [7:0] tlv_len ;
 tlv_types_e tlv_type;
} tlv_word_0_t;
typedef struct packed {
 logic [1:0] tlv_bip2 ;
 logic no_data;
 logic aux_frmd_crc;
 rqe_frame_size_e frame_size;
 logic vf_valid;
 rqe_trace_e trace;
 logic [10:0] unused ;
 logic [10:0] tlv_frame_num ;
 logic [3:0] resv0 ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [7:0] tlv_len ;
 tlv_types_e tlv_type;
} tlv_rqe_word_0_t;
typedef struct packed {
 logic [1:0] tlv_bip2 ;
 logic last_of_command;
 logic [15:0] resv0 ;
 frmd_coding_e coding;
 logic [10:0] tlv_frame_num ;
 logic [3:0] resv1 ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [7:0] tlv_len ;
 tlv_types_e tlv_type;
} tlv_data_word_0_t;
typedef struct packed {
 logic [3:0] pf_number ;
 logic [11:0] vf_number ;
 logic [15:0] scheduler_handle ;
 logic [31:0] src_data_len ;
} tlv_rqe_word_1_t;
typedef struct packed {
 tlvp_corrupt_e tlvp_corrupt;
 cmd_mode_e cmd_mode;
 logic [4:0] module_id ;
 cmd_type_e cmd_type;
 logic [4:0] tlv_num ;
 logic [9:0] byte_num ;
 logic [7:0] byte_msk ;
} cmd_debug_t;
typedef struct packed {
 logic [0:0] rsvd ;
 logic [10:0] on_count ;
 logic [10:0] off_count ;
} bp_debug_t;
typedef struct packed {
 cmd_debug_t debug;
 logic trace;
 logic dst_guid_present;
 logic [6:0] frmd_out_type ;
 cmd_md_op_e md_op;
 cmd_md_type_e md_type;
 logic [6:0] frmd_in_type ;
 logic [5:0] frmd_in_aux ;
 cmd_frmd_crc_in_e frmd_crc_in;
 cmd_guid_present_e src_guid_present;
 cmd_compound_cmd_frm_size_e compound_cmd_frm_size;
} tlv_cmd_word_1_t;
typedef struct packed {
 logic rsvd2;
 aux_key_type_e key_type;
 logic [1:0] rsvd1 ;
 cmd_cipher_pad_e cipher_pad;
 cmd_iv_op_e iv_op;
 logic [7:0] aad_len ;
 cmd_cipher_op_e cipher_op;
 cmd_auth_op_e auth_op, raw_auth_op;
 logic [7:0] rsvd0 ;
 cmd_chu_comp_thrsh_e chu_comp_thrsh;
 cmd_xp10_crc_mode_e xp10_crc_mode;
 logic [5:0] xp10_user_prefix_size ;
 cmd_xp10_prefix_mode_e xp10_prefix_mode;
 cmd_lz77_max_symb_len_e lz77_max_symb_len;
 cmd_lz77_min_match_len_e lz77_min_match_len;
 cmd_lz77_dly_match_win_e lz77_dly_match_win;
 cmd_lz77_win_size_e lz77_win_size;
 cmd_comp_mode_e comp_mode;
} tlv_cmd_word_2_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_key_word1_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_key_word2_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_key_word3_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_key_word4_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} tlv_key_word5_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} tlv_key_word6_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word7_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word8_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word9_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word10_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word11_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word12_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word13_t;
typedef struct packed {
 logic [63:0] dek ;
} tlv_key_word14_t;
typedef struct packed {
 logic [63:0] dak ;
} tlv_key_word15_t;
typedef struct packed {
 logic [63:0] dak ;
} tlv_key_word16_t;
typedef struct packed {
 logic [63:0] dak ;
} tlv_key_word17_t;
typedef struct packed {
 logic [63:0] dak ;
} tlv_key_word18_t;
typedef struct packed {
 logic [55:0] rsvd ;
 zipline_error_e kme_errors;
} tlv_key_word19_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [31:0] crc32 ;
} tlv_key_word20_t;
typedef struct packed {
 logic [63:6] rsvd ;
 logic [5:0] xp10_prefix_sel ;
} tlv_phd_word1_t;
typedef struct packed {
 logic [1:0] tlv_bip2 ;
 logic [11:0] resv0 ;
 logic prefix_src;
 logic [5:0] xp10_prefix_sel ;
 logic [10:0] tlv_frame_num ;
 logic [3:0] resv1 ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [7:0] tlv_len ;
 tlv_types_e tlv_type;
} tlv_pfd_word0_t;
typedef struct packed {
 logic [63:6] rsvd ;
 logic [5:0] xp10_prefix_sel ;
} tlv_pfd_word1_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_guid_word1_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_guid_word2_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_guid_word3_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_guid_word4_t;
typedef struct packed {
 logic [1:0] tlv_bip2 ;
 logic [1:0] rsvd3 ;
 logic [7:0] gen_frmd_out_type ;
 logic [1:0] rsvd2 ;
 frmd_mac_size_e raw_data_mac_size, enc_cmp_data_mac_size;
 frmd_coding_e coding;
 logic rsvd1;
 logic [10:0] tlv_frame_num ;
 logic [3:0] rsvd0 ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [7:0] tlv_len ;
 tlv_types_e tlv_type;
} tlv_ftr_word0_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} tlv_ftr_word1_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} tlv_ftr_word2_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} tlv_ftr_word3_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} tlv_ftr_word4_t;
typedef struct packed {
 logic [63:0] raw_data_cksum ;
} tlv_ftr_word5_t;
typedef struct packed {
 logic [63:0] raw_data_cksum_protocol ;
} tlv_ftr_word6_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} tlv_ftr_word7_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} tlv_ftr_word8_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} tlv_ftr_word9_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} tlv_ftr_word10_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_cksum ;
} tlv_ftr_word11_t;
typedef struct packed {
 logic [15:0] nvme_raw_cksum_crc16t ;
 logic [23:0] bytes_in ;
 logic [23:0] bytes_out ;
} tlv_ftr_word12_t;
typedef struct packed {
 logic [19:0] rsvd1 ;
 logic [23:0] compressed_length ;
 zipline_error_e error_code;
 logic rsvd0;
 logic [10:0] errored_frame_number ;
} tlv_ftr_word13_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_ftr_guid_word0_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_ftr_guid_word1_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_ftr_guid_word2_t;
typedef struct packed {
 logic [63:0] guid ;
} tlv_ftr_guid_word3_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [31:0] iv ;
} tlv_ftr_iv_word0_t;
typedef struct packed {
 logic [63:0] iv ;
} tlv_ftr_iv_word1_t;
typedef struct packed {
 logic [7:0] rsvd1 ;
 logic [23:0] bytes_in ;
 logic [7:0] rsvd0 ;
 logic [23:0] bytes_out ;
} tlv_stats_word1_t;
typedef struct packed {
 logic [30:0] rsvd1 ;
 logic frame_error;
 logic [7:0] rsvd0 ;
 logic [23:0] latency ;
} tlv_stats_word2_t;
typedef struct packed {
 logic [7:0] status_code ;
 logic do_not_resend;
 logic vf_valid;
 logic [1:0] rsvd0 ;
 logic [7:0] error_code ;
 logic [11:0] errored_frame_number ;
 logic [2:0] status_code_type ;
 logic [12:0] stat_cts ;
 logic [3:0] pf_number ;
 logic [11:0] vf_number ;
} tlv_cqe_word1_t;
typedef struct packed {
 logic [47:0] rsvd ;
 logic [15:0] nvme_raw_cksum_crc16t ;
} fmd_user_pi16_word1_t;
typedef struct packed {
 logic [63:0] raw_data_cksum ;
} fmd_user_pi64_word1_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_user_vm_word1_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_user_vm_word2_t;
typedef struct packed {
 logic [63:0] raw_data_cksum ;
} fmd_user_vm_word3_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_user_vm_word4_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_user_vm_word5_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_user_vm_word6_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_user_vm_word7_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [5:0] rsvd0 ;
 frmd_coding_e coding;
 logic [23:0] compressed_length ;
} fmd_int_app_word6_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_cksum ;
} fmd_int_app_word1_t;
typedef struct packed {
 logic [63:0] enc_cmp_mac ;
} fmd_int_app_word2_t;
typedef struct packed {
 logic [63:0] enc_cmp_mac ;
} fmd_int_app_word3_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_int_app_word4_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [31:0] ivtweak ;
} fmd_int_app_word5_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [5:0] rsvd0 ;
 frmd_coding_e coding;
 logic [23:0] compressed_length ;
} fmd_int_sip_word3_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_cksum ;
} fmd_int_sip_word1_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_sip_word2_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [5:0] rsvd0 ;
 frmd_coding_e coding;
 logic [23:0] compressed_length ;
} fmd_int_lip_word6_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_cksum ;
} fmd_int_lip_word1_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_lip_word2_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_lip_word3_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_lip_word4_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_lip_word5_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [5:0] rsvd0 ;
 frmd_coding_e coding;
 logic [23:0] compressed_length ;
} fmd_int_vm_word12_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_cksum ;
} fmd_int_vm_word1_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_word2_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_word3_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_word4_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_word5_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_vm_word6_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_vm_word7_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_vm_word8_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_vm_word9_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_int_vm_word10_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_int_vm_word11_t;
typedef struct packed {
 logic [31:0] rsvd ;
 logic [5:0] rsvd0 ;
 frmd_coding_e coding;
 logic [23:0] compressed_length ;
} fmd_int_vm_short_word9_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_cksum ;
} fmd_int_vm_short_word1_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_short_word2_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_short_word3_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_short_word4_t;
typedef struct packed {
 logic [63:0] enc_cmp_data_mac ;
} fmd_int_vm_short_word5_t;
typedef struct packed {
 logic [63:0] raw_data_mac ;
} fmd_int_vm_short_word6_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_int_vm_short_word7_t;
typedef struct packed {
 logic [63:0] ivtweak ;
} fmd_int_vm_short_word8_t;
typedef struct packed {
 logic predet_mem_mask;
 logic [3:0] predet_mem_id ;
 cmd_comp_mode_e comp_mode;
 cmd_lz77_win_size_e lz77_win_size;
 cmd_lz77_min_match_len_e lz77_min_match_len;
 cmd_xp10_prefix_mode_e xp10_prefix_mode;
 logic [5:0] xp10_user_prefix_size ;
 cmd_xp10_crc_mode_e xp10_crc_mode;
 cmd_chu_comp_thrsh_e chu_comp_thrsh;
 logic [0:0] tid ;
 logic [7:0] tuser ;
 logic [23:0] raw_byte_count ;
 logic [17:0] extra_bit_count ;
 logic [10:0] blk_count ;
 logic blk_last;
 logic pdh_crc_err;
 logic [63:0] raw_crc ;
} s_sm_seq_id_intf;
typedef struct packed {
 cmd_comp_mode_e comp_mode;
 cmd_lz77_win_size_e lz77_win_size;
 cmd_xp10_prefix_mode_e xp10_prefix_mode;
} s_seq_id_type_intf;
typedef struct packed {
 logic [17:0] count_part1 ;
 logic [31:0] count_part0 ;
} counter_50_t;
typedef struct packed {
 logic cqe_out;
 logic cqe_sys_err;
 logic cqe_err_sel;
 logic cqe_eng_err;
} cg_stats_t;
typedef struct packed {
 logic [59:0] rsvd ;
 logic ob_stall;
 logic ob_sys_bp;
 logic pdt_fifo_stall;
 logic dat_fifo_stall;
} osf_stats_t;
typedef struct packed {
 logic [54:0] rsvd ;
 logic aux_cmd_match3;
 logic aux_cmd_match2;
 logic aux_cmd_match1;
 logic aux_cmd_match0;
 logic ob_sys_bp;
 logic ib_sys_stall;
 logic ib_stall;
 logic ib_frame;
 logic ib_cmd;
} isf_stats_t;
typedef struct packed {
 logic [9:0] huff_comp_rsvd ;
 logic lz77_stall_stb;
 logic encrypt_stall_stb;
 logic byte_7_stb;
 logic byte_6_stb;
 logic byte_5_stb;
 logic byte_4_stb;
 logic byte_3_stb;
 logic byte_2_stb;
 logic byte_1_stb;
 logic byte_0_stb;
 logic pass_thru_frm_stb;
 logic df_frm_stb;
 logic df_blk_long_ret_stb;
 logic df_blk_shrt_ret_stb;
 logic df_blk_long_sim_stb;
 logic df_blk_shrt_sim_stb;
 logic df_blk_raw_stb;
 logic df_blk_enc_stb;
 logic chu4_cmd_stb;
 logic chu4_frm_long_pre_stb;
 logic chu4_frm_shrt_pre_stb;
 logic chu4_frm_long_ret_stb;
 logic chu4_frm_shrt_ret_stb;
 logic chu4_frm_long_sim_stb;
 logic chu4_frm_shrt_sim_stb;
 logic chu4_frm_enc_stb;
 logic chu4_frm_raw_stb;
 logic chu8_cmd_stb;
 logic chu8_frm_long_pre_stb;
 logic chu8_frm_shrt_pre_stb;
 logic chu8_frm_long_ret_stb;
 logic chu8_frm_shrt_ret_stb;
 logic chu8_frm_long_sim_stb;
 logic chu8_frm_shrt_sim_stb;
 logic chu8_frm_enc_stb;
 logic chu8_frm_raw_stb;
 logic xp10_frm_stb;
 logic xp10_blk_long_pre_stb;
 logic xp10_blk_shrt_pre_stb;
 logic xp10_blk_long_ret_stb;
 logic xp10_blk_shrt_ret_stb;
 logic xp10_blk_long_sim_stb;
 logic xp10_blk_shrt_sim_stb;
 logic xp10_blk_raw_stb;
 logic xp10_blk_enc_stb;
 logic xp9_blk_long_ret_stb;
 logic xp9_blk_shrt_ret_stb;
 logic xp9_blk_long_sim_stb;
 logic xp9_blk_shrt_sim_stb;
 logic xp9_frm_stb;
 logic xp9_frm_raw_stb;
 logic xp9_blk_enc_stb;
 logic long_map_err_stb;
 logic shrt_map_err_stb;
} huf_comp_stats_t;
typedef struct packed {
 logic [48:0] unused ;
 logic [0:0] cipher_aes_gcm ;
 logic [0:0] cipher_aes_xts ;
 logic [0:0] cipher_aes_xex ;
 logic [0:0] cipher_nop ;
 logic [0:0] auth_aes_gmac ;
 logic [0:0] auth_sha256 ;
 logic [0:0] auth_sha256_hmac ;
 logic [0:0] auth_nop ;
 logic [0:0] gcm_tag_fail ;
 logic [0:0] gmac_tag_fail ;
 logic [0:0] sha256_tag_fail ;
 logic [0:0] hmac_sha256_tag_fail ;
 logic [0:0] seq_id_mismatch ;
 logic [0:0] eng_id_mismatch ;
 logic [0:0] reserved ;
} crypto_stats_t;
typedef struct packed {
 aux_key_op_e dak_key_op;
 logic [13:0] dak_key_ref ;
 aux_kdf_mode_e kdf_mode;
 aux_key_op_e dek_key_op;
 logic [13:0] dek_key_ref ;
} aux_key_ctrl_t;
typedef struct packed {
 logic tvalid;
 logic tlast;
 logic [1:0] tuser ;
 logic [7:0] tdata ;
} axi4s_su_dp_bus_t;
typedef struct packed {
 logic tlvp_err;
 logic uncor_ecc_err;
 logic bimc_int;
} generic_int_t;
typedef struct packed {
 logic uncor_ecc_err;
} ecc_int_t;
typedef struct packed {
 logic tlvp_err;
} tlvp_int_t;
typedef struct packed {
 logic bimc_err;
} bimc_int_t;
typedef struct packed {
 logic seed_expire;
 logic id_mismatch;
 logic tlvp_err;
 logic uncor_ecc_err;
} crypto_int_t;
typedef struct packed {
 logic id_mismatch;
 logic tlvp_err;
} crypto_ckmic_int_t;
typedef struct packed {
 logic tlvp_err;
 logic uncor_ecc_err;
} osf_int_t;
typedef struct packed {
 logic sys_stall;
 logic ovfl;
 logic prot_err;
 logic tlvp_int;
 logic uncor_ecc_err;
} isf_int_t;
typedef struct packed {
 logic tlvp_err;
 logic uncor_ecc_err;
} prefix_attach_int_t;
typedef struct packed {
 zipline_error_e error_code;
 logic [10:0] errored_frame_number ;
} ftr_error_t;
typedef struct packed {
 logic [0:0] valid ;
 logic [2:0] label_index ;
 logic [1:0] ckv_length ;
 logic [14:0] ckv_pointer ;
 logic [3:0] pf_num ;
 logic [11:0] vf_num ;
 logic [0:0] vf_valid ;
} kim_entry_t;
typedef struct packed {
 logic [0:0] guid_size ;
 logic [5:0] label_size ;
 logic [255:0] label ;
 logic [0:0] delimiter_valid ;
 logic [7:0] delimiter ;
} label_t;
typedef struct packed {
 logic [0:0] valid ;
 logic [2:0] label_index ;
 logic [0:0] pf_num ;
 logic [0:0] vf_valid ;
 logic [8:0] vf_num ;
 logic [511:0] ckv_key ;
} kim_ckv_resp_t;
typedef enum logic [3:0] {KME_WORD0=4'b0,KME_DEBUG_KEYHDR=4'b01,KME_IVTWEAK=4'b010,KME_GUID=4'b011,KME_KIM=4'b0100,KME_DEK_CKV0=4'b0101,KME_DEK_CKV1=4'b0110,KME_DAK_CKV=4'b0111,KME_EIV=4'b1000,KME_DEK0=4'b1001,
KME_DEK1=4'b1010,KME_ETAG=4'b1011,KME_AIV=4'b1100,KME_DAK=4'b1101,KME_ATAG=4'b1110,KME_ERROR=4'b1111} kme_internal_id;
typedef enum logic [5:0] {IDX_KME_WORD0=6'b0,IDX_KME_DEBUG_KEYHDR=6'b01,IDX_KME_GUID=6'b010,IDX_KME_IVTWEAK=6'b0110,IDX_KME_KIM=6'b01000,IDX_KME_DEK_CKV0=6'b01010,IDX_KME_DEK_CKV1=6'b01110,IDX_KME_DAK_CKV=6'b010010,IDX_KME_EIV=6'b010110,IDX_KME_DEK0=6'b011000,
IDX_KME_DEK1=6'b011100,IDX_KME_ETAG=6'b100000,IDX_KME_AIV=6'b100010,IDX_KME_DAK=6'b100100,IDX_KME_ATAG=6'b101000,IDX_KME_ERROR=6'b101010} kme_internal_idx;
typedef struct packed {
 logic [0:0] sot ;
 logic [0:0] eoi ;
 logic [0:0] eot ;
 kme_internal_id id;
 logic [63:0] tdata ;
} kme_internal_t;
typedef struct packed {
 logic [1:0] tlv_bip2 ;
 logic [12:0] resv0 ;
 logic [0:0] kdf_dek_iter ;
 logic [0:0] keyless_algos ;
 logic [0:0] needs_dek ;
 logic [0:0] needs_dak ;
 aux_key_type_e key_type;
 logic [10:0] tlv_frame_num ;
 logic [3:0] tlv_eng_id ;
 logic [7:0] tlv_seq_num ;
 logic [7:0] tlv_len ;
 tlv_types_e tlv_type;
} kme_internal_word_0_t;
typedef struct packed {
 kim_entry_t dek_kim_entry;
 logic [5:0] unused ;
 logic [0:0] missing_iv ;
 logic [0:0] missing_guid ;
 logic [0:0] validate_dek ;
 logic [0:0] vf_valid ;
 logic [3:0] pf_num ;
 logic [11:0] vf_num ;
} kme_internal_word_8_t;
typedef struct packed {
 kim_entry_t dak_kim_entry;
 logic [7:0] unused ;
 logic [0:0] validate_dak ;
 logic [0:0] vf_valid ;
 logic [3:0] pf_num ;
 logic [11:0] vf_num ;
} kme_internal_word_9_t;
typedef struct packed {
 logic [0:0] corrupt_crc32 ;
 logic [46:0] unused ;
 zipline_error_e error_code;
} kme_internal_word_42_t;
typedef enum logic [2:0] {PT_CKV=3'b0,PT_KEY_BLOB=3'b01,DECRYPT_DEK256=3'b010,DECRYPT_DEK512=3'b011,DECRYPT_DAK=3'b100,DECRYPT_DEK256_COMB=3'b101,DECRYPT_DEK512_COMB=3'b110,DECRYPT_DAK_COMB=3'b111} gcm_op_e;
typedef struct packed {
 logic [255:0] key0 ;
 logic [255:0] key1 ;
 logic [95:0] iv ;
 gcm_op_e op;
} gcm_cmd_t;
typedef struct packed {
 logic [0:0] tag_mismatch ;
} gcm_status_t;
typedef struct packed {
 logic [0:0] combo_mode ;
} keyfilter_cmd_t;
typedef struct packed {
 logic [0:0] kdf_dek_iter ;
 logic [0:0] combo_mode ;
 aux_key_op_e dek_key_op, dak_key_op;
} kdf_cmd_t;
typedef struct packed {
 logic [0:0] combo_mode ;
 logic [0:0] skip ;
 logic [255:0] guid ;
 logic [2:0] label_index ;
 logic [1:0] num_iter ;
} kdfstream_cmd_t;
// synopsys translate_off
import cr_kmePKG::* ;
// synopsys translate_on
import cr_kme_regfilePKG::* ;
localparam CKV_NUM_ENTRIES = 32768;
localparam CKV_DATA_WIDTH = 64;
localparam KIM_NUM_ENTRIES = 16384;
localparam KIM_DATA_WIDTH = 38;
input  clk;
input  rst_n;
input  disable_debug_cmd_q;
input  always_validate_kim_ref;
output reg stitcher_rd;
input axi4s_dp_bus_t stitcher_out;
input  stitcher_empty;
output  parser_kimreader_valid;
output kme_internal_t parser_kimreader_data;
input  kimreader_parser_ack;
output  tlv_parser_idle;
output  tlv_parser_int_tlv_start_pulse;
typedef struct packed {
 logic [0:0] start ;
 logic [0:0] partial ;
 logic [0:0] endian_swap ;
 kme_internal_id till;
} skip_control;
kme_internal_t fifo_in;
wire  fifo_in_stall;
reg fifo_in_valid;
reg key_blob_region;
reg [5:0] int_tlv_counter ;
reg [4:0] tlv_counter ;
tlv_rqe_word_0_t tlv_word0;
tlv_rqe_word_1_t tlv_word1;
tlv_cmd_word_2_t tlv_word2;
kme_internal_id nxt_fifo_in_id;
tlv_cmd_word_1_t frame_word;
kme_internal_word_0_t kme_internal_word0, nxt_kme_internal_word0;
kme_internal_word_8_t kme_internal_dek_kim_word, nxt_kme_internal_dek_kim_word;
kme_internal_word_9_t kme_internal_dak_kim_word, nxt_kme_internal_dak_kim_word;
tlv_types_e tlv_type, nxt_tlv_type;
aux_key_type_e aux_key_type, nxt_aux_key_type;
cmd_iv_op_e aux_iv_op, nxt_aux_iv_op;
cmd_cipher_op_e aux_cipher_op, nxt_aux_cipher_op;
cmd_auth_op_e aux_auth_op, nxt_aux_auth_op, aux_raw_auth_op, nxt_aux_raw_auth_op;
cmd_debug_t debug_cmd, nxt_debug_cmd;
aux_key_ctrl_t aux_key_header, nxt_aux_key_header;
skip_control skip, nxt_skip;
reg [63:0] guid0 ;
reg [63:0] nxt_guid0 ;
reg [63:0] guid1 ;
reg [63:0] nxt_guid1 ;
reg [63:0] guid2 ;
reg [63:0] nxt_guid2 ;
reg [63:0] guid3 ;
reg [63:0] nxt_guid3 ;
reg [63:0] iv0 ;
reg [63:0] nxt_iv0 ;
reg [63:0] iv1 ;
reg [63:0] nxt_iv1 ;
reg [31:0] buffer ;
reg [31:0] nxt_buffer ;
wire  stitcher_sot;
wire  stitcher_eot;
genvar ii;
genvar jj;
genvar kk;
genvar nn;
genvar qq;
wire  _zy_simnet_stitcher_rd_0_w$;
wire  [0:70] _zy_simnet_parser_kimreader_data_1_w$ ;
wire  [0:70] _zy_simnet_parser_kimreader_data_2_w$ ;
wire  _zy_simnet_dio_3;
wire  _zy_simnet_dio_4;
wire  [0:70] _zy_simnet_fifo_in_5_w$ ;
wire  _zy_simnet_fifo_in_valid_6_w$;
wire  _zy_simnet_cio_7;
wire  _zy_sva_key_type0_line4_1_reset_or;
bit [0:0]  _zy_sva_key_type0_line4_1_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type0_line4_1_ccheck
bit [0:0]  _zy_sva_key_type0_line4_1_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type0_line4_1_cpass
bit _zy_sva_b0;
wire  _zy_sva_key_type0_line5a_2_reset_or;
bit [0:0]  _zy_sva_key_type0_line5a_2_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type0_line5a_2_ccheck
bit [0:0]  _zy_sva_key_type0_line5a_2_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type0_line5a_2_cpass
bit _zy_sva_b1;
wire  _zy_sva_key_type0_line5b_3_reset_or;
bit [0:0]  _zy_sva_key_type0_line5b_3_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type0_line5b_3_ccheck
bit [0:0]  _zy_sva_key_type0_line5b_3_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type0_line5b_3_cpass
bit _zy_sva_b2;
wire  _zy_sva_key_type1_line7a_4_reset_or;
bit [0:0]  _zy_sva_key_type1_line7a_4_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line7a_4_ccheck
bit [0:0]  _zy_sva_key_type1_line7a_4_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line7a_4_cpass
bit _zy_sva_b3;
wire  _zy_sva_key_type1_line7b_5_reset_or;
bit [0:0]  _zy_sva_key_type1_line7b_5_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line7b_5_ccheck
bit [0:0]  _zy_sva_key_type1_line7b_5_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line7b_5_cpass
bit _zy_sva_b4;
wire  _zy_sva_key_type1_line8a_6_reset_or;
bit [0:0]  _zy_sva_key_type1_line8a_6_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line8a_6_ccheck
bit [0:0]  _zy_sva_key_type1_line8a_6_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line8a_6_cpass
bit _zy_sva_b5;
wire  _zy_sva_key_type1_line8b_7_reset_or;
bit [0:0]  _zy_sva_key_type1_line8b_7_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line8b_7_ccheck
bit [0:0]  _zy_sva_key_type1_line8b_7_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line8b_7_cpass
bit _zy_sva_b6;
wire  _zy_sva_key_type1_line9_8_reset_or;
bit [0:0]  _zy_sva_key_type1_line9_8_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line9_8_ccheck
bit [0:0]  _zy_sva_key_type1_line9_8_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line9_8_cpass
bit _zy_sva_b7;
wire  _zy_sva_key_type1_line10_9_reset_or;
bit [0:0]  _zy_sva_key_type1_line10_9_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line10_9_ccheck
bit [0:0]  _zy_sva_key_type1_line10_9_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line10_9_cpass
bit _zy_sva_b8;
wire  _zy_sva_key_type1_line11a_10_reset_or;
bit [0:0]  _zy_sva_key_type1_line11a_10_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11a_10_ccheck
bit [0:0]  _zy_sva_key_type1_line11a_10_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11a_10_cpass
bit _zy_sva_b9;
wire  _zy_sva_key_type1_line11b_11_reset_or;
bit [0:0]  _zy_sva_key_type1_line11b_11_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11b_11_ccheck
bit [0:0]  _zy_sva_key_type1_line11b_11_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11b_11_cpass
bit _zy_sva_b10;
wire  _zy_sva_key_type1_line11c_12_reset_or;
bit [0:0]  _zy_sva_key_type1_line11c_12_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11c_12_ccheck
bit [0:0]  _zy_sva_key_type1_line11c_12_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11c_12_cpass
bit _zy_sva_b11;
wire  _zy_sva_key_type1_line11d_13_reset_or;
bit [0:0]  _zy_sva_key_type1_line11d_13_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11d_13_ccheck
bit [0:0]  _zy_sva_key_type1_line11d_13_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line11d_13_cpass
bit _zy_sva_b12;
wire  _zy_sva_key_type1_line12a_14_reset_or;
bit [0:0]  _zy_sva_key_type1_line12a_14_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line12a_14_ccheck
bit [0:0]  _zy_sva_key_type1_line12a_14_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line12a_14_cpass
bit _zy_sva_b13;
wire  _zy_sva_key_type1_line12b_15_reset_or;
bit [0:0]  _zy_sva_key_type1_line12b_15_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line12b_15_ccheck
bit [0:0]  _zy_sva_key_type1_line12b_15_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type1_line12b_15_cpass
bit _zy_sva_b14;
wire  _zy_sva_key_type9_line14_16_reset_or;
bit [0:0]  _zy_sva_key_type9_line14_16_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line14_16_ccheck
bit [0:0]  _zy_sva_key_type9_line14_16_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line14_16_cpass
bit _zy_sva_b15;
wire  _zy_sva_key_type9_line15_17_reset_or;
bit [0:0]  _zy_sva_key_type9_line15_17_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line15_17_ccheck
bit [0:0]  _zy_sva_key_type9_line15_17_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line15_17_cpass
bit _zy_sva_b16;
wire  _zy_sva_key_type9_line16a_18_reset_or;
bit [0:0]  _zy_sva_key_type9_line16a_18_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line16a_18_ccheck
bit [0:0]  _zy_sva_key_type9_line16a_18_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line16a_18_cpass
bit _zy_sva_b17;
wire  _zy_sva_key_type9_line16b_19_reset_or;
bit [0:0]  _zy_sva_key_type9_line16b_19_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line16b_19_ccheck
bit [0:0]  _zy_sva_key_type9_line16b_19_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line16b_19_cpass
bit _zy_sva_b18;
wire  _zy_sva_key_type9_line17a_20_reset_or;
bit [0:0]  _zy_sva_key_type9_line17a_20_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line17a_20_ccheck
bit [0:0]  _zy_sva_key_type9_line17a_20_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line17a_20_cpass
bit _zy_sva_b19;
wire  _zy_sva_key_type9_line17b_21_reset_or;
bit [0:0]  _zy_sva_key_type9_line17b_21_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line17b_21_ccheck
bit [0:0]  _zy_sva_key_type9_line17b_21_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line17b_21_cpass
bit _zy_sva_b20;
wire  _zy_sva_key_type9_line18a_22_reset_or;
bit [0:0]  _zy_sva_key_type9_line18a_22_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line18a_22_ccheck
bit [0:0]  _zy_sva_key_type9_line18a_22_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line18a_22_cpass
bit _zy_sva_b21;
wire  _zy_sva_key_type9_line18b_23_reset_or;
bit [0:0]  _zy_sva_key_type9_line18b_23_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line18b_23_ccheck
bit [0:0]  _zy_sva_key_type9_line18b_23_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line18b_23_cpass
bit _zy_sva_b22;
wire  _zy_sva_key_type9_line19a_24_reset_or;
bit [0:0]  _zy_sva_key_type9_line19a_24_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19a_24_ccheck
bit [0:0]  _zy_sva_key_type9_line19a_24_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19a_24_cpass
bit _zy_sva_b23;
wire  _zy_sva_key_type9_line19b_25_reset_or;
bit [0:0]  _zy_sva_key_type9_line19b_25_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19b_25_ccheck
bit [0:0]  _zy_sva_key_type9_line19b_25_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19b_25_cpass
bit _zy_sva_b24;
wire  _zy_sva_key_type9_line19c_26_reset_or;
bit [0:0]  _zy_sva_key_type9_line19c_26_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19c_26_ccheck
bit [0:0]  _zy_sva_key_type9_line19c_26_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19c_26_cpass
bit _zy_sva_b25;
wire  _zy_sva_key_type9_line19d_27_reset_or;
bit [0:0]  _zy_sva_key_type9_line19d_27_ccheck = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19d_27_ccheck
bit [0:0]  _zy_sva_key_type9_line19d_27_cpass = 1'b0;
// quickturn keep_net _zy_sva_key_type9_line19d_27_cpass
bit _zy_sva_b26;
wire  _zy_sva_guid_miss_aux_cmd_0_28_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_0_28_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_0_28_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_0_28_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_0_28_cpass
bit _zy_sva_b27;
wire  _zy_sva_guid_miss_aux_cmd_1_29_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_1_29_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_1_29_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_1_29_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_1_29_cpass
bit _zy_sva_b28;
wire  _zy_sva_guid_miss_aux_cmd_2_30_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_2_30_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_2_30_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_2_30_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_2_30_cpass
bit _zy_sva_b29;
wire  _zy_sva_guid_miss_aux_cmd_3_31_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_3_31_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_3_31_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_3_31_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_3_31_cpass
bit _zy_sva_b30;
wire  _zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass
bit _zy_sva_b31;
wire  _zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass
bit _zy_sva_b32;
wire  _zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass
bit _zy_sva_b33;
wire  _zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or;
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck
bit [0:0]  _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass = 1'b0;
// quickturn keep_net _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass
bit _zy_sva_b34;
wire  _zy_sva_iv_miss_aux_cmd_0_36_reset_or;
bit [0:0]  _zy_sva_iv_miss_aux_cmd_0_36_ccheck = 1'b0;
// quickturn keep_net _zy_sva_iv_miss_aux_cmd_0_36_ccheck
bit [0:0]  _zy_sva_iv_miss_aux_cmd_0_36_cpass = 1'b0;
// quickturn keep_net _zy_sva_iv_miss_aux_cmd_0_36_cpass
bit _zy_sva_b35;
wire  _zy_sva_iv_miss_aux_cmd_1_37_reset_or;
bit [0:0]  _zy_sva_iv_miss_aux_cmd_1_37_ccheck = 1'b0;
// quickturn keep_net _zy_sva_iv_miss_aux_cmd_1_37_ccheck
bit [0:0]  _zy_sva_iv_miss_aux_cmd_1_37_cpass = 1'b0;
// quickturn keep_net _zy_sva_iv_miss_aux_cmd_1_37_cpass
bit _zy_sva_b36;
wire  _zy_sva_iv_miss_aux_cmd_guid_38_reset_or;
bit [0:0]  _zy_sva_iv_miss_aux_cmd_guid_38_ccheck = 1'b0;
// quickturn keep_net _zy_sva_iv_miss_aux_cmd_guid_38_ccheck
bit [0:0]  _zy_sva_iv_miss_aux_cmd_guid_38_cpass = 1'b0;
// quickturn keep_net _zy_sva_iv_miss_aux_cmd_guid_38_cpass
bit _zy_sva_b37;
wire  _zy_sva_brcm_aux_cmd_39_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_39_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_39_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_39_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_39_cpass
bit _zy_sva_b38;
wire  _zy_sva_brcm_aux_cmd_iv_40_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_40_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_40_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_40_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_40_cpass
bit _zy_sva_b39;
wire  _zy_sva_brcm_aux_cmd_guid_41_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_41_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_41_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_41_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_41_cpass
bit _zy_sva_b40;
wire  _zy_sva_brcm_aux_cmd_guid_iv_42_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_42_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_42_cpass
bit _zy_sva_b41;
wire  _zy_sva_brcm_key_type_43_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_43_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_43_ccheck
bit [0:0]  _zy_sva_brcm_key_type_43_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_43_cpass
bit _zy_sva_b42;
wire  _zy_sva_brcm_aux_cmd_44_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_44_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_44_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_44_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_44_cpass
bit _zy_sva_b43;
wire  _zy_sva_brcm_aux_cmd_iv_45_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_45_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_45_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_45_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_45_cpass
bit _zy_sva_b44;
wire  _zy_sva_brcm_aux_cmd_guid_46_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_46_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_46_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_46_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_46_cpass
bit _zy_sva_b45;
wire  _zy_sva_brcm_aux_cmd_guid_iv_47_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_47_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_47_cpass
bit _zy_sva_b46;
wire  _zy_sva_brcm_key_type_48_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_48_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_48_ccheck
bit [0:0]  _zy_sva_brcm_key_type_48_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_48_cpass
bit _zy_sva_b47;
wire  _zy_sva_brcm_aux_cmd_49_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_49_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_49_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_49_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_49_cpass
bit _zy_sva_b48;
wire  _zy_sva_brcm_aux_cmd_iv_50_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_50_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_50_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_50_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_50_cpass
bit _zy_sva_b49;
wire  _zy_sva_brcm_aux_cmd_guid_51_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_51_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_51_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_51_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_51_cpass
bit _zy_sva_b50;
wire  _zy_sva_brcm_aux_cmd_guid_iv_52_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_52_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_52_cpass
bit _zy_sva_b51;
wire  _zy_sva_brcm_key_type_53_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_53_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_53_ccheck
bit [0:0]  _zy_sva_brcm_key_type_53_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_53_cpass
bit _zy_sva_b52;
wire  _zy_sva_brcm_aux_cmd_54_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_54_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_54_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_54_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_54_cpass
bit _zy_sva_b53;
wire  _zy_sva_brcm_aux_cmd_iv_55_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_55_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_55_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_55_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_55_cpass
bit _zy_sva_b54;
wire  _zy_sva_brcm_aux_cmd_guid_56_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_56_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_56_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_56_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_56_cpass
bit _zy_sva_b55;
wire  _zy_sva_brcm_aux_cmd_guid_iv_57_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_57_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_57_cpass
bit _zy_sva_b56;
wire  _zy_sva_brcm_key_type_58_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_58_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_58_ccheck
bit [0:0]  _zy_sva_brcm_key_type_58_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_58_cpass
bit _zy_sva_b57;
wire  _zy_sva_brcm_aux_cmd_59_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_59_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_59_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_59_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_59_cpass
bit _zy_sva_b58;
wire  _zy_sva_brcm_aux_cmd_iv_60_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_60_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_60_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_60_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_60_cpass
bit _zy_sva_b59;
wire  _zy_sva_brcm_aux_cmd_guid_61_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_61_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_61_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_61_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_61_cpass
bit _zy_sva_b60;
wire  _zy_sva_brcm_aux_cmd_guid_iv_62_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_62_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_62_cpass
bit _zy_sva_b61;
wire  _zy_sva_brcm_key_type_63_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_63_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_63_ccheck
bit [0:0]  _zy_sva_brcm_key_type_63_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_63_cpass
bit _zy_sva_b62;
wire  _zy_sva_brcm_aux_cmd_64_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_64_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_64_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_64_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_64_cpass
bit _zy_sva_b63;
wire  _zy_sva_brcm_aux_cmd_iv_65_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_65_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_65_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_65_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_65_cpass
bit _zy_sva_b64;
wire  _zy_sva_brcm_aux_cmd_guid_66_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_66_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_66_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_66_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_66_cpass
bit _zy_sva_b65;
wire  _zy_sva_brcm_aux_cmd_guid_iv_67_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_67_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_67_cpass
bit _zy_sva_b66;
wire  _zy_sva_brcm_key_type_68_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_68_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_68_ccheck
bit [0:0]  _zy_sva_brcm_key_type_68_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_68_cpass
bit _zy_sva_b67;
wire  _zy_sva_brcm_aux_cmd_69_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_69_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_69_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_69_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_69_cpass
bit _zy_sva_b68;
wire  _zy_sva_brcm_aux_cmd_iv_70_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_70_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_70_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_70_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_70_cpass
bit _zy_sva_b69;
wire  _zy_sva_brcm_aux_cmd_guid_71_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_71_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_71_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_71_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_71_cpass
bit _zy_sva_b70;
wire  _zy_sva_brcm_aux_cmd_guid_iv_72_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_72_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_72_cpass
bit _zy_sva_b71;
wire  _zy_sva_brcm_key_type_73_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_73_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_73_ccheck
bit [0:0]  _zy_sva_brcm_key_type_73_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_73_cpass
bit _zy_sva_b72;
wire  _zy_sva_brcm_aux_cmd_74_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_74_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_74_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_74_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_74_cpass
bit _zy_sva_b73;
wire  _zy_sva_brcm_aux_cmd_iv_75_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_75_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_75_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_75_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_75_cpass
bit _zy_sva_b74;
wire  _zy_sva_brcm_aux_cmd_guid_76_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_76_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_76_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_76_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_76_cpass
bit _zy_sva_b75;
wire  _zy_sva_brcm_aux_cmd_guid_iv_77_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_77_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_77_cpass
bit _zy_sva_b76;
wire  _zy_sva_brcm_key_type_78_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_78_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_78_ccheck
bit [0:0]  _zy_sva_brcm_key_type_78_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_78_cpass
bit _zy_sva_b77;
wire  _zy_sva_brcm_aux_cmd_79_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_79_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_79_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_79_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_79_cpass
bit _zy_sva_b78;
wire  _zy_sva_brcm_aux_cmd_iv_80_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_80_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_80_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_80_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_80_cpass
bit _zy_sva_b79;
wire  _zy_sva_brcm_aux_cmd_guid_81_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_81_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_81_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_81_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_81_cpass
bit _zy_sva_b80;
wire  _zy_sva_brcm_aux_cmd_guid_iv_82_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_82_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_82_cpass
bit _zy_sva_b81;
wire  _zy_sva_brcm_key_type_83_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_83_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_83_ccheck
bit [0:0]  _zy_sva_brcm_key_type_83_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_83_cpass
bit _zy_sva_b82;
wire  _zy_sva_brcm_aux_cmd_84_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_84_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_84_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_84_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_84_cpass
bit _zy_sva_b83;
wire  _zy_sva_brcm_aux_cmd_iv_85_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_85_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_85_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_85_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_85_cpass
bit _zy_sva_b84;
wire  _zy_sva_brcm_aux_cmd_guid_86_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_86_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_86_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_86_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_86_cpass
bit _zy_sva_b85;
wire  _zy_sva_brcm_aux_cmd_guid_iv_87_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_87_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_87_cpass
bit _zy_sva_b86;
wire  _zy_sva_brcm_key_type_88_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_88_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_88_ccheck
bit [0:0]  _zy_sva_brcm_key_type_88_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_88_cpass
bit _zy_sva_b87;
wire  _zy_sva_brcm_aux_cmd_89_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_89_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_89_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_89_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_89_cpass
bit _zy_sva_b88;
wire  _zy_sva_brcm_aux_cmd_iv_90_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_90_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_90_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_90_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_90_cpass
bit _zy_sva_b89;
wire  _zy_sva_brcm_aux_cmd_guid_91_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_91_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_91_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_91_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_91_cpass
bit _zy_sva_b90;
wire  _zy_sva_brcm_aux_cmd_guid_iv_92_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_92_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_92_cpass
bit _zy_sva_b91;
wire  _zy_sva_brcm_key_type_93_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_93_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_93_ccheck
bit [0:0]  _zy_sva_brcm_key_type_93_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_93_cpass
bit _zy_sva_b92;
wire  _zy_sva_brcm_aux_cmd_94_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_94_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_94_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_94_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_94_cpass
bit _zy_sva_b93;
wire  _zy_sva_brcm_aux_cmd_iv_95_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_95_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_95_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_95_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_95_cpass
bit _zy_sva_b94;
wire  _zy_sva_brcm_aux_cmd_guid_96_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_96_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_96_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_96_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_96_cpass
bit _zy_sva_b95;
wire  _zy_sva_brcm_aux_cmd_guid_iv_97_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_97_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_97_cpass
bit _zy_sva_b96;
wire  _zy_sva_brcm_key_type_98_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_98_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_98_ccheck
bit [0:0]  _zy_sva_brcm_key_type_98_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_98_cpass
bit _zy_sva_b97;
wire  _zy_sva_brcm_aux_cmd_99_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_99_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_99_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_99_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_99_cpass
bit _zy_sva_b98;
wire  _zy_sva_brcm_aux_cmd_iv_100_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_100_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_100_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_100_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_100_cpass
bit _zy_sva_b99;
wire  _zy_sva_brcm_aux_cmd_guid_101_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_101_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_101_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_101_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_101_cpass
bit _zy_sva_b100;
wire  _zy_sva_brcm_aux_cmd_guid_iv_102_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_102_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_102_cpass
bit _zy_sva_b101;
wire  _zy_sva_brcm_key_type_103_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_103_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_103_ccheck
bit [0:0]  _zy_sva_brcm_key_type_103_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_103_cpass
bit _zy_sva_b102;
wire  _zy_sva_brcm_aux_cmd_104_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_104_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_104_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_104_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_104_cpass
bit _zy_sva_b103;
wire  _zy_sva_brcm_aux_cmd_iv_105_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_105_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_105_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_iv_105_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_iv_105_cpass
bit _zy_sva_b104;
wire  _zy_sva_brcm_aux_cmd_guid_106_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_106_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_106_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_106_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_106_cpass
bit _zy_sva_b105;
wire  _zy_sva_brcm_aux_cmd_guid_iv_107_reset_or;
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck
bit [0:0]  _zy_sva_brcm_aux_cmd_guid_iv_107_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_aux_cmd_guid_iv_107_cpass
bit _zy_sva_b106;
wire  _zy_sva_brcm_key_type_108_reset_or;
bit [0:0]  _zy_sva_brcm_key_type_108_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_108_ccheck
bit [0:0]  _zy_sva_brcm_key_type_108_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_key_type_108_cpass
bit _zy_sva_b107;
wire  _zy_sva_brcm_kdf_ops_109_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_109_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_109_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_109_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_109_cpass
bit _zy_sva_b108;
wire  _zy_sva_brcm_kdf_ops_110_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_110_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_110_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_110_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_110_cpass
bit _zy_sva_b109;
wire  _zy_sva_brcm_kdf_ops_111_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_111_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_111_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_111_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_111_cpass
bit _zy_sva_b110;
wire  _zy_sva_brcm_kdf_ops_112_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_112_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_112_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_112_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_112_cpass
bit _zy_sva_b111;
wire  _zy_sva_brcm_kdf_ops_113_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_113_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_113_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_113_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_113_cpass
bit _zy_sva_b112;
wire  _zy_sva_brcm_kdf_ops_114_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_114_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_114_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_114_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_114_cpass
bit _zy_sva_b113;
wire  _zy_sva_brcm_kdf_ops_115_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_115_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_115_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_115_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_115_cpass
bit _zy_sva_b114;
wire  _zy_sva_brcm_kdf_ops_116_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_116_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_116_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_116_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_116_cpass
bit _zy_sva_b115;
wire  _zy_sva_brcm_kdf_ops_117_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_117_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_117_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_117_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_117_cpass
bit _zy_sva_b116;
wire  _zy_sva_brcm_kdf_ops_118_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_118_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_118_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_118_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_118_cpass
bit _zy_sva_b117;
wire  _zy_sva_brcm_kdf_ops_119_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_119_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_119_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_119_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_119_cpass
bit _zy_sva_b118;
wire  _zy_sva_brcm_kdf_ops_120_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_120_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_120_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_120_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_120_cpass
bit _zy_sva_b119;
wire  _zy_sva_brcm_kdf_ops_121_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_121_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_121_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_121_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_121_cpass
bit _zy_sva_b120;
wire  _zy_sva_brcm_kdf_ops_122_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_122_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_122_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_122_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_122_cpass
bit _zy_sva_b121;
wire  _zy_sva_brcm_kdf_ops_123_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_123_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_123_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_123_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_123_cpass
bit _zy_sva_b122;
wire  _zy_sva_brcm_kdf_ops_124_reset_or;
bit [0:0]  _zy_sva_brcm_kdf_ops_124_ccheck = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_124_ccheck
bit [0:0]  _zy_sva_brcm_kdf_ops_124_cpass = 1'b0;
// quickturn keep_net _zy_sva_brcm_kdf_ops_124_cpass
bit _zy_sva_b123;
wire  _zy_sva_null_gcm_125_reset_or;
bit [0:0]  _zy_sva_null_gcm_125_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_125_ccheck
bit [0:0]  _zy_sva_null_gcm_125_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_125_cpass
bit _zy_sva_b124;
wire  _zy_sva_sha_gcm_126_reset_or;
bit [0:0]  _zy_sva_sha_gcm_126_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_126_ccheck
bit [0:0]  _zy_sva_sha_gcm_126_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_126_cpass
bit _zy_sva_b125;
wire  _zy_sva_null_xts_127_reset_or;
bit [0:0]  _zy_sva_null_xts_127_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_xts_127_ccheck
bit [0:0]  _zy_sva_null_xts_127_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_xts_127_cpass
bit _zy_sva_b126;
wire  _zy_sva_sha_xts_128_reset_or;
bit [0:0]  _zy_sva_sha_xts_128_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_128_ccheck
bit [0:0]  _zy_sva_sha_xts_128_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_128_cpass
bit _zy_sva_b127;
wire  _zy_sva_null_null_129_reset_or;
bit [0:0]  _zy_sva_null_null_129_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_null_129_ccheck
bit [0:0]  _zy_sva_null_null_129_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_null_129_cpass
bit _zy_sva_b128;
wire  _zy_sva_sha_null_130_reset_or;
bit [0:0]  _zy_sva_sha_null_130_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_null_130_ccheck
bit [0:0]  _zy_sva_sha_null_130_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_null_130_cpass
bit _zy_sva_b129;
wire  _zy_sva_hmac_gcm_131_reset_or;
bit [0:0]  _zy_sva_hmac_gcm_131_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_131_ccheck
bit [0:0]  _zy_sva_hmac_gcm_131_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_131_cpass
bit _zy_sva_b130;
wire  _zy_sva_hmac_xts_132_reset_or;
bit [0:0]  _zy_sva_hmac_xts_132_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_132_ccheck
bit [0:0]  _zy_sva_hmac_xts_132_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_132_cpass
bit _zy_sva_b131;
wire  _zy_sva_hmac_null_133_reset_or;
bit [0:0]  _zy_sva_hmac_null_133_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_133_ccheck
bit [0:0]  _zy_sva_hmac_null_133_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_133_cpass
bit _zy_sva_b132;
wire  _zy_sva_null_gcm_134_reset_or;
bit [0:0]  _zy_sva_null_gcm_134_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_134_ccheck
bit [0:0]  _zy_sva_null_gcm_134_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_134_cpass
bit _zy_sva_b133;
wire  _zy_sva_sha_gcm_135_reset_or;
bit [0:0]  _zy_sva_sha_gcm_135_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_135_ccheck
bit [0:0]  _zy_sva_sha_gcm_135_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_135_cpass
bit _zy_sva_b134;
wire  _zy_sva_null_xts_136_reset_or;
bit [0:0]  _zy_sva_null_xts_136_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_xts_136_ccheck
bit [0:0]  _zy_sva_null_xts_136_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_xts_136_cpass
bit _zy_sva_b135;
wire  _zy_sva_sha_xts_137_reset_or;
bit [0:0]  _zy_sva_sha_xts_137_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_137_ccheck
bit [0:0]  _zy_sva_sha_xts_137_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_137_cpass
bit _zy_sva_b136;
wire  _zy_sva_null_null_138_reset_or;
bit [0:0]  _zy_sva_null_null_138_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_null_138_ccheck
bit [0:0]  _zy_sva_null_null_138_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_null_138_cpass
bit _zy_sva_b137;
wire  _zy_sva_sha_null_139_reset_or;
bit [0:0]  _zy_sva_sha_null_139_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_null_139_ccheck
bit [0:0]  _zy_sva_sha_null_139_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_null_139_cpass
bit _zy_sva_b138;
wire  _zy_sva_hmac_gcm_140_reset_or;
bit [0:0]  _zy_sva_hmac_gcm_140_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_140_ccheck
bit [0:0]  _zy_sva_hmac_gcm_140_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_140_cpass
bit _zy_sva_b139;
wire  _zy_sva_hmac_xts_141_reset_or;
bit [0:0]  _zy_sva_hmac_xts_141_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_141_ccheck
bit [0:0]  _zy_sva_hmac_xts_141_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_141_cpass
bit _zy_sva_b140;
wire  _zy_sva_hmac_null_142_reset_or;
bit [0:0]  _zy_sva_hmac_null_142_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_142_ccheck
bit [0:0]  _zy_sva_hmac_null_142_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_142_cpass
bit _zy_sva_b141;
wire  _zy_sva_null_gcm_143_reset_or;
bit [0:0]  _zy_sva_null_gcm_143_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_143_ccheck
bit [0:0]  _zy_sva_null_gcm_143_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_143_cpass
bit _zy_sva_b142;
wire  _zy_sva_sha_gcm_144_reset_or;
bit [0:0]  _zy_sva_sha_gcm_144_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_144_ccheck
bit [0:0]  _zy_sva_sha_gcm_144_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_144_cpass
bit _zy_sva_b143;
wire  _zy_sva_null_xts_145_reset_or;
bit [0:0]  _zy_sva_null_xts_145_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_xts_145_ccheck
bit [0:0]  _zy_sva_null_xts_145_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_xts_145_cpass
bit _zy_sva_b144;
wire  _zy_sva_sha_xts_146_reset_or;
bit [0:0]  _zy_sva_sha_xts_146_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_146_ccheck
bit [0:0]  _zy_sva_sha_xts_146_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_146_cpass
bit _zy_sva_b145;
wire  _zy_sva_null_null_147_reset_or;
bit [0:0]  _zy_sva_null_null_147_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_null_147_ccheck
bit [0:0]  _zy_sva_null_null_147_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_null_147_cpass
bit _zy_sva_b146;
wire  _zy_sva_sha_null_148_reset_or;
bit [0:0]  _zy_sva_sha_null_148_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_null_148_ccheck
bit [0:0]  _zy_sva_sha_null_148_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_null_148_cpass
bit _zy_sva_b147;
wire  _zy_sva_hmac_gcm_149_reset_or;
bit [0:0]  _zy_sva_hmac_gcm_149_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_149_ccheck
bit [0:0]  _zy_sva_hmac_gcm_149_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_149_cpass
bit _zy_sva_b148;
wire  _zy_sva_hmac_xts_150_reset_or;
bit [0:0]  _zy_sva_hmac_xts_150_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_150_ccheck
bit [0:0]  _zy_sva_hmac_xts_150_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_150_cpass
bit _zy_sva_b149;
wire  _zy_sva_hmac_null_151_reset_or;
bit [0:0]  _zy_sva_hmac_null_151_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_151_ccheck
bit [0:0]  _zy_sva_hmac_null_151_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_151_cpass
bit _zy_sva_b150;
wire  _zy_sva_null_gcm_152_reset_or;
bit [0:0]  _zy_sva_null_gcm_152_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_152_ccheck
bit [0:0]  _zy_sva_null_gcm_152_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_152_cpass
bit _zy_sva_b151;
wire  _zy_sva_sha_gcm_153_reset_or;
bit [0:0]  _zy_sva_sha_gcm_153_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_153_ccheck
bit [0:0]  _zy_sva_sha_gcm_153_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_153_cpass
bit _zy_sva_b152;
wire  _zy_sva_null_xts_154_reset_or;
bit [0:0]  _zy_sva_null_xts_154_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_xts_154_ccheck
bit [0:0]  _zy_sva_null_xts_154_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_xts_154_cpass
bit _zy_sva_b153;
wire  _zy_sva_sha_xts_155_reset_or;
bit [0:0]  _zy_sva_sha_xts_155_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_155_ccheck
bit [0:0]  _zy_sva_sha_xts_155_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_155_cpass
bit _zy_sva_b154;
wire  _zy_sva_null_null_156_reset_or;
bit [0:0]  _zy_sva_null_null_156_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_null_156_ccheck
bit [0:0]  _zy_sva_null_null_156_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_null_156_cpass
bit _zy_sva_b155;
wire  _zy_sva_sha_null_157_reset_or;
bit [0:0]  _zy_sva_sha_null_157_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_null_157_ccheck
bit [0:0]  _zy_sva_sha_null_157_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_null_157_cpass
bit _zy_sva_b156;
wire  _zy_sva_hmac_gcm_158_reset_or;
bit [0:0]  _zy_sva_hmac_gcm_158_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_158_ccheck
bit [0:0]  _zy_sva_hmac_gcm_158_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_158_cpass
bit _zy_sva_b157;
wire  _zy_sva_hmac_xts_159_reset_or;
bit [0:0]  _zy_sva_hmac_xts_159_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_159_ccheck
bit [0:0]  _zy_sva_hmac_xts_159_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_159_cpass
bit _zy_sva_b158;
wire  _zy_sva_hmac_null_160_reset_or;
bit [0:0]  _zy_sva_hmac_null_160_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_160_ccheck
bit [0:0]  _zy_sva_hmac_null_160_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_160_cpass
bit _zy_sva_b159;
wire  _zy_sva_null_gcm_161_reset_or;
bit [0:0]  _zy_sva_null_gcm_161_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_161_ccheck
bit [0:0]  _zy_sva_null_gcm_161_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_161_cpass
bit _zy_sva_b160;
wire  _zy_sva_sha_gcm_162_reset_or;
bit [0:0]  _zy_sva_sha_gcm_162_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_162_ccheck
bit [0:0]  _zy_sva_sha_gcm_162_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_162_cpass
bit _zy_sva_b161;
wire  _zy_sva_null_xts_163_reset_or;
bit [0:0]  _zy_sva_null_xts_163_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_xts_163_ccheck
bit [0:0]  _zy_sva_null_xts_163_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_xts_163_cpass
bit _zy_sva_b162;
wire  _zy_sva_sha_xts_164_reset_or;
bit [0:0]  _zy_sva_sha_xts_164_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_164_ccheck
bit [0:0]  _zy_sva_sha_xts_164_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_164_cpass
bit _zy_sva_b163;
wire  _zy_sva_null_null_165_reset_or;
bit [0:0]  _zy_sva_null_null_165_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_null_165_ccheck
bit [0:0]  _zy_sva_null_null_165_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_null_165_cpass
bit _zy_sva_b164;
wire  _zy_sva_sha_null_166_reset_or;
bit [0:0]  _zy_sva_sha_null_166_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_null_166_ccheck
bit [0:0]  _zy_sva_sha_null_166_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_null_166_cpass
bit _zy_sva_b165;
wire  _zy_sva_hmac_gcm_167_reset_or;
bit [0:0]  _zy_sva_hmac_gcm_167_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_167_ccheck
bit [0:0]  _zy_sva_hmac_gcm_167_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_167_cpass
bit _zy_sva_b166;
wire  _zy_sva_hmac_xts_168_reset_or;
bit [0:0]  _zy_sva_hmac_xts_168_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_168_ccheck
bit [0:0]  _zy_sva_hmac_xts_168_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_168_cpass
bit _zy_sva_b167;
wire  _zy_sva_hmac_null_169_reset_or;
bit [0:0]  _zy_sva_hmac_null_169_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_169_ccheck
bit [0:0]  _zy_sva_hmac_null_169_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_169_cpass
bit _zy_sva_b168;
wire  _zy_sva_null_gcm_170_reset_or;
bit [0:0]  _zy_sva_null_gcm_170_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_170_ccheck
bit [0:0]  _zy_sva_null_gcm_170_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_gcm_170_cpass
bit _zy_sva_b169;
wire  _zy_sva_sha_gcm_171_reset_or;
bit [0:0]  _zy_sva_sha_gcm_171_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_171_ccheck
bit [0:0]  _zy_sva_sha_gcm_171_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_gcm_171_cpass
bit _zy_sva_b170;
wire  _zy_sva_null_xts_172_reset_or;
bit [0:0]  _zy_sva_null_xts_172_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_xts_172_ccheck
bit [0:0]  _zy_sva_null_xts_172_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_xts_172_cpass
bit _zy_sva_b171;
wire  _zy_sva_sha_xts_173_reset_or;
bit [0:0]  _zy_sva_sha_xts_173_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_173_ccheck
bit [0:0]  _zy_sva_sha_xts_173_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_xts_173_cpass
bit _zy_sva_b172;
wire  _zy_sva_null_null_174_reset_or;
bit [0:0]  _zy_sva_null_null_174_ccheck = 1'b0;
// quickturn keep_net _zy_sva_null_null_174_ccheck
bit [0:0]  _zy_sva_null_null_174_cpass = 1'b0;
// quickturn keep_net _zy_sva_null_null_174_cpass
bit _zy_sva_b173;
wire  _zy_sva_sha_null_175_reset_or;
bit [0:0]  _zy_sva_sha_null_175_ccheck = 1'b0;
// quickturn keep_net _zy_sva_sha_null_175_ccheck
bit [0:0]  _zy_sva_sha_null_175_cpass = 1'b0;
// quickturn keep_net _zy_sva_sha_null_175_cpass
bit _zy_sva_b174;
wire  _zy_sva_hmac_gcm_176_reset_or;
bit [0:0]  _zy_sva_hmac_gcm_176_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_176_ccheck
bit [0:0]  _zy_sva_hmac_gcm_176_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_gcm_176_cpass
bit _zy_sva_b175;
wire  _zy_sva_hmac_xts_177_reset_or;
bit [0:0]  _zy_sva_hmac_xts_177_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_177_ccheck
bit [0:0]  _zy_sva_hmac_xts_177_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_xts_177_cpass
bit _zy_sva_b176;
wire  _zy_sva_hmac_null_178_reset_or;
bit [0:0]  _zy_sva_hmac_null_178_ccheck = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_178_ccheck
bit [0:0]  _zy_sva_hmac_null_178_cpass = 1'b0;
// quickturn keep_net _zy_sva_hmac_null_178_cpass
bit _zy_sva_b177;
// synopsys translate_off
wire  _sva_placeholder_clk;
wire  _sva_placeholder_expr;
// synopsys translate_on
wire  _zy_sva_b0_t;
wire  _zy_sva_b1_t;
wire  _zy_sva_b2_t;
wire  _zy_sva_b3_t;
wire  _zy_sva_b4_t;
wire  _zy_sva_b5_t;
wire  _zy_sva_b6_t;
wire  _zy_sva_b7_t;
wire  _zy_sva_b8_t;
wire  _zy_sva_b9_t;
wire  _zy_sva_b10_t;
wire  _zy_sva_b11_t;
wire  _zy_sva_b12_t;
wire  _zy_sva_b13_t;
wire  _zy_sva_b14_t;
wire  _zy_sva_b15_t;
wire  _zy_sva_b16_t;
wire  _zy_sva_b17_t;
wire  _zy_sva_b18_t;
wire  _zy_sva_b19_t;
wire  _zy_sva_b20_t;
wire  _zy_sva_b21_t;
wire  _zy_sva_b22_t;
wire  _zy_sva_b23_t;
wire  _zy_sva_b24_t;
wire  _zy_sva_b25_t;
wire  _zy_sva_b26_t;
wire  _zy_sva_b27_t;
wire  _zy_sva_b28_t;
wire  _zy_sva_b29_t;
wire  _zy_sva_b30_t;
wire  _zy_sva_b31_t;
wire  _zy_sva_b32_t;
wire  _zy_sva_b33_t;
wire  _zy_sva_b34_t;
wire  _zy_sva_b35_t;
wire  _zy_sva_b36_t;
wire  _zy_sva_b37_t;
wire  _zy_sva_b38_t;
wire  _zy_sva_b39_t;
wire  _zy_sva_b40_t;
wire  _zy_sva_b41_t;
wire  _zy_sva_b42_t;
wire  _zy_sva_b43_t;
wire  _zy_sva_b44_t;
wire  _zy_sva_b45_t;
wire  _zy_sva_b46_t;
wire  _zy_sva_b47_t;
wire  _zy_sva_b48_t;
wire  _zy_sva_b49_t;
wire  _zy_sva_b50_t;
wire  _zy_sva_b51_t;
wire  _zy_sva_b52_t;
wire  _zy_sva_b53_t;
wire  _zy_sva_b54_t;
wire  _zy_sva_b55_t;
wire  _zy_sva_b56_t;
wire  _zy_sva_b57_t;
wire  _zy_sva_b58_t;
wire  _zy_sva_b59_t;
wire  _zy_sva_b60_t;
wire  _zy_sva_b61_t;
wire  _zy_sva_b62_t;
wire  _zy_sva_b63_t;
wire  _zy_sva_b64_t;
wire  _zy_sva_b65_t;
wire  _zy_sva_b66_t;
wire  _zy_sva_b67_t;
wire  _zy_sva_b68_t;
wire  _zy_sva_b69_t;
wire  _zy_sva_b70_t;
wire  _zy_sva_b71_t;
wire  _zy_sva_b72_t;
wire  _zy_sva_b73_t;
wire  _zy_sva_b74_t;
wire  _zy_sva_b75_t;
wire  _zy_sva_b76_t;
wire  _zy_sva_b77_t;
wire  _zy_sva_b78_t;
wire  _zy_sva_b79_t;
wire  _zy_sva_b80_t;
wire  _zy_sva_b81_t;
wire  _zy_sva_b82_t;
wire  _zy_sva_b83_t;
wire  _zy_sva_b84_t;
wire  _zy_sva_b85_t;
wire  _zy_sva_b86_t;
wire  _zy_sva_b87_t;
wire  _zy_sva_b88_t;
wire  _zy_sva_b89_t;
wire  _zy_sva_b90_t;
wire  _zy_sva_b91_t;
wire  _zy_sva_b92_t;
wire  _zy_sva_b93_t;
wire  _zy_sva_b94_t;
wire  _zy_sva_b95_t;
wire  _zy_sva_b96_t;
wire  _zy_sva_b97_t;
wire  _zy_sva_b98_t;
wire  _zy_sva_b99_t;
wire  _zy_sva_b100_t;
wire  _zy_sva_b101_t;
wire  _zy_sva_b102_t;
wire  _zy_sva_b103_t;
wire  _zy_sva_b104_t;
wire  _zy_sva_b105_t;
wire  _zy_sva_b106_t;
wire  _zy_sva_b107_t;
wire  _zy_sva_b108_t;
wire  _zy_sva_b109_t;
wire  _zy_sva_b110_t;
wire  _zy_sva_b111_t;
wire  _zy_sva_b112_t;
wire  _zy_sva_b113_t;
wire  _zy_sva_b114_t;
wire  _zy_sva_b115_t;
wire  _zy_sva_b116_t;
wire  _zy_sva_b117_t;
wire  _zy_sva_b118_t;
wire  _zy_sva_b119_t;
wire  _zy_sva_b120_t;
wire  _zy_sva_b121_t;
wire  _zy_sva_b122_t;
wire  _zy_sva_b123_t;
wire  _zy_sva_b124_t;
wire  _zy_sva_b125_t;
wire  _zy_sva_b126_t;
wire  _zy_sva_b127_t;
wire  _zy_sva_b128_t;
wire  _zy_sva_b129_t;
wire  _zy_sva_b130_t;
wire  _zy_sva_b131_t;
wire  _zy_sva_b132_t;
wire  _zy_sva_b133_t;
wire  _zy_sva_b134_t;
wire  _zy_sva_b135_t;
wire  _zy_sva_b136_t;
wire  _zy_sva_b137_t;
wire  _zy_sva_b138_t;
wire  _zy_sva_b139_t;
wire  _zy_sva_b140_t;
wire  _zy_sva_b141_t;
wire  _zy_sva_b142_t;
wire  _zy_sva_b143_t;
wire  _zy_sva_b144_t;
wire  _zy_sva_b145_t;
wire  _zy_sva_b146_t;
wire  _zy_sva_b147_t;
wire  _zy_sva_b148_t;
wire  _zy_sva_b149_t;
wire  _zy_sva_b150_t;
wire  _zy_sva_b151_t;
wire  _zy_sva_b152_t;
wire  _zy_sva_b153_t;
wire  _zy_sva_b154_t;
wire  _zy_sva_b155_t;
wire  _zy_sva_b156_t;
wire  _zy_sva_b157_t;
wire  _zy_sva_b158_t;
wire  _zy_sva_b159_t;
wire  _zy_sva_b160_t;
wire  _zy_sva_b161_t;
wire  _zy_sva_b162_t;
wire  _zy_sva_b163_t;
wire  _zy_sva_b164_t;
wire  _zy_sva_b165_t;
wire  _zy_sva_b166_t;
wire  _zy_sva_b167_t;
wire  _zy_sva_b168_t;
wire  _zy_sva_b169_t;
wire  _zy_sva_b170_t;
wire  _zy_sva_b171_t;
wire  _zy_sva_b172_t;
wire  _zy_sva_b173_t;
wire  _zy_sva_b174_t;
wire  _zy_sva_b175_t;
wire  _zy_sva_b176_t;
wire  _zy_sva_b177_t;
reg [63:0] _zyL234_tfiRv52 ;
reg _zyL252_tfiRv53;
reg _zyL253_tfiRv54;
reg _zyL254_tfiRv55;
reg _zyL255_tfiRv56;
reg [63:0] _zyL288_tfiRv57 ;
reg [63:0] _zyL293_tfiRv58 ;
reg [63:0] _zyL301_tfiRv59 ;
reg [63:0] _zyL306_tfiRv60 ;
reg [63:0] _zyL313_tfiRv61 ;
reg [63:0] _zyL321_tfiRv62 ;
reg [63:0] _zyL327_tfiRv63 ;
reg [63:0] _zyL337_tfiRv64 ;
reg [63:0] _zyL346_tfiRv65 ;
reg [63:0] _zyL354_tfiRv66 ;
reg [63:0] _zyL359_tfiRv67 ;
reg [63:0] _zyL368_tfiRv68 ;
reg [63:0] _zyL373_tfiRv69 ;
reg [63:0] _zyL382_tfiRv70 ;
reg [63:0] _zyL390_tfiRv71 ;
reg [63:0] _zyL395_tfiRv72 ;
reg [63:0] _zyL410_tfiRv73 ;
reg _zyL485_tfiRv74;
reg _zyL486_tfiRv75;
reg _zyL489_tfiRv76;
reg _zyL489_tfiRv77;
reg _zyL492_tfiRv78;
reg [63:0] _zyL526_tfiRv79 ;
reg [63:0] _zyL527_tfiRv80 ;
reg [63:0] _zyL541_tfiRv81 ;
reg [63:0] _zyL542_tfiRv82 ;
reg [63:0] _zyL555_tfiRv83 ;
reg [63:0] _zyL556_tfiRv84 ;
reg [63:0] _zyL569_tfiRv85 ;
reg [63:0] _zyL570_tfiRv86 ;
assign  stitcher_sot = (stitcher_out.tuser == 8'b01);
assign  stitcher_eot = (stitcher_out.tuser == 8'b010);
assign  tlv_parser_idle = (stitcher_empty & (tlv_counter == 5'b0));
assign  tlv_parser_int_tlv_start_pulse = (fifo_in_valid & fifo_in.sot);
ixc_assign  #(1) _zz_strnp_0 (_zy_simnet_stitcher_rd_0_w$,stitcher_rd);
ixc_assign  #(71) _zz_strnp_1 (_zy_simnet_parser_kimreader_data_1_w$,parser_kimreader_data);
ixc_assign  #(71) _zz_strnp_2 (parser_kimreader_data,_zy_simnet_parser_kimreader_data_2_w$);
ixc_assign  #(71) _zz_strnp_3 (_zy_simnet_fifo_in_5_w$,fifo_in);
ixc_assign  #(1) _zz_strnp_4 (_zy_simnet_fifo_in_valid_6_w$,fifo_in_valid);
assign  _zy_simnet_cio_7 = 1'b0;
assign  _zy_sva_key_type0_line4_1_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type0_line5a_2_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type0_line5b_3_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line7a_4_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line7b_5_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line8a_6_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line8b_7_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line9_8_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line10_9_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line11a_10_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line11b_11_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line11c_12_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line11d_13_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line12a_14_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type1_line12b_15_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line14_16_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line15_17_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line16a_18_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line16b_19_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line17a_20_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line17b_21_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line18a_22_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line18b_23_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line19a_24_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line19b_25_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line19c_26_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_key_type9_line19d_27_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_0_28_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_1_29_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_2_30_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_3_31_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_iv_miss_aux_cmd_0_36_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_iv_miss_aux_cmd_1_37_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_iv_miss_aux_cmd_guid_38_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_39_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_40_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_41_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_42_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_43_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_44_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_45_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_46_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_47_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_48_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_49_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_50_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_51_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_52_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_53_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_54_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_55_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_56_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_57_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_58_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_59_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_60_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_61_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_62_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_63_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_64_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_65_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_66_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_67_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_68_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_69_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_70_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_71_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_72_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_73_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_74_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_75_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_76_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_77_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_78_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_79_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_80_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_81_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_82_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_83_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_84_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_85_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_86_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_87_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_88_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_89_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_90_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_91_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_92_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_93_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_94_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_95_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_96_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_97_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_98_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_99_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_100_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_101_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_102_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_103_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_104_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_iv_105_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_106_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_aux_cmd_guid_iv_107_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_key_type_108_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_109_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_110_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_111_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_112_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_113_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_114_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_115_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_116_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_117_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_118_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_119_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_120_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_121_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_122_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_123_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_brcm_kdf_ops_124_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_gcm_125_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_gcm_126_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_xts_127_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_xts_128_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_null_129_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_null_130_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_gcm_131_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_xts_132_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_null_133_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_gcm_134_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_gcm_135_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_xts_136_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_xts_137_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_null_138_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_null_139_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_gcm_140_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_xts_141_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_null_142_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_gcm_143_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_gcm_144_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_xts_145_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_xts_146_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_null_147_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_null_148_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_gcm_149_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_xts_150_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_null_151_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_gcm_152_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_gcm_153_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_xts_154_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_xts_155_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_null_156_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_null_157_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_gcm_158_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_xts_159_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_null_160_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_gcm_161_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_gcm_162_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_xts_163_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_xts_164_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_null_165_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_null_166_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_gcm_167_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_xts_168_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_null_169_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_gcm_170_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_gcm_171_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_xts_172_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_xts_173_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_null_null_174_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_sha_null_175_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_gcm_176_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_xts_177_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_hmac_null_178_reset_or = (rst_n !== 32'b01);
assign  _zy_sva_b0_t = ((((int_tlv_counter == IDX_KME_IVTWEAK) && ((aux_auth_op == HMAC_SHA2) || (aux_raw_auth_op == HMAC_SHA2))) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == NO_AUX_KEY));
assign  _zy_sva_b1_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op != HMAC_SHA2)) && (aux_raw_auth_op != HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == NO_AUX_KEY));
assign  _zy_sva_b2_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op != HMAC_SHA2)) && (aux_raw_auth_op != HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == NO_AUX_KEY));
assign  _zy_sva_b3_t = (((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == AUX_KEY_ONLY)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_GUID)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_RGUID));
assign  _zy_sva_b4_t = (((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == AUX_KEY_ONLY)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_GUID)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_RGUID));
assign  _zy_sva_b5_t = ((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == AUX_KEY_ONLY)) && ((aux_key_header.kdf_mode == KDF_MODE_COMB_GUID) || (aux_key_header.kdf_mode == KDF_MODE_COMB_RGUID)));
assign  _zy_sva_b6_t = ((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == AUX_KEY_ONLY)) && ((aux_key_header.kdf_mode == KDF_MODE_COMB_GUID) || (aux_key_header.kdf_mode == KDF_MODE_COMB_RGUID)));
assign  _zy_sva_b7_t = (((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == AUX_KEY_ONLY)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_GUID)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_RGUID));
assign  _zy_sva_b8_t = ((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == AUX_KEY_ONLY)) && ((aux_key_header.kdf_mode == KDF_MODE_COMB_GUID) || (aux_key_header.kdf_mode == KDF_MODE_COMB_RGUID)));
assign  _zy_sva_b9_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == AUX_KEY_ONLY));
assign  _zy_sva_b10_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == AUX_KEY_ONLY));
assign  _zy_sva_b11_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == AUX_KEY_ONLY));
assign  _zy_sva_b12_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == AUX_KEY_ONLY));
assign  _zy_sva_b13_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == AUX_KEY_ONLY));
assign  _zy_sva_b14_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == AUX_KEY_ONLY));
assign  _zy_sva_b15_t = (((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == ENC_DAK)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_GUID)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_RGUID));
assign  _zy_sva_b16_t = ((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == ENC_DAK)) && ((aux_key_header.kdf_mode == KDF_MODE_COMB_GUID) || (aux_key_header.kdf_mode == KDF_MODE_COMB_RGUID)));
assign  _zy_sva_b17_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == ENC_DAK));
assign  _zy_sva_b18_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == ENC_DAK));
assign  _zy_sva_b19_t = (((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == ENC_DAK)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_GUID)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_RGUID));
assign  _zy_sva_b20_t = (((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == ENC_DAK)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_GUID)) && (aux_key_header.kdf_mode != KDF_MODE_COMB_RGUID));
assign  _zy_sva_b21_t = ((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == ENC_DAK)) && ((aux_key_header.kdf_mode == KDF_MODE_COMB_GUID) || (aux_key_header.kdf_mode == KDF_MODE_COMB_RGUID)));
assign  _zy_sva_b22_t = ((((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == ENC_DAK)) && ((aux_key_header.kdf_mode == KDF_MODE_COMB_GUID) || (aux_key_header.kdf_mode == KDF_MODE_COMB_RGUID)));
assign  _zy_sva_b23_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == ENC_DAK));
assign  _zy_sva_b24_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == ENC_DAK));
assign  _zy_sva_b25_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == ENC_DAK));
assign  _zy_sva_b26_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == ENC_DAK));
assign  _zy_sva_b27_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD)) && (aux_key_header.kdf_mode == KDF_MODE_GUID)) && (aux_key_header.dek_key_op == KDF)) && (aux_key_header.dak_key_op == NOOP));
assign  _zy_sva_b28_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD)) && (aux_key_header.kdf_mode == KDF_MODE_GUID)) && (aux_key_header.dek_key_op == NOOP)) && (aux_key_header.dak_key_op == KDF));
assign  _zy_sva_b29_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD)) && (aux_key_header.kdf_mode == KDF_MODE_COMB_GUID)) && (aux_key_header.dek_key_op == KDF)) && (aux_key_header.dak_key_op == NOOP));
assign  _zy_sva_b30_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD)) && (aux_key_header.kdf_mode == KDF_MODE_COMB_GUID)) && (aux_key_header.dek_key_op == NOOP)) && (aux_key_header.dak_key_op == KDF));
assign  _zy_sva_b31_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD_IV)) && (aux_key_header.kdf_mode == KDF_MODE_GUID)) && (aux_key_header.dek_key_op == KDF)) && (aux_key_header.dak_key_op == NOOP));
assign  _zy_sva_b32_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD_IV)) && (aux_key_header.kdf_mode == KDF_MODE_GUID)) && (aux_key_header.dek_key_op == NOOP)) && (aux_key_header.dak_key_op == KDF));
assign  _zy_sva_b33_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD_IV)) && (aux_key_header.kdf_mode == KDF_MODE_COMB_GUID)) && (aux_key_header.dek_key_op == KDF)) && (aux_key_header.dak_key_op == NOOP));
assign  _zy_sva_b34_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD_IV)) && (aux_key_header.kdf_mode == KDF_MODE_COMB_GUID)) && (aux_key_header.dek_key_op == NOOP)) && (aux_key_header.dak_key_op == KDF));
assign  _zy_sva_b35_t = ((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD)) && (aux_iv_op == IV_INC)) && (aux_cipher_op == AES_GCM));
assign  _zy_sva_b36_t = ((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD)) && (aux_iv_op == IV_INC)) && (aux_cipher_op == AES_XTS_XEX));
assign  _zy_sva_b37_t = ((((int_tlv_counter == IDX_KME_IVTWEAK) && (tlv_type == AUX_CMD_GUID)) && (aux_iv_op == IV_INC)) && (aux_cipher_op == AES_XTS_XEX));
assign  _zy_sva_b38_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b0));
assign  _zy_sva_b39_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b0));
assign  _zy_sva_b40_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b0));
assign  _zy_sva_b41_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b0));
assign  _zy_sva_b42_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b0));
assign  _zy_sva_b43_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01));
assign  _zy_sva_b44_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01));
assign  _zy_sva_b45_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01));
assign  _zy_sva_b46_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01));
assign  _zy_sva_b47_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01));
assign  _zy_sva_b48_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b010));
assign  _zy_sva_b49_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b010));
assign  _zy_sva_b50_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b010));
assign  _zy_sva_b51_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b010));
assign  _zy_sva_b52_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b010));
assign  _zy_sva_b53_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b011));
assign  _zy_sva_b54_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b011));
assign  _zy_sva_b55_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b011));
assign  _zy_sva_b56_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b011));
assign  _zy_sva_b57_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b011));
assign  _zy_sva_b58_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b0100));
assign  _zy_sva_b59_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b0100));
assign  _zy_sva_b60_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b0100));
assign  _zy_sva_b61_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b0100));
assign  _zy_sva_b62_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b0100));
assign  _zy_sva_b63_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b0101));
assign  _zy_sva_b64_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b0101));
assign  _zy_sva_b65_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b0101));
assign  _zy_sva_b66_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b0101));
assign  _zy_sva_b67_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b0101));
assign  _zy_sva_b68_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b0110));
assign  _zy_sva_b69_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b0110));
assign  _zy_sva_b70_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b0110));
assign  _zy_sva_b71_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b0110));
assign  _zy_sva_b72_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b0110));
assign  _zy_sva_b73_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b0111));
assign  _zy_sva_b74_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b0111));
assign  _zy_sva_b75_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b0111));
assign  _zy_sva_b76_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b0111));
assign  _zy_sva_b77_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b0111));
assign  _zy_sva_b78_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01000));
assign  _zy_sva_b79_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01000));
assign  _zy_sva_b80_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01000));
assign  _zy_sva_b81_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01000));
assign  _zy_sva_b82_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01000));
assign  _zy_sva_b83_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01001));
assign  _zy_sva_b84_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01001));
assign  _zy_sva_b85_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01001));
assign  _zy_sva_b86_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01001));
assign  _zy_sva_b87_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01001));
assign  _zy_sva_b88_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01010));
assign  _zy_sva_b89_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01010));
assign  _zy_sva_b90_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01010));
assign  _zy_sva_b91_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01010));
assign  _zy_sva_b92_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01010));
assign  _zy_sva_b93_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01011));
assign  _zy_sva_b94_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01011));
assign  _zy_sva_b95_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01011));
assign  _zy_sva_b96_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01011));
assign  _zy_sva_b97_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01011));
assign  _zy_sva_b98_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01100));
assign  _zy_sva_b99_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01100));
assign  _zy_sva_b100_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01100));
assign  _zy_sva_b101_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01100));
assign  _zy_sva_b102_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01100));
assign  _zy_sva_b103_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010101)) & (tlv_word2.key_type == 32'b01101));
assign  _zy_sva_b104_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b010111)) & (tlv_word2.key_type == 32'b01101));
assign  _zy_sva_b105_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011000)) & (tlv_word2.key_type == 32'b01101));
assign  _zy_sva_b106_t = (((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_type == 32'b011001)) & (tlv_word2.key_type == 32'b01101));
assign  _zy_sva_b107_t = ((fifo_in_valid & (fifo_in.id == KME_WORD0)) & (tlv_word2.key_type == 32'b01101));
assign  _zy_sva_b108_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b0)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b109_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b0)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b110_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b0)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b111_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b0)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b112_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b01)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b113_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b01)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b114_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b01)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b115_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b01)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b116_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b010)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b117_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b010)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b118_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b010)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b119_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b010)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b120_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b011)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b121_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b011)) & (aux_key_header.dek_key_op == 32'b0)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b122_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b011)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b0));
assign  _zy_sva_b123_t = ((((fifo_in_valid & (fifo_in.id == KME_ERROR)) & (aux_key_header.kdf_mode == 32'b011)) & (aux_key_header.dek_key_op == 32'b01)) & (aux_key_header.dak_key_op == 32'b01));
assign  _zy_sva_b124_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b125_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b126_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b127_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b128_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b129_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b130_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b131_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b132_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b0111));
assign  _zy_sva_b133_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b134_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b135_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b136_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b137_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b138_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b139_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b140_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b141_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01000));
assign  _zy_sva_b142_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b143_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b144_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b145_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b146_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b147_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b148_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b149_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b150_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01010));
assign  _zy_sva_b151_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b152_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b153_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b154_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b155_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b156_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b157_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b158_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b159_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01011));
assign  _zy_sva_b160_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b161_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b162_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b163_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b164_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b165_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b166_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b167_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b168_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01100));
assign  _zy_sva_b169_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b170_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b171_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b172_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b173_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == AUTH_NULL)) && (aux_raw_auth_op == AUTH_NULL)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b174_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == SHA2)) && (aux_raw_auth_op == SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b175_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_GCM)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b176_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == AES_XTS_XEX)) && (aux_key_type == 32'b01101));
assign  _zy_sva_b177_t = (((((int_tlv_counter == IDX_KME_IVTWEAK) && (aux_auth_op == HMAC_SHA2)) && (aux_raw_auth_op == HMAC_SHA2)) && (aux_cipher_op == CPH_NULL)) && (aux_key_type == 32'b01101));
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b0 (_zy_sva_b0,_zy_sva_b0_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b1 (_zy_sva_b1,_zy_sva_b1_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b2 (_zy_sva_b2,_zy_sva_b2_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b3 (_zy_sva_b3,_zy_sva_b3_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b4 (_zy_sva_b4,_zy_sva_b4_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b5 (_zy_sva_b5,_zy_sva_b5_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b6 (_zy_sva_b6,_zy_sva_b6_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b7 (_zy_sva_b7,_zy_sva_b7_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b8 (_zy_sva_b8,_zy_sva_b8_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b9 (_zy_sva_b9,_zy_sva_b9_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b10 (_zy_sva_b10,_zy_sva_b10_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b11 (_zy_sva_b11,_zy_sva_b11_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b12 (_zy_sva_b12,_zy_sva_b12_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b13 (_zy_sva_b13,_zy_sva_b13_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b14 (_zy_sva_b14,_zy_sva_b14_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b15 (_zy_sva_b15,_zy_sva_b15_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b16 (_zy_sva_b16,_zy_sva_b16_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b17 (_zy_sva_b17,_zy_sva_b17_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b18 (_zy_sva_b18,_zy_sva_b18_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b19 (_zy_sva_b19,_zy_sva_b19_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b20 (_zy_sva_b20,_zy_sva_b20_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b21 (_zy_sva_b21,_zy_sva_b21_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b22 (_zy_sva_b22,_zy_sva_b22_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b23 (_zy_sva_b23,_zy_sva_b23_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b24 (_zy_sva_b24,_zy_sva_b24_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b25 (_zy_sva_b25,_zy_sva_b25_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b26 (_zy_sva_b26,_zy_sva_b26_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b27 (_zy_sva_b27,_zy_sva_b27_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b28 (_zy_sva_b28,_zy_sva_b28_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b29 (_zy_sva_b29,_zy_sva_b29_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b30 (_zy_sva_b30,_zy_sva_b30_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b31 (_zy_sva_b31,_zy_sva_b31_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b32 (_zy_sva_b32,_zy_sva_b32_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b33 (_zy_sva_b33,_zy_sva_b33_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b34 (_zy_sva_b34,_zy_sva_b34_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b35 (_zy_sva_b35,_zy_sva_b35_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b36 (_zy_sva_b36,_zy_sva_b36_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b37 (_zy_sva_b37,_zy_sva_b37_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b38 (_zy_sva_b38,_zy_sva_b38_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b39 (_zy_sva_b39,_zy_sva_b39_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b40 (_zy_sva_b40,_zy_sva_b40_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b41 (_zy_sva_b41,_zy_sva_b41_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b42 (_zy_sva_b42,_zy_sva_b42_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b43 (_zy_sva_b43,_zy_sva_b43_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b44 (_zy_sva_b44,_zy_sva_b44_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b45 (_zy_sva_b45,_zy_sva_b45_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b46 (_zy_sva_b46,_zy_sva_b46_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b47 (_zy_sva_b47,_zy_sva_b47_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b48 (_zy_sva_b48,_zy_sva_b48_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b49 (_zy_sva_b49,_zy_sva_b49_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b50 (_zy_sva_b50,_zy_sva_b50_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b51 (_zy_sva_b51,_zy_sva_b51_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b52 (_zy_sva_b52,_zy_sva_b52_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b53 (_zy_sva_b53,_zy_sva_b53_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b54 (_zy_sva_b54,_zy_sva_b54_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b55 (_zy_sva_b55,_zy_sva_b55_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b56 (_zy_sva_b56,_zy_sva_b56_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b57 (_zy_sva_b57,_zy_sva_b57_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b58 (_zy_sva_b58,_zy_sva_b58_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b59 (_zy_sva_b59,_zy_sva_b59_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b60 (_zy_sva_b60,_zy_sva_b60_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b61 (_zy_sva_b61,_zy_sva_b61_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b62 (_zy_sva_b62,_zy_sva_b62_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b63 (_zy_sva_b63,_zy_sva_b63_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b64 (_zy_sva_b64,_zy_sva_b64_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b65 (_zy_sva_b65,_zy_sva_b65_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b66 (_zy_sva_b66,_zy_sva_b66_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b67 (_zy_sva_b67,_zy_sva_b67_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b68 (_zy_sva_b68,_zy_sva_b68_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b69 (_zy_sva_b69,_zy_sva_b69_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b70 (_zy_sva_b70,_zy_sva_b70_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b71 (_zy_sva_b71,_zy_sva_b71_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b72 (_zy_sva_b72,_zy_sva_b72_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b73 (_zy_sva_b73,_zy_sva_b73_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b74 (_zy_sva_b74,_zy_sva_b74_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b75 (_zy_sva_b75,_zy_sva_b75_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b76 (_zy_sva_b76,_zy_sva_b76_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b77 (_zy_sva_b77,_zy_sva_b77_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b78 (_zy_sva_b78,_zy_sva_b78_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b79 (_zy_sva_b79,_zy_sva_b79_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b80 (_zy_sva_b80,_zy_sva_b80_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b81 (_zy_sva_b81,_zy_sva_b81_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b82 (_zy_sva_b82,_zy_sva_b82_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b83 (_zy_sva_b83,_zy_sva_b83_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b84 (_zy_sva_b84,_zy_sva_b84_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b85 (_zy_sva_b85,_zy_sva_b85_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b86 (_zy_sva_b86,_zy_sva_b86_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b87 (_zy_sva_b87,_zy_sva_b87_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b88 (_zy_sva_b88,_zy_sva_b88_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b89 (_zy_sva_b89,_zy_sva_b89_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b90 (_zy_sva_b90,_zy_sva_b90_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b91 (_zy_sva_b91,_zy_sva_b91_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b92 (_zy_sva_b92,_zy_sva_b92_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b93 (_zy_sva_b93,_zy_sva_b93_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b94 (_zy_sva_b94,_zy_sva_b94_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b95 (_zy_sva_b95,_zy_sva_b95_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b96 (_zy_sva_b96,_zy_sva_b96_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b97 (_zy_sva_b97,_zy_sva_b97_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b98 (_zy_sva_b98,_zy_sva_b98_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b99 (_zy_sva_b99,_zy_sva_b99_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b100 (_zy_sva_b100,_zy_sva_b100_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b101 (_zy_sva_b101,_zy_sva_b101_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b102 (_zy_sva_b102,_zy_sva_b102_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b103 (_zy_sva_b103,_zy_sva_b103_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b104 (_zy_sva_b104,_zy_sva_b104_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b105 (_zy_sva_b105,_zy_sva_b105_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b106 (_zy_sva_b106,_zy_sva_b106_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b107 (_zy_sva_b107,_zy_sva_b107_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b108 (_zy_sva_b108,_zy_sva_b108_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b109 (_zy_sva_b109,_zy_sva_b109_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b110 (_zy_sva_b110,_zy_sva_b110_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b111 (_zy_sva_b111,_zy_sva_b111_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b112 (_zy_sva_b112,_zy_sva_b112_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b113 (_zy_sva_b113,_zy_sva_b113_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b114 (_zy_sva_b114,_zy_sva_b114_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b115 (_zy_sva_b115,_zy_sva_b115_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b116 (_zy_sva_b116,_zy_sva_b116_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b117 (_zy_sva_b117,_zy_sva_b117_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b118 (_zy_sva_b118,_zy_sva_b118_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b119 (_zy_sva_b119,_zy_sva_b119_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b120 (_zy_sva_b120,_zy_sva_b120_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b121 (_zy_sva_b121,_zy_sva_b121_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b122 (_zy_sva_b122,_zy_sva_b122_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b123 (_zy_sva_b123,_zy_sva_b123_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b124 (_zy_sva_b124,_zy_sva_b124_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b125 (_zy_sva_b125,_zy_sva_b125_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b126 (_zy_sva_b126,_zy_sva_b126_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b127 (_zy_sva_b127,_zy_sva_b127_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b128 (_zy_sva_b128,_zy_sva_b128_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b129 (_zy_sva_b129,_zy_sva_b129_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b130 (_zy_sva_b130,_zy_sva_b130_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b131 (_zy_sva_b131,_zy_sva_b131_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b132 (_zy_sva_b132,_zy_sva_b132_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b133 (_zy_sva_b133,_zy_sva_b133_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b134 (_zy_sva_b134,_zy_sva_b134_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b135 (_zy_sva_b135,_zy_sva_b135_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b136 (_zy_sva_b136,_zy_sva_b136_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b137 (_zy_sva_b137,_zy_sva_b137_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b138 (_zy_sva_b138,_zy_sva_b138_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b139 (_zy_sva_b139,_zy_sva_b139_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b140 (_zy_sva_b140,_zy_sva_b140_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b141 (_zy_sva_b141,_zy_sva_b141_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b142 (_zy_sva_b142,_zy_sva_b142_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b143 (_zy_sva_b143,_zy_sva_b143_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b144 (_zy_sva_b144,_zy_sva_b144_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b145 (_zy_sva_b145,_zy_sva_b145_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b146 (_zy_sva_b146,_zy_sva_b146_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b147 (_zy_sva_b147,_zy_sva_b147_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b148 (_zy_sva_b148,_zy_sva_b148_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b149 (_zy_sva_b149,_zy_sva_b149_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b150 (_zy_sva_b150,_zy_sva_b150_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b151 (_zy_sva_b151,_zy_sva_b151_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b152 (_zy_sva_b152,_zy_sva_b152_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b153 (_zy_sva_b153,_zy_sva_b153_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b154 (_zy_sva_b154,_zy_sva_b154_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b155 (_zy_sva_b155,_zy_sva_b155_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b156 (_zy_sva_b156,_zy_sva_b156_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b157 (_zy_sva_b157,_zy_sva_b157_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b158 (_zy_sva_b158,_zy_sva_b158_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b159 (_zy_sva_b159,_zy_sva_b159_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b160 (_zy_sva_b160,_zy_sva_b160_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b161 (_zy_sva_b161,_zy_sva_b161_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b162 (_zy_sva_b162,_zy_sva_b162_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b163 (_zy_sva_b163,_zy_sva_b163_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b164 (_zy_sva_b164,_zy_sva_b164_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b165 (_zy_sva_b165,_zy_sva_b165_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b166 (_zy_sva_b166,_zy_sva_b166_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b167 (_zy_sva_b167,_zy_sva_b167_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b168 (_zy_sva_b168,_zy_sva_b168_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b169 (_zy_sva_b169,_zy_sva_b169_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b170 (_zy_sva_b170,_zy_sva_b170_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b171 (_zy_sva_b171,_zy_sva_b171_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b172 (_zy_sva_b172,_zy_sva_b172_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b173 (_zy_sva_b173,_zy_sva_b173_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b174 (_zy_sva_b174,_zy_sva_b174_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b175 (_zy_sva_b175,_zy_sva_b175_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b176 (_zy_sva_b176,_zy_sva_b176_t);
ixc_sample_logic #(32'b01,3)_zz_zy_sva_b177 (_zy_sva_b177,_zy_sva_b177_t);
cr_kme_fifo_xcm57 parser_fifo(
  .fifo_in_stall(fifo_in_stall) ,
  .fifo_out(_zy_simnet_parser_kimreader_data_2_w$) ,
  .fifo_out_valid(parser_kimreader_valid) ,
  .fifo_overflow(_zy_simnet_dio_3) ,
  .fifo_underflow(_zy_simnet_dio_4) ,
  .clk(clk) ,
  .rst_n(rst_n) ,
  .fifo_in(_zy_simnet_fifo_in_5_w$) ,
  .fifo_in_valid(_zy_simnet_fifo_in_valid_6_w$) ,
  .fifo_out_ack(kimreader_parser_ack) ,
  .fifo_in_stall_override(_zy_simnet_cio_7) ); 
always 
 @(posedge clk or posedge _zy_sva_key_type0_line4_1_reset_or)
  begin
   if (_zy_sva_key_type0_line4_1_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_1_1
     bit _zy_sva_nts_1_1_pass;
     _zy_sva_nts_1_1_pass = _zy_sva_b0;
     _zy_sva_key_type0_line4_1_ccheck = 1'b1;
     if (_zy_sva_nts_1_1_pass)
      begin
       _zy_sva_key_type0_line4_1_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type0_line5a_2_reset_or)
  begin
   if (_zy_sva_key_type0_line5a_2_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_2_1
     bit _zy_sva_nts_2_1_pass;
     _zy_sva_nts_2_1_pass = _zy_sva_b1;
     _zy_sva_key_type0_line5a_2_ccheck = 1'b1;
     if (_zy_sva_nts_2_1_pass)
      begin
       _zy_sva_key_type0_line5a_2_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type0_line5b_3_reset_or)
  begin
   if (_zy_sva_key_type0_line5b_3_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_3_1
     bit _zy_sva_nts_3_1_pass;
     _zy_sva_nts_3_1_pass = _zy_sva_b2;
     _zy_sva_key_type0_line5b_3_ccheck = 1'b1;
     if (_zy_sva_nts_3_1_pass)
      begin
       _zy_sva_key_type0_line5b_3_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line7a_4_reset_or)
  begin
   if (_zy_sva_key_type1_line7a_4_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_4_1
     bit _zy_sva_nts_4_1_pass;
     _zy_sva_nts_4_1_pass = _zy_sva_b3;
     _zy_sva_key_type1_line7a_4_ccheck = 1'b1;
     if (_zy_sva_nts_4_1_pass)
      begin
       _zy_sva_key_type1_line7a_4_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line7b_5_reset_or)
  begin
   if (_zy_sva_key_type1_line7b_5_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_5_1
     bit _zy_sva_nts_5_1_pass;
     _zy_sva_nts_5_1_pass = _zy_sva_b4;
     _zy_sva_key_type1_line7b_5_ccheck = 1'b1;
     if (_zy_sva_nts_5_1_pass)
      begin
       _zy_sva_key_type1_line7b_5_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line8a_6_reset_or)
  begin
   if (_zy_sva_key_type1_line8a_6_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_6_1
     bit _zy_sva_nts_6_1_pass;
     _zy_sva_nts_6_1_pass = _zy_sva_b5;
     _zy_sva_key_type1_line8a_6_ccheck = 1'b1;
     if (_zy_sva_nts_6_1_pass)
      begin
       _zy_sva_key_type1_line8a_6_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line8b_7_reset_or)
  begin
   if (_zy_sva_key_type1_line8b_7_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_7_1
     bit _zy_sva_nts_7_1_pass;
     _zy_sva_nts_7_1_pass = _zy_sva_b6;
     _zy_sva_key_type1_line8b_7_ccheck = 1'b1;
     if (_zy_sva_nts_7_1_pass)
      begin
       _zy_sva_key_type1_line8b_7_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line9_8_reset_or)
  begin
   if (_zy_sva_key_type1_line9_8_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_8_1
     bit _zy_sva_nts_8_1_pass;
     _zy_sva_nts_8_1_pass = _zy_sva_b7;
     _zy_sva_key_type1_line9_8_ccheck = 1'b1;
     if (_zy_sva_nts_8_1_pass)
      begin
       _zy_sva_key_type1_line9_8_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line10_9_reset_or)
  begin
   if (_zy_sva_key_type1_line10_9_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_9_1
     bit _zy_sva_nts_9_1_pass;
     _zy_sva_nts_9_1_pass = _zy_sva_b8;
     _zy_sva_key_type1_line10_9_ccheck = 1'b1;
     if (_zy_sva_nts_9_1_pass)
      begin
       _zy_sva_key_type1_line10_9_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line11a_10_reset_or)
  begin
   if (_zy_sva_key_type1_line11a_10_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_10_1
     bit _zy_sva_nts_10_1_pass;
     _zy_sva_nts_10_1_pass = _zy_sva_b9;
     _zy_sva_key_type1_line11a_10_ccheck = 1'b1;
     if (_zy_sva_nts_10_1_pass)
      begin
       _zy_sva_key_type1_line11a_10_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line11b_11_reset_or)
  begin
   if (_zy_sva_key_type1_line11b_11_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_11_1
     bit _zy_sva_nts_11_1_pass;
     _zy_sva_nts_11_1_pass = _zy_sva_b10;
     _zy_sva_key_type1_line11b_11_ccheck = 1'b1;
     if (_zy_sva_nts_11_1_pass)
      begin
       _zy_sva_key_type1_line11b_11_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line11c_12_reset_or)
  begin
   if (_zy_sva_key_type1_line11c_12_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_12_1
     bit _zy_sva_nts_12_1_pass;
     _zy_sva_nts_12_1_pass = _zy_sva_b11;
     _zy_sva_key_type1_line11c_12_ccheck = 1'b1;
     if (_zy_sva_nts_12_1_pass)
      begin
       _zy_sva_key_type1_line11c_12_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line11d_13_reset_or)
  begin
   if (_zy_sva_key_type1_line11d_13_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_13_1
     bit _zy_sva_nts_13_1_pass;
     _zy_sva_nts_13_1_pass = _zy_sva_b12;
     _zy_sva_key_type1_line11d_13_ccheck = 1'b1;
     if (_zy_sva_nts_13_1_pass)
      begin
       _zy_sva_key_type1_line11d_13_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line12a_14_reset_or)
  begin
   if (_zy_sva_key_type1_line12a_14_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_14_1
     bit _zy_sva_nts_14_1_pass;
     _zy_sva_nts_14_1_pass = _zy_sva_b13;
     _zy_sva_key_type1_line12a_14_ccheck = 1'b1;
     if (_zy_sva_nts_14_1_pass)
      begin
       _zy_sva_key_type1_line12a_14_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type1_line12b_15_reset_or)
  begin
   if (_zy_sva_key_type1_line12b_15_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_15_1
     bit _zy_sva_nts_15_1_pass;
     _zy_sva_nts_15_1_pass = _zy_sva_b14;
     _zy_sva_key_type1_line12b_15_ccheck = 1'b1;
     if (_zy_sva_nts_15_1_pass)
      begin
       _zy_sva_key_type1_line12b_15_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line14_16_reset_or)
  begin
   if (_zy_sva_key_type9_line14_16_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_16_1
     bit _zy_sva_nts_16_1_pass;
     _zy_sva_nts_16_1_pass = _zy_sva_b15;
     _zy_sva_key_type9_line14_16_ccheck = 1'b1;
     if (_zy_sva_nts_16_1_pass)
      begin
       _zy_sva_key_type9_line14_16_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line15_17_reset_or)
  begin
   if (_zy_sva_key_type9_line15_17_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_17_1
     bit _zy_sva_nts_17_1_pass;
     _zy_sva_nts_17_1_pass = _zy_sva_b16;
     _zy_sva_key_type9_line15_17_ccheck = 1'b1;
     if (_zy_sva_nts_17_1_pass)
      begin
       _zy_sva_key_type9_line15_17_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line16a_18_reset_or)
  begin
   if (_zy_sva_key_type9_line16a_18_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_18_1
     bit _zy_sva_nts_18_1_pass;
     _zy_sva_nts_18_1_pass = _zy_sva_b17;
     _zy_sva_key_type9_line16a_18_ccheck = 1'b1;
     if (_zy_sva_nts_18_1_pass)
      begin
       _zy_sva_key_type9_line16a_18_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line16b_19_reset_or)
  begin
   if (_zy_sva_key_type9_line16b_19_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_19_1
     bit _zy_sva_nts_19_1_pass;
     _zy_sva_nts_19_1_pass = _zy_sva_b18;
     _zy_sva_key_type9_line16b_19_ccheck = 1'b1;
     if (_zy_sva_nts_19_1_pass)
      begin
       _zy_sva_key_type9_line16b_19_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line17a_20_reset_or)
  begin
   if (_zy_sva_key_type9_line17a_20_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_20_1
     bit _zy_sva_nts_20_1_pass;
     _zy_sva_nts_20_1_pass = _zy_sva_b19;
     _zy_sva_key_type9_line17a_20_ccheck = 1'b1;
     if (_zy_sva_nts_20_1_pass)
      begin
       _zy_sva_key_type9_line17a_20_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line17b_21_reset_or)
  begin
   if (_zy_sva_key_type9_line17b_21_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_21_1
     bit _zy_sva_nts_21_1_pass;
     _zy_sva_nts_21_1_pass = _zy_sva_b20;
     _zy_sva_key_type9_line17b_21_ccheck = 1'b1;
     if (_zy_sva_nts_21_1_pass)
      begin
       _zy_sva_key_type9_line17b_21_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line18a_22_reset_or)
  begin
   if (_zy_sva_key_type9_line18a_22_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_22_1
     bit _zy_sva_nts_22_1_pass;
     _zy_sva_nts_22_1_pass = _zy_sva_b21;
     _zy_sva_key_type9_line18a_22_ccheck = 1'b1;
     if (_zy_sva_nts_22_1_pass)
      begin
       _zy_sva_key_type9_line18a_22_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line18b_23_reset_or)
  begin
   if (_zy_sva_key_type9_line18b_23_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_23_1
     bit _zy_sva_nts_23_1_pass;
     _zy_sva_nts_23_1_pass = _zy_sva_b22;
     _zy_sva_key_type9_line18b_23_ccheck = 1'b1;
     if (_zy_sva_nts_23_1_pass)
      begin
       _zy_sva_key_type9_line18b_23_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line19a_24_reset_or)
  begin
   if (_zy_sva_key_type9_line19a_24_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_24_1
     bit _zy_sva_nts_24_1_pass;
     _zy_sva_nts_24_1_pass = _zy_sva_b23;
     _zy_sva_key_type9_line19a_24_ccheck = 1'b1;
     if (_zy_sva_nts_24_1_pass)
      begin
       _zy_sva_key_type9_line19a_24_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line19b_25_reset_or)
  begin
   if (_zy_sva_key_type9_line19b_25_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_25_1
     bit _zy_sva_nts_25_1_pass;
     _zy_sva_nts_25_1_pass = _zy_sva_b24;
     _zy_sva_key_type9_line19b_25_ccheck = 1'b1;
     if (_zy_sva_nts_25_1_pass)
      begin
       _zy_sva_key_type9_line19b_25_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line19c_26_reset_or)
  begin
   if (_zy_sva_key_type9_line19c_26_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_26_1
     bit _zy_sva_nts_26_1_pass;
     _zy_sva_nts_26_1_pass = _zy_sva_b25;
     _zy_sva_key_type9_line19c_26_ccheck = 1'b1;
     if (_zy_sva_nts_26_1_pass)
      begin
       _zy_sva_key_type9_line19c_26_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_key_type9_line19d_27_reset_or)
  begin
   if (_zy_sva_key_type9_line19d_27_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_27_1
     bit _zy_sva_nts_27_1_pass;
     _zy_sva_nts_27_1_pass = _zy_sva_b26;
     _zy_sva_key_type9_line19d_27_ccheck = 1'b1;
     if (_zy_sva_nts_27_1_pass)
      begin
       _zy_sva_key_type9_line19d_27_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_0_28_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_0_28_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_28_1
     bit _zy_sva_nts_28_1_pass;
     _zy_sva_nts_28_1_pass = _zy_sva_b27;
     _zy_sva_guid_miss_aux_cmd_0_28_ccheck = 1'b1;
     if (_zy_sva_nts_28_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_0_28_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_1_29_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_1_29_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_29_1
     bit _zy_sva_nts_29_1_pass;
     _zy_sva_nts_29_1_pass = _zy_sva_b28;
     _zy_sva_guid_miss_aux_cmd_1_29_ccheck = 1'b1;
     if (_zy_sva_nts_29_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_1_29_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_2_30_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_2_30_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_30_1
     bit _zy_sva_nts_30_1_pass;
     _zy_sva_nts_30_1_pass = _zy_sva_b29;
     _zy_sva_guid_miss_aux_cmd_2_30_ccheck = 1'b1;
     if (_zy_sva_nts_30_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_2_30_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_3_31_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_3_31_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_31_1
     bit _zy_sva_nts_31_1_pass;
     _zy_sva_nts_31_1_pass = _zy_sva_b30;
     _zy_sva_guid_miss_aux_cmd_3_31_ccheck = 1'b1;
     if (_zy_sva_nts_31_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_3_31_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_iv_0_32_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_32_1
     bit _zy_sva_nts_32_1_pass;
     _zy_sva_nts_32_1_pass = _zy_sva_b31;
     _zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck = 1'b1;
     if (_zy_sva_nts_32_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_iv_0_32_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_iv_1_33_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_33_1
     bit _zy_sva_nts_33_1_pass;
     _zy_sva_nts_33_1_pass = _zy_sva_b32;
     _zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck = 1'b1;
     if (_zy_sva_nts_33_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_iv_1_33_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_iv_2_34_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_34_1
     bit _zy_sva_nts_34_1_pass;
     _zy_sva_nts_34_1_pass = _zy_sva_b33;
     _zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck = 1'b1;
     if (_zy_sva_nts_34_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_iv_2_34_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or)
  begin
   if (_zy_sva_guid_miss_aux_cmd_iv_3_35_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_35_1
     bit _zy_sva_nts_35_1_pass;
     _zy_sva_nts_35_1_pass = _zy_sva_b34;
     _zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck = 1'b1;
     if (_zy_sva_nts_35_1_pass)
      begin
       _zy_sva_guid_miss_aux_cmd_iv_3_35_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_iv_miss_aux_cmd_0_36_reset_or)
  begin
   if (_zy_sva_iv_miss_aux_cmd_0_36_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_36_1
     bit _zy_sva_nts_36_1_pass;
     _zy_sva_nts_36_1_pass = _zy_sva_b35;
     _zy_sva_iv_miss_aux_cmd_0_36_ccheck = 1'b1;
     if (_zy_sva_nts_36_1_pass)
      begin
       _zy_sva_iv_miss_aux_cmd_0_36_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_iv_miss_aux_cmd_1_37_reset_or)
  begin
   if (_zy_sva_iv_miss_aux_cmd_1_37_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_37_1
     bit _zy_sva_nts_37_1_pass;
     _zy_sva_nts_37_1_pass = _zy_sva_b36;
     _zy_sva_iv_miss_aux_cmd_1_37_ccheck = 1'b1;
     if (_zy_sva_nts_37_1_pass)
      begin
       _zy_sva_iv_miss_aux_cmd_1_37_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_iv_miss_aux_cmd_guid_38_reset_or)
  begin
   if (_zy_sva_iv_miss_aux_cmd_guid_38_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_38_1
     bit _zy_sva_nts_38_1_pass;
     _zy_sva_nts_38_1_pass = _zy_sva_b37;
     _zy_sva_iv_miss_aux_cmd_guid_38_ccheck = 1'b1;
     if (_zy_sva_nts_38_1_pass)
      begin
       _zy_sva_iv_miss_aux_cmd_guid_38_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_39_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_39_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_39_1
     bit _zy_sva_nts_39_1_pass;
     _zy_sva_nts_39_1_pass = _zy_sva_b38;
     _zy_sva_brcm_aux_cmd_39_ccheck = 1'b1;
     if (_zy_sva_nts_39_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_39_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_40_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_40_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_40_1
     bit _zy_sva_nts_40_1_pass;
     _zy_sva_nts_40_1_pass = _zy_sva_b39;
     _zy_sva_brcm_aux_cmd_iv_40_ccheck = 1'b1;
     if (_zy_sva_nts_40_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_40_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_41_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_41_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_41_1
     bit _zy_sva_nts_41_1_pass;
     _zy_sva_nts_41_1_pass = _zy_sva_b40;
     _zy_sva_brcm_aux_cmd_guid_41_ccheck = 1'b1;
     if (_zy_sva_nts_41_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_41_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_42_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_42_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_42_1
     bit _zy_sva_nts_42_1_pass;
     _zy_sva_nts_42_1_pass = _zy_sva_b41;
     _zy_sva_brcm_aux_cmd_guid_iv_42_ccheck = 1'b1;
     if (_zy_sva_nts_42_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_42_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_43_reset_or)
  begin
   if (_zy_sva_brcm_key_type_43_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_43_1
     bit _zy_sva_nts_43_1_pass;
     _zy_sva_nts_43_1_pass = _zy_sva_b42;
     _zy_sva_brcm_key_type_43_ccheck = 1'b1;
     if (_zy_sva_nts_43_1_pass)
      begin
       _zy_sva_brcm_key_type_43_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_44_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_44_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_44_1
     bit _zy_sva_nts_44_1_pass;
     _zy_sva_nts_44_1_pass = _zy_sva_b43;
     _zy_sva_brcm_aux_cmd_44_ccheck = 1'b1;
     if (_zy_sva_nts_44_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_44_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_45_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_45_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_45_1
     bit _zy_sva_nts_45_1_pass;
     _zy_sva_nts_45_1_pass = _zy_sva_b44;
     _zy_sva_brcm_aux_cmd_iv_45_ccheck = 1'b1;
     if (_zy_sva_nts_45_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_45_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_46_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_46_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_46_1
     bit _zy_sva_nts_46_1_pass;
     _zy_sva_nts_46_1_pass = _zy_sva_b45;
     _zy_sva_brcm_aux_cmd_guid_46_ccheck = 1'b1;
     if (_zy_sva_nts_46_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_46_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_47_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_47_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_47_1
     bit _zy_sva_nts_47_1_pass;
     _zy_sva_nts_47_1_pass = _zy_sva_b46;
     _zy_sva_brcm_aux_cmd_guid_iv_47_ccheck = 1'b1;
     if (_zy_sva_nts_47_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_47_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_48_reset_or)
  begin
   if (_zy_sva_brcm_key_type_48_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_48_1
     bit _zy_sva_nts_48_1_pass;
     _zy_sva_nts_48_1_pass = _zy_sva_b47;
     _zy_sva_brcm_key_type_48_ccheck = 1'b1;
     if (_zy_sva_nts_48_1_pass)
      begin
       _zy_sva_brcm_key_type_48_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_49_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_49_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_49_1
     bit _zy_sva_nts_49_1_pass;
     _zy_sva_nts_49_1_pass = _zy_sva_b48;
     _zy_sva_brcm_aux_cmd_49_ccheck = 1'b1;
     if (_zy_sva_nts_49_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_49_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_50_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_50_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_50_1
     bit _zy_sva_nts_50_1_pass;
     _zy_sva_nts_50_1_pass = _zy_sva_b49;
     _zy_sva_brcm_aux_cmd_iv_50_ccheck = 1'b1;
     if (_zy_sva_nts_50_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_50_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_51_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_51_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_51_1
     bit _zy_sva_nts_51_1_pass;
     _zy_sva_nts_51_1_pass = _zy_sva_b50;
     _zy_sva_brcm_aux_cmd_guid_51_ccheck = 1'b1;
     if (_zy_sva_nts_51_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_51_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_52_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_52_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_52_1
     bit _zy_sva_nts_52_1_pass;
     _zy_sva_nts_52_1_pass = _zy_sva_b51;
     _zy_sva_brcm_aux_cmd_guid_iv_52_ccheck = 1'b1;
     if (_zy_sva_nts_52_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_52_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_53_reset_or)
  begin
   if (_zy_sva_brcm_key_type_53_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_53_1
     bit _zy_sva_nts_53_1_pass;
     _zy_sva_nts_53_1_pass = _zy_sva_b52;
     _zy_sva_brcm_key_type_53_ccheck = 1'b1;
     if (_zy_sva_nts_53_1_pass)
      begin
       _zy_sva_brcm_key_type_53_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_54_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_54_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_54_1
     bit _zy_sva_nts_54_1_pass;
     _zy_sva_nts_54_1_pass = _zy_sva_b53;
     _zy_sva_brcm_aux_cmd_54_ccheck = 1'b1;
     if (_zy_sva_nts_54_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_54_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_55_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_55_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_55_1
     bit _zy_sva_nts_55_1_pass;
     _zy_sva_nts_55_1_pass = _zy_sva_b54;
     _zy_sva_brcm_aux_cmd_iv_55_ccheck = 1'b1;
     if (_zy_sva_nts_55_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_55_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_56_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_56_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_56_1
     bit _zy_sva_nts_56_1_pass;
     _zy_sva_nts_56_1_pass = _zy_sva_b55;
     _zy_sva_brcm_aux_cmd_guid_56_ccheck = 1'b1;
     if (_zy_sva_nts_56_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_56_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_57_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_57_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_57_1
     bit _zy_sva_nts_57_1_pass;
     _zy_sva_nts_57_1_pass = _zy_sva_b56;
     _zy_sva_brcm_aux_cmd_guid_iv_57_ccheck = 1'b1;
     if (_zy_sva_nts_57_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_57_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_58_reset_or)
  begin
   if (_zy_sva_brcm_key_type_58_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_58_1
     bit _zy_sva_nts_58_1_pass;
     _zy_sva_nts_58_1_pass = _zy_sva_b57;
     _zy_sva_brcm_key_type_58_ccheck = 1'b1;
     if (_zy_sva_nts_58_1_pass)
      begin
       _zy_sva_brcm_key_type_58_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_59_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_59_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_59_1
     bit _zy_sva_nts_59_1_pass;
     _zy_sva_nts_59_1_pass = _zy_sva_b58;
     _zy_sva_brcm_aux_cmd_59_ccheck = 1'b1;
     if (_zy_sva_nts_59_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_59_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_60_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_60_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_60_1
     bit _zy_sva_nts_60_1_pass;
     _zy_sva_nts_60_1_pass = _zy_sva_b59;
     _zy_sva_brcm_aux_cmd_iv_60_ccheck = 1'b1;
     if (_zy_sva_nts_60_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_60_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_61_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_61_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_61_1
     bit _zy_sva_nts_61_1_pass;
     _zy_sva_nts_61_1_pass = _zy_sva_b60;
     _zy_sva_brcm_aux_cmd_guid_61_ccheck = 1'b1;
     if (_zy_sva_nts_61_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_61_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_62_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_62_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_62_1
     bit _zy_sva_nts_62_1_pass;
     _zy_sva_nts_62_1_pass = _zy_sva_b61;
     _zy_sva_brcm_aux_cmd_guid_iv_62_ccheck = 1'b1;
     if (_zy_sva_nts_62_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_62_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_63_reset_or)
  begin
   if (_zy_sva_brcm_key_type_63_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_63_1
     bit _zy_sva_nts_63_1_pass;
     _zy_sva_nts_63_1_pass = _zy_sva_b62;
     _zy_sva_brcm_key_type_63_ccheck = 1'b1;
     if (_zy_sva_nts_63_1_pass)
      begin
       _zy_sva_brcm_key_type_63_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_64_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_64_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_64_1
     bit _zy_sva_nts_64_1_pass;
     _zy_sva_nts_64_1_pass = _zy_sva_b63;
     _zy_sva_brcm_aux_cmd_64_ccheck = 1'b1;
     if (_zy_sva_nts_64_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_64_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_65_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_65_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_65_1
     bit _zy_sva_nts_65_1_pass;
     _zy_sva_nts_65_1_pass = _zy_sva_b64;
     _zy_sva_brcm_aux_cmd_iv_65_ccheck = 1'b1;
     if (_zy_sva_nts_65_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_65_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_66_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_66_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_66_1
     bit _zy_sva_nts_66_1_pass;
     _zy_sva_nts_66_1_pass = _zy_sva_b65;
     _zy_sva_brcm_aux_cmd_guid_66_ccheck = 1'b1;
     if (_zy_sva_nts_66_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_66_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_67_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_67_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_67_1
     bit _zy_sva_nts_67_1_pass;
     _zy_sva_nts_67_1_pass = _zy_sva_b66;
     _zy_sva_brcm_aux_cmd_guid_iv_67_ccheck = 1'b1;
     if (_zy_sva_nts_67_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_67_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_68_reset_or)
  begin
   if (_zy_sva_brcm_key_type_68_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_68_1
     bit _zy_sva_nts_68_1_pass;
     _zy_sva_nts_68_1_pass = _zy_sva_b67;
     _zy_sva_brcm_key_type_68_ccheck = 1'b1;
     if (_zy_sva_nts_68_1_pass)
      begin
       _zy_sva_brcm_key_type_68_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_69_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_69_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_69_1
     bit _zy_sva_nts_69_1_pass;
     _zy_sva_nts_69_1_pass = _zy_sva_b68;
     _zy_sva_brcm_aux_cmd_69_ccheck = 1'b1;
     if (_zy_sva_nts_69_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_69_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_70_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_70_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_70_1
     bit _zy_sva_nts_70_1_pass;
     _zy_sva_nts_70_1_pass = _zy_sva_b69;
     _zy_sva_brcm_aux_cmd_iv_70_ccheck = 1'b1;
     if (_zy_sva_nts_70_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_70_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_71_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_71_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_71_1
     bit _zy_sva_nts_71_1_pass;
     _zy_sva_nts_71_1_pass = _zy_sva_b70;
     _zy_sva_brcm_aux_cmd_guid_71_ccheck = 1'b1;
     if (_zy_sva_nts_71_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_71_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_72_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_72_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_72_1
     bit _zy_sva_nts_72_1_pass;
     _zy_sva_nts_72_1_pass = _zy_sva_b71;
     _zy_sva_brcm_aux_cmd_guid_iv_72_ccheck = 1'b1;
     if (_zy_sva_nts_72_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_72_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_73_reset_or)
  begin
   if (_zy_sva_brcm_key_type_73_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_73_1
     bit _zy_sva_nts_73_1_pass;
     _zy_sva_nts_73_1_pass = _zy_sva_b72;
     _zy_sva_brcm_key_type_73_ccheck = 1'b1;
     if (_zy_sva_nts_73_1_pass)
      begin
       _zy_sva_brcm_key_type_73_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_74_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_74_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_74_1
     bit _zy_sva_nts_74_1_pass;
     _zy_sva_nts_74_1_pass = _zy_sva_b73;
     _zy_sva_brcm_aux_cmd_74_ccheck = 1'b1;
     if (_zy_sva_nts_74_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_74_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_75_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_75_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_75_1
     bit _zy_sva_nts_75_1_pass;
     _zy_sva_nts_75_1_pass = _zy_sva_b74;
     _zy_sva_brcm_aux_cmd_iv_75_ccheck = 1'b1;
     if (_zy_sva_nts_75_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_75_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_76_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_76_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_76_1
     bit _zy_sva_nts_76_1_pass;
     _zy_sva_nts_76_1_pass = _zy_sva_b75;
     _zy_sva_brcm_aux_cmd_guid_76_ccheck = 1'b1;
     if (_zy_sva_nts_76_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_76_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_77_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_77_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_77_1
     bit _zy_sva_nts_77_1_pass;
     _zy_sva_nts_77_1_pass = _zy_sva_b76;
     _zy_sva_brcm_aux_cmd_guid_iv_77_ccheck = 1'b1;
     if (_zy_sva_nts_77_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_77_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_78_reset_or)
  begin
   if (_zy_sva_brcm_key_type_78_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_78_1
     bit _zy_sva_nts_78_1_pass;
     _zy_sva_nts_78_1_pass = _zy_sva_b77;
     _zy_sva_brcm_key_type_78_ccheck = 1'b1;
     if (_zy_sva_nts_78_1_pass)
      begin
       _zy_sva_brcm_key_type_78_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_79_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_79_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_79_1
     bit _zy_sva_nts_79_1_pass;
     _zy_sva_nts_79_1_pass = _zy_sva_b78;
     _zy_sva_brcm_aux_cmd_79_ccheck = 1'b1;
     if (_zy_sva_nts_79_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_79_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_80_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_80_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_80_1
     bit _zy_sva_nts_80_1_pass;
     _zy_sva_nts_80_1_pass = _zy_sva_b79;
     _zy_sva_brcm_aux_cmd_iv_80_ccheck = 1'b1;
     if (_zy_sva_nts_80_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_80_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_81_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_81_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_81_1
     bit _zy_sva_nts_81_1_pass;
     _zy_sva_nts_81_1_pass = _zy_sva_b80;
     _zy_sva_brcm_aux_cmd_guid_81_ccheck = 1'b1;
     if (_zy_sva_nts_81_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_81_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_82_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_82_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_82_1
     bit _zy_sva_nts_82_1_pass;
     _zy_sva_nts_82_1_pass = _zy_sva_b81;
     _zy_sva_brcm_aux_cmd_guid_iv_82_ccheck = 1'b1;
     if (_zy_sva_nts_82_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_82_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_83_reset_or)
  begin
   if (_zy_sva_brcm_key_type_83_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_83_1
     bit _zy_sva_nts_83_1_pass;
     _zy_sva_nts_83_1_pass = _zy_sva_b82;
     _zy_sva_brcm_key_type_83_ccheck = 1'b1;
     if (_zy_sva_nts_83_1_pass)
      begin
       _zy_sva_brcm_key_type_83_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_84_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_84_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_84_1
     bit _zy_sva_nts_84_1_pass;
     _zy_sva_nts_84_1_pass = _zy_sva_b83;
     _zy_sva_brcm_aux_cmd_84_ccheck = 1'b1;
     if (_zy_sva_nts_84_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_84_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_85_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_85_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_85_1
     bit _zy_sva_nts_85_1_pass;
     _zy_sva_nts_85_1_pass = _zy_sva_b84;
     _zy_sva_brcm_aux_cmd_iv_85_ccheck = 1'b1;
     if (_zy_sva_nts_85_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_85_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_86_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_86_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_86_1
     bit _zy_sva_nts_86_1_pass;
     _zy_sva_nts_86_1_pass = _zy_sva_b85;
     _zy_sva_brcm_aux_cmd_guid_86_ccheck = 1'b1;
     if (_zy_sva_nts_86_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_86_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_87_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_87_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_87_1
     bit _zy_sva_nts_87_1_pass;
     _zy_sva_nts_87_1_pass = _zy_sva_b86;
     _zy_sva_brcm_aux_cmd_guid_iv_87_ccheck = 1'b1;
     if (_zy_sva_nts_87_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_87_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_88_reset_or)
  begin
   if (_zy_sva_brcm_key_type_88_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_88_1
     bit _zy_sva_nts_88_1_pass;
     _zy_sva_nts_88_1_pass = _zy_sva_b87;
     _zy_sva_brcm_key_type_88_ccheck = 1'b1;
     if (_zy_sva_nts_88_1_pass)
      begin
       _zy_sva_brcm_key_type_88_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_89_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_89_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_89_1
     bit _zy_sva_nts_89_1_pass;
     _zy_sva_nts_89_1_pass = _zy_sva_b88;
     _zy_sva_brcm_aux_cmd_89_ccheck = 1'b1;
     if (_zy_sva_nts_89_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_89_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_90_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_90_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_90_1
     bit _zy_sva_nts_90_1_pass;
     _zy_sva_nts_90_1_pass = _zy_sva_b89;
     _zy_sva_brcm_aux_cmd_iv_90_ccheck = 1'b1;
     if (_zy_sva_nts_90_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_90_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_91_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_91_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_91_1
     bit _zy_sva_nts_91_1_pass;
     _zy_sva_nts_91_1_pass = _zy_sva_b90;
     _zy_sva_brcm_aux_cmd_guid_91_ccheck = 1'b1;
     if (_zy_sva_nts_91_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_91_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_92_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_92_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_92_1
     bit _zy_sva_nts_92_1_pass;
     _zy_sva_nts_92_1_pass = _zy_sva_b91;
     _zy_sva_brcm_aux_cmd_guid_iv_92_ccheck = 1'b1;
     if (_zy_sva_nts_92_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_92_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_93_reset_or)
  begin
   if (_zy_sva_brcm_key_type_93_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_93_1
     bit _zy_sva_nts_93_1_pass;
     _zy_sva_nts_93_1_pass = _zy_sva_b92;
     _zy_sva_brcm_key_type_93_ccheck = 1'b1;
     if (_zy_sva_nts_93_1_pass)
      begin
       _zy_sva_brcm_key_type_93_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_94_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_94_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_94_1
     bit _zy_sva_nts_94_1_pass;
     _zy_sva_nts_94_1_pass = _zy_sva_b93;
     _zy_sva_brcm_aux_cmd_94_ccheck = 1'b1;
     if (_zy_sva_nts_94_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_94_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_95_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_95_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_95_1
     bit _zy_sva_nts_95_1_pass;
     _zy_sva_nts_95_1_pass = _zy_sva_b94;
     _zy_sva_brcm_aux_cmd_iv_95_ccheck = 1'b1;
     if (_zy_sva_nts_95_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_95_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_96_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_96_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_96_1
     bit _zy_sva_nts_96_1_pass;
     _zy_sva_nts_96_1_pass = _zy_sva_b95;
     _zy_sva_brcm_aux_cmd_guid_96_ccheck = 1'b1;
     if (_zy_sva_nts_96_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_96_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_97_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_97_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_97_1
     bit _zy_sva_nts_97_1_pass;
     _zy_sva_nts_97_1_pass = _zy_sva_b96;
     _zy_sva_brcm_aux_cmd_guid_iv_97_ccheck = 1'b1;
     if (_zy_sva_nts_97_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_97_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_98_reset_or)
  begin
   if (_zy_sva_brcm_key_type_98_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_98_1
     bit _zy_sva_nts_98_1_pass;
     _zy_sva_nts_98_1_pass = _zy_sva_b97;
     _zy_sva_brcm_key_type_98_ccheck = 1'b1;
     if (_zy_sva_nts_98_1_pass)
      begin
       _zy_sva_brcm_key_type_98_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_99_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_99_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_99_1
     bit _zy_sva_nts_99_1_pass;
     _zy_sva_nts_99_1_pass = _zy_sva_b98;
     _zy_sva_brcm_aux_cmd_99_ccheck = 1'b1;
     if (_zy_sva_nts_99_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_99_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_100_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_100_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_100_1
     bit _zy_sva_nts_100_1_pass;
     _zy_sva_nts_100_1_pass = _zy_sva_b99;
     _zy_sva_brcm_aux_cmd_iv_100_ccheck = 1'b1;
     if (_zy_sva_nts_100_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_100_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_101_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_101_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_101_1
     bit _zy_sva_nts_101_1_pass;
     _zy_sva_nts_101_1_pass = _zy_sva_b100;
     _zy_sva_brcm_aux_cmd_guid_101_ccheck = 1'b1;
     if (_zy_sva_nts_101_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_101_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_102_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_102_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_102_1
     bit _zy_sva_nts_102_1_pass;
     _zy_sva_nts_102_1_pass = _zy_sva_b101;
     _zy_sva_brcm_aux_cmd_guid_iv_102_ccheck = 1'b1;
     if (_zy_sva_nts_102_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_102_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_103_reset_or)
  begin
   if (_zy_sva_brcm_key_type_103_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_103_1
     bit _zy_sva_nts_103_1_pass;
     _zy_sva_nts_103_1_pass = _zy_sva_b102;
     _zy_sva_brcm_key_type_103_ccheck = 1'b1;
     if (_zy_sva_nts_103_1_pass)
      begin
       _zy_sva_brcm_key_type_103_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_104_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_104_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_104_1
     bit _zy_sva_nts_104_1_pass;
     _zy_sva_nts_104_1_pass = _zy_sva_b103;
     _zy_sva_brcm_aux_cmd_104_ccheck = 1'b1;
     if (_zy_sva_nts_104_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_104_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_iv_105_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_iv_105_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_105_1
     bit _zy_sva_nts_105_1_pass;
     _zy_sva_nts_105_1_pass = _zy_sva_b104;
     _zy_sva_brcm_aux_cmd_iv_105_ccheck = 1'b1;
     if (_zy_sva_nts_105_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_iv_105_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_106_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_106_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_106_1
     bit _zy_sva_nts_106_1_pass;
     _zy_sva_nts_106_1_pass = _zy_sva_b105;
     _zy_sva_brcm_aux_cmd_guid_106_ccheck = 1'b1;
     if (_zy_sva_nts_106_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_106_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_aux_cmd_guid_iv_107_reset_or)
  begin
   if (_zy_sva_brcm_aux_cmd_guid_iv_107_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_107_1
     bit _zy_sva_nts_107_1_pass;
     _zy_sva_nts_107_1_pass = _zy_sva_b106;
     _zy_sva_brcm_aux_cmd_guid_iv_107_ccheck = 1'b1;
     if (_zy_sva_nts_107_1_pass)
      begin
       _zy_sva_brcm_aux_cmd_guid_iv_107_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_key_type_108_reset_or)
  begin
   if (_zy_sva_brcm_key_type_108_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_108_1
     bit _zy_sva_nts_108_1_pass;
     _zy_sva_nts_108_1_pass = _zy_sva_b107;
     _zy_sva_brcm_key_type_108_ccheck = 1'b1;
     if (_zy_sva_nts_108_1_pass)
      begin
       _zy_sva_brcm_key_type_108_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_109_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_109_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_109_1
     bit _zy_sva_nts_109_1_pass;
     _zy_sva_nts_109_1_pass = _zy_sva_b108;
     _zy_sva_brcm_kdf_ops_109_ccheck = 1'b1;
     if (_zy_sva_nts_109_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_109_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_110_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_110_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_110_1
     bit _zy_sva_nts_110_1_pass;
     _zy_sva_nts_110_1_pass = _zy_sva_b109;
     _zy_sva_brcm_kdf_ops_110_ccheck = 1'b1;
     if (_zy_sva_nts_110_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_110_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_111_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_111_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_111_1
     bit _zy_sva_nts_111_1_pass;
     _zy_sva_nts_111_1_pass = _zy_sva_b110;
     _zy_sva_brcm_kdf_ops_111_ccheck = 1'b1;
     if (_zy_sva_nts_111_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_111_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_112_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_112_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_112_1
     bit _zy_sva_nts_112_1_pass;
     _zy_sva_nts_112_1_pass = _zy_sva_b111;
     _zy_sva_brcm_kdf_ops_112_ccheck = 1'b1;
     if (_zy_sva_nts_112_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_112_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_113_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_113_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_113_1
     bit _zy_sva_nts_113_1_pass;
     _zy_sva_nts_113_1_pass = _zy_sva_b112;
     _zy_sva_brcm_kdf_ops_113_ccheck = 1'b1;
     if (_zy_sva_nts_113_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_113_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_114_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_114_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_114_1
     bit _zy_sva_nts_114_1_pass;
     _zy_sva_nts_114_1_pass = _zy_sva_b113;
     _zy_sva_brcm_kdf_ops_114_ccheck = 1'b1;
     if (_zy_sva_nts_114_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_114_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_115_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_115_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_115_1
     bit _zy_sva_nts_115_1_pass;
     _zy_sva_nts_115_1_pass = _zy_sva_b114;
     _zy_sva_brcm_kdf_ops_115_ccheck = 1'b1;
     if (_zy_sva_nts_115_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_115_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_116_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_116_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_116_1
     bit _zy_sva_nts_116_1_pass;
     _zy_sva_nts_116_1_pass = _zy_sva_b115;
     _zy_sva_brcm_kdf_ops_116_ccheck = 1'b1;
     if (_zy_sva_nts_116_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_116_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_117_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_117_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_117_1
     bit _zy_sva_nts_117_1_pass;
     _zy_sva_nts_117_1_pass = _zy_sva_b116;
     _zy_sva_brcm_kdf_ops_117_ccheck = 1'b1;
     if (_zy_sva_nts_117_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_117_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_118_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_118_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_118_1
     bit _zy_sva_nts_118_1_pass;
     _zy_sva_nts_118_1_pass = _zy_sva_b117;
     _zy_sva_brcm_kdf_ops_118_ccheck = 1'b1;
     if (_zy_sva_nts_118_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_118_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_119_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_119_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_119_1
     bit _zy_sva_nts_119_1_pass;
     _zy_sva_nts_119_1_pass = _zy_sva_b118;
     _zy_sva_brcm_kdf_ops_119_ccheck = 1'b1;
     if (_zy_sva_nts_119_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_119_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_120_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_120_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_120_1
     bit _zy_sva_nts_120_1_pass;
     _zy_sva_nts_120_1_pass = _zy_sva_b119;
     _zy_sva_brcm_kdf_ops_120_ccheck = 1'b1;
     if (_zy_sva_nts_120_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_120_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_121_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_121_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_121_1
     bit _zy_sva_nts_121_1_pass;
     _zy_sva_nts_121_1_pass = _zy_sva_b120;
     _zy_sva_brcm_kdf_ops_121_ccheck = 1'b1;
     if (_zy_sva_nts_121_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_121_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_122_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_122_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_122_1
     bit _zy_sva_nts_122_1_pass;
     _zy_sva_nts_122_1_pass = _zy_sva_b121;
     _zy_sva_brcm_kdf_ops_122_ccheck = 1'b1;
     if (_zy_sva_nts_122_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_122_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_123_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_123_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_123_1
     bit _zy_sva_nts_123_1_pass;
     _zy_sva_nts_123_1_pass = _zy_sva_b122;
     _zy_sva_brcm_kdf_ops_123_ccheck = 1'b1;
     if (_zy_sva_nts_123_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_123_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_brcm_kdf_ops_124_reset_or)
  begin
   if (_zy_sva_brcm_kdf_ops_124_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_124_1
     bit _zy_sva_nts_124_1_pass;
     _zy_sva_nts_124_1_pass = _zy_sva_b123;
     _zy_sva_brcm_kdf_ops_124_ccheck = 1'b1;
     if (_zy_sva_nts_124_1_pass)
      begin
       _zy_sva_brcm_kdf_ops_124_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_gcm_125_reset_or)
  begin
   if (_zy_sva_null_gcm_125_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_125_1
     bit _zy_sva_nts_125_1_pass;
     _zy_sva_nts_125_1_pass = _zy_sva_b124;
     _zy_sva_null_gcm_125_ccheck = 1'b1;
     if (_zy_sva_nts_125_1_pass)
      begin
       _zy_sva_null_gcm_125_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_gcm_126_reset_or)
  begin
   if (_zy_sva_sha_gcm_126_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_126_1
     bit _zy_sva_nts_126_1_pass;
     _zy_sva_nts_126_1_pass = _zy_sva_b125;
     _zy_sva_sha_gcm_126_ccheck = 1'b1;
     if (_zy_sva_nts_126_1_pass)
      begin
       _zy_sva_sha_gcm_126_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_xts_127_reset_or)
  begin
   if (_zy_sva_null_xts_127_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_127_1
     bit _zy_sva_nts_127_1_pass;
     _zy_sva_nts_127_1_pass = _zy_sva_b126;
     _zy_sva_null_xts_127_ccheck = 1'b1;
     if (_zy_sva_nts_127_1_pass)
      begin
       _zy_sva_null_xts_127_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_xts_128_reset_or)
  begin
   if (_zy_sva_sha_xts_128_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_128_1
     bit _zy_sva_nts_128_1_pass;
     _zy_sva_nts_128_1_pass = _zy_sva_b127;
     _zy_sva_sha_xts_128_ccheck = 1'b1;
     if (_zy_sva_nts_128_1_pass)
      begin
       _zy_sva_sha_xts_128_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_null_129_reset_or)
  begin
   if (_zy_sva_null_null_129_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_129_1
     bit _zy_sva_nts_129_1_pass;
     _zy_sva_nts_129_1_pass = _zy_sva_b128;
     _zy_sva_null_null_129_ccheck = 1'b1;
     if (_zy_sva_nts_129_1_pass)
      begin
       _zy_sva_null_null_129_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_null_130_reset_or)
  begin
   if (_zy_sva_sha_null_130_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_130_1
     bit _zy_sva_nts_130_1_pass;
     _zy_sva_nts_130_1_pass = _zy_sva_b129;
     _zy_sva_sha_null_130_ccheck = 1'b1;
     if (_zy_sva_nts_130_1_pass)
      begin
       _zy_sva_sha_null_130_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_gcm_131_reset_or)
  begin
   if (_zy_sva_hmac_gcm_131_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_131_1
     bit _zy_sva_nts_131_1_pass;
     _zy_sva_nts_131_1_pass = _zy_sva_b130;
     _zy_sva_hmac_gcm_131_ccheck = 1'b1;
     if (_zy_sva_nts_131_1_pass)
      begin
       _zy_sva_hmac_gcm_131_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_xts_132_reset_or)
  begin
   if (_zy_sva_hmac_xts_132_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_132_1
     bit _zy_sva_nts_132_1_pass;
     _zy_sva_nts_132_1_pass = _zy_sva_b131;
     _zy_sva_hmac_xts_132_ccheck = 1'b1;
     if (_zy_sva_nts_132_1_pass)
      begin
       _zy_sva_hmac_xts_132_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_null_133_reset_or)
  begin
   if (_zy_sva_hmac_null_133_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_133_1
     bit _zy_sva_nts_133_1_pass;
     _zy_sva_nts_133_1_pass = _zy_sva_b132;
     _zy_sva_hmac_null_133_ccheck = 1'b1;
     if (_zy_sva_nts_133_1_pass)
      begin
       _zy_sva_hmac_null_133_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_gcm_134_reset_or)
  begin
   if (_zy_sva_null_gcm_134_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_134_1
     bit _zy_sva_nts_134_1_pass;
     _zy_sva_nts_134_1_pass = _zy_sva_b133;
     _zy_sva_null_gcm_134_ccheck = 1'b1;
     if (_zy_sva_nts_134_1_pass)
      begin
       _zy_sva_null_gcm_134_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_gcm_135_reset_or)
  begin
   if (_zy_sva_sha_gcm_135_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_135_1
     bit _zy_sva_nts_135_1_pass;
     _zy_sva_nts_135_1_pass = _zy_sva_b134;
     _zy_sva_sha_gcm_135_ccheck = 1'b1;
     if (_zy_sva_nts_135_1_pass)
      begin
       _zy_sva_sha_gcm_135_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_xts_136_reset_or)
  begin
   if (_zy_sva_null_xts_136_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_136_1
     bit _zy_sva_nts_136_1_pass;
     _zy_sva_nts_136_1_pass = _zy_sva_b135;
     _zy_sva_null_xts_136_ccheck = 1'b1;
     if (_zy_sva_nts_136_1_pass)
      begin
       _zy_sva_null_xts_136_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_xts_137_reset_or)
  begin
   if (_zy_sva_sha_xts_137_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_137_1
     bit _zy_sva_nts_137_1_pass;
     _zy_sva_nts_137_1_pass = _zy_sva_b136;
     _zy_sva_sha_xts_137_ccheck = 1'b1;
     if (_zy_sva_nts_137_1_pass)
      begin
       _zy_sva_sha_xts_137_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_null_138_reset_or)
  begin
   if (_zy_sva_null_null_138_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_138_1
     bit _zy_sva_nts_138_1_pass;
     _zy_sva_nts_138_1_pass = _zy_sva_b137;
     _zy_sva_null_null_138_ccheck = 1'b1;
     if (_zy_sva_nts_138_1_pass)
      begin
       _zy_sva_null_null_138_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_null_139_reset_or)
  begin
   if (_zy_sva_sha_null_139_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_139_1
     bit _zy_sva_nts_139_1_pass;
     _zy_sva_nts_139_1_pass = _zy_sva_b138;
     _zy_sva_sha_null_139_ccheck = 1'b1;
     if (_zy_sva_nts_139_1_pass)
      begin
       _zy_sva_sha_null_139_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_gcm_140_reset_or)
  begin
   if (_zy_sva_hmac_gcm_140_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_140_1
     bit _zy_sva_nts_140_1_pass;
     _zy_sva_nts_140_1_pass = _zy_sva_b139;
     _zy_sva_hmac_gcm_140_ccheck = 1'b1;
     if (_zy_sva_nts_140_1_pass)
      begin
       _zy_sva_hmac_gcm_140_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_xts_141_reset_or)
  begin
   if (_zy_sva_hmac_xts_141_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_141_1
     bit _zy_sva_nts_141_1_pass;
     _zy_sva_nts_141_1_pass = _zy_sva_b140;
     _zy_sva_hmac_xts_141_ccheck = 1'b1;
     if (_zy_sva_nts_141_1_pass)
      begin
       _zy_sva_hmac_xts_141_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_null_142_reset_or)
  begin
   if (_zy_sva_hmac_null_142_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_142_1
     bit _zy_sva_nts_142_1_pass;
     _zy_sva_nts_142_1_pass = _zy_sva_b141;
     _zy_sva_hmac_null_142_ccheck = 1'b1;
     if (_zy_sva_nts_142_1_pass)
      begin
       _zy_sva_hmac_null_142_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_gcm_143_reset_or)
  begin
   if (_zy_sva_null_gcm_143_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_143_1
     bit _zy_sva_nts_143_1_pass;
     _zy_sva_nts_143_1_pass = _zy_sva_b142;
     _zy_sva_null_gcm_143_ccheck = 1'b1;
     if (_zy_sva_nts_143_1_pass)
      begin
       _zy_sva_null_gcm_143_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_gcm_144_reset_or)
  begin
   if (_zy_sva_sha_gcm_144_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_144_1
     bit _zy_sva_nts_144_1_pass;
     _zy_sva_nts_144_1_pass = _zy_sva_b143;
     _zy_sva_sha_gcm_144_ccheck = 1'b1;
     if (_zy_sva_nts_144_1_pass)
      begin
       _zy_sva_sha_gcm_144_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_xts_145_reset_or)
  begin
   if (_zy_sva_null_xts_145_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_145_1
     bit _zy_sva_nts_145_1_pass;
     _zy_sva_nts_145_1_pass = _zy_sva_b144;
     _zy_sva_null_xts_145_ccheck = 1'b1;
     if (_zy_sva_nts_145_1_pass)
      begin
       _zy_sva_null_xts_145_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_xts_146_reset_or)
  begin
   if (_zy_sva_sha_xts_146_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_146_1
     bit _zy_sva_nts_146_1_pass;
     _zy_sva_nts_146_1_pass = _zy_sva_b145;
     _zy_sva_sha_xts_146_ccheck = 1'b1;
     if (_zy_sva_nts_146_1_pass)
      begin
       _zy_sva_sha_xts_146_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_null_147_reset_or)
  begin
   if (_zy_sva_null_null_147_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_147_1
     bit _zy_sva_nts_147_1_pass;
     _zy_sva_nts_147_1_pass = _zy_sva_b146;
     _zy_sva_null_null_147_ccheck = 1'b1;
     if (_zy_sva_nts_147_1_pass)
      begin
       _zy_sva_null_null_147_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_null_148_reset_or)
  begin
   if (_zy_sva_sha_null_148_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_148_1
     bit _zy_sva_nts_148_1_pass;
     _zy_sva_nts_148_1_pass = _zy_sva_b147;
     _zy_sva_sha_null_148_ccheck = 1'b1;
     if (_zy_sva_nts_148_1_pass)
      begin
       _zy_sva_sha_null_148_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_gcm_149_reset_or)
  begin
   if (_zy_sva_hmac_gcm_149_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_149_1
     bit _zy_sva_nts_149_1_pass;
     _zy_sva_nts_149_1_pass = _zy_sva_b148;
     _zy_sva_hmac_gcm_149_ccheck = 1'b1;
     if (_zy_sva_nts_149_1_pass)
      begin
       _zy_sva_hmac_gcm_149_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_xts_150_reset_or)
  begin
   if (_zy_sva_hmac_xts_150_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_150_1
     bit _zy_sva_nts_150_1_pass;
     _zy_sva_nts_150_1_pass = _zy_sva_b149;
     _zy_sva_hmac_xts_150_ccheck = 1'b1;
     if (_zy_sva_nts_150_1_pass)
      begin
       _zy_sva_hmac_xts_150_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_null_151_reset_or)
  begin
   if (_zy_sva_hmac_null_151_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_151_1
     bit _zy_sva_nts_151_1_pass;
     _zy_sva_nts_151_1_pass = _zy_sva_b150;
     _zy_sva_hmac_null_151_ccheck = 1'b1;
     if (_zy_sva_nts_151_1_pass)
      begin
       _zy_sva_hmac_null_151_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_gcm_152_reset_or)
  begin
   if (_zy_sva_null_gcm_152_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_152_1
     bit _zy_sva_nts_152_1_pass;
     _zy_sva_nts_152_1_pass = _zy_sva_b151;
     _zy_sva_null_gcm_152_ccheck = 1'b1;
     if (_zy_sva_nts_152_1_pass)
      begin
       _zy_sva_null_gcm_152_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_gcm_153_reset_or)
  begin
   if (_zy_sva_sha_gcm_153_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_153_1
     bit _zy_sva_nts_153_1_pass;
     _zy_sva_nts_153_1_pass = _zy_sva_b152;
     _zy_sva_sha_gcm_153_ccheck = 1'b1;
     if (_zy_sva_nts_153_1_pass)
      begin
       _zy_sva_sha_gcm_153_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_xts_154_reset_or)
  begin
   if (_zy_sva_null_xts_154_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_154_1
     bit _zy_sva_nts_154_1_pass;
     _zy_sva_nts_154_1_pass = _zy_sva_b153;
     _zy_sva_null_xts_154_ccheck = 1'b1;
     if (_zy_sva_nts_154_1_pass)
      begin
       _zy_sva_null_xts_154_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_xts_155_reset_or)
  begin
   if (_zy_sva_sha_xts_155_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_155_1
     bit _zy_sva_nts_155_1_pass;
     _zy_sva_nts_155_1_pass = _zy_sva_b154;
     _zy_sva_sha_xts_155_ccheck = 1'b1;
     if (_zy_sva_nts_155_1_pass)
      begin
       _zy_sva_sha_xts_155_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_null_156_reset_or)
  begin
   if (_zy_sva_null_null_156_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_156_1
     bit _zy_sva_nts_156_1_pass;
     _zy_sva_nts_156_1_pass = _zy_sva_b155;
     _zy_sva_null_null_156_ccheck = 1'b1;
     if (_zy_sva_nts_156_1_pass)
      begin
       _zy_sva_null_null_156_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_null_157_reset_or)
  begin
   if (_zy_sva_sha_null_157_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_157_1
     bit _zy_sva_nts_157_1_pass;
     _zy_sva_nts_157_1_pass = _zy_sva_b156;
     _zy_sva_sha_null_157_ccheck = 1'b1;
     if (_zy_sva_nts_157_1_pass)
      begin
       _zy_sva_sha_null_157_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_gcm_158_reset_or)
  begin
   if (_zy_sva_hmac_gcm_158_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_158_1
     bit _zy_sva_nts_158_1_pass;
     _zy_sva_nts_158_1_pass = _zy_sva_b157;
     _zy_sva_hmac_gcm_158_ccheck = 1'b1;
     if (_zy_sva_nts_158_1_pass)
      begin
       _zy_sva_hmac_gcm_158_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_xts_159_reset_or)
  begin
   if (_zy_sva_hmac_xts_159_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_159_1
     bit _zy_sva_nts_159_1_pass;
     _zy_sva_nts_159_1_pass = _zy_sva_b158;
     _zy_sva_hmac_xts_159_ccheck = 1'b1;
     if (_zy_sva_nts_159_1_pass)
      begin
       _zy_sva_hmac_xts_159_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_null_160_reset_or)
  begin
   if (_zy_sva_hmac_null_160_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_160_1
     bit _zy_sva_nts_160_1_pass;
     _zy_sva_nts_160_1_pass = _zy_sva_b159;
     _zy_sva_hmac_null_160_ccheck = 1'b1;
     if (_zy_sva_nts_160_1_pass)
      begin
       _zy_sva_hmac_null_160_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_gcm_161_reset_or)
  begin
   if (_zy_sva_null_gcm_161_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_161_1
     bit _zy_sva_nts_161_1_pass;
     _zy_sva_nts_161_1_pass = _zy_sva_b160;
     _zy_sva_null_gcm_161_ccheck = 1'b1;
     if (_zy_sva_nts_161_1_pass)
      begin
       _zy_sva_null_gcm_161_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_gcm_162_reset_or)
  begin
   if (_zy_sva_sha_gcm_162_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_162_1
     bit _zy_sva_nts_162_1_pass;
     _zy_sva_nts_162_1_pass = _zy_sva_b161;
     _zy_sva_sha_gcm_162_ccheck = 1'b1;
     if (_zy_sva_nts_162_1_pass)
      begin
       _zy_sva_sha_gcm_162_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_xts_163_reset_or)
  begin
   if (_zy_sva_null_xts_163_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_163_1
     bit _zy_sva_nts_163_1_pass;
     _zy_sva_nts_163_1_pass = _zy_sva_b162;
     _zy_sva_null_xts_163_ccheck = 1'b1;
     if (_zy_sva_nts_163_1_pass)
      begin
       _zy_sva_null_xts_163_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_xts_164_reset_or)
  begin
   if (_zy_sva_sha_xts_164_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_164_1
     bit _zy_sva_nts_164_1_pass;
     _zy_sva_nts_164_1_pass = _zy_sva_b163;
     _zy_sva_sha_xts_164_ccheck = 1'b1;
     if (_zy_sva_nts_164_1_pass)
      begin
       _zy_sva_sha_xts_164_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_null_165_reset_or)
  begin
   if (_zy_sva_null_null_165_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_165_1
     bit _zy_sva_nts_165_1_pass;
     _zy_sva_nts_165_1_pass = _zy_sva_b164;
     _zy_sva_null_null_165_ccheck = 1'b1;
     if (_zy_sva_nts_165_1_pass)
      begin
       _zy_sva_null_null_165_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_null_166_reset_or)
  begin
   if (_zy_sva_sha_null_166_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_166_1
     bit _zy_sva_nts_166_1_pass;
     _zy_sva_nts_166_1_pass = _zy_sva_b165;
     _zy_sva_sha_null_166_ccheck = 1'b1;
     if (_zy_sva_nts_166_1_pass)
      begin
       _zy_sva_sha_null_166_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_gcm_167_reset_or)
  begin
   if (_zy_sva_hmac_gcm_167_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_167_1
     bit _zy_sva_nts_167_1_pass;
     _zy_sva_nts_167_1_pass = _zy_sva_b166;
     _zy_sva_hmac_gcm_167_ccheck = 1'b1;
     if (_zy_sva_nts_167_1_pass)
      begin
       _zy_sva_hmac_gcm_167_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_xts_168_reset_or)
  begin
   if (_zy_sva_hmac_xts_168_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_168_1
     bit _zy_sva_nts_168_1_pass;
     _zy_sva_nts_168_1_pass = _zy_sva_b167;
     _zy_sva_hmac_xts_168_ccheck = 1'b1;
     if (_zy_sva_nts_168_1_pass)
      begin
       _zy_sva_hmac_xts_168_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_null_169_reset_or)
  begin
   if (_zy_sva_hmac_null_169_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_169_1
     bit _zy_sva_nts_169_1_pass;
     _zy_sva_nts_169_1_pass = _zy_sva_b168;
     _zy_sva_hmac_null_169_ccheck = 1'b1;
     if (_zy_sva_nts_169_1_pass)
      begin
       _zy_sva_hmac_null_169_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_gcm_170_reset_or)
  begin
   if (_zy_sva_null_gcm_170_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_170_1
     bit _zy_sva_nts_170_1_pass;
     _zy_sva_nts_170_1_pass = _zy_sva_b169;
     _zy_sva_null_gcm_170_ccheck = 1'b1;
     if (_zy_sva_nts_170_1_pass)
      begin
       _zy_sva_null_gcm_170_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_gcm_171_reset_or)
  begin
   if (_zy_sva_sha_gcm_171_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_171_1
     bit _zy_sva_nts_171_1_pass;
     _zy_sva_nts_171_1_pass = _zy_sva_b170;
     _zy_sva_sha_gcm_171_ccheck = 1'b1;
     if (_zy_sva_nts_171_1_pass)
      begin
       _zy_sva_sha_gcm_171_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_xts_172_reset_or)
  begin
   if (_zy_sva_null_xts_172_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_172_1
     bit _zy_sva_nts_172_1_pass;
     _zy_sva_nts_172_1_pass = _zy_sva_b171;
     _zy_sva_null_xts_172_ccheck = 1'b1;
     if (_zy_sva_nts_172_1_pass)
      begin
       _zy_sva_null_xts_172_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_xts_173_reset_or)
  begin
   if (_zy_sva_sha_xts_173_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_173_1
     bit _zy_sva_nts_173_1_pass;
     _zy_sva_nts_173_1_pass = _zy_sva_b172;
     _zy_sva_sha_xts_173_ccheck = 1'b1;
     if (_zy_sva_nts_173_1_pass)
      begin
       _zy_sva_sha_xts_173_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_null_null_174_reset_or)
  begin
   if (_zy_sva_null_null_174_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_174_1
     bit _zy_sva_nts_174_1_pass;
     _zy_sva_nts_174_1_pass = _zy_sva_b173;
     _zy_sva_null_null_174_ccheck = 1'b1;
     if (_zy_sva_nts_174_1_pass)
      begin
       _zy_sva_null_null_174_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_sha_null_175_reset_or)
  begin
   if (_zy_sva_sha_null_175_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_175_1
     bit _zy_sva_nts_175_1_pass;
     _zy_sva_nts_175_1_pass = _zy_sva_b174;
     _zy_sva_sha_null_175_ccheck = 1'b1;
     if (_zy_sva_nts_175_1_pass)
      begin
       _zy_sva_sha_null_175_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_gcm_176_reset_or)
  begin
   if (_zy_sva_hmac_gcm_176_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_176_1
     bit _zy_sva_nts_176_1_pass;
     _zy_sva_nts_176_1_pass = _zy_sva_b175;
     _zy_sva_hmac_gcm_176_ccheck = 1'b1;
     if (_zy_sva_nts_176_1_pass)
      begin
       _zy_sva_hmac_gcm_176_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_xts_177_reset_or)
  begin
   if (_zy_sva_hmac_xts_177_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_177_1
     bit _zy_sva_nts_177_1_pass;
     _zy_sva_nts_177_1_pass = _zy_sva_b176;
     _zy_sva_hmac_xts_177_ccheck = 1'b1;
     if (_zy_sva_nts_177_1_pass)
      begin
       _zy_sva_hmac_xts_177_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or posedge _zy_sva_hmac_null_178_reset_or)
  begin
   if (_zy_sva_hmac_null_178_reset_or)
    begin
    end
   else
    begin:_zy_sva_sblk_178_1
     bit _zy_sva_nts_178_1_pass;
     _zy_sva_nts_178_1_pass = _zy_sva_b177;
     _zy_sva_hmac_null_178_ccheck = 1'b1;
     if (_zy_sva_nts_178_1_pass)
      begin
       _zy_sva_hmac_null_178_cpass = 1'b1;
      end
    end
  end
always 
 @(posedge clk or negedge rst_n)
  begin
   if (( !rst_n ))
    begin
     tlv_counter <= 5'b0;
    end
   else
    if (stitcher_rd)
     begin
      if (stitcher_eot)
       begin
        tlv_counter <= 5'b0;
       end
      else
       begin
        tlv_counter <= (tlv_counter + 5'b01);
       end
     end
  end
always 
 @(posedge clk or negedge rst_n)
  begin
   if (( !rst_n ))
    begin
     tlv_type <= RQE;
     aux_key_type <= NO_AUX_KEY;
     aux_iv_op <= IV_SRC;
     aux_cipher_op <= CPH_NULL;
     aux_auth_op <= AUTH_NULL;
     aux_raw_auth_op <= AUTH_NULL;
     kme_internal_word0 <= 64'b0;
     kme_internal_dek_kim_word <= 64'b0;
     kme_internal_dak_kim_word <= 64'b0;
     debug_cmd <= 32'b0;
     aux_key_header <= 32'b0;
     skip <= 7'b0;
     guid0 <= 64'b0;
     guid1 <= 64'b0;
     guid2 <= 64'b0;
     guid3 <= 64'b0;
     iv0 <= 64'b0;
     iv1 <= 64'b0;
     buffer <= 32'b0;
     fifo_in.id <= KME_WORD0;
    end
   else
    begin
     tlv_type <= nxt_tlv_type;
     aux_key_type <= nxt_aux_key_type;
     aux_iv_op <= nxt_aux_iv_op;
     aux_cipher_op <= nxt_aux_cipher_op;
     aux_auth_op <= nxt_aux_auth_op;
     aux_raw_auth_op <= nxt_aux_raw_auth_op;
     kme_internal_word0 <= nxt_kme_internal_word0;
     kme_internal_dek_kim_word <= nxt_kme_internal_dek_kim_word;
     kme_internal_dak_kim_word <= nxt_kme_internal_dak_kim_word;
     debug_cmd <= nxt_debug_cmd;
     aux_key_header <= nxt_aux_key_header;
     skip <= nxt_skip;
     guid0 <= nxt_guid0;
     guid1 <= nxt_guid1;
     guid2 <= nxt_guid2;
     guid3 <= nxt_guid3;
     iv0 <= nxt_iv0;
     iv1 <= nxt_iv1;
     buffer <= nxt_buffer;
     fifo_in.id <= nxt_fifo_in_id;
    end
  end
always 
 @(*)
  begin
   fifo_in.tdata = 64'b0;
   fifo_in_valid = 1'b0;
   nxt_tlv_type = tlv_type;
   nxt_aux_key_type = aux_key_type;
   nxt_aux_iv_op = aux_iv_op;
   nxt_aux_cipher_op = aux_cipher_op;
   nxt_aux_auth_op = aux_auth_op;
   nxt_aux_raw_auth_op = aux_raw_auth_op;
   nxt_kme_internal_word0 = kme_internal_word0;
   nxt_kme_internal_dek_kim_word = kme_internal_dek_kim_word;
   nxt_kme_internal_dak_kim_word = kme_internal_dak_kim_word;
   nxt_aux_key_header = aux_key_header;
   nxt_debug_cmd = debug_cmd;
   nxt_skip = skip;
   nxt_guid0 = guid0;
   nxt_guid1 = guid1;
   nxt_guid2 = guid2;
   nxt_guid3 = guid3;
   nxt_iv0 = iv0;
   nxt_iv1 = iv1;
   nxt_buffer = buffer;
   tlv_word0 = stitcher_out.tdata;
   tlv_word1 = stitcher_out.tdata;
   tlv_word2 = stitcher_out.tdata;
   frame_word = stitcher_out.tdata;
   stitcher_rd = ((( ~stitcher_empty ) & ( ~fifo_in_stall )) & ( ~skip.start ));
   if (( !fifo_in_stall ))
    begin
     if (skip.start)
      begin
       if ((fifo_in.id == skip.till))
        begin
         nxt_skip.start = 1'b0;
        end
       else
        begin
         fifo_in_valid = 1'b1;
        end
       if (skip.partial)
        begin
         nxt_skip.partial = 1'b0;
         nxt_skip.endian_swap = 1'b0;
         begin:_zypbctfiCscp13_L234_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {32'b0,buffer};
          _zyL234_tfiRv52 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
         end
         fifo_in.tdata = (skip.endian_swap ? _zyL234_tfiRv52 : {buffer,32'b0});
        end
       case (int_tlv_counter)
        6'b010:
         fifo_in.tdata = guid0;
        6'b011:
         fifo_in.tdata = guid1;
        6'b0100:
         fifo_in.tdata = guid2;
        6'b0101:
         fifo_in.tdata = guid3;
        6'b0110:
         fifo_in.tdata = iv0;
        6'b0111:
         fifo_in.tdata = iv1;
        6'b01000:
         fifo_in.tdata = kme_internal_dek_kim_word;
        6'b01001:
         fifo_in.tdata = kme_internal_dak_kim_word;
       endcase
       if ((int_tlv_counter == IDX_KME_IVTWEAK))
        begin
         begin:_zypbctfiCscp14_L252_validate_dek
          reg _zyoff_L753_tfiV2;
          aux_key_type_e _zykey_type_L754_tfiV3;
          cmd_cipher_op_e _zycipher_op_L755_tfiV4;
          aux_kdf_mode_e _zykdf_mode_L756_tfiV5;
          reg _zyL768_tfiRv7;
          reg _zyL768_tfiRv8;
          reg _zyL769_tfiRv9;
          reg _zyL769_tfiRv10;
          _zyoff_L753_tfiV2 = always_validate_kim_ref;
          _zykey_type_L754_tfiV3 = aux_key_type;
          _zycipher_op_L755_tfiV4 = aux_cipher_op;
          _zykdf_mode_L756_tfiV5 = aux_key_header.kdf_mode;
          _zyL252_tfiRv53 = 1'b1;
          if (( !_zyoff_L753_tfiV2 ))
          begin
          case (_zykey_type_L754_tfiV3)
          NO_AUX_KEY:
          _zyL252_tfiRv53 = 1'b0;
          AUX_KEY_ONLY:
          begin
          begin:_zypbctfiCscp0_L768_is_keyless_cipher
          cmd_cipher_op_e _zycipher_op_L845_tfiV11;
          _zycipher_op_L845_tfiV11 = _zycipher_op_L755_tfiV4;
          _zyL768_tfiRv7 = ( ~(((_zycipher_op_L845_tfiV11 == AES_GCM) | (_zycipher_op_L845_tfiV11 == AES_XTS_XEX)) | (_zycipher_op_L845_tfiV11 == AES_GMAC)) );
          end
          begin:_zypbctfiCscp1_L768_is_kdf_non_combo
          aux_kdf_mode_e _zykdf_mode_L862_tfiV13;
          _zykdf_mode_L862_tfiV13 = _zykdf_mode_L756_tfiV5;
          _zyL768_tfiRv8 = ((_zykdf_mode_L862_tfiV13 == KDF_MODE_GUID) | (_zykdf_mode_L862_tfiV13 == KDF_MODE_RGUID));
          end
          if ((_zyL768_tfiRv7 & _zyL768_tfiRv8))
          _zyL252_tfiRv53 = 1'b0;
          end
          ENC_DAK:
          begin
          begin:_zypbctfiCscp2_L769_is_keyless_cipher
          cmd_cipher_op_e _zycipher_op_L845_tfiV11;
          _zycipher_op_L845_tfiV11 = _zycipher_op_L755_tfiV4;
          _zyL769_tfiRv9 = ( ~(((_zycipher_op_L845_tfiV11 == AES_GCM) | (_zycipher_op_L845_tfiV11 == AES_XTS_XEX)) | (_zycipher_op_L845_tfiV11 == AES_GMAC)) );
          end
          begin:_zypbctfiCscp3_L769_is_kdf_non_combo
          aux_kdf_mode_e _zykdf_mode_L862_tfiV13;
          _zykdf_mode_L862_tfiV13 = _zykdf_mode_L756_tfiV5;
          _zyL769_tfiRv10 = ((_zykdf_mode_L862_tfiV13 == KDF_MODE_GUID) | (_zykdf_mode_L862_tfiV13 == KDF_MODE_RGUID));
          end
          if ((_zyL769_tfiRv9 & _zyL769_tfiRv10))
          _zyL252_tfiRv53 = 1'b0;
          end
          endcase
          end
         end
         nxt_kme_internal_dek_kim_word.validate_dek = _zyL252_tfiRv53;
         begin:_zypbctfiCscp15_L253_missing_guid
          tlv_types_e _zyl_tlv_type_L725_tfiV15;
          aux_kdf_mode_e _zykdf_mode_L726_tfiV16;
          aux_key_op_e _zydek_key_op_L727_tfiV17, _zydak_key_op_L728_tfiV18;
          _zyl_tlv_type_L725_tfiV15 = tlv_type;
          _zykdf_mode_L726_tfiV16 = aux_key_header.kdf_mode;
          _zydek_key_op_L727_tfiV17 = aux_key_header.dek_key_op;
          _zydak_key_op_L728_tfiV18 = aux_key_header.dak_key_op;
          _zyL253_tfiRv54 = ((((_zyl_tlv_type_L725_tfiV15 == AUX_CMD) || (_zyl_tlv_type_L725_tfiV15 == AUX_CMD_IV)) && ((_zydek_key_op_L727_tfiV17 == KDF) || (_zydak_key_op_L728_tfiV18 == KDF))) && ((_zykdf_mode_L726_tfiV16 == KDF_MODE_GUID) || (_zykdf_mode_L726_tfiV16 == KDF_MODE_COMB_GUID)));
         end
         nxt_kme_internal_dek_kim_word.missing_guid = _zyL253_tfiRv54;
         begin:_zypbctfiCscp16_L254_missing_iv
          tlv_types_e _zyl_tlv_type_L740_tfiV20;
          cmd_iv_op_e _zyiv_op_L741_tfiV21;
          cmd_cipher_op_e _zycipher_op_L742_tfiV22;
          reg _zyL746_tfiRv24;
          _zyl_tlv_type_L740_tfiV20 = tlv_type;
          _zyiv_op_L741_tfiV21 = aux_iv_op;
          _zycipher_op_L742_tfiV22 = aux_cipher_op;
          begin:_zypbctfiCscp4_L746_is_keyless_cipher
          cmd_cipher_op_e _zycipher_op_L845_tfiV11;
          _zycipher_op_L845_tfiV11 = _zycipher_op_L742_tfiV22;
          _zyL746_tfiRv24 = ( ~(((_zycipher_op_L845_tfiV11 == AES_GCM) | (_zycipher_op_L845_tfiV11 == AES_XTS_XEX)) | (_zycipher_op_L845_tfiV11 == AES_GMAC)) );
          end
          _zyL254_tfiRv55 = ((((_zyl_tlv_type_L740_tfiV20 == AUX_CMD) || (_zyl_tlv_type_L740_tfiV20 == AUX_CMD_GUID)) && (_zyiv_op_L741_tfiV21 == IV_INC)) && ( ~_zyL746_tfiRv24 ));
         end
         nxt_kme_internal_dek_kim_word.missing_iv = _zyL254_tfiRv55;
         begin:_zypbctfiCscp17_L255_validate_dak
          reg _zyoff_L777_tfiV25;
          aux_key_type_e _zykey_type_L778_tfiV26;
          cmd_auth_op_e _zyauth_op_L779_tfiV27, _zyraw_auth_op_L780_tfiV28;
          reg _zyL792_tfiRv30;
          reg _zyL793_tfiRv31;
          reg _zyL794_tfiRv32;
          _zyoff_L777_tfiV25 = always_validate_kim_ref;
          _zykey_type_L778_tfiV26 = aux_key_type;
          _zyauth_op_L779_tfiV27 = aux_auth_op;
          _zyraw_auth_op_L780_tfiV28 = aux_raw_auth_op;
          _zyL255_tfiRv56 = 1'b1;
          if (( !_zyoff_L777_tfiV25 ))
          begin
          case (_zykey_type_L778_tfiV26)
          NO_AUX_KEY:
          _zyL255_tfiRv56 = 1'b0;
          AUX_KEY_ONLY:
          begin
          begin:_zypbctfiCscp5_L792_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = _zyauth_op_L779_tfiV27;
          _zyraw_auth_op_L854_tfiV34 = _zyraw_auth_op_L780_tfiV28;
          _zyL792_tfiRv30 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          if (_zyL792_tfiRv30)
          _zyL255_tfiRv56 = 1'b0;
          end
          ENC_DEK256:
          begin
          begin:_zypbctfiCscp6_L793_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = _zyauth_op_L779_tfiV27;
          _zyraw_auth_op_L854_tfiV34 = _zyraw_auth_op_L780_tfiV28;
          _zyL793_tfiRv31 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          if (_zyL793_tfiRv31)
          _zyL255_tfiRv56 = 1'b0;
          end
          ENC_DEK512:
          begin
          begin:_zypbctfiCscp7_L794_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = _zyauth_op_L779_tfiV27;
          _zyraw_auth_op_L854_tfiV34 = _zyraw_auth_op_L780_tfiV28;
          _zyL794_tfiRv32 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          if (_zyL794_tfiRv32)
          _zyL255_tfiRv56 = 1'b0;
          end
          endcase
          end
         end
         nxt_kme_internal_dak_kim_word.validate_dak = _zyL255_tfiRv56;
        end
      end
    end
   if (stitcher_rd)
    begin
     if (key_blob_region)
      begin
       case (aux_key_type)
        DEK256,
        DEK512,
        DAK:
         begin
          fifo_in_valid = 1'b1;
          begin:_zypbctfiCscp18_L288_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL288_tfiRv57 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL288_tfiRv57;
          nxt_buffer = stitcher_out.tdata[63:32];
          if (stitcher_eot)
          begin
          begin:_zypbctfiCscp19_L293_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL293_tfiRv58 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL293_tfiRv58;
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_WORD0;
          end
         end
        DEK256_DAK,
        DEK512_DAK:
         begin
          fifo_in_valid = 1'b1;
          begin:_zypbctfiCscp20_L301_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL301_tfiRv59 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL301_tfiRv59;
          nxt_buffer = stitcher_out.tdata[63:32];
          if ((int_tlv_counter == 32'b011111))
          begin
          begin:_zypbctfiCscp21_L306_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL306_tfiRv60 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL306_tfiRv60;
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_DAK;
          end
          if (stitcher_eot)
          begin
          begin:_zypbctfiCscp22_L313_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL313_tfiRv61 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL313_tfiRv61;
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_WORD0;
          end
         end
        ENC_DEK256,
        ENC_DEK512,
        ENC_DAK:
         begin
          fifo_in_valid = 1'b1;
          begin:_zypbctfiCscp23_L321_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL321_tfiRv62 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL321_tfiRv62;
          nxt_buffer = stitcher_out.tdata[63:32];
          if ((int_tlv_counter == IDX_KME_EIV))
          begin
          begin:_zypbctfiCscp24_L327_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL327_tfiRv63 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL327_tfiRv63;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          nxt_skip.endian_swap = 1'b1;
          nxt_skip.till = ((aux_key_type == ENC_DEK256) ? KME_DEK1 : KME_DEK0);
          end
          if ((int_tlv_counter == IDX_KME_AIV))
          begin
          begin:_zypbctfiCscp25_L337_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL337_tfiRv64 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL337_tfiRv64;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          nxt_skip.endian_swap = 1'b1;
          nxt_skip.till = KME_DAK;
          end
          if (stitcher_eot)
          begin
          begin:_zypbctfiCscp26_L346_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {32'b0,stitcher_out.tdata[32'sd31:32'sd0]};
          _zyL346_tfiRv65 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL346_tfiRv65;
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_WORD0;
          end
         end
        ENC_DEK256_DAK,
        ENC_DEK512_DAK:
         begin
          fifo_in_valid = 1'b1;
          begin:_zypbctfiCscp27_L354_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL354_tfiRv66 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL354_tfiRv66;
          nxt_buffer = stitcher_out.tdata[63:32];
          if ((int_tlv_counter == IDX_KME_EIV))
          begin
          begin:_zypbctfiCscp28_L359_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL359_tfiRv67 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL359_tfiRv67;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          nxt_skip.endian_swap = 1'b1;
          nxt_skip.till = ((aux_key_type == ENC_DEK256_DAK) ? KME_DEK1 : KME_DEK0);
          end
          if ((int_tlv_counter == 32'b0100001))
          begin
          begin:_zypbctfiCscp29_L368_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {32'b0,stitcher_out.tdata[32'sd31:32'sd0]};
          _zyL368_tfiRv68 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL368_tfiRv68;
          end
          if ((int_tlv_counter == IDX_KME_AIV))
          begin
          begin:_zypbctfiCscp30_L373_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL373_tfiRv69 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL373_tfiRv69;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          nxt_skip.endian_swap = 1'b1;
          nxt_skip.till = KME_DAK;
          end
          if (stitcher_eot)
          begin
          begin:_zypbctfiCscp31_L382_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {32'b0,stitcher_out.tdata[32'sd31:32'sd0]};
          _zyL382_tfiRv70 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL382_tfiRv70;
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_WORD0;
          end
         end
        ENC_DEK256_DAK_COMB,
        ENC_DEK512_DAK_COMB:
         begin
          fifo_in_valid = 1'b1;
          begin:_zypbctfiCscp32_L390_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL390_tfiRv71 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL390_tfiRv71;
          nxt_buffer = stitcher_out.tdata[63:32];
          if ((int_tlv_counter == IDX_KME_EIV))
          begin
          begin:_zypbctfiCscp33_L395_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {stitcher_out.tdata[32'sd31:32'sd0],buffer};
          _zyL395_tfiRv72 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL395_tfiRv72;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          nxt_skip.endian_swap = 1'b1;
          nxt_skip.till = ((aux_key_type == ENC_DEK256_DAK_COMB) ? KME_DEK1 : KME_DEK0);
          end
          if ((int_tlv_counter == 32'b011111))
          begin
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_DAK;
          end
          if (stitcher_eot)
          begin
          begin:_zypbctfiCscp34_L410_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = {32'b0,stitcher_out.tdata[32'sd31:32'sd0]};
          _zyL410_tfiRv73 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          fifo_in.tdata = _zyL410_tfiRv73;
          nxt_skip.start = 1'b1;
          nxt_skip.till = KME_WORD0;
          end
         end
       endcase
      end
     else
      begin
       case (tlv_counter)
        5'b0:
         begin
          nxt_kme_internal_word0 = 64'b0;
          nxt_kme_internal_word0.tlv_type = tlv_word0.tlv_type;
          nxt_kme_internal_word0.tlv_eng_id = tlv_word0.tlv_eng_id;
          nxt_kme_internal_word0.tlv_seq_num = tlv_word0.tlv_seq_num;
          nxt_kme_internal_word0.tlv_frame_num = tlv_word0.tlv_frame_num;
          nxt_tlv_type = tlv_word0.tlv_type;
          if ((tlv_word0.tlv_type == RQE))
          begin
          nxt_kme_internal_dek_kim_word = 64'b0;
          nxt_kme_internal_dak_kim_word = 64'b0;
          nxt_kme_internal_dek_kim_word.vf_valid = tlv_word0.vf_valid;
          nxt_kme_internal_dak_kim_word.vf_valid = tlv_word0.vf_valid;
          end
          nxt_aux_key_type = NO_AUX_KEY;
          nxt_aux_iv_op = IV_SRC;
          nxt_aux_cipher_op = CPH_NULL;
          nxt_aux_auth_op = AUTH_NULL;
          nxt_aux_raw_auth_op = AUTH_NULL;
          nxt_aux_key_header = 32'b0;
          nxt_iv0 = 64'b0;
          nxt_iv1 = 64'b0;
          nxt_guid0 = 64'b0;
          nxt_guid1 = 64'b0;
          nxt_guid2 = 64'b0;
          nxt_guid3 = 64'b0;
         end
        5'b01:
         begin
          if ((tlv_type == RQE))
          begin
          nxt_kme_internal_dek_kim_word.pf_num = tlv_word1.pf_number;
          nxt_kme_internal_dek_kim_word.vf_num = tlv_word1.vf_number;
          nxt_kme_internal_dak_kim_word.pf_num = tlv_word1.pf_number;
          nxt_kme_internal_dak_kim_word.vf_num = tlv_word1.vf_number;
          end
          else
          begin
          case (tlv_type)
          AUX_CMD:
          if ((frame_word.src_guid_present == GUID_PRESENT))
          nxt_tlv_type = AUX_CMD_GUID;
          AUX_CMD_IV:
          if ((frame_word.src_guid_present == GUID_PRESENT))
          nxt_tlv_type = AUX_CMD_GUID_IV;
          endcase
          if (disable_debug_cmd_q)
          begin
          nxt_debug_cmd = 32'b0;
          end
          else
          begin
          nxt_debug_cmd = stitcher_out.tdata[63:32];
          end
          end
         end
        5'b010:
         begin
          nxt_kme_internal_word0.key_type = tlv_word2.key_type;
          begin:_zypbctfiCscp35_L485_needs_dek
          reg _zyoff_L802_tfiV36;
          aux_key_type_e _zykey_type_L803_tfiV37;
          cmd_cipher_op_e _zycipher_op_L804_tfiV38;
          reg _zyL814_tfiRv40;
          reg _zyL815_tfiRv41;
          _zyoff_L802_tfiV36 = always_validate_kim_ref;
          _zykey_type_L803_tfiV37 = tlv_word2.key_type;
          _zycipher_op_L804_tfiV38 = tlv_word2.cipher_op;
          _zyL485_tfiRv74 = 1'b1;
          if (( !_zyoff_L802_tfiV36 ))
          begin
          case (_zykey_type_L803_tfiV37)
          NO_AUX_KEY:
          _zyL485_tfiRv74 = 1'b0;
          AUX_KEY_ONLY:
          begin
          begin:_zypbctfiCscp8_L814_is_keyless_cipher
          cmd_cipher_op_e _zycipher_op_L845_tfiV11;
          _zycipher_op_L845_tfiV11 = _zycipher_op_L804_tfiV38;
          _zyL814_tfiRv40 = ( ~(((_zycipher_op_L845_tfiV11 == AES_GCM) | (_zycipher_op_L845_tfiV11 == AES_XTS_XEX)) | (_zycipher_op_L845_tfiV11 == AES_GMAC)) );
          end
          if (_zyL814_tfiRv40)
          _zyL485_tfiRv74 = 1'b0;
          end
          ENC_DAK:
          begin
          begin:_zypbctfiCscp9_L815_is_keyless_cipher
          cmd_cipher_op_e _zycipher_op_L845_tfiV11;
          _zycipher_op_L845_tfiV11 = _zycipher_op_L804_tfiV38;
          _zyL815_tfiRv41 = ( ~(((_zycipher_op_L845_tfiV11 == AES_GCM) | (_zycipher_op_L845_tfiV11 == AES_XTS_XEX)) | (_zycipher_op_L845_tfiV11 == AES_GMAC)) );
          end
          if (_zyL815_tfiRv41)
          _zyL485_tfiRv74 = 1'b0;
          end
          endcase
          end
          end
          nxt_kme_internal_word0.needs_dek = _zyL485_tfiRv74;
          begin:_zypbctfiCscp36_L486_needs_dak
          reg _zyoff_L823_tfiV42;
          aux_key_type_e _zykey_type_L824_tfiV43;
          cmd_auth_op_e _zyauth_op_L825_tfiV44, _zyraw_auth_op_L826_tfiV45;
          reg _zyL836_tfiRv47;
          reg _zyL837_tfiRv48;
          reg _zyL838_tfiRv49;
          _zyoff_L823_tfiV42 = always_validate_kim_ref;
          _zykey_type_L824_tfiV43 = tlv_word2.key_type;
          _zyauth_op_L825_tfiV44 = tlv_word2.auth_op;
          _zyraw_auth_op_L826_tfiV45 = tlv_word2.raw_auth_op;
          _zyL486_tfiRv75 = 1'b1;
          if (( !_zyoff_L823_tfiV42 ))
          begin
          case (_zykey_type_L824_tfiV43)
          NO_AUX_KEY:
          _zyL486_tfiRv75 = 1'b0;
          AUX_KEY_ONLY:
          begin
          begin:_zypbctfiCscp10_L836_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = _zyauth_op_L825_tfiV44;
          _zyraw_auth_op_L854_tfiV34 = _zyraw_auth_op_L826_tfiV45;
          _zyL836_tfiRv47 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          if (_zyL836_tfiRv47)
          _zyL486_tfiRv75 = 1'b0;
          end
          ENC_DEK256:
          begin
          begin:_zypbctfiCscp11_L837_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = _zyauth_op_L825_tfiV44;
          _zyraw_auth_op_L854_tfiV34 = _zyraw_auth_op_L826_tfiV45;
          _zyL837_tfiRv48 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          if (_zyL837_tfiRv48)
          _zyL486_tfiRv75 = 1'b0;
          end
          ENC_DEK512:
          begin
          begin:_zypbctfiCscp12_L838_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = _zyauth_op_L825_tfiV44;
          _zyraw_auth_op_L854_tfiV34 = _zyraw_auth_op_L826_tfiV45;
          _zyL838_tfiRv49 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          if (_zyL838_tfiRv49)
          _zyL486_tfiRv75 = 1'b0;
          end
          endcase
          end
          end
          nxt_kme_internal_word0.needs_dak = _zyL486_tfiRv75;
          begin:_zypbctfiCscp37_L489_is_keyless_cipher
          cmd_cipher_op_e _zycipher_op_L845_tfiV11;
          _zycipher_op_L845_tfiV11 = tlv_word2.cipher_op;
          _zyL489_tfiRv76 = ( ~(((_zycipher_op_L845_tfiV11 == AES_GCM) | (_zycipher_op_L845_tfiV11 == AES_XTS_XEX)) | (_zycipher_op_L845_tfiV11 == AES_GMAC)) );
          end
          begin:_zypbctfiCscp38_L489_is_keyless_hash
          cmd_auth_op_e _zyauth_op_L853_tfiV33, _zyraw_auth_op_L854_tfiV34;
          _zyauth_op_L853_tfiV33 = tlv_word2.auth_op;
          _zyraw_auth_op_L854_tfiV34 = tlv_word2.raw_auth_op;
          _zyL489_tfiRv77 = ((_zyauth_op_L853_tfiV33 != HMAC_SHA2) & (_zyraw_auth_op_L854_tfiV34 != HMAC_SHA2));
          end
          nxt_kme_internal_word0.keyless_algos = (_zyL489_tfiRv76 & _zyL489_tfiRv77);
          begin:_zypbctfiCscp39_L492_kdf_dek_iter_f
          cmd_cipher_op_e _zycipher_op_L871_tfiV50;
          _zycipher_op_L871_tfiV50 = tlv_word2.cipher_op;
          _zyL492_tfiRv78 = ((_zycipher_op_L871_tfiV50 == AES_XTS_XEX) ? 1'b1 : 1'b0);
          end
          nxt_kme_internal_word0.kdf_dek_iter = _zyL492_tfiRv78;
          nxt_aux_key_type = tlv_word2.key_type;
          nxt_aux_iv_op = tlv_word2.iv_op;
          nxt_aux_cipher_op = tlv_word2.cipher_op;
          nxt_aux_auth_op = tlv_word2.auth_op;
          nxt_aux_raw_auth_op = tlv_word2.raw_auth_op;
          fifo_in_valid = 1'b1;
          fifo_in.tdata = nxt_kme_internal_word0;
          if (stitcher_eot)
          begin
          nxt_buffer = debug_cmd;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          end
         end
        5'b011:
         begin
          case (tlv_type)
          AUX_CMD_GUID:
          begin
          begin:_zypbctfiCscp40_L526_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL526_tfiRv79 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid0 = _zyL526_tfiRv79;
          end
          AUX_CMD_GUID_IV:
          begin
          begin:_zypbctfiCscp41_L527_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL527_tfiRv80 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid0 = _zyL527_tfiRv80;
          end
          AUX_CMD_IV:
          nxt_iv0 = stitcher_out.tdata;
          endcase
          if ((tlv_type == AUX_CMD))
          begin
          {nxt_buffer,nxt_aux_key_header} = stitcher_out.tdata;
          fifo_in_valid = 1'b1;
          fifo_in.tdata = {debug_cmd,nxt_aux_key_header};
          nxt_skip.start = 1'b1;
          end
         end
        5'b0100:
         begin
          case (tlv_type)
          AUX_CMD_GUID:
          begin
          begin:_zypbctfiCscp42_L541_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL541_tfiRv81 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid1 = _zyL541_tfiRv81;
          end
          AUX_CMD_GUID_IV:
          begin
          begin:_zypbctfiCscp43_L542_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL542_tfiRv82 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid1 = _zyL542_tfiRv82;
          end
          AUX_CMD_IV:
          nxt_iv1 = stitcher_out.tdata;
          endcase
          if (stitcher_eot)
          begin
          nxt_buffer = debug_cmd;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          end
         end
        5'b0101:
         begin
          case (tlv_type)
          AUX_CMD_GUID:
          begin
          begin:_zypbctfiCscp44_L555_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL555_tfiRv83 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid2 = _zyL555_tfiRv83;
          end
          AUX_CMD_GUID_IV:
          begin
          begin:_zypbctfiCscp45_L556_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL556_tfiRv84 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid2 = _zyL556_tfiRv84;
          end
          endcase
          if ((tlv_type == AUX_CMD_IV))
          begin
          {nxt_buffer,nxt_aux_key_header} = stitcher_out.tdata;
          fifo_in_valid = 1'b1;
          fifo_in.tdata = {debug_cmd,nxt_aux_key_header};
          nxt_skip.start = 1'b1;
          end
         end
        5'b0110:
         begin
          case (tlv_type)
          AUX_CMD_GUID:
          begin
          begin:_zypbctfiCscp46_L569_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL569_tfiRv85 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid3 = _zyL569_tfiRv85;
          end
          AUX_CMD_GUID_IV:
          begin
          begin:_zypbctfiCscp47_L570_endian_switch
          reg [63:0] _zydata_L20_tfiV0 ;
          _zydata_L20_tfiV0 = stitcher_out.tdata;
          _zyL570_tfiRv86 = {_zydata_L20_tfiV0[32'sd7:32'sd0],_zydata_L20_tfiV0[32'sd15:32'sd8],_zydata_L20_tfiV0[32'sd23:32'sd16],_zydata_L20_tfiV0[32'sd31:32'sd24],_zydata_L20_tfiV0[32'sd39:32'sd32],_zydata_L20_tfiV0[32'sd47:32'sd40],_zydata_L20_tfiV0[32'sd55:32'sd48],_zydata_L20_tfiV0[32'sd63:32'sd56]};
          end
          nxt_guid3 = _zyL570_tfiRv86;
          end
          endcase
          if (stitcher_eot)
          begin
          nxt_buffer = debug_cmd;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          end
         end
        5'b0111:
         begin
          case (tlv_type)
          AUX_CMD_GUID_IV:
          nxt_iv0 = stitcher_out.tdata;
          endcase
          if ((tlv_type == AUX_CMD_GUID))
          begin
          {nxt_buffer,nxt_aux_key_header} = stitcher_out.tdata;
          fifo_in_valid = 1'b1;
          fifo_in.tdata = {debug_cmd,nxt_aux_key_header};
          nxt_skip.start = 1'b1;
          end
         end
        5'b01000:
         begin
          case (tlv_type)
          AUX_CMD_GUID_IV:
          nxt_iv1 = stitcher_out.tdata;
          endcase
          if (stitcher_eot)
          begin
          nxt_buffer = debug_cmd;
          nxt_skip.start = 1'b1;
          nxt_skip.partial = 1'b1;
          end
         end
        5'b01001:
         begin
          {nxt_buffer,nxt_aux_key_header} = stitcher_out.tdata;
          fifo_in_valid = 1'b1;
          fifo_in.tdata = {debug_cmd,nxt_aux_key_header};
          nxt_skip.start = 1'b1;
         end
       endcase
       case (aux_key_type)
        NO_AUX_KEY:
         nxt_skip.till = KME_WORD0;
        AUX_KEY_ONLY:
         nxt_skip.till = KME_WORD0;
        DEK256:
         nxt_skip.till = KME_DEK1;
        DEK512:
         nxt_skip.till = KME_DEK0;
        DAK:
         nxt_skip.till = KME_DAK;
        DEK256_DAK:
         nxt_skip.till = KME_DEK1;
        DEK512_DAK:
         nxt_skip.till = KME_DEK0;
        ENC_DEK256:
         nxt_skip.till = KME_EIV;
        ENC_DEK512:
         nxt_skip.till = KME_EIV;
        ENC_DAK:
         nxt_skip.till = KME_AIV;
        ENC_DEK256_DAK:
         nxt_skip.till = KME_EIV;
        ENC_DEK512_DAK:
         nxt_skip.till = KME_EIV;
        ENC_DEK256_DAK_COMB:
         nxt_skip.till = KME_EIV;
        ENC_DEK512_DAK_COMB:
         nxt_skip.till = KME_EIV;
       endcase
      end
    end
  end
always 
 @(posedge clk or negedge rst_n)
  begin
   if (( !rst_n ))
    begin
     fifo_in.eot <= 1'b0;
     key_blob_region <= 1'b0;
     int_tlv_counter <= 6'b0;
    end
   else
    if (fifo_in_valid)
     begin
      case (int_tlv_counter)
       6'b101001:
        fifo_in.eot <= 1'b1;
       6'b101010:
        fifo_in.eot <= 1'b0;
       default:
        fifo_in.eot <= fifo_in.eot;
      endcase
      case (int_tlv_counter)
       6'b010101:
        key_blob_region <= 1'b1;
       6'b101010:
        key_blob_region <= 1'b0;
       default:
        key_blob_region <= key_blob_region;
      endcase
      case (int_tlv_counter)
       6'b101010:
        int_tlv_counter <= 6'b0;
       default:
        int_tlv_counter <= (int_tlv_counter + 6'b01);
      endcase
     end
  end
always 
 @(*)
  begin
   nxt_fifo_in_id = fifo_in.id;
   fifo_in.sot = (fifo_in_valid & (fifo_in.id == KME_WORD0));
   fifo_in.eoi = 1'b0;
   if (fifo_in_valid)
    begin
     case (int_tlv_counter)
      6'b0:
       begin
        nxt_fifo_in_id = KME_DEBUG_KEYHDR;
        fifo_in.eoi = 1'b1;
       end
      6'b01:
       begin
        nxt_fifo_in_id = KME_GUID;
        fifo_in.eoi = 1'b1;
       end
      6'b0101:
       begin
        nxt_fifo_in_id = KME_IVTWEAK;
        fifo_in.eoi = 1'b1;
       end
      6'b0111:
       begin
        nxt_fifo_in_id = KME_KIM;
        fifo_in.eoi = 1'b1;
       end
      6'b01001:
       begin
        nxt_fifo_in_id = KME_DEK_CKV0;
        fifo_in.eoi = 1'b1;
       end
      6'b01101:
       begin
        nxt_fifo_in_id = KME_DEK_CKV1;
        fifo_in.eoi = 1'b1;
       end
      6'b010001:
       begin
        nxt_fifo_in_id = KME_DAK_CKV;
        fifo_in.eoi = 1'b1;
       end
      6'b010101:
       begin
        nxt_fifo_in_id = KME_EIV;
        fifo_in.eoi = 1'b1;
       end
      6'b010111:
       begin
        nxt_fifo_in_id = KME_DEK0;
        fifo_in.eoi = 1'b1;
       end
      6'b011011:
       begin
        nxt_fifo_in_id = KME_DEK1;
        fifo_in.eoi = 1'b1;
       end
      6'b011111:
       begin
        nxt_fifo_in_id = KME_ETAG;
        fifo_in.eoi = 1'b1;
       end
      6'b100001:
       begin
        nxt_fifo_in_id = KME_AIV;
        fifo_in.eoi = 1'b1;
       end
      6'b100011:
       begin
        nxt_fifo_in_id = KME_DAK;
        fifo_in.eoi = 1'b1;
       end
      6'b100111:
       begin
        nxt_fifo_in_id = KME_ATAG;
        fifo_in.eoi = 1'b1;
       end
      6'b101001:
       begin
        nxt_fifo_in_id = KME_ERROR;
        fifo_in.eoi = 1'b1;
       end
      IDX_KME_ERROR:
       begin
        nxt_fifo_in_id = KME_WORD0;
        fifo_in.eoi = 1'b1;
       end
     endcase
    end
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[0]"
//pragma RTLNAME "key_type[0]" "key_type_0_"
if(1) begin: key_type_0_
 localparam integer jj = 0;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_39_cpass,,_zy_sva_brcm_aux_cmd_39_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_40_cpass,,_zy_sva_brcm_aux_cmd_iv_40_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_41_cpass,,_zy_sva_brcm_aux_cmd_guid_41_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_42_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_42_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_43_cpass,,_zy_sva_brcm_key_type_43_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[1]"
//pragma RTLNAME "key_type[1]" "key_type_1_"
if(1) begin: key_type_1_
 localparam integer jj = 1;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_44_cpass,,_zy_sva_brcm_aux_cmd_44_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_45_cpass,,_zy_sva_brcm_aux_cmd_iv_45_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_46_cpass,,_zy_sva_brcm_aux_cmd_guid_46_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_47_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_47_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_48_cpass,,_zy_sva_brcm_key_type_48_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[2]"
//pragma RTLNAME "key_type[2]" "key_type_2_"
if(1) begin: key_type_2_
 localparam integer jj = 2;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_49_cpass,,_zy_sva_brcm_aux_cmd_49_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_50_cpass,,_zy_sva_brcm_aux_cmd_iv_50_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_51_cpass,,_zy_sva_brcm_aux_cmd_guid_51_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_52_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_52_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_53_cpass,,_zy_sva_brcm_key_type_53_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[3]"
//pragma RTLNAME "key_type[3]" "key_type_3_"
if(1) begin: key_type_3_
 localparam integer jj = 3;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_54_cpass,,_zy_sva_brcm_aux_cmd_54_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_55_cpass,,_zy_sva_brcm_aux_cmd_iv_55_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_56_cpass,,_zy_sva_brcm_aux_cmd_guid_56_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_57_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_57_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_58_cpass,,_zy_sva_brcm_key_type_58_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[4]"
//pragma RTLNAME "key_type[4]" "key_type_4_"
if(1) begin: key_type_4_
 localparam integer jj = 4;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_59_cpass,,_zy_sva_brcm_aux_cmd_59_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_60_cpass,,_zy_sva_brcm_aux_cmd_iv_60_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_61_cpass,,_zy_sva_brcm_aux_cmd_guid_61_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_62_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_62_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_63_cpass,,_zy_sva_brcm_key_type_63_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[5]"
//pragma RTLNAME "key_type[5]" "key_type_5_"
if(1) begin: key_type_5_
 localparam integer jj = 5;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_64_cpass,,_zy_sva_brcm_aux_cmd_64_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_65_cpass,,_zy_sva_brcm_aux_cmd_iv_65_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_66_cpass,,_zy_sva_brcm_aux_cmd_guid_66_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_67_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_67_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_68_cpass,,_zy_sva_brcm_key_type_68_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[6]"
//pragma RTLNAME "key_type[6]" "key_type_6_"
if(1) begin: key_type_6_
 localparam integer jj = 6;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_69_cpass,,_zy_sva_brcm_aux_cmd_69_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_70_cpass,,_zy_sva_brcm_aux_cmd_iv_70_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_71_cpass,,_zy_sva_brcm_aux_cmd_guid_71_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_72_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_72_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_73_cpass,,_zy_sva_brcm_key_type_73_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[7]"
//pragma RTLNAME "key_type[7]" "key_type_7_"
if(1) begin: key_type_7_
 localparam integer jj = 7;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_74_cpass,,_zy_sva_brcm_aux_cmd_74_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_75_cpass,,_zy_sva_brcm_aux_cmd_iv_75_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_76_cpass,,_zy_sva_brcm_aux_cmd_guid_76_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_77_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_77_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_78_cpass,,_zy_sva_brcm_key_type_78_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[8]"
//pragma RTLNAME "key_type[8]" "key_type_8_"
if(1) begin: key_type_8_
 localparam integer jj = 8;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_79_cpass,,_zy_sva_brcm_aux_cmd_79_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_80_cpass,,_zy_sva_brcm_aux_cmd_iv_80_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_81_cpass,,_zy_sva_brcm_aux_cmd_guid_81_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_82_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_82_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_83_cpass,,_zy_sva_brcm_key_type_83_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[9]"
//pragma RTLNAME "key_type[9]" "key_type_9_"
if(1) begin: key_type_9_
 localparam integer jj = 9;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_84_cpass,,_zy_sva_brcm_aux_cmd_84_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_85_cpass,,_zy_sva_brcm_aux_cmd_iv_85_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_86_cpass,,_zy_sva_brcm_aux_cmd_guid_86_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_87_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_87_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_88_cpass,,_zy_sva_brcm_key_type_88_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[10]"
//pragma RTLNAME "key_type[10]" "key_type_10_"
if(1) begin: key_type_10_
 localparam integer jj = 10;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_89_cpass,,_zy_sva_brcm_aux_cmd_89_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_90_cpass,,_zy_sva_brcm_aux_cmd_iv_90_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_91_cpass,,_zy_sva_brcm_aux_cmd_guid_91_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_92_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_92_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_93_cpass,,_zy_sva_brcm_key_type_93_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[11]"
//pragma RTLNAME "key_type[11]" "key_type_11_"
if(1) begin: key_type_11_
 localparam integer jj = 11;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_94_cpass,,_zy_sva_brcm_aux_cmd_94_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_95_cpass,,_zy_sva_brcm_aux_cmd_iv_95_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_96_cpass,,_zy_sva_brcm_aux_cmd_guid_96_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_97_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_97_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_98_cpass,,_zy_sva_brcm_key_type_98_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[12]"
//pragma RTLNAME "key_type[12]" "key_type_12_"
if(1) begin: key_type_12_
 localparam integer jj = 12;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_99_cpass,,_zy_sva_brcm_aux_cmd_99_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_100_cpass,,_zy_sva_brcm_aux_cmd_iv_100_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_101_cpass,,_zy_sva_brcm_aux_cmd_guid_101_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_102_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_102_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_103_cpass,,_zy_sva_brcm_key_type_103_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type[13]"
//pragma RTLNAME "key_type[13]" "key_type_13_"
if(1) begin: key_type_13_
 localparam integer jj = 13;
  axis_assert("brcm_aux_cmd",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_104_cpass,,_zy_sva_brcm_aux_cmd_104_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",889,3'b000);
  axis_assert("brcm_aux_cmd_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_iv_105_cpass,,_zy_sva_brcm_aux_cmd_iv_105_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",890,3'b000);
  axis_assert("brcm_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_106_cpass,,_zy_sva_brcm_aux_cmd_guid_106_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",891,3'b000);
  axis_assert("brcm_aux_cmd_guid_iv",1'b0,2'b10,,,,,,,_zy_sva_brcm_aux_cmd_guid_iv_107_cpass,,_zy_sva_brcm_aux_cmd_guid_iv_107_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",892,3'b000);
  axis_assert("brcm_key_type",1'b0,2'b10,,,,,,,_zy_sva_brcm_key_type_108_cpass,,_zy_sva_brcm_key_type_108_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",893,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0]"
//pragma RTLNAME "kdf_mode[0]" "kdf_mode_0_"
if(1) begin: kdf_mode_0_
 localparam integer ii = 0;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0]"
//pragma RTLNAME "dek_op[0]" "dek_op_0_"
 if(1) begin: dek_op_0_
  localparam integer jj = 0;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_109_cpass,,_zy_sva_brcm_kdf_ops_109_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[0].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_110_cpass,,_zy_sva_brcm_kdf_ops_110_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1]"
//pragma RTLNAME "dek_op[1]" "dek_op_1_"
 if(1) begin: dek_op_1_
  localparam integer jj = 1;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_111_cpass,,_zy_sva_brcm_kdf_ops_111_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[0].dek_op[1].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_112_cpass,,_zy_sva_brcm_kdf_ops_112_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1]"
//pragma RTLNAME "kdf_mode[1]" "kdf_mode_1_"
if(1) begin: kdf_mode_1_
 localparam integer ii = 1;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0]"
//pragma RTLNAME "dek_op[0]" "dek_op_0_"
 if(1) begin: dek_op_0_
  localparam integer jj = 0;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_113_cpass,,_zy_sva_brcm_kdf_ops_113_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[0].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_114_cpass,,_zy_sva_brcm_kdf_ops_114_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1]"
//pragma RTLNAME "dek_op[1]" "dek_op_1_"
 if(1) begin: dek_op_1_
  localparam integer jj = 1;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_115_cpass,,_zy_sva_brcm_kdf_ops_115_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[1].dek_op[1].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_116_cpass,,_zy_sva_brcm_kdf_ops_116_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2]"
//pragma RTLNAME "kdf_mode[2]" "kdf_mode_2_"
if(1) begin: kdf_mode_2_
 localparam integer ii = 2;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0]"
//pragma RTLNAME "dek_op[0]" "dek_op_0_"
 if(1) begin: dek_op_0_
  localparam integer jj = 0;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_117_cpass,,_zy_sva_brcm_kdf_ops_117_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[0].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_118_cpass,,_zy_sva_brcm_kdf_ops_118_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1]"
//pragma RTLNAME "dek_op[1]" "dek_op_1_"
 if(1) begin: dek_op_1_
  localparam integer jj = 1;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_119_cpass,,_zy_sva_brcm_kdf_ops_119_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[2].dek_op[1].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_120_cpass,,_zy_sva_brcm_kdf_ops_120_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3]"
//pragma RTLNAME "kdf_mode[3]" "kdf_mode_3_"
if(1) begin: kdf_mode_3_
 localparam integer ii = 3;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0]"
//pragma RTLNAME "dek_op[0]" "dek_op_0_"
 if(1) begin: dek_op_0_
  localparam integer jj = 0;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_121_cpass,,_zy_sva_brcm_kdf_ops_121_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[0].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_122_cpass,,_zy_sva_brcm_kdf_ops_122_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1]"
//pragma RTLNAME "dek_op[1]" "dek_op_1_"
 if(1) begin: dek_op_1_
  localparam integer jj = 1;
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1].dak_op[0]"
//pragma RTLNAME "dak_op[0]" "dak_op_0_"
  if(1) begin: dak_op_0_
   localparam integer kk = 0;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_123_cpass,,_zy_sva_brcm_kdf_ops_123_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "kdf_mode[3].dek_op[1].dak_op[1]"
//pragma RTLNAME "dak_op[1]" "dak_op_1_"
  if(1) begin: dak_op_1_
   localparam integer kk = 1;
      axis_assert("brcm_kdf_ops",1'b0,2'b10,,,,,,,_zy_sva_brcm_kdf_ops_124_cpass,,_zy_sva_brcm_kdf_ops_124_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",902,3'b000);
  end
 end
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[7]"
//pragma RTLNAME "key_type_enc_dek[7]" "key_type_enc_dek_7_"
if(1) begin: key_type_enc_dek_7_
 localparam integer nn = 7;
  axis_assert("null_gcm",1'b0,2'b10,,,,,,,_zy_sva_null_gcm_125_cpass,,_zy_sva_null_gcm_125_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1114,3'b000);
  axis_assert("sha_gcm",1'b0,2'b10,,,,,,,_zy_sva_sha_gcm_126_cpass,,_zy_sva_sha_gcm_126_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1121,3'b000);
  axis_assert("null_xts",1'b0,2'b10,,,,,,,_zy_sva_null_xts_127_cpass,,_zy_sva_null_xts_127_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1127,3'b000);
  axis_assert("sha_xts",1'b0,2'b10,,,,,,,_zy_sva_sha_xts_128_cpass,,_zy_sva_sha_xts_128_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1133,3'b000);
  axis_assert("null_null",1'b0,2'b10,,,,,,,_zy_sva_null_null_129_cpass,,_zy_sva_null_null_129_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1139,3'b000);
  axis_assert("sha_null",1'b0,2'b10,,,,,,,_zy_sva_sha_null_130_cpass,,_zy_sva_sha_null_130_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1145,3'b000);
  axis_assert("hmac_gcm",1'b0,2'b10,,,,,,,_zy_sva_hmac_gcm_131_cpass,,_zy_sva_hmac_gcm_131_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1152,3'b000);
  axis_assert("hmac_xts",1'b0,2'b10,,,,,,,_zy_sva_hmac_xts_132_cpass,,_zy_sva_hmac_xts_132_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1158,3'b000);
  axis_assert("hmac_null",1'b0,2'b10,,,,,,,_zy_sva_hmac_null_133_cpass,,_zy_sva_hmac_null_133_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1164,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek[8]"
//pragma RTLNAME "key_type_enc_dek[8]" "key_type_enc_dek_8_"
if(1) begin: key_type_enc_dek_8_
 localparam integer nn = 8;
  axis_assert("null_gcm",1'b0,2'b10,,,,,,,_zy_sva_null_gcm_134_cpass,,_zy_sva_null_gcm_134_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1114,3'b000);
  axis_assert("sha_gcm",1'b0,2'b10,,,,,,,_zy_sva_sha_gcm_135_cpass,,_zy_sva_sha_gcm_135_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1121,3'b000);
  axis_assert("null_xts",1'b0,2'b10,,,,,,,_zy_sva_null_xts_136_cpass,,_zy_sva_null_xts_136_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1127,3'b000);
  axis_assert("sha_xts",1'b0,2'b10,,,,,,,_zy_sva_sha_xts_137_cpass,,_zy_sva_sha_xts_137_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1133,3'b000);
  axis_assert("null_null",1'b0,2'b10,,,,,,,_zy_sva_null_null_138_cpass,,_zy_sva_null_null_138_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1139,3'b000);
  axis_assert("sha_null",1'b0,2'b10,,,,,,,_zy_sva_sha_null_139_cpass,,_zy_sva_sha_null_139_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1145,3'b000);
  axis_assert("hmac_gcm",1'b0,2'b10,,,,,,,_zy_sva_hmac_gcm_140_cpass,,_zy_sva_hmac_gcm_140_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1152,3'b000);
  axis_assert("hmac_xts",1'b0,2'b10,,,,,,,_zy_sva_hmac_xts_141_cpass,,_zy_sva_hmac_xts_141_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1158,3'b000);
  axis_assert("hmac_null",1'b0,2'b10,,,,,,,_zy_sva_hmac_null_142_cpass,,_zy_sva_hmac_null_142_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1164,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[10]"
//pragma RTLNAME "key_type_enc_dek_dak[10]" "key_type_enc_dek_dak_10_"
if(1) begin: key_type_enc_dek_dak_10_
 localparam integer qq = 10;
  axis_assert("null_gcm",1'b0,2'b10,,,,,,,_zy_sva_null_gcm_143_cpass,,_zy_sva_null_gcm_143_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1175,3'b000);
  axis_assert("sha_gcm",1'b0,2'b10,,,,,,,_zy_sva_sha_gcm_144_cpass,,_zy_sva_sha_gcm_144_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1182,3'b000);
  axis_assert("null_xts",1'b0,2'b10,,,,,,,_zy_sva_null_xts_145_cpass,,_zy_sva_null_xts_145_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1188,3'b000);
  axis_assert("sha_xts",1'b0,2'b10,,,,,,,_zy_sva_sha_xts_146_cpass,,_zy_sva_sha_xts_146_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1194,3'b000);
  axis_assert("null_null",1'b0,2'b10,,,,,,,_zy_sva_null_null_147_cpass,,_zy_sva_null_null_147_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1200,3'b000);
  axis_assert("sha_null",1'b0,2'b10,,,,,,,_zy_sva_sha_null_148_cpass,,_zy_sva_sha_null_148_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1206,3'b000);
  axis_assert("hmac_gcm",1'b0,2'b10,,,,,,,_zy_sva_hmac_gcm_149_cpass,,_zy_sva_hmac_gcm_149_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1213,3'b000);
  axis_assert("hmac_xts",1'b0,2'b10,,,,,,,_zy_sva_hmac_xts_150_cpass,,_zy_sva_hmac_xts_150_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1219,3'b000);
  axis_assert("hmac_null",1'b0,2'b10,,,,,,,_zy_sva_hmac_null_151_cpass,,_zy_sva_hmac_null_151_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1225,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[11]"
//pragma RTLNAME "key_type_enc_dek_dak[11]" "key_type_enc_dek_dak_11_"
if(1) begin: key_type_enc_dek_dak_11_
 localparam integer qq = 11;
  axis_assert("null_gcm",1'b0,2'b10,,,,,,,_zy_sva_null_gcm_152_cpass,,_zy_sva_null_gcm_152_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1175,3'b000);
  axis_assert("sha_gcm",1'b0,2'b10,,,,,,,_zy_sva_sha_gcm_153_cpass,,_zy_sva_sha_gcm_153_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1182,3'b000);
  axis_assert("null_xts",1'b0,2'b10,,,,,,,_zy_sva_null_xts_154_cpass,,_zy_sva_null_xts_154_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1188,3'b000);
  axis_assert("sha_xts",1'b0,2'b10,,,,,,,_zy_sva_sha_xts_155_cpass,,_zy_sva_sha_xts_155_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1194,3'b000);
  axis_assert("null_null",1'b0,2'b10,,,,,,,_zy_sva_null_null_156_cpass,,_zy_sva_null_null_156_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1200,3'b000);
  axis_assert("sha_null",1'b0,2'b10,,,,,,,_zy_sva_sha_null_157_cpass,,_zy_sva_sha_null_157_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1206,3'b000);
  axis_assert("hmac_gcm",1'b0,2'b10,,,,,,,_zy_sva_hmac_gcm_158_cpass,,_zy_sva_hmac_gcm_158_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1213,3'b000);
  axis_assert("hmac_xts",1'b0,2'b10,,,,,,,_zy_sva_hmac_xts_159_cpass,,_zy_sva_hmac_xts_159_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1219,3'b000);
  axis_assert("hmac_null",1'b0,2'b10,,,,,,,_zy_sva_hmac_null_160_cpass,,_zy_sva_hmac_null_160_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1225,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[12]"
//pragma RTLNAME "key_type_enc_dek_dak[12]" "key_type_enc_dek_dak_12_"
if(1) begin: key_type_enc_dek_dak_12_
 localparam integer qq = 12;
  axis_assert("null_gcm",1'b0,2'b10,,,,,,,_zy_sva_null_gcm_161_cpass,,_zy_sva_null_gcm_161_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1175,3'b000);
  axis_assert("sha_gcm",1'b0,2'b10,,,,,,,_zy_sva_sha_gcm_162_cpass,,_zy_sva_sha_gcm_162_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1182,3'b000);
  axis_assert("null_xts",1'b0,2'b10,,,,,,,_zy_sva_null_xts_163_cpass,,_zy_sva_null_xts_163_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1188,3'b000);
  axis_assert("sha_xts",1'b0,2'b10,,,,,,,_zy_sva_sha_xts_164_cpass,,_zy_sva_sha_xts_164_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1194,3'b000);
  axis_assert("null_null",1'b0,2'b10,,,,,,,_zy_sva_null_null_165_cpass,,_zy_sva_null_null_165_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1200,3'b000);
  axis_assert("sha_null",1'b0,2'b10,,,,,,,_zy_sva_sha_null_166_cpass,,_zy_sva_sha_null_166_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1206,3'b000);
  axis_assert("hmac_gcm",1'b0,2'b10,,,,,,,_zy_sva_hmac_gcm_167_cpass,,_zy_sva_hmac_gcm_167_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1213,3'b000);
  axis_assert("hmac_xts",1'b0,2'b10,,,,,,,_zy_sva_hmac_xts_168_cpass,,_zy_sva_hmac_xts_168_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1219,3'b000);
  axis_assert("hmac_null",1'b0,2'b10,,,,,,,_zy_sva_hmac_null_169_cpass,,_zy_sva_hmac_null_169_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1225,3'b000);
end
//pragma CVASTRPROP MODULE HDLICE cva_for_generate "key_type_enc_dek_dak[13]"
//pragma RTLNAME "key_type_enc_dek_dak[13]" "key_type_enc_dek_dak_13_"
if(1) begin: key_type_enc_dek_dak_13_
 localparam integer qq = 13;
  axis_assert("null_gcm",1'b0,2'b10,,,,,,,_zy_sva_null_gcm_170_cpass,,_zy_sva_null_gcm_170_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1175,3'b000);
  axis_assert("sha_gcm",1'b0,2'b10,,,,,,,_zy_sva_sha_gcm_171_cpass,,_zy_sva_sha_gcm_171_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1182,3'b000);
  axis_assert("null_xts",1'b0,2'b10,,,,,,,_zy_sva_null_xts_172_cpass,,_zy_sva_null_xts_172_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1188,3'b000);
  axis_assert("sha_xts",1'b0,2'b10,,,,,,,_zy_sva_sha_xts_173_cpass,,_zy_sva_sha_xts_173_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1194,3'b000);
  axis_assert("null_null",1'b0,2'b10,,,,,,,_zy_sva_null_null_174_cpass,,_zy_sva_null_null_174_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1200,3'b000);
  axis_assert("sha_null",1'b0,2'b10,,,,,,,_zy_sva_sha_null_175_cpass,,_zy_sva_sha_null_175_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1206,3'b000);
  axis_assert("hmac_gcm",1'b0,2'b10,,,,,,,_zy_sva_hmac_gcm_176_cpass,,_zy_sva_hmac_gcm_176_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1213,3'b000);
  axis_assert("hmac_xts",1'b0,2'b10,,,,,,,_zy_sva_hmac_xts_177_cpass,,_zy_sva_hmac_xts_177_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1219,3'b000);
  axis_assert("hmac_null",1'b0,2'b10,,,,,,,_zy_sva_hmac_null_178_cpass,,_zy_sva_hmac_null_178_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1225,3'b000);
end
axis_assert("key_type0_line4",1'b0,2'b10,,,,,,,_zy_sva_key_type0_line4_1_cpass,,_zy_sva_key_type0_line4_1_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",914,3'b000);
axis_assert("key_type0_line5a",1'b0,2'b10,,,,,,,_zy_sva_key_type0_line5a_2_cpass,,_zy_sva_key_type0_line5a_2_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",920,3'b000);
axis_assert("key_type0_line5b",1'b0,2'b10,,,,,,,_zy_sva_key_type0_line5b_3_cpass,,_zy_sva_key_type0_line5b_3_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",926,3'b000);
axis_assert("key_type1_line7a",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line7a_4_cpass,,_zy_sva_key_type1_line7a_4_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",936,3'b000);
axis_assert("key_type1_line7b",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line7b_5_cpass,,_zy_sva_key_type1_line7b_5_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",944,3'b000);
axis_assert("key_type1_line8a",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line8a_6_cpass,,_zy_sva_key_type1_line8a_6_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",952,3'b000);
axis_assert("key_type1_line8b",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line8b_7_cpass,,_zy_sva_key_type1_line8b_7_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",960,3'b000);
axis_assert("key_type1_line9",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line9_8_cpass,,_zy_sva_key_type1_line9_8_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",969,3'b000);
axis_assert("key_type1_line10",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line10_9_cpass,,_zy_sva_key_type1_line10_9_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",977,3'b000);
axis_assert("key_type1_line11a",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line11a_10_cpass,,_zy_sva_key_type1_line11a_10_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",983,3'b000);
axis_assert("key_type1_line11b",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line11b_11_cpass,,_zy_sva_key_type1_line11b_11_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",989,3'b000);
axis_assert("key_type1_line11c",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line11c_12_cpass,,_zy_sva_key_type1_line11c_12_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",995,3'b000);
axis_assert("key_type1_line11d",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line11d_13_cpass,,_zy_sva_key_type1_line11d_13_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1001,3'b000);
axis_assert("key_type1_line12a",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line12a_14_cpass,,_zy_sva_key_type1_line12a_14_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1007,3'b000);
axis_assert("key_type1_line12b",1'b0,2'b10,,,,,,,_zy_sva_key_type1_line12b_15_cpass,,_zy_sva_key_type1_line12b_15_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1014,3'b000);
axis_assert("key_type9_line14",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line14_16_cpass,,_zy_sva_key_type9_line14_16_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1023,3'b000);
axis_assert("key_type9_line15",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line15_17_cpass,,_zy_sva_key_type9_line15_17_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1030,3'b000);
axis_assert("key_type9_line16a",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line16a_18_cpass,,_zy_sva_key_type9_line16a_18_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1036,3'b000);
axis_assert("key_type9_line16b",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line16b_19_cpass,,_zy_sva_key_type9_line16b_19_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1042,3'b000);
axis_assert("key_type9_line17a",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line17a_20_cpass,,_zy_sva_key_type9_line17a_20_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1050,3'b000);
axis_assert("key_type9_line17b",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line17b_21_cpass,,_zy_sva_key_type9_line17b_21_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1059,3'b000);
axis_assert("key_type9_line18a",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line18a_22_cpass,,_zy_sva_key_type9_line18a_22_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1066,3'b000);
axis_assert("key_type9_line18b",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line18b_23_cpass,,_zy_sva_key_type9_line18b_23_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1074,3'b000);
axis_assert("key_type9_line19a",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line19a_24_cpass,,_zy_sva_key_type9_line19a_24_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1081,3'b000);
axis_assert("key_type9_line19b",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line19b_25_cpass,,_zy_sva_key_type9_line19b_25_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1088,3'b000);
axis_assert("key_type9_line19c",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line19c_26_cpass,,_zy_sva_key_type9_line19c_26_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1094,3'b000);
axis_assert("key_type9_line19d",1'b0,2'b10,,,,,,,_zy_sva_key_type9_line19d_27_cpass,,_zy_sva_key_type9_line19d_27_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1101,3'b000);
axis_assert("guid_miss_aux_cmd_0",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_0_28_cpass,,_zy_sva_guid_miss_aux_cmd_0_28_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1234,3'b000);
axis_assert("guid_miss_aux_cmd_1",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_1_29_cpass,,_zy_sva_guid_miss_aux_cmd_1_29_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1240,3'b000);
axis_assert("guid_miss_aux_cmd_2",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_2_30_cpass,,_zy_sva_guid_miss_aux_cmd_2_30_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1246,3'b000);
axis_assert("guid_miss_aux_cmd_3",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_3_31_cpass,,_zy_sva_guid_miss_aux_cmd_3_31_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1252,3'b000);
axis_assert("guid_miss_aux_cmd_iv_0",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_iv_0_32_cpass,,_zy_sva_guid_miss_aux_cmd_iv_0_32_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1258,3'b000);
axis_assert("guid_miss_aux_cmd_iv_1",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_iv_1_33_cpass,,_zy_sva_guid_miss_aux_cmd_iv_1_33_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1264,3'b000);
axis_assert("guid_miss_aux_cmd_iv_2",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_iv_2_34_cpass,,_zy_sva_guid_miss_aux_cmd_iv_2_34_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1270,3'b000);
axis_assert("guid_miss_aux_cmd_iv_3",1'b0,2'b10,,,,,,,_zy_sva_guid_miss_aux_cmd_iv_3_35_cpass,,_zy_sva_guid_miss_aux_cmd_iv_3_35_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1276,3'b000);
axis_assert("iv_miss_aux_cmd_0",1'b0,2'b10,,,,,,,_zy_sva_iv_miss_aux_cmd_0_36_cpass,,_zy_sva_iv_miss_aux_cmd_0_36_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1282,3'b000);
axis_assert("iv_miss_aux_cmd_1",1'b0,2'b10,,,,,,,_zy_sva_iv_miss_aux_cmd_1_37_cpass,,_zy_sva_iv_miss_aux_cmd_1_37_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1287,3'b000);
axis_assert("iv_miss_aux_cmd_guid",1'b0,2'b10,,,,,,,_zy_sva_iv_miss_aux_cmd_guid_38_cpass,,_zy_sva_iv_miss_aux_cmd_guid_38_ccheck,,"/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_tlv_parser.v",1292,3'b000);
// pragma CVASTRPROP MODULE cr_kme_tlv_parser PROP_RANOFF TRUE
  //pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 key_type 0 13 "
  //pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 kdf_mode 0 3 "
  //pragma CVASTRPROP MODULE HDLICE cva_for_generate_2 "1 dek_op 0 1 "
  //pragma CVASTRPROP MODULE HDLICE cva_for_generate_3 "2 dak_op 0 1 "
  //pragma CVASTRPROP MODULE HDLICE cva_for_generate_4 "-1 key_type_enc_dek 7 8 "
  //pragma CVASTRPROP MODULE HDLICE cva_for_generate_5 "-1 key_type_enc_dek_dak 10 13 "
endmodule

