
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_kdf_stream_gen ( kdfstream_cmdfifo_ack, cmdfifo_hash_valid, 
	cmdfifo_hash_skip, cmdfifo_hash_small_size, hash_len_data_out, 
	hash_len_data_out_valid, in_hash_valid, in_hash_eof, in_hash_eoc, 
	in_hash_num_bytes, in_hash_data, clk, rst_n, cmdfifo_kdfstream_valid, 
	.cmdfifo_kdfstream_cmd( {\cmdfifo_kdfstream_cmd.combo_mode [0], 
	\cmdfifo_kdfstream_cmd.skip [0], \cmdfifo_kdfstream_cmd.guid [255], 
	\cmdfifo_kdfstream_cmd.guid [254], \cmdfifo_kdfstream_cmd.guid [253], 
	\cmdfifo_kdfstream_cmd.guid [252], \cmdfifo_kdfstream_cmd.guid [251], 
	\cmdfifo_kdfstream_cmd.guid [250], \cmdfifo_kdfstream_cmd.guid [249], 
	\cmdfifo_kdfstream_cmd.guid [248], \cmdfifo_kdfstream_cmd.guid [247], 
	\cmdfifo_kdfstream_cmd.guid [246], \cmdfifo_kdfstream_cmd.guid [245], 
	\cmdfifo_kdfstream_cmd.guid [244], \cmdfifo_kdfstream_cmd.guid [243], 
	\cmdfifo_kdfstream_cmd.guid [242], \cmdfifo_kdfstream_cmd.guid [241], 
	\cmdfifo_kdfstream_cmd.guid [240], \cmdfifo_kdfstream_cmd.guid [239], 
	\cmdfifo_kdfstream_cmd.guid [238], \cmdfifo_kdfstream_cmd.guid [237], 
	\cmdfifo_kdfstream_cmd.guid [236], \cmdfifo_kdfstream_cmd.guid [235], 
	\cmdfifo_kdfstream_cmd.guid [234], \cmdfifo_kdfstream_cmd.guid [233], 
	\cmdfifo_kdfstream_cmd.guid [232], \cmdfifo_kdfstream_cmd.guid [231], 
	\cmdfifo_kdfstream_cmd.guid [230], \cmdfifo_kdfstream_cmd.guid [229], 
	\cmdfifo_kdfstream_cmd.guid [228], \cmdfifo_kdfstream_cmd.guid [227], 
	\cmdfifo_kdfstream_cmd.guid [226], \cmdfifo_kdfstream_cmd.guid [225], 
	\cmdfifo_kdfstream_cmd.guid [224], \cmdfifo_kdfstream_cmd.guid [223], 
	\cmdfifo_kdfstream_cmd.guid [222], \cmdfifo_kdfstream_cmd.guid [221], 
	\cmdfifo_kdfstream_cmd.guid [220], \cmdfifo_kdfstream_cmd.guid [219], 
	\cmdfifo_kdfstream_cmd.guid [218], \cmdfifo_kdfstream_cmd.guid [217], 
	\cmdfifo_kdfstream_cmd.guid [216], \cmdfifo_kdfstream_cmd.guid [215], 
	\cmdfifo_kdfstream_cmd.guid [214], \cmdfifo_kdfstream_cmd.guid [213], 
	\cmdfifo_kdfstream_cmd.guid [212], \cmdfifo_kdfstream_cmd.guid [211], 
	\cmdfifo_kdfstream_cmd.guid [210], \cmdfifo_kdfstream_cmd.guid [209], 
	\cmdfifo_kdfstream_cmd.guid [208], \cmdfifo_kdfstream_cmd.guid [207], 
	\cmdfifo_kdfstream_cmd.guid [206], \cmdfifo_kdfstream_cmd.guid [205], 
	\cmdfifo_kdfstream_cmd.guid [204], \cmdfifo_kdfstream_cmd.guid [203], 
	\cmdfifo_kdfstream_cmd.guid [202], \cmdfifo_kdfstream_cmd.guid [201], 
	\cmdfifo_kdfstream_cmd.guid [200], \cmdfifo_kdfstream_cmd.guid [199], 
	\cmdfifo_kdfstream_cmd.guid [198], \cmdfifo_kdfstream_cmd.guid [197], 
	\cmdfifo_kdfstream_cmd.guid [196], \cmdfifo_kdfstream_cmd.guid [195], 
	\cmdfifo_kdfstream_cmd.guid [194], \cmdfifo_kdfstream_cmd.guid [193], 
	\cmdfifo_kdfstream_cmd.guid [192], \cmdfifo_kdfstream_cmd.guid [191], 
	\cmdfifo_kdfstream_cmd.guid [190], \cmdfifo_kdfstream_cmd.guid [189], 
	\cmdfifo_kdfstream_cmd.guid [188], \cmdfifo_kdfstream_cmd.guid [187], 
	\cmdfifo_kdfstream_cmd.guid [186], \cmdfifo_kdfstream_cmd.guid [185], 
	\cmdfifo_kdfstream_cmd.guid [184], \cmdfifo_kdfstream_cmd.guid [183], 
	\cmdfifo_kdfstream_cmd.guid [182], \cmdfifo_kdfstream_cmd.guid [181], 
	\cmdfifo_kdfstream_cmd.guid [180], \cmdfifo_kdfstream_cmd.guid [179], 
	\cmdfifo_kdfstream_cmd.guid [178], \cmdfifo_kdfstream_cmd.guid [177], 
	\cmdfifo_kdfstream_cmd.guid [176], \cmdfifo_kdfstream_cmd.guid [175], 
	\cmdfifo_kdfstream_cmd.guid [174], \cmdfifo_kdfstream_cmd.guid [173], 
	\cmdfifo_kdfstream_cmd.guid [172], \cmdfifo_kdfstream_cmd.guid [171], 
	\cmdfifo_kdfstream_cmd.guid [170], \cmdfifo_kdfstream_cmd.guid [169], 
	\cmdfifo_kdfstream_cmd.guid [168], \cmdfifo_kdfstream_cmd.guid [167], 
	\cmdfifo_kdfstream_cmd.guid [166], \cmdfifo_kdfstream_cmd.guid [165], 
	\cmdfifo_kdfstream_cmd.guid [164], \cmdfifo_kdfstream_cmd.guid [163], 
	\cmdfifo_kdfstream_cmd.guid [162], \cmdfifo_kdfstream_cmd.guid [161], 
	\cmdfifo_kdfstream_cmd.guid [160], \cmdfifo_kdfstream_cmd.guid [159], 
	\cmdfifo_kdfstream_cmd.guid [158], \cmdfifo_kdfstream_cmd.guid [157], 
	\cmdfifo_kdfstream_cmd.guid [156], \cmdfifo_kdfstream_cmd.guid [155], 
	\cmdfifo_kdfstream_cmd.guid [154], \cmdfifo_kdfstream_cmd.guid [153], 
	\cmdfifo_kdfstream_cmd.guid [152], \cmdfifo_kdfstream_cmd.guid [151], 
	\cmdfifo_kdfstream_cmd.guid [150], \cmdfifo_kdfstream_cmd.guid [149], 
	\cmdfifo_kdfstream_cmd.guid [148], \cmdfifo_kdfstream_cmd.guid [147], 
	\cmdfifo_kdfstream_cmd.guid [146], \cmdfifo_kdfstream_cmd.guid [145], 
	\cmdfifo_kdfstream_cmd.guid [144], \cmdfifo_kdfstream_cmd.guid [143], 
	\cmdfifo_kdfstream_cmd.guid [142], \cmdfifo_kdfstream_cmd.guid [141], 
	\cmdfifo_kdfstream_cmd.guid [140], \cmdfifo_kdfstream_cmd.guid [139], 
	\cmdfifo_kdfstream_cmd.guid [138], \cmdfifo_kdfstream_cmd.guid [137], 
	\cmdfifo_kdfstream_cmd.guid [136], \cmdfifo_kdfstream_cmd.guid [135], 
	\cmdfifo_kdfstream_cmd.guid [134], \cmdfifo_kdfstream_cmd.guid [133], 
	\cmdfifo_kdfstream_cmd.guid [132], \cmdfifo_kdfstream_cmd.guid [131], 
	\cmdfifo_kdfstream_cmd.guid [130], \cmdfifo_kdfstream_cmd.guid [129], 
	\cmdfifo_kdfstream_cmd.guid [128], \cmdfifo_kdfstream_cmd.guid [127], 
	\cmdfifo_kdfstream_cmd.guid [126], \cmdfifo_kdfstream_cmd.guid [125], 
	\cmdfifo_kdfstream_cmd.guid [124], \cmdfifo_kdfstream_cmd.guid [123], 
	\cmdfifo_kdfstream_cmd.guid [122], \cmdfifo_kdfstream_cmd.guid [121], 
	\cmdfifo_kdfstream_cmd.guid [120], \cmdfifo_kdfstream_cmd.guid [119], 
	\cmdfifo_kdfstream_cmd.guid [118], \cmdfifo_kdfstream_cmd.guid [117], 
	\cmdfifo_kdfstream_cmd.guid [116], \cmdfifo_kdfstream_cmd.guid [115], 
	\cmdfifo_kdfstream_cmd.guid [114], \cmdfifo_kdfstream_cmd.guid [113], 
	\cmdfifo_kdfstream_cmd.guid [112], \cmdfifo_kdfstream_cmd.guid [111], 
	\cmdfifo_kdfstream_cmd.guid [110], \cmdfifo_kdfstream_cmd.guid [109], 
	\cmdfifo_kdfstream_cmd.guid [108], \cmdfifo_kdfstream_cmd.guid [107], 
	\cmdfifo_kdfstream_cmd.guid [106], \cmdfifo_kdfstream_cmd.guid [105], 
	\cmdfifo_kdfstream_cmd.guid [104], \cmdfifo_kdfstream_cmd.guid [103], 
	\cmdfifo_kdfstream_cmd.guid [102], \cmdfifo_kdfstream_cmd.guid [101], 
	\cmdfifo_kdfstream_cmd.guid [100], \cmdfifo_kdfstream_cmd.guid [99], 
	\cmdfifo_kdfstream_cmd.guid [98], \cmdfifo_kdfstream_cmd.guid [97], 
	\cmdfifo_kdfstream_cmd.guid [96], \cmdfifo_kdfstream_cmd.guid [95], 
	\cmdfifo_kdfstream_cmd.guid [94], \cmdfifo_kdfstream_cmd.guid [93], 
	\cmdfifo_kdfstream_cmd.guid [92], \cmdfifo_kdfstream_cmd.guid [91], 
	\cmdfifo_kdfstream_cmd.guid [90], \cmdfifo_kdfstream_cmd.guid [89], 
	\cmdfifo_kdfstream_cmd.guid [88], \cmdfifo_kdfstream_cmd.guid [87], 
	\cmdfifo_kdfstream_cmd.guid [86], \cmdfifo_kdfstream_cmd.guid [85], 
	\cmdfifo_kdfstream_cmd.guid [84], \cmdfifo_kdfstream_cmd.guid [83], 
	\cmdfifo_kdfstream_cmd.guid [82], \cmdfifo_kdfstream_cmd.guid [81], 
	\cmdfifo_kdfstream_cmd.guid [80], \cmdfifo_kdfstream_cmd.guid [79], 
	\cmdfifo_kdfstream_cmd.guid [78], \cmdfifo_kdfstream_cmd.guid [77], 
	\cmdfifo_kdfstream_cmd.guid [76], \cmdfifo_kdfstream_cmd.guid [75], 
	\cmdfifo_kdfstream_cmd.guid [74], \cmdfifo_kdfstream_cmd.guid [73], 
	\cmdfifo_kdfstream_cmd.guid [72], \cmdfifo_kdfstream_cmd.guid [71], 
	\cmdfifo_kdfstream_cmd.guid [70], \cmdfifo_kdfstream_cmd.guid [69], 
	\cmdfifo_kdfstream_cmd.guid [68], \cmdfifo_kdfstream_cmd.guid [67], 
	\cmdfifo_kdfstream_cmd.guid [66], \cmdfifo_kdfstream_cmd.guid [65], 
	\cmdfifo_kdfstream_cmd.guid [64], \cmdfifo_kdfstream_cmd.guid [63], 
	\cmdfifo_kdfstream_cmd.guid [62], \cmdfifo_kdfstream_cmd.guid [61], 
	\cmdfifo_kdfstream_cmd.guid [60], \cmdfifo_kdfstream_cmd.guid [59], 
	\cmdfifo_kdfstream_cmd.guid [58], \cmdfifo_kdfstream_cmd.guid [57], 
	\cmdfifo_kdfstream_cmd.guid [56], \cmdfifo_kdfstream_cmd.guid [55], 
	\cmdfifo_kdfstream_cmd.guid [54], \cmdfifo_kdfstream_cmd.guid [53], 
	\cmdfifo_kdfstream_cmd.guid [52], \cmdfifo_kdfstream_cmd.guid [51], 
	\cmdfifo_kdfstream_cmd.guid [50], \cmdfifo_kdfstream_cmd.guid [49], 
	\cmdfifo_kdfstream_cmd.guid [48], \cmdfifo_kdfstream_cmd.guid [47], 
	\cmdfifo_kdfstream_cmd.guid [46], \cmdfifo_kdfstream_cmd.guid [45], 
	\cmdfifo_kdfstream_cmd.guid [44], \cmdfifo_kdfstream_cmd.guid [43], 
	\cmdfifo_kdfstream_cmd.guid [42], \cmdfifo_kdfstream_cmd.guid [41], 
	\cmdfifo_kdfstream_cmd.guid [40], \cmdfifo_kdfstream_cmd.guid [39], 
	\cmdfifo_kdfstream_cmd.guid [38], \cmdfifo_kdfstream_cmd.guid [37], 
	\cmdfifo_kdfstream_cmd.guid [36], \cmdfifo_kdfstream_cmd.guid [35], 
	\cmdfifo_kdfstream_cmd.guid [34], \cmdfifo_kdfstream_cmd.guid [33], 
	\cmdfifo_kdfstream_cmd.guid [32], \cmdfifo_kdfstream_cmd.guid [31], 
	\cmdfifo_kdfstream_cmd.guid [30], \cmdfifo_kdfstream_cmd.guid [29], 
	\cmdfifo_kdfstream_cmd.guid [28], \cmdfifo_kdfstream_cmd.guid [27], 
	\cmdfifo_kdfstream_cmd.guid [26], \cmdfifo_kdfstream_cmd.guid [25], 
	\cmdfifo_kdfstream_cmd.guid [24], \cmdfifo_kdfstream_cmd.guid [23], 
	\cmdfifo_kdfstream_cmd.guid [22], \cmdfifo_kdfstream_cmd.guid [21], 
	\cmdfifo_kdfstream_cmd.guid [20], \cmdfifo_kdfstream_cmd.guid [19], 
	\cmdfifo_kdfstream_cmd.guid [18], \cmdfifo_kdfstream_cmd.guid [17], 
	\cmdfifo_kdfstream_cmd.guid [16], \cmdfifo_kdfstream_cmd.guid [15], 
	\cmdfifo_kdfstream_cmd.guid [14], \cmdfifo_kdfstream_cmd.guid [13], 
	\cmdfifo_kdfstream_cmd.guid [12], \cmdfifo_kdfstream_cmd.guid [11], 
	\cmdfifo_kdfstream_cmd.guid [10], \cmdfifo_kdfstream_cmd.guid [9], 
	\cmdfifo_kdfstream_cmd.guid [8], \cmdfifo_kdfstream_cmd.guid [7], 
	\cmdfifo_kdfstream_cmd.guid [6], \cmdfifo_kdfstream_cmd.guid [5], 
	\cmdfifo_kdfstream_cmd.guid [4], \cmdfifo_kdfstream_cmd.guid [3], 
	\cmdfifo_kdfstream_cmd.guid [2], \cmdfifo_kdfstream_cmd.guid [1], 
	\cmdfifo_kdfstream_cmd.guid [0], 
	\cmdfifo_kdfstream_cmd.label_index [2], 
	\cmdfifo_kdfstream_cmd.label_index [1], 
	\cmdfifo_kdfstream_cmd.label_index [0], 
	\cmdfifo_kdfstream_cmd.num_iter [1], 
	\cmdfifo_kdfstream_cmd.num_iter [0]} ), .labels( {
	\labels[7].guid_size[0] , \labels[7].label_size[5] , 
	\labels[7].label_size[4] , \labels[7].label_size[3] , 
	\labels[7].label_size[2] , \labels[7].label_size[1] , 
	\labels[7].label_size[0] , \labels[7].label[255] , 
	\labels[7].label[254] , \labels[7].label[253] , 
	\labels[7].label[252] , \labels[7].label[251] , 
	\labels[7].label[250] , \labels[7].label[249] , 
	\labels[7].label[248] , \labels[7].label[247] , 
	\labels[7].label[246] , \labels[7].label[245] , 
	\labels[7].label[244] , \labels[7].label[243] , 
	\labels[7].label[242] , \labels[7].label[241] , 
	\labels[7].label[240] , \labels[7].label[239] , 
	\labels[7].label[238] , \labels[7].label[237] , 
	\labels[7].label[236] , \labels[7].label[235] , 
	\labels[7].label[234] , \labels[7].label[233] , 
	\labels[7].label[232] , \labels[7].label[231] , 
	\labels[7].label[230] , \labels[7].label[229] , 
	\labels[7].label[228] , \labels[7].label[227] , 
	\labels[7].label[226] , \labels[7].label[225] , 
	\labels[7].label[224] , \labels[7].label[223] , 
	\labels[7].label[222] , \labels[7].label[221] , 
	\labels[7].label[220] , \labels[7].label[219] , 
	\labels[7].label[218] , \labels[7].label[217] , 
	\labels[7].label[216] , \labels[7].label[215] , 
	\labels[7].label[214] , \labels[7].label[213] , 
	\labels[7].label[212] , \labels[7].label[211] , 
	\labels[7].label[210] , \labels[7].label[209] , 
	\labels[7].label[208] , \labels[7].label[207] , 
	\labels[7].label[206] , \labels[7].label[205] , 
	\labels[7].label[204] , \labels[7].label[203] , 
	\labels[7].label[202] , \labels[7].label[201] , 
	\labels[7].label[200] , \labels[7].label[199] , 
	\labels[7].label[198] , \labels[7].label[197] , 
	\labels[7].label[196] , \labels[7].label[195] , 
	\labels[7].label[194] , \labels[7].label[193] , 
	\labels[7].label[192] , \labels[7].label[191] , 
	\labels[7].label[190] , \labels[7].label[189] , 
	\labels[7].label[188] , \labels[7].label[187] , 
	\labels[7].label[186] , \labels[7].label[185] , 
	\labels[7].label[184] , \labels[7].label[183] , 
	\labels[7].label[182] , \labels[7].label[181] , 
	\labels[7].label[180] , \labels[7].label[179] , 
	\labels[7].label[178] , \labels[7].label[177] , 
	\labels[7].label[176] , \labels[7].label[175] , 
	\labels[7].label[174] , \labels[7].label[173] , 
	\labels[7].label[172] , \labels[7].label[171] , 
	\labels[7].label[170] , \labels[7].label[169] , 
	\labels[7].label[168] , \labels[7].label[167] , 
	\labels[7].label[166] , \labels[7].label[165] , 
	\labels[7].label[164] , \labels[7].label[163] , 
	\labels[7].label[162] , \labels[7].label[161] , 
	\labels[7].label[160] , \labels[7].label[159] , 
	\labels[7].label[158] , \labels[7].label[157] , 
	\labels[7].label[156] , \labels[7].label[155] , 
	\labels[7].label[154] , \labels[7].label[153] , 
	\labels[7].label[152] , \labels[7].label[151] , 
	\labels[7].label[150] , \labels[7].label[149] , 
	\labels[7].label[148] , \labels[7].label[147] , 
	\labels[7].label[146] , \labels[7].label[145] , 
	\labels[7].label[144] , \labels[7].label[143] , 
	\labels[7].label[142] , \labels[7].label[141] , 
	\labels[7].label[140] , \labels[7].label[139] , 
	\labels[7].label[138] , \labels[7].label[137] , 
	\labels[7].label[136] , \labels[7].label[135] , 
	\labels[7].label[134] , \labels[7].label[133] , 
	\labels[7].label[132] , \labels[7].label[131] , 
	\labels[7].label[130] , \labels[7].label[129] , 
	\labels[7].label[128] , \labels[7].label[127] , 
	\labels[7].label[126] , \labels[7].label[125] , 
	\labels[7].label[124] , \labels[7].label[123] , 
	\labels[7].label[122] , \labels[7].label[121] , 
	\labels[7].label[120] , \labels[7].label[119] , 
	\labels[7].label[118] , \labels[7].label[117] , 
	\labels[7].label[116] , \labels[7].label[115] , 
	\labels[7].label[114] , \labels[7].label[113] , 
	\labels[7].label[112] , \labels[7].label[111] , 
	\labels[7].label[110] , \labels[7].label[109] , 
	\labels[7].label[108] , \labels[7].label[107] , 
	\labels[7].label[106] , \labels[7].label[105] , 
	\labels[7].label[104] , \labels[7].label[103] , 
	\labels[7].label[102] , \labels[7].label[101] , 
	\labels[7].label[100] , \labels[7].label[99] , \labels[7].label[98] , 
	\labels[7].label[97] , \labels[7].label[96] , \labels[7].label[95] , 
	\labels[7].label[94] , \labels[7].label[93] , \labels[7].label[92] , 
	\labels[7].label[91] , \labels[7].label[90] , \labels[7].label[89] , 
	\labels[7].label[88] , \labels[7].label[87] , \labels[7].label[86] , 
	\labels[7].label[85] , \labels[7].label[84] , \labels[7].label[83] , 
	\labels[7].label[82] , \labels[7].label[81] , \labels[7].label[80] , 
	\labels[7].label[79] , \labels[7].label[78] , \labels[7].label[77] , 
	\labels[7].label[76] , \labels[7].label[75] , \labels[7].label[74] , 
	\labels[7].label[73] , \labels[7].label[72] , \labels[7].label[71] , 
	\labels[7].label[70] , \labels[7].label[69] , \labels[7].label[68] , 
	\labels[7].label[67] , \labels[7].label[66] , \labels[7].label[65] , 
	\labels[7].label[64] , \labels[7].label[63] , \labels[7].label[62] , 
	\labels[7].label[61] , \labels[7].label[60] , \labels[7].label[59] , 
	\labels[7].label[58] , \labels[7].label[57] , \labels[7].label[56] , 
	\labels[7].label[55] , \labels[7].label[54] , \labels[7].label[53] , 
	\labels[7].label[52] , \labels[7].label[51] , \labels[7].label[50] , 
	\labels[7].label[49] , \labels[7].label[48] , \labels[7].label[47] , 
	\labels[7].label[46] , \labels[7].label[45] , \labels[7].label[44] , 
	\labels[7].label[43] , \labels[7].label[42] , \labels[7].label[41] , 
	\labels[7].label[40] , \labels[7].label[39] , \labels[7].label[38] , 
	\labels[7].label[37] , \labels[7].label[36] , \labels[7].label[35] , 
	\labels[7].label[34] , \labels[7].label[33] , \labels[7].label[32] , 
	\labels[7].label[31] , \labels[7].label[30] , \labels[7].label[29] , 
	\labels[7].label[28] , \labels[7].label[27] , \labels[7].label[26] , 
	\labels[7].label[25] , \labels[7].label[24] , \labels[7].label[23] , 
	\labels[7].label[22] , \labels[7].label[21] , \labels[7].label[20] , 
	\labels[7].label[19] , \labels[7].label[18] , \labels[7].label[17] , 
	\labels[7].label[16] , \labels[7].label[15] , \labels[7].label[14] , 
	\labels[7].label[13] , \labels[7].label[12] , \labels[7].label[11] , 
	\labels[7].label[10] , \labels[7].label[9] , \labels[7].label[8] , 
	\labels[7].label[7] , \labels[7].label[6] , \labels[7].label[5] , 
	\labels[7].label[4] , \labels[7].label[3] , \labels[7].label[2] , 
	\labels[7].label[1] , \labels[7].label[0] , 
	\labels[7].delimiter_valid[0] , \labels[7].delimiter[7] , 
	\labels[7].delimiter[6] , \labels[7].delimiter[5] , 
	\labels[7].delimiter[4] , \labels[7].delimiter[3] , 
	\labels[7].delimiter[2] , \labels[7].delimiter[1] , 
	\labels[7].delimiter[0] , \labels[6].guid_size[0] , 
	\labels[6].label_size[5] , \labels[6].label_size[4] , 
	\labels[6].label_size[3] , \labels[6].label_size[2] , 
	\labels[6].label_size[1] , \labels[6].label_size[0] , 
	\labels[6].label[255] , \labels[6].label[254] , 
	\labels[6].label[253] , \labels[6].label[252] , 
	\labels[6].label[251] , \labels[6].label[250] , 
	\labels[6].label[249] , \labels[6].label[248] , 
	\labels[6].label[247] , \labels[6].label[246] , 
	\labels[6].label[245] , \labels[6].label[244] , 
	\labels[6].label[243] , \labels[6].label[242] , 
	\labels[6].label[241] , \labels[6].label[240] , 
	\labels[6].label[239] , \labels[6].label[238] , 
	\labels[6].label[237] , \labels[6].label[236] , 
	\labels[6].label[235] , \labels[6].label[234] , 
	\labels[6].label[233] , \labels[6].label[232] , 
	\labels[6].label[231] , \labels[6].label[230] , 
	\labels[6].label[229] , \labels[6].label[228] , 
	\labels[6].label[227] , \labels[6].label[226] , 
	\labels[6].label[225] , \labels[6].label[224] , 
	\labels[6].label[223] , \labels[6].label[222] , 
	\labels[6].label[221] , \labels[6].label[220] , 
	\labels[6].label[219] , \labels[6].label[218] , 
	\labels[6].label[217] , \labels[6].label[216] , 
	\labels[6].label[215] , \labels[6].label[214] , 
	\labels[6].label[213] , \labels[6].label[212] , 
	\labels[6].label[211] , \labels[6].label[210] , 
	\labels[6].label[209] , \labels[6].label[208] , 
	\labels[6].label[207] , \labels[6].label[206] , 
	\labels[6].label[205] , \labels[6].label[204] , 
	\labels[6].label[203] , \labels[6].label[202] , 
	\labels[6].label[201] , \labels[6].label[200] , 
	\labels[6].label[199] , \labels[6].label[198] , 
	\labels[6].label[197] , \labels[6].label[196] , 
	\labels[6].label[195] , \labels[6].label[194] , 
	\labels[6].label[193] , \labels[6].label[192] , 
	\labels[6].label[191] , \labels[6].label[190] , 
	\labels[6].label[189] , \labels[6].label[188] , 
	\labels[6].label[187] , \labels[6].label[186] , 
	\labels[6].label[185] , \labels[6].label[184] , 
	\labels[6].label[183] , \labels[6].label[182] , 
	\labels[6].label[181] , \labels[6].label[180] , 
	\labels[6].label[179] , \labels[6].label[178] , 
	\labels[6].label[177] , \labels[6].label[176] , 
	\labels[6].label[175] , \labels[6].label[174] , 
	\labels[6].label[173] , \labels[6].label[172] , 
	\labels[6].label[171] , \labels[6].label[170] , 
	\labels[6].label[169] , \labels[6].label[168] , 
	\labels[6].label[167] , \labels[6].label[166] , 
	\labels[6].label[165] , \labels[6].label[164] , 
	\labels[6].label[163] , \labels[6].label[162] , 
	\labels[6].label[161] , \labels[6].label[160] , 
	\labels[6].label[159] , \labels[6].label[158] , 
	\labels[6].label[157] , \labels[6].label[156] , 
	\labels[6].label[155] , \labels[6].label[154] , 
	\labels[6].label[153] , \labels[6].label[152] , 
	\labels[6].label[151] , \labels[6].label[150] , 
	\labels[6].label[149] , \labels[6].label[148] , 
	\labels[6].label[147] , \labels[6].label[146] , 
	\labels[6].label[145] , \labels[6].label[144] , 
	\labels[6].label[143] , \labels[6].label[142] , 
	\labels[6].label[141] , \labels[6].label[140] , 
	\labels[6].label[139] , \labels[6].label[138] , 
	\labels[6].label[137] , \labels[6].label[136] , 
	\labels[6].label[135] , \labels[6].label[134] , 
	\labels[6].label[133] , \labels[6].label[132] , 
	\labels[6].label[131] , \labels[6].label[130] , 
	\labels[6].label[129] , \labels[6].label[128] , 
	\labels[6].label[127] , \labels[6].label[126] , 
	\labels[6].label[125] , \labels[6].label[124] , 
	\labels[6].label[123] , \labels[6].label[122] , 
	\labels[6].label[121] , \labels[6].label[120] , 
	\labels[6].label[119] , \labels[6].label[118] , 
	\labels[6].label[117] , \labels[6].label[116] , 
	\labels[6].label[115] , \labels[6].label[114] , 
	\labels[6].label[113] , \labels[6].label[112] , 
	\labels[6].label[111] , \labels[6].label[110] , 
	\labels[6].label[109] , \labels[6].label[108] , 
	\labels[6].label[107] , \labels[6].label[106] , 
	\labels[6].label[105] , \labels[6].label[104] , 
	\labels[6].label[103] , \labels[6].label[102] , 
	\labels[6].label[101] , \labels[6].label[100] , 
	\labels[6].label[99] , \labels[6].label[98] , \labels[6].label[97] , 
	\labels[6].label[96] , \labels[6].label[95] , \labels[6].label[94] , 
	\labels[6].label[93] , \labels[6].label[92] , \labels[6].label[91] , 
	\labels[6].label[90] , \labels[6].label[89] , \labels[6].label[88] , 
	\labels[6].label[87] , \labels[6].label[86] , \labels[6].label[85] , 
	\labels[6].label[84] , \labels[6].label[83] , \labels[6].label[82] , 
	\labels[6].label[81] , \labels[6].label[80] , \labels[6].label[79] , 
	\labels[6].label[78] , \labels[6].label[77] , \labels[6].label[76] , 
	\labels[6].label[75] , \labels[6].label[74] , \labels[6].label[73] , 
	\labels[6].label[72] , \labels[6].label[71] , \labels[6].label[70] , 
	\labels[6].label[69] , \labels[6].label[68] , \labels[6].label[67] , 
	\labels[6].label[66] , \labels[6].label[65] , \labels[6].label[64] , 
	\labels[6].label[63] , \labels[6].label[62] , \labels[6].label[61] , 
	\labels[6].label[60] , \labels[6].label[59] , \labels[6].label[58] , 
	\labels[6].label[57] , \labels[6].label[56] , \labels[6].label[55] , 
	\labels[6].label[54] , \labels[6].label[53] , \labels[6].label[52] , 
	\labels[6].label[51] , \labels[6].label[50] , \labels[6].label[49] , 
	\labels[6].label[48] , \labels[6].label[47] , \labels[6].label[46] , 
	\labels[6].label[45] , \labels[6].label[44] , \labels[6].label[43] , 
	\labels[6].label[42] , \labels[6].label[41] , \labels[6].label[40] , 
	\labels[6].label[39] , \labels[6].label[38] , \labels[6].label[37] , 
	\labels[6].label[36] , \labels[6].label[35] , \labels[6].label[34] , 
	\labels[6].label[33] , \labels[6].label[32] , \labels[6].label[31] , 
	\labels[6].label[30] , \labels[6].label[29] , \labels[6].label[28] , 
	\labels[6].label[27] , \labels[6].label[26] , \labels[6].label[25] , 
	\labels[6].label[24] , \labels[6].label[23] , \labels[6].label[22] , 
	\labels[6].label[21] , \labels[6].label[20] , \labels[6].label[19] , 
	\labels[6].label[18] , \labels[6].label[17] , \labels[6].label[16] , 
	\labels[6].label[15] , \labels[6].label[14] , \labels[6].label[13] , 
	\labels[6].label[12] , \labels[6].label[11] , \labels[6].label[10] , 
	\labels[6].label[9] , \labels[6].label[8] , \labels[6].label[7] , 
	\labels[6].label[6] , \labels[6].label[5] , \labels[6].label[4] , 
	\labels[6].label[3] , \labels[6].label[2] , \labels[6].label[1] , 
	\labels[6].label[0] , \labels[6].delimiter_valid[0] , 
	\labels[6].delimiter[7] , \labels[6].delimiter[6] , 
	\labels[6].delimiter[5] , \labels[6].delimiter[4] , 
	\labels[6].delimiter[3] , \labels[6].delimiter[2] , 
	\labels[6].delimiter[1] , \labels[6].delimiter[0] , 
	\labels[5].guid_size[0] , \labels[5].label_size[5] , 
	\labels[5].label_size[4] , \labels[5].label_size[3] , 
	\labels[5].label_size[2] , \labels[5].label_size[1] , 
	\labels[5].label_size[0] , \labels[5].label[255] , 
	\labels[5].label[254] , \labels[5].label[253] , 
	\labels[5].label[252] , \labels[5].label[251] , 
	\labels[5].label[250] , \labels[5].label[249] , 
	\labels[5].label[248] , \labels[5].label[247] , 
	\labels[5].label[246] , \labels[5].label[245] , 
	\labels[5].label[244] , \labels[5].label[243] , 
	\labels[5].label[242] , \labels[5].label[241] , 
	\labels[5].label[240] , \labels[5].label[239] , 
	\labels[5].label[238] , \labels[5].label[237] , 
	\labels[5].label[236] , \labels[5].label[235] , 
	\labels[5].label[234] , \labels[5].label[233] , 
	\labels[5].label[232] , \labels[5].label[231] , 
	\labels[5].label[230] , \labels[5].label[229] , 
	\labels[5].label[228] , \labels[5].label[227] , 
	\labels[5].label[226] , \labels[5].label[225] , 
	\labels[5].label[224] , \labels[5].label[223] , 
	\labels[5].label[222] , \labels[5].label[221] , 
	\labels[5].label[220] , \labels[5].label[219] , 
	\labels[5].label[218] , \labels[5].label[217] , 
	\labels[5].label[216] , \labels[5].label[215] , 
	\labels[5].label[214] , \labels[5].label[213] , 
	\labels[5].label[212] , \labels[5].label[211] , 
	\labels[5].label[210] , \labels[5].label[209] , 
	\labels[5].label[208] , \labels[5].label[207] , 
	\labels[5].label[206] , \labels[5].label[205] , 
	\labels[5].label[204] , \labels[5].label[203] , 
	\labels[5].label[202] , \labels[5].label[201] , 
	\labels[5].label[200] , \labels[5].label[199] , 
	\labels[5].label[198] , \labels[5].label[197] , 
	\labels[5].label[196] , \labels[5].label[195] , 
	\labels[5].label[194] , \labels[5].label[193] , 
	\labels[5].label[192] , \labels[5].label[191] , 
	\labels[5].label[190] , \labels[5].label[189] , 
	\labels[5].label[188] , \labels[5].label[187] , 
	\labels[5].label[186] , \labels[5].label[185] , 
	\labels[5].label[184] , \labels[5].label[183] , 
	\labels[5].label[182] , \labels[5].label[181] , 
	\labels[5].label[180] , \labels[5].label[179] , 
	\labels[5].label[178] , \labels[5].label[177] , 
	\labels[5].label[176] , \labels[5].label[175] , 
	\labels[5].label[174] , \labels[5].label[173] , 
	\labels[5].label[172] , \labels[5].label[171] , 
	\labels[5].label[170] , \labels[5].label[169] , 
	\labels[5].label[168] , \labels[5].label[167] , 
	\labels[5].label[166] , \labels[5].label[165] , 
	\labels[5].label[164] , \labels[5].label[163] , 
	\labels[5].label[162] , \labels[5].label[161] , 
	\labels[5].label[160] , \labels[5].label[159] , 
	\labels[5].label[158] , \labels[5].label[157] , 
	\labels[5].label[156] , \labels[5].label[155] , 
	\labels[5].label[154] , \labels[5].label[153] , 
	\labels[5].label[152] , \labels[5].label[151] , 
	\labels[5].label[150] , \labels[5].label[149] , 
	\labels[5].label[148] , \labels[5].label[147] , 
	\labels[5].label[146] , \labels[5].label[145] , 
	\labels[5].label[144] , \labels[5].label[143] , 
	\labels[5].label[142] , \labels[5].label[141] , 
	\labels[5].label[140] , \labels[5].label[139] , 
	\labels[5].label[138] , \labels[5].label[137] , 
	\labels[5].label[136] , \labels[5].label[135] , 
	\labels[5].label[134] , \labels[5].label[133] , 
	\labels[5].label[132] , \labels[5].label[131] , 
	\labels[5].label[130] , \labels[5].label[129] , 
	\labels[5].label[128] , \labels[5].label[127] , 
	\labels[5].label[126] , \labels[5].label[125] , 
	\labels[5].label[124] , \labels[5].label[123] , 
	\labels[5].label[122] , \labels[5].label[121] , 
	\labels[5].label[120] , \labels[5].label[119] , 
	\labels[5].label[118] , \labels[5].label[117] , 
	\labels[5].label[116] , \labels[5].label[115] , 
	\labels[5].label[114] , \labels[5].label[113] , 
	\labels[5].label[112] , \labels[5].label[111] , 
	\labels[5].label[110] , \labels[5].label[109] , 
	\labels[5].label[108] , \labels[5].label[107] , 
	\labels[5].label[106] , \labels[5].label[105] , 
	\labels[5].label[104] , \labels[5].label[103] , 
	\labels[5].label[102] , \labels[5].label[101] , 
	\labels[5].label[100] , \labels[5].label[99] , \labels[5].label[98] , 
	\labels[5].label[97] , \labels[5].label[96] , \labels[5].label[95] , 
	\labels[5].label[94] , \labels[5].label[93] , \labels[5].label[92] , 
	\labels[5].label[91] , \labels[5].label[90] , \labels[5].label[89] , 
	\labels[5].label[88] , \labels[5].label[87] , \labels[5].label[86] , 
	\labels[5].label[85] , \labels[5].label[84] , \labels[5].label[83] , 
	\labels[5].label[82] , \labels[5].label[81] , \labels[5].label[80] , 
	\labels[5].label[79] , \labels[5].label[78] , \labels[5].label[77] , 
	\labels[5].label[76] , \labels[5].label[75] , \labels[5].label[74] , 
	\labels[5].label[73] , \labels[5].label[72] , \labels[5].label[71] , 
	\labels[5].label[70] , \labels[5].label[69] , \labels[5].label[68] , 
	\labels[5].label[67] , \labels[5].label[66] , \labels[5].label[65] , 
	\labels[5].label[64] , \labels[5].label[63] , \labels[5].label[62] , 
	\labels[5].label[61] , \labels[5].label[60] , \labels[5].label[59] , 
	\labels[5].label[58] , \labels[5].label[57] , \labels[5].label[56] , 
	\labels[5].label[55] , \labels[5].label[54] , \labels[5].label[53] , 
	\labels[5].label[52] , \labels[5].label[51] , \labels[5].label[50] , 
	\labels[5].label[49] , \labels[5].label[48] , \labels[5].label[47] , 
	\labels[5].label[46] , \labels[5].label[45] , \labels[5].label[44] , 
	\labels[5].label[43] , \labels[5].label[42] , \labels[5].label[41] , 
	\labels[5].label[40] , \labels[5].label[39] , \labels[5].label[38] , 
	\labels[5].label[37] , \labels[5].label[36] , \labels[5].label[35] , 
	\labels[5].label[34] , \labels[5].label[33] , \labels[5].label[32] , 
	\labels[5].label[31] , \labels[5].label[30] , \labels[5].label[29] , 
	\labels[5].label[28] , \labels[5].label[27] , \labels[5].label[26] , 
	\labels[5].label[25] , \labels[5].label[24] , \labels[5].label[23] , 
	\labels[5].label[22] , \labels[5].label[21] , \labels[5].label[20] , 
	\labels[5].label[19] , \labels[5].label[18] , \labels[5].label[17] , 
	\labels[5].label[16] , \labels[5].label[15] , \labels[5].label[14] , 
	\labels[5].label[13] , \labels[5].label[12] , \labels[5].label[11] , 
	\labels[5].label[10] , \labels[5].label[9] , \labels[5].label[8] , 
	\labels[5].label[7] , \labels[5].label[6] , \labels[5].label[5] , 
	\labels[5].label[4] , \labels[5].label[3] , \labels[5].label[2] , 
	\labels[5].label[1] , \labels[5].label[0] , 
	\labels[5].delimiter_valid[0] , \labels[5].delimiter[7] , 
	\labels[5].delimiter[6] , \labels[5].delimiter[5] , 
	\labels[5].delimiter[4] , \labels[5].delimiter[3] , 
	\labels[5].delimiter[2] , \labels[5].delimiter[1] , 
	\labels[5].delimiter[0] , \labels[4].guid_size[0] , 
	\labels[4].label_size[5] , \labels[4].label_size[4] , 
	\labels[4].label_size[3] , \labels[4].label_size[2] , 
	\labels[4].label_size[1] , \labels[4].label_size[0] , 
	\labels[4].label[255] , \labels[4].label[254] , 
	\labels[4].label[253] , \labels[4].label[252] , 
	\labels[4].label[251] , \labels[4].label[250] , 
	\labels[4].label[249] , \labels[4].label[248] , 
	\labels[4].label[247] , \labels[4].label[246] , 
	\labels[4].label[245] , \labels[4].label[244] , 
	\labels[4].label[243] , \labels[4].label[242] , 
	\labels[4].label[241] , \labels[4].label[240] , 
	\labels[4].label[239] , \labels[4].label[238] , 
	\labels[4].label[237] , \labels[4].label[236] , 
	\labels[4].label[235] , \labels[4].label[234] , 
	\labels[4].label[233] , \labels[4].label[232] , 
	\labels[4].label[231] , \labels[4].label[230] , 
	\labels[4].label[229] , \labels[4].label[228] , 
	\labels[4].label[227] , \labels[4].label[226] , 
	\labels[4].label[225] , \labels[4].label[224] , 
	\labels[4].label[223] , \labels[4].label[222] , 
	\labels[4].label[221] , \labels[4].label[220] , 
	\labels[4].label[219] , \labels[4].label[218] , 
	\labels[4].label[217] , \labels[4].label[216] , 
	\labels[4].label[215] , \labels[4].label[214] , 
	\labels[4].label[213] , \labels[4].label[212] , 
	\labels[4].label[211] , \labels[4].label[210] , 
	\labels[4].label[209] , \labels[4].label[208] , 
	\labels[4].label[207] , \labels[4].label[206] , 
	\labels[4].label[205] , \labels[4].label[204] , 
	\labels[4].label[203] , \labels[4].label[202] , 
	\labels[4].label[201] , \labels[4].label[200] , 
	\labels[4].label[199] , \labels[4].label[198] , 
	\labels[4].label[197] , \labels[4].label[196] , 
	\labels[4].label[195] , \labels[4].label[194] , 
	\labels[4].label[193] , \labels[4].label[192] , 
	\labels[4].label[191] , \labels[4].label[190] , 
	\labels[4].label[189] , \labels[4].label[188] , 
	\labels[4].label[187] , \labels[4].label[186] , 
	\labels[4].label[185] , \labels[4].label[184] , 
	\labels[4].label[183] , \labels[4].label[182] , 
	\labels[4].label[181] , \labels[4].label[180] , 
	\labels[4].label[179] , \labels[4].label[178] , 
	\labels[4].label[177] , \labels[4].label[176] , 
	\labels[4].label[175] , \labels[4].label[174] , 
	\labels[4].label[173] , \labels[4].label[172] , 
	\labels[4].label[171] , \labels[4].label[170] , 
	\labels[4].label[169] , \labels[4].label[168] , 
	\labels[4].label[167] , \labels[4].label[166] , 
	\labels[4].label[165] , \labels[4].label[164] , 
	\labels[4].label[163] , \labels[4].label[162] , 
	\labels[4].label[161] , \labels[4].label[160] , 
	\labels[4].label[159] , \labels[4].label[158] , 
	\labels[4].label[157] , \labels[4].label[156] , 
	\labels[4].label[155] , \labels[4].label[154] , 
	\labels[4].label[153] , \labels[4].label[152] , 
	\labels[4].label[151] , \labels[4].label[150] , 
	\labels[4].label[149] , \labels[4].label[148] , 
	\labels[4].label[147] , \labels[4].label[146] , 
	\labels[4].label[145] , \labels[4].label[144] , 
	\labels[4].label[143] , \labels[4].label[142] , 
	\labels[4].label[141] , \labels[4].label[140] , 
	\labels[4].label[139] , \labels[4].label[138] , 
	\labels[4].label[137] , \labels[4].label[136] , 
	\labels[4].label[135] , \labels[4].label[134] , 
	\labels[4].label[133] , \labels[4].label[132] , 
	\labels[4].label[131] , \labels[4].label[130] , 
	\labels[4].label[129] , \labels[4].label[128] , 
	\labels[4].label[127] , \labels[4].label[126] , 
	\labels[4].label[125] , \labels[4].label[124] , 
	\labels[4].label[123] , \labels[4].label[122] , 
	\labels[4].label[121] , \labels[4].label[120] , 
	\labels[4].label[119] , \labels[4].label[118] , 
	\labels[4].label[117] , \labels[4].label[116] , 
	\labels[4].label[115] , \labels[4].label[114] , 
	\labels[4].label[113] , \labels[4].label[112] , 
	\labels[4].label[111] , \labels[4].label[110] , 
	\labels[4].label[109] , \labels[4].label[108] , 
	\labels[4].label[107] , \labels[4].label[106] , 
	\labels[4].label[105] , \labels[4].label[104] , 
	\labels[4].label[103] , \labels[4].label[102] , 
	\labels[4].label[101] , \labels[4].label[100] , 
	\labels[4].label[99] , \labels[4].label[98] , \labels[4].label[97] , 
	\labels[4].label[96] , \labels[4].label[95] , \labels[4].label[94] , 
	\labels[4].label[93] , \labels[4].label[92] , \labels[4].label[91] , 
	\labels[4].label[90] , \labels[4].label[89] , \labels[4].label[88] , 
	\labels[4].label[87] , \labels[4].label[86] , \labels[4].label[85] , 
	\labels[4].label[84] , \labels[4].label[83] , \labels[4].label[82] , 
	\labels[4].label[81] , \labels[4].label[80] , \labels[4].label[79] , 
	\labels[4].label[78] , \labels[4].label[77] , \labels[4].label[76] , 
	\labels[4].label[75] , \labels[4].label[74] , \labels[4].label[73] , 
	\labels[4].label[72] , \labels[4].label[71] , \labels[4].label[70] , 
	\labels[4].label[69] , \labels[4].label[68] , \labels[4].label[67] , 
	\labels[4].label[66] , \labels[4].label[65] , \labels[4].label[64] , 
	\labels[4].label[63] , \labels[4].label[62] , \labels[4].label[61] , 
	\labels[4].label[60] , \labels[4].label[59] , \labels[4].label[58] , 
	\labels[4].label[57] , \labels[4].label[56] , \labels[4].label[55] , 
	\labels[4].label[54] , \labels[4].label[53] , \labels[4].label[52] , 
	\labels[4].label[51] , \labels[4].label[50] , \labels[4].label[49] , 
	\labels[4].label[48] , \labels[4].label[47] , \labels[4].label[46] , 
	\labels[4].label[45] , \labels[4].label[44] , \labels[4].label[43] , 
	\labels[4].label[42] , \labels[4].label[41] , \labels[4].label[40] , 
	\labels[4].label[39] , \labels[4].label[38] , \labels[4].label[37] , 
	\labels[4].label[36] , \labels[4].label[35] , \labels[4].label[34] , 
	\labels[4].label[33] , \labels[4].label[32] , \labels[4].label[31] , 
	\labels[4].label[30] , \labels[4].label[29] , \labels[4].label[28] , 
	\labels[4].label[27] , \labels[4].label[26] , \labels[4].label[25] , 
	\labels[4].label[24] , \labels[4].label[23] , \labels[4].label[22] , 
	\labels[4].label[21] , \labels[4].label[20] , \labels[4].label[19] , 
	\labels[4].label[18] , \labels[4].label[17] , \labels[4].label[16] , 
	\labels[4].label[15] , \labels[4].label[14] , \labels[4].label[13] , 
	\labels[4].label[12] , \labels[4].label[11] , \labels[4].label[10] , 
	\labels[4].label[9] , \labels[4].label[8] , \labels[4].label[7] , 
	\labels[4].label[6] , \labels[4].label[5] , \labels[4].label[4] , 
	\labels[4].label[3] , \labels[4].label[2] , \labels[4].label[1] , 
	\labels[4].label[0] , \labels[4].delimiter_valid[0] , 
	\labels[4].delimiter[7] , \labels[4].delimiter[6] , 
	\labels[4].delimiter[5] , \labels[4].delimiter[4] , 
	\labels[4].delimiter[3] , \labels[4].delimiter[2] , 
	\labels[4].delimiter[1] , \labels[4].delimiter[0] , 
	\labels[3].guid_size[0] , \labels[3].label_size[5] , 
	\labels[3].label_size[4] , \labels[3].label_size[3] , 
	\labels[3].label_size[2] , \labels[3].label_size[1] , 
	\labels[3].label_size[0] , \labels[3].label[255] , 
	\labels[3].label[254] , \labels[3].label[253] , 
	\labels[3].label[252] , \labels[3].label[251] , 
	\labels[3].label[250] , \labels[3].label[249] , 
	\labels[3].label[248] , \labels[3].label[247] , 
	\labels[3].label[246] , \labels[3].label[245] , 
	\labels[3].label[244] , \labels[3].label[243] , 
	\labels[3].label[242] , \labels[3].label[241] , 
	\labels[3].label[240] , \labels[3].label[239] , 
	\labels[3].label[238] , \labels[3].label[237] , 
	\labels[3].label[236] , \labels[3].label[235] , 
	\labels[3].label[234] , \labels[3].label[233] , 
	\labels[3].label[232] , \labels[3].label[231] , 
	\labels[3].label[230] , \labels[3].label[229] , 
	\labels[3].label[228] , \labels[3].label[227] , 
	\labels[3].label[226] , \labels[3].label[225] , 
	\labels[3].label[224] , \labels[3].label[223] , 
	\labels[3].label[222] , \labels[3].label[221] , 
	\labels[3].label[220] , \labels[3].label[219] , 
	\labels[3].label[218] , \labels[3].label[217] , 
	\labels[3].label[216] , \labels[3].label[215] , 
	\labels[3].label[214] , \labels[3].label[213] , 
	\labels[3].label[212] , \labels[3].label[211] , 
	\labels[3].label[210] , \labels[3].label[209] , 
	\labels[3].label[208] , \labels[3].label[207] , 
	\labels[3].label[206] , \labels[3].label[205] , 
	\labels[3].label[204] , \labels[3].label[203] , 
	\labels[3].label[202] , \labels[3].label[201] , 
	\labels[3].label[200] , \labels[3].label[199] , 
	\labels[3].label[198] , \labels[3].label[197] , 
	\labels[3].label[196] , \labels[3].label[195] , 
	\labels[3].label[194] , \labels[3].label[193] , 
	\labels[3].label[192] , \labels[3].label[191] , 
	\labels[3].label[190] , \labels[3].label[189] , 
	\labels[3].label[188] , \labels[3].label[187] , 
	\labels[3].label[186] , \labels[3].label[185] , 
	\labels[3].label[184] , \labels[3].label[183] , 
	\labels[3].label[182] , \labels[3].label[181] , 
	\labels[3].label[180] , \labels[3].label[179] , 
	\labels[3].label[178] , \labels[3].label[177] , 
	\labels[3].label[176] , \labels[3].label[175] , 
	\labels[3].label[174] , \labels[3].label[173] , 
	\labels[3].label[172] , \labels[3].label[171] , 
	\labels[3].label[170] , \labels[3].label[169] , 
	\labels[3].label[168] , \labels[3].label[167] , 
	\labels[3].label[166] , \labels[3].label[165] , 
	\labels[3].label[164] , \labels[3].label[163] , 
	\labels[3].label[162] , \labels[3].label[161] , 
	\labels[3].label[160] , \labels[3].label[159] , 
	\labels[3].label[158] , \labels[3].label[157] , 
	\labels[3].label[156] , \labels[3].label[155] , 
	\labels[3].label[154] , \labels[3].label[153] , 
	\labels[3].label[152] , \labels[3].label[151] , 
	\labels[3].label[150] , \labels[3].label[149] , 
	\labels[3].label[148] , \labels[3].label[147] , 
	\labels[3].label[146] , \labels[3].label[145] , 
	\labels[3].label[144] , \labels[3].label[143] , 
	\labels[3].label[142] , \labels[3].label[141] , 
	\labels[3].label[140] , \labels[3].label[139] , 
	\labels[3].label[138] , \labels[3].label[137] , 
	\labels[3].label[136] , \labels[3].label[135] , 
	\labels[3].label[134] , \labels[3].label[133] , 
	\labels[3].label[132] , \labels[3].label[131] , 
	\labels[3].label[130] , \labels[3].label[129] , 
	\labels[3].label[128] , \labels[3].label[127] , 
	\labels[3].label[126] , \labels[3].label[125] , 
	\labels[3].label[124] , \labels[3].label[123] , 
	\labels[3].label[122] , \labels[3].label[121] , 
	\labels[3].label[120] , \labels[3].label[119] , 
	\labels[3].label[118] , \labels[3].label[117] , 
	\labels[3].label[116] , \labels[3].label[115] , 
	\labels[3].label[114] , \labels[3].label[113] , 
	\labels[3].label[112] , \labels[3].label[111] , 
	\labels[3].label[110] , \labels[3].label[109] , 
	\labels[3].label[108] , \labels[3].label[107] , 
	\labels[3].label[106] , \labels[3].label[105] , 
	\labels[3].label[104] , \labels[3].label[103] , 
	\labels[3].label[102] , \labels[3].label[101] , 
	\labels[3].label[100] , \labels[3].label[99] , \labels[3].label[98] , 
	\labels[3].label[97] , \labels[3].label[96] , \labels[3].label[95] , 
	\labels[3].label[94] , \labels[3].label[93] , \labels[3].label[92] , 
	\labels[3].label[91] , \labels[3].label[90] , \labels[3].label[89] , 
	\labels[3].label[88] , \labels[3].label[87] , \labels[3].label[86] , 
	\labels[3].label[85] , \labels[3].label[84] , \labels[3].label[83] , 
	\labels[3].label[82] , \labels[3].label[81] , \labels[3].label[80] , 
	\labels[3].label[79] , \labels[3].label[78] , \labels[3].label[77] , 
	\labels[3].label[76] , \labels[3].label[75] , \labels[3].label[74] , 
	\labels[3].label[73] , \labels[3].label[72] , \labels[3].label[71] , 
	\labels[3].label[70] , \labels[3].label[69] , \labels[3].label[68] , 
	\labels[3].label[67] , \labels[3].label[66] , \labels[3].label[65] , 
	\labels[3].label[64] , \labels[3].label[63] , \labels[3].label[62] , 
	\labels[3].label[61] , \labels[3].label[60] , \labels[3].label[59] , 
	\labels[3].label[58] , \labels[3].label[57] , \labels[3].label[56] , 
	\labels[3].label[55] , \labels[3].label[54] , \labels[3].label[53] , 
	\labels[3].label[52] , \labels[3].label[51] , \labels[3].label[50] , 
	\labels[3].label[49] , \labels[3].label[48] , \labels[3].label[47] , 
	\labels[3].label[46] , \labels[3].label[45] , \labels[3].label[44] , 
	\labels[3].label[43] , \labels[3].label[42] , \labels[3].label[41] , 
	\labels[3].label[40] , \labels[3].label[39] , \labels[3].label[38] , 
	\labels[3].label[37] , \labels[3].label[36] , \labels[3].label[35] , 
	\labels[3].label[34] , \labels[3].label[33] , \labels[3].label[32] , 
	\labels[3].label[31] , \labels[3].label[30] , \labels[3].label[29] , 
	\labels[3].label[28] , \labels[3].label[27] , \labels[3].label[26] , 
	\labels[3].label[25] , \labels[3].label[24] , \labels[3].label[23] , 
	\labels[3].label[22] , \labels[3].label[21] , \labels[3].label[20] , 
	\labels[3].label[19] , \labels[3].label[18] , \labels[3].label[17] , 
	\labels[3].label[16] , \labels[3].label[15] , \labels[3].label[14] , 
	\labels[3].label[13] , \labels[3].label[12] , \labels[3].label[11] , 
	\labels[3].label[10] , \labels[3].label[9] , \labels[3].label[8] , 
	\labels[3].label[7] , \labels[3].label[6] , \labels[3].label[5] , 
	\labels[3].label[4] , \labels[3].label[3] , \labels[3].label[2] , 
	\labels[3].label[1] , \labels[3].label[0] , 
	\labels[3].delimiter_valid[0] , \labels[3].delimiter[7] , 
	\labels[3].delimiter[6] , \labels[3].delimiter[5] , 
	\labels[3].delimiter[4] , \labels[3].delimiter[3] , 
	\labels[3].delimiter[2] , \labels[3].delimiter[1] , 
	\labels[3].delimiter[0] , \labels[2].guid_size[0] , 
	\labels[2].label_size[5] , \labels[2].label_size[4] , 
	\labels[2].label_size[3] , \labels[2].label_size[2] , 
	\labels[2].label_size[1] , \labels[2].label_size[0] , 
	\labels[2].label[255] , \labels[2].label[254] , 
	\labels[2].label[253] , \labels[2].label[252] , 
	\labels[2].label[251] , \labels[2].label[250] , 
	\labels[2].label[249] , \labels[2].label[248] , 
	\labels[2].label[247] , \labels[2].label[246] , 
	\labels[2].label[245] , \labels[2].label[244] , 
	\labels[2].label[243] , \labels[2].label[242] , 
	\labels[2].label[241] , \labels[2].label[240] , 
	\labels[2].label[239] , \labels[2].label[238] , 
	\labels[2].label[237] , \labels[2].label[236] , 
	\labels[2].label[235] , \labels[2].label[234] , 
	\labels[2].label[233] , \labels[2].label[232] , 
	\labels[2].label[231] , \labels[2].label[230] , 
	\labels[2].label[229] , \labels[2].label[228] , 
	\labels[2].label[227] , \labels[2].label[226] , 
	\labels[2].label[225] , \labels[2].label[224] , 
	\labels[2].label[223] , \labels[2].label[222] , 
	\labels[2].label[221] , \labels[2].label[220] , 
	\labels[2].label[219] , \labels[2].label[218] , 
	\labels[2].label[217] , \labels[2].label[216] , 
	\labels[2].label[215] , \labels[2].label[214] , 
	\labels[2].label[213] , \labels[2].label[212] , 
	\labels[2].label[211] , \labels[2].label[210] , 
	\labels[2].label[209] , \labels[2].label[208] , 
	\labels[2].label[207] , \labels[2].label[206] , 
	\labels[2].label[205] , \labels[2].label[204] , 
	\labels[2].label[203] , \labels[2].label[202] , 
	\labels[2].label[201] , \labels[2].label[200] , 
	\labels[2].label[199] , \labels[2].label[198] , 
	\labels[2].label[197] , \labels[2].label[196] , 
	\labels[2].label[195] , \labels[2].label[194] , 
	\labels[2].label[193] , \labels[2].label[192] , 
	\labels[2].label[191] , \labels[2].label[190] , 
	\labels[2].label[189] , \labels[2].label[188] , 
	\labels[2].label[187] , \labels[2].label[186] , 
	\labels[2].label[185] , \labels[2].label[184] , 
	\labels[2].label[183] , \labels[2].label[182] , 
	\labels[2].label[181] , \labels[2].label[180] , 
	\labels[2].label[179] , \labels[2].label[178] , 
	\labels[2].label[177] , \labels[2].label[176] , 
	\labels[2].label[175] , \labels[2].label[174] , 
	\labels[2].label[173] , \labels[2].label[172] , 
	\labels[2].label[171] , \labels[2].label[170] , 
	\labels[2].label[169] , \labels[2].label[168] , 
	\labels[2].label[167] , \labels[2].label[166] , 
	\labels[2].label[165] , \labels[2].label[164] , 
	\labels[2].label[163] , \labels[2].label[162] , 
	\labels[2].label[161] , \labels[2].label[160] , 
	\labels[2].label[159] , \labels[2].label[158] , 
	\labels[2].label[157] , \labels[2].label[156] , 
	\labels[2].label[155] , \labels[2].label[154] , 
	\labels[2].label[153] , \labels[2].label[152] , 
	\labels[2].label[151] , \labels[2].label[150] , 
	\labels[2].label[149] , \labels[2].label[148] , 
	\labels[2].label[147] , \labels[2].label[146] , 
	\labels[2].label[145] , \labels[2].label[144] , 
	\labels[2].label[143] , \labels[2].label[142] , 
	\labels[2].label[141] , \labels[2].label[140] , 
	\labels[2].label[139] , \labels[2].label[138] , 
	\labels[2].label[137] , \labels[2].label[136] , 
	\labels[2].label[135] , \labels[2].label[134] , 
	\labels[2].label[133] , \labels[2].label[132] , 
	\labels[2].label[131] , \labels[2].label[130] , 
	\labels[2].label[129] , \labels[2].label[128] , 
	\labels[2].label[127] , \labels[2].label[126] , 
	\labels[2].label[125] , \labels[2].label[124] , 
	\labels[2].label[123] , \labels[2].label[122] , 
	\labels[2].label[121] , \labels[2].label[120] , 
	\labels[2].label[119] , \labels[2].label[118] , 
	\labels[2].label[117] , \labels[2].label[116] , 
	\labels[2].label[115] , \labels[2].label[114] , 
	\labels[2].label[113] , \labels[2].label[112] , 
	\labels[2].label[111] , \labels[2].label[110] , 
	\labels[2].label[109] , \labels[2].label[108] , 
	\labels[2].label[107] , \labels[2].label[106] , 
	\labels[2].label[105] , \labels[2].label[104] , 
	\labels[2].label[103] , \labels[2].label[102] , 
	\labels[2].label[101] , \labels[2].label[100] , 
	\labels[2].label[99] , \labels[2].label[98] , \labels[2].label[97] , 
	\labels[2].label[96] , \labels[2].label[95] , \labels[2].label[94] , 
	\labels[2].label[93] , \labels[2].label[92] , \labels[2].label[91] , 
	\labels[2].label[90] , \labels[2].label[89] , \labels[2].label[88] , 
	\labels[2].label[87] , \labels[2].label[86] , \labels[2].label[85] , 
	\labels[2].label[84] , \labels[2].label[83] , \labels[2].label[82] , 
	\labels[2].label[81] , \labels[2].label[80] , \labels[2].label[79] , 
	\labels[2].label[78] , \labels[2].label[77] , \labels[2].label[76] , 
	\labels[2].label[75] , \labels[2].label[74] , \labels[2].label[73] , 
	\labels[2].label[72] , \labels[2].label[71] , \labels[2].label[70] , 
	\labels[2].label[69] , \labels[2].label[68] , \labels[2].label[67] , 
	\labels[2].label[66] , \labels[2].label[65] , \labels[2].label[64] , 
	\labels[2].label[63] , \labels[2].label[62] , \labels[2].label[61] , 
	\labels[2].label[60] , \labels[2].label[59] , \labels[2].label[58] , 
	\labels[2].label[57] , \labels[2].label[56] , \labels[2].label[55] , 
	\labels[2].label[54] , \labels[2].label[53] , \labels[2].label[52] , 
	\labels[2].label[51] , \labels[2].label[50] , \labels[2].label[49] , 
	\labels[2].label[48] , \labels[2].label[47] , \labels[2].label[46] , 
	\labels[2].label[45] , \labels[2].label[44] , \labels[2].label[43] , 
	\labels[2].label[42] , \labels[2].label[41] , \labels[2].label[40] , 
	\labels[2].label[39] , \labels[2].label[38] , \labels[2].label[37] , 
	\labels[2].label[36] , \labels[2].label[35] , \labels[2].label[34] , 
	\labels[2].label[33] , \labels[2].label[32] , \labels[2].label[31] , 
	\labels[2].label[30] , \labels[2].label[29] , \labels[2].label[28] , 
	\labels[2].label[27] , \labels[2].label[26] , \labels[2].label[25] , 
	\labels[2].label[24] , \labels[2].label[23] , \labels[2].label[22] , 
	\labels[2].label[21] , \labels[2].label[20] , \labels[2].label[19] , 
	\labels[2].label[18] , \labels[2].label[17] , \labels[2].label[16] , 
	\labels[2].label[15] , \labels[2].label[14] , \labels[2].label[13] , 
	\labels[2].label[12] , \labels[2].label[11] , \labels[2].label[10] , 
	\labels[2].label[9] , \labels[2].label[8] , \labels[2].label[7] , 
	\labels[2].label[6] , \labels[2].label[5] , \labels[2].label[4] , 
	\labels[2].label[3] , \labels[2].label[2] , \labels[2].label[1] , 
	\labels[2].label[0] , \labels[2].delimiter_valid[0] , 
	\labels[2].delimiter[7] , \labels[2].delimiter[6] , 
	\labels[2].delimiter[5] , \labels[2].delimiter[4] , 
	\labels[2].delimiter[3] , \labels[2].delimiter[2] , 
	\labels[2].delimiter[1] , \labels[2].delimiter[0] , 
	\labels[1].guid_size[0] , \labels[1].label_size[5] , 
	\labels[1].label_size[4] , \labels[1].label_size[3] , 
	\labels[1].label_size[2] , \labels[1].label_size[1] , 
	\labels[1].label_size[0] , \labels[1].label[255] , 
	\labels[1].label[254] , \labels[1].label[253] , 
	\labels[1].label[252] , \labels[1].label[251] , 
	\labels[1].label[250] , \labels[1].label[249] , 
	\labels[1].label[248] , \labels[1].label[247] , 
	\labels[1].label[246] , \labels[1].label[245] , 
	\labels[1].label[244] , \labels[1].label[243] , 
	\labels[1].label[242] , \labels[1].label[241] , 
	\labels[1].label[240] , \labels[1].label[239] , 
	\labels[1].label[238] , \labels[1].label[237] , 
	\labels[1].label[236] , \labels[1].label[235] , 
	\labels[1].label[234] , \labels[1].label[233] , 
	\labels[1].label[232] , \labels[1].label[231] , 
	\labels[1].label[230] , \labels[1].label[229] , 
	\labels[1].label[228] , \labels[1].label[227] , 
	\labels[1].label[226] , \labels[1].label[225] , 
	\labels[1].label[224] , \labels[1].label[223] , 
	\labels[1].label[222] , \labels[1].label[221] , 
	\labels[1].label[220] , \labels[1].label[219] , 
	\labels[1].label[218] , \labels[1].label[217] , 
	\labels[1].label[216] , \labels[1].label[215] , 
	\labels[1].label[214] , \labels[1].label[213] , 
	\labels[1].label[212] , \labels[1].label[211] , 
	\labels[1].label[210] , \labels[1].label[209] , 
	\labels[1].label[208] , \labels[1].label[207] , 
	\labels[1].label[206] , \labels[1].label[205] , 
	\labels[1].label[204] , \labels[1].label[203] , 
	\labels[1].label[202] , \labels[1].label[201] , 
	\labels[1].label[200] , \labels[1].label[199] , 
	\labels[1].label[198] , \labels[1].label[197] , 
	\labels[1].label[196] , \labels[1].label[195] , 
	\labels[1].label[194] , \labels[1].label[193] , 
	\labels[1].label[192] , \labels[1].label[191] , 
	\labels[1].label[190] , \labels[1].label[189] , 
	\labels[1].label[188] , \labels[1].label[187] , 
	\labels[1].label[186] , \labels[1].label[185] , 
	\labels[1].label[184] , \labels[1].label[183] , 
	\labels[1].label[182] , \labels[1].label[181] , 
	\labels[1].label[180] , \labels[1].label[179] , 
	\labels[1].label[178] , \labels[1].label[177] , 
	\labels[1].label[176] , \labels[1].label[175] , 
	\labels[1].label[174] , \labels[1].label[173] , 
	\labels[1].label[172] , \labels[1].label[171] , 
	\labels[1].label[170] , \labels[1].label[169] , 
	\labels[1].label[168] , \labels[1].label[167] , 
	\labels[1].label[166] , \labels[1].label[165] , 
	\labels[1].label[164] , \labels[1].label[163] , 
	\labels[1].label[162] , \labels[1].label[161] , 
	\labels[1].label[160] , \labels[1].label[159] , 
	\labels[1].label[158] , \labels[1].label[157] , 
	\labels[1].label[156] , \labels[1].label[155] , 
	\labels[1].label[154] , \labels[1].label[153] , 
	\labels[1].label[152] , \labels[1].label[151] , 
	\labels[1].label[150] , \labels[1].label[149] , 
	\labels[1].label[148] , \labels[1].label[147] , 
	\labels[1].label[146] , \labels[1].label[145] , 
	\labels[1].label[144] , \labels[1].label[143] , 
	\labels[1].label[142] , \labels[1].label[141] , 
	\labels[1].label[140] , \labels[1].label[139] , 
	\labels[1].label[138] , \labels[1].label[137] , 
	\labels[1].label[136] , \labels[1].label[135] , 
	\labels[1].label[134] , \labels[1].label[133] , 
	\labels[1].label[132] , \labels[1].label[131] , 
	\labels[1].label[130] , \labels[1].label[129] , 
	\labels[1].label[128] , \labels[1].label[127] , 
	\labels[1].label[126] , \labels[1].label[125] , 
	\labels[1].label[124] , \labels[1].label[123] , 
	\labels[1].label[122] , \labels[1].label[121] , 
	\labels[1].label[120] , \labels[1].label[119] , 
	\labels[1].label[118] , \labels[1].label[117] , 
	\labels[1].label[116] , \labels[1].label[115] , 
	\labels[1].label[114] , \labels[1].label[113] , 
	\labels[1].label[112] , \labels[1].label[111] , 
	\labels[1].label[110] , \labels[1].label[109] , 
	\labels[1].label[108] , \labels[1].label[107] , 
	\labels[1].label[106] , \labels[1].label[105] , 
	\labels[1].label[104] , \labels[1].label[103] , 
	\labels[1].label[102] , \labels[1].label[101] , 
	\labels[1].label[100] , \labels[1].label[99] , \labels[1].label[98] , 
	\labels[1].label[97] , \labels[1].label[96] , \labels[1].label[95] , 
	\labels[1].label[94] , \labels[1].label[93] , \labels[1].label[92] , 
	\labels[1].label[91] , \labels[1].label[90] , \labels[1].label[89] , 
	\labels[1].label[88] , \labels[1].label[87] , \labels[1].label[86] , 
	\labels[1].label[85] , \labels[1].label[84] , \labels[1].label[83] , 
	\labels[1].label[82] , \labels[1].label[81] , \labels[1].label[80] , 
	\labels[1].label[79] , \labels[1].label[78] , \labels[1].label[77] , 
	\labels[1].label[76] , \labels[1].label[75] , \labels[1].label[74] , 
	\labels[1].label[73] , \labels[1].label[72] , \labels[1].label[71] , 
	\labels[1].label[70] , \labels[1].label[69] , \labels[1].label[68] , 
	\labels[1].label[67] , \labels[1].label[66] , \labels[1].label[65] , 
	\labels[1].label[64] , \labels[1].label[63] , \labels[1].label[62] , 
	\labels[1].label[61] , \labels[1].label[60] , \labels[1].label[59] , 
	\labels[1].label[58] , \labels[1].label[57] , \labels[1].label[56] , 
	\labels[1].label[55] , \labels[1].label[54] , \labels[1].label[53] , 
	\labels[1].label[52] , \labels[1].label[51] , \labels[1].label[50] , 
	\labels[1].label[49] , \labels[1].label[48] , \labels[1].label[47] , 
	\labels[1].label[46] , \labels[1].label[45] , \labels[1].label[44] , 
	\labels[1].label[43] , \labels[1].label[42] , \labels[1].label[41] , 
	\labels[1].label[40] , \labels[1].label[39] , \labels[1].label[38] , 
	\labels[1].label[37] , \labels[1].label[36] , \labels[1].label[35] , 
	\labels[1].label[34] , \labels[1].label[33] , \labels[1].label[32] , 
	\labels[1].label[31] , \labels[1].label[30] , \labels[1].label[29] , 
	\labels[1].label[28] , \labels[1].label[27] , \labels[1].label[26] , 
	\labels[1].label[25] , \labels[1].label[24] , \labels[1].label[23] , 
	\labels[1].label[22] , \labels[1].label[21] , \labels[1].label[20] , 
	\labels[1].label[19] , \labels[1].label[18] , \labels[1].label[17] , 
	\labels[1].label[16] , \labels[1].label[15] , \labels[1].label[14] , 
	\labels[1].label[13] , \labels[1].label[12] , \labels[1].label[11] , 
	\labels[1].label[10] , \labels[1].label[9] , \labels[1].label[8] , 
	\labels[1].label[7] , \labels[1].label[6] , \labels[1].label[5] , 
	\labels[1].label[4] , \labels[1].label[3] , \labels[1].label[2] , 
	\labels[1].label[1] , \labels[1].label[0] , 
	\labels[1].delimiter_valid[0] , \labels[1].delimiter[7] , 
	\labels[1].delimiter[6] , \labels[1].delimiter[5] , 
	\labels[1].delimiter[4] , \labels[1].delimiter[3] , 
	\labels[1].delimiter[2] , \labels[1].delimiter[1] , 
	\labels[1].delimiter[0] , \labels[0].guid_size[0] , 
	\labels[0].label_size[5] , \labels[0].label_size[4] , 
	\labels[0].label_size[3] , \labels[0].label_size[2] , 
	\labels[0].label_size[1] , \labels[0].label_size[0] , 
	\labels[0].label[255] , \labels[0].label[254] , 
	\labels[0].label[253] , \labels[0].label[252] , 
	\labels[0].label[251] , \labels[0].label[250] , 
	\labels[0].label[249] , \labels[0].label[248] , 
	\labels[0].label[247] , \labels[0].label[246] , 
	\labels[0].label[245] , \labels[0].label[244] , 
	\labels[0].label[243] , \labels[0].label[242] , 
	\labels[0].label[241] , \labels[0].label[240] , 
	\labels[0].label[239] , \labels[0].label[238] , 
	\labels[0].label[237] , \labels[0].label[236] , 
	\labels[0].label[235] , \labels[0].label[234] , 
	\labels[0].label[233] , \labels[0].label[232] , 
	\labels[0].label[231] , \labels[0].label[230] , 
	\labels[0].label[229] , \labels[0].label[228] , 
	\labels[0].label[227] , \labels[0].label[226] , 
	\labels[0].label[225] , \labels[0].label[224] , 
	\labels[0].label[223] , \labels[0].label[222] , 
	\labels[0].label[221] , \labels[0].label[220] , 
	\labels[0].label[219] , \labels[0].label[218] , 
	\labels[0].label[217] , \labels[0].label[216] , 
	\labels[0].label[215] , \labels[0].label[214] , 
	\labels[0].label[213] , \labels[0].label[212] , 
	\labels[0].label[211] , \labels[0].label[210] , 
	\labels[0].label[209] , \labels[0].label[208] , 
	\labels[0].label[207] , \labels[0].label[206] , 
	\labels[0].label[205] , \labels[0].label[204] , 
	\labels[0].label[203] , \labels[0].label[202] , 
	\labels[0].label[201] , \labels[0].label[200] , 
	\labels[0].label[199] , \labels[0].label[198] , 
	\labels[0].label[197] , \labels[0].label[196] , 
	\labels[0].label[195] , \labels[0].label[194] , 
	\labels[0].label[193] , \labels[0].label[192] , 
	\labels[0].label[191] , \labels[0].label[190] , 
	\labels[0].label[189] , \labels[0].label[188] , 
	\labels[0].label[187] , \labels[0].label[186] , 
	\labels[0].label[185] , \labels[0].label[184] , 
	\labels[0].label[183] , \labels[0].label[182] , 
	\labels[0].label[181] , \labels[0].label[180] , 
	\labels[0].label[179] , \labels[0].label[178] , 
	\labels[0].label[177] , \labels[0].label[176] , 
	\labels[0].label[175] , \labels[0].label[174] , 
	\labels[0].label[173] , \labels[0].label[172] , 
	\labels[0].label[171] , \labels[0].label[170] , 
	\labels[0].label[169] , \labels[0].label[168] , 
	\labels[0].label[167] , \labels[0].label[166] , 
	\labels[0].label[165] , \labels[0].label[164] , 
	\labels[0].label[163] , \labels[0].label[162] , 
	\labels[0].label[161] , \labels[0].label[160] , 
	\labels[0].label[159] , \labels[0].label[158] , 
	\labels[0].label[157] , \labels[0].label[156] , 
	\labels[0].label[155] , \labels[0].label[154] , 
	\labels[0].label[153] , \labels[0].label[152] , 
	\labels[0].label[151] , \labels[0].label[150] , 
	\labels[0].label[149] , \labels[0].label[148] , 
	\labels[0].label[147] , \labels[0].label[146] , 
	\labels[0].label[145] , \labels[0].label[144] , 
	\labels[0].label[143] , \labels[0].label[142] , 
	\labels[0].label[141] , \labels[0].label[140] , 
	\labels[0].label[139] , \labels[0].label[138] , 
	\labels[0].label[137] , \labels[0].label[136] , 
	\labels[0].label[135] , \labels[0].label[134] , 
	\labels[0].label[133] , \labels[0].label[132] , 
	\labels[0].label[131] , \labels[0].label[130] , 
	\labels[0].label[129] , \labels[0].label[128] , 
	\labels[0].label[127] , \labels[0].label[126] , 
	\labels[0].label[125] , \labels[0].label[124] , 
	\labels[0].label[123] , \labels[0].label[122] , 
	\labels[0].label[121] , \labels[0].label[120] , 
	\labels[0].label[119] , \labels[0].label[118] , 
	\labels[0].label[117] , \labels[0].label[116] , 
	\labels[0].label[115] , \labels[0].label[114] , 
	\labels[0].label[113] , \labels[0].label[112] , 
	\labels[0].label[111] , \labels[0].label[110] , 
	\labels[0].label[109] , \labels[0].label[108] , 
	\labels[0].label[107] , \labels[0].label[106] , 
	\labels[0].label[105] , \labels[0].label[104] , 
	\labels[0].label[103] , \labels[0].label[102] , 
	\labels[0].label[101] , \labels[0].label[100] , 
	\labels[0].label[99] , \labels[0].label[98] , \labels[0].label[97] , 
	\labels[0].label[96] , \labels[0].label[95] , \labels[0].label[94] , 
	\labels[0].label[93] , \labels[0].label[92] , \labels[0].label[91] , 
	\labels[0].label[90] , \labels[0].label[89] , \labels[0].label[88] , 
	\labels[0].label[87] , \labels[0].label[86] , \labels[0].label[85] , 
	\labels[0].label[84] , \labels[0].label[83] , \labels[0].label[82] , 
	\labels[0].label[81] , \labels[0].label[80] , \labels[0].label[79] , 
	\labels[0].label[78] , \labels[0].label[77] , \labels[0].label[76] , 
	\labels[0].label[75] , \labels[0].label[74] , \labels[0].label[73] , 
	\labels[0].label[72] , \labels[0].label[71] , \labels[0].label[70] , 
	\labels[0].label[69] , \labels[0].label[68] , \labels[0].label[67] , 
	\labels[0].label[66] , \labels[0].label[65] , \labels[0].label[64] , 
	\labels[0].label[63] , \labels[0].label[62] , \labels[0].label[61] , 
	\labels[0].label[60] , \labels[0].label[59] , \labels[0].label[58] , 
	\labels[0].label[57] , \labels[0].label[56] , \labels[0].label[55] , 
	\labels[0].label[54] , \labels[0].label[53] , \labels[0].label[52] , 
	\labels[0].label[51] , \labels[0].label[50] , \labels[0].label[49] , 
	\labels[0].label[48] , \labels[0].label[47] , \labels[0].label[46] , 
	\labels[0].label[45] , \labels[0].label[44] , \labels[0].label[43] , 
	\labels[0].label[42] , \labels[0].label[41] , \labels[0].label[40] , 
	\labels[0].label[39] , \labels[0].label[38] , \labels[0].label[37] , 
	\labels[0].label[36] , \labels[0].label[35] , \labels[0].label[34] , 
	\labels[0].label[33] , \labels[0].label[32] , \labels[0].label[31] , 
	\labels[0].label[30] , \labels[0].label[29] , \labels[0].label[28] , 
	\labels[0].label[27] , \labels[0].label[26] , \labels[0].label[25] , 
	\labels[0].label[24] , \labels[0].label[23] , \labels[0].label[22] , 
	\labels[0].label[21] , \labels[0].label[20] , \labels[0].label[19] , 
	\labels[0].label[18] , \labels[0].label[17] , \labels[0].label[16] , 
	\labels[0].label[15] , \labels[0].label[14] , \labels[0].label[13] , 
	\labels[0].label[12] , \labels[0].label[11] , \labels[0].label[10] , 
	\labels[0].label[9] , \labels[0].label[8] , \labels[0].label[7] , 
	\labels[0].label[6] , \labels[0].label[5] , \labels[0].label[4] , 
	\labels[0].label[3] , \labels[0].label[2] , \labels[0].label[1] , 
	\labels[0].label[0] , \labels[0].delimiter_valid[0] , 
	\labels[0].delimiter[7] , \labels[0].delimiter[6] , 
	\labels[0].delimiter[5] , \labels[0].delimiter[4] , 
	\labels[0].delimiter[3] , \labels[0].delimiter[2] , 
	\labels[0].delimiter[1] , \labels[0].delimiter[0] } ), 
	hash_cmdfifo_ack, hash_len_data_out_ack, hash_in_stall, 
	kdf_test_key_size, kdf_test_mode_en);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output kdfstream_cmdfifo_ack;
output cmdfifo_hash_valid;
output cmdfifo_hash_skip;
output cmdfifo_hash_small_size;
output [31:0] hash_len_data_out;
output hash_len_data_out_valid;
output in_hash_valid;
output in_hash_eof;
output in_hash_eoc;
output [4:0] in_hash_num_bytes;
output [127:0] in_hash_data;
input clk;
input rst_n;
input cmdfifo_kdfstream_valid;
input [0:0] \cmdfifo_kdfstream_cmd.combo_mode ;
input [0:0] \cmdfifo_kdfstream_cmd.skip ;
input [255:0] \cmdfifo_kdfstream_cmd.guid ;
input [2:0] \cmdfifo_kdfstream_cmd.label_index ;
input [1:0] \cmdfifo_kdfstream_cmd.num_iter ;
wire [262:0] cmdfifo_kdfstream_cmd;
input \labels[7].guid_size[0] ,\labels[7].label_size[5] 
	,\labels[7].label_size[4] ,\labels[7].label_size[3] 
	,\labels[7].label_size[2] ,\labels[7].label_size[1] 
	,\labels[7].label_size[0] ,\labels[7].label[255] 
	,\labels[7].label[254] ,\labels[7].label[253] ,\labels[7].label[252] 
	,\labels[7].label[251] ,\labels[7].label[250] ,\labels[7].label[249] 
	,\labels[7].label[248] ,\labels[7].label[247] ,\labels[7].label[246] 
	,\labels[7].label[245] ,\labels[7].label[244] ,\labels[7].label[243] 
	,\labels[7].label[242] ,\labels[7].label[241] ,\labels[7].label[240] 
	,\labels[7].label[239] ,\labels[7].label[238] ,\labels[7].label[237] 
	,\labels[7].label[236] ,\labels[7].label[235] ,\labels[7].label[234] 
	,\labels[7].label[233] ,\labels[7].label[232] ,\labels[7].label[231] 
	,\labels[7].label[230] ,\labels[7].label[229] ,\labels[7].label[228] 
	,\labels[7].label[227] ,\labels[7].label[226] ,\labels[7].label[225] 
	,\labels[7].label[224] ,\labels[7].label[223] ,\labels[7].label[222] 
	,\labels[7].label[221] ,\labels[7].label[220] ,\labels[7].label[219] 
	,\labels[7].label[218] ,\labels[7].label[217] ,\labels[7].label[216] 
	,\labels[7].label[215] ,\labels[7].label[214] ,\labels[7].label[213] 
	,\labels[7].label[212] ,\labels[7].label[211] ,\labels[7].label[210] 
	,\labels[7].label[209] ,\labels[7].label[208] ,\labels[7].label[207] 
	,\labels[7].label[206] ,\labels[7].label[205] ,\labels[7].label[204] 
	,\labels[7].label[203] ,\labels[7].label[202] ,\labels[7].label[201] 
	,\labels[7].label[200] ,\labels[7].label[199] ,\labels[7].label[198] 
	,\labels[7].label[197] ,\labels[7].label[196] ,\labels[7].label[195] 
	,\labels[7].label[194] ,\labels[7].label[193] ,\labels[7].label[192] 
	,\labels[7].label[191] ,\labels[7].label[190] ,\labels[7].label[189] 
	,\labels[7].label[188] ,\labels[7].label[187] ,\labels[7].label[186] 
	,\labels[7].label[185] ,\labels[7].label[184] ,\labels[7].label[183] 
	,\labels[7].label[182] ,\labels[7].label[181] ,\labels[7].label[180] 
	,\labels[7].label[179] ,\labels[7].label[178] ,\labels[7].label[177] 
	,\labels[7].label[176] ,\labels[7].label[175] ,\labels[7].label[174] 
	,\labels[7].label[173] ,\labels[7].label[172] ,\labels[7].label[171] 
	,\labels[7].label[170] ,\labels[7].label[169] ,\labels[7].label[168] 
	,\labels[7].label[167] ,\labels[7].label[166] ,\labels[7].label[165] 
	,\labels[7].label[164] ,\labels[7].label[163] ,\labels[7].label[162] 
	,\labels[7].label[161] ,\labels[7].label[160] ,\labels[7].label[159] 
	,\labels[7].label[158] ,\labels[7].label[157] ,\labels[7].label[156] 
	,\labels[7].label[155] ,\labels[7].label[154] ,\labels[7].label[153] 
	,\labels[7].label[152] ,\labels[7].label[151] ,\labels[7].label[150] 
	,\labels[7].label[149] ,\labels[7].label[148] ,\labels[7].label[147] 
	,\labels[7].label[146] ,\labels[7].label[145] ,\labels[7].label[144] 
	,\labels[7].label[143] ,\labels[7].label[142] ,\labels[7].label[141] 
	,\labels[7].label[140] ,\labels[7].label[139] ,\labels[7].label[138] 
	,\labels[7].label[137] ,\labels[7].label[136] ,\labels[7].label[135] 
	,\labels[7].label[134] ,\labels[7].label[133] ,\labels[7].label[132] 
	,\labels[7].label[131] ,\labels[7].label[130] ,\labels[7].label[129] 
	,\labels[7].label[128] ,\labels[7].label[127] ,\labels[7].label[126] 
	,\labels[7].label[125] ,\labels[7].label[124] ,\labels[7].label[123] 
	,\labels[7].label[122] ,\labels[7].label[121] ,\labels[7].label[120] 
	,\labels[7].label[119] ,\labels[7].label[118] ,\labels[7].label[117] 
	,\labels[7].label[116] ,\labels[7].label[115] ,\labels[7].label[114] 
	,\labels[7].label[113] ,\labels[7].label[112] ,\labels[7].label[111] 
	,\labels[7].label[110] ,\labels[7].label[109] ,\labels[7].label[108] 
	,\labels[7].label[107] ,\labels[7].label[106] ,\labels[7].label[105] 
	,\labels[7].label[104] ,\labels[7].label[103] ,\labels[7].label[102] 
	,\labels[7].label[101] ,\labels[7].label[100] ,\labels[7].label[99] 
	,\labels[7].label[98] ,\labels[7].label[97] ,\labels[7].label[96] 
	,\labels[7].label[95] ,\labels[7].label[94] ,\labels[7].label[93] 
	,\labels[7].label[92] ,\labels[7].label[91] ,\labels[7].label[90] 
	,\labels[7].label[89] ,\labels[7].label[88] ,\labels[7].label[87] 
	,\labels[7].label[86] ,\labels[7].label[85] ,\labels[7].label[84] 
	,\labels[7].label[83] ,\labels[7].label[82] ,\labels[7].label[81] 
	,\labels[7].label[80] ,\labels[7].label[79] ,\labels[7].label[78] 
	,\labels[7].label[77] ,\labels[7].label[76] ,\labels[7].label[75] 
	,\labels[7].label[74] ,\labels[7].label[73] ,\labels[7].label[72] 
	,\labels[7].label[71] ,\labels[7].label[70] ,\labels[7].label[69] 
	,\labels[7].label[68] ,\labels[7].label[67] ,\labels[7].label[66] 
	,\labels[7].label[65] ,\labels[7].label[64] ,\labels[7].label[63] 
	,\labels[7].label[62] ,\labels[7].label[61] ,\labels[7].label[60] 
	,\labels[7].label[59] ,\labels[7].label[58] ,\labels[7].label[57] 
	,\labels[7].label[56] ,\labels[7].label[55] ,\labels[7].label[54] 
	,\labels[7].label[53] ,\labels[7].label[52] ,\labels[7].label[51] 
	,\labels[7].label[50] ,\labels[7].label[49] ,\labels[7].label[48] 
	,\labels[7].label[47] ,\labels[7].label[46] ,\labels[7].label[45] 
	,\labels[7].label[44] ,\labels[7].label[43] ,\labels[7].label[42] 
	,\labels[7].label[41] ,\labels[7].label[40] ,\labels[7].label[39] 
	,\labels[7].label[38] ,\labels[7].label[37] ,\labels[7].label[36] 
	,\labels[7].label[35] ,\labels[7].label[34] ,\labels[7].label[33] 
	,\labels[7].label[32] ,\labels[7].label[31] ,\labels[7].label[30] 
	,\labels[7].label[29] ,\labels[7].label[28] ,\labels[7].label[27] 
	,\labels[7].label[26] ,\labels[7].label[25] ,\labels[7].label[24] 
	,\labels[7].label[23] ,\labels[7].label[22] ,\labels[7].label[21] 
	,\labels[7].label[20] ,\labels[7].label[19] ,\labels[7].label[18] 
	,\labels[7].label[17] ,\labels[7].label[16] ,\labels[7].label[15] 
	,\labels[7].label[14] ,\labels[7].label[13] ,\labels[7].label[12] 
	,\labels[7].label[11] ,\labels[7].label[10] ,\labels[7].label[9] 
	,\labels[7].label[8] ,\labels[7].label[7] ,\labels[7].label[6] 
	,\labels[7].label[5] ,\labels[7].label[4] ,\labels[7].label[3] 
	,\labels[7].label[2] ,\labels[7].label[1] ,\labels[7].label[0] 
	,\labels[7].delimiter_valid[0] ,\labels[7].delimiter[7] 
	,\labels[7].delimiter[6] ,\labels[7].delimiter[5] 
	,\labels[7].delimiter[4] ,\labels[7].delimiter[3] 
	,\labels[7].delimiter[2] ,\labels[7].delimiter[1] 
	,\labels[7].delimiter[0] ,\labels[6].guid_size[0] 
	,\labels[6].label_size[5] ,\labels[6].label_size[4] 
	,\labels[6].label_size[3] ,\labels[6].label_size[2] 
	,\labels[6].label_size[1] ,\labels[6].label_size[0] 
	,\labels[6].label[255] ,\labels[6].label[254] ,\labels[6].label[253] 
	,\labels[6].label[252] ,\labels[6].label[251] ,\labels[6].label[250] 
	,\labels[6].label[249] ,\labels[6].label[248] ,\labels[6].label[247] 
	,\labels[6].label[246] ,\labels[6].label[245] ,\labels[6].label[244] 
	,\labels[6].label[243] ,\labels[6].label[242] ,\labels[6].label[241] 
	,\labels[6].label[240] ,\labels[6].label[239] ,\labels[6].label[238] 
	,\labels[6].label[237] ,\labels[6].label[236] ,\labels[6].label[235] 
	,\labels[6].label[234] ,\labels[6].label[233] ,\labels[6].label[232] 
	,\labels[6].label[231] ,\labels[6].label[230] ,\labels[6].label[229] 
	,\labels[6].label[228] ,\labels[6].label[227] ,\labels[6].label[226] 
	,\labels[6].label[225] ,\labels[6].label[224] ,\labels[6].label[223] 
	,\labels[6].label[222] ,\labels[6].label[221] ,\labels[6].label[220] 
	,\labels[6].label[219] ,\labels[6].label[218] ,\labels[6].label[217] 
	,\labels[6].label[216] ,\labels[6].label[215] ,\labels[6].label[214] 
	,\labels[6].label[213] ,\labels[6].label[212] ,\labels[6].label[211] 
	,\labels[6].label[210] ,\labels[6].label[209] ,\labels[6].label[208] 
	,\labels[6].label[207] ,\labels[6].label[206] ,\labels[6].label[205] 
	,\labels[6].label[204] ,\labels[6].label[203] ,\labels[6].label[202] 
	,\labels[6].label[201] ,\labels[6].label[200] ,\labels[6].label[199] 
	,\labels[6].label[198] ,\labels[6].label[197] ,\labels[6].label[196] 
	,\labels[6].label[195] ,\labels[6].label[194] ,\labels[6].label[193] 
	,\labels[6].label[192] ,\labels[6].label[191] ,\labels[6].label[190] 
	,\labels[6].label[189] ,\labels[6].label[188] ,\labels[6].label[187] 
	,\labels[6].label[186] ,\labels[6].label[185] ,\labels[6].label[184] 
	,\labels[6].label[183] ,\labels[6].label[182] ,\labels[6].label[181] 
	,\labels[6].label[180] ,\labels[6].label[179] ,\labels[6].label[178] 
	,\labels[6].label[177] ,\labels[6].label[176] ,\labels[6].label[175] 
	,\labels[6].label[174] ,\labels[6].label[173] ,\labels[6].label[172] 
	,\labels[6].label[171] ,\labels[6].label[170] ,\labels[6].label[169] 
	,\labels[6].label[168] ,\labels[6].label[167] ,\labels[6].label[166] 
	,\labels[6].label[165] ,\labels[6].label[164] ,\labels[6].label[163] 
	,\labels[6].label[162] ,\labels[6].label[161] ,\labels[6].label[160] 
	,\labels[6].label[159] ,\labels[6].label[158] ,\labels[6].label[157] 
	,\labels[6].label[156] ,\labels[6].label[155] ,\labels[6].label[154] 
	,\labels[6].label[153] ,\labels[6].label[152] ,\labels[6].label[151] 
	,\labels[6].label[150] ,\labels[6].label[149] ,\labels[6].label[148] 
	,\labels[6].label[147] ,\labels[6].label[146] ,\labels[6].label[145] 
	,\labels[6].label[144] ,\labels[6].label[143] ,\labels[6].label[142] 
	,\labels[6].label[141] ,\labels[6].label[140] ,\labels[6].label[139] 
	,\labels[6].label[138] ,\labels[6].label[137] ,\labels[6].label[136] 
	,\labels[6].label[135] ,\labels[6].label[134] ,\labels[6].label[133] 
	,\labels[6].label[132] ,\labels[6].label[131] ,\labels[6].label[130] 
	,\labels[6].label[129] ,\labels[6].label[128] ,\labels[6].label[127] 
	,\labels[6].label[126] ,\labels[6].label[125] ,\labels[6].label[124] 
	,\labels[6].label[123] ,\labels[6].label[122] ,\labels[6].label[121] 
	,\labels[6].label[120] ,\labels[6].label[119] ,\labels[6].label[118] 
	,\labels[6].label[117] ,\labels[6].label[116] ,\labels[6].label[115] 
	,\labels[6].label[114] ,\labels[6].label[113] ,\labels[6].label[112] 
	,\labels[6].label[111] ,\labels[6].label[110] ,\labels[6].label[109] 
	,\labels[6].label[108] ,\labels[6].label[107] ,\labels[6].label[106] 
	,\labels[6].label[105] ,\labels[6].label[104] ,\labels[6].label[103] 
	,\labels[6].label[102] ,\labels[6].label[101] ,\labels[6].label[100] 
	,\labels[6].label[99] ,\labels[6].label[98] ,\labels[6].label[97] 
	,\labels[6].label[96] ,\labels[6].label[95] ,\labels[6].label[94] 
	,\labels[6].label[93] ,\labels[6].label[92] ,\labels[6].label[91] 
	,\labels[6].label[90] ,\labels[6].label[89] ,\labels[6].label[88] 
	,\labels[6].label[87] ,\labels[6].label[86] ,\labels[6].label[85] 
	,\labels[6].label[84] ,\labels[6].label[83] ,\labels[6].label[82] 
	,\labels[6].label[81] ,\labels[6].label[80] ,\labels[6].label[79] 
	,\labels[6].label[78] ,\labels[6].label[77] ,\labels[6].label[76] 
	,\labels[6].label[75] ,\labels[6].label[74] ,\labels[6].label[73] 
	,\labels[6].label[72] ,\labels[6].label[71] ,\labels[6].label[70] 
	,\labels[6].label[69] ,\labels[6].label[68] ,\labels[6].label[67] 
	,\labels[6].label[66] ,\labels[6].label[65] ,\labels[6].label[64] 
	,\labels[6].label[63] ,\labels[6].label[62] ,\labels[6].label[61] 
	,\labels[6].label[60] ,\labels[6].label[59] ,\labels[6].label[58] 
	,\labels[6].label[57] ,\labels[6].label[56] ,\labels[6].label[55] 
	,\labels[6].label[54] ,\labels[6].label[53] ,\labels[6].label[52] 
	,\labels[6].label[51] ,\labels[6].label[50] ,\labels[6].label[49] 
	,\labels[6].label[48] ,\labels[6].label[47] ,\labels[6].label[46] 
	,\labels[6].label[45] ,\labels[6].label[44] ,\labels[6].label[43] 
	,\labels[6].label[42] ,\labels[6].label[41] ,\labels[6].label[40] 
	,\labels[6].label[39] ,\labels[6].label[38] ,\labels[6].label[37] 
	,\labels[6].label[36] ,\labels[6].label[35] ,\labels[6].label[34] 
	,\labels[6].label[33] ,\labels[6].label[32] ,\labels[6].label[31] 
	,\labels[6].label[30] ,\labels[6].label[29] ,\labels[6].label[28] 
	,\labels[6].label[27] ,\labels[6].label[26] ,\labels[6].label[25] 
	,\labels[6].label[24] ,\labels[6].label[23] ,\labels[6].label[22] 
	,\labels[6].label[21] ,\labels[6].label[20] ,\labels[6].label[19] 
	,\labels[6].label[18] ,\labels[6].label[17] ,\labels[6].label[16] 
	,\labels[6].label[15] ,\labels[6].label[14] ,\labels[6].label[13] 
	,\labels[6].label[12] ,\labels[6].label[11] ,\labels[6].label[10] 
	,\labels[6].label[9] ,\labels[6].label[8] ,\labels[6].label[7] 
	,\labels[6].label[6] ,\labels[6].label[5] ,\labels[6].label[4] 
	,\labels[6].label[3] ,\labels[6].label[2] ,\labels[6].label[1] 
	,\labels[6].label[0] ,\labels[6].delimiter_valid[0] 
	,\labels[6].delimiter[7] ,\labels[6].delimiter[6] 
	,\labels[6].delimiter[5] ,\labels[6].delimiter[4] 
	,\labels[6].delimiter[3] ,\labels[6].delimiter[2] 
	,\labels[6].delimiter[1] ,\labels[6].delimiter[0] 
	,\labels[5].guid_size[0] ,\labels[5].label_size[5] 
	,\labels[5].label_size[4] ,\labels[5].label_size[3] 
	,\labels[5].label_size[2] ,\labels[5].label_size[1] 
	,\labels[5].label_size[0] ,\labels[5].label[255] 
	,\labels[5].label[254] ,\labels[5].label[253] ,\labels[5].label[252] 
	,\labels[5].label[251] ,\labels[5].label[250] ,\labels[5].label[249] 
	,\labels[5].label[248] ,\labels[5].label[247] ,\labels[5].label[246] 
	,\labels[5].label[245] ,\labels[5].label[244] ,\labels[5].label[243] 
	,\labels[5].label[242] ,\labels[5].label[241] ,\labels[5].label[240] 
	,\labels[5].label[239] ,\labels[5].label[238] ,\labels[5].label[237] 
	,\labels[5].label[236] ,\labels[5].label[235] ,\labels[5].label[234] 
	,\labels[5].label[233] ,\labels[5].label[232] ,\labels[5].label[231] 
	,\labels[5].label[230] ,\labels[5].label[229] ,\labels[5].label[228] 
	,\labels[5].label[227] ,\labels[5].label[226] ,\labels[5].label[225] 
	,\labels[5].label[224] ,\labels[5].label[223] ,\labels[5].label[222] 
	,\labels[5].label[221] ,\labels[5].label[220] ,\labels[5].label[219] 
	,\labels[5].label[218] ,\labels[5].label[217] ,\labels[5].label[216] 
	,\labels[5].label[215] ,\labels[5].label[214] ,\labels[5].label[213] 
	,\labels[5].label[212] ,\labels[5].label[211] ,\labels[5].label[210] 
	,\labels[5].label[209] ,\labels[5].label[208] ,\labels[5].label[207] 
	,\labels[5].label[206] ,\labels[5].label[205] ,\labels[5].label[204] 
	,\labels[5].label[203] ,\labels[5].label[202] ,\labels[5].label[201] 
	,\labels[5].label[200] ,\labels[5].label[199] ,\labels[5].label[198] 
	,\labels[5].label[197] ,\labels[5].label[196] ,\labels[5].label[195] 
	,\labels[5].label[194] ,\labels[5].label[193] ,\labels[5].label[192] 
	,\labels[5].label[191] ,\labels[5].label[190] ,\labels[5].label[189] 
	,\labels[5].label[188] ,\labels[5].label[187] ,\labels[5].label[186] 
	,\labels[5].label[185] ,\labels[5].label[184] ,\labels[5].label[183] 
	,\labels[5].label[182] ,\labels[5].label[181] ,\labels[5].label[180] 
	,\labels[5].label[179] ,\labels[5].label[178] ,\labels[5].label[177] 
	,\labels[5].label[176] ,\labels[5].label[175] ,\labels[5].label[174] 
	,\labels[5].label[173] ,\labels[5].label[172] ,\labels[5].label[171] 
	,\labels[5].label[170] ,\labels[5].label[169] ,\labels[5].label[168] 
	,\labels[5].label[167] ,\labels[5].label[166] ,\labels[5].label[165] 
	,\labels[5].label[164] ,\labels[5].label[163] ,\labels[5].label[162] 
	,\labels[5].label[161] ,\labels[5].label[160] ,\labels[5].label[159] 
	,\labels[5].label[158] ,\labels[5].label[157] ,\labels[5].label[156] 
	,\labels[5].label[155] ,\labels[5].label[154] ,\labels[5].label[153] 
	,\labels[5].label[152] ,\labels[5].label[151] ,\labels[5].label[150] 
	,\labels[5].label[149] ,\labels[5].label[148] ,\labels[5].label[147] 
	,\labels[5].label[146] ,\labels[5].label[145] ,\labels[5].label[144] 
	,\labels[5].label[143] ,\labels[5].label[142] ,\labels[5].label[141] 
	,\labels[5].label[140] ,\labels[5].label[139] ,\labels[5].label[138] 
	,\labels[5].label[137] ,\labels[5].label[136] ,\labels[5].label[135] 
	,\labels[5].label[134] ,\labels[5].label[133] ,\labels[5].label[132] 
	,\labels[5].label[131] ,\labels[5].label[130] ,\labels[5].label[129] 
	,\labels[5].label[128] ,\labels[5].label[127] ,\labels[5].label[126] 
	,\labels[5].label[125] ,\labels[5].label[124] ,\labels[5].label[123] 
	,\labels[5].label[122] ,\labels[5].label[121] ,\labels[5].label[120] 
	,\labels[5].label[119] ,\labels[5].label[118] ,\labels[5].label[117] 
	,\labels[5].label[116] ,\labels[5].label[115] ,\labels[5].label[114] 
	,\labels[5].label[113] ,\labels[5].label[112] ,\labels[5].label[111] 
	,\labels[5].label[110] ,\labels[5].label[109] ,\labels[5].label[108] 
	,\labels[5].label[107] ,\labels[5].label[106] ,\labels[5].label[105] 
	,\labels[5].label[104] ,\labels[5].label[103] ,\labels[5].label[102] 
	,\labels[5].label[101] ,\labels[5].label[100] ,\labels[5].label[99] 
	,\labels[5].label[98] ,\labels[5].label[97] ,\labels[5].label[96] 
	,\labels[5].label[95] ,\labels[5].label[94] ,\labels[5].label[93] 
	,\labels[5].label[92] ,\labels[5].label[91] ,\labels[5].label[90] 
	,\labels[5].label[89] ,\labels[5].label[88] ,\labels[5].label[87] 
	,\labels[5].label[86] ,\labels[5].label[85] ,\labels[5].label[84] 
	,\labels[5].label[83] ,\labels[5].label[82] ,\labels[5].label[81] 
	,\labels[5].label[80] ,\labels[5].label[79] ,\labels[5].label[78] 
	,\labels[5].label[77] ,\labels[5].label[76] ,\labels[5].label[75] 
	,\labels[5].label[74] ,\labels[5].label[73] ,\labels[5].label[72] 
	,\labels[5].label[71] ,\labels[5].label[70] ,\labels[5].label[69] 
	,\labels[5].label[68] ,\labels[5].label[67] ,\labels[5].label[66] 
	,\labels[5].label[65] ,\labels[5].label[64] ,\labels[5].label[63] 
	,\labels[5].label[62] ,\labels[5].label[61] ,\labels[5].label[60] 
	,\labels[5].label[59] ,\labels[5].label[58] ,\labels[5].label[57] 
	,\labels[5].label[56] ,\labels[5].label[55] ,\labels[5].label[54] 
	,\labels[5].label[53] ,\labels[5].label[52] ,\labels[5].label[51] 
	,\labels[5].label[50] ,\labels[5].label[49] ,\labels[5].label[48] 
	,\labels[5].label[47] ,\labels[5].label[46] ,\labels[5].label[45] 
	,\labels[5].label[44] ,\labels[5].label[43] ,\labels[5].label[42] 
	,\labels[5].label[41] ,\labels[5].label[40] ,\labels[5].label[39] 
	,\labels[5].label[38] ,\labels[5].label[37] ,\labels[5].label[36] 
	,\labels[5].label[35] ,\labels[5].label[34] ,\labels[5].label[33] 
	,\labels[5].label[32] ,\labels[5].label[31] ,\labels[5].label[30] 
	,\labels[5].label[29] ,\labels[5].label[28] ,\labels[5].label[27] 
	,\labels[5].label[26] ,\labels[5].label[25] ,\labels[5].label[24] 
	,\labels[5].label[23] ,\labels[5].label[22] ,\labels[5].label[21] 
	,\labels[5].label[20] ,\labels[5].label[19] ,\labels[5].label[18] 
	,\labels[5].label[17] ,\labels[5].label[16] ,\labels[5].label[15] 
	,\labels[5].label[14] ,\labels[5].label[13] ,\labels[5].label[12] 
	,\labels[5].label[11] ,\labels[5].label[10] ,\labels[5].label[9] 
	,\labels[5].label[8] ,\labels[5].label[7] ,\labels[5].label[6] 
	,\labels[5].label[5] ,\labels[5].label[4] ,\labels[5].label[3] 
	,\labels[5].label[2] ,\labels[5].label[1] ,\labels[5].label[0] 
	,\labels[5].delimiter_valid[0] ,\labels[5].delimiter[7] 
	,\labels[5].delimiter[6] ,\labels[5].delimiter[5] 
	,\labels[5].delimiter[4] ,\labels[5].delimiter[3] 
	,\labels[5].delimiter[2] ,\labels[5].delimiter[1] 
	,\labels[5].delimiter[0] ,\labels[4].guid_size[0] 
	,\labels[4].label_size[5] ,\labels[4].label_size[4] 
	,\labels[4].label_size[3] ,\labels[4].label_size[2] 
	,\labels[4].label_size[1] ,\labels[4].label_size[0] 
	,\labels[4].label[255] ,\labels[4].label[254] ,\labels[4].label[253] 
	,\labels[4].label[252] ,\labels[4].label[251] ,\labels[4].label[250] 
	,\labels[4].label[249] ,\labels[4].label[248] ,\labels[4].label[247] 
	,\labels[4].label[246] ,\labels[4].label[245] ,\labels[4].label[244] 
	,\labels[4].label[243] ,\labels[4].label[242] ,\labels[4].label[241] 
	,\labels[4].label[240] ,\labels[4].label[239] ,\labels[4].label[238] 
	,\labels[4].label[237] ,\labels[4].label[236] ,\labels[4].label[235] 
	,\labels[4].label[234] ,\labels[4].label[233] ,\labels[4].label[232] 
	,\labels[4].label[231] ,\labels[4].label[230] ,\labels[4].label[229] 
	,\labels[4].label[228] ,\labels[4].label[227] ,\labels[4].label[226] 
	,\labels[4].label[225] ,\labels[4].label[224] ,\labels[4].label[223] 
	,\labels[4].label[222] ,\labels[4].label[221] ,\labels[4].label[220] 
	,\labels[4].label[219] ,\labels[4].label[218] ,\labels[4].label[217] 
	,\labels[4].label[216] ,\labels[4].label[215] ,\labels[4].label[214] 
	,\labels[4].label[213] ,\labels[4].label[212] ,\labels[4].label[211] 
	,\labels[4].label[210] ,\labels[4].label[209] ,\labels[4].label[208] 
	,\labels[4].label[207] ,\labels[4].label[206] ,\labels[4].label[205] 
	,\labels[4].label[204] ,\labels[4].label[203] ,\labels[4].label[202] 
	,\labels[4].label[201] ,\labels[4].label[200] ,\labels[4].label[199] 
	,\labels[4].label[198] ,\labels[4].label[197] ,\labels[4].label[196] 
	,\labels[4].label[195] ,\labels[4].label[194] ,\labels[4].label[193] 
	,\labels[4].label[192] ,\labels[4].label[191] ,\labels[4].label[190] 
	,\labels[4].label[189] ,\labels[4].label[188] ,\labels[4].label[187] 
	,\labels[4].label[186] ,\labels[4].label[185] ,\labels[4].label[184] 
	,\labels[4].label[183] ,\labels[4].label[182] ,\labels[4].label[181] 
	,\labels[4].label[180] ,\labels[4].label[179] ,\labels[4].label[178] 
	,\labels[4].label[177] ,\labels[4].label[176] ,\labels[4].label[175] 
	,\labels[4].label[174] ,\labels[4].label[173] ,\labels[4].label[172] 
	,\labels[4].label[171] ,\labels[4].label[170] ,\labels[4].label[169] 
	,\labels[4].label[168] ,\labels[4].label[167] ,\labels[4].label[166] 
	,\labels[4].label[165] ,\labels[4].label[164] ,\labels[4].label[163] 
	,\labels[4].label[162] ,\labels[4].label[161] ,\labels[4].label[160] 
	,\labels[4].label[159] ,\labels[4].label[158] ,\labels[4].label[157] 
	,\labels[4].label[156] ,\labels[4].label[155] ,\labels[4].label[154] 
	,\labels[4].label[153] ,\labels[4].label[152] ,\labels[4].label[151] 
	,\labels[4].label[150] ,\labels[4].label[149] ,\labels[4].label[148] 
	,\labels[4].label[147] ,\labels[4].label[146] ,\labels[4].label[145] 
	,\labels[4].label[144] ,\labels[4].label[143] ,\labels[4].label[142] 
	,\labels[4].label[141] ,\labels[4].label[140] ,\labels[4].label[139] 
	,\labels[4].label[138] ,\labels[4].label[137] ,\labels[4].label[136] 
	,\labels[4].label[135] ,\labels[4].label[134] ,\labels[4].label[133] 
	,\labels[4].label[132] ,\labels[4].label[131] ,\labels[4].label[130] 
	,\labels[4].label[129] ,\labels[4].label[128] ,\labels[4].label[127] 
	,\labels[4].label[126] ,\labels[4].label[125] ,\labels[4].label[124] 
	,\labels[4].label[123] ,\labels[4].label[122] ,\labels[4].label[121] 
	,\labels[4].label[120] ,\labels[4].label[119] ,\labels[4].label[118] 
	,\labels[4].label[117] ,\labels[4].label[116] ,\labels[4].label[115] 
	,\labels[4].label[114] ,\labels[4].label[113] ,\labels[4].label[112] 
	,\labels[4].label[111] ,\labels[4].label[110] ,\labels[4].label[109] 
	,\labels[4].label[108] ,\labels[4].label[107] ,\labels[4].label[106] 
	,\labels[4].label[105] ,\labels[4].label[104] ,\labels[4].label[103] 
	,\labels[4].label[102] ,\labels[4].label[101] ,\labels[4].label[100] 
	,\labels[4].label[99] ,\labels[4].label[98] ,\labels[4].label[97] 
	,\labels[4].label[96] ,\labels[4].label[95] ,\labels[4].label[94] 
	,\labels[4].label[93] ,\labels[4].label[92] ,\labels[4].label[91] 
	,\labels[4].label[90] ,\labels[4].label[89] ,\labels[4].label[88] 
	,\labels[4].label[87] ,\labels[4].label[86] ,\labels[4].label[85] 
	,\labels[4].label[84] ,\labels[4].label[83] ,\labels[4].label[82] 
	,\labels[4].label[81] ,\labels[4].label[80] ,\labels[4].label[79] 
	,\labels[4].label[78] ,\labels[4].label[77] ,\labels[4].label[76] 
	,\labels[4].label[75] ,\labels[4].label[74] ,\labels[4].label[73] 
	,\labels[4].label[72] ,\labels[4].label[71] ,\labels[4].label[70] 
	,\labels[4].label[69] ,\labels[4].label[68] ,\labels[4].label[67] 
	,\labels[4].label[66] ,\labels[4].label[65] ,\labels[4].label[64] 
	,\labels[4].label[63] ,\labels[4].label[62] ,\labels[4].label[61] 
	,\labels[4].label[60] ,\labels[4].label[59] ,\labels[4].label[58] 
	,\labels[4].label[57] ,\labels[4].label[56] ,\labels[4].label[55] 
	,\labels[4].label[54] ,\labels[4].label[53] ,\labels[4].label[52] 
	,\labels[4].label[51] ,\labels[4].label[50] ,\labels[4].label[49] 
	,\labels[4].label[48] ,\labels[4].label[47] ,\labels[4].label[46] 
	,\labels[4].label[45] ,\labels[4].label[44] ,\labels[4].label[43] 
	,\labels[4].label[42] ,\labels[4].label[41] ,\labels[4].label[40] 
	,\labels[4].label[39] ,\labels[4].label[38] ,\labels[4].label[37] 
	,\labels[4].label[36] ,\labels[4].label[35] ,\labels[4].label[34] 
	,\labels[4].label[33] ,\labels[4].label[32] ,\labels[4].label[31] 
	,\labels[4].label[30] ,\labels[4].label[29] ,\labels[4].label[28] 
	,\labels[4].label[27] ,\labels[4].label[26] ,\labels[4].label[25] 
	,\labels[4].label[24] ,\labels[4].label[23] ,\labels[4].label[22] 
	,\labels[4].label[21] ,\labels[4].label[20] ,\labels[4].label[19] 
	,\labels[4].label[18] ,\labels[4].label[17] ,\labels[4].label[16] 
	,\labels[4].label[15] ,\labels[4].label[14] ,\labels[4].label[13] 
	,\labels[4].label[12] ,\labels[4].label[11] ,\labels[4].label[10] 
	,\labels[4].label[9] ,\labels[4].label[8] ,\labels[4].label[7] 
	,\labels[4].label[6] ,\labels[4].label[5] ,\labels[4].label[4] 
	,\labels[4].label[3] ,\labels[4].label[2] ,\labels[4].label[1] 
	,\labels[4].label[0] ,\labels[4].delimiter_valid[0] 
	,\labels[4].delimiter[7] ,\labels[4].delimiter[6] 
	,\labels[4].delimiter[5] ,\labels[4].delimiter[4] 
	,\labels[4].delimiter[3] ,\labels[4].delimiter[2] 
	,\labels[4].delimiter[1] ,\labels[4].delimiter[0] 
	,\labels[3].guid_size[0] ,\labels[3].label_size[5] 
	,\labels[3].label_size[4] ,\labels[3].label_size[3] 
	,\labels[3].label_size[2] ,\labels[3].label_size[1] 
	,\labels[3].label_size[0] ,\labels[3].label[255] 
	,\labels[3].label[254] ,\labels[3].label[253] ,\labels[3].label[252] 
	,\labels[3].label[251] ,\labels[3].label[250] ,\labels[3].label[249] 
	,\labels[3].label[248] ,\labels[3].label[247] ,\labels[3].label[246] 
	,\labels[3].label[245] ,\labels[3].label[244] ,\labels[3].label[243] 
	,\labels[3].label[242] ,\labels[3].label[241] ,\labels[3].label[240] 
	,\labels[3].label[239] ,\labels[3].label[238] ,\labels[3].label[237] 
	,\labels[3].label[236] ,\labels[3].label[235] ,\labels[3].label[234] 
	,\labels[3].label[233] ,\labels[3].label[232] ,\labels[3].label[231] 
	,\labels[3].label[230] ,\labels[3].label[229] ,\labels[3].label[228] 
	,\labels[3].label[227] ,\labels[3].label[226] ,\labels[3].label[225] 
	,\labels[3].label[224] ,\labels[3].label[223] ,\labels[3].label[222] 
	,\labels[3].label[221] ,\labels[3].label[220] ,\labels[3].label[219] 
	,\labels[3].label[218] ,\labels[3].label[217] ,\labels[3].label[216] 
	,\labels[3].label[215] ,\labels[3].label[214] ,\labels[3].label[213] 
	,\labels[3].label[212] ,\labels[3].label[211] ,\labels[3].label[210] 
	,\labels[3].label[209] ,\labels[3].label[208] ,\labels[3].label[207] 
	,\labels[3].label[206] ,\labels[3].label[205] ,\labels[3].label[204] 
	,\labels[3].label[203] ,\labels[3].label[202] ,\labels[3].label[201] 
	,\labels[3].label[200] ,\labels[3].label[199] ,\labels[3].label[198] 
	,\labels[3].label[197] ,\labels[3].label[196] ,\labels[3].label[195] 
	,\labels[3].label[194] ,\labels[3].label[193] ,\labels[3].label[192] 
	,\labels[3].label[191] ,\labels[3].label[190] ,\labels[3].label[189] 
	,\labels[3].label[188] ,\labels[3].label[187] ,\labels[3].label[186] 
	,\labels[3].label[185] ,\labels[3].label[184] ,\labels[3].label[183] 
	,\labels[3].label[182] ,\labels[3].label[181] ,\labels[3].label[180] 
	,\labels[3].label[179] ,\labels[3].label[178] ,\labels[3].label[177] 
	,\labels[3].label[176] ,\labels[3].label[175] ,\labels[3].label[174] 
	,\labels[3].label[173] ,\labels[3].label[172] ,\labels[3].label[171] 
	,\labels[3].label[170] ,\labels[3].label[169] ,\labels[3].label[168] 
	,\labels[3].label[167] ,\labels[3].label[166] ,\labels[3].label[165] 
	,\labels[3].label[164] ,\labels[3].label[163] ,\labels[3].label[162] 
	,\labels[3].label[161] ,\labels[3].label[160] ,\labels[3].label[159] 
	,\labels[3].label[158] ,\labels[3].label[157] ,\labels[3].label[156] 
	,\labels[3].label[155] ,\labels[3].label[154] ,\labels[3].label[153] 
	,\labels[3].label[152] ,\labels[3].label[151] ,\labels[3].label[150] 
	,\labels[3].label[149] ,\labels[3].label[148] ,\labels[3].label[147] 
	,\labels[3].label[146] ,\labels[3].label[145] ,\labels[3].label[144] 
	,\labels[3].label[143] ,\labels[3].label[142] ,\labels[3].label[141] 
	,\labels[3].label[140] ,\labels[3].label[139] ,\labels[3].label[138] 
	,\labels[3].label[137] ,\labels[3].label[136] ,\labels[3].label[135] 
	,\labels[3].label[134] ,\labels[3].label[133] ,\labels[3].label[132] 
	,\labels[3].label[131] ,\labels[3].label[130] ,\labels[3].label[129] 
	,\labels[3].label[128] ,\labels[3].label[127] ,\labels[3].label[126] 
	,\labels[3].label[125] ,\labels[3].label[124] ,\labels[3].label[123] 
	,\labels[3].label[122] ,\labels[3].label[121] ,\labels[3].label[120] 
	,\labels[3].label[119] ,\labels[3].label[118] ,\labels[3].label[117] 
	,\labels[3].label[116] ,\labels[3].label[115] ,\labels[3].label[114] 
	,\labels[3].label[113] ,\labels[3].label[112] ,\labels[3].label[111] 
	,\labels[3].label[110] ,\labels[3].label[109] ,\labels[3].label[108] 
	,\labels[3].label[107] ,\labels[3].label[106] ,\labels[3].label[105] 
	,\labels[3].label[104] ,\labels[3].label[103] ,\labels[3].label[102] 
	,\labels[3].label[101] ,\labels[3].label[100] ,\labels[3].label[99] 
	,\labels[3].label[98] ,\labels[3].label[97] ,\labels[3].label[96] 
	,\labels[3].label[95] ,\labels[3].label[94] ,\labels[3].label[93] 
	,\labels[3].label[92] ,\labels[3].label[91] ,\labels[3].label[90] 
	,\labels[3].label[89] ,\labels[3].label[88] ,\labels[3].label[87] 
	,\labels[3].label[86] ,\labels[3].label[85] ,\labels[3].label[84] 
	,\labels[3].label[83] ,\labels[3].label[82] ,\labels[3].label[81] 
	,\labels[3].label[80] ,\labels[3].label[79] ,\labels[3].label[78] 
	,\labels[3].label[77] ,\labels[3].label[76] ,\labels[3].label[75] 
	,\labels[3].label[74] ,\labels[3].label[73] ,\labels[3].label[72] 
	,\labels[3].label[71] ,\labels[3].label[70] ,\labels[3].label[69] 
	,\labels[3].label[68] ,\labels[3].label[67] ,\labels[3].label[66] 
	,\labels[3].label[65] ,\labels[3].label[64] ,\labels[3].label[63] 
	,\labels[3].label[62] ,\labels[3].label[61] ,\labels[3].label[60] 
	,\labels[3].label[59] ,\labels[3].label[58] ,\labels[3].label[57] 
	,\labels[3].label[56] ,\labels[3].label[55] ,\labels[3].label[54] 
	,\labels[3].label[53] ,\labels[3].label[52] ,\labels[3].label[51] 
	,\labels[3].label[50] ,\labels[3].label[49] ,\labels[3].label[48] 
	,\labels[3].label[47] ,\labels[3].label[46] ,\labels[3].label[45] 
	,\labels[3].label[44] ,\labels[3].label[43] ,\labels[3].label[42] 
	,\labels[3].label[41] ,\labels[3].label[40] ,\labels[3].label[39] 
	,\labels[3].label[38] ,\labels[3].label[37] ,\labels[3].label[36] 
	,\labels[3].label[35] ,\labels[3].label[34] ,\labels[3].label[33] 
	,\labels[3].label[32] ,\labels[3].label[31] ,\labels[3].label[30] 
	,\labels[3].label[29] ,\labels[3].label[28] ,\labels[3].label[27] 
	,\labels[3].label[26] ,\labels[3].label[25] ,\labels[3].label[24] 
	,\labels[3].label[23] ,\labels[3].label[22] ,\labels[3].label[21] 
	,\labels[3].label[20] ,\labels[3].label[19] ,\labels[3].label[18] 
	,\labels[3].label[17] ,\labels[3].label[16] ,\labels[3].label[15] 
	,\labels[3].label[14] ,\labels[3].label[13] ,\labels[3].label[12] 
	,\labels[3].label[11] ,\labels[3].label[10] ,\labels[3].label[9] 
	,\labels[3].label[8] ,\labels[3].label[7] ,\labels[3].label[6] 
	,\labels[3].label[5] ,\labels[3].label[4] ,\labels[3].label[3] 
	,\labels[3].label[2] ,\labels[3].label[1] ,\labels[3].label[0] 
	,\labels[3].delimiter_valid[0] ,\labels[3].delimiter[7] 
	,\labels[3].delimiter[6] ,\labels[3].delimiter[5] 
	,\labels[3].delimiter[4] ,\labels[3].delimiter[3] 
	,\labels[3].delimiter[2] ,\labels[3].delimiter[1] 
	,\labels[3].delimiter[0] ,\labels[2].guid_size[0] 
	,\labels[2].label_size[5] ,\labels[2].label_size[4] 
	,\labels[2].label_size[3] ,\labels[2].label_size[2] 
	,\labels[2].label_size[1] ,\labels[2].label_size[0] 
	,\labels[2].label[255] ,\labels[2].label[254] ,\labels[2].label[253] 
	,\labels[2].label[252] ,\labels[2].label[251] ,\labels[2].label[250] 
	,\labels[2].label[249] ,\labels[2].label[248] ,\labels[2].label[247] 
	,\labels[2].label[246] ,\labels[2].label[245] ,\labels[2].label[244] 
	,\labels[2].label[243] ,\labels[2].label[242] ,\labels[2].label[241] 
	,\labels[2].label[240] ,\labels[2].label[239] ,\labels[2].label[238] 
	,\labels[2].label[237] ,\labels[2].label[236] ,\labels[2].label[235] 
	,\labels[2].label[234] ,\labels[2].label[233] ,\labels[2].label[232] 
	,\labels[2].label[231] ,\labels[2].label[230] ,\labels[2].label[229] 
	,\labels[2].label[228] ,\labels[2].label[227] ,\labels[2].label[226] 
	,\labels[2].label[225] ,\labels[2].label[224] ,\labels[2].label[223] 
	,\labels[2].label[222] ,\labels[2].label[221] ,\labels[2].label[220] 
	,\labels[2].label[219] ,\labels[2].label[218] ,\labels[2].label[217] 
	,\labels[2].label[216] ,\labels[2].label[215] ,\labels[2].label[214] 
	,\labels[2].label[213] ,\labels[2].label[212] ,\labels[2].label[211] 
	,\labels[2].label[210] ,\labels[2].label[209] ,\labels[2].label[208] 
	,\labels[2].label[207] ,\labels[2].label[206] ,\labels[2].label[205] 
	,\labels[2].label[204] ,\labels[2].label[203] ,\labels[2].label[202] 
	,\labels[2].label[201] ,\labels[2].label[200] ,\labels[2].label[199] 
	,\labels[2].label[198] ,\labels[2].label[197] ,\labels[2].label[196] 
	,\labels[2].label[195] ,\labels[2].label[194] ,\labels[2].label[193] 
	,\labels[2].label[192] ,\labels[2].label[191] ,\labels[2].label[190] 
	,\labels[2].label[189] ,\labels[2].label[188] ,\labels[2].label[187] 
	,\labels[2].label[186] ,\labels[2].label[185] ,\labels[2].label[184] 
	,\labels[2].label[183] ,\labels[2].label[182] ,\labels[2].label[181] 
	,\labels[2].label[180] ,\labels[2].label[179] ,\labels[2].label[178] 
	,\labels[2].label[177] ,\labels[2].label[176] ,\labels[2].label[175] 
	,\labels[2].label[174] ,\labels[2].label[173] ,\labels[2].label[172] 
	,\labels[2].label[171] ,\labels[2].label[170] ,\labels[2].label[169] 
	,\labels[2].label[168] ,\labels[2].label[167] ,\labels[2].label[166] 
	,\labels[2].label[165] ,\labels[2].label[164] ,\labels[2].label[163] 
	,\labels[2].label[162] ,\labels[2].label[161] ,\labels[2].label[160] 
	,\labels[2].label[159] ,\labels[2].label[158] ,\labels[2].label[157] 
	,\labels[2].label[156] ,\labels[2].label[155] ,\labels[2].label[154] 
	,\labels[2].label[153] ,\labels[2].label[152] ,\labels[2].label[151] 
	,\labels[2].label[150] ,\labels[2].label[149] ,\labels[2].label[148] 
	,\labels[2].label[147] ,\labels[2].label[146] ,\labels[2].label[145] 
	,\labels[2].label[144] ,\labels[2].label[143] ,\labels[2].label[142] 
	,\labels[2].label[141] ,\labels[2].label[140] ,\labels[2].label[139] 
	,\labels[2].label[138] ,\labels[2].label[137] ,\labels[2].label[136] 
	,\labels[2].label[135] ,\labels[2].label[134] ,\labels[2].label[133] 
	,\labels[2].label[132] ,\labels[2].label[131] ,\labels[2].label[130] 
	,\labels[2].label[129] ,\labels[2].label[128] ,\labels[2].label[127] 
	,\labels[2].label[126] ,\labels[2].label[125] ,\labels[2].label[124] 
	,\labels[2].label[123] ,\labels[2].label[122] ,\labels[2].label[121] 
	,\labels[2].label[120] ,\labels[2].label[119] ,\labels[2].label[118] 
	,\labels[2].label[117] ,\labels[2].label[116] ,\labels[2].label[115] 
	,\labels[2].label[114] ,\labels[2].label[113] ,\labels[2].label[112] 
	,\labels[2].label[111] ,\labels[2].label[110] ,\labels[2].label[109] 
	,\labels[2].label[108] ,\labels[2].label[107] ,\labels[2].label[106] 
	,\labels[2].label[105] ,\labels[2].label[104] ,\labels[2].label[103] 
	,\labels[2].label[102] ,\labels[2].label[101] ,\labels[2].label[100] 
	,\labels[2].label[99] ,\labels[2].label[98] ,\labels[2].label[97] 
	,\labels[2].label[96] ,\labels[2].label[95] ,\labels[2].label[94] 
	,\labels[2].label[93] ,\labels[2].label[92] ,\labels[2].label[91] 
	,\labels[2].label[90] ,\labels[2].label[89] ,\labels[2].label[88] 
	,\labels[2].label[87] ,\labels[2].label[86] ,\labels[2].label[85] 
	,\labels[2].label[84] ,\labels[2].label[83] ,\labels[2].label[82] 
	,\labels[2].label[81] ,\labels[2].label[80] ,\labels[2].label[79] 
	,\labels[2].label[78] ,\labels[2].label[77] ,\labels[2].label[76] 
	,\labels[2].label[75] ,\labels[2].label[74] ,\labels[2].label[73] 
	,\labels[2].label[72] ,\labels[2].label[71] ,\labels[2].label[70] 
	,\labels[2].label[69] ,\labels[2].label[68] ,\labels[2].label[67] 
	,\labels[2].label[66] ,\labels[2].label[65] ,\labels[2].label[64] 
	,\labels[2].label[63] ,\labels[2].label[62] ,\labels[2].label[61] 
	,\labels[2].label[60] ,\labels[2].label[59] ,\labels[2].label[58] 
	,\labels[2].label[57] ,\labels[2].label[56] ,\labels[2].label[55] 
	,\labels[2].label[54] ,\labels[2].label[53] ,\labels[2].label[52] 
	,\labels[2].label[51] ,\labels[2].label[50] ,\labels[2].label[49] 
	,\labels[2].label[48] ,\labels[2].label[47] ,\labels[2].label[46] 
	,\labels[2].label[45] ,\labels[2].label[44] ,\labels[2].label[43] 
	,\labels[2].label[42] ,\labels[2].label[41] ,\labels[2].label[40] 
	,\labels[2].label[39] ,\labels[2].label[38] ,\labels[2].label[37] 
	,\labels[2].label[36] ,\labels[2].label[35] ,\labels[2].label[34] 
	,\labels[2].label[33] ,\labels[2].label[32] ,\labels[2].label[31] 
	,\labels[2].label[30] ,\labels[2].label[29] ,\labels[2].label[28] 
	,\labels[2].label[27] ,\labels[2].label[26] ,\labels[2].label[25] 
	,\labels[2].label[24] ,\labels[2].label[23] ,\labels[2].label[22] 
	,\labels[2].label[21] ,\labels[2].label[20] ,\labels[2].label[19] 
	,\labels[2].label[18] ,\labels[2].label[17] ,\labels[2].label[16] 
	,\labels[2].label[15] ,\labels[2].label[14] ,\labels[2].label[13] 
	,\labels[2].label[12] ,\labels[2].label[11] ,\labels[2].label[10] 
	,\labels[2].label[9] ,\labels[2].label[8] ,\labels[2].label[7] 
	,\labels[2].label[6] ,\labels[2].label[5] ,\labels[2].label[4] 
	,\labels[2].label[3] ,\labels[2].label[2] ,\labels[2].label[1] 
	,\labels[2].label[0] ,\labels[2].delimiter_valid[0] 
	,\labels[2].delimiter[7] ,\labels[2].delimiter[6] 
	,\labels[2].delimiter[5] ,\labels[2].delimiter[4] 
	,\labels[2].delimiter[3] ,\labels[2].delimiter[2] 
	,\labels[2].delimiter[1] ,\labels[2].delimiter[0] 
	,\labels[1].guid_size[0] ,\labels[1].label_size[5] 
	,\labels[1].label_size[4] ,\labels[1].label_size[3] 
	,\labels[1].label_size[2] ,\labels[1].label_size[1] 
	,\labels[1].label_size[0] ,\labels[1].label[255] 
	,\labels[1].label[254] ,\labels[1].label[253] ,\labels[1].label[252] 
	,\labels[1].label[251] ,\labels[1].label[250] ,\labels[1].label[249] 
	,\labels[1].label[248] ,\labels[1].label[247] ,\labels[1].label[246] 
	,\labels[1].label[245] ,\labels[1].label[244] ,\labels[1].label[243] 
	,\labels[1].label[242] ,\labels[1].label[241] ,\labels[1].label[240] 
	,\labels[1].label[239] ,\labels[1].label[238] ,\labels[1].label[237] 
	,\labels[1].label[236] ,\labels[1].label[235] ,\labels[1].label[234] 
	,\labels[1].label[233] ,\labels[1].label[232] ,\labels[1].label[231] 
	,\labels[1].label[230] ,\labels[1].label[229] ,\labels[1].label[228] 
	,\labels[1].label[227] ,\labels[1].label[226] ,\labels[1].label[225] 
	,\labels[1].label[224] ,\labels[1].label[223] ,\labels[1].label[222] 
	,\labels[1].label[221] ,\labels[1].label[220] ,\labels[1].label[219] 
	,\labels[1].label[218] ,\labels[1].label[217] ,\labels[1].label[216] 
	,\labels[1].label[215] ,\labels[1].label[214] ,\labels[1].label[213] 
	,\labels[1].label[212] ,\labels[1].label[211] ,\labels[1].label[210] 
	,\labels[1].label[209] ,\labels[1].label[208] ,\labels[1].label[207] 
	,\labels[1].label[206] ,\labels[1].label[205] ,\labels[1].label[204] 
	,\labels[1].label[203] ,\labels[1].label[202] ,\labels[1].label[201] 
	,\labels[1].label[200] ,\labels[1].label[199] ,\labels[1].label[198] 
	,\labels[1].label[197] ,\labels[1].label[196] ,\labels[1].label[195] 
	,\labels[1].label[194] ,\labels[1].label[193] ,\labels[1].label[192] 
	,\labels[1].label[191] ,\labels[1].label[190] ,\labels[1].label[189] 
	,\labels[1].label[188] ,\labels[1].label[187] ,\labels[1].label[186] 
	,\labels[1].label[185] ,\labels[1].label[184] ,\labels[1].label[183] 
	,\labels[1].label[182] ,\labels[1].label[181] ,\labels[1].label[180] 
	,\labels[1].label[179] ,\labels[1].label[178] ,\labels[1].label[177] 
	,\labels[1].label[176] ,\labels[1].label[175] ,\labels[1].label[174] 
	,\labels[1].label[173] ,\labels[1].label[172] ,\labels[1].label[171] 
	,\labels[1].label[170] ,\labels[1].label[169] ,\labels[1].label[168] 
	,\labels[1].label[167] ,\labels[1].label[166] ,\labels[1].label[165] 
	,\labels[1].label[164] ,\labels[1].label[163] ,\labels[1].label[162] 
	,\labels[1].label[161] ,\labels[1].label[160] ,\labels[1].label[159] 
	,\labels[1].label[158] ,\labels[1].label[157] ,\labels[1].label[156] 
	,\labels[1].label[155] ,\labels[1].label[154] ,\labels[1].label[153] 
	,\labels[1].label[152] ,\labels[1].label[151] ,\labels[1].label[150] 
	,\labels[1].label[149] ,\labels[1].label[148] ,\labels[1].label[147] 
	,\labels[1].label[146] ,\labels[1].label[145] ,\labels[1].label[144] 
	,\labels[1].label[143] ,\labels[1].label[142] ,\labels[1].label[141] 
	,\labels[1].label[140] ,\labels[1].label[139] ,\labels[1].label[138] 
	,\labels[1].label[137] ,\labels[1].label[136] ,\labels[1].label[135] 
	,\labels[1].label[134] ,\labels[1].label[133] ,\labels[1].label[132] 
	,\labels[1].label[131] ,\labels[1].label[130] ,\labels[1].label[129] 
	,\labels[1].label[128] ,\labels[1].label[127] ,\labels[1].label[126] 
	,\labels[1].label[125] ,\labels[1].label[124] ,\labels[1].label[123] 
	,\labels[1].label[122] ,\labels[1].label[121] ,\labels[1].label[120] 
	,\labels[1].label[119] ,\labels[1].label[118] ,\labels[1].label[117] 
	,\labels[1].label[116] ,\labels[1].label[115] ,\labels[1].label[114] 
	,\labels[1].label[113] ,\labels[1].label[112] ,\labels[1].label[111] 
	,\labels[1].label[110] ,\labels[1].label[109] ,\labels[1].label[108] 
	,\labels[1].label[107] ,\labels[1].label[106] ,\labels[1].label[105] 
	,\labels[1].label[104] ,\labels[1].label[103] ,\labels[1].label[102] 
	,\labels[1].label[101] ,\labels[1].label[100] ,\labels[1].label[99] 
	,\labels[1].label[98] ,\labels[1].label[97] ,\labels[1].label[96] 
	,\labels[1].label[95] ,\labels[1].label[94] ,\labels[1].label[93] 
	,\labels[1].label[92] ,\labels[1].label[91] ,\labels[1].label[90] 
	,\labels[1].label[89] ,\labels[1].label[88] ,\labels[1].label[87] 
	,\labels[1].label[86] ,\labels[1].label[85] ,\labels[1].label[84] 
	,\labels[1].label[83] ,\labels[1].label[82] ,\labels[1].label[81] 
	,\labels[1].label[80] ,\labels[1].label[79] ,\labels[1].label[78] 
	,\labels[1].label[77] ,\labels[1].label[76] ,\labels[1].label[75] 
	,\labels[1].label[74] ,\labels[1].label[73] ,\labels[1].label[72] 
	,\labels[1].label[71] ,\labels[1].label[70] ,\labels[1].label[69] 
	,\labels[1].label[68] ,\labels[1].label[67] ,\labels[1].label[66] 
	,\labels[1].label[65] ,\labels[1].label[64] ,\labels[1].label[63] 
	,\labels[1].label[62] ,\labels[1].label[61] ,\labels[1].label[60] 
	,\labels[1].label[59] ,\labels[1].label[58] ,\labels[1].label[57] 
	,\labels[1].label[56] ,\labels[1].label[55] ,\labels[1].label[54] 
	,\labels[1].label[53] ,\labels[1].label[52] ,\labels[1].label[51] 
	,\labels[1].label[50] ,\labels[1].label[49] ,\labels[1].label[48] 
	,\labels[1].label[47] ,\labels[1].label[46] ,\labels[1].label[45] 
	,\labels[1].label[44] ,\labels[1].label[43] ,\labels[1].label[42] 
	,\labels[1].label[41] ,\labels[1].label[40] ,\labels[1].label[39] 
	,\labels[1].label[38] ,\labels[1].label[37] ,\labels[1].label[36] 
	,\labels[1].label[35] ,\labels[1].label[34] ,\labels[1].label[33] 
	,\labels[1].label[32] ,\labels[1].label[31] ,\labels[1].label[30] 
	,\labels[1].label[29] ,\labels[1].label[28] ,\labels[1].label[27] 
	,\labels[1].label[26] ,\labels[1].label[25] ,\labels[1].label[24] 
	,\labels[1].label[23] ,\labels[1].label[22] ,\labels[1].label[21] 
	,\labels[1].label[20] ,\labels[1].label[19] ,\labels[1].label[18] 
	,\labels[1].label[17] ,\labels[1].label[16] ,\labels[1].label[15] 
	,\labels[1].label[14] ,\labels[1].label[13] ,\labels[1].label[12] 
	,\labels[1].label[11] ,\labels[1].label[10] ,\labels[1].label[9] 
	,\labels[1].label[8] ,\labels[1].label[7] ,\labels[1].label[6] 
	,\labels[1].label[5] ,\labels[1].label[4] ,\labels[1].label[3] 
	,\labels[1].label[2] ,\labels[1].label[1] ,\labels[1].label[0] 
	,\labels[1].delimiter_valid[0] ,\labels[1].delimiter[7] 
	,\labels[1].delimiter[6] ,\labels[1].delimiter[5] 
	,\labels[1].delimiter[4] ,\labels[1].delimiter[3] 
	,\labels[1].delimiter[2] ,\labels[1].delimiter[1] 
	,\labels[1].delimiter[0] ,\labels[0].guid_size[0] 
	,\labels[0].label_size[5] ,\labels[0].label_size[4] 
	,\labels[0].label_size[3] ,\labels[0].label_size[2] 
	,\labels[0].label_size[1] ,\labels[0].label_size[0] 
	,\labels[0].label[255] ,\labels[0].label[254] ,\labels[0].label[253] 
	,\labels[0].label[252] ,\labels[0].label[251] ,\labels[0].label[250] 
	,\labels[0].label[249] ,\labels[0].label[248] ,\labels[0].label[247] 
	,\labels[0].label[246] ,\labels[0].label[245] ,\labels[0].label[244] 
	,\labels[0].label[243] ,\labels[0].label[242] ,\labels[0].label[241] 
	,\labels[0].label[240] ,\labels[0].label[239] ,\labels[0].label[238] 
	,\labels[0].label[237] ,\labels[0].label[236] ,\labels[0].label[235] 
	,\labels[0].label[234] ,\labels[0].label[233] ,\labels[0].label[232] 
	,\labels[0].label[231] ,\labels[0].label[230] ,\labels[0].label[229] 
	,\labels[0].label[228] ,\labels[0].label[227] ,\labels[0].label[226] 
	,\labels[0].label[225] ,\labels[0].label[224] ,\labels[0].label[223] 
	,\labels[0].label[222] ,\labels[0].label[221] ,\labels[0].label[220] 
	,\labels[0].label[219] ,\labels[0].label[218] ,\labels[0].label[217] 
	,\labels[0].label[216] ,\labels[0].label[215] ,\labels[0].label[214] 
	,\labels[0].label[213] ,\labels[0].label[212] ,\labels[0].label[211] 
	,\labels[0].label[210] ,\labels[0].label[209] ,\labels[0].label[208] 
	,\labels[0].label[207] ,\labels[0].label[206] ,\labels[0].label[205] 
	,\labels[0].label[204] ,\labels[0].label[203] ,\labels[0].label[202] 
	,\labels[0].label[201] ,\labels[0].label[200] ,\labels[0].label[199] 
	,\labels[0].label[198] ,\labels[0].label[197] ,\labels[0].label[196] 
	,\labels[0].label[195] ,\labels[0].label[194] ,\labels[0].label[193] 
	,\labels[0].label[192] ,\labels[0].label[191] ,\labels[0].label[190] 
	,\labels[0].label[189] ,\labels[0].label[188] ,\labels[0].label[187] 
	,\labels[0].label[186] ,\labels[0].label[185] ,\labels[0].label[184] 
	,\labels[0].label[183] ,\labels[0].label[182] ,\labels[0].label[181] 
	,\labels[0].label[180] ,\labels[0].label[179] ,\labels[0].label[178] 
	,\labels[0].label[177] ,\labels[0].label[176] ,\labels[0].label[175] 
	,\labels[0].label[174] ,\labels[0].label[173] ,\labels[0].label[172] 
	,\labels[0].label[171] ,\labels[0].label[170] ,\labels[0].label[169] 
	,\labels[0].label[168] ,\labels[0].label[167] ,\labels[0].label[166] 
	,\labels[0].label[165] ,\labels[0].label[164] ,\labels[0].label[163] 
	,\labels[0].label[162] ,\labels[0].label[161] ,\labels[0].label[160] 
	,\labels[0].label[159] ,\labels[0].label[158] ,\labels[0].label[157] 
	,\labels[0].label[156] ,\labels[0].label[155] ,\labels[0].label[154] 
	,\labels[0].label[153] ,\labels[0].label[152] ,\labels[0].label[151] 
	,\labels[0].label[150] ,\labels[0].label[149] ,\labels[0].label[148] 
	,\labels[0].label[147] ,\labels[0].label[146] ,\labels[0].label[145] 
	,\labels[0].label[144] ,\labels[0].label[143] ,\labels[0].label[142] 
	,\labels[0].label[141] ,\labels[0].label[140] ,\labels[0].label[139] 
	,\labels[0].label[138] ,\labels[0].label[137] ,\labels[0].label[136] 
	,\labels[0].label[135] ,\labels[0].label[134] ,\labels[0].label[133] 
	,\labels[0].label[132] ,\labels[0].label[131] ,\labels[0].label[130] 
	,\labels[0].label[129] ,\labels[0].label[128] ,\labels[0].label[127] 
	,\labels[0].label[126] ,\labels[0].label[125] ,\labels[0].label[124] 
	,\labels[0].label[123] ,\labels[0].label[122] ,\labels[0].label[121] 
	,\labels[0].label[120] ,\labels[0].label[119] ,\labels[0].label[118] 
	,\labels[0].label[117] ,\labels[0].label[116] ,\labels[0].label[115] 
	,\labels[0].label[114] ,\labels[0].label[113] ,\labels[0].label[112] 
	,\labels[0].label[111] ,\labels[0].label[110] ,\labels[0].label[109] 
	,\labels[0].label[108] ,\labels[0].label[107] ,\labels[0].label[106] 
	,\labels[0].label[105] ,\labels[0].label[104] ,\labels[0].label[103] 
	,\labels[0].label[102] ,\labels[0].label[101] ,\labels[0].label[100] 
	,\labels[0].label[99] ,\labels[0].label[98] ,\labels[0].label[97] 
	,\labels[0].label[96] ,\labels[0].label[95] ,\labels[0].label[94] 
	,\labels[0].label[93] ,\labels[0].label[92] ,\labels[0].label[91] 
	,\labels[0].label[90] ,\labels[0].label[89] ,\labels[0].label[88] 
	,\labels[0].label[87] ,\labels[0].label[86] ,\labels[0].label[85] 
	,\labels[0].label[84] ,\labels[0].label[83] ,\labels[0].label[82] 
	,\labels[0].label[81] ,\labels[0].label[80] ,\labels[0].label[79] 
	,\labels[0].label[78] ,\labels[0].label[77] ,\labels[0].label[76] 
	,\labels[0].label[75] ,\labels[0].label[74] ,\labels[0].label[73] 
	,\labels[0].label[72] ,\labels[0].label[71] ,\labels[0].label[70] 
	,\labels[0].label[69] ,\labels[0].label[68] ,\labels[0].label[67] 
	,\labels[0].label[66] ,\labels[0].label[65] ,\labels[0].label[64] 
	,\labels[0].label[63] ,\labels[0].label[62] ,\labels[0].label[61] 
	,\labels[0].label[60] ,\labels[0].label[59] ,\labels[0].label[58] 
	,\labels[0].label[57] ,\labels[0].label[56] ,\labels[0].label[55] 
	,\labels[0].label[54] ,\labels[0].label[53] ,\labels[0].label[52] 
	,\labels[0].label[51] ,\labels[0].label[50] ,\labels[0].label[49] 
	,\labels[0].label[48] ,\labels[0].label[47] ,\labels[0].label[46] 
	,\labels[0].label[45] ,\labels[0].label[44] ,\labels[0].label[43] 
	,\labels[0].label[42] ,\labels[0].label[41] ,\labels[0].label[40] 
	,\labels[0].label[39] ,\labels[0].label[38] ,\labels[0].label[37] 
	,\labels[0].label[36] ,\labels[0].label[35] ,\labels[0].label[34] 
	,\labels[0].label[33] ,\labels[0].label[32] ,\labels[0].label[31] 
	,\labels[0].label[30] ,\labels[0].label[29] ,\labels[0].label[28] 
	,\labels[0].label[27] ,\labels[0].label[26] ,\labels[0].label[25] 
	,\labels[0].label[24] ,\labels[0].label[23] ,\labels[0].label[22] 
	,\labels[0].label[21] ,\labels[0].label[20] ,\labels[0].label[19] 
	,\labels[0].label[18] ,\labels[0].label[17] ,\labels[0].label[16] 
	,\labels[0].label[15] ,\labels[0].label[14] ,\labels[0].label[13] 
	,\labels[0].label[12] ,\labels[0].label[11] ,\labels[0].label[10] 
	,\labels[0].label[9] ,\labels[0].label[8] ,\labels[0].label[7] 
	,\labels[0].label[6] ,\labels[0].label[5] ,\labels[0].label[4] 
	,\labels[0].label[3] ,\labels[0].label[2] ,\labels[0].label[1] 
	,\labels[0].label[0] ,\labels[0].delimiter_valid[0] 
	,\labels[0].delimiter[7] ,\labels[0].delimiter[6] 
	,\labels[0].delimiter[5] ,\labels[0].delimiter[4] 
	,\labels[0].delimiter[3] ,\labels[0].delimiter[2] 
	,\labels[0].delimiter[1] ,\labels[0].delimiter[0] ;
input hash_cmdfifo_ack;
input hash_len_data_out_ack;
input hash_in_stall;
input [31:0] kdf_test_key_size;
input kdf_test_mode_en;
wire [0:0] hash_cmd_in_stall;
wire [33:0] fifo_out;
wire [0:0] fifo_out_valid;
wire [0:0] fifo_out_ack;
wire [31:0] iter1_kdf_key_size;
wire [31:0] iter2_kdf_key_size;
wire [31:0] iter3_kdf_key_size;
wire st_tx_data;
wire program_pipes;
wire moving_to_tx_data;
wire is_small_size;
wire [31:0] total_hash_size;
wire _zy_simnet_kdfstream_cmdfifo_ack_0_w$;
wire _zy_simnet_cmdfifo_hash_valid_1_w$;
wire _zy_simnet_cmdfifo_hash_skip_2_w$;
wire _zy_simnet_cmdfifo_hash_small_size_3_w$;
wire [0:31] _zy_simnet_hash_len_data_out_4_w$;
wire _zy_simnet_hash_len_data_out_valid_5_w$;
wire _zy_simnet_in_hash_valid_6_w$;
wire _zy_simnet_in_hash_eof_7_w$;
wire _zy_simnet_in_hash_eoc_8_w$;
wire [0:4] _zy_simnet_in_hash_num_bytes_9_w$;
wire [0:127] _zy_simnet_in_hash_data_10_w$;
wire _zy_simnet_cmd_il_valid_11_w$;
wire [0:5] _zy_simnet_cmd_il_data_size_12_w$;
wire [0:287] _zy_simnet_cmd_il_data_13_w$;
wire _zy_simnet_pipe_array_ack_14_w$;
wire [0:4] _zy_simnet_pipe_array_ack_num_bytes_15_w$;
wire _zy_simnet_cmd_dgl_valid_16_w$;
wire [0:5] _zy_simnet_cmd_dgl_data_size_17_w$;
wire [0:295] _zy_simnet_cmd_dgl_data_18_w$;
wire _zy_simnet_pipe_array_ack_19_w$;
wire [0:4] _zy_simnet_pipe_array_ack_num_bytes_20_w$;
wire _zy_simnet_dio_21;
wire _zy_simnet_dio_22;
wire [0:33] _zy_simnet_hash_cmd_in_23_w$;
wire _zy_simnet_hash_cmd_in_valid_24_w$;
wire _zy_simnet_cio_25;
wire cmd_il_valid;
wire [5:0] cmd_il_data_size;
wire [287:0] cmd_il_data;
wire cmd_dgl_valid;
wire [5:0] cmd_dgl_data_size;
wire [295:0] cmd_dgl_data;
wire [1:0] cur_state;
wire [1:0] nxt_state;
wire [1:0] iter_num;
wire [6:0] num_bytes_remaining;
wire [4:0] num_bytes_to_tx;
wire [4:0] in_hash_byte_accumulator;
wire [33:0] hash_cmd_in;
wire [0:0] hash_cmd_in_valid;
wire [31:0] i;
supply0 n1;
tran (cmdfifo_kdfstream_cmd[262], \cmdfifo_kdfstream_cmd.combo_mode [0]);
tran (cmdfifo_kdfstream_cmd[261], \cmdfifo_kdfstream_cmd.skip [0]);
tran (cmdfifo_kdfstream_cmd[260], \cmdfifo_kdfstream_cmd.guid [255]);
tran (cmdfifo_kdfstream_cmd[259], \cmdfifo_kdfstream_cmd.guid [254]);
tran (cmdfifo_kdfstream_cmd[258], \cmdfifo_kdfstream_cmd.guid [253]);
tran (cmdfifo_kdfstream_cmd[257], \cmdfifo_kdfstream_cmd.guid [252]);
tran (cmdfifo_kdfstream_cmd[256], \cmdfifo_kdfstream_cmd.guid [251]);
tran (cmdfifo_kdfstream_cmd[255], \cmdfifo_kdfstream_cmd.guid [250]);
tran (cmdfifo_kdfstream_cmd[254], \cmdfifo_kdfstream_cmd.guid [249]);
tran (cmdfifo_kdfstream_cmd[253], \cmdfifo_kdfstream_cmd.guid [248]);
tran (cmdfifo_kdfstream_cmd[252], \cmdfifo_kdfstream_cmd.guid [247]);
tran (cmdfifo_kdfstream_cmd[251], \cmdfifo_kdfstream_cmd.guid [246]);
tran (cmdfifo_kdfstream_cmd[250], \cmdfifo_kdfstream_cmd.guid [245]);
tran (cmdfifo_kdfstream_cmd[249], \cmdfifo_kdfstream_cmd.guid [244]);
tran (cmdfifo_kdfstream_cmd[248], \cmdfifo_kdfstream_cmd.guid [243]);
tran (cmdfifo_kdfstream_cmd[247], \cmdfifo_kdfstream_cmd.guid [242]);
tran (cmdfifo_kdfstream_cmd[246], \cmdfifo_kdfstream_cmd.guid [241]);
tran (cmdfifo_kdfstream_cmd[245], \cmdfifo_kdfstream_cmd.guid [240]);
tran (cmdfifo_kdfstream_cmd[244], \cmdfifo_kdfstream_cmd.guid [239]);
tran (cmdfifo_kdfstream_cmd[243], \cmdfifo_kdfstream_cmd.guid [238]);
tran (cmdfifo_kdfstream_cmd[242], \cmdfifo_kdfstream_cmd.guid [237]);
tran (cmdfifo_kdfstream_cmd[241], \cmdfifo_kdfstream_cmd.guid [236]);
tran (cmdfifo_kdfstream_cmd[240], \cmdfifo_kdfstream_cmd.guid [235]);
tran (cmdfifo_kdfstream_cmd[239], \cmdfifo_kdfstream_cmd.guid [234]);
tran (cmdfifo_kdfstream_cmd[238], \cmdfifo_kdfstream_cmd.guid [233]);
tran (cmdfifo_kdfstream_cmd[237], \cmdfifo_kdfstream_cmd.guid [232]);
tran (cmdfifo_kdfstream_cmd[236], \cmdfifo_kdfstream_cmd.guid [231]);
tran (cmdfifo_kdfstream_cmd[235], \cmdfifo_kdfstream_cmd.guid [230]);
tran (cmdfifo_kdfstream_cmd[234], \cmdfifo_kdfstream_cmd.guid [229]);
tran (cmdfifo_kdfstream_cmd[233], \cmdfifo_kdfstream_cmd.guid [228]);
tran (cmdfifo_kdfstream_cmd[232], \cmdfifo_kdfstream_cmd.guid [227]);
tran (cmdfifo_kdfstream_cmd[231], \cmdfifo_kdfstream_cmd.guid [226]);
tran (cmdfifo_kdfstream_cmd[230], \cmdfifo_kdfstream_cmd.guid [225]);
tran (cmdfifo_kdfstream_cmd[229], \cmdfifo_kdfstream_cmd.guid [224]);
tran (cmdfifo_kdfstream_cmd[228], \cmdfifo_kdfstream_cmd.guid [223]);
tran (cmdfifo_kdfstream_cmd[227], \cmdfifo_kdfstream_cmd.guid [222]);
tran (cmdfifo_kdfstream_cmd[226], \cmdfifo_kdfstream_cmd.guid [221]);
tran (cmdfifo_kdfstream_cmd[225], \cmdfifo_kdfstream_cmd.guid [220]);
tran (cmdfifo_kdfstream_cmd[224], \cmdfifo_kdfstream_cmd.guid [219]);
tran (cmdfifo_kdfstream_cmd[223], \cmdfifo_kdfstream_cmd.guid [218]);
tran (cmdfifo_kdfstream_cmd[222], \cmdfifo_kdfstream_cmd.guid [217]);
tran (cmdfifo_kdfstream_cmd[221], \cmdfifo_kdfstream_cmd.guid [216]);
tran (cmdfifo_kdfstream_cmd[220], \cmdfifo_kdfstream_cmd.guid [215]);
tran (cmdfifo_kdfstream_cmd[219], \cmdfifo_kdfstream_cmd.guid [214]);
tran (cmdfifo_kdfstream_cmd[218], \cmdfifo_kdfstream_cmd.guid [213]);
tran (cmdfifo_kdfstream_cmd[217], \cmdfifo_kdfstream_cmd.guid [212]);
tran (cmdfifo_kdfstream_cmd[216], \cmdfifo_kdfstream_cmd.guid [211]);
tran (cmdfifo_kdfstream_cmd[215], \cmdfifo_kdfstream_cmd.guid [210]);
tran (cmdfifo_kdfstream_cmd[214], \cmdfifo_kdfstream_cmd.guid [209]);
tran (cmdfifo_kdfstream_cmd[213], \cmdfifo_kdfstream_cmd.guid [208]);
tran (cmdfifo_kdfstream_cmd[212], \cmdfifo_kdfstream_cmd.guid [207]);
tran (cmdfifo_kdfstream_cmd[211], \cmdfifo_kdfstream_cmd.guid [206]);
tran (cmdfifo_kdfstream_cmd[210], \cmdfifo_kdfstream_cmd.guid [205]);
tran (cmdfifo_kdfstream_cmd[209], \cmdfifo_kdfstream_cmd.guid [204]);
tran (cmdfifo_kdfstream_cmd[208], \cmdfifo_kdfstream_cmd.guid [203]);
tran (cmdfifo_kdfstream_cmd[207], \cmdfifo_kdfstream_cmd.guid [202]);
tran (cmdfifo_kdfstream_cmd[206], \cmdfifo_kdfstream_cmd.guid [201]);
tran (cmdfifo_kdfstream_cmd[205], \cmdfifo_kdfstream_cmd.guid [200]);
tran (cmdfifo_kdfstream_cmd[204], \cmdfifo_kdfstream_cmd.guid [199]);
tran (cmdfifo_kdfstream_cmd[203], \cmdfifo_kdfstream_cmd.guid [198]);
tran (cmdfifo_kdfstream_cmd[202], \cmdfifo_kdfstream_cmd.guid [197]);
tran (cmdfifo_kdfstream_cmd[201], \cmdfifo_kdfstream_cmd.guid [196]);
tran (cmdfifo_kdfstream_cmd[200], \cmdfifo_kdfstream_cmd.guid [195]);
tran (cmdfifo_kdfstream_cmd[199], \cmdfifo_kdfstream_cmd.guid [194]);
tran (cmdfifo_kdfstream_cmd[198], \cmdfifo_kdfstream_cmd.guid [193]);
tran (cmdfifo_kdfstream_cmd[197], \cmdfifo_kdfstream_cmd.guid [192]);
tran (cmdfifo_kdfstream_cmd[196], \cmdfifo_kdfstream_cmd.guid [191]);
tran (cmdfifo_kdfstream_cmd[195], \cmdfifo_kdfstream_cmd.guid [190]);
tran (cmdfifo_kdfstream_cmd[194], \cmdfifo_kdfstream_cmd.guid [189]);
tran (cmdfifo_kdfstream_cmd[193], \cmdfifo_kdfstream_cmd.guid [188]);
tran (cmdfifo_kdfstream_cmd[192], \cmdfifo_kdfstream_cmd.guid [187]);
tran (cmdfifo_kdfstream_cmd[191], \cmdfifo_kdfstream_cmd.guid [186]);
tran (cmdfifo_kdfstream_cmd[190], \cmdfifo_kdfstream_cmd.guid [185]);
tran (cmdfifo_kdfstream_cmd[189], \cmdfifo_kdfstream_cmd.guid [184]);
tran (cmdfifo_kdfstream_cmd[188], \cmdfifo_kdfstream_cmd.guid [183]);
tran (cmdfifo_kdfstream_cmd[187], \cmdfifo_kdfstream_cmd.guid [182]);
tran (cmdfifo_kdfstream_cmd[186], \cmdfifo_kdfstream_cmd.guid [181]);
tran (cmdfifo_kdfstream_cmd[185], \cmdfifo_kdfstream_cmd.guid [180]);
tran (cmdfifo_kdfstream_cmd[184], \cmdfifo_kdfstream_cmd.guid [179]);
tran (cmdfifo_kdfstream_cmd[183], \cmdfifo_kdfstream_cmd.guid [178]);
tran (cmdfifo_kdfstream_cmd[182], \cmdfifo_kdfstream_cmd.guid [177]);
tran (cmdfifo_kdfstream_cmd[181], \cmdfifo_kdfstream_cmd.guid [176]);
tran (cmdfifo_kdfstream_cmd[180], \cmdfifo_kdfstream_cmd.guid [175]);
tran (cmdfifo_kdfstream_cmd[179], \cmdfifo_kdfstream_cmd.guid [174]);
tran (cmdfifo_kdfstream_cmd[178], \cmdfifo_kdfstream_cmd.guid [173]);
tran (cmdfifo_kdfstream_cmd[177], \cmdfifo_kdfstream_cmd.guid [172]);
tran (cmdfifo_kdfstream_cmd[176], \cmdfifo_kdfstream_cmd.guid [171]);
tran (cmdfifo_kdfstream_cmd[175], \cmdfifo_kdfstream_cmd.guid [170]);
tran (cmdfifo_kdfstream_cmd[174], \cmdfifo_kdfstream_cmd.guid [169]);
tran (cmdfifo_kdfstream_cmd[173], \cmdfifo_kdfstream_cmd.guid [168]);
tran (cmdfifo_kdfstream_cmd[172], \cmdfifo_kdfstream_cmd.guid [167]);
tran (cmdfifo_kdfstream_cmd[171], \cmdfifo_kdfstream_cmd.guid [166]);
tran (cmdfifo_kdfstream_cmd[170], \cmdfifo_kdfstream_cmd.guid [165]);
tran (cmdfifo_kdfstream_cmd[169], \cmdfifo_kdfstream_cmd.guid [164]);
tran (cmdfifo_kdfstream_cmd[168], \cmdfifo_kdfstream_cmd.guid [163]);
tran (cmdfifo_kdfstream_cmd[167], \cmdfifo_kdfstream_cmd.guid [162]);
tran (cmdfifo_kdfstream_cmd[166], \cmdfifo_kdfstream_cmd.guid [161]);
tran (cmdfifo_kdfstream_cmd[165], \cmdfifo_kdfstream_cmd.guid [160]);
tran (cmdfifo_kdfstream_cmd[164], \cmdfifo_kdfstream_cmd.guid [159]);
tran (cmdfifo_kdfstream_cmd[163], \cmdfifo_kdfstream_cmd.guid [158]);
tran (cmdfifo_kdfstream_cmd[162], \cmdfifo_kdfstream_cmd.guid [157]);
tran (cmdfifo_kdfstream_cmd[161], \cmdfifo_kdfstream_cmd.guid [156]);
tran (cmdfifo_kdfstream_cmd[160], \cmdfifo_kdfstream_cmd.guid [155]);
tran (cmdfifo_kdfstream_cmd[159], \cmdfifo_kdfstream_cmd.guid [154]);
tran (cmdfifo_kdfstream_cmd[158], \cmdfifo_kdfstream_cmd.guid [153]);
tran (cmdfifo_kdfstream_cmd[157], \cmdfifo_kdfstream_cmd.guid [152]);
tran (cmdfifo_kdfstream_cmd[156], \cmdfifo_kdfstream_cmd.guid [151]);
tran (cmdfifo_kdfstream_cmd[155], \cmdfifo_kdfstream_cmd.guid [150]);
tran (cmdfifo_kdfstream_cmd[154], \cmdfifo_kdfstream_cmd.guid [149]);
tran (cmdfifo_kdfstream_cmd[153], \cmdfifo_kdfstream_cmd.guid [148]);
tran (cmdfifo_kdfstream_cmd[152], \cmdfifo_kdfstream_cmd.guid [147]);
tran (cmdfifo_kdfstream_cmd[151], \cmdfifo_kdfstream_cmd.guid [146]);
tran (cmdfifo_kdfstream_cmd[150], \cmdfifo_kdfstream_cmd.guid [145]);
tran (cmdfifo_kdfstream_cmd[149], \cmdfifo_kdfstream_cmd.guid [144]);
tran (cmdfifo_kdfstream_cmd[148], \cmdfifo_kdfstream_cmd.guid [143]);
tran (cmdfifo_kdfstream_cmd[147], \cmdfifo_kdfstream_cmd.guid [142]);
tran (cmdfifo_kdfstream_cmd[146], \cmdfifo_kdfstream_cmd.guid [141]);
tran (cmdfifo_kdfstream_cmd[145], \cmdfifo_kdfstream_cmd.guid [140]);
tran (cmdfifo_kdfstream_cmd[144], \cmdfifo_kdfstream_cmd.guid [139]);
tran (cmdfifo_kdfstream_cmd[143], \cmdfifo_kdfstream_cmd.guid [138]);
tran (cmdfifo_kdfstream_cmd[142], \cmdfifo_kdfstream_cmd.guid [137]);
tran (cmdfifo_kdfstream_cmd[141], \cmdfifo_kdfstream_cmd.guid [136]);
tran (cmdfifo_kdfstream_cmd[140], \cmdfifo_kdfstream_cmd.guid [135]);
tran (cmdfifo_kdfstream_cmd[139], \cmdfifo_kdfstream_cmd.guid [134]);
tran (cmdfifo_kdfstream_cmd[138], \cmdfifo_kdfstream_cmd.guid [133]);
tran (cmdfifo_kdfstream_cmd[137], \cmdfifo_kdfstream_cmd.guid [132]);
tran (cmdfifo_kdfstream_cmd[136], \cmdfifo_kdfstream_cmd.guid [131]);
tran (cmdfifo_kdfstream_cmd[135], \cmdfifo_kdfstream_cmd.guid [130]);
tran (cmdfifo_kdfstream_cmd[134], \cmdfifo_kdfstream_cmd.guid [129]);
tran (cmdfifo_kdfstream_cmd[133], \cmdfifo_kdfstream_cmd.guid [128]);
tran (cmdfifo_kdfstream_cmd[132], \cmdfifo_kdfstream_cmd.guid [127]);
tran (cmdfifo_kdfstream_cmd[131], \cmdfifo_kdfstream_cmd.guid [126]);
tran (cmdfifo_kdfstream_cmd[130], \cmdfifo_kdfstream_cmd.guid [125]);
tran (cmdfifo_kdfstream_cmd[129], \cmdfifo_kdfstream_cmd.guid [124]);
tran (cmdfifo_kdfstream_cmd[128], \cmdfifo_kdfstream_cmd.guid [123]);
tran (cmdfifo_kdfstream_cmd[127], \cmdfifo_kdfstream_cmd.guid [122]);
tran (cmdfifo_kdfstream_cmd[126], \cmdfifo_kdfstream_cmd.guid [121]);
tran (cmdfifo_kdfstream_cmd[125], \cmdfifo_kdfstream_cmd.guid [120]);
tran (cmdfifo_kdfstream_cmd[124], \cmdfifo_kdfstream_cmd.guid [119]);
tran (cmdfifo_kdfstream_cmd[123], \cmdfifo_kdfstream_cmd.guid [118]);
tran (cmdfifo_kdfstream_cmd[122], \cmdfifo_kdfstream_cmd.guid [117]);
tran (cmdfifo_kdfstream_cmd[121], \cmdfifo_kdfstream_cmd.guid [116]);
tran (cmdfifo_kdfstream_cmd[120], \cmdfifo_kdfstream_cmd.guid [115]);
tran (cmdfifo_kdfstream_cmd[119], \cmdfifo_kdfstream_cmd.guid [114]);
tran (cmdfifo_kdfstream_cmd[118], \cmdfifo_kdfstream_cmd.guid [113]);
tran (cmdfifo_kdfstream_cmd[117], \cmdfifo_kdfstream_cmd.guid [112]);
tran (cmdfifo_kdfstream_cmd[116], \cmdfifo_kdfstream_cmd.guid [111]);
tran (cmdfifo_kdfstream_cmd[115], \cmdfifo_kdfstream_cmd.guid [110]);
tran (cmdfifo_kdfstream_cmd[114], \cmdfifo_kdfstream_cmd.guid [109]);
tran (cmdfifo_kdfstream_cmd[113], \cmdfifo_kdfstream_cmd.guid [108]);
tran (cmdfifo_kdfstream_cmd[112], \cmdfifo_kdfstream_cmd.guid [107]);
tran (cmdfifo_kdfstream_cmd[111], \cmdfifo_kdfstream_cmd.guid [106]);
tran (cmdfifo_kdfstream_cmd[110], \cmdfifo_kdfstream_cmd.guid [105]);
tran (cmdfifo_kdfstream_cmd[109], \cmdfifo_kdfstream_cmd.guid [104]);
tran (cmdfifo_kdfstream_cmd[108], \cmdfifo_kdfstream_cmd.guid [103]);
tran (cmdfifo_kdfstream_cmd[107], \cmdfifo_kdfstream_cmd.guid [102]);
tran (cmdfifo_kdfstream_cmd[106], \cmdfifo_kdfstream_cmd.guid [101]);
tran (cmdfifo_kdfstream_cmd[105], \cmdfifo_kdfstream_cmd.guid [100]);
tran (cmdfifo_kdfstream_cmd[104], \cmdfifo_kdfstream_cmd.guid [99]);
tran (cmdfifo_kdfstream_cmd[103], \cmdfifo_kdfstream_cmd.guid [98]);
tran (cmdfifo_kdfstream_cmd[102], \cmdfifo_kdfstream_cmd.guid [97]);
tran (cmdfifo_kdfstream_cmd[101], \cmdfifo_kdfstream_cmd.guid [96]);
tran (cmdfifo_kdfstream_cmd[100], \cmdfifo_kdfstream_cmd.guid [95]);
tran (cmdfifo_kdfstream_cmd[99], \cmdfifo_kdfstream_cmd.guid [94]);
tran (cmdfifo_kdfstream_cmd[98], \cmdfifo_kdfstream_cmd.guid [93]);
tran (cmdfifo_kdfstream_cmd[97], \cmdfifo_kdfstream_cmd.guid [92]);
tran (cmdfifo_kdfstream_cmd[96], \cmdfifo_kdfstream_cmd.guid [91]);
tran (cmdfifo_kdfstream_cmd[95], \cmdfifo_kdfstream_cmd.guid [90]);
tran (cmdfifo_kdfstream_cmd[94], \cmdfifo_kdfstream_cmd.guid [89]);
tran (cmdfifo_kdfstream_cmd[93], \cmdfifo_kdfstream_cmd.guid [88]);
tran (cmdfifo_kdfstream_cmd[92], \cmdfifo_kdfstream_cmd.guid [87]);
tran (cmdfifo_kdfstream_cmd[91], \cmdfifo_kdfstream_cmd.guid [86]);
tran (cmdfifo_kdfstream_cmd[90], \cmdfifo_kdfstream_cmd.guid [85]);
tran (cmdfifo_kdfstream_cmd[89], \cmdfifo_kdfstream_cmd.guid [84]);
tran (cmdfifo_kdfstream_cmd[88], \cmdfifo_kdfstream_cmd.guid [83]);
tran (cmdfifo_kdfstream_cmd[87], \cmdfifo_kdfstream_cmd.guid [82]);
tran (cmdfifo_kdfstream_cmd[86], \cmdfifo_kdfstream_cmd.guid [81]);
tran (cmdfifo_kdfstream_cmd[85], \cmdfifo_kdfstream_cmd.guid [80]);
tran (cmdfifo_kdfstream_cmd[84], \cmdfifo_kdfstream_cmd.guid [79]);
tran (cmdfifo_kdfstream_cmd[83], \cmdfifo_kdfstream_cmd.guid [78]);
tran (cmdfifo_kdfstream_cmd[82], \cmdfifo_kdfstream_cmd.guid [77]);
tran (cmdfifo_kdfstream_cmd[81], \cmdfifo_kdfstream_cmd.guid [76]);
tran (cmdfifo_kdfstream_cmd[80], \cmdfifo_kdfstream_cmd.guid [75]);
tran (cmdfifo_kdfstream_cmd[79], \cmdfifo_kdfstream_cmd.guid [74]);
tran (cmdfifo_kdfstream_cmd[78], \cmdfifo_kdfstream_cmd.guid [73]);
tran (cmdfifo_kdfstream_cmd[77], \cmdfifo_kdfstream_cmd.guid [72]);
tran (cmdfifo_kdfstream_cmd[76], \cmdfifo_kdfstream_cmd.guid [71]);
tran (cmdfifo_kdfstream_cmd[75], \cmdfifo_kdfstream_cmd.guid [70]);
tran (cmdfifo_kdfstream_cmd[74], \cmdfifo_kdfstream_cmd.guid [69]);
tran (cmdfifo_kdfstream_cmd[73], \cmdfifo_kdfstream_cmd.guid [68]);
tran (cmdfifo_kdfstream_cmd[72], \cmdfifo_kdfstream_cmd.guid [67]);
tran (cmdfifo_kdfstream_cmd[71], \cmdfifo_kdfstream_cmd.guid [66]);
tran (cmdfifo_kdfstream_cmd[70], \cmdfifo_kdfstream_cmd.guid [65]);
tran (cmdfifo_kdfstream_cmd[69], \cmdfifo_kdfstream_cmd.guid [64]);
tran (cmdfifo_kdfstream_cmd[68], \cmdfifo_kdfstream_cmd.guid [63]);
tran (cmdfifo_kdfstream_cmd[67], \cmdfifo_kdfstream_cmd.guid [62]);
tran (cmdfifo_kdfstream_cmd[66], \cmdfifo_kdfstream_cmd.guid [61]);
tran (cmdfifo_kdfstream_cmd[65], \cmdfifo_kdfstream_cmd.guid [60]);
tran (cmdfifo_kdfstream_cmd[64], \cmdfifo_kdfstream_cmd.guid [59]);
tran (cmdfifo_kdfstream_cmd[63], \cmdfifo_kdfstream_cmd.guid [58]);
tran (cmdfifo_kdfstream_cmd[62], \cmdfifo_kdfstream_cmd.guid [57]);
tran (cmdfifo_kdfstream_cmd[61], \cmdfifo_kdfstream_cmd.guid [56]);
tran (cmdfifo_kdfstream_cmd[60], \cmdfifo_kdfstream_cmd.guid [55]);
tran (cmdfifo_kdfstream_cmd[59], \cmdfifo_kdfstream_cmd.guid [54]);
tran (cmdfifo_kdfstream_cmd[58], \cmdfifo_kdfstream_cmd.guid [53]);
tran (cmdfifo_kdfstream_cmd[57], \cmdfifo_kdfstream_cmd.guid [52]);
tran (cmdfifo_kdfstream_cmd[56], \cmdfifo_kdfstream_cmd.guid [51]);
tran (cmdfifo_kdfstream_cmd[55], \cmdfifo_kdfstream_cmd.guid [50]);
tran (cmdfifo_kdfstream_cmd[54], \cmdfifo_kdfstream_cmd.guid [49]);
tran (cmdfifo_kdfstream_cmd[53], \cmdfifo_kdfstream_cmd.guid [48]);
tran (cmdfifo_kdfstream_cmd[52], \cmdfifo_kdfstream_cmd.guid [47]);
tran (cmdfifo_kdfstream_cmd[51], \cmdfifo_kdfstream_cmd.guid [46]);
tran (cmdfifo_kdfstream_cmd[50], \cmdfifo_kdfstream_cmd.guid [45]);
tran (cmdfifo_kdfstream_cmd[49], \cmdfifo_kdfstream_cmd.guid [44]);
tran (cmdfifo_kdfstream_cmd[48], \cmdfifo_kdfstream_cmd.guid [43]);
tran (cmdfifo_kdfstream_cmd[47], \cmdfifo_kdfstream_cmd.guid [42]);
tran (cmdfifo_kdfstream_cmd[46], \cmdfifo_kdfstream_cmd.guid [41]);
tran (cmdfifo_kdfstream_cmd[45], \cmdfifo_kdfstream_cmd.guid [40]);
tran (cmdfifo_kdfstream_cmd[44], \cmdfifo_kdfstream_cmd.guid [39]);
tran (cmdfifo_kdfstream_cmd[43], \cmdfifo_kdfstream_cmd.guid [38]);
tran (cmdfifo_kdfstream_cmd[42], \cmdfifo_kdfstream_cmd.guid [37]);
tran (cmdfifo_kdfstream_cmd[41], \cmdfifo_kdfstream_cmd.guid [36]);
tran (cmdfifo_kdfstream_cmd[40], \cmdfifo_kdfstream_cmd.guid [35]);
tran (cmdfifo_kdfstream_cmd[39], \cmdfifo_kdfstream_cmd.guid [34]);
tran (cmdfifo_kdfstream_cmd[38], \cmdfifo_kdfstream_cmd.guid [33]);
tran (cmdfifo_kdfstream_cmd[37], \cmdfifo_kdfstream_cmd.guid [32]);
tran (cmdfifo_kdfstream_cmd[36], \cmdfifo_kdfstream_cmd.guid [31]);
tran (cmdfifo_kdfstream_cmd[35], \cmdfifo_kdfstream_cmd.guid [30]);
tran (cmdfifo_kdfstream_cmd[34], \cmdfifo_kdfstream_cmd.guid [29]);
tran (cmdfifo_kdfstream_cmd[33], \cmdfifo_kdfstream_cmd.guid [28]);
tran (cmdfifo_kdfstream_cmd[32], \cmdfifo_kdfstream_cmd.guid [27]);
tran (cmdfifo_kdfstream_cmd[31], \cmdfifo_kdfstream_cmd.guid [26]);
tran (cmdfifo_kdfstream_cmd[30], \cmdfifo_kdfstream_cmd.guid [25]);
tran (cmdfifo_kdfstream_cmd[29], \cmdfifo_kdfstream_cmd.guid [24]);
tran (cmdfifo_kdfstream_cmd[28], \cmdfifo_kdfstream_cmd.guid [23]);
tran (cmdfifo_kdfstream_cmd[27], \cmdfifo_kdfstream_cmd.guid [22]);
tran (cmdfifo_kdfstream_cmd[26], \cmdfifo_kdfstream_cmd.guid [21]);
tran (cmdfifo_kdfstream_cmd[25], \cmdfifo_kdfstream_cmd.guid [20]);
tran (cmdfifo_kdfstream_cmd[24], \cmdfifo_kdfstream_cmd.guid [19]);
tran (cmdfifo_kdfstream_cmd[23], \cmdfifo_kdfstream_cmd.guid [18]);
tran (cmdfifo_kdfstream_cmd[22], \cmdfifo_kdfstream_cmd.guid [17]);
tran (cmdfifo_kdfstream_cmd[21], \cmdfifo_kdfstream_cmd.guid [16]);
tran (cmdfifo_kdfstream_cmd[20], \cmdfifo_kdfstream_cmd.guid [15]);
tran (cmdfifo_kdfstream_cmd[19], \cmdfifo_kdfstream_cmd.guid [14]);
tran (cmdfifo_kdfstream_cmd[18], \cmdfifo_kdfstream_cmd.guid [13]);
tran (cmdfifo_kdfstream_cmd[17], \cmdfifo_kdfstream_cmd.guid [12]);
tran (cmdfifo_kdfstream_cmd[16], \cmdfifo_kdfstream_cmd.guid [11]);
tran (cmdfifo_kdfstream_cmd[15], \cmdfifo_kdfstream_cmd.guid [10]);
tran (cmdfifo_kdfstream_cmd[14], \cmdfifo_kdfstream_cmd.guid [9]);
tran (cmdfifo_kdfstream_cmd[13], \cmdfifo_kdfstream_cmd.guid [8]);
tran (cmdfifo_kdfstream_cmd[12], \cmdfifo_kdfstream_cmd.guid [7]);
tran (cmdfifo_kdfstream_cmd[11], \cmdfifo_kdfstream_cmd.guid [6]);
tran (cmdfifo_kdfstream_cmd[10], \cmdfifo_kdfstream_cmd.guid [5]);
tran (cmdfifo_kdfstream_cmd[9], \cmdfifo_kdfstream_cmd.guid [4]);
tran (cmdfifo_kdfstream_cmd[8], \cmdfifo_kdfstream_cmd.guid [3]);
tran (cmdfifo_kdfstream_cmd[7], \cmdfifo_kdfstream_cmd.guid [2]);
tran (cmdfifo_kdfstream_cmd[6], \cmdfifo_kdfstream_cmd.guid [1]);
tran (cmdfifo_kdfstream_cmd[5], \cmdfifo_kdfstream_cmd.guid [0]);
tran (cmdfifo_kdfstream_cmd[4], \cmdfifo_kdfstream_cmd.label_index [2]);
tran (cmdfifo_kdfstream_cmd[3], \cmdfifo_kdfstream_cmd.label_index [1]);
tran (cmdfifo_kdfstream_cmd[2], \cmdfifo_kdfstream_cmd.label_index [0]);
tran (cmdfifo_kdfstream_cmd[1], \cmdfifo_kdfstream_cmd.num_iter [1]);
tran (cmdfifo_kdfstream_cmd[0], \cmdfifo_kdfstream_cmd.num_iter [0]);
tran (\labels[0][0] , \labels[0].delimiter[0] );
tran (\labels[0][1] , \labels[0].delimiter[1] );
tran (\labels[0][2] , \labels[0].delimiter[2] );
tran (\labels[0][3] , \labels[0].delimiter[3] );
tran (\labels[0][4] , \labels[0].delimiter[4] );
tran (\labels[0][5] , \labels[0].delimiter[5] );
tran (\labels[0][6] , \labels[0].delimiter[6] );
tran (\labels[0][7] , \labels[0].delimiter[7] );
tran (\labels[0][8] , \labels[0].delimiter_valid[0] );
tran (\labels[0][9] , \labels[0].label[0] );
tran (\labels[0][10] , \labels[0].label[1] );
tran (\labels[0][11] , \labels[0].label[2] );
tran (\labels[0][12] , \labels[0].label[3] );
tran (\labels[0][13] , \labels[0].label[4] );
tran (\labels[0][14] , \labels[0].label[5] );
tran (\labels[0][15] , \labels[0].label[6] );
tran (\labels[0][16] , \labels[0].label[7] );
tran (\labels[0][17] , \labels[0].label[8] );
tran (\labels[0][18] , \labels[0].label[9] );
tran (\labels[0][19] , \labels[0].label[10] );
tran (\labels[0][20] , \labels[0].label[11] );
tran (\labels[0][21] , \labels[0].label[12] );
tran (\labels[0][22] , \labels[0].label[13] );
tran (\labels[0][23] , \labels[0].label[14] );
tran (\labels[0][24] , \labels[0].label[15] );
tran (\labels[0][25] , \labels[0].label[16] );
tran (\labels[0][26] , \labels[0].label[17] );
tran (\labels[0][27] , \labels[0].label[18] );
tran (\labels[0][28] , \labels[0].label[19] );
tran (\labels[0][29] , \labels[0].label[20] );
tran (\labels[0][30] , \labels[0].label[21] );
tran (\labels[0][31] , \labels[0].label[22] );
tran (\labels[0][32] , \labels[0].label[23] );
tran (\labels[0][33] , \labels[0].label[24] );
tran (\labels[0][34] , \labels[0].label[25] );
tran (\labels[0][35] , \labels[0].label[26] );
tran (\labels[0][36] , \labels[0].label[27] );
tran (\labels[0][37] , \labels[0].label[28] );
tran (\labels[0][38] , \labels[0].label[29] );
tran (\labels[0][39] , \labels[0].label[30] );
tran (\labels[0][40] , \labels[0].label[31] );
tran (\labels[0][41] , \labels[0].label[32] );
tran (\labels[0][42] , \labels[0].label[33] );
tran (\labels[0][43] , \labels[0].label[34] );
tran (\labels[0][44] , \labels[0].label[35] );
tran (\labels[0][45] , \labels[0].label[36] );
tran (\labels[0][46] , \labels[0].label[37] );
tran (\labels[0][47] , \labels[0].label[38] );
tran (\labels[0][48] , \labels[0].label[39] );
tran (\labels[0][49] , \labels[0].label[40] );
tran (\labels[0][50] , \labels[0].label[41] );
tran (\labels[0][51] , \labels[0].label[42] );
tran (\labels[0][52] , \labels[0].label[43] );
tran (\labels[0][53] , \labels[0].label[44] );
tran (\labels[0][54] , \labels[0].label[45] );
tran (\labels[0][55] , \labels[0].label[46] );
tran (\labels[0][56] , \labels[0].label[47] );
tran (\labels[0][57] , \labels[0].label[48] );
tran (\labels[0][58] , \labels[0].label[49] );
tran (\labels[0][59] , \labels[0].label[50] );
tran (\labels[0][60] , \labels[0].label[51] );
tran (\labels[0][61] , \labels[0].label[52] );
tran (\labels[0][62] , \labels[0].label[53] );
tran (\labels[0][63] , \labels[0].label[54] );
tran (\labels[0][64] , \labels[0].label[55] );
tran (\labels[0][65] , \labels[0].label[56] );
tran (\labels[0][66] , \labels[0].label[57] );
tran (\labels[0][67] , \labels[0].label[58] );
tran (\labels[0][68] , \labels[0].label[59] );
tran (\labels[0][69] , \labels[0].label[60] );
tran (\labels[0][70] , \labels[0].label[61] );
tran (\labels[0][71] , \labels[0].label[62] );
tran (\labels[0][72] , \labels[0].label[63] );
tran (\labels[0][73] , \labels[0].label[64] );
tran (\labels[0][74] , \labels[0].label[65] );
tran (\labels[0][75] , \labels[0].label[66] );
tran (\labels[0][76] , \labels[0].label[67] );
tran (\labels[0][77] , \labels[0].label[68] );
tran (\labels[0][78] , \labels[0].label[69] );
tran (\labels[0][79] , \labels[0].label[70] );
tran (\labels[0][80] , \labels[0].label[71] );
tran (\labels[0][81] , \labels[0].label[72] );
tran (\labels[0][82] , \labels[0].label[73] );
tran (\labels[0][83] , \labels[0].label[74] );
tran (\labels[0][84] , \labels[0].label[75] );
tran (\labels[0][85] , \labels[0].label[76] );
tran (\labels[0][86] , \labels[0].label[77] );
tran (\labels[0][87] , \labels[0].label[78] );
tran (\labels[0][88] , \labels[0].label[79] );
tran (\labels[0][89] , \labels[0].label[80] );
tran (\labels[0][90] , \labels[0].label[81] );
tran (\labels[0][91] , \labels[0].label[82] );
tran (\labels[0][92] , \labels[0].label[83] );
tran (\labels[0][93] , \labels[0].label[84] );
tran (\labels[0][94] , \labels[0].label[85] );
tran (\labels[0][95] , \labels[0].label[86] );
tran (\labels[0][96] , \labels[0].label[87] );
tran (\labels[0][97] , \labels[0].label[88] );
tran (\labels[0][98] , \labels[0].label[89] );
tran (\labels[0][99] , \labels[0].label[90] );
tran (\labels[0][100] , \labels[0].label[91] );
tran (\labels[0][101] , \labels[0].label[92] );
tran (\labels[0][102] , \labels[0].label[93] );
tran (\labels[0][103] , \labels[0].label[94] );
tran (\labels[0][104] , \labels[0].label[95] );
tran (\labels[0][105] , \labels[0].label[96] );
tran (\labels[0][106] , \labels[0].label[97] );
tran (\labels[0][107] , \labels[0].label[98] );
tran (\labels[0][108] , \labels[0].label[99] );
tran (\labels[0][109] , \labels[0].label[100] );
tran (\labels[0][110] , \labels[0].label[101] );
tran (\labels[0][111] , \labels[0].label[102] );
tran (\labels[0][112] , \labels[0].label[103] );
tran (\labels[0][113] , \labels[0].label[104] );
tran (\labels[0][114] , \labels[0].label[105] );
tran (\labels[0][115] , \labels[0].label[106] );
tran (\labels[0][116] , \labels[0].label[107] );
tran (\labels[0][117] , \labels[0].label[108] );
tran (\labels[0][118] , \labels[0].label[109] );
tran (\labels[0][119] , \labels[0].label[110] );
tran (\labels[0][120] , \labels[0].label[111] );
tran (\labels[0][121] , \labels[0].label[112] );
tran (\labels[0][122] , \labels[0].label[113] );
tran (\labels[0][123] , \labels[0].label[114] );
tran (\labels[0][124] , \labels[0].label[115] );
tran (\labels[0][125] , \labels[0].label[116] );
tran (\labels[0][126] , \labels[0].label[117] );
tran (\labels[0][127] , \labels[0].label[118] );
tran (\labels[0][128] , \labels[0].label[119] );
tran (\labels[0][129] , \labels[0].label[120] );
tran (\labels[0][130] , \labels[0].label[121] );
tran (\labels[0][131] , \labels[0].label[122] );
tran (\labels[0][132] , \labels[0].label[123] );
tran (\labels[0][133] , \labels[0].label[124] );
tran (\labels[0][134] , \labels[0].label[125] );
tran (\labels[0][135] , \labels[0].label[126] );
tran (\labels[0][136] , \labels[0].label[127] );
tran (\labels[0][137] , \labels[0].label[128] );
tran (\labels[0][138] , \labels[0].label[129] );
tran (\labels[0][139] , \labels[0].label[130] );
tran (\labels[0][140] , \labels[0].label[131] );
tran (\labels[0][141] , \labels[0].label[132] );
tran (\labels[0][142] , \labels[0].label[133] );
tran (\labels[0][143] , \labels[0].label[134] );
tran (\labels[0][144] , \labels[0].label[135] );
tran (\labels[0][145] , \labels[0].label[136] );
tran (\labels[0][146] , \labels[0].label[137] );
tran (\labels[0][147] , \labels[0].label[138] );
tran (\labels[0][148] , \labels[0].label[139] );
tran (\labels[0][149] , \labels[0].label[140] );
tran (\labels[0][150] , \labels[0].label[141] );
tran (\labels[0][151] , \labels[0].label[142] );
tran (\labels[0][152] , \labels[0].label[143] );
tran (\labels[0][153] , \labels[0].label[144] );
tran (\labels[0][154] , \labels[0].label[145] );
tran (\labels[0][155] , \labels[0].label[146] );
tran (\labels[0][156] , \labels[0].label[147] );
tran (\labels[0][157] , \labels[0].label[148] );
tran (\labels[0][158] , \labels[0].label[149] );
tran (\labels[0][159] , \labels[0].label[150] );
tran (\labels[0][160] , \labels[0].label[151] );
tran (\labels[0][161] , \labels[0].label[152] );
tran (\labels[0][162] , \labels[0].label[153] );
tran (\labels[0][163] , \labels[0].label[154] );
tran (\labels[0][164] , \labels[0].label[155] );
tran (\labels[0][165] , \labels[0].label[156] );
tran (\labels[0][166] , \labels[0].label[157] );
tran (\labels[0][167] , \labels[0].label[158] );
tran (\labels[0][168] , \labels[0].label[159] );
tran (\labels[0][169] , \labels[0].label[160] );
tran (\labels[0][170] , \labels[0].label[161] );
tran (\labels[0][171] , \labels[0].label[162] );
tran (\labels[0][172] , \labels[0].label[163] );
tran (\labels[0][173] , \labels[0].label[164] );
tran (\labels[0][174] , \labels[0].label[165] );
tran (\labels[0][175] , \labels[0].label[166] );
tran (\labels[0][176] , \labels[0].label[167] );
tran (\labels[0][177] , \labels[0].label[168] );
tran (\labels[0][178] , \labels[0].label[169] );
tran (\labels[0][179] , \labels[0].label[170] );
tran (\labels[0][180] , \labels[0].label[171] );
tran (\labels[0][181] , \labels[0].label[172] );
tran (\labels[0][182] , \labels[0].label[173] );
tran (\labels[0][183] , \labels[0].label[174] );
tran (\labels[0][184] , \labels[0].label[175] );
tran (\labels[0][185] , \labels[0].label[176] );
tran (\labels[0][186] , \labels[0].label[177] );
tran (\labels[0][187] , \labels[0].label[178] );
tran (\labels[0][188] , \labels[0].label[179] );
tran (\labels[0][189] , \labels[0].label[180] );
tran (\labels[0][190] , \labels[0].label[181] );
tran (\labels[0][191] , \labels[0].label[182] );
tran (\labels[0][192] , \labels[0].label[183] );
tran (\labels[0][193] , \labels[0].label[184] );
tran (\labels[0][194] , \labels[0].label[185] );
tran (\labels[0][195] , \labels[0].label[186] );
tran (\labels[0][196] , \labels[0].label[187] );
tran (\labels[0][197] , \labels[0].label[188] );
tran (\labels[0][198] , \labels[0].label[189] );
tran (\labels[0][199] , \labels[0].label[190] );
tran (\labels[0][200] , \labels[0].label[191] );
tran (\labels[0][201] , \labels[0].label[192] );
tran (\labels[0][202] , \labels[0].label[193] );
tran (\labels[0][203] , \labels[0].label[194] );
tran (\labels[0][204] , \labels[0].label[195] );
tran (\labels[0][205] , \labels[0].label[196] );
tran (\labels[0][206] , \labels[0].label[197] );
tran (\labels[0][207] , \labels[0].label[198] );
tran (\labels[0][208] , \labels[0].label[199] );
tran (\labels[0][209] , \labels[0].label[200] );
tran (\labels[0][210] , \labels[0].label[201] );
tran (\labels[0][211] , \labels[0].label[202] );
tran (\labels[0][212] , \labels[0].label[203] );
tran (\labels[0][213] , \labels[0].label[204] );
tran (\labels[0][214] , \labels[0].label[205] );
tran (\labels[0][215] , \labels[0].label[206] );
tran (\labels[0][216] , \labels[0].label[207] );
tran (\labels[0][217] , \labels[0].label[208] );
tran (\labels[0][218] , \labels[0].label[209] );
tran (\labels[0][219] , \labels[0].label[210] );
tran (\labels[0][220] , \labels[0].label[211] );
tran (\labels[0][221] , \labels[0].label[212] );
tran (\labels[0][222] , \labels[0].label[213] );
tran (\labels[0][223] , \labels[0].label[214] );
tran (\labels[0][224] , \labels[0].label[215] );
tran (\labels[0][225] , \labels[0].label[216] );
tran (\labels[0][226] , \labels[0].label[217] );
tran (\labels[0][227] , \labels[0].label[218] );
tran (\labels[0][228] , \labels[0].label[219] );
tran (\labels[0][229] , \labels[0].label[220] );
tran (\labels[0][230] , \labels[0].label[221] );
tran (\labels[0][231] , \labels[0].label[222] );
tran (\labels[0][232] , \labels[0].label[223] );
tran (\labels[0][233] , \labels[0].label[224] );
tran (\labels[0][234] , \labels[0].label[225] );
tran (\labels[0][235] , \labels[0].label[226] );
tran (\labels[0][236] , \labels[0].label[227] );
tran (\labels[0][237] , \labels[0].label[228] );
tran (\labels[0][238] , \labels[0].label[229] );
tran (\labels[0][239] , \labels[0].label[230] );
tran (\labels[0][240] , \labels[0].label[231] );
tran (\labels[0][241] , \labels[0].label[232] );
tran (\labels[0][242] , \labels[0].label[233] );
tran (\labels[0][243] , \labels[0].label[234] );
tran (\labels[0][244] , \labels[0].label[235] );
tran (\labels[0][245] , \labels[0].label[236] );
tran (\labels[0][246] , \labels[0].label[237] );
tran (\labels[0][247] , \labels[0].label[238] );
tran (\labels[0][248] , \labels[0].label[239] );
tran (\labels[0][249] , \labels[0].label[240] );
tran (\labels[0][250] , \labels[0].label[241] );
tran (\labels[0][251] , \labels[0].label[242] );
tran (\labels[0][252] , \labels[0].label[243] );
tran (\labels[0][253] , \labels[0].label[244] );
tran (\labels[0][254] , \labels[0].label[245] );
tran (\labels[0][255] , \labels[0].label[246] );
tran (\labels[0][256] , \labels[0].label[247] );
tran (\labels[0][257] , \labels[0].label[248] );
tran (\labels[0][258] , \labels[0].label[249] );
tran (\labels[0][259] , \labels[0].label[250] );
tran (\labels[0][260] , \labels[0].label[251] );
tran (\labels[0][261] , \labels[0].label[252] );
tran (\labels[0][262] , \labels[0].label[253] );
tran (\labels[0][263] , \labels[0].label[254] );
tran (\labels[0][264] , \labels[0].label[255] );
tran (\labels[0][265] , \labels[0].label_size[0] );
tran (\labels[0][266] , \labels[0].label_size[1] );
tran (\labels[0][267] , \labels[0].label_size[2] );
tran (\labels[0][268] , \labels[0].label_size[3] );
tran (\labels[0][269] , \labels[0].label_size[4] );
tran (\labels[0][270] , \labels[0].label_size[5] );
tran (\labels[0][271] , \labels[0].guid_size[0] );
tran (\labels[1][0] , \labels[1].delimiter[0] );
tran (\labels[1][1] , \labels[1].delimiter[1] );
tran (\labels[1][2] , \labels[1].delimiter[2] );
tran (\labels[1][3] , \labels[1].delimiter[3] );
tran (\labels[1][4] , \labels[1].delimiter[4] );
tran (\labels[1][5] , \labels[1].delimiter[5] );
tran (\labels[1][6] , \labels[1].delimiter[6] );
tran (\labels[1][7] , \labels[1].delimiter[7] );
tran (\labels[1][8] , \labels[1].delimiter_valid[0] );
tran (\labels[1][9] , \labels[1].label[0] );
tran (\labels[1][10] , \labels[1].label[1] );
tran (\labels[1][11] , \labels[1].label[2] );
tran (\labels[1][12] , \labels[1].label[3] );
tran (\labels[1][13] , \labels[1].label[4] );
tran (\labels[1][14] , \labels[1].label[5] );
tran (\labels[1][15] , \labels[1].label[6] );
tran (\labels[1][16] , \labels[1].label[7] );
tran (\labels[1][17] , \labels[1].label[8] );
tran (\labels[1][18] , \labels[1].label[9] );
tran (\labels[1][19] , \labels[1].label[10] );
tran (\labels[1][20] , \labels[1].label[11] );
tran (\labels[1][21] , \labels[1].label[12] );
tran (\labels[1][22] , \labels[1].label[13] );
tran (\labels[1][23] , \labels[1].label[14] );
tran (\labels[1][24] , \labels[1].label[15] );
tran (\labels[1][25] , \labels[1].label[16] );
tran (\labels[1][26] , \labels[1].label[17] );
tran (\labels[1][27] , \labels[1].label[18] );
tran (\labels[1][28] , \labels[1].label[19] );
tran (\labels[1][29] , \labels[1].label[20] );
tran (\labels[1][30] , \labels[1].label[21] );
tran (\labels[1][31] , \labels[1].label[22] );
tran (\labels[1][32] , \labels[1].label[23] );
tran (\labels[1][33] , \labels[1].label[24] );
tran (\labels[1][34] , \labels[1].label[25] );
tran (\labels[1][35] , \labels[1].label[26] );
tran (\labels[1][36] , \labels[1].label[27] );
tran (\labels[1][37] , \labels[1].label[28] );
tran (\labels[1][38] , \labels[1].label[29] );
tran (\labels[1][39] , \labels[1].label[30] );
tran (\labels[1][40] , \labels[1].label[31] );
tran (\labels[1][41] , \labels[1].label[32] );
tran (\labels[1][42] , \labels[1].label[33] );
tran (\labels[1][43] , \labels[1].label[34] );
tran (\labels[1][44] , \labels[1].label[35] );
tran (\labels[1][45] , \labels[1].label[36] );
tran (\labels[1][46] , \labels[1].label[37] );
tran (\labels[1][47] , \labels[1].label[38] );
tran (\labels[1][48] , \labels[1].label[39] );
tran (\labels[1][49] , \labels[1].label[40] );
tran (\labels[1][50] , \labels[1].label[41] );
tran (\labels[1][51] , \labels[1].label[42] );
tran (\labels[1][52] , \labels[1].label[43] );
tran (\labels[1][53] , \labels[1].label[44] );
tran (\labels[1][54] , \labels[1].label[45] );
tran (\labels[1][55] , \labels[1].label[46] );
tran (\labels[1][56] , \labels[1].label[47] );
tran (\labels[1][57] , \labels[1].label[48] );
tran (\labels[1][58] , \labels[1].label[49] );
tran (\labels[1][59] , \labels[1].label[50] );
tran (\labels[1][60] , \labels[1].label[51] );
tran (\labels[1][61] , \labels[1].label[52] );
tran (\labels[1][62] , \labels[1].label[53] );
tran (\labels[1][63] , \labels[1].label[54] );
tran (\labels[1][64] , \labels[1].label[55] );
tran (\labels[1][65] , \labels[1].label[56] );
tran (\labels[1][66] , \labels[1].label[57] );
tran (\labels[1][67] , \labels[1].label[58] );
tran (\labels[1][68] , \labels[1].label[59] );
tran (\labels[1][69] , \labels[1].label[60] );
tran (\labels[1][70] , \labels[1].label[61] );
tran (\labels[1][71] , \labels[1].label[62] );
tran (\labels[1][72] , \labels[1].label[63] );
tran (\labels[1][73] , \labels[1].label[64] );
tran (\labels[1][74] , \labels[1].label[65] );
tran (\labels[1][75] , \labels[1].label[66] );
tran (\labels[1][76] , \labels[1].label[67] );
tran (\labels[1][77] , \labels[1].label[68] );
tran (\labels[1][78] , \labels[1].label[69] );
tran (\labels[1][79] , \labels[1].label[70] );
tran (\labels[1][80] , \labels[1].label[71] );
tran (\labels[1][81] , \labels[1].label[72] );
tran (\labels[1][82] , \labels[1].label[73] );
tran (\labels[1][83] , \labels[1].label[74] );
tran (\labels[1][84] , \labels[1].label[75] );
tran (\labels[1][85] , \labels[1].label[76] );
tran (\labels[1][86] , \labels[1].label[77] );
tran (\labels[1][87] , \labels[1].label[78] );
tran (\labels[1][88] , \labels[1].label[79] );
tran (\labels[1][89] , \labels[1].label[80] );
tran (\labels[1][90] , \labels[1].label[81] );
tran (\labels[1][91] , \labels[1].label[82] );
tran (\labels[1][92] , \labels[1].label[83] );
tran (\labels[1][93] , \labels[1].label[84] );
tran (\labels[1][94] , \labels[1].label[85] );
tran (\labels[1][95] , \labels[1].label[86] );
tran (\labels[1][96] , \labels[1].label[87] );
tran (\labels[1][97] , \labels[1].label[88] );
tran (\labels[1][98] , \labels[1].label[89] );
tran (\labels[1][99] , \labels[1].label[90] );
tran (\labels[1][100] , \labels[1].label[91] );
tran (\labels[1][101] , \labels[1].label[92] );
tran (\labels[1][102] , \labels[1].label[93] );
tran (\labels[1][103] , \labels[1].label[94] );
tran (\labels[1][104] , \labels[1].label[95] );
tran (\labels[1][105] , \labels[1].label[96] );
tran (\labels[1][106] , \labels[1].label[97] );
tran (\labels[1][107] , \labels[1].label[98] );
tran (\labels[1][108] , \labels[1].label[99] );
tran (\labels[1][109] , \labels[1].label[100] );
tran (\labels[1][110] , \labels[1].label[101] );
tran (\labels[1][111] , \labels[1].label[102] );
tran (\labels[1][112] , \labels[1].label[103] );
tran (\labels[1][113] , \labels[1].label[104] );
tran (\labels[1][114] , \labels[1].label[105] );
tran (\labels[1][115] , \labels[1].label[106] );
tran (\labels[1][116] , \labels[1].label[107] );
tran (\labels[1][117] , \labels[1].label[108] );
tran (\labels[1][118] , \labels[1].label[109] );
tran (\labels[1][119] , \labels[1].label[110] );
tran (\labels[1][120] , \labels[1].label[111] );
tran (\labels[1][121] , \labels[1].label[112] );
tran (\labels[1][122] , \labels[1].label[113] );
tran (\labels[1][123] , \labels[1].label[114] );
tran (\labels[1][124] , \labels[1].label[115] );
tran (\labels[1][125] , \labels[1].label[116] );
tran (\labels[1][126] , \labels[1].label[117] );
tran (\labels[1][127] , \labels[1].label[118] );
tran (\labels[1][128] , \labels[1].label[119] );
tran (\labels[1][129] , \labels[1].label[120] );
tran (\labels[1][130] , \labels[1].label[121] );
tran (\labels[1][131] , \labels[1].label[122] );
tran (\labels[1][132] , \labels[1].label[123] );
tran (\labels[1][133] , \labels[1].label[124] );
tran (\labels[1][134] , \labels[1].label[125] );
tran (\labels[1][135] , \labels[1].label[126] );
tran (\labels[1][136] , \labels[1].label[127] );
tran (\labels[1][137] , \labels[1].label[128] );
tran (\labels[1][138] , \labels[1].label[129] );
tran (\labels[1][139] , \labels[1].label[130] );
tran (\labels[1][140] , \labels[1].label[131] );
tran (\labels[1][141] , \labels[1].label[132] );
tran (\labels[1][142] , \labels[1].label[133] );
tran (\labels[1][143] , \labels[1].label[134] );
tran (\labels[1][144] , \labels[1].label[135] );
tran (\labels[1][145] , \labels[1].label[136] );
tran (\labels[1][146] , \labels[1].label[137] );
tran (\labels[1][147] , \labels[1].label[138] );
tran (\labels[1][148] , \labels[1].label[139] );
tran (\labels[1][149] , \labels[1].label[140] );
tran (\labels[1][150] , \labels[1].label[141] );
tran (\labels[1][151] , \labels[1].label[142] );
tran (\labels[1][152] , \labels[1].label[143] );
tran (\labels[1][153] , \labels[1].label[144] );
tran (\labels[1][154] , \labels[1].label[145] );
tran (\labels[1][155] , \labels[1].label[146] );
tran (\labels[1][156] , \labels[1].label[147] );
tran (\labels[1][157] , \labels[1].label[148] );
tran (\labels[1][158] , \labels[1].label[149] );
tran (\labels[1][159] , \labels[1].label[150] );
tran (\labels[1][160] , \labels[1].label[151] );
tran (\labels[1][161] , \labels[1].label[152] );
tran (\labels[1][162] , \labels[1].label[153] );
tran (\labels[1][163] , \labels[1].label[154] );
tran (\labels[1][164] , \labels[1].label[155] );
tran (\labels[1][165] , \labels[1].label[156] );
tran (\labels[1][166] , \labels[1].label[157] );
tran (\labels[1][167] , \labels[1].label[158] );
tran (\labels[1][168] , \labels[1].label[159] );
tran (\labels[1][169] , \labels[1].label[160] );
tran (\labels[1][170] , \labels[1].label[161] );
tran (\labels[1][171] , \labels[1].label[162] );
tran (\labels[1][172] , \labels[1].label[163] );
tran (\labels[1][173] , \labels[1].label[164] );
tran (\labels[1][174] , \labels[1].label[165] );
tran (\labels[1][175] , \labels[1].label[166] );
tran (\labels[1][176] , \labels[1].label[167] );
tran (\labels[1][177] , \labels[1].label[168] );
tran (\labels[1][178] , \labels[1].label[169] );
tran (\labels[1][179] , \labels[1].label[170] );
tran (\labels[1][180] , \labels[1].label[171] );
tran (\labels[1][181] , \labels[1].label[172] );
tran (\labels[1][182] , \labels[1].label[173] );
tran (\labels[1][183] , \labels[1].label[174] );
tran (\labels[1][184] , \labels[1].label[175] );
tran (\labels[1][185] , \labels[1].label[176] );
tran (\labels[1][186] , \labels[1].label[177] );
tran (\labels[1][187] , \labels[1].label[178] );
tran (\labels[1][188] , \labels[1].label[179] );
tran (\labels[1][189] , \labels[1].label[180] );
tran (\labels[1][190] , \labels[1].label[181] );
tran (\labels[1][191] , \labels[1].label[182] );
tran (\labels[1][192] , \labels[1].label[183] );
tran (\labels[1][193] , \labels[1].label[184] );
tran (\labels[1][194] , \labels[1].label[185] );
tran (\labels[1][195] , \labels[1].label[186] );
tran (\labels[1][196] , \labels[1].label[187] );
tran (\labels[1][197] , \labels[1].label[188] );
tran (\labels[1][198] , \labels[1].label[189] );
tran (\labels[1][199] , \labels[1].label[190] );
tran (\labels[1][200] , \labels[1].label[191] );
tran (\labels[1][201] , \labels[1].label[192] );
tran (\labels[1][202] , \labels[1].label[193] );
tran (\labels[1][203] , \labels[1].label[194] );
tran (\labels[1][204] , \labels[1].label[195] );
tran (\labels[1][205] , \labels[1].label[196] );
tran (\labels[1][206] , \labels[1].label[197] );
tran (\labels[1][207] , \labels[1].label[198] );
tran (\labels[1][208] , \labels[1].label[199] );
tran (\labels[1][209] , \labels[1].label[200] );
tran (\labels[1][210] , \labels[1].label[201] );
tran (\labels[1][211] , \labels[1].label[202] );
tran (\labels[1][212] , \labels[1].label[203] );
tran (\labels[1][213] , \labels[1].label[204] );
tran (\labels[1][214] , \labels[1].label[205] );
tran (\labels[1][215] , \labels[1].label[206] );
tran (\labels[1][216] , \labels[1].label[207] );
tran (\labels[1][217] , \labels[1].label[208] );
tran (\labels[1][218] , \labels[1].label[209] );
tran (\labels[1][219] , \labels[1].label[210] );
tran (\labels[1][220] , \labels[1].label[211] );
tran (\labels[1][221] , \labels[1].label[212] );
tran (\labels[1][222] , \labels[1].label[213] );
tran (\labels[1][223] , \labels[1].label[214] );
tran (\labels[1][224] , \labels[1].label[215] );
tran (\labels[1][225] , \labels[1].label[216] );
tran (\labels[1][226] , \labels[1].label[217] );
tran (\labels[1][227] , \labels[1].label[218] );
tran (\labels[1][228] , \labels[1].label[219] );
tran (\labels[1][229] , \labels[1].label[220] );
tran (\labels[1][230] , \labels[1].label[221] );
tran (\labels[1][231] , \labels[1].label[222] );
tran (\labels[1][232] , \labels[1].label[223] );
tran (\labels[1][233] , \labels[1].label[224] );
tran (\labels[1][234] , \labels[1].label[225] );
tran (\labels[1][235] , \labels[1].label[226] );
tran (\labels[1][236] , \labels[1].label[227] );
tran (\labels[1][237] , \labels[1].label[228] );
tran (\labels[1][238] , \labels[1].label[229] );
tran (\labels[1][239] , \labels[1].label[230] );
tran (\labels[1][240] , \labels[1].label[231] );
tran (\labels[1][241] , \labels[1].label[232] );
tran (\labels[1][242] , \labels[1].label[233] );
tran (\labels[1][243] , \labels[1].label[234] );
tran (\labels[1][244] , \labels[1].label[235] );
tran (\labels[1][245] , \labels[1].label[236] );
tran (\labels[1][246] , \labels[1].label[237] );
tran (\labels[1][247] , \labels[1].label[238] );
tran (\labels[1][248] , \labels[1].label[239] );
tran (\labels[1][249] , \labels[1].label[240] );
tran (\labels[1][250] , \labels[1].label[241] );
tran (\labels[1][251] , \labels[1].label[242] );
tran (\labels[1][252] , \labels[1].label[243] );
tran (\labels[1][253] , \labels[1].label[244] );
tran (\labels[1][254] , \labels[1].label[245] );
tran (\labels[1][255] , \labels[1].label[246] );
tran (\labels[1][256] , \labels[1].label[247] );
tran (\labels[1][257] , \labels[1].label[248] );
tran (\labels[1][258] , \labels[1].label[249] );
tran (\labels[1][259] , \labels[1].label[250] );
tran (\labels[1][260] , \labels[1].label[251] );
tran (\labels[1][261] , \labels[1].label[252] );
tran (\labels[1][262] , \labels[1].label[253] );
tran (\labels[1][263] , \labels[1].label[254] );
tran (\labels[1][264] , \labels[1].label[255] );
tran (\labels[1][265] , \labels[1].label_size[0] );
tran (\labels[1][266] , \labels[1].label_size[1] );
tran (\labels[1][267] , \labels[1].label_size[2] );
tran (\labels[1][268] , \labels[1].label_size[3] );
tran (\labels[1][269] , \labels[1].label_size[4] );
tran (\labels[1][270] , \labels[1].label_size[5] );
tran (\labels[1][271] , \labels[1].guid_size[0] );
tran (\labels[2][0] , \labels[2].delimiter[0] );
tran (\labels[2][1] , \labels[2].delimiter[1] );
tran (\labels[2][2] , \labels[2].delimiter[2] );
tran (\labels[2][3] , \labels[2].delimiter[3] );
tran (\labels[2][4] , \labels[2].delimiter[4] );
tran (\labels[2][5] , \labels[2].delimiter[5] );
tran (\labels[2][6] , \labels[2].delimiter[6] );
tran (\labels[2][7] , \labels[2].delimiter[7] );
tran (\labels[2][8] , \labels[2].delimiter_valid[0] );
tran (\labels[2][9] , \labels[2].label[0] );
tran (\labels[2][10] , \labels[2].label[1] );
tran (\labels[2][11] , \labels[2].label[2] );
tran (\labels[2][12] , \labels[2].label[3] );
tran (\labels[2][13] , \labels[2].label[4] );
tran (\labels[2][14] , \labels[2].label[5] );
tran (\labels[2][15] , \labels[2].label[6] );
tran (\labels[2][16] , \labels[2].label[7] );
tran (\labels[2][17] , \labels[2].label[8] );
tran (\labels[2][18] , \labels[2].label[9] );
tran (\labels[2][19] , \labels[2].label[10] );
tran (\labels[2][20] , \labels[2].label[11] );
tran (\labels[2][21] , \labels[2].label[12] );
tran (\labels[2][22] , \labels[2].label[13] );
tran (\labels[2][23] , \labels[2].label[14] );
tran (\labels[2][24] , \labels[2].label[15] );
tran (\labels[2][25] , \labels[2].label[16] );
tran (\labels[2][26] , \labels[2].label[17] );
tran (\labels[2][27] , \labels[2].label[18] );
tran (\labels[2][28] , \labels[2].label[19] );
tran (\labels[2][29] , \labels[2].label[20] );
tran (\labels[2][30] , \labels[2].label[21] );
tran (\labels[2][31] , \labels[2].label[22] );
tran (\labels[2][32] , \labels[2].label[23] );
tran (\labels[2][33] , \labels[2].label[24] );
tran (\labels[2][34] , \labels[2].label[25] );
tran (\labels[2][35] , \labels[2].label[26] );
tran (\labels[2][36] , \labels[2].label[27] );
tran (\labels[2][37] , \labels[2].label[28] );
tran (\labels[2][38] , \labels[2].label[29] );
tran (\labels[2][39] , \labels[2].label[30] );
tran (\labels[2][40] , \labels[2].label[31] );
tran (\labels[2][41] , \labels[2].label[32] );
tran (\labels[2][42] , \labels[2].label[33] );
tran (\labels[2][43] , \labels[2].label[34] );
tran (\labels[2][44] , \labels[2].label[35] );
tran (\labels[2][45] , \labels[2].label[36] );
tran (\labels[2][46] , \labels[2].label[37] );
tran (\labels[2][47] , \labels[2].label[38] );
tran (\labels[2][48] , \labels[2].label[39] );
tran (\labels[2][49] , \labels[2].label[40] );
tran (\labels[2][50] , \labels[2].label[41] );
tran (\labels[2][51] , \labels[2].label[42] );
tran (\labels[2][52] , \labels[2].label[43] );
tran (\labels[2][53] , \labels[2].label[44] );
tran (\labels[2][54] , \labels[2].label[45] );
tran (\labels[2][55] , \labels[2].label[46] );
tran (\labels[2][56] , \labels[2].label[47] );
tran (\labels[2][57] , \labels[2].label[48] );
tran (\labels[2][58] , \labels[2].label[49] );
tran (\labels[2][59] , \labels[2].label[50] );
tran (\labels[2][60] , \labels[2].label[51] );
tran (\labels[2][61] , \labels[2].label[52] );
tran (\labels[2][62] , \labels[2].label[53] );
tran (\labels[2][63] , \labels[2].label[54] );
tran (\labels[2][64] , \labels[2].label[55] );
tran (\labels[2][65] , \labels[2].label[56] );
tran (\labels[2][66] , \labels[2].label[57] );
tran (\labels[2][67] , \labels[2].label[58] );
tran (\labels[2][68] , \labels[2].label[59] );
tran (\labels[2][69] , \labels[2].label[60] );
tran (\labels[2][70] , \labels[2].label[61] );
tran (\labels[2][71] , \labels[2].label[62] );
tran (\labels[2][72] , \labels[2].label[63] );
tran (\labels[2][73] , \labels[2].label[64] );
tran (\labels[2][74] , \labels[2].label[65] );
tran (\labels[2][75] , \labels[2].label[66] );
tran (\labels[2][76] , \labels[2].label[67] );
tran (\labels[2][77] , \labels[2].label[68] );
tran (\labels[2][78] , \labels[2].label[69] );
tran (\labels[2][79] , \labels[2].label[70] );
tran (\labels[2][80] , \labels[2].label[71] );
tran (\labels[2][81] , \labels[2].label[72] );
tran (\labels[2][82] , \labels[2].label[73] );
tran (\labels[2][83] , \labels[2].label[74] );
tran (\labels[2][84] , \labels[2].label[75] );
tran (\labels[2][85] , \labels[2].label[76] );
tran (\labels[2][86] , \labels[2].label[77] );
tran (\labels[2][87] , \labels[2].label[78] );
tran (\labels[2][88] , \labels[2].label[79] );
tran (\labels[2][89] , \labels[2].label[80] );
tran (\labels[2][90] , \labels[2].label[81] );
tran (\labels[2][91] , \labels[2].label[82] );
tran (\labels[2][92] , \labels[2].label[83] );
tran (\labels[2][93] , \labels[2].label[84] );
tran (\labels[2][94] , \labels[2].label[85] );
tran (\labels[2][95] , \labels[2].label[86] );
tran (\labels[2][96] , \labels[2].label[87] );
tran (\labels[2][97] , \labels[2].label[88] );
tran (\labels[2][98] , \labels[2].label[89] );
tran (\labels[2][99] , \labels[2].label[90] );
tran (\labels[2][100] , \labels[2].label[91] );
tran (\labels[2][101] , \labels[2].label[92] );
tran (\labels[2][102] , \labels[2].label[93] );
tran (\labels[2][103] , \labels[2].label[94] );
tran (\labels[2][104] , \labels[2].label[95] );
tran (\labels[2][105] , \labels[2].label[96] );
tran (\labels[2][106] , \labels[2].label[97] );
tran (\labels[2][107] , \labels[2].label[98] );
tran (\labels[2][108] , \labels[2].label[99] );
tran (\labels[2][109] , \labels[2].label[100] );
tran (\labels[2][110] , \labels[2].label[101] );
tran (\labels[2][111] , \labels[2].label[102] );
tran (\labels[2][112] , \labels[2].label[103] );
tran (\labels[2][113] , \labels[2].label[104] );
tran (\labels[2][114] , \labels[2].label[105] );
tran (\labels[2][115] , \labels[2].label[106] );
tran (\labels[2][116] , \labels[2].label[107] );
tran (\labels[2][117] , \labels[2].label[108] );
tran (\labels[2][118] , \labels[2].label[109] );
tran (\labels[2][119] , \labels[2].label[110] );
tran (\labels[2][120] , \labels[2].label[111] );
tran (\labels[2][121] , \labels[2].label[112] );
tran (\labels[2][122] , \labels[2].label[113] );
tran (\labels[2][123] , \labels[2].label[114] );
tran (\labels[2][124] , \labels[2].label[115] );
tran (\labels[2][125] , \labels[2].label[116] );
tran (\labels[2][126] , \labels[2].label[117] );
tran (\labels[2][127] , \labels[2].label[118] );
tran (\labels[2][128] , \labels[2].label[119] );
tran (\labels[2][129] , \labels[2].label[120] );
tran (\labels[2][130] , \labels[2].label[121] );
tran (\labels[2][131] , \labels[2].label[122] );
tran (\labels[2][132] , \labels[2].label[123] );
tran (\labels[2][133] , \labels[2].label[124] );
tran (\labels[2][134] , \labels[2].label[125] );
tran (\labels[2][135] , \labels[2].label[126] );
tran (\labels[2][136] , \labels[2].label[127] );
tran (\labels[2][137] , \labels[2].label[128] );
tran (\labels[2][138] , \labels[2].label[129] );
tran (\labels[2][139] , \labels[2].label[130] );
tran (\labels[2][140] , \labels[2].label[131] );
tran (\labels[2][141] , \labels[2].label[132] );
tran (\labels[2][142] , \labels[2].label[133] );
tran (\labels[2][143] , \labels[2].label[134] );
tran (\labels[2][144] , \labels[2].label[135] );
tran (\labels[2][145] , \labels[2].label[136] );
tran (\labels[2][146] , \labels[2].label[137] );
tran (\labels[2][147] , \labels[2].label[138] );
tran (\labels[2][148] , \labels[2].label[139] );
tran (\labels[2][149] , \labels[2].label[140] );
tran (\labels[2][150] , \labels[2].label[141] );
tran (\labels[2][151] , \labels[2].label[142] );
tran (\labels[2][152] , \labels[2].label[143] );
tran (\labels[2][153] , \labels[2].label[144] );
tran (\labels[2][154] , \labels[2].label[145] );
tran (\labels[2][155] , \labels[2].label[146] );
tran (\labels[2][156] , \labels[2].label[147] );
tran (\labels[2][157] , \labels[2].label[148] );
tran (\labels[2][158] , \labels[2].label[149] );
tran (\labels[2][159] , \labels[2].label[150] );
tran (\labels[2][160] , \labels[2].label[151] );
tran (\labels[2][161] , \labels[2].label[152] );
tran (\labels[2][162] , \labels[2].label[153] );
tran (\labels[2][163] , \labels[2].label[154] );
tran (\labels[2][164] , \labels[2].label[155] );
tran (\labels[2][165] , \labels[2].label[156] );
tran (\labels[2][166] , \labels[2].label[157] );
tran (\labels[2][167] , \labels[2].label[158] );
tran (\labels[2][168] , \labels[2].label[159] );
tran (\labels[2][169] , \labels[2].label[160] );
tran (\labels[2][170] , \labels[2].label[161] );
tran (\labels[2][171] , \labels[2].label[162] );
tran (\labels[2][172] , \labels[2].label[163] );
tran (\labels[2][173] , \labels[2].label[164] );
tran (\labels[2][174] , \labels[2].label[165] );
tran (\labels[2][175] , \labels[2].label[166] );
tran (\labels[2][176] , \labels[2].label[167] );
tran (\labels[2][177] , \labels[2].label[168] );
tran (\labels[2][178] , \labels[2].label[169] );
tran (\labels[2][179] , \labels[2].label[170] );
tran (\labels[2][180] , \labels[2].label[171] );
tran (\labels[2][181] , \labels[2].label[172] );
tran (\labels[2][182] , \labels[2].label[173] );
tran (\labels[2][183] , \labels[2].label[174] );
tran (\labels[2][184] , \labels[2].label[175] );
tran (\labels[2][185] , \labels[2].label[176] );
tran (\labels[2][186] , \labels[2].label[177] );
tran (\labels[2][187] , \labels[2].label[178] );
tran (\labels[2][188] , \labels[2].label[179] );
tran (\labels[2][189] , \labels[2].label[180] );
tran (\labels[2][190] , \labels[2].label[181] );
tran (\labels[2][191] , \labels[2].label[182] );
tran (\labels[2][192] , \labels[2].label[183] );
tran (\labels[2][193] , \labels[2].label[184] );
tran (\labels[2][194] , \labels[2].label[185] );
tran (\labels[2][195] , \labels[2].label[186] );
tran (\labels[2][196] , \labels[2].label[187] );
tran (\labels[2][197] , \labels[2].label[188] );
tran (\labels[2][198] , \labels[2].label[189] );
tran (\labels[2][199] , \labels[2].label[190] );
tran (\labels[2][200] , \labels[2].label[191] );
tran (\labels[2][201] , \labels[2].label[192] );
tran (\labels[2][202] , \labels[2].label[193] );
tran (\labels[2][203] , \labels[2].label[194] );
tran (\labels[2][204] , \labels[2].label[195] );
tran (\labels[2][205] , \labels[2].label[196] );
tran (\labels[2][206] , \labels[2].label[197] );
tran (\labels[2][207] , \labels[2].label[198] );
tran (\labels[2][208] , \labels[2].label[199] );
tran (\labels[2][209] , \labels[2].label[200] );
tran (\labels[2][210] , \labels[2].label[201] );
tran (\labels[2][211] , \labels[2].label[202] );
tran (\labels[2][212] , \labels[2].label[203] );
tran (\labels[2][213] , \labels[2].label[204] );
tran (\labels[2][214] , \labels[2].label[205] );
tran (\labels[2][215] , \labels[2].label[206] );
tran (\labels[2][216] , \labels[2].label[207] );
tran (\labels[2][217] , \labels[2].label[208] );
tran (\labels[2][218] , \labels[2].label[209] );
tran (\labels[2][219] , \labels[2].label[210] );
tran (\labels[2][220] , \labels[2].label[211] );
tran (\labels[2][221] , \labels[2].label[212] );
tran (\labels[2][222] , \labels[2].label[213] );
tran (\labels[2][223] , \labels[2].label[214] );
tran (\labels[2][224] , \labels[2].label[215] );
tran (\labels[2][225] , \labels[2].label[216] );
tran (\labels[2][226] , \labels[2].label[217] );
tran (\labels[2][227] , \labels[2].label[218] );
tran (\labels[2][228] , \labels[2].label[219] );
tran (\labels[2][229] , \labels[2].label[220] );
tran (\labels[2][230] , \labels[2].label[221] );
tran (\labels[2][231] , \labels[2].label[222] );
tran (\labels[2][232] , \labels[2].label[223] );
tran (\labels[2][233] , \labels[2].label[224] );
tran (\labels[2][234] , \labels[2].label[225] );
tran (\labels[2][235] , \labels[2].label[226] );
tran (\labels[2][236] , \labels[2].label[227] );
tran (\labels[2][237] , \labels[2].label[228] );
tran (\labels[2][238] , \labels[2].label[229] );
tran (\labels[2][239] , \labels[2].label[230] );
tran (\labels[2][240] , \labels[2].label[231] );
tran (\labels[2][241] , \labels[2].label[232] );
tran (\labels[2][242] , \labels[2].label[233] );
tran (\labels[2][243] , \labels[2].label[234] );
tran (\labels[2][244] , \labels[2].label[235] );
tran (\labels[2][245] , \labels[2].label[236] );
tran (\labels[2][246] , \labels[2].label[237] );
tran (\labels[2][247] , \labels[2].label[238] );
tran (\labels[2][248] , \labels[2].label[239] );
tran (\labels[2][249] , \labels[2].label[240] );
tran (\labels[2][250] , \labels[2].label[241] );
tran (\labels[2][251] , \labels[2].label[242] );
tran (\labels[2][252] , \labels[2].label[243] );
tran (\labels[2][253] , \labels[2].label[244] );
tran (\labels[2][254] , \labels[2].label[245] );
tran (\labels[2][255] , \labels[2].label[246] );
tran (\labels[2][256] , \labels[2].label[247] );
tran (\labels[2][257] , \labels[2].label[248] );
tran (\labels[2][258] , \labels[2].label[249] );
tran (\labels[2][259] , \labels[2].label[250] );
tran (\labels[2][260] , \labels[2].label[251] );
tran (\labels[2][261] , \labels[2].label[252] );
tran (\labels[2][262] , \labels[2].label[253] );
tran (\labels[2][263] , \labels[2].label[254] );
tran (\labels[2][264] , \labels[2].label[255] );
tran (\labels[2][265] , \labels[2].label_size[0] );
tran (\labels[2][266] , \labels[2].label_size[1] );
tran (\labels[2][267] , \labels[2].label_size[2] );
tran (\labels[2][268] , \labels[2].label_size[3] );
tran (\labels[2][269] , \labels[2].label_size[4] );
tran (\labels[2][270] , \labels[2].label_size[5] );
tran (\labels[2][271] , \labels[2].guid_size[0] );
tran (\labels[3][0] , \labels[3].delimiter[0] );
tran (\labels[3][1] , \labels[3].delimiter[1] );
tran (\labels[3][2] , \labels[3].delimiter[2] );
tran (\labels[3][3] , \labels[3].delimiter[3] );
tran (\labels[3][4] , \labels[3].delimiter[4] );
tran (\labels[3][5] , \labels[3].delimiter[5] );
tran (\labels[3][6] , \labels[3].delimiter[6] );
tran (\labels[3][7] , \labels[3].delimiter[7] );
tran (\labels[3][8] , \labels[3].delimiter_valid[0] );
tran (\labels[3][9] , \labels[3].label[0] );
tran (\labels[3][10] , \labels[3].label[1] );
tran (\labels[3][11] , \labels[3].label[2] );
tran (\labels[3][12] , \labels[3].label[3] );
tran (\labels[3][13] , \labels[3].label[4] );
tran (\labels[3][14] , \labels[3].label[5] );
tran (\labels[3][15] , \labels[3].label[6] );
tran (\labels[3][16] , \labels[3].label[7] );
tran (\labels[3][17] , \labels[3].label[8] );
tran (\labels[3][18] , \labels[3].label[9] );
tran (\labels[3][19] , \labels[3].label[10] );
tran (\labels[3][20] , \labels[3].label[11] );
tran (\labels[3][21] , \labels[3].label[12] );
tran (\labels[3][22] , \labels[3].label[13] );
tran (\labels[3][23] , \labels[3].label[14] );
tran (\labels[3][24] , \labels[3].label[15] );
tran (\labels[3][25] , \labels[3].label[16] );
tran (\labels[3][26] , \labels[3].label[17] );
tran (\labels[3][27] , \labels[3].label[18] );
tran (\labels[3][28] , \labels[3].label[19] );
tran (\labels[3][29] , \labels[3].label[20] );
tran (\labels[3][30] , \labels[3].label[21] );
tran (\labels[3][31] , \labels[3].label[22] );
tran (\labels[3][32] , \labels[3].label[23] );
tran (\labels[3][33] , \labels[3].label[24] );
tran (\labels[3][34] , \labels[3].label[25] );
tran (\labels[3][35] , \labels[3].label[26] );
tran (\labels[3][36] , \labels[3].label[27] );
tran (\labels[3][37] , \labels[3].label[28] );
tran (\labels[3][38] , \labels[3].label[29] );
tran (\labels[3][39] , \labels[3].label[30] );
tran (\labels[3][40] , \labels[3].label[31] );
tran (\labels[3][41] , \labels[3].label[32] );
tran (\labels[3][42] , \labels[3].label[33] );
tran (\labels[3][43] , \labels[3].label[34] );
tran (\labels[3][44] , \labels[3].label[35] );
tran (\labels[3][45] , \labels[3].label[36] );
tran (\labels[3][46] , \labels[3].label[37] );
tran (\labels[3][47] , \labels[3].label[38] );
tran (\labels[3][48] , \labels[3].label[39] );
tran (\labels[3][49] , \labels[3].label[40] );
tran (\labels[3][50] , \labels[3].label[41] );
tran (\labels[3][51] , \labels[3].label[42] );
tran (\labels[3][52] , \labels[3].label[43] );
tran (\labels[3][53] , \labels[3].label[44] );
tran (\labels[3][54] , \labels[3].label[45] );
tran (\labels[3][55] , \labels[3].label[46] );
tran (\labels[3][56] , \labels[3].label[47] );
tran (\labels[3][57] , \labels[3].label[48] );
tran (\labels[3][58] , \labels[3].label[49] );
tran (\labels[3][59] , \labels[3].label[50] );
tran (\labels[3][60] , \labels[3].label[51] );
tran (\labels[3][61] , \labels[3].label[52] );
tran (\labels[3][62] , \labels[3].label[53] );
tran (\labels[3][63] , \labels[3].label[54] );
tran (\labels[3][64] , \labels[3].label[55] );
tran (\labels[3][65] , \labels[3].label[56] );
tran (\labels[3][66] , \labels[3].label[57] );
tran (\labels[3][67] , \labels[3].label[58] );
tran (\labels[3][68] , \labels[3].label[59] );
tran (\labels[3][69] , \labels[3].label[60] );
tran (\labels[3][70] , \labels[3].label[61] );
tran (\labels[3][71] , \labels[3].label[62] );
tran (\labels[3][72] , \labels[3].label[63] );
tran (\labels[3][73] , \labels[3].label[64] );
tran (\labels[3][74] , \labels[3].label[65] );
tran (\labels[3][75] , \labels[3].label[66] );
tran (\labels[3][76] , \labels[3].label[67] );
tran (\labels[3][77] , \labels[3].label[68] );
tran (\labels[3][78] , \labels[3].label[69] );
tran (\labels[3][79] , \labels[3].label[70] );
tran (\labels[3][80] , \labels[3].label[71] );
tran (\labels[3][81] , \labels[3].label[72] );
tran (\labels[3][82] , \labels[3].label[73] );
tran (\labels[3][83] , \labels[3].label[74] );
tran (\labels[3][84] , \labels[3].label[75] );
tran (\labels[3][85] , \labels[3].label[76] );
tran (\labels[3][86] , \labels[3].label[77] );
tran (\labels[3][87] , \labels[3].label[78] );
tran (\labels[3][88] , \labels[3].label[79] );
tran (\labels[3][89] , \labels[3].label[80] );
tran (\labels[3][90] , \labels[3].label[81] );
tran (\labels[3][91] , \labels[3].label[82] );
tran (\labels[3][92] , \labels[3].label[83] );
tran (\labels[3][93] , \labels[3].label[84] );
tran (\labels[3][94] , \labels[3].label[85] );
tran (\labels[3][95] , \labels[3].label[86] );
tran (\labels[3][96] , \labels[3].label[87] );
tran (\labels[3][97] , \labels[3].label[88] );
tran (\labels[3][98] , \labels[3].label[89] );
tran (\labels[3][99] , \labels[3].label[90] );
tran (\labels[3][100] , \labels[3].label[91] );
tran (\labels[3][101] , \labels[3].label[92] );
tran (\labels[3][102] , \labels[3].label[93] );
tran (\labels[3][103] , \labels[3].label[94] );
tran (\labels[3][104] , \labels[3].label[95] );
tran (\labels[3][105] , \labels[3].label[96] );
tran (\labels[3][106] , \labels[3].label[97] );
tran (\labels[3][107] , \labels[3].label[98] );
tran (\labels[3][108] , \labels[3].label[99] );
tran (\labels[3][109] , \labels[3].label[100] );
tran (\labels[3][110] , \labels[3].label[101] );
tran (\labels[3][111] , \labels[3].label[102] );
tran (\labels[3][112] , \labels[3].label[103] );
tran (\labels[3][113] , \labels[3].label[104] );
tran (\labels[3][114] , \labels[3].label[105] );
tran (\labels[3][115] , \labels[3].label[106] );
tran (\labels[3][116] , \labels[3].label[107] );
tran (\labels[3][117] , \labels[3].label[108] );
tran (\labels[3][118] , \labels[3].label[109] );
tran (\labels[3][119] , \labels[3].label[110] );
tran (\labels[3][120] , \labels[3].label[111] );
tran (\labels[3][121] , \labels[3].label[112] );
tran (\labels[3][122] , \labels[3].label[113] );
tran (\labels[3][123] , \labels[3].label[114] );
tran (\labels[3][124] , \labels[3].label[115] );
tran (\labels[3][125] , \labels[3].label[116] );
tran (\labels[3][126] , \labels[3].label[117] );
tran (\labels[3][127] , \labels[3].label[118] );
tran (\labels[3][128] , \labels[3].label[119] );
tran (\labels[3][129] , \labels[3].label[120] );
tran (\labels[3][130] , \labels[3].label[121] );
tran (\labels[3][131] , \labels[3].label[122] );
tran (\labels[3][132] , \labels[3].label[123] );
tran (\labels[3][133] , \labels[3].label[124] );
tran (\labels[3][134] , \labels[3].label[125] );
tran (\labels[3][135] , \labels[3].label[126] );
tran (\labels[3][136] , \labels[3].label[127] );
tran (\labels[3][137] , \labels[3].label[128] );
tran (\labels[3][138] , \labels[3].label[129] );
tran (\labels[3][139] , \labels[3].label[130] );
tran (\labels[3][140] , \labels[3].label[131] );
tran (\labels[3][141] , \labels[3].label[132] );
tran (\labels[3][142] , \labels[3].label[133] );
tran (\labels[3][143] , \labels[3].label[134] );
tran (\labels[3][144] , \labels[3].label[135] );
tran (\labels[3][145] , \labels[3].label[136] );
tran (\labels[3][146] , \labels[3].label[137] );
tran (\labels[3][147] , \labels[3].label[138] );
tran (\labels[3][148] , \labels[3].label[139] );
tran (\labels[3][149] , \labels[3].label[140] );
tran (\labels[3][150] , \labels[3].label[141] );
tran (\labels[3][151] , \labels[3].label[142] );
tran (\labels[3][152] , \labels[3].label[143] );
tran (\labels[3][153] , \labels[3].label[144] );
tran (\labels[3][154] , \labels[3].label[145] );
tran (\labels[3][155] , \labels[3].label[146] );
tran (\labels[3][156] , \labels[3].label[147] );
tran (\labels[3][157] , \labels[3].label[148] );
tran (\labels[3][158] , \labels[3].label[149] );
tran (\labels[3][159] , \labels[3].label[150] );
tran (\labels[3][160] , \labels[3].label[151] );
tran (\labels[3][161] , \labels[3].label[152] );
tran (\labels[3][162] , \labels[3].label[153] );
tran (\labels[3][163] , \labels[3].label[154] );
tran (\labels[3][164] , \labels[3].label[155] );
tran (\labels[3][165] , \labels[3].label[156] );
tran (\labels[3][166] , \labels[3].label[157] );
tran (\labels[3][167] , \labels[3].label[158] );
tran (\labels[3][168] , \labels[3].label[159] );
tran (\labels[3][169] , \labels[3].label[160] );
tran (\labels[3][170] , \labels[3].label[161] );
tran (\labels[3][171] , \labels[3].label[162] );
tran (\labels[3][172] , \labels[3].label[163] );
tran (\labels[3][173] , \labels[3].label[164] );
tran (\labels[3][174] , \labels[3].label[165] );
tran (\labels[3][175] , \labels[3].label[166] );
tran (\labels[3][176] , \labels[3].label[167] );
tran (\labels[3][177] , \labels[3].label[168] );
tran (\labels[3][178] , \labels[3].label[169] );
tran (\labels[3][179] , \labels[3].label[170] );
tran (\labels[3][180] , \labels[3].label[171] );
tran (\labels[3][181] , \labels[3].label[172] );
tran (\labels[3][182] , \labels[3].label[173] );
tran (\labels[3][183] , \labels[3].label[174] );
tran (\labels[3][184] , \labels[3].label[175] );
tran (\labels[3][185] , \labels[3].label[176] );
tran (\labels[3][186] , \labels[3].label[177] );
tran (\labels[3][187] , \labels[3].label[178] );
tran (\labels[3][188] , \labels[3].label[179] );
tran (\labels[3][189] , \labels[3].label[180] );
tran (\labels[3][190] , \labels[3].label[181] );
tran (\labels[3][191] , \labels[3].label[182] );
tran (\labels[3][192] , \labels[3].label[183] );
tran (\labels[3][193] , \labels[3].label[184] );
tran (\labels[3][194] , \labels[3].label[185] );
tran (\labels[3][195] , \labels[3].label[186] );
tran (\labels[3][196] , \labels[3].label[187] );
tran (\labels[3][197] , \labels[3].label[188] );
tran (\labels[3][198] , \labels[3].label[189] );
tran (\labels[3][199] , \labels[3].label[190] );
tran (\labels[3][200] , \labels[3].label[191] );
tran (\labels[3][201] , \labels[3].label[192] );
tran (\labels[3][202] , \labels[3].label[193] );
tran (\labels[3][203] , \labels[3].label[194] );
tran (\labels[3][204] , \labels[3].label[195] );
tran (\labels[3][205] , \labels[3].label[196] );
tran (\labels[3][206] , \labels[3].label[197] );
tran (\labels[3][207] , \labels[3].label[198] );
tran (\labels[3][208] , \labels[3].label[199] );
tran (\labels[3][209] , \labels[3].label[200] );
tran (\labels[3][210] , \labels[3].label[201] );
tran (\labels[3][211] , \labels[3].label[202] );
tran (\labels[3][212] , \labels[3].label[203] );
tran (\labels[3][213] , \labels[3].label[204] );
tran (\labels[3][214] , \labels[3].label[205] );
tran (\labels[3][215] , \labels[3].label[206] );
tran (\labels[3][216] , \labels[3].label[207] );
tran (\labels[3][217] , \labels[3].label[208] );
tran (\labels[3][218] , \labels[3].label[209] );
tran (\labels[3][219] , \labels[3].label[210] );
tran (\labels[3][220] , \labels[3].label[211] );
tran (\labels[3][221] , \labels[3].label[212] );
tran (\labels[3][222] , \labels[3].label[213] );
tran (\labels[3][223] , \labels[3].label[214] );
tran (\labels[3][224] , \labels[3].label[215] );
tran (\labels[3][225] , \labels[3].label[216] );
tran (\labels[3][226] , \labels[3].label[217] );
tran (\labels[3][227] , \labels[3].label[218] );
tran (\labels[3][228] , \labels[3].label[219] );
tran (\labels[3][229] , \labels[3].label[220] );
tran (\labels[3][230] , \labels[3].label[221] );
tran (\labels[3][231] , \labels[3].label[222] );
tran (\labels[3][232] , \labels[3].label[223] );
tran (\labels[3][233] , \labels[3].label[224] );
tran (\labels[3][234] , \labels[3].label[225] );
tran (\labels[3][235] , \labels[3].label[226] );
tran (\labels[3][236] , \labels[3].label[227] );
tran (\labels[3][237] , \labels[3].label[228] );
tran (\labels[3][238] , \labels[3].label[229] );
tran (\labels[3][239] , \labels[3].label[230] );
tran (\labels[3][240] , \labels[3].label[231] );
tran (\labels[3][241] , \labels[3].label[232] );
tran (\labels[3][242] , \labels[3].label[233] );
tran (\labels[3][243] , \labels[3].label[234] );
tran (\labels[3][244] , \labels[3].label[235] );
tran (\labels[3][245] , \labels[3].label[236] );
tran (\labels[3][246] , \labels[3].label[237] );
tran (\labels[3][247] , \labels[3].label[238] );
tran (\labels[3][248] , \labels[3].label[239] );
tran (\labels[3][249] , \labels[3].label[240] );
tran (\labels[3][250] , \labels[3].label[241] );
tran (\labels[3][251] , \labels[3].label[242] );
tran (\labels[3][252] , \labels[3].label[243] );
tran (\labels[3][253] , \labels[3].label[244] );
tran (\labels[3][254] , \labels[3].label[245] );
tran (\labels[3][255] , \labels[3].label[246] );
tran (\labels[3][256] , \labels[3].label[247] );
tran (\labels[3][257] , \labels[3].label[248] );
tran (\labels[3][258] , \labels[3].label[249] );
tran (\labels[3][259] , \labels[3].label[250] );
tran (\labels[3][260] , \labels[3].label[251] );
tran (\labels[3][261] , \labels[3].label[252] );
tran (\labels[3][262] , \labels[3].label[253] );
tran (\labels[3][263] , \labels[3].label[254] );
tran (\labels[3][264] , \labels[3].label[255] );
tran (\labels[3][265] , \labels[3].label_size[0] );
tran (\labels[3][266] , \labels[3].label_size[1] );
tran (\labels[3][267] , \labels[3].label_size[2] );
tran (\labels[3][268] , \labels[3].label_size[3] );
tran (\labels[3][269] , \labels[3].label_size[4] );
tran (\labels[3][270] , \labels[3].label_size[5] );
tran (\labels[3][271] , \labels[3].guid_size[0] );
tran (\labels[4][0] , \labels[4].delimiter[0] );
tran (\labels[4][1] , \labels[4].delimiter[1] );
tran (\labels[4][2] , \labels[4].delimiter[2] );
tran (\labels[4][3] , \labels[4].delimiter[3] );
tran (\labels[4][4] , \labels[4].delimiter[4] );
tran (\labels[4][5] , \labels[4].delimiter[5] );
tran (\labels[4][6] , \labels[4].delimiter[6] );
tran (\labels[4][7] , \labels[4].delimiter[7] );
tran (\labels[4][8] , \labels[4].delimiter_valid[0] );
tran (\labels[4][9] , \labels[4].label[0] );
tran (\labels[4][10] , \labels[4].label[1] );
tran (\labels[4][11] , \labels[4].label[2] );
tran (\labels[4][12] , \labels[4].label[3] );
tran (\labels[4][13] , \labels[4].label[4] );
tran (\labels[4][14] , \labels[4].label[5] );
tran (\labels[4][15] , \labels[4].label[6] );
tran (\labels[4][16] , \labels[4].label[7] );
tran (\labels[4][17] , \labels[4].label[8] );
tran (\labels[4][18] , \labels[4].label[9] );
tran (\labels[4][19] , \labels[4].label[10] );
tran (\labels[4][20] , \labels[4].label[11] );
tran (\labels[4][21] , \labels[4].label[12] );
tran (\labels[4][22] , \labels[4].label[13] );
tran (\labels[4][23] , \labels[4].label[14] );
tran (\labels[4][24] , \labels[4].label[15] );
tran (\labels[4][25] , \labels[4].label[16] );
tran (\labels[4][26] , \labels[4].label[17] );
tran (\labels[4][27] , \labels[4].label[18] );
tran (\labels[4][28] , \labels[4].label[19] );
tran (\labels[4][29] , \labels[4].label[20] );
tran (\labels[4][30] , \labels[4].label[21] );
tran (\labels[4][31] , \labels[4].label[22] );
tran (\labels[4][32] , \labels[4].label[23] );
tran (\labels[4][33] , \labels[4].label[24] );
tran (\labels[4][34] , \labels[4].label[25] );
tran (\labels[4][35] , \labels[4].label[26] );
tran (\labels[4][36] , \labels[4].label[27] );
tran (\labels[4][37] , \labels[4].label[28] );
tran (\labels[4][38] , \labels[4].label[29] );
tran (\labels[4][39] , \labels[4].label[30] );
tran (\labels[4][40] , \labels[4].label[31] );
tran (\labels[4][41] , \labels[4].label[32] );
tran (\labels[4][42] , \labels[4].label[33] );
tran (\labels[4][43] , \labels[4].label[34] );
tran (\labels[4][44] , \labels[4].label[35] );
tran (\labels[4][45] , \labels[4].label[36] );
tran (\labels[4][46] , \labels[4].label[37] );
tran (\labels[4][47] , \labels[4].label[38] );
tran (\labels[4][48] , \labels[4].label[39] );
tran (\labels[4][49] , \labels[4].label[40] );
tran (\labels[4][50] , \labels[4].label[41] );
tran (\labels[4][51] , \labels[4].label[42] );
tran (\labels[4][52] , \labels[4].label[43] );
tran (\labels[4][53] , \labels[4].label[44] );
tran (\labels[4][54] , \labels[4].label[45] );
tran (\labels[4][55] , \labels[4].label[46] );
tran (\labels[4][56] , \labels[4].label[47] );
tran (\labels[4][57] , \labels[4].label[48] );
tran (\labels[4][58] , \labels[4].label[49] );
tran (\labels[4][59] , \labels[4].label[50] );
tran (\labels[4][60] , \labels[4].label[51] );
tran (\labels[4][61] , \labels[4].label[52] );
tran (\labels[4][62] , \labels[4].label[53] );
tran (\labels[4][63] , \labels[4].label[54] );
tran (\labels[4][64] , \labels[4].label[55] );
tran (\labels[4][65] , \labels[4].label[56] );
tran (\labels[4][66] , \labels[4].label[57] );
tran (\labels[4][67] , \labels[4].label[58] );
tran (\labels[4][68] , \labels[4].label[59] );
tran (\labels[4][69] , \labels[4].label[60] );
tran (\labels[4][70] , \labels[4].label[61] );
tran (\labels[4][71] , \labels[4].label[62] );
tran (\labels[4][72] , \labels[4].label[63] );
tran (\labels[4][73] , \labels[4].label[64] );
tran (\labels[4][74] , \labels[4].label[65] );
tran (\labels[4][75] , \labels[4].label[66] );
tran (\labels[4][76] , \labels[4].label[67] );
tran (\labels[4][77] , \labels[4].label[68] );
tran (\labels[4][78] , \labels[4].label[69] );
tran (\labels[4][79] , \labels[4].label[70] );
tran (\labels[4][80] , \labels[4].label[71] );
tran (\labels[4][81] , \labels[4].label[72] );
tran (\labels[4][82] , \labels[4].label[73] );
tran (\labels[4][83] , \labels[4].label[74] );
tran (\labels[4][84] , \labels[4].label[75] );
tran (\labels[4][85] , \labels[4].label[76] );
tran (\labels[4][86] , \labels[4].label[77] );
tran (\labels[4][87] , \labels[4].label[78] );
tran (\labels[4][88] , \labels[4].label[79] );
tran (\labels[4][89] , \labels[4].label[80] );
tran (\labels[4][90] , \labels[4].label[81] );
tran (\labels[4][91] , \labels[4].label[82] );
tran (\labels[4][92] , \labels[4].label[83] );
tran (\labels[4][93] , \labels[4].label[84] );
tran (\labels[4][94] , \labels[4].label[85] );
tran (\labels[4][95] , \labels[4].label[86] );
tran (\labels[4][96] , \labels[4].label[87] );
tran (\labels[4][97] , \labels[4].label[88] );
tran (\labels[4][98] , \labels[4].label[89] );
tran (\labels[4][99] , \labels[4].label[90] );
tran (\labels[4][100] , \labels[4].label[91] );
tran (\labels[4][101] , \labels[4].label[92] );
tran (\labels[4][102] , \labels[4].label[93] );
tran (\labels[4][103] , \labels[4].label[94] );
tran (\labels[4][104] , \labels[4].label[95] );
tran (\labels[4][105] , \labels[4].label[96] );
tran (\labels[4][106] , \labels[4].label[97] );
tran (\labels[4][107] , \labels[4].label[98] );
tran (\labels[4][108] , \labels[4].label[99] );
tran (\labels[4][109] , \labels[4].label[100] );
tran (\labels[4][110] , \labels[4].label[101] );
tran (\labels[4][111] , \labels[4].label[102] );
tran (\labels[4][112] , \labels[4].label[103] );
tran (\labels[4][113] , \labels[4].label[104] );
tran (\labels[4][114] , \labels[4].label[105] );
tran (\labels[4][115] , \labels[4].label[106] );
tran (\labels[4][116] , \labels[4].label[107] );
tran (\labels[4][117] , \labels[4].label[108] );
tran (\labels[4][118] , \labels[4].label[109] );
tran (\labels[4][119] , \labels[4].label[110] );
tran (\labels[4][120] , \labels[4].label[111] );
tran (\labels[4][121] , \labels[4].label[112] );
tran (\labels[4][122] , \labels[4].label[113] );
tran (\labels[4][123] , \labels[4].label[114] );
tran (\labels[4][124] , \labels[4].label[115] );
tran (\labels[4][125] , \labels[4].label[116] );
tran (\labels[4][126] , \labels[4].label[117] );
tran (\labels[4][127] , \labels[4].label[118] );
tran (\labels[4][128] , \labels[4].label[119] );
tran (\labels[4][129] , \labels[4].label[120] );
tran (\labels[4][130] , \labels[4].label[121] );
tran (\labels[4][131] , \labels[4].label[122] );
tran (\labels[4][132] , \labels[4].label[123] );
tran (\labels[4][133] , \labels[4].label[124] );
tran (\labels[4][134] , \labels[4].label[125] );
tran (\labels[4][135] , \labels[4].label[126] );
tran (\labels[4][136] , \labels[4].label[127] );
tran (\labels[4][137] , \labels[4].label[128] );
tran (\labels[4][138] , \labels[4].label[129] );
tran (\labels[4][139] , \labels[4].label[130] );
tran (\labels[4][140] , \labels[4].label[131] );
tran (\labels[4][141] , \labels[4].label[132] );
tran (\labels[4][142] , \labels[4].label[133] );
tran (\labels[4][143] , \labels[4].label[134] );
tran (\labels[4][144] , \labels[4].label[135] );
tran (\labels[4][145] , \labels[4].label[136] );
tran (\labels[4][146] , \labels[4].label[137] );
tran (\labels[4][147] , \labels[4].label[138] );
tran (\labels[4][148] , \labels[4].label[139] );
tran (\labels[4][149] , \labels[4].label[140] );
tran (\labels[4][150] , \labels[4].label[141] );
tran (\labels[4][151] , \labels[4].label[142] );
tran (\labels[4][152] , \labels[4].label[143] );
tran (\labels[4][153] , \labels[4].label[144] );
tran (\labels[4][154] , \labels[4].label[145] );
tran (\labels[4][155] , \labels[4].label[146] );
tran (\labels[4][156] , \labels[4].label[147] );
tran (\labels[4][157] , \labels[4].label[148] );
tran (\labels[4][158] , \labels[4].label[149] );
tran (\labels[4][159] , \labels[4].label[150] );
tran (\labels[4][160] , \labels[4].label[151] );
tran (\labels[4][161] , \labels[4].label[152] );
tran (\labels[4][162] , \labels[4].label[153] );
tran (\labels[4][163] , \labels[4].label[154] );
tran (\labels[4][164] , \labels[4].label[155] );
tran (\labels[4][165] , \labels[4].label[156] );
tran (\labels[4][166] , \labels[4].label[157] );
tran (\labels[4][167] , \labels[4].label[158] );
tran (\labels[4][168] , \labels[4].label[159] );
tran (\labels[4][169] , \labels[4].label[160] );
tran (\labels[4][170] , \labels[4].label[161] );
tran (\labels[4][171] , \labels[4].label[162] );
tran (\labels[4][172] , \labels[4].label[163] );
tran (\labels[4][173] , \labels[4].label[164] );
tran (\labels[4][174] , \labels[4].label[165] );
tran (\labels[4][175] , \labels[4].label[166] );
tran (\labels[4][176] , \labels[4].label[167] );
tran (\labels[4][177] , \labels[4].label[168] );
tran (\labels[4][178] , \labels[4].label[169] );
tran (\labels[4][179] , \labels[4].label[170] );
tran (\labels[4][180] , \labels[4].label[171] );
tran (\labels[4][181] , \labels[4].label[172] );
tran (\labels[4][182] , \labels[4].label[173] );
tran (\labels[4][183] , \labels[4].label[174] );
tran (\labels[4][184] , \labels[4].label[175] );
tran (\labels[4][185] , \labels[4].label[176] );
tran (\labels[4][186] , \labels[4].label[177] );
tran (\labels[4][187] , \labels[4].label[178] );
tran (\labels[4][188] , \labels[4].label[179] );
tran (\labels[4][189] , \labels[4].label[180] );
tran (\labels[4][190] , \labels[4].label[181] );
tran (\labels[4][191] , \labels[4].label[182] );
tran (\labels[4][192] , \labels[4].label[183] );
tran (\labels[4][193] , \labels[4].label[184] );
tran (\labels[4][194] , \labels[4].label[185] );
tran (\labels[4][195] , \labels[4].label[186] );
tran (\labels[4][196] , \labels[4].label[187] );
tran (\labels[4][197] , \labels[4].label[188] );
tran (\labels[4][198] , \labels[4].label[189] );
tran (\labels[4][199] , \labels[4].label[190] );
tran (\labels[4][200] , \labels[4].label[191] );
tran (\labels[4][201] , \labels[4].label[192] );
tran (\labels[4][202] , \labels[4].label[193] );
tran (\labels[4][203] , \labels[4].label[194] );
tran (\labels[4][204] , \labels[4].label[195] );
tran (\labels[4][205] , \labels[4].label[196] );
tran (\labels[4][206] , \labels[4].label[197] );
tran (\labels[4][207] , \labels[4].label[198] );
tran (\labels[4][208] , \labels[4].label[199] );
tran (\labels[4][209] , \labels[4].label[200] );
tran (\labels[4][210] , \labels[4].label[201] );
tran (\labels[4][211] , \labels[4].label[202] );
tran (\labels[4][212] , \labels[4].label[203] );
tran (\labels[4][213] , \labels[4].label[204] );
tran (\labels[4][214] , \labels[4].label[205] );
tran (\labels[4][215] , \labels[4].label[206] );
tran (\labels[4][216] , \labels[4].label[207] );
tran (\labels[4][217] , \labels[4].label[208] );
tran (\labels[4][218] , \labels[4].label[209] );
tran (\labels[4][219] , \labels[4].label[210] );
tran (\labels[4][220] , \labels[4].label[211] );
tran (\labels[4][221] , \labels[4].label[212] );
tran (\labels[4][222] , \labels[4].label[213] );
tran (\labels[4][223] , \labels[4].label[214] );
tran (\labels[4][224] , \labels[4].label[215] );
tran (\labels[4][225] , \labels[4].label[216] );
tran (\labels[4][226] , \labels[4].label[217] );
tran (\labels[4][227] , \labels[4].label[218] );
tran (\labels[4][228] , \labels[4].label[219] );
tran (\labels[4][229] , \labels[4].label[220] );
tran (\labels[4][230] , \labels[4].label[221] );
tran (\labels[4][231] , \labels[4].label[222] );
tran (\labels[4][232] , \labels[4].label[223] );
tran (\labels[4][233] , \labels[4].label[224] );
tran (\labels[4][234] , \labels[4].label[225] );
tran (\labels[4][235] , \labels[4].label[226] );
tran (\labels[4][236] , \labels[4].label[227] );
tran (\labels[4][237] , \labels[4].label[228] );
tran (\labels[4][238] , \labels[4].label[229] );
tran (\labels[4][239] , \labels[4].label[230] );
tran (\labels[4][240] , \labels[4].label[231] );
tran (\labels[4][241] , \labels[4].label[232] );
tran (\labels[4][242] , \labels[4].label[233] );
tran (\labels[4][243] , \labels[4].label[234] );
tran (\labels[4][244] , \labels[4].label[235] );
tran (\labels[4][245] , \labels[4].label[236] );
tran (\labels[4][246] , \labels[4].label[237] );
tran (\labels[4][247] , \labels[4].label[238] );
tran (\labels[4][248] , \labels[4].label[239] );
tran (\labels[4][249] , \labels[4].label[240] );
tran (\labels[4][250] , \labels[4].label[241] );
tran (\labels[4][251] , \labels[4].label[242] );
tran (\labels[4][252] , \labels[4].label[243] );
tran (\labels[4][253] , \labels[4].label[244] );
tran (\labels[4][254] , \labels[4].label[245] );
tran (\labels[4][255] , \labels[4].label[246] );
tran (\labels[4][256] , \labels[4].label[247] );
tran (\labels[4][257] , \labels[4].label[248] );
tran (\labels[4][258] , \labels[4].label[249] );
tran (\labels[4][259] , \labels[4].label[250] );
tran (\labels[4][260] , \labels[4].label[251] );
tran (\labels[4][261] , \labels[4].label[252] );
tran (\labels[4][262] , \labels[4].label[253] );
tran (\labels[4][263] , \labels[4].label[254] );
tran (\labels[4][264] , \labels[4].label[255] );
tran (\labels[4][265] , \labels[4].label_size[0] );
tran (\labels[4][266] , \labels[4].label_size[1] );
tran (\labels[4][267] , \labels[4].label_size[2] );
tran (\labels[4][268] , \labels[4].label_size[3] );
tran (\labels[4][269] , \labels[4].label_size[4] );
tran (\labels[4][270] , \labels[4].label_size[5] );
tran (\labels[4][271] , \labels[4].guid_size[0] );
tran (\labels[5][0] , \labels[5].delimiter[0] );
tran (\labels[5][1] , \labels[5].delimiter[1] );
tran (\labels[5][2] , \labels[5].delimiter[2] );
tran (\labels[5][3] , \labels[5].delimiter[3] );
tran (\labels[5][4] , \labels[5].delimiter[4] );
tran (\labels[5][5] , \labels[5].delimiter[5] );
tran (\labels[5][6] , \labels[5].delimiter[6] );
tran (\labels[5][7] , \labels[5].delimiter[7] );
tran (\labels[5][8] , \labels[5].delimiter_valid[0] );
tran (\labels[5][9] , \labels[5].label[0] );
tran (\labels[5][10] , \labels[5].label[1] );
tran (\labels[5][11] , \labels[5].label[2] );
tran (\labels[5][12] , \labels[5].label[3] );
tran (\labels[5][13] , \labels[5].label[4] );
tran (\labels[5][14] , \labels[5].label[5] );
tran (\labels[5][15] , \labels[5].label[6] );
tran (\labels[5][16] , \labels[5].label[7] );
tran (\labels[5][17] , \labels[5].label[8] );
tran (\labels[5][18] , \labels[5].label[9] );
tran (\labels[5][19] , \labels[5].label[10] );
tran (\labels[5][20] , \labels[5].label[11] );
tran (\labels[5][21] , \labels[5].label[12] );
tran (\labels[5][22] , \labels[5].label[13] );
tran (\labels[5][23] , \labels[5].label[14] );
tran (\labels[5][24] , \labels[5].label[15] );
tran (\labels[5][25] , \labels[5].label[16] );
tran (\labels[5][26] , \labels[5].label[17] );
tran (\labels[5][27] , \labels[5].label[18] );
tran (\labels[5][28] , \labels[5].label[19] );
tran (\labels[5][29] , \labels[5].label[20] );
tran (\labels[5][30] , \labels[5].label[21] );
tran (\labels[5][31] , \labels[5].label[22] );
tran (\labels[5][32] , \labels[5].label[23] );
tran (\labels[5][33] , \labels[5].label[24] );
tran (\labels[5][34] , \labels[5].label[25] );
tran (\labels[5][35] , \labels[5].label[26] );
tran (\labels[5][36] , \labels[5].label[27] );
tran (\labels[5][37] , \labels[5].label[28] );
tran (\labels[5][38] , \labels[5].label[29] );
tran (\labels[5][39] , \labels[5].label[30] );
tran (\labels[5][40] , \labels[5].label[31] );
tran (\labels[5][41] , \labels[5].label[32] );
tran (\labels[5][42] , \labels[5].label[33] );
tran (\labels[5][43] , \labels[5].label[34] );
tran (\labels[5][44] , \labels[5].label[35] );
tran (\labels[5][45] , \labels[5].label[36] );
tran (\labels[5][46] , \labels[5].label[37] );
tran (\labels[5][47] , \labels[5].label[38] );
tran (\labels[5][48] , \labels[5].label[39] );
tran (\labels[5][49] , \labels[5].label[40] );
tran (\labels[5][50] , \labels[5].label[41] );
tran (\labels[5][51] , \labels[5].label[42] );
tran (\labels[5][52] , \labels[5].label[43] );
tran (\labels[5][53] , \labels[5].label[44] );
tran (\labels[5][54] , \labels[5].label[45] );
tran (\labels[5][55] , \labels[5].label[46] );
tran (\labels[5][56] , \labels[5].label[47] );
tran (\labels[5][57] , \labels[5].label[48] );
tran (\labels[5][58] , \labels[5].label[49] );
tran (\labels[5][59] , \labels[5].label[50] );
tran (\labels[5][60] , \labels[5].label[51] );
tran (\labels[5][61] , \labels[5].label[52] );
tran (\labels[5][62] , \labels[5].label[53] );
tran (\labels[5][63] , \labels[5].label[54] );
tran (\labels[5][64] , \labels[5].label[55] );
tran (\labels[5][65] , \labels[5].label[56] );
tran (\labels[5][66] , \labels[5].label[57] );
tran (\labels[5][67] , \labels[5].label[58] );
tran (\labels[5][68] , \labels[5].label[59] );
tran (\labels[5][69] , \labels[5].label[60] );
tran (\labels[5][70] , \labels[5].label[61] );
tran (\labels[5][71] , \labels[5].label[62] );
tran (\labels[5][72] , \labels[5].label[63] );
tran (\labels[5][73] , \labels[5].label[64] );
tran (\labels[5][74] , \labels[5].label[65] );
tran (\labels[5][75] , \labels[5].label[66] );
tran (\labels[5][76] , \labels[5].label[67] );
tran (\labels[5][77] , \labels[5].label[68] );
tran (\labels[5][78] , \labels[5].label[69] );
tran (\labels[5][79] , \labels[5].label[70] );
tran (\labels[5][80] , \labels[5].label[71] );
tran (\labels[5][81] , \labels[5].label[72] );
tran (\labels[5][82] , \labels[5].label[73] );
tran (\labels[5][83] , \labels[5].label[74] );
tran (\labels[5][84] , \labels[5].label[75] );
tran (\labels[5][85] , \labels[5].label[76] );
tran (\labels[5][86] , \labels[5].label[77] );
tran (\labels[5][87] , \labels[5].label[78] );
tran (\labels[5][88] , \labels[5].label[79] );
tran (\labels[5][89] , \labels[5].label[80] );
tran (\labels[5][90] , \labels[5].label[81] );
tran (\labels[5][91] , \labels[5].label[82] );
tran (\labels[5][92] , \labels[5].label[83] );
tran (\labels[5][93] , \labels[5].label[84] );
tran (\labels[5][94] , \labels[5].label[85] );
tran (\labels[5][95] , \labels[5].label[86] );
tran (\labels[5][96] , \labels[5].label[87] );
tran (\labels[5][97] , \labels[5].label[88] );
tran (\labels[5][98] , \labels[5].label[89] );
tran (\labels[5][99] , \labels[5].label[90] );
tran (\labels[5][100] , \labels[5].label[91] );
tran (\labels[5][101] , \labels[5].label[92] );
tran (\labels[5][102] , \labels[5].label[93] );
tran (\labels[5][103] , \labels[5].label[94] );
tran (\labels[5][104] , \labels[5].label[95] );
tran (\labels[5][105] , \labels[5].label[96] );
tran (\labels[5][106] , \labels[5].label[97] );
tran (\labels[5][107] , \labels[5].label[98] );
tran (\labels[5][108] , \labels[5].label[99] );
tran (\labels[5][109] , \labels[5].label[100] );
tran (\labels[5][110] , \labels[5].label[101] );
tran (\labels[5][111] , \labels[5].label[102] );
tran (\labels[5][112] , \labels[5].label[103] );
tran (\labels[5][113] , \labels[5].label[104] );
tran (\labels[5][114] , \labels[5].label[105] );
tran (\labels[5][115] , \labels[5].label[106] );
tran (\labels[5][116] , \labels[5].label[107] );
tran (\labels[5][117] , \labels[5].label[108] );
tran (\labels[5][118] , \labels[5].label[109] );
tran (\labels[5][119] , \labels[5].label[110] );
tran (\labels[5][120] , \labels[5].label[111] );
tran (\labels[5][121] , \labels[5].label[112] );
tran (\labels[5][122] , \labels[5].label[113] );
tran (\labels[5][123] , \labels[5].label[114] );
tran (\labels[5][124] , \labels[5].label[115] );
tran (\labels[5][125] , \labels[5].label[116] );
tran (\labels[5][126] , \labels[5].label[117] );
tran (\labels[5][127] , \labels[5].label[118] );
tran (\labels[5][128] , \labels[5].label[119] );
tran (\labels[5][129] , \labels[5].label[120] );
tran (\labels[5][130] , \labels[5].label[121] );
tran (\labels[5][131] , \labels[5].label[122] );
tran (\labels[5][132] , \labels[5].label[123] );
tran (\labels[5][133] , \labels[5].label[124] );
tran (\labels[5][134] , \labels[5].label[125] );
tran (\labels[5][135] , \labels[5].label[126] );
tran (\labels[5][136] , \labels[5].label[127] );
tran (\labels[5][137] , \labels[5].label[128] );
tran (\labels[5][138] , \labels[5].label[129] );
tran (\labels[5][139] , \labels[5].label[130] );
tran (\labels[5][140] , \labels[5].label[131] );
tran (\labels[5][141] , \labels[5].label[132] );
tran (\labels[5][142] , \labels[5].label[133] );
tran (\labels[5][143] , \labels[5].label[134] );
tran (\labels[5][144] , \labels[5].label[135] );
tran (\labels[5][145] , \labels[5].label[136] );
tran (\labels[5][146] , \labels[5].label[137] );
tran (\labels[5][147] , \labels[5].label[138] );
tran (\labels[5][148] , \labels[5].label[139] );
tran (\labels[5][149] , \labels[5].label[140] );
tran (\labels[5][150] , \labels[5].label[141] );
tran (\labels[5][151] , \labels[5].label[142] );
tran (\labels[5][152] , \labels[5].label[143] );
tran (\labels[5][153] , \labels[5].label[144] );
tran (\labels[5][154] , \labels[5].label[145] );
tran (\labels[5][155] , \labels[5].label[146] );
tran (\labels[5][156] , \labels[5].label[147] );
tran (\labels[5][157] , \labels[5].label[148] );
tran (\labels[5][158] , \labels[5].label[149] );
tran (\labels[5][159] , \labels[5].label[150] );
tran (\labels[5][160] , \labels[5].label[151] );
tran (\labels[5][161] , \labels[5].label[152] );
tran (\labels[5][162] , \labels[5].label[153] );
tran (\labels[5][163] , \labels[5].label[154] );
tran (\labels[5][164] , \labels[5].label[155] );
tran (\labels[5][165] , \labels[5].label[156] );
tran (\labels[5][166] , \labels[5].label[157] );
tran (\labels[5][167] , \labels[5].label[158] );
tran (\labels[5][168] , \labels[5].label[159] );
tran (\labels[5][169] , \labels[5].label[160] );
tran (\labels[5][170] , \labels[5].label[161] );
tran (\labels[5][171] , \labels[5].label[162] );
tran (\labels[5][172] , \labels[5].label[163] );
tran (\labels[5][173] , \labels[5].label[164] );
tran (\labels[5][174] , \labels[5].label[165] );
tran (\labels[5][175] , \labels[5].label[166] );
tran (\labels[5][176] , \labels[5].label[167] );
tran (\labels[5][177] , \labels[5].label[168] );
tran (\labels[5][178] , \labels[5].label[169] );
tran (\labels[5][179] , \labels[5].label[170] );
tran (\labels[5][180] , \labels[5].label[171] );
tran (\labels[5][181] , \labels[5].label[172] );
tran (\labels[5][182] , \labels[5].label[173] );
tran (\labels[5][183] , \labels[5].label[174] );
tran (\labels[5][184] , \labels[5].label[175] );
tran (\labels[5][185] , \labels[5].label[176] );
tran (\labels[5][186] , \labels[5].label[177] );
tran (\labels[5][187] , \labels[5].label[178] );
tran (\labels[5][188] , \labels[5].label[179] );
tran (\labels[5][189] , \labels[5].label[180] );
tran (\labels[5][190] , \labels[5].label[181] );
tran (\labels[5][191] , \labels[5].label[182] );
tran (\labels[5][192] , \labels[5].label[183] );
tran (\labels[5][193] , \labels[5].label[184] );
tran (\labels[5][194] , \labels[5].label[185] );
tran (\labels[5][195] , \labels[5].label[186] );
tran (\labels[5][196] , \labels[5].label[187] );
tran (\labels[5][197] , \labels[5].label[188] );
tran (\labels[5][198] , \labels[5].label[189] );
tran (\labels[5][199] , \labels[5].label[190] );
tran (\labels[5][200] , \labels[5].label[191] );
tran (\labels[5][201] , \labels[5].label[192] );
tran (\labels[5][202] , \labels[5].label[193] );
tran (\labels[5][203] , \labels[5].label[194] );
tran (\labels[5][204] , \labels[5].label[195] );
tran (\labels[5][205] , \labels[5].label[196] );
tran (\labels[5][206] , \labels[5].label[197] );
tran (\labels[5][207] , \labels[5].label[198] );
tran (\labels[5][208] , \labels[5].label[199] );
tran (\labels[5][209] , \labels[5].label[200] );
tran (\labels[5][210] , \labels[5].label[201] );
tran (\labels[5][211] , \labels[5].label[202] );
tran (\labels[5][212] , \labels[5].label[203] );
tran (\labels[5][213] , \labels[5].label[204] );
tran (\labels[5][214] , \labels[5].label[205] );
tran (\labels[5][215] , \labels[5].label[206] );
tran (\labels[5][216] , \labels[5].label[207] );
tran (\labels[5][217] , \labels[5].label[208] );
tran (\labels[5][218] , \labels[5].label[209] );
tran (\labels[5][219] , \labels[5].label[210] );
tran (\labels[5][220] , \labels[5].label[211] );
tran (\labels[5][221] , \labels[5].label[212] );
tran (\labels[5][222] , \labels[5].label[213] );
tran (\labels[5][223] , \labels[5].label[214] );
tran (\labels[5][224] , \labels[5].label[215] );
tran (\labels[5][225] , \labels[5].label[216] );
tran (\labels[5][226] , \labels[5].label[217] );
tran (\labels[5][227] , \labels[5].label[218] );
tran (\labels[5][228] , \labels[5].label[219] );
tran (\labels[5][229] , \labels[5].label[220] );
tran (\labels[5][230] , \labels[5].label[221] );
tran (\labels[5][231] , \labels[5].label[222] );
tran (\labels[5][232] , \labels[5].label[223] );
tran (\labels[5][233] , \labels[5].label[224] );
tran (\labels[5][234] , \labels[5].label[225] );
tran (\labels[5][235] , \labels[5].label[226] );
tran (\labels[5][236] , \labels[5].label[227] );
tran (\labels[5][237] , \labels[5].label[228] );
tran (\labels[5][238] , \labels[5].label[229] );
tran (\labels[5][239] , \labels[5].label[230] );
tran (\labels[5][240] , \labels[5].label[231] );
tran (\labels[5][241] , \labels[5].label[232] );
tran (\labels[5][242] , \labels[5].label[233] );
tran (\labels[5][243] , \labels[5].label[234] );
tran (\labels[5][244] , \labels[5].label[235] );
tran (\labels[5][245] , \labels[5].label[236] );
tran (\labels[5][246] , \labels[5].label[237] );
tran (\labels[5][247] , \labels[5].label[238] );
tran (\labels[5][248] , \labels[5].label[239] );
tran (\labels[5][249] , \labels[5].label[240] );
tran (\labels[5][250] , \labels[5].label[241] );
tran (\labels[5][251] , \labels[5].label[242] );
tran (\labels[5][252] , \labels[5].label[243] );
tran (\labels[5][253] , \labels[5].label[244] );
tran (\labels[5][254] , \labels[5].label[245] );
tran (\labels[5][255] , \labels[5].label[246] );
tran (\labels[5][256] , \labels[5].label[247] );
tran (\labels[5][257] , \labels[5].label[248] );
tran (\labels[5][258] , \labels[5].label[249] );
tran (\labels[5][259] , \labels[5].label[250] );
tran (\labels[5][260] , \labels[5].label[251] );
tran (\labels[5][261] , \labels[5].label[252] );
tran (\labels[5][262] , \labels[5].label[253] );
tran (\labels[5][263] , \labels[5].label[254] );
tran (\labels[5][264] , \labels[5].label[255] );
tran (\labels[5][265] , \labels[5].label_size[0] );
tran (\labels[5][266] , \labels[5].label_size[1] );
tran (\labels[5][267] , \labels[5].label_size[2] );
tran (\labels[5][268] , \labels[5].label_size[3] );
tran (\labels[5][269] , \labels[5].label_size[4] );
tran (\labels[5][270] , \labels[5].label_size[5] );
tran (\labels[5][271] , \labels[5].guid_size[0] );
tran (\labels[6][0] , \labels[6].delimiter[0] );
tran (\labels[6][1] , \labels[6].delimiter[1] );
tran (\labels[6][2] , \labels[6].delimiter[2] );
tran (\labels[6][3] , \labels[6].delimiter[3] );
tran (\labels[6][4] , \labels[6].delimiter[4] );
tran (\labels[6][5] , \labels[6].delimiter[5] );
tran (\labels[6][6] , \labels[6].delimiter[6] );
tran (\labels[6][7] , \labels[6].delimiter[7] );
tran (\labels[6][8] , \labels[6].delimiter_valid[0] );
tran (\labels[6][9] , \labels[6].label[0] );
tran (\labels[6][10] , \labels[6].label[1] );
tran (\labels[6][11] , \labels[6].label[2] );
tran (\labels[6][12] , \labels[6].label[3] );
tran (\labels[6][13] , \labels[6].label[4] );
tran (\labels[6][14] , \labels[6].label[5] );
tran (\labels[6][15] , \labels[6].label[6] );
tran (\labels[6][16] , \labels[6].label[7] );
tran (\labels[6][17] , \labels[6].label[8] );
tran (\labels[6][18] , \labels[6].label[9] );
tran (\labels[6][19] , \labels[6].label[10] );
tran (\labels[6][20] , \labels[6].label[11] );
tran (\labels[6][21] , \labels[6].label[12] );
tran (\labels[6][22] , \labels[6].label[13] );
tran (\labels[6][23] , \labels[6].label[14] );
tran (\labels[6][24] , \labels[6].label[15] );
tran (\labels[6][25] , \labels[6].label[16] );
tran (\labels[6][26] , \labels[6].label[17] );
tran (\labels[6][27] , \labels[6].label[18] );
tran (\labels[6][28] , \labels[6].label[19] );
tran (\labels[6][29] , \labels[6].label[20] );
tran (\labels[6][30] , \labels[6].label[21] );
tran (\labels[6][31] , \labels[6].label[22] );
tran (\labels[6][32] , \labels[6].label[23] );
tran (\labels[6][33] , \labels[6].label[24] );
tran (\labels[6][34] , \labels[6].label[25] );
tran (\labels[6][35] , \labels[6].label[26] );
tran (\labels[6][36] , \labels[6].label[27] );
tran (\labels[6][37] , \labels[6].label[28] );
tran (\labels[6][38] , \labels[6].label[29] );
tran (\labels[6][39] , \labels[6].label[30] );
tran (\labels[6][40] , \labels[6].label[31] );
tran (\labels[6][41] , \labels[6].label[32] );
tran (\labels[6][42] , \labels[6].label[33] );
tran (\labels[6][43] , \labels[6].label[34] );
tran (\labels[6][44] , \labels[6].label[35] );
tran (\labels[6][45] , \labels[6].label[36] );
tran (\labels[6][46] , \labels[6].label[37] );
tran (\labels[6][47] , \labels[6].label[38] );
tran (\labels[6][48] , \labels[6].label[39] );
tran (\labels[6][49] , \labels[6].label[40] );
tran (\labels[6][50] , \labels[6].label[41] );
tran (\labels[6][51] , \labels[6].label[42] );
tran (\labels[6][52] , \labels[6].label[43] );
tran (\labels[6][53] , \labels[6].label[44] );
tran (\labels[6][54] , \labels[6].label[45] );
tran (\labels[6][55] , \labels[6].label[46] );
tran (\labels[6][56] , \labels[6].label[47] );
tran (\labels[6][57] , \labels[6].label[48] );
tran (\labels[6][58] , \labels[6].label[49] );
tran (\labels[6][59] , \labels[6].label[50] );
tran (\labels[6][60] , \labels[6].label[51] );
tran (\labels[6][61] , \labels[6].label[52] );
tran (\labels[6][62] , \labels[6].label[53] );
tran (\labels[6][63] , \labels[6].label[54] );
tran (\labels[6][64] , \labels[6].label[55] );
tran (\labels[6][65] , \labels[6].label[56] );
tran (\labels[6][66] , \labels[6].label[57] );
tran (\labels[6][67] , \labels[6].label[58] );
tran (\labels[6][68] , \labels[6].label[59] );
tran (\labels[6][69] , \labels[6].label[60] );
tran (\labels[6][70] , \labels[6].label[61] );
tran (\labels[6][71] , \labels[6].label[62] );
tran (\labels[6][72] , \labels[6].label[63] );
tran (\labels[6][73] , \labels[6].label[64] );
tran (\labels[6][74] , \labels[6].label[65] );
tran (\labels[6][75] , \labels[6].label[66] );
tran (\labels[6][76] , \labels[6].label[67] );
tran (\labels[6][77] , \labels[6].label[68] );
tran (\labels[6][78] , \labels[6].label[69] );
tran (\labels[6][79] , \labels[6].label[70] );
tran (\labels[6][80] , \labels[6].label[71] );
tran (\labels[6][81] , \labels[6].label[72] );
tran (\labels[6][82] , \labels[6].label[73] );
tran (\labels[6][83] , \labels[6].label[74] );
tran (\labels[6][84] , \labels[6].label[75] );
tran (\labels[6][85] , \labels[6].label[76] );
tran (\labels[6][86] , \labels[6].label[77] );
tran (\labels[6][87] , \labels[6].label[78] );
tran (\labels[6][88] , \labels[6].label[79] );
tran (\labels[6][89] , \labels[6].label[80] );
tran (\labels[6][90] , \labels[6].label[81] );
tran (\labels[6][91] , \labels[6].label[82] );
tran (\labels[6][92] , \labels[6].label[83] );
tran (\labels[6][93] , \labels[6].label[84] );
tran (\labels[6][94] , \labels[6].label[85] );
tran (\labels[6][95] , \labels[6].label[86] );
tran (\labels[6][96] , \labels[6].label[87] );
tran (\labels[6][97] , \labels[6].label[88] );
tran (\labels[6][98] , \labels[6].label[89] );
tran (\labels[6][99] , \labels[6].label[90] );
tran (\labels[6][100] , \labels[6].label[91] );
tran (\labels[6][101] , \labels[6].label[92] );
tran (\labels[6][102] , \labels[6].label[93] );
tran (\labels[6][103] , \labels[6].label[94] );
tran (\labels[6][104] , \labels[6].label[95] );
tran (\labels[6][105] , \labels[6].label[96] );
tran (\labels[6][106] , \labels[6].label[97] );
tran (\labels[6][107] , \labels[6].label[98] );
tran (\labels[6][108] , \labels[6].label[99] );
tran (\labels[6][109] , \labels[6].label[100] );
tran (\labels[6][110] , \labels[6].label[101] );
tran (\labels[6][111] , \labels[6].label[102] );
tran (\labels[6][112] , \labels[6].label[103] );
tran (\labels[6][113] , \labels[6].label[104] );
tran (\labels[6][114] , \labels[6].label[105] );
tran (\labels[6][115] , \labels[6].label[106] );
tran (\labels[6][116] , \labels[6].label[107] );
tran (\labels[6][117] , \labels[6].label[108] );
tran (\labels[6][118] , \labels[6].label[109] );
tran (\labels[6][119] , \labels[6].label[110] );
tran (\labels[6][120] , \labels[6].label[111] );
tran (\labels[6][121] , \labels[6].label[112] );
tran (\labels[6][122] , \labels[6].label[113] );
tran (\labels[6][123] , \labels[6].label[114] );
tran (\labels[6][124] , \labels[6].label[115] );
tran (\labels[6][125] , \labels[6].label[116] );
tran (\labels[6][126] , \labels[6].label[117] );
tran (\labels[6][127] , \labels[6].label[118] );
tran (\labels[6][128] , \labels[6].label[119] );
tran (\labels[6][129] , \labels[6].label[120] );
tran (\labels[6][130] , \labels[6].label[121] );
tran (\labels[6][131] , \labels[6].label[122] );
tran (\labels[6][132] , \labels[6].label[123] );
tran (\labels[6][133] , \labels[6].label[124] );
tran (\labels[6][134] , \labels[6].label[125] );
tran (\labels[6][135] , \labels[6].label[126] );
tran (\labels[6][136] , \labels[6].label[127] );
tran (\labels[6][137] , \labels[6].label[128] );
tran (\labels[6][138] , \labels[6].label[129] );
tran (\labels[6][139] , \labels[6].label[130] );
tran (\labels[6][140] , \labels[6].label[131] );
tran (\labels[6][141] , \labels[6].label[132] );
tran (\labels[6][142] , \labels[6].label[133] );
tran (\labels[6][143] , \labels[6].label[134] );
tran (\labels[6][144] , \labels[6].label[135] );
tran (\labels[6][145] , \labels[6].label[136] );
tran (\labels[6][146] , \labels[6].label[137] );
tran (\labels[6][147] , \labels[6].label[138] );
tran (\labels[6][148] , \labels[6].label[139] );
tran (\labels[6][149] , \labels[6].label[140] );
tran (\labels[6][150] , \labels[6].label[141] );
tran (\labels[6][151] , \labels[6].label[142] );
tran (\labels[6][152] , \labels[6].label[143] );
tran (\labels[6][153] , \labels[6].label[144] );
tran (\labels[6][154] , \labels[6].label[145] );
tran (\labels[6][155] , \labels[6].label[146] );
tran (\labels[6][156] , \labels[6].label[147] );
tran (\labels[6][157] , \labels[6].label[148] );
tran (\labels[6][158] , \labels[6].label[149] );
tran (\labels[6][159] , \labels[6].label[150] );
tran (\labels[6][160] , \labels[6].label[151] );
tran (\labels[6][161] , \labels[6].label[152] );
tran (\labels[6][162] , \labels[6].label[153] );
tran (\labels[6][163] , \labels[6].label[154] );
tran (\labels[6][164] , \labels[6].label[155] );
tran (\labels[6][165] , \labels[6].label[156] );
tran (\labels[6][166] , \labels[6].label[157] );
tran (\labels[6][167] , \labels[6].label[158] );
tran (\labels[6][168] , \labels[6].label[159] );
tran (\labels[6][169] , \labels[6].label[160] );
tran (\labels[6][170] , \labels[6].label[161] );
tran (\labels[6][171] , \labels[6].label[162] );
tran (\labels[6][172] , \labels[6].label[163] );
tran (\labels[6][173] , \labels[6].label[164] );
tran (\labels[6][174] , \labels[6].label[165] );
tran (\labels[6][175] , \labels[6].label[166] );
tran (\labels[6][176] , \labels[6].label[167] );
tran (\labels[6][177] , \labels[6].label[168] );
tran (\labels[6][178] , \labels[6].label[169] );
tran (\labels[6][179] , \labels[6].label[170] );
tran (\labels[6][180] , \labels[6].label[171] );
tran (\labels[6][181] , \labels[6].label[172] );
tran (\labels[6][182] , \labels[6].label[173] );
tran (\labels[6][183] , \labels[6].label[174] );
tran (\labels[6][184] , \labels[6].label[175] );
tran (\labels[6][185] , \labels[6].label[176] );
tran (\labels[6][186] , \labels[6].label[177] );
tran (\labels[6][187] , \labels[6].label[178] );
tran (\labels[6][188] , \labels[6].label[179] );
tran (\labels[6][189] , \labels[6].label[180] );
tran (\labels[6][190] , \labels[6].label[181] );
tran (\labels[6][191] , \labels[6].label[182] );
tran (\labels[6][192] , \labels[6].label[183] );
tran (\labels[6][193] , \labels[6].label[184] );
tran (\labels[6][194] , \labels[6].label[185] );
tran (\labels[6][195] , \labels[6].label[186] );
tran (\labels[6][196] , \labels[6].label[187] );
tran (\labels[6][197] , \labels[6].label[188] );
tran (\labels[6][198] , \labels[6].label[189] );
tran (\labels[6][199] , \labels[6].label[190] );
tran (\labels[6][200] , \labels[6].label[191] );
tran (\labels[6][201] , \labels[6].label[192] );
tran (\labels[6][202] , \labels[6].label[193] );
tran (\labels[6][203] , \labels[6].label[194] );
tran (\labels[6][204] , \labels[6].label[195] );
tran (\labels[6][205] , \labels[6].label[196] );
tran (\labels[6][206] , \labels[6].label[197] );
tran (\labels[6][207] , \labels[6].label[198] );
tran (\labels[6][208] , \labels[6].label[199] );
tran (\labels[6][209] , \labels[6].label[200] );
tran (\labels[6][210] , \labels[6].label[201] );
tran (\labels[6][211] , \labels[6].label[202] );
tran (\labels[6][212] , \labels[6].label[203] );
tran (\labels[6][213] , \labels[6].label[204] );
tran (\labels[6][214] , \labels[6].label[205] );
tran (\labels[6][215] , \labels[6].label[206] );
tran (\labels[6][216] , \labels[6].label[207] );
tran (\labels[6][217] , \labels[6].label[208] );
tran (\labels[6][218] , \labels[6].label[209] );
tran (\labels[6][219] , \labels[6].label[210] );
tran (\labels[6][220] , \labels[6].label[211] );
tran (\labels[6][221] , \labels[6].label[212] );
tran (\labels[6][222] , \labels[6].label[213] );
tran (\labels[6][223] , \labels[6].label[214] );
tran (\labels[6][224] , \labels[6].label[215] );
tran (\labels[6][225] , \labels[6].label[216] );
tran (\labels[6][226] , \labels[6].label[217] );
tran (\labels[6][227] , \labels[6].label[218] );
tran (\labels[6][228] , \labels[6].label[219] );
tran (\labels[6][229] , \labels[6].label[220] );
tran (\labels[6][230] , \labels[6].label[221] );
tran (\labels[6][231] , \labels[6].label[222] );
tran (\labels[6][232] , \labels[6].label[223] );
tran (\labels[6][233] , \labels[6].label[224] );
tran (\labels[6][234] , \labels[6].label[225] );
tran (\labels[6][235] , \labels[6].label[226] );
tran (\labels[6][236] , \labels[6].label[227] );
tran (\labels[6][237] , \labels[6].label[228] );
tran (\labels[6][238] , \labels[6].label[229] );
tran (\labels[6][239] , \labels[6].label[230] );
tran (\labels[6][240] , \labels[6].label[231] );
tran (\labels[6][241] , \labels[6].label[232] );
tran (\labels[6][242] , \labels[6].label[233] );
tran (\labels[6][243] , \labels[6].label[234] );
tran (\labels[6][244] , \labels[6].label[235] );
tran (\labels[6][245] , \labels[6].label[236] );
tran (\labels[6][246] , \labels[6].label[237] );
tran (\labels[6][247] , \labels[6].label[238] );
tran (\labels[6][248] , \labels[6].label[239] );
tran (\labels[6][249] , \labels[6].label[240] );
tran (\labels[6][250] , \labels[6].label[241] );
tran (\labels[6][251] , \labels[6].label[242] );
tran (\labels[6][252] , \labels[6].label[243] );
tran (\labels[6][253] , \labels[6].label[244] );
tran (\labels[6][254] , \labels[6].label[245] );
tran (\labels[6][255] , \labels[6].label[246] );
tran (\labels[6][256] , \labels[6].label[247] );
tran (\labels[6][257] , \labels[6].label[248] );
tran (\labels[6][258] , \labels[6].label[249] );
tran (\labels[6][259] , \labels[6].label[250] );
tran (\labels[6][260] , \labels[6].label[251] );
tran (\labels[6][261] , \labels[6].label[252] );
tran (\labels[6][262] , \labels[6].label[253] );
tran (\labels[6][263] , \labels[6].label[254] );
tran (\labels[6][264] , \labels[6].label[255] );
tran (\labels[6][265] , \labels[6].label_size[0] );
tran (\labels[6][266] , \labels[6].label_size[1] );
tran (\labels[6][267] , \labels[6].label_size[2] );
tran (\labels[6][268] , \labels[6].label_size[3] );
tran (\labels[6][269] , \labels[6].label_size[4] );
tran (\labels[6][270] , \labels[6].label_size[5] );
tran (\labels[6][271] , \labels[6].guid_size[0] );
tran (\labels[7][0] , \labels[7].delimiter[0] );
tran (\labels[7][1] , \labels[7].delimiter[1] );
tran (\labels[7][2] , \labels[7].delimiter[2] );
tran (\labels[7][3] , \labels[7].delimiter[3] );
tran (\labels[7][4] , \labels[7].delimiter[4] );
tran (\labels[7][5] , \labels[7].delimiter[5] );
tran (\labels[7][6] , \labels[7].delimiter[6] );
tran (\labels[7][7] , \labels[7].delimiter[7] );
tran (\labels[7][8] , \labels[7].delimiter_valid[0] );
tran (\labels[7][9] , \labels[7].label[0] );
tran (\labels[7][10] , \labels[7].label[1] );
tran (\labels[7][11] , \labels[7].label[2] );
tran (\labels[7][12] , \labels[7].label[3] );
tran (\labels[7][13] , \labels[7].label[4] );
tran (\labels[7][14] , \labels[7].label[5] );
tran (\labels[7][15] , \labels[7].label[6] );
tran (\labels[7][16] , \labels[7].label[7] );
tran (\labels[7][17] , \labels[7].label[8] );
tran (\labels[7][18] , \labels[7].label[9] );
tran (\labels[7][19] , \labels[7].label[10] );
tran (\labels[7][20] , \labels[7].label[11] );
tran (\labels[7][21] , \labels[7].label[12] );
tran (\labels[7][22] , \labels[7].label[13] );
tran (\labels[7][23] , \labels[7].label[14] );
tran (\labels[7][24] , \labels[7].label[15] );
tran (\labels[7][25] , \labels[7].label[16] );
tran (\labels[7][26] , \labels[7].label[17] );
tran (\labels[7][27] , \labels[7].label[18] );
tran (\labels[7][28] , \labels[7].label[19] );
tran (\labels[7][29] , \labels[7].label[20] );
tran (\labels[7][30] , \labels[7].label[21] );
tran (\labels[7][31] , \labels[7].label[22] );
tran (\labels[7][32] , \labels[7].label[23] );
tran (\labels[7][33] , \labels[7].label[24] );
tran (\labels[7][34] , \labels[7].label[25] );
tran (\labels[7][35] , \labels[7].label[26] );
tran (\labels[7][36] , \labels[7].label[27] );
tran (\labels[7][37] , \labels[7].label[28] );
tran (\labels[7][38] , \labels[7].label[29] );
tran (\labels[7][39] , \labels[7].label[30] );
tran (\labels[7][40] , \labels[7].label[31] );
tran (\labels[7][41] , \labels[7].label[32] );
tran (\labels[7][42] , \labels[7].label[33] );
tran (\labels[7][43] , \labels[7].label[34] );
tran (\labels[7][44] , \labels[7].label[35] );
tran (\labels[7][45] , \labels[7].label[36] );
tran (\labels[7][46] , \labels[7].label[37] );
tran (\labels[7][47] , \labels[7].label[38] );
tran (\labels[7][48] , \labels[7].label[39] );
tran (\labels[7][49] , \labels[7].label[40] );
tran (\labels[7][50] , \labels[7].label[41] );
tran (\labels[7][51] , \labels[7].label[42] );
tran (\labels[7][52] , \labels[7].label[43] );
tran (\labels[7][53] , \labels[7].label[44] );
tran (\labels[7][54] , \labels[7].label[45] );
tran (\labels[7][55] , \labels[7].label[46] );
tran (\labels[7][56] , \labels[7].label[47] );
tran (\labels[7][57] , \labels[7].label[48] );
tran (\labels[7][58] , \labels[7].label[49] );
tran (\labels[7][59] , \labels[7].label[50] );
tran (\labels[7][60] , \labels[7].label[51] );
tran (\labels[7][61] , \labels[7].label[52] );
tran (\labels[7][62] , \labels[7].label[53] );
tran (\labels[7][63] , \labels[7].label[54] );
tran (\labels[7][64] , \labels[7].label[55] );
tran (\labels[7][65] , \labels[7].label[56] );
tran (\labels[7][66] , \labels[7].label[57] );
tran (\labels[7][67] , \labels[7].label[58] );
tran (\labels[7][68] , \labels[7].label[59] );
tran (\labels[7][69] , \labels[7].label[60] );
tran (\labels[7][70] , \labels[7].label[61] );
tran (\labels[7][71] , \labels[7].label[62] );
tran (\labels[7][72] , \labels[7].label[63] );
tran (\labels[7][73] , \labels[7].label[64] );
tran (\labels[7][74] , \labels[7].label[65] );
tran (\labels[7][75] , \labels[7].label[66] );
tran (\labels[7][76] , \labels[7].label[67] );
tran (\labels[7][77] , \labels[7].label[68] );
tran (\labels[7][78] , \labels[7].label[69] );
tran (\labels[7][79] , \labels[7].label[70] );
tran (\labels[7][80] , \labels[7].label[71] );
tran (\labels[7][81] , \labels[7].label[72] );
tran (\labels[7][82] , \labels[7].label[73] );
tran (\labels[7][83] , \labels[7].label[74] );
tran (\labels[7][84] , \labels[7].label[75] );
tran (\labels[7][85] , \labels[7].label[76] );
tran (\labels[7][86] , \labels[7].label[77] );
tran (\labels[7][87] , \labels[7].label[78] );
tran (\labels[7][88] , \labels[7].label[79] );
tran (\labels[7][89] , \labels[7].label[80] );
tran (\labels[7][90] , \labels[7].label[81] );
tran (\labels[7][91] , \labels[7].label[82] );
tran (\labels[7][92] , \labels[7].label[83] );
tran (\labels[7][93] , \labels[7].label[84] );
tran (\labels[7][94] , \labels[7].label[85] );
tran (\labels[7][95] , \labels[7].label[86] );
tran (\labels[7][96] , \labels[7].label[87] );
tran (\labels[7][97] , \labels[7].label[88] );
tran (\labels[7][98] , \labels[7].label[89] );
tran (\labels[7][99] , \labels[7].label[90] );
tran (\labels[7][100] , \labels[7].label[91] );
tran (\labels[7][101] , \labels[7].label[92] );
tran (\labels[7][102] , \labels[7].label[93] );
tran (\labels[7][103] , \labels[7].label[94] );
tran (\labels[7][104] , \labels[7].label[95] );
tran (\labels[7][105] , \labels[7].label[96] );
tran (\labels[7][106] , \labels[7].label[97] );
tran (\labels[7][107] , \labels[7].label[98] );
tran (\labels[7][108] , \labels[7].label[99] );
tran (\labels[7][109] , \labels[7].label[100] );
tran (\labels[7][110] , \labels[7].label[101] );
tran (\labels[7][111] , \labels[7].label[102] );
tran (\labels[7][112] , \labels[7].label[103] );
tran (\labels[7][113] , \labels[7].label[104] );
tran (\labels[7][114] , \labels[7].label[105] );
tran (\labels[7][115] , \labels[7].label[106] );
tran (\labels[7][116] , \labels[7].label[107] );
tran (\labels[7][117] , \labels[7].label[108] );
tran (\labels[7][118] , \labels[7].label[109] );
tran (\labels[7][119] , \labels[7].label[110] );
tran (\labels[7][120] , \labels[7].label[111] );
tran (\labels[7][121] , \labels[7].label[112] );
tran (\labels[7][122] , \labels[7].label[113] );
tran (\labels[7][123] , \labels[7].label[114] );
tran (\labels[7][124] , \labels[7].label[115] );
tran (\labels[7][125] , \labels[7].label[116] );
tran (\labels[7][126] , \labels[7].label[117] );
tran (\labels[7][127] , \labels[7].label[118] );
tran (\labels[7][128] , \labels[7].label[119] );
tran (\labels[7][129] , \labels[7].label[120] );
tran (\labels[7][130] , \labels[7].label[121] );
tran (\labels[7][131] , \labels[7].label[122] );
tran (\labels[7][132] , \labels[7].label[123] );
tran (\labels[7][133] , \labels[7].label[124] );
tran (\labels[7][134] , \labels[7].label[125] );
tran (\labels[7][135] , \labels[7].label[126] );
tran (\labels[7][136] , \labels[7].label[127] );
tran (\labels[7][137] , \labels[7].label[128] );
tran (\labels[7][138] , \labels[7].label[129] );
tran (\labels[7][139] , \labels[7].label[130] );
tran (\labels[7][140] , \labels[7].label[131] );
tran (\labels[7][141] , \labels[7].label[132] );
tran (\labels[7][142] , \labels[7].label[133] );
tran (\labels[7][143] , \labels[7].label[134] );
tran (\labels[7][144] , \labels[7].label[135] );
tran (\labels[7][145] , \labels[7].label[136] );
tran (\labels[7][146] , \labels[7].label[137] );
tran (\labels[7][147] , \labels[7].label[138] );
tran (\labels[7][148] , \labels[7].label[139] );
tran (\labels[7][149] , \labels[7].label[140] );
tran (\labels[7][150] , \labels[7].label[141] );
tran (\labels[7][151] , \labels[7].label[142] );
tran (\labels[7][152] , \labels[7].label[143] );
tran (\labels[7][153] , \labels[7].label[144] );
tran (\labels[7][154] , \labels[7].label[145] );
tran (\labels[7][155] , \labels[7].label[146] );
tran (\labels[7][156] , \labels[7].label[147] );
tran (\labels[7][157] , \labels[7].label[148] );
tran (\labels[7][158] , \labels[7].label[149] );
tran (\labels[7][159] , \labels[7].label[150] );
tran (\labels[7][160] , \labels[7].label[151] );
tran (\labels[7][161] , \labels[7].label[152] );
tran (\labels[7][162] , \labels[7].label[153] );
tran (\labels[7][163] , \labels[7].label[154] );
tran (\labels[7][164] , \labels[7].label[155] );
tran (\labels[7][165] , \labels[7].label[156] );
tran (\labels[7][166] , \labels[7].label[157] );
tran (\labels[7][167] , \labels[7].label[158] );
tran (\labels[7][168] , \labels[7].label[159] );
tran (\labels[7][169] , \labels[7].label[160] );
tran (\labels[7][170] , \labels[7].label[161] );
tran (\labels[7][171] , \labels[7].label[162] );
tran (\labels[7][172] , \labels[7].label[163] );
tran (\labels[7][173] , \labels[7].label[164] );
tran (\labels[7][174] , \labels[7].label[165] );
tran (\labels[7][175] , \labels[7].label[166] );
tran (\labels[7][176] , \labels[7].label[167] );
tran (\labels[7][177] , \labels[7].label[168] );
tran (\labels[7][178] , \labels[7].label[169] );
tran (\labels[7][179] , \labels[7].label[170] );
tran (\labels[7][180] , \labels[7].label[171] );
tran (\labels[7][181] , \labels[7].label[172] );
tran (\labels[7][182] , \labels[7].label[173] );
tran (\labels[7][183] , \labels[7].label[174] );
tran (\labels[7][184] , \labels[7].label[175] );
tran (\labels[7][185] , \labels[7].label[176] );
tran (\labels[7][186] , \labels[7].label[177] );
tran (\labels[7][187] , \labels[7].label[178] );
tran (\labels[7][188] , \labels[7].label[179] );
tran (\labels[7][189] , \labels[7].label[180] );
tran (\labels[7][190] , \labels[7].label[181] );
tran (\labels[7][191] , \labels[7].label[182] );
tran (\labels[7][192] , \labels[7].label[183] );
tran (\labels[7][193] , \labels[7].label[184] );
tran (\labels[7][194] , \labels[7].label[185] );
tran (\labels[7][195] , \labels[7].label[186] );
tran (\labels[7][196] , \labels[7].label[187] );
tran (\labels[7][197] , \labels[7].label[188] );
tran (\labels[7][198] , \labels[7].label[189] );
tran (\labels[7][199] , \labels[7].label[190] );
tran (\labels[7][200] , \labels[7].label[191] );
tran (\labels[7][201] , \labels[7].label[192] );
tran (\labels[7][202] , \labels[7].label[193] );
tran (\labels[7][203] , \labels[7].label[194] );
tran (\labels[7][204] , \labels[7].label[195] );
tran (\labels[7][205] , \labels[7].label[196] );
tran (\labels[7][206] , \labels[7].label[197] );
tran (\labels[7][207] , \labels[7].label[198] );
tran (\labels[7][208] , \labels[7].label[199] );
tran (\labels[7][209] , \labels[7].label[200] );
tran (\labels[7][210] , \labels[7].label[201] );
tran (\labels[7][211] , \labels[7].label[202] );
tran (\labels[7][212] , \labels[7].label[203] );
tran (\labels[7][213] , \labels[7].label[204] );
tran (\labels[7][214] , \labels[7].label[205] );
tran (\labels[7][215] , \labels[7].label[206] );
tran (\labels[7][216] , \labels[7].label[207] );
tran (\labels[7][217] , \labels[7].label[208] );
tran (\labels[7][218] , \labels[7].label[209] );
tran (\labels[7][219] , \labels[7].label[210] );
tran (\labels[7][220] , \labels[7].label[211] );
tran (\labels[7][221] , \labels[7].label[212] );
tran (\labels[7][222] , \labels[7].label[213] );
tran (\labels[7][223] , \labels[7].label[214] );
tran (\labels[7][224] , \labels[7].label[215] );
tran (\labels[7][225] , \labels[7].label[216] );
tran (\labels[7][226] , \labels[7].label[217] );
tran (\labels[7][227] , \labels[7].label[218] );
tran (\labels[7][228] , \labels[7].label[219] );
tran (\labels[7][229] , \labels[7].label[220] );
tran (\labels[7][230] , \labels[7].label[221] );
tran (\labels[7][231] , \labels[7].label[222] );
tran (\labels[7][232] , \labels[7].label[223] );
tran (\labels[7][233] , \labels[7].label[224] );
tran (\labels[7][234] , \labels[7].label[225] );
tran (\labels[7][235] , \labels[7].label[226] );
tran (\labels[7][236] , \labels[7].label[227] );
tran (\labels[7][237] , \labels[7].label[228] );
tran (\labels[7][238] , \labels[7].label[229] );
tran (\labels[7][239] , \labels[7].label[230] );
tran (\labels[7][240] , \labels[7].label[231] );
tran (\labels[7][241] , \labels[7].label[232] );
tran (\labels[7][242] , \labels[7].label[233] );
tran (\labels[7][243] , \labels[7].label[234] );
tran (\labels[7][244] , \labels[7].label[235] );
tran (\labels[7][245] , \labels[7].label[236] );
tran (\labels[7][246] , \labels[7].label[237] );
tran (\labels[7][247] , \labels[7].label[238] );
tran (\labels[7][248] , \labels[7].label[239] );
tran (\labels[7][249] , \labels[7].label[240] );
tran (\labels[7][250] , \labels[7].label[241] );
tran (\labels[7][251] , \labels[7].label[242] );
tran (\labels[7][252] , \labels[7].label[243] );
tran (\labels[7][253] , \labels[7].label[244] );
tran (\labels[7][254] , \labels[7].label[245] );
tran (\labels[7][255] , \labels[7].label[246] );
tran (\labels[7][256] , \labels[7].label[247] );
tran (\labels[7][257] , \labels[7].label[248] );
tran (\labels[7][258] , \labels[7].label[249] );
tran (\labels[7][259] , \labels[7].label[250] );
tran (\labels[7][260] , \labels[7].label[251] );
tran (\labels[7][261] , \labels[7].label[252] );
tran (\labels[7][262] , \labels[7].label[253] );
tran (\labels[7][263] , \labels[7].label[254] );
tran (\labels[7][264] , \labels[7].label[255] );
tran (\labels[7][265] , \labels[7].label_size[0] );
tran (\labels[7][266] , \labels[7].label_size[1] );
tran (\labels[7][267] , \labels[7].label_size[2] );
tran (\labels[7][268] , \labels[7].label_size[3] );
tran (\labels[7][269] , \labels[7].label_size[4] );
tran (\labels[7][270] , \labels[7].label_size[5] );
tran (\labels[7][271] , \labels[7].guid_size[0] );
Q_BUF U0 ( .A(n1), .Z(cmd_il_data[287]));
Q_BUF U1 ( .A(n1), .Z(cmd_il_data[286]));
Q_BUF U2 ( .A(n1), .Z(cmd_il_data[285]));
Q_BUF U3 ( .A(n1), .Z(cmd_il_data[284]));
Q_BUF U4 ( .A(n1), .Z(cmd_il_data[283]));
Q_BUF U5 ( .A(n1), .Z(cmd_il_data[282]));
Q_BUF U6 ( .A(n1), .Z(cmd_il_data[281]));
Q_BUF U7 ( .A(n1), .Z(cmd_il_data[280]));
Q_BUF U8 ( .A(n1), .Z(cmd_il_data[279]));
Q_BUF U9 ( .A(n1), .Z(cmd_il_data[278]));
Q_BUF U10 ( .A(n1), .Z(cmd_il_data[277]));
Q_BUF U11 ( .A(n1), .Z(cmd_il_data[276]));
Q_BUF U12 ( .A(n1), .Z(cmd_il_data[275]));
Q_BUF U13 ( .A(n1), .Z(cmd_il_data[274]));
Q_BUF U14 ( .A(n1), .Z(cmd_il_data[273]));
Q_BUF U15 ( .A(n1), .Z(cmd_il_data[272]));
Q_BUF U16 ( .A(n1), .Z(cmd_il_data[271]));
Q_BUF U17 ( .A(n1), .Z(cmd_il_data[270]));
Q_BUF U18 ( .A(n1), .Z(cmd_il_data[269]));
Q_BUF U19 ( .A(n1), .Z(cmd_il_data[268]));
Q_BUF U20 ( .A(n1), .Z(cmd_il_data[267]));
Q_BUF U21 ( .A(n1), .Z(cmd_il_data[266]));
Q_BUF U22 ( .A(n1), .Z(cmd_il_data[265]));
Q_BUF U23 ( .A(n1), .Z(cmd_il_data[264]));
Q_BUF U24 ( .A(n1), .Z(cmd_il_data[263]));
Q_BUF U25 ( .A(n1), .Z(cmd_il_data[262]));
Q_BUF U26 ( .A(n1), .Z(cmd_il_data[261]));
Q_BUF U27 ( .A(n1), .Z(cmd_il_data[260]));
Q_BUF U28 ( .A(n1), .Z(cmd_il_data[259]));
Q_BUF U29 ( .A(n1), .Z(cmd_il_data[258]));
Q_BUF U30 ( .A(n1), .Z(cmd_dgl_data_size[3]));
Q_BUF U31 ( .A(n1), .Z(cmd_dgl_data_size[1]));
Q_BUF U32 ( .A(n1), .Z(hash_cmd_in[32]));
Q_BUF U33 ( .A(n1), .Z(hash_cmd_in[31]));
Q_BUF U34 ( .A(n1), .Z(hash_cmd_in[30]));
Q_BUF U35 ( .A(n1), .Z(hash_cmd_in[29]));
Q_BUF U36 ( .A(n1), .Z(hash_cmd_in[28]));
Q_BUF U37 ( .A(n1), .Z(hash_cmd_in[27]));
Q_BUF U38 ( .A(n1), .Z(hash_cmd_in[26]));
Q_BUF U39 ( .A(n1), .Z(hash_cmd_in[25]));
Q_BUF U40 ( .A(n1), .Z(hash_cmd_in[24]));
Q_BUF U41 ( .A(n1), .Z(hash_cmd_in[23]));
Q_BUF U42 ( .A(n1), .Z(hash_cmd_in[22]));
Q_BUF U43 ( .A(n1), .Z(hash_cmd_in[21]));
Q_BUF U44 ( .A(n1), .Z(hash_cmd_in[20]));
Q_BUF U45 ( .A(n1), .Z(hash_cmd_in[19]));
Q_BUF U46 ( .A(n1), .Z(hash_cmd_in[18]));
Q_BUF U47 ( .A(n1), .Z(hash_cmd_in[17]));
Q_BUF U48 ( .A(n1), .Z(hash_cmd_in[16]));
Q_BUF U49 ( .A(n1), .Z(hash_cmd_in[15]));
Q_BUF U50 ( .A(n1), .Z(hash_cmd_in[14]));
Q_BUF U51 ( .A(n1), .Z(hash_cmd_in[13]));
Q_BUF U52 ( .A(n1), .Z(hash_cmd_in[12]));
Q_BUF U53 ( .A(n1), .Z(hash_cmd_in[3]));
Q_BUF U54 ( .A(n1), .Z(hash_cmd_in[2]));
Q_BUF U55 ( .A(n1), .Z(hash_cmd_in[1]));
Q_BUF U56 ( .A(n1), .Z(_zy_simnet_cio_25));
Q_BUF U57 ( .A(n1), .Z(total_hash_size[31]));
Q_BUF U58 ( .A(n1), .Z(total_hash_size[30]));
Q_BUF U59 ( .A(n1), .Z(total_hash_size[29]));
Q_BUF U60 ( .A(n1), .Z(total_hash_size[28]));
Q_BUF U61 ( .A(n1), .Z(total_hash_size[27]));
Q_BUF U62 ( .A(n1), .Z(total_hash_size[26]));
Q_BUF U63 ( .A(n1), .Z(total_hash_size[25]));
Q_BUF U64 ( .A(n1), .Z(total_hash_size[24]));
Q_BUF U65 ( .A(n1), .Z(total_hash_size[23]));
Q_BUF U66 ( .A(n1), .Z(total_hash_size[22]));
Q_BUF U67 ( .A(n1), .Z(total_hash_size[21]));
Q_BUF U68 ( .A(n1), .Z(total_hash_size[20]));
Q_BUF U69 ( .A(n1), .Z(total_hash_size[19]));
Q_BUF U70 ( .A(n1), .Z(total_hash_size[18]));
Q_BUF U71 ( .A(n1), .Z(total_hash_size[17]));
Q_BUF U72 ( .A(n1), .Z(total_hash_size[16]));
Q_BUF U73 ( .A(n1), .Z(total_hash_size[15]));
Q_BUF U74 ( .A(n1), .Z(total_hash_size[14]));
Q_BUF U75 ( .A(n1), .Z(total_hash_size[13]));
Q_BUF U76 ( .A(n1), .Z(total_hash_size[12]));
Q_BUF U77 ( .A(n1), .Z(total_hash_size[11]));
Q_BUF U78 ( .A(n1), .Z(total_hash_size[10]));
Q_BUF U79 ( .A(n1), .Z(total_hash_size[9]));
Q_BUF U80 ( .A(n1), .Z(total_hash_size[8]));
Q_BUF U81 ( .A(n1), .Z(total_hash_size[7]));
Q_BUF U82 ( .A(iter1_kdf_key_size[31]), .Z(iter3_kdf_key_size[31]));
Q_BUF U83 ( .A(iter2_kdf_key_size[31]), .Z(iter1_kdf_key_size[31]));
Q_BUF U84 ( .A(iter1_kdf_key_size[30]), .Z(iter3_kdf_key_size[30]));
Q_BUF U85 ( .A(iter2_kdf_key_size[30]), .Z(iter1_kdf_key_size[30]));
Q_BUF U86 ( .A(iter1_kdf_key_size[29]), .Z(iter3_kdf_key_size[29]));
Q_BUF U87 ( .A(iter2_kdf_key_size[29]), .Z(iter1_kdf_key_size[29]));
Q_BUF U88 ( .A(iter1_kdf_key_size[28]), .Z(iter3_kdf_key_size[28]));
Q_BUF U89 ( .A(iter2_kdf_key_size[28]), .Z(iter1_kdf_key_size[28]));
Q_BUF U90 ( .A(iter1_kdf_key_size[27]), .Z(iter3_kdf_key_size[27]));
Q_BUF U91 ( .A(iter2_kdf_key_size[27]), .Z(iter1_kdf_key_size[27]));
Q_BUF U92 ( .A(iter1_kdf_key_size[26]), .Z(iter3_kdf_key_size[26]));
Q_BUF U93 ( .A(iter2_kdf_key_size[26]), .Z(iter1_kdf_key_size[26]));
Q_BUF U94 ( .A(iter1_kdf_key_size[25]), .Z(iter3_kdf_key_size[25]));
Q_BUF U95 ( .A(iter2_kdf_key_size[25]), .Z(iter1_kdf_key_size[25]));
Q_BUF U96 ( .A(iter1_kdf_key_size[24]), .Z(iter3_kdf_key_size[24]));
Q_BUF U97 ( .A(iter2_kdf_key_size[24]), .Z(iter1_kdf_key_size[24]));
Q_BUF U98 ( .A(iter2_kdf_key_size[23]), .Z(iter3_kdf_key_size[23]));
Q_BUF U99 ( .A(iter1_kdf_key_size[23]), .Z(iter2_kdf_key_size[23]));
Q_BUF U100 ( .A(iter1_kdf_key_size[22]), .Z(iter3_kdf_key_size[22]));
Q_BUF U101 ( .A(iter2_kdf_key_size[22]), .Z(iter1_kdf_key_size[22]));
Q_BUF U102 ( .A(iter2_kdf_key_size[21]), .Z(iter3_kdf_key_size[21]));
Q_BUF U103 ( .A(iter1_kdf_key_size[21]), .Z(iter2_kdf_key_size[21]));
Q_BUF U104 ( .A(iter2_kdf_key_size[20]), .Z(iter3_kdf_key_size[20]));
Q_BUF U105 ( .A(iter1_kdf_key_size[20]), .Z(iter2_kdf_key_size[20]));
Q_BUF U106 ( .A(iter2_kdf_key_size[19]), .Z(iter3_kdf_key_size[19]));
Q_BUF U107 ( .A(iter1_kdf_key_size[19]), .Z(iter2_kdf_key_size[19]));
Q_BUF U108 ( .A(iter2_kdf_key_size[18]), .Z(iter3_kdf_key_size[18]));
Q_BUF U109 ( .A(iter1_kdf_key_size[18]), .Z(iter2_kdf_key_size[18]));
Q_BUF U110 ( .A(iter1_kdf_key_size[17]), .Z(iter3_kdf_key_size[17]));
Q_BUF U111 ( .A(iter2_kdf_key_size[17]), .Z(iter1_kdf_key_size[17]));
Q_BUF U112 ( .A(iter1_kdf_key_size[16]), .Z(iter3_kdf_key_size[16]));
Q_BUF U113 ( .A(iter2_kdf_key_size[16]), .Z(iter1_kdf_key_size[16]));
Q_BUF U114 ( .A(iter2_kdf_key_size[15]), .Z(iter3_kdf_key_size[15]));
Q_BUF U115 ( .A(iter1_kdf_key_size[15]), .Z(iter2_kdf_key_size[15]));
Q_BUF U116 ( .A(iter1_kdf_key_size[14]), .Z(iter3_kdf_key_size[14]));
Q_BUF U117 ( .A(iter2_kdf_key_size[14]), .Z(iter1_kdf_key_size[14]));
Q_BUF U118 ( .A(iter2_kdf_key_size[13]), .Z(iter3_kdf_key_size[13]));
Q_BUF U119 ( .A(iter1_kdf_key_size[13]), .Z(iter2_kdf_key_size[13]));
Q_BUF U120 ( .A(iter1_kdf_key_size[12]), .Z(iter3_kdf_key_size[12]));
Q_BUF U121 ( .A(iter2_kdf_key_size[12]), .Z(iter1_kdf_key_size[12]));
Q_BUF U122 ( .A(iter1_kdf_key_size[11]), .Z(iter3_kdf_key_size[11]));
Q_BUF U123 ( .A(iter2_kdf_key_size[11]), .Z(iter1_kdf_key_size[11]));
Q_BUF U124 ( .A(iter2_kdf_key_size[10]), .Z(iter3_kdf_key_size[10]));
Q_BUF U125 ( .A(iter1_kdf_key_size[10]), .Z(iter2_kdf_key_size[10]));
Q_BUF U126 ( .A(iter2_kdf_key_size[9]), .Z(iter3_kdf_key_size[9]));
Q_BUF U127 ( .A(iter1_kdf_key_size[8]), .Z(iter3_kdf_key_size[8]));
Q_BUF U128 ( .A(iter1_kdf_key_size[7]), .Z(iter3_kdf_key_size[7]));
Q_BUF U129 ( .A(iter2_kdf_key_size[7]), .Z(iter1_kdf_key_size[7]));
Q_BUF U130 ( .A(iter1_kdf_key_size[6]), .Z(iter3_kdf_key_size[6]));
Q_BUF U131 ( .A(iter2_kdf_key_size[6]), .Z(iter1_kdf_key_size[6]));
Q_BUF U132 ( .A(iter2_kdf_key_size[5]), .Z(iter3_kdf_key_size[5]));
Q_BUF U133 ( .A(iter1_kdf_key_size[5]), .Z(iter2_kdf_key_size[5]));
Q_BUF U134 ( .A(iter2_kdf_key_size[4]), .Z(iter3_kdf_key_size[4]));
Q_BUF U135 ( .A(iter1_kdf_key_size[4]), .Z(iter2_kdf_key_size[4]));
Q_BUF U136 ( .A(iter1_kdf_key_size[3]), .Z(iter3_kdf_key_size[3]));
Q_BUF U137 ( .A(iter2_kdf_key_size[3]), .Z(iter1_kdf_key_size[3]));
Q_BUF U138 ( .A(iter1_kdf_key_size[2]), .Z(iter3_kdf_key_size[2]));
Q_BUF U139 ( .A(iter2_kdf_key_size[2]), .Z(iter1_kdf_key_size[2]));
Q_BUF U140 ( .A(iter2_kdf_key_size[1]), .Z(iter3_kdf_key_size[1]));
Q_BUF U141 ( .A(iter1_kdf_key_size[1]), .Z(iter2_kdf_key_size[1]));
Q_BUF U142 ( .A(iter1_kdf_key_size[0]), .Z(iter3_kdf_key_size[0]));
Q_BUF U143 ( .A(iter2_kdf_key_size[0]), .Z(iter1_kdf_key_size[0]));
Q_ASSIGN U144 ( .B(cmdfifo_kdfstream_cmd[261]), .A(hash_cmd_in[33]));
Q_BUF U145 ( .A(is_small_size), .Z(hash_cmd_in[0]));
Q_BUF U146 ( .A(moving_to_tx_data), .Z(hash_cmd_in_valid[0]));
Q_BUF U147 ( .A(total_hash_size[0]), .Z(hash_cmd_in[4]));
Q_BUF U148 ( .A(total_hash_size[1]), .Z(hash_cmd_in[5]));
Q_BUF U149 ( .A(total_hash_size[2]), .Z(hash_cmd_in[6]));
Q_BUF U150 ( .A(total_hash_size[3]), .Z(hash_cmd_in[7]));
Q_BUF U151 ( .A(total_hash_size[4]), .Z(hash_cmd_in[8]));
Q_BUF U152 ( .A(total_hash_size[5]), .Z(hash_cmd_in[9]));
Q_BUF U153 ( .A(total_hash_size[6]), .Z(hash_cmd_in[11]));
Q_BUF U154 ( .A(cmd_dgl_valid), .Z(cmd_il_valid));
Q_BUF U155 ( .A(cmd_dgl_data_size[2]), .Z(cmd_dgl_valid));
Q_BUF U156 ( .A(program_pipes), .Z(cmd_dgl_data_size[2]));
Q_BUF U157 ( .A(kdfstream_cmdfifo_ack), .Z(in_hash_eoc));
Q_AN02 U158 ( .A0(n1197), .A1(n3), .Z(n2));
Q_INV U159 ( .A(n1188), .Z(n3));
Q_AN02 U160 ( .A0(n1964), .A1(cmd_il_data_size[1]), .Z(n1963));
Q_XOR2 U161 ( .A0(n1964), .A1(cmd_il_data_size[1]), .Z(total_hash_size[1]));
Q_MX08 U162 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][271] ), .A1(\labels[1][271] ), .A2(\labels[2][271] ), .A3(\labels[3][271] ), .A4(\labels[4][271] ), .A5(\labels[5][271] ), .A6(\labels[6][271] ), .A7(\labels[7][271] ), .Z(n1188));
Q_MX08 U163 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][270] ), .A1(\labels[1][270] ), .A2(\labels[2][270] ), .A3(\labels[3][270] ), .A4(\labels[4][270] ), .A5(\labels[5][270] ), .A6(\labels[6][270] ), .A7(\labels[7][270] ), .Z(n4));
Q_MX08 U164 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][269] ), .A1(\labels[1][269] ), .A2(\labels[2][269] ), .A3(\labels[3][269] ), .A4(\labels[4][269] ), .A5(\labels[5][269] ), .A6(\labels[6][269] ), .A7(\labels[7][269] ), .Z(n5));
Q_MX08 U165 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][268] ), .A1(\labels[1][268] ), .A2(\labels[2][268] ), .A3(\labels[3][268] ), .A4(\labels[4][268] ), .A5(\labels[5][268] ), .A6(\labels[6][268] ), .A7(\labels[7][268] ), .Z(n6));
Q_MX08 U166 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][267] ), .A1(\labels[1][267] ), .A2(\labels[2][267] ), .A3(\labels[3][267] ), .A4(\labels[4][267] ), .A5(\labels[5][267] ), .A6(\labels[6][267] ), .A7(\labels[7][267] ), .Z(n7));
Q_MX08 U167 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][266] ), .A1(\labels[1][266] ), .A2(\labels[2][266] ), .A3(\labels[3][266] ), .A4(\labels[4][266] ), .A5(\labels[5][266] ), .A6(\labels[6][266] ), .A7(\labels[7][266] ), .Z(n8));
Q_MX08 U168 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][265] ), .A1(\labels[1][265] ), .A2(\labels[2][265] ), .A3(\labels[3][265] ), .A4(\labels[4][265] ), .A5(\labels[5][265] ), .A6(\labels[6][265] ), .A7(\labels[7][265] ), .Z(n9));
Q_MX08 U169 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][264] ), .A1(\labels[1][264] ), .A2(\labels[2][264] ), .A3(\labels[3][264] ), .A4(\labels[4][264] ), .A5(\labels[5][264] ), .A6(\labels[6][264] ), .A7(\labels[7][264] ), .Z(n10));
Q_MX08 U170 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][263] ), .A1(\labels[1][263] ), .A2(\labels[2][263] ), .A3(\labels[3][263] ), .A4(\labels[4][263] ), .A5(\labels[5][263] ), .A6(\labels[6][263] ), .A7(\labels[7][263] ), .Z(n11));
Q_MX08 U171 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][262] ), .A1(\labels[1][262] ), .A2(\labels[2][262] ), .A3(\labels[3][262] ), .A4(\labels[4][262] ), .A5(\labels[5][262] ), .A6(\labels[6][262] ), .A7(\labels[7][262] ), .Z(n12));
Q_MX08 U172 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][261] ), .A1(\labels[1][261] ), .A2(\labels[2][261] ), .A3(\labels[3][261] ), .A4(\labels[4][261] ), .A5(\labels[5][261] ), .A6(\labels[6][261] ), .A7(\labels[7][261] ), .Z(n13));
Q_MX08 U173 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][260] ), .A1(\labels[1][260] ), .A2(\labels[2][260] ), .A3(\labels[3][260] ), .A4(\labels[4][260] ), .A5(\labels[5][260] ), .A6(\labels[6][260] ), .A7(\labels[7][260] ), .Z(n14));
Q_MX08 U174 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][259] ), .A1(\labels[1][259] ), .A2(\labels[2][259] ), .A3(\labels[3][259] ), .A4(\labels[4][259] ), .A5(\labels[5][259] ), .A6(\labels[6][259] ), .A7(\labels[7][259] ), .Z(n15));
Q_MX08 U175 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][258] ), .A1(\labels[1][258] ), .A2(\labels[2][258] ), .A3(\labels[3][258] ), .A4(\labels[4][258] ), .A5(\labels[5][258] ), .A6(\labels[6][258] ), .A7(\labels[7][258] ), .Z(n16));
Q_MX08 U176 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][257] ), .A1(\labels[1][257] ), .A2(\labels[2][257] ), .A3(\labels[3][257] ), .A4(\labels[4][257] ), .A5(\labels[5][257] ), .A6(\labels[6][257] ), .A7(\labels[7][257] ), .Z(n17));
Q_MX08 U177 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][256] ), .A1(\labels[1][256] ), .A2(\labels[2][256] ), .A3(\labels[3][256] ), .A4(\labels[4][256] ), .A5(\labels[5][256] ), .A6(\labels[6][256] ), .A7(\labels[7][256] ), .Z(n18));
Q_MX08 U178 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][255] ), .A1(\labels[1][255] ), .A2(\labels[2][255] ), .A3(\labels[3][255] ), .A4(\labels[4][255] ), .A5(\labels[5][255] ), .A6(\labels[6][255] ), .A7(\labels[7][255] ), .Z(n19));
Q_MX08 U179 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][254] ), .A1(\labels[1][254] ), .A2(\labels[2][254] ), .A3(\labels[3][254] ), .A4(\labels[4][254] ), .A5(\labels[5][254] ), .A6(\labels[6][254] ), .A7(\labels[7][254] ), .Z(n20));
Q_MX08 U180 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][253] ), .A1(\labels[1][253] ), .A2(\labels[2][253] ), .A3(\labels[3][253] ), .A4(\labels[4][253] ), .A5(\labels[5][253] ), .A6(\labels[6][253] ), .A7(\labels[7][253] ), .Z(n21));
Q_MX08 U181 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][252] ), .A1(\labels[1][252] ), .A2(\labels[2][252] ), .A3(\labels[3][252] ), .A4(\labels[4][252] ), .A5(\labels[5][252] ), .A6(\labels[6][252] ), .A7(\labels[7][252] ), .Z(n22));
Q_MX08 U182 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][251] ), .A1(\labels[1][251] ), .A2(\labels[2][251] ), .A3(\labels[3][251] ), .A4(\labels[4][251] ), .A5(\labels[5][251] ), .A6(\labels[6][251] ), .A7(\labels[7][251] ), .Z(n23));
Q_MX08 U183 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][250] ), .A1(\labels[1][250] ), .A2(\labels[2][250] ), .A3(\labels[3][250] ), .A4(\labels[4][250] ), .A5(\labels[5][250] ), .A6(\labels[6][250] ), .A7(\labels[7][250] ), .Z(n24));
Q_MX08 U184 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][249] ), .A1(\labels[1][249] ), .A2(\labels[2][249] ), .A3(\labels[3][249] ), .A4(\labels[4][249] ), .A5(\labels[5][249] ), .A6(\labels[6][249] ), .A7(\labels[7][249] ), .Z(n25));
Q_MX08 U185 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][248] ), .A1(\labels[1][248] ), .A2(\labels[2][248] ), .A3(\labels[3][248] ), .A4(\labels[4][248] ), .A5(\labels[5][248] ), .A6(\labels[6][248] ), .A7(\labels[7][248] ), .Z(n26));
Q_MX08 U186 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][247] ), .A1(\labels[1][247] ), .A2(\labels[2][247] ), .A3(\labels[3][247] ), .A4(\labels[4][247] ), .A5(\labels[5][247] ), .A6(\labels[6][247] ), .A7(\labels[7][247] ), .Z(n27));
Q_MX08 U187 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][246] ), .A1(\labels[1][246] ), .A2(\labels[2][246] ), .A3(\labels[3][246] ), .A4(\labels[4][246] ), .A5(\labels[5][246] ), .A6(\labels[6][246] ), .A7(\labels[7][246] ), .Z(n28));
Q_MX08 U188 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][245] ), .A1(\labels[1][245] ), .A2(\labels[2][245] ), .A3(\labels[3][245] ), .A4(\labels[4][245] ), .A5(\labels[5][245] ), .A6(\labels[6][245] ), .A7(\labels[7][245] ), .Z(n29));
Q_MX08 U189 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][244] ), .A1(\labels[1][244] ), .A2(\labels[2][244] ), .A3(\labels[3][244] ), .A4(\labels[4][244] ), .A5(\labels[5][244] ), .A6(\labels[6][244] ), .A7(\labels[7][244] ), .Z(n30));
Q_MX08 U190 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][243] ), .A1(\labels[1][243] ), .A2(\labels[2][243] ), .A3(\labels[3][243] ), .A4(\labels[4][243] ), .A5(\labels[5][243] ), .A6(\labels[6][243] ), .A7(\labels[7][243] ), .Z(n31));
Q_MX08 U191 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][242] ), .A1(\labels[1][242] ), .A2(\labels[2][242] ), .A3(\labels[3][242] ), .A4(\labels[4][242] ), .A5(\labels[5][242] ), .A6(\labels[6][242] ), .A7(\labels[7][242] ), .Z(n32));
Q_MX08 U192 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][241] ), .A1(\labels[1][241] ), .A2(\labels[2][241] ), .A3(\labels[3][241] ), .A4(\labels[4][241] ), .A5(\labels[5][241] ), .A6(\labels[6][241] ), .A7(\labels[7][241] ), .Z(n33));
Q_MX08 U193 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][240] ), .A1(\labels[1][240] ), .A2(\labels[2][240] ), .A3(\labels[3][240] ), .A4(\labels[4][240] ), .A5(\labels[5][240] ), .A6(\labels[6][240] ), .A7(\labels[7][240] ), .Z(n34));
Q_MX08 U194 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][239] ), .A1(\labels[1][239] ), .A2(\labels[2][239] ), .A3(\labels[3][239] ), .A4(\labels[4][239] ), .A5(\labels[5][239] ), .A6(\labels[6][239] ), .A7(\labels[7][239] ), .Z(n35));
Q_MX08 U195 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][238] ), .A1(\labels[1][238] ), .A2(\labels[2][238] ), .A3(\labels[3][238] ), .A4(\labels[4][238] ), .A5(\labels[5][238] ), .A6(\labels[6][238] ), .A7(\labels[7][238] ), .Z(n36));
Q_MX08 U196 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][237] ), .A1(\labels[1][237] ), .A2(\labels[2][237] ), .A3(\labels[3][237] ), .A4(\labels[4][237] ), .A5(\labels[5][237] ), .A6(\labels[6][237] ), .A7(\labels[7][237] ), .Z(n37));
Q_MX08 U197 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][236] ), .A1(\labels[1][236] ), .A2(\labels[2][236] ), .A3(\labels[3][236] ), .A4(\labels[4][236] ), .A5(\labels[5][236] ), .A6(\labels[6][236] ), .A7(\labels[7][236] ), .Z(n38));
Q_MX08 U198 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][235] ), .A1(\labels[1][235] ), .A2(\labels[2][235] ), .A3(\labels[3][235] ), .A4(\labels[4][235] ), .A5(\labels[5][235] ), .A6(\labels[6][235] ), .A7(\labels[7][235] ), .Z(n39));
Q_MX08 U199 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][234] ), .A1(\labels[1][234] ), .A2(\labels[2][234] ), .A3(\labels[3][234] ), .A4(\labels[4][234] ), .A5(\labels[5][234] ), .A6(\labels[6][234] ), .A7(\labels[7][234] ), .Z(n40));
Q_MX08 U200 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][233] ), .A1(\labels[1][233] ), .A2(\labels[2][233] ), .A3(\labels[3][233] ), .A4(\labels[4][233] ), .A5(\labels[5][233] ), .A6(\labels[6][233] ), .A7(\labels[7][233] ), .Z(n41));
Q_MX08 U201 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][232] ), .A1(\labels[1][232] ), .A2(\labels[2][232] ), .A3(\labels[3][232] ), .A4(\labels[4][232] ), .A5(\labels[5][232] ), .A6(\labels[6][232] ), .A7(\labels[7][232] ), .Z(n42));
Q_MX08 U202 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][231] ), .A1(\labels[1][231] ), .A2(\labels[2][231] ), .A3(\labels[3][231] ), .A4(\labels[4][231] ), .A5(\labels[5][231] ), .A6(\labels[6][231] ), .A7(\labels[7][231] ), .Z(n43));
Q_MX08 U203 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][230] ), .A1(\labels[1][230] ), .A2(\labels[2][230] ), .A3(\labels[3][230] ), .A4(\labels[4][230] ), .A5(\labels[5][230] ), .A6(\labels[6][230] ), .A7(\labels[7][230] ), .Z(n44));
Q_MX08 U204 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][229] ), .A1(\labels[1][229] ), .A2(\labels[2][229] ), .A3(\labels[3][229] ), .A4(\labels[4][229] ), .A5(\labels[5][229] ), .A6(\labels[6][229] ), .A7(\labels[7][229] ), .Z(n45));
Q_MX08 U205 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][228] ), .A1(\labels[1][228] ), .A2(\labels[2][228] ), .A3(\labels[3][228] ), .A4(\labels[4][228] ), .A5(\labels[5][228] ), .A6(\labels[6][228] ), .A7(\labels[7][228] ), .Z(n46));
Q_MX08 U206 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][227] ), .A1(\labels[1][227] ), .A2(\labels[2][227] ), .A3(\labels[3][227] ), .A4(\labels[4][227] ), .A5(\labels[5][227] ), .A6(\labels[6][227] ), .A7(\labels[7][227] ), .Z(n47));
Q_MX08 U207 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][226] ), .A1(\labels[1][226] ), .A2(\labels[2][226] ), .A3(\labels[3][226] ), .A4(\labels[4][226] ), .A5(\labels[5][226] ), .A6(\labels[6][226] ), .A7(\labels[7][226] ), .Z(n48));
Q_MX08 U208 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][225] ), .A1(\labels[1][225] ), .A2(\labels[2][225] ), .A3(\labels[3][225] ), .A4(\labels[4][225] ), .A5(\labels[5][225] ), .A6(\labels[6][225] ), .A7(\labels[7][225] ), .Z(n49));
Q_MX08 U209 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][224] ), .A1(\labels[1][224] ), .A2(\labels[2][224] ), .A3(\labels[3][224] ), .A4(\labels[4][224] ), .A5(\labels[5][224] ), .A6(\labels[6][224] ), .A7(\labels[7][224] ), .Z(n50));
Q_MX08 U210 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][223] ), .A1(\labels[1][223] ), .A2(\labels[2][223] ), .A3(\labels[3][223] ), .A4(\labels[4][223] ), .A5(\labels[5][223] ), .A6(\labels[6][223] ), .A7(\labels[7][223] ), .Z(n51));
Q_MX08 U211 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][222] ), .A1(\labels[1][222] ), .A2(\labels[2][222] ), .A3(\labels[3][222] ), .A4(\labels[4][222] ), .A5(\labels[5][222] ), .A6(\labels[6][222] ), .A7(\labels[7][222] ), .Z(n52));
Q_MX08 U212 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][221] ), .A1(\labels[1][221] ), .A2(\labels[2][221] ), .A3(\labels[3][221] ), .A4(\labels[4][221] ), .A5(\labels[5][221] ), .A6(\labels[6][221] ), .A7(\labels[7][221] ), .Z(n53));
Q_MX08 U213 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][220] ), .A1(\labels[1][220] ), .A2(\labels[2][220] ), .A3(\labels[3][220] ), .A4(\labels[4][220] ), .A5(\labels[5][220] ), .A6(\labels[6][220] ), .A7(\labels[7][220] ), .Z(n54));
Q_MX08 U214 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][219] ), .A1(\labels[1][219] ), .A2(\labels[2][219] ), .A3(\labels[3][219] ), .A4(\labels[4][219] ), .A5(\labels[5][219] ), .A6(\labels[6][219] ), .A7(\labels[7][219] ), .Z(n55));
Q_MX08 U215 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][218] ), .A1(\labels[1][218] ), .A2(\labels[2][218] ), .A3(\labels[3][218] ), .A4(\labels[4][218] ), .A5(\labels[5][218] ), .A6(\labels[6][218] ), .A7(\labels[7][218] ), .Z(n56));
Q_MX08 U216 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][217] ), .A1(\labels[1][217] ), .A2(\labels[2][217] ), .A3(\labels[3][217] ), .A4(\labels[4][217] ), .A5(\labels[5][217] ), .A6(\labels[6][217] ), .A7(\labels[7][217] ), .Z(n57));
Q_MX08 U217 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][216] ), .A1(\labels[1][216] ), .A2(\labels[2][216] ), .A3(\labels[3][216] ), .A4(\labels[4][216] ), .A5(\labels[5][216] ), .A6(\labels[6][216] ), .A7(\labels[7][216] ), .Z(n58));
Q_MX08 U218 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][215] ), .A1(\labels[1][215] ), .A2(\labels[2][215] ), .A3(\labels[3][215] ), .A4(\labels[4][215] ), .A5(\labels[5][215] ), .A6(\labels[6][215] ), .A7(\labels[7][215] ), .Z(n59));
Q_MX08 U219 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][214] ), .A1(\labels[1][214] ), .A2(\labels[2][214] ), .A3(\labels[3][214] ), .A4(\labels[4][214] ), .A5(\labels[5][214] ), .A6(\labels[6][214] ), .A7(\labels[7][214] ), .Z(n60));
Q_MX08 U220 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][213] ), .A1(\labels[1][213] ), .A2(\labels[2][213] ), .A3(\labels[3][213] ), .A4(\labels[4][213] ), .A5(\labels[5][213] ), .A6(\labels[6][213] ), .A7(\labels[7][213] ), .Z(n61));
Q_MX08 U221 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][212] ), .A1(\labels[1][212] ), .A2(\labels[2][212] ), .A3(\labels[3][212] ), .A4(\labels[4][212] ), .A5(\labels[5][212] ), .A6(\labels[6][212] ), .A7(\labels[7][212] ), .Z(n62));
Q_MX08 U222 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][211] ), .A1(\labels[1][211] ), .A2(\labels[2][211] ), .A3(\labels[3][211] ), .A4(\labels[4][211] ), .A5(\labels[5][211] ), .A6(\labels[6][211] ), .A7(\labels[7][211] ), .Z(n63));
Q_MX08 U223 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][210] ), .A1(\labels[1][210] ), .A2(\labels[2][210] ), .A3(\labels[3][210] ), .A4(\labels[4][210] ), .A5(\labels[5][210] ), .A6(\labels[6][210] ), .A7(\labels[7][210] ), .Z(n64));
Q_MX08 U224 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][209] ), .A1(\labels[1][209] ), .A2(\labels[2][209] ), .A3(\labels[3][209] ), .A4(\labels[4][209] ), .A5(\labels[5][209] ), .A6(\labels[6][209] ), .A7(\labels[7][209] ), .Z(n65));
Q_MX08 U225 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][208] ), .A1(\labels[1][208] ), .A2(\labels[2][208] ), .A3(\labels[3][208] ), .A4(\labels[4][208] ), .A5(\labels[5][208] ), .A6(\labels[6][208] ), .A7(\labels[7][208] ), .Z(n66));
Q_MX08 U226 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][207] ), .A1(\labels[1][207] ), .A2(\labels[2][207] ), .A3(\labels[3][207] ), .A4(\labels[4][207] ), .A5(\labels[5][207] ), .A6(\labels[6][207] ), .A7(\labels[7][207] ), .Z(n67));
Q_MX08 U227 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][206] ), .A1(\labels[1][206] ), .A2(\labels[2][206] ), .A3(\labels[3][206] ), .A4(\labels[4][206] ), .A5(\labels[5][206] ), .A6(\labels[6][206] ), .A7(\labels[7][206] ), .Z(n68));
Q_MX08 U228 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][205] ), .A1(\labels[1][205] ), .A2(\labels[2][205] ), .A3(\labels[3][205] ), .A4(\labels[4][205] ), .A5(\labels[5][205] ), .A6(\labels[6][205] ), .A7(\labels[7][205] ), .Z(n69));
Q_MX08 U229 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][204] ), .A1(\labels[1][204] ), .A2(\labels[2][204] ), .A3(\labels[3][204] ), .A4(\labels[4][204] ), .A5(\labels[5][204] ), .A6(\labels[6][204] ), .A7(\labels[7][204] ), .Z(n70));
Q_MX08 U230 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][203] ), .A1(\labels[1][203] ), .A2(\labels[2][203] ), .A3(\labels[3][203] ), .A4(\labels[4][203] ), .A5(\labels[5][203] ), .A6(\labels[6][203] ), .A7(\labels[7][203] ), .Z(n71));
Q_MX08 U231 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][202] ), .A1(\labels[1][202] ), .A2(\labels[2][202] ), .A3(\labels[3][202] ), .A4(\labels[4][202] ), .A5(\labels[5][202] ), .A6(\labels[6][202] ), .A7(\labels[7][202] ), .Z(n72));
Q_MX08 U232 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][201] ), .A1(\labels[1][201] ), .A2(\labels[2][201] ), .A3(\labels[3][201] ), .A4(\labels[4][201] ), .A5(\labels[5][201] ), .A6(\labels[6][201] ), .A7(\labels[7][201] ), .Z(n73));
Q_MX08 U233 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][200] ), .A1(\labels[1][200] ), .A2(\labels[2][200] ), .A3(\labels[3][200] ), .A4(\labels[4][200] ), .A5(\labels[5][200] ), .A6(\labels[6][200] ), .A7(\labels[7][200] ), .Z(n74));
Q_MX08 U234 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][199] ), .A1(\labels[1][199] ), .A2(\labels[2][199] ), .A3(\labels[3][199] ), .A4(\labels[4][199] ), .A5(\labels[5][199] ), .A6(\labels[6][199] ), .A7(\labels[7][199] ), .Z(n75));
Q_MX08 U235 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][198] ), .A1(\labels[1][198] ), .A2(\labels[2][198] ), .A3(\labels[3][198] ), .A4(\labels[4][198] ), .A5(\labels[5][198] ), .A6(\labels[6][198] ), .A7(\labels[7][198] ), .Z(n76));
Q_MX08 U236 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][197] ), .A1(\labels[1][197] ), .A2(\labels[2][197] ), .A3(\labels[3][197] ), .A4(\labels[4][197] ), .A5(\labels[5][197] ), .A6(\labels[6][197] ), .A7(\labels[7][197] ), .Z(n77));
Q_MX08 U237 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][196] ), .A1(\labels[1][196] ), .A2(\labels[2][196] ), .A3(\labels[3][196] ), .A4(\labels[4][196] ), .A5(\labels[5][196] ), .A6(\labels[6][196] ), .A7(\labels[7][196] ), .Z(n78));
Q_MX08 U238 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][195] ), .A1(\labels[1][195] ), .A2(\labels[2][195] ), .A3(\labels[3][195] ), .A4(\labels[4][195] ), .A5(\labels[5][195] ), .A6(\labels[6][195] ), .A7(\labels[7][195] ), .Z(n79));
Q_MX08 U239 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][194] ), .A1(\labels[1][194] ), .A2(\labels[2][194] ), .A3(\labels[3][194] ), .A4(\labels[4][194] ), .A5(\labels[5][194] ), .A6(\labels[6][194] ), .A7(\labels[7][194] ), .Z(n80));
Q_MX08 U240 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][193] ), .A1(\labels[1][193] ), .A2(\labels[2][193] ), .A3(\labels[3][193] ), .A4(\labels[4][193] ), .A5(\labels[5][193] ), .A6(\labels[6][193] ), .A7(\labels[7][193] ), .Z(n81));
Q_MX08 U241 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][192] ), .A1(\labels[1][192] ), .A2(\labels[2][192] ), .A3(\labels[3][192] ), .A4(\labels[4][192] ), .A5(\labels[5][192] ), .A6(\labels[6][192] ), .A7(\labels[7][192] ), .Z(n82));
Q_MX08 U242 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][191] ), .A1(\labels[1][191] ), .A2(\labels[2][191] ), .A3(\labels[3][191] ), .A4(\labels[4][191] ), .A5(\labels[5][191] ), .A6(\labels[6][191] ), .A7(\labels[7][191] ), .Z(n83));
Q_MX08 U243 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][190] ), .A1(\labels[1][190] ), .A2(\labels[2][190] ), .A3(\labels[3][190] ), .A4(\labels[4][190] ), .A5(\labels[5][190] ), .A6(\labels[6][190] ), .A7(\labels[7][190] ), .Z(n84));
Q_MX08 U244 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][189] ), .A1(\labels[1][189] ), .A2(\labels[2][189] ), .A3(\labels[3][189] ), .A4(\labels[4][189] ), .A5(\labels[5][189] ), .A6(\labels[6][189] ), .A7(\labels[7][189] ), .Z(n85));
Q_MX08 U245 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][188] ), .A1(\labels[1][188] ), .A2(\labels[2][188] ), .A3(\labels[3][188] ), .A4(\labels[4][188] ), .A5(\labels[5][188] ), .A6(\labels[6][188] ), .A7(\labels[7][188] ), .Z(n86));
Q_MX08 U246 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][187] ), .A1(\labels[1][187] ), .A2(\labels[2][187] ), .A3(\labels[3][187] ), .A4(\labels[4][187] ), .A5(\labels[5][187] ), .A6(\labels[6][187] ), .A7(\labels[7][187] ), .Z(n87));
Q_MX08 U247 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][186] ), .A1(\labels[1][186] ), .A2(\labels[2][186] ), .A3(\labels[3][186] ), .A4(\labels[4][186] ), .A5(\labels[5][186] ), .A6(\labels[6][186] ), .A7(\labels[7][186] ), .Z(n88));
Q_MX08 U248 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][185] ), .A1(\labels[1][185] ), .A2(\labels[2][185] ), .A3(\labels[3][185] ), .A4(\labels[4][185] ), .A5(\labels[5][185] ), .A6(\labels[6][185] ), .A7(\labels[7][185] ), .Z(n89));
Q_MX08 U249 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][184] ), .A1(\labels[1][184] ), .A2(\labels[2][184] ), .A3(\labels[3][184] ), .A4(\labels[4][184] ), .A5(\labels[5][184] ), .A6(\labels[6][184] ), .A7(\labels[7][184] ), .Z(n90));
Q_MX08 U250 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][183] ), .A1(\labels[1][183] ), .A2(\labels[2][183] ), .A3(\labels[3][183] ), .A4(\labels[4][183] ), .A5(\labels[5][183] ), .A6(\labels[6][183] ), .A7(\labels[7][183] ), .Z(n91));
Q_MX08 U251 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][182] ), .A1(\labels[1][182] ), .A2(\labels[2][182] ), .A3(\labels[3][182] ), .A4(\labels[4][182] ), .A5(\labels[5][182] ), .A6(\labels[6][182] ), .A7(\labels[7][182] ), .Z(n92));
Q_MX08 U252 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][181] ), .A1(\labels[1][181] ), .A2(\labels[2][181] ), .A3(\labels[3][181] ), .A4(\labels[4][181] ), .A5(\labels[5][181] ), .A6(\labels[6][181] ), .A7(\labels[7][181] ), .Z(n93));
Q_MX08 U253 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][180] ), .A1(\labels[1][180] ), .A2(\labels[2][180] ), .A3(\labels[3][180] ), .A4(\labels[4][180] ), .A5(\labels[5][180] ), .A6(\labels[6][180] ), .A7(\labels[7][180] ), .Z(n94));
Q_MX08 U254 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][179] ), .A1(\labels[1][179] ), .A2(\labels[2][179] ), .A3(\labels[3][179] ), .A4(\labels[4][179] ), .A5(\labels[5][179] ), .A6(\labels[6][179] ), .A7(\labels[7][179] ), .Z(n95));
Q_MX08 U255 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][178] ), .A1(\labels[1][178] ), .A2(\labels[2][178] ), .A3(\labels[3][178] ), .A4(\labels[4][178] ), .A5(\labels[5][178] ), .A6(\labels[6][178] ), .A7(\labels[7][178] ), .Z(n96));
Q_MX08 U256 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][177] ), .A1(\labels[1][177] ), .A2(\labels[2][177] ), .A3(\labels[3][177] ), .A4(\labels[4][177] ), .A5(\labels[5][177] ), .A6(\labels[6][177] ), .A7(\labels[7][177] ), .Z(n97));
Q_MX08 U257 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][176] ), .A1(\labels[1][176] ), .A2(\labels[2][176] ), .A3(\labels[3][176] ), .A4(\labels[4][176] ), .A5(\labels[5][176] ), .A6(\labels[6][176] ), .A7(\labels[7][176] ), .Z(n98));
Q_MX08 U258 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][175] ), .A1(\labels[1][175] ), .A2(\labels[2][175] ), .A3(\labels[3][175] ), .A4(\labels[4][175] ), .A5(\labels[5][175] ), .A6(\labels[6][175] ), .A7(\labels[7][175] ), .Z(n99));
Q_MX08 U259 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][174] ), .A1(\labels[1][174] ), .A2(\labels[2][174] ), .A3(\labels[3][174] ), .A4(\labels[4][174] ), .A5(\labels[5][174] ), .A6(\labels[6][174] ), .A7(\labels[7][174] ), .Z(n100));
Q_MX08 U260 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][173] ), .A1(\labels[1][173] ), .A2(\labels[2][173] ), .A3(\labels[3][173] ), .A4(\labels[4][173] ), .A5(\labels[5][173] ), .A6(\labels[6][173] ), .A7(\labels[7][173] ), .Z(n101));
Q_MX08 U261 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][172] ), .A1(\labels[1][172] ), .A2(\labels[2][172] ), .A3(\labels[3][172] ), .A4(\labels[4][172] ), .A5(\labels[5][172] ), .A6(\labels[6][172] ), .A7(\labels[7][172] ), .Z(n102));
Q_MX08 U262 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][171] ), .A1(\labels[1][171] ), .A2(\labels[2][171] ), .A3(\labels[3][171] ), .A4(\labels[4][171] ), .A5(\labels[5][171] ), .A6(\labels[6][171] ), .A7(\labels[7][171] ), .Z(n103));
Q_MX08 U263 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][170] ), .A1(\labels[1][170] ), .A2(\labels[2][170] ), .A3(\labels[3][170] ), .A4(\labels[4][170] ), .A5(\labels[5][170] ), .A6(\labels[6][170] ), .A7(\labels[7][170] ), .Z(n104));
Q_MX08 U264 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][169] ), .A1(\labels[1][169] ), .A2(\labels[2][169] ), .A3(\labels[3][169] ), .A4(\labels[4][169] ), .A5(\labels[5][169] ), .A6(\labels[6][169] ), .A7(\labels[7][169] ), .Z(n105));
Q_MX08 U265 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][168] ), .A1(\labels[1][168] ), .A2(\labels[2][168] ), .A3(\labels[3][168] ), .A4(\labels[4][168] ), .A5(\labels[5][168] ), .A6(\labels[6][168] ), .A7(\labels[7][168] ), .Z(n106));
Q_MX08 U266 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][167] ), .A1(\labels[1][167] ), .A2(\labels[2][167] ), .A3(\labels[3][167] ), .A4(\labels[4][167] ), .A5(\labels[5][167] ), .A6(\labels[6][167] ), .A7(\labels[7][167] ), .Z(n107));
Q_MX08 U267 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][166] ), .A1(\labels[1][166] ), .A2(\labels[2][166] ), .A3(\labels[3][166] ), .A4(\labels[4][166] ), .A5(\labels[5][166] ), .A6(\labels[6][166] ), .A7(\labels[7][166] ), .Z(n108));
Q_MX08 U268 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][165] ), .A1(\labels[1][165] ), .A2(\labels[2][165] ), .A3(\labels[3][165] ), .A4(\labels[4][165] ), .A5(\labels[5][165] ), .A6(\labels[6][165] ), .A7(\labels[7][165] ), .Z(n109));
Q_MX08 U269 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][164] ), .A1(\labels[1][164] ), .A2(\labels[2][164] ), .A3(\labels[3][164] ), .A4(\labels[4][164] ), .A5(\labels[5][164] ), .A6(\labels[6][164] ), .A7(\labels[7][164] ), .Z(n110));
Q_MX08 U270 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][163] ), .A1(\labels[1][163] ), .A2(\labels[2][163] ), .A3(\labels[3][163] ), .A4(\labels[4][163] ), .A5(\labels[5][163] ), .A6(\labels[6][163] ), .A7(\labels[7][163] ), .Z(n111));
Q_MX08 U271 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][162] ), .A1(\labels[1][162] ), .A2(\labels[2][162] ), .A3(\labels[3][162] ), .A4(\labels[4][162] ), .A5(\labels[5][162] ), .A6(\labels[6][162] ), .A7(\labels[7][162] ), .Z(n112));
Q_MX08 U272 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][161] ), .A1(\labels[1][161] ), .A2(\labels[2][161] ), .A3(\labels[3][161] ), .A4(\labels[4][161] ), .A5(\labels[5][161] ), .A6(\labels[6][161] ), .A7(\labels[7][161] ), .Z(n113));
Q_MX08 U273 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][160] ), .A1(\labels[1][160] ), .A2(\labels[2][160] ), .A3(\labels[3][160] ), .A4(\labels[4][160] ), .A5(\labels[5][160] ), .A6(\labels[6][160] ), .A7(\labels[7][160] ), .Z(n114));
Q_MX08 U274 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][159] ), .A1(\labels[1][159] ), .A2(\labels[2][159] ), .A3(\labels[3][159] ), .A4(\labels[4][159] ), .A5(\labels[5][159] ), .A6(\labels[6][159] ), .A7(\labels[7][159] ), .Z(n115));
Q_MX08 U275 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][158] ), .A1(\labels[1][158] ), .A2(\labels[2][158] ), .A3(\labels[3][158] ), .A4(\labels[4][158] ), .A5(\labels[5][158] ), .A6(\labels[6][158] ), .A7(\labels[7][158] ), .Z(n116));
Q_MX08 U276 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][157] ), .A1(\labels[1][157] ), .A2(\labels[2][157] ), .A3(\labels[3][157] ), .A4(\labels[4][157] ), .A5(\labels[5][157] ), .A6(\labels[6][157] ), .A7(\labels[7][157] ), .Z(n117));
Q_MX08 U277 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][156] ), .A1(\labels[1][156] ), .A2(\labels[2][156] ), .A3(\labels[3][156] ), .A4(\labels[4][156] ), .A5(\labels[5][156] ), .A6(\labels[6][156] ), .A7(\labels[7][156] ), .Z(n118));
Q_MX08 U278 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][155] ), .A1(\labels[1][155] ), .A2(\labels[2][155] ), .A3(\labels[3][155] ), .A4(\labels[4][155] ), .A5(\labels[5][155] ), .A6(\labels[6][155] ), .A7(\labels[7][155] ), .Z(n119));
Q_MX08 U279 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][154] ), .A1(\labels[1][154] ), .A2(\labels[2][154] ), .A3(\labels[3][154] ), .A4(\labels[4][154] ), .A5(\labels[5][154] ), .A6(\labels[6][154] ), .A7(\labels[7][154] ), .Z(n120));
Q_MX08 U280 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][153] ), .A1(\labels[1][153] ), .A2(\labels[2][153] ), .A3(\labels[3][153] ), .A4(\labels[4][153] ), .A5(\labels[5][153] ), .A6(\labels[6][153] ), .A7(\labels[7][153] ), .Z(n121));
Q_MX08 U281 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][152] ), .A1(\labels[1][152] ), .A2(\labels[2][152] ), .A3(\labels[3][152] ), .A4(\labels[4][152] ), .A5(\labels[5][152] ), .A6(\labels[6][152] ), .A7(\labels[7][152] ), .Z(n122));
Q_MX08 U282 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][151] ), .A1(\labels[1][151] ), .A2(\labels[2][151] ), .A3(\labels[3][151] ), .A4(\labels[4][151] ), .A5(\labels[5][151] ), .A6(\labels[6][151] ), .A7(\labels[7][151] ), .Z(n123));
Q_MX08 U283 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][150] ), .A1(\labels[1][150] ), .A2(\labels[2][150] ), .A3(\labels[3][150] ), .A4(\labels[4][150] ), .A5(\labels[5][150] ), .A6(\labels[6][150] ), .A7(\labels[7][150] ), .Z(n124));
Q_MX08 U284 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][149] ), .A1(\labels[1][149] ), .A2(\labels[2][149] ), .A3(\labels[3][149] ), .A4(\labels[4][149] ), .A5(\labels[5][149] ), .A6(\labels[6][149] ), .A7(\labels[7][149] ), .Z(n125));
Q_MX08 U285 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][148] ), .A1(\labels[1][148] ), .A2(\labels[2][148] ), .A3(\labels[3][148] ), .A4(\labels[4][148] ), .A5(\labels[5][148] ), .A6(\labels[6][148] ), .A7(\labels[7][148] ), .Z(n126));
Q_MX08 U286 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][147] ), .A1(\labels[1][147] ), .A2(\labels[2][147] ), .A3(\labels[3][147] ), .A4(\labels[4][147] ), .A5(\labels[5][147] ), .A6(\labels[6][147] ), .A7(\labels[7][147] ), .Z(n127));
Q_MX08 U287 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][146] ), .A1(\labels[1][146] ), .A2(\labels[2][146] ), .A3(\labels[3][146] ), .A4(\labels[4][146] ), .A5(\labels[5][146] ), .A6(\labels[6][146] ), .A7(\labels[7][146] ), .Z(n128));
Q_MX08 U288 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][145] ), .A1(\labels[1][145] ), .A2(\labels[2][145] ), .A3(\labels[3][145] ), .A4(\labels[4][145] ), .A5(\labels[5][145] ), .A6(\labels[6][145] ), .A7(\labels[7][145] ), .Z(n129));
Q_MX08 U289 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][144] ), .A1(\labels[1][144] ), .A2(\labels[2][144] ), .A3(\labels[3][144] ), .A4(\labels[4][144] ), .A5(\labels[5][144] ), .A6(\labels[6][144] ), .A7(\labels[7][144] ), .Z(n130));
Q_MX08 U290 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][143] ), .A1(\labels[1][143] ), .A2(\labels[2][143] ), .A3(\labels[3][143] ), .A4(\labels[4][143] ), .A5(\labels[5][143] ), .A6(\labels[6][143] ), .A7(\labels[7][143] ), .Z(n131));
Q_MX08 U291 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][142] ), .A1(\labels[1][142] ), .A2(\labels[2][142] ), .A3(\labels[3][142] ), .A4(\labels[4][142] ), .A5(\labels[5][142] ), .A6(\labels[6][142] ), .A7(\labels[7][142] ), .Z(n132));
Q_MX08 U292 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][141] ), .A1(\labels[1][141] ), .A2(\labels[2][141] ), .A3(\labels[3][141] ), .A4(\labels[4][141] ), .A5(\labels[5][141] ), .A6(\labels[6][141] ), .A7(\labels[7][141] ), .Z(n133));
Q_MX08 U293 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][140] ), .A1(\labels[1][140] ), .A2(\labels[2][140] ), .A3(\labels[3][140] ), .A4(\labels[4][140] ), .A5(\labels[5][140] ), .A6(\labels[6][140] ), .A7(\labels[7][140] ), .Z(n134));
Q_MX08 U294 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][139] ), .A1(\labels[1][139] ), .A2(\labels[2][139] ), .A3(\labels[3][139] ), .A4(\labels[4][139] ), .A5(\labels[5][139] ), .A6(\labels[6][139] ), .A7(\labels[7][139] ), .Z(n135));
Q_MX08 U295 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][138] ), .A1(\labels[1][138] ), .A2(\labels[2][138] ), .A3(\labels[3][138] ), .A4(\labels[4][138] ), .A5(\labels[5][138] ), .A6(\labels[6][138] ), .A7(\labels[7][138] ), .Z(n136));
Q_MX08 U296 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][137] ), .A1(\labels[1][137] ), .A2(\labels[2][137] ), .A3(\labels[3][137] ), .A4(\labels[4][137] ), .A5(\labels[5][137] ), .A6(\labels[6][137] ), .A7(\labels[7][137] ), .Z(n137));
Q_MX08 U297 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][136] ), .A1(\labels[1][136] ), .A2(\labels[2][136] ), .A3(\labels[3][136] ), .A4(\labels[4][136] ), .A5(\labels[5][136] ), .A6(\labels[6][136] ), .A7(\labels[7][136] ), .Z(n138));
Q_MX08 U298 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][135] ), .A1(\labels[1][135] ), .A2(\labels[2][135] ), .A3(\labels[3][135] ), .A4(\labels[4][135] ), .A5(\labels[5][135] ), .A6(\labels[6][135] ), .A7(\labels[7][135] ), .Z(n139));
Q_MX08 U299 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][134] ), .A1(\labels[1][134] ), .A2(\labels[2][134] ), .A3(\labels[3][134] ), .A4(\labels[4][134] ), .A5(\labels[5][134] ), .A6(\labels[6][134] ), .A7(\labels[7][134] ), .Z(n140));
Q_MX08 U300 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][133] ), .A1(\labels[1][133] ), .A2(\labels[2][133] ), .A3(\labels[3][133] ), .A4(\labels[4][133] ), .A5(\labels[5][133] ), .A6(\labels[6][133] ), .A7(\labels[7][133] ), .Z(n141));
Q_MX08 U301 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][132] ), .A1(\labels[1][132] ), .A2(\labels[2][132] ), .A3(\labels[3][132] ), .A4(\labels[4][132] ), .A5(\labels[5][132] ), .A6(\labels[6][132] ), .A7(\labels[7][132] ), .Z(n142));
Q_MX08 U302 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][131] ), .A1(\labels[1][131] ), .A2(\labels[2][131] ), .A3(\labels[3][131] ), .A4(\labels[4][131] ), .A5(\labels[5][131] ), .A6(\labels[6][131] ), .A7(\labels[7][131] ), .Z(n143));
Q_MX08 U303 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][130] ), .A1(\labels[1][130] ), .A2(\labels[2][130] ), .A3(\labels[3][130] ), .A4(\labels[4][130] ), .A5(\labels[5][130] ), .A6(\labels[6][130] ), .A7(\labels[7][130] ), .Z(n144));
Q_MX08 U304 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][129] ), .A1(\labels[1][129] ), .A2(\labels[2][129] ), .A3(\labels[3][129] ), .A4(\labels[4][129] ), .A5(\labels[5][129] ), .A6(\labels[6][129] ), .A7(\labels[7][129] ), .Z(n145));
Q_MX08 U305 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][128] ), .A1(\labels[1][128] ), .A2(\labels[2][128] ), .A3(\labels[3][128] ), .A4(\labels[4][128] ), .A5(\labels[5][128] ), .A6(\labels[6][128] ), .A7(\labels[7][128] ), .Z(n146));
Q_MX08 U306 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][127] ), .A1(\labels[1][127] ), .A2(\labels[2][127] ), .A3(\labels[3][127] ), .A4(\labels[4][127] ), .A5(\labels[5][127] ), .A6(\labels[6][127] ), .A7(\labels[7][127] ), .Z(n147));
Q_MX08 U307 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][126] ), .A1(\labels[1][126] ), .A2(\labels[2][126] ), .A3(\labels[3][126] ), .A4(\labels[4][126] ), .A5(\labels[5][126] ), .A6(\labels[6][126] ), .A7(\labels[7][126] ), .Z(n148));
Q_MX08 U308 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][125] ), .A1(\labels[1][125] ), .A2(\labels[2][125] ), .A3(\labels[3][125] ), .A4(\labels[4][125] ), .A5(\labels[5][125] ), .A6(\labels[6][125] ), .A7(\labels[7][125] ), .Z(n149));
Q_MX08 U309 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][124] ), .A1(\labels[1][124] ), .A2(\labels[2][124] ), .A3(\labels[3][124] ), .A4(\labels[4][124] ), .A5(\labels[5][124] ), .A6(\labels[6][124] ), .A7(\labels[7][124] ), .Z(n150));
Q_MX08 U310 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][123] ), .A1(\labels[1][123] ), .A2(\labels[2][123] ), .A3(\labels[3][123] ), .A4(\labels[4][123] ), .A5(\labels[5][123] ), .A6(\labels[6][123] ), .A7(\labels[7][123] ), .Z(n151));
Q_MX08 U311 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][122] ), .A1(\labels[1][122] ), .A2(\labels[2][122] ), .A3(\labels[3][122] ), .A4(\labels[4][122] ), .A5(\labels[5][122] ), .A6(\labels[6][122] ), .A7(\labels[7][122] ), .Z(n152));
Q_MX08 U312 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][121] ), .A1(\labels[1][121] ), .A2(\labels[2][121] ), .A3(\labels[3][121] ), .A4(\labels[4][121] ), .A5(\labels[5][121] ), .A6(\labels[6][121] ), .A7(\labels[7][121] ), .Z(n153));
Q_MX08 U313 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][120] ), .A1(\labels[1][120] ), .A2(\labels[2][120] ), .A3(\labels[3][120] ), .A4(\labels[4][120] ), .A5(\labels[5][120] ), .A6(\labels[6][120] ), .A7(\labels[7][120] ), .Z(n154));
Q_MX08 U314 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][119] ), .A1(\labels[1][119] ), .A2(\labels[2][119] ), .A3(\labels[3][119] ), .A4(\labels[4][119] ), .A5(\labels[5][119] ), .A6(\labels[6][119] ), .A7(\labels[7][119] ), .Z(n155));
Q_MX08 U315 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][118] ), .A1(\labels[1][118] ), .A2(\labels[2][118] ), .A3(\labels[3][118] ), .A4(\labels[4][118] ), .A5(\labels[5][118] ), .A6(\labels[6][118] ), .A7(\labels[7][118] ), .Z(n156));
Q_MX08 U316 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][117] ), .A1(\labels[1][117] ), .A2(\labels[2][117] ), .A3(\labels[3][117] ), .A4(\labels[4][117] ), .A5(\labels[5][117] ), .A6(\labels[6][117] ), .A7(\labels[7][117] ), .Z(n157));
Q_MX08 U317 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][116] ), .A1(\labels[1][116] ), .A2(\labels[2][116] ), .A3(\labels[3][116] ), .A4(\labels[4][116] ), .A5(\labels[5][116] ), .A6(\labels[6][116] ), .A7(\labels[7][116] ), .Z(n158));
Q_MX08 U318 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][115] ), .A1(\labels[1][115] ), .A2(\labels[2][115] ), .A3(\labels[3][115] ), .A4(\labels[4][115] ), .A5(\labels[5][115] ), .A6(\labels[6][115] ), .A7(\labels[7][115] ), .Z(n159));
Q_MX08 U319 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][114] ), .A1(\labels[1][114] ), .A2(\labels[2][114] ), .A3(\labels[3][114] ), .A4(\labels[4][114] ), .A5(\labels[5][114] ), .A6(\labels[6][114] ), .A7(\labels[7][114] ), .Z(n160));
Q_MX08 U320 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][113] ), .A1(\labels[1][113] ), .A2(\labels[2][113] ), .A3(\labels[3][113] ), .A4(\labels[4][113] ), .A5(\labels[5][113] ), .A6(\labels[6][113] ), .A7(\labels[7][113] ), .Z(n161));
Q_MX08 U321 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][112] ), .A1(\labels[1][112] ), .A2(\labels[2][112] ), .A3(\labels[3][112] ), .A4(\labels[4][112] ), .A5(\labels[5][112] ), .A6(\labels[6][112] ), .A7(\labels[7][112] ), .Z(n162));
Q_MX08 U322 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][111] ), .A1(\labels[1][111] ), .A2(\labels[2][111] ), .A3(\labels[3][111] ), .A4(\labels[4][111] ), .A5(\labels[5][111] ), .A6(\labels[6][111] ), .A7(\labels[7][111] ), .Z(n163));
Q_MX08 U323 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][110] ), .A1(\labels[1][110] ), .A2(\labels[2][110] ), .A3(\labels[3][110] ), .A4(\labels[4][110] ), .A5(\labels[5][110] ), .A6(\labels[6][110] ), .A7(\labels[7][110] ), .Z(n164));
Q_MX08 U324 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][109] ), .A1(\labels[1][109] ), .A2(\labels[2][109] ), .A3(\labels[3][109] ), .A4(\labels[4][109] ), .A5(\labels[5][109] ), .A6(\labels[6][109] ), .A7(\labels[7][109] ), .Z(n165));
Q_MX08 U325 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][108] ), .A1(\labels[1][108] ), .A2(\labels[2][108] ), .A3(\labels[3][108] ), .A4(\labels[4][108] ), .A5(\labels[5][108] ), .A6(\labels[6][108] ), .A7(\labels[7][108] ), .Z(n166));
Q_MX08 U326 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][107] ), .A1(\labels[1][107] ), .A2(\labels[2][107] ), .A3(\labels[3][107] ), .A4(\labels[4][107] ), .A5(\labels[5][107] ), .A6(\labels[6][107] ), .A7(\labels[7][107] ), .Z(n167));
Q_MX08 U327 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][106] ), .A1(\labels[1][106] ), .A2(\labels[2][106] ), .A3(\labels[3][106] ), .A4(\labels[4][106] ), .A5(\labels[5][106] ), .A6(\labels[6][106] ), .A7(\labels[7][106] ), .Z(n168));
Q_MX08 U328 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][105] ), .A1(\labels[1][105] ), .A2(\labels[2][105] ), .A3(\labels[3][105] ), .A4(\labels[4][105] ), .A5(\labels[5][105] ), .A6(\labels[6][105] ), .A7(\labels[7][105] ), .Z(n169));
Q_MX08 U329 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][104] ), .A1(\labels[1][104] ), .A2(\labels[2][104] ), .A3(\labels[3][104] ), .A4(\labels[4][104] ), .A5(\labels[5][104] ), .A6(\labels[6][104] ), .A7(\labels[7][104] ), .Z(n170));
Q_MX08 U330 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][103] ), .A1(\labels[1][103] ), .A2(\labels[2][103] ), .A3(\labels[3][103] ), .A4(\labels[4][103] ), .A5(\labels[5][103] ), .A6(\labels[6][103] ), .A7(\labels[7][103] ), .Z(n171));
Q_MX08 U331 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][102] ), .A1(\labels[1][102] ), .A2(\labels[2][102] ), .A3(\labels[3][102] ), .A4(\labels[4][102] ), .A5(\labels[5][102] ), .A6(\labels[6][102] ), .A7(\labels[7][102] ), .Z(n172));
Q_MX08 U332 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][101] ), .A1(\labels[1][101] ), .A2(\labels[2][101] ), .A3(\labels[3][101] ), .A4(\labels[4][101] ), .A5(\labels[5][101] ), .A6(\labels[6][101] ), .A7(\labels[7][101] ), .Z(n173));
Q_MX08 U333 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][100] ), .A1(\labels[1][100] ), .A2(\labels[2][100] ), .A3(\labels[3][100] ), .A4(\labels[4][100] ), .A5(\labels[5][100] ), .A6(\labels[6][100] ), .A7(\labels[7][100] ), .Z(n174));
Q_MX08 U334 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][99] ), .A1(\labels[1][99] ), .A2(\labels[2][99] ), .A3(\labels[3][99] ), .A4(\labels[4][99] ), .A5(\labels[5][99] ), .A6(\labels[6][99] ), .A7(\labels[7][99] ), .Z(n175));
Q_MX08 U335 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][98] ), .A1(\labels[1][98] ), .A2(\labels[2][98] ), .A3(\labels[3][98] ), .A4(\labels[4][98] ), .A5(\labels[5][98] ), .A6(\labels[6][98] ), .A7(\labels[7][98] ), .Z(n176));
Q_MX08 U336 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][97] ), .A1(\labels[1][97] ), .A2(\labels[2][97] ), .A3(\labels[3][97] ), .A4(\labels[4][97] ), .A5(\labels[5][97] ), .A6(\labels[6][97] ), .A7(\labels[7][97] ), .Z(n177));
Q_MX08 U337 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][96] ), .A1(\labels[1][96] ), .A2(\labels[2][96] ), .A3(\labels[3][96] ), .A4(\labels[4][96] ), .A5(\labels[5][96] ), .A6(\labels[6][96] ), .A7(\labels[7][96] ), .Z(n178));
Q_MX08 U338 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][95] ), .A1(\labels[1][95] ), .A2(\labels[2][95] ), .A3(\labels[3][95] ), .A4(\labels[4][95] ), .A5(\labels[5][95] ), .A6(\labels[6][95] ), .A7(\labels[7][95] ), .Z(n179));
Q_MX08 U339 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][94] ), .A1(\labels[1][94] ), .A2(\labels[2][94] ), .A3(\labels[3][94] ), .A4(\labels[4][94] ), .A5(\labels[5][94] ), .A6(\labels[6][94] ), .A7(\labels[7][94] ), .Z(n180));
Q_MX08 U340 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][93] ), .A1(\labels[1][93] ), .A2(\labels[2][93] ), .A3(\labels[3][93] ), .A4(\labels[4][93] ), .A5(\labels[5][93] ), .A6(\labels[6][93] ), .A7(\labels[7][93] ), .Z(n181));
Q_MX08 U341 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][92] ), .A1(\labels[1][92] ), .A2(\labels[2][92] ), .A3(\labels[3][92] ), .A4(\labels[4][92] ), .A5(\labels[5][92] ), .A6(\labels[6][92] ), .A7(\labels[7][92] ), .Z(n182));
Q_MX08 U342 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][91] ), .A1(\labels[1][91] ), .A2(\labels[2][91] ), .A3(\labels[3][91] ), .A4(\labels[4][91] ), .A5(\labels[5][91] ), .A6(\labels[6][91] ), .A7(\labels[7][91] ), .Z(n183));
Q_MX08 U343 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][90] ), .A1(\labels[1][90] ), .A2(\labels[2][90] ), .A3(\labels[3][90] ), .A4(\labels[4][90] ), .A5(\labels[5][90] ), .A6(\labels[6][90] ), .A7(\labels[7][90] ), .Z(n184));
Q_MX08 U344 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][89] ), .A1(\labels[1][89] ), .A2(\labels[2][89] ), .A3(\labels[3][89] ), .A4(\labels[4][89] ), .A5(\labels[5][89] ), .A6(\labels[6][89] ), .A7(\labels[7][89] ), .Z(n185));
Q_MX08 U345 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][88] ), .A1(\labels[1][88] ), .A2(\labels[2][88] ), .A3(\labels[3][88] ), .A4(\labels[4][88] ), .A5(\labels[5][88] ), .A6(\labels[6][88] ), .A7(\labels[7][88] ), .Z(n186));
Q_MX08 U346 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][87] ), .A1(\labels[1][87] ), .A2(\labels[2][87] ), .A3(\labels[3][87] ), .A4(\labels[4][87] ), .A5(\labels[5][87] ), .A6(\labels[6][87] ), .A7(\labels[7][87] ), .Z(n187));
Q_MX08 U347 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][86] ), .A1(\labels[1][86] ), .A2(\labels[2][86] ), .A3(\labels[3][86] ), .A4(\labels[4][86] ), .A5(\labels[5][86] ), .A6(\labels[6][86] ), .A7(\labels[7][86] ), .Z(n188));
Q_MX08 U348 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][85] ), .A1(\labels[1][85] ), .A2(\labels[2][85] ), .A3(\labels[3][85] ), .A4(\labels[4][85] ), .A5(\labels[5][85] ), .A6(\labels[6][85] ), .A7(\labels[7][85] ), .Z(n189));
Q_MX08 U349 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][84] ), .A1(\labels[1][84] ), .A2(\labels[2][84] ), .A3(\labels[3][84] ), .A4(\labels[4][84] ), .A5(\labels[5][84] ), .A6(\labels[6][84] ), .A7(\labels[7][84] ), .Z(n190));
Q_MX08 U350 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][83] ), .A1(\labels[1][83] ), .A2(\labels[2][83] ), .A3(\labels[3][83] ), .A4(\labels[4][83] ), .A5(\labels[5][83] ), .A6(\labels[6][83] ), .A7(\labels[7][83] ), .Z(n191));
Q_MX08 U351 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][82] ), .A1(\labels[1][82] ), .A2(\labels[2][82] ), .A3(\labels[3][82] ), .A4(\labels[4][82] ), .A5(\labels[5][82] ), .A6(\labels[6][82] ), .A7(\labels[7][82] ), .Z(n192));
Q_MX08 U352 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][81] ), .A1(\labels[1][81] ), .A2(\labels[2][81] ), .A3(\labels[3][81] ), .A4(\labels[4][81] ), .A5(\labels[5][81] ), .A6(\labels[6][81] ), .A7(\labels[7][81] ), .Z(n193));
Q_MX08 U353 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][80] ), .A1(\labels[1][80] ), .A2(\labels[2][80] ), .A3(\labels[3][80] ), .A4(\labels[4][80] ), .A5(\labels[5][80] ), .A6(\labels[6][80] ), .A7(\labels[7][80] ), .Z(n194));
Q_MX08 U354 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][79] ), .A1(\labels[1][79] ), .A2(\labels[2][79] ), .A3(\labels[3][79] ), .A4(\labels[4][79] ), .A5(\labels[5][79] ), .A6(\labels[6][79] ), .A7(\labels[7][79] ), .Z(n195));
Q_MX08 U355 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][78] ), .A1(\labels[1][78] ), .A2(\labels[2][78] ), .A3(\labels[3][78] ), .A4(\labels[4][78] ), .A5(\labels[5][78] ), .A6(\labels[6][78] ), .A7(\labels[7][78] ), .Z(n196));
Q_MX08 U356 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][77] ), .A1(\labels[1][77] ), .A2(\labels[2][77] ), .A3(\labels[3][77] ), .A4(\labels[4][77] ), .A5(\labels[5][77] ), .A6(\labels[6][77] ), .A7(\labels[7][77] ), .Z(n197));
Q_MX08 U357 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][76] ), .A1(\labels[1][76] ), .A2(\labels[2][76] ), .A3(\labels[3][76] ), .A4(\labels[4][76] ), .A5(\labels[5][76] ), .A6(\labels[6][76] ), .A7(\labels[7][76] ), .Z(n198));
Q_MX08 U358 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][75] ), .A1(\labels[1][75] ), .A2(\labels[2][75] ), .A3(\labels[3][75] ), .A4(\labels[4][75] ), .A5(\labels[5][75] ), .A6(\labels[6][75] ), .A7(\labels[7][75] ), .Z(n199));
Q_MX08 U359 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][74] ), .A1(\labels[1][74] ), .A2(\labels[2][74] ), .A3(\labels[3][74] ), .A4(\labels[4][74] ), .A5(\labels[5][74] ), .A6(\labels[6][74] ), .A7(\labels[7][74] ), .Z(n200));
Q_MX08 U360 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][73] ), .A1(\labels[1][73] ), .A2(\labels[2][73] ), .A3(\labels[3][73] ), .A4(\labels[4][73] ), .A5(\labels[5][73] ), .A6(\labels[6][73] ), .A7(\labels[7][73] ), .Z(n201));
Q_MX08 U361 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][72] ), .A1(\labels[1][72] ), .A2(\labels[2][72] ), .A3(\labels[3][72] ), .A4(\labels[4][72] ), .A5(\labels[5][72] ), .A6(\labels[6][72] ), .A7(\labels[7][72] ), .Z(n202));
Q_MX08 U362 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][71] ), .A1(\labels[1][71] ), .A2(\labels[2][71] ), .A3(\labels[3][71] ), .A4(\labels[4][71] ), .A5(\labels[5][71] ), .A6(\labels[6][71] ), .A7(\labels[7][71] ), .Z(n203));
Q_MX08 U363 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][70] ), .A1(\labels[1][70] ), .A2(\labels[2][70] ), .A3(\labels[3][70] ), .A4(\labels[4][70] ), .A5(\labels[5][70] ), .A6(\labels[6][70] ), .A7(\labels[7][70] ), .Z(n204));
Q_MX08 U364 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][69] ), .A1(\labels[1][69] ), .A2(\labels[2][69] ), .A3(\labels[3][69] ), .A4(\labels[4][69] ), .A5(\labels[5][69] ), .A6(\labels[6][69] ), .A7(\labels[7][69] ), .Z(n205));
Q_MX08 U365 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][68] ), .A1(\labels[1][68] ), .A2(\labels[2][68] ), .A3(\labels[3][68] ), .A4(\labels[4][68] ), .A5(\labels[5][68] ), .A6(\labels[6][68] ), .A7(\labels[7][68] ), .Z(n206));
Q_MX08 U366 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][67] ), .A1(\labels[1][67] ), .A2(\labels[2][67] ), .A3(\labels[3][67] ), .A4(\labels[4][67] ), .A5(\labels[5][67] ), .A6(\labels[6][67] ), .A7(\labels[7][67] ), .Z(n207));
Q_MX08 U367 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][66] ), .A1(\labels[1][66] ), .A2(\labels[2][66] ), .A3(\labels[3][66] ), .A4(\labels[4][66] ), .A5(\labels[5][66] ), .A6(\labels[6][66] ), .A7(\labels[7][66] ), .Z(n208));
Q_MX08 U368 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][65] ), .A1(\labels[1][65] ), .A2(\labels[2][65] ), .A3(\labels[3][65] ), .A4(\labels[4][65] ), .A5(\labels[5][65] ), .A6(\labels[6][65] ), .A7(\labels[7][65] ), .Z(n209));
Q_MX08 U369 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][64] ), .A1(\labels[1][64] ), .A2(\labels[2][64] ), .A3(\labels[3][64] ), .A4(\labels[4][64] ), .A5(\labels[5][64] ), .A6(\labels[6][64] ), .A7(\labels[7][64] ), .Z(n210));
Q_MX08 U370 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][63] ), .A1(\labels[1][63] ), .A2(\labels[2][63] ), .A3(\labels[3][63] ), .A4(\labels[4][63] ), .A5(\labels[5][63] ), .A6(\labels[6][63] ), .A7(\labels[7][63] ), .Z(n211));
Q_MX08 U371 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][62] ), .A1(\labels[1][62] ), .A2(\labels[2][62] ), .A3(\labels[3][62] ), .A4(\labels[4][62] ), .A5(\labels[5][62] ), .A6(\labels[6][62] ), .A7(\labels[7][62] ), .Z(n212));
Q_MX08 U372 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][61] ), .A1(\labels[1][61] ), .A2(\labels[2][61] ), .A3(\labels[3][61] ), .A4(\labels[4][61] ), .A5(\labels[5][61] ), .A6(\labels[6][61] ), .A7(\labels[7][61] ), .Z(n213));
Q_MX08 U373 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][60] ), .A1(\labels[1][60] ), .A2(\labels[2][60] ), .A3(\labels[3][60] ), .A4(\labels[4][60] ), .A5(\labels[5][60] ), .A6(\labels[6][60] ), .A7(\labels[7][60] ), .Z(n214));
Q_MX08 U374 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][59] ), .A1(\labels[1][59] ), .A2(\labels[2][59] ), .A3(\labels[3][59] ), .A4(\labels[4][59] ), .A5(\labels[5][59] ), .A6(\labels[6][59] ), .A7(\labels[7][59] ), .Z(n215));
Q_MX08 U375 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][58] ), .A1(\labels[1][58] ), .A2(\labels[2][58] ), .A3(\labels[3][58] ), .A4(\labels[4][58] ), .A5(\labels[5][58] ), .A6(\labels[6][58] ), .A7(\labels[7][58] ), .Z(n216));
Q_MX08 U376 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][57] ), .A1(\labels[1][57] ), .A2(\labels[2][57] ), .A3(\labels[3][57] ), .A4(\labels[4][57] ), .A5(\labels[5][57] ), .A6(\labels[6][57] ), .A7(\labels[7][57] ), .Z(n217));
Q_MX08 U377 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][56] ), .A1(\labels[1][56] ), .A2(\labels[2][56] ), .A3(\labels[3][56] ), .A4(\labels[4][56] ), .A5(\labels[5][56] ), .A6(\labels[6][56] ), .A7(\labels[7][56] ), .Z(n218));
Q_MX08 U378 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][55] ), .A1(\labels[1][55] ), .A2(\labels[2][55] ), .A3(\labels[3][55] ), .A4(\labels[4][55] ), .A5(\labels[5][55] ), .A6(\labels[6][55] ), .A7(\labels[7][55] ), .Z(n219));
Q_MX08 U379 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][54] ), .A1(\labels[1][54] ), .A2(\labels[2][54] ), .A3(\labels[3][54] ), .A4(\labels[4][54] ), .A5(\labels[5][54] ), .A6(\labels[6][54] ), .A7(\labels[7][54] ), .Z(n220));
Q_MX08 U380 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][53] ), .A1(\labels[1][53] ), .A2(\labels[2][53] ), .A3(\labels[3][53] ), .A4(\labels[4][53] ), .A5(\labels[5][53] ), .A6(\labels[6][53] ), .A7(\labels[7][53] ), .Z(n221));
Q_MX08 U381 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][52] ), .A1(\labels[1][52] ), .A2(\labels[2][52] ), .A3(\labels[3][52] ), .A4(\labels[4][52] ), .A5(\labels[5][52] ), .A6(\labels[6][52] ), .A7(\labels[7][52] ), .Z(n222));
Q_MX08 U382 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][51] ), .A1(\labels[1][51] ), .A2(\labels[2][51] ), .A3(\labels[3][51] ), .A4(\labels[4][51] ), .A5(\labels[5][51] ), .A6(\labels[6][51] ), .A7(\labels[7][51] ), .Z(n223));
Q_MX08 U383 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][50] ), .A1(\labels[1][50] ), .A2(\labels[2][50] ), .A3(\labels[3][50] ), .A4(\labels[4][50] ), .A5(\labels[5][50] ), .A6(\labels[6][50] ), .A7(\labels[7][50] ), .Z(n224));
Q_MX08 U384 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][49] ), .A1(\labels[1][49] ), .A2(\labels[2][49] ), .A3(\labels[3][49] ), .A4(\labels[4][49] ), .A5(\labels[5][49] ), .A6(\labels[6][49] ), .A7(\labels[7][49] ), .Z(n225));
Q_MX08 U385 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][48] ), .A1(\labels[1][48] ), .A2(\labels[2][48] ), .A3(\labels[3][48] ), .A4(\labels[4][48] ), .A5(\labels[5][48] ), .A6(\labels[6][48] ), .A7(\labels[7][48] ), .Z(n226));
Q_MX08 U386 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][47] ), .A1(\labels[1][47] ), .A2(\labels[2][47] ), .A3(\labels[3][47] ), .A4(\labels[4][47] ), .A5(\labels[5][47] ), .A6(\labels[6][47] ), .A7(\labels[7][47] ), .Z(n227));
Q_MX08 U387 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][46] ), .A1(\labels[1][46] ), .A2(\labels[2][46] ), .A3(\labels[3][46] ), .A4(\labels[4][46] ), .A5(\labels[5][46] ), .A6(\labels[6][46] ), .A7(\labels[7][46] ), .Z(n228));
Q_MX08 U388 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][45] ), .A1(\labels[1][45] ), .A2(\labels[2][45] ), .A3(\labels[3][45] ), .A4(\labels[4][45] ), .A5(\labels[5][45] ), .A6(\labels[6][45] ), .A7(\labels[7][45] ), .Z(n229));
Q_MX08 U389 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][44] ), .A1(\labels[1][44] ), .A2(\labels[2][44] ), .A3(\labels[3][44] ), .A4(\labels[4][44] ), .A5(\labels[5][44] ), .A6(\labels[6][44] ), .A7(\labels[7][44] ), .Z(n230));
Q_MX08 U390 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][43] ), .A1(\labels[1][43] ), .A2(\labels[2][43] ), .A3(\labels[3][43] ), .A4(\labels[4][43] ), .A5(\labels[5][43] ), .A6(\labels[6][43] ), .A7(\labels[7][43] ), .Z(n231));
Q_MX08 U391 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][42] ), .A1(\labels[1][42] ), .A2(\labels[2][42] ), .A3(\labels[3][42] ), .A4(\labels[4][42] ), .A5(\labels[5][42] ), .A6(\labels[6][42] ), .A7(\labels[7][42] ), .Z(n232));
Q_MX08 U392 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][41] ), .A1(\labels[1][41] ), .A2(\labels[2][41] ), .A3(\labels[3][41] ), .A4(\labels[4][41] ), .A5(\labels[5][41] ), .A6(\labels[6][41] ), .A7(\labels[7][41] ), .Z(n233));
Q_MX08 U393 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][40] ), .A1(\labels[1][40] ), .A2(\labels[2][40] ), .A3(\labels[3][40] ), .A4(\labels[4][40] ), .A5(\labels[5][40] ), .A6(\labels[6][40] ), .A7(\labels[7][40] ), .Z(n234));
Q_MX08 U394 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][39] ), .A1(\labels[1][39] ), .A2(\labels[2][39] ), .A3(\labels[3][39] ), .A4(\labels[4][39] ), .A5(\labels[5][39] ), .A6(\labels[6][39] ), .A7(\labels[7][39] ), .Z(n235));
Q_MX08 U395 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][38] ), .A1(\labels[1][38] ), .A2(\labels[2][38] ), .A3(\labels[3][38] ), .A4(\labels[4][38] ), .A5(\labels[5][38] ), .A6(\labels[6][38] ), .A7(\labels[7][38] ), .Z(n236));
Q_MX08 U396 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][37] ), .A1(\labels[1][37] ), .A2(\labels[2][37] ), .A3(\labels[3][37] ), .A4(\labels[4][37] ), .A5(\labels[5][37] ), .A6(\labels[6][37] ), .A7(\labels[7][37] ), .Z(n237));
Q_MX08 U397 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][36] ), .A1(\labels[1][36] ), .A2(\labels[2][36] ), .A3(\labels[3][36] ), .A4(\labels[4][36] ), .A5(\labels[5][36] ), .A6(\labels[6][36] ), .A7(\labels[7][36] ), .Z(n238));
Q_MX08 U398 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][35] ), .A1(\labels[1][35] ), .A2(\labels[2][35] ), .A3(\labels[3][35] ), .A4(\labels[4][35] ), .A5(\labels[5][35] ), .A6(\labels[6][35] ), .A7(\labels[7][35] ), .Z(n239));
Q_MX08 U399 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][34] ), .A1(\labels[1][34] ), .A2(\labels[2][34] ), .A3(\labels[3][34] ), .A4(\labels[4][34] ), .A5(\labels[5][34] ), .A6(\labels[6][34] ), .A7(\labels[7][34] ), .Z(n240));
Q_MX08 U400 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][33] ), .A1(\labels[1][33] ), .A2(\labels[2][33] ), .A3(\labels[3][33] ), .A4(\labels[4][33] ), .A5(\labels[5][33] ), .A6(\labels[6][33] ), .A7(\labels[7][33] ), .Z(n241));
Q_MX08 U401 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][32] ), .A1(\labels[1][32] ), .A2(\labels[2][32] ), .A3(\labels[3][32] ), .A4(\labels[4][32] ), .A5(\labels[5][32] ), .A6(\labels[6][32] ), .A7(\labels[7][32] ), .Z(n242));
Q_MX08 U402 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][31] ), .A1(\labels[1][31] ), .A2(\labels[2][31] ), .A3(\labels[3][31] ), .A4(\labels[4][31] ), .A5(\labels[5][31] ), .A6(\labels[6][31] ), .A7(\labels[7][31] ), .Z(n243));
Q_MX08 U403 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][30] ), .A1(\labels[1][30] ), .A2(\labels[2][30] ), .A3(\labels[3][30] ), .A4(\labels[4][30] ), .A5(\labels[5][30] ), .A6(\labels[6][30] ), .A7(\labels[7][30] ), .Z(n244));
Q_MX08 U404 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][29] ), .A1(\labels[1][29] ), .A2(\labels[2][29] ), .A3(\labels[3][29] ), .A4(\labels[4][29] ), .A5(\labels[5][29] ), .A6(\labels[6][29] ), .A7(\labels[7][29] ), .Z(n245));
Q_MX08 U405 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][28] ), .A1(\labels[1][28] ), .A2(\labels[2][28] ), .A3(\labels[3][28] ), .A4(\labels[4][28] ), .A5(\labels[5][28] ), .A6(\labels[6][28] ), .A7(\labels[7][28] ), .Z(n246));
Q_MX08 U406 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][27] ), .A1(\labels[1][27] ), .A2(\labels[2][27] ), .A3(\labels[3][27] ), .A4(\labels[4][27] ), .A5(\labels[5][27] ), .A6(\labels[6][27] ), .A7(\labels[7][27] ), .Z(n247));
Q_MX08 U407 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][26] ), .A1(\labels[1][26] ), .A2(\labels[2][26] ), .A3(\labels[3][26] ), .A4(\labels[4][26] ), .A5(\labels[5][26] ), .A6(\labels[6][26] ), .A7(\labels[7][26] ), .Z(n248));
Q_MX08 U408 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][25] ), .A1(\labels[1][25] ), .A2(\labels[2][25] ), .A3(\labels[3][25] ), .A4(\labels[4][25] ), .A5(\labels[5][25] ), .A6(\labels[6][25] ), .A7(\labels[7][25] ), .Z(n249));
Q_MX08 U409 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][24] ), .A1(\labels[1][24] ), .A2(\labels[2][24] ), .A3(\labels[3][24] ), .A4(\labels[4][24] ), .A5(\labels[5][24] ), .A6(\labels[6][24] ), .A7(\labels[7][24] ), .Z(n250));
Q_MX08 U410 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][23] ), .A1(\labels[1][23] ), .A2(\labels[2][23] ), .A3(\labels[3][23] ), .A4(\labels[4][23] ), .A5(\labels[5][23] ), .A6(\labels[6][23] ), .A7(\labels[7][23] ), .Z(n251));
Q_MX08 U411 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][22] ), .A1(\labels[1][22] ), .A2(\labels[2][22] ), .A3(\labels[3][22] ), .A4(\labels[4][22] ), .A5(\labels[5][22] ), .A6(\labels[6][22] ), .A7(\labels[7][22] ), .Z(n252));
Q_MX08 U412 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][21] ), .A1(\labels[1][21] ), .A2(\labels[2][21] ), .A3(\labels[3][21] ), .A4(\labels[4][21] ), .A5(\labels[5][21] ), .A6(\labels[6][21] ), .A7(\labels[7][21] ), .Z(n253));
Q_MX08 U413 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][20] ), .A1(\labels[1][20] ), .A2(\labels[2][20] ), .A3(\labels[3][20] ), .A4(\labels[4][20] ), .A5(\labels[5][20] ), .A6(\labels[6][20] ), .A7(\labels[7][20] ), .Z(n254));
Q_MX08 U414 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][19] ), .A1(\labels[1][19] ), .A2(\labels[2][19] ), .A3(\labels[3][19] ), .A4(\labels[4][19] ), .A5(\labels[5][19] ), .A6(\labels[6][19] ), .A7(\labels[7][19] ), .Z(n255));
Q_MX08 U415 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][18] ), .A1(\labels[1][18] ), .A2(\labels[2][18] ), .A3(\labels[3][18] ), .A4(\labels[4][18] ), .A5(\labels[5][18] ), .A6(\labels[6][18] ), .A7(\labels[7][18] ), .Z(n256));
Q_MX08 U416 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][17] ), .A1(\labels[1][17] ), .A2(\labels[2][17] ), .A3(\labels[3][17] ), .A4(\labels[4][17] ), .A5(\labels[5][17] ), .A6(\labels[6][17] ), .A7(\labels[7][17] ), .Z(n257));
Q_MX08 U417 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][16] ), .A1(\labels[1][16] ), .A2(\labels[2][16] ), .A3(\labels[3][16] ), .A4(\labels[4][16] ), .A5(\labels[5][16] ), .A6(\labels[6][16] ), .A7(\labels[7][16] ), .Z(n258));
Q_MX08 U418 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][15] ), .A1(\labels[1][15] ), .A2(\labels[2][15] ), .A3(\labels[3][15] ), .A4(\labels[4][15] ), .A5(\labels[5][15] ), .A6(\labels[6][15] ), .A7(\labels[7][15] ), .Z(n259));
Q_MX08 U419 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][14] ), .A1(\labels[1][14] ), .A2(\labels[2][14] ), .A3(\labels[3][14] ), .A4(\labels[4][14] ), .A5(\labels[5][14] ), .A6(\labels[6][14] ), .A7(\labels[7][14] ), .Z(n260));
Q_MX08 U420 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][13] ), .A1(\labels[1][13] ), .A2(\labels[2][13] ), .A3(\labels[3][13] ), .A4(\labels[4][13] ), .A5(\labels[5][13] ), .A6(\labels[6][13] ), .A7(\labels[7][13] ), .Z(n261));
Q_MX08 U421 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][12] ), .A1(\labels[1][12] ), .A2(\labels[2][12] ), .A3(\labels[3][12] ), .A4(\labels[4][12] ), .A5(\labels[5][12] ), .A6(\labels[6][12] ), .A7(\labels[7][12] ), .Z(n262));
Q_MX08 U422 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][11] ), .A1(\labels[1][11] ), .A2(\labels[2][11] ), .A3(\labels[3][11] ), .A4(\labels[4][11] ), .A5(\labels[5][11] ), .A6(\labels[6][11] ), .A7(\labels[7][11] ), .Z(n263));
Q_MX08 U423 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][10] ), .A1(\labels[1][10] ), .A2(\labels[2][10] ), .A3(\labels[3][10] ), .A4(\labels[4][10] ), .A5(\labels[5][10] ), .A6(\labels[6][10] ), .A7(\labels[7][10] ), .Z(n264));
Q_MX08 U424 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][9] ), .A1(\labels[1][9] ), .A2(\labels[2][9] ), .A3(\labels[3][9] ), .A4(\labels[4][9] ), .A5(\labels[5][9] ), .A6(\labels[6][9] ), .A7(\labels[7][9] ), .Z(n265));
Q_MX08 U425 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][8] ), .A1(\labels[1][8] ), .A2(\labels[2][8] ), .A3(\labels[3][8] ), .A4(\labels[4][8] ), .A5(\labels[5][8] ), .A6(\labels[6][8] ), .A7(\labels[7][8] ), .Z(n1187));
Q_MX08 U426 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][7] ), .A1(\labels[1][7] ), .A2(\labels[2][7] ), .A3(\labels[3][7] ), .A4(\labels[4][7] ), .A5(\labels[5][7] ), .A6(\labels[6][7] ), .A7(\labels[7][7] ), .Z(n266));
Q_MX08 U427 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][6] ), .A1(\labels[1][6] ), .A2(\labels[2][6] ), .A3(\labels[3][6] ), .A4(\labels[4][6] ), .A5(\labels[5][6] ), .A6(\labels[6][6] ), .A7(\labels[7][6] ), .Z(n267));
Q_MX08 U428 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][5] ), .A1(\labels[1][5] ), .A2(\labels[2][5] ), .A3(\labels[3][5] ), .A4(\labels[4][5] ), .A5(\labels[5][5] ), .A6(\labels[6][5] ), .A7(\labels[7][5] ), .Z(n268));
Q_MX08 U429 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][4] ), .A1(\labels[1][4] ), .A2(\labels[2][4] ), .A3(\labels[3][4] ), .A4(\labels[4][4] ), .A5(\labels[5][4] ), .A6(\labels[6][4] ), .A7(\labels[7][4] ), .Z(n269));
Q_MX08 U430 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][3] ), .A1(\labels[1][3] ), .A2(\labels[2][3] ), .A3(\labels[3][3] ), .A4(\labels[4][3] ), .A5(\labels[5][3] ), .A6(\labels[6][3] ), .A7(\labels[7][3] ), .Z(n270));
Q_MX08 U431 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][2] ), .A1(\labels[1][2] ), .A2(\labels[2][2] ), .A3(\labels[3][2] ), .A4(\labels[4][2] ), .A5(\labels[5][2] ), .A6(\labels[6][2] ), .A7(\labels[7][2] ), .Z(n271));
Q_MX08 U432 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][1] ), .A1(\labels[1][1] ), .A2(\labels[2][1] ), .A3(\labels[3][1] ), .A4(\labels[4][1] ), .A5(\labels[5][1] ), .A6(\labels[6][1] ), .A7(\labels[7][1] ), .Z(n272));
Q_MX08 U433 ( .S0(cmdfifo_kdfstream_cmd[2]), .S1(cmdfifo_kdfstream_cmd[3]), .S2(cmdfifo_kdfstream_cmd[4]), .A0(\labels[0][0] ), .A1(\labels[1][0] ), .A2(\labels[2][0] ), .A3(\labels[3][0] ), .A4(\labels[4][0] ), .A5(\labels[5][0] ), .A6(\labels[6][0] ), .A7(\labels[7][0] ), .Z(n273));
Q_MX02 U434 ( .S(\pipe_array_ack[1][0] ), .A0(n881), .A1(n274), .Z(in_hash_byte_accumulator[4]));
Q_MX02 U435 ( .S(\pipe_array_ack[1][0] ), .A0(n882), .A1(n276), .Z(in_hash_byte_accumulator[3]));
Q_MX02 U436 ( .S(\pipe_array_ack[1][0] ), .A0(n883), .A1(n277), .Z(in_hash_byte_accumulator[2]));
Q_MX02 U437 ( .S(\pipe_array_ack[1][0] ), .A0(n884), .A1(n279), .Z(in_hash_byte_accumulator[1]));
Q_MX02 U438 ( .S(\pipe_array_ack[1][0] ), .A0(n885), .A1(n281), .Z(in_hash_byte_accumulator[0]));
Q_AD02 U439 ( .CI(n278), .A0(\pipe_array_ack_num_bytes[1][2] ), .A1(\pipe_array_ack_num_bytes[1][3] ), .B0(n883), .B1(n882), .S0(n277), .S1(n276), .CO(n275));
Q_AD01 U440 ( .CI(n884), .A0(\pipe_array_ack_num_bytes[1][1] ), .B0(n280), .S(n279), .CO(n278));
Q_XOR3 U441 ( .A0(\pipe_array_ack_num_bytes[1][4] ), .A1(n881), .A2(n275), .Z(n274));
Q_AD01HF U442 ( .A0(\pipe_array_ack_num_bytes[1][0] ), .B0(n885), .S(n281), .CO(n280));
Q_OR02 U443 ( .A0(n950), .A1(n2036), .Z(in_hash_data[63]));
Q_OR02 U444 ( .A0(n951), .A1(n2035), .Z(in_hash_data[62]));
Q_OR02 U445 ( .A0(n952), .A1(n2034), .Z(in_hash_data[61]));
Q_OR02 U446 ( .A0(n953), .A1(n2033), .Z(in_hash_data[60]));
Q_OR02 U447 ( .A0(n954), .A1(n2032), .Z(in_hash_data[59]));
Q_OR02 U448 ( .A0(n955), .A1(n2031), .Z(in_hash_data[58]));
Q_OR02 U449 ( .A0(n956), .A1(n2030), .Z(in_hash_data[57]));
Q_OR02 U450 ( .A0(n957), .A1(n2029), .Z(in_hash_data[56]));
Q_OR02 U451 ( .A0(n958), .A1(n2028), .Z(in_hash_data[55]));
Q_OR02 U452 ( .A0(n959), .A1(n2027), .Z(in_hash_data[54]));
Q_OR02 U453 ( .A0(n960), .A1(n2026), .Z(in_hash_data[53]));
Q_OR02 U454 ( .A0(n961), .A1(n2025), .Z(in_hash_data[52]));
Q_OR02 U455 ( .A0(n962), .A1(n2024), .Z(in_hash_data[51]));
Q_OR02 U456 ( .A0(n963), .A1(n2023), .Z(in_hash_data[50]));
Q_OR02 U457 ( .A0(n964), .A1(n2022), .Z(in_hash_data[49]));
Q_OR02 U458 ( .A0(n965), .A1(n2021), .Z(in_hash_data[48]));
Q_OR02 U459 ( .A0(n966), .A1(n2020), .Z(in_hash_data[47]));
Q_OR02 U460 ( .A0(n967), .A1(n2019), .Z(in_hash_data[46]));
Q_OR02 U461 ( .A0(n968), .A1(n2018), .Z(in_hash_data[45]));
Q_OR02 U462 ( .A0(n969), .A1(n2017), .Z(in_hash_data[44]));
Q_OR02 U463 ( .A0(n970), .A1(n2016), .Z(in_hash_data[43]));
Q_OR02 U464 ( .A0(n971), .A1(n2015), .Z(in_hash_data[42]));
Q_OR02 U465 ( .A0(n972), .A1(n2014), .Z(in_hash_data[41]));
Q_OR02 U466 ( .A0(n973), .A1(n2013), .Z(in_hash_data[40]));
Q_OR02 U467 ( .A0(n974), .A1(n2012), .Z(in_hash_data[39]));
Q_OR02 U468 ( .A0(n975), .A1(n2011), .Z(in_hash_data[38]));
Q_OR02 U469 ( .A0(n976), .A1(n2010), .Z(in_hash_data[37]));
Q_OR02 U470 ( .A0(n977), .A1(n2009), .Z(in_hash_data[36]));
Q_OR02 U471 ( .A0(n978), .A1(n2008), .Z(in_hash_data[35]));
Q_OR02 U472 ( .A0(n979), .A1(n2007), .Z(in_hash_data[34]));
Q_OR02 U473 ( .A0(n980), .A1(n2006), .Z(in_hash_data[33]));
Q_OR02 U474 ( .A0(n981), .A1(n2005), .Z(in_hash_data[32]));
Q_OR02 U475 ( .A0(n982), .A1(n2004), .Z(in_hash_data[31]));
Q_OR02 U476 ( .A0(n983), .A1(n2003), .Z(in_hash_data[30]));
Q_OR02 U477 ( .A0(n984), .A1(n2002), .Z(in_hash_data[29]));
Q_OR02 U478 ( .A0(n985), .A1(n2001), .Z(in_hash_data[28]));
Q_OR02 U479 ( .A0(n986), .A1(n2000), .Z(in_hash_data[27]));
Q_OR02 U480 ( .A0(n987), .A1(n1999), .Z(in_hash_data[26]));
Q_OR02 U481 ( .A0(n988), .A1(n1998), .Z(in_hash_data[25]));
Q_OR02 U482 ( .A0(n989), .A1(n1997), .Z(in_hash_data[24]));
Q_OR02 U483 ( .A0(n990), .A1(n1996), .Z(in_hash_data[23]));
Q_OR02 U484 ( .A0(n991), .A1(n1995), .Z(in_hash_data[22]));
Q_OR02 U485 ( .A0(n992), .A1(n1994), .Z(in_hash_data[21]));
Q_OR02 U486 ( .A0(n993), .A1(n1993), .Z(in_hash_data[20]));
Q_OR02 U487 ( .A0(n994), .A1(n1992), .Z(in_hash_data[19]));
Q_OR02 U488 ( .A0(n995), .A1(n1991), .Z(in_hash_data[18]));
Q_OR02 U489 ( .A0(n996), .A1(n1990), .Z(in_hash_data[17]));
Q_OR02 U490 ( .A0(n997), .A1(n1989), .Z(in_hash_data[16]));
Q_OR02 U491 ( .A0(n998), .A1(n1988), .Z(in_hash_data[15]));
Q_OR02 U492 ( .A0(n999), .A1(n1987), .Z(in_hash_data[14]));
Q_OR02 U493 ( .A0(n1000), .A1(n1986), .Z(in_hash_data[13]));
Q_OR02 U494 ( .A0(n1001), .A1(n1985), .Z(in_hash_data[12]));
Q_OR02 U495 ( .A0(n1002), .A1(n1984), .Z(in_hash_data[11]));
Q_OR02 U496 ( .A0(n1003), .A1(n1983), .Z(in_hash_data[10]));
Q_OR02 U497 ( .A0(n1004), .A1(n1982), .Z(in_hash_data[9]));
Q_OR02 U498 ( .A0(n1005), .A1(n1981), .Z(in_hash_data[8]));
Q_OR02 U499 ( .A0(n1006), .A1(n1980), .Z(in_hash_data[7]));
Q_OR02 U500 ( .A0(n1007), .A1(n1979), .Z(in_hash_data[6]));
Q_OR02 U501 ( .A0(n1008), .A1(n1978), .Z(in_hash_data[5]));
Q_OR02 U502 ( .A0(n1009), .A1(n1977), .Z(in_hash_data[4]));
Q_OR02 U503 ( .A0(n1010), .A1(n1976), .Z(in_hash_data[3]));
Q_OR02 U504 ( .A0(n1011), .A1(n1975), .Z(in_hash_data[2]));
Q_OR02 U505 ( .A0(n1012), .A1(n1974), .Z(in_hash_data[1]));
Q_OR02 U506 ( .A0(n1013), .A1(n1973), .Z(in_hash_data[0]));
Q_AN03 U507 ( .A0(n346), .A1(n348), .A2(\pipe_array_ack[1][0] ), .Z(n2036));
Q_AN03 U508 ( .A0(n346), .A1(n349), .A2(\pipe_array_ack[1][0] ), .Z(n2035));
Q_AN03 U509 ( .A0(n346), .A1(n350), .A2(\pipe_array_ack[1][0] ), .Z(n2034));
Q_AN03 U510 ( .A0(n346), .A1(n351), .A2(\pipe_array_ack[1][0] ), .Z(n2033));
Q_AN03 U511 ( .A0(n346), .A1(n352), .A2(\pipe_array_ack[1][0] ), .Z(n2032));
Q_AN03 U512 ( .A0(n346), .A1(n353), .A2(\pipe_array_ack[1][0] ), .Z(n2031));
Q_AN03 U513 ( .A0(n346), .A1(n354), .A2(\pipe_array_ack[1][0] ), .Z(n2030));
Q_AN03 U514 ( .A0(n346), .A1(n355), .A2(\pipe_array_ack[1][0] ), .Z(n2029));
Q_AN03 U515 ( .A0(n346), .A1(n356), .A2(\pipe_array_ack[1][0] ), .Z(n2028));
Q_AN03 U516 ( .A0(n346), .A1(n357), .A2(\pipe_array_ack[1][0] ), .Z(n2027));
Q_AN03 U517 ( .A0(n346), .A1(n358), .A2(\pipe_array_ack[1][0] ), .Z(n2026));
Q_AN03 U518 ( .A0(n346), .A1(n359), .A2(\pipe_array_ack[1][0] ), .Z(n2025));
Q_AN03 U519 ( .A0(n346), .A1(n360), .A2(\pipe_array_ack[1][0] ), .Z(n2024));
Q_AN03 U520 ( .A0(n346), .A1(n361), .A2(\pipe_array_ack[1][0] ), .Z(n2023));
Q_AN03 U521 ( .A0(n346), .A1(n362), .A2(\pipe_array_ack[1][0] ), .Z(n2022));
Q_AN03 U522 ( .A0(n346), .A1(n363), .A2(\pipe_array_ack[1][0] ), .Z(n2021));
Q_AN03 U523 ( .A0(n346), .A1(n364), .A2(\pipe_array_ack[1][0] ), .Z(n2020));
Q_AN03 U524 ( .A0(n346), .A1(n365), .A2(\pipe_array_ack[1][0] ), .Z(n2019));
Q_AN03 U525 ( .A0(n346), .A1(n366), .A2(\pipe_array_ack[1][0] ), .Z(n2018));
Q_AN03 U526 ( .A0(n346), .A1(n367), .A2(\pipe_array_ack[1][0] ), .Z(n2017));
Q_AN03 U527 ( .A0(n346), .A1(n368), .A2(\pipe_array_ack[1][0] ), .Z(n2016));
Q_AN03 U528 ( .A0(n346), .A1(n369), .A2(\pipe_array_ack[1][0] ), .Z(n2015));
Q_AN03 U529 ( .A0(n346), .A1(n370), .A2(\pipe_array_ack[1][0] ), .Z(n2014));
Q_AN03 U530 ( .A0(n346), .A1(n371), .A2(\pipe_array_ack[1][0] ), .Z(n2013));
Q_AN03 U531 ( .A0(n346), .A1(n372), .A2(\pipe_array_ack[1][0] ), .Z(n2012));
Q_AN03 U532 ( .A0(n346), .A1(n373), .A2(\pipe_array_ack[1][0] ), .Z(n2011));
Q_AN03 U533 ( .A0(n346), .A1(n374), .A2(\pipe_array_ack[1][0] ), .Z(n2010));
Q_AN03 U534 ( .A0(n346), .A1(n375), .A2(\pipe_array_ack[1][0] ), .Z(n2009));
Q_AN03 U535 ( .A0(n346), .A1(n376), .A2(\pipe_array_ack[1][0] ), .Z(n2008));
Q_AN03 U536 ( .A0(n346), .A1(n377), .A2(\pipe_array_ack[1][0] ), .Z(n2007));
Q_AN03 U537 ( .A0(n346), .A1(n378), .A2(\pipe_array_ack[1][0] ), .Z(n2006));
Q_AN03 U538 ( .A0(n346), .A1(n379), .A2(\pipe_array_ack[1][0] ), .Z(n2005));
Q_AN03 U539 ( .A0(n346), .A1(n380), .A2(\pipe_array_ack[1][0] ), .Z(n2004));
Q_AN03 U540 ( .A0(n346), .A1(n381), .A2(\pipe_array_ack[1][0] ), .Z(n2003));
Q_AN03 U541 ( .A0(n346), .A1(n382), .A2(\pipe_array_ack[1][0] ), .Z(n2002));
Q_AN03 U542 ( .A0(n346), .A1(n383), .A2(\pipe_array_ack[1][0] ), .Z(n2001));
Q_AN03 U543 ( .A0(n346), .A1(n384), .A2(\pipe_array_ack[1][0] ), .Z(n2000));
Q_AN03 U544 ( .A0(n346), .A1(n385), .A2(\pipe_array_ack[1][0] ), .Z(n1999));
Q_AN03 U545 ( .A0(n346), .A1(n386), .A2(\pipe_array_ack[1][0] ), .Z(n1998));
Q_AN03 U546 ( .A0(n346), .A1(n387), .A2(\pipe_array_ack[1][0] ), .Z(n1997));
Q_AN03 U547 ( .A0(n346), .A1(n388), .A2(\pipe_array_ack[1][0] ), .Z(n1996));
Q_AN03 U548 ( .A0(n346), .A1(n389), .A2(\pipe_array_ack[1][0] ), .Z(n1995));
Q_AN03 U549 ( .A0(n346), .A1(n390), .A2(\pipe_array_ack[1][0] ), .Z(n1994));
Q_AN03 U550 ( .A0(n346), .A1(n391), .A2(\pipe_array_ack[1][0] ), .Z(n1993));
Q_AN03 U551 ( .A0(n346), .A1(n392), .A2(\pipe_array_ack[1][0] ), .Z(n1992));
Q_AN03 U552 ( .A0(n346), .A1(n393), .A2(\pipe_array_ack[1][0] ), .Z(n1991));
Q_AN03 U553 ( .A0(n346), .A1(n394), .A2(\pipe_array_ack[1][0] ), .Z(n1990));
Q_AN03 U554 ( .A0(n346), .A1(n395), .A2(\pipe_array_ack[1][0] ), .Z(n1989));
Q_AN03 U555 ( .A0(n346), .A1(n396), .A2(\pipe_array_ack[1][0] ), .Z(n1988));
Q_AN03 U556 ( .A0(n346), .A1(n397), .A2(\pipe_array_ack[1][0] ), .Z(n1987));
Q_AN03 U557 ( .A0(n346), .A1(n398), .A2(\pipe_array_ack[1][0] ), .Z(n1986));
Q_AN03 U558 ( .A0(n346), .A1(n399), .A2(\pipe_array_ack[1][0] ), .Z(n1985));
Q_AN03 U559 ( .A0(n346), .A1(n400), .A2(\pipe_array_ack[1][0] ), .Z(n1984));
Q_AN03 U560 ( .A0(n346), .A1(n401), .A2(\pipe_array_ack[1][0] ), .Z(n1983));
Q_AN03 U561 ( .A0(n346), .A1(n402), .A2(\pipe_array_ack[1][0] ), .Z(n1982));
Q_AN03 U562 ( .A0(n346), .A1(n403), .A2(\pipe_array_ack[1][0] ), .Z(n1981));
Q_AN03 U563 ( .A0(n346), .A1(n404), .A2(\pipe_array_ack[1][0] ), .Z(n1980));
Q_AN03 U564 ( .A0(n346), .A1(n405), .A2(\pipe_array_ack[1][0] ), .Z(n1979));
Q_AN03 U565 ( .A0(n346), .A1(n406), .A2(\pipe_array_ack[1][0] ), .Z(n1978));
Q_AN03 U566 ( .A0(n346), .A1(n407), .A2(\pipe_array_ack[1][0] ), .Z(n1977));
Q_AN03 U567 ( .A0(n346), .A1(n408), .A2(\pipe_array_ack[1][0] ), .Z(n1976));
Q_AN03 U568 ( .A0(n346), .A1(n409), .A2(\pipe_array_ack[1][0] ), .Z(n1975));
Q_AN03 U569 ( .A0(n346), .A1(n410), .A2(\pipe_array_ack[1][0] ), .Z(n1974));
Q_AN03 U570 ( .A0(n346), .A1(n411), .A2(\pipe_array_ack[1][0] ), .Z(n1973));
Q_INV U571 ( .A(n881), .Z(n346));
Q_AN03 U572 ( .A0(n347), .A1(n412), .A2(n346), .Z(n282));
Q_AN03 U573 ( .A0(n347), .A1(n413), .A2(n346), .Z(n283));
Q_AN03 U574 ( .A0(n347), .A1(n414), .A2(n346), .Z(n284));
Q_AN03 U575 ( .A0(n347), .A1(n415), .A2(n346), .Z(n285));
Q_AN03 U576 ( .A0(n347), .A1(n416), .A2(n346), .Z(n286));
Q_AN03 U577 ( .A0(n347), .A1(n417), .A2(n346), .Z(n287));
Q_AN03 U578 ( .A0(n347), .A1(n418), .A2(n346), .Z(n288));
Q_AN03 U579 ( .A0(n347), .A1(n419), .A2(n346), .Z(n289));
Q_AN03 U580 ( .A0(n347), .A1(n420), .A2(n346), .Z(n290));
Q_AN03 U581 ( .A0(n347), .A1(n421), .A2(n346), .Z(n291));
Q_AN03 U582 ( .A0(n347), .A1(n422), .A2(n346), .Z(n292));
Q_AN03 U583 ( .A0(n347), .A1(n423), .A2(n346), .Z(n293));
Q_AN03 U584 ( .A0(n347), .A1(n424), .A2(n346), .Z(n294));
Q_AN03 U585 ( .A0(n347), .A1(n425), .A2(n346), .Z(n295));
Q_AN03 U586 ( .A0(n347), .A1(n426), .A2(n346), .Z(n296));
Q_AN03 U587 ( .A0(n347), .A1(n427), .A2(n346), .Z(n297));
Q_AN03 U588 ( .A0(n347), .A1(n428), .A2(n346), .Z(n298));
Q_AN03 U589 ( .A0(n347), .A1(n429), .A2(n346), .Z(n299));
Q_AN03 U590 ( .A0(n347), .A1(n430), .A2(n346), .Z(n300));
Q_AN03 U591 ( .A0(n347), .A1(n431), .A2(n346), .Z(n301));
Q_AN03 U592 ( .A0(n347), .A1(n432), .A2(n346), .Z(n302));
Q_AN03 U593 ( .A0(n347), .A1(n433), .A2(n346), .Z(n303));
Q_AN03 U594 ( .A0(n347), .A1(n434), .A2(n346), .Z(n304));
Q_AN03 U595 ( .A0(n347), .A1(n435), .A2(n346), .Z(n305));
Q_AN03 U596 ( .A0(n347), .A1(n436), .A2(n346), .Z(n306));
Q_AN03 U597 ( .A0(n347), .A1(n437), .A2(n346), .Z(n307));
Q_AN03 U598 ( .A0(n347), .A1(n438), .A2(n346), .Z(n308));
Q_AN03 U599 ( .A0(n347), .A1(n439), .A2(n346), .Z(n309));
Q_AN03 U600 ( .A0(n347), .A1(n440), .A2(n346), .Z(n310));
Q_AN03 U601 ( .A0(n347), .A1(n441), .A2(n346), .Z(n311));
Q_AN03 U602 ( .A0(n347), .A1(n442), .A2(n346), .Z(n312));
Q_AN03 U603 ( .A0(n347), .A1(n443), .A2(n346), .Z(n313));
Q_AN03 U604 ( .A0(n347), .A1(n445), .A2(n346), .Z(n314));
Q_AN03 U605 ( .A0(n347), .A1(n446), .A2(n346), .Z(n315));
Q_AN03 U606 ( .A0(n347), .A1(n447), .A2(n346), .Z(n316));
Q_AN03 U607 ( .A0(n347), .A1(n448), .A2(n346), .Z(n317));
Q_AN03 U608 ( .A0(n347), .A1(n449), .A2(n346), .Z(n318));
Q_AN03 U609 ( .A0(n347), .A1(n450), .A2(n346), .Z(n319));
Q_AN03 U610 ( .A0(n347), .A1(n451), .A2(n346), .Z(n320));
Q_AN03 U611 ( .A0(n347), .A1(n452), .A2(n346), .Z(n321));
Q_AN03 U612 ( .A0(n347), .A1(n453), .A2(n346), .Z(n322));
Q_AN03 U613 ( .A0(n347), .A1(n454), .A2(n346), .Z(n323));
Q_AN03 U614 ( .A0(n347), .A1(n455), .A2(n346), .Z(n324));
Q_AN03 U615 ( .A0(n347), .A1(n456), .A2(n346), .Z(n325));
Q_AN03 U616 ( .A0(n347), .A1(n457), .A2(n346), .Z(n326));
Q_AN03 U617 ( .A0(n347), .A1(n458), .A2(n346), .Z(n327));
Q_AN03 U618 ( .A0(n347), .A1(n459), .A2(n346), .Z(n328));
Q_AN03 U619 ( .A0(n347), .A1(n460), .A2(n346), .Z(n329));
Q_AN03 U620 ( .A0(n347), .A1(n461), .A2(n346), .Z(n330));
Q_AN03 U621 ( .A0(n347), .A1(n462), .A2(n346), .Z(n331));
Q_AN03 U622 ( .A0(n347), .A1(n463), .A2(n346), .Z(n332));
Q_AN03 U623 ( .A0(n347), .A1(n464), .A2(n346), .Z(n333));
Q_AN03 U624 ( .A0(n347), .A1(n465), .A2(n346), .Z(n334));
Q_AN03 U625 ( .A0(n347), .A1(n466), .A2(n346), .Z(n335));
Q_AN03 U626 ( .A0(n347), .A1(n467), .A2(n346), .Z(n336));
Q_AN03 U627 ( .A0(n347), .A1(n468), .A2(n346), .Z(n337));
Q_AN03 U628 ( .A0(n347), .A1(n469), .A2(n346), .Z(n338));
Q_AN03 U629 ( .A0(n347), .A1(n470), .A2(n346), .Z(n339));
Q_AN03 U630 ( .A0(n347), .A1(n471), .A2(n346), .Z(n340));
Q_AN03 U631 ( .A0(n347), .A1(n472), .A2(n346), .Z(n341));
Q_AN03 U632 ( .A0(n347), .A1(n473), .A2(n346), .Z(n342));
Q_AN03 U633 ( .A0(n347), .A1(n474), .A2(n346), .Z(n343));
Q_AN03 U634 ( .A0(n347), .A1(n475), .A2(n346), .Z(n344));
Q_AN03 U635 ( .A0(n347), .A1(n476), .A2(n346), .Z(n345));
Q_INV U636 ( .A(n882), .Z(n347));
Q_MX03 U637 ( .S0(n883), .S1(n882), .A0(n558), .A1(n526), .A2(n412), .Z(n348));
Q_MX03 U638 ( .S0(n883), .S1(n882), .A0(n559), .A1(n527), .A2(n413), .Z(n349));
Q_MX03 U639 ( .S0(n883), .S1(n882), .A0(n560), .A1(n528), .A2(n414), .Z(n350));
Q_MX03 U640 ( .S0(n883), .S1(n882), .A0(n561), .A1(n529), .A2(n415), .Z(n351));
Q_MX03 U641 ( .S0(n883), .S1(n882), .A0(n562), .A1(n530), .A2(n416), .Z(n352));
Q_MX03 U642 ( .S0(n883), .S1(n882), .A0(n563), .A1(n531), .A2(n417), .Z(n353));
Q_MX03 U643 ( .S0(n883), .S1(n882), .A0(n564), .A1(n532), .A2(n418), .Z(n354));
Q_MX03 U644 ( .S0(n883), .S1(n882), .A0(n565), .A1(n533), .A2(n419), .Z(n355));
Q_MX03 U645 ( .S0(n883), .S1(n882), .A0(n566), .A1(n534), .A2(n420), .Z(n356));
Q_MX03 U646 ( .S0(n883), .S1(n882), .A0(n567), .A1(n535), .A2(n421), .Z(n357));
Q_MX03 U647 ( .S0(n883), .S1(n882), .A0(n568), .A1(n536), .A2(n422), .Z(n358));
Q_MX03 U648 ( .S0(n883), .S1(n882), .A0(n569), .A1(n537), .A2(n423), .Z(n359));
Q_MX03 U649 ( .S0(n883), .S1(n882), .A0(n570), .A1(n538), .A2(n424), .Z(n360));
Q_MX03 U650 ( .S0(n883), .S1(n882), .A0(n571), .A1(n539), .A2(n425), .Z(n361));
Q_MX03 U651 ( .S0(n883), .S1(n882), .A0(n572), .A1(n540), .A2(n426), .Z(n362));
Q_MX03 U652 ( .S0(n883), .S1(n882), .A0(n573), .A1(n541), .A2(n427), .Z(n363));
Q_MX03 U653 ( .S0(n883), .S1(n882), .A0(n574), .A1(n542), .A2(n428), .Z(n364));
Q_MX03 U654 ( .S0(n883), .S1(n882), .A0(n575), .A1(n543), .A2(n429), .Z(n365));
Q_MX03 U655 ( .S0(n883), .S1(n882), .A0(n576), .A1(n544), .A2(n430), .Z(n366));
Q_MX03 U656 ( .S0(n883), .S1(n882), .A0(n577), .A1(n545), .A2(n431), .Z(n367));
Q_MX03 U657 ( .S0(n883), .S1(n882), .A0(n578), .A1(n546), .A2(n432), .Z(n368));
Q_MX03 U658 ( .S0(n883), .S1(n882), .A0(n579), .A1(n547), .A2(n433), .Z(n369));
Q_MX03 U659 ( .S0(n883), .S1(n882), .A0(n580), .A1(n548), .A2(n434), .Z(n370));
Q_MX03 U660 ( .S0(n883), .S1(n882), .A0(n581), .A1(n549), .A2(n435), .Z(n371));
Q_MX03 U661 ( .S0(n883), .S1(n882), .A0(n582), .A1(n550), .A2(n436), .Z(n372));
Q_MX03 U662 ( .S0(n883), .S1(n882), .A0(n583), .A1(n551), .A2(n437), .Z(n373));
Q_MX03 U663 ( .S0(n883), .S1(n882), .A0(n584), .A1(n552), .A2(n438), .Z(n374));
Q_MX03 U664 ( .S0(n883), .S1(n882), .A0(n585), .A1(n553), .A2(n439), .Z(n375));
Q_MX03 U665 ( .S0(n883), .S1(n882), .A0(n586), .A1(n554), .A2(n440), .Z(n376));
Q_MX03 U666 ( .S0(n883), .S1(n882), .A0(n587), .A1(n555), .A2(n441), .Z(n377));
Q_MX03 U667 ( .S0(n883), .S1(n882), .A0(n588), .A1(n556), .A2(n442), .Z(n378));
Q_MX03 U668 ( .S0(n883), .S1(n882), .A0(n589), .A1(n557), .A2(n443), .Z(n379));
Q_MX02 U669 ( .S(n882), .A0(n477), .A1(n445), .Z(n380));
Q_MX02 U670 ( .S(n882), .A0(n478), .A1(n446), .Z(n381));
Q_MX02 U671 ( .S(n882), .A0(n479), .A1(n447), .Z(n382));
Q_MX02 U672 ( .S(n882), .A0(n480), .A1(n448), .Z(n383));
Q_MX02 U673 ( .S(n882), .A0(n481), .A1(n449), .Z(n384));
Q_MX02 U674 ( .S(n882), .A0(n482), .A1(n450), .Z(n385));
Q_MX02 U675 ( .S(n882), .A0(n483), .A1(n451), .Z(n386));
Q_MX02 U676 ( .S(n882), .A0(n484), .A1(n452), .Z(n387));
Q_MX02 U677 ( .S(n882), .A0(n485), .A1(n453), .Z(n388));
Q_MX02 U678 ( .S(n882), .A0(n486), .A1(n454), .Z(n389));
Q_MX02 U679 ( .S(n882), .A0(n487), .A1(n455), .Z(n390));
Q_MX02 U680 ( .S(n882), .A0(n488), .A1(n456), .Z(n391));
Q_MX02 U681 ( .S(n882), .A0(n489), .A1(n457), .Z(n392));
Q_MX02 U682 ( .S(n882), .A0(n490), .A1(n458), .Z(n393));
Q_MX02 U683 ( .S(n882), .A0(n491), .A1(n459), .Z(n394));
Q_MX02 U684 ( .S(n882), .A0(n492), .A1(n460), .Z(n395));
Q_MX03 U685 ( .S0(n883), .S1(n882), .A0(n590), .A1(n574), .A2(n461), .Z(n396));
Q_MX03 U686 ( .S0(n883), .S1(n882), .A0(n591), .A1(n575), .A2(n462), .Z(n397));
Q_MX03 U687 ( .S0(n883), .S1(n882), .A0(n592), .A1(n576), .A2(n463), .Z(n398));
Q_MX03 U688 ( .S0(n883), .S1(n882), .A0(n593), .A1(n577), .A2(n464), .Z(n399));
Q_MX03 U689 ( .S0(n883), .S1(n882), .A0(n594), .A1(n578), .A2(n465), .Z(n400));
Q_MX03 U690 ( .S0(n883), .S1(n882), .A0(n595), .A1(n579), .A2(n466), .Z(n401));
Q_MX03 U691 ( .S0(n883), .S1(n882), .A0(n596), .A1(n580), .A2(n467), .Z(n402));
Q_MX03 U692 ( .S0(n883), .S1(n882), .A0(n597), .A1(n581), .A2(n468), .Z(n403));
Q_MX03 U693 ( .S0(n883), .S1(n882), .A0(n598), .A1(n582), .A2(n469), .Z(n404));
Q_MX03 U694 ( .S0(n883), .S1(n882), .A0(n599), .A1(n583), .A2(n470), .Z(n405));
Q_MX03 U695 ( .S0(n883), .S1(n882), .A0(n600), .A1(n584), .A2(n471), .Z(n406));
Q_MX03 U696 ( .S0(n883), .S1(n882), .A0(n601), .A1(n585), .A2(n472), .Z(n407));
Q_MX03 U697 ( .S0(n883), .S1(n882), .A0(n602), .A1(n586), .A2(n473), .Z(n408));
Q_MX03 U698 ( .S0(n883), .S1(n882), .A0(n603), .A1(n587), .A2(n474), .Z(n409));
Q_MX03 U699 ( .S0(n883), .S1(n882), .A0(n604), .A1(n588), .A2(n475), .Z(n410));
Q_MX03 U700 ( .S0(n883), .S1(n882), .A0(n605), .A1(n589), .A2(n476), .Z(n411));
Q_AN02 U701 ( .A0(n444), .A1(n493), .Z(n412));
Q_AN02 U702 ( .A0(n444), .A1(n494), .Z(n413));
Q_AN02 U703 ( .A0(n444), .A1(n495), .Z(n414));
Q_AN02 U704 ( .A0(n444), .A1(n496), .Z(n415));
Q_AN02 U705 ( .A0(n444), .A1(n497), .Z(n416));
Q_AN02 U706 ( .A0(n444), .A1(n498), .Z(n417));
Q_AN02 U707 ( .A0(n444), .A1(n499), .Z(n418));
Q_AN02 U708 ( .A0(n444), .A1(n500), .Z(n419));
Q_AN02 U709 ( .A0(n444), .A1(n501), .Z(n420));
Q_AN02 U710 ( .A0(n444), .A1(n502), .Z(n421));
Q_AN02 U711 ( .A0(n444), .A1(n503), .Z(n422));
Q_AN02 U712 ( .A0(n444), .A1(n504), .Z(n423));
Q_AN02 U713 ( .A0(n444), .A1(n505), .Z(n424));
Q_AN02 U714 ( .A0(n444), .A1(n506), .Z(n425));
Q_AN02 U715 ( .A0(n444), .A1(n507), .Z(n426));
Q_AN02 U716 ( .A0(n444), .A1(n508), .Z(n427));
Q_AN02 U717 ( .A0(n444), .A1(n510), .Z(n428));
Q_AN02 U718 ( .A0(n444), .A1(n511), .Z(n429));
Q_AN02 U719 ( .A0(n444), .A1(n512), .Z(n430));
Q_AN02 U720 ( .A0(n444), .A1(n513), .Z(n431));
Q_AN02 U721 ( .A0(n444), .A1(n514), .Z(n432));
Q_AN02 U722 ( .A0(n444), .A1(n515), .Z(n433));
Q_AN02 U723 ( .A0(n444), .A1(n516), .Z(n434));
Q_AN02 U724 ( .A0(n444), .A1(n517), .Z(n435));
Q_AN02 U725 ( .A0(n444), .A1(n518), .Z(n436));
Q_AN02 U726 ( .A0(n444), .A1(n519), .Z(n437));
Q_AN02 U727 ( .A0(n444), .A1(n520), .Z(n438));
Q_AN02 U728 ( .A0(n444), .A1(n521), .Z(n439));
Q_AN02 U729 ( .A0(n444), .A1(n522), .Z(n440));
Q_AN02 U730 ( .A0(n444), .A1(n523), .Z(n441));
Q_AN02 U731 ( .A0(n444), .A1(n524), .Z(n442));
Q_AN02 U732 ( .A0(n444), .A1(n525), .Z(n443));
Q_INV U733 ( .A(n883), .Z(n444));
Q_MX02 U734 ( .S(n883), .A0(n526), .A1(n493), .Z(n445));
Q_MX02 U735 ( .S(n883), .A0(n527), .A1(n494), .Z(n446));
Q_MX02 U736 ( .S(n883), .A0(n528), .A1(n495), .Z(n447));
Q_MX02 U737 ( .S(n883), .A0(n529), .A1(n496), .Z(n448));
Q_MX02 U738 ( .S(n883), .A0(n530), .A1(n497), .Z(n449));
Q_MX02 U739 ( .S(n883), .A0(n531), .A1(n498), .Z(n450));
Q_MX02 U740 ( .S(n883), .A0(n532), .A1(n499), .Z(n451));
Q_MX02 U741 ( .S(n883), .A0(n533), .A1(n500), .Z(n452));
Q_MX02 U742 ( .S(n883), .A0(n534), .A1(n501), .Z(n453));
Q_MX02 U743 ( .S(n883), .A0(n535), .A1(n502), .Z(n454));
Q_MX02 U744 ( .S(n883), .A0(n536), .A1(n503), .Z(n455));
Q_MX02 U745 ( .S(n883), .A0(n537), .A1(n504), .Z(n456));
Q_MX02 U746 ( .S(n883), .A0(n538), .A1(n505), .Z(n457));
Q_MX02 U747 ( .S(n883), .A0(n539), .A1(n506), .Z(n458));
Q_MX02 U748 ( .S(n883), .A0(n540), .A1(n507), .Z(n459));
Q_MX02 U749 ( .S(n883), .A0(n541), .A1(n508), .Z(n460));
Q_MX02 U750 ( .S(n883), .A0(n542), .A1(n510), .Z(n461));
Q_MX02 U751 ( .S(n883), .A0(n543), .A1(n511), .Z(n462));
Q_MX02 U752 ( .S(n883), .A0(n544), .A1(n512), .Z(n463));
Q_MX02 U753 ( .S(n883), .A0(n545), .A1(n513), .Z(n464));
Q_MX02 U754 ( .S(n883), .A0(n546), .A1(n514), .Z(n465));
Q_MX02 U755 ( .S(n883), .A0(n547), .A1(n515), .Z(n466));
Q_MX02 U756 ( .S(n883), .A0(n548), .A1(n516), .Z(n467));
Q_MX02 U757 ( .S(n883), .A0(n549), .A1(n517), .Z(n468));
Q_MX02 U758 ( .S(n883), .A0(n550), .A1(n518), .Z(n469));
Q_MX02 U759 ( .S(n883), .A0(n551), .A1(n519), .Z(n470));
Q_MX02 U760 ( .S(n883), .A0(n552), .A1(n520), .Z(n471));
Q_MX02 U761 ( .S(n883), .A0(n553), .A1(n521), .Z(n472));
Q_MX02 U762 ( .S(n883), .A0(n554), .A1(n522), .Z(n473));
Q_MX02 U763 ( .S(n883), .A0(n555), .A1(n523), .Z(n474));
Q_MX02 U764 ( .S(n883), .A0(n556), .A1(n524), .Z(n475));
Q_MX02 U765 ( .S(n883), .A0(n557), .A1(n525), .Z(n476));
Q_MX03 U766 ( .S0(n884), .S1(n883), .A0(n703), .A1(n687), .A2(n558), .Z(n477));
Q_MX03 U767 ( .S0(n884), .S1(n883), .A0(n704), .A1(n688), .A2(n559), .Z(n478));
Q_MX03 U768 ( .S0(n884), .S1(n883), .A0(n705), .A1(n689), .A2(n560), .Z(n479));
Q_MX03 U769 ( .S0(n884), .S1(n883), .A0(n706), .A1(n690), .A2(n561), .Z(n480));
Q_MX03 U770 ( .S0(n884), .S1(n883), .A0(n707), .A1(n691), .A2(n562), .Z(n481));
Q_MX03 U771 ( .S0(n884), .S1(n883), .A0(n708), .A1(n692), .A2(n563), .Z(n482));
Q_MX03 U772 ( .S0(n884), .S1(n883), .A0(n709), .A1(n693), .A2(n564), .Z(n483));
Q_MX03 U773 ( .S0(n884), .S1(n883), .A0(n710), .A1(n694), .A2(n565), .Z(n484));
Q_MX03 U774 ( .S0(n884), .S1(n883), .A0(n711), .A1(n695), .A2(n566), .Z(n485));
Q_MX03 U775 ( .S0(n884), .S1(n883), .A0(n712), .A1(n696), .A2(n567), .Z(n486));
Q_MX03 U776 ( .S0(n884), .S1(n883), .A0(n713), .A1(n697), .A2(n568), .Z(n487));
Q_MX03 U777 ( .S0(n884), .S1(n883), .A0(n714), .A1(n698), .A2(n569), .Z(n488));
Q_MX03 U778 ( .S0(n884), .S1(n883), .A0(n715), .A1(n699), .A2(n570), .Z(n489));
Q_MX03 U779 ( .S0(n884), .S1(n883), .A0(n716), .A1(n700), .A2(n571), .Z(n490));
Q_MX03 U780 ( .S0(n884), .S1(n883), .A0(n717), .A1(n701), .A2(n572), .Z(n491));
Q_MX03 U781 ( .S0(n884), .S1(n883), .A0(n718), .A1(n702), .A2(n573), .Z(n492));
Q_AN02 U782 ( .A0(n509), .A1(n606), .Z(n493));
Q_AN02 U783 ( .A0(n509), .A1(n607), .Z(n494));
Q_AN02 U784 ( .A0(n509), .A1(n608), .Z(n495));
Q_AN02 U785 ( .A0(n509), .A1(n609), .Z(n496));
Q_AN02 U786 ( .A0(n509), .A1(n610), .Z(n497));
Q_AN02 U787 ( .A0(n509), .A1(n611), .Z(n498));
Q_AN02 U788 ( .A0(n509), .A1(n612), .Z(n499));
Q_AN02 U789 ( .A0(n509), .A1(n613), .Z(n500));
Q_AN02 U790 ( .A0(n509), .A1(n615), .Z(n501));
Q_AN02 U791 ( .A0(n509), .A1(n616), .Z(n502));
Q_AN02 U792 ( .A0(n509), .A1(n617), .Z(n503));
Q_AN02 U793 ( .A0(n509), .A1(n618), .Z(n504));
Q_AN02 U794 ( .A0(n509), .A1(n619), .Z(n505));
Q_AN02 U795 ( .A0(n509), .A1(n620), .Z(n506));
Q_AN02 U796 ( .A0(n509), .A1(n621), .Z(n507));
Q_AN02 U797 ( .A0(n509), .A1(n622), .Z(n508));
Q_INV U798 ( .A(n884), .Z(n509));
Q_MX02 U799 ( .S(n884), .A0(n623), .A1(n606), .Z(n510));
Q_MX02 U800 ( .S(n884), .A0(n624), .A1(n607), .Z(n511));
Q_MX02 U801 ( .S(n884), .A0(n625), .A1(n608), .Z(n512));
Q_MX02 U802 ( .S(n884), .A0(n626), .A1(n609), .Z(n513));
Q_MX02 U803 ( .S(n884), .A0(n627), .A1(n610), .Z(n514));
Q_MX02 U804 ( .S(n884), .A0(n628), .A1(n611), .Z(n515));
Q_MX02 U805 ( .S(n884), .A0(n629), .A1(n612), .Z(n516));
Q_MX02 U806 ( .S(n884), .A0(n630), .A1(n613), .Z(n517));
Q_MX02 U807 ( .S(n884), .A0(n631), .A1(n615), .Z(n518));
Q_MX02 U808 ( .S(n884), .A0(n632), .A1(n616), .Z(n519));
Q_MX02 U809 ( .S(n884), .A0(n633), .A1(n617), .Z(n520));
Q_MX02 U810 ( .S(n884), .A0(n634), .A1(n618), .Z(n521));
Q_MX02 U811 ( .S(n884), .A0(n635), .A1(n619), .Z(n522));
Q_MX02 U812 ( .S(n884), .A0(n636), .A1(n620), .Z(n523));
Q_MX02 U813 ( .S(n884), .A0(n637), .A1(n621), .Z(n524));
Q_MX02 U814 ( .S(n884), .A0(n638), .A1(n622), .Z(n525));
Q_MX02 U815 ( .S(n884), .A0(n639), .A1(n623), .Z(n526));
Q_MX02 U816 ( .S(n884), .A0(n640), .A1(n624), .Z(n527));
Q_MX02 U817 ( .S(n884), .A0(n641), .A1(n625), .Z(n528));
Q_MX02 U818 ( .S(n884), .A0(n642), .A1(n626), .Z(n529));
Q_MX02 U819 ( .S(n884), .A0(n643), .A1(n627), .Z(n530));
Q_MX02 U820 ( .S(n884), .A0(n644), .A1(n628), .Z(n531));
Q_MX02 U821 ( .S(n884), .A0(n645), .A1(n629), .Z(n532));
Q_MX02 U822 ( .S(n884), .A0(n646), .A1(n630), .Z(n533));
Q_MX02 U823 ( .S(n884), .A0(n647), .A1(n631), .Z(n534));
Q_MX02 U824 ( .S(n884), .A0(n648), .A1(n632), .Z(n535));
Q_MX02 U825 ( .S(n884), .A0(n649), .A1(n633), .Z(n536));
Q_MX02 U826 ( .S(n884), .A0(n650), .A1(n634), .Z(n537));
Q_MX02 U827 ( .S(n884), .A0(n651), .A1(n635), .Z(n538));
Q_MX02 U828 ( .S(n884), .A0(n652), .A1(n636), .Z(n539));
Q_MX02 U829 ( .S(n884), .A0(n653), .A1(n637), .Z(n540));
Q_MX02 U830 ( .S(n884), .A0(n654), .A1(n638), .Z(n541));
Q_MX02 U831 ( .S(n884), .A0(n655), .A1(n639), .Z(n542));
Q_MX02 U832 ( .S(n884), .A0(n656), .A1(n640), .Z(n543));
Q_MX02 U833 ( .S(n884), .A0(n657), .A1(n641), .Z(n544));
Q_MX02 U834 ( .S(n884), .A0(n658), .A1(n642), .Z(n545));
Q_MX02 U835 ( .S(n884), .A0(n659), .A1(n643), .Z(n546));
Q_MX02 U836 ( .S(n884), .A0(n660), .A1(n644), .Z(n547));
Q_MX02 U837 ( .S(n884), .A0(n661), .A1(n645), .Z(n548));
Q_MX02 U838 ( .S(n884), .A0(n662), .A1(n646), .Z(n549));
Q_MX02 U839 ( .S(n884), .A0(n663), .A1(n647), .Z(n550));
Q_MX02 U840 ( .S(n884), .A0(n664), .A1(n648), .Z(n551));
Q_MX02 U841 ( .S(n884), .A0(n665), .A1(n649), .Z(n552));
Q_MX02 U842 ( .S(n884), .A0(n666), .A1(n650), .Z(n553));
Q_MX02 U843 ( .S(n884), .A0(n667), .A1(n651), .Z(n554));
Q_MX02 U844 ( .S(n884), .A0(n668), .A1(n652), .Z(n555));
Q_MX02 U845 ( .S(n884), .A0(n669), .A1(n653), .Z(n556));
Q_MX02 U846 ( .S(n884), .A0(n670), .A1(n654), .Z(n557));
Q_MX02 U847 ( .S(n884), .A0(n671), .A1(n655), .Z(n558));
Q_MX02 U848 ( .S(n884), .A0(n672), .A1(n656), .Z(n559));
Q_MX02 U849 ( .S(n884), .A0(n673), .A1(n657), .Z(n560));
Q_MX02 U850 ( .S(n884), .A0(n674), .A1(n658), .Z(n561));
Q_MX02 U851 ( .S(n884), .A0(n675), .A1(n659), .Z(n562));
Q_MX02 U852 ( .S(n884), .A0(n676), .A1(n660), .Z(n563));
Q_MX02 U853 ( .S(n884), .A0(n677), .A1(n661), .Z(n564));
Q_MX02 U854 ( .S(n884), .A0(n678), .A1(n662), .Z(n565));
Q_MX02 U855 ( .S(n884), .A0(n679), .A1(n663), .Z(n566));
Q_MX02 U856 ( .S(n884), .A0(n680), .A1(n664), .Z(n567));
Q_MX02 U857 ( .S(n884), .A0(n681), .A1(n665), .Z(n568));
Q_MX02 U858 ( .S(n884), .A0(n682), .A1(n666), .Z(n569));
Q_MX02 U859 ( .S(n884), .A0(n683), .A1(n667), .Z(n570));
Q_MX02 U860 ( .S(n884), .A0(n684), .A1(n668), .Z(n571));
Q_MX02 U861 ( .S(n884), .A0(n685), .A1(n669), .Z(n572));
Q_MX02 U862 ( .S(n884), .A0(n686), .A1(n670), .Z(n573));
Q_MX02 U863 ( .S(n884), .A0(n687), .A1(n671), .Z(n574));
Q_MX02 U864 ( .S(n884), .A0(n688), .A1(n672), .Z(n575));
Q_MX02 U865 ( .S(n884), .A0(n689), .A1(n673), .Z(n576));
Q_MX02 U866 ( .S(n884), .A0(n690), .A1(n674), .Z(n577));
Q_MX02 U867 ( .S(n884), .A0(n691), .A1(n675), .Z(n578));
Q_MX02 U868 ( .S(n884), .A0(n692), .A1(n676), .Z(n579));
Q_MX02 U869 ( .S(n884), .A0(n693), .A1(n677), .Z(n580));
Q_MX02 U870 ( .S(n884), .A0(n694), .A1(n678), .Z(n581));
Q_MX02 U871 ( .S(n884), .A0(n695), .A1(n679), .Z(n582));
Q_MX02 U872 ( .S(n884), .A0(n696), .A1(n680), .Z(n583));
Q_MX02 U873 ( .S(n884), .A0(n697), .A1(n681), .Z(n584));
Q_MX02 U874 ( .S(n884), .A0(n698), .A1(n682), .Z(n585));
Q_MX02 U875 ( .S(n884), .A0(n699), .A1(n683), .Z(n586));
Q_MX02 U876 ( .S(n884), .A0(n700), .A1(n684), .Z(n587));
Q_MX02 U877 ( .S(n884), .A0(n701), .A1(n685), .Z(n588));
Q_MX02 U878 ( .S(n884), .A0(n702), .A1(n686), .Z(n589));
Q_MX03 U879 ( .S0(n885), .S1(n884), .A0(n831), .A1(n823), .A2(n703), .Z(n590));
Q_MX03 U880 ( .S0(n885), .S1(n884), .A0(n832), .A1(n824), .A2(n704), .Z(n591));
Q_MX03 U881 ( .S0(n885), .S1(n884), .A0(n833), .A1(n825), .A2(n705), .Z(n592));
Q_MX03 U882 ( .S0(n885), .S1(n884), .A0(n834), .A1(n826), .A2(n706), .Z(n593));
Q_MX03 U883 ( .S0(n885), .S1(n884), .A0(n835), .A1(n827), .A2(n707), .Z(n594));
Q_MX03 U884 ( .S0(n885), .S1(n884), .A0(n836), .A1(n828), .A2(n708), .Z(n595));
Q_MX03 U885 ( .S0(n885), .S1(n884), .A0(n837), .A1(n829), .A2(n709), .Z(n596));
Q_MX03 U886 ( .S0(n885), .S1(n884), .A0(n838), .A1(n830), .A2(n710), .Z(n597));
Q_MX03 U887 ( .S0(n885), .S1(n884), .A0(n839), .A1(n831), .A2(n711), .Z(n598));
Q_MX03 U888 ( .S0(n885), .S1(n884), .A0(n840), .A1(n832), .A2(n712), .Z(n599));
Q_MX03 U889 ( .S0(n885), .S1(n884), .A0(n841), .A1(n833), .A2(n713), .Z(n600));
Q_MX03 U890 ( .S0(n885), .S1(n884), .A0(n842), .A1(n834), .A2(n714), .Z(n601));
Q_MX03 U891 ( .S0(n885), .S1(n884), .A0(n843), .A1(n835), .A2(n715), .Z(n602));
Q_MX03 U892 ( .S0(n885), .S1(n884), .A0(n844), .A1(n836), .A2(n716), .Z(n603));
Q_MX03 U893 ( .S0(n885), .S1(n884), .A0(n845), .A1(n837), .A2(n717), .Z(n604));
Q_MX03 U894 ( .S0(n885), .S1(n884), .A0(n846), .A1(n838), .A2(n718), .Z(n605));
Q_AN02 U895 ( .A0(n614), .A1(n719), .Z(n606));
Q_AN02 U896 ( .A0(n614), .A1(n720), .Z(n607));
Q_AN02 U897 ( .A0(n614), .A1(n721), .Z(n608));
Q_AN02 U898 ( .A0(n614), .A1(n722), .Z(n609));
Q_AN02 U899 ( .A0(n614), .A1(n723), .Z(n610));
Q_AN02 U900 ( .A0(n614), .A1(n724), .Z(n611));
Q_AN02 U901 ( .A0(n614), .A1(n725), .Z(n612));
Q_AN02 U902 ( .A0(n614), .A1(n726), .Z(n613));
Q_INV U903 ( .A(n885), .Z(n614));
Q_MX02 U904 ( .S(n885), .A0(n727), .A1(n719), .Z(n615));
Q_MX02 U905 ( .S(n885), .A0(n728), .A1(n720), .Z(n616));
Q_MX02 U906 ( .S(n885), .A0(n729), .A1(n721), .Z(n617));
Q_MX02 U907 ( .S(n885), .A0(n730), .A1(n722), .Z(n618));
Q_MX02 U908 ( .S(n885), .A0(n731), .A1(n723), .Z(n619));
Q_MX02 U909 ( .S(n885), .A0(n732), .A1(n724), .Z(n620));
Q_MX02 U910 ( .S(n885), .A0(n733), .A1(n725), .Z(n621));
Q_MX02 U911 ( .S(n885), .A0(n734), .A1(n726), .Z(n622));
Q_MX02 U912 ( .S(n885), .A0(n735), .A1(n727), .Z(n623));
Q_MX02 U913 ( .S(n885), .A0(n736), .A1(n728), .Z(n624));
Q_MX02 U914 ( .S(n885), .A0(n737), .A1(n729), .Z(n625));
Q_MX02 U915 ( .S(n885), .A0(n738), .A1(n730), .Z(n626));
Q_MX02 U916 ( .S(n885), .A0(n739), .A1(n731), .Z(n627));
Q_MX02 U917 ( .S(n885), .A0(n740), .A1(n732), .Z(n628));
Q_MX02 U918 ( .S(n885), .A0(n741), .A1(n733), .Z(n629));
Q_MX02 U919 ( .S(n885), .A0(n742), .A1(n734), .Z(n630));
Q_MX02 U920 ( .S(n885), .A0(n743), .A1(n735), .Z(n631));
Q_MX02 U921 ( .S(n885), .A0(n744), .A1(n736), .Z(n632));
Q_MX02 U922 ( .S(n885), .A0(n745), .A1(n737), .Z(n633));
Q_MX02 U923 ( .S(n885), .A0(n746), .A1(n738), .Z(n634));
Q_MX02 U924 ( .S(n885), .A0(n747), .A1(n739), .Z(n635));
Q_MX02 U925 ( .S(n885), .A0(n748), .A1(n740), .Z(n636));
Q_MX02 U926 ( .S(n885), .A0(n749), .A1(n741), .Z(n637));
Q_MX02 U927 ( .S(n885), .A0(n750), .A1(n742), .Z(n638));
Q_MX02 U928 ( .S(n885), .A0(n751), .A1(n743), .Z(n639));
Q_MX02 U929 ( .S(n885), .A0(n752), .A1(n744), .Z(n640));
Q_MX02 U930 ( .S(n885), .A0(n753), .A1(n745), .Z(n641));
Q_MX02 U931 ( .S(n885), .A0(n754), .A1(n746), .Z(n642));
Q_MX02 U932 ( .S(n885), .A0(n755), .A1(n747), .Z(n643));
Q_MX02 U933 ( .S(n885), .A0(n756), .A1(n748), .Z(n644));
Q_MX02 U934 ( .S(n885), .A0(n757), .A1(n749), .Z(n645));
Q_MX02 U935 ( .S(n885), .A0(n758), .A1(n750), .Z(n646));
Q_MX02 U936 ( .S(n885), .A0(n759), .A1(n751), .Z(n647));
Q_MX02 U937 ( .S(n885), .A0(n760), .A1(n752), .Z(n648));
Q_MX02 U938 ( .S(n885), .A0(n761), .A1(n753), .Z(n649));
Q_MX02 U939 ( .S(n885), .A0(n762), .A1(n754), .Z(n650));
Q_MX02 U940 ( .S(n885), .A0(n763), .A1(n755), .Z(n651));
Q_MX02 U941 ( .S(n885), .A0(n764), .A1(n756), .Z(n652));
Q_MX02 U942 ( .S(n885), .A0(n765), .A1(n757), .Z(n653));
Q_MX02 U943 ( .S(n885), .A0(n766), .A1(n758), .Z(n654));
Q_MX02 U944 ( .S(n885), .A0(n767), .A1(n759), .Z(n655));
Q_MX02 U945 ( .S(n885), .A0(n768), .A1(n760), .Z(n656));
Q_MX02 U946 ( .S(n885), .A0(n769), .A1(n761), .Z(n657));
Q_MX02 U947 ( .S(n885), .A0(n770), .A1(n762), .Z(n658));
Q_MX02 U948 ( .S(n885), .A0(n771), .A1(n763), .Z(n659));
Q_MX02 U949 ( .S(n885), .A0(n772), .A1(n764), .Z(n660));
Q_MX02 U950 ( .S(n885), .A0(n773), .A1(n765), .Z(n661));
Q_MX02 U951 ( .S(n885), .A0(n774), .A1(n766), .Z(n662));
Q_MX02 U952 ( .S(n885), .A0(n775), .A1(n767), .Z(n663));
Q_MX02 U953 ( .S(n885), .A0(n776), .A1(n768), .Z(n664));
Q_MX02 U954 ( .S(n885), .A0(n777), .A1(n769), .Z(n665));
Q_MX02 U955 ( .S(n885), .A0(n778), .A1(n770), .Z(n666));
Q_MX02 U956 ( .S(n885), .A0(n779), .A1(n771), .Z(n667));
Q_MX02 U957 ( .S(n885), .A0(n780), .A1(n772), .Z(n668));
Q_MX02 U958 ( .S(n885), .A0(n781), .A1(n773), .Z(n669));
Q_MX02 U959 ( .S(n885), .A0(n782), .A1(n774), .Z(n670));
Q_MX02 U960 ( .S(n885), .A0(n783), .A1(n775), .Z(n671));
Q_MX02 U961 ( .S(n885), .A0(n784), .A1(n776), .Z(n672));
Q_MX02 U962 ( .S(n885), .A0(n785), .A1(n777), .Z(n673));
Q_MX02 U963 ( .S(n885), .A0(n786), .A1(n778), .Z(n674));
Q_MX02 U964 ( .S(n885), .A0(n787), .A1(n779), .Z(n675));
Q_MX02 U965 ( .S(n885), .A0(n788), .A1(n780), .Z(n676));
Q_MX02 U966 ( .S(n885), .A0(n789), .A1(n781), .Z(n677));
Q_MX02 U967 ( .S(n885), .A0(n790), .A1(n782), .Z(n678));
Q_MX02 U968 ( .S(n885), .A0(n791), .A1(n783), .Z(n679));
Q_MX02 U969 ( .S(n885), .A0(n792), .A1(n784), .Z(n680));
Q_MX02 U970 ( .S(n885), .A0(n793), .A1(n785), .Z(n681));
Q_MX02 U971 ( .S(n885), .A0(n794), .A1(n786), .Z(n682));
Q_MX02 U972 ( .S(n885), .A0(n795), .A1(n787), .Z(n683));
Q_MX02 U973 ( .S(n885), .A0(n796), .A1(n788), .Z(n684));
Q_MX02 U974 ( .S(n885), .A0(n797), .A1(n789), .Z(n685));
Q_MX02 U975 ( .S(n885), .A0(n798), .A1(n790), .Z(n686));
Q_MX02 U976 ( .S(n885), .A0(n799), .A1(n791), .Z(n687));
Q_MX02 U977 ( .S(n885), .A0(n800), .A1(n792), .Z(n688));
Q_MX02 U978 ( .S(n885), .A0(n801), .A1(n793), .Z(n689));
Q_MX02 U979 ( .S(n885), .A0(n802), .A1(n794), .Z(n690));
Q_MX02 U980 ( .S(n885), .A0(n803), .A1(n795), .Z(n691));
Q_MX02 U981 ( .S(n885), .A0(n804), .A1(n796), .Z(n692));
Q_MX02 U982 ( .S(n885), .A0(n805), .A1(n797), .Z(n693));
Q_MX02 U983 ( .S(n885), .A0(n806), .A1(n798), .Z(n694));
Q_MX02 U984 ( .S(n885), .A0(n807), .A1(n799), .Z(n695));
Q_MX02 U985 ( .S(n885), .A0(n808), .A1(n800), .Z(n696));
Q_MX02 U986 ( .S(n885), .A0(n809), .A1(n801), .Z(n697));
Q_MX02 U987 ( .S(n885), .A0(n810), .A1(n802), .Z(n698));
Q_MX02 U988 ( .S(n885), .A0(n811), .A1(n803), .Z(n699));
Q_MX02 U989 ( .S(n885), .A0(n812), .A1(n804), .Z(n700));
Q_MX02 U990 ( .S(n885), .A0(n813), .A1(n805), .Z(n701));
Q_MX02 U991 ( .S(n885), .A0(n814), .A1(n806), .Z(n702));
Q_MX02 U992 ( .S(n885), .A0(n815), .A1(n807), .Z(n703));
Q_MX02 U993 ( .S(n885), .A0(n816), .A1(n808), .Z(n704));
Q_MX02 U994 ( .S(n885), .A0(n817), .A1(n809), .Z(n705));
Q_MX02 U995 ( .S(n885), .A0(n818), .A1(n810), .Z(n706));
Q_MX02 U996 ( .S(n885), .A0(n819), .A1(n811), .Z(n707));
Q_MX02 U997 ( .S(n885), .A0(n820), .A1(n812), .Z(n708));
Q_MX02 U998 ( .S(n885), .A0(n821), .A1(n813), .Z(n709));
Q_MX02 U999 ( .S(n885), .A0(n822), .A1(n814), .Z(n710));
Q_MX02 U1000 ( .S(n885), .A0(n823), .A1(n815), .Z(n711));
Q_MX02 U1001 ( .S(n885), .A0(n824), .A1(n816), .Z(n712));
Q_MX02 U1002 ( .S(n885), .A0(n825), .A1(n817), .Z(n713));
Q_MX02 U1003 ( .S(n885), .A0(n826), .A1(n818), .Z(n714));
Q_MX02 U1004 ( .S(n885), .A0(n827), .A1(n819), .Z(n715));
Q_MX02 U1005 ( .S(n885), .A0(n828), .A1(n820), .Z(n716));
Q_MX02 U1006 ( .S(n885), .A0(n829), .A1(n821), .Z(n717));
Q_MX02 U1007 ( .S(n885), .A0(n830), .A1(n822), .Z(n718));
Q_AN02 U1008 ( .A0(\pipe_array_data[1][127] ), .A1(n853), .Z(n719));
Q_AN02 U1009 ( .A0(\pipe_array_data[1][126] ), .A1(n853), .Z(n720));
Q_AN02 U1010 ( .A0(\pipe_array_data[1][125] ), .A1(n853), .Z(n721));
Q_AN02 U1011 ( .A0(\pipe_array_data[1][124] ), .A1(n853), .Z(n722));
Q_AN02 U1012 ( .A0(\pipe_array_data[1][123] ), .A1(n853), .Z(n723));
Q_AN02 U1013 ( .A0(\pipe_array_data[1][122] ), .A1(n853), .Z(n724));
Q_AN02 U1014 ( .A0(\pipe_array_data[1][121] ), .A1(n853), .Z(n725));
Q_AN02 U1015 ( .A0(\pipe_array_data[1][120] ), .A1(n853), .Z(n726));
Q_AN02 U1016 ( .A0(\pipe_array_data[1][119] ), .A1(n854), .Z(n727));
Q_AN02 U1017 ( .A0(\pipe_array_data[1][118] ), .A1(n854), .Z(n728));
Q_AN02 U1018 ( .A0(\pipe_array_data[1][117] ), .A1(n854), .Z(n729));
Q_AN02 U1019 ( .A0(\pipe_array_data[1][116] ), .A1(n854), .Z(n730));
Q_AN02 U1020 ( .A0(\pipe_array_data[1][115] ), .A1(n854), .Z(n731));
Q_AN02 U1021 ( .A0(\pipe_array_data[1][114] ), .A1(n854), .Z(n732));
Q_AN02 U1022 ( .A0(\pipe_array_data[1][113] ), .A1(n854), .Z(n733));
Q_AN02 U1023 ( .A0(\pipe_array_data[1][112] ), .A1(n854), .Z(n734));
Q_AN02 U1024 ( .A0(\pipe_array_data[1][111] ), .A1(n855), .Z(n735));
Q_AN02 U1025 ( .A0(\pipe_array_data[1][110] ), .A1(n855), .Z(n736));
Q_AN02 U1026 ( .A0(\pipe_array_data[1][109] ), .A1(n855), .Z(n737));
Q_AN02 U1027 ( .A0(\pipe_array_data[1][108] ), .A1(n855), .Z(n738));
Q_AN02 U1028 ( .A0(\pipe_array_data[1][107] ), .A1(n855), .Z(n739));
Q_AN02 U1029 ( .A0(\pipe_array_data[1][106] ), .A1(n855), .Z(n740));
Q_AN02 U1030 ( .A0(\pipe_array_data[1][105] ), .A1(n855), .Z(n741));
Q_AN02 U1031 ( .A0(\pipe_array_data[1][104] ), .A1(n855), .Z(n742));
Q_AN02 U1032 ( .A0(\pipe_array_data[1][103] ), .A1(n856), .Z(n743));
Q_AN02 U1033 ( .A0(\pipe_array_data[1][102] ), .A1(n856), .Z(n744));
Q_AN02 U1034 ( .A0(\pipe_array_data[1][101] ), .A1(n856), .Z(n745));
Q_AN02 U1035 ( .A0(\pipe_array_data[1][100] ), .A1(n856), .Z(n746));
Q_AN02 U1036 ( .A0(\pipe_array_data[1][99] ), .A1(n856), .Z(n747));
Q_AN02 U1037 ( .A0(\pipe_array_data[1][98] ), .A1(n856), .Z(n748));
Q_AN02 U1038 ( .A0(\pipe_array_data[1][97] ), .A1(n856), .Z(n749));
Q_AN02 U1039 ( .A0(\pipe_array_data[1][96] ), .A1(n856), .Z(n750));
Q_AN02 U1040 ( .A0(\pipe_array_data[1][95] ), .A1(n857), .Z(n751));
Q_AN02 U1041 ( .A0(\pipe_array_data[1][94] ), .A1(n857), .Z(n752));
Q_AN02 U1042 ( .A0(\pipe_array_data[1][93] ), .A1(n857), .Z(n753));
Q_AN02 U1043 ( .A0(\pipe_array_data[1][92] ), .A1(n857), .Z(n754));
Q_AN02 U1044 ( .A0(\pipe_array_data[1][91] ), .A1(n857), .Z(n755));
Q_AN02 U1045 ( .A0(\pipe_array_data[1][90] ), .A1(n857), .Z(n756));
Q_AN02 U1046 ( .A0(\pipe_array_data[1][89] ), .A1(n857), .Z(n757));
Q_AN02 U1047 ( .A0(\pipe_array_data[1][88] ), .A1(n857), .Z(n758));
Q_AN02 U1048 ( .A0(\pipe_array_data[1][87] ), .A1(n858), .Z(n759));
Q_AN02 U1049 ( .A0(\pipe_array_data[1][86] ), .A1(n858), .Z(n760));
Q_AN02 U1050 ( .A0(\pipe_array_data[1][85] ), .A1(n858), .Z(n761));
Q_AN02 U1051 ( .A0(\pipe_array_data[1][84] ), .A1(n858), .Z(n762));
Q_AN02 U1052 ( .A0(\pipe_array_data[1][83] ), .A1(n858), .Z(n763));
Q_AN02 U1053 ( .A0(\pipe_array_data[1][82] ), .A1(n858), .Z(n764));
Q_AN02 U1054 ( .A0(\pipe_array_data[1][81] ), .A1(n858), .Z(n765));
Q_AN02 U1055 ( .A0(\pipe_array_data[1][80] ), .A1(n858), .Z(n766));
Q_AN02 U1056 ( .A0(\pipe_array_data[1][79] ), .A1(n859), .Z(n767));
Q_AN02 U1057 ( .A0(\pipe_array_data[1][78] ), .A1(n859), .Z(n768));
Q_AN02 U1058 ( .A0(\pipe_array_data[1][77] ), .A1(n859), .Z(n769));
Q_AN02 U1059 ( .A0(\pipe_array_data[1][76] ), .A1(n859), .Z(n770));
Q_AN02 U1060 ( .A0(\pipe_array_data[1][75] ), .A1(n859), .Z(n771));
Q_AN02 U1061 ( .A0(\pipe_array_data[1][74] ), .A1(n859), .Z(n772));
Q_AN02 U1062 ( .A0(\pipe_array_data[1][73] ), .A1(n859), .Z(n773));
Q_AN02 U1063 ( .A0(\pipe_array_data[1][72] ), .A1(n859), .Z(n774));
Q_AN02 U1064 ( .A0(\pipe_array_data[1][71] ), .A1(n860), .Z(n775));
Q_AN02 U1065 ( .A0(\pipe_array_data[1][70] ), .A1(n860), .Z(n776));
Q_AN02 U1066 ( .A0(\pipe_array_data[1][69] ), .A1(n860), .Z(n777));
Q_AN02 U1067 ( .A0(\pipe_array_data[1][68] ), .A1(n860), .Z(n778));
Q_AN02 U1068 ( .A0(\pipe_array_data[1][67] ), .A1(n860), .Z(n779));
Q_AN02 U1069 ( .A0(\pipe_array_data[1][66] ), .A1(n860), .Z(n780));
Q_AN02 U1070 ( .A0(\pipe_array_data[1][65] ), .A1(n860), .Z(n781));
Q_AN02 U1071 ( .A0(\pipe_array_data[1][64] ), .A1(n860), .Z(n782));
Q_AN02 U1072 ( .A0(\pipe_array_data[1][63] ), .A1(n847), .Z(n783));
Q_AN02 U1073 ( .A0(\pipe_array_data[1][62] ), .A1(n847), .Z(n784));
Q_AN02 U1074 ( .A0(\pipe_array_data[1][61] ), .A1(n847), .Z(n785));
Q_AN02 U1075 ( .A0(\pipe_array_data[1][60] ), .A1(n847), .Z(n786));
Q_AN02 U1076 ( .A0(\pipe_array_data[1][59] ), .A1(n847), .Z(n787));
Q_AN02 U1077 ( .A0(\pipe_array_data[1][58] ), .A1(n847), .Z(n788));
Q_AN02 U1078 ( .A0(\pipe_array_data[1][57] ), .A1(n847), .Z(n789));
Q_AN02 U1079 ( .A0(\pipe_array_data[1][56] ), .A1(n847), .Z(n790));
Q_AN02 U1080 ( .A0(\pipe_array_data[1][55] ), .A1(n848), .Z(n791));
Q_AN02 U1081 ( .A0(\pipe_array_data[1][54] ), .A1(n848), .Z(n792));
Q_AN02 U1082 ( .A0(\pipe_array_data[1][53] ), .A1(n848), .Z(n793));
Q_AN02 U1083 ( .A0(\pipe_array_data[1][52] ), .A1(n848), .Z(n794));
Q_AN02 U1084 ( .A0(\pipe_array_data[1][51] ), .A1(n848), .Z(n795));
Q_AN02 U1085 ( .A0(\pipe_array_data[1][50] ), .A1(n848), .Z(n796));
Q_AN02 U1086 ( .A0(\pipe_array_data[1][49] ), .A1(n848), .Z(n797));
Q_AN02 U1087 ( .A0(\pipe_array_data[1][48] ), .A1(n848), .Z(n798));
Q_AN02 U1088 ( .A0(\pipe_array_data[1][47] ), .A1(n849), .Z(n799));
Q_AN02 U1089 ( .A0(\pipe_array_data[1][46] ), .A1(n849), .Z(n800));
Q_AN02 U1090 ( .A0(\pipe_array_data[1][45] ), .A1(n849), .Z(n801));
Q_AN02 U1091 ( .A0(\pipe_array_data[1][44] ), .A1(n849), .Z(n802));
Q_AN02 U1092 ( .A0(\pipe_array_data[1][43] ), .A1(n849), .Z(n803));
Q_AN02 U1093 ( .A0(\pipe_array_data[1][42] ), .A1(n849), .Z(n804));
Q_AN02 U1094 ( .A0(\pipe_array_data[1][41] ), .A1(n849), .Z(n805));
Q_AN02 U1095 ( .A0(\pipe_array_data[1][40] ), .A1(n849), .Z(n806));
Q_AN02 U1096 ( .A0(\pipe_array_data[1][39] ), .A1(n864), .Z(n807));
Q_AN02 U1097 ( .A0(\pipe_array_data[1][38] ), .A1(n864), .Z(n808));
Q_AN02 U1098 ( .A0(\pipe_array_data[1][37] ), .A1(n864), .Z(n809));
Q_AN02 U1099 ( .A0(\pipe_array_data[1][36] ), .A1(n864), .Z(n810));
Q_AN02 U1100 ( .A0(\pipe_array_data[1][35] ), .A1(n864), .Z(n811));
Q_AN02 U1101 ( .A0(\pipe_array_data[1][34] ), .A1(n864), .Z(n812));
Q_AN02 U1102 ( .A0(\pipe_array_data[1][33] ), .A1(n864), .Z(n813));
Q_AN02 U1103 ( .A0(\pipe_array_data[1][32] ), .A1(n864), .Z(n814));
Q_AN02 U1104 ( .A0(\pipe_array_data[1][31] ), .A1(n850), .Z(n815));
Q_AN02 U1105 ( .A0(\pipe_array_data[1][30] ), .A1(n850), .Z(n816));
Q_AN02 U1106 ( .A0(\pipe_array_data[1][29] ), .A1(n850), .Z(n817));
Q_AN02 U1107 ( .A0(\pipe_array_data[1][28] ), .A1(n850), .Z(n818));
Q_AN02 U1108 ( .A0(\pipe_array_data[1][27] ), .A1(n850), .Z(n819));
Q_AN02 U1109 ( .A0(\pipe_array_data[1][26] ), .A1(n850), .Z(n820));
Q_AN02 U1110 ( .A0(\pipe_array_data[1][25] ), .A1(n850), .Z(n821));
Q_AN02 U1111 ( .A0(\pipe_array_data[1][24] ), .A1(n850), .Z(n822));
Q_AN02 U1112 ( .A0(\pipe_array_data[1][23] ), .A1(n851), .Z(n823));
Q_AN02 U1113 ( .A0(\pipe_array_data[1][22] ), .A1(n851), .Z(n824));
Q_AN02 U1114 ( .A0(\pipe_array_data[1][21] ), .A1(n851), .Z(n825));
Q_AN02 U1115 ( .A0(\pipe_array_data[1][20] ), .A1(n851), .Z(n826));
Q_AN02 U1116 ( .A0(\pipe_array_data[1][19] ), .A1(n851), .Z(n827));
Q_AN02 U1117 ( .A0(\pipe_array_data[1][18] ), .A1(n851), .Z(n828));
Q_AN02 U1118 ( .A0(\pipe_array_data[1][17] ), .A1(n851), .Z(n829));
Q_AN02 U1119 ( .A0(\pipe_array_data[1][16] ), .A1(n851), .Z(n830));
Q_AN02 U1120 ( .A0(\pipe_array_data[1][15] ), .A1(n852), .Z(n831));
Q_AN02 U1121 ( .A0(\pipe_array_data[1][14] ), .A1(n852), .Z(n832));
Q_AN02 U1122 ( .A0(\pipe_array_data[1][13] ), .A1(n852), .Z(n833));
Q_AN02 U1123 ( .A0(\pipe_array_data[1][12] ), .A1(n852), .Z(n834));
Q_AN02 U1124 ( .A0(\pipe_array_data[1][11] ), .A1(n852), .Z(n835));
Q_AN02 U1125 ( .A0(\pipe_array_data[1][10] ), .A1(n852), .Z(n836));
Q_AN02 U1126 ( .A0(\pipe_array_data[1][9] ), .A1(n852), .Z(n837));
Q_AN02 U1127 ( .A0(\pipe_array_data[1][8] ), .A1(n852), .Z(n838));
Q_AN02 U1128 ( .A0(\pipe_array_data[1][7] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n839));
Q_AN02 U1129 ( .A0(\pipe_array_data[1][6] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n840));
Q_AN02 U1130 ( .A0(\pipe_array_data[1][5] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n841));
Q_AN02 U1131 ( .A0(\pipe_array_data[1][4] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n842));
Q_AN02 U1132 ( .A0(\pipe_array_data[1][3] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n843));
Q_AN02 U1133 ( .A0(\pipe_array_data[1][2] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n844));
Q_AN02 U1134 ( .A0(\pipe_array_data[1][1] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n845));
Q_AN02 U1135 ( .A0(\pipe_array_data[1][0] ), .A1(\pipe_array_ack_num_bytes[1][4] ), .Z(n846));
Q_INV U1136 ( .A(n861), .Z(n847));
Q_INV U1137 ( .A(n862), .Z(n848));
Q_INV U1138 ( .A(n863), .Z(n849));
Q_INV U1139 ( .A(n865), .Z(n850));
Q_INV U1140 ( .A(n866), .Z(n851));
Q_INV U1141 ( .A(n867), .Z(n852));
Q_ND02 U1142 ( .A0(n868), .A1(n869), .Z(n856));
Q_OR02 U1143 ( .A0(\pipe_array_ack_num_bytes[1][4] ), .A1(\pipe_array_ack_num_bytes[1][3] ), .Z(n860));
Q_ND02 U1144 ( .A0(n868), .A1(n870), .Z(n864));
Q_INV U1145 ( .A(\pipe_array_ack_num_bytes[1][4] ), .Z(n868));
Q_ND03 U1146 ( .A0(n871), .A1(n872), .A2(n868), .Z(n853));
Q_ND03 U1147 ( .A0(n871), .A1(n873), .A2(n868), .Z(n854));
Q_ND03 U1148 ( .A0(n871), .A1(n874), .A2(n868), .Z(n855));
Q_NR02 U1149 ( .A0(\pipe_array_ack_num_bytes[1][3] ), .A1(\pipe_array_ack_num_bytes[1][2] ), .Z(n869));
Q_ND03 U1150 ( .A0(n871), .A1(n875), .A2(n868), .Z(n857));
Q_ND03 U1151 ( .A0(n871), .A1(n876), .A2(n868), .Z(n858));
Q_ND03 U1152 ( .A0(n871), .A1(n877), .A2(n868), .Z(n859));
Q_OA21 U1153 ( .A0(n871), .A1(n872), .B0(n868), .Z(n861));
Q_OA21 U1154 ( .A0(n871), .A1(n873), .B0(n868), .Z(n862));
Q_OA21 U1155 ( .A0(n871), .A1(n874), .B0(n868), .Z(n863));
Q_ND02 U1156 ( .A0(\pipe_array_ack_num_bytes[1][3] ), .A1(\pipe_array_ack_num_bytes[1][2] ), .Z(n870));
Q_OA21 U1157 ( .A0(n871), .A1(n875), .B0(n868), .Z(n865));
Q_OA21 U1158 ( .A0(n871), .A1(n876), .B0(n868), .Z(n866));
Q_OA21 U1159 ( .A0(n871), .A1(n877), .B0(n868), .Z(n867));
Q_INV U1160 ( .A(\pipe_array_ack_num_bytes[1][3] ), .Z(n871));
Q_AN02 U1161 ( .A0(n878), .A1(n879), .Z(n872));
Q_NR02 U1162 ( .A0(\pipe_array_ack_num_bytes[1][2] ), .A1(\pipe_array_ack_num_bytes[1][1] ), .Z(n873));
Q_AN02 U1163 ( .A0(n878), .A1(n880), .Z(n874));
Q_OR02 U1164 ( .A0(n878), .A1(n879), .Z(n875));
Q_ND02 U1165 ( .A0(\pipe_array_ack_num_bytes[1][2] ), .A1(\pipe_array_ack_num_bytes[1][1] ), .Z(n876));
Q_OR02 U1166 ( .A0(n878), .A1(n880), .Z(n877));
Q_INV U1167 ( .A(\pipe_array_ack_num_bytes[1][2] ), .Z(n878));
Q_NR02 U1168 ( .A0(\pipe_array_ack_num_bytes[1][1] ), .A1(\pipe_array_ack_num_bytes[1][0] ), .Z(n879));
Q_ND02 U1169 ( .A0(\pipe_array_ack_num_bytes[1][1] ), .A1(\pipe_array_ack_num_bytes[1][0] ), .Z(n880));
Q_AN02 U1170 ( .A0(\pipe_array_ack[0][0] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .Z(n881));
Q_AN02 U1171 ( .A0(\pipe_array_ack[0][0] ), .A1(\pipe_array_ack_num_bytes[0][3] ), .Z(n882));
Q_AN02 U1172 ( .A0(\pipe_array_ack[0][0] ), .A1(\pipe_array_ack_num_bytes[0][2] ), .Z(n883));
Q_AN02 U1173 ( .A0(\pipe_array_ack[0][0] ), .A1(\pipe_array_ack_num_bytes[0][1] ), .Z(n884));
Q_AN02 U1174 ( .A0(\pipe_array_ack[0][0] ), .A1(\pipe_array_ack_num_bytes[0][0] ), .Z(n885));
Q_AN03 U1175 ( .A0(\pipe_array_data[0][127] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n886));
Q_AN03 U1176 ( .A0(\pipe_array_data[0][126] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n887));
Q_AN03 U1177 ( .A0(\pipe_array_data[0][125] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n888));
Q_AN03 U1178 ( .A0(\pipe_array_data[0][124] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n889));
Q_AN03 U1179 ( .A0(\pipe_array_data[0][123] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n890));
Q_AN03 U1180 ( .A0(\pipe_array_data[0][122] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n891));
Q_AN03 U1181 ( .A0(\pipe_array_data[0][121] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n892));
Q_AN03 U1182 ( .A0(\pipe_array_data[0][120] ), .A1(n1020), .A2(\pipe_array_ack[0][0] ), .Z(n893));
Q_AN03 U1183 ( .A0(\pipe_array_data[0][119] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n894));
Q_AN03 U1184 ( .A0(\pipe_array_data[0][118] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n895));
Q_AN03 U1185 ( .A0(\pipe_array_data[0][117] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n896));
Q_AN03 U1186 ( .A0(\pipe_array_data[0][116] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n897));
Q_AN03 U1187 ( .A0(\pipe_array_data[0][115] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n898));
Q_AN03 U1188 ( .A0(\pipe_array_data[0][114] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n899));
Q_AN03 U1189 ( .A0(\pipe_array_data[0][113] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n900));
Q_AN03 U1190 ( .A0(\pipe_array_data[0][112] ), .A1(n1021), .A2(\pipe_array_ack[0][0] ), .Z(n901));
Q_AN03 U1191 ( .A0(\pipe_array_data[0][111] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n902));
Q_AN03 U1192 ( .A0(\pipe_array_data[0][110] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n903));
Q_AN03 U1193 ( .A0(\pipe_array_data[0][109] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n904));
Q_AN03 U1194 ( .A0(\pipe_array_data[0][108] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n905));
Q_AN03 U1195 ( .A0(\pipe_array_data[0][107] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n906));
Q_AN03 U1196 ( .A0(\pipe_array_data[0][106] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n907));
Q_AN03 U1197 ( .A0(\pipe_array_data[0][105] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n908));
Q_AN03 U1198 ( .A0(\pipe_array_data[0][104] ), .A1(n1022), .A2(\pipe_array_ack[0][0] ), .Z(n909));
Q_AN03 U1199 ( .A0(\pipe_array_data[0][103] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n910));
Q_AN03 U1200 ( .A0(\pipe_array_data[0][102] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n911));
Q_AN03 U1201 ( .A0(\pipe_array_data[0][101] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n912));
Q_AN03 U1202 ( .A0(\pipe_array_data[0][100] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n913));
Q_AN03 U1203 ( .A0(\pipe_array_data[0][99] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n914));
Q_AN03 U1204 ( .A0(\pipe_array_data[0][98] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n915));
Q_AN03 U1205 ( .A0(\pipe_array_data[0][97] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n916));
Q_AN03 U1206 ( .A0(\pipe_array_data[0][96] ), .A1(n1023), .A2(\pipe_array_ack[0][0] ), .Z(n917));
Q_AN03 U1207 ( .A0(\pipe_array_data[0][95] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n918));
Q_AN03 U1208 ( .A0(\pipe_array_data[0][94] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n919));
Q_AN03 U1209 ( .A0(\pipe_array_data[0][93] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n920));
Q_AN03 U1210 ( .A0(\pipe_array_data[0][92] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n921));
Q_AN03 U1211 ( .A0(\pipe_array_data[0][91] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n922));
Q_AN03 U1212 ( .A0(\pipe_array_data[0][90] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n923));
Q_AN03 U1213 ( .A0(\pipe_array_data[0][89] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n924));
Q_AN03 U1214 ( .A0(\pipe_array_data[0][88] ), .A1(n1024), .A2(\pipe_array_ack[0][0] ), .Z(n925));
Q_AN03 U1215 ( .A0(\pipe_array_data[0][87] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n926));
Q_AN03 U1216 ( .A0(\pipe_array_data[0][86] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n927));
Q_AN03 U1217 ( .A0(\pipe_array_data[0][85] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n928));
Q_AN03 U1218 ( .A0(\pipe_array_data[0][84] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n929));
Q_AN03 U1219 ( .A0(\pipe_array_data[0][83] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n930));
Q_AN03 U1220 ( .A0(\pipe_array_data[0][82] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n931));
Q_AN03 U1221 ( .A0(\pipe_array_data[0][81] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n932));
Q_AN03 U1222 ( .A0(\pipe_array_data[0][80] ), .A1(n1025), .A2(\pipe_array_ack[0][0] ), .Z(n933));
Q_AN03 U1223 ( .A0(\pipe_array_data[0][79] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n934));
Q_AN03 U1224 ( .A0(\pipe_array_data[0][78] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n935));
Q_AN03 U1225 ( .A0(\pipe_array_data[0][77] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n936));
Q_AN03 U1226 ( .A0(\pipe_array_data[0][76] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n937));
Q_AN03 U1227 ( .A0(\pipe_array_data[0][75] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n938));
Q_AN03 U1228 ( .A0(\pipe_array_data[0][74] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n939));
Q_AN03 U1229 ( .A0(\pipe_array_data[0][73] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n940));
Q_AN03 U1230 ( .A0(\pipe_array_data[0][72] ), .A1(n1026), .A2(\pipe_array_ack[0][0] ), .Z(n941));
Q_AN03 U1231 ( .A0(\pipe_array_data[0][71] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n942));
Q_AN03 U1232 ( .A0(\pipe_array_data[0][70] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n943));
Q_AN03 U1233 ( .A0(\pipe_array_data[0][69] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n944));
Q_AN03 U1234 ( .A0(\pipe_array_data[0][68] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n945));
Q_AN03 U1235 ( .A0(\pipe_array_data[0][67] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n946));
Q_AN03 U1236 ( .A0(\pipe_array_data[0][66] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n947));
Q_AN03 U1237 ( .A0(\pipe_array_data[0][65] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n948));
Q_AN03 U1238 ( .A0(\pipe_array_data[0][64] ), .A1(n1027), .A2(\pipe_array_ack[0][0] ), .Z(n949));
Q_AN03 U1239 ( .A0(\pipe_array_data[0][63] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n950));
Q_AN03 U1240 ( .A0(\pipe_array_data[0][62] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n951));
Q_AN03 U1241 ( .A0(\pipe_array_data[0][61] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n952));
Q_AN03 U1242 ( .A0(\pipe_array_data[0][60] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n953));
Q_AN03 U1243 ( .A0(\pipe_array_data[0][59] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n954));
Q_AN03 U1244 ( .A0(\pipe_array_data[0][58] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n955));
Q_AN03 U1245 ( .A0(\pipe_array_data[0][57] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n956));
Q_AN03 U1246 ( .A0(\pipe_array_data[0][56] ), .A1(n1014), .A2(\pipe_array_ack[0][0] ), .Z(n957));
Q_AN03 U1247 ( .A0(\pipe_array_data[0][55] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n958));
Q_AN03 U1248 ( .A0(\pipe_array_data[0][54] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n959));
Q_AN03 U1249 ( .A0(\pipe_array_data[0][53] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n960));
Q_AN03 U1250 ( .A0(\pipe_array_data[0][52] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n961));
Q_AN03 U1251 ( .A0(\pipe_array_data[0][51] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n962));
Q_AN03 U1252 ( .A0(\pipe_array_data[0][50] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n963));
Q_AN03 U1253 ( .A0(\pipe_array_data[0][49] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n964));
Q_AN03 U1254 ( .A0(\pipe_array_data[0][48] ), .A1(n1015), .A2(\pipe_array_ack[0][0] ), .Z(n965));
Q_AN03 U1255 ( .A0(\pipe_array_data[0][47] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n966));
Q_AN03 U1256 ( .A0(\pipe_array_data[0][46] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n967));
Q_AN03 U1257 ( .A0(\pipe_array_data[0][45] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n968));
Q_AN03 U1258 ( .A0(\pipe_array_data[0][44] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n969));
Q_AN03 U1259 ( .A0(\pipe_array_data[0][43] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n970));
Q_AN03 U1260 ( .A0(\pipe_array_data[0][42] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n971));
Q_AN03 U1261 ( .A0(\pipe_array_data[0][41] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n972));
Q_AN03 U1262 ( .A0(\pipe_array_data[0][40] ), .A1(n1016), .A2(\pipe_array_ack[0][0] ), .Z(n973));
Q_AN03 U1263 ( .A0(\pipe_array_data[0][39] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n974));
Q_AN03 U1264 ( .A0(\pipe_array_data[0][38] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n975));
Q_AN03 U1265 ( .A0(\pipe_array_data[0][37] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n976));
Q_AN03 U1266 ( .A0(\pipe_array_data[0][36] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n977));
Q_AN03 U1267 ( .A0(\pipe_array_data[0][35] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n978));
Q_AN03 U1268 ( .A0(\pipe_array_data[0][34] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n979));
Q_AN03 U1269 ( .A0(\pipe_array_data[0][33] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n980));
Q_AN03 U1270 ( .A0(\pipe_array_data[0][32] ), .A1(n1031), .A2(\pipe_array_ack[0][0] ), .Z(n981));
Q_AN03 U1271 ( .A0(\pipe_array_data[0][31] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n982));
Q_AN03 U1272 ( .A0(\pipe_array_data[0][30] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n983));
Q_AN03 U1273 ( .A0(\pipe_array_data[0][29] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n984));
Q_AN03 U1274 ( .A0(\pipe_array_data[0][28] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n985));
Q_AN03 U1275 ( .A0(\pipe_array_data[0][27] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n986));
Q_AN03 U1276 ( .A0(\pipe_array_data[0][26] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n987));
Q_AN03 U1277 ( .A0(\pipe_array_data[0][25] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n988));
Q_AN03 U1278 ( .A0(\pipe_array_data[0][24] ), .A1(n1017), .A2(\pipe_array_ack[0][0] ), .Z(n989));
Q_AN03 U1279 ( .A0(\pipe_array_data[0][23] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n990));
Q_AN03 U1280 ( .A0(\pipe_array_data[0][22] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n991));
Q_AN03 U1281 ( .A0(\pipe_array_data[0][21] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n992));
Q_AN03 U1282 ( .A0(\pipe_array_data[0][20] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n993));
Q_AN03 U1283 ( .A0(\pipe_array_data[0][19] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n994));
Q_AN03 U1284 ( .A0(\pipe_array_data[0][18] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n995));
Q_AN03 U1285 ( .A0(\pipe_array_data[0][17] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n996));
Q_AN03 U1286 ( .A0(\pipe_array_data[0][16] ), .A1(n1018), .A2(\pipe_array_ack[0][0] ), .Z(n997));
Q_AN03 U1287 ( .A0(\pipe_array_data[0][15] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n998));
Q_AN03 U1288 ( .A0(\pipe_array_data[0][14] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n999));
Q_AN03 U1289 ( .A0(\pipe_array_data[0][13] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n1000));
Q_AN03 U1290 ( .A0(\pipe_array_data[0][12] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n1001));
Q_AN03 U1291 ( .A0(\pipe_array_data[0][11] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n1002));
Q_AN03 U1292 ( .A0(\pipe_array_data[0][10] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n1003));
Q_AN03 U1293 ( .A0(\pipe_array_data[0][9] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n1004));
Q_AN03 U1294 ( .A0(\pipe_array_data[0][8] ), .A1(n1019), .A2(\pipe_array_ack[0][0] ), .Z(n1005));
Q_AN03 U1295 ( .A0(\pipe_array_data[0][7] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1006));
Q_AN03 U1296 ( .A0(\pipe_array_data[0][6] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1007));
Q_AN03 U1297 ( .A0(\pipe_array_data[0][5] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1008));
Q_AN03 U1298 ( .A0(\pipe_array_data[0][4] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1009));
Q_AN03 U1299 ( .A0(\pipe_array_data[0][3] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1010));
Q_AN03 U1300 ( .A0(\pipe_array_data[0][2] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1011));
Q_AN03 U1301 ( .A0(\pipe_array_data[0][1] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1012));
Q_AN03 U1302 ( .A0(\pipe_array_data[0][0] ), .A1(\pipe_array_ack_num_bytes[0][4] ), .A2(\pipe_array_ack[0][0] ), .Z(n1013));
Q_INV U1303 ( .A(n1028), .Z(n1014));
Q_INV U1304 ( .A(n1029), .Z(n1015));
Q_INV U1305 ( .A(n1030), .Z(n1016));
Q_INV U1306 ( .A(n1032), .Z(n1017));
Q_INV U1307 ( .A(n1033), .Z(n1018));
Q_INV U1308 ( .A(n1034), .Z(n1019));
Q_ND02 U1309 ( .A0(n1035), .A1(n1036), .Z(n1023));
Q_OR02 U1310 ( .A0(\pipe_array_ack_num_bytes[0][4] ), .A1(\pipe_array_ack_num_bytes[0][3] ), .Z(n1027));
Q_ND02 U1311 ( .A0(n1035), .A1(n1037), .Z(n1031));
Q_INV U1312 ( .A(\pipe_array_ack_num_bytes[0][4] ), .Z(n1035));
Q_ND03 U1313 ( .A0(n1038), .A1(n1039), .A2(n1035), .Z(n1020));
Q_ND03 U1314 ( .A0(n1038), .A1(n1040), .A2(n1035), .Z(n1021));
Q_ND03 U1315 ( .A0(n1038), .A1(n1041), .A2(n1035), .Z(n1022));
Q_NR02 U1316 ( .A0(\pipe_array_ack_num_bytes[0][3] ), .A1(\pipe_array_ack_num_bytes[0][2] ), .Z(n1036));
Q_ND03 U1317 ( .A0(n1038), .A1(n1042), .A2(n1035), .Z(n1024));
Q_ND03 U1318 ( .A0(n1038), .A1(n1043), .A2(n1035), .Z(n1025));
Q_ND03 U1319 ( .A0(n1038), .A1(n1044), .A2(n1035), .Z(n1026));
Q_OA21 U1320 ( .A0(n1038), .A1(n1039), .B0(n1035), .Z(n1028));
Q_OA21 U1321 ( .A0(n1038), .A1(n1040), .B0(n1035), .Z(n1029));
Q_OA21 U1322 ( .A0(n1038), .A1(n1041), .B0(n1035), .Z(n1030));
Q_ND02 U1323 ( .A0(\pipe_array_ack_num_bytes[0][3] ), .A1(\pipe_array_ack_num_bytes[0][2] ), .Z(n1037));
Q_OA21 U1324 ( .A0(n1038), .A1(n1042), .B0(n1035), .Z(n1032));
Q_OA21 U1325 ( .A0(n1038), .A1(n1043), .B0(n1035), .Z(n1033));
Q_OA21 U1326 ( .A0(n1038), .A1(n1044), .B0(n1035), .Z(n1034));
Q_INV U1327 ( .A(\pipe_array_ack_num_bytes[0][3] ), .Z(n1038));
Q_AN02 U1328 ( .A0(n1045), .A1(n1046), .Z(n1039));
Q_NR02 U1329 ( .A0(\pipe_array_ack_num_bytes[0][2] ), .A1(\pipe_array_ack_num_bytes[0][1] ), .Z(n1040));
Q_AN02 U1330 ( .A0(n1045), .A1(n1047), .Z(n1041));
Q_OR02 U1331 ( .A0(n1045), .A1(n1046), .Z(n1042));
Q_ND02 U1332 ( .A0(\pipe_array_ack_num_bytes[0][2] ), .A1(\pipe_array_ack_num_bytes[0][1] ), .Z(n1043));
Q_OR02 U1333 ( .A0(n1045), .A1(n1047), .Z(n1044));
Q_INV U1334 ( .A(\pipe_array_ack_num_bytes[0][2] ), .Z(n1045));
Q_NR02 U1335 ( .A0(\pipe_array_ack_num_bytes[0][1] ), .A1(\pipe_array_ack_num_bytes[0][0] ), .Z(n1046));
Q_ND02 U1336 ( .A0(\pipe_array_ack_num_bytes[0][1] ), .A1(\pipe_array_ack_num_bytes[0][0] ), .Z(n1047));
Q_INV U1337 ( .A(in_hash_valid), .Z(n1060));
Q_OR02 U1338 ( .A0(n1054), .A1(n1053), .Z(n1067));
Q_OR03 U1339 ( .A0(n1056), .A1(n1055), .A2(n1067), .Z(n1068));
Q_OA21 U1340 ( .A0(n1057), .A1(n1068), .B0(\pipe_array_valid[0][0] ), .Z(n1076));
Q_AN02 U1341 ( .A0(n1059), .A1(n1076), .Z(n1063));
Q_AN02 U1342 ( .A0(in_hash_valid), .A1(n1063), .Z(n1061));
Q_INV U1343 ( .A(n1076), .Z(n1064));
Q_ND02 U1344 ( .A0(in_hash_valid), .A1(n1135), .Z(n1069));
Q_NR02 U1345 ( .A0(n1069), .A1(n1064), .Z(n1070));
Q_INV U1346 ( .A(n1052), .Z(n1071));
Q_OR02 U1347 ( .A0(n1048), .A1(n1049), .Z(n1072));
Q_OR02 U1348 ( .A0(n1050), .A1(n1051), .Z(n1073));
Q_OA21 U1349 ( .A0(n1073), .A1(n1072), .B0(\pipe_array_valid[1][0] ), .Z(n1074));
Q_MX02 U1350 ( .S(n1052), .A0(n1074), .A1(\pipe_array_valid[1][0] ), .Z(n1077));
Q_AN02 U1351 ( .A0(in_hash_valid), .A1(n1077), .Z(\pipe_array_ack[1][0] ));
Q_AN02 U1352 ( .A0(n1058), .A1(\pipe_array_ack[1][0] ), .Z(n1062));
Q_AN02 U1353 ( .A0(n1099), .A1(\pipe_array_ack[1][0] ), .Z(n1075));
Q_AN02 U1354 ( .A0(in_hash_valid), .A1(n1076), .Z(\pipe_array_ack[0][0] ));
Q_NR02 U1355 ( .A0(n1060), .A1(n1077), .Z(n1078));
Q_MX02 U1356 ( .S(n1062), .A0(n1079), .A1(n1084), .Z(num_bytes_to_tx[4]));
Q_AN02 U1357 ( .A0(n1078), .A1(n1048), .Z(n1079));
Q_MX02 U1358 ( .S(n1062), .A0(n1080), .A1(n1086), .Z(num_bytes_to_tx[3]));
Q_AN02 U1359 ( .A0(n1078), .A1(n1049), .Z(n1080));
Q_MX02 U1360 ( .S(n1062), .A0(n1081), .A1(n1087), .Z(num_bytes_to_tx[2]));
Q_AN02 U1361 ( .A0(n1078), .A1(n1050), .Z(n1081));
Q_MX02 U1362 ( .S(n1062), .A0(n1082), .A1(n1089), .Z(num_bytes_to_tx[1]));
Q_AN02 U1363 ( .A0(n1078), .A1(n1051), .Z(n1082));
Q_MX02 U1364 ( .S(n1062), .A0(n1083), .A1(n1090), .Z(num_bytes_to_tx[0]));
Q_AN02 U1365 ( .A0(n1078), .A1(n1052), .Z(n1083));
Q_AD02 U1366 ( .CI(n1088), .A0(n1092), .A1(n1091), .B0(n1050), .B1(n1049), .S0(n1087), .S1(n1086), .CO(n1085));
Q_AD01 U1367 ( .CI(n1051), .A0(n1093), .B0(n1970), .S(n1089), .CO(n1088));
Q_XOR2 U1368 ( .A0(\pipe_array_byte_count[1][0] ), .A1(n1052), .Z(n1090));
Q_XNR3 U1369 ( .A0(\pipe_array_byte_count[1][4] ), .A1(n1048), .A2(n1085), .Z(n1084));
Q_INV U1370 ( .A(\pipe_array_byte_count[1][3] ), .Z(n1091));
Q_INV U1371 ( .A(\pipe_array_byte_count[1][2] ), .Z(n1092));
Q_INV U1372 ( .A(\pipe_array_byte_count[1][1] ), .Z(n1093));
Q_MX02 U1373 ( .S(n1062), .A0(n1094), .A1(\pipe_array_byte_count[1][4] ), .Z(\pipe_array_ack_num_bytes[1][4] ));
Q_AN02 U1374 ( .A0(n1075), .A1(n1048), .Z(n1094));
Q_MX02 U1375 ( .S(n1062), .A0(n1095), .A1(\pipe_array_byte_count[1][3] ), .Z(\pipe_array_ack_num_bytes[1][3] ));
Q_AN02 U1376 ( .A0(n1075), .A1(n1049), .Z(n1095));
Q_MX02 U1377 ( .S(n1062), .A0(n1096), .A1(\pipe_array_byte_count[1][2] ), .Z(\pipe_array_ack_num_bytes[1][2] ));
Q_AN02 U1378 ( .A0(n1075), .A1(n1050), .Z(n1096));
Q_MX02 U1379 ( .S(n1062), .A0(n1097), .A1(\pipe_array_byte_count[1][1] ), .Z(\pipe_array_ack_num_bytes[1][1] ));
Q_AN02 U1380 ( .A0(n1075), .A1(n1051), .Z(n1097));
Q_MX02 U1381 ( .S(n1062), .A0(n1098), .A1(\pipe_array_byte_count[1][0] ), .Z(\pipe_array_ack_num_bytes[1][0] ));
Q_AN02 U1382 ( .A0(n1075), .A1(n1052), .Z(n1098));
Q_INV U1383 ( .A(n1099), .Z(n1058));
Q_AO21 U1384 ( .A0(n1105), .A1(n1100), .B0(n1106), .Z(n1099));
Q_AO21 U1385 ( .A0(n1102), .A1(n1101), .B0(n1103), .Z(n1100));
Q_AN02 U1386 ( .A0(\pipe_array_byte_count[1][0] ), .A1(n1071), .Z(n1101));
Q_OR02 U1387 ( .A0(\pipe_array_byte_count[1][1] ), .A1(n1104), .Z(n1102));
Q_AN02 U1388 ( .A0(\pipe_array_byte_count[1][1] ), .A1(n1104), .Z(n1103));
Q_INV U1389 ( .A(n1051), .Z(n1104));
Q_OR03 U1390 ( .A0(n1108), .A1(n1109), .A2(n1107), .Z(n1106));
Q_OA21 U1391 ( .A0(\pipe_array_byte_count[1][2] ), .A1(n1111), .B0(n1110), .Z(n1105));
Q_AN03 U1392 ( .A0(\pipe_array_byte_count[1][2] ), .A1(n1111), .A2(n1110), .Z(n1109));
Q_INV U1393 ( .A(n1050), .Z(n1111));
Q_OA21 U1394 ( .A0(\pipe_array_byte_count[1][3] ), .A1(n1112), .B0(n1113), .Z(n1110));
Q_AN03 U1395 ( .A0(\pipe_array_byte_count[1][3] ), .A1(n1112), .A2(n1113), .Z(n1108));
Q_INV U1396 ( .A(n1049), .Z(n1112));
Q_OR02 U1397 ( .A0(\pipe_array_byte_count[1][4] ), .A1(n1114), .Z(n1113));
Q_AO21 U1398 ( .A0(\pipe_array_byte_count[1][4] ), .A1(n1114), .B0(\pipe_array_byte_count[1][5] ), .Z(n1107));
Q_INV U1399 ( .A(n1048), .Z(n1114));
Q_MX02 U1400 ( .S(n1063), .A0(n1115), .A1(n1120), .Z(n1048));
Q_AN02 U1401 ( .A0(n1064), .A1(n1053), .Z(n1115));
Q_MX02 U1402 ( .S(n1063), .A0(n1116), .A1(n1122), .Z(n1049));
Q_AN02 U1403 ( .A0(n1064), .A1(n1054), .Z(n1116));
Q_MX02 U1404 ( .S(n1063), .A0(n1117), .A1(n1123), .Z(n1050));
Q_AN02 U1405 ( .A0(n1064), .A1(n1055), .Z(n1117));
Q_MX02 U1406 ( .S(n1063), .A0(n1118), .A1(n1124), .Z(n1051));
Q_AN02 U1407 ( .A0(n1064), .A1(n1056), .Z(n1118));
Q_MX02 U1408 ( .S(n1063), .A0(n1119), .A1(n1126), .Z(n1052));
Q_AN02 U1409 ( .A0(n1064), .A1(n1057), .Z(n1119));
Q_AD02 U1410 ( .CI(n1971), .A0(n1128), .A1(n1127), .B0(n1055), .B1(n1054), .S0(n1123), .S1(n1122), .CO(n1121));
Q_OR02 U1411 ( .A0(n1129), .A1(n1057), .Z(n1125));
Q_XNR2 U1412 ( .A0(n1129), .A1(n1057), .Z(n1126));
Q_XNR3 U1413 ( .A0(\pipe_array_byte_count[0][4] ), .A1(n1053), .A2(n1121), .Z(n1120));
Q_INV U1414 ( .A(\pipe_array_byte_count[0][3] ), .Z(n1127));
Q_INV U1415 ( .A(\pipe_array_byte_count[0][2] ), .Z(n1128));
Q_INV U1416 ( .A(\pipe_array_byte_count[0][0] ), .Z(n1129));
Q_MX02 U1417 ( .S(n1061), .A0(n1130), .A1(\pipe_array_byte_count[0][4] ), .Z(\pipe_array_ack_num_bytes[0][4] ));
Q_AN02 U1418 ( .A0(n1070), .A1(n1053), .Z(n1130));
Q_MX02 U1419 ( .S(n1061), .A0(n1131), .A1(\pipe_array_byte_count[0][3] ), .Z(\pipe_array_ack_num_bytes[0][3] ));
Q_AN02 U1420 ( .A0(n1070), .A1(n1054), .Z(n1131));
Q_MX02 U1421 ( .S(n1061), .A0(n1132), .A1(\pipe_array_byte_count[0][2] ), .Z(\pipe_array_ack_num_bytes[0][2] ));
Q_AN02 U1422 ( .A0(n1070), .A1(n1055), .Z(n1132));
Q_MX02 U1423 ( .S(n1061), .A0(n1133), .A1(\pipe_array_byte_count[0][1] ), .Z(\pipe_array_ack_num_bytes[0][1] ));
Q_AN02 U1424 ( .A0(n1070), .A1(n1056), .Z(n1133));
Q_MX02 U1425 ( .S(n1061), .A0(n1134), .A1(\pipe_array_byte_count[0][0] ), .Z(\pipe_array_ack_num_bytes[0][0] ));
Q_AN02 U1426 ( .A0(n1070), .A1(n1057), .Z(n1134));
Q_AN02 U1427 ( .A0(in_hash_valid), .A1(n1066), .Z(in_hash_eof));
Q_INV U1428 ( .A(n1135), .Z(n1059));
Q_AO21 U1429 ( .A0(n1142), .A1(n1136), .B0(n1143), .Z(n1135));
Q_AO21 U1430 ( .A0(n1139), .A1(n1137), .B0(n1140), .Z(n1136));
Q_AN02 U1431 ( .A0(\pipe_array_byte_count[0][0] ), .A1(n1138), .Z(n1137));
Q_INV U1432 ( .A(n1057), .Z(n1138));
Q_OR02 U1433 ( .A0(\pipe_array_byte_count[0][1] ), .A1(n1141), .Z(n1139));
Q_AN02 U1434 ( .A0(\pipe_array_byte_count[0][1] ), .A1(n1141), .Z(n1140));
Q_INV U1435 ( .A(n1056), .Z(n1141));
Q_OR03 U1436 ( .A0(n1145), .A1(n1146), .A2(n1144), .Z(n1143));
Q_OA21 U1437 ( .A0(\pipe_array_byte_count[0][2] ), .A1(n1148), .B0(n1147), .Z(n1142));
Q_AN03 U1438 ( .A0(\pipe_array_byte_count[0][2] ), .A1(n1148), .A2(n1147), .Z(n1146));
Q_INV U1439 ( .A(n1055), .Z(n1148));
Q_OA21 U1440 ( .A0(\pipe_array_byte_count[0][3] ), .A1(n1149), .B0(n1150), .Z(n1147));
Q_AN03 U1441 ( .A0(\pipe_array_byte_count[0][3] ), .A1(n1149), .A2(n1150), .Z(n1145));
Q_INV U1442 ( .A(n1054), .Z(n1149));
Q_OR02 U1443 ( .A0(\pipe_array_byte_count[0][4] ), .A1(n1151), .Z(n1150));
Q_AO21 U1444 ( .A0(\pipe_array_byte_count[0][4] ), .A1(n1151), .B0(\pipe_array_byte_count[0][5] ), .Z(n1144));
Q_INV U1445 ( .A(n1053), .Z(n1151));
Q_OR02 U1446 ( .A0(n1152), .A1(num_bytes_remaining[4]), .Z(n1053));
Q_INV U1447 ( .A(n1065), .Z(n1152));
Q_AN02 U1448 ( .A0(n1065), .A1(num_bytes_remaining[3]), .Z(n1054));
Q_AN02 U1449 ( .A0(n1065), .A1(num_bytes_remaining[2]), .Z(n1055));
Q_AN02 U1450 ( .A0(n1065), .A1(num_bytes_remaining[1]), .Z(n1056));
Q_AN02 U1451 ( .A0(n1065), .A1(num_bytes_remaining[0]), .Z(n1057));
Q_OA21 U1452 ( .A0(n1156), .A1(num_bytes_remaining[4]), .B0(in_hash_valid), .Z(in_hash_num_bytes[4]));
Q_AN03 U1453 ( .A0(n1066), .A1(num_bytes_remaining[3]), .A2(in_hash_valid), .Z(in_hash_num_bytes[3]));
Q_AN03 U1454 ( .A0(n1066), .A1(num_bytes_remaining[2]), .A2(in_hash_valid), .Z(in_hash_num_bytes[2]));
Q_AN03 U1455 ( .A0(n1066), .A1(num_bytes_remaining[1]), .A2(in_hash_valid), .Z(in_hash_num_bytes[1]));
Q_AN03 U1456 ( .A0(n1066), .A1(num_bytes_remaining[0]), .A2(in_hash_valid), .Z(in_hash_num_bytes[0]));
Q_AN03 U1457 ( .A0(n1066), .A1(n1153), .A2(in_hash_valid), .Z(kdfstream_cmdfifo_ack));
Q_NR02 U1458 ( .A0(n1155), .A1(n1154), .Z(n1153));
Q_XOR2 U1459 ( .A0(iter_num[1]), .A1(cmdfifo_kdfstream_cmd[1]), .Z(n1154));
Q_XOR2 U1460 ( .A0(iter_num[0]), .A1(cmdfifo_kdfstream_cmd[0]), .Z(n1155));
Q_INV U1461 ( .A(n1156), .Z(n1066));
Q_AO21 U1462 ( .A0(num_bytes_remaining[4]), .A1(n1157), .B0(n1158), .Z(n1156));
Q_OR03 U1463 ( .A0(num_bytes_remaining[2]), .A1(num_bytes_remaining[1]), .A2(num_bytes_remaining[0]), .Z(n1157));
Q_OR02 U1464 ( .A0(num_bytes_remaining[6]), .A1(num_bytes_remaining[5]), .Z(n1159));
Q_AO21 U1465 ( .A0(num_bytes_remaining[4]), .A1(num_bytes_remaining[3]), .B0(n1159), .Z(n1158));
Q_AN02 U1466 ( .A0(n1160), .A1(n1161), .Z(n1065));
Q_NR02 U1467 ( .A0(num_bytes_remaining[6]), .A1(num_bytes_remaining[5]), .Z(n1160));
Q_AN02 U1468 ( .A0(st_tx_data), .A1(n1162), .Z(in_hash_valid));
Q_INV U1469 ( .A(hash_in_stall), .Z(n1162));
Q_INV U1470 ( .A(st_tx_data), .Z(program_pipes));
Q_FDP1 \num_bytes_remaining_REG[0] ( .CK(clk), .R(rst_n), .D(n1163), .Q(num_bytes_remaining[0]), .QN( ));
Q_FDP1 \num_bytes_remaining_REG[1] ( .CK(clk), .R(rst_n), .D(n1164), .Q(num_bytes_remaining[1]), .QN( ));
Q_FDP1 \num_bytes_remaining_REG[2] ( .CK(clk), .R(rst_n), .D(n1165), .Q(num_bytes_remaining[2]), .QN( ));
Q_FDP1 \num_bytes_remaining_REG[3] ( .CK(clk), .R(rst_n), .D(n1166), .Q(num_bytes_remaining[3]), .QN( ));
Q_FDP1 \num_bytes_remaining_REG[4] ( .CK(clk), .R(rst_n), .D(n1167), .Q(num_bytes_remaining[4]), .QN(n1161));
Q_FDP1 \num_bytes_remaining_REG[5] ( .CK(clk), .R(rst_n), .D(n1168), .Q(num_bytes_remaining[5]), .QN( ));
Q_FDP1 \num_bytes_remaining_REG[6] ( .CK(clk), .R(rst_n), .D(n1169), .Q(num_bytes_remaining[6]), .QN( ));
Q_MX02 U1478 ( .S(st_tx_data), .A0(hash_cmd_in[11]), .A1(n1170), .Z(n1169));
Q_MX02 U1479 ( .S(st_tx_data), .A0(hash_cmd_in[9]), .A1(n1172), .Z(n1168));
Q_MX02 U1480 ( .S(st_tx_data), .A0(hash_cmd_in[8]), .A1(n1174), .Z(n1167));
Q_MX02 U1481 ( .S(st_tx_data), .A0(hash_cmd_in[7]), .A1(n1176), .Z(n1166));
Q_MX02 U1482 ( .S(st_tx_data), .A0(hash_cmd_in[6]), .A1(n1177), .Z(n1165));
Q_MX02 U1483 ( .S(st_tx_data), .A0(hash_cmd_in[5]), .A1(n1179), .Z(n1164));
Q_MX02 U1484 ( .S(st_tx_data), .A0(hash_cmd_in[4]), .A1(n1181), .Z(n1163));
Q_XNR2 U1485 ( .A0(num_bytes_remaining[6]), .A1(n1171), .Z(n1170));
Q_OR02 U1486 ( .A0(num_bytes_remaining[5]), .A1(n1173), .Z(n1171));
Q_XNR2 U1487 ( .A0(num_bytes_remaining[5]), .A1(n1173), .Z(n1172));
Q_AD01 U1488 ( .CI(n1175), .A0(num_bytes_remaining[4]), .B0(n1182), .S(n1174), .CO(n1173));
Q_AD02 U1489 ( .CI(n1178), .A0(num_bytes_remaining[2]), .A1(num_bytes_remaining[3]), .B0(n1184), .B1(n1183), .S0(n1177), .S1(n1176), .CO(n1175));
Q_AD01 U1490 ( .CI(n1180), .A0(num_bytes_remaining[1]), .B0(n1185), .S(n1179), .CO(n1178));
Q_OR02 U1491 ( .A0(num_bytes_remaining[0]), .A1(n1186), .Z(n1180));
Q_XNR2 U1492 ( .A0(num_bytes_remaining[0]), .A1(n1186), .Z(n1181));
Q_INV U1493 ( .A(in_hash_num_bytes[4]), .Z(n1182));
Q_INV U1494 ( .A(in_hash_num_bytes[3]), .Z(n1183));
Q_INV U1495 ( .A(in_hash_num_bytes[2]), .Z(n1184));
Q_INV U1496 ( .A(in_hash_num_bytes[1]), .Z(n1185));
Q_INV U1497 ( .A(in_hash_num_bytes[0]), .Z(n1186));
Q_AN02 U1498 ( .A0(cmd_il_valid), .A1(n1187), .Z(cmd_dgl_data_size[0]));
Q_NR02 U1499 ( .A0(st_tx_data), .A1(n1187), .Z(n1189));
Q_INV U1500 ( .A(cmdfifo_kdfstream_cmd[0]), .Z(n1195));
Q_INV U1501 ( .A(cmdfifo_kdfstream_cmd[1]), .Z(n1194));
Q_AN02 U1502 ( .A0(n1194), .A1(cmdfifo_kdfstream_cmd[0]), .Z(n1196));
Q_OR02 U1503 ( .A0(cmdfifo_kdfstream_cmd[1]), .A1(n1196), .Z(n1199));
Q_AN02 U1504 ( .A0(n1188), .A1(n1199), .Z(n1192));
Q_AN02 U1505 ( .A0(cmdfifo_kdfstream_cmd[1]), .A1(n1195), .Z(n1197));
Q_OR02 U1506 ( .A0(n2), .A1(n1196), .Z(n1190));
Q_MX02 U1507 ( .S(n1188), .A0(cmdfifo_kdfstream_cmd[0]), .A1(n1197), .Z(n1191));
Q_INV U1508 ( .A(n1192), .Z(n1198));
Q_AN02 U1509 ( .A0(n1199), .A1(n1198), .Z(n1193));
Q_AN02 U1510 ( .A0(cmd_il_valid), .A1(n1188), .Z(cmd_dgl_data_size[5]));
Q_NR02 U1511 ( .A0(st_tx_data), .A1(n1188), .Z(cmd_dgl_data_size[4]));
Q_AN02 U1512 ( .A0(cmd_il_valid), .A1(n1200), .Z(cmd_il_data_size[5]));
Q_AN02 U1513 ( .A0(cmd_il_valid), .A1(n1202), .Z(cmd_il_data_size[4]));
Q_AN02 U1514 ( .A0(cmd_il_valid), .A1(n1204), .Z(cmd_il_data_size[3]));
Q_NR02 U1515 ( .A0(st_tx_data), .A1(n7), .Z(cmd_il_data_size[2]));
Q_AN02 U1516 ( .A0(cmd_il_valid), .A1(n8), .Z(cmd_il_data_size[1]));
Q_AN02 U1517 ( .A0(cmd_il_valid), .A1(n9), .Z(cmd_il_data_size[0]));
Q_AN02 U1518 ( .A0(cmd_il_valid), .A1(iter_num[1]), .Z(cmd_il_data[257]));
Q_AN02 U1519 ( .A0(cmd_il_valid), .A1(iter_num[0]), .Z(cmd_il_data[256]));
Q_AN02 U1520 ( .A0(cmd_il_valid), .A1(n10), .Z(cmd_il_data[255]));
Q_AN02 U1521 ( .A0(cmd_il_valid), .A1(n11), .Z(cmd_il_data[254]));
Q_AN02 U1522 ( .A0(cmd_il_valid), .A1(n12), .Z(cmd_il_data[253]));
Q_AN02 U1523 ( .A0(cmd_il_valid), .A1(n13), .Z(cmd_il_data[252]));
Q_AN02 U1524 ( .A0(cmd_il_valid), .A1(n14), .Z(cmd_il_data[251]));
Q_AN02 U1525 ( .A0(cmd_il_valid), .A1(n15), .Z(cmd_il_data[250]));
Q_AN02 U1526 ( .A0(cmd_il_valid), .A1(n16), .Z(cmd_il_data[249]));
Q_AN02 U1527 ( .A0(cmd_il_valid), .A1(n17), .Z(cmd_il_data[248]));
Q_AN02 U1528 ( .A0(cmd_il_valid), .A1(n18), .Z(cmd_il_data[247]));
Q_AN02 U1529 ( .A0(cmd_il_valid), .A1(n19), .Z(cmd_il_data[246]));
Q_AN02 U1530 ( .A0(cmd_il_valid), .A1(n20), .Z(cmd_il_data[245]));
Q_AN02 U1531 ( .A0(cmd_il_valid), .A1(n21), .Z(cmd_il_data[244]));
Q_AN02 U1532 ( .A0(cmd_il_valid), .A1(n22), .Z(cmd_il_data[243]));
Q_AN02 U1533 ( .A0(cmd_il_valid), .A1(n23), .Z(cmd_il_data[242]));
Q_AN02 U1534 ( .A0(cmd_il_valid), .A1(n24), .Z(cmd_il_data[241]));
Q_AN02 U1535 ( .A0(cmd_il_valid), .A1(n25), .Z(cmd_il_data[240]));
Q_AN02 U1536 ( .A0(cmd_il_valid), .A1(n26), .Z(cmd_il_data[239]));
Q_AN02 U1537 ( .A0(cmd_il_valid), .A1(n27), .Z(cmd_il_data[238]));
Q_AN02 U1538 ( .A0(cmd_il_valid), .A1(n28), .Z(cmd_il_data[237]));
Q_AN02 U1539 ( .A0(cmd_il_valid), .A1(n29), .Z(cmd_il_data[236]));
Q_AN02 U1540 ( .A0(cmd_il_valid), .A1(n30), .Z(cmd_il_data[235]));
Q_AN02 U1541 ( .A0(cmd_il_valid), .A1(n31), .Z(cmd_il_data[234]));
Q_AN02 U1542 ( .A0(cmd_il_valid), .A1(n32), .Z(cmd_il_data[233]));
Q_AN02 U1543 ( .A0(cmd_il_valid), .A1(n33), .Z(cmd_il_data[232]));
Q_AN02 U1544 ( .A0(cmd_il_valid), .A1(n34), .Z(cmd_il_data[231]));
Q_AN02 U1545 ( .A0(cmd_il_valid), .A1(n35), .Z(cmd_il_data[230]));
Q_AN02 U1546 ( .A0(cmd_il_valid), .A1(n36), .Z(cmd_il_data[229]));
Q_AN02 U1547 ( .A0(cmd_il_valid), .A1(n37), .Z(cmd_il_data[228]));
Q_AN02 U1548 ( .A0(cmd_il_valid), .A1(n38), .Z(cmd_il_data[227]));
Q_AN02 U1549 ( .A0(cmd_il_valid), .A1(n39), .Z(cmd_il_data[226]));
Q_AN02 U1550 ( .A0(cmd_il_valid), .A1(n40), .Z(cmd_il_data[225]));
Q_AN02 U1551 ( .A0(cmd_il_valid), .A1(n41), .Z(cmd_il_data[224]));
Q_AN02 U1552 ( .A0(cmd_il_valid), .A1(n42), .Z(cmd_il_data[223]));
Q_AN02 U1553 ( .A0(cmd_il_valid), .A1(n43), .Z(cmd_il_data[222]));
Q_AN02 U1554 ( .A0(cmd_il_valid), .A1(n44), .Z(cmd_il_data[221]));
Q_AN02 U1555 ( .A0(cmd_il_valid), .A1(n45), .Z(cmd_il_data[220]));
Q_AN02 U1556 ( .A0(cmd_il_valid), .A1(n46), .Z(cmd_il_data[219]));
Q_AN02 U1557 ( .A0(cmd_il_valid), .A1(n47), .Z(cmd_il_data[218]));
Q_AN02 U1558 ( .A0(cmd_il_valid), .A1(n48), .Z(cmd_il_data[217]));
Q_AN02 U1559 ( .A0(cmd_il_valid), .A1(n49), .Z(cmd_il_data[216]));
Q_AN02 U1560 ( .A0(cmd_il_valid), .A1(n50), .Z(cmd_il_data[215]));
Q_AN02 U1561 ( .A0(cmd_il_valid), .A1(n51), .Z(cmd_il_data[214]));
Q_AN02 U1562 ( .A0(cmd_il_valid), .A1(n52), .Z(cmd_il_data[213]));
Q_AN02 U1563 ( .A0(cmd_il_valid), .A1(n53), .Z(cmd_il_data[212]));
Q_AN02 U1564 ( .A0(cmd_il_valid), .A1(n54), .Z(cmd_il_data[211]));
Q_AN02 U1565 ( .A0(cmd_il_valid), .A1(n55), .Z(cmd_il_data[210]));
Q_AN02 U1566 ( .A0(cmd_il_valid), .A1(n56), .Z(cmd_il_data[209]));
Q_AN02 U1567 ( .A0(cmd_il_valid), .A1(n57), .Z(cmd_il_data[208]));
Q_AN02 U1568 ( .A0(cmd_il_valid), .A1(n58), .Z(cmd_il_data[207]));
Q_AN02 U1569 ( .A0(cmd_il_valid), .A1(n59), .Z(cmd_il_data[206]));
Q_AN02 U1570 ( .A0(cmd_il_valid), .A1(n60), .Z(cmd_il_data[205]));
Q_AN02 U1571 ( .A0(cmd_il_valid), .A1(n61), .Z(cmd_il_data[204]));
Q_AN02 U1572 ( .A0(cmd_il_valid), .A1(n62), .Z(cmd_il_data[203]));
Q_AN02 U1573 ( .A0(cmd_il_valid), .A1(n63), .Z(cmd_il_data[202]));
Q_AN02 U1574 ( .A0(cmd_il_valid), .A1(n64), .Z(cmd_il_data[201]));
Q_AN02 U1575 ( .A0(cmd_il_valid), .A1(n65), .Z(cmd_il_data[200]));
Q_AN02 U1576 ( .A0(cmd_il_valid), .A1(n66), .Z(cmd_il_data[199]));
Q_AN02 U1577 ( .A0(cmd_il_valid), .A1(n67), .Z(cmd_il_data[198]));
Q_AN02 U1578 ( .A0(cmd_il_valid), .A1(n68), .Z(cmd_il_data[197]));
Q_AN02 U1579 ( .A0(cmd_il_valid), .A1(n69), .Z(cmd_il_data[196]));
Q_AN02 U1580 ( .A0(cmd_il_valid), .A1(n70), .Z(cmd_il_data[195]));
Q_AN02 U1581 ( .A0(cmd_il_valid), .A1(n71), .Z(cmd_il_data[194]));
Q_AN02 U1582 ( .A0(cmd_il_valid), .A1(n72), .Z(cmd_il_data[193]));
Q_AN02 U1583 ( .A0(cmd_il_valid), .A1(n73), .Z(cmd_il_data[192]));
Q_AN02 U1584 ( .A0(cmd_il_valid), .A1(n74), .Z(cmd_il_data[191]));
Q_AN02 U1585 ( .A0(cmd_il_valid), .A1(n75), .Z(cmd_il_data[190]));
Q_AN02 U1586 ( .A0(cmd_il_valid), .A1(n76), .Z(cmd_il_data[189]));
Q_AN02 U1587 ( .A0(cmd_il_valid), .A1(n77), .Z(cmd_il_data[188]));
Q_AN02 U1588 ( .A0(cmd_il_valid), .A1(n78), .Z(cmd_il_data[187]));
Q_AN02 U1589 ( .A0(cmd_il_valid), .A1(n79), .Z(cmd_il_data[186]));
Q_AN02 U1590 ( .A0(cmd_il_valid), .A1(n80), .Z(cmd_il_data[185]));
Q_AN02 U1591 ( .A0(cmd_il_valid), .A1(n81), .Z(cmd_il_data[184]));
Q_AN02 U1592 ( .A0(cmd_il_valid), .A1(n82), .Z(cmd_il_data[183]));
Q_AN02 U1593 ( .A0(cmd_il_valid), .A1(n83), .Z(cmd_il_data[182]));
Q_AN02 U1594 ( .A0(cmd_il_valid), .A1(n84), .Z(cmd_il_data[181]));
Q_AN02 U1595 ( .A0(cmd_il_valid), .A1(n85), .Z(cmd_il_data[180]));
Q_AN02 U1596 ( .A0(cmd_il_valid), .A1(n86), .Z(cmd_il_data[179]));
Q_AN02 U1597 ( .A0(cmd_il_valid), .A1(n87), .Z(cmd_il_data[178]));
Q_AN02 U1598 ( .A0(cmd_il_valid), .A1(n88), .Z(cmd_il_data[177]));
Q_AN02 U1599 ( .A0(cmd_il_valid), .A1(n89), .Z(cmd_il_data[176]));
Q_AN02 U1600 ( .A0(cmd_il_valid), .A1(n90), .Z(cmd_il_data[175]));
Q_AN02 U1601 ( .A0(cmd_il_valid), .A1(n91), .Z(cmd_il_data[174]));
Q_AN02 U1602 ( .A0(cmd_il_valid), .A1(n92), .Z(cmd_il_data[173]));
Q_AN02 U1603 ( .A0(cmd_il_valid), .A1(n93), .Z(cmd_il_data[172]));
Q_AN02 U1604 ( .A0(cmd_il_valid), .A1(n94), .Z(cmd_il_data[171]));
Q_AN02 U1605 ( .A0(cmd_il_valid), .A1(n95), .Z(cmd_il_data[170]));
Q_AN02 U1606 ( .A0(cmd_il_valid), .A1(n96), .Z(cmd_il_data[169]));
Q_AN02 U1607 ( .A0(cmd_il_valid), .A1(n97), .Z(cmd_il_data[168]));
Q_AN02 U1608 ( .A0(cmd_il_valid), .A1(n98), .Z(cmd_il_data[167]));
Q_AN02 U1609 ( .A0(cmd_il_valid), .A1(n99), .Z(cmd_il_data[166]));
Q_AN02 U1610 ( .A0(cmd_il_valid), .A1(n100), .Z(cmd_il_data[165]));
Q_AN02 U1611 ( .A0(cmd_il_valid), .A1(n101), .Z(cmd_il_data[164]));
Q_AN02 U1612 ( .A0(cmd_il_valid), .A1(n102), .Z(cmd_il_data[163]));
Q_AN02 U1613 ( .A0(cmd_il_valid), .A1(n103), .Z(cmd_il_data[162]));
Q_AN02 U1614 ( .A0(cmd_il_valid), .A1(n104), .Z(cmd_il_data[161]));
Q_AN02 U1615 ( .A0(cmd_il_valid), .A1(n105), .Z(cmd_il_data[160]));
Q_AN02 U1616 ( .A0(cmd_il_valid), .A1(n106), .Z(cmd_il_data[159]));
Q_AN02 U1617 ( .A0(cmd_il_valid), .A1(n107), .Z(cmd_il_data[158]));
Q_AN02 U1618 ( .A0(cmd_il_valid), .A1(n108), .Z(cmd_il_data[157]));
Q_AN02 U1619 ( .A0(cmd_il_valid), .A1(n109), .Z(cmd_il_data[156]));
Q_AN02 U1620 ( .A0(cmd_il_valid), .A1(n110), .Z(cmd_il_data[155]));
Q_AN02 U1621 ( .A0(cmd_il_valid), .A1(n111), .Z(cmd_il_data[154]));
Q_AN02 U1622 ( .A0(cmd_il_valid), .A1(n112), .Z(cmd_il_data[153]));
Q_AN02 U1623 ( .A0(cmd_il_valid), .A1(n113), .Z(cmd_il_data[152]));
Q_AN02 U1624 ( .A0(cmd_il_valid), .A1(n114), .Z(cmd_il_data[151]));
Q_AN02 U1625 ( .A0(cmd_il_valid), .A1(n115), .Z(cmd_il_data[150]));
Q_AN02 U1626 ( .A0(cmd_il_valid), .A1(n116), .Z(cmd_il_data[149]));
Q_AN02 U1627 ( .A0(cmd_il_valid), .A1(n117), .Z(cmd_il_data[148]));
Q_AN02 U1628 ( .A0(cmd_il_valid), .A1(n118), .Z(cmd_il_data[147]));
Q_AN02 U1629 ( .A0(cmd_il_valid), .A1(n119), .Z(cmd_il_data[146]));
Q_AN02 U1630 ( .A0(cmd_il_valid), .A1(n120), .Z(cmd_il_data[145]));
Q_AN02 U1631 ( .A0(cmd_il_valid), .A1(n121), .Z(cmd_il_data[144]));
Q_AN02 U1632 ( .A0(cmd_il_valid), .A1(n122), .Z(cmd_il_data[143]));
Q_AN02 U1633 ( .A0(cmd_il_valid), .A1(n123), .Z(cmd_il_data[142]));
Q_AN02 U1634 ( .A0(cmd_il_valid), .A1(n124), .Z(cmd_il_data[141]));
Q_AN02 U1635 ( .A0(cmd_il_valid), .A1(n125), .Z(cmd_il_data[140]));
Q_AN02 U1636 ( .A0(cmd_il_valid), .A1(n126), .Z(cmd_il_data[139]));
Q_AN02 U1637 ( .A0(cmd_il_valid), .A1(n127), .Z(cmd_il_data[138]));
Q_AN02 U1638 ( .A0(cmd_il_valid), .A1(n128), .Z(cmd_il_data[137]));
Q_AN02 U1639 ( .A0(cmd_il_valid), .A1(n129), .Z(cmd_il_data[136]));
Q_AN02 U1640 ( .A0(cmd_il_valid), .A1(n130), .Z(cmd_il_data[135]));
Q_AN02 U1641 ( .A0(cmd_il_valid), .A1(n131), .Z(cmd_il_data[134]));
Q_AN02 U1642 ( .A0(cmd_il_valid), .A1(n132), .Z(cmd_il_data[133]));
Q_AN02 U1643 ( .A0(cmd_il_valid), .A1(n133), .Z(cmd_il_data[132]));
Q_AN02 U1644 ( .A0(cmd_il_valid), .A1(n134), .Z(cmd_il_data[131]));
Q_AN02 U1645 ( .A0(cmd_il_valid), .A1(n135), .Z(cmd_il_data[130]));
Q_AN02 U1646 ( .A0(cmd_il_valid), .A1(n136), .Z(cmd_il_data[129]));
Q_AN02 U1647 ( .A0(cmd_il_valid), .A1(n137), .Z(cmd_il_data[128]));
Q_AN02 U1648 ( .A0(cmd_il_valid), .A1(n138), .Z(cmd_il_data[127]));
Q_AN02 U1649 ( .A0(cmd_il_valid), .A1(n139), .Z(cmd_il_data[126]));
Q_AN02 U1650 ( .A0(cmd_il_valid), .A1(n140), .Z(cmd_il_data[125]));
Q_AN02 U1651 ( .A0(cmd_il_valid), .A1(n141), .Z(cmd_il_data[124]));
Q_AN02 U1652 ( .A0(cmd_il_valid), .A1(n142), .Z(cmd_il_data[123]));
Q_AN02 U1653 ( .A0(cmd_il_valid), .A1(n143), .Z(cmd_il_data[122]));
Q_AN02 U1654 ( .A0(cmd_il_valid), .A1(n144), .Z(cmd_il_data[121]));
Q_AN02 U1655 ( .A0(cmd_il_valid), .A1(n145), .Z(cmd_il_data[120]));
Q_AN02 U1656 ( .A0(cmd_il_valid), .A1(n146), .Z(cmd_il_data[119]));
Q_AN02 U1657 ( .A0(cmd_il_valid), .A1(n147), .Z(cmd_il_data[118]));
Q_AN02 U1658 ( .A0(cmd_il_valid), .A1(n148), .Z(cmd_il_data[117]));
Q_AN02 U1659 ( .A0(cmd_il_valid), .A1(n149), .Z(cmd_il_data[116]));
Q_AN02 U1660 ( .A0(cmd_il_valid), .A1(n150), .Z(cmd_il_data[115]));
Q_AN02 U1661 ( .A0(cmd_il_valid), .A1(n151), .Z(cmd_il_data[114]));
Q_AN02 U1662 ( .A0(cmd_il_valid), .A1(n152), .Z(cmd_il_data[113]));
Q_AN02 U1663 ( .A0(cmd_il_valid), .A1(n153), .Z(cmd_il_data[112]));
Q_AN02 U1664 ( .A0(cmd_il_valid), .A1(n154), .Z(cmd_il_data[111]));
Q_AN02 U1665 ( .A0(cmd_il_valid), .A1(n155), .Z(cmd_il_data[110]));
Q_AN02 U1666 ( .A0(cmd_il_valid), .A1(n156), .Z(cmd_il_data[109]));
Q_AN02 U1667 ( .A0(cmd_il_valid), .A1(n157), .Z(cmd_il_data[108]));
Q_AN02 U1668 ( .A0(cmd_il_valid), .A1(n158), .Z(cmd_il_data[107]));
Q_AN02 U1669 ( .A0(cmd_il_valid), .A1(n159), .Z(cmd_il_data[106]));
Q_AN02 U1670 ( .A0(cmd_il_valid), .A1(n160), .Z(cmd_il_data[105]));
Q_AN02 U1671 ( .A0(cmd_il_valid), .A1(n161), .Z(cmd_il_data[104]));
Q_AN02 U1672 ( .A0(cmd_il_valid), .A1(n162), .Z(cmd_il_data[103]));
Q_AN02 U1673 ( .A0(cmd_il_valid), .A1(n163), .Z(cmd_il_data[102]));
Q_AN02 U1674 ( .A0(cmd_il_valid), .A1(n164), .Z(cmd_il_data[101]));
Q_AN02 U1675 ( .A0(cmd_il_valid), .A1(n165), .Z(cmd_il_data[100]));
Q_AN02 U1676 ( .A0(cmd_il_valid), .A1(n166), .Z(cmd_il_data[99]));
Q_AN02 U1677 ( .A0(cmd_il_valid), .A1(n167), .Z(cmd_il_data[98]));
Q_AN02 U1678 ( .A0(cmd_il_valid), .A1(n168), .Z(cmd_il_data[97]));
Q_AN02 U1679 ( .A0(cmd_il_valid), .A1(n169), .Z(cmd_il_data[96]));
Q_AN02 U1680 ( .A0(cmd_il_valid), .A1(n170), .Z(cmd_il_data[95]));
Q_AN02 U1681 ( .A0(cmd_il_valid), .A1(n171), .Z(cmd_il_data[94]));
Q_AN02 U1682 ( .A0(cmd_il_valid), .A1(n172), .Z(cmd_il_data[93]));
Q_AN02 U1683 ( .A0(cmd_il_valid), .A1(n173), .Z(cmd_il_data[92]));
Q_AN02 U1684 ( .A0(cmd_il_valid), .A1(n174), .Z(cmd_il_data[91]));
Q_AN02 U1685 ( .A0(cmd_il_valid), .A1(n175), .Z(cmd_il_data[90]));
Q_AN02 U1686 ( .A0(cmd_il_valid), .A1(n176), .Z(cmd_il_data[89]));
Q_AN02 U1687 ( .A0(cmd_il_valid), .A1(n177), .Z(cmd_il_data[88]));
Q_AN02 U1688 ( .A0(cmd_il_valid), .A1(n178), .Z(cmd_il_data[87]));
Q_AN02 U1689 ( .A0(cmd_il_valid), .A1(n179), .Z(cmd_il_data[86]));
Q_AN02 U1690 ( .A0(cmd_il_valid), .A1(n180), .Z(cmd_il_data[85]));
Q_AN02 U1691 ( .A0(cmd_il_valid), .A1(n181), .Z(cmd_il_data[84]));
Q_AN02 U1692 ( .A0(cmd_il_valid), .A1(n182), .Z(cmd_il_data[83]));
Q_AN02 U1693 ( .A0(cmd_il_valid), .A1(n183), .Z(cmd_il_data[82]));
Q_AN02 U1694 ( .A0(cmd_il_valid), .A1(n184), .Z(cmd_il_data[81]));
Q_AN02 U1695 ( .A0(cmd_il_valid), .A1(n185), .Z(cmd_il_data[80]));
Q_AN02 U1696 ( .A0(cmd_il_valid), .A1(n186), .Z(cmd_il_data[79]));
Q_AN02 U1697 ( .A0(cmd_il_valid), .A1(n187), .Z(cmd_il_data[78]));
Q_AN02 U1698 ( .A0(cmd_il_valid), .A1(n188), .Z(cmd_il_data[77]));
Q_AN02 U1699 ( .A0(cmd_il_valid), .A1(n189), .Z(cmd_il_data[76]));
Q_AN02 U1700 ( .A0(cmd_il_valid), .A1(n190), .Z(cmd_il_data[75]));
Q_AN02 U1701 ( .A0(cmd_il_valid), .A1(n191), .Z(cmd_il_data[74]));
Q_AN02 U1702 ( .A0(cmd_il_valid), .A1(n192), .Z(cmd_il_data[73]));
Q_AN02 U1703 ( .A0(cmd_il_valid), .A1(n193), .Z(cmd_il_data[72]));
Q_AN02 U1704 ( .A0(cmd_il_valid), .A1(n194), .Z(cmd_il_data[71]));
Q_AN02 U1705 ( .A0(cmd_il_valid), .A1(n195), .Z(cmd_il_data[70]));
Q_AN02 U1706 ( .A0(cmd_il_valid), .A1(n196), .Z(cmd_il_data[69]));
Q_AN02 U1707 ( .A0(cmd_il_valid), .A1(n197), .Z(cmd_il_data[68]));
Q_AN02 U1708 ( .A0(cmd_il_valid), .A1(n198), .Z(cmd_il_data[67]));
Q_AN02 U1709 ( .A0(cmd_il_valid), .A1(n199), .Z(cmd_il_data[66]));
Q_AN02 U1710 ( .A0(cmd_il_valid), .A1(n200), .Z(cmd_il_data[65]));
Q_AN02 U1711 ( .A0(cmd_il_valid), .A1(n201), .Z(cmd_il_data[64]));
Q_AN02 U1712 ( .A0(cmd_il_valid), .A1(n202), .Z(cmd_il_data[63]));
Q_AN02 U1713 ( .A0(cmd_il_valid), .A1(n203), .Z(cmd_il_data[62]));
Q_AN02 U1714 ( .A0(cmd_il_valid), .A1(n204), .Z(cmd_il_data[61]));
Q_AN02 U1715 ( .A0(cmd_il_valid), .A1(n205), .Z(cmd_il_data[60]));
Q_AN02 U1716 ( .A0(cmd_il_valid), .A1(n206), .Z(cmd_il_data[59]));
Q_AN02 U1717 ( .A0(cmd_il_valid), .A1(n207), .Z(cmd_il_data[58]));
Q_AN02 U1718 ( .A0(cmd_il_valid), .A1(n208), .Z(cmd_il_data[57]));
Q_AN02 U1719 ( .A0(cmd_il_valid), .A1(n209), .Z(cmd_il_data[56]));
Q_AN02 U1720 ( .A0(cmd_il_valid), .A1(n210), .Z(cmd_il_data[55]));
Q_AN02 U1721 ( .A0(cmd_il_valid), .A1(n211), .Z(cmd_il_data[54]));
Q_AN02 U1722 ( .A0(cmd_il_valid), .A1(n212), .Z(cmd_il_data[53]));
Q_AN02 U1723 ( .A0(cmd_il_valid), .A1(n213), .Z(cmd_il_data[52]));
Q_AN02 U1724 ( .A0(cmd_il_valid), .A1(n214), .Z(cmd_il_data[51]));
Q_AN02 U1725 ( .A0(cmd_il_valid), .A1(n215), .Z(cmd_il_data[50]));
Q_AN02 U1726 ( .A0(cmd_il_valid), .A1(n216), .Z(cmd_il_data[49]));
Q_AN02 U1727 ( .A0(cmd_il_valid), .A1(n217), .Z(cmd_il_data[48]));
Q_AN02 U1728 ( .A0(cmd_il_valid), .A1(n218), .Z(cmd_il_data[47]));
Q_AN02 U1729 ( .A0(cmd_il_valid), .A1(n219), .Z(cmd_il_data[46]));
Q_AN02 U1730 ( .A0(cmd_il_valid), .A1(n220), .Z(cmd_il_data[45]));
Q_AN02 U1731 ( .A0(cmd_il_valid), .A1(n221), .Z(cmd_il_data[44]));
Q_AN02 U1732 ( .A0(cmd_il_valid), .A1(n222), .Z(cmd_il_data[43]));
Q_AN02 U1733 ( .A0(cmd_il_valid), .A1(n223), .Z(cmd_il_data[42]));
Q_AN02 U1734 ( .A0(cmd_il_valid), .A1(n224), .Z(cmd_il_data[41]));
Q_AN02 U1735 ( .A0(cmd_il_valid), .A1(n225), .Z(cmd_il_data[40]));
Q_AN02 U1736 ( .A0(cmd_il_valid), .A1(n226), .Z(cmd_il_data[39]));
Q_AN02 U1737 ( .A0(cmd_il_valid), .A1(n227), .Z(cmd_il_data[38]));
Q_AN02 U1738 ( .A0(cmd_il_valid), .A1(n228), .Z(cmd_il_data[37]));
Q_AN02 U1739 ( .A0(cmd_il_valid), .A1(n229), .Z(cmd_il_data[36]));
Q_AN02 U1740 ( .A0(cmd_il_valid), .A1(n230), .Z(cmd_il_data[35]));
Q_AN02 U1741 ( .A0(cmd_il_valid), .A1(n231), .Z(cmd_il_data[34]));
Q_AN02 U1742 ( .A0(cmd_il_valid), .A1(n232), .Z(cmd_il_data[33]));
Q_AN02 U1743 ( .A0(cmd_il_valid), .A1(n233), .Z(cmd_il_data[32]));
Q_AN02 U1744 ( .A0(cmd_il_valid), .A1(n234), .Z(cmd_il_data[31]));
Q_AN02 U1745 ( .A0(cmd_il_valid), .A1(n235), .Z(cmd_il_data[30]));
Q_AN02 U1746 ( .A0(cmd_il_valid), .A1(n236), .Z(cmd_il_data[29]));
Q_AN02 U1747 ( .A0(cmd_il_valid), .A1(n237), .Z(cmd_il_data[28]));
Q_AN02 U1748 ( .A0(cmd_il_valid), .A1(n238), .Z(cmd_il_data[27]));
Q_AN02 U1749 ( .A0(cmd_il_valid), .A1(n239), .Z(cmd_il_data[26]));
Q_AN02 U1750 ( .A0(cmd_il_valid), .A1(n240), .Z(cmd_il_data[25]));
Q_AN02 U1751 ( .A0(cmd_il_valid), .A1(n241), .Z(cmd_il_data[24]));
Q_AN02 U1752 ( .A0(cmd_il_valid), .A1(n242), .Z(cmd_il_data[23]));
Q_AN02 U1753 ( .A0(cmd_il_valid), .A1(n243), .Z(cmd_il_data[22]));
Q_AN02 U1754 ( .A0(cmd_il_valid), .A1(n244), .Z(cmd_il_data[21]));
Q_AN02 U1755 ( .A0(cmd_il_valid), .A1(n245), .Z(cmd_il_data[20]));
Q_AN02 U1756 ( .A0(cmd_il_valid), .A1(n246), .Z(cmd_il_data[19]));
Q_AN02 U1757 ( .A0(cmd_il_valid), .A1(n247), .Z(cmd_il_data[18]));
Q_AN02 U1758 ( .A0(cmd_il_valid), .A1(n248), .Z(cmd_il_data[17]));
Q_AN02 U1759 ( .A0(cmd_il_valid), .A1(n249), .Z(cmd_il_data[16]));
Q_AN02 U1760 ( .A0(cmd_il_valid), .A1(n250), .Z(cmd_il_data[15]));
Q_AN02 U1761 ( .A0(cmd_il_valid), .A1(n251), .Z(cmd_il_data[14]));
Q_AN02 U1762 ( .A0(cmd_il_valid), .A1(n252), .Z(cmd_il_data[13]));
Q_AN02 U1763 ( .A0(cmd_il_valid), .A1(n253), .Z(cmd_il_data[12]));
Q_AN02 U1764 ( .A0(cmd_il_valid), .A1(n254), .Z(cmd_il_data[11]));
Q_AN02 U1765 ( .A0(cmd_il_valid), .A1(n255), .Z(cmd_il_data[10]));
Q_AN02 U1766 ( .A0(cmd_il_valid), .A1(n256), .Z(cmd_il_data[9]));
Q_AN02 U1767 ( .A0(cmd_il_valid), .A1(n257), .Z(cmd_il_data[8]));
Q_AN02 U1768 ( .A0(cmd_il_valid), .A1(n258), .Z(cmd_il_data[7]));
Q_AN02 U1769 ( .A0(cmd_il_valid), .A1(n259), .Z(cmd_il_data[6]));
Q_AN02 U1770 ( .A0(cmd_il_valid), .A1(n260), .Z(cmd_il_data[5]));
Q_AN02 U1771 ( .A0(cmd_il_valid), .A1(n261), .Z(cmd_il_data[4]));
Q_AN02 U1772 ( .A0(cmd_il_valid), .A1(n262), .Z(cmd_il_data[3]));
Q_AN02 U1773 ( .A0(cmd_il_valid), .A1(n263), .Z(cmd_il_data[2]));
Q_AN02 U1774 ( .A0(cmd_il_valid), .A1(n264), .Z(cmd_il_data[1]));
Q_AN02 U1775 ( .A0(cmd_il_valid), .A1(n265), .Z(cmd_il_data[0]));
Q_XOR2 U1776 ( .A0(n4), .A1(n1201), .Z(n1200));
Q_AD01HF U1777 ( .A0(n5), .B0(n1203), .S(n1202), .CO(n1201));
Q_AD01HF U1778 ( .A0(n6), .B0(n7), .S(n1204), .CO(n1203));
Q_INV U1779 ( .A(hash_cmd_in[11]), .Z(hash_cmd_in[10]));
Q_MX02 U1780 ( .S(cmd_dgl_data_size[0]), .A0(n1205), .A1(n1929), .Z(cmd_dgl_data[287]));
Q_AN02 U1781 ( .A0(n1189), .A1(n1493), .Z(n1205));
Q_MX02 U1782 ( .S(cmd_dgl_data_size[0]), .A0(n1206), .A1(n1931), .Z(cmd_dgl_data[286]));
Q_AN02 U1783 ( .A0(n1189), .A1(n1495), .Z(n1206));
Q_MX02 U1784 ( .S(cmd_dgl_data_size[0]), .A0(n1207), .A1(n1933), .Z(cmd_dgl_data[285]));
Q_AN02 U1785 ( .A0(n1189), .A1(n1497), .Z(n1207));
Q_MX02 U1786 ( .S(cmd_dgl_data_size[0]), .A0(n1208), .A1(n1935), .Z(cmd_dgl_data[284]));
Q_AN02 U1787 ( .A0(n1189), .A1(n1499), .Z(n1208));
Q_MX02 U1788 ( .S(cmd_dgl_data_size[0]), .A0(n1209), .A1(n1937), .Z(cmd_dgl_data[283]));
Q_AN02 U1789 ( .A0(n1189), .A1(n1501), .Z(n1209));
Q_MX02 U1790 ( .S(cmd_dgl_data_size[0]), .A0(n1210), .A1(n1939), .Z(cmd_dgl_data[282]));
Q_AN02 U1791 ( .A0(n1189), .A1(n1503), .Z(n1210));
Q_MX02 U1792 ( .S(cmd_dgl_data_size[0]), .A0(n1211), .A1(n1941), .Z(cmd_dgl_data[281]));
Q_AN02 U1793 ( .A0(n1189), .A1(n1505), .Z(n1211));
Q_MX02 U1794 ( .S(cmd_dgl_data_size[0]), .A0(n1212), .A1(n1943), .Z(cmd_dgl_data[280]));
Q_AN02 U1795 ( .A0(n1189), .A1(n1507), .Z(n1212));
Q_MX02 U1796 ( .S(cmd_dgl_data_size[0]), .A0(n1213), .A1(n1493), .Z(cmd_dgl_data[279]));
Q_AN02 U1797 ( .A0(n1189), .A1(n1509), .Z(n1213));
Q_MX02 U1798 ( .S(cmd_dgl_data_size[0]), .A0(n1214), .A1(n1495), .Z(cmd_dgl_data[278]));
Q_AN02 U1799 ( .A0(n1189), .A1(n1511), .Z(n1214));
Q_MX02 U1800 ( .S(cmd_dgl_data_size[0]), .A0(n1215), .A1(n1497), .Z(cmd_dgl_data[277]));
Q_AN02 U1801 ( .A0(n1189), .A1(n1513), .Z(n1215));
Q_MX02 U1802 ( .S(cmd_dgl_data_size[0]), .A0(n1216), .A1(n1499), .Z(cmd_dgl_data[276]));
Q_AN02 U1803 ( .A0(n1189), .A1(n1515), .Z(n1216));
Q_MX02 U1804 ( .S(cmd_dgl_data_size[0]), .A0(n1217), .A1(n1501), .Z(cmd_dgl_data[275]));
Q_AN02 U1805 ( .A0(n1189), .A1(n1517), .Z(n1217));
Q_MX02 U1806 ( .S(cmd_dgl_data_size[0]), .A0(n1218), .A1(n1503), .Z(cmd_dgl_data[274]));
Q_AN02 U1807 ( .A0(n1189), .A1(n1519), .Z(n1218));
Q_MX02 U1808 ( .S(cmd_dgl_data_size[0]), .A0(n1219), .A1(n1505), .Z(cmd_dgl_data[273]));
Q_AN02 U1809 ( .A0(n1189), .A1(n1521), .Z(n1219));
Q_MX02 U1810 ( .S(cmd_dgl_data_size[0]), .A0(n1220), .A1(n1507), .Z(cmd_dgl_data[272]));
Q_AN02 U1811 ( .A0(n1189), .A1(n1523), .Z(n1220));
Q_MX02 U1812 ( .S(cmd_dgl_data_size[0]), .A0(n1221), .A1(n1509), .Z(cmd_dgl_data[271]));
Q_AN02 U1813 ( .A0(n1189), .A1(n1525), .Z(n1221));
Q_MX02 U1814 ( .S(cmd_dgl_data_size[0]), .A0(n1222), .A1(n1511), .Z(cmd_dgl_data[270]));
Q_AN02 U1815 ( .A0(n1189), .A1(n1527), .Z(n1222));
Q_MX02 U1816 ( .S(cmd_dgl_data_size[0]), .A0(n1223), .A1(n1513), .Z(cmd_dgl_data[269]));
Q_AN02 U1817 ( .A0(n1189), .A1(n1529), .Z(n1223));
Q_MX02 U1818 ( .S(cmd_dgl_data_size[0]), .A0(n1224), .A1(n1515), .Z(cmd_dgl_data[268]));
Q_AN02 U1819 ( .A0(n1189), .A1(n1531), .Z(n1224));
Q_MX02 U1820 ( .S(cmd_dgl_data_size[0]), .A0(n1225), .A1(n1517), .Z(cmd_dgl_data[267]));
Q_AN02 U1821 ( .A0(n1189), .A1(n1533), .Z(n1225));
Q_MX02 U1822 ( .S(cmd_dgl_data_size[0]), .A0(n1226), .A1(n1519), .Z(cmd_dgl_data[266]));
Q_AN02 U1823 ( .A0(n1189), .A1(n1535), .Z(n1226));
Q_MX02 U1824 ( .S(cmd_dgl_data_size[0]), .A0(n1227), .A1(n1521), .Z(cmd_dgl_data[265]));
Q_AN02 U1825 ( .A0(n1189), .A1(n1537), .Z(n1227));
Q_MX02 U1826 ( .S(cmd_dgl_data_size[0]), .A0(n1228), .A1(n1523), .Z(cmd_dgl_data[264]));
Q_AN02 U1827 ( .A0(n1189), .A1(n1539), .Z(n1228));
Q_MX02 U1828 ( .S(cmd_dgl_data_size[0]), .A0(n1229), .A1(n1525), .Z(cmd_dgl_data[263]));
Q_AN02 U1829 ( .A0(n1189), .A1(n1541), .Z(n1229));
Q_MX02 U1830 ( .S(cmd_dgl_data_size[0]), .A0(n1230), .A1(n1527), .Z(cmd_dgl_data[262]));
Q_AN02 U1831 ( .A0(n1189), .A1(n1543), .Z(n1230));
Q_MX02 U1832 ( .S(cmd_dgl_data_size[0]), .A0(n1231), .A1(n1529), .Z(cmd_dgl_data[261]));
Q_AN02 U1833 ( .A0(n1189), .A1(n1545), .Z(n1231));
Q_MX02 U1834 ( .S(cmd_dgl_data_size[0]), .A0(n1232), .A1(n1531), .Z(cmd_dgl_data[260]));
Q_AN02 U1835 ( .A0(n1189), .A1(n1547), .Z(n1232));
Q_MX02 U1836 ( .S(cmd_dgl_data_size[0]), .A0(n1233), .A1(n1533), .Z(cmd_dgl_data[259]));
Q_AN02 U1837 ( .A0(n1189), .A1(n1549), .Z(n1233));
Q_MX02 U1838 ( .S(cmd_dgl_data_size[0]), .A0(n1234), .A1(n1535), .Z(cmd_dgl_data[258]));
Q_AN02 U1839 ( .A0(n1189), .A1(n1551), .Z(n1234));
Q_MX02 U1840 ( .S(cmd_dgl_data_size[0]), .A0(n1235), .A1(n1537), .Z(cmd_dgl_data[257]));
Q_AN02 U1841 ( .A0(n1189), .A1(n1553), .Z(n1235));
Q_MX02 U1842 ( .S(cmd_dgl_data_size[0]), .A0(n1236), .A1(n1539), .Z(cmd_dgl_data[256]));
Q_AN02 U1843 ( .A0(n1189), .A1(n1555), .Z(n1236));
Q_MX02 U1844 ( .S(cmd_dgl_data_size[0]), .A0(n1237), .A1(n1541), .Z(cmd_dgl_data[255]));
Q_AN02 U1845 ( .A0(n1189), .A1(n1557), .Z(n1237));
Q_MX02 U1846 ( .S(cmd_dgl_data_size[0]), .A0(n1238), .A1(n1543), .Z(cmd_dgl_data[254]));
Q_AN02 U1847 ( .A0(n1189), .A1(n1559), .Z(n1238));
Q_MX02 U1848 ( .S(cmd_dgl_data_size[0]), .A0(n1239), .A1(n1545), .Z(cmd_dgl_data[253]));
Q_AN02 U1849 ( .A0(n1189), .A1(n1561), .Z(n1239));
Q_MX02 U1850 ( .S(cmd_dgl_data_size[0]), .A0(n1240), .A1(n1547), .Z(cmd_dgl_data[252]));
Q_AN02 U1851 ( .A0(n1189), .A1(n1563), .Z(n1240));
Q_MX02 U1852 ( .S(cmd_dgl_data_size[0]), .A0(n1241), .A1(n1549), .Z(cmd_dgl_data[251]));
Q_AN02 U1853 ( .A0(n1189), .A1(n1565), .Z(n1241));
Q_MX02 U1854 ( .S(cmd_dgl_data_size[0]), .A0(n1242), .A1(n1551), .Z(cmd_dgl_data[250]));
Q_AN02 U1855 ( .A0(n1189), .A1(n1567), .Z(n1242));
Q_MX02 U1856 ( .S(cmd_dgl_data_size[0]), .A0(n1243), .A1(n1553), .Z(cmd_dgl_data[249]));
Q_AN02 U1857 ( .A0(n1189), .A1(n1569), .Z(n1243));
Q_MX02 U1858 ( .S(cmd_dgl_data_size[0]), .A0(n1244), .A1(n1555), .Z(cmd_dgl_data[248]));
Q_AN02 U1859 ( .A0(n1189), .A1(n1571), .Z(n1244));
Q_MX02 U1860 ( .S(cmd_dgl_data_size[0]), .A0(n1245), .A1(n1557), .Z(cmd_dgl_data[247]));
Q_AN02 U1861 ( .A0(n1189), .A1(n1573), .Z(n1245));
Q_MX02 U1862 ( .S(cmd_dgl_data_size[0]), .A0(n1246), .A1(n1559), .Z(cmd_dgl_data[246]));
Q_AN02 U1863 ( .A0(n1189), .A1(n1575), .Z(n1246));
Q_MX02 U1864 ( .S(cmd_dgl_data_size[0]), .A0(n1247), .A1(n1561), .Z(cmd_dgl_data[245]));
Q_AN02 U1865 ( .A0(n1189), .A1(n1577), .Z(n1247));
Q_MX02 U1866 ( .S(cmd_dgl_data_size[0]), .A0(n1248), .A1(n1563), .Z(cmd_dgl_data[244]));
Q_AN02 U1867 ( .A0(n1189), .A1(n1579), .Z(n1248));
Q_MX02 U1868 ( .S(cmd_dgl_data_size[0]), .A0(n1249), .A1(n1565), .Z(cmd_dgl_data[243]));
Q_AN02 U1869 ( .A0(n1189), .A1(n1581), .Z(n1249));
Q_MX02 U1870 ( .S(cmd_dgl_data_size[0]), .A0(n1250), .A1(n1567), .Z(cmd_dgl_data[242]));
Q_AN02 U1871 ( .A0(n1189), .A1(n1583), .Z(n1250));
Q_MX02 U1872 ( .S(cmd_dgl_data_size[0]), .A0(n1251), .A1(n1569), .Z(cmd_dgl_data[241]));
Q_AN02 U1873 ( .A0(n1189), .A1(n1585), .Z(n1251));
Q_MX02 U1874 ( .S(cmd_dgl_data_size[0]), .A0(n1252), .A1(n1571), .Z(cmd_dgl_data[240]));
Q_AN02 U1875 ( .A0(n1189), .A1(n1587), .Z(n1252));
Q_MX02 U1876 ( .S(cmd_dgl_data_size[0]), .A0(n1253), .A1(n1573), .Z(cmd_dgl_data[239]));
Q_AN02 U1877 ( .A0(n1189), .A1(n1589), .Z(n1253));
Q_MX02 U1878 ( .S(cmd_dgl_data_size[0]), .A0(n1254), .A1(n1575), .Z(cmd_dgl_data[238]));
Q_AN02 U1879 ( .A0(n1189), .A1(n1591), .Z(n1254));
Q_MX02 U1880 ( .S(cmd_dgl_data_size[0]), .A0(n1255), .A1(n1577), .Z(cmd_dgl_data[237]));
Q_AN02 U1881 ( .A0(n1189), .A1(n1593), .Z(n1255));
Q_MX02 U1882 ( .S(cmd_dgl_data_size[0]), .A0(n1256), .A1(n1579), .Z(cmd_dgl_data[236]));
Q_AN02 U1883 ( .A0(n1189), .A1(n1595), .Z(n1256));
Q_MX02 U1884 ( .S(cmd_dgl_data_size[0]), .A0(n1257), .A1(n1581), .Z(cmd_dgl_data[235]));
Q_AN02 U1885 ( .A0(n1189), .A1(n1597), .Z(n1257));
Q_MX02 U1886 ( .S(cmd_dgl_data_size[0]), .A0(n1258), .A1(n1583), .Z(cmd_dgl_data[234]));
Q_AN02 U1887 ( .A0(n1189), .A1(n1599), .Z(n1258));
Q_MX02 U1888 ( .S(cmd_dgl_data_size[0]), .A0(n1259), .A1(n1585), .Z(cmd_dgl_data[233]));
Q_AN02 U1889 ( .A0(n1189), .A1(n1601), .Z(n1259));
Q_MX02 U1890 ( .S(cmd_dgl_data_size[0]), .A0(n1260), .A1(n1587), .Z(cmd_dgl_data[232]));
Q_AN02 U1891 ( .A0(n1189), .A1(n1603), .Z(n1260));
Q_MX02 U1892 ( .S(cmd_dgl_data_size[0]), .A0(n1261), .A1(n1589), .Z(cmd_dgl_data[231]));
Q_AN02 U1893 ( .A0(n1189), .A1(n1605), .Z(n1261));
Q_MX02 U1894 ( .S(cmd_dgl_data_size[0]), .A0(n1262), .A1(n1591), .Z(cmd_dgl_data[230]));
Q_AN02 U1895 ( .A0(n1189), .A1(n1607), .Z(n1262));
Q_MX02 U1896 ( .S(cmd_dgl_data_size[0]), .A0(n1263), .A1(n1593), .Z(cmd_dgl_data[229]));
Q_AN02 U1897 ( .A0(n1189), .A1(n1609), .Z(n1263));
Q_MX02 U1898 ( .S(cmd_dgl_data_size[0]), .A0(n1264), .A1(n1595), .Z(cmd_dgl_data[228]));
Q_AN02 U1899 ( .A0(n1189), .A1(n1611), .Z(n1264));
Q_MX02 U1900 ( .S(cmd_dgl_data_size[0]), .A0(n1265), .A1(n1597), .Z(cmd_dgl_data[227]));
Q_AN02 U1901 ( .A0(n1189), .A1(n1613), .Z(n1265));
Q_MX02 U1902 ( .S(cmd_dgl_data_size[0]), .A0(n1266), .A1(n1599), .Z(cmd_dgl_data[226]));
Q_AN02 U1903 ( .A0(n1189), .A1(n1615), .Z(n1266));
Q_MX02 U1904 ( .S(cmd_dgl_data_size[0]), .A0(n1267), .A1(n1601), .Z(cmd_dgl_data[225]));
Q_AN02 U1905 ( .A0(n1189), .A1(n1617), .Z(n1267));
Q_MX02 U1906 ( .S(cmd_dgl_data_size[0]), .A0(n1268), .A1(n1603), .Z(cmd_dgl_data[224]));
Q_AN02 U1907 ( .A0(n1189), .A1(n1619), .Z(n1268));
Q_MX02 U1908 ( .S(cmd_dgl_data_size[0]), .A0(n1269), .A1(n1605), .Z(cmd_dgl_data[223]));
Q_AN02 U1909 ( .A0(n1189), .A1(n1621), .Z(n1269));
Q_MX02 U1910 ( .S(cmd_dgl_data_size[0]), .A0(n1270), .A1(n1607), .Z(cmd_dgl_data[222]));
Q_AN02 U1911 ( .A0(n1189), .A1(n1623), .Z(n1270));
Q_MX02 U1912 ( .S(cmd_dgl_data_size[0]), .A0(n1271), .A1(n1609), .Z(cmd_dgl_data[221]));
Q_AN02 U1913 ( .A0(n1189), .A1(n1625), .Z(n1271));
Q_MX02 U1914 ( .S(cmd_dgl_data_size[0]), .A0(n1272), .A1(n1611), .Z(cmd_dgl_data[220]));
Q_AN02 U1915 ( .A0(n1189), .A1(n1627), .Z(n1272));
Q_MX02 U1916 ( .S(cmd_dgl_data_size[0]), .A0(n1273), .A1(n1613), .Z(cmd_dgl_data[219]));
Q_AN02 U1917 ( .A0(n1189), .A1(n1629), .Z(n1273));
Q_MX02 U1918 ( .S(cmd_dgl_data_size[0]), .A0(n1274), .A1(n1615), .Z(cmd_dgl_data[218]));
Q_AN02 U1919 ( .A0(n1189), .A1(n1631), .Z(n1274));
Q_MX02 U1920 ( .S(cmd_dgl_data_size[0]), .A0(n1275), .A1(n1617), .Z(cmd_dgl_data[217]));
Q_AN02 U1921 ( .A0(n1189), .A1(n1633), .Z(n1275));
Q_MX02 U1922 ( .S(cmd_dgl_data_size[0]), .A0(n1276), .A1(n1619), .Z(cmd_dgl_data[216]));
Q_AN02 U1923 ( .A0(n1189), .A1(n1635), .Z(n1276));
Q_MX02 U1924 ( .S(cmd_dgl_data_size[0]), .A0(n1277), .A1(n1621), .Z(cmd_dgl_data[215]));
Q_AN02 U1925 ( .A0(n1189), .A1(n1637), .Z(n1277));
Q_MX02 U1926 ( .S(cmd_dgl_data_size[0]), .A0(n1278), .A1(n1623), .Z(cmd_dgl_data[214]));
Q_AN02 U1927 ( .A0(n1189), .A1(n1639), .Z(n1278));
Q_MX02 U1928 ( .S(cmd_dgl_data_size[0]), .A0(n1279), .A1(n1625), .Z(cmd_dgl_data[213]));
Q_AN02 U1929 ( .A0(n1189), .A1(n1641), .Z(n1279));
Q_MX02 U1930 ( .S(cmd_dgl_data_size[0]), .A0(n1280), .A1(n1627), .Z(cmd_dgl_data[212]));
Q_AN02 U1931 ( .A0(n1189), .A1(n1643), .Z(n1280));
Q_MX02 U1932 ( .S(cmd_dgl_data_size[0]), .A0(n1281), .A1(n1629), .Z(cmd_dgl_data[211]));
Q_AN02 U1933 ( .A0(n1189), .A1(n1645), .Z(n1281));
Q_MX02 U1934 ( .S(cmd_dgl_data_size[0]), .A0(n1282), .A1(n1631), .Z(cmd_dgl_data[210]));
Q_AN02 U1935 ( .A0(n1189), .A1(n1647), .Z(n1282));
Q_MX02 U1936 ( .S(cmd_dgl_data_size[0]), .A0(n1283), .A1(n1633), .Z(cmd_dgl_data[209]));
Q_AN02 U1937 ( .A0(n1189), .A1(n1649), .Z(n1283));
Q_MX02 U1938 ( .S(cmd_dgl_data_size[0]), .A0(n1284), .A1(n1635), .Z(cmd_dgl_data[208]));
Q_AN02 U1939 ( .A0(n1189), .A1(n1651), .Z(n1284));
Q_MX02 U1940 ( .S(cmd_dgl_data_size[0]), .A0(n1285), .A1(n1637), .Z(cmd_dgl_data[207]));
Q_AN02 U1941 ( .A0(n1189), .A1(n1653), .Z(n1285));
Q_MX02 U1942 ( .S(cmd_dgl_data_size[0]), .A0(n1286), .A1(n1639), .Z(cmd_dgl_data[206]));
Q_AN02 U1943 ( .A0(n1189), .A1(n1655), .Z(n1286));
Q_MX02 U1944 ( .S(cmd_dgl_data_size[0]), .A0(n1287), .A1(n1641), .Z(cmd_dgl_data[205]));
Q_AN02 U1945 ( .A0(n1189), .A1(n1657), .Z(n1287));
Q_MX02 U1946 ( .S(cmd_dgl_data_size[0]), .A0(n1288), .A1(n1643), .Z(cmd_dgl_data[204]));
Q_AN02 U1947 ( .A0(n1189), .A1(n1659), .Z(n1288));
Q_MX02 U1948 ( .S(cmd_dgl_data_size[0]), .A0(n1289), .A1(n1645), .Z(cmd_dgl_data[203]));
Q_AN02 U1949 ( .A0(n1189), .A1(n1661), .Z(n1289));
Q_MX02 U1950 ( .S(cmd_dgl_data_size[0]), .A0(n1290), .A1(n1647), .Z(cmd_dgl_data[202]));
Q_AN02 U1951 ( .A0(n1189), .A1(n1663), .Z(n1290));
Q_MX02 U1952 ( .S(cmd_dgl_data_size[0]), .A0(n1291), .A1(n1649), .Z(cmd_dgl_data[201]));
Q_AN02 U1953 ( .A0(n1189), .A1(n1665), .Z(n1291));
Q_MX02 U1954 ( .S(cmd_dgl_data_size[0]), .A0(n1292), .A1(n1651), .Z(cmd_dgl_data[200]));
Q_AN02 U1955 ( .A0(n1189), .A1(n1667), .Z(n1292));
Q_MX02 U1956 ( .S(cmd_dgl_data_size[0]), .A0(n1293), .A1(n1653), .Z(cmd_dgl_data[199]));
Q_AN02 U1957 ( .A0(n1189), .A1(n1669), .Z(n1293));
Q_MX02 U1958 ( .S(cmd_dgl_data_size[0]), .A0(n1294), .A1(n1655), .Z(cmd_dgl_data[198]));
Q_AN02 U1959 ( .A0(n1189), .A1(n1671), .Z(n1294));
Q_MX02 U1960 ( .S(cmd_dgl_data_size[0]), .A0(n1295), .A1(n1657), .Z(cmd_dgl_data[197]));
Q_AN02 U1961 ( .A0(n1189), .A1(n1673), .Z(n1295));
Q_MX02 U1962 ( .S(cmd_dgl_data_size[0]), .A0(n1296), .A1(n1659), .Z(cmd_dgl_data[196]));
Q_AN02 U1963 ( .A0(n1189), .A1(n1675), .Z(n1296));
Q_MX02 U1964 ( .S(cmd_dgl_data_size[0]), .A0(n1297), .A1(n1661), .Z(cmd_dgl_data[195]));
Q_AN02 U1965 ( .A0(n1189), .A1(n1677), .Z(n1297));
Q_MX02 U1966 ( .S(cmd_dgl_data_size[0]), .A0(n1298), .A1(n1663), .Z(cmd_dgl_data[194]));
Q_AN02 U1967 ( .A0(n1189), .A1(n1679), .Z(n1298));
Q_MX02 U1968 ( .S(cmd_dgl_data_size[0]), .A0(n1299), .A1(n1665), .Z(cmd_dgl_data[193]));
Q_AN02 U1969 ( .A0(n1189), .A1(n1681), .Z(n1299));
Q_MX02 U1970 ( .S(cmd_dgl_data_size[0]), .A0(n1300), .A1(n1667), .Z(cmd_dgl_data[192]));
Q_AN02 U1971 ( .A0(n1189), .A1(n1683), .Z(n1300));
Q_MX02 U1972 ( .S(cmd_dgl_data_size[0]), .A0(n1301), .A1(n1669), .Z(cmd_dgl_data[191]));
Q_AN02 U1973 ( .A0(n1189), .A1(n1685), .Z(n1301));
Q_MX02 U1974 ( .S(cmd_dgl_data_size[0]), .A0(n1302), .A1(n1671), .Z(cmd_dgl_data[190]));
Q_AN02 U1975 ( .A0(n1189), .A1(n1687), .Z(n1302));
Q_MX02 U1976 ( .S(cmd_dgl_data_size[0]), .A0(n1303), .A1(n1673), .Z(cmd_dgl_data[189]));
Q_AN02 U1977 ( .A0(n1189), .A1(n1689), .Z(n1303));
Q_MX02 U1978 ( .S(cmd_dgl_data_size[0]), .A0(n1304), .A1(n1675), .Z(cmd_dgl_data[188]));
Q_AN02 U1979 ( .A0(n1189), .A1(n1691), .Z(n1304));
Q_MX02 U1980 ( .S(cmd_dgl_data_size[0]), .A0(n1305), .A1(n1677), .Z(cmd_dgl_data[187]));
Q_AN02 U1981 ( .A0(n1189), .A1(n1693), .Z(n1305));
Q_MX02 U1982 ( .S(cmd_dgl_data_size[0]), .A0(n1306), .A1(n1679), .Z(cmd_dgl_data[186]));
Q_AN02 U1983 ( .A0(n1189), .A1(n1695), .Z(n1306));
Q_MX02 U1984 ( .S(cmd_dgl_data_size[0]), .A0(n1307), .A1(n1681), .Z(cmd_dgl_data[185]));
Q_AN02 U1985 ( .A0(n1189), .A1(n1697), .Z(n1307));
Q_MX02 U1986 ( .S(cmd_dgl_data_size[0]), .A0(n1308), .A1(n1683), .Z(cmd_dgl_data[184]));
Q_AN02 U1987 ( .A0(n1189), .A1(n1699), .Z(n1308));
Q_MX02 U1988 ( .S(cmd_dgl_data_size[0]), .A0(n1309), .A1(n1685), .Z(cmd_dgl_data[183]));
Q_AN02 U1989 ( .A0(n1189), .A1(n1701), .Z(n1309));
Q_MX02 U1990 ( .S(cmd_dgl_data_size[0]), .A0(n1310), .A1(n1687), .Z(cmd_dgl_data[182]));
Q_AN02 U1991 ( .A0(n1189), .A1(n1703), .Z(n1310));
Q_MX02 U1992 ( .S(cmd_dgl_data_size[0]), .A0(n1311), .A1(n1689), .Z(cmd_dgl_data[181]));
Q_AN02 U1993 ( .A0(n1189), .A1(n1705), .Z(n1311));
Q_MX02 U1994 ( .S(cmd_dgl_data_size[0]), .A0(n1312), .A1(n1691), .Z(cmd_dgl_data[180]));
Q_AN02 U1995 ( .A0(n1189), .A1(n1707), .Z(n1312));
Q_MX02 U1996 ( .S(cmd_dgl_data_size[0]), .A0(n1313), .A1(n1693), .Z(cmd_dgl_data[179]));
Q_AN02 U1997 ( .A0(n1189), .A1(n1709), .Z(n1313));
Q_MX02 U1998 ( .S(cmd_dgl_data_size[0]), .A0(n1314), .A1(n1695), .Z(cmd_dgl_data[178]));
Q_AN02 U1999 ( .A0(n1189), .A1(n1711), .Z(n1314));
Q_MX02 U2000 ( .S(cmd_dgl_data_size[0]), .A0(n1315), .A1(n1697), .Z(cmd_dgl_data[177]));
Q_AN02 U2001 ( .A0(n1189), .A1(n1713), .Z(n1315));
Q_MX02 U2002 ( .S(cmd_dgl_data_size[0]), .A0(n1316), .A1(n1699), .Z(cmd_dgl_data[176]));
Q_AN02 U2003 ( .A0(n1189), .A1(n1715), .Z(n1316));
Q_MX02 U2004 ( .S(cmd_dgl_data_size[0]), .A0(n1317), .A1(n1701), .Z(cmd_dgl_data[175]));
Q_AN02 U2005 ( .A0(n1189), .A1(n1717), .Z(n1317));
Q_MX02 U2006 ( .S(cmd_dgl_data_size[0]), .A0(n1318), .A1(n1703), .Z(cmd_dgl_data[174]));
Q_AN02 U2007 ( .A0(n1189), .A1(n1719), .Z(n1318));
Q_MX02 U2008 ( .S(cmd_dgl_data_size[0]), .A0(n1319), .A1(n1705), .Z(cmd_dgl_data[173]));
Q_AN02 U2009 ( .A0(n1189), .A1(n1721), .Z(n1319));
Q_MX02 U2010 ( .S(cmd_dgl_data_size[0]), .A0(n1320), .A1(n1707), .Z(cmd_dgl_data[172]));
Q_AN02 U2011 ( .A0(n1189), .A1(n1723), .Z(n1320));
Q_MX02 U2012 ( .S(cmd_dgl_data_size[0]), .A0(n1321), .A1(n1709), .Z(cmd_dgl_data[171]));
Q_AN02 U2013 ( .A0(n1189), .A1(n1725), .Z(n1321));
Q_MX02 U2014 ( .S(cmd_dgl_data_size[0]), .A0(n1322), .A1(n1711), .Z(cmd_dgl_data[170]));
Q_AN02 U2015 ( .A0(n1189), .A1(n1727), .Z(n1322));
Q_MX02 U2016 ( .S(cmd_dgl_data_size[0]), .A0(n1323), .A1(n1713), .Z(cmd_dgl_data[169]));
Q_AN02 U2017 ( .A0(n1189), .A1(n1729), .Z(n1323));
Q_MX02 U2018 ( .S(cmd_dgl_data_size[0]), .A0(n1324), .A1(n1715), .Z(cmd_dgl_data[168]));
Q_AN02 U2019 ( .A0(n1189), .A1(n1731), .Z(n1324));
Q_MX02 U2020 ( .S(cmd_dgl_data_size[0]), .A0(n1325), .A1(n1717), .Z(cmd_dgl_data[167]));
Q_AN02 U2021 ( .A0(n1189), .A1(n1733), .Z(n1325));
Q_MX02 U2022 ( .S(cmd_dgl_data_size[0]), .A0(n1326), .A1(n1719), .Z(cmd_dgl_data[166]));
Q_AN02 U2023 ( .A0(n1189), .A1(n1735), .Z(n1326));
Q_MX02 U2024 ( .S(cmd_dgl_data_size[0]), .A0(n1327), .A1(n1721), .Z(cmd_dgl_data[165]));
Q_AN02 U2025 ( .A0(n1189), .A1(n1737), .Z(n1327));
Q_MX02 U2026 ( .S(cmd_dgl_data_size[0]), .A0(n1328), .A1(n1723), .Z(cmd_dgl_data[164]));
Q_AN02 U2027 ( .A0(n1189), .A1(n1739), .Z(n1328));
Q_MX02 U2028 ( .S(cmd_dgl_data_size[0]), .A0(n1329), .A1(n1725), .Z(cmd_dgl_data[163]));
Q_AN02 U2029 ( .A0(n1189), .A1(n1741), .Z(n1329));
Q_MX02 U2030 ( .S(cmd_dgl_data_size[0]), .A0(n1330), .A1(n1727), .Z(cmd_dgl_data[162]));
Q_AN02 U2031 ( .A0(n1189), .A1(n1743), .Z(n1330));
Q_MX02 U2032 ( .S(cmd_dgl_data_size[0]), .A0(n1331), .A1(n1729), .Z(cmd_dgl_data[161]));
Q_AN02 U2033 ( .A0(n1189), .A1(n1745), .Z(n1331));
Q_MX02 U2034 ( .S(cmd_dgl_data_size[0]), .A0(n1332), .A1(n1731), .Z(cmd_dgl_data[160]));
Q_AN02 U2035 ( .A0(n1189), .A1(n1747), .Z(n1332));
Q_MX02 U2036 ( .S(cmd_dgl_data_size[0]), .A0(n1333), .A1(n1733), .Z(cmd_dgl_data[159]));
Q_AN02 U2037 ( .A0(n1189), .A1(n1749), .Z(n1333));
Q_MX02 U2038 ( .S(cmd_dgl_data_size[0]), .A0(n1334), .A1(n1735), .Z(cmd_dgl_data[158]));
Q_AN02 U2039 ( .A0(n1189), .A1(n1751), .Z(n1334));
Q_MX02 U2040 ( .S(cmd_dgl_data_size[0]), .A0(n1335), .A1(n1737), .Z(cmd_dgl_data[157]));
Q_AN02 U2041 ( .A0(n1189), .A1(n1753), .Z(n1335));
Q_MX02 U2042 ( .S(cmd_dgl_data_size[0]), .A0(n1336), .A1(n1739), .Z(cmd_dgl_data[156]));
Q_AN02 U2043 ( .A0(n1189), .A1(n1755), .Z(n1336));
Q_MX02 U2044 ( .S(cmd_dgl_data_size[0]), .A0(n1337), .A1(n1741), .Z(cmd_dgl_data[155]));
Q_AN02 U2045 ( .A0(n1189), .A1(n1757), .Z(n1337));
Q_MX02 U2046 ( .S(cmd_dgl_data_size[0]), .A0(n1338), .A1(n1743), .Z(cmd_dgl_data[154]));
Q_AN02 U2047 ( .A0(n1189), .A1(n1759), .Z(n1338));
Q_MX02 U2048 ( .S(cmd_dgl_data_size[0]), .A0(n1339), .A1(n1745), .Z(cmd_dgl_data[153]));
Q_AN02 U2049 ( .A0(n1189), .A1(n1761), .Z(n1339));
Q_MX02 U2050 ( .S(cmd_dgl_data_size[0]), .A0(n1340), .A1(n1747), .Z(cmd_dgl_data[152]));
Q_AN02 U2051 ( .A0(n1189), .A1(n1763), .Z(n1340));
Q_MX02 U2052 ( .S(cmd_dgl_data_size[0]), .A0(n1341), .A1(n1749), .Z(cmd_dgl_data[151]));
Q_AN02 U2053 ( .A0(n1189), .A1(n1765), .Z(n1341));
Q_MX02 U2054 ( .S(cmd_dgl_data_size[0]), .A0(n1342), .A1(n1751), .Z(cmd_dgl_data[150]));
Q_AN02 U2055 ( .A0(n1189), .A1(n1767), .Z(n1342));
Q_MX02 U2056 ( .S(cmd_dgl_data_size[0]), .A0(n1343), .A1(n1753), .Z(cmd_dgl_data[149]));
Q_AN02 U2057 ( .A0(n1189), .A1(n1769), .Z(n1343));
Q_MX02 U2058 ( .S(cmd_dgl_data_size[0]), .A0(n1344), .A1(n1755), .Z(cmd_dgl_data[148]));
Q_AN02 U2059 ( .A0(n1189), .A1(n1771), .Z(n1344));
Q_MX02 U2060 ( .S(cmd_dgl_data_size[0]), .A0(n1345), .A1(n1757), .Z(cmd_dgl_data[147]));
Q_AN02 U2061 ( .A0(n1189), .A1(n1773), .Z(n1345));
Q_MX02 U2062 ( .S(cmd_dgl_data_size[0]), .A0(n1346), .A1(n1759), .Z(cmd_dgl_data[146]));
Q_AN02 U2063 ( .A0(n1189), .A1(n1775), .Z(n1346));
Q_MX02 U2064 ( .S(cmd_dgl_data_size[0]), .A0(n1347), .A1(n1761), .Z(cmd_dgl_data[145]));
Q_AN02 U2065 ( .A0(n1189), .A1(n1777), .Z(n1347));
Q_MX02 U2066 ( .S(cmd_dgl_data_size[0]), .A0(n1348), .A1(n1763), .Z(cmd_dgl_data[144]));
Q_AN02 U2067 ( .A0(n1189), .A1(n1780), .Z(n1348));
Q_MX02 U2068 ( .S(cmd_dgl_data_size[0]), .A0(n1349), .A1(n1765), .Z(cmd_dgl_data[143]));
Q_AN02 U2069 ( .A0(n1189), .A1(n1783), .Z(n1349));
Q_MX02 U2070 ( .S(cmd_dgl_data_size[0]), .A0(n1350), .A1(n1767), .Z(cmd_dgl_data[142]));
Q_AN02 U2071 ( .A0(n1189), .A1(n1785), .Z(n1350));
Q_MX02 U2072 ( .S(cmd_dgl_data_size[0]), .A0(n1351), .A1(n1769), .Z(cmd_dgl_data[141]));
Q_AN02 U2073 ( .A0(n1189), .A1(n1787), .Z(n1351));
Q_MX02 U2074 ( .S(cmd_dgl_data_size[0]), .A0(n1352), .A1(n1771), .Z(cmd_dgl_data[140]));
Q_AN02 U2075 ( .A0(n1189), .A1(n1789), .Z(n1352));
Q_MX02 U2076 ( .S(cmd_dgl_data_size[0]), .A0(n1353), .A1(n1773), .Z(cmd_dgl_data[139]));
Q_AN02 U2077 ( .A0(n1189), .A1(n1791), .Z(n1353));
Q_MX02 U2078 ( .S(cmd_dgl_data_size[0]), .A0(n1354), .A1(n1775), .Z(cmd_dgl_data[138]));
Q_AN02 U2079 ( .A0(n1189), .A1(n1793), .Z(n1354));
Q_MX02 U2080 ( .S(cmd_dgl_data_size[0]), .A0(n1355), .A1(n1777), .Z(cmd_dgl_data[137]));
Q_AN02 U2081 ( .A0(n1189), .A1(n1795), .Z(n1355));
Q_MX02 U2082 ( .S(cmd_dgl_data_size[0]), .A0(n1356), .A1(n1780), .Z(cmd_dgl_data[136]));
Q_AN02 U2083 ( .A0(n1189), .A1(n1797), .Z(n1356));
Q_MX02 U2084 ( .S(cmd_dgl_data_size[0]), .A0(n1357), .A1(n1783), .Z(cmd_dgl_data[135]));
Q_AN02 U2085 ( .A0(n1189), .A1(n1799), .Z(n1357));
Q_MX02 U2086 ( .S(cmd_dgl_data_size[0]), .A0(n1358), .A1(n1785), .Z(cmd_dgl_data[134]));
Q_AN02 U2087 ( .A0(n1189), .A1(n1800), .Z(n1358));
Q_MX02 U2088 ( .S(cmd_dgl_data_size[0]), .A0(n1359), .A1(n1787), .Z(cmd_dgl_data[133]));
Q_AN02 U2089 ( .A0(n1189), .A1(n1801), .Z(n1359));
Q_MX02 U2090 ( .S(cmd_dgl_data_size[0]), .A0(n1360), .A1(n1789), .Z(cmd_dgl_data[132]));
Q_AN02 U2091 ( .A0(n1189), .A1(n1802), .Z(n1360));
Q_MX02 U2092 ( .S(cmd_dgl_data_size[0]), .A0(n1361), .A1(n1791), .Z(cmd_dgl_data[131]));
Q_AN02 U2093 ( .A0(n1189), .A1(n1803), .Z(n1361));
Q_MX02 U2094 ( .S(cmd_dgl_data_size[0]), .A0(n1362), .A1(n1793), .Z(cmd_dgl_data[130]));
Q_AN02 U2095 ( .A0(n1189), .A1(n1804), .Z(n1362));
Q_MX02 U2096 ( .S(cmd_dgl_data_size[0]), .A0(n1363), .A1(n1795), .Z(cmd_dgl_data[129]));
Q_AN02 U2097 ( .A0(n1189), .A1(n1805), .Z(n1363));
Q_MX02 U2098 ( .S(cmd_dgl_data_size[0]), .A0(n1364), .A1(n1797), .Z(cmd_dgl_data[128]));
Q_AN02 U2099 ( .A0(n1189), .A1(n1806), .Z(n1364));
Q_MX02 U2100 ( .S(cmd_dgl_data_size[0]), .A0(n1365), .A1(n1799), .Z(cmd_dgl_data[127]));
Q_AN02 U2101 ( .A0(n1189), .A1(n1807), .Z(n1365));
Q_MX02 U2102 ( .S(cmd_dgl_data_size[0]), .A0(n1366), .A1(n1800), .Z(cmd_dgl_data[126]));
Q_AN02 U2103 ( .A0(n1189), .A1(n1808), .Z(n1366));
Q_MX02 U2104 ( .S(cmd_dgl_data_size[0]), .A0(n1367), .A1(n1801), .Z(cmd_dgl_data[125]));
Q_AN02 U2105 ( .A0(n1189), .A1(n1809), .Z(n1367));
Q_MX02 U2106 ( .S(cmd_dgl_data_size[0]), .A0(n1368), .A1(n1802), .Z(cmd_dgl_data[124]));
Q_AN02 U2107 ( .A0(n1189), .A1(n1810), .Z(n1368));
Q_MX02 U2108 ( .S(cmd_dgl_data_size[0]), .A0(n1369), .A1(n1803), .Z(cmd_dgl_data[123]));
Q_AN02 U2109 ( .A0(n1189), .A1(n1811), .Z(n1369));
Q_MX02 U2110 ( .S(cmd_dgl_data_size[0]), .A0(n1370), .A1(n1804), .Z(cmd_dgl_data[122]));
Q_AN02 U2111 ( .A0(n1189), .A1(n1812), .Z(n1370));
Q_MX02 U2112 ( .S(cmd_dgl_data_size[0]), .A0(n1371), .A1(n1805), .Z(cmd_dgl_data[121]));
Q_AN02 U2113 ( .A0(n1189), .A1(n1813), .Z(n1371));
Q_MX02 U2114 ( .S(cmd_dgl_data_size[0]), .A0(n1372), .A1(n1806), .Z(cmd_dgl_data[120]));
Q_AN02 U2115 ( .A0(n1189), .A1(n1814), .Z(n1372));
Q_MX02 U2116 ( .S(cmd_dgl_data_size[0]), .A0(n1373), .A1(n1807), .Z(cmd_dgl_data[119]));
Q_AN02 U2117 ( .A0(n1189), .A1(n1815), .Z(n1373));
Q_MX02 U2118 ( .S(cmd_dgl_data_size[0]), .A0(n1374), .A1(n1808), .Z(cmd_dgl_data[118]));
Q_AN02 U2119 ( .A0(n1189), .A1(n1816), .Z(n1374));
Q_MX02 U2120 ( .S(cmd_dgl_data_size[0]), .A0(n1375), .A1(n1809), .Z(cmd_dgl_data[117]));
Q_AN02 U2121 ( .A0(n1189), .A1(n1817), .Z(n1375));
Q_MX02 U2122 ( .S(cmd_dgl_data_size[0]), .A0(n1376), .A1(n1810), .Z(cmd_dgl_data[116]));
Q_AN02 U2123 ( .A0(n1189), .A1(n1818), .Z(n1376));
Q_MX02 U2124 ( .S(cmd_dgl_data_size[0]), .A0(n1377), .A1(n1811), .Z(cmd_dgl_data[115]));
Q_AN02 U2125 ( .A0(n1189), .A1(n1819), .Z(n1377));
Q_MX02 U2126 ( .S(cmd_dgl_data_size[0]), .A0(n1378), .A1(n1812), .Z(cmd_dgl_data[114]));
Q_AN02 U2127 ( .A0(n1189), .A1(n1820), .Z(n1378));
Q_MX02 U2128 ( .S(cmd_dgl_data_size[0]), .A0(n1379), .A1(n1813), .Z(cmd_dgl_data[113]));
Q_AN02 U2129 ( .A0(n1189), .A1(n1821), .Z(n1379));
Q_MX02 U2130 ( .S(cmd_dgl_data_size[0]), .A0(n1380), .A1(n1814), .Z(cmd_dgl_data[112]));
Q_AN02 U2131 ( .A0(n1189), .A1(n1822), .Z(n1380));
Q_MX02 U2132 ( .S(cmd_dgl_data_size[0]), .A0(n1381), .A1(n1815), .Z(cmd_dgl_data[111]));
Q_AN02 U2133 ( .A0(n1189), .A1(n1823), .Z(n1381));
Q_MX02 U2134 ( .S(cmd_dgl_data_size[0]), .A0(n1382), .A1(n1816), .Z(cmd_dgl_data[110]));
Q_AN02 U2135 ( .A0(n1189), .A1(n1824), .Z(n1382));
Q_MX02 U2136 ( .S(cmd_dgl_data_size[0]), .A0(n1383), .A1(n1817), .Z(cmd_dgl_data[109]));
Q_AN02 U2137 ( .A0(n1189), .A1(n1825), .Z(n1383));
Q_MX02 U2138 ( .S(cmd_dgl_data_size[0]), .A0(n1384), .A1(n1818), .Z(cmd_dgl_data[108]));
Q_AN02 U2139 ( .A0(n1189), .A1(n1826), .Z(n1384));
Q_MX02 U2140 ( .S(cmd_dgl_data_size[0]), .A0(n1385), .A1(n1819), .Z(cmd_dgl_data[107]));
Q_AN02 U2141 ( .A0(n1189), .A1(n1827), .Z(n1385));
Q_MX02 U2142 ( .S(cmd_dgl_data_size[0]), .A0(n1386), .A1(n1820), .Z(cmd_dgl_data[106]));
Q_AN02 U2143 ( .A0(n1189), .A1(n1828), .Z(n1386));
Q_MX02 U2144 ( .S(cmd_dgl_data_size[0]), .A0(n1387), .A1(n1821), .Z(cmd_dgl_data[105]));
Q_AN02 U2145 ( .A0(n1189), .A1(n1829), .Z(n1387));
Q_MX02 U2146 ( .S(cmd_dgl_data_size[0]), .A0(n1388), .A1(n1822), .Z(cmd_dgl_data[104]));
Q_AN02 U2147 ( .A0(n1189), .A1(n1830), .Z(n1388));
Q_MX02 U2148 ( .S(cmd_dgl_data_size[0]), .A0(n1389), .A1(n1823), .Z(cmd_dgl_data[103]));
Q_AN02 U2149 ( .A0(n1189), .A1(n1831), .Z(n1389));
Q_MX02 U2150 ( .S(cmd_dgl_data_size[0]), .A0(n1390), .A1(n1824), .Z(cmd_dgl_data[102]));
Q_AN02 U2151 ( .A0(n1189), .A1(n1832), .Z(n1390));
Q_MX02 U2152 ( .S(cmd_dgl_data_size[0]), .A0(n1391), .A1(n1825), .Z(cmd_dgl_data[101]));
Q_AN02 U2153 ( .A0(n1189), .A1(n1833), .Z(n1391));
Q_MX02 U2154 ( .S(cmd_dgl_data_size[0]), .A0(n1392), .A1(n1826), .Z(cmd_dgl_data[100]));
Q_AN02 U2155 ( .A0(n1189), .A1(n1834), .Z(n1392));
Q_MX02 U2156 ( .S(cmd_dgl_data_size[0]), .A0(n1393), .A1(n1827), .Z(cmd_dgl_data[99]));
Q_AN02 U2157 ( .A0(n1189), .A1(n1835), .Z(n1393));
Q_MX02 U2158 ( .S(cmd_dgl_data_size[0]), .A0(n1394), .A1(n1828), .Z(cmd_dgl_data[98]));
Q_AN02 U2159 ( .A0(n1189), .A1(n1836), .Z(n1394));
Q_MX02 U2160 ( .S(cmd_dgl_data_size[0]), .A0(n1395), .A1(n1829), .Z(cmd_dgl_data[97]));
Q_AN02 U2161 ( .A0(n1189), .A1(n1837), .Z(n1395));
Q_MX02 U2162 ( .S(cmd_dgl_data_size[0]), .A0(n1396), .A1(n1830), .Z(cmd_dgl_data[96]));
Q_AN02 U2163 ( .A0(n1189), .A1(n1838), .Z(n1396));
Q_MX02 U2164 ( .S(cmd_dgl_data_size[0]), .A0(n1397), .A1(n1831), .Z(cmd_dgl_data[95]));
Q_AN02 U2165 ( .A0(n1189), .A1(n1839), .Z(n1397));
Q_MX02 U2166 ( .S(cmd_dgl_data_size[0]), .A0(n1398), .A1(n1832), .Z(cmd_dgl_data[94]));
Q_AN02 U2167 ( .A0(n1189), .A1(n1840), .Z(n1398));
Q_MX02 U2168 ( .S(cmd_dgl_data_size[0]), .A0(n1399), .A1(n1833), .Z(cmd_dgl_data[93]));
Q_AN02 U2169 ( .A0(n1189), .A1(n1841), .Z(n1399));
Q_MX02 U2170 ( .S(cmd_dgl_data_size[0]), .A0(n1400), .A1(n1834), .Z(cmd_dgl_data[92]));
Q_AN02 U2171 ( .A0(n1189), .A1(n1842), .Z(n1400));
Q_MX02 U2172 ( .S(cmd_dgl_data_size[0]), .A0(n1401), .A1(n1835), .Z(cmd_dgl_data[91]));
Q_AN02 U2173 ( .A0(n1189), .A1(n1843), .Z(n1401));
Q_MX02 U2174 ( .S(cmd_dgl_data_size[0]), .A0(n1402), .A1(n1836), .Z(cmd_dgl_data[90]));
Q_AN02 U2175 ( .A0(n1189), .A1(n1844), .Z(n1402));
Q_MX02 U2176 ( .S(cmd_dgl_data_size[0]), .A0(n1403), .A1(n1837), .Z(cmd_dgl_data[89]));
Q_AN02 U2177 ( .A0(n1189), .A1(n1845), .Z(n1403));
Q_MX02 U2178 ( .S(cmd_dgl_data_size[0]), .A0(n1404), .A1(n1838), .Z(cmd_dgl_data[88]));
Q_AN02 U2179 ( .A0(n1189), .A1(n1846), .Z(n1404));
Q_MX02 U2180 ( .S(cmd_dgl_data_size[0]), .A0(n1405), .A1(n1839), .Z(cmd_dgl_data[87]));
Q_AN02 U2181 ( .A0(n1189), .A1(n1847), .Z(n1405));
Q_MX02 U2182 ( .S(cmd_dgl_data_size[0]), .A0(n1406), .A1(n1840), .Z(cmd_dgl_data[86]));
Q_AN02 U2183 ( .A0(n1189), .A1(n1848), .Z(n1406));
Q_MX02 U2184 ( .S(cmd_dgl_data_size[0]), .A0(n1407), .A1(n1841), .Z(cmd_dgl_data[85]));
Q_AN02 U2185 ( .A0(n1189), .A1(n1849), .Z(n1407));
Q_MX02 U2186 ( .S(cmd_dgl_data_size[0]), .A0(n1408), .A1(n1842), .Z(cmd_dgl_data[84]));
Q_AN02 U2187 ( .A0(n1189), .A1(n1850), .Z(n1408));
Q_MX02 U2188 ( .S(cmd_dgl_data_size[0]), .A0(n1409), .A1(n1843), .Z(cmd_dgl_data[83]));
Q_AN02 U2189 ( .A0(n1189), .A1(n1851), .Z(n1409));
Q_MX02 U2190 ( .S(cmd_dgl_data_size[0]), .A0(n1410), .A1(n1844), .Z(cmd_dgl_data[82]));
Q_AN02 U2191 ( .A0(n1189), .A1(n1852), .Z(n1410));
Q_MX02 U2192 ( .S(cmd_dgl_data_size[0]), .A0(n1411), .A1(n1845), .Z(cmd_dgl_data[81]));
Q_AN02 U2193 ( .A0(n1189), .A1(n1853), .Z(n1411));
Q_MX02 U2194 ( .S(cmd_dgl_data_size[0]), .A0(n1412), .A1(n1846), .Z(cmd_dgl_data[80]));
Q_AN02 U2195 ( .A0(n1189), .A1(n1854), .Z(n1412));
Q_MX02 U2196 ( .S(cmd_dgl_data_size[0]), .A0(n1413), .A1(n1847), .Z(cmd_dgl_data[79]));
Q_AN02 U2197 ( .A0(n1189), .A1(n1855), .Z(n1413));
Q_MX02 U2198 ( .S(cmd_dgl_data_size[0]), .A0(n1414), .A1(n1848), .Z(cmd_dgl_data[78]));
Q_AN02 U2199 ( .A0(n1189), .A1(n1856), .Z(n1414));
Q_MX02 U2200 ( .S(cmd_dgl_data_size[0]), .A0(n1415), .A1(n1849), .Z(cmd_dgl_data[77]));
Q_AN02 U2201 ( .A0(n1189), .A1(n1857), .Z(n1415));
Q_MX02 U2202 ( .S(cmd_dgl_data_size[0]), .A0(n1416), .A1(n1850), .Z(cmd_dgl_data[76]));
Q_AN02 U2203 ( .A0(n1189), .A1(n1858), .Z(n1416));
Q_MX02 U2204 ( .S(cmd_dgl_data_size[0]), .A0(n1417), .A1(n1851), .Z(cmd_dgl_data[75]));
Q_AN02 U2205 ( .A0(n1189), .A1(n1859), .Z(n1417));
Q_MX02 U2206 ( .S(cmd_dgl_data_size[0]), .A0(n1418), .A1(n1852), .Z(cmd_dgl_data[74]));
Q_AN02 U2207 ( .A0(n1189), .A1(n1860), .Z(n1418));
Q_MX02 U2208 ( .S(cmd_dgl_data_size[0]), .A0(n1419), .A1(n1853), .Z(cmd_dgl_data[73]));
Q_AN02 U2209 ( .A0(n1189), .A1(n1861), .Z(n1419));
Q_MX02 U2210 ( .S(cmd_dgl_data_size[0]), .A0(n1420), .A1(n1854), .Z(cmd_dgl_data[72]));
Q_AN02 U2211 ( .A0(n1189), .A1(n1862), .Z(n1420));
Q_MX02 U2212 ( .S(cmd_dgl_data_size[0]), .A0(n1421), .A1(n1855), .Z(cmd_dgl_data[71]));
Q_AN02 U2213 ( .A0(n1189), .A1(n1863), .Z(n1421));
Q_MX02 U2214 ( .S(cmd_dgl_data_size[0]), .A0(n1422), .A1(n1856), .Z(cmd_dgl_data[70]));
Q_AN02 U2215 ( .A0(n1189), .A1(n1864), .Z(n1422));
Q_MX02 U2216 ( .S(cmd_dgl_data_size[0]), .A0(n1423), .A1(n1857), .Z(cmd_dgl_data[69]));
Q_AN02 U2217 ( .A0(n1189), .A1(n1865), .Z(n1423));
Q_MX02 U2218 ( .S(cmd_dgl_data_size[0]), .A0(n1424), .A1(n1858), .Z(cmd_dgl_data[68]));
Q_AN02 U2219 ( .A0(n1189), .A1(n1866), .Z(n1424));
Q_MX02 U2220 ( .S(cmd_dgl_data_size[0]), .A0(n1425), .A1(n1859), .Z(cmd_dgl_data[67]));
Q_AN02 U2221 ( .A0(n1189), .A1(n1867), .Z(n1425));
Q_MX02 U2222 ( .S(cmd_dgl_data_size[0]), .A0(n1426), .A1(n1860), .Z(cmd_dgl_data[66]));
Q_AN02 U2223 ( .A0(n1189), .A1(n1868), .Z(n1426));
Q_MX02 U2224 ( .S(cmd_dgl_data_size[0]), .A0(n1427), .A1(n1861), .Z(cmd_dgl_data[65]));
Q_AN02 U2225 ( .A0(n1189), .A1(n1869), .Z(n1427));
Q_MX02 U2226 ( .S(cmd_dgl_data_size[0]), .A0(n1428), .A1(n1862), .Z(cmd_dgl_data[64]));
Q_AN02 U2227 ( .A0(n1189), .A1(n1870), .Z(n1428));
Q_MX02 U2228 ( .S(cmd_dgl_data_size[0]), .A0(n1429), .A1(n1863), .Z(cmd_dgl_data[63]));
Q_AN02 U2229 ( .A0(n1189), .A1(n1871), .Z(n1429));
Q_MX02 U2230 ( .S(cmd_dgl_data_size[0]), .A0(n1430), .A1(n1864), .Z(cmd_dgl_data[62]));
Q_AN02 U2231 ( .A0(n1189), .A1(n1872), .Z(n1430));
Q_MX02 U2232 ( .S(cmd_dgl_data_size[0]), .A0(n1431), .A1(n1865), .Z(cmd_dgl_data[61]));
Q_AN02 U2233 ( .A0(n1189), .A1(n1873), .Z(n1431));
Q_MX02 U2234 ( .S(cmd_dgl_data_size[0]), .A0(n1432), .A1(n1866), .Z(cmd_dgl_data[60]));
Q_AN02 U2235 ( .A0(n1189), .A1(n1874), .Z(n1432));
Q_MX02 U2236 ( .S(cmd_dgl_data_size[0]), .A0(n1433), .A1(n1867), .Z(cmd_dgl_data[59]));
Q_AN02 U2237 ( .A0(n1189), .A1(n1875), .Z(n1433));
Q_MX02 U2238 ( .S(cmd_dgl_data_size[0]), .A0(n1434), .A1(n1868), .Z(cmd_dgl_data[58]));
Q_AN02 U2239 ( .A0(n1189), .A1(n1876), .Z(n1434));
Q_MX02 U2240 ( .S(cmd_dgl_data_size[0]), .A0(n1435), .A1(n1869), .Z(cmd_dgl_data[57]));
Q_AN02 U2241 ( .A0(n1189), .A1(n1877), .Z(n1435));
Q_MX02 U2242 ( .S(cmd_dgl_data_size[0]), .A0(n1436), .A1(n1870), .Z(cmd_dgl_data[56]));
Q_AN02 U2243 ( .A0(n1189), .A1(n1878), .Z(n1436));
Q_MX02 U2244 ( .S(cmd_dgl_data_size[0]), .A0(n1437), .A1(n1871), .Z(cmd_dgl_data[55]));
Q_AN02 U2245 ( .A0(n1189), .A1(n1879), .Z(n1437));
Q_MX02 U2246 ( .S(cmd_dgl_data_size[0]), .A0(n1438), .A1(n1872), .Z(cmd_dgl_data[54]));
Q_AN02 U2247 ( .A0(n1189), .A1(n1880), .Z(n1438));
Q_MX02 U2248 ( .S(cmd_dgl_data_size[0]), .A0(n1439), .A1(n1873), .Z(cmd_dgl_data[53]));
Q_AN02 U2249 ( .A0(n1189), .A1(n1881), .Z(n1439));
Q_MX02 U2250 ( .S(cmd_dgl_data_size[0]), .A0(n1440), .A1(n1874), .Z(cmd_dgl_data[52]));
Q_AN02 U2251 ( .A0(n1189), .A1(n1882), .Z(n1440));
Q_MX02 U2252 ( .S(cmd_dgl_data_size[0]), .A0(n1441), .A1(n1875), .Z(cmd_dgl_data[51]));
Q_AN02 U2253 ( .A0(n1189), .A1(n1883), .Z(n1441));
Q_MX02 U2254 ( .S(cmd_dgl_data_size[0]), .A0(n1442), .A1(n1876), .Z(cmd_dgl_data[50]));
Q_AN02 U2255 ( .A0(n1189), .A1(n1884), .Z(n1442));
Q_MX02 U2256 ( .S(cmd_dgl_data_size[0]), .A0(n1443), .A1(n1877), .Z(cmd_dgl_data[49]));
Q_AN02 U2257 ( .A0(n1189), .A1(n1885), .Z(n1443));
Q_MX02 U2258 ( .S(cmd_dgl_data_size[0]), .A0(n1444), .A1(n1878), .Z(cmd_dgl_data[48]));
Q_AN02 U2259 ( .A0(n1189), .A1(n1886), .Z(n1444));
Q_MX02 U2260 ( .S(cmd_dgl_data_size[0]), .A0(n1445), .A1(n1879), .Z(cmd_dgl_data[47]));
Q_AN02 U2261 ( .A0(n1189), .A1(n1887), .Z(n1445));
Q_MX02 U2262 ( .S(cmd_dgl_data_size[0]), .A0(n1446), .A1(n1880), .Z(cmd_dgl_data[46]));
Q_AN02 U2263 ( .A0(n1189), .A1(n1888), .Z(n1446));
Q_MX02 U2264 ( .S(cmd_dgl_data_size[0]), .A0(n1447), .A1(n1881), .Z(cmd_dgl_data[45]));
Q_AN02 U2265 ( .A0(n1189), .A1(n1889), .Z(n1447));
Q_MX02 U2266 ( .S(cmd_dgl_data_size[0]), .A0(n1448), .A1(n1882), .Z(cmd_dgl_data[44]));
Q_AN02 U2267 ( .A0(n1189), .A1(n1890), .Z(n1448));
Q_MX02 U2268 ( .S(cmd_dgl_data_size[0]), .A0(n1449), .A1(n1883), .Z(cmd_dgl_data[43]));
Q_AN02 U2269 ( .A0(n1189), .A1(n1891), .Z(n1449));
Q_MX02 U2270 ( .S(cmd_dgl_data_size[0]), .A0(n1450), .A1(n1884), .Z(cmd_dgl_data[42]));
Q_AN02 U2271 ( .A0(n1189), .A1(n1892), .Z(n1450));
Q_MX02 U2272 ( .S(cmd_dgl_data_size[0]), .A0(n1451), .A1(n1885), .Z(cmd_dgl_data[41]));
Q_AN02 U2273 ( .A0(n1189), .A1(n1893), .Z(n1451));
Q_MX02 U2274 ( .S(cmd_dgl_data_size[0]), .A0(n1452), .A1(n1886), .Z(cmd_dgl_data[40]));
Q_AN02 U2275 ( .A0(n1189), .A1(n1894), .Z(n1452));
Q_MX02 U2276 ( .S(cmd_dgl_data_size[0]), .A0(n1453), .A1(n1887), .Z(cmd_dgl_data[39]));
Q_AN02 U2277 ( .A0(n1189), .A1(n1895), .Z(n1453));
Q_MX02 U2278 ( .S(cmd_dgl_data_size[0]), .A0(n1454), .A1(n1888), .Z(cmd_dgl_data[38]));
Q_AN02 U2279 ( .A0(n1189), .A1(n1896), .Z(n1454));
Q_MX02 U2280 ( .S(cmd_dgl_data_size[0]), .A0(n1455), .A1(n1889), .Z(cmd_dgl_data[37]));
Q_AN02 U2281 ( .A0(n1189), .A1(n1897), .Z(n1455));
Q_MX02 U2282 ( .S(cmd_dgl_data_size[0]), .A0(n1456), .A1(n1890), .Z(cmd_dgl_data[36]));
Q_AN02 U2283 ( .A0(n1189), .A1(n1898), .Z(n1456));
Q_MX02 U2284 ( .S(cmd_dgl_data_size[0]), .A0(n1457), .A1(n1891), .Z(cmd_dgl_data[35]));
Q_AN02 U2285 ( .A0(n1189), .A1(n1899), .Z(n1457));
Q_MX02 U2286 ( .S(cmd_dgl_data_size[0]), .A0(n1458), .A1(n1892), .Z(cmd_dgl_data[34]));
Q_AN02 U2287 ( .A0(n1189), .A1(n1900), .Z(n1458));
Q_MX02 U2288 ( .S(cmd_dgl_data_size[0]), .A0(n1459), .A1(n1893), .Z(cmd_dgl_data[33]));
Q_AN02 U2289 ( .A0(n1189), .A1(n1901), .Z(n1459));
Q_MX02 U2290 ( .S(cmd_dgl_data_size[0]), .A0(n1460), .A1(n1894), .Z(cmd_dgl_data[32]));
Q_AN02 U2291 ( .A0(n1189), .A1(n1902), .Z(n1460));
Q_MX02 U2292 ( .S(cmd_dgl_data_size[0]), .A0(n1461), .A1(n1895), .Z(cmd_dgl_data[31]));
Q_AN02 U2293 ( .A0(n1189), .A1(n1903), .Z(n1461));
Q_MX02 U2294 ( .S(cmd_dgl_data_size[0]), .A0(n1462), .A1(n1896), .Z(cmd_dgl_data[30]));
Q_AN02 U2295 ( .A0(n1189), .A1(n1904), .Z(n1462));
Q_MX02 U2296 ( .S(cmd_dgl_data_size[0]), .A0(n1463), .A1(n1897), .Z(cmd_dgl_data[29]));
Q_AN02 U2297 ( .A0(n1189), .A1(n1905), .Z(n1463));
Q_MX02 U2298 ( .S(cmd_dgl_data_size[0]), .A0(n1464), .A1(n1898), .Z(cmd_dgl_data[28]));
Q_AN02 U2299 ( .A0(n1189), .A1(n1906), .Z(n1464));
Q_MX02 U2300 ( .S(cmd_dgl_data_size[0]), .A0(n1465), .A1(n1899), .Z(cmd_dgl_data[27]));
Q_AN02 U2301 ( .A0(n1189), .A1(n1907), .Z(n1465));
Q_MX02 U2302 ( .S(cmd_dgl_data_size[0]), .A0(n1466), .A1(n1900), .Z(cmd_dgl_data[26]));
Q_AN02 U2303 ( .A0(n1189), .A1(n1908), .Z(n1466));
Q_MX02 U2304 ( .S(cmd_dgl_data_size[0]), .A0(n1467), .A1(n1901), .Z(cmd_dgl_data[25]));
Q_AN02 U2305 ( .A0(n1189), .A1(n1909), .Z(n1467));
Q_MX02 U2306 ( .S(cmd_dgl_data_size[0]), .A0(n1468), .A1(n1902), .Z(cmd_dgl_data[24]));
Q_AN02 U2307 ( .A0(n1189), .A1(n1910), .Z(n1468));
Q_MX02 U2308 ( .S(cmd_dgl_data_size[0]), .A0(n1469), .A1(n1903), .Z(cmd_dgl_data[23]));
Q_AN02 U2309 ( .A0(n1189), .A1(n1911), .Z(n1469));
Q_MX02 U2310 ( .S(cmd_dgl_data_size[0]), .A0(n1470), .A1(n1904), .Z(cmd_dgl_data[22]));
Q_AN02 U2311 ( .A0(n1189), .A1(n1912), .Z(n1470));
Q_MX02 U2312 ( .S(cmd_dgl_data_size[0]), .A0(n1471), .A1(n1905), .Z(cmd_dgl_data[21]));
Q_AN02 U2313 ( .A0(n1189), .A1(n1913), .Z(n1471));
Q_MX02 U2314 ( .S(cmd_dgl_data_size[0]), .A0(n1472), .A1(n1906), .Z(cmd_dgl_data[20]));
Q_AN02 U2315 ( .A0(n1189), .A1(n1914), .Z(n1472));
Q_MX02 U2316 ( .S(cmd_dgl_data_size[0]), .A0(n1473), .A1(n1907), .Z(cmd_dgl_data[19]));
Q_AN02 U2317 ( .A0(n1189), .A1(n1915), .Z(n1473));
Q_MX02 U2318 ( .S(cmd_dgl_data_size[0]), .A0(n1474), .A1(n1908), .Z(cmd_dgl_data[18]));
Q_AN02 U2319 ( .A0(n1189), .A1(n1916), .Z(n1474));
Q_MX02 U2320 ( .S(cmd_dgl_data_size[0]), .A0(n1475), .A1(n1909), .Z(cmd_dgl_data[17]));
Q_AN02 U2321 ( .A0(n1189), .A1(n1917), .Z(n1475));
Q_MX02 U2322 ( .S(cmd_dgl_data_size[0]), .A0(n1476), .A1(n1910), .Z(cmd_dgl_data[16]));
Q_AN02 U2323 ( .A0(n1189), .A1(n1919), .Z(n1476));
Q_MX02 U2324 ( .S(cmd_dgl_data_size[0]), .A0(n1477), .A1(n1911), .Z(cmd_dgl_data[15]));
Q_AN02 U2325 ( .A0(n1189), .A1(n1921), .Z(n1477));
Q_MX02 U2326 ( .S(cmd_dgl_data_size[0]), .A0(n1478), .A1(n1912), .Z(cmd_dgl_data[14]));
Q_AN02 U2327 ( .A0(n1189), .A1(n1922), .Z(n1478));
Q_MX02 U2328 ( .S(cmd_dgl_data_size[0]), .A0(n1479), .A1(n1913), .Z(cmd_dgl_data[13]));
Q_AN02 U2329 ( .A0(n1189), .A1(n1923), .Z(n1479));
Q_MX02 U2330 ( .S(cmd_dgl_data_size[0]), .A0(n1480), .A1(n1914), .Z(cmd_dgl_data[12]));
Q_AN02 U2331 ( .A0(n1189), .A1(n1924), .Z(n1480));
Q_MX02 U2332 ( .S(cmd_dgl_data_size[0]), .A0(n1481), .A1(n1915), .Z(cmd_dgl_data[11]));
Q_AN02 U2333 ( .A0(n1189), .A1(n1925), .Z(n1481));
Q_MX02 U2334 ( .S(cmd_dgl_data_size[0]), .A0(n1482), .A1(n1916), .Z(cmd_dgl_data[10]));
Q_AN02 U2335 ( .A0(n1189), .A1(n1926), .Z(n1482));
Q_MX02 U2336 ( .S(cmd_dgl_data_size[0]), .A0(n1483), .A1(n1917), .Z(cmd_dgl_data[9]));
Q_AN02 U2337 ( .A0(n1189), .A1(n1927), .Z(n1483));
Q_MX02 U2338 ( .S(cmd_dgl_data_size[0]), .A0(n1484), .A1(n1919), .Z(cmd_dgl_data[8]));
Q_AN02 U2339 ( .A0(n1189), .A1(n1928), .Z(n1484));
Q_AN02 U2340 ( .A0(cmd_dgl_data_size[0]), .A1(n1921), .Z(cmd_dgl_data[7]));
Q_AN02 U2341 ( .A0(cmd_dgl_data_size[0]), .A1(n1922), .Z(cmd_dgl_data[6]));
Q_AN02 U2342 ( .A0(cmd_dgl_data_size[0]), .A1(n1923), .Z(cmd_dgl_data[5]));
Q_AN02 U2343 ( .A0(cmd_dgl_data_size[0]), .A1(n1924), .Z(cmd_dgl_data[4]));
Q_AN02 U2344 ( .A0(cmd_dgl_data_size[0]), .A1(n1925), .Z(cmd_dgl_data[3]));
Q_AN02 U2345 ( .A0(cmd_dgl_data_size[0]), .A1(n1926), .Z(cmd_dgl_data[2]));
Q_AN02 U2346 ( .A0(cmd_dgl_data_size[0]), .A1(n1927), .Z(cmd_dgl_data[1]));
Q_AN02 U2347 ( .A0(cmd_dgl_data_size[0]), .A1(n1928), .Z(cmd_dgl_data[0]));
Q_MX02 U2348 ( .S(cmd_dgl_data_size[0]), .A0(n1485), .A1(n266), .Z(cmd_dgl_data[295]));
Q_AN02 U2349 ( .A0(n1189), .A1(n1929), .Z(n1485));
Q_MX02 U2350 ( .S(cmd_dgl_data_size[0]), .A0(n1486), .A1(n267), .Z(cmd_dgl_data[294]));
Q_AN02 U2351 ( .A0(n1189), .A1(n1931), .Z(n1486));
Q_MX02 U2352 ( .S(cmd_dgl_data_size[0]), .A0(n1487), .A1(n268), .Z(cmd_dgl_data[293]));
Q_AN02 U2353 ( .A0(n1189), .A1(n1933), .Z(n1487));
Q_MX02 U2354 ( .S(cmd_dgl_data_size[0]), .A0(n1488), .A1(n269), .Z(cmd_dgl_data[292]));
Q_AN02 U2355 ( .A0(n1189), .A1(n1935), .Z(n1488));
Q_MX02 U2356 ( .S(cmd_dgl_data_size[0]), .A0(n1489), .A1(n270), .Z(cmd_dgl_data[291]));
Q_AN02 U2357 ( .A0(n1189), .A1(n1937), .Z(n1489));
Q_MX02 U2358 ( .S(cmd_dgl_data_size[0]), .A0(n1490), .A1(n271), .Z(cmd_dgl_data[290]));
Q_AN02 U2359 ( .A0(n1189), .A1(n1939), .Z(n1490));
Q_MX02 U2360 ( .S(cmd_dgl_data_size[0]), .A0(n1491), .A1(n272), .Z(cmd_dgl_data[289]));
Q_AN02 U2361 ( .A0(n1189), .A1(n1941), .Z(n1491));
Q_MX02 U2362 ( .S(cmd_dgl_data_size[0]), .A0(n1492), .A1(n273), .Z(cmd_dgl_data[288]));
Q_AN02 U2363 ( .A0(n1189), .A1(n1943), .Z(n1492));
Q_MX02 U2364 ( .S(n1192), .A0(n1494), .A1(cmdfifo_kdfstream_cmd[252]), .Z(n1493));
Q_AN02 U2365 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[124]), .Z(n1494));
Q_MX02 U2366 ( .S(n1192), .A0(n1496), .A1(cmdfifo_kdfstream_cmd[251]), .Z(n1495));
Q_AN02 U2367 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[123]), .Z(n1496));
Q_MX02 U2368 ( .S(n1192), .A0(n1498), .A1(cmdfifo_kdfstream_cmd[250]), .Z(n1497));
Q_AN02 U2369 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[122]), .Z(n1498));
Q_MX02 U2370 ( .S(n1192), .A0(n1500), .A1(cmdfifo_kdfstream_cmd[249]), .Z(n1499));
Q_AN02 U2371 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[121]), .Z(n1500));
Q_MX02 U2372 ( .S(n1192), .A0(n1502), .A1(cmdfifo_kdfstream_cmd[248]), .Z(n1501));
Q_AN02 U2373 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[120]), .Z(n1502));
Q_MX02 U2374 ( .S(n1192), .A0(n1504), .A1(cmdfifo_kdfstream_cmd[247]), .Z(n1503));
Q_AN02 U2375 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[119]), .Z(n1504));
Q_MX02 U2376 ( .S(n1192), .A0(n1506), .A1(cmdfifo_kdfstream_cmd[246]), .Z(n1505));
Q_AN02 U2377 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[118]), .Z(n1506));
Q_MX02 U2378 ( .S(n1192), .A0(n1508), .A1(cmdfifo_kdfstream_cmd[245]), .Z(n1507));
Q_AN02 U2379 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[117]), .Z(n1508));
Q_MX02 U2380 ( .S(n1192), .A0(n1510), .A1(cmdfifo_kdfstream_cmd[244]), .Z(n1509));
Q_AN02 U2381 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[116]), .Z(n1510));
Q_MX02 U2382 ( .S(n1192), .A0(n1512), .A1(cmdfifo_kdfstream_cmd[243]), .Z(n1511));
Q_AN02 U2383 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[115]), .Z(n1512));
Q_MX02 U2384 ( .S(n1192), .A0(n1514), .A1(cmdfifo_kdfstream_cmd[242]), .Z(n1513));
Q_AN02 U2385 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[114]), .Z(n1514));
Q_MX02 U2386 ( .S(n1192), .A0(n1516), .A1(cmdfifo_kdfstream_cmd[241]), .Z(n1515));
Q_AN02 U2387 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[113]), .Z(n1516));
Q_MX02 U2388 ( .S(n1192), .A0(n1518), .A1(cmdfifo_kdfstream_cmd[240]), .Z(n1517));
Q_AN02 U2389 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[112]), .Z(n1518));
Q_MX02 U2390 ( .S(n1192), .A0(n1520), .A1(cmdfifo_kdfstream_cmd[239]), .Z(n1519));
Q_AN02 U2391 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[111]), .Z(n1520));
Q_MX02 U2392 ( .S(n1192), .A0(n1522), .A1(cmdfifo_kdfstream_cmd[238]), .Z(n1521));
Q_AN02 U2393 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[110]), .Z(n1522));
Q_MX02 U2394 ( .S(n1192), .A0(n1524), .A1(cmdfifo_kdfstream_cmd[237]), .Z(n1523));
Q_AN02 U2395 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[109]), .Z(n1524));
Q_MX02 U2396 ( .S(n1192), .A0(n1526), .A1(cmdfifo_kdfstream_cmd[236]), .Z(n1525));
Q_AN02 U2397 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[108]), .Z(n1526));
Q_MX02 U2398 ( .S(n1192), .A0(n1528), .A1(cmdfifo_kdfstream_cmd[235]), .Z(n1527));
Q_AN02 U2399 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[107]), .Z(n1528));
Q_MX02 U2400 ( .S(n1192), .A0(n1530), .A1(cmdfifo_kdfstream_cmd[234]), .Z(n1529));
Q_AN02 U2401 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[106]), .Z(n1530));
Q_MX02 U2402 ( .S(n1192), .A0(n1532), .A1(cmdfifo_kdfstream_cmd[233]), .Z(n1531));
Q_AN02 U2403 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[105]), .Z(n1532));
Q_MX02 U2404 ( .S(n1192), .A0(n1534), .A1(cmdfifo_kdfstream_cmd[232]), .Z(n1533));
Q_AN02 U2405 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[104]), .Z(n1534));
Q_MX02 U2406 ( .S(n1192), .A0(n1536), .A1(cmdfifo_kdfstream_cmd[231]), .Z(n1535));
Q_AN02 U2407 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[103]), .Z(n1536));
Q_MX02 U2408 ( .S(n1192), .A0(n1538), .A1(cmdfifo_kdfstream_cmd[230]), .Z(n1537));
Q_AN02 U2409 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[102]), .Z(n1538));
Q_MX02 U2410 ( .S(n1192), .A0(n1540), .A1(cmdfifo_kdfstream_cmd[229]), .Z(n1539));
Q_AN02 U2411 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[101]), .Z(n1540));
Q_MX02 U2412 ( .S(n1192), .A0(n1542), .A1(cmdfifo_kdfstream_cmd[228]), .Z(n1541));
Q_AN02 U2413 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[100]), .Z(n1542));
Q_MX02 U2414 ( .S(n1192), .A0(n1544), .A1(cmdfifo_kdfstream_cmd[227]), .Z(n1543));
Q_AN02 U2415 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[99]), .Z(n1544));
Q_MX02 U2416 ( .S(n1192), .A0(n1546), .A1(cmdfifo_kdfstream_cmd[226]), .Z(n1545));
Q_AN02 U2417 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[98]), .Z(n1546));
Q_MX02 U2418 ( .S(n1192), .A0(n1548), .A1(cmdfifo_kdfstream_cmd[225]), .Z(n1547));
Q_AN02 U2419 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[97]), .Z(n1548));
Q_MX02 U2420 ( .S(n1192), .A0(n1550), .A1(cmdfifo_kdfstream_cmd[224]), .Z(n1549));
Q_AN02 U2421 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[96]), .Z(n1550));
Q_MX02 U2422 ( .S(n1192), .A0(n1552), .A1(cmdfifo_kdfstream_cmd[223]), .Z(n1551));
Q_AN02 U2423 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[95]), .Z(n1552));
Q_MX02 U2424 ( .S(n1192), .A0(n1554), .A1(cmdfifo_kdfstream_cmd[222]), .Z(n1553));
Q_AN02 U2425 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[94]), .Z(n1554));
Q_MX02 U2426 ( .S(n1192), .A0(n1556), .A1(cmdfifo_kdfstream_cmd[221]), .Z(n1555));
Q_AN02 U2427 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[93]), .Z(n1556));
Q_MX02 U2428 ( .S(n1192), .A0(n1558), .A1(cmdfifo_kdfstream_cmd[220]), .Z(n1557));
Q_AN02 U2429 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[92]), .Z(n1558));
Q_MX02 U2430 ( .S(n1192), .A0(n1560), .A1(cmdfifo_kdfstream_cmd[219]), .Z(n1559));
Q_AN02 U2431 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[91]), .Z(n1560));
Q_MX02 U2432 ( .S(n1192), .A0(n1562), .A1(cmdfifo_kdfstream_cmd[218]), .Z(n1561));
Q_AN02 U2433 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[90]), .Z(n1562));
Q_MX02 U2434 ( .S(n1192), .A0(n1564), .A1(cmdfifo_kdfstream_cmd[217]), .Z(n1563));
Q_AN02 U2435 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[89]), .Z(n1564));
Q_MX02 U2436 ( .S(n1192), .A0(n1566), .A1(cmdfifo_kdfstream_cmd[216]), .Z(n1565));
Q_AN02 U2437 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[88]), .Z(n1566));
Q_MX02 U2438 ( .S(n1192), .A0(n1568), .A1(cmdfifo_kdfstream_cmd[215]), .Z(n1567));
Q_AN02 U2439 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[87]), .Z(n1568));
Q_MX02 U2440 ( .S(n1192), .A0(n1570), .A1(cmdfifo_kdfstream_cmd[214]), .Z(n1569));
Q_AN02 U2441 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[86]), .Z(n1570));
Q_MX02 U2442 ( .S(n1192), .A0(n1572), .A1(cmdfifo_kdfstream_cmd[213]), .Z(n1571));
Q_AN02 U2443 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[85]), .Z(n1572));
Q_MX02 U2444 ( .S(n1192), .A0(n1574), .A1(cmdfifo_kdfstream_cmd[212]), .Z(n1573));
Q_AN02 U2445 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[84]), .Z(n1574));
Q_MX02 U2446 ( .S(n1192), .A0(n1576), .A1(cmdfifo_kdfstream_cmd[211]), .Z(n1575));
Q_AN02 U2447 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[83]), .Z(n1576));
Q_MX02 U2448 ( .S(n1192), .A0(n1578), .A1(cmdfifo_kdfstream_cmd[210]), .Z(n1577));
Q_AN02 U2449 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[82]), .Z(n1578));
Q_MX02 U2450 ( .S(n1192), .A0(n1580), .A1(cmdfifo_kdfstream_cmd[209]), .Z(n1579));
Q_AN02 U2451 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[81]), .Z(n1580));
Q_MX02 U2452 ( .S(n1192), .A0(n1582), .A1(cmdfifo_kdfstream_cmd[208]), .Z(n1581));
Q_AN02 U2453 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[80]), .Z(n1582));
Q_MX02 U2454 ( .S(n1192), .A0(n1584), .A1(cmdfifo_kdfstream_cmd[207]), .Z(n1583));
Q_AN02 U2455 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[79]), .Z(n1584));
Q_MX02 U2456 ( .S(n1192), .A0(n1586), .A1(cmdfifo_kdfstream_cmd[206]), .Z(n1585));
Q_AN02 U2457 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[78]), .Z(n1586));
Q_MX02 U2458 ( .S(n1192), .A0(n1588), .A1(cmdfifo_kdfstream_cmd[205]), .Z(n1587));
Q_AN02 U2459 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[77]), .Z(n1588));
Q_MX02 U2460 ( .S(n1192), .A0(n1590), .A1(cmdfifo_kdfstream_cmd[204]), .Z(n1589));
Q_AN02 U2461 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[76]), .Z(n1590));
Q_MX02 U2462 ( .S(n1192), .A0(n1592), .A1(cmdfifo_kdfstream_cmd[203]), .Z(n1591));
Q_AN02 U2463 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[75]), .Z(n1592));
Q_MX02 U2464 ( .S(n1192), .A0(n1594), .A1(cmdfifo_kdfstream_cmd[202]), .Z(n1593));
Q_AN02 U2465 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[74]), .Z(n1594));
Q_MX02 U2466 ( .S(n1192), .A0(n1596), .A1(cmdfifo_kdfstream_cmd[201]), .Z(n1595));
Q_AN02 U2467 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[73]), .Z(n1596));
Q_MX02 U2468 ( .S(n1192), .A0(n1598), .A1(cmdfifo_kdfstream_cmd[200]), .Z(n1597));
Q_AN02 U2469 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[72]), .Z(n1598));
Q_MX02 U2470 ( .S(n1192), .A0(n1600), .A1(cmdfifo_kdfstream_cmd[199]), .Z(n1599));
Q_AN02 U2471 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[71]), .Z(n1600));
Q_MX02 U2472 ( .S(n1192), .A0(n1602), .A1(cmdfifo_kdfstream_cmd[198]), .Z(n1601));
Q_AN02 U2473 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[70]), .Z(n1602));
Q_MX02 U2474 ( .S(n1192), .A0(n1604), .A1(cmdfifo_kdfstream_cmd[197]), .Z(n1603));
Q_AN02 U2475 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[69]), .Z(n1604));
Q_MX02 U2476 ( .S(n1192), .A0(n1606), .A1(cmdfifo_kdfstream_cmd[196]), .Z(n1605));
Q_AN02 U2477 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[68]), .Z(n1606));
Q_MX02 U2478 ( .S(n1192), .A0(n1608), .A1(cmdfifo_kdfstream_cmd[195]), .Z(n1607));
Q_AN02 U2479 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[67]), .Z(n1608));
Q_MX02 U2480 ( .S(n1192), .A0(n1610), .A1(cmdfifo_kdfstream_cmd[194]), .Z(n1609));
Q_AN02 U2481 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[66]), .Z(n1610));
Q_MX02 U2482 ( .S(n1192), .A0(n1612), .A1(cmdfifo_kdfstream_cmd[193]), .Z(n1611));
Q_AN02 U2483 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[65]), .Z(n1612));
Q_MX02 U2484 ( .S(n1192), .A0(n1614), .A1(cmdfifo_kdfstream_cmd[192]), .Z(n1613));
Q_AN02 U2485 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[64]), .Z(n1614));
Q_MX02 U2486 ( .S(n1192), .A0(n1616), .A1(cmdfifo_kdfstream_cmd[191]), .Z(n1615));
Q_AN02 U2487 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[63]), .Z(n1616));
Q_MX02 U2488 ( .S(n1192), .A0(n1618), .A1(cmdfifo_kdfstream_cmd[190]), .Z(n1617));
Q_AN02 U2489 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[62]), .Z(n1618));
Q_MX02 U2490 ( .S(n1192), .A0(n1620), .A1(cmdfifo_kdfstream_cmd[189]), .Z(n1619));
Q_AN02 U2491 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[61]), .Z(n1620));
Q_MX02 U2492 ( .S(n1192), .A0(n1622), .A1(cmdfifo_kdfstream_cmd[188]), .Z(n1621));
Q_AN02 U2493 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[60]), .Z(n1622));
Q_MX02 U2494 ( .S(n1192), .A0(n1624), .A1(cmdfifo_kdfstream_cmd[187]), .Z(n1623));
Q_AN02 U2495 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[59]), .Z(n1624));
Q_MX02 U2496 ( .S(n1192), .A0(n1626), .A1(cmdfifo_kdfstream_cmd[186]), .Z(n1625));
Q_AN02 U2497 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[58]), .Z(n1626));
Q_MX02 U2498 ( .S(n1192), .A0(n1628), .A1(cmdfifo_kdfstream_cmd[185]), .Z(n1627));
Q_AN02 U2499 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[57]), .Z(n1628));
Q_MX02 U2500 ( .S(n1192), .A0(n1630), .A1(cmdfifo_kdfstream_cmd[184]), .Z(n1629));
Q_AN02 U2501 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[56]), .Z(n1630));
Q_MX02 U2502 ( .S(n1192), .A0(n1632), .A1(cmdfifo_kdfstream_cmd[183]), .Z(n1631));
Q_AN02 U2503 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[55]), .Z(n1632));
Q_MX02 U2504 ( .S(n1192), .A0(n1634), .A1(cmdfifo_kdfstream_cmd[182]), .Z(n1633));
Q_AN02 U2505 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[54]), .Z(n1634));
Q_MX02 U2506 ( .S(n1192), .A0(n1636), .A1(cmdfifo_kdfstream_cmd[181]), .Z(n1635));
Q_AN02 U2507 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[53]), .Z(n1636));
Q_MX02 U2508 ( .S(n1192), .A0(n1638), .A1(cmdfifo_kdfstream_cmd[180]), .Z(n1637));
Q_AN02 U2509 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[52]), .Z(n1638));
Q_MX02 U2510 ( .S(n1192), .A0(n1640), .A1(cmdfifo_kdfstream_cmd[179]), .Z(n1639));
Q_AN02 U2511 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[51]), .Z(n1640));
Q_MX02 U2512 ( .S(n1192), .A0(n1642), .A1(cmdfifo_kdfstream_cmd[178]), .Z(n1641));
Q_AN02 U2513 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[50]), .Z(n1642));
Q_MX02 U2514 ( .S(n1192), .A0(n1644), .A1(cmdfifo_kdfstream_cmd[177]), .Z(n1643));
Q_AN02 U2515 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[49]), .Z(n1644));
Q_MX02 U2516 ( .S(n1192), .A0(n1646), .A1(cmdfifo_kdfstream_cmd[176]), .Z(n1645));
Q_AN02 U2517 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[48]), .Z(n1646));
Q_MX02 U2518 ( .S(n1192), .A0(n1648), .A1(cmdfifo_kdfstream_cmd[175]), .Z(n1647));
Q_AN02 U2519 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[47]), .Z(n1648));
Q_MX02 U2520 ( .S(n1192), .A0(n1650), .A1(cmdfifo_kdfstream_cmd[174]), .Z(n1649));
Q_AN02 U2521 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[46]), .Z(n1650));
Q_MX02 U2522 ( .S(n1192), .A0(n1652), .A1(cmdfifo_kdfstream_cmd[173]), .Z(n1651));
Q_AN02 U2523 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[45]), .Z(n1652));
Q_MX02 U2524 ( .S(n1192), .A0(n1654), .A1(cmdfifo_kdfstream_cmd[172]), .Z(n1653));
Q_AN02 U2525 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[44]), .Z(n1654));
Q_MX02 U2526 ( .S(n1192), .A0(n1656), .A1(cmdfifo_kdfstream_cmd[171]), .Z(n1655));
Q_AN02 U2527 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[43]), .Z(n1656));
Q_MX02 U2528 ( .S(n1192), .A0(n1658), .A1(cmdfifo_kdfstream_cmd[170]), .Z(n1657));
Q_AN02 U2529 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[42]), .Z(n1658));
Q_MX02 U2530 ( .S(n1192), .A0(n1660), .A1(cmdfifo_kdfstream_cmd[169]), .Z(n1659));
Q_AN02 U2531 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[41]), .Z(n1660));
Q_MX02 U2532 ( .S(n1192), .A0(n1662), .A1(cmdfifo_kdfstream_cmd[168]), .Z(n1661));
Q_AN02 U2533 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[40]), .Z(n1662));
Q_MX02 U2534 ( .S(n1192), .A0(n1664), .A1(cmdfifo_kdfstream_cmd[167]), .Z(n1663));
Q_AN02 U2535 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[39]), .Z(n1664));
Q_MX02 U2536 ( .S(n1192), .A0(n1666), .A1(cmdfifo_kdfstream_cmd[166]), .Z(n1665));
Q_AN02 U2537 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[38]), .Z(n1666));
Q_MX02 U2538 ( .S(n1192), .A0(n1668), .A1(cmdfifo_kdfstream_cmd[165]), .Z(n1667));
Q_AN02 U2539 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[37]), .Z(n1668));
Q_MX02 U2540 ( .S(n1192), .A0(n1670), .A1(cmdfifo_kdfstream_cmd[164]), .Z(n1669));
Q_AN02 U2541 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[36]), .Z(n1670));
Q_MX02 U2542 ( .S(n1192), .A0(n1672), .A1(cmdfifo_kdfstream_cmd[163]), .Z(n1671));
Q_AN02 U2543 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[35]), .Z(n1672));
Q_MX02 U2544 ( .S(n1192), .A0(n1674), .A1(cmdfifo_kdfstream_cmd[162]), .Z(n1673));
Q_AN02 U2545 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[34]), .Z(n1674));
Q_MX02 U2546 ( .S(n1192), .A0(n1676), .A1(cmdfifo_kdfstream_cmd[161]), .Z(n1675));
Q_AN02 U2547 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[33]), .Z(n1676));
Q_MX02 U2548 ( .S(n1192), .A0(n1678), .A1(cmdfifo_kdfstream_cmd[160]), .Z(n1677));
Q_AN02 U2549 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[32]), .Z(n1678));
Q_MX02 U2550 ( .S(n1192), .A0(n1680), .A1(cmdfifo_kdfstream_cmd[159]), .Z(n1679));
Q_AN02 U2551 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[31]), .Z(n1680));
Q_MX02 U2552 ( .S(n1192), .A0(n1682), .A1(cmdfifo_kdfstream_cmd[158]), .Z(n1681));
Q_AN02 U2553 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[30]), .Z(n1682));
Q_MX02 U2554 ( .S(n1192), .A0(n1684), .A1(cmdfifo_kdfstream_cmd[157]), .Z(n1683));
Q_AN02 U2555 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[29]), .Z(n1684));
Q_MX02 U2556 ( .S(n1192), .A0(n1686), .A1(cmdfifo_kdfstream_cmd[156]), .Z(n1685));
Q_AN02 U2557 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[28]), .Z(n1686));
Q_MX02 U2558 ( .S(n1192), .A0(n1688), .A1(cmdfifo_kdfstream_cmd[155]), .Z(n1687));
Q_AN02 U2559 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[27]), .Z(n1688));
Q_MX02 U2560 ( .S(n1192), .A0(n1690), .A1(cmdfifo_kdfstream_cmd[154]), .Z(n1689));
Q_AN02 U2561 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[26]), .Z(n1690));
Q_MX02 U2562 ( .S(n1192), .A0(n1692), .A1(cmdfifo_kdfstream_cmd[153]), .Z(n1691));
Q_AN02 U2563 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[25]), .Z(n1692));
Q_MX02 U2564 ( .S(n1192), .A0(n1694), .A1(cmdfifo_kdfstream_cmd[152]), .Z(n1693));
Q_AN02 U2565 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[24]), .Z(n1694));
Q_MX02 U2566 ( .S(n1192), .A0(n1696), .A1(cmdfifo_kdfstream_cmd[151]), .Z(n1695));
Q_AN02 U2567 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[23]), .Z(n1696));
Q_MX02 U2568 ( .S(n1192), .A0(n1698), .A1(cmdfifo_kdfstream_cmd[150]), .Z(n1697));
Q_AN02 U2569 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[22]), .Z(n1698));
Q_MX02 U2570 ( .S(n1192), .A0(n1700), .A1(cmdfifo_kdfstream_cmd[149]), .Z(n1699));
Q_AN02 U2571 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[21]), .Z(n1700));
Q_MX02 U2572 ( .S(n1192), .A0(n1702), .A1(cmdfifo_kdfstream_cmd[148]), .Z(n1701));
Q_AN02 U2573 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[20]), .Z(n1702));
Q_MX02 U2574 ( .S(n1192), .A0(n1704), .A1(cmdfifo_kdfstream_cmd[147]), .Z(n1703));
Q_AN02 U2575 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[19]), .Z(n1704));
Q_MX02 U2576 ( .S(n1192), .A0(n1706), .A1(cmdfifo_kdfstream_cmd[146]), .Z(n1705));
Q_AN02 U2577 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[18]), .Z(n1706));
Q_MX02 U2578 ( .S(n1192), .A0(n1708), .A1(cmdfifo_kdfstream_cmd[145]), .Z(n1707));
Q_AN02 U2579 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[17]), .Z(n1708));
Q_MX02 U2580 ( .S(n1192), .A0(n1710), .A1(cmdfifo_kdfstream_cmd[144]), .Z(n1709));
Q_AN02 U2581 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[16]), .Z(n1710));
Q_MX02 U2582 ( .S(n1192), .A0(n1712), .A1(cmdfifo_kdfstream_cmd[143]), .Z(n1711));
Q_AN02 U2583 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[15]), .Z(n1712));
Q_MX02 U2584 ( .S(n1192), .A0(n1714), .A1(cmdfifo_kdfstream_cmd[142]), .Z(n1713));
Q_AN02 U2585 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[14]), .Z(n1714));
Q_MX02 U2586 ( .S(n1192), .A0(n1716), .A1(cmdfifo_kdfstream_cmd[141]), .Z(n1715));
Q_AN02 U2587 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[13]), .Z(n1716));
Q_MX02 U2588 ( .S(n1192), .A0(n1718), .A1(cmdfifo_kdfstream_cmd[140]), .Z(n1717));
Q_AN02 U2589 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[12]), .Z(n1718));
Q_MX02 U2590 ( .S(n1192), .A0(n1720), .A1(cmdfifo_kdfstream_cmd[139]), .Z(n1719));
Q_AN02 U2591 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[11]), .Z(n1720));
Q_MX02 U2592 ( .S(n1192), .A0(n1722), .A1(cmdfifo_kdfstream_cmd[138]), .Z(n1721));
Q_AN02 U2593 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[10]), .Z(n1722));
Q_MX02 U2594 ( .S(n1192), .A0(n1724), .A1(cmdfifo_kdfstream_cmd[137]), .Z(n1723));
Q_AN02 U2595 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[9]), .Z(n1724));
Q_MX02 U2596 ( .S(n1192), .A0(n1726), .A1(cmdfifo_kdfstream_cmd[136]), .Z(n1725));
Q_AN02 U2597 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[8]), .Z(n1726));
Q_MX02 U2598 ( .S(n1192), .A0(n1728), .A1(cmdfifo_kdfstream_cmd[135]), .Z(n1727));
Q_AN02 U2599 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[7]), .Z(n1728));
Q_MX02 U2600 ( .S(n1192), .A0(n1730), .A1(cmdfifo_kdfstream_cmd[134]), .Z(n1729));
Q_AN02 U2601 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[6]), .Z(n1730));
Q_MX02 U2602 ( .S(n1192), .A0(n1732), .A1(cmdfifo_kdfstream_cmd[133]), .Z(n1731));
Q_AN02 U2603 ( .A0(n1972), .A1(cmdfifo_kdfstream_cmd[5]), .Z(n1732));
Q_MX02 U2604 ( .S(n1192), .A0(n1734), .A1(cmdfifo_kdfstream_cmd[132]), .Z(n1733));
Q_AN02 U2605 ( .A0(n1972), .A1(iter3_kdf_key_size[31]), .Z(n1734));
Q_MX02 U2606 ( .S(n1192), .A0(n1736), .A1(cmdfifo_kdfstream_cmd[131]), .Z(n1735));
Q_AN02 U2607 ( .A0(n1972), .A1(iter3_kdf_key_size[30]), .Z(n1736));
Q_MX02 U2608 ( .S(n1192), .A0(n1738), .A1(cmdfifo_kdfstream_cmd[130]), .Z(n1737));
Q_AN02 U2609 ( .A0(n1972), .A1(iter3_kdf_key_size[29]), .Z(n1738));
Q_MX02 U2610 ( .S(n1192), .A0(n1740), .A1(cmdfifo_kdfstream_cmd[129]), .Z(n1739));
Q_AN02 U2611 ( .A0(n1972), .A1(iter3_kdf_key_size[28]), .Z(n1740));
Q_MX02 U2612 ( .S(n1192), .A0(n1742), .A1(cmdfifo_kdfstream_cmd[128]), .Z(n1741));
Q_AN02 U2613 ( .A0(n1972), .A1(iter3_kdf_key_size[27]), .Z(n1742));
Q_MX02 U2614 ( .S(n1192), .A0(n1744), .A1(cmdfifo_kdfstream_cmd[127]), .Z(n1743));
Q_AN02 U2615 ( .A0(n1972), .A1(iter3_kdf_key_size[26]), .Z(n1744));
Q_MX02 U2616 ( .S(n1192), .A0(n1746), .A1(cmdfifo_kdfstream_cmd[126]), .Z(n1745));
Q_AN02 U2617 ( .A0(n1972), .A1(iter3_kdf_key_size[25]), .Z(n1746));
Q_MX02 U2618 ( .S(n1192), .A0(n1748), .A1(cmdfifo_kdfstream_cmd[125]), .Z(n1747));
Q_AN02 U2619 ( .A0(n1972), .A1(iter3_kdf_key_size[24]), .Z(n1748));
Q_MX02 U2620 ( .S(n1192), .A0(n1750), .A1(cmdfifo_kdfstream_cmd[124]), .Z(n1749));
Q_AN02 U2621 ( .A0(n1972), .A1(iter3_kdf_key_size[23]), .Z(n1750));
Q_MX02 U2622 ( .S(n1192), .A0(n1752), .A1(cmdfifo_kdfstream_cmd[123]), .Z(n1751));
Q_AN02 U2623 ( .A0(n1972), .A1(iter3_kdf_key_size[22]), .Z(n1752));
Q_MX02 U2624 ( .S(n1192), .A0(n1754), .A1(cmdfifo_kdfstream_cmd[122]), .Z(n1753));
Q_AN02 U2625 ( .A0(n1972), .A1(iter3_kdf_key_size[21]), .Z(n1754));
Q_MX02 U2626 ( .S(n1192), .A0(n1756), .A1(cmdfifo_kdfstream_cmd[121]), .Z(n1755));
Q_AN02 U2627 ( .A0(n1972), .A1(iter3_kdf_key_size[20]), .Z(n1756));
Q_MX02 U2628 ( .S(n1192), .A0(n1758), .A1(cmdfifo_kdfstream_cmd[120]), .Z(n1757));
Q_AN02 U2629 ( .A0(n1972), .A1(iter3_kdf_key_size[19]), .Z(n1758));
Q_MX02 U2630 ( .S(n1192), .A0(n1760), .A1(cmdfifo_kdfstream_cmd[119]), .Z(n1759));
Q_AN02 U2631 ( .A0(n1972), .A1(iter3_kdf_key_size[18]), .Z(n1760));
Q_MX02 U2632 ( .S(n1192), .A0(n1762), .A1(cmdfifo_kdfstream_cmd[118]), .Z(n1761));
Q_AN02 U2633 ( .A0(n1972), .A1(iter3_kdf_key_size[17]), .Z(n1762));
Q_MX02 U2634 ( .S(n1192), .A0(n1764), .A1(cmdfifo_kdfstream_cmd[117]), .Z(n1763));
Q_AN02 U2635 ( .A0(n1972), .A1(iter3_kdf_key_size[16]), .Z(n1764));
Q_MX02 U2636 ( .S(n1192), .A0(n1766), .A1(cmdfifo_kdfstream_cmd[116]), .Z(n1765));
Q_AN02 U2637 ( .A0(n1972), .A1(iter3_kdf_key_size[15]), .Z(n1766));
Q_MX02 U2638 ( .S(n1192), .A0(n1768), .A1(cmdfifo_kdfstream_cmd[115]), .Z(n1767));
Q_AN02 U2639 ( .A0(n1972), .A1(iter3_kdf_key_size[14]), .Z(n1768));
Q_MX02 U2640 ( .S(n1192), .A0(n1770), .A1(cmdfifo_kdfstream_cmd[114]), .Z(n1769));
Q_AN02 U2641 ( .A0(n1972), .A1(iter3_kdf_key_size[13]), .Z(n1770));
Q_MX02 U2642 ( .S(n1192), .A0(n1772), .A1(cmdfifo_kdfstream_cmd[113]), .Z(n1771));
Q_AN02 U2643 ( .A0(n1972), .A1(iter3_kdf_key_size[12]), .Z(n1772));
Q_MX02 U2644 ( .S(n1192), .A0(n1774), .A1(cmdfifo_kdfstream_cmd[112]), .Z(n1773));
Q_AN02 U2645 ( .A0(n1972), .A1(iter3_kdf_key_size[11]), .Z(n1774));
Q_MX02 U2646 ( .S(n1192), .A0(n1776), .A1(cmdfifo_kdfstream_cmd[111]), .Z(n1775));
Q_AN02 U2647 ( .A0(n1972), .A1(iter3_kdf_key_size[10]), .Z(n1776));
Q_MX03 U2648 ( .S0(n1190), .S1(n1192), .A0(n1778), .A1(n1779), .A2(cmdfifo_kdfstream_cmd[110]), .Z(n1777));
Q_AN02 U2649 ( .A0(n1191), .A1(iter3_kdf_key_size[9]), .Z(n1778));
Q_MX02 U2650 ( .S(n1191), .A0(iter3_kdf_key_size[9]), .A1(iter1_kdf_key_size[9]), .Z(n1779));
Q_MX03 U2651 ( .S0(n1190), .S1(n1192), .A0(n1781), .A1(n1782), .A2(cmdfifo_kdfstream_cmd[109]), .Z(n1780));
Q_AN02 U2652 ( .A0(n1191), .A1(iter3_kdf_key_size[8]), .Z(n1781));
Q_MX02 U2653 ( .S(n1191), .A0(iter2_kdf_key_size[8]), .A1(iter3_kdf_key_size[8]), .Z(n1782));
Q_MX02 U2654 ( .S(n1192), .A0(n1784), .A1(cmdfifo_kdfstream_cmd[108]), .Z(n1783));
Q_AN02 U2655 ( .A0(n1972), .A1(iter3_kdf_key_size[7]), .Z(n1784));
Q_MX02 U2656 ( .S(n1192), .A0(n1786), .A1(cmdfifo_kdfstream_cmd[107]), .Z(n1785));
Q_AN02 U2657 ( .A0(n1972), .A1(iter3_kdf_key_size[6]), .Z(n1786));
Q_MX02 U2658 ( .S(n1192), .A0(n1788), .A1(cmdfifo_kdfstream_cmd[106]), .Z(n1787));
Q_AN02 U2659 ( .A0(n1972), .A1(iter3_kdf_key_size[5]), .Z(n1788));
Q_MX02 U2660 ( .S(n1192), .A0(n1790), .A1(cmdfifo_kdfstream_cmd[105]), .Z(n1789));
Q_AN02 U2661 ( .A0(n1972), .A1(iter3_kdf_key_size[4]), .Z(n1790));
Q_MX02 U2662 ( .S(n1192), .A0(n1792), .A1(cmdfifo_kdfstream_cmd[104]), .Z(n1791));
Q_AN02 U2663 ( .A0(n1972), .A1(iter3_kdf_key_size[3]), .Z(n1792));
Q_MX02 U2664 ( .S(n1192), .A0(n1794), .A1(cmdfifo_kdfstream_cmd[103]), .Z(n1793));
Q_AN02 U2665 ( .A0(n1972), .A1(iter3_kdf_key_size[2]), .Z(n1794));
Q_MX02 U2666 ( .S(n1192), .A0(n1796), .A1(cmdfifo_kdfstream_cmd[102]), .Z(n1795));
Q_AN02 U2667 ( .A0(n1972), .A1(iter3_kdf_key_size[1]), .Z(n1796));
Q_MX02 U2668 ( .S(n1192), .A0(n1798), .A1(cmdfifo_kdfstream_cmd[101]), .Z(n1797));
Q_AN02 U2669 ( .A0(n1972), .A1(iter3_kdf_key_size[0]), .Z(n1798));
Q_AN02 U2670 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[100]), .Z(n1799));
Q_AN02 U2671 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[99]), .Z(n1800));
Q_AN02 U2672 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[98]), .Z(n1801));
Q_AN02 U2673 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[97]), .Z(n1802));
Q_AN02 U2674 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[96]), .Z(n1803));
Q_AN02 U2675 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[95]), .Z(n1804));
Q_AN02 U2676 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[94]), .Z(n1805));
Q_AN02 U2677 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[93]), .Z(n1806));
Q_AN02 U2678 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[92]), .Z(n1807));
Q_AN02 U2679 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[91]), .Z(n1808));
Q_AN02 U2680 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[90]), .Z(n1809));
Q_AN02 U2681 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[89]), .Z(n1810));
Q_AN02 U2682 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[88]), .Z(n1811));
Q_AN02 U2683 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[87]), .Z(n1812));
Q_AN02 U2684 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[86]), .Z(n1813));
Q_AN02 U2685 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[85]), .Z(n1814));
Q_AN02 U2686 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[84]), .Z(n1815));
Q_AN02 U2687 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[83]), .Z(n1816));
Q_AN02 U2688 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[82]), .Z(n1817));
Q_AN02 U2689 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[81]), .Z(n1818));
Q_AN02 U2690 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[80]), .Z(n1819));
Q_AN02 U2691 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[79]), .Z(n1820));
Q_AN02 U2692 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[78]), .Z(n1821));
Q_AN02 U2693 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[77]), .Z(n1822));
Q_AN02 U2694 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[76]), .Z(n1823));
Q_AN02 U2695 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[75]), .Z(n1824));
Q_AN02 U2696 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[74]), .Z(n1825));
Q_AN02 U2697 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[73]), .Z(n1826));
Q_AN02 U2698 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[72]), .Z(n1827));
Q_AN02 U2699 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[71]), .Z(n1828));
Q_AN02 U2700 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[70]), .Z(n1829));
Q_AN02 U2701 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[69]), .Z(n1830));
Q_AN02 U2702 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[68]), .Z(n1831));
Q_AN02 U2703 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[67]), .Z(n1832));
Q_AN02 U2704 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[66]), .Z(n1833));
Q_AN02 U2705 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[65]), .Z(n1834));
Q_AN02 U2706 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[64]), .Z(n1835));
Q_AN02 U2707 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[63]), .Z(n1836));
Q_AN02 U2708 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[62]), .Z(n1837));
Q_AN02 U2709 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[61]), .Z(n1838));
Q_AN02 U2710 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[60]), .Z(n1839));
Q_AN02 U2711 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[59]), .Z(n1840));
Q_AN02 U2712 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[58]), .Z(n1841));
Q_AN02 U2713 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[57]), .Z(n1842));
Q_AN02 U2714 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[56]), .Z(n1843));
Q_AN02 U2715 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[55]), .Z(n1844));
Q_AN02 U2716 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[54]), .Z(n1845));
Q_AN02 U2717 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[53]), .Z(n1846));
Q_AN02 U2718 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[52]), .Z(n1847));
Q_AN02 U2719 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[51]), .Z(n1848));
Q_AN02 U2720 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[50]), .Z(n1849));
Q_AN02 U2721 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[49]), .Z(n1850));
Q_AN02 U2722 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[48]), .Z(n1851));
Q_AN02 U2723 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[47]), .Z(n1852));
Q_AN02 U2724 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[46]), .Z(n1853));
Q_AN02 U2725 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[45]), .Z(n1854));
Q_AN02 U2726 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[44]), .Z(n1855));
Q_AN02 U2727 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[43]), .Z(n1856));
Q_AN02 U2728 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[42]), .Z(n1857));
Q_AN02 U2729 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[41]), .Z(n1858));
Q_AN02 U2730 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[40]), .Z(n1859));
Q_AN02 U2731 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[39]), .Z(n1860));
Q_AN02 U2732 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[38]), .Z(n1861));
Q_AN02 U2733 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[37]), .Z(n1862));
Q_AN02 U2734 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[36]), .Z(n1863));
Q_AN02 U2735 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[35]), .Z(n1864));
Q_AN02 U2736 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[34]), .Z(n1865));
Q_AN02 U2737 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[33]), .Z(n1866));
Q_AN02 U2738 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[32]), .Z(n1867));
Q_AN02 U2739 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[31]), .Z(n1868));
Q_AN02 U2740 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[30]), .Z(n1869));
Q_AN02 U2741 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[29]), .Z(n1870));
Q_AN02 U2742 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[28]), .Z(n1871));
Q_AN02 U2743 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[27]), .Z(n1872));
Q_AN02 U2744 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[26]), .Z(n1873));
Q_AN02 U2745 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[25]), .Z(n1874));
Q_AN02 U2746 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[24]), .Z(n1875));
Q_AN02 U2747 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[23]), .Z(n1876));
Q_AN02 U2748 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[22]), .Z(n1877));
Q_AN02 U2749 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[21]), .Z(n1878));
Q_AN02 U2750 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[20]), .Z(n1879));
Q_AN02 U2751 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[19]), .Z(n1880));
Q_AN02 U2752 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[18]), .Z(n1881));
Q_AN02 U2753 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[17]), .Z(n1882));
Q_AN02 U2754 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[16]), .Z(n1883));
Q_AN02 U2755 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[15]), .Z(n1884));
Q_AN02 U2756 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[14]), .Z(n1885));
Q_AN02 U2757 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[13]), .Z(n1886));
Q_AN02 U2758 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[12]), .Z(n1887));
Q_AN02 U2759 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[11]), .Z(n1888));
Q_AN02 U2760 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[10]), .Z(n1889));
Q_AN02 U2761 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[9]), .Z(n1890));
Q_AN02 U2762 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[8]), .Z(n1891));
Q_AN02 U2763 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[7]), .Z(n1892));
Q_AN02 U2764 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[6]), .Z(n1893));
Q_AN02 U2765 ( .A0(n1192), .A1(cmdfifo_kdfstream_cmd[5]), .Z(n1894));
Q_AN02 U2766 ( .A0(n1192), .A1(iter3_kdf_key_size[31]), .Z(n1895));
Q_AN02 U2767 ( .A0(n1192), .A1(iter3_kdf_key_size[30]), .Z(n1896));
Q_AN02 U2768 ( .A0(n1192), .A1(iter3_kdf_key_size[29]), .Z(n1897));
Q_AN02 U2769 ( .A0(n1192), .A1(iter3_kdf_key_size[28]), .Z(n1898));
Q_AN02 U2770 ( .A0(n1192), .A1(iter3_kdf_key_size[27]), .Z(n1899));
Q_AN02 U2771 ( .A0(n1192), .A1(iter3_kdf_key_size[26]), .Z(n1900));
Q_AN02 U2772 ( .A0(n1192), .A1(iter3_kdf_key_size[25]), .Z(n1901));
Q_AN02 U2773 ( .A0(n1192), .A1(iter3_kdf_key_size[24]), .Z(n1902));
Q_AN02 U2774 ( .A0(n1192), .A1(iter3_kdf_key_size[23]), .Z(n1903));
Q_AN02 U2775 ( .A0(n1192), .A1(iter3_kdf_key_size[22]), .Z(n1904));
Q_AN02 U2776 ( .A0(n1192), .A1(iter3_kdf_key_size[21]), .Z(n1905));
Q_AN02 U2777 ( .A0(n1192), .A1(iter3_kdf_key_size[20]), .Z(n1906));
Q_AN02 U2778 ( .A0(n1192), .A1(iter3_kdf_key_size[19]), .Z(n1907));
Q_AN02 U2779 ( .A0(n1192), .A1(iter3_kdf_key_size[18]), .Z(n1908));
Q_AN02 U2780 ( .A0(n1192), .A1(iter3_kdf_key_size[17]), .Z(n1909));
Q_AN02 U2781 ( .A0(n1192), .A1(iter3_kdf_key_size[16]), .Z(n1910));
Q_AN02 U2782 ( .A0(n1192), .A1(iter3_kdf_key_size[15]), .Z(n1911));
Q_AN02 U2783 ( .A0(n1192), .A1(iter3_kdf_key_size[14]), .Z(n1912));
Q_AN02 U2784 ( .A0(n1192), .A1(iter3_kdf_key_size[13]), .Z(n1913));
Q_AN02 U2785 ( .A0(n1192), .A1(iter3_kdf_key_size[12]), .Z(n1914));
Q_AN02 U2786 ( .A0(n1192), .A1(iter3_kdf_key_size[11]), .Z(n1915));
Q_AN02 U2787 ( .A0(n1192), .A1(iter3_kdf_key_size[10]), .Z(n1916));
Q_AN02 U2788 ( .A0(n1192), .A1(n1918), .Z(n1917));
Q_MX02 U2789 ( .S(n1190), .A0(iter3_kdf_key_size[9]), .A1(iter1_kdf_key_size[9]), .Z(n1918));
Q_AN02 U2790 ( .A0(n1192), .A1(n1920), .Z(n1919));
Q_MX02 U2791 ( .S(n2038), .A0(iter2_kdf_key_size[8]), .A1(iter3_kdf_key_size[8]), .Z(n1920));
Q_AN02 U2792 ( .A0(n1192), .A1(iter3_kdf_key_size[7]), .Z(n1921));
Q_AN02 U2793 ( .A0(n1192), .A1(iter3_kdf_key_size[6]), .Z(n1922));
Q_AN02 U2794 ( .A0(n1192), .A1(iter3_kdf_key_size[5]), .Z(n1923));
Q_AN02 U2795 ( .A0(n1192), .A1(iter3_kdf_key_size[4]), .Z(n1924));
Q_AN02 U2796 ( .A0(n1192), .A1(iter3_kdf_key_size[3]), .Z(n1925));
Q_AN02 U2797 ( .A0(n1192), .A1(iter3_kdf_key_size[2]), .Z(n1926));
Q_AN02 U2798 ( .A0(n1192), .A1(iter3_kdf_key_size[1]), .Z(n1927));
Q_AN02 U2799 ( .A0(n1192), .A1(iter3_kdf_key_size[0]), .Z(n1928));
Q_MX02 U2800 ( .S(n1192), .A0(n1930), .A1(cmdfifo_kdfstream_cmd[260]), .Z(n1929));
Q_AN02 U2801 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[132]), .Z(n1930));
Q_MX02 U2802 ( .S(n1192), .A0(n1932), .A1(cmdfifo_kdfstream_cmd[259]), .Z(n1931));
Q_AN02 U2803 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[131]), .Z(n1932));
Q_MX02 U2804 ( .S(n1192), .A0(n1934), .A1(cmdfifo_kdfstream_cmd[258]), .Z(n1933));
Q_AN02 U2805 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[130]), .Z(n1934));
Q_MX02 U2806 ( .S(n1192), .A0(n1936), .A1(cmdfifo_kdfstream_cmd[257]), .Z(n1935));
Q_AN02 U2807 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[129]), .Z(n1936));
Q_MX02 U2808 ( .S(n1192), .A0(n1938), .A1(cmdfifo_kdfstream_cmd[256]), .Z(n1937));
Q_AN02 U2809 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[128]), .Z(n1938));
Q_MX02 U2810 ( .S(n1192), .A0(n1940), .A1(cmdfifo_kdfstream_cmd[255]), .Z(n1939));
Q_AN02 U2811 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[127]), .Z(n1940));
Q_MX02 U2812 ( .S(n1192), .A0(n1942), .A1(cmdfifo_kdfstream_cmd[254]), .Z(n1941));
Q_AN02 U2813 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[126]), .Z(n1942));
Q_MX02 U2814 ( .S(n1192), .A0(n1944), .A1(cmdfifo_kdfstream_cmd[253]), .Z(n1943));
Q_AN02 U2815 ( .A0(n1193), .A1(cmdfifo_kdfstream_cmd[125]), .Z(n1944));
Q_OR02 U2816 ( .A0(nxt_state[0]), .A1(nxt_state[1]), .Z(n1945));
Q_INV U2817 ( .A(in_hash_eof), .Z(n1946));
Q_ND02 U2818 ( .A0(n1946), .A1(n1945), .Z(n1947));
Q_AN02 U2819 ( .A0(n1945), .A1(n1950), .Z(n1948));
Q_ND02 U2820 ( .A0(n1945), .A1(iter_num[0]), .Z(n1949));
Q_XOR2 U2821 ( .A0(iter_num[1]), .A1(iter_num[0]), .Z(n1950));
Q_INV U2822 ( .A(kdfstream_cmdfifo_ack), .Z(n1952));
Q_AN02 U2823 ( .A0(n1952), .A1(in_hash_eof), .Z(n1956));
Q_OR02 U2824 ( .A0(n1956), .A1(kdfstream_cmdfifo_ack), .Z(n1954));
Q_AN02 U2825 ( .A0(n1953), .A1(cur_state[0]), .Z(st_tx_data));
Q_ND02 U2826 ( .A0(st_tx_data), .A1(n1954), .Z(n1955));
Q_OA21 U2827 ( .A0(cur_state[1]), .A1(cmdfifo_kdfstream_valid), .B0(n1957), .Z(n1958));
Q_AO21 U2828 ( .A0(st_tx_data), .A1(n1956), .B0(n1958), .Z(n1959));
Q_NR02 U2829 ( .A0(cur_state[0]), .A1(hash_cmd_in_stall[0]), .Z(n1957));
Q_INV U2830 ( .A(n1959), .Z(n1951));
Q_MX02 U2831 ( .S(n1955), .A0(n1959), .A1(n1960), .Z(nxt_state[1]));
Q_AN02 U2832 ( .A0(n1951), .A1(cur_state[1]), .Z(n1960));
Q_OA21 U2833 ( .A0(n1959), .A1(cur_state[0]), .B0(n1955), .Z(nxt_state[0]));
Q_FDP1 \cur_state_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_state[1]), .Q(cur_state[1]), .QN(n1953));
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN( ));
Q_AN02 U2836 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[31]), .Z(iter2_kdf_key_size[31]));
Q_AN02 U2837 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[30]), .Z(iter2_kdf_key_size[30]));
Q_AN02 U2838 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[29]), .Z(iter2_kdf_key_size[29]));
Q_AN02 U2839 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[28]), .Z(iter2_kdf_key_size[28]));
Q_AN02 U2840 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[27]), .Z(iter2_kdf_key_size[27]));
Q_AN02 U2841 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[26]), .Z(iter2_kdf_key_size[26]));
Q_AN02 U2842 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[25]), .Z(iter2_kdf_key_size[25]));
Q_AN02 U2843 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[24]), .Z(iter2_kdf_key_size[24]));
Q_AN02 U2844 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[23]), .Z(iter1_kdf_key_size[23]));
Q_AN02 U2845 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[22]), .Z(iter2_kdf_key_size[22]));
Q_AN02 U2846 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[21]), .Z(iter1_kdf_key_size[21]));
Q_AN02 U2847 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[20]), .Z(iter1_kdf_key_size[20]));
Q_AN02 U2848 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[19]), .Z(iter1_kdf_key_size[19]));
Q_AN02 U2849 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[18]), .Z(iter1_kdf_key_size[18]));
Q_AN02 U2850 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[17]), .Z(iter2_kdf_key_size[17]));
Q_AN02 U2851 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[16]), .Z(iter2_kdf_key_size[16]));
Q_AN02 U2852 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[15]), .Z(iter1_kdf_key_size[15]));
Q_AN02 U2853 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[14]), .Z(iter2_kdf_key_size[14]));
Q_AN02 U2854 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[13]), .Z(iter1_kdf_key_size[13]));
Q_AN02 U2855 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[12]), .Z(iter2_kdf_key_size[12]));
Q_AN02 U2856 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[11]), .Z(iter2_kdf_key_size[11]));
Q_AN02 U2857 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[10]), .Z(iter1_kdf_key_size[10]));
Q_OR02 U2858 ( .A0(n1961), .A1(kdf_test_key_size[9]), .Z(iter2_kdf_key_size[9]));
Q_OR02 U2859 ( .A0(n1961), .A1(kdf_test_key_size[8]), .Z(iter1_kdf_key_size[8]));
Q_INV U2860 ( .A(kdf_test_mode_en), .Z(n1961));
Q_AN02 U2861 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[7]), .Z(iter2_kdf_key_size[7]));
Q_AN02 U2862 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[6]), .Z(iter2_kdf_key_size[6]));
Q_AN02 U2863 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[5]), .Z(iter1_kdf_key_size[5]));
Q_AN02 U2864 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[4]), .Z(iter1_kdf_key_size[4]));
Q_AN02 U2865 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[3]), .Z(iter2_kdf_key_size[3]));
Q_AN02 U2866 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[2]), .Z(iter2_kdf_key_size[2]));
Q_AN02 U2867 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[1]), .Z(iter1_kdf_key_size[1]));
Q_AN02 U2868 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[0]), .Z(iter2_kdf_key_size[0]));
Q_AN02 U2869 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[8]), .Z(iter2_kdf_key_size[8]));
Q_AN02 U2870 ( .A0(kdf_test_mode_en), .A1(kdf_test_key_size[9]), .Z(iter1_kdf_key_size[9]));
Q_INV U2871 ( .A(nxt_state[1]), .Z(n1969));
Q_AN03 U2872 ( .A0(nxt_state[0]), .A1(n1969), .A2(cmd_il_valid), .Z(moving_to_tx_data));
Q_AD02 U2873 ( .CI(n1962), .A0(cmd_il_data_size[4]), .A1(cmd_il_data_size[5]), .B0(cmd_dgl_data_size[4]), .B1(cmd_dgl_data_size[5]), .S0(total_hash_size[4]), .S1(total_hash_size[5]), .CO(total_hash_size[6]));
Q_OA21 U2874 ( .A0(hash_cmd_in[8]), .A1(hash_cmd_in[7]), .B0(hash_cmd_in[11]), .Z(n1968));
Q_AO21 U2875 ( .A0(hash_cmd_in[11]), .A1(hash_cmd_in[9]), .B0(n1968), .Z(n1967));
Q_OR03 U2876 ( .A0(hash_cmd_in[6]), .A1(hash_cmd_in[5]), .A2(hash_cmd_in[4]), .Z(n1966));
Q_AO21 U2877 ( .A0(hash_cmd_in[11]), .A1(n1966), .B0(n1967), .Z(n1965));
Q_INV U2878 ( .A(n1965), .Z(is_small_size));
Q_AD02 U2879 ( .CI(n1963), .A0(cmd_il_data_size[2]), .A1(cmd_il_data_size[3]), .B0(cmd_il_valid), .B1(cmd_dgl_data_size[3]), .S0(total_hash_size[2]), .S1(total_hash_size[3]), .CO(n1962));
ixc_assign _zz_strnp_0 ( cmdfifo_hash_valid, fifo_out_valid[0]);
ixc_assign _zz_strnp_1 ( cmdfifo_hash_skip, fifo_out[33]);
ixc_assign _zz_strnp_2 ( cmdfifo_hash_small_size, fifo_out[0]);
ixc_assign _zz_strnp_3 ( hash_len_data_out_valid, fifo_out_valid[0]);
ixc_assign_32 _zz_strnp_4 ( hash_len_data_out[31:0], fifo_out[32:1]);
ixc_assign _zz_strnp_5 ( fifo_out_ack[0], hash_cmdfifo_ack);
ixc_assign _zz_strnp_6 ( _zy_simnet_kdfstream_cmdfifo_ack_0_w$, 
	kdfstream_cmdfifo_ack);
ixc_assign _zz_strnp_7 ( _zy_simnet_cmdfifo_hash_valid_1_w$, 
	cmdfifo_hash_valid);
ixc_assign _zz_strnp_8 ( _zy_simnet_cmdfifo_hash_skip_2_w$, cmdfifo_hash_skip);
ixc_assign _zz_strnp_9 ( _zy_simnet_cmdfifo_hash_small_size_3_w$, 
	cmdfifo_hash_small_size);
ixc_assign_32 _zz_strnp_10 ( _zy_simnet_hash_len_data_out_4_w$[0:31], 
	hash_len_data_out[31:0]);
ixc_assign _zz_strnp_11 ( _zy_simnet_hash_len_data_out_valid_5_w$, 
	hash_len_data_out_valid);
ixc_assign _zz_strnp_12 ( _zy_simnet_in_hash_valid_6_w$, in_hash_valid);
ixc_assign _zz_strnp_13 ( _zy_simnet_in_hash_eof_7_w$, in_hash_eof);
ixc_assign _zz_strnp_14 ( _zy_simnet_in_hash_eoc_8_w$, kdfstream_cmdfifo_ack);
ixc_assign_5 _zz_strnp_15 ( _zy_simnet_in_hash_num_bytes_9_w$[0:4], 
	in_hash_num_bytes[4:0]);
ixc_assign_128 _zz_strnp_16 ( _zy_simnet_in_hash_data_10_w$[0:127], 
	in_hash_data[127:0]);
ixc_assign _zz_strnp_17 ( _zy_simnet_cmd_il_valid_11_w$, cmd_il_valid);
ixc_assign_6 _zz_strnp_18 ( _zy_simnet_cmd_il_data_size_12_w$[0:5], 
	cmd_il_data_size[5:0]);
ixc_assign_288 _zz_strnp_19 ( _zy_simnet_cmd_il_data_13_w$[0:287], 
	cmd_il_data[287:0]);
ixc_assign _zz_strnp_20 ( _zy_simnet_pipe_array_ack_14_w$, 
	\pipe_array_ack[0][0] );
ixc_assign_5 _zz_strnp_21 ( _zy_simnet_pipe_array_ack_num_bytes_15_w$[0:4], { 
	\pipe_array_ack_num_bytes[0][4] , \pipe_array_ack_num_bytes[0][3] , 
	\pipe_array_ack_num_bytes[0][2] , \pipe_array_ack_num_bytes[0][1] , 
	\pipe_array_ack_num_bytes[0][0] });
ixc_assign _zz_strnp_22 ( _zy_simnet_cmd_dgl_valid_16_w$, cmd_il_valid);
ixc_assign_6 _zz_strnp_23 ( _zy_simnet_cmd_dgl_data_size_17_w$[0:5], { 
	cmd_dgl_data_size[5], cmd_dgl_data_size[4], cmd_dgl_data_size[3], 
	cmd_il_valid, cmd_dgl_data_size[1], cmd_dgl_data_size[0]});
ixc_assign_296 _zz_strnp_24 ( _zy_simnet_cmd_dgl_data_18_w$[0:295], 
	cmd_dgl_data[295:0]);
ixc_assign _zz_strnp_25 ( _zy_simnet_pipe_array_ack_19_w$, 
	\pipe_array_ack[1][0] );
ixc_assign_5 _zz_strnp_26 ( _zy_simnet_pipe_array_ack_num_bytes_20_w$[0:4], { 
	\pipe_array_ack_num_bytes[1][4] , \pipe_array_ack_num_bytes[1][3] , 
	\pipe_array_ack_num_bytes[1][2] , \pipe_array_ack_num_bytes[1][1] , 
	\pipe_array_ack_num_bytes[1][0] });
ixc_assign_34 _zz_strnp_27 ( _zy_simnet_hash_cmd_in_23_w$[0:33], 
	hash_cmd_in[33:0]);
ixc_assign _zz_strnp_28 ( _zy_simnet_hash_cmd_in_valid_24_w$, 
	hash_cmd_in_valid[0]);
cr_kme_kop_kdf_stream_pipe_xcm79 il_var ( .pipe_valid( 
	\pipe_array_valid[0][0] ), .pipe_data( { \pipe_array_data[0][127] , 
	\pipe_array_data[0][126] , \pipe_array_data[0][125] , 
	\pipe_array_data[0][124] , \pipe_array_data[0][123] , 
	\pipe_array_data[0][122] , \pipe_array_data[0][121] , 
	\pipe_array_data[0][120] , \pipe_array_data[0][119] , 
	\pipe_array_data[0][118] , \pipe_array_data[0][117] , 
	\pipe_array_data[0][116] , \pipe_array_data[0][115] , 
	\pipe_array_data[0][114] , \pipe_array_data[0][113] , 
	\pipe_array_data[0][112] , \pipe_array_data[0][111] , 
	\pipe_array_data[0][110] , \pipe_array_data[0][109] , 
	\pipe_array_data[0][108] , \pipe_array_data[0][107] , 
	\pipe_array_data[0][106] , \pipe_array_data[0][105] , 
	\pipe_array_data[0][104] , \pipe_array_data[0][103] , 
	\pipe_array_data[0][102] , \pipe_array_data[0][101] , 
	\pipe_array_data[0][100] , \pipe_array_data[0][99] , 
	\pipe_array_data[0][98] , \pipe_array_data[0][97] , 
	\pipe_array_data[0][96] , \pipe_array_data[0][95] , 
	\pipe_array_data[0][94] , \pipe_array_data[0][93] , 
	\pipe_array_data[0][92] , \pipe_array_data[0][91] , 
	\pipe_array_data[0][90] , \pipe_array_data[0][89] , 
	\pipe_array_data[0][88] , \pipe_array_data[0][87] , 
	\pipe_array_data[0][86] , \pipe_array_data[0][85] , 
	\pipe_array_data[0][84] , \pipe_array_data[0][83] , 
	\pipe_array_data[0][82] , \pipe_array_data[0][81] , 
	\pipe_array_data[0][80] , \pipe_array_data[0][79] , 
	\pipe_array_data[0][78] , \pipe_array_data[0][77] , 
	\pipe_array_data[0][76] , \pipe_array_data[0][75] , 
	\pipe_array_data[0][74] , \pipe_array_data[0][73] , 
	\pipe_array_data[0][72] , \pipe_array_data[0][71] , 
	\pipe_array_data[0][70] , \pipe_array_data[0][69] , 
	\pipe_array_data[0][68] , \pipe_array_data[0][67] , 
	\pipe_array_data[0][66] , \pipe_array_data[0][65] , 
	\pipe_array_data[0][64] , \pipe_array_data[0][63] , 
	\pipe_array_data[0][62] , \pipe_array_data[0][61] , 
	\pipe_array_data[0][60] , \pipe_array_data[0][59] , 
	\pipe_array_data[0][58] , \pipe_array_data[0][57] , 
	\pipe_array_data[0][56] , \pipe_array_data[0][55] , 
	\pipe_array_data[0][54] , \pipe_array_data[0][53] , 
	\pipe_array_data[0][52] , \pipe_array_data[0][51] , 
	\pipe_array_data[0][50] , \pipe_array_data[0][49] , 
	\pipe_array_data[0][48] , \pipe_array_data[0][47] , 
	\pipe_array_data[0][46] , \pipe_array_data[0][45] , 
	\pipe_array_data[0][44] , \pipe_array_data[0][43] , 
	\pipe_array_data[0][42] , \pipe_array_data[0][41] , 
	\pipe_array_data[0][40] , \pipe_array_data[0][39] , 
	\pipe_array_data[0][38] , \pipe_array_data[0][37] , 
	\pipe_array_data[0][36] , \pipe_array_data[0][35] , 
	\pipe_array_data[0][34] , \pipe_array_data[0][33] , 
	\pipe_array_data[0][32] , \pipe_array_data[0][31] , 
	\pipe_array_data[0][30] , \pipe_array_data[0][29] , 
	\pipe_array_data[0][28] , \pipe_array_data[0][27] , 
	\pipe_array_data[0][26] , \pipe_array_data[0][25] , 
	\pipe_array_data[0][24] , \pipe_array_data[0][23] , 
	\pipe_array_data[0][22] , \pipe_array_data[0][21] , 
	\pipe_array_data[0][20] , \pipe_array_data[0][19] , 
	\pipe_array_data[0][18] , \pipe_array_data[0][17] , 
	\pipe_array_data[0][16] , \pipe_array_data[0][15] , 
	\pipe_array_data[0][14] , \pipe_array_data[0][13] , 
	\pipe_array_data[0][12] , \pipe_array_data[0][11] , 
	\pipe_array_data[0][10] , \pipe_array_data[0][9] , 
	\pipe_array_data[0][8] , \pipe_array_data[0][7] , 
	\pipe_array_data[0][6] , \pipe_array_data[0][5] , 
	\pipe_array_data[0][4] , \pipe_array_data[0][3] , 
	\pipe_array_data[0][2] , \pipe_array_data[0][1] , 
	\pipe_array_data[0][0] }), .pipe_byte_count( { 
	\pipe_array_byte_count[0][5] , \pipe_array_byte_count[0][4] , 
	\pipe_array_byte_count[0][3] , \pipe_array_byte_count[0][2] , 
	\pipe_array_byte_count[0][1] , \pipe_array_byte_count[0][0] }), 
	.clk( clk), .rst_n( rst_n), .cmd_valid( 
	_zy_simnet_cmd_il_valid_11_w$), .cmd_data_size( 
	_zy_simnet_cmd_il_data_size_12_w$[0:5]), .cmd_data( 
	_zy_simnet_cmd_il_data_13_w$[0:287]), .pipe_ack( 
	_zy_simnet_pipe_array_ack_14_w$), .pipe_ack_num_bytes( 
	_zy_simnet_pipe_array_ack_num_bytes_15_w$[0:4]));
cr_kme_kop_kdf_stream_pipe_xcm78 dgl_var ( .pipe_valid( 
	\pipe_array_valid[1][0] ), .pipe_data( { \pipe_array_data[1][127] , 
	\pipe_array_data[1][126] , \pipe_array_data[1][125] , 
	\pipe_array_data[1][124] , \pipe_array_data[1][123] , 
	\pipe_array_data[1][122] , \pipe_array_data[1][121] , 
	\pipe_array_data[1][120] , \pipe_array_data[1][119] , 
	\pipe_array_data[1][118] , \pipe_array_data[1][117] , 
	\pipe_array_data[1][116] , \pipe_array_data[1][115] , 
	\pipe_array_data[1][114] , \pipe_array_data[1][113] , 
	\pipe_array_data[1][112] , \pipe_array_data[1][111] , 
	\pipe_array_data[1][110] , \pipe_array_data[1][109] , 
	\pipe_array_data[1][108] , \pipe_array_data[1][107] , 
	\pipe_array_data[1][106] , \pipe_array_data[1][105] , 
	\pipe_array_data[1][104] , \pipe_array_data[1][103] , 
	\pipe_array_data[1][102] , \pipe_array_data[1][101] , 
	\pipe_array_data[1][100] , \pipe_array_data[1][99] , 
	\pipe_array_data[1][98] , \pipe_array_data[1][97] , 
	\pipe_array_data[1][96] , \pipe_array_data[1][95] , 
	\pipe_array_data[1][94] , \pipe_array_data[1][93] , 
	\pipe_array_data[1][92] , \pipe_array_data[1][91] , 
	\pipe_array_data[1][90] , \pipe_array_data[1][89] , 
	\pipe_array_data[1][88] , \pipe_array_data[1][87] , 
	\pipe_array_data[1][86] , \pipe_array_data[1][85] , 
	\pipe_array_data[1][84] , \pipe_array_data[1][83] , 
	\pipe_array_data[1][82] , \pipe_array_data[1][81] , 
	\pipe_array_data[1][80] , \pipe_array_data[1][79] , 
	\pipe_array_data[1][78] , \pipe_array_data[1][77] , 
	\pipe_array_data[1][76] , \pipe_array_data[1][75] , 
	\pipe_array_data[1][74] , \pipe_array_data[1][73] , 
	\pipe_array_data[1][72] , \pipe_array_data[1][71] , 
	\pipe_array_data[1][70] , \pipe_array_data[1][69] , 
	\pipe_array_data[1][68] , \pipe_array_data[1][67] , 
	\pipe_array_data[1][66] , \pipe_array_data[1][65] , 
	\pipe_array_data[1][64] , \pipe_array_data[1][63] , 
	\pipe_array_data[1][62] , \pipe_array_data[1][61] , 
	\pipe_array_data[1][60] , \pipe_array_data[1][59] , 
	\pipe_array_data[1][58] , \pipe_array_data[1][57] , 
	\pipe_array_data[1][56] , \pipe_array_data[1][55] , 
	\pipe_array_data[1][54] , \pipe_array_data[1][53] , 
	\pipe_array_data[1][52] , \pipe_array_data[1][51] , 
	\pipe_array_data[1][50] , \pipe_array_data[1][49] , 
	\pipe_array_data[1][48] , \pipe_array_data[1][47] , 
	\pipe_array_data[1][46] , \pipe_array_data[1][45] , 
	\pipe_array_data[1][44] , \pipe_array_data[1][43] , 
	\pipe_array_data[1][42] , \pipe_array_data[1][41] , 
	\pipe_array_data[1][40] , \pipe_array_data[1][39] , 
	\pipe_array_data[1][38] , \pipe_array_data[1][37] , 
	\pipe_array_data[1][36] , \pipe_array_data[1][35] , 
	\pipe_array_data[1][34] , \pipe_array_data[1][33] , 
	\pipe_array_data[1][32] , \pipe_array_data[1][31] , 
	\pipe_array_data[1][30] , \pipe_array_data[1][29] , 
	\pipe_array_data[1][28] , \pipe_array_data[1][27] , 
	\pipe_array_data[1][26] , \pipe_array_data[1][25] , 
	\pipe_array_data[1][24] , \pipe_array_data[1][23] , 
	\pipe_array_data[1][22] , \pipe_array_data[1][21] , 
	\pipe_array_data[1][20] , \pipe_array_data[1][19] , 
	\pipe_array_data[1][18] , \pipe_array_data[1][17] , 
	\pipe_array_data[1][16] , \pipe_array_data[1][15] , 
	\pipe_array_data[1][14] , \pipe_array_data[1][13] , 
	\pipe_array_data[1][12] , \pipe_array_data[1][11] , 
	\pipe_array_data[1][10] , \pipe_array_data[1][9] , 
	\pipe_array_data[1][8] , \pipe_array_data[1][7] , 
	\pipe_array_data[1][6] , \pipe_array_data[1][5] , 
	\pipe_array_data[1][4] , \pipe_array_data[1][3] , 
	\pipe_array_data[1][2] , \pipe_array_data[1][1] , 
	\pipe_array_data[1][0] }), .pipe_byte_count( { 
	\pipe_array_byte_count[1][5] , \pipe_array_byte_count[1][4] , 
	\pipe_array_byte_count[1][3] , \pipe_array_byte_count[1][2] , 
	\pipe_array_byte_count[1][1] , \pipe_array_byte_count[1][0] }), 
	.clk( clk), .rst_n( rst_n), .cmd_valid( 
	_zy_simnet_cmd_dgl_valid_16_w$), .cmd_data_size( 
	_zy_simnet_cmd_dgl_data_size_17_w$[0:5]), .cmd_data( 
	_zy_simnet_cmd_dgl_data_18_w$[0:295]), .pipe_ack( 
	_zy_simnet_pipe_array_ack_19_w$), .pipe_ack_num_bytes( 
	_zy_simnet_pipe_array_ack_num_bytes_20_w$[0:4]));
cr_kme_fifo_xcm52 parser_fifo ( .fifo_in_stall( hash_cmd_in_stall[0]), 
	.fifo_out( fifo_out[33:0]), .fifo_out_valid( fifo_out_valid[0]), 
	.fifo_overflow( _zy_simnet_dio_21), .fifo_underflow( 
	_zy_simnet_dio_22), .clk( clk), .rst_n( rst_n), .fifo_in( 
	_zy_simnet_hash_cmd_in_23_w$[0:33]), .fifo_in_valid( 
	_zy_simnet_hash_cmd_in_valid_24_w$), .fifo_out_ack( fifo_out_ack[0]), 
	.fifo_in_stall_override( _zy_simnet_cio_25));
Q_INV U2912 ( .A(n1101), .Z(n1970));
Q_INV U2913 ( .A(n1136), .Z(n1971));
Q_OR02 U2914 ( .A0(n1191), .A1(n1190), .Z(n1972));
Q_AO21 U2915 ( .A0(n345), .A1(\pipe_array_ack[1][0] ), .B0(n949), .Z(in_hash_data[64]));
Q_AO21 U2916 ( .A0(n344), .A1(\pipe_array_ack[1][0] ), .B0(n948), .Z(in_hash_data[65]));
Q_AO21 U2917 ( .A0(n343), .A1(\pipe_array_ack[1][0] ), .B0(n947), .Z(in_hash_data[66]));
Q_AO21 U2918 ( .A0(n342), .A1(\pipe_array_ack[1][0] ), .B0(n946), .Z(in_hash_data[67]));
Q_AO21 U2919 ( .A0(n341), .A1(\pipe_array_ack[1][0] ), .B0(n945), .Z(in_hash_data[68]));
Q_AO21 U2920 ( .A0(n340), .A1(\pipe_array_ack[1][0] ), .B0(n944), .Z(in_hash_data[69]));
Q_AO21 U2921 ( .A0(n339), .A1(\pipe_array_ack[1][0] ), .B0(n943), .Z(in_hash_data[70]));
Q_AO21 U2922 ( .A0(n338), .A1(\pipe_array_ack[1][0] ), .B0(n942), .Z(in_hash_data[71]));
Q_AO21 U2923 ( .A0(n337), .A1(\pipe_array_ack[1][0] ), .B0(n941), .Z(in_hash_data[72]));
Q_AO21 U2924 ( .A0(n336), .A1(\pipe_array_ack[1][0] ), .B0(n940), .Z(in_hash_data[73]));
Q_AO21 U2925 ( .A0(n335), .A1(\pipe_array_ack[1][0] ), .B0(n939), .Z(in_hash_data[74]));
Q_AO21 U2926 ( .A0(n334), .A1(\pipe_array_ack[1][0] ), .B0(n938), .Z(in_hash_data[75]));
Q_AO21 U2927 ( .A0(n333), .A1(\pipe_array_ack[1][0] ), .B0(n937), .Z(in_hash_data[76]));
Q_AO21 U2928 ( .A0(n332), .A1(\pipe_array_ack[1][0] ), .B0(n936), .Z(in_hash_data[77]));
Q_AO21 U2929 ( .A0(n331), .A1(\pipe_array_ack[1][0] ), .B0(n935), .Z(in_hash_data[78]));
Q_AO21 U2930 ( .A0(n330), .A1(\pipe_array_ack[1][0] ), .B0(n934), .Z(in_hash_data[79]));
Q_AO21 U2931 ( .A0(n329), .A1(\pipe_array_ack[1][0] ), .B0(n933), .Z(in_hash_data[80]));
Q_AO21 U2932 ( .A0(n328), .A1(\pipe_array_ack[1][0] ), .B0(n932), .Z(in_hash_data[81]));
Q_AO21 U2933 ( .A0(n327), .A1(\pipe_array_ack[1][0] ), .B0(n931), .Z(in_hash_data[82]));
Q_AO21 U2934 ( .A0(n326), .A1(\pipe_array_ack[1][0] ), .B0(n930), .Z(in_hash_data[83]));
Q_AO21 U2935 ( .A0(n325), .A1(\pipe_array_ack[1][0] ), .B0(n929), .Z(in_hash_data[84]));
Q_AO21 U2936 ( .A0(n324), .A1(\pipe_array_ack[1][0] ), .B0(n928), .Z(in_hash_data[85]));
Q_AO21 U2937 ( .A0(n323), .A1(\pipe_array_ack[1][0] ), .B0(n927), .Z(in_hash_data[86]));
Q_AO21 U2938 ( .A0(n322), .A1(\pipe_array_ack[1][0] ), .B0(n926), .Z(in_hash_data[87]));
Q_AO21 U2939 ( .A0(n321), .A1(\pipe_array_ack[1][0] ), .B0(n925), .Z(in_hash_data[88]));
Q_AO21 U2940 ( .A0(n320), .A1(\pipe_array_ack[1][0] ), .B0(n924), .Z(in_hash_data[89]));
Q_AO21 U2941 ( .A0(n319), .A1(\pipe_array_ack[1][0] ), .B0(n923), .Z(in_hash_data[90]));
Q_AO21 U2942 ( .A0(n318), .A1(\pipe_array_ack[1][0] ), .B0(n922), .Z(in_hash_data[91]));
Q_AO21 U2943 ( .A0(n317), .A1(\pipe_array_ack[1][0] ), .B0(n921), .Z(in_hash_data[92]));
Q_AO21 U2944 ( .A0(n316), .A1(\pipe_array_ack[1][0] ), .B0(n920), .Z(in_hash_data[93]));
Q_AO21 U2945 ( .A0(n315), .A1(\pipe_array_ack[1][0] ), .B0(n919), .Z(in_hash_data[94]));
Q_AO21 U2946 ( .A0(n314), .A1(\pipe_array_ack[1][0] ), .B0(n918), .Z(in_hash_data[95]));
Q_AO21 U2947 ( .A0(n313), .A1(\pipe_array_ack[1][0] ), .B0(n917), .Z(in_hash_data[96]));
Q_AO21 U2948 ( .A0(n312), .A1(\pipe_array_ack[1][0] ), .B0(n916), .Z(in_hash_data[97]));
Q_AO21 U2949 ( .A0(n311), .A1(\pipe_array_ack[1][0] ), .B0(n915), .Z(in_hash_data[98]));
Q_AO21 U2950 ( .A0(n310), .A1(\pipe_array_ack[1][0] ), .B0(n914), .Z(in_hash_data[99]));
Q_AO21 U2951 ( .A0(n309), .A1(\pipe_array_ack[1][0] ), .B0(n913), .Z(in_hash_data[100]));
Q_AO21 U2952 ( .A0(n308), .A1(\pipe_array_ack[1][0] ), .B0(n912), .Z(in_hash_data[101]));
Q_AO21 U2953 ( .A0(n307), .A1(\pipe_array_ack[1][0] ), .B0(n911), .Z(in_hash_data[102]));
Q_AO21 U2954 ( .A0(n306), .A1(\pipe_array_ack[1][0] ), .B0(n910), .Z(in_hash_data[103]));
Q_AO21 U2955 ( .A0(n305), .A1(\pipe_array_ack[1][0] ), .B0(n909), .Z(in_hash_data[104]));
Q_AO21 U2956 ( .A0(n304), .A1(\pipe_array_ack[1][0] ), .B0(n908), .Z(in_hash_data[105]));
Q_AO21 U2957 ( .A0(n303), .A1(\pipe_array_ack[1][0] ), .B0(n907), .Z(in_hash_data[106]));
Q_AO21 U2958 ( .A0(n302), .A1(\pipe_array_ack[1][0] ), .B0(n906), .Z(in_hash_data[107]));
Q_AO21 U2959 ( .A0(n301), .A1(\pipe_array_ack[1][0] ), .B0(n905), .Z(in_hash_data[108]));
Q_AO21 U2960 ( .A0(n300), .A1(\pipe_array_ack[1][0] ), .B0(n904), .Z(in_hash_data[109]));
Q_AO21 U2961 ( .A0(n299), .A1(\pipe_array_ack[1][0] ), .B0(n903), .Z(in_hash_data[110]));
Q_AO21 U2962 ( .A0(n298), .A1(\pipe_array_ack[1][0] ), .B0(n902), .Z(in_hash_data[111]));
Q_AO21 U2963 ( .A0(n297), .A1(\pipe_array_ack[1][0] ), .B0(n901), .Z(in_hash_data[112]));
Q_AO21 U2964 ( .A0(n296), .A1(\pipe_array_ack[1][0] ), .B0(n900), .Z(in_hash_data[113]));
Q_AO21 U2965 ( .A0(n295), .A1(\pipe_array_ack[1][0] ), .B0(n899), .Z(in_hash_data[114]));
Q_AO21 U2966 ( .A0(n294), .A1(\pipe_array_ack[1][0] ), .B0(n898), .Z(in_hash_data[115]));
Q_AO21 U2967 ( .A0(n293), .A1(\pipe_array_ack[1][0] ), .B0(n897), .Z(in_hash_data[116]));
Q_AO21 U2968 ( .A0(n292), .A1(\pipe_array_ack[1][0] ), .B0(n896), .Z(in_hash_data[117]));
Q_AO21 U2969 ( .A0(n291), .A1(\pipe_array_ack[1][0] ), .B0(n895), .Z(in_hash_data[118]));
Q_AO21 U2970 ( .A0(n290), .A1(\pipe_array_ack[1][0] ), .B0(n894), .Z(in_hash_data[119]));
Q_AO21 U2971 ( .A0(n289), .A1(\pipe_array_ack[1][0] ), .B0(n893), .Z(in_hash_data[120]));
Q_AO21 U2972 ( .A0(n288), .A1(\pipe_array_ack[1][0] ), .B0(n892), .Z(in_hash_data[121]));
Q_AO21 U2973 ( .A0(n287), .A1(\pipe_array_ack[1][0] ), .B0(n891), .Z(in_hash_data[122]));
Q_AO21 U2974 ( .A0(n286), .A1(\pipe_array_ack[1][0] ), .B0(n890), .Z(in_hash_data[123]));
Q_AO21 U2975 ( .A0(n285), .A1(\pipe_array_ack[1][0] ), .B0(n889), .Z(in_hash_data[124]));
Q_AO21 U2976 ( .A0(n284), .A1(\pipe_array_ack[1][0] ), .B0(n888), .Z(in_hash_data[125]));
Q_AO21 U2977 ( .A0(n283), .A1(\pipe_array_ack[1][0] ), .B0(n887), .Z(in_hash_data[126]));
Q_AO21 U2978 ( .A0(n282), .A1(\pipe_array_ack[1][0] ), .B0(n886), .Z(in_hash_data[127]));
Q_INV U2979 ( .A(n1191), .Z(n2037));
Q_OR02 U2980 ( .A0(n2037), .A1(n1190), .Z(n2038));
Q_AN02 U2981 ( .A0(cmd_il_data_size[0]), .A1(cmd_dgl_data_size[0]), .Z(n1964));
Q_XOR2 U2982 ( .A0(cmd_il_data_size[0]), .A1(cmd_dgl_data_size[0]), .Z(total_hash_size[0]));
Q_XNR3 U2983 ( .A0(n1125), .A1(\pipe_array_byte_count[0][1] ), .A2(n1056), .Z(n1124));
Q_FDP4EP \iter_num_REG[1] ( .CK(clk), .CE(n1947), .R(n2039), .D(n1948), .Q(iter_num[1]));
Q_INV U2985 ( .A(rst_n), .Z(n2039));
Q_FDP4EP \iter_num_REG[0] ( .CK(clk), .CE(n1947), .R(n2039), .D(n1949), .Q(iter_num[0]));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "pipe_array_valid 1 0 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "pipe_array_data 1 127 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "pipe_array_byte_count 1 5 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m4 "pipe_array_ack 1 0 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m5 "pipe_array_ack_num_bytes 1 4 0 1 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "5"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\cmdfifo_kdfstream_cmd.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\cmdfifo_kdfstream_cmd.skip  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\cmdfifo_kdfstream_cmd.guid  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\cmdfifo_kdfstream_cmd.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\cmdfifo_kdfstream_cmd.num_iter  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\labels%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\labels%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\labels%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\labels%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\labels%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "labels (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "11"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "cmdfifo_kdfstream_cmd 5 \cmdfifo_kdfstream_cmd.combo_mode  \cmdfifo_kdfstream_cmd.skip  \cmdfifo_kdfstream_cmd.guid  \cmdfifo_kdfstream_cmd.label_index  \cmdfifo_kdfstream_cmd.num_iter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "labels%s 5 \labels%s.guid_size  \labels%s.label_size  \labels%s.label  \labels%s.delimiter_valid  \labels%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "2"
endmodule
