
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module apb_xactor ( psel, penable, paddr, pwdata, pwrite, clk, reset_n, prdata, 
	pready, pslverr);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output psel;
output penable;
output [19:0] paddr;
output [31:0] pwdata;
output pwrite;
input clk;
input reset_n;
input [31:0] prdata;
input pready;
input pslverr;
wire _zy_simnet_psel_0_w$;
wire _zy_simnet_penable_1_w$;
wire [0:19] _zy_simnet_paddr_2_w$;
wire [0:31] _zy_simnet_pwdata_3_w$;
wire _zy_simnet_pwrite_4_w$;
wire _zyL94_iscX1c0_s;
wire [63:0] _zyL94_iscX1c0_i0;
wire _zyL61_iscX2c0_s;
wire [63:0] _zyL61_iscX2c0_i0;
wire [31:0] _zyL61_iscX2c0_i1;
wire _zyM3L94_pbcMevClk4;
wire _zyM3L94_pbcReq4;
wire _zyM3L94_pbcBusy4;
wire _zyM3L94_pbcWait4;
wire _zyM3L61_pbcMevClk9;
wire _zyM3L61_pbcReq9;
wire _zyM3L61_pbcBusy9;
wire _zyM3L61_pbcWait9;
wire _zzpready_M3L25_bcSv0;
wire [31:0] _zzprdata_M3L24_bcSv1;
wire _zzpslverr_M3L26_bcSv2;
wire _zzM3L46_bcP0_EnDNxt;
wire _zzM3L46_bcP0_DOn;
wire _zzM3L94_bcP1_EnDNxt;
wire _zzM3L94_bcP1_DOn;
wire _zzM3L61_bcP2_EnDNxt;
wire _zzM3L61_bcP2_DOn;
wire _zzbcOne;
wire _zzM3_bcBehEvalClk;
wire _zzM3_bcBehHalt;
wire _zzmdxOne;
wire _zzM3L46_mdxP0_EnNxt;
wire _zzM3L46_mdxP0_On;
wire _zzM3L94_mdxP1_EnNxt;
wire _zzM3L94_mdxP1_On;
wire _zzM3L61_mdxP2_EnNxt;
wire _zzM3L61_mdxP2_On;
wire [7:0] bus_timer;
wire _zyL94_iscX1c0_f;
wire _zyL94_iscX1c0_n;
wire [31:0] _zyL94_iscX1c0_o1;
wire _zyL94_iscX1c0_o2;
wire _zyL61_iscX2c0_f;
wire _zyL61_iscX2c0_n;
wire _zyL61_iscX2c0_o2;
wire [63:0] _zyaddr_L95_tfiV0_M3_pbcG0;
wire [31:0] _zydata_L96_tfiV1_M3_pbcG1;
wire _zyresponse_L97_tfiV2_M3_pbcG2;
wire [63:0] _zyaddr_L62_tfiV3_M3_pbcG3;
wire [31:0] _zydata_L63_tfiV4_M3_pbcG4;
wire _zyresponse_L64_tfiV5_M3_pbcG5;
wire _zyM3L94_pbcCapEn0;
wire _zyM3L104_pbcCapEn1;
wire _zyM3L110_pbcCapEn2;
wire _zyM3L121_pbcCapEn3;
wire _zyM3L61_pbcCapEn5;
wire _zyM3L73_pbcCapEn6;
wire _zyM3L79_pbcCapEn7;
wire _zyM3L90_pbcCapEn8;
wire [2:0] _zyM3L94_pbcFsm0_s;
wire _zyM3L94_pbcEn10;
wire [2:0] _zyM3L61_pbcFsm2_s;
wire _zyM3L61_pbcEn11;
wire _zzM3L46_bcP0_EnD;
wire [7:0] _zzM3L46_bcP0_bus_timer_wr0;
wire _zzM3L46_bcP0_bus_timer_Dwen0;
wire _zzM3L46_bcP0_bus_timer_DwenOn0;
wire [7:0] _zzM3L29_bus_timer_nbaTmp3;
wire _zzM3L94_bcP1_EnD;
wire [7:0] _zzM3L94_bcP1_bus_timer_wr0;
wire _zzM3L94_bcP1_bus_timer_Dwen0;
wire _zzM3L94_bcP1_bus_timer_DwenOn0;
wire [31:0] _zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1;
wire _zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_Dwen1;
wire _zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1;
wire [31:0] _zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4;
wire _zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_wr2;
wire _zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_Dwen2;
wire _zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_DwenOn2;
wire _zzM3L97__zyresponse_L97_tfiV2_M3_pbcG2_nbaTmp5;
wire _zzM3L61_bcP2_EnD;
wire [7:0] _zzM3L61_bcP2_bus_timer_wr0;
wire _zzM3L61_bcP2_bus_timer_Dwen0;
wire _zzM3L61_bcP2_bus_timer_DwenOn0;
wire _zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_wr1;
wire _zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_Dwen1;
wire _zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_DwenOn1;
wire _zzM3L64__zyresponse_L64_tfiV5_M3_pbcG5_nbaTmp6;
wire [7:0] _zzbus_timer_M3L29_bcSvLt7;
wire [31:0] _zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8;
wire _zz_zyresponse_L97_tfiV2_M3_pbcG2_M3_bcSvLt9;
wire _zz_zyresponse_L64_tfiV5_M3_pbcG5_M3_bcSvLt10;
wire [31:0] _zzM3_bcBehEval;
wire _zzM3L19_psel_mdxTmp0;
wire _zzM3L20_penable_mdxTmp1;
wire _zzM3L23_pwrite_mdxTmp2;
wire [19:0] _zzM3L21_paddr_mdxTmp3;
wire [31:0] _zzM3L22_pwdata_mdxTmp4;
wire _zzM3L46_mdxP0_En;
wire _zzM3L46_mdxP0_psel_wr0;
wire _zzM3L46_mdxP0_psel_Dwen0;
wire _zzM3L46_mdxP0_psel_DwenOn0;
wire _zzM3L46_mdxP0_penable_wr1;
wire _zzM3L46_mdxP0_penable_Dwen1;
wire _zzM3L46_mdxP0_penable_DwenOn1;
wire _zzM3L46_mdxP0_pwrite_wr2;
wire _zzM3L46_mdxP0_pwrite_Dwen2;
wire _zzM3L46_mdxP0_pwrite_DwenOn2;
wire [19:0] _zzM3L46_mdxP0_paddr_wr3;
wire _zzM3L46_mdxP0_paddr_Dwen3;
wire _zzM3L46_mdxP0_paddr_DwenOn3;
wire [31:0] _zzM3L46_mdxP0_pwdata_wr4;
wire _zzM3L46_mdxP0_pwdata_Dwen4;
wire _zzM3L46_mdxP0_pwdata_DwenOn4;
wire _zzM3L94_mdxP1_En;
wire _zzM3L94_mdxP1_psel_wr0;
wire _zzM3L94_mdxP1_psel_Dwen0;
wire _zzM3L94_mdxP1_psel_DwenOn0;
wire _zzM3L94_mdxP1_penable_wr1;
wire _zzM3L94_mdxP1_penable_Dwen1;
wire _zzM3L94_mdxP1_penable_DwenOn1;
wire _zzM3L94_mdxP1_pwrite_wr2;
wire _zzM3L94_mdxP1_pwrite_Dwen2;
wire _zzM3L94_mdxP1_pwrite_DwenOn2;
wire [19:0] _zzM3L94_mdxP1_paddr_wr3;
wire _zzM3L94_mdxP1_paddr_Dwen3;
wire _zzM3L94_mdxP1_paddr_DwenOn3;
wire _zzM3L61_mdxP2_En;
wire _zzM3L61_mdxP2_psel_wr0;
wire _zzM3L61_mdxP2_psel_Dwen0;
wire _zzM3L61_mdxP2_psel_DwenOn0;
wire _zzM3L61_mdxP2_penable_wr1;
wire _zzM3L61_mdxP2_penable_Dwen1;
wire _zzM3L61_mdxP2_penable_DwenOn1;
wire _zzM3L61_mdxP2_pwrite_wr2;
wire _zzM3L61_mdxP2_pwrite_Dwen2;
wire _zzM3L61_mdxP2_pwrite_DwenOn2;
wire [19:0] _zzM3L61_mdxP2_paddr_wr3;
wire _zzM3L61_mdxP2_paddr_Dwen3;
wire _zzM3L61_mdxP2_paddr_DwenOn3;
wire [31:0] _zzM3L61_mdxP2_pwdata_wr4;
wire _zzM3L61_mdxP2_pwdata_Dwen4;
wire _zzM3L61_mdxP2_pwdata_DwenOn4;
wire _zzpsel_M3L19_mdxSvLt5;
wire _zzpenable_M3L20_mdxSvLt6;
wire _zzpwrite_M3L23_mdxSvLt7;
wire [19:0] _zzpaddr_M3L21_mdxSvLt8;
wire [31:0] _zzpwdata_M3L22_mdxSvLt9;
supply1 n317;
supply1 n318;
supply0 n319;
supply0 n320;
supply0 n321;
supply0 n323;
supply0 n324;
Q_BUF U0 ( .A(n319), .Z(n1));
Q_AN02 U1 ( .A0(n23), .A1(n21), .Z(n2));
Q_INV U2 ( .A(_zzM3L61_mdxP2_pwdata_DwenOn4), .Z(n4));
Q_AN02 U3 ( .A0(_zzM3L46_mdxP0_pwdata_DwenOn4), .A1(n4), .Z(n3));
Q_LDP0 \pwdata_REG[0] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[0]), .Q(pwdata[0]), .QN( ));
Q_LDP0 \pwdata_REG[1] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[1]), .Q(pwdata[1]), .QN( ));
Q_LDP0 \pwdata_REG[2] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[2]), .Q(pwdata[2]), .QN( ));
Q_LDP0 \pwdata_REG[3] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[3]), .Q(pwdata[3]), .QN( ));
Q_LDP0 \pwdata_REG[4] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[4]), .Q(pwdata[4]), .QN( ));
Q_LDP0 \pwdata_REG[5] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[5]), .Q(pwdata[5]), .QN( ));
Q_LDP0 \pwdata_REG[6] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[6]), .Q(pwdata[6]), .QN( ));
Q_LDP0 \pwdata_REG[7] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[7]), .Q(pwdata[7]), .QN( ));
Q_LDP0 \pwdata_REG[8] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[8]), .Q(pwdata[8]), .QN( ));
Q_LDP0 \pwdata_REG[9] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[9]), .Q(pwdata[9]), .QN( ));
Q_LDP0 \pwdata_REG[10] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[10]), .Q(pwdata[10]), .QN( ));
Q_LDP0 \pwdata_REG[11] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[11]), .Q(pwdata[11]), .QN( ));
Q_LDP0 \pwdata_REG[12] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[12]), .Q(pwdata[12]), .QN( ));
Q_LDP0 \pwdata_REG[13] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[13]), .Q(pwdata[13]), .QN( ));
Q_LDP0 \pwdata_REG[14] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[14]), .Q(pwdata[14]), .QN( ));
Q_LDP0 \pwdata_REG[15] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[15]), .Q(pwdata[15]), .QN( ));
Q_LDP0 \pwdata_REG[16] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[16]), .Q(pwdata[16]), .QN( ));
Q_LDP0 \pwdata_REG[17] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[17]), .Q(pwdata[17]), .QN( ));
Q_LDP0 \pwdata_REG[18] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[18]), .Q(pwdata[18]), .QN( ));
Q_LDP0 \pwdata_REG[19] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[19]), .Q(pwdata[19]), .QN( ));
Q_LDP0 \pwdata_REG[20] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[20]), .Q(pwdata[20]), .QN( ));
Q_LDP0 \pwdata_REG[21] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[21]), .Q(pwdata[21]), .QN( ));
Q_LDP0 \pwdata_REG[22] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[22]), .Q(pwdata[22]), .QN( ));
Q_LDP0 \pwdata_REG[23] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[23]), .Q(pwdata[23]), .QN( ));
Q_LDP0 \pwdata_REG[24] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[24]), .Q(pwdata[24]), .QN( ));
Q_LDP0 \pwdata_REG[25] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[25]), .Q(pwdata[25]), .QN( ));
Q_LDP0 \pwdata_REG[26] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[26]), .Q(pwdata[26]), .QN( ));
Q_LDP0 \pwdata_REG[27] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[27]), .Q(pwdata[27]), .QN( ));
Q_LDP0 \pwdata_REG[28] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[28]), .Q(pwdata[28]), .QN( ));
Q_LDP0 \pwdata_REG[29] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[29]), .Q(pwdata[29]), .QN( ));
Q_LDP0 \pwdata_REG[30] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[30]), .Q(pwdata[30]), .QN( ));
Q_LDP0 \pwdata_REG[31] ( .G(_zzmdxOne), .D(_zzM3L22_pwdata_mdxTmp4[31]), .Q(pwdata[31]), .QN( ));
Q_MX03 U36 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[31]), .A1(_zzM3L46_mdxP0_pwdata_wr4[31]), .A2(_zzM3L61_mdxP2_pwdata_wr4[31]), .Z(_zzM3L22_pwdata_mdxTmp4[31]));
Q_MX03 U37 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[30]), .A1(_zzM3L46_mdxP0_pwdata_wr4[30]), .A2(_zzM3L61_mdxP2_pwdata_wr4[30]), .Z(_zzM3L22_pwdata_mdxTmp4[30]));
Q_MX03 U38 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[29]), .A1(_zzM3L46_mdxP0_pwdata_wr4[29]), .A2(_zzM3L61_mdxP2_pwdata_wr4[29]), .Z(_zzM3L22_pwdata_mdxTmp4[29]));
Q_MX03 U39 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[28]), .A1(_zzM3L46_mdxP0_pwdata_wr4[28]), .A2(_zzM3L61_mdxP2_pwdata_wr4[28]), .Z(_zzM3L22_pwdata_mdxTmp4[28]));
Q_MX03 U40 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[27]), .A1(_zzM3L46_mdxP0_pwdata_wr4[27]), .A2(_zzM3L61_mdxP2_pwdata_wr4[27]), .Z(_zzM3L22_pwdata_mdxTmp4[27]));
Q_MX03 U41 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[26]), .A1(_zzM3L46_mdxP0_pwdata_wr4[26]), .A2(_zzM3L61_mdxP2_pwdata_wr4[26]), .Z(_zzM3L22_pwdata_mdxTmp4[26]));
Q_MX03 U42 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[25]), .A1(_zzM3L46_mdxP0_pwdata_wr4[25]), .A2(_zzM3L61_mdxP2_pwdata_wr4[25]), .Z(_zzM3L22_pwdata_mdxTmp4[25]));
Q_MX03 U43 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[24]), .A1(_zzM3L46_mdxP0_pwdata_wr4[24]), .A2(_zzM3L61_mdxP2_pwdata_wr4[24]), .Z(_zzM3L22_pwdata_mdxTmp4[24]));
Q_MX03 U44 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[23]), .A1(_zzM3L46_mdxP0_pwdata_wr4[23]), .A2(_zzM3L61_mdxP2_pwdata_wr4[23]), .Z(_zzM3L22_pwdata_mdxTmp4[23]));
Q_MX03 U45 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[22]), .A1(_zzM3L46_mdxP0_pwdata_wr4[22]), .A2(_zzM3L61_mdxP2_pwdata_wr4[22]), .Z(_zzM3L22_pwdata_mdxTmp4[22]));
Q_MX03 U46 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[21]), .A1(_zzM3L46_mdxP0_pwdata_wr4[21]), .A2(_zzM3L61_mdxP2_pwdata_wr4[21]), .Z(_zzM3L22_pwdata_mdxTmp4[21]));
Q_MX03 U47 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[20]), .A1(_zzM3L46_mdxP0_pwdata_wr4[20]), .A2(_zzM3L61_mdxP2_pwdata_wr4[20]), .Z(_zzM3L22_pwdata_mdxTmp4[20]));
Q_MX03 U48 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[19]), .A1(_zzM3L46_mdxP0_pwdata_wr4[19]), .A2(_zzM3L61_mdxP2_pwdata_wr4[19]), .Z(_zzM3L22_pwdata_mdxTmp4[19]));
Q_MX03 U49 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[18]), .A1(_zzM3L46_mdxP0_pwdata_wr4[18]), .A2(_zzM3L61_mdxP2_pwdata_wr4[18]), .Z(_zzM3L22_pwdata_mdxTmp4[18]));
Q_MX03 U50 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[17]), .A1(_zzM3L46_mdxP0_pwdata_wr4[17]), .A2(_zzM3L61_mdxP2_pwdata_wr4[17]), .Z(_zzM3L22_pwdata_mdxTmp4[17]));
Q_MX03 U51 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[16]), .A1(_zzM3L46_mdxP0_pwdata_wr4[16]), .A2(_zzM3L61_mdxP2_pwdata_wr4[16]), .Z(_zzM3L22_pwdata_mdxTmp4[16]));
Q_MX03 U52 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[15]), .A1(_zzM3L46_mdxP0_pwdata_wr4[15]), .A2(_zzM3L61_mdxP2_pwdata_wr4[15]), .Z(_zzM3L22_pwdata_mdxTmp4[15]));
Q_MX03 U53 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[14]), .A1(_zzM3L46_mdxP0_pwdata_wr4[14]), .A2(_zzM3L61_mdxP2_pwdata_wr4[14]), .Z(_zzM3L22_pwdata_mdxTmp4[14]));
Q_MX03 U54 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[13]), .A1(_zzM3L46_mdxP0_pwdata_wr4[13]), .A2(_zzM3L61_mdxP2_pwdata_wr4[13]), .Z(_zzM3L22_pwdata_mdxTmp4[13]));
Q_MX03 U55 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[12]), .A1(_zzM3L46_mdxP0_pwdata_wr4[12]), .A2(_zzM3L61_mdxP2_pwdata_wr4[12]), .Z(_zzM3L22_pwdata_mdxTmp4[12]));
Q_MX03 U56 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[11]), .A1(_zzM3L46_mdxP0_pwdata_wr4[11]), .A2(_zzM3L61_mdxP2_pwdata_wr4[11]), .Z(_zzM3L22_pwdata_mdxTmp4[11]));
Q_MX03 U57 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[10]), .A1(_zzM3L46_mdxP0_pwdata_wr4[10]), .A2(_zzM3L61_mdxP2_pwdata_wr4[10]), .Z(_zzM3L22_pwdata_mdxTmp4[10]));
Q_MX03 U58 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[9]), .A1(_zzM3L46_mdxP0_pwdata_wr4[9]), .A2(_zzM3L61_mdxP2_pwdata_wr4[9]), .Z(_zzM3L22_pwdata_mdxTmp4[9]));
Q_MX03 U59 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[8]), .A1(_zzM3L46_mdxP0_pwdata_wr4[8]), .A2(_zzM3L61_mdxP2_pwdata_wr4[8]), .Z(_zzM3L22_pwdata_mdxTmp4[8]));
Q_MX03 U60 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[7]), .A1(_zzM3L46_mdxP0_pwdata_wr4[7]), .A2(_zzM3L61_mdxP2_pwdata_wr4[7]), .Z(_zzM3L22_pwdata_mdxTmp4[7]));
Q_MX03 U61 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[6]), .A1(_zzM3L46_mdxP0_pwdata_wr4[6]), .A2(_zzM3L61_mdxP2_pwdata_wr4[6]), .Z(_zzM3L22_pwdata_mdxTmp4[6]));
Q_MX03 U62 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[5]), .A1(_zzM3L46_mdxP0_pwdata_wr4[5]), .A2(_zzM3L61_mdxP2_pwdata_wr4[5]), .Z(_zzM3L22_pwdata_mdxTmp4[5]));
Q_MX03 U63 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[4]), .A1(_zzM3L46_mdxP0_pwdata_wr4[4]), .A2(_zzM3L61_mdxP2_pwdata_wr4[4]), .Z(_zzM3L22_pwdata_mdxTmp4[4]));
Q_MX03 U64 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[3]), .A1(_zzM3L46_mdxP0_pwdata_wr4[3]), .A2(_zzM3L61_mdxP2_pwdata_wr4[3]), .Z(_zzM3L22_pwdata_mdxTmp4[3]));
Q_MX03 U65 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[2]), .A1(_zzM3L46_mdxP0_pwdata_wr4[2]), .A2(_zzM3L61_mdxP2_pwdata_wr4[2]), .Z(_zzM3L22_pwdata_mdxTmp4[2]));
Q_MX03 U66 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[1]), .A1(_zzM3L46_mdxP0_pwdata_wr4[1]), .A2(_zzM3L61_mdxP2_pwdata_wr4[1]), .Z(_zzM3L22_pwdata_mdxTmp4[1]));
Q_MX03 U67 ( .S0(n3), .S1(_zzM3L61_mdxP2_pwdata_DwenOn4), .A0(_zzpwdata_M3L22_mdxSvLt9[0]), .A1(_zzM3L46_mdxP0_pwdata_wr4[0]), .A2(_zzM3L61_mdxP2_pwdata_wr4[0]), .Z(_zzM3L22_pwdata_mdxTmp4[0]));
Q_AN02 U68 ( .A0(_zzM3L61_mdxP2_On), .A1(_zzM3L61_mdxP2_pwdata_Dwen4), .Z(_zzM3L61_mdxP2_pwdata_DwenOn4));
Q_AN02 U69 ( .A0(_zzM3L46_mdxP0_On), .A1(_zzM3L46_mdxP0_pwdata_Dwen4), .Z(_zzM3L46_mdxP0_pwdata_DwenOn4));
Q_OR02 U70 ( .A0(_zzM3L61_mdxP2_paddr_DwenOn3), .A1(_zzM3L94_mdxP1_paddr_DwenOn3), .Z(n5));
Q_INV U71 ( .A(_zzM3L46_mdxP0_paddr_DwenOn3), .Z(n7));
Q_NR02 U72 ( .A0(_zzM3L94_mdxP1_paddr_DwenOn3), .A1(n7), .Z(n8));
Q_OR02 U73 ( .A0(_zzM3L61_mdxP2_paddr_DwenOn3), .A1(n8), .Z(n6));
Q_LDP0 \paddr_REG[0] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[0]), .Q(paddr[0]), .QN( ));
Q_LDP0 \paddr_REG[1] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[1]), .Q(paddr[1]), .QN( ));
Q_LDP0 \paddr_REG[2] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[2]), .Q(paddr[2]), .QN( ));
Q_LDP0 \paddr_REG[3] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[3]), .Q(paddr[3]), .QN( ));
Q_LDP0 \paddr_REG[4] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[4]), .Q(paddr[4]), .QN( ));
Q_LDP0 \paddr_REG[5] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[5]), .Q(paddr[5]), .QN( ));
Q_LDP0 \paddr_REG[6] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[6]), .Q(paddr[6]), .QN( ));
Q_LDP0 \paddr_REG[7] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[7]), .Q(paddr[7]), .QN( ));
Q_LDP0 \paddr_REG[8] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[8]), .Q(paddr[8]), .QN( ));
Q_LDP0 \paddr_REG[9] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[9]), .Q(paddr[9]), .QN( ));
Q_LDP0 \paddr_REG[10] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[10]), .Q(paddr[10]), .QN( ));
Q_LDP0 \paddr_REG[11] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[11]), .Q(paddr[11]), .QN( ));
Q_LDP0 \paddr_REG[12] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[12]), .Q(paddr[12]), .QN( ));
Q_LDP0 \paddr_REG[13] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[13]), .Q(paddr[13]), .QN( ));
Q_LDP0 \paddr_REG[14] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[14]), .Q(paddr[14]), .QN( ));
Q_LDP0 \paddr_REG[15] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[15]), .Q(paddr[15]), .QN( ));
Q_LDP0 \paddr_REG[16] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[16]), .Q(paddr[16]), .QN( ));
Q_LDP0 \paddr_REG[17] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[17]), .Q(paddr[17]), .QN( ));
Q_LDP0 \paddr_REG[18] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[18]), .Q(paddr[18]), .QN( ));
Q_LDP0 \paddr_REG[19] ( .G(_zzmdxOne), .D(_zzM3L21_paddr_mdxTmp3[19]), .Q(paddr[19]), .QN( ));
Q_MX04 U94 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[19]), .A1(_zzM3L46_mdxP0_paddr_wr3[19]), .A2(_zzM3L94_mdxP1_paddr_wr3[19]), .A3(_zzM3L61_mdxP2_paddr_wr3[19]), .Z(_zzM3L21_paddr_mdxTmp3[19]));
Q_MX04 U95 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[18]), .A1(_zzM3L46_mdxP0_paddr_wr3[18]), .A2(_zzM3L94_mdxP1_paddr_wr3[18]), .A3(_zzM3L61_mdxP2_paddr_wr3[18]), .Z(_zzM3L21_paddr_mdxTmp3[18]));
Q_MX04 U96 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[17]), .A1(_zzM3L46_mdxP0_paddr_wr3[17]), .A2(_zzM3L94_mdxP1_paddr_wr3[17]), .A3(_zzM3L61_mdxP2_paddr_wr3[17]), .Z(_zzM3L21_paddr_mdxTmp3[17]));
Q_MX04 U97 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[16]), .A1(_zzM3L46_mdxP0_paddr_wr3[16]), .A2(_zzM3L94_mdxP1_paddr_wr3[16]), .A3(_zzM3L61_mdxP2_paddr_wr3[16]), .Z(_zzM3L21_paddr_mdxTmp3[16]));
Q_MX04 U98 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[15]), .A1(_zzM3L46_mdxP0_paddr_wr3[15]), .A2(_zzM3L94_mdxP1_paddr_wr3[15]), .A3(_zzM3L61_mdxP2_paddr_wr3[15]), .Z(_zzM3L21_paddr_mdxTmp3[15]));
Q_MX04 U99 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[14]), .A1(_zzM3L46_mdxP0_paddr_wr3[14]), .A2(_zzM3L94_mdxP1_paddr_wr3[14]), .A3(_zzM3L61_mdxP2_paddr_wr3[14]), .Z(_zzM3L21_paddr_mdxTmp3[14]));
Q_MX04 U100 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[13]), .A1(_zzM3L46_mdxP0_paddr_wr3[13]), .A2(_zzM3L94_mdxP1_paddr_wr3[13]), .A3(_zzM3L61_mdxP2_paddr_wr3[13]), .Z(_zzM3L21_paddr_mdxTmp3[13]));
Q_MX04 U101 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[12]), .A1(_zzM3L46_mdxP0_paddr_wr3[12]), .A2(_zzM3L94_mdxP1_paddr_wr3[12]), .A3(_zzM3L61_mdxP2_paddr_wr3[12]), .Z(_zzM3L21_paddr_mdxTmp3[12]));
Q_MX04 U102 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[11]), .A1(_zzM3L46_mdxP0_paddr_wr3[11]), .A2(_zzM3L94_mdxP1_paddr_wr3[11]), .A3(_zzM3L61_mdxP2_paddr_wr3[11]), .Z(_zzM3L21_paddr_mdxTmp3[11]));
Q_MX04 U103 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[10]), .A1(_zzM3L46_mdxP0_paddr_wr3[10]), .A2(_zzM3L94_mdxP1_paddr_wr3[10]), .A3(_zzM3L61_mdxP2_paddr_wr3[10]), .Z(_zzM3L21_paddr_mdxTmp3[10]));
Q_MX04 U104 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[9]), .A1(_zzM3L46_mdxP0_paddr_wr3[9]), .A2(_zzM3L94_mdxP1_paddr_wr3[9]), .A3(_zzM3L61_mdxP2_paddr_wr3[9]), .Z(_zzM3L21_paddr_mdxTmp3[9]));
Q_MX04 U105 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[8]), .A1(_zzM3L46_mdxP0_paddr_wr3[8]), .A2(_zzM3L94_mdxP1_paddr_wr3[8]), .A3(_zzM3L61_mdxP2_paddr_wr3[8]), .Z(_zzM3L21_paddr_mdxTmp3[8]));
Q_MX04 U106 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[7]), .A1(_zzM3L46_mdxP0_paddr_wr3[7]), .A2(_zzM3L94_mdxP1_paddr_wr3[7]), .A3(_zzM3L61_mdxP2_paddr_wr3[7]), .Z(_zzM3L21_paddr_mdxTmp3[7]));
Q_MX04 U107 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[6]), .A1(_zzM3L46_mdxP0_paddr_wr3[6]), .A2(_zzM3L94_mdxP1_paddr_wr3[6]), .A3(_zzM3L61_mdxP2_paddr_wr3[6]), .Z(_zzM3L21_paddr_mdxTmp3[6]));
Q_MX04 U108 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[5]), .A1(_zzM3L46_mdxP0_paddr_wr3[5]), .A2(_zzM3L94_mdxP1_paddr_wr3[5]), .A3(_zzM3L61_mdxP2_paddr_wr3[5]), .Z(_zzM3L21_paddr_mdxTmp3[5]));
Q_MX04 U109 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[4]), .A1(_zzM3L46_mdxP0_paddr_wr3[4]), .A2(_zzM3L94_mdxP1_paddr_wr3[4]), .A3(_zzM3L61_mdxP2_paddr_wr3[4]), .Z(_zzM3L21_paddr_mdxTmp3[4]));
Q_MX04 U110 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[3]), .A1(_zzM3L46_mdxP0_paddr_wr3[3]), .A2(_zzM3L94_mdxP1_paddr_wr3[3]), .A3(_zzM3L61_mdxP2_paddr_wr3[3]), .Z(_zzM3L21_paddr_mdxTmp3[3]));
Q_MX04 U111 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[2]), .A1(_zzM3L46_mdxP0_paddr_wr3[2]), .A2(_zzM3L94_mdxP1_paddr_wr3[2]), .A3(_zzM3L61_mdxP2_paddr_wr3[2]), .Z(_zzM3L21_paddr_mdxTmp3[2]));
Q_MX04 U112 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[1]), .A1(_zzM3L46_mdxP0_paddr_wr3[1]), .A2(_zzM3L94_mdxP1_paddr_wr3[1]), .A3(_zzM3L61_mdxP2_paddr_wr3[1]), .Z(_zzM3L21_paddr_mdxTmp3[1]));
Q_MX04 U113 ( .S0(n6), .S1(n5), .A0(_zzpaddr_M3L21_mdxSvLt8[0]), .A1(_zzM3L46_mdxP0_paddr_wr3[0]), .A2(_zzM3L94_mdxP1_paddr_wr3[0]), .A3(_zzM3L61_mdxP2_paddr_wr3[0]), .Z(_zzM3L21_paddr_mdxTmp3[0]));
Q_AN02 U114 ( .A0(_zzM3L61_mdxP2_On), .A1(_zzM3L61_mdxP2_paddr_Dwen3), .Z(_zzM3L61_mdxP2_paddr_DwenOn3));
Q_AN02 U115 ( .A0(_zzM3L94_mdxP1_On), .A1(_zzM3L94_mdxP1_paddr_Dwen3), .Z(_zzM3L94_mdxP1_paddr_DwenOn3));
Q_AN02 U116 ( .A0(_zzM3L46_mdxP0_On), .A1(_zzM3L46_mdxP0_paddr_Dwen3), .Z(_zzM3L46_mdxP0_paddr_DwenOn3));
Q_OR02 U117 ( .A0(_zzM3L61_mdxP2_pwrite_DwenOn2), .A1(_zzM3L94_mdxP1_pwrite_DwenOn2), .Z(n9));
Q_INV U118 ( .A(_zzM3L46_mdxP0_pwrite_DwenOn2), .Z(n11));
Q_NR02 U119 ( .A0(_zzM3L94_mdxP1_pwrite_DwenOn2), .A1(n11), .Z(n12));
Q_OR02 U120 ( .A0(_zzM3L61_mdxP2_pwrite_DwenOn2), .A1(n12), .Z(n10));
Q_LDP0 pwrite_REG  ( .G(_zzmdxOne), .D(_zzM3L23_pwrite_mdxTmp2), .Q(pwrite), .QN( ));
Q_MX04 U122 ( .S0(n10), .S1(n9), .A0(_zzpwrite_M3L23_mdxSvLt7), .A1(_zzM3L46_mdxP0_pwrite_wr2), .A2(_zzM3L94_mdxP1_pwrite_wr2), .A3(_zzM3L61_mdxP2_pwrite_wr2), .Z(_zzM3L23_pwrite_mdxTmp2));
Q_AN02 U123 ( .A0(_zzM3L61_mdxP2_On), .A1(_zzM3L61_mdxP2_pwrite_Dwen2), .Z(_zzM3L61_mdxP2_pwrite_DwenOn2));
Q_AN02 U124 ( .A0(_zzM3L94_mdxP1_On), .A1(_zzM3L94_mdxP1_pwrite_Dwen2), .Z(_zzM3L94_mdxP1_pwrite_DwenOn2));
Q_AN02 U125 ( .A0(_zzM3L46_mdxP0_On), .A1(_zzM3L46_mdxP0_pwrite_Dwen2), .Z(_zzM3L46_mdxP0_pwrite_DwenOn2));
Q_OR02 U126 ( .A0(_zzM3L61_mdxP2_penable_DwenOn1), .A1(_zzM3L94_mdxP1_penable_DwenOn1), .Z(n13));
Q_INV U127 ( .A(_zzM3L46_mdxP0_penable_DwenOn1), .Z(n15));
Q_NR02 U128 ( .A0(_zzM3L94_mdxP1_penable_DwenOn1), .A1(n15), .Z(n16));
Q_OR02 U129 ( .A0(_zzM3L61_mdxP2_penable_DwenOn1), .A1(n16), .Z(n14));
Q_LDP0 penable_REG  ( .G(_zzmdxOne), .D(_zzM3L20_penable_mdxTmp1), .Q(penable), .QN( ));
Q_MX04 U131 ( .S0(n14), .S1(n13), .A0(_zzpenable_M3L20_mdxSvLt6), .A1(_zzM3L46_mdxP0_penable_wr1), .A2(_zzM3L94_mdxP1_penable_wr1), .A3(_zzM3L61_mdxP2_penable_wr1), .Z(_zzM3L20_penable_mdxTmp1));
Q_AN02 U132 ( .A0(_zzM3L61_mdxP2_On), .A1(_zzM3L61_mdxP2_penable_Dwen1), .Z(_zzM3L61_mdxP2_penable_DwenOn1));
Q_AN02 U133 ( .A0(_zzM3L94_mdxP1_On), .A1(_zzM3L94_mdxP1_penable_Dwen1), .Z(_zzM3L94_mdxP1_penable_DwenOn1));
Q_AN02 U134 ( .A0(_zzM3L46_mdxP0_On), .A1(_zzM3L46_mdxP0_penable_Dwen1), .Z(_zzM3L46_mdxP0_penable_DwenOn1));
Q_OR02 U135 ( .A0(_zzM3L61_mdxP2_psel_DwenOn0), .A1(_zzM3L94_mdxP1_psel_DwenOn0), .Z(n17));
Q_INV U136 ( .A(_zzM3L46_mdxP0_psel_DwenOn0), .Z(n19));
Q_NR02 U137 ( .A0(_zzM3L94_mdxP1_psel_DwenOn0), .A1(n19), .Z(n20));
Q_OR02 U138 ( .A0(_zzM3L61_mdxP2_psel_DwenOn0), .A1(n20), .Z(n18));
Q_LDP0 psel_REG  ( .G(_zzmdxOne), .D(_zzM3L19_psel_mdxTmp0), .Q(psel), .QN( ));
Q_MX04 U140 ( .S0(n18), .S1(n17), .A0(_zzpsel_M3L19_mdxSvLt5), .A1(_zzM3L46_mdxP0_psel_wr0), .A2(_zzM3L94_mdxP1_psel_wr0), .A3(_zzM3L61_mdxP2_psel_wr0), .Z(_zzM3L19_psel_mdxTmp0));
Q_AN02 U141 ( .A0(_zzM3L61_mdxP2_On), .A1(_zzM3L61_mdxP2_psel_Dwen0), .Z(_zzM3L61_mdxP2_psel_DwenOn0));
Q_AN02 U142 ( .A0(_zzM3L94_mdxP1_On), .A1(_zzM3L94_mdxP1_psel_Dwen0), .Z(_zzM3L94_mdxP1_psel_DwenOn0));
Q_AN02 U143 ( .A0(_zzM3L46_mdxP0_On), .A1(_zzM3L46_mdxP0_psel_Dwen0), .Z(_zzM3L46_mdxP0_psel_DwenOn0));
Q_AN02 U144 ( .A0(n22), .A1(n81), .Z(n21));
Q_AD01HF U145 ( .A0(_zzM3_bcBehEval[29]), .B0(n25), .S(n24), .CO(n23));
Q_AD01HF U146 ( .A0(_zzM3_bcBehEval[28]), .B0(n27), .S(n26), .CO(n25));
Q_AD01HF U147 ( .A0(_zzM3_bcBehEval[27]), .B0(n29), .S(n28), .CO(n27));
Q_AD01HF U148 ( .A0(_zzM3_bcBehEval[26]), .B0(n31), .S(n30), .CO(n29));
Q_AD01HF U149 ( .A0(_zzM3_bcBehEval[25]), .B0(n33), .S(n32), .CO(n31));
Q_AD01HF U150 ( .A0(_zzM3_bcBehEval[24]), .B0(n35), .S(n34), .CO(n33));
Q_AD01HF U151 ( .A0(_zzM3_bcBehEval[23]), .B0(n37), .S(n36), .CO(n35));
Q_AD01HF U152 ( .A0(_zzM3_bcBehEval[22]), .B0(n39), .S(n38), .CO(n37));
Q_AD01HF U153 ( .A0(_zzM3_bcBehEval[21]), .B0(n41), .S(n40), .CO(n39));
Q_AD01HF U154 ( .A0(_zzM3_bcBehEval[20]), .B0(n43), .S(n42), .CO(n41));
Q_AD01HF U155 ( .A0(_zzM3_bcBehEval[19]), .B0(n45), .S(n44), .CO(n43));
Q_AD01HF U156 ( .A0(_zzM3_bcBehEval[18]), .B0(n47), .S(n46), .CO(n45));
Q_AD01HF U157 ( .A0(_zzM3_bcBehEval[17]), .B0(n49), .S(n48), .CO(n47));
Q_AD01HF U158 ( .A0(_zzM3_bcBehEval[16]), .B0(n51), .S(n50), .CO(n49));
Q_AD01HF U159 ( .A0(_zzM3_bcBehEval[15]), .B0(n53), .S(n52), .CO(n51));
Q_AD01HF U160 ( .A0(_zzM3_bcBehEval[14]), .B0(n55), .S(n54), .CO(n53));
Q_AD01HF U161 ( .A0(_zzM3_bcBehEval[13]), .B0(n57), .S(n56), .CO(n55));
Q_AD01HF U162 ( .A0(_zzM3_bcBehEval[12]), .B0(n59), .S(n58), .CO(n57));
Q_AD01HF U163 ( .A0(_zzM3_bcBehEval[11]), .B0(n61), .S(n60), .CO(n59));
Q_AD01HF U164 ( .A0(_zzM3_bcBehEval[10]), .B0(n63), .S(n62), .CO(n61));
Q_AD01HF U165 ( .A0(_zzM3_bcBehEval[9]), .B0(n65), .S(n64), .CO(n63));
Q_AD01HF U166 ( .A0(_zzM3_bcBehEval[8]), .B0(n67), .S(n66), .CO(n65));
Q_AD01HF U167 ( .A0(_zzM3_bcBehEval[7]), .B0(n69), .S(n68), .CO(n67));
Q_AD01HF U168 ( .A0(_zzM3_bcBehEval[6]), .B0(n71), .S(n70), .CO(n69));
Q_AD01HF U169 ( .A0(_zzM3_bcBehEval[5]), .B0(n73), .S(n72), .CO(n71));
Q_AD01HF U170 ( .A0(_zzM3_bcBehEval[4]), .B0(n75), .S(n74), .CO(n73));
Q_AD01HF U171 ( .A0(_zzM3_bcBehEval[3]), .B0(n77), .S(n76), .CO(n75));
Q_AD01HF U172 ( .A0(_zzM3_bcBehEval[2]), .B0(n79), .S(n78), .CO(n77));
Q_AD01HF U173 ( .A0(_zzM3_bcBehEval[1]), .B0(_zzM3_bcBehEval[0]), .S(n80), .CO(n79));
Q_OR02 U174 ( .A0(_zyM3L94_pbcWait4), .A1(_zyM3L61_pbcWait9), .Z(n22));
Q_ND03 U175 ( .A0(n84), .A1(n83), .A2(n82), .Z(n81));
Q_AN03 U176 ( .A0(n87), .A1(n86), .A2(n85), .Z(n82));
Q_AN03 U177 ( .A0(n90), .A1(n89), .A2(n88), .Z(n83));
Q_AN03 U178 ( .A0(n93), .A1(n92), .A2(n91), .Z(n84));
Q_AN03 U179 ( .A0(_zzM3_bcBehEval[0]), .A1(n95), .A2(n94), .Z(n85));
Q_AN03 U180 ( .A0(_zzM3_bcBehEval[3]), .A1(_zzM3_bcBehEval[2]), .A2(_zzM3_bcBehEval[1]), .Z(n86));
Q_AN03 U181 ( .A0(_zzM3_bcBehEval[6]), .A1(_zzM3_bcBehEval[5]), .A2(_zzM3_bcBehEval[4]), .Z(n87));
Q_AN03 U182 ( .A0(_zzM3_bcBehEval[9]), .A1(_zzM3_bcBehEval[8]), .A2(_zzM3_bcBehEval[7]), .Z(n88));
Q_AN03 U183 ( .A0(_zzM3_bcBehEval[12]), .A1(_zzM3_bcBehEval[11]), .A2(_zzM3_bcBehEval[10]), .Z(n89));
Q_AN03 U184 ( .A0(_zzM3_bcBehEval[15]), .A1(_zzM3_bcBehEval[14]), .A2(_zzM3_bcBehEval[13]), .Z(n90));
Q_AN03 U185 ( .A0(_zzM3_bcBehEval[18]), .A1(_zzM3_bcBehEval[17]), .A2(_zzM3_bcBehEval[16]), .Z(n91));
Q_AN03 U186 ( .A0(_zzM3_bcBehEval[21]), .A1(_zzM3_bcBehEval[20]), .A2(_zzM3_bcBehEval[19]), .Z(n92));
Q_AN03 U187 ( .A0(_zzM3_bcBehEval[24]), .A1(_zzM3_bcBehEval[23]), .A2(_zzM3_bcBehEval[22]), .Z(n93));
Q_AN03 U188 ( .A0(_zzM3_bcBehEval[27]), .A1(_zzM3_bcBehEval[26]), .A2(_zzM3_bcBehEval[25]), .Z(n94));
Q_AN03 U189 ( .A0(_zzM3_bcBehEval[30]), .A1(_zzM3_bcBehEval[29]), .A2(_zzM3_bcBehEval[28]), .Z(n95));
Q_LDP0 _zyresponse_L64_tfiV5_M3_pbcG5_REG  ( .G(_zzbcOne), .D(_zzM3L64__zyresponse_L64_tfiV5_M3_pbcG5_nbaTmp6), .Q(_zyresponse_L64_tfiV5_M3_pbcG5), .QN( ));
Q_MX02 U191 ( .S(_zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_DwenOn1), .A0(_zz_zyresponse_L64_tfiV5_M3_pbcG5_M3_bcSvLt10), .A1(_zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_wr1), .Z(_zzM3L64__zyresponse_L64_tfiV5_M3_pbcG5_nbaTmp6));
Q_AN02 U192 ( .A0(_zzM3L61_bcP2_DOn), .A1(_zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_Dwen1), .Z(_zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_DwenOn1));
Q_LDP0 _zyresponse_L97_tfiV2_M3_pbcG2_REG  ( .G(_zzbcOne), .D(_zzM3L97__zyresponse_L97_tfiV2_M3_pbcG2_nbaTmp5), .Q(_zyresponse_L97_tfiV2_M3_pbcG2), .QN( ));
Q_MX02 U194 ( .S(_zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_DwenOn2), .A0(_zz_zyresponse_L97_tfiV2_M3_pbcG2_M3_bcSvLt9), .A1(_zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_wr2), .Z(_zzM3L97__zyresponse_L97_tfiV2_M3_pbcG2_nbaTmp5));
Q_AN02 U195 ( .A0(_zzM3L94_bcP1_DOn), .A1(_zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_Dwen2), .Z(_zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_DwenOn2));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[0] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[0]), .Q(_zydata_L96_tfiV1_M3_pbcG1[0]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[1] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[1]), .Q(_zydata_L96_tfiV1_M3_pbcG1[1]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[2] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[2]), .Q(_zydata_L96_tfiV1_M3_pbcG1[2]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[3] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[3]), .Q(_zydata_L96_tfiV1_M3_pbcG1[3]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[4] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[4]), .Q(_zydata_L96_tfiV1_M3_pbcG1[4]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[5] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[5]), .Q(_zydata_L96_tfiV1_M3_pbcG1[5]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[6] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[6]), .Q(_zydata_L96_tfiV1_M3_pbcG1[6]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[7] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[7]), .Q(_zydata_L96_tfiV1_M3_pbcG1[7]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[8] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[8]), .Q(_zydata_L96_tfiV1_M3_pbcG1[8]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[9] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[9]), .Q(_zydata_L96_tfiV1_M3_pbcG1[9]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[10] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[10]), .Q(_zydata_L96_tfiV1_M3_pbcG1[10]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[11] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[11]), .Q(_zydata_L96_tfiV1_M3_pbcG1[11]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[12] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[12]), .Q(_zydata_L96_tfiV1_M3_pbcG1[12]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[13] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[13]), .Q(_zydata_L96_tfiV1_M3_pbcG1[13]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[14] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[14]), .Q(_zydata_L96_tfiV1_M3_pbcG1[14]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[15] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[15]), .Q(_zydata_L96_tfiV1_M3_pbcG1[15]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[16] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[16]), .Q(_zydata_L96_tfiV1_M3_pbcG1[16]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[17] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[17]), .Q(_zydata_L96_tfiV1_M3_pbcG1[17]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[18] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[18]), .Q(_zydata_L96_tfiV1_M3_pbcG1[18]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[19] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[19]), .Q(_zydata_L96_tfiV1_M3_pbcG1[19]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[20] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[20]), .Q(_zydata_L96_tfiV1_M3_pbcG1[20]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[21] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[21]), .Q(_zydata_L96_tfiV1_M3_pbcG1[21]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[22] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[22]), .Q(_zydata_L96_tfiV1_M3_pbcG1[22]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[23] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[23]), .Q(_zydata_L96_tfiV1_M3_pbcG1[23]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[24] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[24]), .Q(_zydata_L96_tfiV1_M3_pbcG1[24]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[25] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[25]), .Q(_zydata_L96_tfiV1_M3_pbcG1[25]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[26] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[26]), .Q(_zydata_L96_tfiV1_M3_pbcG1[26]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[27] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[27]), .Q(_zydata_L96_tfiV1_M3_pbcG1[27]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[28] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[28]), .Q(_zydata_L96_tfiV1_M3_pbcG1[28]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[29] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[29]), .Q(_zydata_L96_tfiV1_M3_pbcG1[29]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[30] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[30]), .Q(_zydata_L96_tfiV1_M3_pbcG1[30]), .QN( ));
Q_LDP0 \_zydata_L96_tfiV1_M3_pbcG1_REG[31] ( .G(_zzbcOne), .D(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[31]), .Q(_zydata_L96_tfiV1_M3_pbcG1[31]), .QN( ));
Q_MX02 U228 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[31]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[31]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[31]));
Q_MX02 U229 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[30]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[30]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[30]));
Q_MX02 U230 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[29]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[29]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[29]));
Q_MX02 U231 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[28]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[28]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[28]));
Q_MX02 U232 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[27]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[27]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[27]));
Q_MX02 U233 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[26]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[26]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[26]));
Q_MX02 U234 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[25]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[25]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[25]));
Q_MX02 U235 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[24]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[24]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[24]));
Q_MX02 U236 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[23]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[23]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[23]));
Q_MX02 U237 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[22]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[22]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[22]));
Q_MX02 U238 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[21]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[21]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[21]));
Q_MX02 U239 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[20]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[20]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[20]));
Q_MX02 U240 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[19]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[19]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[19]));
Q_MX02 U241 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[18]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[18]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[18]));
Q_MX02 U242 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[17]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[17]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[17]));
Q_MX02 U243 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[16]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[16]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[16]));
Q_MX02 U244 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[15]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[15]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[15]));
Q_MX02 U245 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[14]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[14]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[14]));
Q_MX02 U246 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[13]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[13]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[13]));
Q_MX02 U247 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[12]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[12]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[12]));
Q_MX02 U248 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[11]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[11]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[11]));
Q_MX02 U249 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[10]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[10]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[10]));
Q_MX02 U250 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[9]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[9]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[9]));
Q_MX02 U251 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[8]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[8]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[8]));
Q_MX02 U252 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[7]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[7]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[7]));
Q_MX02 U253 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[6]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[6]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[6]));
Q_MX02 U254 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[5]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[5]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[5]));
Q_MX02 U255 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[4]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[4]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[4]));
Q_MX02 U256 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[3]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[3]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[3]));
Q_MX02 U257 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[2]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[2]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[2]));
Q_MX02 U258 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[1]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[1]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[1]));
Q_MX02 U259 ( .S(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1), .A0(_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[0]), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[0]), .Z(_zzM3L96__zydata_L96_tfiV1_M3_pbcG1_nbaTmp4[0]));
Q_AN02 U260 ( .A0(_zzM3L94_bcP1_DOn), .A1(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_Dwen1), .Z(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_DwenOn1));
Q_OR02 U261 ( .A0(_zzM3L61_bcP2_bus_timer_DwenOn0), .A1(_zzM3L94_bcP1_bus_timer_DwenOn0), .Z(n96));
Q_INV U262 ( .A(_zzM3L46_bcP0_bus_timer_DwenOn0), .Z(n98));
Q_NR02 U263 ( .A0(_zzM3L94_bcP1_bus_timer_DwenOn0), .A1(n98), .Z(n99));
Q_OR02 U264 ( .A0(_zzM3L61_bcP2_bus_timer_DwenOn0), .A1(n99), .Z(n97));
Q_LDP0 \bus_timer_REG[0] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[0]), .Q(bus_timer[0]), .QN(n297));
Q_LDP0 \bus_timer_REG[1] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[1]), .Q(bus_timer[1]), .QN( ));
Q_LDP0 \bus_timer_REG[2] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[2]), .Q(bus_timer[2]), .QN(n305));
Q_LDP0 \bus_timer_REG[3] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[3]), .Q(bus_timer[3]), .QN( ));
Q_LDP0 \bus_timer_REG[4] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[4]), .Q(bus_timer[4]), .QN(n309));
Q_LDP0 \bus_timer_REG[5] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[5]), .Q(bus_timer[5]), .QN(n310));
Q_LDP0 \bus_timer_REG[6] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[6]), .Q(bus_timer[6]), .QN(n311));
Q_LDP0 \bus_timer_REG[7] ( .G(_zzbcOne), .D(_zzM3L29_bus_timer_nbaTmp3[7]), .Q(bus_timer[7]), .QN(n312));
Q_MX04 U273 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[7]), .A1(_zzM3L46_bcP0_bus_timer_wr0[7]), .A2(_zzM3L94_bcP1_bus_timer_wr0[7]), .A3(_zzM3L61_bcP2_bus_timer_wr0[7]), .Z(_zzM3L29_bus_timer_nbaTmp3[7]));
Q_MX04 U274 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[6]), .A1(_zzM3L46_bcP0_bus_timer_wr0[6]), .A2(_zzM3L94_bcP1_bus_timer_wr0[6]), .A3(_zzM3L61_bcP2_bus_timer_wr0[6]), .Z(_zzM3L29_bus_timer_nbaTmp3[6]));
Q_MX04 U275 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[5]), .A1(_zzM3L46_bcP0_bus_timer_wr0[5]), .A2(_zzM3L94_bcP1_bus_timer_wr0[5]), .A3(_zzM3L61_bcP2_bus_timer_wr0[5]), .Z(_zzM3L29_bus_timer_nbaTmp3[5]));
Q_MX04 U276 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[4]), .A1(_zzM3L46_bcP0_bus_timer_wr0[4]), .A2(_zzM3L94_bcP1_bus_timer_wr0[4]), .A3(_zzM3L61_bcP2_bus_timer_wr0[4]), .Z(_zzM3L29_bus_timer_nbaTmp3[4]));
Q_MX04 U277 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[3]), .A1(_zzM3L46_bcP0_bus_timer_wr0[3]), .A2(_zzM3L94_bcP1_bus_timer_wr0[3]), .A3(_zzM3L61_bcP2_bus_timer_wr0[3]), .Z(_zzM3L29_bus_timer_nbaTmp3[3]));
Q_MX04 U278 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[2]), .A1(_zzM3L46_bcP0_bus_timer_wr0[2]), .A2(_zzM3L94_bcP1_bus_timer_wr0[2]), .A3(_zzM3L61_bcP2_bus_timer_wr0[2]), .Z(_zzM3L29_bus_timer_nbaTmp3[2]));
Q_MX04 U279 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[1]), .A1(_zzM3L46_bcP0_bus_timer_wr0[1]), .A2(_zzM3L94_bcP1_bus_timer_wr0[1]), .A3(_zzM3L61_bcP2_bus_timer_wr0[1]), .Z(_zzM3L29_bus_timer_nbaTmp3[1]));
Q_MX04 U280 ( .S0(n97), .S1(n96), .A0(_zzbus_timer_M3L29_bcSvLt7[0]), .A1(_zzM3L46_bcP0_bus_timer_wr0[0]), .A2(_zzM3L94_bcP1_bus_timer_wr0[0]), .A3(_zzM3L61_bcP2_bus_timer_wr0[0]), .Z(_zzM3L29_bus_timer_nbaTmp3[0]));
Q_AN02 U281 ( .A0(_zzM3L61_bcP2_DOn), .A1(_zzM3L61_bcP2_bus_timer_Dwen0), .Z(_zzM3L61_bcP2_bus_timer_DwenOn0));
Q_AN02 U282 ( .A0(_zzM3L94_bcP1_DOn), .A1(_zzM3L94_bcP1_bus_timer_Dwen0), .Z(_zzM3L94_bcP1_bus_timer_DwenOn0));
Q_AN02 U283 ( .A0(_zzM3L46_bcP0_DOn), .A1(_zzM3L46_bcP0_bus_timer_Dwen0), .Z(_zzM3L46_bcP0_bus_timer_DwenOn0));
Q_AN02 U284 ( .A0(n133), .A1(_zyM3L61_pbcFsm2_s[0]), .Z(n130));
Q_AN02 U285 ( .A0(_zyM3L61_pbcFsm2_s[1]), .A1(n110), .Z(n131));
Q_OR02 U286 ( .A0(n130), .A1(n131), .Z(n136));
Q_AN02 U287 ( .A0(n103), .A1(n136), .Z(n115));
Q_OR02 U288 ( .A0(_zyM3L61_pbcFsm2_s[1]), .A1(_zyM3L61_pbcFsm2_s[0]), .Z(n109));
Q_INV U289 ( .A(_zzpready_M3L25_bcSv0), .Z(n122));
Q_AN02 U290 ( .A0(n122), .A1(n100), .Z(n138));
Q_AO21 U291 ( .A0(n109), .A1(n138), .B0(n135), .Z(n137));
Q_AN02 U292 ( .A0(_zyM3L61_pbcFsm2_s[1]), .A1(_zyM3L61_pbcFsm2_s[0]), .Z(n135));
Q_OR02 U293 ( .A0(n137), .A1(_zyM3L61_pbcFsm2_s[2]), .Z(n123));
Q_INV U294 ( .A(n123), .Z(n120));
Q_OA21 U295 ( .A0(n138), .A1(_zyM3L61_pbcFsm2_s[0]), .B0(_zyM3L61_pbcFsm2_s[1]), .Z(n124));
Q_OR02 U296 ( .A0(n124), .A1(_zyM3L61_pbcFsm2_s[2]), .Z(n125));
Q_INV U297 ( .A(n125), .Z(n118));
Q_INV U298 ( .A(n109), .Z(n119));
Q_OR02 U299 ( .A0(n119), .A1(n138), .Z(n126));
Q_OR03 U300 ( .A0(n135), .A1(_zyM3L61_pbcFsm2_s[2]), .A2(n126), .Z(n128));
Q_AN02 U301 ( .A0(n229), .A1(n128), .Z(n127));
Q_INV U302 ( .A(n128), .Z(n116));
Q_OR02 U303 ( .A0(n101), .A1(n115), .Z(n102));
Q_INV U304 ( .A(n135), .Z(n111));
Q_AO21 U305 ( .A0(n111), .A1(n138), .B0(n119), .Z(n113));
Q_OR02 U306 ( .A0(n113), .A1(_zyM3L61_pbcFsm2_s[2]), .Z(n129));
Q_AO21 U307 ( .A0(n130), .A1(n138), .B0(n131), .Z(n132));
Q_AN02 U308 ( .A0(n103), .A1(n132), .Z(n104));
Q_AN02 U309 ( .A0(n103), .A1(n133), .Z(n105));
Q_INV U310 ( .A(n136), .Z(n134));
Q_AN02 U311 ( .A0(n103), .A1(n134), .Z(n106));
Q_AN02 U312 ( .A0(n103), .A1(n135), .Z(n107));
Q_AN02 U313 ( .A0(n103), .A1(n119), .Z(n108));
Q_AN02 U314 ( .A0(n138), .A1(n136), .Z(n114));
Q_INV U315 ( .A(n137), .Z(n112));
Q_AN02 U316 ( .A0(_zyM3L61_pbcFsm2_s[0]), .A1(n138), .Z(n117));
Q_INV U317 ( .A(n114), .Z(n121));
Q_FDP0 _zzM3L61_mdxP2_pwdata_Dwen4_REG  ( .CK(_zyM3L61_pbcMevClk9), .D(n120), .Q(_zzM3L61_mdxP2_pwdata_Dwen4), .QN( ));
Q_FDP0 _zzM3L61_mdxP2_paddr_Dwen3_REG  ( .CK(_zyM3L61_pbcMevClk9), .D(n120), .Q(_zzM3L61_mdxP2_paddr_Dwen3), .QN( ));
Q_FDP0 _zzM3L61_mdxP2_pwrite_Dwen2_REG  ( .CK(_zyM3L61_pbcMevClk9), .D(n120), .Q(_zzM3L61_mdxP2_pwrite_Dwen2), .QN( ));
Q_FDP0 _zzM3L61_mdxP2_penable_Dwen1_REG  ( .CK(_zyM3L61_pbcMevClk9), .D(n118), .Q(_zzM3L61_mdxP2_penable_Dwen1), .QN( ));
Q_FDP0 _zzM3L61_mdxP2_psel_Dwen0_REG  ( .CK(_zyM3L61_pbcMevClk9), .D(n120), .Q(_zzM3L61_mdxP2_psel_Dwen0), .QN( ));
Q_FDP0 \_zyM3L61_pbcFsm2_s_REG[2] ( .CK(_zyM3L61_pbcMevClk9), .D(_zyM3L61_pbcFsm2_s[2]), .Q(_zyM3L61_pbcFsm2_s[2]), .QN(n103));
Q_XNR2 U324 ( .A0(n113), .A1(n137), .Z(n139));
Q_AN02 U325 ( .A0(n114), .A1(n200), .Z(n140));
Q_AN02 U326 ( .A0(n114), .A1(n202), .Z(n141));
Q_AN02 U327 ( .A0(n114), .A1(n204), .Z(n142));
Q_AN02 U328 ( .A0(n114), .A1(n206), .Z(n143));
Q_AN02 U329 ( .A0(n114), .A1(n208), .Z(n144));
Q_AN02 U330 ( .A0(n114), .A1(n210), .Z(n145));
Q_AN02 U331 ( .A0(n114), .A1(n212), .Z(n146));
Q_AN02 U332 ( .A0(n114), .A1(n213), .Z(n147));
Q_AN02 U333 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[19]), .Z(n148));
Q_AN02 U334 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[18]), .Z(n149));
Q_AN02 U335 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[17]), .Z(n150));
Q_AN02 U336 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[16]), .Z(n151));
Q_AN02 U337 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[15]), .Z(n152));
Q_AN02 U338 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[14]), .Z(n153));
Q_AN02 U339 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[13]), .Z(n154));
Q_AN02 U340 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[12]), .Z(n155));
Q_AN02 U341 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[11]), .Z(n156));
Q_AN02 U342 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[10]), .Z(n157));
Q_AN02 U343 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[9]), .Z(n158));
Q_AN02 U344 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[8]), .Z(n159));
Q_AN02 U345 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[7]), .Z(n160));
Q_AN02 U346 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[6]), .Z(n161));
Q_AN02 U347 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[5]), .Z(n162));
Q_AN02 U348 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[4]), .Z(n163));
Q_AN02 U349 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[3]), .Z(n164));
Q_AN02 U350 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[2]), .Z(n165));
Q_AN02 U351 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[1]), .Z(n166));
Q_AN02 U352 ( .A0(n119), .A1(_zyL61_iscX2c0_i0[0]), .Z(n167));
Q_AN02 U353 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[31]), .Z(n168));
Q_AN02 U354 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[30]), .Z(n169));
Q_AN02 U355 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[29]), .Z(n170));
Q_AN02 U356 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[28]), .Z(n171));
Q_AN02 U357 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[27]), .Z(n172));
Q_AN02 U358 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[26]), .Z(n173));
Q_AN02 U359 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[25]), .Z(n174));
Q_AN02 U360 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[24]), .Z(n175));
Q_AN02 U361 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[23]), .Z(n176));
Q_AN02 U362 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[22]), .Z(n177));
Q_AN02 U363 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[21]), .Z(n178));
Q_AN02 U364 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[20]), .Z(n179));
Q_AN02 U365 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[19]), .Z(n180));
Q_AN02 U366 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[18]), .Z(n181));
Q_AN02 U367 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[17]), .Z(n182));
Q_AN02 U368 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[16]), .Z(n183));
Q_AN02 U369 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[15]), .Z(n184));
Q_AN02 U370 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[14]), .Z(n185));
Q_AN02 U371 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[13]), .Z(n186));
Q_AN02 U372 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[12]), .Z(n187));
Q_AN02 U373 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[11]), .Z(n188));
Q_AN02 U374 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[10]), .Z(n189));
Q_AN02 U375 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[9]), .Z(n190));
Q_AN02 U376 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[8]), .Z(n191));
Q_AN02 U377 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[7]), .Z(n192));
Q_AN02 U378 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[6]), .Z(n193));
Q_AN02 U379 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[5]), .Z(n194));
Q_AN02 U380 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[4]), .Z(n195));
Q_AN02 U381 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[3]), .Z(n196));
Q_AN02 U382 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[2]), .Z(n197));
Q_AN02 U383 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[1]), .Z(n198));
Q_AN02 U384 ( .A0(n119), .A1(_zyL61_iscX2c0_i1[0]), .Z(n199));
Q_XOR2 U385 ( .A0(bus_timer[7]), .A1(n201), .Z(n200));
Q_AD01HF U386 ( .A0(bus_timer[6]), .B0(n203), .S(n202), .CO(n201));
Q_AD01HF U387 ( .A0(bus_timer[5]), .B0(n205), .S(n204), .CO(n203));
Q_AD01HF U388 ( .A0(bus_timer[4]), .B0(n207), .S(n206), .CO(n205));
Q_AD01HF U389 ( .A0(bus_timer[3]), .B0(n209), .S(n208), .CO(n207));
Q_AD01HF U390 ( .A0(bus_timer[2]), .B0(n211), .S(n210), .CO(n209));
Q_AD01HF U391 ( .A0(bus_timer[1]), .B0(bus_timer[0]), .S(n212), .CO(n211));
Q_INV U392 ( .A(bus_timer[0]), .Z(n213));
Q_OR02 U393 ( .A0(_zzpslverr_M3L26_bcSv2), .A1(n215), .Z(n214));
Q_NR02 U394 ( .A0(n217), .A1(n216), .Z(n215));
Q_OR03 U395 ( .A0(bus_timer[1]), .A1(bus_timer[0]), .A2(n218), .Z(n216));
Q_OR03 U396 ( .A0(bus_timer[4]), .A1(bus_timer[3]), .A2(n221), .Z(n217));
Q_OR03 U397 ( .A0(bus_timer[7]), .A1(n219), .A2(n220), .Z(n218));
Q_INV U398 ( .A(bus_timer[6]), .Z(n219));
Q_INV U399 ( .A(bus_timer[5]), .Z(n220));
Q_INV U400 ( .A(bus_timer[2]), .Z(n221));
Q_AO21 U401 ( .A0(n223), .A1(n222), .B0(n224), .Z(n100));
Q_NR02 U402 ( .A0(bus_timer[3]), .A1(bus_timer[2]), .Z(n222));
Q_AN02 U403 ( .A0(n228), .A1(n225), .Z(n223));
Q_OA21 U404 ( .A0(n227), .A1(n226), .B0(n228), .Z(n224));
Q_INV U405 ( .A(bus_timer[4]), .Z(n225));
Q_INV U406 ( .A(bus_timer[5]), .Z(n226));
Q_INV U407 ( .A(bus_timer[6]), .Z(n227));
Q_INV U408 ( .A(bus_timer[7]), .Z(n228));
Q_INV U409 ( .A(n229), .Z(n101));
Q_XNR2 U410 ( .A0(_zzM3L61_bcP2_EnD), .A1(_zzM3L61_bcP2_EnDNxt), .Z(n229));
Q_AN02 U411 ( .A0(n262), .A1(_zyM3L94_pbcFsm0_s[0]), .Z(n259));
Q_AN02 U412 ( .A0(_zyM3L94_pbcFsm0_s[1]), .A1(n240), .Z(n260));
Q_OR02 U413 ( .A0(n259), .A1(n260), .Z(n265));
Q_AN02 U414 ( .A0(n233), .A1(n265), .Z(n245));
Q_OR02 U415 ( .A0(_zyM3L94_pbcFsm0_s[1]), .A1(_zyM3L94_pbcFsm0_s[0]), .Z(n239));
Q_AN02 U416 ( .A0(n122), .A1(n230), .Z(n267));
Q_AO21 U417 ( .A0(n239), .A1(n267), .B0(n264), .Z(n266));
Q_AN02 U418 ( .A0(_zyM3L94_pbcFsm0_s[1]), .A1(_zyM3L94_pbcFsm0_s[0]), .Z(n264));
Q_OR02 U419 ( .A0(n266), .A1(_zyM3L94_pbcFsm0_s[2]), .Z(n252));
Q_INV U420 ( .A(n252), .Z(n250));
Q_OA21 U421 ( .A0(n267), .A1(_zyM3L94_pbcFsm0_s[0]), .B0(_zyM3L94_pbcFsm0_s[1]), .Z(n253));
Q_OR02 U422 ( .A0(n253), .A1(_zyM3L94_pbcFsm0_s[2]), .Z(n254));
Q_INV U423 ( .A(n254), .Z(n248));
Q_INV U424 ( .A(n239), .Z(n249));
Q_OR02 U425 ( .A0(n249), .A1(n267), .Z(n255));
Q_OR03 U426 ( .A0(n264), .A1(_zyM3L94_pbcFsm0_s[2]), .A2(n255), .Z(n257));
Q_AN02 U427 ( .A0(n313), .A1(n257), .Z(n256));
Q_INV U428 ( .A(n257), .Z(n246));
Q_OR02 U429 ( .A0(n231), .A1(n245), .Z(n232));
Q_INV U430 ( .A(n264), .Z(n241));
Q_AO21 U431 ( .A0(n241), .A1(n267), .B0(n249), .Z(n243));
Q_OR02 U432 ( .A0(n243), .A1(_zyM3L94_pbcFsm0_s[2]), .Z(n258));
Q_AO21 U433 ( .A0(n259), .A1(n267), .B0(n260), .Z(n261));
Q_AN02 U434 ( .A0(n233), .A1(n261), .Z(n234));
Q_AN02 U435 ( .A0(n233), .A1(n262), .Z(n235));
Q_INV U436 ( .A(n265), .Z(n263));
Q_AN02 U437 ( .A0(n233), .A1(n263), .Z(n236));
Q_AN02 U438 ( .A0(n233), .A1(n264), .Z(n237));
Q_AN02 U439 ( .A0(n233), .A1(n249), .Z(n238));
Q_AN02 U440 ( .A0(n267), .A1(n265), .Z(n244));
Q_INV U441 ( .A(n266), .Z(n242));
Q_AN02 U442 ( .A0(_zyM3L94_pbcFsm0_s[0]), .A1(n267), .Z(n247));
Q_INV U443 ( .A(n244), .Z(n251));
Q_FDP0 _zzM3L94_mdxP1_paddr_Dwen3_REG  ( .CK(_zyM3L94_pbcMevClk4), .D(n250), .Q(_zzM3L94_mdxP1_paddr_Dwen3), .QN( ));
Q_FDP0 _zzM3L94_mdxP1_pwrite_Dwen2_REG  ( .CK(_zyM3L94_pbcMevClk4), .D(n250), .Q(_zzM3L94_mdxP1_pwrite_Dwen2), .QN( ));
Q_FDP0 _zzM3L94_mdxP1_penable_Dwen1_REG  ( .CK(_zyM3L94_pbcMevClk4), .D(n248), .Q(_zzM3L94_mdxP1_penable_Dwen1), .QN( ));
Q_FDP0 _zzM3L94_mdxP1_psel_Dwen0_REG  ( .CK(_zyM3L94_pbcMevClk4), .D(n250), .Q(_zzM3L94_mdxP1_psel_Dwen0), .QN( ));
Q_FDP0 \_zyM3L94_pbcFsm0_s_REG[2] ( .CK(_zyM3L94_pbcMevClk4), .D(_zyM3L94_pbcFsm0_s[2]), .Q(_zyM3L94_pbcFsm0_s[2]), .QN(n233));
Q_XNR2 U449 ( .A0(n243), .A1(n266), .Z(n268));
Q_AN02 U450 ( .A0(n244), .A1(n200), .Z(n269));
Q_AN02 U451 ( .A0(n244), .A1(n202), .Z(n270));
Q_AN02 U452 ( .A0(n244), .A1(n204), .Z(n271));
Q_AN02 U453 ( .A0(n244), .A1(n206), .Z(n272));
Q_AN02 U454 ( .A0(n244), .A1(n208), .Z(n273));
Q_AN02 U455 ( .A0(n244), .A1(n210), .Z(n274));
Q_AN02 U456 ( .A0(n244), .A1(n212), .Z(n275));
Q_AN02 U457 ( .A0(n244), .A1(n297), .Z(n276));
Q_AN02 U458 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[19]), .Z(n277));
Q_AN02 U459 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[18]), .Z(n278));
Q_AN02 U460 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[17]), .Z(n279));
Q_AN02 U461 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[16]), .Z(n280));
Q_AN02 U462 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[15]), .Z(n281));
Q_AN02 U463 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[14]), .Z(n282));
Q_AN02 U464 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[13]), .Z(n283));
Q_AN02 U465 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[12]), .Z(n284));
Q_AN02 U466 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[11]), .Z(n285));
Q_AN02 U467 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[10]), .Z(n286));
Q_AN02 U468 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[9]), .Z(n287));
Q_AN02 U469 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[8]), .Z(n288));
Q_AN02 U470 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[7]), .Z(n289));
Q_AN02 U471 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[6]), .Z(n290));
Q_AN02 U472 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[5]), .Z(n291));
Q_AN02 U473 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[4]), .Z(n292));
Q_AN02 U474 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[3]), .Z(n293));
Q_AN02 U475 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[2]), .Z(n294));
Q_AN02 U476 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[1]), .Z(n295));
Q_AN02 U477 ( .A0(n249), .A1(_zyL94_iscX1c0_i0[0]), .Z(n296));
Q_OR02 U478 ( .A0(_zzpslverr_M3L26_bcSv2), .A1(n299), .Z(n298));
Q_NR02 U479 ( .A0(n301), .A1(n300), .Z(n299));
Q_OR03 U480 ( .A0(bus_timer[1]), .A1(bus_timer[0]), .A2(n302), .Z(n300));
Q_OR03 U481 ( .A0(bus_timer[4]), .A1(bus_timer[3]), .A2(n305), .Z(n301));
Q_OR03 U482 ( .A0(bus_timer[7]), .A1(n303), .A2(n304), .Z(n302));
Q_INV U483 ( .A(bus_timer[6]), .Z(n303));
Q_INV U484 ( .A(bus_timer[5]), .Z(n304));
Q_AO21 U485 ( .A0(n307), .A1(n306), .B0(n308), .Z(n230));
Q_NR02 U486 ( .A0(bus_timer[3]), .A1(bus_timer[2]), .Z(n306));
Q_AN02 U487 ( .A0(n312), .A1(n309), .Z(n307));
Q_OA21 U488 ( .A0(n311), .A1(n310), .B0(n312), .Z(n308));
Q_INV U489 ( .A(n313), .Z(n231));
Q_XNR2 U490 ( .A0(_zzM3L94_bcP1_EnD), .A1(_zzM3L94_bcP1_EnDNxt), .Z(n313));
Q_INV U491 ( .A(reset_n), .Z(n314));
Q_AN02 U492 ( .A0(n316), .A1(reset_n), .Z(n315));
Q_FDP0 _zzM3L46_mdxP0_pwdata_Dwen4_REG  ( .CK(clk), .D(n314), .Q(_zzM3L46_mdxP0_pwdata_Dwen4), .QN( ));
Q_FDP0 _zzM3L46_mdxP0_paddr_Dwen3_REG  ( .CK(clk), .D(n314), .Q(_zzM3L46_mdxP0_paddr_Dwen3), .QN( ));
Q_FDP0 _zzM3L46_mdxP0_pwrite_Dwen2_REG  ( .CK(clk), .D(n314), .Q(_zzM3L46_mdxP0_pwrite_Dwen2), .QN( ));
Q_FDP0 _zzM3L46_mdxP0_penable_Dwen1_REG  ( .CK(clk), .D(n314), .Q(_zzM3L46_mdxP0_penable_Dwen1), .QN( ));
Q_FDP0 _zzM3L46_mdxP0_psel_Dwen0_REG  ( .CK(clk), .D(n314), .Q(_zzM3L46_mdxP0_psel_Dwen0), .QN( ));
Q_XNR2 U498 ( .A0(_zzM3L46_bcP0_EnD), .A1(_zzM3L46_bcP0_EnDNxt), .Z(n316));
Q_NOT_TOUCH _zzqnt ( .sig());
ixc_assign _zz_strnp_0 ( _zy_simnet_psel_0_w$, psel);
ixc_assign _zz_strnp_1 ( _zy_simnet_penable_1_w$, penable);
ixc_assign_20 _zz_strnp_2 ( _zy_simnet_paddr_2_w$[0:19], paddr[19:0]);
ixc_assign_32 _zz_strnp_3 ( _zy_simnet_pwdata_3_w$[0:31], pwdata[31:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_pwrite_4_w$, pwrite);
Q_OR03 U505 ( .A0(_zyM3L104_pbcCapEn1), .A1(_zyM3L110_pbcCapEn2), .A2(_zyM3L121_pbcCapEn3), .Z(n325));
ixc_mevClk_2_0_0_1_0_2 _zzM3L94_pbcMevClk4 ( _zyM3L94_pbcMevClk4, { 
	_zyL94_iscX1c0_s, clk}, { _zyM3L94_pbcCapEn0, n325}, n324, n323, 
	_zyM3L94_pbcReq4, _zyM3L94_pbcBusy4, _zyM3L94_pbcWait4);
Q_OR03 U507 ( .A0(_zyM3L73_pbcCapEn6), .A1(_zyM3L79_pbcCapEn7), .A2(_zyM3L90_pbcCapEn8), .Z(n322));
ixc_mevClk_2_0_0_1_0_2 _zzM3L61_pbcMevClk9 ( _zyM3L61_pbcMevClk9, { 
	_zyL61_iscX2c0_s, clk}, { _zyM3L61_pbcCapEn5, n322}, n321, n320, 
	_zyM3L61_pbcReq9, _zyM3L61_pbcBusy9, _zyM3L61_pbcWait9);
ixc_sample_logic _zzpready_M3L25_bcSp0 ( _zzpready_M3L25_bcSv0, pready);
ixc_sample_logic_32 _zzprdata_M3L24_bcSp1 ( _zzprdata_M3L24_bcSv1[31:0], 
	prdata[31:0]);
ixc_sample_logic _zzpslverr_M3L26_bcSp2 ( _zzpslverr_M3L26_bcSv2, pslverr);
ixc_nba2BpD _zzM3L46_bcP0_DOnP ( _zzM3L46_bcP0_DOn, _zzM3L46_bcP0_EnDNxt, 
	_zzM3L46_bcP0_EnD);
ixc_nba2BpD _zzM3L94_bcP1_DOnP ( _zzM3L94_bcP1_DOn, _zzM3L94_bcP1_EnDNxt, 
	_zzM3L94_bcP1_EnD);
ixc_nba2BpD _zzM3L61_bcP2_DOnP ( _zzM3L61_bcP2_DOn, _zzM3L61_bcP2_EnDNxt, 
	_zzM3L61_bcP2_EnD);
ixc_sampleLT_8 _zzbus_timer_M3L29_bcSpLt7 ( _zzbus_timer_M3L29_bcSvLt7[7:0], 
	bus_timer[7:0]);
ixc_sampleLT_32 _zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSpLt8 ( 
	_zz_zydata_L96_tfiV1_M3_pbcG1_M3_bcSvLt8[31:0], 
	_zydata_L96_tfiV1_M3_pbcG1[31:0]);
ixc_sampleLT _zz_zyresponse_L97_tfiV2_M3_pbcG2_M3_bcSpLt9 ( 
	_zz_zyresponse_L97_tfiV2_M3_pbcG2_M3_bcSvLt9, 
	_zyresponse_L97_tfiV2_M3_pbcG2);
ixc_sampleLT _zz_zyresponse_L64_tfiV5_M3_pbcG5_M3_bcSpLt10 ( 
	_zz_zyresponse_L64_tfiV5_M3_pbcG5_M3_bcSvLt10, 
	_zyresponse_L64_tfiV5_M3_pbcG5);
ixc_capLoopXp _zzM3L10_bcBehEvalP0 ( _zzM3_bcBehEvalClk, n1,, _zzM3_bcBehHalt);
ixc_mdrOn _zzM3L46_mdxP0_OnP ( _zzM3L46_mdxP0_On, _zzM3L46_mdxP0_EnNxt, 
	_zzM3L46_mdxP0_En);
ixc_mdrOn _zzM3L94_mdxP1_OnP ( _zzM3L94_mdxP1_On, _zzM3L94_mdxP1_EnNxt, 
	_zzM3L94_mdxP1_En);
ixc_mdrOn _zzM3L61_mdxP2_OnP ( _zzM3L61_mdxP2_On, _zzM3L61_mdxP2_EnNxt, 
	_zzM3L61_mdxP2_En);
ixc_sampleLT _zzpsel_M3L19_mdxSpLt5 ( _zzpsel_M3L19_mdxSvLt5, psel);
ixc_sampleLT _zzpenable_M3L20_mdxSpLt6 ( _zzpenable_M3L20_mdxSvLt6, penable);
ixc_sampleLT _zzpwrite_M3L23_mdxSpLt7 ( _zzpwrite_M3L23_mdxSvLt7, pwrite);
ixc_sampleLT_20 _zzpaddr_M3L21_mdxSpLt8 ( _zzpaddr_M3L21_mdxSvLt8[19:0], 
	paddr[19:0]);
ixc_sampleLT_32 _zzpwdata_M3L22_mdxSpLt9 ( _zzpwdata_M3L22_mdxSvLt9[31:0], 
	pwdata[31:0]);
ixc_assign _zzmdx1 ( _zzmdxOne, n318);
ixc_assign _zzbc1 ( _zzbcOne, n317);
Q_FDP4EP _zzM3L46_bcP0_EnD_REG  ( .CK(clk), .CE(n314), .R(n319), .D(_zzM3L46_bcP0_EnDNxt), .Q(_zzM3L46_bcP0_EnD));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[7] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[7]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[6] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[6]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[5] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[5]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[4] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[4]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[3] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[3]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[2] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[2]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[1] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[1]));
Q_FDP4EP \_zzM3L46_bcP0_bus_timer_wr0_REG[0] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_bcP0_bus_timer_wr0[0]));
Q_FDP4EP _zzM3L46_mdxP0_En_REG  ( .CK(clk), .CE(n314), .R(n319), .D(_zzM3L46_mdxP0_EnNxt), .Q(_zzM3L46_mdxP0_En));
Q_FDP4EP _zzM3L46_mdxP0_psel_wr0_REG  ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_psel_wr0));
Q_FDP4EP _zzM3L46_mdxP0_penable_wr1_REG  ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_penable_wr1));
Q_FDP4EP _zzM3L46_mdxP0_pwrite_wr2_REG  ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwrite_wr2));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[19] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[19]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[18] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[18]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[17] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[17]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[16] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[16]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[15] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[15]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[14] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[14]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[13] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[13]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[12] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[12]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[11] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[11]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[10] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[10]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[9] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[9]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[8] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[8]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[7] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[7]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[6] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[6]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[5] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[5]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[4] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[4]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[3] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[3]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[2] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[2]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[1] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[1]));
Q_FDP4EP \_zzM3L46_mdxP0_paddr_wr3_REG[0] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_paddr_wr3[0]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[31] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[31]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[30] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[30]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[29] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[29]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[28] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[28]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[27] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[27]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[26] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[26]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[25] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[25]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[24] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[24]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[23] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[23]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[22] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[22]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[21] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[21]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[20] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[20]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[19] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[19]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[18] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[18]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[17] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[17]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[16] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[16]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[15] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[15]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[14] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[14]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[13] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[13]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[12] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[12]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[11] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[11]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[10] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[10]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[9] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[9]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[8] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[8]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[7] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[7]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[6] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[6]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[5] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[5]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[4] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[4]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[3] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[3]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[2] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[2]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[1] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[1]));
Q_FDP4EP \_zzM3L46_mdxP0_pwdata_wr4_REG[0] ( .CK(clk), .CE(n314), .R(n319), .D(n319), .Q(_zzM3L46_mdxP0_pwdata_wr4[0]));
Q_INV U595 ( .A(n315), .Z(n327));
Q_FDP4EP _zzM3L46_bcP0_bus_timer_Dwen0_REG  ( .CK(clk), .CE(n327), .R(n319), .D(n314), .Q(_zzM3L46_bcP0_bus_timer_Dwen0));
Q_FDP4EP _zyL94_iscX1c0_f_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zyL94_iscX1c0_n), .Q(_zyL94_iscX1c0_f));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[31] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[31]), .Q(_zyL94_iscX1c0_o1[31]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[30] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[30]), .Q(_zyL94_iscX1c0_o1[30]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[29] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[29]), .Q(_zyL94_iscX1c0_o1[29]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[28] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[28]), .Q(_zyL94_iscX1c0_o1[28]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[27] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[27]), .Q(_zyL94_iscX1c0_o1[27]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[26] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[26]), .Q(_zyL94_iscX1c0_o1[26]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[25] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[25]), .Q(_zyL94_iscX1c0_o1[25]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[24] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[24]), .Q(_zyL94_iscX1c0_o1[24]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[23] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[23]), .Q(_zyL94_iscX1c0_o1[23]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[22] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[22]), .Q(_zyL94_iscX1c0_o1[22]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[21] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[21]), .Q(_zyL94_iscX1c0_o1[21]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[20] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[20]), .Q(_zyL94_iscX1c0_o1[20]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[19] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[19]), .Q(_zyL94_iscX1c0_o1[19]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[18] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[18]), .Q(_zyL94_iscX1c0_o1[18]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[17] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[17]), .Q(_zyL94_iscX1c0_o1[17]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[16] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[16]), .Q(_zyL94_iscX1c0_o1[16]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[15] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[15]), .Q(_zyL94_iscX1c0_o1[15]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[14] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[14]), .Q(_zyL94_iscX1c0_o1[14]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[13] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[13]), .Q(_zyL94_iscX1c0_o1[13]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[12] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[12]), .Q(_zyL94_iscX1c0_o1[12]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[11] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[11]), .Q(_zyL94_iscX1c0_o1[11]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[10] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[10]), .Q(_zyL94_iscX1c0_o1[10]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[9] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[9]), .Q(_zyL94_iscX1c0_o1[9]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[8] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[8]), .Q(_zyL94_iscX1c0_o1[8]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[7] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[7]), .Q(_zyL94_iscX1c0_o1[7]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[6] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[6]), .Q(_zyL94_iscX1c0_o1[6]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[5] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[5]), .Q(_zyL94_iscX1c0_o1[5]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[4] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[4]), .Q(_zyL94_iscX1c0_o1[4]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[3] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[3]), .Q(_zyL94_iscX1c0_o1[3]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[2] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[2]), .Q(_zyL94_iscX1c0_o1[2]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[1] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[1]), .Q(_zyL94_iscX1c0_o1[1]));
Q_FDP4EP \_zyL94_iscX1c0_o1_REG[0] ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zydata_L96_tfiV1_M3_pbcG1[0]), .Q(_zyL94_iscX1c0_o1[0]));
Q_FDP4EP _zyL94_iscX1c0_o2_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(_zyresponse_L97_tfiV2_M3_pbcG2), .Q(_zyL94_iscX1c0_o2));
Q_FDP4EP _zzM3L94_bcP1_EnD_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(_zzM3L94_bcP1_EnDNxt), .Q(_zzM3L94_bcP1_EnD));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[31] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[31]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[31]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[30] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[30]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[30]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[29] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[29]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[29]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[28] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[28]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[28]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[27] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[27]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[27]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[26] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[26]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[26]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[25] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[25]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[25]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[24] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[24]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[24]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[23] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[23]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[23]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[22] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[22]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[22]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[21] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[21]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[21]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[20] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[20]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[20]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[19] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[19]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[19]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[18] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[18]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[18]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[17] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[17]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[17]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[16] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[16]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[16]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[15] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[15]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[15]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[14] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[14]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[14]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[13] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[13]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[13]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[12] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[12]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[12]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[11] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[11]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[11]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[10] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[10]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[10]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[9] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[9]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[9]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[8] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[8]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[8]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[7] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[7]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[7]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[6] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[6]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[6]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[5] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[5]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[5]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[4] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[4]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[4]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[3] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[3]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[3]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[2] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[2]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[2]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[1] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[1]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[1]));
Q_FDP4EP \_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1_REG[0] ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(_zzprdata_M3L24_bcSv1[0]), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_wr1[0]));
Q_FDP4EP _zzM3L94_mdxP1_En_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n248), .R(n319), .D(_zzM3L94_mdxP1_EnNxt), .Q(_zzM3L94_mdxP1_En));
Q_FDP4EP _zzM3L94_mdxP1_pwrite_wr2_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n319), .Q(_zzM3L94_mdxP1_pwrite_wr2));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[63] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[63]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[63]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[62] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[62]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[62]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[61] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[61]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[61]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[60] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[60]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[60]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[59] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[59]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[59]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[58] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[58]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[58]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[57] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[57]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[57]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[56] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[56]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[56]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[55] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[55]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[55]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[54] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[54]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[54]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[53] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[53]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[53]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[52] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[52]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[52]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[51] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[51]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[51]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[50] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[50]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[50]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[49] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[49]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[49]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[48] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[48]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[48]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[47] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[47]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[47]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[46] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[46]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[46]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[45] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[45]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[45]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[44] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[44]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[44]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[43] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[43]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[43]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[42] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[42]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[42]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[41] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[41]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[41]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[40] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[40]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[40]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[39] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[39]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[39]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[38] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[38]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[38]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[37] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[37]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[37]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[36] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[36]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[36]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[35] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[35]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[35]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[34] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[34]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[34]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[33] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[33]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[33]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[32] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[32]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[32]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[31] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[31]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[31]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[30] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[30]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[30]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[29] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[29]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[29]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[28] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[28]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[28]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[27] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[27]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[27]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[26] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[26]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[26]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[25] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[25]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[25]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[24] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[24]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[24]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[23] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[23]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[23]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[22] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[22]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[22]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[21] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[21]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[21]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[20] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[20]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[20]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[19] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[19]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[19]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[18] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[18]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[18]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[17] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[17]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[17]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[16] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[16]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[16]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[15] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[15]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[15]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[14] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[14]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[14]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[13] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[13]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[13]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[12] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[12]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[12]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[11] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[11]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[11]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[10] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[10]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[10]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[9] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[9]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[9]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[8] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[8]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[8]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[7] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[7]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[7]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[6] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[6]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[6]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[5] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[5]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[5]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[4] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[4]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[4]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[3] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[3]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[3]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[2] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[2]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[2]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[1] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[1]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[1]));
Q_FDP4EP \_zyaddr_L95_tfiV0_M3_pbcG0_REG[0] ( .CK(_zyM3L94_pbcMevClk4), .CE(n238), .R(n319), .D(_zyL94_iscX1c0_i0[0]), .Q(_zyaddr_L95_tfiV0_M3_pbcG0[0]));
Q_INV U730 ( .A(_zyL94_iscX1c0_n), .Z(n328));
Q_FDP4EP _zyL94_iscX1c0_n_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n237), .R(n319), .D(n328), .Q(_zyL94_iscX1c0_n));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[7] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n269), .Q(_zzM3L94_bcP1_bus_timer_wr0[7]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[6] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n270), .Q(_zzM3L94_bcP1_bus_timer_wr0[6]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[5] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n271), .Q(_zzM3L94_bcP1_bus_timer_wr0[5]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[4] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n272), .Q(_zzM3L94_bcP1_bus_timer_wr0[4]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[3] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n273), .Q(_zzM3L94_bcP1_bus_timer_wr0[3]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[2] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n274), .Q(_zzM3L94_bcP1_bus_timer_wr0[2]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[1] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n275), .Q(_zzM3L94_bcP1_bus_timer_wr0[1]));
Q_FDP4EP \_zzM3L94_bcP1_bus_timer_wr0_REG[0] ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n276), .Q(_zzM3L94_bcP1_bus_timer_wr0[0]));
Q_FDP4EP _zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_wr2_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n246), .R(n319), .D(n298), .Q(_zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_wr2));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[19] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n277), .Q(_zzM3L94_mdxP1_paddr_wr3[19]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[18] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n278), .Q(_zzM3L94_mdxP1_paddr_wr3[18]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[17] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n279), .Q(_zzM3L94_mdxP1_paddr_wr3[17]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[16] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n280), .Q(_zzM3L94_mdxP1_paddr_wr3[16]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[15] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n281), .Q(_zzM3L94_mdxP1_paddr_wr3[15]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[14] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n282), .Q(_zzM3L94_mdxP1_paddr_wr3[14]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[13] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n283), .Q(_zzM3L94_mdxP1_paddr_wr3[13]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[12] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n284), .Q(_zzM3L94_mdxP1_paddr_wr3[12]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[11] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n285), .Q(_zzM3L94_mdxP1_paddr_wr3[11]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[10] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n286), .Q(_zzM3L94_mdxP1_paddr_wr3[10]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[9] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n287), .Q(_zzM3L94_mdxP1_paddr_wr3[9]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[8] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n288), .Q(_zzM3L94_mdxP1_paddr_wr3[8]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[7] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n289), .Q(_zzM3L94_mdxP1_paddr_wr3[7]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[6] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n290), .Q(_zzM3L94_mdxP1_paddr_wr3[6]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[5] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n291), .Q(_zzM3L94_mdxP1_paddr_wr3[5]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[4] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n292), .Q(_zzM3L94_mdxP1_paddr_wr3[4]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[3] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n293), .Q(_zzM3L94_mdxP1_paddr_wr3[3]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[2] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n294), .Q(_zzM3L94_mdxP1_paddr_wr3[2]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[1] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n295), .Q(_zzM3L94_mdxP1_paddr_wr3[1]));
Q_FDP4EP \_zzM3L94_mdxP1_paddr_wr3_REG[0] ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n296), .Q(_zzM3L94_mdxP1_paddr_wr3[0]));
Q_FDP4EP _zyM3L94_pbcCapEn0_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n236), .R(n319), .D(n239), .Q(_zyM3L94_pbcCapEn0));
Q_FDP4EP _zyM3L104_pbcCapEn1_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n235), .R(n319), .D(n240), .Q(_zyM3L104_pbcCapEn1));
Q_FDP4EP _zyM3L110_pbcCapEn2_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n234), .R(n319), .D(n244), .Q(_zyM3L110_pbcCapEn2));
Q_INV U764 ( .A(n258), .Z(n329));
Q_FDP4EP _zyM3L121_pbcCapEn3_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n329), .R(n319), .D(n241), .Q(_zyM3L121_pbcCapEn3));
Q_FDP4EP \_zyM3L94_pbcFsm0_s_REG[1] ( .CK(_zyM3L94_pbcMevClk4), .CE(n233), .R(n319), .D(n268), .Q(_zyM3L94_pbcFsm0_s[1]));
Q_INV U767 ( .A(_zyM3L94_pbcFsm0_s[1]), .Z(n262));
Q_FDP4EP \_zyM3L94_pbcFsm0_s_REG[0] ( .CK(_zyM3L94_pbcMevClk4), .CE(n233), .R(n319), .D(n242), .Q(_zyM3L94_pbcFsm0_s[0]));
Q_INV U769 ( .A(_zyM3L94_pbcFsm0_s[0]), .Z(n240));
Q_FDP4EP _zzM3L94_bcP1_bus_timer_Dwen0_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n232), .R(n319), .D(n245), .Q(_zzM3L94_bcP1_bus_timer_Dwen0));
Q_INV U771 ( .A(n256), .Z(n330));
Q_FDP4EP _zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_Dwen1_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n330), .R(n319), .D(n246), .Q(_zzM3L94_bcP1__zydata_L96_tfiV1_M3_pbcG1_Dwen1));
Q_FDP4EP _zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_Dwen2_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n330), .R(n319), .D(n246), .Q(_zzM3L94_bcP1__zyresponse_L97_tfiV2_M3_pbcG2_Dwen2));
Q_FDP4EP _zzM3L94_mdxP1_psel_wr0_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n250), .R(n319), .D(n249), .Q(_zzM3L94_mdxP1_psel_wr0));
Q_FDP4EP _zzM3L94_mdxP1_penable_wr1_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n248), .R(n319), .D(n247), .Q(_zzM3L94_mdxP1_penable_wr1));
Q_FDP4EP _zyM3L94_pbcEn10_REG  ( .CK(_zyM3L94_pbcMevClk4), .CE(n245), .R(n319), .D(n251), .Q(_zyM3L94_pbcEn10));
Q_FDP4EP _zyL61_iscX2c0_f_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n107), .R(n319), .D(_zyL61_iscX2c0_n), .Q(_zyL61_iscX2c0_f));
Q_FDP4EP _zyL61_iscX2c0_o2_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n107), .R(n319), .D(_zyresponse_L64_tfiV5_M3_pbcG5), .Q(_zyL61_iscX2c0_o2));
Q_FDP4EP _zzM3L61_bcP2_EnD_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(_zzM3L61_bcP2_EnDNxt), .Q(_zzM3L61_bcP2_EnD));
Q_FDP4EP _zzM3L61_mdxP2_En_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n118), .R(n319), .D(_zzM3L61_mdxP2_EnNxt), .Q(_zzM3L61_mdxP2_En));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[63] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[63]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[63]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[62] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[62]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[62]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[61] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[61]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[61]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[60] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[60]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[60]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[59] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[59]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[59]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[58] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[58]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[58]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[57] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[57]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[57]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[56] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[56]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[56]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[55] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[55]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[55]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[54] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[54]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[54]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[53] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[53]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[53]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[52] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[52]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[52]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[51] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[51]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[51]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[50] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[50]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[50]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[49] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[49]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[49]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[48] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[48]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[48]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[47] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[47]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[47]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[46] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[46]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[46]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[45] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[45]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[45]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[44] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[44]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[44]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[43] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[43]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[43]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[42] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[42]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[42]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[41] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[41]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[41]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[40] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[40]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[40]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[39] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[39]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[39]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[38] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[38]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[38]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[37] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[37]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[37]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[36] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[36]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[36]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[35] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[35]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[35]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[34] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[34]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[34]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[33] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[33]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[33]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[32] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[32]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[32]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[31] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[31]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[31]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[30] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[30]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[30]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[29] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[29]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[29]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[28] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[28]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[28]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[27] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[27]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[27]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[26] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[26]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[26]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[25] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[25]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[25]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[24] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[24]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[24]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[23] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[23]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[23]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[22] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[22]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[22]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[21] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[21]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[21]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[20] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[20]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[20]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[19] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[19]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[19]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[18] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[18]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[18]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[17] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[17]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[17]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[16] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[16]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[16]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[15] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[15]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[15]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[14] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[14]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[14]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[13] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[13]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[13]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[12] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[12]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[12]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[11] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[11]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[11]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[10] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[10]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[10]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[9] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[9]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[9]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[8] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[8]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[8]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[7] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[7]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[7]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[6] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[6]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[6]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[5] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[5]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[5]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[4] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[4]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[4]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[3] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[3]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[3]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[2] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[2]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[2]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[1] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[1]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[1]));
Q_FDP4EP \_zyaddr_L62_tfiV3_M3_pbcG3_REG[0] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i0[0]), .Q(_zyaddr_L62_tfiV3_M3_pbcG3[0]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[31] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[31]), .Q(_zydata_L63_tfiV4_M3_pbcG4[31]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[30] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[30]), .Q(_zydata_L63_tfiV4_M3_pbcG4[30]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[29] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[29]), .Q(_zydata_L63_tfiV4_M3_pbcG4[29]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[28] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[28]), .Q(_zydata_L63_tfiV4_M3_pbcG4[28]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[27] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[27]), .Q(_zydata_L63_tfiV4_M3_pbcG4[27]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[26] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[26]), .Q(_zydata_L63_tfiV4_M3_pbcG4[26]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[25] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[25]), .Q(_zydata_L63_tfiV4_M3_pbcG4[25]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[24] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[24]), .Q(_zydata_L63_tfiV4_M3_pbcG4[24]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[23] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[23]), .Q(_zydata_L63_tfiV4_M3_pbcG4[23]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[22] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[22]), .Q(_zydata_L63_tfiV4_M3_pbcG4[22]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[21] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[21]), .Q(_zydata_L63_tfiV4_M3_pbcG4[21]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[20] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[20]), .Q(_zydata_L63_tfiV4_M3_pbcG4[20]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[19] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[19]), .Q(_zydata_L63_tfiV4_M3_pbcG4[19]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[18] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[18]), .Q(_zydata_L63_tfiV4_M3_pbcG4[18]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[17] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[17]), .Q(_zydata_L63_tfiV4_M3_pbcG4[17]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[16] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[16]), .Q(_zydata_L63_tfiV4_M3_pbcG4[16]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[15] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[15]), .Q(_zydata_L63_tfiV4_M3_pbcG4[15]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[14] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[14]), .Q(_zydata_L63_tfiV4_M3_pbcG4[14]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[13] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[13]), .Q(_zydata_L63_tfiV4_M3_pbcG4[13]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[12] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[12]), .Q(_zydata_L63_tfiV4_M3_pbcG4[12]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[11] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[11]), .Q(_zydata_L63_tfiV4_M3_pbcG4[11]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[10] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[10]), .Q(_zydata_L63_tfiV4_M3_pbcG4[10]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[9] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[9]), .Q(_zydata_L63_tfiV4_M3_pbcG4[9]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[8] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[8]), .Q(_zydata_L63_tfiV4_M3_pbcG4[8]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[7] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[7]), .Q(_zydata_L63_tfiV4_M3_pbcG4[7]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[6] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[6]), .Q(_zydata_L63_tfiV4_M3_pbcG4[6]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[5] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[5]), .Q(_zydata_L63_tfiV4_M3_pbcG4[5]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[4] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[4]), .Q(_zydata_L63_tfiV4_M3_pbcG4[4]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[3] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[3]), .Q(_zydata_L63_tfiV4_M3_pbcG4[3]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[2] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[2]), .Q(_zydata_L63_tfiV4_M3_pbcG4[2]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[1] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[1]), .Q(_zydata_L63_tfiV4_M3_pbcG4[1]));
Q_FDP4EP \_zydata_L63_tfiV4_M3_pbcG4_REG[0] ( .CK(_zyM3L61_pbcMevClk9), .CE(n108), .R(n319), .D(_zyL61_iscX2c0_i1[0]), .Q(_zydata_L63_tfiV4_M3_pbcG4[0]));
Q_INV U877 ( .A(_zyL61_iscX2c0_n), .Z(n331));
Q_FDP4EP _zyL61_iscX2c0_n_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n107), .R(n319), .D(n331), .Q(_zyL61_iscX2c0_n));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[7] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n140), .Q(_zzM3L61_bcP2_bus_timer_wr0[7]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[6] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n141), .Q(_zzM3L61_bcP2_bus_timer_wr0[6]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[5] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n142), .Q(_zzM3L61_bcP2_bus_timer_wr0[5]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[4] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n143), .Q(_zzM3L61_bcP2_bus_timer_wr0[4]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[3] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n144), .Q(_zzM3L61_bcP2_bus_timer_wr0[3]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[2] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n145), .Q(_zzM3L61_bcP2_bus_timer_wr0[2]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[1] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n146), .Q(_zzM3L61_bcP2_bus_timer_wr0[1]));
Q_FDP4EP \_zzM3L61_bcP2_bus_timer_wr0_REG[0] ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n147), .Q(_zzM3L61_bcP2_bus_timer_wr0[0]));
Q_FDP4EP _zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_wr1_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n116), .R(n319), .D(n214), .Q(_zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_wr1));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[19] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n148), .Q(_zzM3L61_mdxP2_paddr_wr3[19]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[18] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n149), .Q(_zzM3L61_mdxP2_paddr_wr3[18]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[17] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n150), .Q(_zzM3L61_mdxP2_paddr_wr3[17]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[16] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n151), .Q(_zzM3L61_mdxP2_paddr_wr3[16]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[15] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n152), .Q(_zzM3L61_mdxP2_paddr_wr3[15]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[14] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n153), .Q(_zzM3L61_mdxP2_paddr_wr3[14]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[13] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n154), .Q(_zzM3L61_mdxP2_paddr_wr3[13]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[12] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n155), .Q(_zzM3L61_mdxP2_paddr_wr3[12]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[11] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n156), .Q(_zzM3L61_mdxP2_paddr_wr3[11]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[10] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n157), .Q(_zzM3L61_mdxP2_paddr_wr3[10]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[9] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n158), .Q(_zzM3L61_mdxP2_paddr_wr3[9]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[8] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n159), .Q(_zzM3L61_mdxP2_paddr_wr3[8]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[7] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n160), .Q(_zzM3L61_mdxP2_paddr_wr3[7]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[6] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n161), .Q(_zzM3L61_mdxP2_paddr_wr3[6]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[5] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n162), .Q(_zzM3L61_mdxP2_paddr_wr3[5]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[4] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n163), .Q(_zzM3L61_mdxP2_paddr_wr3[4]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[3] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n164), .Q(_zzM3L61_mdxP2_paddr_wr3[3]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[2] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n165), .Q(_zzM3L61_mdxP2_paddr_wr3[2]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[1] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n166), .Q(_zzM3L61_mdxP2_paddr_wr3[1]));
Q_FDP4EP \_zzM3L61_mdxP2_paddr_wr3_REG[0] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n167), .Q(_zzM3L61_mdxP2_paddr_wr3[0]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[31] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n168), .Q(_zzM3L61_mdxP2_pwdata_wr4[31]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[30] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n169), .Q(_zzM3L61_mdxP2_pwdata_wr4[30]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[29] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n170), .Q(_zzM3L61_mdxP2_pwdata_wr4[29]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[28] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n171), .Q(_zzM3L61_mdxP2_pwdata_wr4[28]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[27] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n172), .Q(_zzM3L61_mdxP2_pwdata_wr4[27]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[26] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n173), .Q(_zzM3L61_mdxP2_pwdata_wr4[26]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[25] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n174), .Q(_zzM3L61_mdxP2_pwdata_wr4[25]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[24] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n175), .Q(_zzM3L61_mdxP2_pwdata_wr4[24]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[23] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n176), .Q(_zzM3L61_mdxP2_pwdata_wr4[23]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[22] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n177), .Q(_zzM3L61_mdxP2_pwdata_wr4[22]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[21] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n178), .Q(_zzM3L61_mdxP2_pwdata_wr4[21]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[20] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n179), .Q(_zzM3L61_mdxP2_pwdata_wr4[20]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[19] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n180), .Q(_zzM3L61_mdxP2_pwdata_wr4[19]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[18] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n181), .Q(_zzM3L61_mdxP2_pwdata_wr4[18]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[17] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n182), .Q(_zzM3L61_mdxP2_pwdata_wr4[17]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[16] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n183), .Q(_zzM3L61_mdxP2_pwdata_wr4[16]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[15] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n184), .Q(_zzM3L61_mdxP2_pwdata_wr4[15]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[14] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n185), .Q(_zzM3L61_mdxP2_pwdata_wr4[14]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[13] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n186), .Q(_zzM3L61_mdxP2_pwdata_wr4[13]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[12] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n187), .Q(_zzM3L61_mdxP2_pwdata_wr4[12]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[11] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n188), .Q(_zzM3L61_mdxP2_pwdata_wr4[11]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[10] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n189), .Q(_zzM3L61_mdxP2_pwdata_wr4[10]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[9] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n190), .Q(_zzM3L61_mdxP2_pwdata_wr4[9]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[8] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n191), .Q(_zzM3L61_mdxP2_pwdata_wr4[8]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[7] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n192), .Q(_zzM3L61_mdxP2_pwdata_wr4[7]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[6] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n193), .Q(_zzM3L61_mdxP2_pwdata_wr4[6]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[5] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n194), .Q(_zzM3L61_mdxP2_pwdata_wr4[5]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[4] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n195), .Q(_zzM3L61_mdxP2_pwdata_wr4[4]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[3] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n196), .Q(_zzM3L61_mdxP2_pwdata_wr4[3]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[2] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n197), .Q(_zzM3L61_mdxP2_pwdata_wr4[2]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[1] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n198), .Q(_zzM3L61_mdxP2_pwdata_wr4[1]));
Q_FDP4EP \_zzM3L61_mdxP2_pwdata_wr4_REG[0] ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n199), .Q(_zzM3L61_mdxP2_pwdata_wr4[0]));
Q_FDP4EP _zyM3L61_pbcCapEn5_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n106), .R(n319), .D(n109), .Q(_zyM3L61_pbcCapEn5));
Q_FDP4EP _zyM3L73_pbcCapEn6_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n105), .R(n319), .D(n110), .Q(_zyM3L73_pbcCapEn6));
Q_FDP4EP _zyM3L79_pbcCapEn7_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n104), .R(n319), .D(n114), .Q(_zyM3L79_pbcCapEn7));
Q_INV U943 ( .A(n129), .Z(n332));
Q_FDP4EP _zyM3L90_pbcCapEn8_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n332), .R(n319), .D(n111), .Q(_zyM3L90_pbcCapEn8));
Q_FDP4EP \_zyM3L61_pbcFsm2_s_REG[1] ( .CK(_zyM3L61_pbcMevClk9), .CE(n103), .R(n319), .D(n139), .Q(_zyM3L61_pbcFsm2_s[1]));
Q_INV U946 ( .A(_zyM3L61_pbcFsm2_s[1]), .Z(n133));
Q_FDP4EP \_zyM3L61_pbcFsm2_s_REG[0] ( .CK(_zyM3L61_pbcMevClk9), .CE(n103), .R(n319), .D(n112), .Q(_zyM3L61_pbcFsm2_s[0]));
Q_INV U948 ( .A(_zyM3L61_pbcFsm2_s[0]), .Z(n110));
Q_FDP4EP _zzM3L61_bcP2_bus_timer_Dwen0_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n102), .R(n319), .D(n115), .Q(_zzM3L61_bcP2_bus_timer_Dwen0));
Q_INV U950 ( .A(n127), .Z(n333));
Q_FDP4EP _zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_Dwen1_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n333), .R(n319), .D(n116), .Q(_zzM3L61_bcP2__zyresponse_L64_tfiV5_M3_pbcG5_Dwen1));
Q_FDP4EP _zzM3L61_mdxP2_psel_wr0_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n119), .Q(_zzM3L61_mdxP2_psel_wr0));
Q_FDP4EP _zzM3L61_mdxP2_penable_wr1_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n118), .R(n319), .D(n117), .Q(_zzM3L61_mdxP2_penable_wr1));
Q_FDP4EP _zzM3L61_mdxP2_pwrite_wr2_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n120), .R(n319), .D(n119), .Q(_zzM3L61_mdxP2_pwrite_wr2));
Q_FDP4EP _zyM3L61_pbcEn11_REG  ( .CK(_zyM3L61_pbcMevClk9), .CE(n115), .R(n319), .D(n121), .Q(_zyM3L61_pbcEn11));
Q_FDP4EP \_zzM3_bcBehEval_REG[31] ( .CK(_zzM3_bcBehEvalClk), .CE(n22), .R(n319), .D(_zzM3_bcBehHalt), .Q(_zzM3_bcBehEval[31]));
Q_INV U957 ( .A(_zzM3_bcBehEval[30]), .Z(n334));
Q_FDP4EP \_zzM3_bcBehEval_REG[30] ( .CK(_zzM3_bcBehEvalClk), .CE(n2), .R(n319), .D(n334), .Q(_zzM3_bcBehEval[30]));
Q_FDP4EP \_zzM3_bcBehEval_REG[29] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n24), .Q(_zzM3_bcBehEval[29]));
Q_FDP4EP \_zzM3_bcBehEval_REG[28] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n26), .Q(_zzM3_bcBehEval[28]));
Q_FDP4EP \_zzM3_bcBehEval_REG[27] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n28), .Q(_zzM3_bcBehEval[27]));
Q_FDP4EP \_zzM3_bcBehEval_REG[26] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n30), .Q(_zzM3_bcBehEval[26]));
Q_FDP4EP \_zzM3_bcBehEval_REG[25] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n32), .Q(_zzM3_bcBehEval[25]));
Q_FDP4EP \_zzM3_bcBehEval_REG[24] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n34), .Q(_zzM3_bcBehEval[24]));
Q_FDP4EP \_zzM3_bcBehEval_REG[23] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n36), .Q(_zzM3_bcBehEval[23]));
Q_FDP4EP \_zzM3_bcBehEval_REG[22] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n38), .Q(_zzM3_bcBehEval[22]));
Q_FDP4EP \_zzM3_bcBehEval_REG[21] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n40), .Q(_zzM3_bcBehEval[21]));
Q_FDP4EP \_zzM3_bcBehEval_REG[20] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n42), .Q(_zzM3_bcBehEval[20]));
Q_FDP4EP \_zzM3_bcBehEval_REG[19] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n44), .Q(_zzM3_bcBehEval[19]));
Q_FDP4EP \_zzM3_bcBehEval_REG[18] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n46), .Q(_zzM3_bcBehEval[18]));
Q_FDP4EP \_zzM3_bcBehEval_REG[17] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n48), .Q(_zzM3_bcBehEval[17]));
Q_FDP4EP \_zzM3_bcBehEval_REG[16] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n50), .Q(_zzM3_bcBehEval[16]));
Q_FDP4EP \_zzM3_bcBehEval_REG[15] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n52), .Q(_zzM3_bcBehEval[15]));
Q_FDP4EP \_zzM3_bcBehEval_REG[14] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n54), .Q(_zzM3_bcBehEval[14]));
Q_FDP4EP \_zzM3_bcBehEval_REG[13] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n56), .Q(_zzM3_bcBehEval[13]));
Q_FDP4EP \_zzM3_bcBehEval_REG[12] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n58), .Q(_zzM3_bcBehEval[12]));
Q_FDP4EP \_zzM3_bcBehEval_REG[11] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n60), .Q(_zzM3_bcBehEval[11]));
Q_FDP4EP \_zzM3_bcBehEval_REG[10] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n62), .Q(_zzM3_bcBehEval[10]));
Q_FDP4EP \_zzM3_bcBehEval_REG[9] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n64), .Q(_zzM3_bcBehEval[9]));
Q_FDP4EP \_zzM3_bcBehEval_REG[8] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n66), .Q(_zzM3_bcBehEval[8]));
Q_FDP4EP \_zzM3_bcBehEval_REG[7] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n68), .Q(_zzM3_bcBehEval[7]));
Q_FDP4EP \_zzM3_bcBehEval_REG[6] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n70), .Q(_zzM3_bcBehEval[6]));
Q_FDP4EP \_zzM3_bcBehEval_REG[5] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n72), .Q(_zzM3_bcBehEval[5]));
Q_FDP4EP \_zzM3_bcBehEval_REG[4] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n74), .Q(_zzM3_bcBehEval[4]));
Q_FDP4EP \_zzM3_bcBehEval_REG[3] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n76), .Q(_zzM3_bcBehEval[3]));
Q_FDP4EP \_zzM3_bcBehEval_REG[2] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n78), .Q(_zzM3_bcBehEval[2]));
Q_FDP4EP \_zzM3_bcBehEval_REG[1] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n80), .Q(_zzM3_bcBehEval[1]));
Q_INV U988 ( .A(_zzM3_bcBehEval[0]), .Z(n335));
Q_FDP4EP \_zzM3_bcBehEval_REG[0] ( .CK(_zzM3_bcBehEvalClk), .CE(n21), .R(n319), .D(n335), .Q(_zzM3_bcBehEval[0]));
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
