
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module IXC_SV_GFIFO_VXE_256 ( rdCnt);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input [63:0] rdCnt;
wire hasMultiLevelGFIFO;
wire GFreq;
wire [19:0] GFcbid;
wire [11:0] GFlen;
wire [511:0] GFidata;
wire GFtsReq;
wire GFfull;
wire LBreq;
wire LBempty;
wire LBfull;
wire flushTbc;
wire [63:0] timeStampPkt;
wire svGFbusy1;
wire svGFbusy2;
`_2_ wire GFtsAdd;
wire [3:0] LBrd;
wire [3:0] LBwr;
wire [3:0] LBwrI;
wire [3:0] LBfill;
`_2_ wire [11:0] argLen;
`_2_ wire [18:0] wLen;
`_2_ wire [17:0] rLen;
`_2_ wire wSync;
`_2_ wire rSync;
`_2_ wire [543:0] xdata;
`_2_ wire [63:0] wrtCnt;
`_2_ wire [63:0] wrtCntD;
wire [7:0] ackId;
wire [7:0] ackIdNew;
wire ackClk;
wire [17:0] ackLen;
`_2_ wire [14:0] ofifoAddr0;
`_2_ wire [14:0] ofifoAddr0N;
`_2_ wire [14:0] ofifoAddr1;
`_2_ wire [14:0] ofifoAddr1N;
`_2_ wire [14:0] ofifoAddr2;
`_2_ wire [14:0] ofifoAddr2N;
`_2_ wire [767:0] ofifoData;
`_2_ wire [767:0] ofifoDataN;
`_2_ wire [5:0] writeLen;
`_2_ wire reqD;
`_2_ wire GFfullD;
`_2_ wire [4:0] oFill;
`_2_ wire [4:0] oFillN;
`_2_ wire [14:0] ofifoWptr;
`_2_ wire [14:0] ofifoWptrN;
`_2_ wire [7:0] shiftCount;
`_2_ wire [767:0] shiftedXdata;
wire gfTsReqO;
wire [63:0] gfTsValO;
wire gfTsEn;
Q_RDN U0 ( .Z(GFcbid[19]));
Q_RDN U1 ( .Z(GFcbid[18]));
Q_RDN U2 ( .Z(GFcbid[17]));
Q_RDN U3 ( .Z(GFcbid[16]));
Q_RDN U4 ( .Z(GFcbid[15]));
Q_RDN U5 ( .Z(GFcbid[14]));
Q_RDN U6 ( .Z(GFcbid[13]));
Q_RDN U7 ( .Z(GFcbid[12]));
Q_RDN U8 ( .Z(GFcbid[11]));
Q_RDN U9 ( .Z(GFcbid[10]));
Q_RDN U10 ( .Z(GFcbid[9]));
Q_RDN U11 ( .Z(GFcbid[8]));
Q_RDN U12 ( .Z(GFcbid[7]));
Q_RDN U13 ( .Z(GFcbid[6]));
Q_RDN U14 ( .Z(GFcbid[5]));
Q_RDN U15 ( .Z(GFcbid[4]));
Q_RDN U16 ( .Z(GFcbid[3]));
Q_RDN U17 ( .Z(GFcbid[2]));
Q_RDN U18 ( .Z(GFcbid[1]));
Q_RDN U19 ( .Z(GFcbid[0]));
Q_RDN U20 ( .Z(GFlen[11]));
Q_RDN U21 ( .Z(GFlen[10]));
Q_RDN U22 ( .Z(GFlen[9]));
Q_RDN U23 ( .Z(GFlen[8]));
Q_RDN U24 ( .Z(GFlen[7]));
Q_RDN U25 ( .Z(GFlen[6]));
Q_RDN U26 ( .Z(GFlen[5]));
Q_RDN U27 ( .Z(GFlen[4]));
Q_RDN U28 ( .Z(GFlen[3]));
Q_RDN U29 ( .Z(GFlen[2]));
Q_RDN U30 ( .Z(GFlen[1]));
Q_RDN U31 ( .Z(GFlen[0]));
Q_RDN U32 ( .Z(GFidata[511]));
Q_RDN U33 ( .Z(GFidata[510]));
Q_RDN U34 ( .Z(GFidata[509]));
Q_RDN U35 ( .Z(GFidata[508]));
Q_RDN U36 ( .Z(GFidata[507]));
Q_RDN U37 ( .Z(GFidata[506]));
Q_RDN U38 ( .Z(GFidata[505]));
Q_RDN U39 ( .Z(GFidata[504]));
Q_RDN U40 ( .Z(GFidata[503]));
Q_RDN U41 ( .Z(GFidata[502]));
Q_RDN U42 ( .Z(GFidata[501]));
Q_RDN U43 ( .Z(GFidata[500]));
Q_RDN U44 ( .Z(GFidata[499]));
Q_RDN U45 ( .Z(GFidata[498]));
Q_RDN U46 ( .Z(GFidata[497]));
Q_RDN U47 ( .Z(GFidata[496]));
Q_RDN U48 ( .Z(GFidata[495]));
Q_RDN U49 ( .Z(GFidata[494]));
Q_RDN U50 ( .Z(GFidata[493]));
Q_RDN U51 ( .Z(GFidata[492]));
Q_RDN U52 ( .Z(GFidata[491]));
Q_RDN U53 ( .Z(GFidata[490]));
Q_RDN U54 ( .Z(GFidata[489]));
Q_RDN U55 ( .Z(GFidata[488]));
Q_RDN U56 ( .Z(GFidata[487]));
Q_RDN U57 ( .Z(GFidata[486]));
Q_RDN U58 ( .Z(GFidata[485]));
Q_RDN U59 ( .Z(GFidata[484]));
Q_RDN U60 ( .Z(GFidata[483]));
Q_RDN U61 ( .Z(GFidata[482]));
Q_RDN U62 ( .Z(GFidata[481]));
Q_RDN U63 ( .Z(GFidata[480]));
Q_RDN U64 ( .Z(GFidata[479]));
Q_RDN U65 ( .Z(GFidata[478]));
Q_RDN U66 ( .Z(GFidata[477]));
Q_RDN U67 ( .Z(GFidata[476]));
Q_RDN U68 ( .Z(GFidata[475]));
Q_RDN U69 ( .Z(GFidata[474]));
Q_RDN U70 ( .Z(GFidata[473]));
Q_RDN U71 ( .Z(GFidata[472]));
Q_RDN U72 ( .Z(GFidata[471]));
Q_RDN U73 ( .Z(GFidata[470]));
Q_RDN U74 ( .Z(GFidata[469]));
Q_RDN U75 ( .Z(GFidata[468]));
Q_RDN U76 ( .Z(GFidata[467]));
Q_RDN U77 ( .Z(GFidata[466]));
Q_RDN U78 ( .Z(GFidata[465]));
Q_RDN U79 ( .Z(GFidata[464]));
Q_RDN U80 ( .Z(GFidata[463]));
Q_RDN U81 ( .Z(GFidata[462]));
Q_RDN U82 ( .Z(GFidata[461]));
Q_RDN U83 ( .Z(GFidata[460]));
Q_RDN U84 ( .Z(GFidata[459]));
Q_RDN U85 ( .Z(GFidata[458]));
Q_RDN U86 ( .Z(GFidata[457]));
Q_RDN U87 ( .Z(GFidata[456]));
Q_RDN U88 ( .Z(GFidata[455]));
Q_RDN U89 ( .Z(GFidata[454]));
Q_RDN U90 ( .Z(GFidata[453]));
Q_RDN U91 ( .Z(GFidata[452]));
Q_RDN U92 ( .Z(GFidata[451]));
Q_RDN U93 ( .Z(GFidata[450]));
Q_RDN U94 ( .Z(GFidata[449]));
Q_RDN U95 ( .Z(GFidata[448]));
Q_RDN U96 ( .Z(GFidata[447]));
Q_RDN U97 ( .Z(GFidata[446]));
Q_RDN U98 ( .Z(GFidata[445]));
Q_RDN U99 ( .Z(GFidata[444]));
Q_RDN U100 ( .Z(GFidata[443]));
Q_RDN U101 ( .Z(GFidata[442]));
Q_RDN U102 ( .Z(GFidata[441]));
Q_RDN U103 ( .Z(GFidata[440]));
Q_RDN U104 ( .Z(GFidata[439]));
Q_RDN U105 ( .Z(GFidata[438]));
Q_RDN U106 ( .Z(GFidata[437]));
Q_RDN U107 ( .Z(GFidata[436]));
Q_RDN U108 ( .Z(GFidata[435]));
Q_RDN U109 ( .Z(GFidata[434]));
Q_RDN U110 ( .Z(GFidata[433]));
Q_RDN U111 ( .Z(GFidata[432]));
Q_RDN U112 ( .Z(GFidata[431]));
Q_RDN U113 ( .Z(GFidata[430]));
Q_RDN U114 ( .Z(GFidata[429]));
Q_RDN U115 ( .Z(GFidata[428]));
Q_RDN U116 ( .Z(GFidata[427]));
Q_RDN U117 ( .Z(GFidata[426]));
Q_RDN U118 ( .Z(GFidata[425]));
Q_RDN U119 ( .Z(GFidata[424]));
Q_RDN U120 ( .Z(GFidata[423]));
Q_RDN U121 ( .Z(GFidata[422]));
Q_RDN U122 ( .Z(GFidata[421]));
Q_RDN U123 ( .Z(GFidata[420]));
Q_RDN U124 ( .Z(GFidata[419]));
Q_RDN U125 ( .Z(GFidata[418]));
Q_RDN U126 ( .Z(GFidata[417]));
Q_RDN U127 ( .Z(GFidata[416]));
Q_RDN U128 ( .Z(GFidata[415]));
Q_RDN U129 ( .Z(GFidata[414]));
Q_RDN U130 ( .Z(GFidata[413]));
Q_RDN U131 ( .Z(GFidata[412]));
Q_RDN U132 ( .Z(GFidata[411]));
Q_RDN U133 ( .Z(GFidata[410]));
Q_RDN U134 ( .Z(GFidata[409]));
Q_RDN U135 ( .Z(GFidata[408]));
Q_RDN U136 ( .Z(GFidata[407]));
Q_RDN U137 ( .Z(GFidata[406]));
Q_RDN U138 ( .Z(GFidata[405]));
Q_RDN U139 ( .Z(GFidata[404]));
Q_RDN U140 ( .Z(GFidata[403]));
Q_RDN U141 ( .Z(GFidata[402]));
Q_RDN U142 ( .Z(GFidata[401]));
Q_RDN U143 ( .Z(GFidata[400]));
Q_RDN U144 ( .Z(GFidata[399]));
Q_RDN U145 ( .Z(GFidata[398]));
Q_RDN U146 ( .Z(GFidata[397]));
Q_RDN U147 ( .Z(GFidata[396]));
Q_RDN U148 ( .Z(GFidata[395]));
Q_RDN U149 ( .Z(GFidata[394]));
Q_RDN U150 ( .Z(GFidata[393]));
Q_RDN U151 ( .Z(GFidata[392]));
Q_RDN U152 ( .Z(GFidata[391]));
Q_RDN U153 ( .Z(GFidata[390]));
Q_RDN U154 ( .Z(GFidata[389]));
Q_RDN U155 ( .Z(GFidata[388]));
Q_RDN U156 ( .Z(GFidata[387]));
Q_RDN U157 ( .Z(GFidata[386]));
Q_RDN U158 ( .Z(GFidata[385]));
Q_RDN U159 ( .Z(GFidata[384]));
Q_RDN U160 ( .Z(GFidata[383]));
Q_RDN U161 ( .Z(GFidata[382]));
Q_RDN U162 ( .Z(GFidata[381]));
Q_RDN U163 ( .Z(GFidata[380]));
Q_RDN U164 ( .Z(GFidata[379]));
Q_RDN U165 ( .Z(GFidata[378]));
Q_RDN U166 ( .Z(GFidata[377]));
Q_RDN U167 ( .Z(GFidata[376]));
Q_RDN U168 ( .Z(GFidata[375]));
Q_RDN U169 ( .Z(GFidata[374]));
Q_RDN U170 ( .Z(GFidata[373]));
Q_RDN U171 ( .Z(GFidata[372]));
Q_RDN U172 ( .Z(GFidata[371]));
Q_RDN U173 ( .Z(GFidata[370]));
Q_RDN U174 ( .Z(GFidata[369]));
Q_RDN U175 ( .Z(GFidata[368]));
Q_RDN U176 ( .Z(GFidata[367]));
Q_RDN U177 ( .Z(GFidata[366]));
Q_RDN U178 ( .Z(GFidata[365]));
Q_RDN U179 ( .Z(GFidata[364]));
Q_RDN U180 ( .Z(GFidata[363]));
Q_RDN U181 ( .Z(GFidata[362]));
Q_RDN U182 ( .Z(GFidata[361]));
Q_RDN U183 ( .Z(GFidata[360]));
Q_RDN U184 ( .Z(GFidata[359]));
Q_RDN U185 ( .Z(GFidata[358]));
Q_RDN U186 ( .Z(GFidata[357]));
Q_RDN U187 ( .Z(GFidata[356]));
Q_RDN U188 ( .Z(GFidata[355]));
Q_RDN U189 ( .Z(GFidata[354]));
Q_RDN U190 ( .Z(GFidata[353]));
Q_RDN U191 ( .Z(GFidata[352]));
Q_RDN U192 ( .Z(GFidata[351]));
Q_RDN U193 ( .Z(GFidata[350]));
Q_RDN U194 ( .Z(GFidata[349]));
Q_RDN U195 ( .Z(GFidata[348]));
Q_RDN U196 ( .Z(GFidata[347]));
Q_RDN U197 ( .Z(GFidata[346]));
Q_RDN U198 ( .Z(GFidata[345]));
Q_RDN U199 ( .Z(GFidata[344]));
Q_RDN U200 ( .Z(GFidata[343]));
Q_RDN U201 ( .Z(GFidata[342]));
Q_RDN U202 ( .Z(GFidata[341]));
Q_RDN U203 ( .Z(GFidata[340]));
Q_RDN U204 ( .Z(GFidata[339]));
Q_RDN U205 ( .Z(GFidata[338]));
Q_RDN U206 ( .Z(GFidata[337]));
Q_RDN U207 ( .Z(GFidata[336]));
Q_RDN U208 ( .Z(GFidata[335]));
Q_RDN U209 ( .Z(GFidata[334]));
Q_RDN U210 ( .Z(GFidata[333]));
Q_RDN U211 ( .Z(GFidata[332]));
Q_RDN U212 ( .Z(GFidata[331]));
Q_RDN U213 ( .Z(GFidata[330]));
Q_RDN U214 ( .Z(GFidata[329]));
Q_RDN U215 ( .Z(GFidata[328]));
Q_RDN U216 ( .Z(GFidata[327]));
Q_RDN U217 ( .Z(GFidata[326]));
Q_RDN U218 ( .Z(GFidata[325]));
Q_RDN U219 ( .Z(GFidata[324]));
Q_RDN U220 ( .Z(GFidata[323]));
Q_RDN U221 ( .Z(GFidata[322]));
Q_RDN U222 ( .Z(GFidata[321]));
Q_RDN U223 ( .Z(GFidata[320]));
Q_RDN U224 ( .Z(GFidata[319]));
Q_RDN U225 ( .Z(GFidata[318]));
Q_RDN U226 ( .Z(GFidata[317]));
Q_RDN U227 ( .Z(GFidata[316]));
Q_RDN U228 ( .Z(GFidata[315]));
Q_RDN U229 ( .Z(GFidata[314]));
Q_RDN U230 ( .Z(GFidata[313]));
Q_RDN U231 ( .Z(GFidata[312]));
Q_RDN U232 ( .Z(GFidata[311]));
Q_RDN U233 ( .Z(GFidata[310]));
Q_RDN U234 ( .Z(GFidata[309]));
Q_RDN U235 ( .Z(GFidata[308]));
Q_RDN U236 ( .Z(GFidata[307]));
Q_RDN U237 ( .Z(GFidata[306]));
Q_RDN U238 ( .Z(GFidata[305]));
Q_RDN U239 ( .Z(GFidata[304]));
Q_RDN U240 ( .Z(GFidata[303]));
Q_RDN U241 ( .Z(GFidata[302]));
Q_RDN U242 ( .Z(GFidata[301]));
Q_RDN U243 ( .Z(GFidata[300]));
Q_RDN U244 ( .Z(GFidata[299]));
Q_RDN U245 ( .Z(GFidata[298]));
Q_RDN U246 ( .Z(GFidata[297]));
Q_RDN U247 ( .Z(GFidata[296]));
Q_RDN U248 ( .Z(GFidata[295]));
Q_RDN U249 ( .Z(GFidata[294]));
Q_RDN U250 ( .Z(GFidata[293]));
Q_RDN U251 ( .Z(GFidata[292]));
Q_RDN U252 ( .Z(GFidata[291]));
Q_RDN U253 ( .Z(GFidata[290]));
Q_RDN U254 ( .Z(GFidata[289]));
Q_RDN U255 ( .Z(GFidata[288]));
Q_RDN U256 ( .Z(GFidata[287]));
Q_RDN U257 ( .Z(GFidata[286]));
Q_RDN U258 ( .Z(GFidata[285]));
Q_RDN U259 ( .Z(GFidata[284]));
Q_RDN U260 ( .Z(GFidata[283]));
Q_RDN U261 ( .Z(GFidata[282]));
Q_RDN U262 ( .Z(GFidata[281]));
Q_RDN U263 ( .Z(GFidata[280]));
Q_RDN U264 ( .Z(GFidata[279]));
Q_RDN U265 ( .Z(GFidata[278]));
Q_RDN U266 ( .Z(GFidata[277]));
Q_RDN U267 ( .Z(GFidata[276]));
Q_RDN U268 ( .Z(GFidata[275]));
Q_RDN U269 ( .Z(GFidata[274]));
Q_RDN U270 ( .Z(GFidata[273]));
Q_RDN U271 ( .Z(GFidata[272]));
Q_RDN U272 ( .Z(GFidata[271]));
Q_RDN U273 ( .Z(GFidata[270]));
Q_RDN U274 ( .Z(GFidata[269]));
Q_RDN U275 ( .Z(GFidata[268]));
Q_RDN U276 ( .Z(GFidata[267]));
Q_RDN U277 ( .Z(GFidata[266]));
Q_RDN U278 ( .Z(GFidata[265]));
Q_RDN U279 ( .Z(GFidata[264]));
Q_RDN U280 ( .Z(GFidata[263]));
Q_RDN U281 ( .Z(GFidata[262]));
Q_RDN U282 ( .Z(GFidata[261]));
Q_RDN U283 ( .Z(GFidata[260]));
Q_RDN U284 ( .Z(GFidata[259]));
Q_RDN U285 ( .Z(GFidata[258]));
Q_RDN U286 ( .Z(GFidata[257]));
Q_RDN U287 ( .Z(GFidata[256]));
Q_RDN U288 ( .Z(GFidata[255]));
Q_RDN U289 ( .Z(GFidata[254]));
Q_RDN U290 ( .Z(GFidata[253]));
Q_RDN U291 ( .Z(GFidata[252]));
Q_RDN U292 ( .Z(GFidata[251]));
Q_RDN U293 ( .Z(GFidata[250]));
Q_RDN U294 ( .Z(GFidata[249]));
Q_RDN U295 ( .Z(GFidata[248]));
Q_RDN U296 ( .Z(GFidata[247]));
Q_RDN U297 ( .Z(GFidata[246]));
Q_RDN U298 ( .Z(GFidata[245]));
Q_RDN U299 ( .Z(GFidata[244]));
Q_RDN U300 ( .Z(GFidata[243]));
Q_RDN U301 ( .Z(GFidata[242]));
Q_RDN U302 ( .Z(GFidata[241]));
Q_RDN U303 ( .Z(GFidata[240]));
Q_RDN U304 ( .Z(GFidata[239]));
Q_RDN U305 ( .Z(GFidata[238]));
Q_RDN U306 ( .Z(GFidata[237]));
Q_RDN U307 ( .Z(GFidata[236]));
Q_RDN U308 ( .Z(GFidata[235]));
Q_RDN U309 ( .Z(GFidata[234]));
Q_RDN U310 ( .Z(GFidata[233]));
Q_RDN U311 ( .Z(GFidata[232]));
Q_RDN U312 ( .Z(GFidata[231]));
Q_RDN U313 ( .Z(GFidata[230]));
Q_RDN U314 ( .Z(GFidata[229]));
Q_RDN U315 ( .Z(GFidata[228]));
Q_RDN U316 ( .Z(GFidata[227]));
Q_RDN U317 ( .Z(GFidata[226]));
Q_RDN U318 ( .Z(GFidata[225]));
Q_RDN U319 ( .Z(GFidata[224]));
Q_RDN U320 ( .Z(GFidata[223]));
Q_RDN U321 ( .Z(GFidata[222]));
Q_RDN U322 ( .Z(GFidata[221]));
Q_RDN U323 ( .Z(GFidata[220]));
Q_RDN U324 ( .Z(GFidata[219]));
Q_RDN U325 ( .Z(GFidata[218]));
Q_RDN U326 ( .Z(GFidata[217]));
Q_RDN U327 ( .Z(GFidata[216]));
Q_RDN U328 ( .Z(GFidata[215]));
Q_RDN U329 ( .Z(GFidata[214]));
Q_RDN U330 ( .Z(GFidata[213]));
Q_RDN U331 ( .Z(GFidata[212]));
Q_RDN U332 ( .Z(GFidata[211]));
Q_RDN U333 ( .Z(GFidata[210]));
Q_RDN U334 ( .Z(GFidata[209]));
Q_RDN U335 ( .Z(GFidata[208]));
Q_RDN U336 ( .Z(GFidata[207]));
Q_RDN U337 ( .Z(GFidata[206]));
Q_RDN U338 ( .Z(GFidata[205]));
Q_RDN U339 ( .Z(GFidata[204]));
Q_RDN U340 ( .Z(GFidata[203]));
Q_RDN U341 ( .Z(GFidata[202]));
Q_RDN U342 ( .Z(GFidata[201]));
Q_RDN U343 ( .Z(GFidata[200]));
Q_RDN U344 ( .Z(GFidata[199]));
Q_RDN U345 ( .Z(GFidata[198]));
Q_RDN U346 ( .Z(GFidata[197]));
Q_RDN U347 ( .Z(GFidata[196]));
Q_RDN U348 ( .Z(GFidata[195]));
Q_RDN U349 ( .Z(GFidata[194]));
Q_RDN U350 ( .Z(GFidata[193]));
Q_RDN U351 ( .Z(GFidata[192]));
Q_RDN U352 ( .Z(GFidata[191]));
Q_RDN U353 ( .Z(GFidata[190]));
Q_RDN U354 ( .Z(GFidata[189]));
Q_RDN U355 ( .Z(GFidata[188]));
Q_RDN U356 ( .Z(GFidata[187]));
Q_RDN U357 ( .Z(GFidata[186]));
Q_RDN U358 ( .Z(GFidata[185]));
Q_RDN U359 ( .Z(GFidata[184]));
Q_RDN U360 ( .Z(GFidata[183]));
Q_RDN U361 ( .Z(GFidata[182]));
Q_RDN U362 ( .Z(GFidata[181]));
Q_RDN U363 ( .Z(GFidata[180]));
Q_RDN U364 ( .Z(GFidata[179]));
Q_RDN U365 ( .Z(GFidata[178]));
Q_RDN U366 ( .Z(GFidata[177]));
Q_RDN U367 ( .Z(GFidata[176]));
Q_RDN U368 ( .Z(GFidata[175]));
Q_RDN U369 ( .Z(GFidata[174]));
Q_RDN U370 ( .Z(GFidata[173]));
Q_RDN U371 ( .Z(GFidata[172]));
Q_RDN U372 ( .Z(GFidata[171]));
Q_RDN U373 ( .Z(GFidata[170]));
Q_RDN U374 ( .Z(GFidata[169]));
Q_RDN U375 ( .Z(GFidata[168]));
Q_RDN U376 ( .Z(GFidata[167]));
Q_RDN U377 ( .Z(GFidata[166]));
Q_RDN U378 ( .Z(GFidata[165]));
Q_RDN U379 ( .Z(GFidata[164]));
Q_RDN U380 ( .Z(GFidata[163]));
Q_RDN U381 ( .Z(GFidata[162]));
Q_RDN U382 ( .Z(GFidata[161]));
Q_RDN U383 ( .Z(GFidata[160]));
Q_RDN U384 ( .Z(GFidata[159]));
Q_RDN U385 ( .Z(GFidata[158]));
Q_RDN U386 ( .Z(GFidata[157]));
Q_RDN U387 ( .Z(GFidata[156]));
Q_RDN U388 ( .Z(GFidata[155]));
Q_RDN U389 ( .Z(GFidata[154]));
Q_RDN U390 ( .Z(GFidata[153]));
Q_RDN U391 ( .Z(GFidata[152]));
Q_RDN U392 ( .Z(GFidata[151]));
Q_RDN U393 ( .Z(GFidata[150]));
Q_RDN U394 ( .Z(GFidata[149]));
Q_RDN U395 ( .Z(GFidata[148]));
Q_RDN U396 ( .Z(GFidata[147]));
Q_RDN U397 ( .Z(GFidata[146]));
Q_RDN U398 ( .Z(GFidata[145]));
Q_RDN U399 ( .Z(GFidata[144]));
Q_RDN U400 ( .Z(GFidata[143]));
Q_RDN U401 ( .Z(GFidata[142]));
Q_RDN U402 ( .Z(GFidata[141]));
Q_RDN U403 ( .Z(GFidata[140]));
Q_RDN U404 ( .Z(GFidata[139]));
Q_RDN U405 ( .Z(GFidata[138]));
Q_RDN U406 ( .Z(GFidata[137]));
Q_RDN U407 ( .Z(GFidata[136]));
Q_RDN U408 ( .Z(GFidata[135]));
Q_RDN U409 ( .Z(GFidata[134]));
Q_RDN U410 ( .Z(GFidata[133]));
Q_RDN U411 ( .Z(GFidata[132]));
Q_RDN U412 ( .Z(GFidata[131]));
Q_RDN U413 ( .Z(GFidata[130]));
Q_RDN U414 ( .Z(GFidata[129]));
Q_RDN U415 ( .Z(GFidata[128]));
Q_RDN U416 ( .Z(GFidata[127]));
Q_RDN U417 ( .Z(GFidata[126]));
Q_RDN U418 ( .Z(GFidata[125]));
Q_RDN U419 ( .Z(GFidata[124]));
Q_RDN U420 ( .Z(GFidata[123]));
Q_RDN U421 ( .Z(GFidata[122]));
Q_RDN U422 ( .Z(GFidata[121]));
Q_RDN U423 ( .Z(GFidata[120]));
Q_RDN U424 ( .Z(GFidata[119]));
Q_RDN U425 ( .Z(GFidata[118]));
Q_RDN U426 ( .Z(GFidata[117]));
Q_RDN U427 ( .Z(GFidata[116]));
Q_RDN U428 ( .Z(GFidata[115]));
Q_RDN U429 ( .Z(GFidata[114]));
Q_RDN U430 ( .Z(GFidata[113]));
Q_RDN U431 ( .Z(GFidata[112]));
Q_RDN U432 ( .Z(GFidata[111]));
Q_RDN U433 ( .Z(GFidata[110]));
Q_RDN U434 ( .Z(GFidata[109]));
Q_RDN U435 ( .Z(GFidata[108]));
Q_RDN U436 ( .Z(GFidata[107]));
Q_RDN U437 ( .Z(GFidata[106]));
Q_RDN U438 ( .Z(GFidata[105]));
Q_RDN U439 ( .Z(GFidata[104]));
Q_RDN U440 ( .Z(GFidata[103]));
Q_RDN U441 ( .Z(GFidata[102]));
Q_RDN U442 ( .Z(GFidata[101]));
Q_RDN U443 ( .Z(GFidata[100]));
Q_RDN U444 ( .Z(GFidata[99]));
Q_RDN U445 ( .Z(GFidata[98]));
Q_RDN U446 ( .Z(GFidata[97]));
Q_RDN U447 ( .Z(GFidata[96]));
Q_RDN U448 ( .Z(GFidata[95]));
Q_RDN U449 ( .Z(GFidata[94]));
Q_RDN U450 ( .Z(GFidata[93]));
Q_RDN U451 ( .Z(GFidata[92]));
Q_RDN U452 ( .Z(GFidata[91]));
Q_RDN U453 ( .Z(GFidata[90]));
Q_RDN U454 ( .Z(GFidata[89]));
Q_RDN U455 ( .Z(GFidata[88]));
Q_RDN U456 ( .Z(GFidata[87]));
Q_RDN U457 ( .Z(GFidata[86]));
Q_RDN U458 ( .Z(GFidata[85]));
Q_RDN U459 ( .Z(GFidata[84]));
Q_RDN U460 ( .Z(GFidata[83]));
Q_RDN U461 ( .Z(GFidata[82]));
Q_RDN U462 ( .Z(GFidata[81]));
Q_RDN U463 ( .Z(GFidata[80]));
Q_RDN U464 ( .Z(GFidata[79]));
Q_RDN U465 ( .Z(GFidata[78]));
Q_RDN U466 ( .Z(GFidata[77]));
Q_RDN U467 ( .Z(GFidata[76]));
Q_RDN U468 ( .Z(GFidata[75]));
Q_RDN U469 ( .Z(GFidata[74]));
Q_RDN U470 ( .Z(GFidata[73]));
Q_RDN U471 ( .Z(GFidata[72]));
Q_RDN U472 ( .Z(GFidata[71]));
Q_RDN U473 ( .Z(GFidata[70]));
Q_RDN U474 ( .Z(GFidata[69]));
Q_RDN U475 ( .Z(GFidata[68]));
Q_RDN U476 ( .Z(GFidata[67]));
Q_RDN U477 ( .Z(GFidata[66]));
Q_RDN U478 ( .Z(GFidata[65]));
Q_RDN U479 ( .Z(GFidata[64]));
Q_RDN U480 ( .Z(GFidata[63]));
Q_RDN U481 ( .Z(GFidata[62]));
Q_RDN U482 ( .Z(GFidata[61]));
Q_RDN U483 ( .Z(GFidata[60]));
Q_RDN U484 ( .Z(GFidata[59]));
Q_RDN U485 ( .Z(GFidata[58]));
Q_RDN U486 ( .Z(GFidata[57]));
Q_RDN U487 ( .Z(GFidata[56]));
Q_RDN U488 ( .Z(GFidata[55]));
Q_RDN U489 ( .Z(GFidata[54]));
Q_RDN U490 ( .Z(GFidata[53]));
Q_RDN U491 ( .Z(GFidata[52]));
Q_RDN U492 ( .Z(GFidata[51]));
Q_RDN U493 ( .Z(GFidata[50]));
Q_RDN U494 ( .Z(GFidata[49]));
Q_RDN U495 ( .Z(GFidata[48]));
Q_RDN U496 ( .Z(GFidata[47]));
Q_RDN U497 ( .Z(GFidata[46]));
Q_RDN U498 ( .Z(GFidata[45]));
Q_RDN U499 ( .Z(GFidata[44]));
Q_RDN U500 ( .Z(GFidata[43]));
Q_RDN U501 ( .Z(GFidata[42]));
Q_RDN U502 ( .Z(GFidata[41]));
Q_RDN U503 ( .Z(GFidata[40]));
Q_RDN U504 ( .Z(GFidata[39]));
Q_RDN U505 ( .Z(GFidata[38]));
Q_RDN U506 ( .Z(GFidata[37]));
Q_RDN U507 ( .Z(GFidata[36]));
Q_RDN U508 ( .Z(GFidata[35]));
Q_RDN U509 ( .Z(GFidata[34]));
Q_RDN U510 ( .Z(GFidata[33]));
Q_RDN U511 ( .Z(GFidata[32]));
Q_RDN U512 ( .Z(GFidata[31]));
Q_RDN U513 ( .Z(GFidata[30]));
Q_RDN U514 ( .Z(GFidata[29]));
Q_RDN U515 ( .Z(GFidata[28]));
Q_RDN U516 ( .Z(GFidata[27]));
Q_RDN U517 ( .Z(GFidata[26]));
Q_RDN U518 ( .Z(GFidata[25]));
Q_RDN U519 ( .Z(GFidata[24]));
Q_RDN U520 ( .Z(GFidata[23]));
Q_RDN U521 ( .Z(GFidata[22]));
Q_RDN U522 ( .Z(GFidata[21]));
Q_RDN U523 ( .Z(GFidata[20]));
Q_RDN U524 ( .Z(GFidata[19]));
Q_RDN U525 ( .Z(GFidata[18]));
Q_RDN U526 ( .Z(GFidata[17]));
Q_RDN U527 ( .Z(GFidata[16]));
Q_RDN U528 ( .Z(GFidata[15]));
Q_RDN U529 ( .Z(GFidata[14]));
Q_RDN U530 ( .Z(GFidata[13]));
Q_RDN U531 ( .Z(GFidata[12]));
Q_RDN U532 ( .Z(GFidata[11]));
Q_RDN U533 ( .Z(GFidata[10]));
Q_RDN U534 ( .Z(GFidata[9]));
Q_RDN U535 ( .Z(GFidata[8]));
Q_RDN U536 ( .Z(GFidata[7]));
Q_RDN U537 ( .Z(GFidata[6]));
Q_RDN U538 ( .Z(GFidata[5]));
Q_RDN U539 ( .Z(GFidata[4]));
Q_RDN U540 ( .Z(GFidata[3]));
Q_RDN U541 ( .Z(GFidata[2]));
Q_RDN U542 ( .Z(GFidata[1]));
Q_RDN U543 ( .Z(GFidata[0]));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_RDN U545 ( .Z(GFtsReq));
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
