
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_xcm117 ( clk, rst_n, wr_stb, reg_addr, cmnd_op, 
	cmnd_addr, cmnd_table_id, stat_code, stat_datawords, stat_addr, 
	stat_table_id, capability_lst, capability_type, enable, .addr_limit( {
	\addr_limit[0][8] , \addr_limit[0][7] , \addr_limit[0][6] , 
	\addr_limit[0][5] , \addr_limit[0][4] , \addr_limit[0][3] , 
	\addr_limit[0][2] , \addr_limit[0][1] , \addr_limit[0][0] } ), 
	wr_dat, rd_dat, sw_cs, sw_ce, sw_we, sw_add, sw_wdat, sw_rdat, 
	sw_match, sw_aindex, grant, yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [8:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [8:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][8] ;
input \addr_limit[0][7] ;
input \addr_limit[0][6] ;
input \addr_limit[0][5] ;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [95:0] wr_dat;
output [95:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [8:0] sw_add;
output [95:0] sw_wdat;
input [95:0] sw_rdat;
input sw_match;
input [7:0] sw_aindex;
input grant;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:8] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:95] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:8] _zy_simnet_sw_add_11_w$;
wire [0:95] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [8:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [5:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [8:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(n1), .Z(stat_datawords[0]));
Q_BUF U1 ( .A(n2), .Z(stat_datawords[1]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U5 ( .A(n1), .Z(capability_type[0]));
Q_BUF U6 ( .A(n1), .Z(capability_type[1]));
Q_BUF U7 ( .A(n1), .Z(capability_type[2]));
Q_BUF U8 ( .A(n1), .Z(capability_type[3]));
Q_BUF U9 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[2]));
Q_BUF U12 ( .A(n2), .Z(capability_lst[3]));
Q_BUF U13 ( .A(n2), .Z(capability_lst[4]));
Q_BUF U14 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[6]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U17 ( .A(n2), .Z(capability_lst[8]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U23 ( .A(n2), .Z(capability_lst[14]));
Q_BUF U24 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U25 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_or_ini_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_96 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:95], sw_wdat[95:0]);
ixc_assign_9 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:8], sw_add[8:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_96 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:95], rd_dat[95:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n1, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n2, 
	n1, n1, n1, n1, n1, n2, n1, n2, n2, n2, n2, n2, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_9 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:8], stat_addr[8:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n2, n1});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_9 _zz_strnp_6 ( stat_addr[8:0], maxaddr[8:0]);
Q_AN02 U46 ( .A0(n36), .A1(grant), .Z(igrant));
Q_AN02 U47 ( .A0(cmnd_issued), .A1(n35), .Z(badaddr));
Q_OR03 U48 ( .A0(n16), .A1(n34), .A2(n33), .Z(n35));
Q_AN02 U49 ( .A0(n17), .A1(n29), .Z(n34));
Q_AN02 U50 ( .A0(n17), .A1(n30), .Z(n32));
Q_AN03 U51 ( .A0(cmnd_addr[0]), .A1(n31), .A2(n32), .Z(n33));
Q_INV U52 ( .A(maxaddr[0]), .Z(n31));
Q_OR03 U53 ( .A0(n26), .A1(n25), .A2(n28), .Z(n29));
Q_OA21 U54 ( .A0(cmnd_addr[1]), .A1(n22), .B0(n24), .Z(n30));
Q_AN03 U55 ( .A0(cmnd_addr[1]), .A1(n22), .A2(n24), .Z(n25));
Q_INV U56 ( .A(maxaddr[1]), .Z(n22));
Q_OA21 U57 ( .A0(cmnd_addr[2]), .A1(n21), .B0(n23), .Z(n24));
Q_AN03 U58 ( .A0(cmnd_addr[2]), .A1(n21), .A2(n23), .Z(n26));
Q_INV U59 ( .A(maxaddr[2]), .Z(n21));
Q_OA21 U60 ( .A0(cmnd_addr[3]), .A1(n20), .B0(n19), .Z(n23));
Q_AN03 U61 ( .A0(cmnd_addr[3]), .A1(n20), .A2(n19), .Z(n27));
Q_INV U62 ( .A(maxaddr[3]), .Z(n20));
Q_OR02 U63 ( .A0(cmnd_addr[4]), .A1(n18), .Z(n19));
Q_AO21 U64 ( .A0(cmnd_addr[4]), .A1(n18), .B0(n27), .Z(n28));
Q_INV U65 ( .A(maxaddr[4]), .Z(n18));
Q_OR03 U66 ( .A0(n13), .A1(n12), .A2(n15), .Z(n16));
Q_OA21 U67 ( .A0(cmnd_addr[5]), .A1(n9), .B0(n11), .Z(n17));
Q_AN03 U68 ( .A0(cmnd_addr[5]), .A1(n9), .A2(n11), .Z(n12));
Q_INV U69 ( .A(maxaddr[5]), .Z(n9));
Q_OA21 U70 ( .A0(cmnd_addr[6]), .A1(n8), .B0(n10), .Z(n11));
Q_AN03 U71 ( .A0(cmnd_addr[6]), .A1(n8), .A2(n10), .Z(n13));
Q_INV U72 ( .A(maxaddr[6]), .Z(n8));
Q_OA21 U73 ( .A0(cmnd_addr[7]), .A1(n7), .B0(n6), .Z(n10));
Q_AN03 U74 ( .A0(cmnd_addr[7]), .A1(n7), .A2(n6), .Z(n14));
Q_INV U75 ( .A(maxaddr[7]), .Z(n7));
Q_OR02 U76 ( .A0(cmnd_addr[8]), .A1(n5), .Z(n6));
Q_AO21 U77 ( .A0(cmnd_addr[8]), .A1(n5), .B0(n14), .Z(n15));
Q_INV U78 ( .A(maxaddr[8]), .Z(n5));
Q_AN02 U79 ( .A0(n3), .A1(n4), .Z(timeout));
Q_AN03 U80 ( .A0(timer_r[2]), .A1(timer_r[1]), .A2(timer_r[0]), .Z(n4));
Q_AN03 U81 ( .A0(timer_r[5]), .A1(timer_r[4]), .A2(timer_r[3]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timer_r[5]);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U86 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U87 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U88 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U89 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U90 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_MX02 U91 ( .S(rst_or_ini_r), .A0(cmnd_addr[5]), .A1(rst_addr_r[5]), .Z(sw_add[5]));
Q_MX02 U92 ( .S(rst_or_ini_r), .A0(cmnd_addr[6]), .A1(rst_addr_r[6]), .Z(sw_add[6]));
Q_MX02 U93 ( .S(rst_or_ini_r), .A0(cmnd_addr[7]), .A1(rst_addr_r[7]), .Z(sw_add[7]));
Q_MX02 U94 ( .S(rst_or_ini_r), .A0(cmnd_addr[8]), .A1(rst_addr_r[8]), .Z(sw_add[8]));
Q_AN02 U95 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U96 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U97 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U98 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U99 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_AN02 U100 ( .A0(enable), .A1(\addr_limit[0][5] ), .Z(maxaddr[5]));
Q_AN02 U101 ( .A0(enable), .A1(\addr_limit[0][6] ), .Z(maxaddr[6]));
Q_AN02 U102 ( .A0(enable), .A1(\addr_limit[0][7] ), .Z(maxaddr[7]));
Q_AN02 U103 ( .A0(enable), .A1(\addr_limit[0][8] ), .Z(maxaddr[8]));
Q_OR03 U104 ( .A0(reg_addr[10]), .A1(reg_addr[9]), .A2(reg_addr[8]), .Z(n37));
Q_ND03 U105 ( .A0(reg_addr[7]), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n38));
Q_OR03 U106 ( .A0(reg_addr[4]), .A1(reg_addr[3]), .A2(reg_addr[2]), .Z(n39));
Q_OR03 U107 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n37), .Z(n40));
Q_NR03 U108 ( .A0(n38), .A1(n39), .A2(n40), .Z(n41));
Q_AN02 U109 ( .A0(wr_stb), .A1(n41), .Z(n65));
Q_INV U110 ( .A(n60), .Z(cmnd_issued));
Q_INV U111 ( .A(unsupported_op), .Z(n59));
Q_OA21 U112 ( .A0(n43), .A1(n44), .B0(n42), .Z(unsupported_op));
Q_AN02 U113 ( .A0(n42), .A1(n45), .Z(ack_error));
Q_AO21 U114 ( .A0(n47), .A1(n48), .B0(n46), .Z(n60));
Q_INV U115 ( .A(n65), .Z(n46));
Q_MX02 U116 ( .S(cmnd[3]), .A0(n51), .A1(n49), .Z(n47));
Q_INV U117 ( .A(cmnd_cmp_stb), .Z(n61));
Q_AN02 U118 ( .A0(n42), .A1(n52), .Z(cmnd_cmp_stb));
Q_AN02 U119 ( .A0(n42), .A1(n53), .Z(cmnd_tmo_stb));
Q_AN03 U120 ( .A0(n42), .A1(n48), .A2(n51), .Z(cmnd_sis_stb));
Q_AN02 U121 ( .A0(n65), .A1(cmnd[3]), .Z(n42));
Q_AN02 U122 ( .A0(n54), .A1(n45), .Z(cmnd_inc_stb));
Q_AN02 U123 ( .A0(n49), .A1(cmnd[0]), .Z(n45));
Q_AN02 U124 ( .A0(n54), .A1(n53), .Z(cmnd_ini_stb));
Q_AN02 U125 ( .A0(n49), .A1(n48), .Z(n53));
Q_AN02 U126 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n49));
Q_INV U127 ( .A(cmnd_rst_stb), .Z(n62));
Q_AN02 U128 ( .A0(n44), .A1(n55), .Z(cmnd_rst_stb));
Q_AN02 U129 ( .A0(n54), .A1(cmnd[0]), .Z(n55));
Q_AN02 U130 ( .A0(n44), .A1(n56), .Z(cmnd_dis_stb));
Q_AN02 U131 ( .A0(n54), .A1(n48), .Z(n56));
Q_AN02 U132 ( .A0(cmnd[2]), .A1(n57), .Z(n44));
Q_AN02 U133 ( .A0(n43), .A1(n55), .Z(cmnd_ena_stb));
Q_INV U134 ( .A(cmnd_wr_stb), .Z(n63));
Q_AN02 U135 ( .A0(n43), .A1(n56), .Z(cmnd_wr_stb));
Q_INV U136 ( .A(cmnd[0]), .Z(n48));
Q_AN02 U137 ( .A0(n58), .A1(cmnd[1]), .Z(n43));
Q_INV U138 ( .A(cmnd_rd_stb), .Z(n64));
Q_AN02 U139 ( .A0(n54), .A1(n52), .Z(cmnd_rd_stb));
Q_AN02 U140 ( .A0(n51), .A1(cmnd[0]), .Z(n52));
Q_NR02 U141 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n51));
Q_INV U142 ( .A(cmnd[1]), .Z(n57));
Q_INV U143 ( .A(cmnd[2]), .Z(n58));
Q_AN02 U144 ( .A0(n65), .A1(n50), .Z(n54));
Q_INV U145 ( .A(cmnd[3]), .Z(n50));
Q_OR02 U146 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n513));
Q_XNR2 U147 ( .A0(rst_addr_r[0]), .A1(maxaddr[0]), .Z(n66));
Q_XNR2 U148 ( .A0(rst_addr_r[1]), .A1(maxaddr[1]), .Z(n67));
Q_XNR2 U149 ( .A0(rst_addr_r[2]), .A1(maxaddr[2]), .Z(n68));
Q_XNR2 U150 ( .A0(rst_addr_r[3]), .A1(maxaddr[3]), .Z(n69));
Q_XNR2 U151 ( .A0(rst_addr_r[4]), .A1(maxaddr[4]), .Z(n70));
Q_XNR2 U152 ( .A0(rst_addr_r[5]), .A1(maxaddr[5]), .Z(n71));
Q_XNR2 U153 ( .A0(rst_addr_r[6]), .A1(maxaddr[6]), .Z(n72));
Q_XNR2 U154 ( .A0(rst_addr_r[7]), .A1(maxaddr[7]), .Z(n73));
Q_XNR2 U155 ( .A0(rst_addr_r[8]), .A1(maxaddr[8]), .Z(n74));
Q_AN03 U156 ( .A0(n74), .A1(n73), .A2(n72), .Z(n75));
Q_AN03 U157 ( .A0(n71), .A1(n70), .A2(n69), .Z(n76));
Q_AN03 U158 ( .A0(n68), .A1(n67), .A2(n66), .Z(n77));
Q_AN03 U159 ( .A0(n75), .A1(n76), .A2(n77), .Z(n514));
Q_XNR2 U160 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n78));
Q_XNR2 U161 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n79));
Q_XNR2 U162 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n80));
Q_XNR2 U163 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n81));
Q_XNR2 U164 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n82));
Q_XNR2 U165 ( .A0(rst_addr_r[5]), .A1(cmnd_addr[5]), .Z(n83));
Q_XNR2 U166 ( .A0(rst_addr_r[6]), .A1(cmnd_addr[6]), .Z(n84));
Q_XNR2 U167 ( .A0(rst_addr_r[7]), .A1(cmnd_addr[7]), .Z(n85));
Q_XNR2 U168 ( .A0(rst_addr_r[8]), .A1(cmnd_addr[8]), .Z(n86));
Q_AN03 U169 ( .A0(n86), .A1(n85), .A2(n84), .Z(n87));
Q_AN03 U170 ( .A0(n83), .A1(n82), .A2(n81), .Z(n88));
Q_AN03 U171 ( .A0(n80), .A1(n79), .A2(n78), .Z(n89));
Q_AN03 U172 ( .A0(n87), .A1(n88), .A2(n89), .Z(n515));
Q_AN02 U173 ( .A0(init_inc_r), .A1(igrant), .Z(n90));
Q_XOR2 U174 ( .A0(inc_r[0]), .A1(n90), .Z(n91));
Q_AD01HF U175 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n92), .CO(n93));
Q_AD01HF U176 ( .A0(rst_addr_r[1]), .B0(n93), .S(n94), .CO(n95));
Q_AD01HF U177 ( .A0(rst_addr_r[2]), .B0(n95), .S(n96), .CO(n97));
Q_AD01HF U178 ( .A0(rst_addr_r[3]), .B0(n97), .S(n98), .CO(n99));
Q_AD01HF U179 ( .A0(rst_addr_r[4]), .B0(n99), .S(n100), .CO(n101));
Q_AD01HF U180 ( .A0(rst_addr_r[5]), .B0(n101), .S(n102), .CO(n103));
Q_AD01HF U181 ( .A0(rst_addr_r[6]), .B0(n103), .S(n104), .CO(n105));
Q_AD01HF U182 ( .A0(rst_addr_r[7]), .B0(n105), .S(n106), .CO(n107));
Q_XOR2 U183 ( .A0(rst_addr_r[8]), .A1(n107), .Z(n108));
Q_AD01HF U184 ( .A0(timer_r[1]), .B0(timer_r[0]), .S(n110), .CO(n111));
Q_AD01HF U185 ( .A0(timer_r[2]), .B0(n111), .S(n112), .CO(n113));
Q_AD01HF U186 ( .A0(timer_r[3]), .B0(n113), .S(n114), .CO(n115));
Q_AD01HF U187 ( .A0(timer_r[4]), .B0(n115), .S(n116), .CO(n117));
Q_XOR2 U188 ( .A0(timer_r[5]), .A1(n117), .Z(n118));
Q_MX02 U189 ( .S(n432), .A0(n124), .A1(n120), .Z(n119));
Q_ND02 U190 ( .A0(n121), .A1(n122), .Z(n120));
Q_ND02 U191 ( .A0(n490), .A1(n396), .Z(n122));
Q_OR02 U192 ( .A0(n123), .A1(n396), .Z(n121));
Q_OR02 U193 ( .A0(n396), .A1(n492), .Z(n124));
Q_INV U194 ( .A(n125), .Z(n126));
Q_MX02 U195 ( .S(n432), .A0(n121), .A1(n127), .Z(n125));
Q_INV U196 ( .A(n128), .Z(n127));
Q_INV U197 ( .A(n129), .Z(n130));
Q_MX02 U198 ( .S(n432), .A0(n136), .A1(n131), .Z(n129));
Q_INV U199 ( .A(n132), .Z(n131));
Q_MX02 U200 ( .S(n396), .A0(n128), .A1(n133), .Z(n132));
Q_INV U201 ( .A(n134), .Z(n133));
Q_XOR2 U202 ( .A0(n490), .A1(n135), .Z(n128));
Q_OR02 U203 ( .A0(n491), .A1(n123), .Z(n136));
Q_OR02 U204 ( .A0(n490), .A1(n492), .Z(n123));
Q_NR02 U205 ( .A0(n493), .A1(n138), .Z(n137));
Q_MX02 U206 ( .S(n396), .A0(n134), .A1(n492), .Z(n138));
Q_OR02 U207 ( .A0(n490), .A1(n135), .Z(n134));
Q_INV U208 ( .A(n492), .Z(n135));
Q_AN03 U209 ( .A0(n491), .A1(n490), .A2(n493), .Z(n139));
Q_AO21 U210 ( .A0(n139), .A1(state_r[3]), .B0(n137), .Z(n519));
Q_AO21 U211 ( .A0(n139), .A1(state_r[2]), .B0(n130), .Z(n518));
Q_AO21 U212 ( .A0(n139), .A1(state_r[1]), .B0(n126), .Z(n517));
Q_AO21 U213 ( .A0(n139), .A1(state_r[0]), .B0(n119), .Z(n516));
Q_AN02 U214 ( .A0(n494), .A1(n109), .Z(n140));
Q_AN02 U215 ( .A0(n494), .A1(n110), .Z(n141));
Q_AN02 U216 ( .A0(n494), .A1(n112), .Z(n142));
Q_AN02 U217 ( .A0(n494), .A1(n114), .Z(n143));
Q_AN02 U218 ( .A0(n494), .A1(n116), .Z(n144));
Q_AN02 U219 ( .A0(n494), .A1(n118), .Z(n145));
Q_AN02 U220 ( .A0(n496), .A1(cmnd_addr[0]), .Z(n146));
Q_MX02 U221 ( .S(n497), .A0(n146), .A1(n92), .Z(n147));
Q_AN02 U222 ( .A0(n496), .A1(cmnd_addr[1]), .Z(n148));
Q_MX02 U223 ( .S(n497), .A0(n148), .A1(n94), .Z(n149));
Q_AN02 U224 ( .A0(n496), .A1(cmnd_addr[2]), .Z(n150));
Q_MX02 U225 ( .S(n497), .A0(n150), .A1(n96), .Z(n151));
Q_AN02 U226 ( .A0(n496), .A1(cmnd_addr[3]), .Z(n152));
Q_MX02 U227 ( .S(n497), .A0(n152), .A1(n98), .Z(n153));
Q_AN02 U228 ( .A0(n496), .A1(cmnd_addr[4]), .Z(n154));
Q_MX02 U229 ( .S(n497), .A0(n154), .A1(n100), .Z(n155));
Q_AN02 U230 ( .A0(n496), .A1(cmnd_addr[5]), .Z(n156));
Q_MX02 U231 ( .S(n497), .A0(n156), .A1(n102), .Z(n157));
Q_AN02 U232 ( .A0(n496), .A1(cmnd_addr[6]), .Z(n158));
Q_MX02 U233 ( .S(n497), .A0(n158), .A1(n104), .Z(n159));
Q_AN02 U234 ( .A0(n496), .A1(cmnd_addr[7]), .Z(n160));
Q_MX02 U235 ( .S(n497), .A0(n160), .A1(n106), .Z(n161));
Q_AN02 U236 ( .A0(n496), .A1(cmnd_addr[8]), .Z(n162));
Q_MX02 U237 ( .S(n497), .A0(n162), .A1(n108), .Z(n163));
Q_AN02 U238 ( .A0(n502), .A1(n91), .Z(n164));
Q_MX03 U239 ( .S0(n504), .S1(n505), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n165));
Q_MX03 U240 ( .S0(n504), .S1(n505), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n166));
Q_MX03 U241 ( .S0(n504), .S1(n505), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n167));
Q_MX03 U242 ( .S0(n504), .S1(n505), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n168));
Q_MX03 U243 ( .S0(n504), .S1(n505), .A0(sw_aindex[4]), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n169));
Q_MX03 U244 ( .S0(n504), .S1(n505), .A0(sw_aindex[5]), .A1(wr_dat[5]), .A2(sw_rdat[5]), .Z(n170));
Q_MX03 U245 ( .S0(n504), .S1(n505), .A0(sw_aindex[6]), .A1(wr_dat[6]), .A2(sw_rdat[6]), .Z(n171));
Q_MX03 U246 ( .S0(n504), .S1(n505), .A0(sw_aindex[7]), .A1(wr_dat[7]), .A2(sw_rdat[7]), .Z(n172));
Q_MX03 U247 ( .S0(n504), .S1(n505), .A0(sw_match), .A1(wr_dat[8]), .A2(sw_rdat[8]), .Z(n173));
Q_AN02 U248 ( .A0(n504), .A1(wr_dat[9]), .Z(n174));
Q_MX02 U249 ( .S(n505), .A0(n174), .A1(sw_rdat[9]), .Z(n175));
Q_AN02 U250 ( .A0(n504), .A1(wr_dat[10]), .Z(n176));
Q_MX02 U251 ( .S(n505), .A0(n176), .A1(sw_rdat[10]), .Z(n177));
Q_AN02 U252 ( .A0(n504), .A1(wr_dat[11]), .Z(n178));
Q_MX02 U253 ( .S(n505), .A0(n178), .A1(sw_rdat[11]), .Z(n179));
Q_AN02 U254 ( .A0(n504), .A1(wr_dat[12]), .Z(n180));
Q_MX02 U255 ( .S(n505), .A0(n180), .A1(sw_rdat[12]), .Z(n181));
Q_AN02 U256 ( .A0(n504), .A1(wr_dat[13]), .Z(n182));
Q_MX02 U257 ( .S(n505), .A0(n182), .A1(sw_rdat[13]), .Z(n183));
Q_AN02 U258 ( .A0(n504), .A1(wr_dat[14]), .Z(n184));
Q_MX02 U259 ( .S(n505), .A0(n184), .A1(sw_rdat[14]), .Z(n185));
Q_AN02 U260 ( .A0(n504), .A1(wr_dat[15]), .Z(n186));
Q_MX02 U261 ( .S(n505), .A0(n186), .A1(sw_rdat[15]), .Z(n187));
Q_AN02 U262 ( .A0(n504), .A1(wr_dat[16]), .Z(n188));
Q_MX02 U263 ( .S(n505), .A0(n188), .A1(sw_rdat[16]), .Z(n189));
Q_AN02 U264 ( .A0(n504), .A1(wr_dat[17]), .Z(n190));
Q_MX02 U265 ( .S(n505), .A0(n190), .A1(sw_rdat[17]), .Z(n191));
Q_AN02 U266 ( .A0(n504), .A1(wr_dat[18]), .Z(n192));
Q_MX02 U267 ( .S(n505), .A0(n192), .A1(sw_rdat[18]), .Z(n193));
Q_AN02 U268 ( .A0(n504), .A1(wr_dat[19]), .Z(n194));
Q_MX02 U269 ( .S(n505), .A0(n194), .A1(sw_rdat[19]), .Z(n195));
Q_AN02 U270 ( .A0(n504), .A1(wr_dat[20]), .Z(n196));
Q_MX02 U271 ( .S(n505), .A0(n196), .A1(sw_rdat[20]), .Z(n197));
Q_AN02 U272 ( .A0(n504), .A1(wr_dat[21]), .Z(n198));
Q_MX02 U273 ( .S(n505), .A0(n198), .A1(sw_rdat[21]), .Z(n199));
Q_AN02 U274 ( .A0(n504), .A1(wr_dat[22]), .Z(n200));
Q_MX02 U275 ( .S(n505), .A0(n200), .A1(sw_rdat[22]), .Z(n201));
Q_AN02 U276 ( .A0(n504), .A1(wr_dat[23]), .Z(n202));
Q_MX02 U277 ( .S(n505), .A0(n202), .A1(sw_rdat[23]), .Z(n203));
Q_AN02 U278 ( .A0(n504), .A1(wr_dat[24]), .Z(n204));
Q_MX02 U279 ( .S(n505), .A0(n204), .A1(sw_rdat[24]), .Z(n205));
Q_AN02 U280 ( .A0(n504), .A1(wr_dat[25]), .Z(n206));
Q_MX02 U281 ( .S(n505), .A0(n206), .A1(sw_rdat[25]), .Z(n207));
Q_AN02 U282 ( .A0(n504), .A1(wr_dat[26]), .Z(n208));
Q_MX02 U283 ( .S(n505), .A0(n208), .A1(sw_rdat[26]), .Z(n209));
Q_AN02 U284 ( .A0(n504), .A1(wr_dat[27]), .Z(n210));
Q_MX02 U285 ( .S(n505), .A0(n210), .A1(sw_rdat[27]), .Z(n211));
Q_AN02 U286 ( .A0(n504), .A1(wr_dat[28]), .Z(n212));
Q_MX02 U287 ( .S(n505), .A0(n212), .A1(sw_rdat[28]), .Z(n213));
Q_AN02 U288 ( .A0(n504), .A1(wr_dat[29]), .Z(n214));
Q_MX02 U289 ( .S(n505), .A0(n214), .A1(sw_rdat[29]), .Z(n215));
Q_AN02 U290 ( .A0(n504), .A1(wr_dat[30]), .Z(n216));
Q_MX02 U291 ( .S(n505), .A0(n216), .A1(sw_rdat[30]), .Z(n217));
Q_AN02 U292 ( .A0(n504), .A1(wr_dat[31]), .Z(n218));
Q_MX02 U293 ( .S(n505), .A0(n218), .A1(sw_rdat[31]), .Z(n219));
Q_AN02 U294 ( .A0(n504), .A1(wr_dat[32]), .Z(n220));
Q_MX02 U295 ( .S(n505), .A0(n220), .A1(sw_rdat[32]), .Z(n221));
Q_AN02 U296 ( .A0(n504), .A1(wr_dat[33]), .Z(n222));
Q_MX02 U297 ( .S(n505), .A0(n222), .A1(sw_rdat[33]), .Z(n223));
Q_AN02 U298 ( .A0(n504), .A1(wr_dat[34]), .Z(n224));
Q_MX02 U299 ( .S(n505), .A0(n224), .A1(sw_rdat[34]), .Z(n225));
Q_AN02 U300 ( .A0(n504), .A1(wr_dat[35]), .Z(n226));
Q_MX02 U301 ( .S(n505), .A0(n226), .A1(sw_rdat[35]), .Z(n227));
Q_AN02 U302 ( .A0(n504), .A1(wr_dat[36]), .Z(n228));
Q_MX02 U303 ( .S(n505), .A0(n228), .A1(sw_rdat[36]), .Z(n229));
Q_AN02 U304 ( .A0(n504), .A1(wr_dat[37]), .Z(n230));
Q_MX02 U305 ( .S(n505), .A0(n230), .A1(sw_rdat[37]), .Z(n231));
Q_AN02 U306 ( .A0(n504), .A1(wr_dat[38]), .Z(n232));
Q_MX02 U307 ( .S(n505), .A0(n232), .A1(sw_rdat[38]), .Z(n233));
Q_AN02 U308 ( .A0(n504), .A1(wr_dat[39]), .Z(n234));
Q_MX02 U309 ( .S(n505), .A0(n234), .A1(sw_rdat[39]), .Z(n235));
Q_AN02 U310 ( .A0(n504), .A1(wr_dat[40]), .Z(n236));
Q_MX02 U311 ( .S(n505), .A0(n236), .A1(sw_rdat[40]), .Z(n237));
Q_AN02 U312 ( .A0(n504), .A1(wr_dat[41]), .Z(n238));
Q_MX02 U313 ( .S(n505), .A0(n238), .A1(sw_rdat[41]), .Z(n239));
Q_AN02 U314 ( .A0(n504), .A1(wr_dat[42]), .Z(n240));
Q_MX02 U315 ( .S(n505), .A0(n240), .A1(sw_rdat[42]), .Z(n241));
Q_AN02 U316 ( .A0(n504), .A1(wr_dat[43]), .Z(n242));
Q_MX02 U317 ( .S(n505), .A0(n242), .A1(sw_rdat[43]), .Z(n243));
Q_AN02 U318 ( .A0(n504), .A1(wr_dat[44]), .Z(n244));
Q_MX02 U319 ( .S(n505), .A0(n244), .A1(sw_rdat[44]), .Z(n245));
Q_AN02 U320 ( .A0(n504), .A1(wr_dat[45]), .Z(n246));
Q_MX02 U321 ( .S(n505), .A0(n246), .A1(sw_rdat[45]), .Z(n247));
Q_AN02 U322 ( .A0(n504), .A1(wr_dat[46]), .Z(n248));
Q_MX02 U323 ( .S(n505), .A0(n248), .A1(sw_rdat[46]), .Z(n249));
Q_AN02 U324 ( .A0(n504), .A1(wr_dat[47]), .Z(n250));
Q_MX02 U325 ( .S(n505), .A0(n250), .A1(sw_rdat[47]), .Z(n251));
Q_AN02 U326 ( .A0(n504), .A1(wr_dat[48]), .Z(n252));
Q_MX02 U327 ( .S(n505), .A0(n252), .A1(sw_rdat[48]), .Z(n253));
Q_AN02 U328 ( .A0(n504), .A1(wr_dat[49]), .Z(n254));
Q_MX02 U329 ( .S(n505), .A0(n254), .A1(sw_rdat[49]), .Z(n255));
Q_AN02 U330 ( .A0(n504), .A1(wr_dat[50]), .Z(n256));
Q_MX02 U331 ( .S(n505), .A0(n256), .A1(sw_rdat[50]), .Z(n257));
Q_AN02 U332 ( .A0(n504), .A1(wr_dat[51]), .Z(n258));
Q_MX02 U333 ( .S(n505), .A0(n258), .A1(sw_rdat[51]), .Z(n259));
Q_AN02 U334 ( .A0(n504), .A1(wr_dat[52]), .Z(n260));
Q_MX02 U335 ( .S(n505), .A0(n260), .A1(sw_rdat[52]), .Z(n261));
Q_AN02 U336 ( .A0(n504), .A1(wr_dat[53]), .Z(n262));
Q_MX02 U337 ( .S(n505), .A0(n262), .A1(sw_rdat[53]), .Z(n263));
Q_AN02 U338 ( .A0(n504), .A1(wr_dat[54]), .Z(n264));
Q_MX02 U339 ( .S(n505), .A0(n264), .A1(sw_rdat[54]), .Z(n265));
Q_AN02 U340 ( .A0(n504), .A1(wr_dat[55]), .Z(n266));
Q_MX02 U341 ( .S(n505), .A0(n266), .A1(sw_rdat[55]), .Z(n267));
Q_AN02 U342 ( .A0(n504), .A1(wr_dat[56]), .Z(n268));
Q_MX02 U343 ( .S(n505), .A0(n268), .A1(sw_rdat[56]), .Z(n269));
Q_AN02 U344 ( .A0(n504), .A1(wr_dat[57]), .Z(n270));
Q_MX02 U345 ( .S(n505), .A0(n270), .A1(sw_rdat[57]), .Z(n271));
Q_AN02 U346 ( .A0(n504), .A1(wr_dat[58]), .Z(n272));
Q_MX02 U347 ( .S(n505), .A0(n272), .A1(sw_rdat[58]), .Z(n273));
Q_AN02 U348 ( .A0(n504), .A1(wr_dat[59]), .Z(n274));
Q_MX02 U349 ( .S(n505), .A0(n274), .A1(sw_rdat[59]), .Z(n275));
Q_AN02 U350 ( .A0(n504), .A1(wr_dat[60]), .Z(n276));
Q_MX02 U351 ( .S(n505), .A0(n276), .A1(sw_rdat[60]), .Z(n277));
Q_AN02 U352 ( .A0(n504), .A1(wr_dat[61]), .Z(n278));
Q_MX02 U353 ( .S(n505), .A0(n278), .A1(sw_rdat[61]), .Z(n279));
Q_AN02 U354 ( .A0(n504), .A1(wr_dat[62]), .Z(n280));
Q_MX02 U355 ( .S(n505), .A0(n280), .A1(sw_rdat[62]), .Z(n281));
Q_AN02 U356 ( .A0(n504), .A1(wr_dat[63]), .Z(n282));
Q_MX02 U357 ( .S(n505), .A0(n282), .A1(sw_rdat[63]), .Z(n283));
Q_AN02 U358 ( .A0(n504), .A1(wr_dat[64]), .Z(n284));
Q_MX02 U359 ( .S(n505), .A0(n284), .A1(sw_rdat[64]), .Z(n285));
Q_AN02 U360 ( .A0(n504), .A1(wr_dat[65]), .Z(n286));
Q_MX02 U361 ( .S(n505), .A0(n286), .A1(sw_rdat[65]), .Z(n287));
Q_AN02 U362 ( .A0(n504), .A1(wr_dat[66]), .Z(n288));
Q_MX02 U363 ( .S(n505), .A0(n288), .A1(sw_rdat[66]), .Z(n289));
Q_AN02 U364 ( .A0(n504), .A1(wr_dat[67]), .Z(n290));
Q_MX02 U365 ( .S(n505), .A0(n290), .A1(sw_rdat[67]), .Z(n291));
Q_AN02 U366 ( .A0(n504), .A1(wr_dat[68]), .Z(n292));
Q_MX02 U367 ( .S(n505), .A0(n292), .A1(sw_rdat[68]), .Z(n293));
Q_AN02 U368 ( .A0(n504), .A1(wr_dat[69]), .Z(n294));
Q_MX02 U369 ( .S(n505), .A0(n294), .A1(sw_rdat[69]), .Z(n295));
Q_AN02 U370 ( .A0(n504), .A1(wr_dat[70]), .Z(n296));
Q_MX02 U371 ( .S(n505), .A0(n296), .A1(sw_rdat[70]), .Z(n297));
Q_AN02 U372 ( .A0(n504), .A1(wr_dat[71]), .Z(n298));
Q_MX02 U373 ( .S(n505), .A0(n298), .A1(sw_rdat[71]), .Z(n299));
Q_AN02 U374 ( .A0(n504), .A1(wr_dat[72]), .Z(n300));
Q_MX02 U375 ( .S(n505), .A0(n300), .A1(sw_rdat[72]), .Z(n301));
Q_AN02 U376 ( .A0(n504), .A1(wr_dat[73]), .Z(n302));
Q_MX02 U377 ( .S(n505), .A0(n302), .A1(sw_rdat[73]), .Z(n303));
Q_AN02 U378 ( .A0(n504), .A1(wr_dat[74]), .Z(n304));
Q_MX02 U379 ( .S(n505), .A0(n304), .A1(sw_rdat[74]), .Z(n305));
Q_AN02 U380 ( .A0(n504), .A1(wr_dat[75]), .Z(n306));
Q_MX02 U381 ( .S(n505), .A0(n306), .A1(sw_rdat[75]), .Z(n307));
Q_AN02 U382 ( .A0(n504), .A1(wr_dat[76]), .Z(n308));
Q_MX02 U383 ( .S(n505), .A0(n308), .A1(sw_rdat[76]), .Z(n309));
Q_AN02 U384 ( .A0(n504), .A1(wr_dat[77]), .Z(n310));
Q_MX02 U385 ( .S(n505), .A0(n310), .A1(sw_rdat[77]), .Z(n311));
Q_AN02 U386 ( .A0(n504), .A1(wr_dat[78]), .Z(n312));
Q_MX02 U387 ( .S(n505), .A0(n312), .A1(sw_rdat[78]), .Z(n313));
Q_AN02 U388 ( .A0(n504), .A1(wr_dat[79]), .Z(n314));
Q_MX02 U389 ( .S(n505), .A0(n314), .A1(sw_rdat[79]), .Z(n315));
Q_AN02 U390 ( .A0(n504), .A1(wr_dat[80]), .Z(n316));
Q_MX02 U391 ( .S(n505), .A0(n316), .A1(sw_rdat[80]), .Z(n317));
Q_AN02 U392 ( .A0(n504), .A1(wr_dat[81]), .Z(n318));
Q_MX02 U393 ( .S(n505), .A0(n318), .A1(sw_rdat[81]), .Z(n319));
Q_AN02 U394 ( .A0(n504), .A1(wr_dat[82]), .Z(n320));
Q_MX02 U395 ( .S(n505), .A0(n320), .A1(sw_rdat[82]), .Z(n321));
Q_AN02 U396 ( .A0(n504), .A1(wr_dat[83]), .Z(n322));
Q_MX02 U397 ( .S(n505), .A0(n322), .A1(sw_rdat[83]), .Z(n323));
Q_AN02 U398 ( .A0(n504), .A1(wr_dat[84]), .Z(n324));
Q_MX02 U399 ( .S(n505), .A0(n324), .A1(sw_rdat[84]), .Z(n325));
Q_AN02 U400 ( .A0(n504), .A1(wr_dat[85]), .Z(n326));
Q_MX02 U401 ( .S(n505), .A0(n326), .A1(sw_rdat[85]), .Z(n327));
Q_AN02 U402 ( .A0(n504), .A1(wr_dat[86]), .Z(n328));
Q_MX02 U403 ( .S(n505), .A0(n328), .A1(sw_rdat[86]), .Z(n329));
Q_AN02 U404 ( .A0(n504), .A1(wr_dat[87]), .Z(n330));
Q_MX02 U405 ( .S(n505), .A0(n330), .A1(sw_rdat[87]), .Z(n331));
Q_AN02 U406 ( .A0(n504), .A1(wr_dat[88]), .Z(n332));
Q_MX02 U407 ( .S(n505), .A0(n332), .A1(sw_rdat[88]), .Z(n333));
Q_AN02 U408 ( .A0(n504), .A1(wr_dat[89]), .Z(n334));
Q_MX02 U409 ( .S(n505), .A0(n334), .A1(sw_rdat[89]), .Z(n335));
Q_AN02 U410 ( .A0(n504), .A1(wr_dat[90]), .Z(n336));
Q_MX02 U411 ( .S(n505), .A0(n336), .A1(sw_rdat[90]), .Z(n337));
Q_AN02 U412 ( .A0(n504), .A1(wr_dat[91]), .Z(n338));
Q_MX02 U413 ( .S(n505), .A0(n338), .A1(sw_rdat[91]), .Z(n339));
Q_AN02 U414 ( .A0(n504), .A1(wr_dat[92]), .Z(n340));
Q_MX02 U415 ( .S(n505), .A0(n340), .A1(sw_rdat[92]), .Z(n341));
Q_AN02 U416 ( .A0(n504), .A1(wr_dat[93]), .Z(n342));
Q_MX02 U417 ( .S(n505), .A0(n342), .A1(sw_rdat[93]), .Z(n343));
Q_AN02 U418 ( .A0(n504), .A1(wr_dat[94]), .Z(n344));
Q_MX02 U419 ( .S(n505), .A0(n344), .A1(sw_rdat[94]), .Z(n345));
Q_AN02 U420 ( .A0(n504), .A1(wr_dat[95]), .Z(n346));
Q_MX02 U421 ( .S(n505), .A0(n346), .A1(sw_rdat[95]), .Z(n347));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n519), .Q(state_r[3]), .QN(n405));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n518), .Q(state_r[2]), .QN(n406));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n517), .Q(state_r[1]), .QN(n408));
Q_FDP1 \state_r_REG[0] ( .CK(clk), .R(rst_n), .D(n516), .Q(state_r[0]), .QN(n377));
Q_FDP1 \timer_r_REG[5] ( .CK(clk), .R(rst_n), .D(n145), .Q(timer_r[5]), .QN( ));
Q_FDP1 \timer_r_REG[4] ( .CK(clk), .R(rst_n), .D(n144), .Q(timer_r[4]), .QN( ));
Q_FDP1 \timer_r_REG[3] ( .CK(clk), .R(rst_n), .D(n143), .Q(timer_r[3]), .QN( ));
Q_FDP1 \timer_r_REG[2] ( .CK(clk), .R(rst_n), .D(n142), .Q(timer_r[2]), .QN( ));
Q_FDP1 \timer_r_REG[1] ( .CK(clk), .R(rst_n), .D(n141), .Q(timer_r[1]), .QN( ));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n140), .Q(timer_r[0]), .QN(n109));
Q_ND02 U432 ( .A0(n349), .A1(n350), .Z(n348));
Q_ND02 U433 ( .A0(n351), .A1(n463), .Z(n350));
Q_OR02 U434 ( .A0(n352), .A1(n507), .Z(n351));
Q_INV U435 ( .A(n506), .Z(n352));
Q_ND02 U436 ( .A0(n349), .A1(n354), .Z(n353));
Q_ND02 U437 ( .A0(n506), .A1(n463), .Z(n354));
Q_OR03 U438 ( .A0(n506), .A1(n507), .A2(n463), .Z(n349));
Q_MX02 U439 ( .S(n463), .A0(n506), .A1(n507), .Z(n355));
Q_FDP2 \stat_code_REG[2] ( .CK(clk), .S(rst_n), .D(n356), .Q(stat_code[2]), .QN( ));
Q_MX02 U441 ( .S(n478), .A0(stat_code[2]), .A1(n355), .Z(n356));
Q_FDP2 \stat_code_REG[1] ( .CK(clk), .S(rst_n), .D(n357), .Q(stat_code[1]), .QN( ));
Q_MX02 U443 ( .S(n478), .A0(stat_code[1]), .A1(n353), .Z(n357));
Q_FDP2 \stat_code_REG[0] ( .CK(clk), .S(rst_n), .D(n358), .Q(stat_code[0]), .QN( ));
Q_MX02 U445 ( .S(n478), .A0(stat_code[0]), .A1(n348), .Z(n358));
Q_FDP2 init_r_REG  ( .CK(clk), .S(rst_n), .D(n359), .Q(init_r), .QN(enable));
Q_MX02 U447 ( .S(n509), .A0(init_r), .A1(n503), .Z(n359));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n501), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n500), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n499), .Q(rst_r), .QN(n520));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n498), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n495), .Q(sw_we_r), .QN( ));
Q_OA21 U453 ( .A0(n361), .A1(n362), .B0(n360), .Z(n490));
Q_OR03 U454 ( .A0(n364), .A1(n365), .A2(n363), .Z(n362));
Q_AN03 U455 ( .A0(state_r[0]), .A1(n368), .A2(n366), .Z(n367));
Q_AN02 U456 ( .A0(n63), .A1(cmnd_rd_stb), .Z(n368));
Q_AN02 U457 ( .A0(n371), .A1(n60), .Z(n372));
Q_AN03 U458 ( .A0(n373), .A1(n372), .A2(n369), .Z(n370));
Q_AN02 U459 ( .A0(n374), .A1(state_r[0]), .Z(n373));
Q_OR03 U460 ( .A0(n370), .A1(n375), .A2(n367), .Z(n365));
Q_AN02 U461 ( .A0(n366), .A1(n376), .Z(n375));
Q_NR02 U462 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n376));
Q_OA21 U463 ( .A0(n379), .A1(n380), .B0(n378), .Z(n364));
Q_AN02 U464 ( .A0(n381), .A1(n382), .Z(n380));
Q_NR02 U465 ( .A0(state_r[0]), .A1(igrant), .Z(n382));
Q_OA21 U466 ( .A0(n385), .A1(n386), .B0(n384), .Z(n379));
Q_AN02 U467 ( .A0(n387), .A1(n383), .Z(n386));
Q_NR02 U468 ( .A0(n388), .A1(n515), .Z(n385));
Q_INV U469 ( .A(n389), .Z(n371));
Q_AN03 U470 ( .A0(cmnd_rst_stb), .A1(n366), .A2(n391), .Z(n392));
Q_OR03 U471 ( .A0(n393), .A1(n392), .A2(n390), .Z(n361));
Q_AN03 U472 ( .A0(n377), .A1(n395), .A2(n394), .Z(n393));
Q_INV U473 ( .A(n396), .Z(n491));
Q_OA21 U474 ( .A0(n397), .A1(n363), .B0(n360), .Z(n396));
Q_AO21 U475 ( .A0(n366), .A1(n400), .B0(n399), .Z(n397));
Q_AN02 U476 ( .A0(state_r[0]), .A1(cmnd_wr_stb), .Z(n400));
Q_AN03 U477 ( .A0(n404), .A1(n377), .A2(n402), .Z(n403));
Q_NR02 U478 ( .A0(state_r[3]), .A1(state_r[2]), .Z(n404));
Q_MX02 U479 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n407), .Z(n402));
Q_OR03 U480 ( .A0(n409), .A1(n403), .A2(n401), .Z(n363));
Q_AN02 U481 ( .A0(n410), .A1(n378), .Z(n401));
Q_AN02 U482 ( .A0(n374), .A1(n60), .Z(n378));
Q_AN02 U483 ( .A0(n411), .A1(n412), .Z(n409));
Q_NR02 U484 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n412));
Q_MX02 U485 ( .S(state_r[3]), .A0(n414), .A1(n413), .Z(n410));
Q_AN02 U486 ( .A0(n449), .A1(n407), .Z(n415));
Q_AN02 U487 ( .A0(ack_error), .A1(enable), .Z(n407));
Q_AO21 U488 ( .A0(n416), .A1(n377), .B0(n415), .Z(n413));
Q_AN02 U489 ( .A0(state_r[2]), .A1(igrant), .Z(n418));
Q_AO21 U490 ( .A0(n419), .A1(n420), .B0(n417), .Z(n414));
Q_OA21 U491 ( .A0(state_r[0]), .A1(n421), .B0(n418), .Z(n417));
Q_AN02 U492 ( .A0(n408), .A1(n515), .Z(n421));
Q_OR02 U493 ( .A0(state_r[2]), .A1(n389), .Z(n419));
Q_AN02 U494 ( .A0(igrant), .A1(n514), .Z(n389));
Q_OA21 U495 ( .A0(n422), .A1(n423), .B0(n398), .Z(n399));
Q_AN03 U496 ( .A0(n424), .A1(n405), .A2(n391), .Z(n423));
Q_AN02 U497 ( .A0(n425), .A1(n426), .Z(n422));
Q_AN03 U498 ( .A0(n428), .A1(n429), .A2(n427), .Z(n492));
Q_AO21 U499 ( .A0(n424), .A1(n431), .B0(n430), .Z(n427));
Q_INV U500 ( .A(n430), .Z(n431));
Q_INV U501 ( .A(n432), .Z(n493));
Q_OA21 U502 ( .A0(n433), .A1(n390), .B0(n360), .Z(n432));
Q_AN03 U503 ( .A0(n430), .A1(n429), .A2(n366), .Z(n434));
Q_AN02 U504 ( .A0(state_r[0]), .A1(n63), .Z(n429));
Q_AO21 U505 ( .A0(n64), .A1(cmnd_cmp_stb), .B0(cmnd_rd_stb), .Z(n430));
Q_AN03 U506 ( .A0(n424), .A1(n366), .A2(n391), .Z(n435));
Q_AN02 U507 ( .A0(n436), .A1(n61), .Z(n391));
Q_AO21 U508 ( .A0(n62), .A1(n513), .B0(cmnd_rst_stb), .Z(n424));
Q_AN03 U509 ( .A0(n425), .A1(n60), .A2(n394), .Z(n438));
Q_AN02 U510 ( .A0(n374), .A1(n381), .Z(n394));
Q_AN02 U511 ( .A0(state_r[3]), .A1(n398), .Z(n381));
Q_OR03 U512 ( .A0(n438), .A1(n437), .A2(n434), .Z(n433));
Q_AO21 U513 ( .A0(n439), .A1(n440), .B0(n435), .Z(n437));
Q_AN02 U514 ( .A0(igrant), .A1(n60), .Z(n395));
Q_AN02 U515 ( .A0(n441), .A1(n395), .Z(n439));
Q_NR02 U516 ( .A0(timeout), .A1(state_r[0]), .Z(n441));
Q_AN02 U517 ( .A0(ack_error), .A1(init_r), .Z(n443));
Q_AO21 U518 ( .A0(n411), .A1(cmnd_dis_stb), .B0(n442), .Z(n390));
Q_AN02 U519 ( .A0(n436), .A1(n445), .Z(n444));
Q_NR02 U520 ( .A0(cmnd_cmp_stb), .A1(n513), .Z(n445));
Q_AN02 U521 ( .A0(state_r[0]), .A1(n446), .Z(n436));
Q_NR02 U522 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n446));
Q_AN03 U523 ( .A0(n62), .A1(n366), .A2(n444), .Z(n411));
Q_OA21 U524 ( .A0(n447), .A1(n448), .B0(n443), .Z(n442));
Q_AN02 U525 ( .A0(n449), .A1(n426), .Z(n447));
Q_AN03 U526 ( .A0(n374), .A1(state_r[3]), .A2(n60), .Z(n426));
Q_INV U527 ( .A(n387), .Z(n420));
Q_AO21 U528 ( .A0(n377), .A1(igrant), .B0(state_r[0]), .Z(n425));
Q_AN02 U529 ( .A0(n383), .A1(n501), .Z(n494));
Q_INV U530 ( .A(igrant), .Z(n383));
Q_OA21 U531 ( .A0(n451), .A1(n452), .B0(n450), .Z(n495));
Q_AN02 U532 ( .A0(n518), .A1(n453), .Z(n452));
Q_AN02 U533 ( .A0(cmnd_sis_stb), .A1(n454), .Z(n496));
Q_INV U534 ( .A(n497), .Z(n454));
Q_ND02 U535 ( .A0(n387), .A1(n406), .Z(n449));
Q_OR02 U536 ( .A0(state_r[0]), .A1(state_r[1]), .Z(n388));
Q_ND02 U537 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n387));
Q_OA21 U538 ( .A0(n451), .A1(n455), .B0(n450), .Z(n498));
Q_AN02 U539 ( .A0(n518), .A1(n456), .Z(n455));
Q_AN02 U540 ( .A0(n457), .A1(n458), .Z(n451));
Q_AN02 U541 ( .A0(n459), .A1(n458), .Z(n499));
Q_OR03 U542 ( .A0(n460), .A1(n500), .A2(n499), .Z(n501));
Q_AN03 U543 ( .A0(n519), .A1(n457), .A2(n456), .Z(n500));
Q_AN03 U544 ( .A0(n450), .A1(n518), .A2(n461), .Z(n460));
Q_INV U545 ( .A(n458), .Z(n461));
Q_INV U546 ( .A(n462), .Z(n502));
Q_AN02 U547 ( .A0(n440), .A1(state_r[0]), .Z(n505));
Q_AN03 U548 ( .A0(state_r[2]), .A1(state_r[1]), .A2(n405), .Z(n440));
Q_AN02 U549 ( .A0(n465), .A1(n466), .Z(n467));
Q_INV U550 ( .A(n468), .Z(n465));
Q_OR03 U551 ( .A0(n469), .A1(n467), .A2(n464), .Z(n463));
Q_AN03 U552 ( .A0(n471), .A1(n59), .A2(n470), .Z(n464));
Q_OR02 U553 ( .A0(n458), .A1(n472), .Z(n469));
Q_AN02 U554 ( .A0(n517), .A1(n516), .Z(n458));
Q_INV U555 ( .A(n459), .Z(n472));
Q_AN02 U556 ( .A0(n459), .A1(n473), .Z(n466));
Q_OA21 U557 ( .A0(n474), .A1(n453), .B0(n466), .Z(n506));
Q_AN02 U558 ( .A0(n59), .A1(n517), .Z(n468));
Q_OA21 U559 ( .A0(n471), .A1(badaddr), .B0(n468), .Z(n474));
Q_AN02 U560 ( .A0(timeout), .A1(n360), .Z(n471));
Q_OA21 U561 ( .A0(n475), .A1(n476), .B0(n459), .Z(n507));
Q_AO21 U562 ( .A0(n453), .A1(n516), .B0(n456), .Z(n476));
Q_AN02 U563 ( .A0(unsupported_op), .A1(n477), .Z(n475));
Q_ND02 U564 ( .A0(n448), .A1(n470), .Z(n478));
Q_AN02 U565 ( .A0(n459), .A1(n477), .Z(n470));
Q_AN02 U566 ( .A0(n517), .A1(n473), .Z(n477));
Q_AN02 U567 ( .A0(n369), .A1(n377), .Z(n448));
Q_AN02 U568 ( .A0(n405), .A1(n416), .Z(n369));
Q_OA21 U569 ( .A0(n504), .A1(n479), .B0(n360), .Z(n508));
Q_AN02 U570 ( .A0(n480), .A1(state_r[1]), .Z(n479));
Q_INV U571 ( .A(n503), .Z(n504));
Q_AN02 U572 ( .A0(n405), .A1(n398), .Z(n366));
Q_MX02 U573 ( .S(state_r[0]), .A0(n481), .A1(n384), .Z(n480));
Q_AN02 U574 ( .A0(state_r[3]), .A1(n406), .Z(n481));
Q_AN02 U575 ( .A0(n405), .A1(state_r[2]), .Z(n384));
Q_AN03 U576 ( .A0(n459), .A1(n456), .A2(n503), .Z(n482));
Q_NR02 U577 ( .A0(n517), .A1(n516), .Z(n456));
Q_INV U578 ( .A(n516), .Z(n473));
Q_INV U579 ( .A(n517), .Z(n453));
Q_NR02 U580 ( .A0(n519), .A1(n518), .Z(n459));
Q_INV U581 ( .A(n518), .Z(n457));
Q_INV U582 ( .A(n519), .Z(n450));
Q_AO21 U583 ( .A0(n428), .A1(n483), .B0(n482), .Z(n509));
Q_AN02 U584 ( .A0(n377), .A1(cmnd_ena_stb), .Z(n483));
Q_OR02 U585 ( .A0(state_r[3]), .A1(state_r[1]), .Z(n484));
Q_OR03 U586 ( .A0(state_r[2]), .A1(state_r[0]), .A2(n484), .Z(n503));
Q_AN03 U587 ( .A0(n486), .A1(n408), .A2(n485), .Z(n510));
Q_AO21 U588 ( .A0(state_r[2]), .A1(n377), .B0(n462), .Z(n485));
Q_AN02 U589 ( .A0(n406), .A1(state_r[0]), .Z(n462));
Q_ND02 U590 ( .A0(n428), .A1(state_r[0]), .Z(n511));
Q_AN02 U591 ( .A0(n486), .A1(n398), .Z(n428));
Q_NR02 U592 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n398));
Q_AN02 U593 ( .A0(n487), .A1(n486), .Z(n497));
Q_NR02 U594 ( .A0(badaddr), .A1(state_r[3]), .Z(n486));
Q_INV U595 ( .A(badaddr), .Z(n360));
Q_OR03 U596 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n497), .Z(n512));
Q_MX02 U597 ( .S(state_r[0]), .A0(n488), .A1(n416), .Z(n487));
Q_AN02 U598 ( .A0(state_r[2]), .A1(n408), .Z(n488));
Q_AN02 U599 ( .A0(n406), .A1(state_r[1]), .Z(n416));
Q_OR02 U600 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n489));
Q_INV U601 ( .A(timeout), .Z(n374));
Q_AN02 U602 ( .A0(n520), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U603 ( .A0(n520), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U604 ( .A0(n520), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U605 ( .A0(n520), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U606 ( .A0(n520), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U607 ( .A0(n520), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U608 ( .A0(n520), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U609 ( .A0(n520), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U610 ( .A0(n520), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U611 ( .A0(n520), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U612 ( .A0(n520), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U613 ( .A0(n520), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U614 ( .A0(n520), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U615 ( .A0(n520), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U616 ( .A0(n520), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U617 ( .A0(n520), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U618 ( .A0(n520), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U619 ( .A0(n520), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U620 ( .A0(n520), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U621 ( .A0(n520), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U622 ( .A0(n520), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U623 ( .A0(n520), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U624 ( .A0(n520), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U625 ( .A0(n520), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U626 ( .A0(n520), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U627 ( .A0(n520), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U628 ( .A0(n520), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U629 ( .A0(n520), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U630 ( .A0(n520), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U631 ( .A0(n520), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U632 ( .A0(n520), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U633 ( .A0(n520), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_AN02 U634 ( .A0(n520), .A1(wr_dat[32]), .Z(sw_wdat[32]));
Q_AN02 U635 ( .A0(n520), .A1(wr_dat[33]), .Z(sw_wdat[33]));
Q_AN02 U636 ( .A0(n520), .A1(wr_dat[34]), .Z(sw_wdat[34]));
Q_AN02 U637 ( .A0(n520), .A1(wr_dat[35]), .Z(sw_wdat[35]));
Q_AN02 U638 ( .A0(n520), .A1(wr_dat[36]), .Z(sw_wdat[36]));
Q_AN02 U639 ( .A0(n520), .A1(wr_dat[37]), .Z(sw_wdat[37]));
Q_AN02 U640 ( .A0(n520), .A1(wr_dat[38]), .Z(sw_wdat[38]));
Q_AN02 U641 ( .A0(n520), .A1(wr_dat[39]), .Z(sw_wdat[39]));
Q_AN02 U642 ( .A0(n520), .A1(wr_dat[40]), .Z(sw_wdat[40]));
Q_AN02 U643 ( .A0(n520), .A1(wr_dat[41]), .Z(sw_wdat[41]));
Q_AN02 U644 ( .A0(n520), .A1(wr_dat[42]), .Z(sw_wdat[42]));
Q_AN02 U645 ( .A0(n520), .A1(wr_dat[43]), .Z(sw_wdat[43]));
Q_AN02 U646 ( .A0(n520), .A1(wr_dat[44]), .Z(sw_wdat[44]));
Q_AN02 U647 ( .A0(n520), .A1(wr_dat[45]), .Z(sw_wdat[45]));
Q_AN02 U648 ( .A0(n520), .A1(wr_dat[46]), .Z(sw_wdat[46]));
Q_AN02 U649 ( .A0(n520), .A1(wr_dat[47]), .Z(sw_wdat[47]));
Q_AN02 U650 ( .A0(n520), .A1(wr_dat[48]), .Z(sw_wdat[48]));
Q_AN02 U651 ( .A0(n520), .A1(wr_dat[49]), .Z(sw_wdat[49]));
Q_AN02 U652 ( .A0(n520), .A1(wr_dat[50]), .Z(sw_wdat[50]));
Q_AN02 U653 ( .A0(n520), .A1(wr_dat[51]), .Z(sw_wdat[51]));
Q_AN02 U654 ( .A0(n520), .A1(wr_dat[52]), .Z(sw_wdat[52]));
Q_AN02 U655 ( .A0(n520), .A1(wr_dat[53]), .Z(sw_wdat[53]));
Q_AN02 U656 ( .A0(n520), .A1(wr_dat[54]), .Z(sw_wdat[54]));
Q_AN02 U657 ( .A0(n520), .A1(wr_dat[55]), .Z(sw_wdat[55]));
Q_AN02 U658 ( .A0(n520), .A1(wr_dat[56]), .Z(sw_wdat[56]));
Q_AN02 U659 ( .A0(n520), .A1(wr_dat[57]), .Z(sw_wdat[57]));
Q_AN02 U660 ( .A0(n520), .A1(wr_dat[58]), .Z(sw_wdat[58]));
Q_AN02 U661 ( .A0(n520), .A1(wr_dat[59]), .Z(sw_wdat[59]));
Q_AN02 U662 ( .A0(n520), .A1(wr_dat[60]), .Z(sw_wdat[60]));
Q_AN02 U663 ( .A0(n520), .A1(wr_dat[61]), .Z(sw_wdat[61]));
Q_AN02 U664 ( .A0(n520), .A1(wr_dat[62]), .Z(sw_wdat[62]));
Q_AN02 U665 ( .A0(n520), .A1(wr_dat[63]), .Z(sw_wdat[63]));
Q_AN02 U666 ( .A0(n520), .A1(wr_dat[64]), .Z(sw_wdat[64]));
Q_AN02 U667 ( .A0(n520), .A1(wr_dat[65]), .Z(sw_wdat[65]));
Q_AN02 U668 ( .A0(n520), .A1(wr_dat[66]), .Z(sw_wdat[66]));
Q_AN02 U669 ( .A0(n520), .A1(wr_dat[67]), .Z(sw_wdat[67]));
Q_AN02 U670 ( .A0(n520), .A1(wr_dat[68]), .Z(sw_wdat[68]));
Q_AN02 U671 ( .A0(n520), .A1(wr_dat[69]), .Z(sw_wdat[69]));
Q_AN02 U672 ( .A0(n520), .A1(wr_dat[70]), .Z(sw_wdat[70]));
Q_AN02 U673 ( .A0(n520), .A1(wr_dat[71]), .Z(sw_wdat[71]));
Q_AN02 U674 ( .A0(n520), .A1(wr_dat[72]), .Z(sw_wdat[72]));
Q_AN02 U675 ( .A0(n520), .A1(wr_dat[73]), .Z(sw_wdat[73]));
Q_AN02 U676 ( .A0(n520), .A1(wr_dat[74]), .Z(sw_wdat[74]));
Q_AN02 U677 ( .A0(n520), .A1(wr_dat[75]), .Z(sw_wdat[75]));
Q_AN02 U678 ( .A0(n520), .A1(wr_dat[76]), .Z(sw_wdat[76]));
Q_AN02 U679 ( .A0(n520), .A1(wr_dat[77]), .Z(sw_wdat[77]));
Q_AN02 U680 ( .A0(n520), .A1(wr_dat[78]), .Z(sw_wdat[78]));
Q_AN02 U681 ( .A0(n520), .A1(wr_dat[79]), .Z(sw_wdat[79]));
Q_AN02 U682 ( .A0(n520), .A1(wr_dat[80]), .Z(sw_wdat[80]));
Q_AN02 U683 ( .A0(n520), .A1(wr_dat[81]), .Z(sw_wdat[81]));
Q_AN02 U684 ( .A0(n520), .A1(wr_dat[82]), .Z(sw_wdat[82]));
Q_AN02 U685 ( .A0(n520), .A1(wr_dat[83]), .Z(sw_wdat[83]));
Q_AN02 U686 ( .A0(n520), .A1(wr_dat[84]), .Z(sw_wdat[84]));
Q_AN02 U687 ( .A0(n520), .A1(wr_dat[85]), .Z(sw_wdat[85]));
Q_AN02 U688 ( .A0(n520), .A1(wr_dat[86]), .Z(sw_wdat[86]));
Q_AN02 U689 ( .A0(n520), .A1(wr_dat[87]), .Z(sw_wdat[87]));
Q_AN02 U690 ( .A0(n520), .A1(wr_dat[88]), .Z(sw_wdat[88]));
Q_AN02 U691 ( .A0(n520), .A1(wr_dat[89]), .Z(sw_wdat[89]));
Q_AN02 U692 ( .A0(n520), .A1(wr_dat[90]), .Z(sw_wdat[90]));
Q_AN02 U693 ( .A0(n520), .A1(wr_dat[91]), .Z(sw_wdat[91]));
Q_AN02 U694 ( .A0(n520), .A1(wr_dat[92]), .Z(sw_wdat[92]));
Q_AN02 U695 ( .A0(n520), .A1(wr_dat[93]), .Z(sw_wdat[93]));
Q_AN02 U696 ( .A0(n520), .A1(wr_dat[94]), .Z(sw_wdat[94]));
Q_AN02 U697 ( .A0(n520), .A1(wr_dat[95]), .Z(sw_wdat[95]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n489), .R(n521), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U699 ( .A(rst_n), .Z(n521));
Q_INV U700 ( .A(sim_tmo_r), .Z(n36));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n512), .R(n521), .D(n147), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n512), .R(n521), .D(n149), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n512), .R(n521), .D(n151), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n512), .R(n521), .D(n153), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n512), .R(n521), .D(n155), .Q(rst_addr_r[4]));
Q_FDP4EP \rst_addr_r_REG[5] ( .CK(clk), .CE(n512), .R(n521), .D(n157), .Q(rst_addr_r[5]));
Q_FDP4EP \rst_addr_r_REG[6] ( .CK(clk), .CE(n512), .R(n521), .D(n159), .Q(rst_addr_r[6]));
Q_FDP4EP \rst_addr_r_REG[7] ( .CK(clk), .CE(n512), .R(n521), .D(n161), .Q(rst_addr_r[7]));
Q_FDP4EP \rst_addr_r_REG[8] ( .CK(clk), .CE(n512), .R(n521), .D(n163), .Q(rst_addr_r[8]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n510), .R(n521), .D(n164), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n508), .R(n521), .D(n165), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n508), .R(n521), .D(n166), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n508), .R(n521), .D(n167), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n508), .R(n521), .D(n168), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n508), .R(n521), .D(n169), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n508), .R(n521), .D(n170), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n508), .R(n521), .D(n171), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n508), .R(n521), .D(n172), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n508), .R(n521), .D(n173), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n508), .R(n521), .D(n175), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n508), .R(n521), .D(n177), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n508), .R(n521), .D(n179), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n508), .R(n521), .D(n181), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n508), .R(n521), .D(n183), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n508), .R(n521), .D(n185), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n508), .R(n521), .D(n187), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n508), .R(n521), .D(n189), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n508), .R(n521), .D(n191), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n508), .R(n521), .D(n193), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n508), .R(n521), .D(n195), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n508), .R(n521), .D(n197), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n508), .R(n521), .D(n199), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n508), .R(n521), .D(n201), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n508), .R(n521), .D(n203), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n508), .R(n521), .D(n205), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n508), .R(n521), .D(n207), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n508), .R(n521), .D(n209), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n508), .R(n521), .D(n211), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n508), .R(n521), .D(n213), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n508), .R(n521), .D(n215), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n508), .R(n521), .D(n217), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n508), .R(n521), .D(n219), .Q(rd_dat[31]));
Q_FDP4EP \rd_dat_REG[32] ( .CK(clk), .CE(n508), .R(n521), .D(n221), .Q(rd_dat[32]));
Q_FDP4EP \rd_dat_REG[33] ( .CK(clk), .CE(n508), .R(n521), .D(n223), .Q(rd_dat[33]));
Q_FDP4EP \rd_dat_REG[34] ( .CK(clk), .CE(n508), .R(n521), .D(n225), .Q(rd_dat[34]));
Q_FDP4EP \rd_dat_REG[35] ( .CK(clk), .CE(n508), .R(n521), .D(n227), .Q(rd_dat[35]));
Q_FDP4EP \rd_dat_REG[36] ( .CK(clk), .CE(n508), .R(n521), .D(n229), .Q(rd_dat[36]));
Q_FDP4EP \rd_dat_REG[37] ( .CK(clk), .CE(n508), .R(n521), .D(n231), .Q(rd_dat[37]));
Q_FDP4EP \rd_dat_REG[38] ( .CK(clk), .CE(n508), .R(n521), .D(n233), .Q(rd_dat[38]));
Q_FDP4EP \rd_dat_REG[39] ( .CK(clk), .CE(n508), .R(n521), .D(n235), .Q(rd_dat[39]));
Q_FDP4EP \rd_dat_REG[40] ( .CK(clk), .CE(n508), .R(n521), .D(n237), .Q(rd_dat[40]));
Q_FDP4EP \rd_dat_REG[41] ( .CK(clk), .CE(n508), .R(n521), .D(n239), .Q(rd_dat[41]));
Q_FDP4EP \rd_dat_REG[42] ( .CK(clk), .CE(n508), .R(n521), .D(n241), .Q(rd_dat[42]));
Q_FDP4EP \rd_dat_REG[43] ( .CK(clk), .CE(n508), .R(n521), .D(n243), .Q(rd_dat[43]));
Q_FDP4EP \rd_dat_REG[44] ( .CK(clk), .CE(n508), .R(n521), .D(n245), .Q(rd_dat[44]));
Q_FDP4EP \rd_dat_REG[45] ( .CK(clk), .CE(n508), .R(n521), .D(n247), .Q(rd_dat[45]));
Q_FDP4EP \rd_dat_REG[46] ( .CK(clk), .CE(n508), .R(n521), .D(n249), .Q(rd_dat[46]));
Q_FDP4EP \rd_dat_REG[47] ( .CK(clk), .CE(n508), .R(n521), .D(n251), .Q(rd_dat[47]));
Q_FDP4EP \rd_dat_REG[48] ( .CK(clk), .CE(n508), .R(n521), .D(n253), .Q(rd_dat[48]));
Q_FDP4EP \rd_dat_REG[49] ( .CK(clk), .CE(n508), .R(n521), .D(n255), .Q(rd_dat[49]));
Q_FDP4EP \rd_dat_REG[50] ( .CK(clk), .CE(n508), .R(n521), .D(n257), .Q(rd_dat[50]));
Q_FDP4EP \rd_dat_REG[51] ( .CK(clk), .CE(n508), .R(n521), .D(n259), .Q(rd_dat[51]));
Q_FDP4EP \rd_dat_REG[52] ( .CK(clk), .CE(n508), .R(n521), .D(n261), .Q(rd_dat[52]));
Q_FDP4EP \rd_dat_REG[53] ( .CK(clk), .CE(n508), .R(n521), .D(n263), .Q(rd_dat[53]));
Q_FDP4EP \rd_dat_REG[54] ( .CK(clk), .CE(n508), .R(n521), .D(n265), .Q(rd_dat[54]));
Q_FDP4EP \rd_dat_REG[55] ( .CK(clk), .CE(n508), .R(n521), .D(n267), .Q(rd_dat[55]));
Q_FDP4EP \rd_dat_REG[56] ( .CK(clk), .CE(n508), .R(n521), .D(n269), .Q(rd_dat[56]));
Q_FDP4EP \rd_dat_REG[57] ( .CK(clk), .CE(n508), .R(n521), .D(n271), .Q(rd_dat[57]));
Q_FDP4EP \rd_dat_REG[58] ( .CK(clk), .CE(n508), .R(n521), .D(n273), .Q(rd_dat[58]));
Q_FDP4EP \rd_dat_REG[59] ( .CK(clk), .CE(n508), .R(n521), .D(n275), .Q(rd_dat[59]));
Q_FDP4EP \rd_dat_REG[60] ( .CK(clk), .CE(n508), .R(n521), .D(n277), .Q(rd_dat[60]));
Q_FDP4EP \rd_dat_REG[61] ( .CK(clk), .CE(n508), .R(n521), .D(n279), .Q(rd_dat[61]));
Q_FDP4EP \rd_dat_REG[62] ( .CK(clk), .CE(n508), .R(n521), .D(n281), .Q(rd_dat[62]));
Q_FDP4EP \rd_dat_REG[63] ( .CK(clk), .CE(n508), .R(n521), .D(n283), .Q(rd_dat[63]));
Q_FDP4EP \rd_dat_REG[64] ( .CK(clk), .CE(n508), .R(n521), .D(n285), .Q(rd_dat[64]));
Q_FDP4EP \rd_dat_REG[65] ( .CK(clk), .CE(n508), .R(n521), .D(n287), .Q(rd_dat[65]));
Q_FDP4EP \rd_dat_REG[66] ( .CK(clk), .CE(n508), .R(n521), .D(n289), .Q(rd_dat[66]));
Q_FDP4EP \rd_dat_REG[67] ( .CK(clk), .CE(n508), .R(n521), .D(n291), .Q(rd_dat[67]));
Q_FDP4EP \rd_dat_REG[68] ( .CK(clk), .CE(n508), .R(n521), .D(n293), .Q(rd_dat[68]));
Q_FDP4EP \rd_dat_REG[69] ( .CK(clk), .CE(n508), .R(n521), .D(n295), .Q(rd_dat[69]));
Q_FDP4EP \rd_dat_REG[70] ( .CK(clk), .CE(n508), .R(n521), .D(n297), .Q(rd_dat[70]));
Q_FDP4EP \rd_dat_REG[71] ( .CK(clk), .CE(n508), .R(n521), .D(n299), .Q(rd_dat[71]));
Q_FDP4EP \rd_dat_REG[72] ( .CK(clk), .CE(n508), .R(n521), .D(n301), .Q(rd_dat[72]));
Q_FDP4EP \rd_dat_REG[73] ( .CK(clk), .CE(n508), .R(n521), .D(n303), .Q(rd_dat[73]));
Q_FDP4EP \rd_dat_REG[74] ( .CK(clk), .CE(n508), .R(n521), .D(n305), .Q(rd_dat[74]));
Q_FDP4EP \rd_dat_REG[75] ( .CK(clk), .CE(n508), .R(n521), .D(n307), .Q(rd_dat[75]));
Q_FDP4EP \rd_dat_REG[76] ( .CK(clk), .CE(n508), .R(n521), .D(n309), .Q(rd_dat[76]));
Q_FDP4EP \rd_dat_REG[77] ( .CK(clk), .CE(n508), .R(n521), .D(n311), .Q(rd_dat[77]));
Q_FDP4EP \rd_dat_REG[78] ( .CK(clk), .CE(n508), .R(n521), .D(n313), .Q(rd_dat[78]));
Q_FDP4EP \rd_dat_REG[79] ( .CK(clk), .CE(n508), .R(n521), .D(n315), .Q(rd_dat[79]));
Q_FDP4EP \rd_dat_REG[80] ( .CK(clk), .CE(n508), .R(n521), .D(n317), .Q(rd_dat[80]));
Q_FDP4EP \rd_dat_REG[81] ( .CK(clk), .CE(n508), .R(n521), .D(n319), .Q(rd_dat[81]));
Q_FDP4EP \rd_dat_REG[82] ( .CK(clk), .CE(n508), .R(n521), .D(n321), .Q(rd_dat[82]));
Q_FDP4EP \rd_dat_REG[83] ( .CK(clk), .CE(n508), .R(n521), .D(n323), .Q(rd_dat[83]));
Q_FDP4EP \rd_dat_REG[84] ( .CK(clk), .CE(n508), .R(n521), .D(n325), .Q(rd_dat[84]));
Q_FDP4EP \rd_dat_REG[85] ( .CK(clk), .CE(n508), .R(n521), .D(n327), .Q(rd_dat[85]));
Q_FDP4EP \rd_dat_REG[86] ( .CK(clk), .CE(n508), .R(n521), .D(n329), .Q(rd_dat[86]));
Q_FDP4EP \rd_dat_REG[87] ( .CK(clk), .CE(n508), .R(n521), .D(n331), .Q(rd_dat[87]));
Q_FDP4EP \rd_dat_REG[88] ( .CK(clk), .CE(n508), .R(n521), .D(n333), .Q(rd_dat[88]));
Q_FDP4EP \rd_dat_REG[89] ( .CK(clk), .CE(n508), .R(n521), .D(n335), .Q(rd_dat[89]));
Q_FDP4EP \rd_dat_REG[90] ( .CK(clk), .CE(n508), .R(n521), .D(n337), .Q(rd_dat[90]));
Q_FDP4EP \rd_dat_REG[91] ( .CK(clk), .CE(n508), .R(n521), .D(n339), .Q(rd_dat[91]));
Q_FDP4EP \rd_dat_REG[92] ( .CK(clk), .CE(n508), .R(n521), .D(n341), .Q(rd_dat[92]));
Q_FDP4EP \rd_dat_REG[93] ( .CK(clk), .CE(n508), .R(n521), .D(n343), .Q(rd_dat[93]));
Q_FDP4EP \rd_dat_REG[94] ( .CK(clk), .CE(n508), .R(n521), .D(n345), .Q(rd_dat[94]));
Q_FDP4EP \rd_dat_REG[95] ( .CK(clk), .CE(n508), .R(n521), .D(n347), .Q(rd_dat[95]));
Q_INV U807 ( .A(n511), .Z(n522));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n522), .R(n521), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 8 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
