library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity xcva_top is
  attribute _2_state_: integer;
end xcva_top ;
