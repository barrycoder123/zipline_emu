
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_gfifo_port_280_2_0 ( tkout, tkin, ireq, cbid, len, idata, CGFtsReq, 
	CGFcbid, CGFlen, CGFidata, CGFfull, CLBreq, CLBrd, CLBwr, CLBfull, 
	Rtkin);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output tkout;
input tkin;
input ireq;
input [19:0] cbid;
input [11:0] len;
input [279:0] idata;
output CGFtsReq;
output [19:0] CGFcbid;
output [11:0] CGFlen;
output [511:0] CGFidata;
input CGFfull;
output CLBreq;
input [3:0] CLBrd;
input [3:0] CLBwr;
input CLBfull;
input Rtkin;
wire fclk;
wire enq;
wire CLBreqWhileFull;
`_2_ wire en;
`_2_ wire ack;
`_2_ wire [279:0] odata;
`_2_ wire oreq;
`_2_ wire [19:0] ocbid;
`_2_ wire [19:0] xcbid;
`_2_ wire [11:0] olen;
`_2_ wire [11:0] xlen;
`_2_ wire [0:0] sel;
`_2_ wire [279:0] xdata;
wire [31:0] i;
`_2_ wire ireqR;
supply1 n5;
Q_ASSIGN U0 ( .B(len[0]), .A(xlen[0]));
Q_ASSIGN U1 ( .B(len[0]), .A(olen[0]));
Q_ASSIGN U2 ( .B(len[1]), .A(xlen[1]));
Q_ASSIGN U3 ( .B(len[1]), .A(olen[1]));
Q_ASSIGN U4 ( .B(len[2]), .A(xlen[2]));
Q_ASSIGN U5 ( .B(len[2]), .A(olen[2]));
Q_ASSIGN U6 ( .B(len[3]), .A(xlen[3]));
Q_ASSIGN U7 ( .B(len[3]), .A(olen[3]));
Q_ASSIGN U8 ( .B(len[4]), .A(xlen[4]));
Q_ASSIGN U9 ( .B(len[4]), .A(olen[4]));
Q_ASSIGN U10 ( .B(len[5]), .A(xlen[5]));
Q_ASSIGN U11 ( .B(len[5]), .A(olen[5]));
Q_ASSIGN U12 ( .B(len[6]), .A(xlen[6]));
Q_ASSIGN U13 ( .B(len[6]), .A(olen[6]));
Q_ASSIGN U14 ( .B(len[7]), .A(xlen[7]));
Q_ASSIGN U15 ( .B(len[7]), .A(olen[7]));
Q_ASSIGN U16 ( .B(len[8]), .A(xlen[8]));
Q_ASSIGN U17 ( .B(len[8]), .A(olen[8]));
Q_ASSIGN U18 ( .B(len[9]), .A(xlen[9]));
Q_ASSIGN U19 ( .B(len[9]), .A(olen[9]));
Q_ASSIGN U20 ( .B(len[10]), .A(xlen[10]));
Q_ASSIGN U21 ( .B(len[10]), .A(olen[10]));
Q_ASSIGN U22 ( .B(len[11]), .A(xlen[11]));
Q_ASSIGN U23 ( .B(len[11]), .A(olen[11]));
Q_BUF U24 ( .A(ocbid[0]), .Z(xcbid[0]));
Q_BUF U25 ( .A(ocbid[1]), .Z(xcbid[1]));
Q_BUF U26 ( .A(ocbid[2]), .Z(xcbid[2]));
Q_BUF U27 ( .A(ocbid[3]), .Z(xcbid[3]));
Q_BUF U28 ( .A(ocbid[4]), .Z(xcbid[4]));
Q_BUF U29 ( .A(ocbid[5]), .Z(xcbid[5]));
Q_BUF U30 ( .A(ocbid[6]), .Z(xcbid[6]));
Q_BUF U31 ( .A(ocbid[7]), .Z(xcbid[7]));
Q_BUF U32 ( .A(ocbid[8]), .Z(xcbid[8]));
Q_BUF U33 ( .A(ocbid[9]), .Z(xcbid[9]));
Q_BUF U34 ( .A(ocbid[10]), .Z(xcbid[10]));
Q_BUF U35 ( .A(ocbid[11]), .Z(xcbid[11]));
Q_BUF U36 ( .A(ocbid[12]), .Z(xcbid[12]));
Q_BUF U37 ( .A(ocbid[13]), .Z(xcbid[13]));
Q_BUF U38 ( .A(ocbid[14]), .Z(xcbid[14]));
Q_BUF U39 ( .A(ocbid[15]), .Z(xcbid[15]));
Q_BUF U40 ( .A(ocbid[16]), .Z(xcbid[16]));
Q_BUF U41 ( .A(ocbid[17]), .Z(xcbid[17]));
Q_BUF U42 ( .A(ocbid[18]), .Z(xcbid[18]));
Q_BUF U43 ( .A(ocbid[19]), .Z(xcbid[19]));
Q_BUF U44 ( .A(odata[0]), .Z(xdata[0]));
Q_BUF U45 ( .A(odata[1]), .Z(xdata[1]));
Q_BUF U46 ( .A(odata[2]), .Z(xdata[2]));
Q_BUF U47 ( .A(odata[3]), .Z(xdata[3]));
Q_BUF U48 ( .A(odata[4]), .Z(xdata[4]));
Q_BUF U49 ( .A(odata[5]), .Z(xdata[5]));
Q_BUF U50 ( .A(odata[6]), .Z(xdata[6]));
Q_BUF U51 ( .A(odata[7]), .Z(xdata[7]));
Q_BUF U52 ( .A(odata[8]), .Z(xdata[8]));
Q_BUF U53 ( .A(odata[9]), .Z(xdata[9]));
Q_BUF U54 ( .A(odata[10]), .Z(xdata[10]));
Q_BUF U55 ( .A(odata[11]), .Z(xdata[11]));
Q_BUF U56 ( .A(odata[12]), .Z(xdata[12]));
Q_BUF U57 ( .A(odata[13]), .Z(xdata[13]));
Q_BUF U58 ( .A(odata[14]), .Z(xdata[14]));
Q_BUF U59 ( .A(odata[15]), .Z(xdata[15]));
Q_BUF U60 ( .A(odata[16]), .Z(xdata[16]));
Q_BUF U61 ( .A(odata[17]), .Z(xdata[17]));
Q_BUF U62 ( .A(odata[18]), .Z(xdata[18]));
Q_BUF U63 ( .A(odata[19]), .Z(xdata[19]));
Q_BUF U64 ( .A(odata[20]), .Z(xdata[20]));
Q_BUF U65 ( .A(odata[21]), .Z(xdata[21]));
Q_BUF U66 ( .A(odata[22]), .Z(xdata[22]));
Q_BUF U67 ( .A(odata[23]), .Z(xdata[23]));
Q_BUF U68 ( .A(odata[24]), .Z(xdata[24]));
Q_BUF U69 ( .A(odata[25]), .Z(xdata[25]));
Q_BUF U70 ( .A(odata[26]), .Z(xdata[26]));
Q_BUF U71 ( .A(odata[27]), .Z(xdata[27]));
Q_BUF U72 ( .A(odata[28]), .Z(xdata[28]));
Q_BUF U73 ( .A(odata[29]), .Z(xdata[29]));
Q_BUF U74 ( .A(odata[30]), .Z(xdata[30]));
Q_BUF U75 ( .A(odata[31]), .Z(xdata[31]));
Q_BUF U76 ( .A(odata[32]), .Z(xdata[32]));
Q_BUF U77 ( .A(odata[33]), .Z(xdata[33]));
Q_BUF U78 ( .A(odata[34]), .Z(xdata[34]));
Q_BUF U79 ( .A(odata[35]), .Z(xdata[35]));
Q_BUF U80 ( .A(odata[36]), .Z(xdata[36]));
Q_BUF U81 ( .A(odata[37]), .Z(xdata[37]));
Q_BUF U82 ( .A(odata[38]), .Z(xdata[38]));
Q_BUF U83 ( .A(odata[39]), .Z(xdata[39]));
Q_BUF U84 ( .A(odata[40]), .Z(xdata[40]));
Q_BUF U85 ( .A(odata[41]), .Z(xdata[41]));
Q_BUF U86 ( .A(odata[42]), .Z(xdata[42]));
Q_BUF U87 ( .A(odata[43]), .Z(xdata[43]));
Q_BUF U88 ( .A(odata[44]), .Z(xdata[44]));
Q_BUF U89 ( .A(odata[45]), .Z(xdata[45]));
Q_BUF U90 ( .A(odata[46]), .Z(xdata[46]));
Q_BUF U91 ( .A(odata[47]), .Z(xdata[47]));
Q_BUF U92 ( .A(odata[48]), .Z(xdata[48]));
Q_BUF U93 ( .A(odata[49]), .Z(xdata[49]));
Q_BUF U94 ( .A(odata[50]), .Z(xdata[50]));
Q_BUF U95 ( .A(odata[51]), .Z(xdata[51]));
Q_BUF U96 ( .A(odata[52]), .Z(xdata[52]));
Q_BUF U97 ( .A(odata[53]), .Z(xdata[53]));
Q_BUF U98 ( .A(odata[54]), .Z(xdata[54]));
Q_BUF U99 ( .A(odata[55]), .Z(xdata[55]));
Q_BUF U100 ( .A(odata[56]), .Z(xdata[56]));
Q_BUF U101 ( .A(odata[57]), .Z(xdata[57]));
Q_BUF U102 ( .A(odata[58]), .Z(xdata[58]));
Q_BUF U103 ( .A(odata[59]), .Z(xdata[59]));
Q_BUF U104 ( .A(odata[60]), .Z(xdata[60]));
Q_BUF U105 ( .A(odata[61]), .Z(xdata[61]));
Q_BUF U106 ( .A(odata[62]), .Z(xdata[62]));
Q_BUF U107 ( .A(odata[63]), .Z(xdata[63]));
Q_BUF U108 ( .A(odata[64]), .Z(xdata[64]));
Q_BUF U109 ( .A(odata[65]), .Z(xdata[65]));
Q_BUF U110 ( .A(odata[66]), .Z(xdata[66]));
Q_BUF U111 ( .A(odata[67]), .Z(xdata[67]));
Q_BUF U112 ( .A(odata[68]), .Z(xdata[68]));
Q_BUF U113 ( .A(odata[69]), .Z(xdata[69]));
Q_BUF U114 ( .A(odata[70]), .Z(xdata[70]));
Q_BUF U115 ( .A(odata[71]), .Z(xdata[71]));
Q_BUF U116 ( .A(odata[72]), .Z(xdata[72]));
Q_BUF U117 ( .A(odata[73]), .Z(xdata[73]));
Q_BUF U118 ( .A(odata[74]), .Z(xdata[74]));
Q_BUF U119 ( .A(odata[75]), .Z(xdata[75]));
Q_BUF U120 ( .A(odata[76]), .Z(xdata[76]));
Q_BUF U121 ( .A(odata[77]), .Z(xdata[77]));
Q_BUF U122 ( .A(odata[78]), .Z(xdata[78]));
Q_BUF U123 ( .A(odata[79]), .Z(xdata[79]));
Q_BUF U124 ( .A(odata[80]), .Z(xdata[80]));
Q_BUF U125 ( .A(odata[81]), .Z(xdata[81]));
Q_BUF U126 ( .A(odata[82]), .Z(xdata[82]));
Q_BUF U127 ( .A(odata[83]), .Z(xdata[83]));
Q_BUF U128 ( .A(odata[84]), .Z(xdata[84]));
Q_BUF U129 ( .A(odata[85]), .Z(xdata[85]));
Q_BUF U130 ( .A(odata[86]), .Z(xdata[86]));
Q_BUF U131 ( .A(odata[87]), .Z(xdata[87]));
Q_BUF U132 ( .A(odata[88]), .Z(xdata[88]));
Q_BUF U133 ( .A(odata[89]), .Z(xdata[89]));
Q_BUF U134 ( .A(odata[90]), .Z(xdata[90]));
Q_BUF U135 ( .A(odata[91]), .Z(xdata[91]));
Q_BUF U136 ( .A(odata[92]), .Z(xdata[92]));
Q_BUF U137 ( .A(odata[93]), .Z(xdata[93]));
Q_BUF U138 ( .A(odata[94]), .Z(xdata[94]));
Q_BUF U139 ( .A(odata[95]), .Z(xdata[95]));
Q_BUF U140 ( .A(odata[96]), .Z(xdata[96]));
Q_BUF U141 ( .A(odata[97]), .Z(xdata[97]));
Q_BUF U142 ( .A(odata[98]), .Z(xdata[98]));
Q_BUF U143 ( .A(odata[99]), .Z(xdata[99]));
Q_BUF U144 ( .A(odata[100]), .Z(xdata[100]));
Q_BUF U145 ( .A(odata[101]), .Z(xdata[101]));
Q_BUF U146 ( .A(odata[102]), .Z(xdata[102]));
Q_BUF U147 ( .A(odata[103]), .Z(xdata[103]));
Q_BUF U148 ( .A(odata[104]), .Z(xdata[104]));
Q_BUF U149 ( .A(odata[105]), .Z(xdata[105]));
Q_BUF U150 ( .A(odata[106]), .Z(xdata[106]));
Q_BUF U151 ( .A(odata[107]), .Z(xdata[107]));
Q_BUF U152 ( .A(odata[108]), .Z(xdata[108]));
Q_BUF U153 ( .A(odata[109]), .Z(xdata[109]));
Q_BUF U154 ( .A(odata[110]), .Z(xdata[110]));
Q_BUF U155 ( .A(odata[111]), .Z(xdata[111]));
Q_BUF U156 ( .A(odata[112]), .Z(xdata[112]));
Q_BUF U157 ( .A(odata[113]), .Z(xdata[113]));
Q_BUF U158 ( .A(odata[114]), .Z(xdata[114]));
Q_BUF U159 ( .A(odata[115]), .Z(xdata[115]));
Q_BUF U160 ( .A(odata[116]), .Z(xdata[116]));
Q_BUF U161 ( .A(odata[117]), .Z(xdata[117]));
Q_BUF U162 ( .A(odata[118]), .Z(xdata[118]));
Q_BUF U163 ( .A(odata[119]), .Z(xdata[119]));
Q_BUF U164 ( .A(odata[120]), .Z(xdata[120]));
Q_BUF U165 ( .A(odata[121]), .Z(xdata[121]));
Q_BUF U166 ( .A(odata[122]), .Z(xdata[122]));
Q_BUF U167 ( .A(odata[123]), .Z(xdata[123]));
Q_BUF U168 ( .A(odata[124]), .Z(xdata[124]));
Q_BUF U169 ( .A(odata[125]), .Z(xdata[125]));
Q_BUF U170 ( .A(odata[126]), .Z(xdata[126]));
Q_BUF U171 ( .A(odata[127]), .Z(xdata[127]));
Q_BUF U172 ( .A(odata[128]), .Z(xdata[128]));
Q_BUF U173 ( .A(odata[129]), .Z(xdata[129]));
Q_BUF U174 ( .A(odata[130]), .Z(xdata[130]));
Q_BUF U175 ( .A(odata[131]), .Z(xdata[131]));
Q_BUF U176 ( .A(odata[132]), .Z(xdata[132]));
Q_BUF U177 ( .A(odata[133]), .Z(xdata[133]));
Q_BUF U178 ( .A(odata[134]), .Z(xdata[134]));
Q_BUF U179 ( .A(odata[135]), .Z(xdata[135]));
Q_BUF U180 ( .A(odata[136]), .Z(xdata[136]));
Q_BUF U181 ( .A(odata[137]), .Z(xdata[137]));
Q_BUF U182 ( .A(odata[138]), .Z(xdata[138]));
Q_BUF U183 ( .A(odata[139]), .Z(xdata[139]));
Q_BUF U184 ( .A(odata[140]), .Z(xdata[140]));
Q_BUF U185 ( .A(odata[141]), .Z(xdata[141]));
Q_BUF U186 ( .A(odata[142]), .Z(xdata[142]));
Q_BUF U187 ( .A(odata[143]), .Z(xdata[143]));
Q_BUF U188 ( .A(odata[144]), .Z(xdata[144]));
Q_BUF U189 ( .A(odata[145]), .Z(xdata[145]));
Q_BUF U190 ( .A(odata[146]), .Z(xdata[146]));
Q_BUF U191 ( .A(odata[147]), .Z(xdata[147]));
Q_BUF U192 ( .A(odata[148]), .Z(xdata[148]));
Q_BUF U193 ( .A(odata[149]), .Z(xdata[149]));
Q_BUF U194 ( .A(odata[150]), .Z(xdata[150]));
Q_BUF U195 ( .A(odata[151]), .Z(xdata[151]));
Q_BUF U196 ( .A(odata[152]), .Z(xdata[152]));
Q_BUF U197 ( .A(odata[153]), .Z(xdata[153]));
Q_BUF U198 ( .A(odata[154]), .Z(xdata[154]));
Q_BUF U199 ( .A(odata[155]), .Z(xdata[155]));
Q_BUF U200 ( .A(odata[156]), .Z(xdata[156]));
Q_BUF U201 ( .A(odata[157]), .Z(xdata[157]));
Q_BUF U202 ( .A(odata[158]), .Z(xdata[158]));
Q_BUF U203 ( .A(odata[159]), .Z(xdata[159]));
Q_BUF U204 ( .A(odata[160]), .Z(xdata[160]));
Q_BUF U205 ( .A(odata[161]), .Z(xdata[161]));
Q_BUF U206 ( .A(odata[162]), .Z(xdata[162]));
Q_BUF U207 ( .A(odata[163]), .Z(xdata[163]));
Q_BUF U208 ( .A(odata[164]), .Z(xdata[164]));
Q_BUF U209 ( .A(odata[165]), .Z(xdata[165]));
Q_BUF U210 ( .A(odata[166]), .Z(xdata[166]));
Q_BUF U211 ( .A(odata[167]), .Z(xdata[167]));
Q_BUF U212 ( .A(odata[168]), .Z(xdata[168]));
Q_BUF U213 ( .A(odata[169]), .Z(xdata[169]));
Q_BUF U214 ( .A(odata[170]), .Z(xdata[170]));
Q_BUF U215 ( .A(odata[171]), .Z(xdata[171]));
Q_BUF U216 ( .A(odata[172]), .Z(xdata[172]));
Q_BUF U217 ( .A(odata[173]), .Z(xdata[173]));
Q_BUF U218 ( .A(odata[174]), .Z(xdata[174]));
Q_BUF U219 ( .A(odata[175]), .Z(xdata[175]));
Q_BUF U220 ( .A(odata[176]), .Z(xdata[176]));
Q_BUF U221 ( .A(odata[177]), .Z(xdata[177]));
Q_BUF U222 ( .A(odata[178]), .Z(xdata[178]));
Q_BUF U223 ( .A(odata[179]), .Z(xdata[179]));
Q_BUF U224 ( .A(odata[180]), .Z(xdata[180]));
Q_BUF U225 ( .A(odata[181]), .Z(xdata[181]));
Q_BUF U226 ( .A(odata[182]), .Z(xdata[182]));
Q_BUF U227 ( .A(odata[183]), .Z(xdata[183]));
Q_BUF U228 ( .A(odata[184]), .Z(xdata[184]));
Q_BUF U229 ( .A(odata[185]), .Z(xdata[185]));
Q_BUF U230 ( .A(odata[186]), .Z(xdata[186]));
Q_BUF U231 ( .A(odata[187]), .Z(xdata[187]));
Q_BUF U232 ( .A(odata[188]), .Z(xdata[188]));
Q_BUF U233 ( .A(odata[189]), .Z(xdata[189]));
Q_BUF U234 ( .A(odata[190]), .Z(xdata[190]));
Q_BUF U235 ( .A(odata[191]), .Z(xdata[191]));
Q_BUF U236 ( .A(odata[192]), .Z(xdata[192]));
Q_BUF U237 ( .A(odata[193]), .Z(xdata[193]));
Q_BUF U238 ( .A(odata[194]), .Z(xdata[194]));
Q_BUF U239 ( .A(odata[195]), .Z(xdata[195]));
Q_BUF U240 ( .A(odata[196]), .Z(xdata[196]));
Q_BUF U241 ( .A(odata[197]), .Z(xdata[197]));
Q_BUF U242 ( .A(odata[198]), .Z(xdata[198]));
Q_BUF U243 ( .A(odata[199]), .Z(xdata[199]));
Q_BUF U244 ( .A(odata[200]), .Z(xdata[200]));
Q_BUF U245 ( .A(odata[201]), .Z(xdata[201]));
Q_BUF U246 ( .A(odata[202]), .Z(xdata[202]));
Q_BUF U247 ( .A(odata[203]), .Z(xdata[203]));
Q_BUF U248 ( .A(odata[204]), .Z(xdata[204]));
Q_BUF U249 ( .A(odata[205]), .Z(xdata[205]));
Q_BUF U250 ( .A(odata[206]), .Z(xdata[206]));
Q_BUF U251 ( .A(odata[207]), .Z(xdata[207]));
Q_BUF U252 ( .A(odata[208]), .Z(xdata[208]));
Q_BUF U253 ( .A(odata[209]), .Z(xdata[209]));
Q_BUF U254 ( .A(odata[210]), .Z(xdata[210]));
Q_BUF U255 ( .A(odata[211]), .Z(xdata[211]));
Q_BUF U256 ( .A(odata[212]), .Z(xdata[212]));
Q_BUF U257 ( .A(odata[213]), .Z(xdata[213]));
Q_BUF U258 ( .A(odata[214]), .Z(xdata[214]));
Q_BUF U259 ( .A(odata[215]), .Z(xdata[215]));
Q_BUF U260 ( .A(odata[216]), .Z(xdata[216]));
Q_BUF U261 ( .A(odata[217]), .Z(xdata[217]));
Q_BUF U262 ( .A(odata[218]), .Z(xdata[218]));
Q_BUF U263 ( .A(odata[219]), .Z(xdata[219]));
Q_BUF U264 ( .A(odata[220]), .Z(xdata[220]));
Q_BUF U265 ( .A(odata[221]), .Z(xdata[221]));
Q_BUF U266 ( .A(odata[222]), .Z(xdata[222]));
Q_BUF U267 ( .A(odata[223]), .Z(xdata[223]));
Q_BUF U268 ( .A(odata[224]), .Z(xdata[224]));
Q_BUF U269 ( .A(odata[225]), .Z(xdata[225]));
Q_BUF U270 ( .A(odata[226]), .Z(xdata[226]));
Q_BUF U271 ( .A(odata[227]), .Z(xdata[227]));
Q_BUF U272 ( .A(odata[228]), .Z(xdata[228]));
Q_BUF U273 ( .A(odata[229]), .Z(xdata[229]));
Q_BUF U274 ( .A(odata[230]), .Z(xdata[230]));
Q_BUF U275 ( .A(odata[231]), .Z(xdata[231]));
Q_BUF U276 ( .A(odata[232]), .Z(xdata[232]));
Q_BUF U277 ( .A(odata[233]), .Z(xdata[233]));
Q_BUF U278 ( .A(odata[234]), .Z(xdata[234]));
Q_BUF U279 ( .A(odata[235]), .Z(xdata[235]));
Q_BUF U280 ( .A(odata[236]), .Z(xdata[236]));
Q_BUF U281 ( .A(odata[237]), .Z(xdata[237]));
Q_BUF U282 ( .A(odata[238]), .Z(xdata[238]));
Q_BUF U283 ( .A(odata[239]), .Z(xdata[239]));
Q_BUF U284 ( .A(odata[240]), .Z(xdata[240]));
Q_BUF U285 ( .A(odata[241]), .Z(xdata[241]));
Q_BUF U286 ( .A(odata[242]), .Z(xdata[242]));
Q_BUF U287 ( .A(odata[243]), .Z(xdata[243]));
Q_BUF U288 ( .A(odata[244]), .Z(xdata[244]));
Q_BUF U289 ( .A(odata[245]), .Z(xdata[245]));
Q_BUF U290 ( .A(odata[246]), .Z(xdata[246]));
Q_BUF U291 ( .A(odata[247]), .Z(xdata[247]));
Q_BUF U292 ( .A(odata[248]), .Z(xdata[248]));
Q_BUF U293 ( .A(odata[249]), .Z(xdata[249]));
Q_BUF U294 ( .A(odata[250]), .Z(xdata[250]));
Q_BUF U295 ( .A(odata[251]), .Z(xdata[251]));
Q_BUF U296 ( .A(odata[252]), .Z(xdata[252]));
Q_BUF U297 ( .A(odata[253]), .Z(xdata[253]));
Q_BUF U298 ( .A(odata[254]), .Z(xdata[254]));
Q_BUF U299 ( .A(odata[255]), .Z(xdata[255]));
Q_BUF U300 ( .A(odata[256]), .Z(xdata[256]));
Q_BUF U301 ( .A(odata[257]), .Z(xdata[257]));
Q_BUF U302 ( .A(odata[258]), .Z(xdata[258]));
Q_BUF U303 ( .A(odata[259]), .Z(xdata[259]));
Q_BUF U304 ( .A(odata[260]), .Z(xdata[260]));
Q_BUF U305 ( .A(odata[261]), .Z(xdata[261]));
Q_BUF U306 ( .A(odata[262]), .Z(xdata[262]));
Q_BUF U307 ( .A(odata[263]), .Z(xdata[263]));
Q_BUF U308 ( .A(odata[264]), .Z(xdata[264]));
Q_BUF U309 ( .A(odata[265]), .Z(xdata[265]));
Q_BUF U310 ( .A(odata[266]), .Z(xdata[266]));
Q_BUF U311 ( .A(odata[267]), .Z(xdata[267]));
Q_BUF U312 ( .A(odata[268]), .Z(xdata[268]));
Q_BUF U313 ( .A(odata[269]), .Z(xdata[269]));
Q_BUF U314 ( .A(odata[270]), .Z(xdata[270]));
Q_BUF U315 ( .A(odata[271]), .Z(xdata[271]));
Q_BUF U316 ( .A(odata[272]), .Z(xdata[272]));
Q_BUF U317 ( .A(odata[273]), .Z(xdata[273]));
Q_BUF U318 ( .A(odata[274]), .Z(xdata[274]));
Q_BUF U319 ( .A(odata[275]), .Z(xdata[275]));
Q_BUF U320 ( .A(odata[276]), .Z(xdata[276]));
Q_BUF U321 ( .A(odata[277]), .Z(xdata[277]));
Q_BUF U322 ( .A(odata[278]), .Z(xdata[278]));
Q_BUF U323 ( .A(odata[279]), .Z(xdata[279]));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_EV_WOR_START qi ( .A(CLBreqWhileFull));
Q_INV U326 ( .A(n4), .Z(tkout));
Q_XNR2 U327 ( .A0(oreq), .A1(ack), .Z(n4));
Q_CCLKCHK cchk ( .sig(ireq));
Q_AN02 U329 ( .A0(enq), .A1(CLBfull), .Z(CLBreqWhileFull));
Q_AN02 U330 ( .A0(n2), .A1(n3), .Z(enq));
Q_INV U331 ( .A(xc_top.GFLock2), .Z(n3));
Q_XOR2 U332 ( .A0(ireq), .A1(ireqR), .Z(n2));
Q_BUFZP U333 ( .OE(CLBreqWhileFull), .A(n5), .Z(xc_top.GFLBfull));
Q_BUFZP U334 ( .OE(en), .A(xcbid[0]), .Z(CGFcbid[0]));
Q_BUFZP U335 ( .OE(en), .A(xcbid[1]), .Z(CGFcbid[1]));
Q_BUFZP U336 ( .OE(en), .A(xcbid[2]), .Z(CGFcbid[2]));
Q_BUFZP U337 ( .OE(en), .A(xcbid[3]), .Z(CGFcbid[3]));
Q_BUFZP U338 ( .OE(en), .A(xcbid[4]), .Z(CGFcbid[4]));
Q_BUFZP U339 ( .OE(en), .A(xcbid[5]), .Z(CGFcbid[5]));
Q_BUFZP U340 ( .OE(en), .A(xcbid[6]), .Z(CGFcbid[6]));
Q_BUFZP U341 ( .OE(en), .A(xcbid[7]), .Z(CGFcbid[7]));
Q_BUFZP U342 ( .OE(en), .A(xcbid[8]), .Z(CGFcbid[8]));
Q_BUFZP U343 ( .OE(en), .A(xcbid[9]), .Z(CGFcbid[9]));
Q_BUFZP U344 ( .OE(en), .A(xcbid[10]), .Z(CGFcbid[10]));
Q_BUFZP U345 ( .OE(en), .A(xcbid[11]), .Z(CGFcbid[11]));
Q_BUFZP U346 ( .OE(en), .A(xcbid[12]), .Z(CGFcbid[12]));
Q_BUFZP U347 ( .OE(en), .A(xcbid[13]), .Z(CGFcbid[13]));
Q_BUFZP U348 ( .OE(en), .A(xcbid[14]), .Z(CGFcbid[14]));
Q_BUFZP U349 ( .OE(en), .A(xcbid[15]), .Z(CGFcbid[15]));
Q_BUFZP U350 ( .OE(en), .A(xcbid[16]), .Z(CGFcbid[16]));
Q_BUFZP U351 ( .OE(en), .A(xcbid[17]), .Z(CGFcbid[17]));
Q_BUFZP U352 ( .OE(en), .A(xcbid[18]), .Z(CGFcbid[18]));
Q_BUFZP U353 ( .OE(en), .A(xcbid[19]), .Z(CGFcbid[19]));
Q_BUFZP U354 ( .OE(en), .A(len[0]), .Z(CGFlen[0]));
Q_BUFZP U355 ( .OE(en), .A(len[1]), .Z(CGFlen[1]));
Q_BUFZP U356 ( .OE(en), .A(len[2]), .Z(CGFlen[2]));
Q_BUFZP U357 ( .OE(en), .A(len[3]), .Z(CGFlen[3]));
Q_BUFZP U358 ( .OE(en), .A(len[4]), .Z(CGFlen[4]));
Q_BUFZP U359 ( .OE(en), .A(len[5]), .Z(CGFlen[5]));
Q_BUFZP U360 ( .OE(en), .A(len[6]), .Z(CGFlen[6]));
Q_BUFZP U361 ( .OE(en), .A(len[7]), .Z(CGFlen[7]));
Q_BUFZP U362 ( .OE(en), .A(len[8]), .Z(CGFlen[8]));
Q_BUFZP U363 ( .OE(en), .A(len[9]), .Z(CGFlen[9]));
Q_BUFZP U364 ( .OE(en), .A(len[10]), .Z(CGFlen[10]));
Q_BUFZP U365 ( .OE(en), .A(len[11]), .Z(CGFlen[11]));
Q_BUFZP U366 ( .OE(en), .A(xdata[0]), .Z(CGFidata[0]));
Q_BUFZP U367 ( .OE(en), .A(xdata[1]), .Z(CGFidata[1]));
Q_BUFZP U368 ( .OE(en), .A(xdata[2]), .Z(CGFidata[2]));
Q_BUFZP U369 ( .OE(en), .A(xdata[3]), .Z(CGFidata[3]));
Q_BUFZP U370 ( .OE(en), .A(xdata[4]), .Z(CGFidata[4]));
Q_BUFZP U371 ( .OE(en), .A(xdata[5]), .Z(CGFidata[5]));
Q_BUFZP U372 ( .OE(en), .A(xdata[6]), .Z(CGFidata[6]));
Q_BUFZP U373 ( .OE(en), .A(xdata[7]), .Z(CGFidata[7]));
Q_BUFZP U374 ( .OE(en), .A(xdata[8]), .Z(CGFidata[8]));
Q_BUFZP U375 ( .OE(en), .A(xdata[9]), .Z(CGFidata[9]));
Q_BUFZP U376 ( .OE(en), .A(xdata[10]), .Z(CGFidata[10]));
Q_BUFZP U377 ( .OE(en), .A(xdata[11]), .Z(CGFidata[11]));
Q_BUFZP U378 ( .OE(en), .A(xdata[12]), .Z(CGFidata[12]));
Q_BUFZP U379 ( .OE(en), .A(xdata[13]), .Z(CGFidata[13]));
Q_BUFZP U380 ( .OE(en), .A(xdata[14]), .Z(CGFidata[14]));
Q_BUFZP U381 ( .OE(en), .A(xdata[15]), .Z(CGFidata[15]));
Q_BUFZP U382 ( .OE(en), .A(xdata[16]), .Z(CGFidata[16]));
Q_BUFZP U383 ( .OE(en), .A(xdata[17]), .Z(CGFidata[17]));
Q_BUFZP U384 ( .OE(en), .A(xdata[18]), .Z(CGFidata[18]));
Q_BUFZP U385 ( .OE(en), .A(xdata[19]), .Z(CGFidata[19]));
Q_BUFZP U386 ( .OE(en), .A(xdata[20]), .Z(CGFidata[20]));
Q_BUFZP U387 ( .OE(en), .A(xdata[21]), .Z(CGFidata[21]));
Q_BUFZP U388 ( .OE(en), .A(xdata[22]), .Z(CGFidata[22]));
Q_BUFZP U389 ( .OE(en), .A(xdata[23]), .Z(CGFidata[23]));
Q_BUFZP U390 ( .OE(en), .A(xdata[24]), .Z(CGFidata[24]));
Q_BUFZP U391 ( .OE(en), .A(xdata[25]), .Z(CGFidata[25]));
Q_BUFZP U392 ( .OE(en), .A(xdata[26]), .Z(CGFidata[26]));
Q_BUFZP U393 ( .OE(en), .A(xdata[27]), .Z(CGFidata[27]));
Q_BUFZP U394 ( .OE(en), .A(xdata[28]), .Z(CGFidata[28]));
Q_BUFZP U395 ( .OE(en), .A(xdata[29]), .Z(CGFidata[29]));
Q_BUFZP U396 ( .OE(en), .A(xdata[30]), .Z(CGFidata[30]));
Q_BUFZP U397 ( .OE(en), .A(xdata[31]), .Z(CGFidata[31]));
Q_BUFZP U398 ( .OE(en), .A(xdata[32]), .Z(CGFidata[32]));
Q_BUFZP U399 ( .OE(en), .A(xdata[33]), .Z(CGFidata[33]));
Q_BUFZP U400 ( .OE(en), .A(xdata[34]), .Z(CGFidata[34]));
Q_BUFZP U401 ( .OE(en), .A(xdata[35]), .Z(CGFidata[35]));
Q_BUFZP U402 ( .OE(en), .A(xdata[36]), .Z(CGFidata[36]));
Q_BUFZP U403 ( .OE(en), .A(xdata[37]), .Z(CGFidata[37]));
Q_BUFZP U404 ( .OE(en), .A(xdata[38]), .Z(CGFidata[38]));
Q_BUFZP U405 ( .OE(en), .A(xdata[39]), .Z(CGFidata[39]));
Q_BUFZP U406 ( .OE(en), .A(xdata[40]), .Z(CGFidata[40]));
Q_BUFZP U407 ( .OE(en), .A(xdata[41]), .Z(CGFidata[41]));
Q_BUFZP U408 ( .OE(en), .A(xdata[42]), .Z(CGFidata[42]));
Q_BUFZP U409 ( .OE(en), .A(xdata[43]), .Z(CGFidata[43]));
Q_BUFZP U410 ( .OE(en), .A(xdata[44]), .Z(CGFidata[44]));
Q_BUFZP U411 ( .OE(en), .A(xdata[45]), .Z(CGFidata[45]));
Q_BUFZP U412 ( .OE(en), .A(xdata[46]), .Z(CGFidata[46]));
Q_BUFZP U413 ( .OE(en), .A(xdata[47]), .Z(CGFidata[47]));
Q_BUFZP U414 ( .OE(en), .A(xdata[48]), .Z(CGFidata[48]));
Q_BUFZP U415 ( .OE(en), .A(xdata[49]), .Z(CGFidata[49]));
Q_BUFZP U416 ( .OE(en), .A(xdata[50]), .Z(CGFidata[50]));
Q_BUFZP U417 ( .OE(en), .A(xdata[51]), .Z(CGFidata[51]));
Q_BUFZP U418 ( .OE(en), .A(xdata[52]), .Z(CGFidata[52]));
Q_BUFZP U419 ( .OE(en), .A(xdata[53]), .Z(CGFidata[53]));
Q_BUFZP U420 ( .OE(en), .A(xdata[54]), .Z(CGFidata[54]));
Q_BUFZP U421 ( .OE(en), .A(xdata[55]), .Z(CGFidata[55]));
Q_BUFZP U422 ( .OE(en), .A(xdata[56]), .Z(CGFidata[56]));
Q_BUFZP U423 ( .OE(en), .A(xdata[57]), .Z(CGFidata[57]));
Q_BUFZP U424 ( .OE(en), .A(xdata[58]), .Z(CGFidata[58]));
Q_BUFZP U425 ( .OE(en), .A(xdata[59]), .Z(CGFidata[59]));
Q_BUFZP U426 ( .OE(en), .A(xdata[60]), .Z(CGFidata[60]));
Q_BUFZP U427 ( .OE(en), .A(xdata[61]), .Z(CGFidata[61]));
Q_BUFZP U428 ( .OE(en), .A(xdata[62]), .Z(CGFidata[62]));
Q_BUFZP U429 ( .OE(en), .A(xdata[63]), .Z(CGFidata[63]));
Q_BUFZP U430 ( .OE(en), .A(xdata[64]), .Z(CGFidata[64]));
Q_BUFZP U431 ( .OE(en), .A(xdata[65]), .Z(CGFidata[65]));
Q_BUFZP U432 ( .OE(en), .A(xdata[66]), .Z(CGFidata[66]));
Q_BUFZP U433 ( .OE(en), .A(xdata[67]), .Z(CGFidata[67]));
Q_BUFZP U434 ( .OE(en), .A(xdata[68]), .Z(CGFidata[68]));
Q_BUFZP U435 ( .OE(en), .A(xdata[69]), .Z(CGFidata[69]));
Q_BUFZP U436 ( .OE(en), .A(xdata[70]), .Z(CGFidata[70]));
Q_BUFZP U437 ( .OE(en), .A(xdata[71]), .Z(CGFidata[71]));
Q_BUFZP U438 ( .OE(en), .A(xdata[72]), .Z(CGFidata[72]));
Q_BUFZP U439 ( .OE(en), .A(xdata[73]), .Z(CGFidata[73]));
Q_BUFZP U440 ( .OE(en), .A(xdata[74]), .Z(CGFidata[74]));
Q_BUFZP U441 ( .OE(en), .A(xdata[75]), .Z(CGFidata[75]));
Q_BUFZP U442 ( .OE(en), .A(xdata[76]), .Z(CGFidata[76]));
Q_BUFZP U443 ( .OE(en), .A(xdata[77]), .Z(CGFidata[77]));
Q_BUFZP U444 ( .OE(en), .A(xdata[78]), .Z(CGFidata[78]));
Q_BUFZP U445 ( .OE(en), .A(xdata[79]), .Z(CGFidata[79]));
Q_BUFZP U446 ( .OE(en), .A(xdata[80]), .Z(CGFidata[80]));
Q_BUFZP U447 ( .OE(en), .A(xdata[81]), .Z(CGFidata[81]));
Q_BUFZP U448 ( .OE(en), .A(xdata[82]), .Z(CGFidata[82]));
Q_BUFZP U449 ( .OE(en), .A(xdata[83]), .Z(CGFidata[83]));
Q_BUFZP U450 ( .OE(en), .A(xdata[84]), .Z(CGFidata[84]));
Q_BUFZP U451 ( .OE(en), .A(xdata[85]), .Z(CGFidata[85]));
Q_BUFZP U452 ( .OE(en), .A(xdata[86]), .Z(CGFidata[86]));
Q_BUFZP U453 ( .OE(en), .A(xdata[87]), .Z(CGFidata[87]));
Q_BUFZP U454 ( .OE(en), .A(xdata[88]), .Z(CGFidata[88]));
Q_BUFZP U455 ( .OE(en), .A(xdata[89]), .Z(CGFidata[89]));
Q_BUFZP U456 ( .OE(en), .A(xdata[90]), .Z(CGFidata[90]));
Q_BUFZP U457 ( .OE(en), .A(xdata[91]), .Z(CGFidata[91]));
Q_BUFZP U458 ( .OE(en), .A(xdata[92]), .Z(CGFidata[92]));
Q_BUFZP U459 ( .OE(en), .A(xdata[93]), .Z(CGFidata[93]));
Q_BUFZP U460 ( .OE(en), .A(xdata[94]), .Z(CGFidata[94]));
Q_BUFZP U461 ( .OE(en), .A(xdata[95]), .Z(CGFidata[95]));
Q_BUFZP U462 ( .OE(en), .A(xdata[96]), .Z(CGFidata[96]));
Q_BUFZP U463 ( .OE(en), .A(xdata[97]), .Z(CGFidata[97]));
Q_BUFZP U464 ( .OE(en), .A(xdata[98]), .Z(CGFidata[98]));
Q_BUFZP U465 ( .OE(en), .A(xdata[99]), .Z(CGFidata[99]));
Q_BUFZP U466 ( .OE(en), .A(xdata[100]), .Z(CGFidata[100]));
Q_BUFZP U467 ( .OE(en), .A(xdata[101]), .Z(CGFidata[101]));
Q_BUFZP U468 ( .OE(en), .A(xdata[102]), .Z(CGFidata[102]));
Q_BUFZP U469 ( .OE(en), .A(xdata[103]), .Z(CGFidata[103]));
Q_BUFZP U470 ( .OE(en), .A(xdata[104]), .Z(CGFidata[104]));
Q_BUFZP U471 ( .OE(en), .A(xdata[105]), .Z(CGFidata[105]));
Q_BUFZP U472 ( .OE(en), .A(xdata[106]), .Z(CGFidata[106]));
Q_BUFZP U473 ( .OE(en), .A(xdata[107]), .Z(CGFidata[107]));
Q_BUFZP U474 ( .OE(en), .A(xdata[108]), .Z(CGFidata[108]));
Q_BUFZP U475 ( .OE(en), .A(xdata[109]), .Z(CGFidata[109]));
Q_BUFZP U476 ( .OE(en), .A(xdata[110]), .Z(CGFidata[110]));
Q_BUFZP U477 ( .OE(en), .A(xdata[111]), .Z(CGFidata[111]));
Q_BUFZP U478 ( .OE(en), .A(xdata[112]), .Z(CGFidata[112]));
Q_BUFZP U479 ( .OE(en), .A(xdata[113]), .Z(CGFidata[113]));
Q_BUFZP U480 ( .OE(en), .A(xdata[114]), .Z(CGFidata[114]));
Q_BUFZP U481 ( .OE(en), .A(xdata[115]), .Z(CGFidata[115]));
Q_BUFZP U482 ( .OE(en), .A(xdata[116]), .Z(CGFidata[116]));
Q_BUFZP U483 ( .OE(en), .A(xdata[117]), .Z(CGFidata[117]));
Q_BUFZP U484 ( .OE(en), .A(xdata[118]), .Z(CGFidata[118]));
Q_BUFZP U485 ( .OE(en), .A(xdata[119]), .Z(CGFidata[119]));
Q_BUFZP U486 ( .OE(en), .A(xdata[120]), .Z(CGFidata[120]));
Q_BUFZP U487 ( .OE(en), .A(xdata[121]), .Z(CGFidata[121]));
Q_BUFZP U488 ( .OE(en), .A(xdata[122]), .Z(CGFidata[122]));
Q_BUFZP U489 ( .OE(en), .A(xdata[123]), .Z(CGFidata[123]));
Q_BUFZP U490 ( .OE(en), .A(xdata[124]), .Z(CGFidata[124]));
Q_BUFZP U491 ( .OE(en), .A(xdata[125]), .Z(CGFidata[125]));
Q_BUFZP U492 ( .OE(en), .A(xdata[126]), .Z(CGFidata[126]));
Q_BUFZP U493 ( .OE(en), .A(xdata[127]), .Z(CGFidata[127]));
Q_BUFZP U494 ( .OE(en), .A(xdata[128]), .Z(CGFidata[128]));
Q_BUFZP U495 ( .OE(en), .A(xdata[129]), .Z(CGFidata[129]));
Q_BUFZP U496 ( .OE(en), .A(xdata[130]), .Z(CGFidata[130]));
Q_BUFZP U497 ( .OE(en), .A(xdata[131]), .Z(CGFidata[131]));
Q_BUFZP U498 ( .OE(en), .A(xdata[132]), .Z(CGFidata[132]));
Q_BUFZP U499 ( .OE(en), .A(xdata[133]), .Z(CGFidata[133]));
Q_BUFZP U500 ( .OE(en), .A(xdata[134]), .Z(CGFidata[134]));
Q_BUFZP U501 ( .OE(en), .A(xdata[135]), .Z(CGFidata[135]));
Q_BUFZP U502 ( .OE(en), .A(xdata[136]), .Z(CGFidata[136]));
Q_BUFZP U503 ( .OE(en), .A(xdata[137]), .Z(CGFidata[137]));
Q_BUFZP U504 ( .OE(en), .A(xdata[138]), .Z(CGFidata[138]));
Q_BUFZP U505 ( .OE(en), .A(xdata[139]), .Z(CGFidata[139]));
Q_BUFZP U506 ( .OE(en), .A(xdata[140]), .Z(CGFidata[140]));
Q_BUFZP U507 ( .OE(en), .A(xdata[141]), .Z(CGFidata[141]));
Q_BUFZP U508 ( .OE(en), .A(xdata[142]), .Z(CGFidata[142]));
Q_BUFZP U509 ( .OE(en), .A(xdata[143]), .Z(CGFidata[143]));
Q_BUFZP U510 ( .OE(en), .A(xdata[144]), .Z(CGFidata[144]));
Q_BUFZP U511 ( .OE(en), .A(xdata[145]), .Z(CGFidata[145]));
Q_BUFZP U512 ( .OE(en), .A(xdata[146]), .Z(CGFidata[146]));
Q_BUFZP U513 ( .OE(en), .A(xdata[147]), .Z(CGFidata[147]));
Q_BUFZP U514 ( .OE(en), .A(xdata[148]), .Z(CGFidata[148]));
Q_BUFZP U515 ( .OE(en), .A(xdata[149]), .Z(CGFidata[149]));
Q_BUFZP U516 ( .OE(en), .A(xdata[150]), .Z(CGFidata[150]));
Q_BUFZP U517 ( .OE(en), .A(xdata[151]), .Z(CGFidata[151]));
Q_BUFZP U518 ( .OE(en), .A(xdata[152]), .Z(CGFidata[152]));
Q_BUFZP U519 ( .OE(en), .A(xdata[153]), .Z(CGFidata[153]));
Q_BUFZP U520 ( .OE(en), .A(xdata[154]), .Z(CGFidata[154]));
Q_BUFZP U521 ( .OE(en), .A(xdata[155]), .Z(CGFidata[155]));
Q_BUFZP U522 ( .OE(en), .A(xdata[156]), .Z(CGFidata[156]));
Q_BUFZP U523 ( .OE(en), .A(xdata[157]), .Z(CGFidata[157]));
Q_BUFZP U524 ( .OE(en), .A(xdata[158]), .Z(CGFidata[158]));
Q_BUFZP U525 ( .OE(en), .A(xdata[159]), .Z(CGFidata[159]));
Q_BUFZP U526 ( .OE(en), .A(xdata[160]), .Z(CGFidata[160]));
Q_BUFZP U527 ( .OE(en), .A(xdata[161]), .Z(CGFidata[161]));
Q_BUFZP U528 ( .OE(en), .A(xdata[162]), .Z(CGFidata[162]));
Q_BUFZP U529 ( .OE(en), .A(xdata[163]), .Z(CGFidata[163]));
Q_BUFZP U530 ( .OE(en), .A(xdata[164]), .Z(CGFidata[164]));
Q_BUFZP U531 ( .OE(en), .A(xdata[165]), .Z(CGFidata[165]));
Q_BUFZP U532 ( .OE(en), .A(xdata[166]), .Z(CGFidata[166]));
Q_BUFZP U533 ( .OE(en), .A(xdata[167]), .Z(CGFidata[167]));
Q_BUFZP U534 ( .OE(en), .A(xdata[168]), .Z(CGFidata[168]));
Q_BUFZP U535 ( .OE(en), .A(xdata[169]), .Z(CGFidata[169]));
Q_BUFZP U536 ( .OE(en), .A(xdata[170]), .Z(CGFidata[170]));
Q_BUFZP U537 ( .OE(en), .A(xdata[171]), .Z(CGFidata[171]));
Q_BUFZP U538 ( .OE(en), .A(xdata[172]), .Z(CGFidata[172]));
Q_BUFZP U539 ( .OE(en), .A(xdata[173]), .Z(CGFidata[173]));
Q_BUFZP U540 ( .OE(en), .A(xdata[174]), .Z(CGFidata[174]));
Q_BUFZP U541 ( .OE(en), .A(xdata[175]), .Z(CGFidata[175]));
Q_BUFZP U542 ( .OE(en), .A(xdata[176]), .Z(CGFidata[176]));
Q_BUFZP U543 ( .OE(en), .A(xdata[177]), .Z(CGFidata[177]));
Q_BUFZP U544 ( .OE(en), .A(xdata[178]), .Z(CGFidata[178]));
Q_BUFZP U545 ( .OE(en), .A(xdata[179]), .Z(CGFidata[179]));
Q_BUFZP U546 ( .OE(en), .A(xdata[180]), .Z(CGFidata[180]));
Q_BUFZP U547 ( .OE(en), .A(xdata[181]), .Z(CGFidata[181]));
Q_BUFZP U548 ( .OE(en), .A(xdata[182]), .Z(CGFidata[182]));
Q_BUFZP U549 ( .OE(en), .A(xdata[183]), .Z(CGFidata[183]));
Q_BUFZP U550 ( .OE(en), .A(xdata[184]), .Z(CGFidata[184]));
Q_BUFZP U551 ( .OE(en), .A(xdata[185]), .Z(CGFidata[185]));
Q_BUFZP U552 ( .OE(en), .A(xdata[186]), .Z(CGFidata[186]));
Q_BUFZP U553 ( .OE(en), .A(xdata[187]), .Z(CGFidata[187]));
Q_BUFZP U554 ( .OE(en), .A(xdata[188]), .Z(CGFidata[188]));
Q_BUFZP U555 ( .OE(en), .A(xdata[189]), .Z(CGFidata[189]));
Q_BUFZP U556 ( .OE(en), .A(xdata[190]), .Z(CGFidata[190]));
Q_BUFZP U557 ( .OE(en), .A(xdata[191]), .Z(CGFidata[191]));
Q_BUFZP U558 ( .OE(en), .A(xdata[192]), .Z(CGFidata[192]));
Q_BUFZP U559 ( .OE(en), .A(xdata[193]), .Z(CGFidata[193]));
Q_BUFZP U560 ( .OE(en), .A(xdata[194]), .Z(CGFidata[194]));
Q_BUFZP U561 ( .OE(en), .A(xdata[195]), .Z(CGFidata[195]));
Q_BUFZP U562 ( .OE(en), .A(xdata[196]), .Z(CGFidata[196]));
Q_BUFZP U563 ( .OE(en), .A(xdata[197]), .Z(CGFidata[197]));
Q_BUFZP U564 ( .OE(en), .A(xdata[198]), .Z(CGFidata[198]));
Q_BUFZP U565 ( .OE(en), .A(xdata[199]), .Z(CGFidata[199]));
Q_BUFZP U566 ( .OE(en), .A(xdata[200]), .Z(CGFidata[200]));
Q_BUFZP U567 ( .OE(en), .A(xdata[201]), .Z(CGFidata[201]));
Q_BUFZP U568 ( .OE(en), .A(xdata[202]), .Z(CGFidata[202]));
Q_BUFZP U569 ( .OE(en), .A(xdata[203]), .Z(CGFidata[203]));
Q_BUFZP U570 ( .OE(en), .A(xdata[204]), .Z(CGFidata[204]));
Q_BUFZP U571 ( .OE(en), .A(xdata[205]), .Z(CGFidata[205]));
Q_BUFZP U572 ( .OE(en), .A(xdata[206]), .Z(CGFidata[206]));
Q_BUFZP U573 ( .OE(en), .A(xdata[207]), .Z(CGFidata[207]));
Q_BUFZP U574 ( .OE(en), .A(xdata[208]), .Z(CGFidata[208]));
Q_BUFZP U575 ( .OE(en), .A(xdata[209]), .Z(CGFidata[209]));
Q_BUFZP U576 ( .OE(en), .A(xdata[210]), .Z(CGFidata[210]));
Q_BUFZP U577 ( .OE(en), .A(xdata[211]), .Z(CGFidata[211]));
Q_BUFZP U578 ( .OE(en), .A(xdata[212]), .Z(CGFidata[212]));
Q_BUFZP U579 ( .OE(en), .A(xdata[213]), .Z(CGFidata[213]));
Q_BUFZP U580 ( .OE(en), .A(xdata[214]), .Z(CGFidata[214]));
Q_BUFZP U581 ( .OE(en), .A(xdata[215]), .Z(CGFidata[215]));
Q_BUFZP U582 ( .OE(en), .A(xdata[216]), .Z(CGFidata[216]));
Q_BUFZP U583 ( .OE(en), .A(xdata[217]), .Z(CGFidata[217]));
Q_BUFZP U584 ( .OE(en), .A(xdata[218]), .Z(CGFidata[218]));
Q_BUFZP U585 ( .OE(en), .A(xdata[219]), .Z(CGFidata[219]));
Q_BUFZP U586 ( .OE(en), .A(xdata[220]), .Z(CGFidata[220]));
Q_BUFZP U587 ( .OE(en), .A(xdata[221]), .Z(CGFidata[221]));
Q_BUFZP U588 ( .OE(en), .A(xdata[222]), .Z(CGFidata[222]));
Q_BUFZP U589 ( .OE(en), .A(xdata[223]), .Z(CGFidata[223]));
Q_BUFZP U590 ( .OE(en), .A(xdata[224]), .Z(CGFidata[224]));
Q_BUFZP U591 ( .OE(en), .A(xdata[225]), .Z(CGFidata[225]));
Q_BUFZP U592 ( .OE(en), .A(xdata[226]), .Z(CGFidata[226]));
Q_BUFZP U593 ( .OE(en), .A(xdata[227]), .Z(CGFidata[227]));
Q_BUFZP U594 ( .OE(en), .A(xdata[228]), .Z(CGFidata[228]));
Q_BUFZP U595 ( .OE(en), .A(xdata[229]), .Z(CGFidata[229]));
Q_BUFZP U596 ( .OE(en), .A(xdata[230]), .Z(CGFidata[230]));
Q_BUFZP U597 ( .OE(en), .A(xdata[231]), .Z(CGFidata[231]));
Q_BUFZP U598 ( .OE(en), .A(xdata[232]), .Z(CGFidata[232]));
Q_BUFZP U599 ( .OE(en), .A(xdata[233]), .Z(CGFidata[233]));
Q_BUFZP U600 ( .OE(en), .A(xdata[234]), .Z(CGFidata[234]));
Q_BUFZP U601 ( .OE(en), .A(xdata[235]), .Z(CGFidata[235]));
Q_BUFZP U602 ( .OE(en), .A(xdata[236]), .Z(CGFidata[236]));
Q_BUFZP U603 ( .OE(en), .A(xdata[237]), .Z(CGFidata[237]));
Q_BUFZP U604 ( .OE(en), .A(xdata[238]), .Z(CGFidata[238]));
Q_BUFZP U605 ( .OE(en), .A(xdata[239]), .Z(CGFidata[239]));
Q_BUFZP U606 ( .OE(en), .A(xdata[240]), .Z(CGFidata[240]));
Q_BUFZP U607 ( .OE(en), .A(xdata[241]), .Z(CGFidata[241]));
Q_BUFZP U608 ( .OE(en), .A(xdata[242]), .Z(CGFidata[242]));
Q_BUFZP U609 ( .OE(en), .A(xdata[243]), .Z(CGFidata[243]));
Q_BUFZP U610 ( .OE(en), .A(xdata[244]), .Z(CGFidata[244]));
Q_BUFZP U611 ( .OE(en), .A(xdata[245]), .Z(CGFidata[245]));
Q_BUFZP U612 ( .OE(en), .A(xdata[246]), .Z(CGFidata[246]));
Q_BUFZP U613 ( .OE(en), .A(xdata[247]), .Z(CGFidata[247]));
Q_BUFZP U614 ( .OE(en), .A(xdata[248]), .Z(CGFidata[248]));
Q_BUFZP U615 ( .OE(en), .A(xdata[249]), .Z(CGFidata[249]));
Q_BUFZP U616 ( .OE(en), .A(xdata[250]), .Z(CGFidata[250]));
Q_BUFZP U617 ( .OE(en), .A(xdata[251]), .Z(CGFidata[251]));
Q_BUFZP U618 ( .OE(en), .A(xdata[252]), .Z(CGFidata[252]));
Q_BUFZP U619 ( .OE(en), .A(xdata[253]), .Z(CGFidata[253]));
Q_BUFZP U620 ( .OE(en), .A(xdata[254]), .Z(CGFidata[254]));
Q_BUFZP U621 ( .OE(en), .A(xdata[255]), .Z(CGFidata[255]));
Q_BUFZP U622 ( .OE(en), .A(xdata[256]), .Z(CGFidata[256]));
Q_BUFZP U623 ( .OE(en), .A(xdata[257]), .Z(CGFidata[257]));
Q_BUFZP U624 ( .OE(en), .A(xdata[258]), .Z(CGFidata[258]));
Q_BUFZP U625 ( .OE(en), .A(xdata[259]), .Z(CGFidata[259]));
Q_BUFZP U626 ( .OE(en), .A(xdata[260]), .Z(CGFidata[260]));
Q_BUFZP U627 ( .OE(en), .A(xdata[261]), .Z(CGFidata[261]));
Q_BUFZP U628 ( .OE(en), .A(xdata[262]), .Z(CGFidata[262]));
Q_BUFZP U629 ( .OE(en), .A(xdata[263]), .Z(CGFidata[263]));
Q_BUFZP U630 ( .OE(en), .A(xdata[264]), .Z(CGFidata[264]));
Q_BUFZP U631 ( .OE(en), .A(xdata[265]), .Z(CGFidata[265]));
Q_BUFZP U632 ( .OE(en), .A(xdata[266]), .Z(CGFidata[266]));
Q_BUFZP U633 ( .OE(en), .A(xdata[267]), .Z(CGFidata[267]));
Q_BUFZP U634 ( .OE(en), .A(xdata[268]), .Z(CGFidata[268]));
Q_BUFZP U635 ( .OE(en), .A(xdata[269]), .Z(CGFidata[269]));
Q_BUFZP U636 ( .OE(en), .A(xdata[270]), .Z(CGFidata[270]));
Q_BUFZP U637 ( .OE(en), .A(xdata[271]), .Z(CGFidata[271]));
Q_BUFZP U638 ( .OE(en), .A(xdata[272]), .Z(CGFidata[272]));
Q_BUFZP U639 ( .OE(en), .A(xdata[273]), .Z(CGFidata[273]));
Q_BUFZP U640 ( .OE(en), .A(xdata[274]), .Z(CGFidata[274]));
Q_BUFZP U641 ( .OE(en), .A(xdata[275]), .Z(CGFidata[275]));
Q_BUFZP U642 ( .OE(en), .A(xdata[276]), .Z(CGFidata[276]));
Q_BUFZP U643 ( .OE(en), .A(xdata[277]), .Z(CGFidata[277]));
Q_BUFZP U644 ( .OE(en), .A(xdata[278]), .Z(CGFidata[278]));
Q_BUFZP U645 ( .OE(en), .A(xdata[279]), .Z(CGFidata[279]));
Q_BUFZP U646 ( .OE(enq), .A(n5), .Z(CLBreq));
Q_INV U647 ( .A(CLBwr[2]), .Z(n6));
ixc_bind \genblk3.b5 ( CLBfull, IXC_GFIFO.O.O.LBfull);
ixc_bind_4 \genblk3.b4 ( CLBwr[3:0], IXC_GFIFO.O.O.LBwr[3:0]);
ixc_bind_4 \genblk3.b3 ( CLBrd[3:0], IXC_GFIFO.O.O.LBrd[3:0]);
ixc_bind \genblk3.b2 ( CLBreq, IXC_GFIFO.O.O.LBreq);
ixc_bind \genblk3.b1 ( CGFfull, IXC_GFIFO.O.O.GFfull);
ixc_bind \genblk3.b0 ( CGFtsReq, IXC_GFIFO.O.O.GFtsReq);
Q_MX02 U654 ( .S(xc_top.GFLock2), .A0(oreq), .A1(ireq), .Z(n8));
Q_FDP0UA U655 ( .D(n9), .QTFCLK( ), .Q(ack));
Q_MX02 U656 ( .S(n14), .A0(ack), .A1(n8), .Z(n9));
Q_FDP0UA U657 ( .D(n10), .QTFCLK( ), .Q(en));
Q_NR02 U658 ( .A0(xc_top.GFLock2), .A1(n11), .Z(n10));
Q_OR02 U659 ( .A0(xc_top.GFLock2), .A1(n12), .Z(n14));
Q_INV U660 ( .A(n11), .Z(n12));
Q_OR03 U661 ( .A0(n4), .A1(tkin), .A2(n13), .Z(n11));
Q_OR02 U662 ( .A0(Rtkin), .A1(CGFfull), .Z(n13));
Q_MX02 U663 ( .S(CLBfull), .A0(ireq), .A1(ireqR), .Z(n15));
Q_FDP0UA U664 ( .D(n15), .QTFCLK( ), .Q(ireqR));
Q_AN02 U665 ( .A0(CLBwr[0]), .A1(n6), .Z(n16));
Q_AN02 U666 ( .A0(CLBwr[1]), .A1(n6), .Z(n17));
Q_INV U667 ( .A(n16), .Z(n18));
Q_INV U668 ( .A(n17), .Z(n19));
Q_NR02 U669 ( .A0(n17), .A1(n16), .Z(n20));
Q_AN02 U670 ( .A0(n19), .A1(n16), .Z(n21));
Q_AN02 U671 ( .A0(n17), .A1(n18), .Z(n22));
Q_AN02 U672 ( .A0(n17), .A1(n16), .Z(n23));
Q_AN02 U673 ( .A0(n20), .A1(n6), .Z(n24));
Q_LDP0 \_zzLB_REG[0][0] ( .G(n24), .D(cbid[0]), .Q(\_zzLB[0][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][1] ( .G(n24), .D(cbid[1]), .Q(\_zzLB[0][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][2] ( .G(n24), .D(cbid[2]), .Q(\_zzLB[0][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][3] ( .G(n24), .D(cbid[3]), .Q(\_zzLB[0][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][4] ( .G(n24), .D(cbid[4]), .Q(\_zzLB[0][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][5] ( .G(n24), .D(cbid[5]), .Q(\_zzLB[0][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][6] ( .G(n24), .D(cbid[6]), .Q(\_zzLB[0][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][7] ( .G(n24), .D(cbid[7]), .Q(\_zzLB[0][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][8] ( .G(n24), .D(cbid[8]), .Q(\_zzLB[0][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][9] ( .G(n24), .D(cbid[9]), .Q(\_zzLB[0][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][10] ( .G(n24), .D(cbid[10]), .Q(\_zzLB[0][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][11] ( .G(n24), .D(cbid[11]), .Q(\_zzLB[0][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][12] ( .G(n24), .D(cbid[12]), .Q(\_zzLB[0][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][13] ( .G(n24), .D(cbid[13]), .Q(\_zzLB[0][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][14] ( .G(n24), .D(cbid[14]), .Q(\_zzLB[0][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][15] ( .G(n24), .D(cbid[15]), .Q(\_zzLB[0][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][16] ( .G(n24), .D(cbid[16]), .Q(\_zzLB[0][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][17] ( .G(n24), .D(cbid[17]), .Q(\_zzLB[0][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][18] ( .G(n24), .D(cbid[18]), .Q(\_zzLB[0][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][19] ( .G(n24), .D(cbid[19]), .Q(\_zzLB[0][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][20] ( .G(n24), .D(idata[0]), .Q(\_zzLB[0][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][21] ( .G(n24), .D(idata[1]), .Q(\_zzLB[0][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][22] ( .G(n24), .D(idata[2]), .Q(\_zzLB[0][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][23] ( .G(n24), .D(idata[3]), .Q(\_zzLB[0][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][24] ( .G(n24), .D(idata[4]), .Q(\_zzLB[0][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][25] ( .G(n24), .D(idata[5]), .Q(\_zzLB[0][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][26] ( .G(n24), .D(idata[6]), .Q(\_zzLB[0][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][27] ( .G(n24), .D(idata[7]), .Q(\_zzLB[0][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][28] ( .G(n24), .D(idata[8]), .Q(\_zzLB[0][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][29] ( .G(n24), .D(idata[9]), .Q(\_zzLB[0][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][30] ( .G(n24), .D(idata[10]), .Q(\_zzLB[0][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][31] ( .G(n24), .D(idata[11]), .Q(\_zzLB[0][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][32] ( .G(n24), .D(idata[12]), .Q(\_zzLB[0][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][33] ( .G(n24), .D(idata[13]), .Q(\_zzLB[0][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][34] ( .G(n24), .D(idata[14]), .Q(\_zzLB[0][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][35] ( .G(n24), .D(idata[15]), .Q(\_zzLB[0][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][36] ( .G(n24), .D(idata[16]), .Q(\_zzLB[0][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][37] ( .G(n24), .D(idata[17]), .Q(\_zzLB[0][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][38] ( .G(n24), .D(idata[18]), .Q(\_zzLB[0][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][39] ( .G(n24), .D(idata[19]), .Q(\_zzLB[0][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][40] ( .G(n24), .D(idata[20]), .Q(\_zzLB[0][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][41] ( .G(n24), .D(idata[21]), .Q(\_zzLB[0][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][42] ( .G(n24), .D(idata[22]), .Q(\_zzLB[0][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][43] ( .G(n24), .D(idata[23]), .Q(\_zzLB[0][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][44] ( .G(n24), .D(idata[24]), .Q(\_zzLB[0][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][45] ( .G(n24), .D(idata[25]), .Q(\_zzLB[0][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][46] ( .G(n24), .D(idata[26]), .Q(\_zzLB[0][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][47] ( .G(n24), .D(idata[27]), .Q(\_zzLB[0][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][48] ( .G(n24), .D(idata[28]), .Q(\_zzLB[0][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][49] ( .G(n24), .D(idata[29]), .Q(\_zzLB[0][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][50] ( .G(n24), .D(idata[30]), .Q(\_zzLB[0][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][51] ( .G(n24), .D(idata[31]), .Q(\_zzLB[0][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][52] ( .G(n24), .D(idata[32]), .Q(\_zzLB[0][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][53] ( .G(n24), .D(idata[33]), .Q(\_zzLB[0][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][54] ( .G(n24), .D(idata[34]), .Q(\_zzLB[0][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][55] ( .G(n24), .D(idata[35]), .Q(\_zzLB[0][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][56] ( .G(n24), .D(idata[36]), .Q(\_zzLB[0][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][57] ( .G(n24), .D(idata[37]), .Q(\_zzLB[0][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][58] ( .G(n24), .D(idata[38]), .Q(\_zzLB[0][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][59] ( .G(n24), .D(idata[39]), .Q(\_zzLB[0][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][60] ( .G(n24), .D(idata[40]), .Q(\_zzLB[0][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][61] ( .G(n24), .D(idata[41]), .Q(\_zzLB[0][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][62] ( .G(n24), .D(idata[42]), .Q(\_zzLB[0][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][63] ( .G(n24), .D(idata[43]), .Q(\_zzLB[0][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][64] ( .G(n24), .D(idata[44]), .Q(\_zzLB[0][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][65] ( .G(n24), .D(idata[45]), .Q(\_zzLB[0][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][66] ( .G(n24), .D(idata[46]), .Q(\_zzLB[0][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][67] ( .G(n24), .D(idata[47]), .Q(\_zzLB[0][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][68] ( .G(n24), .D(idata[48]), .Q(\_zzLB[0][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][69] ( .G(n24), .D(idata[49]), .Q(\_zzLB[0][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][70] ( .G(n24), .D(idata[50]), .Q(\_zzLB[0][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][71] ( .G(n24), .D(idata[51]), .Q(\_zzLB[0][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][72] ( .G(n24), .D(idata[52]), .Q(\_zzLB[0][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][73] ( .G(n24), .D(idata[53]), .Q(\_zzLB[0][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][74] ( .G(n24), .D(idata[54]), .Q(\_zzLB[0][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][75] ( .G(n24), .D(idata[55]), .Q(\_zzLB[0][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][76] ( .G(n24), .D(idata[56]), .Q(\_zzLB[0][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][77] ( .G(n24), .D(idata[57]), .Q(\_zzLB[0][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][78] ( .G(n24), .D(idata[58]), .Q(\_zzLB[0][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][79] ( .G(n24), .D(idata[59]), .Q(\_zzLB[0][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][80] ( .G(n24), .D(idata[60]), .Q(\_zzLB[0][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][81] ( .G(n24), .D(idata[61]), .Q(\_zzLB[0][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][82] ( .G(n24), .D(idata[62]), .Q(\_zzLB[0][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][83] ( .G(n24), .D(idata[63]), .Q(\_zzLB[0][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][84] ( .G(n24), .D(idata[64]), .Q(\_zzLB[0][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][85] ( .G(n24), .D(idata[65]), .Q(\_zzLB[0][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][86] ( .G(n24), .D(idata[66]), .Q(\_zzLB[0][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][87] ( .G(n24), .D(idata[67]), .Q(\_zzLB[0][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][88] ( .G(n24), .D(idata[68]), .Q(\_zzLB[0][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][89] ( .G(n24), .D(idata[69]), .Q(\_zzLB[0][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][90] ( .G(n24), .D(idata[70]), .Q(\_zzLB[0][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][91] ( .G(n24), .D(idata[71]), .Q(\_zzLB[0][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][92] ( .G(n24), .D(idata[72]), .Q(\_zzLB[0][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][93] ( .G(n24), .D(idata[73]), .Q(\_zzLB[0][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][94] ( .G(n24), .D(idata[74]), .Q(\_zzLB[0][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][95] ( .G(n24), .D(idata[75]), .Q(\_zzLB[0][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][96] ( .G(n24), .D(idata[76]), .Q(\_zzLB[0][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][97] ( .G(n24), .D(idata[77]), .Q(\_zzLB[0][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][98] ( .G(n24), .D(idata[78]), .Q(\_zzLB[0][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][99] ( .G(n24), .D(idata[79]), .Q(\_zzLB[0][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][100] ( .G(n24), .D(idata[80]), .Q(\_zzLB[0][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][101] ( .G(n24), .D(idata[81]), .Q(\_zzLB[0][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][102] ( .G(n24), .D(idata[82]), .Q(\_zzLB[0][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][103] ( .G(n24), .D(idata[83]), .Q(\_zzLB[0][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][104] ( .G(n24), .D(idata[84]), .Q(\_zzLB[0][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][105] ( .G(n24), .D(idata[85]), .Q(\_zzLB[0][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][106] ( .G(n24), .D(idata[86]), .Q(\_zzLB[0][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][107] ( .G(n24), .D(idata[87]), .Q(\_zzLB[0][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][108] ( .G(n24), .D(idata[88]), .Q(\_zzLB[0][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][109] ( .G(n24), .D(idata[89]), .Q(\_zzLB[0][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][110] ( .G(n24), .D(idata[90]), .Q(\_zzLB[0][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][111] ( .G(n24), .D(idata[91]), .Q(\_zzLB[0][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][112] ( .G(n24), .D(idata[92]), .Q(\_zzLB[0][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][113] ( .G(n24), .D(idata[93]), .Q(\_zzLB[0][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][114] ( .G(n24), .D(idata[94]), .Q(\_zzLB[0][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][115] ( .G(n24), .D(idata[95]), .Q(\_zzLB[0][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][116] ( .G(n24), .D(idata[96]), .Q(\_zzLB[0][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][117] ( .G(n24), .D(idata[97]), .Q(\_zzLB[0][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][118] ( .G(n24), .D(idata[98]), .Q(\_zzLB[0][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][119] ( .G(n24), .D(idata[99]), .Q(\_zzLB[0][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][120] ( .G(n24), .D(idata[100]), .Q(\_zzLB[0][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][121] ( .G(n24), .D(idata[101]), .Q(\_zzLB[0][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][122] ( .G(n24), .D(idata[102]), .Q(\_zzLB[0][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][123] ( .G(n24), .D(idata[103]), .Q(\_zzLB[0][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][124] ( .G(n24), .D(idata[104]), .Q(\_zzLB[0][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][125] ( .G(n24), .D(idata[105]), .Q(\_zzLB[0][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][126] ( .G(n24), .D(idata[106]), .Q(\_zzLB[0][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][127] ( .G(n24), .D(idata[107]), .Q(\_zzLB[0][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][128] ( .G(n24), .D(idata[108]), .Q(\_zzLB[0][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][129] ( .G(n24), .D(idata[109]), .Q(\_zzLB[0][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][130] ( .G(n24), .D(idata[110]), .Q(\_zzLB[0][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][131] ( .G(n24), .D(idata[111]), .Q(\_zzLB[0][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][132] ( .G(n24), .D(idata[112]), .Q(\_zzLB[0][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][133] ( .G(n24), .D(idata[113]), .Q(\_zzLB[0][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][134] ( .G(n24), .D(idata[114]), .Q(\_zzLB[0][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][135] ( .G(n24), .D(idata[115]), .Q(\_zzLB[0][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][136] ( .G(n24), .D(idata[116]), .Q(\_zzLB[0][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][137] ( .G(n24), .D(idata[117]), .Q(\_zzLB[0][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][138] ( .G(n24), .D(idata[118]), .Q(\_zzLB[0][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][139] ( .G(n24), .D(idata[119]), .Q(\_zzLB[0][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][140] ( .G(n24), .D(idata[120]), .Q(\_zzLB[0][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][141] ( .G(n24), .D(idata[121]), .Q(\_zzLB[0][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][142] ( .G(n24), .D(idata[122]), .Q(\_zzLB[0][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][143] ( .G(n24), .D(idata[123]), .Q(\_zzLB[0][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][144] ( .G(n24), .D(idata[124]), .Q(\_zzLB[0][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][145] ( .G(n24), .D(idata[125]), .Q(\_zzLB[0][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][146] ( .G(n24), .D(idata[126]), .Q(\_zzLB[0][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][147] ( .G(n24), .D(idata[127]), .Q(\_zzLB[0][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][148] ( .G(n24), .D(idata[128]), .Q(\_zzLB[0][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][149] ( .G(n24), .D(idata[129]), .Q(\_zzLB[0][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][150] ( .G(n24), .D(idata[130]), .Q(\_zzLB[0][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][151] ( .G(n24), .D(idata[131]), .Q(\_zzLB[0][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][152] ( .G(n24), .D(idata[132]), .Q(\_zzLB[0][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][153] ( .G(n24), .D(idata[133]), .Q(\_zzLB[0][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][154] ( .G(n24), .D(idata[134]), .Q(\_zzLB[0][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][155] ( .G(n24), .D(idata[135]), .Q(\_zzLB[0][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][156] ( .G(n24), .D(idata[136]), .Q(\_zzLB[0][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][157] ( .G(n24), .D(idata[137]), .Q(\_zzLB[0][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][158] ( .G(n24), .D(idata[138]), .Q(\_zzLB[0][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][159] ( .G(n24), .D(idata[139]), .Q(\_zzLB[0][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][160] ( .G(n24), .D(idata[140]), .Q(\_zzLB[0][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][161] ( .G(n24), .D(idata[141]), .Q(\_zzLB[0][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][162] ( .G(n24), .D(idata[142]), .Q(\_zzLB[0][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][163] ( .G(n24), .D(idata[143]), .Q(\_zzLB[0][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][164] ( .G(n24), .D(idata[144]), .Q(\_zzLB[0][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][165] ( .G(n24), .D(idata[145]), .Q(\_zzLB[0][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][166] ( .G(n24), .D(idata[146]), .Q(\_zzLB[0][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][167] ( .G(n24), .D(idata[147]), .Q(\_zzLB[0][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][168] ( .G(n24), .D(idata[148]), .Q(\_zzLB[0][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][169] ( .G(n24), .D(idata[149]), .Q(\_zzLB[0][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][170] ( .G(n24), .D(idata[150]), .Q(\_zzLB[0][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][171] ( .G(n24), .D(idata[151]), .Q(\_zzLB[0][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][172] ( .G(n24), .D(idata[152]), .Q(\_zzLB[0][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][173] ( .G(n24), .D(idata[153]), .Q(\_zzLB[0][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][174] ( .G(n24), .D(idata[154]), .Q(\_zzLB[0][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][175] ( .G(n24), .D(idata[155]), .Q(\_zzLB[0][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][176] ( .G(n24), .D(idata[156]), .Q(\_zzLB[0][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][177] ( .G(n24), .D(idata[157]), .Q(\_zzLB[0][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][178] ( .G(n24), .D(idata[158]), .Q(\_zzLB[0][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][179] ( .G(n24), .D(idata[159]), .Q(\_zzLB[0][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][180] ( .G(n24), .D(idata[160]), .Q(\_zzLB[0][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][181] ( .G(n24), .D(idata[161]), .Q(\_zzLB[0][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][182] ( .G(n24), .D(idata[162]), .Q(\_zzLB[0][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][183] ( .G(n24), .D(idata[163]), .Q(\_zzLB[0][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][184] ( .G(n24), .D(idata[164]), .Q(\_zzLB[0][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][185] ( .G(n24), .D(idata[165]), .Q(\_zzLB[0][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][186] ( .G(n24), .D(idata[166]), .Q(\_zzLB[0][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][187] ( .G(n24), .D(idata[167]), .Q(\_zzLB[0][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][188] ( .G(n24), .D(idata[168]), .Q(\_zzLB[0][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][189] ( .G(n24), .D(idata[169]), .Q(\_zzLB[0][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][190] ( .G(n24), .D(idata[170]), .Q(\_zzLB[0][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][191] ( .G(n24), .D(idata[171]), .Q(\_zzLB[0][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][192] ( .G(n24), .D(idata[172]), .Q(\_zzLB[0][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][193] ( .G(n24), .D(idata[173]), .Q(\_zzLB[0][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][194] ( .G(n24), .D(idata[174]), .Q(\_zzLB[0][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][195] ( .G(n24), .D(idata[175]), .Q(\_zzLB[0][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][196] ( .G(n24), .D(idata[176]), .Q(\_zzLB[0][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][197] ( .G(n24), .D(idata[177]), .Q(\_zzLB[0][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][198] ( .G(n24), .D(idata[178]), .Q(\_zzLB[0][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][199] ( .G(n24), .D(idata[179]), .Q(\_zzLB[0][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][200] ( .G(n24), .D(idata[180]), .Q(\_zzLB[0][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][201] ( .G(n24), .D(idata[181]), .Q(\_zzLB[0][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][202] ( .G(n24), .D(idata[182]), .Q(\_zzLB[0][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][203] ( .G(n24), .D(idata[183]), .Q(\_zzLB[0][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][204] ( .G(n24), .D(idata[184]), .Q(\_zzLB[0][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][205] ( .G(n24), .D(idata[185]), .Q(\_zzLB[0][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][206] ( .G(n24), .D(idata[186]), .Q(\_zzLB[0][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][207] ( .G(n24), .D(idata[187]), .Q(\_zzLB[0][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][208] ( .G(n24), .D(idata[188]), .Q(\_zzLB[0][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][209] ( .G(n24), .D(idata[189]), .Q(\_zzLB[0][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][210] ( .G(n24), .D(idata[190]), .Q(\_zzLB[0][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][211] ( .G(n24), .D(idata[191]), .Q(\_zzLB[0][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][212] ( .G(n24), .D(idata[192]), .Q(\_zzLB[0][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][213] ( .G(n24), .D(idata[193]), .Q(\_zzLB[0][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][214] ( .G(n24), .D(idata[194]), .Q(\_zzLB[0][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][215] ( .G(n24), .D(idata[195]), .Q(\_zzLB[0][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][216] ( .G(n24), .D(idata[196]), .Q(\_zzLB[0][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][217] ( .G(n24), .D(idata[197]), .Q(\_zzLB[0][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][218] ( .G(n24), .D(idata[198]), .Q(\_zzLB[0][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][219] ( .G(n24), .D(idata[199]), .Q(\_zzLB[0][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][220] ( .G(n24), .D(idata[200]), .Q(\_zzLB[0][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][221] ( .G(n24), .D(idata[201]), .Q(\_zzLB[0][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][222] ( .G(n24), .D(idata[202]), .Q(\_zzLB[0][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][223] ( .G(n24), .D(idata[203]), .Q(\_zzLB[0][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][224] ( .G(n24), .D(idata[204]), .Q(\_zzLB[0][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][225] ( .G(n24), .D(idata[205]), .Q(\_zzLB[0][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][226] ( .G(n24), .D(idata[206]), .Q(\_zzLB[0][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][227] ( .G(n24), .D(idata[207]), .Q(\_zzLB[0][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][228] ( .G(n24), .D(idata[208]), .Q(\_zzLB[0][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][229] ( .G(n24), .D(idata[209]), .Q(\_zzLB[0][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][230] ( .G(n24), .D(idata[210]), .Q(\_zzLB[0][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][231] ( .G(n24), .D(idata[211]), .Q(\_zzLB[0][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][232] ( .G(n24), .D(idata[212]), .Q(\_zzLB[0][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][233] ( .G(n24), .D(idata[213]), .Q(\_zzLB[0][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][234] ( .G(n24), .D(idata[214]), .Q(\_zzLB[0][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][235] ( .G(n24), .D(idata[215]), .Q(\_zzLB[0][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][236] ( .G(n24), .D(idata[216]), .Q(\_zzLB[0][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][237] ( .G(n24), .D(idata[217]), .Q(\_zzLB[0][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][238] ( .G(n24), .D(idata[218]), .Q(\_zzLB[0][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][239] ( .G(n24), .D(idata[219]), .Q(\_zzLB[0][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][240] ( .G(n24), .D(idata[220]), .Q(\_zzLB[0][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][241] ( .G(n24), .D(idata[221]), .Q(\_zzLB[0][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][242] ( .G(n24), .D(idata[222]), .Q(\_zzLB[0][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][243] ( .G(n24), .D(idata[223]), .Q(\_zzLB[0][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][244] ( .G(n24), .D(idata[224]), .Q(\_zzLB[0][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][245] ( .G(n24), .D(idata[225]), .Q(\_zzLB[0][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][246] ( .G(n24), .D(idata[226]), .Q(\_zzLB[0][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][247] ( .G(n24), .D(idata[227]), .Q(\_zzLB[0][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][248] ( .G(n24), .D(idata[228]), .Q(\_zzLB[0][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][249] ( .G(n24), .D(idata[229]), .Q(\_zzLB[0][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][250] ( .G(n24), .D(idata[230]), .Q(\_zzLB[0][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][251] ( .G(n24), .D(idata[231]), .Q(\_zzLB[0][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][252] ( .G(n24), .D(idata[232]), .Q(\_zzLB[0][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][253] ( .G(n24), .D(idata[233]), .Q(\_zzLB[0][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][254] ( .G(n24), .D(idata[234]), .Q(\_zzLB[0][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][255] ( .G(n24), .D(idata[235]), .Q(\_zzLB[0][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][256] ( .G(n24), .D(idata[236]), .Q(\_zzLB[0][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][257] ( .G(n24), .D(idata[237]), .Q(\_zzLB[0][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][258] ( .G(n24), .D(idata[238]), .Q(\_zzLB[0][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][259] ( .G(n24), .D(idata[239]), .Q(\_zzLB[0][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][260] ( .G(n24), .D(idata[240]), .Q(\_zzLB[0][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][261] ( .G(n24), .D(idata[241]), .Q(\_zzLB[0][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][262] ( .G(n24), .D(idata[242]), .Q(\_zzLB[0][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][263] ( .G(n24), .D(idata[243]), .Q(\_zzLB[0][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][264] ( .G(n24), .D(idata[244]), .Q(\_zzLB[0][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][265] ( .G(n24), .D(idata[245]), .Q(\_zzLB[0][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][266] ( .G(n24), .D(idata[246]), .Q(\_zzLB[0][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][267] ( .G(n24), .D(idata[247]), .Q(\_zzLB[0][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][268] ( .G(n24), .D(idata[248]), .Q(\_zzLB[0][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][269] ( .G(n24), .D(idata[249]), .Q(\_zzLB[0][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][270] ( .G(n24), .D(idata[250]), .Q(\_zzLB[0][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][271] ( .G(n24), .D(idata[251]), .Q(\_zzLB[0][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][272] ( .G(n24), .D(idata[252]), .Q(\_zzLB[0][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][273] ( .G(n24), .D(idata[253]), .Q(\_zzLB[0][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][274] ( .G(n24), .D(idata[254]), .Q(\_zzLB[0][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][275] ( .G(n24), .D(idata[255]), .Q(\_zzLB[0][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][276] ( .G(n24), .D(idata[256]), .Q(\_zzLB[0][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][277] ( .G(n24), .D(idata[257]), .Q(\_zzLB[0][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][278] ( .G(n24), .D(idata[258]), .Q(\_zzLB[0][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][279] ( .G(n24), .D(idata[259]), .Q(\_zzLB[0][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][280] ( .G(n24), .D(idata[260]), .Q(\_zzLB[0][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][281] ( .G(n24), .D(idata[261]), .Q(\_zzLB[0][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][282] ( .G(n24), .D(idata[262]), .Q(\_zzLB[0][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][283] ( .G(n24), .D(idata[263]), .Q(\_zzLB[0][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][284] ( .G(n24), .D(idata[264]), .Q(\_zzLB[0][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][285] ( .G(n24), .D(idata[265]), .Q(\_zzLB[0][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][286] ( .G(n24), .D(idata[266]), .Q(\_zzLB[0][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][287] ( .G(n24), .D(idata[267]), .Q(\_zzLB[0][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][288] ( .G(n24), .D(idata[268]), .Q(\_zzLB[0][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][289] ( .G(n24), .D(idata[269]), .Q(\_zzLB[0][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][290] ( .G(n24), .D(idata[270]), .Q(\_zzLB[0][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][291] ( .G(n24), .D(idata[271]), .Q(\_zzLB[0][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][292] ( .G(n24), .D(idata[272]), .Q(\_zzLB[0][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][293] ( .G(n24), .D(idata[273]), .Q(\_zzLB[0][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][294] ( .G(n24), .D(idata[274]), .Q(\_zzLB[0][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][295] ( .G(n24), .D(idata[275]), .Q(\_zzLB[0][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][296] ( .G(n24), .D(idata[276]), .Q(\_zzLB[0][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][297] ( .G(n24), .D(idata[277]), .Q(\_zzLB[0][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][298] ( .G(n24), .D(idata[278]), .Q(\_zzLB[0][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][299] ( .G(n24), .D(idata[279]), .Q(\_zzLB[0][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[0][300] ( .G(n24), .D(ireq), .Q(\_zzLB[0][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][0] ( .G(n21), .D(cbid[0]), .Q(\_zzLB[1][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][1] ( .G(n21), .D(cbid[1]), .Q(\_zzLB[1][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][2] ( .G(n21), .D(cbid[2]), .Q(\_zzLB[1][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][3] ( .G(n21), .D(cbid[3]), .Q(\_zzLB[1][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][4] ( .G(n21), .D(cbid[4]), .Q(\_zzLB[1][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][5] ( .G(n21), .D(cbid[5]), .Q(\_zzLB[1][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][6] ( .G(n21), .D(cbid[6]), .Q(\_zzLB[1][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][7] ( .G(n21), .D(cbid[7]), .Q(\_zzLB[1][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][8] ( .G(n21), .D(cbid[8]), .Q(\_zzLB[1][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][9] ( .G(n21), .D(cbid[9]), .Q(\_zzLB[1][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][10] ( .G(n21), .D(cbid[10]), .Q(\_zzLB[1][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][11] ( .G(n21), .D(cbid[11]), .Q(\_zzLB[1][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][12] ( .G(n21), .D(cbid[12]), .Q(\_zzLB[1][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][13] ( .G(n21), .D(cbid[13]), .Q(\_zzLB[1][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][14] ( .G(n21), .D(cbid[14]), .Q(\_zzLB[1][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][15] ( .G(n21), .D(cbid[15]), .Q(\_zzLB[1][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][16] ( .G(n21), .D(cbid[16]), .Q(\_zzLB[1][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][17] ( .G(n21), .D(cbid[17]), .Q(\_zzLB[1][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][18] ( .G(n21), .D(cbid[18]), .Q(\_zzLB[1][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][19] ( .G(n21), .D(cbid[19]), .Q(\_zzLB[1][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][20] ( .G(n21), .D(idata[0]), .Q(\_zzLB[1][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][21] ( .G(n21), .D(idata[1]), .Q(\_zzLB[1][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][22] ( .G(n21), .D(idata[2]), .Q(\_zzLB[1][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][23] ( .G(n21), .D(idata[3]), .Q(\_zzLB[1][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][24] ( .G(n21), .D(idata[4]), .Q(\_zzLB[1][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][25] ( .G(n21), .D(idata[5]), .Q(\_zzLB[1][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][26] ( .G(n21), .D(idata[6]), .Q(\_zzLB[1][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][27] ( .G(n21), .D(idata[7]), .Q(\_zzLB[1][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][28] ( .G(n21), .D(idata[8]), .Q(\_zzLB[1][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][29] ( .G(n21), .D(idata[9]), .Q(\_zzLB[1][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][30] ( .G(n21), .D(idata[10]), .Q(\_zzLB[1][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][31] ( .G(n21), .D(idata[11]), .Q(\_zzLB[1][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][32] ( .G(n21), .D(idata[12]), .Q(\_zzLB[1][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][33] ( .G(n21), .D(idata[13]), .Q(\_zzLB[1][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][34] ( .G(n21), .D(idata[14]), .Q(\_zzLB[1][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][35] ( .G(n21), .D(idata[15]), .Q(\_zzLB[1][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][36] ( .G(n21), .D(idata[16]), .Q(\_zzLB[1][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][37] ( .G(n21), .D(idata[17]), .Q(\_zzLB[1][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][38] ( .G(n21), .D(idata[18]), .Q(\_zzLB[1][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][39] ( .G(n21), .D(idata[19]), .Q(\_zzLB[1][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][40] ( .G(n21), .D(idata[20]), .Q(\_zzLB[1][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][41] ( .G(n21), .D(idata[21]), .Q(\_zzLB[1][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][42] ( .G(n21), .D(idata[22]), .Q(\_zzLB[1][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][43] ( .G(n21), .D(idata[23]), .Q(\_zzLB[1][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][44] ( .G(n21), .D(idata[24]), .Q(\_zzLB[1][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][45] ( .G(n21), .D(idata[25]), .Q(\_zzLB[1][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][46] ( .G(n21), .D(idata[26]), .Q(\_zzLB[1][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][47] ( .G(n21), .D(idata[27]), .Q(\_zzLB[1][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][48] ( .G(n21), .D(idata[28]), .Q(\_zzLB[1][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][49] ( .G(n21), .D(idata[29]), .Q(\_zzLB[1][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][50] ( .G(n21), .D(idata[30]), .Q(\_zzLB[1][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][51] ( .G(n21), .D(idata[31]), .Q(\_zzLB[1][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][52] ( .G(n21), .D(idata[32]), .Q(\_zzLB[1][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][53] ( .G(n21), .D(idata[33]), .Q(\_zzLB[1][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][54] ( .G(n21), .D(idata[34]), .Q(\_zzLB[1][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][55] ( .G(n21), .D(idata[35]), .Q(\_zzLB[1][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][56] ( .G(n21), .D(idata[36]), .Q(\_zzLB[1][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][57] ( .G(n21), .D(idata[37]), .Q(\_zzLB[1][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][58] ( .G(n21), .D(idata[38]), .Q(\_zzLB[1][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][59] ( .G(n21), .D(idata[39]), .Q(\_zzLB[1][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][60] ( .G(n21), .D(idata[40]), .Q(\_zzLB[1][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][61] ( .G(n21), .D(idata[41]), .Q(\_zzLB[1][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][62] ( .G(n21), .D(idata[42]), .Q(\_zzLB[1][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][63] ( .G(n21), .D(idata[43]), .Q(\_zzLB[1][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][64] ( .G(n21), .D(idata[44]), .Q(\_zzLB[1][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][65] ( .G(n21), .D(idata[45]), .Q(\_zzLB[1][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][66] ( .G(n21), .D(idata[46]), .Q(\_zzLB[1][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][67] ( .G(n21), .D(idata[47]), .Q(\_zzLB[1][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][68] ( .G(n21), .D(idata[48]), .Q(\_zzLB[1][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][69] ( .G(n21), .D(idata[49]), .Q(\_zzLB[1][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][70] ( .G(n21), .D(idata[50]), .Q(\_zzLB[1][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][71] ( .G(n21), .D(idata[51]), .Q(\_zzLB[1][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][72] ( .G(n21), .D(idata[52]), .Q(\_zzLB[1][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][73] ( .G(n21), .D(idata[53]), .Q(\_zzLB[1][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][74] ( .G(n21), .D(idata[54]), .Q(\_zzLB[1][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][75] ( .G(n21), .D(idata[55]), .Q(\_zzLB[1][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][76] ( .G(n21), .D(idata[56]), .Q(\_zzLB[1][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][77] ( .G(n21), .D(idata[57]), .Q(\_zzLB[1][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][78] ( .G(n21), .D(idata[58]), .Q(\_zzLB[1][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][79] ( .G(n21), .D(idata[59]), .Q(\_zzLB[1][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][80] ( .G(n21), .D(idata[60]), .Q(\_zzLB[1][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][81] ( .G(n21), .D(idata[61]), .Q(\_zzLB[1][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][82] ( .G(n21), .D(idata[62]), .Q(\_zzLB[1][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][83] ( .G(n21), .D(idata[63]), .Q(\_zzLB[1][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][84] ( .G(n21), .D(idata[64]), .Q(\_zzLB[1][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][85] ( .G(n21), .D(idata[65]), .Q(\_zzLB[1][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][86] ( .G(n21), .D(idata[66]), .Q(\_zzLB[1][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][87] ( .G(n21), .D(idata[67]), .Q(\_zzLB[1][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][88] ( .G(n21), .D(idata[68]), .Q(\_zzLB[1][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][89] ( .G(n21), .D(idata[69]), .Q(\_zzLB[1][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][90] ( .G(n21), .D(idata[70]), .Q(\_zzLB[1][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][91] ( .G(n21), .D(idata[71]), .Q(\_zzLB[1][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][92] ( .G(n21), .D(idata[72]), .Q(\_zzLB[1][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][93] ( .G(n21), .D(idata[73]), .Q(\_zzLB[1][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][94] ( .G(n21), .D(idata[74]), .Q(\_zzLB[1][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][95] ( .G(n21), .D(idata[75]), .Q(\_zzLB[1][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][96] ( .G(n21), .D(idata[76]), .Q(\_zzLB[1][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][97] ( .G(n21), .D(idata[77]), .Q(\_zzLB[1][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][98] ( .G(n21), .D(idata[78]), .Q(\_zzLB[1][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][99] ( .G(n21), .D(idata[79]), .Q(\_zzLB[1][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][100] ( .G(n21), .D(idata[80]), .Q(\_zzLB[1][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][101] ( .G(n21), .D(idata[81]), .Q(\_zzLB[1][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][102] ( .G(n21), .D(idata[82]), .Q(\_zzLB[1][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][103] ( .G(n21), .D(idata[83]), .Q(\_zzLB[1][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][104] ( .G(n21), .D(idata[84]), .Q(\_zzLB[1][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][105] ( .G(n21), .D(idata[85]), .Q(\_zzLB[1][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][106] ( .G(n21), .D(idata[86]), .Q(\_zzLB[1][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][107] ( .G(n21), .D(idata[87]), .Q(\_zzLB[1][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][108] ( .G(n21), .D(idata[88]), .Q(\_zzLB[1][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][109] ( .G(n21), .D(idata[89]), .Q(\_zzLB[1][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][110] ( .G(n21), .D(idata[90]), .Q(\_zzLB[1][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][111] ( .G(n21), .D(idata[91]), .Q(\_zzLB[1][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][112] ( .G(n21), .D(idata[92]), .Q(\_zzLB[1][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][113] ( .G(n21), .D(idata[93]), .Q(\_zzLB[1][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][114] ( .G(n21), .D(idata[94]), .Q(\_zzLB[1][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][115] ( .G(n21), .D(idata[95]), .Q(\_zzLB[1][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][116] ( .G(n21), .D(idata[96]), .Q(\_zzLB[1][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][117] ( .G(n21), .D(idata[97]), .Q(\_zzLB[1][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][118] ( .G(n21), .D(idata[98]), .Q(\_zzLB[1][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][119] ( .G(n21), .D(idata[99]), .Q(\_zzLB[1][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][120] ( .G(n21), .D(idata[100]), .Q(\_zzLB[1][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][121] ( .G(n21), .D(idata[101]), .Q(\_zzLB[1][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][122] ( .G(n21), .D(idata[102]), .Q(\_zzLB[1][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][123] ( .G(n21), .D(idata[103]), .Q(\_zzLB[1][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][124] ( .G(n21), .D(idata[104]), .Q(\_zzLB[1][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][125] ( .G(n21), .D(idata[105]), .Q(\_zzLB[1][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][126] ( .G(n21), .D(idata[106]), .Q(\_zzLB[1][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][127] ( .G(n21), .D(idata[107]), .Q(\_zzLB[1][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][128] ( .G(n21), .D(idata[108]), .Q(\_zzLB[1][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][129] ( .G(n21), .D(idata[109]), .Q(\_zzLB[1][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][130] ( .G(n21), .D(idata[110]), .Q(\_zzLB[1][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][131] ( .G(n21), .D(idata[111]), .Q(\_zzLB[1][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][132] ( .G(n21), .D(idata[112]), .Q(\_zzLB[1][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][133] ( .G(n21), .D(idata[113]), .Q(\_zzLB[1][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][134] ( .G(n21), .D(idata[114]), .Q(\_zzLB[1][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][135] ( .G(n21), .D(idata[115]), .Q(\_zzLB[1][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][136] ( .G(n21), .D(idata[116]), .Q(\_zzLB[1][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][137] ( .G(n21), .D(idata[117]), .Q(\_zzLB[1][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][138] ( .G(n21), .D(idata[118]), .Q(\_zzLB[1][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][139] ( .G(n21), .D(idata[119]), .Q(\_zzLB[1][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][140] ( .G(n21), .D(idata[120]), .Q(\_zzLB[1][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][141] ( .G(n21), .D(idata[121]), .Q(\_zzLB[1][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][142] ( .G(n21), .D(idata[122]), .Q(\_zzLB[1][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][143] ( .G(n21), .D(idata[123]), .Q(\_zzLB[1][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][144] ( .G(n21), .D(idata[124]), .Q(\_zzLB[1][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][145] ( .G(n21), .D(idata[125]), .Q(\_zzLB[1][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][146] ( .G(n21), .D(idata[126]), .Q(\_zzLB[1][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][147] ( .G(n21), .D(idata[127]), .Q(\_zzLB[1][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][148] ( .G(n21), .D(idata[128]), .Q(\_zzLB[1][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][149] ( .G(n21), .D(idata[129]), .Q(\_zzLB[1][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][150] ( .G(n21), .D(idata[130]), .Q(\_zzLB[1][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][151] ( .G(n21), .D(idata[131]), .Q(\_zzLB[1][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][152] ( .G(n21), .D(idata[132]), .Q(\_zzLB[1][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][153] ( .G(n21), .D(idata[133]), .Q(\_zzLB[1][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][154] ( .G(n21), .D(idata[134]), .Q(\_zzLB[1][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][155] ( .G(n21), .D(idata[135]), .Q(\_zzLB[1][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][156] ( .G(n21), .D(idata[136]), .Q(\_zzLB[1][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][157] ( .G(n21), .D(idata[137]), .Q(\_zzLB[1][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][158] ( .G(n21), .D(idata[138]), .Q(\_zzLB[1][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][159] ( .G(n21), .D(idata[139]), .Q(\_zzLB[1][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][160] ( .G(n21), .D(idata[140]), .Q(\_zzLB[1][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][161] ( .G(n21), .D(idata[141]), .Q(\_zzLB[1][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][162] ( .G(n21), .D(idata[142]), .Q(\_zzLB[1][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][163] ( .G(n21), .D(idata[143]), .Q(\_zzLB[1][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][164] ( .G(n21), .D(idata[144]), .Q(\_zzLB[1][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][165] ( .G(n21), .D(idata[145]), .Q(\_zzLB[1][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][166] ( .G(n21), .D(idata[146]), .Q(\_zzLB[1][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][167] ( .G(n21), .D(idata[147]), .Q(\_zzLB[1][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][168] ( .G(n21), .D(idata[148]), .Q(\_zzLB[1][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][169] ( .G(n21), .D(idata[149]), .Q(\_zzLB[1][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][170] ( .G(n21), .D(idata[150]), .Q(\_zzLB[1][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][171] ( .G(n21), .D(idata[151]), .Q(\_zzLB[1][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][172] ( .G(n21), .D(idata[152]), .Q(\_zzLB[1][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][173] ( .G(n21), .D(idata[153]), .Q(\_zzLB[1][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][174] ( .G(n21), .D(idata[154]), .Q(\_zzLB[1][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][175] ( .G(n21), .D(idata[155]), .Q(\_zzLB[1][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][176] ( .G(n21), .D(idata[156]), .Q(\_zzLB[1][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][177] ( .G(n21), .D(idata[157]), .Q(\_zzLB[1][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][178] ( .G(n21), .D(idata[158]), .Q(\_zzLB[1][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][179] ( .G(n21), .D(idata[159]), .Q(\_zzLB[1][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][180] ( .G(n21), .D(idata[160]), .Q(\_zzLB[1][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][181] ( .G(n21), .D(idata[161]), .Q(\_zzLB[1][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][182] ( .G(n21), .D(idata[162]), .Q(\_zzLB[1][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][183] ( .G(n21), .D(idata[163]), .Q(\_zzLB[1][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][184] ( .G(n21), .D(idata[164]), .Q(\_zzLB[1][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][185] ( .G(n21), .D(idata[165]), .Q(\_zzLB[1][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][186] ( .G(n21), .D(idata[166]), .Q(\_zzLB[1][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][187] ( .G(n21), .D(idata[167]), .Q(\_zzLB[1][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][188] ( .G(n21), .D(idata[168]), .Q(\_zzLB[1][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][189] ( .G(n21), .D(idata[169]), .Q(\_zzLB[1][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][190] ( .G(n21), .D(idata[170]), .Q(\_zzLB[1][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][191] ( .G(n21), .D(idata[171]), .Q(\_zzLB[1][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][192] ( .G(n21), .D(idata[172]), .Q(\_zzLB[1][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][193] ( .G(n21), .D(idata[173]), .Q(\_zzLB[1][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][194] ( .G(n21), .D(idata[174]), .Q(\_zzLB[1][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][195] ( .G(n21), .D(idata[175]), .Q(\_zzLB[1][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][196] ( .G(n21), .D(idata[176]), .Q(\_zzLB[1][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][197] ( .G(n21), .D(idata[177]), .Q(\_zzLB[1][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][198] ( .G(n21), .D(idata[178]), .Q(\_zzLB[1][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][199] ( .G(n21), .D(idata[179]), .Q(\_zzLB[1][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][200] ( .G(n21), .D(idata[180]), .Q(\_zzLB[1][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][201] ( .G(n21), .D(idata[181]), .Q(\_zzLB[1][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][202] ( .G(n21), .D(idata[182]), .Q(\_zzLB[1][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][203] ( .G(n21), .D(idata[183]), .Q(\_zzLB[1][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][204] ( .G(n21), .D(idata[184]), .Q(\_zzLB[1][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][205] ( .G(n21), .D(idata[185]), .Q(\_zzLB[1][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][206] ( .G(n21), .D(idata[186]), .Q(\_zzLB[1][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][207] ( .G(n21), .D(idata[187]), .Q(\_zzLB[1][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][208] ( .G(n21), .D(idata[188]), .Q(\_zzLB[1][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][209] ( .G(n21), .D(idata[189]), .Q(\_zzLB[1][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][210] ( .G(n21), .D(idata[190]), .Q(\_zzLB[1][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][211] ( .G(n21), .D(idata[191]), .Q(\_zzLB[1][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][212] ( .G(n21), .D(idata[192]), .Q(\_zzLB[1][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][213] ( .G(n21), .D(idata[193]), .Q(\_zzLB[1][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][214] ( .G(n21), .D(idata[194]), .Q(\_zzLB[1][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][215] ( .G(n21), .D(idata[195]), .Q(\_zzLB[1][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][216] ( .G(n21), .D(idata[196]), .Q(\_zzLB[1][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][217] ( .G(n21), .D(idata[197]), .Q(\_zzLB[1][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][218] ( .G(n21), .D(idata[198]), .Q(\_zzLB[1][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][219] ( .G(n21), .D(idata[199]), .Q(\_zzLB[1][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][220] ( .G(n21), .D(idata[200]), .Q(\_zzLB[1][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][221] ( .G(n21), .D(idata[201]), .Q(\_zzLB[1][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][222] ( .G(n21), .D(idata[202]), .Q(\_zzLB[1][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][223] ( .G(n21), .D(idata[203]), .Q(\_zzLB[1][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][224] ( .G(n21), .D(idata[204]), .Q(\_zzLB[1][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][225] ( .G(n21), .D(idata[205]), .Q(\_zzLB[1][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][226] ( .G(n21), .D(idata[206]), .Q(\_zzLB[1][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][227] ( .G(n21), .D(idata[207]), .Q(\_zzLB[1][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][228] ( .G(n21), .D(idata[208]), .Q(\_zzLB[1][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][229] ( .G(n21), .D(idata[209]), .Q(\_zzLB[1][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][230] ( .G(n21), .D(idata[210]), .Q(\_zzLB[1][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][231] ( .G(n21), .D(idata[211]), .Q(\_zzLB[1][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][232] ( .G(n21), .D(idata[212]), .Q(\_zzLB[1][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][233] ( .G(n21), .D(idata[213]), .Q(\_zzLB[1][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][234] ( .G(n21), .D(idata[214]), .Q(\_zzLB[1][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][235] ( .G(n21), .D(idata[215]), .Q(\_zzLB[1][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][236] ( .G(n21), .D(idata[216]), .Q(\_zzLB[1][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][237] ( .G(n21), .D(idata[217]), .Q(\_zzLB[1][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][238] ( .G(n21), .D(idata[218]), .Q(\_zzLB[1][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][239] ( .G(n21), .D(idata[219]), .Q(\_zzLB[1][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][240] ( .G(n21), .D(idata[220]), .Q(\_zzLB[1][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][241] ( .G(n21), .D(idata[221]), .Q(\_zzLB[1][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][242] ( .G(n21), .D(idata[222]), .Q(\_zzLB[1][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][243] ( .G(n21), .D(idata[223]), .Q(\_zzLB[1][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][244] ( .G(n21), .D(idata[224]), .Q(\_zzLB[1][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][245] ( .G(n21), .D(idata[225]), .Q(\_zzLB[1][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][246] ( .G(n21), .D(idata[226]), .Q(\_zzLB[1][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][247] ( .G(n21), .D(idata[227]), .Q(\_zzLB[1][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][248] ( .G(n21), .D(idata[228]), .Q(\_zzLB[1][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][249] ( .G(n21), .D(idata[229]), .Q(\_zzLB[1][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][250] ( .G(n21), .D(idata[230]), .Q(\_zzLB[1][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][251] ( .G(n21), .D(idata[231]), .Q(\_zzLB[1][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][252] ( .G(n21), .D(idata[232]), .Q(\_zzLB[1][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][253] ( .G(n21), .D(idata[233]), .Q(\_zzLB[1][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][254] ( .G(n21), .D(idata[234]), .Q(\_zzLB[1][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][255] ( .G(n21), .D(idata[235]), .Q(\_zzLB[1][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][256] ( .G(n21), .D(idata[236]), .Q(\_zzLB[1][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][257] ( .G(n21), .D(idata[237]), .Q(\_zzLB[1][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][258] ( .G(n21), .D(idata[238]), .Q(\_zzLB[1][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][259] ( .G(n21), .D(idata[239]), .Q(\_zzLB[1][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][260] ( .G(n21), .D(idata[240]), .Q(\_zzLB[1][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][261] ( .G(n21), .D(idata[241]), .Q(\_zzLB[1][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][262] ( .G(n21), .D(idata[242]), .Q(\_zzLB[1][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][263] ( .G(n21), .D(idata[243]), .Q(\_zzLB[1][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][264] ( .G(n21), .D(idata[244]), .Q(\_zzLB[1][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][265] ( .G(n21), .D(idata[245]), .Q(\_zzLB[1][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][266] ( .G(n21), .D(idata[246]), .Q(\_zzLB[1][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][267] ( .G(n21), .D(idata[247]), .Q(\_zzLB[1][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][268] ( .G(n21), .D(idata[248]), .Q(\_zzLB[1][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][269] ( .G(n21), .D(idata[249]), .Q(\_zzLB[1][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][270] ( .G(n21), .D(idata[250]), .Q(\_zzLB[1][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][271] ( .G(n21), .D(idata[251]), .Q(\_zzLB[1][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][272] ( .G(n21), .D(idata[252]), .Q(\_zzLB[1][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][273] ( .G(n21), .D(idata[253]), .Q(\_zzLB[1][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][274] ( .G(n21), .D(idata[254]), .Q(\_zzLB[1][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][275] ( .G(n21), .D(idata[255]), .Q(\_zzLB[1][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][276] ( .G(n21), .D(idata[256]), .Q(\_zzLB[1][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][277] ( .G(n21), .D(idata[257]), .Q(\_zzLB[1][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][278] ( .G(n21), .D(idata[258]), .Q(\_zzLB[1][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][279] ( .G(n21), .D(idata[259]), .Q(\_zzLB[1][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][280] ( .G(n21), .D(idata[260]), .Q(\_zzLB[1][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][281] ( .G(n21), .D(idata[261]), .Q(\_zzLB[1][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][282] ( .G(n21), .D(idata[262]), .Q(\_zzLB[1][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][283] ( .G(n21), .D(idata[263]), .Q(\_zzLB[1][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][284] ( .G(n21), .D(idata[264]), .Q(\_zzLB[1][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][285] ( .G(n21), .D(idata[265]), .Q(\_zzLB[1][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][286] ( .G(n21), .D(idata[266]), .Q(\_zzLB[1][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][287] ( .G(n21), .D(idata[267]), .Q(\_zzLB[1][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][288] ( .G(n21), .D(idata[268]), .Q(\_zzLB[1][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][289] ( .G(n21), .D(idata[269]), .Q(\_zzLB[1][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][290] ( .G(n21), .D(idata[270]), .Q(\_zzLB[1][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][291] ( .G(n21), .D(idata[271]), .Q(\_zzLB[1][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][292] ( .G(n21), .D(idata[272]), .Q(\_zzLB[1][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][293] ( .G(n21), .D(idata[273]), .Q(\_zzLB[1][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][294] ( .G(n21), .D(idata[274]), .Q(\_zzLB[1][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][295] ( .G(n21), .D(idata[275]), .Q(\_zzLB[1][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][296] ( .G(n21), .D(idata[276]), .Q(\_zzLB[1][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][297] ( .G(n21), .D(idata[277]), .Q(\_zzLB[1][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][298] ( .G(n21), .D(idata[278]), .Q(\_zzLB[1][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][299] ( .G(n21), .D(idata[279]), .Q(\_zzLB[1][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[1][300] ( .G(n21), .D(ireq), .Q(\_zzLB[1][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][0] ( .G(n22), .D(cbid[0]), .Q(\_zzLB[2][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][1] ( .G(n22), .D(cbid[1]), .Q(\_zzLB[2][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][2] ( .G(n22), .D(cbid[2]), .Q(\_zzLB[2][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][3] ( .G(n22), .D(cbid[3]), .Q(\_zzLB[2][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][4] ( .G(n22), .D(cbid[4]), .Q(\_zzLB[2][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][5] ( .G(n22), .D(cbid[5]), .Q(\_zzLB[2][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][6] ( .G(n22), .D(cbid[6]), .Q(\_zzLB[2][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][7] ( .G(n22), .D(cbid[7]), .Q(\_zzLB[2][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][8] ( .G(n22), .D(cbid[8]), .Q(\_zzLB[2][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][9] ( .G(n22), .D(cbid[9]), .Q(\_zzLB[2][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][10] ( .G(n22), .D(cbid[10]), .Q(\_zzLB[2][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][11] ( .G(n22), .D(cbid[11]), .Q(\_zzLB[2][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][12] ( .G(n22), .D(cbid[12]), .Q(\_zzLB[2][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][13] ( .G(n22), .D(cbid[13]), .Q(\_zzLB[2][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][14] ( .G(n22), .D(cbid[14]), .Q(\_zzLB[2][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][15] ( .G(n22), .D(cbid[15]), .Q(\_zzLB[2][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][16] ( .G(n22), .D(cbid[16]), .Q(\_zzLB[2][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][17] ( .G(n22), .D(cbid[17]), .Q(\_zzLB[2][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][18] ( .G(n22), .D(cbid[18]), .Q(\_zzLB[2][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][19] ( .G(n22), .D(cbid[19]), .Q(\_zzLB[2][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][20] ( .G(n22), .D(idata[0]), .Q(\_zzLB[2][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][21] ( .G(n22), .D(idata[1]), .Q(\_zzLB[2][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][22] ( .G(n22), .D(idata[2]), .Q(\_zzLB[2][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][23] ( .G(n22), .D(idata[3]), .Q(\_zzLB[2][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][24] ( .G(n22), .D(idata[4]), .Q(\_zzLB[2][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][25] ( .G(n22), .D(idata[5]), .Q(\_zzLB[2][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][26] ( .G(n22), .D(idata[6]), .Q(\_zzLB[2][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][27] ( .G(n22), .D(idata[7]), .Q(\_zzLB[2][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][28] ( .G(n22), .D(idata[8]), .Q(\_zzLB[2][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][29] ( .G(n22), .D(idata[9]), .Q(\_zzLB[2][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][30] ( .G(n22), .D(idata[10]), .Q(\_zzLB[2][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][31] ( .G(n22), .D(idata[11]), .Q(\_zzLB[2][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][32] ( .G(n22), .D(idata[12]), .Q(\_zzLB[2][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][33] ( .G(n22), .D(idata[13]), .Q(\_zzLB[2][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][34] ( .G(n22), .D(idata[14]), .Q(\_zzLB[2][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][35] ( .G(n22), .D(idata[15]), .Q(\_zzLB[2][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][36] ( .G(n22), .D(idata[16]), .Q(\_zzLB[2][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][37] ( .G(n22), .D(idata[17]), .Q(\_zzLB[2][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][38] ( .G(n22), .D(idata[18]), .Q(\_zzLB[2][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][39] ( .G(n22), .D(idata[19]), .Q(\_zzLB[2][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][40] ( .G(n22), .D(idata[20]), .Q(\_zzLB[2][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][41] ( .G(n22), .D(idata[21]), .Q(\_zzLB[2][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][42] ( .G(n22), .D(idata[22]), .Q(\_zzLB[2][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][43] ( .G(n22), .D(idata[23]), .Q(\_zzLB[2][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][44] ( .G(n22), .D(idata[24]), .Q(\_zzLB[2][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][45] ( .G(n22), .D(idata[25]), .Q(\_zzLB[2][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][46] ( .G(n22), .D(idata[26]), .Q(\_zzLB[2][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][47] ( .G(n22), .D(idata[27]), .Q(\_zzLB[2][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][48] ( .G(n22), .D(idata[28]), .Q(\_zzLB[2][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][49] ( .G(n22), .D(idata[29]), .Q(\_zzLB[2][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][50] ( .G(n22), .D(idata[30]), .Q(\_zzLB[2][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][51] ( .G(n22), .D(idata[31]), .Q(\_zzLB[2][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][52] ( .G(n22), .D(idata[32]), .Q(\_zzLB[2][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][53] ( .G(n22), .D(idata[33]), .Q(\_zzLB[2][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][54] ( .G(n22), .D(idata[34]), .Q(\_zzLB[2][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][55] ( .G(n22), .D(idata[35]), .Q(\_zzLB[2][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][56] ( .G(n22), .D(idata[36]), .Q(\_zzLB[2][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][57] ( .G(n22), .D(idata[37]), .Q(\_zzLB[2][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][58] ( .G(n22), .D(idata[38]), .Q(\_zzLB[2][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][59] ( .G(n22), .D(idata[39]), .Q(\_zzLB[2][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][60] ( .G(n22), .D(idata[40]), .Q(\_zzLB[2][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][61] ( .G(n22), .D(idata[41]), .Q(\_zzLB[2][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][62] ( .G(n22), .D(idata[42]), .Q(\_zzLB[2][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][63] ( .G(n22), .D(idata[43]), .Q(\_zzLB[2][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][64] ( .G(n22), .D(idata[44]), .Q(\_zzLB[2][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][65] ( .G(n22), .D(idata[45]), .Q(\_zzLB[2][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][66] ( .G(n22), .D(idata[46]), .Q(\_zzLB[2][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][67] ( .G(n22), .D(idata[47]), .Q(\_zzLB[2][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][68] ( .G(n22), .D(idata[48]), .Q(\_zzLB[2][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][69] ( .G(n22), .D(idata[49]), .Q(\_zzLB[2][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][70] ( .G(n22), .D(idata[50]), .Q(\_zzLB[2][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][71] ( .G(n22), .D(idata[51]), .Q(\_zzLB[2][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][72] ( .G(n22), .D(idata[52]), .Q(\_zzLB[2][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][73] ( .G(n22), .D(idata[53]), .Q(\_zzLB[2][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][74] ( .G(n22), .D(idata[54]), .Q(\_zzLB[2][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][75] ( .G(n22), .D(idata[55]), .Q(\_zzLB[2][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][76] ( .G(n22), .D(idata[56]), .Q(\_zzLB[2][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][77] ( .G(n22), .D(idata[57]), .Q(\_zzLB[2][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][78] ( .G(n22), .D(idata[58]), .Q(\_zzLB[2][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][79] ( .G(n22), .D(idata[59]), .Q(\_zzLB[2][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][80] ( .G(n22), .D(idata[60]), .Q(\_zzLB[2][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][81] ( .G(n22), .D(idata[61]), .Q(\_zzLB[2][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][82] ( .G(n22), .D(idata[62]), .Q(\_zzLB[2][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][83] ( .G(n22), .D(idata[63]), .Q(\_zzLB[2][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][84] ( .G(n22), .D(idata[64]), .Q(\_zzLB[2][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][85] ( .G(n22), .D(idata[65]), .Q(\_zzLB[2][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][86] ( .G(n22), .D(idata[66]), .Q(\_zzLB[2][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][87] ( .G(n22), .D(idata[67]), .Q(\_zzLB[2][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][88] ( .G(n22), .D(idata[68]), .Q(\_zzLB[2][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][89] ( .G(n22), .D(idata[69]), .Q(\_zzLB[2][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][90] ( .G(n22), .D(idata[70]), .Q(\_zzLB[2][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][91] ( .G(n22), .D(idata[71]), .Q(\_zzLB[2][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][92] ( .G(n22), .D(idata[72]), .Q(\_zzLB[2][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][93] ( .G(n22), .D(idata[73]), .Q(\_zzLB[2][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][94] ( .G(n22), .D(idata[74]), .Q(\_zzLB[2][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][95] ( .G(n22), .D(idata[75]), .Q(\_zzLB[2][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][96] ( .G(n22), .D(idata[76]), .Q(\_zzLB[2][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][97] ( .G(n22), .D(idata[77]), .Q(\_zzLB[2][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][98] ( .G(n22), .D(idata[78]), .Q(\_zzLB[2][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][99] ( .G(n22), .D(idata[79]), .Q(\_zzLB[2][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][100] ( .G(n22), .D(idata[80]), .Q(\_zzLB[2][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][101] ( .G(n22), .D(idata[81]), .Q(\_zzLB[2][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][102] ( .G(n22), .D(idata[82]), .Q(\_zzLB[2][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][103] ( .G(n22), .D(idata[83]), .Q(\_zzLB[2][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][104] ( .G(n22), .D(idata[84]), .Q(\_zzLB[2][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][105] ( .G(n22), .D(idata[85]), .Q(\_zzLB[2][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][106] ( .G(n22), .D(idata[86]), .Q(\_zzLB[2][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][107] ( .G(n22), .D(idata[87]), .Q(\_zzLB[2][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][108] ( .G(n22), .D(idata[88]), .Q(\_zzLB[2][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][109] ( .G(n22), .D(idata[89]), .Q(\_zzLB[2][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][110] ( .G(n22), .D(idata[90]), .Q(\_zzLB[2][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][111] ( .G(n22), .D(idata[91]), .Q(\_zzLB[2][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][112] ( .G(n22), .D(idata[92]), .Q(\_zzLB[2][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][113] ( .G(n22), .D(idata[93]), .Q(\_zzLB[2][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][114] ( .G(n22), .D(idata[94]), .Q(\_zzLB[2][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][115] ( .G(n22), .D(idata[95]), .Q(\_zzLB[2][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][116] ( .G(n22), .D(idata[96]), .Q(\_zzLB[2][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][117] ( .G(n22), .D(idata[97]), .Q(\_zzLB[2][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][118] ( .G(n22), .D(idata[98]), .Q(\_zzLB[2][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][119] ( .G(n22), .D(idata[99]), .Q(\_zzLB[2][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][120] ( .G(n22), .D(idata[100]), .Q(\_zzLB[2][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][121] ( .G(n22), .D(idata[101]), .Q(\_zzLB[2][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][122] ( .G(n22), .D(idata[102]), .Q(\_zzLB[2][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][123] ( .G(n22), .D(idata[103]), .Q(\_zzLB[2][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][124] ( .G(n22), .D(idata[104]), .Q(\_zzLB[2][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][125] ( .G(n22), .D(idata[105]), .Q(\_zzLB[2][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][126] ( .G(n22), .D(idata[106]), .Q(\_zzLB[2][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][127] ( .G(n22), .D(idata[107]), .Q(\_zzLB[2][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][128] ( .G(n22), .D(idata[108]), .Q(\_zzLB[2][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][129] ( .G(n22), .D(idata[109]), .Q(\_zzLB[2][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][130] ( .G(n22), .D(idata[110]), .Q(\_zzLB[2][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][131] ( .G(n22), .D(idata[111]), .Q(\_zzLB[2][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][132] ( .G(n22), .D(idata[112]), .Q(\_zzLB[2][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][133] ( .G(n22), .D(idata[113]), .Q(\_zzLB[2][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][134] ( .G(n22), .D(idata[114]), .Q(\_zzLB[2][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][135] ( .G(n22), .D(idata[115]), .Q(\_zzLB[2][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][136] ( .G(n22), .D(idata[116]), .Q(\_zzLB[2][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][137] ( .G(n22), .D(idata[117]), .Q(\_zzLB[2][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][138] ( .G(n22), .D(idata[118]), .Q(\_zzLB[2][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][139] ( .G(n22), .D(idata[119]), .Q(\_zzLB[2][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][140] ( .G(n22), .D(idata[120]), .Q(\_zzLB[2][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][141] ( .G(n22), .D(idata[121]), .Q(\_zzLB[2][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][142] ( .G(n22), .D(idata[122]), .Q(\_zzLB[2][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][143] ( .G(n22), .D(idata[123]), .Q(\_zzLB[2][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][144] ( .G(n22), .D(idata[124]), .Q(\_zzLB[2][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][145] ( .G(n22), .D(idata[125]), .Q(\_zzLB[2][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][146] ( .G(n22), .D(idata[126]), .Q(\_zzLB[2][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][147] ( .G(n22), .D(idata[127]), .Q(\_zzLB[2][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][148] ( .G(n22), .D(idata[128]), .Q(\_zzLB[2][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][149] ( .G(n22), .D(idata[129]), .Q(\_zzLB[2][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][150] ( .G(n22), .D(idata[130]), .Q(\_zzLB[2][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][151] ( .G(n22), .D(idata[131]), .Q(\_zzLB[2][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][152] ( .G(n22), .D(idata[132]), .Q(\_zzLB[2][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][153] ( .G(n22), .D(idata[133]), .Q(\_zzLB[2][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][154] ( .G(n22), .D(idata[134]), .Q(\_zzLB[2][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][155] ( .G(n22), .D(idata[135]), .Q(\_zzLB[2][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][156] ( .G(n22), .D(idata[136]), .Q(\_zzLB[2][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][157] ( .G(n22), .D(idata[137]), .Q(\_zzLB[2][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][158] ( .G(n22), .D(idata[138]), .Q(\_zzLB[2][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][159] ( .G(n22), .D(idata[139]), .Q(\_zzLB[2][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][160] ( .G(n22), .D(idata[140]), .Q(\_zzLB[2][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][161] ( .G(n22), .D(idata[141]), .Q(\_zzLB[2][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][162] ( .G(n22), .D(idata[142]), .Q(\_zzLB[2][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][163] ( .G(n22), .D(idata[143]), .Q(\_zzLB[2][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][164] ( .G(n22), .D(idata[144]), .Q(\_zzLB[2][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][165] ( .G(n22), .D(idata[145]), .Q(\_zzLB[2][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][166] ( .G(n22), .D(idata[146]), .Q(\_zzLB[2][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][167] ( .G(n22), .D(idata[147]), .Q(\_zzLB[2][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][168] ( .G(n22), .D(idata[148]), .Q(\_zzLB[2][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][169] ( .G(n22), .D(idata[149]), .Q(\_zzLB[2][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][170] ( .G(n22), .D(idata[150]), .Q(\_zzLB[2][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][171] ( .G(n22), .D(idata[151]), .Q(\_zzLB[2][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][172] ( .G(n22), .D(idata[152]), .Q(\_zzLB[2][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][173] ( .G(n22), .D(idata[153]), .Q(\_zzLB[2][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][174] ( .G(n22), .D(idata[154]), .Q(\_zzLB[2][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][175] ( .G(n22), .D(idata[155]), .Q(\_zzLB[2][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][176] ( .G(n22), .D(idata[156]), .Q(\_zzLB[2][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][177] ( .G(n22), .D(idata[157]), .Q(\_zzLB[2][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][178] ( .G(n22), .D(idata[158]), .Q(\_zzLB[2][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][179] ( .G(n22), .D(idata[159]), .Q(\_zzLB[2][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][180] ( .G(n22), .D(idata[160]), .Q(\_zzLB[2][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][181] ( .G(n22), .D(idata[161]), .Q(\_zzLB[2][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][182] ( .G(n22), .D(idata[162]), .Q(\_zzLB[2][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][183] ( .G(n22), .D(idata[163]), .Q(\_zzLB[2][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][184] ( .G(n22), .D(idata[164]), .Q(\_zzLB[2][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][185] ( .G(n22), .D(idata[165]), .Q(\_zzLB[2][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][186] ( .G(n22), .D(idata[166]), .Q(\_zzLB[2][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][187] ( .G(n22), .D(idata[167]), .Q(\_zzLB[2][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][188] ( .G(n22), .D(idata[168]), .Q(\_zzLB[2][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][189] ( .G(n22), .D(idata[169]), .Q(\_zzLB[2][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][190] ( .G(n22), .D(idata[170]), .Q(\_zzLB[2][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][191] ( .G(n22), .D(idata[171]), .Q(\_zzLB[2][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][192] ( .G(n22), .D(idata[172]), .Q(\_zzLB[2][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][193] ( .G(n22), .D(idata[173]), .Q(\_zzLB[2][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][194] ( .G(n22), .D(idata[174]), .Q(\_zzLB[2][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][195] ( .G(n22), .D(idata[175]), .Q(\_zzLB[2][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][196] ( .G(n22), .D(idata[176]), .Q(\_zzLB[2][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][197] ( .G(n22), .D(idata[177]), .Q(\_zzLB[2][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][198] ( .G(n22), .D(idata[178]), .Q(\_zzLB[2][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][199] ( .G(n22), .D(idata[179]), .Q(\_zzLB[2][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][200] ( .G(n22), .D(idata[180]), .Q(\_zzLB[2][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][201] ( .G(n22), .D(idata[181]), .Q(\_zzLB[2][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][202] ( .G(n22), .D(idata[182]), .Q(\_zzLB[2][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][203] ( .G(n22), .D(idata[183]), .Q(\_zzLB[2][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][204] ( .G(n22), .D(idata[184]), .Q(\_zzLB[2][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][205] ( .G(n22), .D(idata[185]), .Q(\_zzLB[2][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][206] ( .G(n22), .D(idata[186]), .Q(\_zzLB[2][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][207] ( .G(n22), .D(idata[187]), .Q(\_zzLB[2][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][208] ( .G(n22), .D(idata[188]), .Q(\_zzLB[2][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][209] ( .G(n22), .D(idata[189]), .Q(\_zzLB[2][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][210] ( .G(n22), .D(idata[190]), .Q(\_zzLB[2][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][211] ( .G(n22), .D(idata[191]), .Q(\_zzLB[2][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][212] ( .G(n22), .D(idata[192]), .Q(\_zzLB[2][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][213] ( .G(n22), .D(idata[193]), .Q(\_zzLB[2][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][214] ( .G(n22), .D(idata[194]), .Q(\_zzLB[2][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][215] ( .G(n22), .D(idata[195]), .Q(\_zzLB[2][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][216] ( .G(n22), .D(idata[196]), .Q(\_zzLB[2][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][217] ( .G(n22), .D(idata[197]), .Q(\_zzLB[2][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][218] ( .G(n22), .D(idata[198]), .Q(\_zzLB[2][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][219] ( .G(n22), .D(idata[199]), .Q(\_zzLB[2][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][220] ( .G(n22), .D(idata[200]), .Q(\_zzLB[2][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][221] ( .G(n22), .D(idata[201]), .Q(\_zzLB[2][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][222] ( .G(n22), .D(idata[202]), .Q(\_zzLB[2][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][223] ( .G(n22), .D(idata[203]), .Q(\_zzLB[2][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][224] ( .G(n22), .D(idata[204]), .Q(\_zzLB[2][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][225] ( .G(n22), .D(idata[205]), .Q(\_zzLB[2][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][226] ( .G(n22), .D(idata[206]), .Q(\_zzLB[2][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][227] ( .G(n22), .D(idata[207]), .Q(\_zzLB[2][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][228] ( .G(n22), .D(idata[208]), .Q(\_zzLB[2][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][229] ( .G(n22), .D(idata[209]), .Q(\_zzLB[2][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][230] ( .G(n22), .D(idata[210]), .Q(\_zzLB[2][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][231] ( .G(n22), .D(idata[211]), .Q(\_zzLB[2][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][232] ( .G(n22), .D(idata[212]), .Q(\_zzLB[2][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][233] ( .G(n22), .D(idata[213]), .Q(\_zzLB[2][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][234] ( .G(n22), .D(idata[214]), .Q(\_zzLB[2][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][235] ( .G(n22), .D(idata[215]), .Q(\_zzLB[2][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][236] ( .G(n22), .D(idata[216]), .Q(\_zzLB[2][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][237] ( .G(n22), .D(idata[217]), .Q(\_zzLB[2][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][238] ( .G(n22), .D(idata[218]), .Q(\_zzLB[2][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][239] ( .G(n22), .D(idata[219]), .Q(\_zzLB[2][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][240] ( .G(n22), .D(idata[220]), .Q(\_zzLB[2][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][241] ( .G(n22), .D(idata[221]), .Q(\_zzLB[2][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][242] ( .G(n22), .D(idata[222]), .Q(\_zzLB[2][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][243] ( .G(n22), .D(idata[223]), .Q(\_zzLB[2][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][244] ( .G(n22), .D(idata[224]), .Q(\_zzLB[2][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][245] ( .G(n22), .D(idata[225]), .Q(\_zzLB[2][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][246] ( .G(n22), .D(idata[226]), .Q(\_zzLB[2][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][247] ( .G(n22), .D(idata[227]), .Q(\_zzLB[2][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][248] ( .G(n22), .D(idata[228]), .Q(\_zzLB[2][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][249] ( .G(n22), .D(idata[229]), .Q(\_zzLB[2][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][250] ( .G(n22), .D(idata[230]), .Q(\_zzLB[2][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][251] ( .G(n22), .D(idata[231]), .Q(\_zzLB[2][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][252] ( .G(n22), .D(idata[232]), .Q(\_zzLB[2][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][253] ( .G(n22), .D(idata[233]), .Q(\_zzLB[2][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][254] ( .G(n22), .D(idata[234]), .Q(\_zzLB[2][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][255] ( .G(n22), .D(idata[235]), .Q(\_zzLB[2][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][256] ( .G(n22), .D(idata[236]), .Q(\_zzLB[2][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][257] ( .G(n22), .D(idata[237]), .Q(\_zzLB[2][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][258] ( .G(n22), .D(idata[238]), .Q(\_zzLB[2][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][259] ( .G(n22), .D(idata[239]), .Q(\_zzLB[2][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][260] ( .G(n22), .D(idata[240]), .Q(\_zzLB[2][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][261] ( .G(n22), .D(idata[241]), .Q(\_zzLB[2][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][262] ( .G(n22), .D(idata[242]), .Q(\_zzLB[2][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][263] ( .G(n22), .D(idata[243]), .Q(\_zzLB[2][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][264] ( .G(n22), .D(idata[244]), .Q(\_zzLB[2][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][265] ( .G(n22), .D(idata[245]), .Q(\_zzLB[2][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][266] ( .G(n22), .D(idata[246]), .Q(\_zzLB[2][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][267] ( .G(n22), .D(idata[247]), .Q(\_zzLB[2][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][268] ( .G(n22), .D(idata[248]), .Q(\_zzLB[2][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][269] ( .G(n22), .D(idata[249]), .Q(\_zzLB[2][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][270] ( .G(n22), .D(idata[250]), .Q(\_zzLB[2][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][271] ( .G(n22), .D(idata[251]), .Q(\_zzLB[2][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][272] ( .G(n22), .D(idata[252]), .Q(\_zzLB[2][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][273] ( .G(n22), .D(idata[253]), .Q(\_zzLB[2][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][274] ( .G(n22), .D(idata[254]), .Q(\_zzLB[2][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][275] ( .G(n22), .D(idata[255]), .Q(\_zzLB[2][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][276] ( .G(n22), .D(idata[256]), .Q(\_zzLB[2][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][277] ( .G(n22), .D(idata[257]), .Q(\_zzLB[2][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][278] ( .G(n22), .D(idata[258]), .Q(\_zzLB[2][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][279] ( .G(n22), .D(idata[259]), .Q(\_zzLB[2][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][280] ( .G(n22), .D(idata[260]), .Q(\_zzLB[2][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][281] ( .G(n22), .D(idata[261]), .Q(\_zzLB[2][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][282] ( .G(n22), .D(idata[262]), .Q(\_zzLB[2][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][283] ( .G(n22), .D(idata[263]), .Q(\_zzLB[2][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][284] ( .G(n22), .D(idata[264]), .Q(\_zzLB[2][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][285] ( .G(n22), .D(idata[265]), .Q(\_zzLB[2][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][286] ( .G(n22), .D(idata[266]), .Q(\_zzLB[2][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][287] ( .G(n22), .D(idata[267]), .Q(\_zzLB[2][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][288] ( .G(n22), .D(idata[268]), .Q(\_zzLB[2][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][289] ( .G(n22), .D(idata[269]), .Q(\_zzLB[2][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][290] ( .G(n22), .D(idata[270]), .Q(\_zzLB[2][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][291] ( .G(n22), .D(idata[271]), .Q(\_zzLB[2][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][292] ( .G(n22), .D(idata[272]), .Q(\_zzLB[2][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][293] ( .G(n22), .D(idata[273]), .Q(\_zzLB[2][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][294] ( .G(n22), .D(idata[274]), .Q(\_zzLB[2][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][295] ( .G(n22), .D(idata[275]), .Q(\_zzLB[2][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][296] ( .G(n22), .D(idata[276]), .Q(\_zzLB[2][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][297] ( .G(n22), .D(idata[277]), .Q(\_zzLB[2][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][298] ( .G(n22), .D(idata[278]), .Q(\_zzLB[2][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][299] ( .G(n22), .D(idata[279]), .Q(\_zzLB[2][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[2][300] ( .G(n22), .D(ireq), .Q(\_zzLB[2][300] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][0] ( .G(n23), .D(cbid[0]), .Q(\_zzLB[3][0] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][1] ( .G(n23), .D(cbid[1]), .Q(\_zzLB[3][1] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][2] ( .G(n23), .D(cbid[2]), .Q(\_zzLB[3][2] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][3] ( .G(n23), .D(cbid[3]), .Q(\_zzLB[3][3] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][4] ( .G(n23), .D(cbid[4]), .Q(\_zzLB[3][4] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][5] ( .G(n23), .D(cbid[5]), .Q(\_zzLB[3][5] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][6] ( .G(n23), .D(cbid[6]), .Q(\_zzLB[3][6] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][7] ( .G(n23), .D(cbid[7]), .Q(\_zzLB[3][7] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][8] ( .G(n23), .D(cbid[8]), .Q(\_zzLB[3][8] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][9] ( .G(n23), .D(cbid[9]), .Q(\_zzLB[3][9] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][10] ( .G(n23), .D(cbid[10]), .Q(\_zzLB[3][10] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][11] ( .G(n23), .D(cbid[11]), .Q(\_zzLB[3][11] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][12] ( .G(n23), .D(cbid[12]), .Q(\_zzLB[3][12] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][13] ( .G(n23), .D(cbid[13]), .Q(\_zzLB[3][13] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][14] ( .G(n23), .D(cbid[14]), .Q(\_zzLB[3][14] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][15] ( .G(n23), .D(cbid[15]), .Q(\_zzLB[3][15] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][16] ( .G(n23), .D(cbid[16]), .Q(\_zzLB[3][16] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][17] ( .G(n23), .D(cbid[17]), .Q(\_zzLB[3][17] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][18] ( .G(n23), .D(cbid[18]), .Q(\_zzLB[3][18] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][19] ( .G(n23), .D(cbid[19]), .Q(\_zzLB[3][19] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][20] ( .G(n23), .D(idata[0]), .Q(\_zzLB[3][20] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][21] ( .G(n23), .D(idata[1]), .Q(\_zzLB[3][21] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][22] ( .G(n23), .D(idata[2]), .Q(\_zzLB[3][22] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][23] ( .G(n23), .D(idata[3]), .Q(\_zzLB[3][23] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][24] ( .G(n23), .D(idata[4]), .Q(\_zzLB[3][24] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][25] ( .G(n23), .D(idata[5]), .Q(\_zzLB[3][25] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][26] ( .G(n23), .D(idata[6]), .Q(\_zzLB[3][26] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][27] ( .G(n23), .D(idata[7]), .Q(\_zzLB[3][27] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][28] ( .G(n23), .D(idata[8]), .Q(\_zzLB[3][28] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][29] ( .G(n23), .D(idata[9]), .Q(\_zzLB[3][29] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][30] ( .G(n23), .D(idata[10]), .Q(\_zzLB[3][30] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][31] ( .G(n23), .D(idata[11]), .Q(\_zzLB[3][31] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][32] ( .G(n23), .D(idata[12]), .Q(\_zzLB[3][32] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][33] ( .G(n23), .D(idata[13]), .Q(\_zzLB[3][33] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][34] ( .G(n23), .D(idata[14]), .Q(\_zzLB[3][34] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][35] ( .G(n23), .D(idata[15]), .Q(\_zzLB[3][35] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][36] ( .G(n23), .D(idata[16]), .Q(\_zzLB[3][36] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][37] ( .G(n23), .D(idata[17]), .Q(\_zzLB[3][37] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][38] ( .G(n23), .D(idata[18]), .Q(\_zzLB[3][38] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][39] ( .G(n23), .D(idata[19]), .Q(\_zzLB[3][39] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][40] ( .G(n23), .D(idata[20]), .Q(\_zzLB[3][40] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][41] ( .G(n23), .D(idata[21]), .Q(\_zzLB[3][41] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][42] ( .G(n23), .D(idata[22]), .Q(\_zzLB[3][42] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][43] ( .G(n23), .D(idata[23]), .Q(\_zzLB[3][43] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][44] ( .G(n23), .D(idata[24]), .Q(\_zzLB[3][44] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][45] ( .G(n23), .D(idata[25]), .Q(\_zzLB[3][45] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][46] ( .G(n23), .D(idata[26]), .Q(\_zzLB[3][46] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][47] ( .G(n23), .D(idata[27]), .Q(\_zzLB[3][47] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][48] ( .G(n23), .D(idata[28]), .Q(\_zzLB[3][48] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][49] ( .G(n23), .D(idata[29]), .Q(\_zzLB[3][49] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][50] ( .G(n23), .D(idata[30]), .Q(\_zzLB[3][50] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][51] ( .G(n23), .D(idata[31]), .Q(\_zzLB[3][51] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][52] ( .G(n23), .D(idata[32]), .Q(\_zzLB[3][52] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][53] ( .G(n23), .D(idata[33]), .Q(\_zzLB[3][53] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][54] ( .G(n23), .D(idata[34]), .Q(\_zzLB[3][54] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][55] ( .G(n23), .D(idata[35]), .Q(\_zzLB[3][55] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][56] ( .G(n23), .D(idata[36]), .Q(\_zzLB[3][56] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][57] ( .G(n23), .D(idata[37]), .Q(\_zzLB[3][57] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][58] ( .G(n23), .D(idata[38]), .Q(\_zzLB[3][58] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][59] ( .G(n23), .D(idata[39]), .Q(\_zzLB[3][59] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][60] ( .G(n23), .D(idata[40]), .Q(\_zzLB[3][60] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][61] ( .G(n23), .D(idata[41]), .Q(\_zzLB[3][61] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][62] ( .G(n23), .D(idata[42]), .Q(\_zzLB[3][62] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][63] ( .G(n23), .D(idata[43]), .Q(\_zzLB[3][63] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][64] ( .G(n23), .D(idata[44]), .Q(\_zzLB[3][64] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][65] ( .G(n23), .D(idata[45]), .Q(\_zzLB[3][65] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][66] ( .G(n23), .D(idata[46]), .Q(\_zzLB[3][66] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][67] ( .G(n23), .D(idata[47]), .Q(\_zzLB[3][67] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][68] ( .G(n23), .D(idata[48]), .Q(\_zzLB[3][68] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][69] ( .G(n23), .D(idata[49]), .Q(\_zzLB[3][69] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][70] ( .G(n23), .D(idata[50]), .Q(\_zzLB[3][70] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][71] ( .G(n23), .D(idata[51]), .Q(\_zzLB[3][71] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][72] ( .G(n23), .D(idata[52]), .Q(\_zzLB[3][72] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][73] ( .G(n23), .D(idata[53]), .Q(\_zzLB[3][73] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][74] ( .G(n23), .D(idata[54]), .Q(\_zzLB[3][74] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][75] ( .G(n23), .D(idata[55]), .Q(\_zzLB[3][75] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][76] ( .G(n23), .D(idata[56]), .Q(\_zzLB[3][76] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][77] ( .G(n23), .D(idata[57]), .Q(\_zzLB[3][77] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][78] ( .G(n23), .D(idata[58]), .Q(\_zzLB[3][78] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][79] ( .G(n23), .D(idata[59]), .Q(\_zzLB[3][79] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][80] ( .G(n23), .D(idata[60]), .Q(\_zzLB[3][80] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][81] ( .G(n23), .D(idata[61]), .Q(\_zzLB[3][81] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][82] ( .G(n23), .D(idata[62]), .Q(\_zzLB[3][82] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][83] ( .G(n23), .D(idata[63]), .Q(\_zzLB[3][83] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][84] ( .G(n23), .D(idata[64]), .Q(\_zzLB[3][84] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][85] ( .G(n23), .D(idata[65]), .Q(\_zzLB[3][85] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][86] ( .G(n23), .D(idata[66]), .Q(\_zzLB[3][86] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][87] ( .G(n23), .D(idata[67]), .Q(\_zzLB[3][87] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][88] ( .G(n23), .D(idata[68]), .Q(\_zzLB[3][88] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][89] ( .G(n23), .D(idata[69]), .Q(\_zzLB[3][89] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][90] ( .G(n23), .D(idata[70]), .Q(\_zzLB[3][90] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][91] ( .G(n23), .D(idata[71]), .Q(\_zzLB[3][91] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][92] ( .G(n23), .D(idata[72]), .Q(\_zzLB[3][92] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][93] ( .G(n23), .D(idata[73]), .Q(\_zzLB[3][93] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][94] ( .G(n23), .D(idata[74]), .Q(\_zzLB[3][94] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][95] ( .G(n23), .D(idata[75]), .Q(\_zzLB[3][95] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][96] ( .G(n23), .D(idata[76]), .Q(\_zzLB[3][96] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][97] ( .G(n23), .D(idata[77]), .Q(\_zzLB[3][97] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][98] ( .G(n23), .D(idata[78]), .Q(\_zzLB[3][98] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][99] ( .G(n23), .D(idata[79]), .Q(\_zzLB[3][99] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][100] ( .G(n23), .D(idata[80]), .Q(\_zzLB[3][100] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][101] ( .G(n23), .D(idata[81]), .Q(\_zzLB[3][101] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][102] ( .G(n23), .D(idata[82]), .Q(\_zzLB[3][102] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][103] ( .G(n23), .D(idata[83]), .Q(\_zzLB[3][103] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][104] ( .G(n23), .D(idata[84]), .Q(\_zzLB[3][104] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][105] ( .G(n23), .D(idata[85]), .Q(\_zzLB[3][105] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][106] ( .G(n23), .D(idata[86]), .Q(\_zzLB[3][106] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][107] ( .G(n23), .D(idata[87]), .Q(\_zzLB[3][107] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][108] ( .G(n23), .D(idata[88]), .Q(\_zzLB[3][108] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][109] ( .G(n23), .D(idata[89]), .Q(\_zzLB[3][109] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][110] ( .G(n23), .D(idata[90]), .Q(\_zzLB[3][110] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][111] ( .G(n23), .D(idata[91]), .Q(\_zzLB[3][111] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][112] ( .G(n23), .D(idata[92]), .Q(\_zzLB[3][112] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][113] ( .G(n23), .D(idata[93]), .Q(\_zzLB[3][113] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][114] ( .G(n23), .D(idata[94]), .Q(\_zzLB[3][114] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][115] ( .G(n23), .D(idata[95]), .Q(\_zzLB[3][115] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][116] ( .G(n23), .D(idata[96]), .Q(\_zzLB[3][116] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][117] ( .G(n23), .D(idata[97]), .Q(\_zzLB[3][117] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][118] ( .G(n23), .D(idata[98]), .Q(\_zzLB[3][118] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][119] ( .G(n23), .D(idata[99]), .Q(\_zzLB[3][119] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][120] ( .G(n23), .D(idata[100]), .Q(\_zzLB[3][120] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][121] ( .G(n23), .D(idata[101]), .Q(\_zzLB[3][121] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][122] ( .G(n23), .D(idata[102]), .Q(\_zzLB[3][122] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][123] ( .G(n23), .D(idata[103]), .Q(\_zzLB[3][123] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][124] ( .G(n23), .D(idata[104]), .Q(\_zzLB[3][124] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][125] ( .G(n23), .D(idata[105]), .Q(\_zzLB[3][125] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][126] ( .G(n23), .D(idata[106]), .Q(\_zzLB[3][126] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][127] ( .G(n23), .D(idata[107]), .Q(\_zzLB[3][127] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][128] ( .G(n23), .D(idata[108]), .Q(\_zzLB[3][128] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][129] ( .G(n23), .D(idata[109]), .Q(\_zzLB[3][129] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][130] ( .G(n23), .D(idata[110]), .Q(\_zzLB[3][130] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][131] ( .G(n23), .D(idata[111]), .Q(\_zzLB[3][131] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][132] ( .G(n23), .D(idata[112]), .Q(\_zzLB[3][132] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][133] ( .G(n23), .D(idata[113]), .Q(\_zzLB[3][133] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][134] ( .G(n23), .D(idata[114]), .Q(\_zzLB[3][134] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][135] ( .G(n23), .D(idata[115]), .Q(\_zzLB[3][135] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][136] ( .G(n23), .D(idata[116]), .Q(\_zzLB[3][136] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][137] ( .G(n23), .D(idata[117]), .Q(\_zzLB[3][137] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][138] ( .G(n23), .D(idata[118]), .Q(\_zzLB[3][138] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][139] ( .G(n23), .D(idata[119]), .Q(\_zzLB[3][139] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][140] ( .G(n23), .D(idata[120]), .Q(\_zzLB[3][140] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][141] ( .G(n23), .D(idata[121]), .Q(\_zzLB[3][141] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][142] ( .G(n23), .D(idata[122]), .Q(\_zzLB[3][142] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][143] ( .G(n23), .D(idata[123]), .Q(\_zzLB[3][143] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][144] ( .G(n23), .D(idata[124]), .Q(\_zzLB[3][144] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][145] ( .G(n23), .D(idata[125]), .Q(\_zzLB[3][145] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][146] ( .G(n23), .D(idata[126]), .Q(\_zzLB[3][146] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][147] ( .G(n23), .D(idata[127]), .Q(\_zzLB[3][147] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][148] ( .G(n23), .D(idata[128]), .Q(\_zzLB[3][148] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][149] ( .G(n23), .D(idata[129]), .Q(\_zzLB[3][149] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][150] ( .G(n23), .D(idata[130]), .Q(\_zzLB[3][150] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][151] ( .G(n23), .D(idata[131]), .Q(\_zzLB[3][151] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][152] ( .G(n23), .D(idata[132]), .Q(\_zzLB[3][152] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][153] ( .G(n23), .D(idata[133]), .Q(\_zzLB[3][153] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][154] ( .G(n23), .D(idata[134]), .Q(\_zzLB[3][154] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][155] ( .G(n23), .D(idata[135]), .Q(\_zzLB[3][155] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][156] ( .G(n23), .D(idata[136]), .Q(\_zzLB[3][156] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][157] ( .G(n23), .D(idata[137]), .Q(\_zzLB[3][157] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][158] ( .G(n23), .D(idata[138]), .Q(\_zzLB[3][158] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][159] ( .G(n23), .D(idata[139]), .Q(\_zzLB[3][159] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][160] ( .G(n23), .D(idata[140]), .Q(\_zzLB[3][160] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][161] ( .G(n23), .D(idata[141]), .Q(\_zzLB[3][161] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][162] ( .G(n23), .D(idata[142]), .Q(\_zzLB[3][162] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][163] ( .G(n23), .D(idata[143]), .Q(\_zzLB[3][163] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][164] ( .G(n23), .D(idata[144]), .Q(\_zzLB[3][164] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][165] ( .G(n23), .D(idata[145]), .Q(\_zzLB[3][165] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][166] ( .G(n23), .D(idata[146]), .Q(\_zzLB[3][166] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][167] ( .G(n23), .D(idata[147]), .Q(\_zzLB[3][167] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][168] ( .G(n23), .D(idata[148]), .Q(\_zzLB[3][168] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][169] ( .G(n23), .D(idata[149]), .Q(\_zzLB[3][169] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][170] ( .G(n23), .D(idata[150]), .Q(\_zzLB[3][170] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][171] ( .G(n23), .D(idata[151]), .Q(\_zzLB[3][171] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][172] ( .G(n23), .D(idata[152]), .Q(\_zzLB[3][172] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][173] ( .G(n23), .D(idata[153]), .Q(\_zzLB[3][173] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][174] ( .G(n23), .D(idata[154]), .Q(\_zzLB[3][174] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][175] ( .G(n23), .D(idata[155]), .Q(\_zzLB[3][175] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][176] ( .G(n23), .D(idata[156]), .Q(\_zzLB[3][176] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][177] ( .G(n23), .D(idata[157]), .Q(\_zzLB[3][177] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][178] ( .G(n23), .D(idata[158]), .Q(\_zzLB[3][178] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][179] ( .G(n23), .D(idata[159]), .Q(\_zzLB[3][179] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][180] ( .G(n23), .D(idata[160]), .Q(\_zzLB[3][180] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][181] ( .G(n23), .D(idata[161]), .Q(\_zzLB[3][181] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][182] ( .G(n23), .D(idata[162]), .Q(\_zzLB[3][182] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][183] ( .G(n23), .D(idata[163]), .Q(\_zzLB[3][183] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][184] ( .G(n23), .D(idata[164]), .Q(\_zzLB[3][184] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][185] ( .G(n23), .D(idata[165]), .Q(\_zzLB[3][185] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][186] ( .G(n23), .D(idata[166]), .Q(\_zzLB[3][186] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][187] ( .G(n23), .D(idata[167]), .Q(\_zzLB[3][187] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][188] ( .G(n23), .D(idata[168]), .Q(\_zzLB[3][188] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][189] ( .G(n23), .D(idata[169]), .Q(\_zzLB[3][189] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][190] ( .G(n23), .D(idata[170]), .Q(\_zzLB[3][190] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][191] ( .G(n23), .D(idata[171]), .Q(\_zzLB[3][191] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][192] ( .G(n23), .D(idata[172]), .Q(\_zzLB[3][192] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][193] ( .G(n23), .D(idata[173]), .Q(\_zzLB[3][193] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][194] ( .G(n23), .D(idata[174]), .Q(\_zzLB[3][194] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][195] ( .G(n23), .D(idata[175]), .Q(\_zzLB[3][195] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][196] ( .G(n23), .D(idata[176]), .Q(\_zzLB[3][196] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][197] ( .G(n23), .D(idata[177]), .Q(\_zzLB[3][197] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][198] ( .G(n23), .D(idata[178]), .Q(\_zzLB[3][198] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][199] ( .G(n23), .D(idata[179]), .Q(\_zzLB[3][199] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][200] ( .G(n23), .D(idata[180]), .Q(\_zzLB[3][200] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][201] ( .G(n23), .D(idata[181]), .Q(\_zzLB[3][201] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][202] ( .G(n23), .D(idata[182]), .Q(\_zzLB[3][202] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][203] ( .G(n23), .D(idata[183]), .Q(\_zzLB[3][203] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][204] ( .G(n23), .D(idata[184]), .Q(\_zzLB[3][204] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][205] ( .G(n23), .D(idata[185]), .Q(\_zzLB[3][205] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][206] ( .G(n23), .D(idata[186]), .Q(\_zzLB[3][206] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][207] ( .G(n23), .D(idata[187]), .Q(\_zzLB[3][207] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][208] ( .G(n23), .D(idata[188]), .Q(\_zzLB[3][208] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][209] ( .G(n23), .D(idata[189]), .Q(\_zzLB[3][209] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][210] ( .G(n23), .D(idata[190]), .Q(\_zzLB[3][210] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][211] ( .G(n23), .D(idata[191]), .Q(\_zzLB[3][211] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][212] ( .G(n23), .D(idata[192]), .Q(\_zzLB[3][212] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][213] ( .G(n23), .D(idata[193]), .Q(\_zzLB[3][213] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][214] ( .G(n23), .D(idata[194]), .Q(\_zzLB[3][214] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][215] ( .G(n23), .D(idata[195]), .Q(\_zzLB[3][215] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][216] ( .G(n23), .D(idata[196]), .Q(\_zzLB[3][216] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][217] ( .G(n23), .D(idata[197]), .Q(\_zzLB[3][217] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][218] ( .G(n23), .D(idata[198]), .Q(\_zzLB[3][218] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][219] ( .G(n23), .D(idata[199]), .Q(\_zzLB[3][219] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][220] ( .G(n23), .D(idata[200]), .Q(\_zzLB[3][220] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][221] ( .G(n23), .D(idata[201]), .Q(\_zzLB[3][221] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][222] ( .G(n23), .D(idata[202]), .Q(\_zzLB[3][222] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][223] ( .G(n23), .D(idata[203]), .Q(\_zzLB[3][223] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][224] ( .G(n23), .D(idata[204]), .Q(\_zzLB[3][224] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][225] ( .G(n23), .D(idata[205]), .Q(\_zzLB[3][225] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][226] ( .G(n23), .D(idata[206]), .Q(\_zzLB[3][226] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][227] ( .G(n23), .D(idata[207]), .Q(\_zzLB[3][227] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][228] ( .G(n23), .D(idata[208]), .Q(\_zzLB[3][228] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][229] ( .G(n23), .D(idata[209]), .Q(\_zzLB[3][229] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][230] ( .G(n23), .D(idata[210]), .Q(\_zzLB[3][230] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][231] ( .G(n23), .D(idata[211]), .Q(\_zzLB[3][231] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][232] ( .G(n23), .D(idata[212]), .Q(\_zzLB[3][232] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][233] ( .G(n23), .D(idata[213]), .Q(\_zzLB[3][233] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][234] ( .G(n23), .D(idata[214]), .Q(\_zzLB[3][234] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][235] ( .G(n23), .D(idata[215]), .Q(\_zzLB[3][235] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][236] ( .G(n23), .D(idata[216]), .Q(\_zzLB[3][236] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][237] ( .G(n23), .D(idata[217]), .Q(\_zzLB[3][237] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][238] ( .G(n23), .D(idata[218]), .Q(\_zzLB[3][238] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][239] ( .G(n23), .D(idata[219]), .Q(\_zzLB[3][239] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][240] ( .G(n23), .D(idata[220]), .Q(\_zzLB[3][240] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][241] ( .G(n23), .D(idata[221]), .Q(\_zzLB[3][241] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][242] ( .G(n23), .D(idata[222]), .Q(\_zzLB[3][242] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][243] ( .G(n23), .D(idata[223]), .Q(\_zzLB[3][243] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][244] ( .G(n23), .D(idata[224]), .Q(\_zzLB[3][244] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][245] ( .G(n23), .D(idata[225]), .Q(\_zzLB[3][245] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][246] ( .G(n23), .D(idata[226]), .Q(\_zzLB[3][246] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][247] ( .G(n23), .D(idata[227]), .Q(\_zzLB[3][247] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][248] ( .G(n23), .D(idata[228]), .Q(\_zzLB[3][248] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][249] ( .G(n23), .D(idata[229]), .Q(\_zzLB[3][249] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][250] ( .G(n23), .D(idata[230]), .Q(\_zzLB[3][250] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][251] ( .G(n23), .D(idata[231]), .Q(\_zzLB[3][251] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][252] ( .G(n23), .D(idata[232]), .Q(\_zzLB[3][252] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][253] ( .G(n23), .D(idata[233]), .Q(\_zzLB[3][253] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][254] ( .G(n23), .D(idata[234]), .Q(\_zzLB[3][254] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][255] ( .G(n23), .D(idata[235]), .Q(\_zzLB[3][255] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][256] ( .G(n23), .D(idata[236]), .Q(\_zzLB[3][256] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][257] ( .G(n23), .D(idata[237]), .Q(\_zzLB[3][257] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][258] ( .G(n23), .D(idata[238]), .Q(\_zzLB[3][258] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][259] ( .G(n23), .D(idata[239]), .Q(\_zzLB[3][259] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][260] ( .G(n23), .D(idata[240]), .Q(\_zzLB[3][260] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][261] ( .G(n23), .D(idata[241]), .Q(\_zzLB[3][261] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][262] ( .G(n23), .D(idata[242]), .Q(\_zzLB[3][262] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][263] ( .G(n23), .D(idata[243]), .Q(\_zzLB[3][263] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][264] ( .G(n23), .D(idata[244]), .Q(\_zzLB[3][264] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][265] ( .G(n23), .D(idata[245]), .Q(\_zzLB[3][265] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][266] ( .G(n23), .D(idata[246]), .Q(\_zzLB[3][266] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][267] ( .G(n23), .D(idata[247]), .Q(\_zzLB[3][267] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][268] ( .G(n23), .D(idata[248]), .Q(\_zzLB[3][268] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][269] ( .G(n23), .D(idata[249]), .Q(\_zzLB[3][269] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][270] ( .G(n23), .D(idata[250]), .Q(\_zzLB[3][270] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][271] ( .G(n23), .D(idata[251]), .Q(\_zzLB[3][271] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][272] ( .G(n23), .D(idata[252]), .Q(\_zzLB[3][272] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][273] ( .G(n23), .D(idata[253]), .Q(\_zzLB[3][273] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][274] ( .G(n23), .D(idata[254]), .Q(\_zzLB[3][274] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][275] ( .G(n23), .D(idata[255]), .Q(\_zzLB[3][275] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][276] ( .G(n23), .D(idata[256]), .Q(\_zzLB[3][276] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][277] ( .G(n23), .D(idata[257]), .Q(\_zzLB[3][277] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][278] ( .G(n23), .D(idata[258]), .Q(\_zzLB[3][278] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][279] ( .G(n23), .D(idata[259]), .Q(\_zzLB[3][279] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][280] ( .G(n23), .D(idata[260]), .Q(\_zzLB[3][280] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][281] ( .G(n23), .D(idata[261]), .Q(\_zzLB[3][281] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][282] ( .G(n23), .D(idata[262]), .Q(\_zzLB[3][282] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][283] ( .G(n23), .D(idata[263]), .Q(\_zzLB[3][283] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][284] ( .G(n23), .D(idata[264]), .Q(\_zzLB[3][284] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][285] ( .G(n23), .D(idata[265]), .Q(\_zzLB[3][285] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][286] ( .G(n23), .D(idata[266]), .Q(\_zzLB[3][286] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][287] ( .G(n23), .D(idata[267]), .Q(\_zzLB[3][287] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][288] ( .G(n23), .D(idata[268]), .Q(\_zzLB[3][288] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][289] ( .G(n23), .D(idata[269]), .Q(\_zzLB[3][289] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][290] ( .G(n23), .D(idata[270]), .Q(\_zzLB[3][290] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][291] ( .G(n23), .D(idata[271]), .Q(\_zzLB[3][291] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][292] ( .G(n23), .D(idata[272]), .Q(\_zzLB[3][292] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][293] ( .G(n23), .D(idata[273]), .Q(\_zzLB[3][293] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][294] ( .G(n23), .D(idata[274]), .Q(\_zzLB[3][294] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][295] ( .G(n23), .D(idata[275]), .Q(\_zzLB[3][295] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][296] ( .G(n23), .D(idata[276]), .Q(\_zzLB[3][296] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][297] ( .G(n23), .D(idata[277]), .Q(\_zzLB[3][297] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][298] ( .G(n23), .D(idata[278]), .Q(\_zzLB[3][298] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][299] ( .G(n23), .D(idata[279]), .Q(\_zzLB[3][299] ), .QN( ));
Q_LDP0 \_zzLB_REG[3][300] ( .G(n23), .D(ireq), .Q(\_zzLB[3][300] ), .QN( ));
Q_MX04 U1878 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][0] ), .A1(\_zzLB[1][0] ), .A2(\_zzLB[2][0] ), .A3(\_zzLB[3][0] ), .Z(ocbid[0]));
Q_MX04 U1879 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][1] ), .A1(\_zzLB[1][1] ), .A2(\_zzLB[2][1] ), .A3(\_zzLB[3][1] ), .Z(ocbid[1]));
Q_MX04 U1880 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][2] ), .A1(\_zzLB[1][2] ), .A2(\_zzLB[2][2] ), .A3(\_zzLB[3][2] ), .Z(ocbid[2]));
Q_MX04 U1881 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][3] ), .A1(\_zzLB[1][3] ), .A2(\_zzLB[2][3] ), .A3(\_zzLB[3][3] ), .Z(ocbid[3]));
Q_MX04 U1882 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][4] ), .A1(\_zzLB[1][4] ), .A2(\_zzLB[2][4] ), .A3(\_zzLB[3][4] ), .Z(ocbid[4]));
Q_MX04 U1883 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][5] ), .A1(\_zzLB[1][5] ), .A2(\_zzLB[2][5] ), .A3(\_zzLB[3][5] ), .Z(ocbid[5]));
Q_MX04 U1884 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][6] ), .A1(\_zzLB[1][6] ), .A2(\_zzLB[2][6] ), .A3(\_zzLB[3][6] ), .Z(ocbid[6]));
Q_MX04 U1885 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][7] ), .A1(\_zzLB[1][7] ), .A2(\_zzLB[2][7] ), .A3(\_zzLB[3][7] ), .Z(ocbid[7]));
Q_MX04 U1886 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][8] ), .A1(\_zzLB[1][8] ), .A2(\_zzLB[2][8] ), .A3(\_zzLB[3][8] ), .Z(ocbid[8]));
Q_MX04 U1887 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][9] ), .A1(\_zzLB[1][9] ), .A2(\_zzLB[2][9] ), .A3(\_zzLB[3][9] ), .Z(ocbid[9]));
Q_MX04 U1888 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][10] ), .A1(\_zzLB[1][10] ), .A2(\_zzLB[2][10] ), .A3(\_zzLB[3][10] ), .Z(ocbid[10]));
Q_MX04 U1889 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][11] ), .A1(\_zzLB[1][11] ), .A2(\_zzLB[2][11] ), .A3(\_zzLB[3][11] ), .Z(ocbid[11]));
Q_MX04 U1890 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][12] ), .A1(\_zzLB[1][12] ), .A2(\_zzLB[2][12] ), .A3(\_zzLB[3][12] ), .Z(ocbid[12]));
Q_MX04 U1891 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][13] ), .A1(\_zzLB[1][13] ), .A2(\_zzLB[2][13] ), .A3(\_zzLB[3][13] ), .Z(ocbid[13]));
Q_MX04 U1892 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][14] ), .A1(\_zzLB[1][14] ), .A2(\_zzLB[2][14] ), .A3(\_zzLB[3][14] ), .Z(ocbid[14]));
Q_MX04 U1893 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][15] ), .A1(\_zzLB[1][15] ), .A2(\_zzLB[2][15] ), .A3(\_zzLB[3][15] ), .Z(ocbid[15]));
Q_MX04 U1894 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][16] ), .A1(\_zzLB[1][16] ), .A2(\_zzLB[2][16] ), .A3(\_zzLB[3][16] ), .Z(ocbid[16]));
Q_MX04 U1895 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][17] ), .A1(\_zzLB[1][17] ), .A2(\_zzLB[2][17] ), .A3(\_zzLB[3][17] ), .Z(ocbid[17]));
Q_MX04 U1896 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][18] ), .A1(\_zzLB[1][18] ), .A2(\_zzLB[2][18] ), .A3(\_zzLB[3][18] ), .Z(ocbid[18]));
Q_MX04 U1897 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][19] ), .A1(\_zzLB[1][19] ), .A2(\_zzLB[2][19] ), .A3(\_zzLB[3][19] ), .Z(ocbid[19]));
Q_MX04 U1898 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][20] ), .A1(\_zzLB[1][20] ), .A2(\_zzLB[2][20] ), .A3(\_zzLB[3][20] ), .Z(odata[0]));
Q_MX04 U1899 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][21] ), .A1(\_zzLB[1][21] ), .A2(\_zzLB[2][21] ), .A3(\_zzLB[3][21] ), .Z(odata[1]));
Q_MX04 U1900 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][22] ), .A1(\_zzLB[1][22] ), .A2(\_zzLB[2][22] ), .A3(\_zzLB[3][22] ), .Z(odata[2]));
Q_MX04 U1901 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][23] ), .A1(\_zzLB[1][23] ), .A2(\_zzLB[2][23] ), .A3(\_zzLB[3][23] ), .Z(odata[3]));
Q_MX04 U1902 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][24] ), .A1(\_zzLB[1][24] ), .A2(\_zzLB[2][24] ), .A3(\_zzLB[3][24] ), .Z(odata[4]));
Q_MX04 U1903 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][25] ), .A1(\_zzLB[1][25] ), .A2(\_zzLB[2][25] ), .A3(\_zzLB[3][25] ), .Z(odata[5]));
Q_MX04 U1904 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][26] ), .A1(\_zzLB[1][26] ), .A2(\_zzLB[2][26] ), .A3(\_zzLB[3][26] ), .Z(odata[6]));
Q_MX04 U1905 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][27] ), .A1(\_zzLB[1][27] ), .A2(\_zzLB[2][27] ), .A3(\_zzLB[3][27] ), .Z(odata[7]));
Q_MX04 U1906 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][28] ), .A1(\_zzLB[1][28] ), .A2(\_zzLB[2][28] ), .A3(\_zzLB[3][28] ), .Z(odata[8]));
Q_MX04 U1907 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][29] ), .A1(\_zzLB[1][29] ), .A2(\_zzLB[2][29] ), .A3(\_zzLB[3][29] ), .Z(odata[9]));
Q_MX04 U1908 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][30] ), .A1(\_zzLB[1][30] ), .A2(\_zzLB[2][30] ), .A3(\_zzLB[3][30] ), .Z(odata[10]));
Q_MX04 U1909 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][31] ), .A1(\_zzLB[1][31] ), .A2(\_zzLB[2][31] ), .A3(\_zzLB[3][31] ), .Z(odata[11]));
Q_MX04 U1910 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][32] ), .A1(\_zzLB[1][32] ), .A2(\_zzLB[2][32] ), .A3(\_zzLB[3][32] ), .Z(odata[12]));
Q_MX04 U1911 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][33] ), .A1(\_zzLB[1][33] ), .A2(\_zzLB[2][33] ), .A3(\_zzLB[3][33] ), .Z(odata[13]));
Q_MX04 U1912 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][34] ), .A1(\_zzLB[1][34] ), .A2(\_zzLB[2][34] ), .A3(\_zzLB[3][34] ), .Z(odata[14]));
Q_MX04 U1913 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][35] ), .A1(\_zzLB[1][35] ), .A2(\_zzLB[2][35] ), .A3(\_zzLB[3][35] ), .Z(odata[15]));
Q_MX04 U1914 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][36] ), .A1(\_zzLB[1][36] ), .A2(\_zzLB[2][36] ), .A3(\_zzLB[3][36] ), .Z(odata[16]));
Q_MX04 U1915 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][37] ), .A1(\_zzLB[1][37] ), .A2(\_zzLB[2][37] ), .A3(\_zzLB[3][37] ), .Z(odata[17]));
Q_MX04 U1916 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][38] ), .A1(\_zzLB[1][38] ), .A2(\_zzLB[2][38] ), .A3(\_zzLB[3][38] ), .Z(odata[18]));
Q_MX04 U1917 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][39] ), .A1(\_zzLB[1][39] ), .A2(\_zzLB[2][39] ), .A3(\_zzLB[3][39] ), .Z(odata[19]));
Q_MX04 U1918 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][40] ), .A1(\_zzLB[1][40] ), .A2(\_zzLB[2][40] ), .A3(\_zzLB[3][40] ), .Z(odata[20]));
Q_MX04 U1919 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][41] ), .A1(\_zzLB[1][41] ), .A2(\_zzLB[2][41] ), .A3(\_zzLB[3][41] ), .Z(odata[21]));
Q_MX04 U1920 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][42] ), .A1(\_zzLB[1][42] ), .A2(\_zzLB[2][42] ), .A3(\_zzLB[3][42] ), .Z(odata[22]));
Q_MX04 U1921 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][43] ), .A1(\_zzLB[1][43] ), .A2(\_zzLB[2][43] ), .A3(\_zzLB[3][43] ), .Z(odata[23]));
Q_MX04 U1922 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][44] ), .A1(\_zzLB[1][44] ), .A2(\_zzLB[2][44] ), .A3(\_zzLB[3][44] ), .Z(odata[24]));
Q_MX04 U1923 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][45] ), .A1(\_zzLB[1][45] ), .A2(\_zzLB[2][45] ), .A3(\_zzLB[3][45] ), .Z(odata[25]));
Q_MX04 U1924 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][46] ), .A1(\_zzLB[1][46] ), .A2(\_zzLB[2][46] ), .A3(\_zzLB[3][46] ), .Z(odata[26]));
Q_MX04 U1925 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][47] ), .A1(\_zzLB[1][47] ), .A2(\_zzLB[2][47] ), .A3(\_zzLB[3][47] ), .Z(odata[27]));
Q_MX04 U1926 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][48] ), .A1(\_zzLB[1][48] ), .A2(\_zzLB[2][48] ), .A3(\_zzLB[3][48] ), .Z(odata[28]));
Q_MX04 U1927 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][49] ), .A1(\_zzLB[1][49] ), .A2(\_zzLB[2][49] ), .A3(\_zzLB[3][49] ), .Z(odata[29]));
Q_MX04 U1928 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][50] ), .A1(\_zzLB[1][50] ), .A2(\_zzLB[2][50] ), .A3(\_zzLB[3][50] ), .Z(odata[30]));
Q_MX04 U1929 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][51] ), .A1(\_zzLB[1][51] ), .A2(\_zzLB[2][51] ), .A3(\_zzLB[3][51] ), .Z(odata[31]));
Q_MX04 U1930 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][52] ), .A1(\_zzLB[1][52] ), .A2(\_zzLB[2][52] ), .A3(\_zzLB[3][52] ), .Z(odata[32]));
Q_MX04 U1931 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][53] ), .A1(\_zzLB[1][53] ), .A2(\_zzLB[2][53] ), .A3(\_zzLB[3][53] ), .Z(odata[33]));
Q_MX04 U1932 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][54] ), .A1(\_zzLB[1][54] ), .A2(\_zzLB[2][54] ), .A3(\_zzLB[3][54] ), .Z(odata[34]));
Q_MX04 U1933 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][55] ), .A1(\_zzLB[1][55] ), .A2(\_zzLB[2][55] ), .A3(\_zzLB[3][55] ), .Z(odata[35]));
Q_MX04 U1934 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][56] ), .A1(\_zzLB[1][56] ), .A2(\_zzLB[2][56] ), .A3(\_zzLB[3][56] ), .Z(odata[36]));
Q_MX04 U1935 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][57] ), .A1(\_zzLB[1][57] ), .A2(\_zzLB[2][57] ), .A3(\_zzLB[3][57] ), .Z(odata[37]));
Q_MX04 U1936 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][58] ), .A1(\_zzLB[1][58] ), .A2(\_zzLB[2][58] ), .A3(\_zzLB[3][58] ), .Z(odata[38]));
Q_MX04 U1937 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][59] ), .A1(\_zzLB[1][59] ), .A2(\_zzLB[2][59] ), .A3(\_zzLB[3][59] ), .Z(odata[39]));
Q_MX04 U1938 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][60] ), .A1(\_zzLB[1][60] ), .A2(\_zzLB[2][60] ), .A3(\_zzLB[3][60] ), .Z(odata[40]));
Q_MX04 U1939 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][61] ), .A1(\_zzLB[1][61] ), .A2(\_zzLB[2][61] ), .A3(\_zzLB[3][61] ), .Z(odata[41]));
Q_MX04 U1940 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][62] ), .A1(\_zzLB[1][62] ), .A2(\_zzLB[2][62] ), .A3(\_zzLB[3][62] ), .Z(odata[42]));
Q_MX04 U1941 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][63] ), .A1(\_zzLB[1][63] ), .A2(\_zzLB[2][63] ), .A3(\_zzLB[3][63] ), .Z(odata[43]));
Q_MX04 U1942 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][64] ), .A1(\_zzLB[1][64] ), .A2(\_zzLB[2][64] ), .A3(\_zzLB[3][64] ), .Z(odata[44]));
Q_MX04 U1943 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][65] ), .A1(\_zzLB[1][65] ), .A2(\_zzLB[2][65] ), .A3(\_zzLB[3][65] ), .Z(odata[45]));
Q_MX04 U1944 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][66] ), .A1(\_zzLB[1][66] ), .A2(\_zzLB[2][66] ), .A3(\_zzLB[3][66] ), .Z(odata[46]));
Q_MX04 U1945 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][67] ), .A1(\_zzLB[1][67] ), .A2(\_zzLB[2][67] ), .A3(\_zzLB[3][67] ), .Z(odata[47]));
Q_MX04 U1946 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][68] ), .A1(\_zzLB[1][68] ), .A2(\_zzLB[2][68] ), .A3(\_zzLB[3][68] ), .Z(odata[48]));
Q_MX04 U1947 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][69] ), .A1(\_zzLB[1][69] ), .A2(\_zzLB[2][69] ), .A3(\_zzLB[3][69] ), .Z(odata[49]));
Q_MX04 U1948 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][70] ), .A1(\_zzLB[1][70] ), .A2(\_zzLB[2][70] ), .A3(\_zzLB[3][70] ), .Z(odata[50]));
Q_MX04 U1949 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][71] ), .A1(\_zzLB[1][71] ), .A2(\_zzLB[2][71] ), .A3(\_zzLB[3][71] ), .Z(odata[51]));
Q_MX04 U1950 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][72] ), .A1(\_zzLB[1][72] ), .A2(\_zzLB[2][72] ), .A3(\_zzLB[3][72] ), .Z(odata[52]));
Q_MX04 U1951 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][73] ), .A1(\_zzLB[1][73] ), .A2(\_zzLB[2][73] ), .A3(\_zzLB[3][73] ), .Z(odata[53]));
Q_MX04 U1952 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][74] ), .A1(\_zzLB[1][74] ), .A2(\_zzLB[2][74] ), .A3(\_zzLB[3][74] ), .Z(odata[54]));
Q_MX04 U1953 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][75] ), .A1(\_zzLB[1][75] ), .A2(\_zzLB[2][75] ), .A3(\_zzLB[3][75] ), .Z(odata[55]));
Q_MX04 U1954 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][76] ), .A1(\_zzLB[1][76] ), .A2(\_zzLB[2][76] ), .A3(\_zzLB[3][76] ), .Z(odata[56]));
Q_MX04 U1955 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][77] ), .A1(\_zzLB[1][77] ), .A2(\_zzLB[2][77] ), .A3(\_zzLB[3][77] ), .Z(odata[57]));
Q_MX04 U1956 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][78] ), .A1(\_zzLB[1][78] ), .A2(\_zzLB[2][78] ), .A3(\_zzLB[3][78] ), .Z(odata[58]));
Q_MX04 U1957 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][79] ), .A1(\_zzLB[1][79] ), .A2(\_zzLB[2][79] ), .A3(\_zzLB[3][79] ), .Z(odata[59]));
Q_MX04 U1958 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][80] ), .A1(\_zzLB[1][80] ), .A2(\_zzLB[2][80] ), .A3(\_zzLB[3][80] ), .Z(odata[60]));
Q_MX04 U1959 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][81] ), .A1(\_zzLB[1][81] ), .A2(\_zzLB[2][81] ), .A3(\_zzLB[3][81] ), .Z(odata[61]));
Q_MX04 U1960 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][82] ), .A1(\_zzLB[1][82] ), .A2(\_zzLB[2][82] ), .A3(\_zzLB[3][82] ), .Z(odata[62]));
Q_MX04 U1961 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][83] ), .A1(\_zzLB[1][83] ), .A2(\_zzLB[2][83] ), .A3(\_zzLB[3][83] ), .Z(odata[63]));
Q_MX04 U1962 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][84] ), .A1(\_zzLB[1][84] ), .A2(\_zzLB[2][84] ), .A3(\_zzLB[3][84] ), .Z(odata[64]));
Q_MX04 U1963 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][85] ), .A1(\_zzLB[1][85] ), .A2(\_zzLB[2][85] ), .A3(\_zzLB[3][85] ), .Z(odata[65]));
Q_MX04 U1964 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][86] ), .A1(\_zzLB[1][86] ), .A2(\_zzLB[2][86] ), .A3(\_zzLB[3][86] ), .Z(odata[66]));
Q_MX04 U1965 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][87] ), .A1(\_zzLB[1][87] ), .A2(\_zzLB[2][87] ), .A3(\_zzLB[3][87] ), .Z(odata[67]));
Q_MX04 U1966 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][88] ), .A1(\_zzLB[1][88] ), .A2(\_zzLB[2][88] ), .A3(\_zzLB[3][88] ), .Z(odata[68]));
Q_MX04 U1967 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][89] ), .A1(\_zzLB[1][89] ), .A2(\_zzLB[2][89] ), .A3(\_zzLB[3][89] ), .Z(odata[69]));
Q_MX04 U1968 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][90] ), .A1(\_zzLB[1][90] ), .A2(\_zzLB[2][90] ), .A3(\_zzLB[3][90] ), .Z(odata[70]));
Q_MX04 U1969 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][91] ), .A1(\_zzLB[1][91] ), .A2(\_zzLB[2][91] ), .A3(\_zzLB[3][91] ), .Z(odata[71]));
Q_MX04 U1970 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][92] ), .A1(\_zzLB[1][92] ), .A2(\_zzLB[2][92] ), .A3(\_zzLB[3][92] ), .Z(odata[72]));
Q_MX04 U1971 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][93] ), .A1(\_zzLB[1][93] ), .A2(\_zzLB[2][93] ), .A3(\_zzLB[3][93] ), .Z(odata[73]));
Q_MX04 U1972 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][94] ), .A1(\_zzLB[1][94] ), .A2(\_zzLB[2][94] ), .A3(\_zzLB[3][94] ), .Z(odata[74]));
Q_MX04 U1973 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][95] ), .A1(\_zzLB[1][95] ), .A2(\_zzLB[2][95] ), .A3(\_zzLB[3][95] ), .Z(odata[75]));
Q_MX04 U1974 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][96] ), .A1(\_zzLB[1][96] ), .A2(\_zzLB[2][96] ), .A3(\_zzLB[3][96] ), .Z(odata[76]));
Q_MX04 U1975 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][97] ), .A1(\_zzLB[1][97] ), .A2(\_zzLB[2][97] ), .A3(\_zzLB[3][97] ), .Z(odata[77]));
Q_MX04 U1976 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][98] ), .A1(\_zzLB[1][98] ), .A2(\_zzLB[2][98] ), .A3(\_zzLB[3][98] ), .Z(odata[78]));
Q_MX04 U1977 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][99] ), .A1(\_zzLB[1][99] ), .A2(\_zzLB[2][99] ), .A3(\_zzLB[3][99] ), .Z(odata[79]));
Q_MX04 U1978 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][100] ), .A1(\_zzLB[1][100] ), .A2(\_zzLB[2][100] ), .A3(\_zzLB[3][100] ), .Z(odata[80]));
Q_MX04 U1979 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][101] ), .A1(\_zzLB[1][101] ), .A2(\_zzLB[2][101] ), .A3(\_zzLB[3][101] ), .Z(odata[81]));
Q_MX04 U1980 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][102] ), .A1(\_zzLB[1][102] ), .A2(\_zzLB[2][102] ), .A3(\_zzLB[3][102] ), .Z(odata[82]));
Q_MX04 U1981 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][103] ), .A1(\_zzLB[1][103] ), .A2(\_zzLB[2][103] ), .A3(\_zzLB[3][103] ), .Z(odata[83]));
Q_MX04 U1982 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][104] ), .A1(\_zzLB[1][104] ), .A2(\_zzLB[2][104] ), .A3(\_zzLB[3][104] ), .Z(odata[84]));
Q_MX04 U1983 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][105] ), .A1(\_zzLB[1][105] ), .A2(\_zzLB[2][105] ), .A3(\_zzLB[3][105] ), .Z(odata[85]));
Q_MX04 U1984 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][106] ), .A1(\_zzLB[1][106] ), .A2(\_zzLB[2][106] ), .A3(\_zzLB[3][106] ), .Z(odata[86]));
Q_MX04 U1985 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][107] ), .A1(\_zzLB[1][107] ), .A2(\_zzLB[2][107] ), .A3(\_zzLB[3][107] ), .Z(odata[87]));
Q_MX04 U1986 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][108] ), .A1(\_zzLB[1][108] ), .A2(\_zzLB[2][108] ), .A3(\_zzLB[3][108] ), .Z(odata[88]));
Q_MX04 U1987 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][109] ), .A1(\_zzLB[1][109] ), .A2(\_zzLB[2][109] ), .A3(\_zzLB[3][109] ), .Z(odata[89]));
Q_MX04 U1988 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][110] ), .A1(\_zzLB[1][110] ), .A2(\_zzLB[2][110] ), .A3(\_zzLB[3][110] ), .Z(odata[90]));
Q_MX04 U1989 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][111] ), .A1(\_zzLB[1][111] ), .A2(\_zzLB[2][111] ), .A3(\_zzLB[3][111] ), .Z(odata[91]));
Q_MX04 U1990 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][112] ), .A1(\_zzLB[1][112] ), .A2(\_zzLB[2][112] ), .A3(\_zzLB[3][112] ), .Z(odata[92]));
Q_MX04 U1991 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][113] ), .A1(\_zzLB[1][113] ), .A2(\_zzLB[2][113] ), .A3(\_zzLB[3][113] ), .Z(odata[93]));
Q_MX04 U1992 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][114] ), .A1(\_zzLB[1][114] ), .A2(\_zzLB[2][114] ), .A3(\_zzLB[3][114] ), .Z(odata[94]));
Q_MX04 U1993 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][115] ), .A1(\_zzLB[1][115] ), .A2(\_zzLB[2][115] ), .A3(\_zzLB[3][115] ), .Z(odata[95]));
Q_MX04 U1994 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][116] ), .A1(\_zzLB[1][116] ), .A2(\_zzLB[2][116] ), .A3(\_zzLB[3][116] ), .Z(odata[96]));
Q_MX04 U1995 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][117] ), .A1(\_zzLB[1][117] ), .A2(\_zzLB[2][117] ), .A3(\_zzLB[3][117] ), .Z(odata[97]));
Q_MX04 U1996 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][118] ), .A1(\_zzLB[1][118] ), .A2(\_zzLB[2][118] ), .A3(\_zzLB[3][118] ), .Z(odata[98]));
Q_MX04 U1997 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][119] ), .A1(\_zzLB[1][119] ), .A2(\_zzLB[2][119] ), .A3(\_zzLB[3][119] ), .Z(odata[99]));
Q_MX04 U1998 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][120] ), .A1(\_zzLB[1][120] ), .A2(\_zzLB[2][120] ), .A3(\_zzLB[3][120] ), .Z(odata[100]));
Q_MX04 U1999 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][121] ), .A1(\_zzLB[1][121] ), .A2(\_zzLB[2][121] ), .A3(\_zzLB[3][121] ), .Z(odata[101]));
Q_MX04 U2000 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][122] ), .A1(\_zzLB[1][122] ), .A2(\_zzLB[2][122] ), .A3(\_zzLB[3][122] ), .Z(odata[102]));
Q_MX04 U2001 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][123] ), .A1(\_zzLB[1][123] ), .A2(\_zzLB[2][123] ), .A3(\_zzLB[3][123] ), .Z(odata[103]));
Q_MX04 U2002 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][124] ), .A1(\_zzLB[1][124] ), .A2(\_zzLB[2][124] ), .A3(\_zzLB[3][124] ), .Z(odata[104]));
Q_MX04 U2003 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][125] ), .A1(\_zzLB[1][125] ), .A2(\_zzLB[2][125] ), .A3(\_zzLB[3][125] ), .Z(odata[105]));
Q_MX04 U2004 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][126] ), .A1(\_zzLB[1][126] ), .A2(\_zzLB[2][126] ), .A3(\_zzLB[3][126] ), .Z(odata[106]));
Q_MX04 U2005 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][127] ), .A1(\_zzLB[1][127] ), .A2(\_zzLB[2][127] ), .A3(\_zzLB[3][127] ), .Z(odata[107]));
Q_MX04 U2006 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][128] ), .A1(\_zzLB[1][128] ), .A2(\_zzLB[2][128] ), .A3(\_zzLB[3][128] ), .Z(odata[108]));
Q_MX04 U2007 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][129] ), .A1(\_zzLB[1][129] ), .A2(\_zzLB[2][129] ), .A3(\_zzLB[3][129] ), .Z(odata[109]));
Q_MX04 U2008 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][130] ), .A1(\_zzLB[1][130] ), .A2(\_zzLB[2][130] ), .A3(\_zzLB[3][130] ), .Z(odata[110]));
Q_MX04 U2009 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][131] ), .A1(\_zzLB[1][131] ), .A2(\_zzLB[2][131] ), .A3(\_zzLB[3][131] ), .Z(odata[111]));
Q_MX04 U2010 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][132] ), .A1(\_zzLB[1][132] ), .A2(\_zzLB[2][132] ), .A3(\_zzLB[3][132] ), .Z(odata[112]));
Q_MX04 U2011 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][133] ), .A1(\_zzLB[1][133] ), .A2(\_zzLB[2][133] ), .A3(\_zzLB[3][133] ), .Z(odata[113]));
Q_MX04 U2012 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][134] ), .A1(\_zzLB[1][134] ), .A2(\_zzLB[2][134] ), .A3(\_zzLB[3][134] ), .Z(odata[114]));
Q_MX04 U2013 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][135] ), .A1(\_zzLB[1][135] ), .A2(\_zzLB[2][135] ), .A3(\_zzLB[3][135] ), .Z(odata[115]));
Q_MX04 U2014 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][136] ), .A1(\_zzLB[1][136] ), .A2(\_zzLB[2][136] ), .A3(\_zzLB[3][136] ), .Z(odata[116]));
Q_MX04 U2015 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][137] ), .A1(\_zzLB[1][137] ), .A2(\_zzLB[2][137] ), .A3(\_zzLB[3][137] ), .Z(odata[117]));
Q_MX04 U2016 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][138] ), .A1(\_zzLB[1][138] ), .A2(\_zzLB[2][138] ), .A3(\_zzLB[3][138] ), .Z(odata[118]));
Q_MX04 U2017 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][139] ), .A1(\_zzLB[1][139] ), .A2(\_zzLB[2][139] ), .A3(\_zzLB[3][139] ), .Z(odata[119]));
Q_MX04 U2018 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][140] ), .A1(\_zzLB[1][140] ), .A2(\_zzLB[2][140] ), .A3(\_zzLB[3][140] ), .Z(odata[120]));
Q_MX04 U2019 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][141] ), .A1(\_zzLB[1][141] ), .A2(\_zzLB[2][141] ), .A3(\_zzLB[3][141] ), .Z(odata[121]));
Q_MX04 U2020 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][142] ), .A1(\_zzLB[1][142] ), .A2(\_zzLB[2][142] ), .A3(\_zzLB[3][142] ), .Z(odata[122]));
Q_MX04 U2021 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][143] ), .A1(\_zzLB[1][143] ), .A2(\_zzLB[2][143] ), .A3(\_zzLB[3][143] ), .Z(odata[123]));
Q_MX04 U2022 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][144] ), .A1(\_zzLB[1][144] ), .A2(\_zzLB[2][144] ), .A3(\_zzLB[3][144] ), .Z(odata[124]));
Q_MX04 U2023 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][145] ), .A1(\_zzLB[1][145] ), .A2(\_zzLB[2][145] ), .A3(\_zzLB[3][145] ), .Z(odata[125]));
Q_MX04 U2024 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][146] ), .A1(\_zzLB[1][146] ), .A2(\_zzLB[2][146] ), .A3(\_zzLB[3][146] ), .Z(odata[126]));
Q_MX04 U2025 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][147] ), .A1(\_zzLB[1][147] ), .A2(\_zzLB[2][147] ), .A3(\_zzLB[3][147] ), .Z(odata[127]));
Q_MX04 U2026 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][148] ), .A1(\_zzLB[1][148] ), .A2(\_zzLB[2][148] ), .A3(\_zzLB[3][148] ), .Z(odata[128]));
Q_MX04 U2027 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][149] ), .A1(\_zzLB[1][149] ), .A2(\_zzLB[2][149] ), .A3(\_zzLB[3][149] ), .Z(odata[129]));
Q_MX04 U2028 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][150] ), .A1(\_zzLB[1][150] ), .A2(\_zzLB[2][150] ), .A3(\_zzLB[3][150] ), .Z(odata[130]));
Q_MX04 U2029 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][151] ), .A1(\_zzLB[1][151] ), .A2(\_zzLB[2][151] ), .A3(\_zzLB[3][151] ), .Z(odata[131]));
Q_MX04 U2030 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][152] ), .A1(\_zzLB[1][152] ), .A2(\_zzLB[2][152] ), .A3(\_zzLB[3][152] ), .Z(odata[132]));
Q_MX04 U2031 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][153] ), .A1(\_zzLB[1][153] ), .A2(\_zzLB[2][153] ), .A3(\_zzLB[3][153] ), .Z(odata[133]));
Q_MX04 U2032 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][154] ), .A1(\_zzLB[1][154] ), .A2(\_zzLB[2][154] ), .A3(\_zzLB[3][154] ), .Z(odata[134]));
Q_MX04 U2033 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][155] ), .A1(\_zzLB[1][155] ), .A2(\_zzLB[2][155] ), .A3(\_zzLB[3][155] ), .Z(odata[135]));
Q_MX04 U2034 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][156] ), .A1(\_zzLB[1][156] ), .A2(\_zzLB[2][156] ), .A3(\_zzLB[3][156] ), .Z(odata[136]));
Q_MX04 U2035 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][157] ), .A1(\_zzLB[1][157] ), .A2(\_zzLB[2][157] ), .A3(\_zzLB[3][157] ), .Z(odata[137]));
Q_MX04 U2036 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][158] ), .A1(\_zzLB[1][158] ), .A2(\_zzLB[2][158] ), .A3(\_zzLB[3][158] ), .Z(odata[138]));
Q_MX04 U2037 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][159] ), .A1(\_zzLB[1][159] ), .A2(\_zzLB[2][159] ), .A3(\_zzLB[3][159] ), .Z(odata[139]));
Q_MX04 U2038 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][160] ), .A1(\_zzLB[1][160] ), .A2(\_zzLB[2][160] ), .A3(\_zzLB[3][160] ), .Z(odata[140]));
Q_MX04 U2039 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][161] ), .A1(\_zzLB[1][161] ), .A2(\_zzLB[2][161] ), .A3(\_zzLB[3][161] ), .Z(odata[141]));
Q_MX04 U2040 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][162] ), .A1(\_zzLB[1][162] ), .A2(\_zzLB[2][162] ), .A3(\_zzLB[3][162] ), .Z(odata[142]));
Q_MX04 U2041 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][163] ), .A1(\_zzLB[1][163] ), .A2(\_zzLB[2][163] ), .A3(\_zzLB[3][163] ), .Z(odata[143]));
Q_MX04 U2042 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][164] ), .A1(\_zzLB[1][164] ), .A2(\_zzLB[2][164] ), .A3(\_zzLB[3][164] ), .Z(odata[144]));
Q_MX04 U2043 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][165] ), .A1(\_zzLB[1][165] ), .A2(\_zzLB[2][165] ), .A3(\_zzLB[3][165] ), .Z(odata[145]));
Q_MX04 U2044 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][166] ), .A1(\_zzLB[1][166] ), .A2(\_zzLB[2][166] ), .A3(\_zzLB[3][166] ), .Z(odata[146]));
Q_MX04 U2045 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][167] ), .A1(\_zzLB[1][167] ), .A2(\_zzLB[2][167] ), .A3(\_zzLB[3][167] ), .Z(odata[147]));
Q_MX04 U2046 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][168] ), .A1(\_zzLB[1][168] ), .A2(\_zzLB[2][168] ), .A3(\_zzLB[3][168] ), .Z(odata[148]));
Q_MX04 U2047 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][169] ), .A1(\_zzLB[1][169] ), .A2(\_zzLB[2][169] ), .A3(\_zzLB[3][169] ), .Z(odata[149]));
Q_MX04 U2048 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][170] ), .A1(\_zzLB[1][170] ), .A2(\_zzLB[2][170] ), .A3(\_zzLB[3][170] ), .Z(odata[150]));
Q_MX04 U2049 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][171] ), .A1(\_zzLB[1][171] ), .A2(\_zzLB[2][171] ), .A3(\_zzLB[3][171] ), .Z(odata[151]));
Q_MX04 U2050 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][172] ), .A1(\_zzLB[1][172] ), .A2(\_zzLB[2][172] ), .A3(\_zzLB[3][172] ), .Z(odata[152]));
Q_MX04 U2051 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][173] ), .A1(\_zzLB[1][173] ), .A2(\_zzLB[2][173] ), .A3(\_zzLB[3][173] ), .Z(odata[153]));
Q_MX04 U2052 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][174] ), .A1(\_zzLB[1][174] ), .A2(\_zzLB[2][174] ), .A3(\_zzLB[3][174] ), .Z(odata[154]));
Q_MX04 U2053 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][175] ), .A1(\_zzLB[1][175] ), .A2(\_zzLB[2][175] ), .A3(\_zzLB[3][175] ), .Z(odata[155]));
Q_MX04 U2054 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][176] ), .A1(\_zzLB[1][176] ), .A2(\_zzLB[2][176] ), .A3(\_zzLB[3][176] ), .Z(odata[156]));
Q_MX04 U2055 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][177] ), .A1(\_zzLB[1][177] ), .A2(\_zzLB[2][177] ), .A3(\_zzLB[3][177] ), .Z(odata[157]));
Q_MX04 U2056 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][178] ), .A1(\_zzLB[1][178] ), .A2(\_zzLB[2][178] ), .A3(\_zzLB[3][178] ), .Z(odata[158]));
Q_MX04 U2057 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][179] ), .A1(\_zzLB[1][179] ), .A2(\_zzLB[2][179] ), .A3(\_zzLB[3][179] ), .Z(odata[159]));
Q_MX04 U2058 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][180] ), .A1(\_zzLB[1][180] ), .A2(\_zzLB[2][180] ), .A3(\_zzLB[3][180] ), .Z(odata[160]));
Q_MX04 U2059 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][181] ), .A1(\_zzLB[1][181] ), .A2(\_zzLB[2][181] ), .A3(\_zzLB[3][181] ), .Z(odata[161]));
Q_MX04 U2060 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][182] ), .A1(\_zzLB[1][182] ), .A2(\_zzLB[2][182] ), .A3(\_zzLB[3][182] ), .Z(odata[162]));
Q_MX04 U2061 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][183] ), .A1(\_zzLB[1][183] ), .A2(\_zzLB[2][183] ), .A3(\_zzLB[3][183] ), .Z(odata[163]));
Q_MX04 U2062 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][184] ), .A1(\_zzLB[1][184] ), .A2(\_zzLB[2][184] ), .A3(\_zzLB[3][184] ), .Z(odata[164]));
Q_MX04 U2063 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][185] ), .A1(\_zzLB[1][185] ), .A2(\_zzLB[2][185] ), .A3(\_zzLB[3][185] ), .Z(odata[165]));
Q_MX04 U2064 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][186] ), .A1(\_zzLB[1][186] ), .A2(\_zzLB[2][186] ), .A3(\_zzLB[3][186] ), .Z(odata[166]));
Q_MX04 U2065 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][187] ), .A1(\_zzLB[1][187] ), .A2(\_zzLB[2][187] ), .A3(\_zzLB[3][187] ), .Z(odata[167]));
Q_MX04 U2066 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][188] ), .A1(\_zzLB[1][188] ), .A2(\_zzLB[2][188] ), .A3(\_zzLB[3][188] ), .Z(odata[168]));
Q_MX04 U2067 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][189] ), .A1(\_zzLB[1][189] ), .A2(\_zzLB[2][189] ), .A3(\_zzLB[3][189] ), .Z(odata[169]));
Q_MX04 U2068 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][190] ), .A1(\_zzLB[1][190] ), .A2(\_zzLB[2][190] ), .A3(\_zzLB[3][190] ), .Z(odata[170]));
Q_MX04 U2069 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][191] ), .A1(\_zzLB[1][191] ), .A2(\_zzLB[2][191] ), .A3(\_zzLB[3][191] ), .Z(odata[171]));
Q_MX04 U2070 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][192] ), .A1(\_zzLB[1][192] ), .A2(\_zzLB[2][192] ), .A3(\_zzLB[3][192] ), .Z(odata[172]));
Q_MX04 U2071 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][193] ), .A1(\_zzLB[1][193] ), .A2(\_zzLB[2][193] ), .A3(\_zzLB[3][193] ), .Z(odata[173]));
Q_MX04 U2072 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][194] ), .A1(\_zzLB[1][194] ), .A2(\_zzLB[2][194] ), .A3(\_zzLB[3][194] ), .Z(odata[174]));
Q_MX04 U2073 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][195] ), .A1(\_zzLB[1][195] ), .A2(\_zzLB[2][195] ), .A3(\_zzLB[3][195] ), .Z(odata[175]));
Q_MX04 U2074 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][196] ), .A1(\_zzLB[1][196] ), .A2(\_zzLB[2][196] ), .A3(\_zzLB[3][196] ), .Z(odata[176]));
Q_MX04 U2075 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][197] ), .A1(\_zzLB[1][197] ), .A2(\_zzLB[2][197] ), .A3(\_zzLB[3][197] ), .Z(odata[177]));
Q_MX04 U2076 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][198] ), .A1(\_zzLB[1][198] ), .A2(\_zzLB[2][198] ), .A3(\_zzLB[3][198] ), .Z(odata[178]));
Q_MX04 U2077 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][199] ), .A1(\_zzLB[1][199] ), .A2(\_zzLB[2][199] ), .A3(\_zzLB[3][199] ), .Z(odata[179]));
Q_MX04 U2078 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][200] ), .A1(\_zzLB[1][200] ), .A2(\_zzLB[2][200] ), .A3(\_zzLB[3][200] ), .Z(odata[180]));
Q_MX04 U2079 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][201] ), .A1(\_zzLB[1][201] ), .A2(\_zzLB[2][201] ), .A3(\_zzLB[3][201] ), .Z(odata[181]));
Q_MX04 U2080 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][202] ), .A1(\_zzLB[1][202] ), .A2(\_zzLB[2][202] ), .A3(\_zzLB[3][202] ), .Z(odata[182]));
Q_MX04 U2081 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][203] ), .A1(\_zzLB[1][203] ), .A2(\_zzLB[2][203] ), .A3(\_zzLB[3][203] ), .Z(odata[183]));
Q_MX04 U2082 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][204] ), .A1(\_zzLB[1][204] ), .A2(\_zzLB[2][204] ), .A3(\_zzLB[3][204] ), .Z(odata[184]));
Q_MX04 U2083 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][205] ), .A1(\_zzLB[1][205] ), .A2(\_zzLB[2][205] ), .A3(\_zzLB[3][205] ), .Z(odata[185]));
Q_MX04 U2084 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][206] ), .A1(\_zzLB[1][206] ), .A2(\_zzLB[2][206] ), .A3(\_zzLB[3][206] ), .Z(odata[186]));
Q_MX04 U2085 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][207] ), .A1(\_zzLB[1][207] ), .A2(\_zzLB[2][207] ), .A3(\_zzLB[3][207] ), .Z(odata[187]));
Q_MX04 U2086 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][208] ), .A1(\_zzLB[1][208] ), .A2(\_zzLB[2][208] ), .A3(\_zzLB[3][208] ), .Z(odata[188]));
Q_MX04 U2087 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][209] ), .A1(\_zzLB[1][209] ), .A2(\_zzLB[2][209] ), .A3(\_zzLB[3][209] ), .Z(odata[189]));
Q_MX04 U2088 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][210] ), .A1(\_zzLB[1][210] ), .A2(\_zzLB[2][210] ), .A3(\_zzLB[3][210] ), .Z(odata[190]));
Q_MX04 U2089 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][211] ), .A1(\_zzLB[1][211] ), .A2(\_zzLB[2][211] ), .A3(\_zzLB[3][211] ), .Z(odata[191]));
Q_MX04 U2090 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][212] ), .A1(\_zzLB[1][212] ), .A2(\_zzLB[2][212] ), .A3(\_zzLB[3][212] ), .Z(odata[192]));
Q_MX04 U2091 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][213] ), .A1(\_zzLB[1][213] ), .A2(\_zzLB[2][213] ), .A3(\_zzLB[3][213] ), .Z(odata[193]));
Q_MX04 U2092 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][214] ), .A1(\_zzLB[1][214] ), .A2(\_zzLB[2][214] ), .A3(\_zzLB[3][214] ), .Z(odata[194]));
Q_MX04 U2093 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][215] ), .A1(\_zzLB[1][215] ), .A2(\_zzLB[2][215] ), .A3(\_zzLB[3][215] ), .Z(odata[195]));
Q_MX04 U2094 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][216] ), .A1(\_zzLB[1][216] ), .A2(\_zzLB[2][216] ), .A3(\_zzLB[3][216] ), .Z(odata[196]));
Q_MX04 U2095 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][217] ), .A1(\_zzLB[1][217] ), .A2(\_zzLB[2][217] ), .A3(\_zzLB[3][217] ), .Z(odata[197]));
Q_MX04 U2096 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][218] ), .A1(\_zzLB[1][218] ), .A2(\_zzLB[2][218] ), .A3(\_zzLB[3][218] ), .Z(odata[198]));
Q_MX04 U2097 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][219] ), .A1(\_zzLB[1][219] ), .A2(\_zzLB[2][219] ), .A3(\_zzLB[3][219] ), .Z(odata[199]));
Q_MX04 U2098 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][220] ), .A1(\_zzLB[1][220] ), .A2(\_zzLB[2][220] ), .A3(\_zzLB[3][220] ), .Z(odata[200]));
Q_MX04 U2099 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][221] ), .A1(\_zzLB[1][221] ), .A2(\_zzLB[2][221] ), .A3(\_zzLB[3][221] ), .Z(odata[201]));
Q_MX04 U2100 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][222] ), .A1(\_zzLB[1][222] ), .A2(\_zzLB[2][222] ), .A3(\_zzLB[3][222] ), .Z(odata[202]));
Q_MX04 U2101 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][223] ), .A1(\_zzLB[1][223] ), .A2(\_zzLB[2][223] ), .A3(\_zzLB[3][223] ), .Z(odata[203]));
Q_MX04 U2102 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][224] ), .A1(\_zzLB[1][224] ), .A2(\_zzLB[2][224] ), .A3(\_zzLB[3][224] ), .Z(odata[204]));
Q_MX04 U2103 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][225] ), .A1(\_zzLB[1][225] ), .A2(\_zzLB[2][225] ), .A3(\_zzLB[3][225] ), .Z(odata[205]));
Q_MX04 U2104 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][226] ), .A1(\_zzLB[1][226] ), .A2(\_zzLB[2][226] ), .A3(\_zzLB[3][226] ), .Z(odata[206]));
Q_MX04 U2105 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][227] ), .A1(\_zzLB[1][227] ), .A2(\_zzLB[2][227] ), .A3(\_zzLB[3][227] ), .Z(odata[207]));
Q_MX04 U2106 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][228] ), .A1(\_zzLB[1][228] ), .A2(\_zzLB[2][228] ), .A3(\_zzLB[3][228] ), .Z(odata[208]));
Q_MX04 U2107 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][229] ), .A1(\_zzLB[1][229] ), .A2(\_zzLB[2][229] ), .A3(\_zzLB[3][229] ), .Z(odata[209]));
Q_MX04 U2108 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][230] ), .A1(\_zzLB[1][230] ), .A2(\_zzLB[2][230] ), .A3(\_zzLB[3][230] ), .Z(odata[210]));
Q_MX04 U2109 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][231] ), .A1(\_zzLB[1][231] ), .A2(\_zzLB[2][231] ), .A3(\_zzLB[3][231] ), .Z(odata[211]));
Q_MX04 U2110 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][232] ), .A1(\_zzLB[1][232] ), .A2(\_zzLB[2][232] ), .A3(\_zzLB[3][232] ), .Z(odata[212]));
Q_MX04 U2111 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][233] ), .A1(\_zzLB[1][233] ), .A2(\_zzLB[2][233] ), .A3(\_zzLB[3][233] ), .Z(odata[213]));
Q_MX04 U2112 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][234] ), .A1(\_zzLB[1][234] ), .A2(\_zzLB[2][234] ), .A3(\_zzLB[3][234] ), .Z(odata[214]));
Q_MX04 U2113 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][235] ), .A1(\_zzLB[1][235] ), .A2(\_zzLB[2][235] ), .A3(\_zzLB[3][235] ), .Z(odata[215]));
Q_MX04 U2114 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][236] ), .A1(\_zzLB[1][236] ), .A2(\_zzLB[2][236] ), .A3(\_zzLB[3][236] ), .Z(odata[216]));
Q_MX04 U2115 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][237] ), .A1(\_zzLB[1][237] ), .A2(\_zzLB[2][237] ), .A3(\_zzLB[3][237] ), .Z(odata[217]));
Q_MX04 U2116 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][238] ), .A1(\_zzLB[1][238] ), .A2(\_zzLB[2][238] ), .A3(\_zzLB[3][238] ), .Z(odata[218]));
Q_MX04 U2117 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][239] ), .A1(\_zzLB[1][239] ), .A2(\_zzLB[2][239] ), .A3(\_zzLB[3][239] ), .Z(odata[219]));
Q_MX04 U2118 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][240] ), .A1(\_zzLB[1][240] ), .A2(\_zzLB[2][240] ), .A3(\_zzLB[3][240] ), .Z(odata[220]));
Q_MX04 U2119 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][241] ), .A1(\_zzLB[1][241] ), .A2(\_zzLB[2][241] ), .A3(\_zzLB[3][241] ), .Z(odata[221]));
Q_MX04 U2120 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][242] ), .A1(\_zzLB[1][242] ), .A2(\_zzLB[2][242] ), .A3(\_zzLB[3][242] ), .Z(odata[222]));
Q_MX04 U2121 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][243] ), .A1(\_zzLB[1][243] ), .A2(\_zzLB[2][243] ), .A3(\_zzLB[3][243] ), .Z(odata[223]));
Q_MX04 U2122 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][244] ), .A1(\_zzLB[1][244] ), .A2(\_zzLB[2][244] ), .A3(\_zzLB[3][244] ), .Z(odata[224]));
Q_MX04 U2123 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][245] ), .A1(\_zzLB[1][245] ), .A2(\_zzLB[2][245] ), .A3(\_zzLB[3][245] ), .Z(odata[225]));
Q_MX04 U2124 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][246] ), .A1(\_zzLB[1][246] ), .A2(\_zzLB[2][246] ), .A3(\_zzLB[3][246] ), .Z(odata[226]));
Q_MX04 U2125 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][247] ), .A1(\_zzLB[1][247] ), .A2(\_zzLB[2][247] ), .A3(\_zzLB[3][247] ), .Z(odata[227]));
Q_MX04 U2126 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][248] ), .A1(\_zzLB[1][248] ), .A2(\_zzLB[2][248] ), .A3(\_zzLB[3][248] ), .Z(odata[228]));
Q_MX04 U2127 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][249] ), .A1(\_zzLB[1][249] ), .A2(\_zzLB[2][249] ), .A3(\_zzLB[3][249] ), .Z(odata[229]));
Q_MX04 U2128 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][250] ), .A1(\_zzLB[1][250] ), .A2(\_zzLB[2][250] ), .A3(\_zzLB[3][250] ), .Z(odata[230]));
Q_MX04 U2129 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][251] ), .A1(\_zzLB[1][251] ), .A2(\_zzLB[2][251] ), .A3(\_zzLB[3][251] ), .Z(odata[231]));
Q_MX04 U2130 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][252] ), .A1(\_zzLB[1][252] ), .A2(\_zzLB[2][252] ), .A3(\_zzLB[3][252] ), .Z(odata[232]));
Q_MX04 U2131 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][253] ), .A1(\_zzLB[1][253] ), .A2(\_zzLB[2][253] ), .A3(\_zzLB[3][253] ), .Z(odata[233]));
Q_MX04 U2132 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][254] ), .A1(\_zzLB[1][254] ), .A2(\_zzLB[2][254] ), .A3(\_zzLB[3][254] ), .Z(odata[234]));
Q_MX04 U2133 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][255] ), .A1(\_zzLB[1][255] ), .A2(\_zzLB[2][255] ), .A3(\_zzLB[3][255] ), .Z(odata[235]));
Q_MX04 U2134 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][256] ), .A1(\_zzLB[1][256] ), .A2(\_zzLB[2][256] ), .A3(\_zzLB[3][256] ), .Z(odata[236]));
Q_MX04 U2135 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][257] ), .A1(\_zzLB[1][257] ), .A2(\_zzLB[2][257] ), .A3(\_zzLB[3][257] ), .Z(odata[237]));
Q_MX04 U2136 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][258] ), .A1(\_zzLB[1][258] ), .A2(\_zzLB[2][258] ), .A3(\_zzLB[3][258] ), .Z(odata[238]));
Q_MX04 U2137 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][259] ), .A1(\_zzLB[1][259] ), .A2(\_zzLB[2][259] ), .A3(\_zzLB[3][259] ), .Z(odata[239]));
Q_MX04 U2138 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][260] ), .A1(\_zzLB[1][260] ), .A2(\_zzLB[2][260] ), .A3(\_zzLB[3][260] ), .Z(odata[240]));
Q_MX04 U2139 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][261] ), .A1(\_zzLB[1][261] ), .A2(\_zzLB[2][261] ), .A3(\_zzLB[3][261] ), .Z(odata[241]));
Q_MX04 U2140 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][262] ), .A1(\_zzLB[1][262] ), .A2(\_zzLB[2][262] ), .A3(\_zzLB[3][262] ), .Z(odata[242]));
Q_MX04 U2141 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][263] ), .A1(\_zzLB[1][263] ), .A2(\_zzLB[2][263] ), .A3(\_zzLB[3][263] ), .Z(odata[243]));
Q_MX04 U2142 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][264] ), .A1(\_zzLB[1][264] ), .A2(\_zzLB[2][264] ), .A3(\_zzLB[3][264] ), .Z(odata[244]));
Q_MX04 U2143 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][265] ), .A1(\_zzLB[1][265] ), .A2(\_zzLB[2][265] ), .A3(\_zzLB[3][265] ), .Z(odata[245]));
Q_MX04 U2144 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][266] ), .A1(\_zzLB[1][266] ), .A2(\_zzLB[2][266] ), .A3(\_zzLB[3][266] ), .Z(odata[246]));
Q_MX04 U2145 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][267] ), .A1(\_zzLB[1][267] ), .A2(\_zzLB[2][267] ), .A3(\_zzLB[3][267] ), .Z(odata[247]));
Q_MX04 U2146 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][268] ), .A1(\_zzLB[1][268] ), .A2(\_zzLB[2][268] ), .A3(\_zzLB[3][268] ), .Z(odata[248]));
Q_MX04 U2147 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][269] ), .A1(\_zzLB[1][269] ), .A2(\_zzLB[2][269] ), .A3(\_zzLB[3][269] ), .Z(odata[249]));
Q_MX04 U2148 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][270] ), .A1(\_zzLB[1][270] ), .A2(\_zzLB[2][270] ), .A3(\_zzLB[3][270] ), .Z(odata[250]));
Q_MX04 U2149 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][271] ), .A1(\_zzLB[1][271] ), .A2(\_zzLB[2][271] ), .A3(\_zzLB[3][271] ), .Z(odata[251]));
Q_MX04 U2150 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][272] ), .A1(\_zzLB[1][272] ), .A2(\_zzLB[2][272] ), .A3(\_zzLB[3][272] ), .Z(odata[252]));
Q_MX04 U2151 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][273] ), .A1(\_zzLB[1][273] ), .A2(\_zzLB[2][273] ), .A3(\_zzLB[3][273] ), .Z(odata[253]));
Q_MX04 U2152 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][274] ), .A1(\_zzLB[1][274] ), .A2(\_zzLB[2][274] ), .A3(\_zzLB[3][274] ), .Z(odata[254]));
Q_MX04 U2153 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][275] ), .A1(\_zzLB[1][275] ), .A2(\_zzLB[2][275] ), .A3(\_zzLB[3][275] ), .Z(odata[255]));
Q_MX04 U2154 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][276] ), .A1(\_zzLB[1][276] ), .A2(\_zzLB[2][276] ), .A3(\_zzLB[3][276] ), .Z(odata[256]));
Q_MX04 U2155 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][277] ), .A1(\_zzLB[1][277] ), .A2(\_zzLB[2][277] ), .A3(\_zzLB[3][277] ), .Z(odata[257]));
Q_MX04 U2156 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][278] ), .A1(\_zzLB[1][278] ), .A2(\_zzLB[2][278] ), .A3(\_zzLB[3][278] ), .Z(odata[258]));
Q_MX04 U2157 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][279] ), .A1(\_zzLB[1][279] ), .A2(\_zzLB[2][279] ), .A3(\_zzLB[3][279] ), .Z(odata[259]));
Q_MX04 U2158 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][280] ), .A1(\_zzLB[1][280] ), .A2(\_zzLB[2][280] ), .A3(\_zzLB[3][280] ), .Z(odata[260]));
Q_MX04 U2159 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][281] ), .A1(\_zzLB[1][281] ), .A2(\_zzLB[2][281] ), .A3(\_zzLB[3][281] ), .Z(odata[261]));
Q_MX04 U2160 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][282] ), .A1(\_zzLB[1][282] ), .A2(\_zzLB[2][282] ), .A3(\_zzLB[3][282] ), .Z(odata[262]));
Q_MX04 U2161 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][283] ), .A1(\_zzLB[1][283] ), .A2(\_zzLB[2][283] ), .A3(\_zzLB[3][283] ), .Z(odata[263]));
Q_MX04 U2162 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][284] ), .A1(\_zzLB[1][284] ), .A2(\_zzLB[2][284] ), .A3(\_zzLB[3][284] ), .Z(odata[264]));
Q_MX04 U2163 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][285] ), .A1(\_zzLB[1][285] ), .A2(\_zzLB[2][285] ), .A3(\_zzLB[3][285] ), .Z(odata[265]));
Q_MX04 U2164 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][286] ), .A1(\_zzLB[1][286] ), .A2(\_zzLB[2][286] ), .A3(\_zzLB[3][286] ), .Z(odata[266]));
Q_MX04 U2165 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][287] ), .A1(\_zzLB[1][287] ), .A2(\_zzLB[2][287] ), .A3(\_zzLB[3][287] ), .Z(odata[267]));
Q_MX04 U2166 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][288] ), .A1(\_zzLB[1][288] ), .A2(\_zzLB[2][288] ), .A3(\_zzLB[3][288] ), .Z(odata[268]));
Q_MX04 U2167 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][289] ), .A1(\_zzLB[1][289] ), .A2(\_zzLB[2][289] ), .A3(\_zzLB[3][289] ), .Z(odata[269]));
Q_MX04 U2168 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][290] ), .A1(\_zzLB[1][290] ), .A2(\_zzLB[2][290] ), .A3(\_zzLB[3][290] ), .Z(odata[270]));
Q_MX04 U2169 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][291] ), .A1(\_zzLB[1][291] ), .A2(\_zzLB[2][291] ), .A3(\_zzLB[3][291] ), .Z(odata[271]));
Q_MX04 U2170 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][292] ), .A1(\_zzLB[1][292] ), .A2(\_zzLB[2][292] ), .A3(\_zzLB[3][292] ), .Z(odata[272]));
Q_MX04 U2171 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][293] ), .A1(\_zzLB[1][293] ), .A2(\_zzLB[2][293] ), .A3(\_zzLB[3][293] ), .Z(odata[273]));
Q_MX04 U2172 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][294] ), .A1(\_zzLB[1][294] ), .A2(\_zzLB[2][294] ), .A3(\_zzLB[3][294] ), .Z(odata[274]));
Q_MX04 U2173 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][295] ), .A1(\_zzLB[1][295] ), .A2(\_zzLB[2][295] ), .A3(\_zzLB[3][295] ), .Z(odata[275]));
Q_MX04 U2174 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][296] ), .A1(\_zzLB[1][296] ), .A2(\_zzLB[2][296] ), .A3(\_zzLB[3][296] ), .Z(odata[276]));
Q_MX04 U2175 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][297] ), .A1(\_zzLB[1][297] ), .A2(\_zzLB[2][297] ), .A3(\_zzLB[3][297] ), .Z(odata[277]));
Q_MX04 U2176 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][298] ), .A1(\_zzLB[1][298] ), .A2(\_zzLB[2][298] ), .A3(\_zzLB[3][298] ), .Z(odata[278]));
Q_MX04 U2177 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][299] ), .A1(\_zzLB[1][299] ), .A2(\_zzLB[2][299] ), .A3(\_zzLB[3][299] ), .Z(odata[279]));
Q_MX04 U2178 ( .S0(CLBrd[0]), .S1(CLBrd[1]), .A0(\_zzLB[0][300] ), .A1(\_zzLB[1][300] ), .A2(\_zzLB[2][300] ), .A3(\_zzLB[3][300] ), .Z(oreq));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "_zzLB 1 300 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_gfifo_port"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
