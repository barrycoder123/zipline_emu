
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_tlv_inspector_xcm69 ( kme_internal_out_ack, .gcm_cmd_in( {
	\gcm_cmd_in.key0 [255], \gcm_cmd_in.key0 [254], 
	\gcm_cmd_in.key0 [253], \gcm_cmd_in.key0 [252], 
	\gcm_cmd_in.key0 [251], \gcm_cmd_in.key0 [250], 
	\gcm_cmd_in.key0 [249], \gcm_cmd_in.key0 [248], 
	\gcm_cmd_in.key0 [247], \gcm_cmd_in.key0 [246], 
	\gcm_cmd_in.key0 [245], \gcm_cmd_in.key0 [244], 
	\gcm_cmd_in.key0 [243], \gcm_cmd_in.key0 [242], 
	\gcm_cmd_in.key0 [241], \gcm_cmd_in.key0 [240], 
	\gcm_cmd_in.key0 [239], \gcm_cmd_in.key0 [238], 
	\gcm_cmd_in.key0 [237], \gcm_cmd_in.key0 [236], 
	\gcm_cmd_in.key0 [235], \gcm_cmd_in.key0 [234], 
	\gcm_cmd_in.key0 [233], \gcm_cmd_in.key0 [232], 
	\gcm_cmd_in.key0 [231], \gcm_cmd_in.key0 [230], 
	\gcm_cmd_in.key0 [229], \gcm_cmd_in.key0 [228], 
	\gcm_cmd_in.key0 [227], \gcm_cmd_in.key0 [226], 
	\gcm_cmd_in.key0 [225], \gcm_cmd_in.key0 [224], 
	\gcm_cmd_in.key0 [223], \gcm_cmd_in.key0 [222], 
	\gcm_cmd_in.key0 [221], \gcm_cmd_in.key0 [220], 
	\gcm_cmd_in.key0 [219], \gcm_cmd_in.key0 [218], 
	\gcm_cmd_in.key0 [217], \gcm_cmd_in.key0 [216], 
	\gcm_cmd_in.key0 [215], \gcm_cmd_in.key0 [214], 
	\gcm_cmd_in.key0 [213], \gcm_cmd_in.key0 [212], 
	\gcm_cmd_in.key0 [211], \gcm_cmd_in.key0 [210], 
	\gcm_cmd_in.key0 [209], \gcm_cmd_in.key0 [208], 
	\gcm_cmd_in.key0 [207], \gcm_cmd_in.key0 [206], 
	\gcm_cmd_in.key0 [205], \gcm_cmd_in.key0 [204], 
	\gcm_cmd_in.key0 [203], \gcm_cmd_in.key0 [202], 
	\gcm_cmd_in.key0 [201], \gcm_cmd_in.key0 [200], 
	\gcm_cmd_in.key0 [199], \gcm_cmd_in.key0 [198], 
	\gcm_cmd_in.key0 [197], \gcm_cmd_in.key0 [196], 
	\gcm_cmd_in.key0 [195], \gcm_cmd_in.key0 [194], 
	\gcm_cmd_in.key0 [193], \gcm_cmd_in.key0 [192], 
	\gcm_cmd_in.key0 [191], \gcm_cmd_in.key0 [190], 
	\gcm_cmd_in.key0 [189], \gcm_cmd_in.key0 [188], 
	\gcm_cmd_in.key0 [187], \gcm_cmd_in.key0 [186], 
	\gcm_cmd_in.key0 [185], \gcm_cmd_in.key0 [184], 
	\gcm_cmd_in.key0 [183], \gcm_cmd_in.key0 [182], 
	\gcm_cmd_in.key0 [181], \gcm_cmd_in.key0 [180], 
	\gcm_cmd_in.key0 [179], \gcm_cmd_in.key0 [178], 
	\gcm_cmd_in.key0 [177], \gcm_cmd_in.key0 [176], 
	\gcm_cmd_in.key0 [175], \gcm_cmd_in.key0 [174], 
	\gcm_cmd_in.key0 [173], \gcm_cmd_in.key0 [172], 
	\gcm_cmd_in.key0 [171], \gcm_cmd_in.key0 [170], 
	\gcm_cmd_in.key0 [169], \gcm_cmd_in.key0 [168], 
	\gcm_cmd_in.key0 [167], \gcm_cmd_in.key0 [166], 
	\gcm_cmd_in.key0 [165], \gcm_cmd_in.key0 [164], 
	\gcm_cmd_in.key0 [163], \gcm_cmd_in.key0 [162], 
	\gcm_cmd_in.key0 [161], \gcm_cmd_in.key0 [160], 
	\gcm_cmd_in.key0 [159], \gcm_cmd_in.key0 [158], 
	\gcm_cmd_in.key0 [157], \gcm_cmd_in.key0 [156], 
	\gcm_cmd_in.key0 [155], \gcm_cmd_in.key0 [154], 
	\gcm_cmd_in.key0 [153], \gcm_cmd_in.key0 [152], 
	\gcm_cmd_in.key0 [151], \gcm_cmd_in.key0 [150], 
	\gcm_cmd_in.key0 [149], \gcm_cmd_in.key0 [148], 
	\gcm_cmd_in.key0 [147], \gcm_cmd_in.key0 [146], 
	\gcm_cmd_in.key0 [145], \gcm_cmd_in.key0 [144], 
	\gcm_cmd_in.key0 [143], \gcm_cmd_in.key0 [142], 
	\gcm_cmd_in.key0 [141], \gcm_cmd_in.key0 [140], 
	\gcm_cmd_in.key0 [139], \gcm_cmd_in.key0 [138], 
	\gcm_cmd_in.key0 [137], \gcm_cmd_in.key0 [136], 
	\gcm_cmd_in.key0 [135], \gcm_cmd_in.key0 [134], 
	\gcm_cmd_in.key0 [133], \gcm_cmd_in.key0 [132], 
	\gcm_cmd_in.key0 [131], \gcm_cmd_in.key0 [130], 
	\gcm_cmd_in.key0 [129], \gcm_cmd_in.key0 [128], 
	\gcm_cmd_in.key0 [127], \gcm_cmd_in.key0 [126], 
	\gcm_cmd_in.key0 [125], \gcm_cmd_in.key0 [124], 
	\gcm_cmd_in.key0 [123], \gcm_cmd_in.key0 [122], 
	\gcm_cmd_in.key0 [121], \gcm_cmd_in.key0 [120], 
	\gcm_cmd_in.key0 [119], \gcm_cmd_in.key0 [118], 
	\gcm_cmd_in.key0 [117], \gcm_cmd_in.key0 [116], 
	\gcm_cmd_in.key0 [115], \gcm_cmd_in.key0 [114], 
	\gcm_cmd_in.key0 [113], \gcm_cmd_in.key0 [112], 
	\gcm_cmd_in.key0 [111], \gcm_cmd_in.key0 [110], 
	\gcm_cmd_in.key0 [109], \gcm_cmd_in.key0 [108], 
	\gcm_cmd_in.key0 [107], \gcm_cmd_in.key0 [106], 
	\gcm_cmd_in.key0 [105], \gcm_cmd_in.key0 [104], 
	\gcm_cmd_in.key0 [103], \gcm_cmd_in.key0 [102], 
	\gcm_cmd_in.key0 [101], \gcm_cmd_in.key0 [100], 
	\gcm_cmd_in.key0 [99], \gcm_cmd_in.key0 [98], \gcm_cmd_in.key0 [97], 
	\gcm_cmd_in.key0 [96], \gcm_cmd_in.key0 [95], \gcm_cmd_in.key0 [94], 
	\gcm_cmd_in.key0 [93], \gcm_cmd_in.key0 [92], \gcm_cmd_in.key0 [91], 
	\gcm_cmd_in.key0 [90], \gcm_cmd_in.key0 [89], \gcm_cmd_in.key0 [88], 
	\gcm_cmd_in.key0 [87], \gcm_cmd_in.key0 [86], \gcm_cmd_in.key0 [85], 
	\gcm_cmd_in.key0 [84], \gcm_cmd_in.key0 [83], \gcm_cmd_in.key0 [82], 
	\gcm_cmd_in.key0 [81], \gcm_cmd_in.key0 [80], \gcm_cmd_in.key0 [79], 
	\gcm_cmd_in.key0 [78], \gcm_cmd_in.key0 [77], \gcm_cmd_in.key0 [76], 
	\gcm_cmd_in.key0 [75], \gcm_cmd_in.key0 [74], \gcm_cmd_in.key0 [73], 
	\gcm_cmd_in.key0 [72], \gcm_cmd_in.key0 [71], \gcm_cmd_in.key0 [70], 
	\gcm_cmd_in.key0 [69], \gcm_cmd_in.key0 [68], \gcm_cmd_in.key0 [67], 
	\gcm_cmd_in.key0 [66], \gcm_cmd_in.key0 [65], \gcm_cmd_in.key0 [64], 
	\gcm_cmd_in.key0 [63], \gcm_cmd_in.key0 [62], \gcm_cmd_in.key0 [61], 
	\gcm_cmd_in.key0 [60], \gcm_cmd_in.key0 [59], \gcm_cmd_in.key0 [58], 
	\gcm_cmd_in.key0 [57], \gcm_cmd_in.key0 [56], \gcm_cmd_in.key0 [55], 
	\gcm_cmd_in.key0 [54], \gcm_cmd_in.key0 [53], \gcm_cmd_in.key0 [52], 
	\gcm_cmd_in.key0 [51], \gcm_cmd_in.key0 [50], \gcm_cmd_in.key0 [49], 
	\gcm_cmd_in.key0 [48], \gcm_cmd_in.key0 [47], \gcm_cmd_in.key0 [46], 
	\gcm_cmd_in.key0 [45], \gcm_cmd_in.key0 [44], \gcm_cmd_in.key0 [43], 
	\gcm_cmd_in.key0 [42], \gcm_cmd_in.key0 [41], \gcm_cmd_in.key0 [40], 
	\gcm_cmd_in.key0 [39], \gcm_cmd_in.key0 [38], \gcm_cmd_in.key0 [37], 
	\gcm_cmd_in.key0 [36], \gcm_cmd_in.key0 [35], \gcm_cmd_in.key0 [34], 
	\gcm_cmd_in.key0 [33], \gcm_cmd_in.key0 [32], \gcm_cmd_in.key0 [31], 
	\gcm_cmd_in.key0 [30], \gcm_cmd_in.key0 [29], \gcm_cmd_in.key0 [28], 
	\gcm_cmd_in.key0 [27], \gcm_cmd_in.key0 [26], \gcm_cmd_in.key0 [25], 
	\gcm_cmd_in.key0 [24], \gcm_cmd_in.key0 [23], \gcm_cmd_in.key0 [22], 
	\gcm_cmd_in.key0 [21], \gcm_cmd_in.key0 [20], \gcm_cmd_in.key0 [19], 
	\gcm_cmd_in.key0 [18], \gcm_cmd_in.key0 [17], \gcm_cmd_in.key0 [16], 
	\gcm_cmd_in.key0 [15], \gcm_cmd_in.key0 [14], \gcm_cmd_in.key0 [13], 
	\gcm_cmd_in.key0 [12], \gcm_cmd_in.key0 [11], \gcm_cmd_in.key0 [10], 
	\gcm_cmd_in.key0 [9], \gcm_cmd_in.key0 [8], \gcm_cmd_in.key0 [7], 
	\gcm_cmd_in.key0 [6], \gcm_cmd_in.key0 [5], \gcm_cmd_in.key0 [4], 
	\gcm_cmd_in.key0 [3], \gcm_cmd_in.key0 [2], \gcm_cmd_in.key0 [1], 
	\gcm_cmd_in.key0 [0], \gcm_cmd_in.key1 [255], \gcm_cmd_in.key1 [254], 
	\gcm_cmd_in.key1 [253], \gcm_cmd_in.key1 [252], 
	\gcm_cmd_in.key1 [251], \gcm_cmd_in.key1 [250], 
	\gcm_cmd_in.key1 [249], \gcm_cmd_in.key1 [248], 
	\gcm_cmd_in.key1 [247], \gcm_cmd_in.key1 [246], 
	\gcm_cmd_in.key1 [245], \gcm_cmd_in.key1 [244], 
	\gcm_cmd_in.key1 [243], \gcm_cmd_in.key1 [242], 
	\gcm_cmd_in.key1 [241], \gcm_cmd_in.key1 [240], 
	\gcm_cmd_in.key1 [239], \gcm_cmd_in.key1 [238], 
	\gcm_cmd_in.key1 [237], \gcm_cmd_in.key1 [236], 
	\gcm_cmd_in.key1 [235], \gcm_cmd_in.key1 [234], 
	\gcm_cmd_in.key1 [233], \gcm_cmd_in.key1 [232], 
	\gcm_cmd_in.key1 [231], \gcm_cmd_in.key1 [230], 
	\gcm_cmd_in.key1 [229], \gcm_cmd_in.key1 [228], 
	\gcm_cmd_in.key1 [227], \gcm_cmd_in.key1 [226], 
	\gcm_cmd_in.key1 [225], \gcm_cmd_in.key1 [224], 
	\gcm_cmd_in.key1 [223], \gcm_cmd_in.key1 [222], 
	\gcm_cmd_in.key1 [221], \gcm_cmd_in.key1 [220], 
	\gcm_cmd_in.key1 [219], \gcm_cmd_in.key1 [218], 
	\gcm_cmd_in.key1 [217], \gcm_cmd_in.key1 [216], 
	\gcm_cmd_in.key1 [215], \gcm_cmd_in.key1 [214], 
	\gcm_cmd_in.key1 [213], \gcm_cmd_in.key1 [212], 
	\gcm_cmd_in.key1 [211], \gcm_cmd_in.key1 [210], 
	\gcm_cmd_in.key1 [209], \gcm_cmd_in.key1 [208], 
	\gcm_cmd_in.key1 [207], \gcm_cmd_in.key1 [206], 
	\gcm_cmd_in.key1 [205], \gcm_cmd_in.key1 [204], 
	\gcm_cmd_in.key1 [203], \gcm_cmd_in.key1 [202], 
	\gcm_cmd_in.key1 [201], \gcm_cmd_in.key1 [200], 
	\gcm_cmd_in.key1 [199], \gcm_cmd_in.key1 [198], 
	\gcm_cmd_in.key1 [197], \gcm_cmd_in.key1 [196], 
	\gcm_cmd_in.key1 [195], \gcm_cmd_in.key1 [194], 
	\gcm_cmd_in.key1 [193], \gcm_cmd_in.key1 [192], 
	\gcm_cmd_in.key1 [191], \gcm_cmd_in.key1 [190], 
	\gcm_cmd_in.key1 [189], \gcm_cmd_in.key1 [188], 
	\gcm_cmd_in.key1 [187], \gcm_cmd_in.key1 [186], 
	\gcm_cmd_in.key1 [185], \gcm_cmd_in.key1 [184], 
	\gcm_cmd_in.key1 [183], \gcm_cmd_in.key1 [182], 
	\gcm_cmd_in.key1 [181], \gcm_cmd_in.key1 [180], 
	\gcm_cmd_in.key1 [179], \gcm_cmd_in.key1 [178], 
	\gcm_cmd_in.key1 [177], \gcm_cmd_in.key1 [176], 
	\gcm_cmd_in.key1 [175], \gcm_cmd_in.key1 [174], 
	\gcm_cmd_in.key1 [173], \gcm_cmd_in.key1 [172], 
	\gcm_cmd_in.key1 [171], \gcm_cmd_in.key1 [170], 
	\gcm_cmd_in.key1 [169], \gcm_cmd_in.key1 [168], 
	\gcm_cmd_in.key1 [167], \gcm_cmd_in.key1 [166], 
	\gcm_cmd_in.key1 [165], \gcm_cmd_in.key1 [164], 
	\gcm_cmd_in.key1 [163], \gcm_cmd_in.key1 [162], 
	\gcm_cmd_in.key1 [161], \gcm_cmd_in.key1 [160], 
	\gcm_cmd_in.key1 [159], \gcm_cmd_in.key1 [158], 
	\gcm_cmd_in.key1 [157], \gcm_cmd_in.key1 [156], 
	\gcm_cmd_in.key1 [155], \gcm_cmd_in.key1 [154], 
	\gcm_cmd_in.key1 [153], \gcm_cmd_in.key1 [152], 
	\gcm_cmd_in.key1 [151], \gcm_cmd_in.key1 [150], 
	\gcm_cmd_in.key1 [149], \gcm_cmd_in.key1 [148], 
	\gcm_cmd_in.key1 [147], \gcm_cmd_in.key1 [146], 
	\gcm_cmd_in.key1 [145], \gcm_cmd_in.key1 [144], 
	\gcm_cmd_in.key1 [143], \gcm_cmd_in.key1 [142], 
	\gcm_cmd_in.key1 [141], \gcm_cmd_in.key1 [140], 
	\gcm_cmd_in.key1 [139], \gcm_cmd_in.key1 [138], 
	\gcm_cmd_in.key1 [137], \gcm_cmd_in.key1 [136], 
	\gcm_cmd_in.key1 [135], \gcm_cmd_in.key1 [134], 
	\gcm_cmd_in.key1 [133], \gcm_cmd_in.key1 [132], 
	\gcm_cmd_in.key1 [131], \gcm_cmd_in.key1 [130], 
	\gcm_cmd_in.key1 [129], \gcm_cmd_in.key1 [128], 
	\gcm_cmd_in.key1 [127], \gcm_cmd_in.key1 [126], 
	\gcm_cmd_in.key1 [125], \gcm_cmd_in.key1 [124], 
	\gcm_cmd_in.key1 [123], \gcm_cmd_in.key1 [122], 
	\gcm_cmd_in.key1 [121], \gcm_cmd_in.key1 [120], 
	\gcm_cmd_in.key1 [119], \gcm_cmd_in.key1 [118], 
	\gcm_cmd_in.key1 [117], \gcm_cmd_in.key1 [116], 
	\gcm_cmd_in.key1 [115], \gcm_cmd_in.key1 [114], 
	\gcm_cmd_in.key1 [113], \gcm_cmd_in.key1 [112], 
	\gcm_cmd_in.key1 [111], \gcm_cmd_in.key1 [110], 
	\gcm_cmd_in.key1 [109], \gcm_cmd_in.key1 [108], 
	\gcm_cmd_in.key1 [107], \gcm_cmd_in.key1 [106], 
	\gcm_cmd_in.key1 [105], \gcm_cmd_in.key1 [104], 
	\gcm_cmd_in.key1 [103], \gcm_cmd_in.key1 [102], 
	\gcm_cmd_in.key1 [101], \gcm_cmd_in.key1 [100], 
	\gcm_cmd_in.key1 [99], \gcm_cmd_in.key1 [98], \gcm_cmd_in.key1 [97], 
	\gcm_cmd_in.key1 [96], \gcm_cmd_in.key1 [95], \gcm_cmd_in.key1 [94], 
	\gcm_cmd_in.key1 [93], \gcm_cmd_in.key1 [92], \gcm_cmd_in.key1 [91], 
	\gcm_cmd_in.key1 [90], \gcm_cmd_in.key1 [89], \gcm_cmd_in.key1 [88], 
	\gcm_cmd_in.key1 [87], \gcm_cmd_in.key1 [86], \gcm_cmd_in.key1 [85], 
	\gcm_cmd_in.key1 [84], \gcm_cmd_in.key1 [83], \gcm_cmd_in.key1 [82], 
	\gcm_cmd_in.key1 [81], \gcm_cmd_in.key1 [80], \gcm_cmd_in.key1 [79], 
	\gcm_cmd_in.key1 [78], \gcm_cmd_in.key1 [77], \gcm_cmd_in.key1 [76], 
	\gcm_cmd_in.key1 [75], \gcm_cmd_in.key1 [74], \gcm_cmd_in.key1 [73], 
	\gcm_cmd_in.key1 [72], \gcm_cmd_in.key1 [71], \gcm_cmd_in.key1 [70], 
	\gcm_cmd_in.key1 [69], \gcm_cmd_in.key1 [68], \gcm_cmd_in.key1 [67], 
	\gcm_cmd_in.key1 [66], \gcm_cmd_in.key1 [65], \gcm_cmd_in.key1 [64], 
	\gcm_cmd_in.key1 [63], \gcm_cmd_in.key1 [62], \gcm_cmd_in.key1 [61], 
	\gcm_cmd_in.key1 [60], \gcm_cmd_in.key1 [59], \gcm_cmd_in.key1 [58], 
	\gcm_cmd_in.key1 [57], \gcm_cmd_in.key1 [56], \gcm_cmd_in.key1 [55], 
	\gcm_cmd_in.key1 [54], \gcm_cmd_in.key1 [53], \gcm_cmd_in.key1 [52], 
	\gcm_cmd_in.key1 [51], \gcm_cmd_in.key1 [50], \gcm_cmd_in.key1 [49], 
	\gcm_cmd_in.key1 [48], \gcm_cmd_in.key1 [47], \gcm_cmd_in.key1 [46], 
	\gcm_cmd_in.key1 [45], \gcm_cmd_in.key1 [44], \gcm_cmd_in.key1 [43], 
	\gcm_cmd_in.key1 [42], \gcm_cmd_in.key1 [41], \gcm_cmd_in.key1 [40], 
	\gcm_cmd_in.key1 [39], \gcm_cmd_in.key1 [38], \gcm_cmd_in.key1 [37], 
	\gcm_cmd_in.key1 [36], \gcm_cmd_in.key1 [35], \gcm_cmd_in.key1 [34], 
	\gcm_cmd_in.key1 [33], \gcm_cmd_in.key1 [32], \gcm_cmd_in.key1 [31], 
	\gcm_cmd_in.key1 [30], \gcm_cmd_in.key1 [29], \gcm_cmd_in.key1 [28], 
	\gcm_cmd_in.key1 [27], \gcm_cmd_in.key1 [26], \gcm_cmd_in.key1 [25], 
	\gcm_cmd_in.key1 [24], \gcm_cmd_in.key1 [23], \gcm_cmd_in.key1 [22], 
	\gcm_cmd_in.key1 [21], \gcm_cmd_in.key1 [20], \gcm_cmd_in.key1 [19], 
	\gcm_cmd_in.key1 [18], \gcm_cmd_in.key1 [17], \gcm_cmd_in.key1 [16], 
	\gcm_cmd_in.key1 [15], \gcm_cmd_in.key1 [14], \gcm_cmd_in.key1 [13], 
	\gcm_cmd_in.key1 [12], \gcm_cmd_in.key1 [11], \gcm_cmd_in.key1 [10], 
	\gcm_cmd_in.key1 [9], \gcm_cmd_in.key1 [8], \gcm_cmd_in.key1 [7], 
	\gcm_cmd_in.key1 [6], \gcm_cmd_in.key1 [5], \gcm_cmd_in.key1 [4], 
	\gcm_cmd_in.key1 [3], \gcm_cmd_in.key1 [2], \gcm_cmd_in.key1 [1], 
	\gcm_cmd_in.key1 [0], \gcm_cmd_in.iv [95], \gcm_cmd_in.iv [94], 
	\gcm_cmd_in.iv [93], \gcm_cmd_in.iv [92], \gcm_cmd_in.iv [91], 
	\gcm_cmd_in.iv [90], \gcm_cmd_in.iv [89], \gcm_cmd_in.iv [88], 
	\gcm_cmd_in.iv [87], \gcm_cmd_in.iv [86], \gcm_cmd_in.iv [85], 
	\gcm_cmd_in.iv [84], \gcm_cmd_in.iv [83], \gcm_cmd_in.iv [82], 
	\gcm_cmd_in.iv [81], \gcm_cmd_in.iv [80], \gcm_cmd_in.iv [79], 
	\gcm_cmd_in.iv [78], \gcm_cmd_in.iv [77], \gcm_cmd_in.iv [76], 
	\gcm_cmd_in.iv [75], \gcm_cmd_in.iv [74], \gcm_cmd_in.iv [73], 
	\gcm_cmd_in.iv [72], \gcm_cmd_in.iv [71], \gcm_cmd_in.iv [70], 
	\gcm_cmd_in.iv [69], \gcm_cmd_in.iv [68], \gcm_cmd_in.iv [67], 
	\gcm_cmd_in.iv [66], \gcm_cmd_in.iv [65], \gcm_cmd_in.iv [64], 
	\gcm_cmd_in.iv [63], \gcm_cmd_in.iv [62], \gcm_cmd_in.iv [61], 
	\gcm_cmd_in.iv [60], \gcm_cmd_in.iv [59], \gcm_cmd_in.iv [58], 
	\gcm_cmd_in.iv [57], \gcm_cmd_in.iv [56], \gcm_cmd_in.iv [55], 
	\gcm_cmd_in.iv [54], \gcm_cmd_in.iv [53], \gcm_cmd_in.iv [52], 
	\gcm_cmd_in.iv [51], \gcm_cmd_in.iv [50], \gcm_cmd_in.iv [49], 
	\gcm_cmd_in.iv [48], \gcm_cmd_in.iv [47], \gcm_cmd_in.iv [46], 
	\gcm_cmd_in.iv [45], \gcm_cmd_in.iv [44], \gcm_cmd_in.iv [43], 
	\gcm_cmd_in.iv [42], \gcm_cmd_in.iv [41], \gcm_cmd_in.iv [40], 
	\gcm_cmd_in.iv [39], \gcm_cmd_in.iv [38], \gcm_cmd_in.iv [37], 
	\gcm_cmd_in.iv [36], \gcm_cmd_in.iv [35], \gcm_cmd_in.iv [34], 
	\gcm_cmd_in.iv [33], \gcm_cmd_in.iv [32], \gcm_cmd_in.iv [31], 
	\gcm_cmd_in.iv [30], \gcm_cmd_in.iv [29], \gcm_cmd_in.iv [28], 
	\gcm_cmd_in.iv [27], \gcm_cmd_in.iv [26], \gcm_cmd_in.iv [25], 
	\gcm_cmd_in.iv [24], \gcm_cmd_in.iv [23], \gcm_cmd_in.iv [22], 
	\gcm_cmd_in.iv [21], \gcm_cmd_in.iv [20], \gcm_cmd_in.iv [19], 
	\gcm_cmd_in.iv [18], \gcm_cmd_in.iv [17], \gcm_cmd_in.iv [16], 
	\gcm_cmd_in.iv [15], \gcm_cmd_in.iv [14], \gcm_cmd_in.iv [13], 
	\gcm_cmd_in.iv [12], \gcm_cmd_in.iv [11], \gcm_cmd_in.iv [10], 
	\gcm_cmd_in.iv [9], \gcm_cmd_in.iv [8], \gcm_cmd_in.iv [7], 
	\gcm_cmd_in.iv [6], \gcm_cmd_in.iv [5], \gcm_cmd_in.iv [4], 
	\gcm_cmd_in.iv [3], \gcm_cmd_in.iv [2], \gcm_cmd_in.iv [1], 
	\gcm_cmd_in.iv [0], \gcm_cmd_in.op [2], \gcm_cmd_in.op [1], 
	\gcm_cmd_in.op [0]} ), gcm_cmd_in_valid, gcm_tag_data_in, 
	gcm_tag_data_in_valid, inspector_upsizer_valid, 
	inspector_upsizer_eof, inspector_upsizer_data, .keyfilter_cmd_in( {
	\keyfilter_cmd_in.combo_mode [0]} ), keyfilter_cmd_in_valid, 
	.kdfstream_cmd_in( {\kdfstream_cmd_in.combo_mode [0], 
	\kdfstream_cmd_in.skip [0], \kdfstream_cmd_in.guid [255], 
	\kdfstream_cmd_in.guid [254], \kdfstream_cmd_in.guid [253], 
	\kdfstream_cmd_in.guid [252], \kdfstream_cmd_in.guid [251], 
	\kdfstream_cmd_in.guid [250], \kdfstream_cmd_in.guid [249], 
	\kdfstream_cmd_in.guid [248], \kdfstream_cmd_in.guid [247], 
	\kdfstream_cmd_in.guid [246], \kdfstream_cmd_in.guid [245], 
	\kdfstream_cmd_in.guid [244], \kdfstream_cmd_in.guid [243], 
	\kdfstream_cmd_in.guid [242], \kdfstream_cmd_in.guid [241], 
	\kdfstream_cmd_in.guid [240], \kdfstream_cmd_in.guid [239], 
	\kdfstream_cmd_in.guid [238], \kdfstream_cmd_in.guid [237], 
	\kdfstream_cmd_in.guid [236], \kdfstream_cmd_in.guid [235], 
	\kdfstream_cmd_in.guid [234], \kdfstream_cmd_in.guid [233], 
	\kdfstream_cmd_in.guid [232], \kdfstream_cmd_in.guid [231], 
	\kdfstream_cmd_in.guid [230], \kdfstream_cmd_in.guid [229], 
	\kdfstream_cmd_in.guid [228], \kdfstream_cmd_in.guid [227], 
	\kdfstream_cmd_in.guid [226], \kdfstream_cmd_in.guid [225], 
	\kdfstream_cmd_in.guid [224], \kdfstream_cmd_in.guid [223], 
	\kdfstream_cmd_in.guid [222], \kdfstream_cmd_in.guid [221], 
	\kdfstream_cmd_in.guid [220], \kdfstream_cmd_in.guid [219], 
	\kdfstream_cmd_in.guid [218], \kdfstream_cmd_in.guid [217], 
	\kdfstream_cmd_in.guid [216], \kdfstream_cmd_in.guid [215], 
	\kdfstream_cmd_in.guid [214], \kdfstream_cmd_in.guid [213], 
	\kdfstream_cmd_in.guid [212], \kdfstream_cmd_in.guid [211], 
	\kdfstream_cmd_in.guid [210], \kdfstream_cmd_in.guid [209], 
	\kdfstream_cmd_in.guid [208], \kdfstream_cmd_in.guid [207], 
	\kdfstream_cmd_in.guid [206], \kdfstream_cmd_in.guid [205], 
	\kdfstream_cmd_in.guid [204], \kdfstream_cmd_in.guid [203], 
	\kdfstream_cmd_in.guid [202], \kdfstream_cmd_in.guid [201], 
	\kdfstream_cmd_in.guid [200], \kdfstream_cmd_in.guid [199], 
	\kdfstream_cmd_in.guid [198], \kdfstream_cmd_in.guid [197], 
	\kdfstream_cmd_in.guid [196], \kdfstream_cmd_in.guid [195], 
	\kdfstream_cmd_in.guid [194], \kdfstream_cmd_in.guid [193], 
	\kdfstream_cmd_in.guid [192], \kdfstream_cmd_in.guid [191], 
	\kdfstream_cmd_in.guid [190], \kdfstream_cmd_in.guid [189], 
	\kdfstream_cmd_in.guid [188], \kdfstream_cmd_in.guid [187], 
	\kdfstream_cmd_in.guid [186], \kdfstream_cmd_in.guid [185], 
	\kdfstream_cmd_in.guid [184], \kdfstream_cmd_in.guid [183], 
	\kdfstream_cmd_in.guid [182], \kdfstream_cmd_in.guid [181], 
	\kdfstream_cmd_in.guid [180], \kdfstream_cmd_in.guid [179], 
	\kdfstream_cmd_in.guid [178], \kdfstream_cmd_in.guid [177], 
	\kdfstream_cmd_in.guid [176], \kdfstream_cmd_in.guid [175], 
	\kdfstream_cmd_in.guid [174], \kdfstream_cmd_in.guid [173], 
	\kdfstream_cmd_in.guid [172], \kdfstream_cmd_in.guid [171], 
	\kdfstream_cmd_in.guid [170], \kdfstream_cmd_in.guid [169], 
	\kdfstream_cmd_in.guid [168], \kdfstream_cmd_in.guid [167], 
	\kdfstream_cmd_in.guid [166], \kdfstream_cmd_in.guid [165], 
	\kdfstream_cmd_in.guid [164], \kdfstream_cmd_in.guid [163], 
	\kdfstream_cmd_in.guid [162], \kdfstream_cmd_in.guid [161], 
	\kdfstream_cmd_in.guid [160], \kdfstream_cmd_in.guid [159], 
	\kdfstream_cmd_in.guid [158], \kdfstream_cmd_in.guid [157], 
	\kdfstream_cmd_in.guid [156], \kdfstream_cmd_in.guid [155], 
	\kdfstream_cmd_in.guid [154], \kdfstream_cmd_in.guid [153], 
	\kdfstream_cmd_in.guid [152], \kdfstream_cmd_in.guid [151], 
	\kdfstream_cmd_in.guid [150], \kdfstream_cmd_in.guid [149], 
	\kdfstream_cmd_in.guid [148], \kdfstream_cmd_in.guid [147], 
	\kdfstream_cmd_in.guid [146], \kdfstream_cmd_in.guid [145], 
	\kdfstream_cmd_in.guid [144], \kdfstream_cmd_in.guid [143], 
	\kdfstream_cmd_in.guid [142], \kdfstream_cmd_in.guid [141], 
	\kdfstream_cmd_in.guid [140], \kdfstream_cmd_in.guid [139], 
	\kdfstream_cmd_in.guid [138], \kdfstream_cmd_in.guid [137], 
	\kdfstream_cmd_in.guid [136], \kdfstream_cmd_in.guid [135], 
	\kdfstream_cmd_in.guid [134], \kdfstream_cmd_in.guid [133], 
	\kdfstream_cmd_in.guid [132], \kdfstream_cmd_in.guid [131], 
	\kdfstream_cmd_in.guid [130], \kdfstream_cmd_in.guid [129], 
	\kdfstream_cmd_in.guid [128], \kdfstream_cmd_in.guid [127], 
	\kdfstream_cmd_in.guid [126], \kdfstream_cmd_in.guid [125], 
	\kdfstream_cmd_in.guid [124], \kdfstream_cmd_in.guid [123], 
	\kdfstream_cmd_in.guid [122], \kdfstream_cmd_in.guid [121], 
	\kdfstream_cmd_in.guid [120], \kdfstream_cmd_in.guid [119], 
	\kdfstream_cmd_in.guid [118], \kdfstream_cmd_in.guid [117], 
	\kdfstream_cmd_in.guid [116], \kdfstream_cmd_in.guid [115], 
	\kdfstream_cmd_in.guid [114], \kdfstream_cmd_in.guid [113], 
	\kdfstream_cmd_in.guid [112], \kdfstream_cmd_in.guid [111], 
	\kdfstream_cmd_in.guid [110], \kdfstream_cmd_in.guid [109], 
	\kdfstream_cmd_in.guid [108], \kdfstream_cmd_in.guid [107], 
	\kdfstream_cmd_in.guid [106], \kdfstream_cmd_in.guid [105], 
	\kdfstream_cmd_in.guid [104], \kdfstream_cmd_in.guid [103], 
	\kdfstream_cmd_in.guid [102], \kdfstream_cmd_in.guid [101], 
	\kdfstream_cmd_in.guid [100], \kdfstream_cmd_in.guid [99], 
	\kdfstream_cmd_in.guid [98], \kdfstream_cmd_in.guid [97], 
	\kdfstream_cmd_in.guid [96], \kdfstream_cmd_in.guid [95], 
	\kdfstream_cmd_in.guid [94], \kdfstream_cmd_in.guid [93], 
	\kdfstream_cmd_in.guid [92], \kdfstream_cmd_in.guid [91], 
	\kdfstream_cmd_in.guid [90], \kdfstream_cmd_in.guid [89], 
	\kdfstream_cmd_in.guid [88], \kdfstream_cmd_in.guid [87], 
	\kdfstream_cmd_in.guid [86], \kdfstream_cmd_in.guid [85], 
	\kdfstream_cmd_in.guid [84], \kdfstream_cmd_in.guid [83], 
	\kdfstream_cmd_in.guid [82], \kdfstream_cmd_in.guid [81], 
	\kdfstream_cmd_in.guid [80], \kdfstream_cmd_in.guid [79], 
	\kdfstream_cmd_in.guid [78], \kdfstream_cmd_in.guid [77], 
	\kdfstream_cmd_in.guid [76], \kdfstream_cmd_in.guid [75], 
	\kdfstream_cmd_in.guid [74], \kdfstream_cmd_in.guid [73], 
	\kdfstream_cmd_in.guid [72], \kdfstream_cmd_in.guid [71], 
	\kdfstream_cmd_in.guid [70], \kdfstream_cmd_in.guid [69], 
	\kdfstream_cmd_in.guid [68], \kdfstream_cmd_in.guid [67], 
	\kdfstream_cmd_in.guid [66], \kdfstream_cmd_in.guid [65], 
	\kdfstream_cmd_in.guid [64], \kdfstream_cmd_in.guid [63], 
	\kdfstream_cmd_in.guid [62], \kdfstream_cmd_in.guid [61], 
	\kdfstream_cmd_in.guid [60], \kdfstream_cmd_in.guid [59], 
	\kdfstream_cmd_in.guid [58], \kdfstream_cmd_in.guid [57], 
	\kdfstream_cmd_in.guid [56], \kdfstream_cmd_in.guid [55], 
	\kdfstream_cmd_in.guid [54], \kdfstream_cmd_in.guid [53], 
	\kdfstream_cmd_in.guid [52], \kdfstream_cmd_in.guid [51], 
	\kdfstream_cmd_in.guid [50], \kdfstream_cmd_in.guid [49], 
	\kdfstream_cmd_in.guid [48], \kdfstream_cmd_in.guid [47], 
	\kdfstream_cmd_in.guid [46], \kdfstream_cmd_in.guid [45], 
	\kdfstream_cmd_in.guid [44], \kdfstream_cmd_in.guid [43], 
	\kdfstream_cmd_in.guid [42], \kdfstream_cmd_in.guid [41], 
	\kdfstream_cmd_in.guid [40], \kdfstream_cmd_in.guid [39], 
	\kdfstream_cmd_in.guid [38], \kdfstream_cmd_in.guid [37], 
	\kdfstream_cmd_in.guid [36], \kdfstream_cmd_in.guid [35], 
	\kdfstream_cmd_in.guid [34], \kdfstream_cmd_in.guid [33], 
	\kdfstream_cmd_in.guid [32], \kdfstream_cmd_in.guid [31], 
	\kdfstream_cmd_in.guid [30], \kdfstream_cmd_in.guid [29], 
	\kdfstream_cmd_in.guid [28], \kdfstream_cmd_in.guid [27], 
	\kdfstream_cmd_in.guid [26], \kdfstream_cmd_in.guid [25], 
	\kdfstream_cmd_in.guid [24], \kdfstream_cmd_in.guid [23], 
	\kdfstream_cmd_in.guid [22], \kdfstream_cmd_in.guid [21], 
	\kdfstream_cmd_in.guid [20], \kdfstream_cmd_in.guid [19], 
	\kdfstream_cmd_in.guid [18], \kdfstream_cmd_in.guid [17], 
	\kdfstream_cmd_in.guid [16], \kdfstream_cmd_in.guid [15], 
	\kdfstream_cmd_in.guid [14], \kdfstream_cmd_in.guid [13], 
	\kdfstream_cmd_in.guid [12], \kdfstream_cmd_in.guid [11], 
	\kdfstream_cmd_in.guid [10], \kdfstream_cmd_in.guid [9], 
	\kdfstream_cmd_in.guid [8], \kdfstream_cmd_in.guid [7], 
	\kdfstream_cmd_in.guid [6], \kdfstream_cmd_in.guid [5], 
	\kdfstream_cmd_in.guid [4], \kdfstream_cmd_in.guid [3], 
	\kdfstream_cmd_in.guid [2], \kdfstream_cmd_in.guid [1], 
	\kdfstream_cmd_in.guid [0], \kdfstream_cmd_in.label_index [2], 
	\kdfstream_cmd_in.label_index [1], \kdfstream_cmd_in.label_index [0], 
	\kdfstream_cmd_in.num_iter [1], \kdfstream_cmd_in.num_iter [0]} ), 
	kdfstream_cmd_in_valid, .kdf_cmd_in( {\kdf_cmd_in.kdf_dek_iter [0], 
	\kdf_cmd_in.combo_mode [0], \kdf_cmd_in.dek_key_op [0], 
	\kdf_cmd_in.dak_key_op [0]} ), kdf_cmd_in_valid, tlv_sb_data_in, 
	tlv_sb_data_in_valid, clk, rst_n, .labels( {
	\labels[7].guid_size[0] , \labels[7].label_size[5] , 
	\labels[7].label_size[4] , \labels[7].label_size[3] , 
	\labels[7].label_size[2] , \labels[7].label_size[1] , 
	\labels[7].label_size[0] , \labels[7].label[255] , 
	\labels[7].label[254] , \labels[7].label[253] , 
	\labels[7].label[252] , \labels[7].label[251] , 
	\labels[7].label[250] , \labels[7].label[249] , 
	\labels[7].label[248] , \labels[7].label[247] , 
	\labels[7].label[246] , \labels[7].label[245] , 
	\labels[7].label[244] , \labels[7].label[243] , 
	\labels[7].label[242] , \labels[7].label[241] , 
	\labels[7].label[240] , \labels[7].label[239] , 
	\labels[7].label[238] , \labels[7].label[237] , 
	\labels[7].label[236] , \labels[7].label[235] , 
	\labels[7].label[234] , \labels[7].label[233] , 
	\labels[7].label[232] , \labels[7].label[231] , 
	\labels[7].label[230] , \labels[7].label[229] , 
	\labels[7].label[228] , \labels[7].label[227] , 
	\labels[7].label[226] , \labels[7].label[225] , 
	\labels[7].label[224] , \labels[7].label[223] , 
	\labels[7].label[222] , \labels[7].label[221] , 
	\labels[7].label[220] , \labels[7].label[219] , 
	\labels[7].label[218] , \labels[7].label[217] , 
	\labels[7].label[216] , \labels[7].label[215] , 
	\labels[7].label[214] , \labels[7].label[213] , 
	\labels[7].label[212] , \labels[7].label[211] , 
	\labels[7].label[210] , \labels[7].label[209] , 
	\labels[7].label[208] , \labels[7].label[207] , 
	\labels[7].label[206] , \labels[7].label[205] , 
	\labels[7].label[204] , \labels[7].label[203] , 
	\labels[7].label[202] , \labels[7].label[201] , 
	\labels[7].label[200] , \labels[7].label[199] , 
	\labels[7].label[198] , \labels[7].label[197] , 
	\labels[7].label[196] , \labels[7].label[195] , 
	\labels[7].label[194] , \labels[7].label[193] , 
	\labels[7].label[192] , \labels[7].label[191] , 
	\labels[7].label[190] , \labels[7].label[189] , 
	\labels[7].label[188] , \labels[7].label[187] , 
	\labels[7].label[186] , \labels[7].label[185] , 
	\labels[7].label[184] , \labels[7].label[183] , 
	\labels[7].label[182] , \labels[7].label[181] , 
	\labels[7].label[180] , \labels[7].label[179] , 
	\labels[7].label[178] , \labels[7].label[177] , 
	\labels[7].label[176] , \labels[7].label[175] , 
	\labels[7].label[174] , \labels[7].label[173] , 
	\labels[7].label[172] , \labels[7].label[171] , 
	\labels[7].label[170] , \labels[7].label[169] , 
	\labels[7].label[168] , \labels[7].label[167] , 
	\labels[7].label[166] , \labels[7].label[165] , 
	\labels[7].label[164] , \labels[7].label[163] , 
	\labels[7].label[162] , \labels[7].label[161] , 
	\labels[7].label[160] , \labels[7].label[159] , 
	\labels[7].label[158] , \labels[7].label[157] , 
	\labels[7].label[156] , \labels[7].label[155] , 
	\labels[7].label[154] , \labels[7].label[153] , 
	\labels[7].label[152] , \labels[7].label[151] , 
	\labels[7].label[150] , \labels[7].label[149] , 
	\labels[7].label[148] , \labels[7].label[147] , 
	\labels[7].label[146] , \labels[7].label[145] , 
	\labels[7].label[144] , \labels[7].label[143] , 
	\labels[7].label[142] , \labels[7].label[141] , 
	\labels[7].label[140] , \labels[7].label[139] , 
	\labels[7].label[138] , \labels[7].label[137] , 
	\labels[7].label[136] , \labels[7].label[135] , 
	\labels[7].label[134] , \labels[7].label[133] , 
	\labels[7].label[132] , \labels[7].label[131] , 
	\labels[7].label[130] , \labels[7].label[129] , 
	\labels[7].label[128] , \labels[7].label[127] , 
	\labels[7].label[126] , \labels[7].label[125] , 
	\labels[7].label[124] , \labels[7].label[123] , 
	\labels[7].label[122] , \labels[7].label[121] , 
	\labels[7].label[120] , \labels[7].label[119] , 
	\labels[7].label[118] , \labels[7].label[117] , 
	\labels[7].label[116] , \labels[7].label[115] , 
	\labels[7].label[114] , \labels[7].label[113] , 
	\labels[7].label[112] , \labels[7].label[111] , 
	\labels[7].label[110] , \labels[7].label[109] , 
	\labels[7].label[108] , \labels[7].label[107] , 
	\labels[7].label[106] , \labels[7].label[105] , 
	\labels[7].label[104] , \labels[7].label[103] , 
	\labels[7].label[102] , \labels[7].label[101] , 
	\labels[7].label[100] , \labels[7].label[99] , \labels[7].label[98] , 
	\labels[7].label[97] , \labels[7].label[96] , \labels[7].label[95] , 
	\labels[7].label[94] , \labels[7].label[93] , \labels[7].label[92] , 
	\labels[7].label[91] , \labels[7].label[90] , \labels[7].label[89] , 
	\labels[7].label[88] , \labels[7].label[87] , \labels[7].label[86] , 
	\labels[7].label[85] , \labels[7].label[84] , \labels[7].label[83] , 
	\labels[7].label[82] , \labels[7].label[81] , \labels[7].label[80] , 
	\labels[7].label[79] , \labels[7].label[78] , \labels[7].label[77] , 
	\labels[7].label[76] , \labels[7].label[75] , \labels[7].label[74] , 
	\labels[7].label[73] , \labels[7].label[72] , \labels[7].label[71] , 
	\labels[7].label[70] , \labels[7].label[69] , \labels[7].label[68] , 
	\labels[7].label[67] , \labels[7].label[66] , \labels[7].label[65] , 
	\labels[7].label[64] , \labels[7].label[63] , \labels[7].label[62] , 
	\labels[7].label[61] , \labels[7].label[60] , \labels[7].label[59] , 
	\labels[7].label[58] , \labels[7].label[57] , \labels[7].label[56] , 
	\labels[7].label[55] , \labels[7].label[54] , \labels[7].label[53] , 
	\labels[7].label[52] , \labels[7].label[51] , \labels[7].label[50] , 
	\labels[7].label[49] , \labels[7].label[48] , \labels[7].label[47] , 
	\labels[7].label[46] , \labels[7].label[45] , \labels[7].label[44] , 
	\labels[7].label[43] , \labels[7].label[42] , \labels[7].label[41] , 
	\labels[7].label[40] , \labels[7].label[39] , \labels[7].label[38] , 
	\labels[7].label[37] , \labels[7].label[36] , \labels[7].label[35] , 
	\labels[7].label[34] , \labels[7].label[33] , \labels[7].label[32] , 
	\labels[7].label[31] , \labels[7].label[30] , \labels[7].label[29] , 
	\labels[7].label[28] , \labels[7].label[27] , \labels[7].label[26] , 
	\labels[7].label[25] , \labels[7].label[24] , \labels[7].label[23] , 
	\labels[7].label[22] , \labels[7].label[21] , \labels[7].label[20] , 
	\labels[7].label[19] , \labels[7].label[18] , \labels[7].label[17] , 
	\labels[7].label[16] , \labels[7].label[15] , \labels[7].label[14] , 
	\labels[7].label[13] , \labels[7].label[12] , \labels[7].label[11] , 
	\labels[7].label[10] , \labels[7].label[9] , \labels[7].label[8] , 
	\labels[7].label[7] , \labels[7].label[6] , \labels[7].label[5] , 
	\labels[7].label[4] , \labels[7].label[3] , \labels[7].label[2] , 
	\labels[7].label[1] , \labels[7].label[0] , 
	\labels[7].delimiter_valid[0] , \labels[7].delimiter[7] , 
	\labels[7].delimiter[6] , \labels[7].delimiter[5] , 
	\labels[7].delimiter[4] , \labels[7].delimiter[3] , 
	\labels[7].delimiter[2] , \labels[7].delimiter[1] , 
	\labels[7].delimiter[0] , \labels[6].guid_size[0] , 
	\labels[6].label_size[5] , \labels[6].label_size[4] , 
	\labels[6].label_size[3] , \labels[6].label_size[2] , 
	\labels[6].label_size[1] , \labels[6].label_size[0] , 
	\labels[6].label[255] , \labels[6].label[254] , 
	\labels[6].label[253] , \labels[6].label[252] , 
	\labels[6].label[251] , \labels[6].label[250] , 
	\labels[6].label[249] , \labels[6].label[248] , 
	\labels[6].label[247] , \labels[6].label[246] , 
	\labels[6].label[245] , \labels[6].label[244] , 
	\labels[6].label[243] , \labels[6].label[242] , 
	\labels[6].label[241] , \labels[6].label[240] , 
	\labels[6].label[239] , \labels[6].label[238] , 
	\labels[6].label[237] , \labels[6].label[236] , 
	\labels[6].label[235] , \labels[6].label[234] , 
	\labels[6].label[233] , \labels[6].label[232] , 
	\labels[6].label[231] , \labels[6].label[230] , 
	\labels[6].label[229] , \labels[6].label[228] , 
	\labels[6].label[227] , \labels[6].label[226] , 
	\labels[6].label[225] , \labels[6].label[224] , 
	\labels[6].label[223] , \labels[6].label[222] , 
	\labels[6].label[221] , \labels[6].label[220] , 
	\labels[6].label[219] , \labels[6].label[218] , 
	\labels[6].label[217] , \labels[6].label[216] , 
	\labels[6].label[215] , \labels[6].label[214] , 
	\labels[6].label[213] , \labels[6].label[212] , 
	\labels[6].label[211] , \labels[6].label[210] , 
	\labels[6].label[209] , \labels[6].label[208] , 
	\labels[6].label[207] , \labels[6].label[206] , 
	\labels[6].label[205] , \labels[6].label[204] , 
	\labels[6].label[203] , \labels[6].label[202] , 
	\labels[6].label[201] , \labels[6].label[200] , 
	\labels[6].label[199] , \labels[6].label[198] , 
	\labels[6].label[197] , \labels[6].label[196] , 
	\labels[6].label[195] , \labels[6].label[194] , 
	\labels[6].label[193] , \labels[6].label[192] , 
	\labels[6].label[191] , \labels[6].label[190] , 
	\labels[6].label[189] , \labels[6].label[188] , 
	\labels[6].label[187] , \labels[6].label[186] , 
	\labels[6].label[185] , \labels[6].label[184] , 
	\labels[6].label[183] , \labels[6].label[182] , 
	\labels[6].label[181] , \labels[6].label[180] , 
	\labels[6].label[179] , \labels[6].label[178] , 
	\labels[6].label[177] , \labels[6].label[176] , 
	\labels[6].label[175] , \labels[6].label[174] , 
	\labels[6].label[173] , \labels[6].label[172] , 
	\labels[6].label[171] , \labels[6].label[170] , 
	\labels[6].label[169] , \labels[6].label[168] , 
	\labels[6].label[167] , \labels[6].label[166] , 
	\labels[6].label[165] , \labels[6].label[164] , 
	\labels[6].label[163] , \labels[6].label[162] , 
	\labels[6].label[161] , \labels[6].label[160] , 
	\labels[6].label[159] , \labels[6].label[158] , 
	\labels[6].label[157] , \labels[6].label[156] , 
	\labels[6].label[155] , \labels[6].label[154] , 
	\labels[6].label[153] , \labels[6].label[152] , 
	\labels[6].label[151] , \labels[6].label[150] , 
	\labels[6].label[149] , \labels[6].label[148] , 
	\labels[6].label[147] , \labels[6].label[146] , 
	\labels[6].label[145] , \labels[6].label[144] , 
	\labels[6].label[143] , \labels[6].label[142] , 
	\labels[6].label[141] , \labels[6].label[140] , 
	\labels[6].label[139] , \labels[6].label[138] , 
	\labels[6].label[137] , \labels[6].label[136] , 
	\labels[6].label[135] , \labels[6].label[134] , 
	\labels[6].label[133] , \labels[6].label[132] , 
	\labels[6].label[131] , \labels[6].label[130] , 
	\labels[6].label[129] , \labels[6].label[128] , 
	\labels[6].label[127] , \labels[6].label[126] , 
	\labels[6].label[125] , \labels[6].label[124] , 
	\labels[6].label[123] , \labels[6].label[122] , 
	\labels[6].label[121] , \labels[6].label[120] , 
	\labels[6].label[119] , \labels[6].label[118] , 
	\labels[6].label[117] , \labels[6].label[116] , 
	\labels[6].label[115] , \labels[6].label[114] , 
	\labels[6].label[113] , \labels[6].label[112] , 
	\labels[6].label[111] , \labels[6].label[110] , 
	\labels[6].label[109] , \labels[6].label[108] , 
	\labels[6].label[107] , \labels[6].label[106] , 
	\labels[6].label[105] , \labels[6].label[104] , 
	\labels[6].label[103] , \labels[6].label[102] , 
	\labels[6].label[101] , \labels[6].label[100] , 
	\labels[6].label[99] , \labels[6].label[98] , \labels[6].label[97] , 
	\labels[6].label[96] , \labels[6].label[95] , \labels[6].label[94] , 
	\labels[6].label[93] , \labels[6].label[92] , \labels[6].label[91] , 
	\labels[6].label[90] , \labels[6].label[89] , \labels[6].label[88] , 
	\labels[6].label[87] , \labels[6].label[86] , \labels[6].label[85] , 
	\labels[6].label[84] , \labels[6].label[83] , \labels[6].label[82] , 
	\labels[6].label[81] , \labels[6].label[80] , \labels[6].label[79] , 
	\labels[6].label[78] , \labels[6].label[77] , \labels[6].label[76] , 
	\labels[6].label[75] , \labels[6].label[74] , \labels[6].label[73] , 
	\labels[6].label[72] , \labels[6].label[71] , \labels[6].label[70] , 
	\labels[6].label[69] , \labels[6].label[68] , \labels[6].label[67] , 
	\labels[6].label[66] , \labels[6].label[65] , \labels[6].label[64] , 
	\labels[6].label[63] , \labels[6].label[62] , \labels[6].label[61] , 
	\labels[6].label[60] , \labels[6].label[59] , \labels[6].label[58] , 
	\labels[6].label[57] , \labels[6].label[56] , \labels[6].label[55] , 
	\labels[6].label[54] , \labels[6].label[53] , \labels[6].label[52] , 
	\labels[6].label[51] , \labels[6].label[50] , \labels[6].label[49] , 
	\labels[6].label[48] , \labels[6].label[47] , \labels[6].label[46] , 
	\labels[6].label[45] , \labels[6].label[44] , \labels[6].label[43] , 
	\labels[6].label[42] , \labels[6].label[41] , \labels[6].label[40] , 
	\labels[6].label[39] , \labels[6].label[38] , \labels[6].label[37] , 
	\labels[6].label[36] , \labels[6].label[35] , \labels[6].label[34] , 
	\labels[6].label[33] , \labels[6].label[32] , \labels[6].label[31] , 
	\labels[6].label[30] , \labels[6].label[29] , \labels[6].label[28] , 
	\labels[6].label[27] , \labels[6].label[26] , \labels[6].label[25] , 
	\labels[6].label[24] , \labels[6].label[23] , \labels[6].label[22] , 
	\labels[6].label[21] , \labels[6].label[20] , \labels[6].label[19] , 
	\labels[6].label[18] , \labels[6].label[17] , \labels[6].label[16] , 
	\labels[6].label[15] , \labels[6].label[14] , \labels[6].label[13] , 
	\labels[6].label[12] , \labels[6].label[11] , \labels[6].label[10] , 
	\labels[6].label[9] , \labels[6].label[8] , \labels[6].label[7] , 
	\labels[6].label[6] , \labels[6].label[5] , \labels[6].label[4] , 
	\labels[6].label[3] , \labels[6].label[2] , \labels[6].label[1] , 
	\labels[6].label[0] , \labels[6].delimiter_valid[0] , 
	\labels[6].delimiter[7] , \labels[6].delimiter[6] , 
	\labels[6].delimiter[5] , \labels[6].delimiter[4] , 
	\labels[6].delimiter[3] , \labels[6].delimiter[2] , 
	\labels[6].delimiter[1] , \labels[6].delimiter[0] , 
	\labels[5].guid_size[0] , \labels[5].label_size[5] , 
	\labels[5].label_size[4] , \labels[5].label_size[3] , 
	\labels[5].label_size[2] , \labels[5].label_size[1] , 
	\labels[5].label_size[0] , \labels[5].label[255] , 
	\labels[5].label[254] , \labels[5].label[253] , 
	\labels[5].label[252] , \labels[5].label[251] , 
	\labels[5].label[250] , \labels[5].label[249] , 
	\labels[5].label[248] , \labels[5].label[247] , 
	\labels[5].label[246] , \labels[5].label[245] , 
	\labels[5].label[244] , \labels[5].label[243] , 
	\labels[5].label[242] , \labels[5].label[241] , 
	\labels[5].label[240] , \labels[5].label[239] , 
	\labels[5].label[238] , \labels[5].label[237] , 
	\labels[5].label[236] , \labels[5].label[235] , 
	\labels[5].label[234] , \labels[5].label[233] , 
	\labels[5].label[232] , \labels[5].label[231] , 
	\labels[5].label[230] , \labels[5].label[229] , 
	\labels[5].label[228] , \labels[5].label[227] , 
	\labels[5].label[226] , \labels[5].label[225] , 
	\labels[5].label[224] , \labels[5].label[223] , 
	\labels[5].label[222] , \labels[5].label[221] , 
	\labels[5].label[220] , \labels[5].label[219] , 
	\labels[5].label[218] , \labels[5].label[217] , 
	\labels[5].label[216] , \labels[5].label[215] , 
	\labels[5].label[214] , \labels[5].label[213] , 
	\labels[5].label[212] , \labels[5].label[211] , 
	\labels[5].label[210] , \labels[5].label[209] , 
	\labels[5].label[208] , \labels[5].label[207] , 
	\labels[5].label[206] , \labels[5].label[205] , 
	\labels[5].label[204] , \labels[5].label[203] , 
	\labels[5].label[202] , \labels[5].label[201] , 
	\labels[5].label[200] , \labels[5].label[199] , 
	\labels[5].label[198] , \labels[5].label[197] , 
	\labels[5].label[196] , \labels[5].label[195] , 
	\labels[5].label[194] , \labels[5].label[193] , 
	\labels[5].label[192] , \labels[5].label[191] , 
	\labels[5].label[190] , \labels[5].label[189] , 
	\labels[5].label[188] , \labels[5].label[187] , 
	\labels[5].label[186] , \labels[5].label[185] , 
	\labels[5].label[184] , \labels[5].label[183] , 
	\labels[5].label[182] , \labels[5].label[181] , 
	\labels[5].label[180] , \labels[5].label[179] , 
	\labels[5].label[178] , \labels[5].label[177] , 
	\labels[5].label[176] , \labels[5].label[175] , 
	\labels[5].label[174] , \labels[5].label[173] , 
	\labels[5].label[172] , \labels[5].label[171] , 
	\labels[5].label[170] , \labels[5].label[169] , 
	\labels[5].label[168] , \labels[5].label[167] , 
	\labels[5].label[166] , \labels[5].label[165] , 
	\labels[5].label[164] , \labels[5].label[163] , 
	\labels[5].label[162] , \labels[5].label[161] , 
	\labels[5].label[160] , \labels[5].label[159] , 
	\labels[5].label[158] , \labels[5].label[157] , 
	\labels[5].label[156] , \labels[5].label[155] , 
	\labels[5].label[154] , \labels[5].label[153] , 
	\labels[5].label[152] , \labels[5].label[151] , 
	\labels[5].label[150] , \labels[5].label[149] , 
	\labels[5].label[148] , \labels[5].label[147] , 
	\labels[5].label[146] , \labels[5].label[145] , 
	\labels[5].label[144] , \labels[5].label[143] , 
	\labels[5].label[142] , \labels[5].label[141] , 
	\labels[5].label[140] , \labels[5].label[139] , 
	\labels[5].label[138] , \labels[5].label[137] , 
	\labels[5].label[136] , \labels[5].label[135] , 
	\labels[5].label[134] , \labels[5].label[133] , 
	\labels[5].label[132] , \labels[5].label[131] , 
	\labels[5].label[130] , \labels[5].label[129] , 
	\labels[5].label[128] , \labels[5].label[127] , 
	\labels[5].label[126] , \labels[5].label[125] , 
	\labels[5].label[124] , \labels[5].label[123] , 
	\labels[5].label[122] , \labels[5].label[121] , 
	\labels[5].label[120] , \labels[5].label[119] , 
	\labels[5].label[118] , \labels[5].label[117] , 
	\labels[5].label[116] , \labels[5].label[115] , 
	\labels[5].label[114] , \labels[5].label[113] , 
	\labels[5].label[112] , \labels[5].label[111] , 
	\labels[5].label[110] , \labels[5].label[109] , 
	\labels[5].label[108] , \labels[5].label[107] , 
	\labels[5].label[106] , \labels[5].label[105] , 
	\labels[5].label[104] , \labels[5].label[103] , 
	\labels[5].label[102] , \labels[5].label[101] , 
	\labels[5].label[100] , \labels[5].label[99] , \labels[5].label[98] , 
	\labels[5].label[97] , \labels[5].label[96] , \labels[5].label[95] , 
	\labels[5].label[94] , \labels[5].label[93] , \labels[5].label[92] , 
	\labels[5].label[91] , \labels[5].label[90] , \labels[5].label[89] , 
	\labels[5].label[88] , \labels[5].label[87] , \labels[5].label[86] , 
	\labels[5].label[85] , \labels[5].label[84] , \labels[5].label[83] , 
	\labels[5].label[82] , \labels[5].label[81] , \labels[5].label[80] , 
	\labels[5].label[79] , \labels[5].label[78] , \labels[5].label[77] , 
	\labels[5].label[76] , \labels[5].label[75] , \labels[5].label[74] , 
	\labels[5].label[73] , \labels[5].label[72] , \labels[5].label[71] , 
	\labels[5].label[70] , \labels[5].label[69] , \labels[5].label[68] , 
	\labels[5].label[67] , \labels[5].label[66] , \labels[5].label[65] , 
	\labels[5].label[64] , \labels[5].label[63] , \labels[5].label[62] , 
	\labels[5].label[61] , \labels[5].label[60] , \labels[5].label[59] , 
	\labels[5].label[58] , \labels[5].label[57] , \labels[5].label[56] , 
	\labels[5].label[55] , \labels[5].label[54] , \labels[5].label[53] , 
	\labels[5].label[52] , \labels[5].label[51] , \labels[5].label[50] , 
	\labels[5].label[49] , \labels[5].label[48] , \labels[5].label[47] , 
	\labels[5].label[46] , \labels[5].label[45] , \labels[5].label[44] , 
	\labels[5].label[43] , \labels[5].label[42] , \labels[5].label[41] , 
	\labels[5].label[40] , \labels[5].label[39] , \labels[5].label[38] , 
	\labels[5].label[37] , \labels[5].label[36] , \labels[5].label[35] , 
	\labels[5].label[34] , \labels[5].label[33] , \labels[5].label[32] , 
	\labels[5].label[31] , \labels[5].label[30] , \labels[5].label[29] , 
	\labels[5].label[28] , \labels[5].label[27] , \labels[5].label[26] , 
	\labels[5].label[25] , \labels[5].label[24] , \labels[5].label[23] , 
	\labels[5].label[22] , \labels[5].label[21] , \labels[5].label[20] , 
	\labels[5].label[19] , \labels[5].label[18] , \labels[5].label[17] , 
	\labels[5].label[16] , \labels[5].label[15] , \labels[5].label[14] , 
	\labels[5].label[13] , \labels[5].label[12] , \labels[5].label[11] , 
	\labels[5].label[10] , \labels[5].label[9] , \labels[5].label[8] , 
	\labels[5].label[7] , \labels[5].label[6] , \labels[5].label[5] , 
	\labels[5].label[4] , \labels[5].label[3] , \labels[5].label[2] , 
	\labels[5].label[1] , \labels[5].label[0] , 
	\labels[5].delimiter_valid[0] , \labels[5].delimiter[7] , 
	\labels[5].delimiter[6] , \labels[5].delimiter[5] , 
	\labels[5].delimiter[4] , \labels[5].delimiter[3] , 
	\labels[5].delimiter[2] , \labels[5].delimiter[1] , 
	\labels[5].delimiter[0] , \labels[4].guid_size[0] , 
	\labels[4].label_size[5] , \labels[4].label_size[4] , 
	\labels[4].label_size[3] , \labels[4].label_size[2] , 
	\labels[4].label_size[1] , \labels[4].label_size[0] , 
	\labels[4].label[255] , \labels[4].label[254] , 
	\labels[4].label[253] , \labels[4].label[252] , 
	\labels[4].label[251] , \labels[4].label[250] , 
	\labels[4].label[249] , \labels[4].label[248] , 
	\labels[4].label[247] , \labels[4].label[246] , 
	\labels[4].label[245] , \labels[4].label[244] , 
	\labels[4].label[243] , \labels[4].label[242] , 
	\labels[4].label[241] , \labels[4].label[240] , 
	\labels[4].label[239] , \labels[4].label[238] , 
	\labels[4].label[237] , \labels[4].label[236] , 
	\labels[4].label[235] , \labels[4].label[234] , 
	\labels[4].label[233] , \labels[4].label[232] , 
	\labels[4].label[231] , \labels[4].label[230] , 
	\labels[4].label[229] , \labels[4].label[228] , 
	\labels[4].label[227] , \labels[4].label[226] , 
	\labels[4].label[225] , \labels[4].label[224] , 
	\labels[4].label[223] , \labels[4].label[222] , 
	\labels[4].label[221] , \labels[4].label[220] , 
	\labels[4].label[219] , \labels[4].label[218] , 
	\labels[4].label[217] , \labels[4].label[216] , 
	\labels[4].label[215] , \labels[4].label[214] , 
	\labels[4].label[213] , \labels[4].label[212] , 
	\labels[4].label[211] , \labels[4].label[210] , 
	\labels[4].label[209] , \labels[4].label[208] , 
	\labels[4].label[207] , \labels[4].label[206] , 
	\labels[4].label[205] , \labels[4].label[204] , 
	\labels[4].label[203] , \labels[4].label[202] , 
	\labels[4].label[201] , \labels[4].label[200] , 
	\labels[4].label[199] , \labels[4].label[198] , 
	\labels[4].label[197] , \labels[4].label[196] , 
	\labels[4].label[195] , \labels[4].label[194] , 
	\labels[4].label[193] , \labels[4].label[192] , 
	\labels[4].label[191] , \labels[4].label[190] , 
	\labels[4].label[189] , \labels[4].label[188] , 
	\labels[4].label[187] , \labels[4].label[186] , 
	\labels[4].label[185] , \labels[4].label[184] , 
	\labels[4].label[183] , \labels[4].label[182] , 
	\labels[4].label[181] , \labels[4].label[180] , 
	\labels[4].label[179] , \labels[4].label[178] , 
	\labels[4].label[177] , \labels[4].label[176] , 
	\labels[4].label[175] , \labels[4].label[174] , 
	\labels[4].label[173] , \labels[4].label[172] , 
	\labels[4].label[171] , \labels[4].label[170] , 
	\labels[4].label[169] , \labels[4].label[168] , 
	\labels[4].label[167] , \labels[4].label[166] , 
	\labels[4].label[165] , \labels[4].label[164] , 
	\labels[4].label[163] , \labels[4].label[162] , 
	\labels[4].label[161] , \labels[4].label[160] , 
	\labels[4].label[159] , \labels[4].label[158] , 
	\labels[4].label[157] , \labels[4].label[156] , 
	\labels[4].label[155] , \labels[4].label[154] , 
	\labels[4].label[153] , \labels[4].label[152] , 
	\labels[4].label[151] , \labels[4].label[150] , 
	\labels[4].label[149] , \labels[4].label[148] , 
	\labels[4].label[147] , \labels[4].label[146] , 
	\labels[4].label[145] , \labels[4].label[144] , 
	\labels[4].label[143] , \labels[4].label[142] , 
	\labels[4].label[141] , \labels[4].label[140] , 
	\labels[4].label[139] , \labels[4].label[138] , 
	\labels[4].label[137] , \labels[4].label[136] , 
	\labels[4].label[135] , \labels[4].label[134] , 
	\labels[4].label[133] , \labels[4].label[132] , 
	\labels[4].label[131] , \labels[4].label[130] , 
	\labels[4].label[129] , \labels[4].label[128] , 
	\labels[4].label[127] , \labels[4].label[126] , 
	\labels[4].label[125] , \labels[4].label[124] , 
	\labels[4].label[123] , \labels[4].label[122] , 
	\labels[4].label[121] , \labels[4].label[120] , 
	\labels[4].label[119] , \labels[4].label[118] , 
	\labels[4].label[117] , \labels[4].label[116] , 
	\labels[4].label[115] , \labels[4].label[114] , 
	\labels[4].label[113] , \labels[4].label[112] , 
	\labels[4].label[111] , \labels[4].label[110] , 
	\labels[4].label[109] , \labels[4].label[108] , 
	\labels[4].label[107] , \labels[4].label[106] , 
	\labels[4].label[105] , \labels[4].label[104] , 
	\labels[4].label[103] , \labels[4].label[102] , 
	\labels[4].label[101] , \labels[4].label[100] , 
	\labels[4].label[99] , \labels[4].label[98] , \labels[4].label[97] , 
	\labels[4].label[96] , \labels[4].label[95] , \labels[4].label[94] , 
	\labels[4].label[93] , \labels[4].label[92] , \labels[4].label[91] , 
	\labels[4].label[90] , \labels[4].label[89] , \labels[4].label[88] , 
	\labels[4].label[87] , \labels[4].label[86] , \labels[4].label[85] , 
	\labels[4].label[84] , \labels[4].label[83] , \labels[4].label[82] , 
	\labels[4].label[81] , \labels[4].label[80] , \labels[4].label[79] , 
	\labels[4].label[78] , \labels[4].label[77] , \labels[4].label[76] , 
	\labels[4].label[75] , \labels[4].label[74] , \labels[4].label[73] , 
	\labels[4].label[72] , \labels[4].label[71] , \labels[4].label[70] , 
	\labels[4].label[69] , \labels[4].label[68] , \labels[4].label[67] , 
	\labels[4].label[66] , \labels[4].label[65] , \labels[4].label[64] , 
	\labels[4].label[63] , \labels[4].label[62] , \labels[4].label[61] , 
	\labels[4].label[60] , \labels[4].label[59] , \labels[4].label[58] , 
	\labels[4].label[57] , \labels[4].label[56] , \labels[4].label[55] , 
	\labels[4].label[54] , \labels[4].label[53] , \labels[4].label[52] , 
	\labels[4].label[51] , \labels[4].label[50] , \labels[4].label[49] , 
	\labels[4].label[48] , \labels[4].label[47] , \labels[4].label[46] , 
	\labels[4].label[45] , \labels[4].label[44] , \labels[4].label[43] , 
	\labels[4].label[42] , \labels[4].label[41] , \labels[4].label[40] , 
	\labels[4].label[39] , \labels[4].label[38] , \labels[4].label[37] , 
	\labels[4].label[36] , \labels[4].label[35] , \labels[4].label[34] , 
	\labels[4].label[33] , \labels[4].label[32] , \labels[4].label[31] , 
	\labels[4].label[30] , \labels[4].label[29] , \labels[4].label[28] , 
	\labels[4].label[27] , \labels[4].label[26] , \labels[4].label[25] , 
	\labels[4].label[24] , \labels[4].label[23] , \labels[4].label[22] , 
	\labels[4].label[21] , \labels[4].label[20] , \labels[4].label[19] , 
	\labels[4].label[18] , \labels[4].label[17] , \labels[4].label[16] , 
	\labels[4].label[15] , \labels[4].label[14] , \labels[4].label[13] , 
	\labels[4].label[12] , \labels[4].label[11] , \labels[4].label[10] , 
	\labels[4].label[9] , \labels[4].label[8] , \labels[4].label[7] , 
	\labels[4].label[6] , \labels[4].label[5] , \labels[4].label[4] , 
	\labels[4].label[3] , \labels[4].label[2] , \labels[4].label[1] , 
	\labels[4].label[0] , \labels[4].delimiter_valid[0] , 
	\labels[4].delimiter[7] , \labels[4].delimiter[6] , 
	\labels[4].delimiter[5] , \labels[4].delimiter[4] , 
	\labels[4].delimiter[3] , \labels[4].delimiter[2] , 
	\labels[4].delimiter[1] , \labels[4].delimiter[0] , 
	\labels[3].guid_size[0] , \labels[3].label_size[5] , 
	\labels[3].label_size[4] , \labels[3].label_size[3] , 
	\labels[3].label_size[2] , \labels[3].label_size[1] , 
	\labels[3].label_size[0] , \labels[3].label[255] , 
	\labels[3].label[254] , \labels[3].label[253] , 
	\labels[3].label[252] , \labels[3].label[251] , 
	\labels[3].label[250] , \labels[3].label[249] , 
	\labels[3].label[248] , \labels[3].label[247] , 
	\labels[3].label[246] , \labels[3].label[245] , 
	\labels[3].label[244] , \labels[3].label[243] , 
	\labels[3].label[242] , \labels[3].label[241] , 
	\labels[3].label[240] , \labels[3].label[239] , 
	\labels[3].label[238] , \labels[3].label[237] , 
	\labels[3].label[236] , \labels[3].label[235] , 
	\labels[3].label[234] , \labels[3].label[233] , 
	\labels[3].label[232] , \labels[3].label[231] , 
	\labels[3].label[230] , \labels[3].label[229] , 
	\labels[3].label[228] , \labels[3].label[227] , 
	\labels[3].label[226] , \labels[3].label[225] , 
	\labels[3].label[224] , \labels[3].label[223] , 
	\labels[3].label[222] , \labels[3].label[221] , 
	\labels[3].label[220] , \labels[3].label[219] , 
	\labels[3].label[218] , \labels[3].label[217] , 
	\labels[3].label[216] , \labels[3].label[215] , 
	\labels[3].label[214] , \labels[3].label[213] , 
	\labels[3].label[212] , \labels[3].label[211] , 
	\labels[3].label[210] , \labels[3].label[209] , 
	\labels[3].label[208] , \labels[3].label[207] , 
	\labels[3].label[206] , \labels[3].label[205] , 
	\labels[3].label[204] , \labels[3].label[203] , 
	\labels[3].label[202] , \labels[3].label[201] , 
	\labels[3].label[200] , \labels[3].label[199] , 
	\labels[3].label[198] , \labels[3].label[197] , 
	\labels[3].label[196] , \labels[3].label[195] , 
	\labels[3].label[194] , \labels[3].label[193] , 
	\labels[3].label[192] , \labels[3].label[191] , 
	\labels[3].label[190] , \labels[3].label[189] , 
	\labels[3].label[188] , \labels[3].label[187] , 
	\labels[3].label[186] , \labels[3].label[185] , 
	\labels[3].label[184] , \labels[3].label[183] , 
	\labels[3].label[182] , \labels[3].label[181] , 
	\labels[3].label[180] , \labels[3].label[179] , 
	\labels[3].label[178] , \labels[3].label[177] , 
	\labels[3].label[176] , \labels[3].label[175] , 
	\labels[3].label[174] , \labels[3].label[173] , 
	\labels[3].label[172] , \labels[3].label[171] , 
	\labels[3].label[170] , \labels[3].label[169] , 
	\labels[3].label[168] , \labels[3].label[167] , 
	\labels[3].label[166] , \labels[3].label[165] , 
	\labels[3].label[164] , \labels[3].label[163] , 
	\labels[3].label[162] , \labels[3].label[161] , 
	\labels[3].label[160] , \labels[3].label[159] , 
	\labels[3].label[158] , \labels[3].label[157] , 
	\labels[3].label[156] , \labels[3].label[155] , 
	\labels[3].label[154] , \labels[3].label[153] , 
	\labels[3].label[152] , \labels[3].label[151] , 
	\labels[3].label[150] , \labels[3].label[149] , 
	\labels[3].label[148] , \labels[3].label[147] , 
	\labels[3].label[146] , \labels[3].label[145] , 
	\labels[3].label[144] , \labels[3].label[143] , 
	\labels[3].label[142] , \labels[3].label[141] , 
	\labels[3].label[140] , \labels[3].label[139] , 
	\labels[3].label[138] , \labels[3].label[137] , 
	\labels[3].label[136] , \labels[3].label[135] , 
	\labels[3].label[134] , \labels[3].label[133] , 
	\labels[3].label[132] , \labels[3].label[131] , 
	\labels[3].label[130] , \labels[3].label[129] , 
	\labels[3].label[128] , \labels[3].label[127] , 
	\labels[3].label[126] , \labels[3].label[125] , 
	\labels[3].label[124] , \labels[3].label[123] , 
	\labels[3].label[122] , \labels[3].label[121] , 
	\labels[3].label[120] , \labels[3].label[119] , 
	\labels[3].label[118] , \labels[3].label[117] , 
	\labels[3].label[116] , \labels[3].label[115] , 
	\labels[3].label[114] , \labels[3].label[113] , 
	\labels[3].label[112] , \labels[3].label[111] , 
	\labels[3].label[110] , \labels[3].label[109] , 
	\labels[3].label[108] , \labels[3].label[107] , 
	\labels[3].label[106] , \labels[3].label[105] , 
	\labels[3].label[104] , \labels[3].label[103] , 
	\labels[3].label[102] , \labels[3].label[101] , 
	\labels[3].label[100] , \labels[3].label[99] , \labels[3].label[98] , 
	\labels[3].label[97] , \labels[3].label[96] , \labels[3].label[95] , 
	\labels[3].label[94] , \labels[3].label[93] , \labels[3].label[92] , 
	\labels[3].label[91] , \labels[3].label[90] , \labels[3].label[89] , 
	\labels[3].label[88] , \labels[3].label[87] , \labels[3].label[86] , 
	\labels[3].label[85] , \labels[3].label[84] , \labels[3].label[83] , 
	\labels[3].label[82] , \labels[3].label[81] , \labels[3].label[80] , 
	\labels[3].label[79] , \labels[3].label[78] , \labels[3].label[77] , 
	\labels[3].label[76] , \labels[3].label[75] , \labels[3].label[74] , 
	\labels[3].label[73] , \labels[3].label[72] , \labels[3].label[71] , 
	\labels[3].label[70] , \labels[3].label[69] , \labels[3].label[68] , 
	\labels[3].label[67] , \labels[3].label[66] , \labels[3].label[65] , 
	\labels[3].label[64] , \labels[3].label[63] , \labels[3].label[62] , 
	\labels[3].label[61] , \labels[3].label[60] , \labels[3].label[59] , 
	\labels[3].label[58] , \labels[3].label[57] , \labels[3].label[56] , 
	\labels[3].label[55] , \labels[3].label[54] , \labels[3].label[53] , 
	\labels[3].label[52] , \labels[3].label[51] , \labels[3].label[50] , 
	\labels[3].label[49] , \labels[3].label[48] , \labels[3].label[47] , 
	\labels[3].label[46] , \labels[3].label[45] , \labels[3].label[44] , 
	\labels[3].label[43] , \labels[3].label[42] , \labels[3].label[41] , 
	\labels[3].label[40] , \labels[3].label[39] , \labels[3].label[38] , 
	\labels[3].label[37] , \labels[3].label[36] , \labels[3].label[35] , 
	\labels[3].label[34] , \labels[3].label[33] , \labels[3].label[32] , 
	\labels[3].label[31] , \labels[3].label[30] , \labels[3].label[29] , 
	\labels[3].label[28] , \labels[3].label[27] , \labels[3].label[26] , 
	\labels[3].label[25] , \labels[3].label[24] , \labels[3].label[23] , 
	\labels[3].label[22] , \labels[3].label[21] , \labels[3].label[20] , 
	\labels[3].label[19] , \labels[3].label[18] , \labels[3].label[17] , 
	\labels[3].label[16] , \labels[3].label[15] , \labels[3].label[14] , 
	\labels[3].label[13] , \labels[3].label[12] , \labels[3].label[11] , 
	\labels[3].label[10] , \labels[3].label[9] , \labels[3].label[8] , 
	\labels[3].label[7] , \labels[3].label[6] , \labels[3].label[5] , 
	\labels[3].label[4] , \labels[3].label[3] , \labels[3].label[2] , 
	\labels[3].label[1] , \labels[3].label[0] , 
	\labels[3].delimiter_valid[0] , \labels[3].delimiter[7] , 
	\labels[3].delimiter[6] , \labels[3].delimiter[5] , 
	\labels[3].delimiter[4] , \labels[3].delimiter[3] , 
	\labels[3].delimiter[2] , \labels[3].delimiter[1] , 
	\labels[3].delimiter[0] , \labels[2].guid_size[0] , 
	\labels[2].label_size[5] , \labels[2].label_size[4] , 
	\labels[2].label_size[3] , \labels[2].label_size[2] , 
	\labels[2].label_size[1] , \labels[2].label_size[0] , 
	\labels[2].label[255] , \labels[2].label[254] , 
	\labels[2].label[253] , \labels[2].label[252] , 
	\labels[2].label[251] , \labels[2].label[250] , 
	\labels[2].label[249] , \labels[2].label[248] , 
	\labels[2].label[247] , \labels[2].label[246] , 
	\labels[2].label[245] , \labels[2].label[244] , 
	\labels[2].label[243] , \labels[2].label[242] , 
	\labels[2].label[241] , \labels[2].label[240] , 
	\labels[2].label[239] , \labels[2].label[238] , 
	\labels[2].label[237] , \labels[2].label[236] , 
	\labels[2].label[235] , \labels[2].label[234] , 
	\labels[2].label[233] , \labels[2].label[232] , 
	\labels[2].label[231] , \labels[2].label[230] , 
	\labels[2].label[229] , \labels[2].label[228] , 
	\labels[2].label[227] , \labels[2].label[226] , 
	\labels[2].label[225] , \labels[2].label[224] , 
	\labels[2].label[223] , \labels[2].label[222] , 
	\labels[2].label[221] , \labels[2].label[220] , 
	\labels[2].label[219] , \labels[2].label[218] , 
	\labels[2].label[217] , \labels[2].label[216] , 
	\labels[2].label[215] , \labels[2].label[214] , 
	\labels[2].label[213] , \labels[2].label[212] , 
	\labels[2].label[211] , \labels[2].label[210] , 
	\labels[2].label[209] , \labels[2].label[208] , 
	\labels[2].label[207] , \labels[2].label[206] , 
	\labels[2].label[205] , \labels[2].label[204] , 
	\labels[2].label[203] , \labels[2].label[202] , 
	\labels[2].label[201] , \labels[2].label[200] , 
	\labels[2].label[199] , \labels[2].label[198] , 
	\labels[2].label[197] , \labels[2].label[196] , 
	\labels[2].label[195] , \labels[2].label[194] , 
	\labels[2].label[193] , \labels[2].label[192] , 
	\labels[2].label[191] , \labels[2].label[190] , 
	\labels[2].label[189] , \labels[2].label[188] , 
	\labels[2].label[187] , \labels[2].label[186] , 
	\labels[2].label[185] , \labels[2].label[184] , 
	\labels[2].label[183] , \labels[2].label[182] , 
	\labels[2].label[181] , \labels[2].label[180] , 
	\labels[2].label[179] , \labels[2].label[178] , 
	\labels[2].label[177] , \labels[2].label[176] , 
	\labels[2].label[175] , \labels[2].label[174] , 
	\labels[2].label[173] , \labels[2].label[172] , 
	\labels[2].label[171] , \labels[2].label[170] , 
	\labels[2].label[169] , \labels[2].label[168] , 
	\labels[2].label[167] , \labels[2].label[166] , 
	\labels[2].label[165] , \labels[2].label[164] , 
	\labels[2].label[163] , \labels[2].label[162] , 
	\labels[2].label[161] , \labels[2].label[160] , 
	\labels[2].label[159] , \labels[2].label[158] , 
	\labels[2].label[157] , \labels[2].label[156] , 
	\labels[2].label[155] , \labels[2].label[154] , 
	\labels[2].label[153] , \labels[2].label[152] , 
	\labels[2].label[151] , \labels[2].label[150] , 
	\labels[2].label[149] , \labels[2].label[148] , 
	\labels[2].label[147] , \labels[2].label[146] , 
	\labels[2].label[145] , \labels[2].label[144] , 
	\labels[2].label[143] , \labels[2].label[142] , 
	\labels[2].label[141] , \labels[2].label[140] , 
	\labels[2].label[139] , \labels[2].label[138] , 
	\labels[2].label[137] , \labels[2].label[136] , 
	\labels[2].label[135] , \labels[2].label[134] , 
	\labels[2].label[133] , \labels[2].label[132] , 
	\labels[2].label[131] , \labels[2].label[130] , 
	\labels[2].label[129] , \labels[2].label[128] , 
	\labels[2].label[127] , \labels[2].label[126] , 
	\labels[2].label[125] , \labels[2].label[124] , 
	\labels[2].label[123] , \labels[2].label[122] , 
	\labels[2].label[121] , \labels[2].label[120] , 
	\labels[2].label[119] , \labels[2].label[118] , 
	\labels[2].label[117] , \labels[2].label[116] , 
	\labels[2].label[115] , \labels[2].label[114] , 
	\labels[2].label[113] , \labels[2].label[112] , 
	\labels[2].label[111] , \labels[2].label[110] , 
	\labels[2].label[109] , \labels[2].label[108] , 
	\labels[2].label[107] , \labels[2].label[106] , 
	\labels[2].label[105] , \labels[2].label[104] , 
	\labels[2].label[103] , \labels[2].label[102] , 
	\labels[2].label[101] , \labels[2].label[100] , 
	\labels[2].label[99] , \labels[2].label[98] , \labels[2].label[97] , 
	\labels[2].label[96] , \labels[2].label[95] , \labels[2].label[94] , 
	\labels[2].label[93] , \labels[2].label[92] , \labels[2].label[91] , 
	\labels[2].label[90] , \labels[2].label[89] , \labels[2].label[88] , 
	\labels[2].label[87] , \labels[2].label[86] , \labels[2].label[85] , 
	\labels[2].label[84] , \labels[2].label[83] , \labels[2].label[82] , 
	\labels[2].label[81] , \labels[2].label[80] , \labels[2].label[79] , 
	\labels[2].label[78] , \labels[2].label[77] , \labels[2].label[76] , 
	\labels[2].label[75] , \labels[2].label[74] , \labels[2].label[73] , 
	\labels[2].label[72] , \labels[2].label[71] , \labels[2].label[70] , 
	\labels[2].label[69] , \labels[2].label[68] , \labels[2].label[67] , 
	\labels[2].label[66] , \labels[2].label[65] , \labels[2].label[64] , 
	\labels[2].label[63] , \labels[2].label[62] , \labels[2].label[61] , 
	\labels[2].label[60] , \labels[2].label[59] , \labels[2].label[58] , 
	\labels[2].label[57] , \labels[2].label[56] , \labels[2].label[55] , 
	\labels[2].label[54] , \labels[2].label[53] , \labels[2].label[52] , 
	\labels[2].label[51] , \labels[2].label[50] , \labels[2].label[49] , 
	\labels[2].label[48] , \labels[2].label[47] , \labels[2].label[46] , 
	\labels[2].label[45] , \labels[2].label[44] , \labels[2].label[43] , 
	\labels[2].label[42] , \labels[2].label[41] , \labels[2].label[40] , 
	\labels[2].label[39] , \labels[2].label[38] , \labels[2].label[37] , 
	\labels[2].label[36] , \labels[2].label[35] , \labels[2].label[34] , 
	\labels[2].label[33] , \labels[2].label[32] , \labels[2].label[31] , 
	\labels[2].label[30] , \labels[2].label[29] , \labels[2].label[28] , 
	\labels[2].label[27] , \labels[2].label[26] , \labels[2].label[25] , 
	\labels[2].label[24] , \labels[2].label[23] , \labels[2].label[22] , 
	\labels[2].label[21] , \labels[2].label[20] , \labels[2].label[19] , 
	\labels[2].label[18] , \labels[2].label[17] , \labels[2].label[16] , 
	\labels[2].label[15] , \labels[2].label[14] , \labels[2].label[13] , 
	\labels[2].label[12] , \labels[2].label[11] , \labels[2].label[10] , 
	\labels[2].label[9] , \labels[2].label[8] , \labels[2].label[7] , 
	\labels[2].label[6] , \labels[2].label[5] , \labels[2].label[4] , 
	\labels[2].label[3] , \labels[2].label[2] , \labels[2].label[1] , 
	\labels[2].label[0] , \labels[2].delimiter_valid[0] , 
	\labels[2].delimiter[7] , \labels[2].delimiter[6] , 
	\labels[2].delimiter[5] , \labels[2].delimiter[4] , 
	\labels[2].delimiter[3] , \labels[2].delimiter[2] , 
	\labels[2].delimiter[1] , \labels[2].delimiter[0] , 
	\labels[1].guid_size[0] , \labels[1].label_size[5] , 
	\labels[1].label_size[4] , \labels[1].label_size[3] , 
	\labels[1].label_size[2] , \labels[1].label_size[1] , 
	\labels[1].label_size[0] , \labels[1].label[255] , 
	\labels[1].label[254] , \labels[1].label[253] , 
	\labels[1].label[252] , \labels[1].label[251] , 
	\labels[1].label[250] , \labels[1].label[249] , 
	\labels[1].label[248] , \labels[1].label[247] , 
	\labels[1].label[246] , \labels[1].label[245] , 
	\labels[1].label[244] , \labels[1].label[243] , 
	\labels[1].label[242] , \labels[1].label[241] , 
	\labels[1].label[240] , \labels[1].label[239] , 
	\labels[1].label[238] , \labels[1].label[237] , 
	\labels[1].label[236] , \labels[1].label[235] , 
	\labels[1].label[234] , \labels[1].label[233] , 
	\labels[1].label[232] , \labels[1].label[231] , 
	\labels[1].label[230] , \labels[1].label[229] , 
	\labels[1].label[228] , \labels[1].label[227] , 
	\labels[1].label[226] , \labels[1].label[225] , 
	\labels[1].label[224] , \labels[1].label[223] , 
	\labels[1].label[222] , \labels[1].label[221] , 
	\labels[1].label[220] , \labels[1].label[219] , 
	\labels[1].label[218] , \labels[1].label[217] , 
	\labels[1].label[216] , \labels[1].label[215] , 
	\labels[1].label[214] , \labels[1].label[213] , 
	\labels[1].label[212] , \labels[1].label[211] , 
	\labels[1].label[210] , \labels[1].label[209] , 
	\labels[1].label[208] , \labels[1].label[207] , 
	\labels[1].label[206] , \labels[1].label[205] , 
	\labels[1].label[204] , \labels[1].label[203] , 
	\labels[1].label[202] , \labels[1].label[201] , 
	\labels[1].label[200] , \labels[1].label[199] , 
	\labels[1].label[198] , \labels[1].label[197] , 
	\labels[1].label[196] , \labels[1].label[195] , 
	\labels[1].label[194] , \labels[1].label[193] , 
	\labels[1].label[192] , \labels[1].label[191] , 
	\labels[1].label[190] , \labels[1].label[189] , 
	\labels[1].label[188] , \labels[1].label[187] , 
	\labels[1].label[186] , \labels[1].label[185] , 
	\labels[1].label[184] , \labels[1].label[183] , 
	\labels[1].label[182] , \labels[1].label[181] , 
	\labels[1].label[180] , \labels[1].label[179] , 
	\labels[1].label[178] , \labels[1].label[177] , 
	\labels[1].label[176] , \labels[1].label[175] , 
	\labels[1].label[174] , \labels[1].label[173] , 
	\labels[1].label[172] , \labels[1].label[171] , 
	\labels[1].label[170] , \labels[1].label[169] , 
	\labels[1].label[168] , \labels[1].label[167] , 
	\labels[1].label[166] , \labels[1].label[165] , 
	\labels[1].label[164] , \labels[1].label[163] , 
	\labels[1].label[162] , \labels[1].label[161] , 
	\labels[1].label[160] , \labels[1].label[159] , 
	\labels[1].label[158] , \labels[1].label[157] , 
	\labels[1].label[156] , \labels[1].label[155] , 
	\labels[1].label[154] , \labels[1].label[153] , 
	\labels[1].label[152] , \labels[1].label[151] , 
	\labels[1].label[150] , \labels[1].label[149] , 
	\labels[1].label[148] , \labels[1].label[147] , 
	\labels[1].label[146] , \labels[1].label[145] , 
	\labels[1].label[144] , \labels[1].label[143] , 
	\labels[1].label[142] , \labels[1].label[141] , 
	\labels[1].label[140] , \labels[1].label[139] , 
	\labels[1].label[138] , \labels[1].label[137] , 
	\labels[1].label[136] , \labels[1].label[135] , 
	\labels[1].label[134] , \labels[1].label[133] , 
	\labels[1].label[132] , \labels[1].label[131] , 
	\labels[1].label[130] , \labels[1].label[129] , 
	\labels[1].label[128] , \labels[1].label[127] , 
	\labels[1].label[126] , \labels[1].label[125] , 
	\labels[1].label[124] , \labels[1].label[123] , 
	\labels[1].label[122] , \labels[1].label[121] , 
	\labels[1].label[120] , \labels[1].label[119] , 
	\labels[1].label[118] , \labels[1].label[117] , 
	\labels[1].label[116] , \labels[1].label[115] , 
	\labels[1].label[114] , \labels[1].label[113] , 
	\labels[1].label[112] , \labels[1].label[111] , 
	\labels[1].label[110] , \labels[1].label[109] , 
	\labels[1].label[108] , \labels[1].label[107] , 
	\labels[1].label[106] , \labels[1].label[105] , 
	\labels[1].label[104] , \labels[1].label[103] , 
	\labels[1].label[102] , \labels[1].label[101] , 
	\labels[1].label[100] , \labels[1].label[99] , \labels[1].label[98] , 
	\labels[1].label[97] , \labels[1].label[96] , \labels[1].label[95] , 
	\labels[1].label[94] , \labels[1].label[93] , \labels[1].label[92] , 
	\labels[1].label[91] , \labels[1].label[90] , \labels[1].label[89] , 
	\labels[1].label[88] , \labels[1].label[87] , \labels[1].label[86] , 
	\labels[1].label[85] , \labels[1].label[84] , \labels[1].label[83] , 
	\labels[1].label[82] , \labels[1].label[81] , \labels[1].label[80] , 
	\labels[1].label[79] , \labels[1].label[78] , \labels[1].label[77] , 
	\labels[1].label[76] , \labels[1].label[75] , \labels[1].label[74] , 
	\labels[1].label[73] , \labels[1].label[72] , \labels[1].label[71] , 
	\labels[1].label[70] , \labels[1].label[69] , \labels[1].label[68] , 
	\labels[1].label[67] , \labels[1].label[66] , \labels[1].label[65] , 
	\labels[1].label[64] , \labels[1].label[63] , \labels[1].label[62] , 
	\labels[1].label[61] , \labels[1].label[60] , \labels[1].label[59] , 
	\labels[1].label[58] , \labels[1].label[57] , \labels[1].label[56] , 
	\labels[1].label[55] , \labels[1].label[54] , \labels[1].label[53] , 
	\labels[1].label[52] , \labels[1].label[51] , \labels[1].label[50] , 
	\labels[1].label[49] , \labels[1].label[48] , \labels[1].label[47] , 
	\labels[1].label[46] , \labels[1].label[45] , \labels[1].label[44] , 
	\labels[1].label[43] , \labels[1].label[42] , \labels[1].label[41] , 
	\labels[1].label[40] , \labels[1].label[39] , \labels[1].label[38] , 
	\labels[1].label[37] , \labels[1].label[36] , \labels[1].label[35] , 
	\labels[1].label[34] , \labels[1].label[33] , \labels[1].label[32] , 
	\labels[1].label[31] , \labels[1].label[30] , \labels[1].label[29] , 
	\labels[1].label[28] , \labels[1].label[27] , \labels[1].label[26] , 
	\labels[1].label[25] , \labels[1].label[24] , \labels[1].label[23] , 
	\labels[1].label[22] , \labels[1].label[21] , \labels[1].label[20] , 
	\labels[1].label[19] , \labels[1].label[18] , \labels[1].label[17] , 
	\labels[1].label[16] , \labels[1].label[15] , \labels[1].label[14] , 
	\labels[1].label[13] , \labels[1].label[12] , \labels[1].label[11] , 
	\labels[1].label[10] , \labels[1].label[9] , \labels[1].label[8] , 
	\labels[1].label[7] , \labels[1].label[6] , \labels[1].label[5] , 
	\labels[1].label[4] , \labels[1].label[3] , \labels[1].label[2] , 
	\labels[1].label[1] , \labels[1].label[0] , 
	\labels[1].delimiter_valid[0] , \labels[1].delimiter[7] , 
	\labels[1].delimiter[6] , \labels[1].delimiter[5] , 
	\labels[1].delimiter[4] , \labels[1].delimiter[3] , 
	\labels[1].delimiter[2] , \labels[1].delimiter[1] , 
	\labels[1].delimiter[0] , \labels[0].guid_size[0] , 
	\labels[0].label_size[5] , \labels[0].label_size[4] , 
	\labels[0].label_size[3] , \labels[0].label_size[2] , 
	\labels[0].label_size[1] , \labels[0].label_size[0] , 
	\labels[0].label[255] , \labels[0].label[254] , 
	\labels[0].label[253] , \labels[0].label[252] , 
	\labels[0].label[251] , \labels[0].label[250] , 
	\labels[0].label[249] , \labels[0].label[248] , 
	\labels[0].label[247] , \labels[0].label[246] , 
	\labels[0].label[245] , \labels[0].label[244] , 
	\labels[0].label[243] , \labels[0].label[242] , 
	\labels[0].label[241] , \labels[0].label[240] , 
	\labels[0].label[239] , \labels[0].label[238] , 
	\labels[0].label[237] , \labels[0].label[236] , 
	\labels[0].label[235] , \labels[0].label[234] , 
	\labels[0].label[233] , \labels[0].label[232] , 
	\labels[0].label[231] , \labels[0].label[230] , 
	\labels[0].label[229] , \labels[0].label[228] , 
	\labels[0].label[227] , \labels[0].label[226] , 
	\labels[0].label[225] , \labels[0].label[224] , 
	\labels[0].label[223] , \labels[0].label[222] , 
	\labels[0].label[221] , \labels[0].label[220] , 
	\labels[0].label[219] , \labels[0].label[218] , 
	\labels[0].label[217] , \labels[0].label[216] , 
	\labels[0].label[215] , \labels[0].label[214] , 
	\labels[0].label[213] , \labels[0].label[212] , 
	\labels[0].label[211] , \labels[0].label[210] , 
	\labels[0].label[209] , \labels[0].label[208] , 
	\labels[0].label[207] , \labels[0].label[206] , 
	\labels[0].label[205] , \labels[0].label[204] , 
	\labels[0].label[203] , \labels[0].label[202] , 
	\labels[0].label[201] , \labels[0].label[200] , 
	\labels[0].label[199] , \labels[0].label[198] , 
	\labels[0].label[197] , \labels[0].label[196] , 
	\labels[0].label[195] , \labels[0].label[194] , 
	\labels[0].label[193] , \labels[0].label[192] , 
	\labels[0].label[191] , \labels[0].label[190] , 
	\labels[0].label[189] , \labels[0].label[188] , 
	\labels[0].label[187] , \labels[0].label[186] , 
	\labels[0].label[185] , \labels[0].label[184] , 
	\labels[0].label[183] , \labels[0].label[182] , 
	\labels[0].label[181] , \labels[0].label[180] , 
	\labels[0].label[179] , \labels[0].label[178] , 
	\labels[0].label[177] , \labels[0].label[176] , 
	\labels[0].label[175] , \labels[0].label[174] , 
	\labels[0].label[173] , \labels[0].label[172] , 
	\labels[0].label[171] , \labels[0].label[170] , 
	\labels[0].label[169] , \labels[0].label[168] , 
	\labels[0].label[167] , \labels[0].label[166] , 
	\labels[0].label[165] , \labels[0].label[164] , 
	\labels[0].label[163] , \labels[0].label[162] , 
	\labels[0].label[161] , \labels[0].label[160] , 
	\labels[0].label[159] , \labels[0].label[158] , 
	\labels[0].label[157] , \labels[0].label[156] , 
	\labels[0].label[155] , \labels[0].label[154] , 
	\labels[0].label[153] , \labels[0].label[152] , 
	\labels[0].label[151] , \labels[0].label[150] , 
	\labels[0].label[149] , \labels[0].label[148] , 
	\labels[0].label[147] , \labels[0].label[146] , 
	\labels[0].label[145] , \labels[0].label[144] , 
	\labels[0].label[143] , \labels[0].label[142] , 
	\labels[0].label[141] , \labels[0].label[140] , 
	\labels[0].label[139] , \labels[0].label[138] , 
	\labels[0].label[137] , \labels[0].label[136] , 
	\labels[0].label[135] , \labels[0].label[134] , 
	\labels[0].label[133] , \labels[0].label[132] , 
	\labels[0].label[131] , \labels[0].label[130] , 
	\labels[0].label[129] , \labels[0].label[128] , 
	\labels[0].label[127] , \labels[0].label[126] , 
	\labels[0].label[125] , \labels[0].label[124] , 
	\labels[0].label[123] , \labels[0].label[122] , 
	\labels[0].label[121] , \labels[0].label[120] , 
	\labels[0].label[119] , \labels[0].label[118] , 
	\labels[0].label[117] , \labels[0].label[116] , 
	\labels[0].label[115] , \labels[0].label[114] , 
	\labels[0].label[113] , \labels[0].label[112] , 
	\labels[0].label[111] , \labels[0].label[110] , 
	\labels[0].label[109] , \labels[0].label[108] , 
	\labels[0].label[107] , \labels[0].label[106] , 
	\labels[0].label[105] , \labels[0].label[104] , 
	\labels[0].label[103] , \labels[0].label[102] , 
	\labels[0].label[101] , \labels[0].label[100] , 
	\labels[0].label[99] , \labels[0].label[98] , \labels[0].label[97] , 
	\labels[0].label[96] , \labels[0].label[95] , \labels[0].label[94] , 
	\labels[0].label[93] , \labels[0].label[92] , \labels[0].label[91] , 
	\labels[0].label[90] , \labels[0].label[89] , \labels[0].label[88] , 
	\labels[0].label[87] , \labels[0].label[86] , \labels[0].label[85] , 
	\labels[0].label[84] , \labels[0].label[83] , \labels[0].label[82] , 
	\labels[0].label[81] , \labels[0].label[80] , \labels[0].label[79] , 
	\labels[0].label[78] , \labels[0].label[77] , \labels[0].label[76] , 
	\labels[0].label[75] , \labels[0].label[74] , \labels[0].label[73] , 
	\labels[0].label[72] , \labels[0].label[71] , \labels[0].label[70] , 
	\labels[0].label[69] , \labels[0].label[68] , \labels[0].label[67] , 
	\labels[0].label[66] , \labels[0].label[65] , \labels[0].label[64] , 
	\labels[0].label[63] , \labels[0].label[62] , \labels[0].label[61] , 
	\labels[0].label[60] , \labels[0].label[59] , \labels[0].label[58] , 
	\labels[0].label[57] , \labels[0].label[56] , \labels[0].label[55] , 
	\labels[0].label[54] , \labels[0].label[53] , \labels[0].label[52] , 
	\labels[0].label[51] , \labels[0].label[50] , \labels[0].label[49] , 
	\labels[0].label[48] , \labels[0].label[47] , \labels[0].label[46] , 
	\labels[0].label[45] , \labels[0].label[44] , \labels[0].label[43] , 
	\labels[0].label[42] , \labels[0].label[41] , \labels[0].label[40] , 
	\labels[0].label[39] , \labels[0].label[38] , \labels[0].label[37] , 
	\labels[0].label[36] , \labels[0].label[35] , \labels[0].label[34] , 
	\labels[0].label[33] , \labels[0].label[32] , \labels[0].label[31] , 
	\labels[0].label[30] , \labels[0].label[29] , \labels[0].label[28] , 
	\labels[0].label[27] , \labels[0].label[26] , \labels[0].label[25] , 
	\labels[0].label[24] , \labels[0].label[23] , \labels[0].label[22] , 
	\labels[0].label[21] , \labels[0].label[20] , \labels[0].label[19] , 
	\labels[0].label[18] , \labels[0].label[17] , \labels[0].label[16] , 
	\labels[0].label[15] , \labels[0].label[14] , \labels[0].label[13] , 
	\labels[0].label[12] , \labels[0].label[11] , \labels[0].label[10] , 
	\labels[0].label[9] , \labels[0].label[8] , \labels[0].label[7] , 
	\labels[0].label[6] , \labels[0].label[5] , \labels[0].label[4] , 
	\labels[0].label[3] , \labels[0].label[2] , \labels[0].label[1] , 
	\labels[0].label[0] , \labels[0].delimiter_valid[0] , 
	\labels[0].delimiter[7] , \labels[0].delimiter[6] , 
	\labels[0].delimiter[5] , \labels[0].delimiter[4] , 
	\labels[0].delimiter[3] , \labels[0].delimiter[2] , 
	\labels[0].delimiter[1] , \labels[0].delimiter[0] } ), 
	.kme_internal_out( {\kme_internal_out.sot [0], 
	\kme_internal_out.eoi [0], \kme_internal_out.eot [0], 
	\kme_internal_out.id [3], \kme_internal_out.id [2], 
	\kme_internal_out.id [1], \kme_internal_out.id [0], 
	\kme_internal_out.tdata [63], \kme_internal_out.tdata [62], 
	\kme_internal_out.tdata [61], \kme_internal_out.tdata [60], 
	\kme_internal_out.tdata [59], \kme_internal_out.tdata [58], 
	\kme_internal_out.tdata [57], \kme_internal_out.tdata [56], 
	\kme_internal_out.tdata [55], \kme_internal_out.tdata [54], 
	\kme_internal_out.tdata [53], \kme_internal_out.tdata [52], 
	\kme_internal_out.tdata [51], \kme_internal_out.tdata [50], 
	\kme_internal_out.tdata [49], \kme_internal_out.tdata [48], 
	\kme_internal_out.tdata [47], \kme_internal_out.tdata [46], 
	\kme_internal_out.tdata [45], \kme_internal_out.tdata [44], 
	\kme_internal_out.tdata [43], \kme_internal_out.tdata [42], 
	\kme_internal_out.tdata [41], \kme_internal_out.tdata [40], 
	\kme_internal_out.tdata [39], \kme_internal_out.tdata [38], 
	\kme_internal_out.tdata [37], \kme_internal_out.tdata [36], 
	\kme_internal_out.tdata [35], \kme_internal_out.tdata [34], 
	\kme_internal_out.tdata [33], \kme_internal_out.tdata [32], 
	\kme_internal_out.tdata [31], \kme_internal_out.tdata [30], 
	\kme_internal_out.tdata [29], \kme_internal_out.tdata [28], 
	\kme_internal_out.tdata [27], \kme_internal_out.tdata [26], 
	\kme_internal_out.tdata [25], \kme_internal_out.tdata [24], 
	\kme_internal_out.tdata [23], \kme_internal_out.tdata [22], 
	\kme_internal_out.tdata [21], \kme_internal_out.tdata [20], 
	\kme_internal_out.tdata [19], \kme_internal_out.tdata [18], 
	\kme_internal_out.tdata [17], \kme_internal_out.tdata [16], 
	\kme_internal_out.tdata [15], \kme_internal_out.tdata [14], 
	\kme_internal_out.tdata [13], \kme_internal_out.tdata [12], 
	\kme_internal_out.tdata [11], \kme_internal_out.tdata [10], 
	\kme_internal_out.tdata [9], \kme_internal_out.tdata [8], 
	\kme_internal_out.tdata [7], \kme_internal_out.tdata [6], 
	\kme_internal_out.tdata [5], \kme_internal_out.tdata [4], 
	\kme_internal_out.tdata [3], \kme_internal_out.tdata [2], 
	\kme_internal_out.tdata [1], \kme_internal_out.tdata [0]} ), 
	kme_internal_out_valid, gcm_cmd_in_stall, gcm_tag_data_in_stall, 
	upsizer_inspector_stall, keyfilter_cmd_in_stall, 
	kdfstream_cmd_in_stall, kdf_cmd_in_stall, tlv_sb_data_in_stall);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output kme_internal_out_ack;
output [255:0] \gcm_cmd_in.key0 ;
output [255:0] \gcm_cmd_in.key1 ;
output [95:0] \gcm_cmd_in.iv ;
output [2:0] \gcm_cmd_in.op ;
wire [610:0] gcm_cmd_in;
output gcm_cmd_in_valid;
output [95:0] gcm_tag_data_in;
output gcm_tag_data_in_valid;
output inspector_upsizer_valid;
output inspector_upsizer_eof;
output [63:0] inspector_upsizer_data;
output [0:0] \keyfilter_cmd_in.combo_mode ;
wire [0:0] keyfilter_cmd_in;
output keyfilter_cmd_in_valid;
output [0:0] \kdfstream_cmd_in.combo_mode ;
output [0:0] \kdfstream_cmd_in.skip ;
output [255:0] \kdfstream_cmd_in.guid ;
output [2:0] \kdfstream_cmd_in.label_index ;
output [1:0] \kdfstream_cmd_in.num_iter ;
wire [262:0] kdfstream_cmd_in;
output kdfstream_cmd_in_valid;
output [0:0] \kdf_cmd_in.kdf_dek_iter ;
output [0:0] \kdf_cmd_in.combo_mode ;
output [0:0] \kdf_cmd_in.dek_key_op ;
output [0:0] \kdf_cmd_in.dak_key_op ;
wire [3:0] kdf_cmd_in;
output kdf_cmd_in_valid;
output [63:0] tlv_sb_data_in;
output tlv_sb_data_in_valid;
input clk;
input rst_n;
input \labels[7].guid_size[0] ,\labels[7].label_size[5] 
	,\labels[7].label_size[4] ,\labels[7].label_size[3] 
	,\labels[7].label_size[2] ,\labels[7].label_size[1] 
	,\labels[7].label_size[0] ,\labels[7].label[255] 
	,\labels[7].label[254] ,\labels[7].label[253] ,\labels[7].label[252] 
	,\labels[7].label[251] ,\labels[7].label[250] ,\labels[7].label[249] 
	,\labels[7].label[248] ,\labels[7].label[247] ,\labels[7].label[246] 
	,\labels[7].label[245] ,\labels[7].label[244] ,\labels[7].label[243] 
	,\labels[7].label[242] ,\labels[7].label[241] ,\labels[7].label[240] 
	,\labels[7].label[239] ,\labels[7].label[238] ,\labels[7].label[237] 
	,\labels[7].label[236] ,\labels[7].label[235] ,\labels[7].label[234] 
	,\labels[7].label[233] ,\labels[7].label[232] ,\labels[7].label[231] 
	,\labels[7].label[230] ,\labels[7].label[229] ,\labels[7].label[228] 
	,\labels[7].label[227] ,\labels[7].label[226] ,\labels[7].label[225] 
	,\labels[7].label[224] ,\labels[7].label[223] ,\labels[7].label[222] 
	,\labels[7].label[221] ,\labels[7].label[220] ,\labels[7].label[219] 
	,\labels[7].label[218] ,\labels[7].label[217] ,\labels[7].label[216] 
	,\labels[7].label[215] ,\labels[7].label[214] ,\labels[7].label[213] 
	,\labels[7].label[212] ,\labels[7].label[211] ,\labels[7].label[210] 
	,\labels[7].label[209] ,\labels[7].label[208] ,\labels[7].label[207] 
	,\labels[7].label[206] ,\labels[7].label[205] ,\labels[7].label[204] 
	,\labels[7].label[203] ,\labels[7].label[202] ,\labels[7].label[201] 
	,\labels[7].label[200] ,\labels[7].label[199] ,\labels[7].label[198] 
	,\labels[7].label[197] ,\labels[7].label[196] ,\labels[7].label[195] 
	,\labels[7].label[194] ,\labels[7].label[193] ,\labels[7].label[192] 
	,\labels[7].label[191] ,\labels[7].label[190] ,\labels[7].label[189] 
	,\labels[7].label[188] ,\labels[7].label[187] ,\labels[7].label[186] 
	,\labels[7].label[185] ,\labels[7].label[184] ,\labels[7].label[183] 
	,\labels[7].label[182] ,\labels[7].label[181] ,\labels[7].label[180] 
	,\labels[7].label[179] ,\labels[7].label[178] ,\labels[7].label[177] 
	,\labels[7].label[176] ,\labels[7].label[175] ,\labels[7].label[174] 
	,\labels[7].label[173] ,\labels[7].label[172] ,\labels[7].label[171] 
	,\labels[7].label[170] ,\labels[7].label[169] ,\labels[7].label[168] 
	,\labels[7].label[167] ,\labels[7].label[166] ,\labels[7].label[165] 
	,\labels[7].label[164] ,\labels[7].label[163] ,\labels[7].label[162] 
	,\labels[7].label[161] ,\labels[7].label[160] ,\labels[7].label[159] 
	,\labels[7].label[158] ,\labels[7].label[157] ,\labels[7].label[156] 
	,\labels[7].label[155] ,\labels[7].label[154] ,\labels[7].label[153] 
	,\labels[7].label[152] ,\labels[7].label[151] ,\labels[7].label[150] 
	,\labels[7].label[149] ,\labels[7].label[148] ,\labels[7].label[147] 
	,\labels[7].label[146] ,\labels[7].label[145] ,\labels[7].label[144] 
	,\labels[7].label[143] ,\labels[7].label[142] ,\labels[7].label[141] 
	,\labels[7].label[140] ,\labels[7].label[139] ,\labels[7].label[138] 
	,\labels[7].label[137] ,\labels[7].label[136] ,\labels[7].label[135] 
	,\labels[7].label[134] ,\labels[7].label[133] ,\labels[7].label[132] 
	,\labels[7].label[131] ,\labels[7].label[130] ,\labels[7].label[129] 
	,\labels[7].label[128] ,\labels[7].label[127] ,\labels[7].label[126] 
	,\labels[7].label[125] ,\labels[7].label[124] ,\labels[7].label[123] 
	,\labels[7].label[122] ,\labels[7].label[121] ,\labels[7].label[120] 
	,\labels[7].label[119] ,\labels[7].label[118] ,\labels[7].label[117] 
	,\labels[7].label[116] ,\labels[7].label[115] ,\labels[7].label[114] 
	,\labels[7].label[113] ,\labels[7].label[112] ,\labels[7].label[111] 
	,\labels[7].label[110] ,\labels[7].label[109] ,\labels[7].label[108] 
	,\labels[7].label[107] ,\labels[7].label[106] ,\labels[7].label[105] 
	,\labels[7].label[104] ,\labels[7].label[103] ,\labels[7].label[102] 
	,\labels[7].label[101] ,\labels[7].label[100] ,\labels[7].label[99] 
	,\labels[7].label[98] ,\labels[7].label[97] ,\labels[7].label[96] 
	,\labels[7].label[95] ,\labels[7].label[94] ,\labels[7].label[93] 
	,\labels[7].label[92] ,\labels[7].label[91] ,\labels[7].label[90] 
	,\labels[7].label[89] ,\labels[7].label[88] ,\labels[7].label[87] 
	,\labels[7].label[86] ,\labels[7].label[85] ,\labels[7].label[84] 
	,\labels[7].label[83] ,\labels[7].label[82] ,\labels[7].label[81] 
	,\labels[7].label[80] ,\labels[7].label[79] ,\labels[7].label[78] 
	,\labels[7].label[77] ,\labels[7].label[76] ,\labels[7].label[75] 
	,\labels[7].label[74] ,\labels[7].label[73] ,\labels[7].label[72] 
	,\labels[7].label[71] ,\labels[7].label[70] ,\labels[7].label[69] 
	,\labels[7].label[68] ,\labels[7].label[67] ,\labels[7].label[66] 
	,\labels[7].label[65] ,\labels[7].label[64] ,\labels[7].label[63] 
	,\labels[7].label[62] ,\labels[7].label[61] ,\labels[7].label[60] 
	,\labels[7].label[59] ,\labels[7].label[58] ,\labels[7].label[57] 
	,\labels[7].label[56] ,\labels[7].label[55] ,\labels[7].label[54] 
	,\labels[7].label[53] ,\labels[7].label[52] ,\labels[7].label[51] 
	,\labels[7].label[50] ,\labels[7].label[49] ,\labels[7].label[48] 
	,\labels[7].label[47] ,\labels[7].label[46] ,\labels[7].label[45] 
	,\labels[7].label[44] ,\labels[7].label[43] ,\labels[7].label[42] 
	,\labels[7].label[41] ,\labels[7].label[40] ,\labels[7].label[39] 
	,\labels[7].label[38] ,\labels[7].label[37] ,\labels[7].label[36] 
	,\labels[7].label[35] ,\labels[7].label[34] ,\labels[7].label[33] 
	,\labels[7].label[32] ,\labels[7].label[31] ,\labels[7].label[30] 
	,\labels[7].label[29] ,\labels[7].label[28] ,\labels[7].label[27] 
	,\labels[7].label[26] ,\labels[7].label[25] ,\labels[7].label[24] 
	,\labels[7].label[23] ,\labels[7].label[22] ,\labels[7].label[21] 
	,\labels[7].label[20] ,\labels[7].label[19] ,\labels[7].label[18] 
	,\labels[7].label[17] ,\labels[7].label[16] ,\labels[7].label[15] 
	,\labels[7].label[14] ,\labels[7].label[13] ,\labels[7].label[12] 
	,\labels[7].label[11] ,\labels[7].label[10] ,\labels[7].label[9] 
	,\labels[7].label[8] ,\labels[7].label[7] ,\labels[7].label[6] 
	,\labels[7].label[5] ,\labels[7].label[4] ,\labels[7].label[3] 
	,\labels[7].label[2] ,\labels[7].label[1] ,\labels[7].label[0] 
	,\labels[7].delimiter_valid[0] ,\labels[7].delimiter[7] 
	,\labels[7].delimiter[6] ,\labels[7].delimiter[5] 
	,\labels[7].delimiter[4] ,\labels[7].delimiter[3] 
	,\labels[7].delimiter[2] ,\labels[7].delimiter[1] 
	,\labels[7].delimiter[0] ,\labels[6].guid_size[0] 
	,\labels[6].label_size[5] ,\labels[6].label_size[4] 
	,\labels[6].label_size[3] ,\labels[6].label_size[2] 
	,\labels[6].label_size[1] ,\labels[6].label_size[0] 
	,\labels[6].label[255] ,\labels[6].label[254] ,\labels[6].label[253] 
	,\labels[6].label[252] ,\labels[6].label[251] ,\labels[6].label[250] 
	,\labels[6].label[249] ,\labels[6].label[248] ,\labels[6].label[247] 
	,\labels[6].label[246] ,\labels[6].label[245] ,\labels[6].label[244] 
	,\labels[6].label[243] ,\labels[6].label[242] ,\labels[6].label[241] 
	,\labels[6].label[240] ,\labels[6].label[239] ,\labels[6].label[238] 
	,\labels[6].label[237] ,\labels[6].label[236] ,\labels[6].label[235] 
	,\labels[6].label[234] ,\labels[6].label[233] ,\labels[6].label[232] 
	,\labels[6].label[231] ,\labels[6].label[230] ,\labels[6].label[229] 
	,\labels[6].label[228] ,\labels[6].label[227] ,\labels[6].label[226] 
	,\labels[6].label[225] ,\labels[6].label[224] ,\labels[6].label[223] 
	,\labels[6].label[222] ,\labels[6].label[221] ,\labels[6].label[220] 
	,\labels[6].label[219] ,\labels[6].label[218] ,\labels[6].label[217] 
	,\labels[6].label[216] ,\labels[6].label[215] ,\labels[6].label[214] 
	,\labels[6].label[213] ,\labels[6].label[212] ,\labels[6].label[211] 
	,\labels[6].label[210] ,\labels[6].label[209] ,\labels[6].label[208] 
	,\labels[6].label[207] ,\labels[6].label[206] ,\labels[6].label[205] 
	,\labels[6].label[204] ,\labels[6].label[203] ,\labels[6].label[202] 
	,\labels[6].label[201] ,\labels[6].label[200] ,\labels[6].label[199] 
	,\labels[6].label[198] ,\labels[6].label[197] ,\labels[6].label[196] 
	,\labels[6].label[195] ,\labels[6].label[194] ,\labels[6].label[193] 
	,\labels[6].label[192] ,\labels[6].label[191] ,\labels[6].label[190] 
	,\labels[6].label[189] ,\labels[6].label[188] ,\labels[6].label[187] 
	,\labels[6].label[186] ,\labels[6].label[185] ,\labels[6].label[184] 
	,\labels[6].label[183] ,\labels[6].label[182] ,\labels[6].label[181] 
	,\labels[6].label[180] ,\labels[6].label[179] ,\labels[6].label[178] 
	,\labels[6].label[177] ,\labels[6].label[176] ,\labels[6].label[175] 
	,\labels[6].label[174] ,\labels[6].label[173] ,\labels[6].label[172] 
	,\labels[6].label[171] ,\labels[6].label[170] ,\labels[6].label[169] 
	,\labels[6].label[168] ,\labels[6].label[167] ,\labels[6].label[166] 
	,\labels[6].label[165] ,\labels[6].label[164] ,\labels[6].label[163] 
	,\labels[6].label[162] ,\labels[6].label[161] ,\labels[6].label[160] 
	,\labels[6].label[159] ,\labels[6].label[158] ,\labels[6].label[157] 
	,\labels[6].label[156] ,\labels[6].label[155] ,\labels[6].label[154] 
	,\labels[6].label[153] ,\labels[6].label[152] ,\labels[6].label[151] 
	,\labels[6].label[150] ,\labels[6].label[149] ,\labels[6].label[148] 
	,\labels[6].label[147] ,\labels[6].label[146] ,\labels[6].label[145] 
	,\labels[6].label[144] ,\labels[6].label[143] ,\labels[6].label[142] 
	,\labels[6].label[141] ,\labels[6].label[140] ,\labels[6].label[139] 
	,\labels[6].label[138] ,\labels[6].label[137] ,\labels[6].label[136] 
	,\labels[6].label[135] ,\labels[6].label[134] ,\labels[6].label[133] 
	,\labels[6].label[132] ,\labels[6].label[131] ,\labels[6].label[130] 
	,\labels[6].label[129] ,\labels[6].label[128] ,\labels[6].label[127] 
	,\labels[6].label[126] ,\labels[6].label[125] ,\labels[6].label[124] 
	,\labels[6].label[123] ,\labels[6].label[122] ,\labels[6].label[121] 
	,\labels[6].label[120] ,\labels[6].label[119] ,\labels[6].label[118] 
	,\labels[6].label[117] ,\labels[6].label[116] ,\labels[6].label[115] 
	,\labels[6].label[114] ,\labels[6].label[113] ,\labels[6].label[112] 
	,\labels[6].label[111] ,\labels[6].label[110] ,\labels[6].label[109] 
	,\labels[6].label[108] ,\labels[6].label[107] ,\labels[6].label[106] 
	,\labels[6].label[105] ,\labels[6].label[104] ,\labels[6].label[103] 
	,\labels[6].label[102] ,\labels[6].label[101] ,\labels[6].label[100] 
	,\labels[6].label[99] ,\labels[6].label[98] ,\labels[6].label[97] 
	,\labels[6].label[96] ,\labels[6].label[95] ,\labels[6].label[94] 
	,\labels[6].label[93] ,\labels[6].label[92] ,\labels[6].label[91] 
	,\labels[6].label[90] ,\labels[6].label[89] ,\labels[6].label[88] 
	,\labels[6].label[87] ,\labels[6].label[86] ,\labels[6].label[85] 
	,\labels[6].label[84] ,\labels[6].label[83] ,\labels[6].label[82] 
	,\labels[6].label[81] ,\labels[6].label[80] ,\labels[6].label[79] 
	,\labels[6].label[78] ,\labels[6].label[77] ,\labels[6].label[76] 
	,\labels[6].label[75] ,\labels[6].label[74] ,\labels[6].label[73] 
	,\labels[6].label[72] ,\labels[6].label[71] ,\labels[6].label[70] 
	,\labels[6].label[69] ,\labels[6].label[68] ,\labels[6].label[67] 
	,\labels[6].label[66] ,\labels[6].label[65] ,\labels[6].label[64] 
	,\labels[6].label[63] ,\labels[6].label[62] ,\labels[6].label[61] 
	,\labels[6].label[60] ,\labels[6].label[59] ,\labels[6].label[58] 
	,\labels[6].label[57] ,\labels[6].label[56] ,\labels[6].label[55] 
	,\labels[6].label[54] ,\labels[6].label[53] ,\labels[6].label[52] 
	,\labels[6].label[51] ,\labels[6].label[50] ,\labels[6].label[49] 
	,\labels[6].label[48] ,\labels[6].label[47] ,\labels[6].label[46] 
	,\labels[6].label[45] ,\labels[6].label[44] ,\labels[6].label[43] 
	,\labels[6].label[42] ,\labels[6].label[41] ,\labels[6].label[40] 
	,\labels[6].label[39] ,\labels[6].label[38] ,\labels[6].label[37] 
	,\labels[6].label[36] ,\labels[6].label[35] ,\labels[6].label[34] 
	,\labels[6].label[33] ,\labels[6].label[32] ,\labels[6].label[31] 
	,\labels[6].label[30] ,\labels[6].label[29] ,\labels[6].label[28] 
	,\labels[6].label[27] ,\labels[6].label[26] ,\labels[6].label[25] 
	,\labels[6].label[24] ,\labels[6].label[23] ,\labels[6].label[22] 
	,\labels[6].label[21] ,\labels[6].label[20] ,\labels[6].label[19] 
	,\labels[6].label[18] ,\labels[6].label[17] ,\labels[6].label[16] 
	,\labels[6].label[15] ,\labels[6].label[14] ,\labels[6].label[13] 
	,\labels[6].label[12] ,\labels[6].label[11] ,\labels[6].label[10] 
	,\labels[6].label[9] ,\labels[6].label[8] ,\labels[6].label[7] 
	,\labels[6].label[6] ,\labels[6].label[5] ,\labels[6].label[4] 
	,\labels[6].label[3] ,\labels[6].label[2] ,\labels[6].label[1] 
	,\labels[6].label[0] ,\labels[6].delimiter_valid[0] 
	,\labels[6].delimiter[7] ,\labels[6].delimiter[6] 
	,\labels[6].delimiter[5] ,\labels[6].delimiter[4] 
	,\labels[6].delimiter[3] ,\labels[6].delimiter[2] 
	,\labels[6].delimiter[1] ,\labels[6].delimiter[0] 
	,\labels[5].guid_size[0] ,\labels[5].label_size[5] 
	,\labels[5].label_size[4] ,\labels[5].label_size[3] 
	,\labels[5].label_size[2] ,\labels[5].label_size[1] 
	,\labels[5].label_size[0] ,\labels[5].label[255] 
	,\labels[5].label[254] ,\labels[5].label[253] ,\labels[5].label[252] 
	,\labels[5].label[251] ,\labels[5].label[250] ,\labels[5].label[249] 
	,\labels[5].label[248] ,\labels[5].label[247] ,\labels[5].label[246] 
	,\labels[5].label[245] ,\labels[5].label[244] ,\labels[5].label[243] 
	,\labels[5].label[242] ,\labels[5].label[241] ,\labels[5].label[240] 
	,\labels[5].label[239] ,\labels[5].label[238] ,\labels[5].label[237] 
	,\labels[5].label[236] ,\labels[5].label[235] ,\labels[5].label[234] 
	,\labels[5].label[233] ,\labels[5].label[232] ,\labels[5].label[231] 
	,\labels[5].label[230] ,\labels[5].label[229] ,\labels[5].label[228] 
	,\labels[5].label[227] ,\labels[5].label[226] ,\labels[5].label[225] 
	,\labels[5].label[224] ,\labels[5].label[223] ,\labels[5].label[222] 
	,\labels[5].label[221] ,\labels[5].label[220] ,\labels[5].label[219] 
	,\labels[5].label[218] ,\labels[5].label[217] ,\labels[5].label[216] 
	,\labels[5].label[215] ,\labels[5].label[214] ,\labels[5].label[213] 
	,\labels[5].label[212] ,\labels[5].label[211] ,\labels[5].label[210] 
	,\labels[5].label[209] ,\labels[5].label[208] ,\labels[5].label[207] 
	,\labels[5].label[206] ,\labels[5].label[205] ,\labels[5].label[204] 
	,\labels[5].label[203] ,\labels[5].label[202] ,\labels[5].label[201] 
	,\labels[5].label[200] ,\labels[5].label[199] ,\labels[5].label[198] 
	,\labels[5].label[197] ,\labels[5].label[196] ,\labels[5].label[195] 
	,\labels[5].label[194] ,\labels[5].label[193] ,\labels[5].label[192] 
	,\labels[5].label[191] ,\labels[5].label[190] ,\labels[5].label[189] 
	,\labels[5].label[188] ,\labels[5].label[187] ,\labels[5].label[186] 
	,\labels[5].label[185] ,\labels[5].label[184] ,\labels[5].label[183] 
	,\labels[5].label[182] ,\labels[5].label[181] ,\labels[5].label[180] 
	,\labels[5].label[179] ,\labels[5].label[178] ,\labels[5].label[177] 
	,\labels[5].label[176] ,\labels[5].label[175] ,\labels[5].label[174] 
	,\labels[5].label[173] ,\labels[5].label[172] ,\labels[5].label[171] 
	,\labels[5].label[170] ,\labels[5].label[169] ,\labels[5].label[168] 
	,\labels[5].label[167] ,\labels[5].label[166] ,\labels[5].label[165] 
	,\labels[5].label[164] ,\labels[5].label[163] ,\labels[5].label[162] 
	,\labels[5].label[161] ,\labels[5].label[160] ,\labels[5].label[159] 
	,\labels[5].label[158] ,\labels[5].label[157] ,\labels[5].label[156] 
	,\labels[5].label[155] ,\labels[5].label[154] ,\labels[5].label[153] 
	,\labels[5].label[152] ,\labels[5].label[151] ,\labels[5].label[150] 
	,\labels[5].label[149] ,\labels[5].label[148] ,\labels[5].label[147] 
	,\labels[5].label[146] ,\labels[5].label[145] ,\labels[5].label[144] 
	,\labels[5].label[143] ,\labels[5].label[142] ,\labels[5].label[141] 
	,\labels[5].label[140] ,\labels[5].label[139] ,\labels[5].label[138] 
	,\labels[5].label[137] ,\labels[5].label[136] ,\labels[5].label[135] 
	,\labels[5].label[134] ,\labels[5].label[133] ,\labels[5].label[132] 
	,\labels[5].label[131] ,\labels[5].label[130] ,\labels[5].label[129] 
	,\labels[5].label[128] ,\labels[5].label[127] ,\labels[5].label[126] 
	,\labels[5].label[125] ,\labels[5].label[124] ,\labels[5].label[123] 
	,\labels[5].label[122] ,\labels[5].label[121] ,\labels[5].label[120] 
	,\labels[5].label[119] ,\labels[5].label[118] ,\labels[5].label[117] 
	,\labels[5].label[116] ,\labels[5].label[115] ,\labels[5].label[114] 
	,\labels[5].label[113] ,\labels[5].label[112] ,\labels[5].label[111] 
	,\labels[5].label[110] ,\labels[5].label[109] ,\labels[5].label[108] 
	,\labels[5].label[107] ,\labels[5].label[106] ,\labels[5].label[105] 
	,\labels[5].label[104] ,\labels[5].label[103] ,\labels[5].label[102] 
	,\labels[5].label[101] ,\labels[5].label[100] ,\labels[5].label[99] 
	,\labels[5].label[98] ,\labels[5].label[97] ,\labels[5].label[96] 
	,\labels[5].label[95] ,\labels[5].label[94] ,\labels[5].label[93] 
	,\labels[5].label[92] ,\labels[5].label[91] ,\labels[5].label[90] 
	,\labels[5].label[89] ,\labels[5].label[88] ,\labels[5].label[87] 
	,\labels[5].label[86] ,\labels[5].label[85] ,\labels[5].label[84] 
	,\labels[5].label[83] ,\labels[5].label[82] ,\labels[5].label[81] 
	,\labels[5].label[80] ,\labels[5].label[79] ,\labels[5].label[78] 
	,\labels[5].label[77] ,\labels[5].label[76] ,\labels[5].label[75] 
	,\labels[5].label[74] ,\labels[5].label[73] ,\labels[5].label[72] 
	,\labels[5].label[71] ,\labels[5].label[70] ,\labels[5].label[69] 
	,\labels[5].label[68] ,\labels[5].label[67] ,\labels[5].label[66] 
	,\labels[5].label[65] ,\labels[5].label[64] ,\labels[5].label[63] 
	,\labels[5].label[62] ,\labels[5].label[61] ,\labels[5].label[60] 
	,\labels[5].label[59] ,\labels[5].label[58] ,\labels[5].label[57] 
	,\labels[5].label[56] ,\labels[5].label[55] ,\labels[5].label[54] 
	,\labels[5].label[53] ,\labels[5].label[52] ,\labels[5].label[51] 
	,\labels[5].label[50] ,\labels[5].label[49] ,\labels[5].label[48] 
	,\labels[5].label[47] ,\labels[5].label[46] ,\labels[5].label[45] 
	,\labels[5].label[44] ,\labels[5].label[43] ,\labels[5].label[42] 
	,\labels[5].label[41] ,\labels[5].label[40] ,\labels[5].label[39] 
	,\labels[5].label[38] ,\labels[5].label[37] ,\labels[5].label[36] 
	,\labels[5].label[35] ,\labels[5].label[34] ,\labels[5].label[33] 
	,\labels[5].label[32] ,\labels[5].label[31] ,\labels[5].label[30] 
	,\labels[5].label[29] ,\labels[5].label[28] ,\labels[5].label[27] 
	,\labels[5].label[26] ,\labels[5].label[25] ,\labels[5].label[24] 
	,\labels[5].label[23] ,\labels[5].label[22] ,\labels[5].label[21] 
	,\labels[5].label[20] ,\labels[5].label[19] ,\labels[5].label[18] 
	,\labels[5].label[17] ,\labels[5].label[16] ,\labels[5].label[15] 
	,\labels[5].label[14] ,\labels[5].label[13] ,\labels[5].label[12] 
	,\labels[5].label[11] ,\labels[5].label[10] ,\labels[5].label[9] 
	,\labels[5].label[8] ,\labels[5].label[7] ,\labels[5].label[6] 
	,\labels[5].label[5] ,\labels[5].label[4] ,\labels[5].label[3] 
	,\labels[5].label[2] ,\labels[5].label[1] ,\labels[5].label[0] 
	,\labels[5].delimiter_valid[0] ,\labels[5].delimiter[7] 
	,\labels[5].delimiter[6] ,\labels[5].delimiter[5] 
	,\labels[5].delimiter[4] ,\labels[5].delimiter[3] 
	,\labels[5].delimiter[2] ,\labels[5].delimiter[1] 
	,\labels[5].delimiter[0] ,\labels[4].guid_size[0] 
	,\labels[4].label_size[5] ,\labels[4].label_size[4] 
	,\labels[4].label_size[3] ,\labels[4].label_size[2] 
	,\labels[4].label_size[1] ,\labels[4].label_size[0] 
	,\labels[4].label[255] ,\labels[4].label[254] ,\labels[4].label[253] 
	,\labels[4].label[252] ,\labels[4].label[251] ,\labels[4].label[250] 
	,\labels[4].label[249] ,\labels[4].label[248] ,\labels[4].label[247] 
	,\labels[4].label[246] ,\labels[4].label[245] ,\labels[4].label[244] 
	,\labels[4].label[243] ,\labels[4].label[242] ,\labels[4].label[241] 
	,\labels[4].label[240] ,\labels[4].label[239] ,\labels[4].label[238] 
	,\labels[4].label[237] ,\labels[4].label[236] ,\labels[4].label[235] 
	,\labels[4].label[234] ,\labels[4].label[233] ,\labels[4].label[232] 
	,\labels[4].label[231] ,\labels[4].label[230] ,\labels[4].label[229] 
	,\labels[4].label[228] ,\labels[4].label[227] ,\labels[4].label[226] 
	,\labels[4].label[225] ,\labels[4].label[224] ,\labels[4].label[223] 
	,\labels[4].label[222] ,\labels[4].label[221] ,\labels[4].label[220] 
	,\labels[4].label[219] ,\labels[4].label[218] ,\labels[4].label[217] 
	,\labels[4].label[216] ,\labels[4].label[215] ,\labels[4].label[214] 
	,\labels[4].label[213] ,\labels[4].label[212] ,\labels[4].label[211] 
	,\labels[4].label[210] ,\labels[4].label[209] ,\labels[4].label[208] 
	,\labels[4].label[207] ,\labels[4].label[206] ,\labels[4].label[205] 
	,\labels[4].label[204] ,\labels[4].label[203] ,\labels[4].label[202] 
	,\labels[4].label[201] ,\labels[4].label[200] ,\labels[4].label[199] 
	,\labels[4].label[198] ,\labels[4].label[197] ,\labels[4].label[196] 
	,\labels[4].label[195] ,\labels[4].label[194] ,\labels[4].label[193] 
	,\labels[4].label[192] ,\labels[4].label[191] ,\labels[4].label[190] 
	,\labels[4].label[189] ,\labels[4].label[188] ,\labels[4].label[187] 
	,\labels[4].label[186] ,\labels[4].label[185] ,\labels[4].label[184] 
	,\labels[4].label[183] ,\labels[4].label[182] ,\labels[4].label[181] 
	,\labels[4].label[180] ,\labels[4].label[179] ,\labels[4].label[178] 
	,\labels[4].label[177] ,\labels[4].label[176] ,\labels[4].label[175] 
	,\labels[4].label[174] ,\labels[4].label[173] ,\labels[4].label[172] 
	,\labels[4].label[171] ,\labels[4].label[170] ,\labels[4].label[169] 
	,\labels[4].label[168] ,\labels[4].label[167] ,\labels[4].label[166] 
	,\labels[4].label[165] ,\labels[4].label[164] ,\labels[4].label[163] 
	,\labels[4].label[162] ,\labels[4].label[161] ,\labels[4].label[160] 
	,\labels[4].label[159] ,\labels[4].label[158] ,\labels[4].label[157] 
	,\labels[4].label[156] ,\labels[4].label[155] ,\labels[4].label[154] 
	,\labels[4].label[153] ,\labels[4].label[152] ,\labels[4].label[151] 
	,\labels[4].label[150] ,\labels[4].label[149] ,\labels[4].label[148] 
	,\labels[4].label[147] ,\labels[4].label[146] ,\labels[4].label[145] 
	,\labels[4].label[144] ,\labels[4].label[143] ,\labels[4].label[142] 
	,\labels[4].label[141] ,\labels[4].label[140] ,\labels[4].label[139] 
	,\labels[4].label[138] ,\labels[4].label[137] ,\labels[4].label[136] 
	,\labels[4].label[135] ,\labels[4].label[134] ,\labels[4].label[133] 
	,\labels[4].label[132] ,\labels[4].label[131] ,\labels[4].label[130] 
	,\labels[4].label[129] ,\labels[4].label[128] ,\labels[4].label[127] 
	,\labels[4].label[126] ,\labels[4].label[125] ,\labels[4].label[124] 
	,\labels[4].label[123] ,\labels[4].label[122] ,\labels[4].label[121] 
	,\labels[4].label[120] ,\labels[4].label[119] ,\labels[4].label[118] 
	,\labels[4].label[117] ,\labels[4].label[116] ,\labels[4].label[115] 
	,\labels[4].label[114] ,\labels[4].label[113] ,\labels[4].label[112] 
	,\labels[4].label[111] ,\labels[4].label[110] ,\labels[4].label[109] 
	,\labels[4].label[108] ,\labels[4].label[107] ,\labels[4].label[106] 
	,\labels[4].label[105] ,\labels[4].label[104] ,\labels[4].label[103] 
	,\labels[4].label[102] ,\labels[4].label[101] ,\labels[4].label[100] 
	,\labels[4].label[99] ,\labels[4].label[98] ,\labels[4].label[97] 
	,\labels[4].label[96] ,\labels[4].label[95] ,\labels[4].label[94] 
	,\labels[4].label[93] ,\labels[4].label[92] ,\labels[4].label[91] 
	,\labels[4].label[90] ,\labels[4].label[89] ,\labels[4].label[88] 
	,\labels[4].label[87] ,\labels[4].label[86] ,\labels[4].label[85] 
	,\labels[4].label[84] ,\labels[4].label[83] ,\labels[4].label[82] 
	,\labels[4].label[81] ,\labels[4].label[80] ,\labels[4].label[79] 
	,\labels[4].label[78] ,\labels[4].label[77] ,\labels[4].label[76] 
	,\labels[4].label[75] ,\labels[4].label[74] ,\labels[4].label[73] 
	,\labels[4].label[72] ,\labels[4].label[71] ,\labels[4].label[70] 
	,\labels[4].label[69] ,\labels[4].label[68] ,\labels[4].label[67] 
	,\labels[4].label[66] ,\labels[4].label[65] ,\labels[4].label[64] 
	,\labels[4].label[63] ,\labels[4].label[62] ,\labels[4].label[61] 
	,\labels[4].label[60] ,\labels[4].label[59] ,\labels[4].label[58] 
	,\labels[4].label[57] ,\labels[4].label[56] ,\labels[4].label[55] 
	,\labels[4].label[54] ,\labels[4].label[53] ,\labels[4].label[52] 
	,\labels[4].label[51] ,\labels[4].label[50] ,\labels[4].label[49] 
	,\labels[4].label[48] ,\labels[4].label[47] ,\labels[4].label[46] 
	,\labels[4].label[45] ,\labels[4].label[44] ,\labels[4].label[43] 
	,\labels[4].label[42] ,\labels[4].label[41] ,\labels[4].label[40] 
	,\labels[4].label[39] ,\labels[4].label[38] ,\labels[4].label[37] 
	,\labels[4].label[36] ,\labels[4].label[35] ,\labels[4].label[34] 
	,\labels[4].label[33] ,\labels[4].label[32] ,\labels[4].label[31] 
	,\labels[4].label[30] ,\labels[4].label[29] ,\labels[4].label[28] 
	,\labels[4].label[27] ,\labels[4].label[26] ,\labels[4].label[25] 
	,\labels[4].label[24] ,\labels[4].label[23] ,\labels[4].label[22] 
	,\labels[4].label[21] ,\labels[4].label[20] ,\labels[4].label[19] 
	,\labels[4].label[18] ,\labels[4].label[17] ,\labels[4].label[16] 
	,\labels[4].label[15] ,\labels[4].label[14] ,\labels[4].label[13] 
	,\labels[4].label[12] ,\labels[4].label[11] ,\labels[4].label[10] 
	,\labels[4].label[9] ,\labels[4].label[8] ,\labels[4].label[7] 
	,\labels[4].label[6] ,\labels[4].label[5] ,\labels[4].label[4] 
	,\labels[4].label[3] ,\labels[4].label[2] ,\labels[4].label[1] 
	,\labels[4].label[0] ,\labels[4].delimiter_valid[0] 
	,\labels[4].delimiter[7] ,\labels[4].delimiter[6] 
	,\labels[4].delimiter[5] ,\labels[4].delimiter[4] 
	,\labels[4].delimiter[3] ,\labels[4].delimiter[2] 
	,\labels[4].delimiter[1] ,\labels[4].delimiter[0] 
	,\labels[3].guid_size[0] ,\labels[3].label_size[5] 
	,\labels[3].label_size[4] ,\labels[3].label_size[3] 
	,\labels[3].label_size[2] ,\labels[3].label_size[1] 
	,\labels[3].label_size[0] ,\labels[3].label[255] 
	,\labels[3].label[254] ,\labels[3].label[253] ,\labels[3].label[252] 
	,\labels[3].label[251] ,\labels[3].label[250] ,\labels[3].label[249] 
	,\labels[3].label[248] ,\labels[3].label[247] ,\labels[3].label[246] 
	,\labels[3].label[245] ,\labels[3].label[244] ,\labels[3].label[243] 
	,\labels[3].label[242] ,\labels[3].label[241] ,\labels[3].label[240] 
	,\labels[3].label[239] ,\labels[3].label[238] ,\labels[3].label[237] 
	,\labels[3].label[236] ,\labels[3].label[235] ,\labels[3].label[234] 
	,\labels[3].label[233] ,\labels[3].label[232] ,\labels[3].label[231] 
	,\labels[3].label[230] ,\labels[3].label[229] ,\labels[3].label[228] 
	,\labels[3].label[227] ,\labels[3].label[226] ,\labels[3].label[225] 
	,\labels[3].label[224] ,\labels[3].label[223] ,\labels[3].label[222] 
	,\labels[3].label[221] ,\labels[3].label[220] ,\labels[3].label[219] 
	,\labels[3].label[218] ,\labels[3].label[217] ,\labels[3].label[216] 
	,\labels[3].label[215] ,\labels[3].label[214] ,\labels[3].label[213] 
	,\labels[3].label[212] ,\labels[3].label[211] ,\labels[3].label[210] 
	,\labels[3].label[209] ,\labels[3].label[208] ,\labels[3].label[207] 
	,\labels[3].label[206] ,\labels[3].label[205] ,\labels[3].label[204] 
	,\labels[3].label[203] ,\labels[3].label[202] ,\labels[3].label[201] 
	,\labels[3].label[200] ,\labels[3].label[199] ,\labels[3].label[198] 
	,\labels[3].label[197] ,\labels[3].label[196] ,\labels[3].label[195] 
	,\labels[3].label[194] ,\labels[3].label[193] ,\labels[3].label[192] 
	,\labels[3].label[191] ,\labels[3].label[190] ,\labels[3].label[189] 
	,\labels[3].label[188] ,\labels[3].label[187] ,\labels[3].label[186] 
	,\labels[3].label[185] ,\labels[3].label[184] ,\labels[3].label[183] 
	,\labels[3].label[182] ,\labels[3].label[181] ,\labels[3].label[180] 
	,\labels[3].label[179] ,\labels[3].label[178] ,\labels[3].label[177] 
	,\labels[3].label[176] ,\labels[3].label[175] ,\labels[3].label[174] 
	,\labels[3].label[173] ,\labels[3].label[172] ,\labels[3].label[171] 
	,\labels[3].label[170] ,\labels[3].label[169] ,\labels[3].label[168] 
	,\labels[3].label[167] ,\labels[3].label[166] ,\labels[3].label[165] 
	,\labels[3].label[164] ,\labels[3].label[163] ,\labels[3].label[162] 
	,\labels[3].label[161] ,\labels[3].label[160] ,\labels[3].label[159] 
	,\labels[3].label[158] ,\labels[3].label[157] ,\labels[3].label[156] 
	,\labels[3].label[155] ,\labels[3].label[154] ,\labels[3].label[153] 
	,\labels[3].label[152] ,\labels[3].label[151] ,\labels[3].label[150] 
	,\labels[3].label[149] ,\labels[3].label[148] ,\labels[3].label[147] 
	,\labels[3].label[146] ,\labels[3].label[145] ,\labels[3].label[144] 
	,\labels[3].label[143] ,\labels[3].label[142] ,\labels[3].label[141] 
	,\labels[3].label[140] ,\labels[3].label[139] ,\labels[3].label[138] 
	,\labels[3].label[137] ,\labels[3].label[136] ,\labels[3].label[135] 
	,\labels[3].label[134] ,\labels[3].label[133] ,\labels[3].label[132] 
	,\labels[3].label[131] ,\labels[3].label[130] ,\labels[3].label[129] 
	,\labels[3].label[128] ,\labels[3].label[127] ,\labels[3].label[126] 
	,\labels[3].label[125] ,\labels[3].label[124] ,\labels[3].label[123] 
	,\labels[3].label[122] ,\labels[3].label[121] ,\labels[3].label[120] 
	,\labels[3].label[119] ,\labels[3].label[118] ,\labels[3].label[117] 
	,\labels[3].label[116] ,\labels[3].label[115] ,\labels[3].label[114] 
	,\labels[3].label[113] ,\labels[3].label[112] ,\labels[3].label[111] 
	,\labels[3].label[110] ,\labels[3].label[109] ,\labels[3].label[108] 
	,\labels[3].label[107] ,\labels[3].label[106] ,\labels[3].label[105] 
	,\labels[3].label[104] ,\labels[3].label[103] ,\labels[3].label[102] 
	,\labels[3].label[101] ,\labels[3].label[100] ,\labels[3].label[99] 
	,\labels[3].label[98] ,\labels[3].label[97] ,\labels[3].label[96] 
	,\labels[3].label[95] ,\labels[3].label[94] ,\labels[3].label[93] 
	,\labels[3].label[92] ,\labels[3].label[91] ,\labels[3].label[90] 
	,\labels[3].label[89] ,\labels[3].label[88] ,\labels[3].label[87] 
	,\labels[3].label[86] ,\labels[3].label[85] ,\labels[3].label[84] 
	,\labels[3].label[83] ,\labels[3].label[82] ,\labels[3].label[81] 
	,\labels[3].label[80] ,\labels[3].label[79] ,\labels[3].label[78] 
	,\labels[3].label[77] ,\labels[3].label[76] ,\labels[3].label[75] 
	,\labels[3].label[74] ,\labels[3].label[73] ,\labels[3].label[72] 
	,\labels[3].label[71] ,\labels[3].label[70] ,\labels[3].label[69] 
	,\labels[3].label[68] ,\labels[3].label[67] ,\labels[3].label[66] 
	,\labels[3].label[65] ,\labels[3].label[64] ,\labels[3].label[63] 
	,\labels[3].label[62] ,\labels[3].label[61] ,\labels[3].label[60] 
	,\labels[3].label[59] ,\labels[3].label[58] ,\labels[3].label[57] 
	,\labels[3].label[56] ,\labels[3].label[55] ,\labels[3].label[54] 
	,\labels[3].label[53] ,\labels[3].label[52] ,\labels[3].label[51] 
	,\labels[3].label[50] ,\labels[3].label[49] ,\labels[3].label[48] 
	,\labels[3].label[47] ,\labels[3].label[46] ,\labels[3].label[45] 
	,\labels[3].label[44] ,\labels[3].label[43] ,\labels[3].label[42] 
	,\labels[3].label[41] ,\labels[3].label[40] ,\labels[3].label[39] 
	,\labels[3].label[38] ,\labels[3].label[37] ,\labels[3].label[36] 
	,\labels[3].label[35] ,\labels[3].label[34] ,\labels[3].label[33] 
	,\labels[3].label[32] ,\labels[3].label[31] ,\labels[3].label[30] 
	,\labels[3].label[29] ,\labels[3].label[28] ,\labels[3].label[27] 
	,\labels[3].label[26] ,\labels[3].label[25] ,\labels[3].label[24] 
	,\labels[3].label[23] ,\labels[3].label[22] ,\labels[3].label[21] 
	,\labels[3].label[20] ,\labels[3].label[19] ,\labels[3].label[18] 
	,\labels[3].label[17] ,\labels[3].label[16] ,\labels[3].label[15] 
	,\labels[3].label[14] ,\labels[3].label[13] ,\labels[3].label[12] 
	,\labels[3].label[11] ,\labels[3].label[10] ,\labels[3].label[9] 
	,\labels[3].label[8] ,\labels[3].label[7] ,\labels[3].label[6] 
	,\labels[3].label[5] ,\labels[3].label[4] ,\labels[3].label[3] 
	,\labels[3].label[2] ,\labels[3].label[1] ,\labels[3].label[0] 
	,\labels[3].delimiter_valid[0] ,\labels[3].delimiter[7] 
	,\labels[3].delimiter[6] ,\labels[3].delimiter[5] 
	,\labels[3].delimiter[4] ,\labels[3].delimiter[3] 
	,\labels[3].delimiter[2] ,\labels[3].delimiter[1] 
	,\labels[3].delimiter[0] ,\labels[2].guid_size[0] 
	,\labels[2].label_size[5] ,\labels[2].label_size[4] 
	,\labels[2].label_size[3] ,\labels[2].label_size[2] 
	,\labels[2].label_size[1] ,\labels[2].label_size[0] 
	,\labels[2].label[255] ,\labels[2].label[254] ,\labels[2].label[253] 
	,\labels[2].label[252] ,\labels[2].label[251] ,\labels[2].label[250] 
	,\labels[2].label[249] ,\labels[2].label[248] ,\labels[2].label[247] 
	,\labels[2].label[246] ,\labels[2].label[245] ,\labels[2].label[244] 
	,\labels[2].label[243] ,\labels[2].label[242] ,\labels[2].label[241] 
	,\labels[2].label[240] ,\labels[2].label[239] ,\labels[2].label[238] 
	,\labels[2].label[237] ,\labels[2].label[236] ,\labels[2].label[235] 
	,\labels[2].label[234] ,\labels[2].label[233] ,\labels[2].label[232] 
	,\labels[2].label[231] ,\labels[2].label[230] ,\labels[2].label[229] 
	,\labels[2].label[228] ,\labels[2].label[227] ,\labels[2].label[226] 
	,\labels[2].label[225] ,\labels[2].label[224] ,\labels[2].label[223] 
	,\labels[2].label[222] ,\labels[2].label[221] ,\labels[2].label[220] 
	,\labels[2].label[219] ,\labels[2].label[218] ,\labels[2].label[217] 
	,\labels[2].label[216] ,\labels[2].label[215] ,\labels[2].label[214] 
	,\labels[2].label[213] ,\labels[2].label[212] ,\labels[2].label[211] 
	,\labels[2].label[210] ,\labels[2].label[209] ,\labels[2].label[208] 
	,\labels[2].label[207] ,\labels[2].label[206] ,\labels[2].label[205] 
	,\labels[2].label[204] ,\labels[2].label[203] ,\labels[2].label[202] 
	,\labels[2].label[201] ,\labels[2].label[200] ,\labels[2].label[199] 
	,\labels[2].label[198] ,\labels[2].label[197] ,\labels[2].label[196] 
	,\labels[2].label[195] ,\labels[2].label[194] ,\labels[2].label[193] 
	,\labels[2].label[192] ,\labels[2].label[191] ,\labels[2].label[190] 
	,\labels[2].label[189] ,\labels[2].label[188] ,\labels[2].label[187] 
	,\labels[2].label[186] ,\labels[2].label[185] ,\labels[2].label[184] 
	,\labels[2].label[183] ,\labels[2].label[182] ,\labels[2].label[181] 
	,\labels[2].label[180] ,\labels[2].label[179] ,\labels[2].label[178] 
	,\labels[2].label[177] ,\labels[2].label[176] ,\labels[2].label[175] 
	,\labels[2].label[174] ,\labels[2].label[173] ,\labels[2].label[172] 
	,\labels[2].label[171] ,\labels[2].label[170] ,\labels[2].label[169] 
	,\labels[2].label[168] ,\labels[2].label[167] ,\labels[2].label[166] 
	,\labels[2].label[165] ,\labels[2].label[164] ,\labels[2].label[163] 
	,\labels[2].label[162] ,\labels[2].label[161] ,\labels[2].label[160] 
	,\labels[2].label[159] ,\labels[2].label[158] ,\labels[2].label[157] 
	,\labels[2].label[156] ,\labels[2].label[155] ,\labels[2].label[154] 
	,\labels[2].label[153] ,\labels[2].label[152] ,\labels[2].label[151] 
	,\labels[2].label[150] ,\labels[2].label[149] ,\labels[2].label[148] 
	,\labels[2].label[147] ,\labels[2].label[146] ,\labels[2].label[145] 
	,\labels[2].label[144] ,\labels[2].label[143] ,\labels[2].label[142] 
	,\labels[2].label[141] ,\labels[2].label[140] ,\labels[2].label[139] 
	,\labels[2].label[138] ,\labels[2].label[137] ,\labels[2].label[136] 
	,\labels[2].label[135] ,\labels[2].label[134] ,\labels[2].label[133] 
	,\labels[2].label[132] ,\labels[2].label[131] ,\labels[2].label[130] 
	,\labels[2].label[129] ,\labels[2].label[128] ,\labels[2].label[127] 
	,\labels[2].label[126] ,\labels[2].label[125] ,\labels[2].label[124] 
	,\labels[2].label[123] ,\labels[2].label[122] ,\labels[2].label[121] 
	,\labels[2].label[120] ,\labels[2].label[119] ,\labels[2].label[118] 
	,\labels[2].label[117] ,\labels[2].label[116] ,\labels[2].label[115] 
	,\labels[2].label[114] ,\labels[2].label[113] ,\labels[2].label[112] 
	,\labels[2].label[111] ,\labels[2].label[110] ,\labels[2].label[109] 
	,\labels[2].label[108] ,\labels[2].label[107] ,\labels[2].label[106] 
	,\labels[2].label[105] ,\labels[2].label[104] ,\labels[2].label[103] 
	,\labels[2].label[102] ,\labels[2].label[101] ,\labels[2].label[100] 
	,\labels[2].label[99] ,\labels[2].label[98] ,\labels[2].label[97] 
	,\labels[2].label[96] ,\labels[2].label[95] ,\labels[2].label[94] 
	,\labels[2].label[93] ,\labels[2].label[92] ,\labels[2].label[91] 
	,\labels[2].label[90] ,\labels[2].label[89] ,\labels[2].label[88] 
	,\labels[2].label[87] ,\labels[2].label[86] ,\labels[2].label[85] 
	,\labels[2].label[84] ,\labels[2].label[83] ,\labels[2].label[82] 
	,\labels[2].label[81] ,\labels[2].label[80] ,\labels[2].label[79] 
	,\labels[2].label[78] ,\labels[2].label[77] ,\labels[2].label[76] 
	,\labels[2].label[75] ,\labels[2].label[74] ,\labels[2].label[73] 
	,\labels[2].label[72] ,\labels[2].label[71] ,\labels[2].label[70] 
	,\labels[2].label[69] ,\labels[2].label[68] ,\labels[2].label[67] 
	,\labels[2].label[66] ,\labels[2].label[65] ,\labels[2].label[64] 
	,\labels[2].label[63] ,\labels[2].label[62] ,\labels[2].label[61] 
	,\labels[2].label[60] ,\labels[2].label[59] ,\labels[2].label[58] 
	,\labels[2].label[57] ,\labels[2].label[56] ,\labels[2].label[55] 
	,\labels[2].label[54] ,\labels[2].label[53] ,\labels[2].label[52] 
	,\labels[2].label[51] ,\labels[2].label[50] ,\labels[2].label[49] 
	,\labels[2].label[48] ,\labels[2].label[47] ,\labels[2].label[46] 
	,\labels[2].label[45] ,\labels[2].label[44] ,\labels[2].label[43] 
	,\labels[2].label[42] ,\labels[2].label[41] ,\labels[2].label[40] 
	,\labels[2].label[39] ,\labels[2].label[38] ,\labels[2].label[37] 
	,\labels[2].label[36] ,\labels[2].label[35] ,\labels[2].label[34] 
	,\labels[2].label[33] ,\labels[2].label[32] ,\labels[2].label[31] 
	,\labels[2].label[30] ,\labels[2].label[29] ,\labels[2].label[28] 
	,\labels[2].label[27] ,\labels[2].label[26] ,\labels[2].label[25] 
	,\labels[2].label[24] ,\labels[2].label[23] ,\labels[2].label[22] 
	,\labels[2].label[21] ,\labels[2].label[20] ,\labels[2].label[19] 
	,\labels[2].label[18] ,\labels[2].label[17] ,\labels[2].label[16] 
	,\labels[2].label[15] ,\labels[2].label[14] ,\labels[2].label[13] 
	,\labels[2].label[12] ,\labels[2].label[11] ,\labels[2].label[10] 
	,\labels[2].label[9] ,\labels[2].label[8] ,\labels[2].label[7] 
	,\labels[2].label[6] ,\labels[2].label[5] ,\labels[2].label[4] 
	,\labels[2].label[3] ,\labels[2].label[2] ,\labels[2].label[1] 
	,\labels[2].label[0] ,\labels[2].delimiter_valid[0] 
	,\labels[2].delimiter[7] ,\labels[2].delimiter[6] 
	,\labels[2].delimiter[5] ,\labels[2].delimiter[4] 
	,\labels[2].delimiter[3] ,\labels[2].delimiter[2] 
	,\labels[2].delimiter[1] ,\labels[2].delimiter[0] 
	,\labels[1].guid_size[0] ,\labels[1].label_size[5] 
	,\labels[1].label_size[4] ,\labels[1].label_size[3] 
	,\labels[1].label_size[2] ,\labels[1].label_size[1] 
	,\labels[1].label_size[0] ,\labels[1].label[255] 
	,\labels[1].label[254] ,\labels[1].label[253] ,\labels[1].label[252] 
	,\labels[1].label[251] ,\labels[1].label[250] ,\labels[1].label[249] 
	,\labels[1].label[248] ,\labels[1].label[247] ,\labels[1].label[246] 
	,\labels[1].label[245] ,\labels[1].label[244] ,\labels[1].label[243] 
	,\labels[1].label[242] ,\labels[1].label[241] ,\labels[1].label[240] 
	,\labels[1].label[239] ,\labels[1].label[238] ,\labels[1].label[237] 
	,\labels[1].label[236] ,\labels[1].label[235] ,\labels[1].label[234] 
	,\labels[1].label[233] ,\labels[1].label[232] ,\labels[1].label[231] 
	,\labels[1].label[230] ,\labels[1].label[229] ,\labels[1].label[228] 
	,\labels[1].label[227] ,\labels[1].label[226] ,\labels[1].label[225] 
	,\labels[1].label[224] ,\labels[1].label[223] ,\labels[1].label[222] 
	,\labels[1].label[221] ,\labels[1].label[220] ,\labels[1].label[219] 
	,\labels[1].label[218] ,\labels[1].label[217] ,\labels[1].label[216] 
	,\labels[1].label[215] ,\labels[1].label[214] ,\labels[1].label[213] 
	,\labels[1].label[212] ,\labels[1].label[211] ,\labels[1].label[210] 
	,\labels[1].label[209] ,\labels[1].label[208] ,\labels[1].label[207] 
	,\labels[1].label[206] ,\labels[1].label[205] ,\labels[1].label[204] 
	,\labels[1].label[203] ,\labels[1].label[202] ,\labels[1].label[201] 
	,\labels[1].label[200] ,\labels[1].label[199] ,\labels[1].label[198] 
	,\labels[1].label[197] ,\labels[1].label[196] ,\labels[1].label[195] 
	,\labels[1].label[194] ,\labels[1].label[193] ,\labels[1].label[192] 
	,\labels[1].label[191] ,\labels[1].label[190] ,\labels[1].label[189] 
	,\labels[1].label[188] ,\labels[1].label[187] ,\labels[1].label[186] 
	,\labels[1].label[185] ,\labels[1].label[184] ,\labels[1].label[183] 
	,\labels[1].label[182] ,\labels[1].label[181] ,\labels[1].label[180] 
	,\labels[1].label[179] ,\labels[1].label[178] ,\labels[1].label[177] 
	,\labels[1].label[176] ,\labels[1].label[175] ,\labels[1].label[174] 
	,\labels[1].label[173] ,\labels[1].label[172] ,\labels[1].label[171] 
	,\labels[1].label[170] ,\labels[1].label[169] ,\labels[1].label[168] 
	,\labels[1].label[167] ,\labels[1].label[166] ,\labels[1].label[165] 
	,\labels[1].label[164] ,\labels[1].label[163] ,\labels[1].label[162] 
	,\labels[1].label[161] ,\labels[1].label[160] ,\labels[1].label[159] 
	,\labels[1].label[158] ,\labels[1].label[157] ,\labels[1].label[156] 
	,\labels[1].label[155] ,\labels[1].label[154] ,\labels[1].label[153] 
	,\labels[1].label[152] ,\labels[1].label[151] ,\labels[1].label[150] 
	,\labels[1].label[149] ,\labels[1].label[148] ,\labels[1].label[147] 
	,\labels[1].label[146] ,\labels[1].label[145] ,\labels[1].label[144] 
	,\labels[1].label[143] ,\labels[1].label[142] ,\labels[1].label[141] 
	,\labels[1].label[140] ,\labels[1].label[139] ,\labels[1].label[138] 
	,\labels[1].label[137] ,\labels[1].label[136] ,\labels[1].label[135] 
	,\labels[1].label[134] ,\labels[1].label[133] ,\labels[1].label[132] 
	,\labels[1].label[131] ,\labels[1].label[130] ,\labels[1].label[129] 
	,\labels[1].label[128] ,\labels[1].label[127] ,\labels[1].label[126] 
	,\labels[1].label[125] ,\labels[1].label[124] ,\labels[1].label[123] 
	,\labels[1].label[122] ,\labels[1].label[121] ,\labels[1].label[120] 
	,\labels[1].label[119] ,\labels[1].label[118] ,\labels[1].label[117] 
	,\labels[1].label[116] ,\labels[1].label[115] ,\labels[1].label[114] 
	,\labels[1].label[113] ,\labels[1].label[112] ,\labels[1].label[111] 
	,\labels[1].label[110] ,\labels[1].label[109] ,\labels[1].label[108] 
	,\labels[1].label[107] ,\labels[1].label[106] ,\labels[1].label[105] 
	,\labels[1].label[104] ,\labels[1].label[103] ,\labels[1].label[102] 
	,\labels[1].label[101] ,\labels[1].label[100] ,\labels[1].label[99] 
	,\labels[1].label[98] ,\labels[1].label[97] ,\labels[1].label[96] 
	,\labels[1].label[95] ,\labels[1].label[94] ,\labels[1].label[93] 
	,\labels[1].label[92] ,\labels[1].label[91] ,\labels[1].label[90] 
	,\labels[1].label[89] ,\labels[1].label[88] ,\labels[1].label[87] 
	,\labels[1].label[86] ,\labels[1].label[85] ,\labels[1].label[84] 
	,\labels[1].label[83] ,\labels[1].label[82] ,\labels[1].label[81] 
	,\labels[1].label[80] ,\labels[1].label[79] ,\labels[1].label[78] 
	,\labels[1].label[77] ,\labels[1].label[76] ,\labels[1].label[75] 
	,\labels[1].label[74] ,\labels[1].label[73] ,\labels[1].label[72] 
	,\labels[1].label[71] ,\labels[1].label[70] ,\labels[1].label[69] 
	,\labels[1].label[68] ,\labels[1].label[67] ,\labels[1].label[66] 
	,\labels[1].label[65] ,\labels[1].label[64] ,\labels[1].label[63] 
	,\labels[1].label[62] ,\labels[1].label[61] ,\labels[1].label[60] 
	,\labels[1].label[59] ,\labels[1].label[58] ,\labels[1].label[57] 
	,\labels[1].label[56] ,\labels[1].label[55] ,\labels[1].label[54] 
	,\labels[1].label[53] ,\labels[1].label[52] ,\labels[1].label[51] 
	,\labels[1].label[50] ,\labels[1].label[49] ,\labels[1].label[48] 
	,\labels[1].label[47] ,\labels[1].label[46] ,\labels[1].label[45] 
	,\labels[1].label[44] ,\labels[1].label[43] ,\labels[1].label[42] 
	,\labels[1].label[41] ,\labels[1].label[40] ,\labels[1].label[39] 
	,\labels[1].label[38] ,\labels[1].label[37] ,\labels[1].label[36] 
	,\labels[1].label[35] ,\labels[1].label[34] ,\labels[1].label[33] 
	,\labels[1].label[32] ,\labels[1].label[31] ,\labels[1].label[30] 
	,\labels[1].label[29] ,\labels[1].label[28] ,\labels[1].label[27] 
	,\labels[1].label[26] ,\labels[1].label[25] ,\labels[1].label[24] 
	,\labels[1].label[23] ,\labels[1].label[22] ,\labels[1].label[21] 
	,\labels[1].label[20] ,\labels[1].label[19] ,\labels[1].label[18] 
	,\labels[1].label[17] ,\labels[1].label[16] ,\labels[1].label[15] 
	,\labels[1].label[14] ,\labels[1].label[13] ,\labels[1].label[12] 
	,\labels[1].label[11] ,\labels[1].label[10] ,\labels[1].label[9] 
	,\labels[1].label[8] ,\labels[1].label[7] ,\labels[1].label[6] 
	,\labels[1].label[5] ,\labels[1].label[4] ,\labels[1].label[3] 
	,\labels[1].label[2] ,\labels[1].label[1] ,\labels[1].label[0] 
	,\labels[1].delimiter_valid[0] ,\labels[1].delimiter[7] 
	,\labels[1].delimiter[6] ,\labels[1].delimiter[5] 
	,\labels[1].delimiter[4] ,\labels[1].delimiter[3] 
	,\labels[1].delimiter[2] ,\labels[1].delimiter[1] 
	,\labels[1].delimiter[0] ,\labels[0].guid_size[0] 
	,\labels[0].label_size[5] ,\labels[0].label_size[4] 
	,\labels[0].label_size[3] ,\labels[0].label_size[2] 
	,\labels[0].label_size[1] ,\labels[0].label_size[0] 
	,\labels[0].label[255] ,\labels[0].label[254] ,\labels[0].label[253] 
	,\labels[0].label[252] ,\labels[0].label[251] ,\labels[0].label[250] 
	,\labels[0].label[249] ,\labels[0].label[248] ,\labels[0].label[247] 
	,\labels[0].label[246] ,\labels[0].label[245] ,\labels[0].label[244] 
	,\labels[0].label[243] ,\labels[0].label[242] ,\labels[0].label[241] 
	,\labels[0].label[240] ,\labels[0].label[239] ,\labels[0].label[238] 
	,\labels[0].label[237] ,\labels[0].label[236] ,\labels[0].label[235] 
	,\labels[0].label[234] ,\labels[0].label[233] ,\labels[0].label[232] 
	,\labels[0].label[231] ,\labels[0].label[230] ,\labels[0].label[229] 
	,\labels[0].label[228] ,\labels[0].label[227] ,\labels[0].label[226] 
	,\labels[0].label[225] ,\labels[0].label[224] ,\labels[0].label[223] 
	,\labels[0].label[222] ,\labels[0].label[221] ,\labels[0].label[220] 
	,\labels[0].label[219] ,\labels[0].label[218] ,\labels[0].label[217] 
	,\labels[0].label[216] ,\labels[0].label[215] ,\labels[0].label[214] 
	,\labels[0].label[213] ,\labels[0].label[212] ,\labels[0].label[211] 
	,\labels[0].label[210] ,\labels[0].label[209] ,\labels[0].label[208] 
	,\labels[0].label[207] ,\labels[0].label[206] ,\labels[0].label[205] 
	,\labels[0].label[204] ,\labels[0].label[203] ,\labels[0].label[202] 
	,\labels[0].label[201] ,\labels[0].label[200] ,\labels[0].label[199] 
	,\labels[0].label[198] ,\labels[0].label[197] ,\labels[0].label[196] 
	,\labels[0].label[195] ,\labels[0].label[194] ,\labels[0].label[193] 
	,\labels[0].label[192] ,\labels[0].label[191] ,\labels[0].label[190] 
	,\labels[0].label[189] ,\labels[0].label[188] ,\labels[0].label[187] 
	,\labels[0].label[186] ,\labels[0].label[185] ,\labels[0].label[184] 
	,\labels[0].label[183] ,\labels[0].label[182] ,\labels[0].label[181] 
	,\labels[0].label[180] ,\labels[0].label[179] ,\labels[0].label[178] 
	,\labels[0].label[177] ,\labels[0].label[176] ,\labels[0].label[175] 
	,\labels[0].label[174] ,\labels[0].label[173] ,\labels[0].label[172] 
	,\labels[0].label[171] ,\labels[0].label[170] ,\labels[0].label[169] 
	,\labels[0].label[168] ,\labels[0].label[167] ,\labels[0].label[166] 
	,\labels[0].label[165] ,\labels[0].label[164] ,\labels[0].label[163] 
	,\labels[0].label[162] ,\labels[0].label[161] ,\labels[0].label[160] 
	,\labels[0].label[159] ,\labels[0].label[158] ,\labels[0].label[157] 
	,\labels[0].label[156] ,\labels[0].label[155] ,\labels[0].label[154] 
	,\labels[0].label[153] ,\labels[0].label[152] ,\labels[0].label[151] 
	,\labels[0].label[150] ,\labels[0].label[149] ,\labels[0].label[148] 
	,\labels[0].label[147] ,\labels[0].label[146] ,\labels[0].label[145] 
	,\labels[0].label[144] ,\labels[0].label[143] ,\labels[0].label[142] 
	,\labels[0].label[141] ,\labels[0].label[140] ,\labels[0].label[139] 
	,\labels[0].label[138] ,\labels[0].label[137] ,\labels[0].label[136] 
	,\labels[0].label[135] ,\labels[0].label[134] ,\labels[0].label[133] 
	,\labels[0].label[132] ,\labels[0].label[131] ,\labels[0].label[130] 
	,\labels[0].label[129] ,\labels[0].label[128] ,\labels[0].label[127] 
	,\labels[0].label[126] ,\labels[0].label[125] ,\labels[0].label[124] 
	,\labels[0].label[123] ,\labels[0].label[122] ,\labels[0].label[121] 
	,\labels[0].label[120] ,\labels[0].label[119] ,\labels[0].label[118] 
	,\labels[0].label[117] ,\labels[0].label[116] ,\labels[0].label[115] 
	,\labels[0].label[114] ,\labels[0].label[113] ,\labels[0].label[112] 
	,\labels[0].label[111] ,\labels[0].label[110] ,\labels[0].label[109] 
	,\labels[0].label[108] ,\labels[0].label[107] ,\labels[0].label[106] 
	,\labels[0].label[105] ,\labels[0].label[104] ,\labels[0].label[103] 
	,\labels[0].label[102] ,\labels[0].label[101] ,\labels[0].label[100] 
	,\labels[0].label[99] ,\labels[0].label[98] ,\labels[0].label[97] 
	,\labels[0].label[96] ,\labels[0].label[95] ,\labels[0].label[94] 
	,\labels[0].label[93] ,\labels[0].label[92] ,\labels[0].label[91] 
	,\labels[0].label[90] ,\labels[0].label[89] ,\labels[0].label[88] 
	,\labels[0].label[87] ,\labels[0].label[86] ,\labels[0].label[85] 
	,\labels[0].label[84] ,\labels[0].label[83] ,\labels[0].label[82] 
	,\labels[0].label[81] ,\labels[0].label[80] ,\labels[0].label[79] 
	,\labels[0].label[78] ,\labels[0].label[77] ,\labels[0].label[76] 
	,\labels[0].label[75] ,\labels[0].label[74] ,\labels[0].label[73] 
	,\labels[0].label[72] ,\labels[0].label[71] ,\labels[0].label[70] 
	,\labels[0].label[69] ,\labels[0].label[68] ,\labels[0].label[67] 
	,\labels[0].label[66] ,\labels[0].label[65] ,\labels[0].label[64] 
	,\labels[0].label[63] ,\labels[0].label[62] ,\labels[0].label[61] 
	,\labels[0].label[60] ,\labels[0].label[59] ,\labels[0].label[58] 
	,\labels[0].label[57] ,\labels[0].label[56] ,\labels[0].label[55] 
	,\labels[0].label[54] ,\labels[0].label[53] ,\labels[0].label[52] 
	,\labels[0].label[51] ,\labels[0].label[50] ,\labels[0].label[49] 
	,\labels[0].label[48] ,\labels[0].label[47] ,\labels[0].label[46] 
	,\labels[0].label[45] ,\labels[0].label[44] ,\labels[0].label[43] 
	,\labels[0].label[42] ,\labels[0].label[41] ,\labels[0].label[40] 
	,\labels[0].label[39] ,\labels[0].label[38] ,\labels[0].label[37] 
	,\labels[0].label[36] ,\labels[0].label[35] ,\labels[0].label[34] 
	,\labels[0].label[33] ,\labels[0].label[32] ,\labels[0].label[31] 
	,\labels[0].label[30] ,\labels[0].label[29] ,\labels[0].label[28] 
	,\labels[0].label[27] ,\labels[0].label[26] ,\labels[0].label[25] 
	,\labels[0].label[24] ,\labels[0].label[23] ,\labels[0].label[22] 
	,\labels[0].label[21] ,\labels[0].label[20] ,\labels[0].label[19] 
	,\labels[0].label[18] ,\labels[0].label[17] ,\labels[0].label[16] 
	,\labels[0].label[15] ,\labels[0].label[14] ,\labels[0].label[13] 
	,\labels[0].label[12] ,\labels[0].label[11] ,\labels[0].label[10] 
	,\labels[0].label[9] ,\labels[0].label[8] ,\labels[0].label[7] 
	,\labels[0].label[6] ,\labels[0].label[5] ,\labels[0].label[4] 
	,\labels[0].label[3] ,\labels[0].label[2] ,\labels[0].label[1] 
	,\labels[0].label[0] ,\labels[0].delimiter_valid[0] 
	,\labels[0].delimiter[7] ,\labels[0].delimiter[6] 
	,\labels[0].delimiter[5] ,\labels[0].delimiter[4] 
	,\labels[0].delimiter[3] ,\labels[0].delimiter[2] 
	,\labels[0].delimiter[1] ,\labels[0].delimiter[0] ;
input [0:0] \kme_internal_out.sot ;
input [0:0] \kme_internal_out.eoi ;
input [0:0] \kme_internal_out.eot ;
input [3:0] \kme_internal_out.id ;
input [63:0] \kme_internal_out.tdata ;
wire [70:0] kme_internal_out;
input kme_internal_out_valid;
input gcm_cmd_in_stall;
input gcm_tag_data_in_stall;
input upsizer_inspector_stall;
input keyfilter_cmd_in_stall;
input kdfstream_cmd_in_stall;
input kdf_cmd_in_stall;
input tlv_sb_data_in_stall;
wire _zy_simnet_kme_internal_out_ack_0_w$;
wire [0:610] _zy_simnet_gcm_cmd_in_1_w$;
wire _zy_simnet_gcm_cmd_in_valid_2_w$;
wire [0:95] _zy_simnet_gcm_tag_data_in_3_w$;
wire _zy_simnet_gcm_tag_data_in_valid_4_w$;
wire _zy_simnet_inspector_upsizer_valid_5_w$;
wire _zy_simnet_inspector_upsizer_eof_6_w$;
wire [0:63] _zy_simnet_inspector_upsizer_data_7_w$;
wire _zy_simnet_keyfilter_cmd_in_8_w$;
wire _zy_simnet_keyfilter_cmd_in_valid_9_w$;
wire [0:262] _zy_simnet_kdfstream_cmd_in_10_w$;
wire _zy_simnet_kdfstream_cmd_in_valid_11_w$;
wire [0:3] _zy_simnet_kdf_cmd_in_12_w$;
wire _zy_simnet_kdf_cmd_in_valid_13_w$;
wire [0:63] _zy_simnet_tlv_sb_data_in_14_w$;
wire _zy_simnet_tlv_sb_data_in_valid_15_w$;
wire _zy_sva_brcm_gcm_dek256_with_512bit_key_1_reset_or;
wire _zy_sva_brcm_gcm_dek512_with_512bit_key_2_reset_or;
wire _zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_reset_or;
wire _zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_reset_or;
wire _zy_sva_brcm_gcm_enc_dek256_no_kbk_5_reset_or;
wire _zy_sva_brcm_gcm_enc_dek512_no_kbk_6_reset_or;
wire _zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_reset_or;
wire _zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_reset_or;
wire _zy_sva_brcm_tlv_sb_stall_on_guid_9_reset_or;
wire _zy_sva_brcm_gcm_10_reset_or;
wire _zy_sva_brcm_gcm_11_reset_or;
wire _zy_sva_brcm_gcm_12_reset_or;
wire _zy_sva_brcm_gcm_13_reset_or;
wire _zy_sva_brcm_gcm_14_reset_or;
wire _zy_sva_brcm_gcm_15_reset_or;
wire _zy_sva_brcm_gcm_16_reset_or;
wire _zy_sva_brcm_gcm_17_reset_or;
wire _zy_sva_brcm_kdf_label0_8_18_reset_or;
wire _zy_sva_brcm_kdf_label9_16_19_reset_or;
wire _zy_sva_brcm_kdf_label17_24_20_reset_or;
wire _zy_sva_brcm_kdf_label25_32_21_reset_or;
wire _zy_sva_brcm_kdf_label0_8_22_reset_or;
wire _zy_sva_brcm_kdf_label9_16_23_reset_or;
wire _zy_sva_brcm_kdf_label17_24_24_reset_or;
wire _zy_sva_brcm_kdf_label25_32_25_reset_or;
wire _zy_sva_brcm_kdf_label0_8_26_reset_or;
wire _zy_sva_brcm_kdf_label9_16_27_reset_or;
wire _zy_sva_brcm_kdf_label17_24_28_reset_or;
wire _zy_sva_brcm_kdf_label25_32_29_reset_or;
wire _zy_sva_brcm_kdf_label0_8_30_reset_or;
wire _zy_sva_brcm_kdf_label9_16_31_reset_or;
wire _zy_sva_brcm_kdf_label17_24_32_reset_or;
wire _zy_sva_brcm_kdf_label25_32_33_reset_or;
wire _zy_sva_b0_t;
wire _zy_sva_b1_t;
wire _zy_sva_b2_t;
wire _zy_sva_b3_t;
wire _zy_sva_b4_t;
wire _zy_sva_b5_t;
wire _zy_sva_b6_t;
wire _zy_sva_b7_t;
wire _zy_sva_b8_t;
wire _zy_sva_b9_t;
wire _zy_sva_b10_t;
wire _zy_sva_b11_t;
wire _zy_sva_b12_t;
wire _zy_sva_b13_t;
wire _zy_sva_b14_t;
wire _zy_sva_b15_t;
wire _zy_sva_b16_t;
wire _zy_sva_b17_t;
wire _zy_sva_b18_t;
wire _zy_sva_b19_t;
wire _zy_sva_b20_t;
wire _zy_sva_b21_t;
wire _zy_sva_b22_t;
wire _zy_sva_b23_t;
wire _zy_sva_b24_t;
wire _zy_sva_b25_t;
wire _zy_sva_b26_t;
wire _zy_sva_b27_t;
wire _zy_sva_b28_t;
wire _zy_sva_b29_t;
wire _zy_sva_b30_t;
wire _zy_sva_b31_t;
wire _zy_sva_b32_t;
wire [31:0] debug_cmd;
wire [63:0] int_tlv_word0;
wire [63:0] int_tlv_word8;
wire [63:0] int_tlv_word9;
wire [55:0] int_tlv_word42;
wire [31:0] key_header;
wire [262:0] stream_cmd_in;
wire [262:0] stream_cmd_in_nxt;
wire [610:0] gcm_dek_cmd_in;
wire [610:0] gcm_dek_cmd_in_nxt;
wire [610:0] gcm_dak_cmd_in;
wire [610:0] gcm_dak_cmd_in_nxt;
wire skip_dek_kdf;
wire skip_dek_kdf_nxt;
wire skip_dak_kdf;
wire skip_dak_kdf_nxt;
wire [95:0] gcm_dek_tag;
wire [95:0] gcm_dek_tag_nxt;
wire [95:0] gcm_dak_tag;
wire [95:0] gcm_dak_tag_nxt;
wire corrupt_kme_error_bit_0;
wire rst_corrupt_kme_error_bit_0;
wire corrupt_crc32;
wire rst_corrupt_crc32;
wire kdf_dek_iter_nxt;
wire kdf_dek_iter;
wire [1:0] dek_ckv_length_q;
wire kek_tag_q;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek256_with_512bit_key_1_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek256_with_512bit_key_1_cpass;
`_2_ wire _zy_sva_b0;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek512_with_512bit_key_2_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek512_with_512bit_key_2_cpass;
`_2_ wire _zy_sva_b1;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_cpass;
`_2_ wire _zy_sva_b2;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_cpass;
`_2_ wire _zy_sva_b3;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek256_no_kbk_5_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek256_no_kbk_5_cpass;
`_2_ wire _zy_sva_b4;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek512_no_kbk_6_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek512_no_kbk_6_cpass;
`_2_ wire _zy_sva_b5;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_cpass;
`_2_ wire _zy_sva_b6;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_cpass;
`_2_ wire _zy_sva_b7;
`_2_ wire [0:0] _zy_sva_brcm_tlv_sb_stall_on_guid_9_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_tlv_sb_stall_on_guid_9_cpass;
`_2_ wire _zy_sva_b8;
`_2_ wire [0:0] _zy_sva_brcm_gcm_10_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_10_cpass;
`_2_ wire _zy_sva_b9;
`_2_ wire [0:0] _zy_sva_brcm_gcm_11_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_11_cpass;
`_2_ wire _zy_sva_b10;
`_2_ wire [0:0] _zy_sva_brcm_gcm_12_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_12_cpass;
`_2_ wire _zy_sva_b11;
`_2_ wire [0:0] _zy_sva_brcm_gcm_13_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_13_cpass;
`_2_ wire _zy_sva_b12;
`_2_ wire [0:0] _zy_sva_brcm_gcm_14_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_14_cpass;
`_2_ wire _zy_sva_b13;
`_2_ wire [0:0] _zy_sva_brcm_gcm_15_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_15_cpass;
`_2_ wire _zy_sva_b14;
`_2_ wire [0:0] _zy_sva_brcm_gcm_16_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_16_cpass;
`_2_ wire _zy_sva_b15;
`_2_ wire [0:0] _zy_sva_brcm_gcm_17_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_gcm_17_cpass;
`_2_ wire _zy_sva_b16;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_18_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_18_cpass;
`_2_ wire _zy_sva_b17;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_19_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_19_cpass;
`_2_ wire _zy_sva_b18;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_20_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_20_cpass;
`_2_ wire _zy_sva_b19;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_21_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_21_cpass;
`_2_ wire _zy_sva_b20;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_22_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_22_cpass;
`_2_ wire _zy_sva_b21;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_23_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_23_cpass;
`_2_ wire _zy_sva_b22;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_24_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_24_cpass;
`_2_ wire _zy_sva_b23;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_25_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_25_cpass;
`_2_ wire _zy_sva_b24;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_26_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_26_cpass;
`_2_ wire _zy_sva_b25;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_27_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_27_cpass;
`_2_ wire _zy_sva_b26;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_28_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_28_cpass;
`_2_ wire _zy_sva_b27;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_29_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_29_cpass;
`_2_ wire _zy_sva_b28;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_30_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label0_8_30_cpass;
`_2_ wire _zy_sva_b29;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_31_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label9_16_31_cpass;
`_2_ wire _zy_sva_b30;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_32_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label17_24_32_cpass;
`_2_ wire _zy_sva_b31;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_33_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_kdf_label25_32_33_cpass;
`_2_ wire _zy_sva_b32;
supply1 n2850;
supply0 n2851;
wire [0:0] \debug_cmd.tlvp_corrupt ;
wire [1:0] \debug_cmd.cmd_mode ;
wire [4:0] \debug_cmd.module_id ;
wire [0:0] \debug_cmd.cmd_type ;
wire [4:0] \debug_cmd.tlv_num ;
wire [9:0] \debug_cmd.byte_num ;
wire [7:0] \debug_cmd.byte_msk ;
wire [1:0] \int_tlv_word0.tlv_bip2 ;
wire [12:0] \int_tlv_word0.resv0 ;
wire [0:0] \int_tlv_word0.kdf_dek_iter ;
wire [0:0] \int_tlv_word0.keyless_algos ;
wire [0:0] \int_tlv_word0.needs_dek ;
wire [0:0] \int_tlv_word0.needs_dak ;
wire [5:0] \int_tlv_word0.key_type ;
wire [10:0] \int_tlv_word0.tlv_frame_num ;
wire [3:0] \int_tlv_word0.tlv_eng_id ;
wire [7:0] \int_tlv_word0.tlv_seq_num ;
wire [7:0] \int_tlv_word0.tlv_len ;
wire [7:0] \int_tlv_word0.tlv_type ;
wire [0:0] \int_tlv_word8.dek_kim_entry.valid ;
wire [2:0] \int_tlv_word8.dek_kim_entry.label_index ;
wire [1:0] \int_tlv_word8.dek_kim_entry.ckv_length ;
wire [14:0] \int_tlv_word8.dek_kim_entry.ckv_pointer ;
wire [3:0] \int_tlv_word8.dek_kim_entry.pf_num ;
wire [11:0] \int_tlv_word8.dek_kim_entry.vf_num ;
wire [0:0] \int_tlv_word8.dek_kim_entry.vf_valid ;
wire [5:0] \int_tlv_word8.unused ;
wire [0:0] \int_tlv_word8.missing_iv ;
wire [0:0] \int_tlv_word8.missing_guid ;
wire [0:0] \int_tlv_word8.validate_dek ;
wire [0:0] \int_tlv_word8.vf_valid ;
wire [3:0] \int_tlv_word8.pf_num ;
wire [11:0] \int_tlv_word8.vf_num ;
wire [0:0] \int_tlv_word9.dak_kim_entry.valid ;
wire [2:0] \int_tlv_word9.dak_kim_entry.label_index ;
wire [1:0] \int_tlv_word9.dak_kim_entry.ckv_length ;
wire [14:0] \int_tlv_word9.dak_kim_entry.ckv_pointer ;
wire [3:0] \int_tlv_word9.dak_kim_entry.pf_num ;
wire [11:0] \int_tlv_word9.dak_kim_entry.vf_num ;
wire [0:0] \int_tlv_word9.dak_kim_entry.vf_valid ;
wire [7:0] \int_tlv_word9.unused ;
wire [0:0] \int_tlv_word9.validate_dak ;
wire [0:0] \int_tlv_word9.vf_valid ;
wire [3:0] \int_tlv_word9.pf_num ;
wire [11:0] \int_tlv_word9.vf_num ;
wire [0:0] \int_tlv_word42.corrupt_crc32 ;
wire [46:0] \int_tlv_word42.unused ;
wire [7:0] \int_tlv_word42.error_code ;
wire [0:0] \key_header.dak_key_op ;
wire [13:0] \key_header.dak_key_ref ;
wire [1:0] \key_header.kdf_mode ;
wire [0:0] \key_header.dek_key_op ;
wire [13:0] \key_header.dek_key_ref ;
wire [0:0] \stream_cmd_in.combo_mode ;
wire [0:0] \stream_cmd_in.skip ;
wire [255:0] \stream_cmd_in.guid ;
wire [2:0] \stream_cmd_in.label_index ;
wire [1:0] \stream_cmd_in.num_iter ;
wire [0:0] \stream_cmd_in_nxt.combo_mode ;
wire [0:0] \stream_cmd_in_nxt.skip ;
wire [255:0] \stream_cmd_in_nxt.guid ;
wire [2:0] \stream_cmd_in_nxt.label_index ;
wire [1:0] \stream_cmd_in_nxt.num_iter ;
wire [255:0] \gcm_dek_cmd_in.key0 ;
wire [255:0] \gcm_dek_cmd_in.key1 ;
wire [95:0] \gcm_dek_cmd_in.iv ;
wire [2:0] \gcm_dek_cmd_in.op ;
wire [255:0] \gcm_dek_cmd_in_nxt.key0 ;
wire [255:0] \gcm_dek_cmd_in_nxt.key1 ;
wire [95:0] \gcm_dek_cmd_in_nxt.iv ;
wire [2:0] \gcm_dek_cmd_in_nxt.op ;
wire [255:0] \gcm_dak_cmd_in.key0 ;
wire [255:0] \gcm_dak_cmd_in.key1 ;
wire [95:0] \gcm_dak_cmd_in.iv ;
wire [2:0] \gcm_dak_cmd_in.op ;
wire [255:0] \gcm_dak_cmd_in_nxt.key0 ;
wire [255:0] \gcm_dak_cmd_in_nxt.key1 ;
wire [95:0] \gcm_dak_cmd_in_nxt.iv ;
wire [2:0] \gcm_dak_cmd_in_nxt.op ;
tran (gcm_cmd_in[610], \gcm_cmd_in.key0 [255]);
tran (gcm_cmd_in[609], \gcm_cmd_in.key0 [254]);
tran (gcm_cmd_in[608], \gcm_cmd_in.key0 [253]);
tran (gcm_cmd_in[607], \gcm_cmd_in.key0 [252]);
tran (gcm_cmd_in[606], \gcm_cmd_in.key0 [251]);
tran (gcm_cmd_in[605], \gcm_cmd_in.key0 [250]);
tran (gcm_cmd_in[604], \gcm_cmd_in.key0 [249]);
tran (gcm_cmd_in[603], \gcm_cmd_in.key0 [248]);
tran (gcm_cmd_in[602], \gcm_cmd_in.key0 [247]);
tran (gcm_cmd_in[601], \gcm_cmd_in.key0 [246]);
tran (gcm_cmd_in[600], \gcm_cmd_in.key0 [245]);
tran (gcm_cmd_in[599], \gcm_cmd_in.key0 [244]);
tran (gcm_cmd_in[598], \gcm_cmd_in.key0 [243]);
tran (gcm_cmd_in[597], \gcm_cmd_in.key0 [242]);
tran (gcm_cmd_in[596], \gcm_cmd_in.key0 [241]);
tran (gcm_cmd_in[595], \gcm_cmd_in.key0 [240]);
tran (gcm_cmd_in[594], \gcm_cmd_in.key0 [239]);
tran (gcm_cmd_in[593], \gcm_cmd_in.key0 [238]);
tran (gcm_cmd_in[592], \gcm_cmd_in.key0 [237]);
tran (gcm_cmd_in[591], \gcm_cmd_in.key0 [236]);
tran (gcm_cmd_in[590], \gcm_cmd_in.key0 [235]);
tran (gcm_cmd_in[589], \gcm_cmd_in.key0 [234]);
tran (gcm_cmd_in[588], \gcm_cmd_in.key0 [233]);
tran (gcm_cmd_in[587], \gcm_cmd_in.key0 [232]);
tran (gcm_cmd_in[586], \gcm_cmd_in.key0 [231]);
tran (gcm_cmd_in[585], \gcm_cmd_in.key0 [230]);
tran (gcm_cmd_in[584], \gcm_cmd_in.key0 [229]);
tran (gcm_cmd_in[583], \gcm_cmd_in.key0 [228]);
tran (gcm_cmd_in[582], \gcm_cmd_in.key0 [227]);
tran (gcm_cmd_in[581], \gcm_cmd_in.key0 [226]);
tran (gcm_cmd_in[580], \gcm_cmd_in.key0 [225]);
tran (gcm_cmd_in[579], \gcm_cmd_in.key0 [224]);
tran (gcm_cmd_in[578], \gcm_cmd_in.key0 [223]);
tran (gcm_cmd_in[577], \gcm_cmd_in.key0 [222]);
tran (gcm_cmd_in[576], \gcm_cmd_in.key0 [221]);
tran (gcm_cmd_in[575], \gcm_cmd_in.key0 [220]);
tran (gcm_cmd_in[574], \gcm_cmd_in.key0 [219]);
tran (gcm_cmd_in[573], \gcm_cmd_in.key0 [218]);
tran (gcm_cmd_in[572], \gcm_cmd_in.key0 [217]);
tran (gcm_cmd_in[571], \gcm_cmd_in.key0 [216]);
tran (gcm_cmd_in[570], \gcm_cmd_in.key0 [215]);
tran (gcm_cmd_in[569], \gcm_cmd_in.key0 [214]);
tran (gcm_cmd_in[568], \gcm_cmd_in.key0 [213]);
tran (gcm_cmd_in[567], \gcm_cmd_in.key0 [212]);
tran (gcm_cmd_in[566], \gcm_cmd_in.key0 [211]);
tran (gcm_cmd_in[565], \gcm_cmd_in.key0 [210]);
tran (gcm_cmd_in[564], \gcm_cmd_in.key0 [209]);
tran (gcm_cmd_in[563], \gcm_cmd_in.key0 [208]);
tran (gcm_cmd_in[562], \gcm_cmd_in.key0 [207]);
tran (gcm_cmd_in[561], \gcm_cmd_in.key0 [206]);
tran (gcm_cmd_in[560], \gcm_cmd_in.key0 [205]);
tran (gcm_cmd_in[559], \gcm_cmd_in.key0 [204]);
tran (gcm_cmd_in[558], \gcm_cmd_in.key0 [203]);
tran (gcm_cmd_in[557], \gcm_cmd_in.key0 [202]);
tran (gcm_cmd_in[556], \gcm_cmd_in.key0 [201]);
tran (gcm_cmd_in[555], \gcm_cmd_in.key0 [200]);
tran (gcm_cmd_in[554], \gcm_cmd_in.key0 [199]);
tran (gcm_cmd_in[553], \gcm_cmd_in.key0 [198]);
tran (gcm_cmd_in[552], \gcm_cmd_in.key0 [197]);
tran (gcm_cmd_in[551], \gcm_cmd_in.key0 [196]);
tran (gcm_cmd_in[550], \gcm_cmd_in.key0 [195]);
tran (gcm_cmd_in[549], \gcm_cmd_in.key0 [194]);
tran (gcm_cmd_in[548], \gcm_cmd_in.key0 [193]);
tran (gcm_cmd_in[547], \gcm_cmd_in.key0 [192]);
tran (gcm_cmd_in[546], \gcm_cmd_in.key0 [191]);
tran (gcm_cmd_in[545], \gcm_cmd_in.key0 [190]);
tran (gcm_cmd_in[544], \gcm_cmd_in.key0 [189]);
tran (gcm_cmd_in[543], \gcm_cmd_in.key0 [188]);
tran (gcm_cmd_in[542], \gcm_cmd_in.key0 [187]);
tran (gcm_cmd_in[541], \gcm_cmd_in.key0 [186]);
tran (gcm_cmd_in[540], \gcm_cmd_in.key0 [185]);
tran (gcm_cmd_in[539], \gcm_cmd_in.key0 [184]);
tran (gcm_cmd_in[538], \gcm_cmd_in.key0 [183]);
tran (gcm_cmd_in[537], \gcm_cmd_in.key0 [182]);
tran (gcm_cmd_in[536], \gcm_cmd_in.key0 [181]);
tran (gcm_cmd_in[535], \gcm_cmd_in.key0 [180]);
tran (gcm_cmd_in[534], \gcm_cmd_in.key0 [179]);
tran (gcm_cmd_in[533], \gcm_cmd_in.key0 [178]);
tran (gcm_cmd_in[532], \gcm_cmd_in.key0 [177]);
tran (gcm_cmd_in[531], \gcm_cmd_in.key0 [176]);
tran (gcm_cmd_in[530], \gcm_cmd_in.key0 [175]);
tran (gcm_cmd_in[529], \gcm_cmd_in.key0 [174]);
tran (gcm_cmd_in[528], \gcm_cmd_in.key0 [173]);
tran (gcm_cmd_in[527], \gcm_cmd_in.key0 [172]);
tran (gcm_cmd_in[526], \gcm_cmd_in.key0 [171]);
tran (gcm_cmd_in[525], \gcm_cmd_in.key0 [170]);
tran (gcm_cmd_in[524], \gcm_cmd_in.key0 [169]);
tran (gcm_cmd_in[523], \gcm_cmd_in.key0 [168]);
tran (gcm_cmd_in[522], \gcm_cmd_in.key0 [167]);
tran (gcm_cmd_in[521], \gcm_cmd_in.key0 [166]);
tran (gcm_cmd_in[520], \gcm_cmd_in.key0 [165]);
tran (gcm_cmd_in[519], \gcm_cmd_in.key0 [164]);
tran (gcm_cmd_in[518], \gcm_cmd_in.key0 [163]);
tran (gcm_cmd_in[517], \gcm_cmd_in.key0 [162]);
tran (gcm_cmd_in[516], \gcm_cmd_in.key0 [161]);
tran (gcm_cmd_in[515], \gcm_cmd_in.key0 [160]);
tran (gcm_cmd_in[514], \gcm_cmd_in.key0 [159]);
tran (gcm_cmd_in[513], \gcm_cmd_in.key0 [158]);
tran (gcm_cmd_in[512], \gcm_cmd_in.key0 [157]);
tran (gcm_cmd_in[511], \gcm_cmd_in.key0 [156]);
tran (gcm_cmd_in[510], \gcm_cmd_in.key0 [155]);
tran (gcm_cmd_in[509], \gcm_cmd_in.key0 [154]);
tran (gcm_cmd_in[508], \gcm_cmd_in.key0 [153]);
tran (gcm_cmd_in[507], \gcm_cmd_in.key0 [152]);
tran (gcm_cmd_in[506], \gcm_cmd_in.key0 [151]);
tran (gcm_cmd_in[505], \gcm_cmd_in.key0 [150]);
tran (gcm_cmd_in[504], \gcm_cmd_in.key0 [149]);
tran (gcm_cmd_in[503], \gcm_cmd_in.key0 [148]);
tran (gcm_cmd_in[502], \gcm_cmd_in.key0 [147]);
tran (gcm_cmd_in[501], \gcm_cmd_in.key0 [146]);
tran (gcm_cmd_in[500], \gcm_cmd_in.key0 [145]);
tran (gcm_cmd_in[499], \gcm_cmd_in.key0 [144]);
tran (gcm_cmd_in[498], \gcm_cmd_in.key0 [143]);
tran (gcm_cmd_in[497], \gcm_cmd_in.key0 [142]);
tran (gcm_cmd_in[496], \gcm_cmd_in.key0 [141]);
tran (gcm_cmd_in[495], \gcm_cmd_in.key0 [140]);
tran (gcm_cmd_in[494], \gcm_cmd_in.key0 [139]);
tran (gcm_cmd_in[493], \gcm_cmd_in.key0 [138]);
tran (gcm_cmd_in[492], \gcm_cmd_in.key0 [137]);
tran (gcm_cmd_in[491], \gcm_cmd_in.key0 [136]);
tran (gcm_cmd_in[490], \gcm_cmd_in.key0 [135]);
tran (gcm_cmd_in[489], \gcm_cmd_in.key0 [134]);
tran (gcm_cmd_in[488], \gcm_cmd_in.key0 [133]);
tran (gcm_cmd_in[487], \gcm_cmd_in.key0 [132]);
tran (gcm_cmd_in[486], \gcm_cmd_in.key0 [131]);
tran (gcm_cmd_in[485], \gcm_cmd_in.key0 [130]);
tran (gcm_cmd_in[484], \gcm_cmd_in.key0 [129]);
tran (gcm_cmd_in[483], \gcm_cmd_in.key0 [128]);
tran (gcm_cmd_in[482], \gcm_cmd_in.key0 [127]);
tran (gcm_cmd_in[481], \gcm_cmd_in.key0 [126]);
tran (gcm_cmd_in[480], \gcm_cmd_in.key0 [125]);
tran (gcm_cmd_in[479], \gcm_cmd_in.key0 [124]);
tran (gcm_cmd_in[478], \gcm_cmd_in.key0 [123]);
tran (gcm_cmd_in[477], \gcm_cmd_in.key0 [122]);
tran (gcm_cmd_in[476], \gcm_cmd_in.key0 [121]);
tran (gcm_cmd_in[475], \gcm_cmd_in.key0 [120]);
tran (gcm_cmd_in[474], \gcm_cmd_in.key0 [119]);
tran (gcm_cmd_in[473], \gcm_cmd_in.key0 [118]);
tran (gcm_cmd_in[472], \gcm_cmd_in.key0 [117]);
tran (gcm_cmd_in[471], \gcm_cmd_in.key0 [116]);
tran (gcm_cmd_in[470], \gcm_cmd_in.key0 [115]);
tran (gcm_cmd_in[469], \gcm_cmd_in.key0 [114]);
tran (gcm_cmd_in[468], \gcm_cmd_in.key0 [113]);
tran (gcm_cmd_in[467], \gcm_cmd_in.key0 [112]);
tran (gcm_cmd_in[466], \gcm_cmd_in.key0 [111]);
tran (gcm_cmd_in[465], \gcm_cmd_in.key0 [110]);
tran (gcm_cmd_in[464], \gcm_cmd_in.key0 [109]);
tran (gcm_cmd_in[463], \gcm_cmd_in.key0 [108]);
tran (gcm_cmd_in[462], \gcm_cmd_in.key0 [107]);
tran (gcm_cmd_in[461], \gcm_cmd_in.key0 [106]);
tran (gcm_cmd_in[460], \gcm_cmd_in.key0 [105]);
tran (gcm_cmd_in[459], \gcm_cmd_in.key0 [104]);
tran (gcm_cmd_in[458], \gcm_cmd_in.key0 [103]);
tran (gcm_cmd_in[457], \gcm_cmd_in.key0 [102]);
tran (gcm_cmd_in[456], \gcm_cmd_in.key0 [101]);
tran (gcm_cmd_in[455], \gcm_cmd_in.key0 [100]);
tran (gcm_cmd_in[454], \gcm_cmd_in.key0 [99]);
tran (gcm_cmd_in[453], \gcm_cmd_in.key0 [98]);
tran (gcm_cmd_in[452], \gcm_cmd_in.key0 [97]);
tran (gcm_cmd_in[451], \gcm_cmd_in.key0 [96]);
tran (gcm_cmd_in[450], \gcm_cmd_in.key0 [95]);
tran (gcm_cmd_in[449], \gcm_cmd_in.key0 [94]);
tran (gcm_cmd_in[448], \gcm_cmd_in.key0 [93]);
tran (gcm_cmd_in[447], \gcm_cmd_in.key0 [92]);
tran (gcm_cmd_in[446], \gcm_cmd_in.key0 [91]);
tran (gcm_cmd_in[445], \gcm_cmd_in.key0 [90]);
tran (gcm_cmd_in[444], \gcm_cmd_in.key0 [89]);
tran (gcm_cmd_in[443], \gcm_cmd_in.key0 [88]);
tran (gcm_cmd_in[442], \gcm_cmd_in.key0 [87]);
tran (gcm_cmd_in[441], \gcm_cmd_in.key0 [86]);
tran (gcm_cmd_in[440], \gcm_cmd_in.key0 [85]);
tran (gcm_cmd_in[439], \gcm_cmd_in.key0 [84]);
tran (gcm_cmd_in[438], \gcm_cmd_in.key0 [83]);
tran (gcm_cmd_in[437], \gcm_cmd_in.key0 [82]);
tran (gcm_cmd_in[436], \gcm_cmd_in.key0 [81]);
tran (gcm_cmd_in[435], \gcm_cmd_in.key0 [80]);
tran (gcm_cmd_in[434], \gcm_cmd_in.key0 [79]);
tran (gcm_cmd_in[433], \gcm_cmd_in.key0 [78]);
tran (gcm_cmd_in[432], \gcm_cmd_in.key0 [77]);
tran (gcm_cmd_in[431], \gcm_cmd_in.key0 [76]);
tran (gcm_cmd_in[430], \gcm_cmd_in.key0 [75]);
tran (gcm_cmd_in[429], \gcm_cmd_in.key0 [74]);
tran (gcm_cmd_in[428], \gcm_cmd_in.key0 [73]);
tran (gcm_cmd_in[427], \gcm_cmd_in.key0 [72]);
tran (gcm_cmd_in[426], \gcm_cmd_in.key0 [71]);
tran (gcm_cmd_in[425], \gcm_cmd_in.key0 [70]);
tran (gcm_cmd_in[424], \gcm_cmd_in.key0 [69]);
tran (gcm_cmd_in[423], \gcm_cmd_in.key0 [68]);
tran (gcm_cmd_in[422], \gcm_cmd_in.key0 [67]);
tran (gcm_cmd_in[421], \gcm_cmd_in.key0 [66]);
tran (gcm_cmd_in[420], \gcm_cmd_in.key0 [65]);
tran (gcm_cmd_in[419], \gcm_cmd_in.key0 [64]);
tran (gcm_cmd_in[418], \gcm_cmd_in.key0 [63]);
tran (gcm_cmd_in[417], \gcm_cmd_in.key0 [62]);
tran (gcm_cmd_in[416], \gcm_cmd_in.key0 [61]);
tran (gcm_cmd_in[415], \gcm_cmd_in.key0 [60]);
tran (gcm_cmd_in[414], \gcm_cmd_in.key0 [59]);
tran (gcm_cmd_in[413], \gcm_cmd_in.key0 [58]);
tran (gcm_cmd_in[412], \gcm_cmd_in.key0 [57]);
tran (gcm_cmd_in[411], \gcm_cmd_in.key0 [56]);
tran (gcm_cmd_in[410], \gcm_cmd_in.key0 [55]);
tran (gcm_cmd_in[409], \gcm_cmd_in.key0 [54]);
tran (gcm_cmd_in[408], \gcm_cmd_in.key0 [53]);
tran (gcm_cmd_in[407], \gcm_cmd_in.key0 [52]);
tran (gcm_cmd_in[406], \gcm_cmd_in.key0 [51]);
tran (gcm_cmd_in[405], \gcm_cmd_in.key0 [50]);
tran (gcm_cmd_in[404], \gcm_cmd_in.key0 [49]);
tran (gcm_cmd_in[403], \gcm_cmd_in.key0 [48]);
tran (gcm_cmd_in[402], \gcm_cmd_in.key0 [47]);
tran (gcm_cmd_in[401], \gcm_cmd_in.key0 [46]);
tran (gcm_cmd_in[400], \gcm_cmd_in.key0 [45]);
tran (gcm_cmd_in[399], \gcm_cmd_in.key0 [44]);
tran (gcm_cmd_in[398], \gcm_cmd_in.key0 [43]);
tran (gcm_cmd_in[397], \gcm_cmd_in.key0 [42]);
tran (gcm_cmd_in[396], \gcm_cmd_in.key0 [41]);
tran (gcm_cmd_in[395], \gcm_cmd_in.key0 [40]);
tran (gcm_cmd_in[394], \gcm_cmd_in.key0 [39]);
tran (gcm_cmd_in[393], \gcm_cmd_in.key0 [38]);
tran (gcm_cmd_in[392], \gcm_cmd_in.key0 [37]);
tran (gcm_cmd_in[391], \gcm_cmd_in.key0 [36]);
tran (gcm_cmd_in[390], \gcm_cmd_in.key0 [35]);
tran (gcm_cmd_in[389], \gcm_cmd_in.key0 [34]);
tran (gcm_cmd_in[388], \gcm_cmd_in.key0 [33]);
tran (gcm_cmd_in[387], \gcm_cmd_in.key0 [32]);
tran (gcm_cmd_in[386], \gcm_cmd_in.key0 [31]);
tran (gcm_cmd_in[385], \gcm_cmd_in.key0 [30]);
tran (gcm_cmd_in[384], \gcm_cmd_in.key0 [29]);
tran (gcm_cmd_in[383], \gcm_cmd_in.key0 [28]);
tran (gcm_cmd_in[382], \gcm_cmd_in.key0 [27]);
tran (gcm_cmd_in[381], \gcm_cmd_in.key0 [26]);
tran (gcm_cmd_in[380], \gcm_cmd_in.key0 [25]);
tran (gcm_cmd_in[379], \gcm_cmd_in.key0 [24]);
tran (gcm_cmd_in[378], \gcm_cmd_in.key0 [23]);
tran (gcm_cmd_in[377], \gcm_cmd_in.key0 [22]);
tran (gcm_cmd_in[376], \gcm_cmd_in.key0 [21]);
tran (gcm_cmd_in[375], \gcm_cmd_in.key0 [20]);
tran (gcm_cmd_in[374], \gcm_cmd_in.key0 [19]);
tran (gcm_cmd_in[373], \gcm_cmd_in.key0 [18]);
tran (gcm_cmd_in[372], \gcm_cmd_in.key0 [17]);
tran (gcm_cmd_in[371], \gcm_cmd_in.key0 [16]);
tran (gcm_cmd_in[370], \gcm_cmd_in.key0 [15]);
tran (gcm_cmd_in[369], \gcm_cmd_in.key0 [14]);
tran (gcm_cmd_in[368], \gcm_cmd_in.key0 [13]);
tran (gcm_cmd_in[367], \gcm_cmd_in.key0 [12]);
tran (gcm_cmd_in[366], \gcm_cmd_in.key0 [11]);
tran (gcm_cmd_in[365], \gcm_cmd_in.key0 [10]);
tran (gcm_cmd_in[364], \gcm_cmd_in.key0 [9]);
tran (gcm_cmd_in[363], \gcm_cmd_in.key0 [8]);
tran (gcm_cmd_in[362], \gcm_cmd_in.key0 [7]);
tran (gcm_cmd_in[361], \gcm_cmd_in.key0 [6]);
tran (gcm_cmd_in[360], \gcm_cmd_in.key0 [5]);
tran (gcm_cmd_in[359], \gcm_cmd_in.key0 [4]);
tran (gcm_cmd_in[358], \gcm_cmd_in.key0 [3]);
tran (gcm_cmd_in[357], \gcm_cmd_in.key0 [2]);
tran (gcm_cmd_in[356], \gcm_cmd_in.key0 [1]);
tran (gcm_cmd_in[355], \gcm_cmd_in.key0 [0]);
tran (gcm_cmd_in[354], \gcm_cmd_in.key1 [255]);
tran (gcm_cmd_in[353], \gcm_cmd_in.key1 [254]);
tran (gcm_cmd_in[352], \gcm_cmd_in.key1 [253]);
tran (gcm_cmd_in[351], \gcm_cmd_in.key1 [252]);
tran (gcm_cmd_in[350], \gcm_cmd_in.key1 [251]);
tran (gcm_cmd_in[349], \gcm_cmd_in.key1 [250]);
tran (gcm_cmd_in[348], \gcm_cmd_in.key1 [249]);
tran (gcm_cmd_in[347], \gcm_cmd_in.key1 [248]);
tran (gcm_cmd_in[346], \gcm_cmd_in.key1 [247]);
tran (gcm_cmd_in[345], \gcm_cmd_in.key1 [246]);
tran (gcm_cmd_in[344], \gcm_cmd_in.key1 [245]);
tran (gcm_cmd_in[343], \gcm_cmd_in.key1 [244]);
tran (gcm_cmd_in[342], \gcm_cmd_in.key1 [243]);
tran (gcm_cmd_in[341], \gcm_cmd_in.key1 [242]);
tran (gcm_cmd_in[340], \gcm_cmd_in.key1 [241]);
tran (gcm_cmd_in[339], \gcm_cmd_in.key1 [240]);
tran (gcm_cmd_in[338], \gcm_cmd_in.key1 [239]);
tran (gcm_cmd_in[337], \gcm_cmd_in.key1 [238]);
tran (gcm_cmd_in[336], \gcm_cmd_in.key1 [237]);
tran (gcm_cmd_in[335], \gcm_cmd_in.key1 [236]);
tran (gcm_cmd_in[334], \gcm_cmd_in.key1 [235]);
tran (gcm_cmd_in[333], \gcm_cmd_in.key1 [234]);
tran (gcm_cmd_in[332], \gcm_cmd_in.key1 [233]);
tran (gcm_cmd_in[331], \gcm_cmd_in.key1 [232]);
tran (gcm_cmd_in[330], \gcm_cmd_in.key1 [231]);
tran (gcm_cmd_in[329], \gcm_cmd_in.key1 [230]);
tran (gcm_cmd_in[328], \gcm_cmd_in.key1 [229]);
tran (gcm_cmd_in[327], \gcm_cmd_in.key1 [228]);
tran (gcm_cmd_in[326], \gcm_cmd_in.key1 [227]);
tran (gcm_cmd_in[325], \gcm_cmd_in.key1 [226]);
tran (gcm_cmd_in[324], \gcm_cmd_in.key1 [225]);
tran (gcm_cmd_in[323], \gcm_cmd_in.key1 [224]);
tran (gcm_cmd_in[322], \gcm_cmd_in.key1 [223]);
tran (gcm_cmd_in[321], \gcm_cmd_in.key1 [222]);
tran (gcm_cmd_in[320], \gcm_cmd_in.key1 [221]);
tran (gcm_cmd_in[319], \gcm_cmd_in.key1 [220]);
tran (gcm_cmd_in[318], \gcm_cmd_in.key1 [219]);
tran (gcm_cmd_in[317], \gcm_cmd_in.key1 [218]);
tran (gcm_cmd_in[316], \gcm_cmd_in.key1 [217]);
tran (gcm_cmd_in[315], \gcm_cmd_in.key1 [216]);
tran (gcm_cmd_in[314], \gcm_cmd_in.key1 [215]);
tran (gcm_cmd_in[313], \gcm_cmd_in.key1 [214]);
tran (gcm_cmd_in[312], \gcm_cmd_in.key1 [213]);
tran (gcm_cmd_in[311], \gcm_cmd_in.key1 [212]);
tran (gcm_cmd_in[310], \gcm_cmd_in.key1 [211]);
tran (gcm_cmd_in[309], \gcm_cmd_in.key1 [210]);
tran (gcm_cmd_in[308], \gcm_cmd_in.key1 [209]);
tran (gcm_cmd_in[307], \gcm_cmd_in.key1 [208]);
tran (gcm_cmd_in[306], \gcm_cmd_in.key1 [207]);
tran (gcm_cmd_in[305], \gcm_cmd_in.key1 [206]);
tran (gcm_cmd_in[304], \gcm_cmd_in.key1 [205]);
tran (gcm_cmd_in[303], \gcm_cmd_in.key1 [204]);
tran (gcm_cmd_in[302], \gcm_cmd_in.key1 [203]);
tran (gcm_cmd_in[301], \gcm_cmd_in.key1 [202]);
tran (gcm_cmd_in[300], \gcm_cmd_in.key1 [201]);
tran (gcm_cmd_in[299], \gcm_cmd_in.key1 [200]);
tran (gcm_cmd_in[298], \gcm_cmd_in.key1 [199]);
tran (gcm_cmd_in[297], \gcm_cmd_in.key1 [198]);
tran (gcm_cmd_in[296], \gcm_cmd_in.key1 [197]);
tran (gcm_cmd_in[295], \gcm_cmd_in.key1 [196]);
tran (gcm_cmd_in[294], \gcm_cmd_in.key1 [195]);
tran (gcm_cmd_in[293], \gcm_cmd_in.key1 [194]);
tran (gcm_cmd_in[292], \gcm_cmd_in.key1 [193]);
tran (gcm_cmd_in[291], \gcm_cmd_in.key1 [192]);
tran (gcm_cmd_in[290], \gcm_cmd_in.key1 [191]);
tran (gcm_cmd_in[289], \gcm_cmd_in.key1 [190]);
tran (gcm_cmd_in[288], \gcm_cmd_in.key1 [189]);
tran (gcm_cmd_in[287], \gcm_cmd_in.key1 [188]);
tran (gcm_cmd_in[286], \gcm_cmd_in.key1 [187]);
tran (gcm_cmd_in[285], \gcm_cmd_in.key1 [186]);
tran (gcm_cmd_in[284], \gcm_cmd_in.key1 [185]);
tran (gcm_cmd_in[283], \gcm_cmd_in.key1 [184]);
tran (gcm_cmd_in[282], \gcm_cmd_in.key1 [183]);
tran (gcm_cmd_in[281], \gcm_cmd_in.key1 [182]);
tran (gcm_cmd_in[280], \gcm_cmd_in.key1 [181]);
tran (gcm_cmd_in[279], \gcm_cmd_in.key1 [180]);
tran (gcm_cmd_in[278], \gcm_cmd_in.key1 [179]);
tran (gcm_cmd_in[277], \gcm_cmd_in.key1 [178]);
tran (gcm_cmd_in[276], \gcm_cmd_in.key1 [177]);
tran (gcm_cmd_in[275], \gcm_cmd_in.key1 [176]);
tran (gcm_cmd_in[274], \gcm_cmd_in.key1 [175]);
tran (gcm_cmd_in[273], \gcm_cmd_in.key1 [174]);
tran (gcm_cmd_in[272], \gcm_cmd_in.key1 [173]);
tran (gcm_cmd_in[271], \gcm_cmd_in.key1 [172]);
tran (gcm_cmd_in[270], \gcm_cmd_in.key1 [171]);
tran (gcm_cmd_in[269], \gcm_cmd_in.key1 [170]);
tran (gcm_cmd_in[268], \gcm_cmd_in.key1 [169]);
tran (gcm_cmd_in[267], \gcm_cmd_in.key1 [168]);
tran (gcm_cmd_in[266], \gcm_cmd_in.key1 [167]);
tran (gcm_cmd_in[265], \gcm_cmd_in.key1 [166]);
tran (gcm_cmd_in[264], \gcm_cmd_in.key1 [165]);
tran (gcm_cmd_in[263], \gcm_cmd_in.key1 [164]);
tran (gcm_cmd_in[262], \gcm_cmd_in.key1 [163]);
tran (gcm_cmd_in[261], \gcm_cmd_in.key1 [162]);
tran (gcm_cmd_in[260], \gcm_cmd_in.key1 [161]);
tran (gcm_cmd_in[259], \gcm_cmd_in.key1 [160]);
tran (gcm_cmd_in[258], \gcm_cmd_in.key1 [159]);
tran (gcm_cmd_in[257], \gcm_cmd_in.key1 [158]);
tran (gcm_cmd_in[256], \gcm_cmd_in.key1 [157]);
tran (gcm_cmd_in[255], \gcm_cmd_in.key1 [156]);
tran (gcm_cmd_in[254], \gcm_cmd_in.key1 [155]);
tran (gcm_cmd_in[253], \gcm_cmd_in.key1 [154]);
tran (gcm_cmd_in[252], \gcm_cmd_in.key1 [153]);
tran (gcm_cmd_in[251], \gcm_cmd_in.key1 [152]);
tran (gcm_cmd_in[250], \gcm_cmd_in.key1 [151]);
tran (gcm_cmd_in[249], \gcm_cmd_in.key1 [150]);
tran (gcm_cmd_in[248], \gcm_cmd_in.key1 [149]);
tran (gcm_cmd_in[247], \gcm_cmd_in.key1 [148]);
tran (gcm_cmd_in[246], \gcm_cmd_in.key1 [147]);
tran (gcm_cmd_in[245], \gcm_cmd_in.key1 [146]);
tran (gcm_cmd_in[244], \gcm_cmd_in.key1 [145]);
tran (gcm_cmd_in[243], \gcm_cmd_in.key1 [144]);
tran (gcm_cmd_in[242], \gcm_cmd_in.key1 [143]);
tran (gcm_cmd_in[241], \gcm_cmd_in.key1 [142]);
tran (gcm_cmd_in[240], \gcm_cmd_in.key1 [141]);
tran (gcm_cmd_in[239], \gcm_cmd_in.key1 [140]);
tran (gcm_cmd_in[238], \gcm_cmd_in.key1 [139]);
tran (gcm_cmd_in[237], \gcm_cmd_in.key1 [138]);
tran (gcm_cmd_in[236], \gcm_cmd_in.key1 [137]);
tran (gcm_cmd_in[235], \gcm_cmd_in.key1 [136]);
tran (gcm_cmd_in[234], \gcm_cmd_in.key1 [135]);
tran (gcm_cmd_in[233], \gcm_cmd_in.key1 [134]);
tran (gcm_cmd_in[232], \gcm_cmd_in.key1 [133]);
tran (gcm_cmd_in[231], \gcm_cmd_in.key1 [132]);
tran (gcm_cmd_in[230], \gcm_cmd_in.key1 [131]);
tran (gcm_cmd_in[229], \gcm_cmd_in.key1 [130]);
tran (gcm_cmd_in[228], \gcm_cmd_in.key1 [129]);
tran (gcm_cmd_in[227], \gcm_cmd_in.key1 [128]);
tran (gcm_cmd_in[226], \gcm_cmd_in.key1 [127]);
tran (gcm_cmd_in[225], \gcm_cmd_in.key1 [126]);
tran (gcm_cmd_in[224], \gcm_cmd_in.key1 [125]);
tran (gcm_cmd_in[223], \gcm_cmd_in.key1 [124]);
tran (gcm_cmd_in[222], \gcm_cmd_in.key1 [123]);
tran (gcm_cmd_in[221], \gcm_cmd_in.key1 [122]);
tran (gcm_cmd_in[220], \gcm_cmd_in.key1 [121]);
tran (gcm_cmd_in[219], \gcm_cmd_in.key1 [120]);
tran (gcm_cmd_in[218], \gcm_cmd_in.key1 [119]);
tran (gcm_cmd_in[217], \gcm_cmd_in.key1 [118]);
tran (gcm_cmd_in[216], \gcm_cmd_in.key1 [117]);
tran (gcm_cmd_in[215], \gcm_cmd_in.key1 [116]);
tran (gcm_cmd_in[214], \gcm_cmd_in.key1 [115]);
tran (gcm_cmd_in[213], \gcm_cmd_in.key1 [114]);
tran (gcm_cmd_in[212], \gcm_cmd_in.key1 [113]);
tran (gcm_cmd_in[211], \gcm_cmd_in.key1 [112]);
tran (gcm_cmd_in[210], \gcm_cmd_in.key1 [111]);
tran (gcm_cmd_in[209], \gcm_cmd_in.key1 [110]);
tran (gcm_cmd_in[208], \gcm_cmd_in.key1 [109]);
tran (gcm_cmd_in[207], \gcm_cmd_in.key1 [108]);
tran (gcm_cmd_in[206], \gcm_cmd_in.key1 [107]);
tran (gcm_cmd_in[205], \gcm_cmd_in.key1 [106]);
tran (gcm_cmd_in[204], \gcm_cmd_in.key1 [105]);
tran (gcm_cmd_in[203], \gcm_cmd_in.key1 [104]);
tran (gcm_cmd_in[202], \gcm_cmd_in.key1 [103]);
tran (gcm_cmd_in[201], \gcm_cmd_in.key1 [102]);
tran (gcm_cmd_in[200], \gcm_cmd_in.key1 [101]);
tran (gcm_cmd_in[199], \gcm_cmd_in.key1 [100]);
tran (gcm_cmd_in[198], \gcm_cmd_in.key1 [99]);
tran (gcm_cmd_in[197], \gcm_cmd_in.key1 [98]);
tran (gcm_cmd_in[196], \gcm_cmd_in.key1 [97]);
tran (gcm_cmd_in[195], \gcm_cmd_in.key1 [96]);
tran (gcm_cmd_in[194], \gcm_cmd_in.key1 [95]);
tran (gcm_cmd_in[193], \gcm_cmd_in.key1 [94]);
tran (gcm_cmd_in[192], \gcm_cmd_in.key1 [93]);
tran (gcm_cmd_in[191], \gcm_cmd_in.key1 [92]);
tran (gcm_cmd_in[190], \gcm_cmd_in.key1 [91]);
tran (gcm_cmd_in[189], \gcm_cmd_in.key1 [90]);
tran (gcm_cmd_in[188], \gcm_cmd_in.key1 [89]);
tran (gcm_cmd_in[187], \gcm_cmd_in.key1 [88]);
tran (gcm_cmd_in[186], \gcm_cmd_in.key1 [87]);
tran (gcm_cmd_in[185], \gcm_cmd_in.key1 [86]);
tran (gcm_cmd_in[184], \gcm_cmd_in.key1 [85]);
tran (gcm_cmd_in[183], \gcm_cmd_in.key1 [84]);
tran (gcm_cmd_in[182], \gcm_cmd_in.key1 [83]);
tran (gcm_cmd_in[181], \gcm_cmd_in.key1 [82]);
tran (gcm_cmd_in[180], \gcm_cmd_in.key1 [81]);
tran (gcm_cmd_in[179], \gcm_cmd_in.key1 [80]);
tran (gcm_cmd_in[178], \gcm_cmd_in.key1 [79]);
tran (gcm_cmd_in[177], \gcm_cmd_in.key1 [78]);
tran (gcm_cmd_in[176], \gcm_cmd_in.key1 [77]);
tran (gcm_cmd_in[175], \gcm_cmd_in.key1 [76]);
tran (gcm_cmd_in[174], \gcm_cmd_in.key1 [75]);
tran (gcm_cmd_in[173], \gcm_cmd_in.key1 [74]);
tran (gcm_cmd_in[172], \gcm_cmd_in.key1 [73]);
tran (gcm_cmd_in[171], \gcm_cmd_in.key1 [72]);
tran (gcm_cmd_in[170], \gcm_cmd_in.key1 [71]);
tran (gcm_cmd_in[169], \gcm_cmd_in.key1 [70]);
tran (gcm_cmd_in[168], \gcm_cmd_in.key1 [69]);
tran (gcm_cmd_in[167], \gcm_cmd_in.key1 [68]);
tran (gcm_cmd_in[166], \gcm_cmd_in.key1 [67]);
tran (gcm_cmd_in[165], \gcm_cmd_in.key1 [66]);
tran (gcm_cmd_in[164], \gcm_cmd_in.key1 [65]);
tran (gcm_cmd_in[163], \gcm_cmd_in.key1 [64]);
tran (gcm_cmd_in[162], \gcm_cmd_in.key1 [63]);
tran (gcm_cmd_in[161], \gcm_cmd_in.key1 [62]);
tran (gcm_cmd_in[160], \gcm_cmd_in.key1 [61]);
tran (gcm_cmd_in[159], \gcm_cmd_in.key1 [60]);
tran (gcm_cmd_in[158], \gcm_cmd_in.key1 [59]);
tran (gcm_cmd_in[157], \gcm_cmd_in.key1 [58]);
tran (gcm_cmd_in[156], \gcm_cmd_in.key1 [57]);
tran (gcm_cmd_in[155], \gcm_cmd_in.key1 [56]);
tran (gcm_cmd_in[154], \gcm_cmd_in.key1 [55]);
tran (gcm_cmd_in[153], \gcm_cmd_in.key1 [54]);
tran (gcm_cmd_in[152], \gcm_cmd_in.key1 [53]);
tran (gcm_cmd_in[151], \gcm_cmd_in.key1 [52]);
tran (gcm_cmd_in[150], \gcm_cmd_in.key1 [51]);
tran (gcm_cmd_in[149], \gcm_cmd_in.key1 [50]);
tran (gcm_cmd_in[148], \gcm_cmd_in.key1 [49]);
tran (gcm_cmd_in[147], \gcm_cmd_in.key1 [48]);
tran (gcm_cmd_in[146], \gcm_cmd_in.key1 [47]);
tran (gcm_cmd_in[145], \gcm_cmd_in.key1 [46]);
tran (gcm_cmd_in[144], \gcm_cmd_in.key1 [45]);
tran (gcm_cmd_in[143], \gcm_cmd_in.key1 [44]);
tran (gcm_cmd_in[142], \gcm_cmd_in.key1 [43]);
tran (gcm_cmd_in[141], \gcm_cmd_in.key1 [42]);
tran (gcm_cmd_in[140], \gcm_cmd_in.key1 [41]);
tran (gcm_cmd_in[139], \gcm_cmd_in.key1 [40]);
tran (gcm_cmd_in[138], \gcm_cmd_in.key1 [39]);
tran (gcm_cmd_in[137], \gcm_cmd_in.key1 [38]);
tran (gcm_cmd_in[136], \gcm_cmd_in.key1 [37]);
tran (gcm_cmd_in[135], \gcm_cmd_in.key1 [36]);
tran (gcm_cmd_in[134], \gcm_cmd_in.key1 [35]);
tran (gcm_cmd_in[133], \gcm_cmd_in.key1 [34]);
tran (gcm_cmd_in[132], \gcm_cmd_in.key1 [33]);
tran (gcm_cmd_in[131], \gcm_cmd_in.key1 [32]);
tran (gcm_cmd_in[130], \gcm_cmd_in.key1 [31]);
tran (gcm_cmd_in[129], \gcm_cmd_in.key1 [30]);
tran (gcm_cmd_in[128], \gcm_cmd_in.key1 [29]);
tran (gcm_cmd_in[127], \gcm_cmd_in.key1 [28]);
tran (gcm_cmd_in[126], \gcm_cmd_in.key1 [27]);
tran (gcm_cmd_in[125], \gcm_cmd_in.key1 [26]);
tran (gcm_cmd_in[124], \gcm_cmd_in.key1 [25]);
tran (gcm_cmd_in[123], \gcm_cmd_in.key1 [24]);
tran (gcm_cmd_in[122], \gcm_cmd_in.key1 [23]);
tran (gcm_cmd_in[121], \gcm_cmd_in.key1 [22]);
tran (gcm_cmd_in[120], \gcm_cmd_in.key1 [21]);
tran (gcm_cmd_in[119], \gcm_cmd_in.key1 [20]);
tran (gcm_cmd_in[118], \gcm_cmd_in.key1 [19]);
tran (gcm_cmd_in[117], \gcm_cmd_in.key1 [18]);
tran (gcm_cmd_in[116], \gcm_cmd_in.key1 [17]);
tran (gcm_cmd_in[115], \gcm_cmd_in.key1 [16]);
tran (gcm_cmd_in[114], \gcm_cmd_in.key1 [15]);
tran (gcm_cmd_in[113], \gcm_cmd_in.key1 [14]);
tran (gcm_cmd_in[112], \gcm_cmd_in.key1 [13]);
tran (gcm_cmd_in[111], \gcm_cmd_in.key1 [12]);
tran (gcm_cmd_in[110], \gcm_cmd_in.key1 [11]);
tran (gcm_cmd_in[109], \gcm_cmd_in.key1 [10]);
tran (gcm_cmd_in[108], \gcm_cmd_in.key1 [9]);
tran (gcm_cmd_in[107], \gcm_cmd_in.key1 [8]);
tran (gcm_cmd_in[106], \gcm_cmd_in.key1 [7]);
tran (gcm_cmd_in[105], \gcm_cmd_in.key1 [6]);
tran (gcm_cmd_in[104], \gcm_cmd_in.key1 [5]);
tran (gcm_cmd_in[103], \gcm_cmd_in.key1 [4]);
tran (gcm_cmd_in[102], \gcm_cmd_in.key1 [3]);
tran (gcm_cmd_in[101], \gcm_cmd_in.key1 [2]);
tran (gcm_cmd_in[100], \gcm_cmd_in.key1 [1]);
tran (gcm_cmd_in[99], \gcm_cmd_in.key1 [0]);
tran (gcm_cmd_in[98], \gcm_cmd_in.iv [95]);
tran (gcm_cmd_in[97], \gcm_cmd_in.iv [94]);
tran (gcm_cmd_in[96], \gcm_cmd_in.iv [93]);
tran (gcm_cmd_in[95], \gcm_cmd_in.iv [92]);
tran (gcm_cmd_in[94], \gcm_cmd_in.iv [91]);
tran (gcm_cmd_in[93], \gcm_cmd_in.iv [90]);
tran (gcm_cmd_in[92], \gcm_cmd_in.iv [89]);
tran (gcm_cmd_in[91], \gcm_cmd_in.iv [88]);
tran (gcm_cmd_in[90], \gcm_cmd_in.iv [87]);
tran (gcm_cmd_in[89], \gcm_cmd_in.iv [86]);
tran (gcm_cmd_in[88], \gcm_cmd_in.iv [85]);
tran (gcm_cmd_in[87], \gcm_cmd_in.iv [84]);
tran (gcm_cmd_in[86], \gcm_cmd_in.iv [83]);
tran (gcm_cmd_in[85], \gcm_cmd_in.iv [82]);
tran (gcm_cmd_in[84], \gcm_cmd_in.iv [81]);
tran (gcm_cmd_in[83], \gcm_cmd_in.iv [80]);
tran (gcm_cmd_in[82], \gcm_cmd_in.iv [79]);
tran (gcm_cmd_in[81], \gcm_cmd_in.iv [78]);
tran (gcm_cmd_in[80], \gcm_cmd_in.iv [77]);
tran (gcm_cmd_in[79], \gcm_cmd_in.iv [76]);
tran (gcm_cmd_in[78], \gcm_cmd_in.iv [75]);
tran (gcm_cmd_in[77], \gcm_cmd_in.iv [74]);
tran (gcm_cmd_in[76], \gcm_cmd_in.iv [73]);
tran (gcm_cmd_in[75], \gcm_cmd_in.iv [72]);
tran (gcm_cmd_in[74], \gcm_cmd_in.iv [71]);
tran (gcm_cmd_in[73], \gcm_cmd_in.iv [70]);
tran (gcm_cmd_in[72], \gcm_cmd_in.iv [69]);
tran (gcm_cmd_in[71], \gcm_cmd_in.iv [68]);
tran (gcm_cmd_in[70], \gcm_cmd_in.iv [67]);
tran (gcm_cmd_in[69], \gcm_cmd_in.iv [66]);
tran (gcm_cmd_in[68], \gcm_cmd_in.iv [65]);
tran (gcm_cmd_in[67], \gcm_cmd_in.iv [64]);
tran (gcm_cmd_in[66], \gcm_cmd_in.iv [63]);
tran (gcm_cmd_in[65], \gcm_cmd_in.iv [62]);
tran (gcm_cmd_in[64], \gcm_cmd_in.iv [61]);
tran (gcm_cmd_in[63], \gcm_cmd_in.iv [60]);
tran (gcm_cmd_in[62], \gcm_cmd_in.iv [59]);
tran (gcm_cmd_in[61], \gcm_cmd_in.iv [58]);
tran (gcm_cmd_in[60], \gcm_cmd_in.iv [57]);
tran (gcm_cmd_in[59], \gcm_cmd_in.iv [56]);
tran (gcm_cmd_in[58], \gcm_cmd_in.iv [55]);
tran (gcm_cmd_in[57], \gcm_cmd_in.iv [54]);
tran (gcm_cmd_in[56], \gcm_cmd_in.iv [53]);
tran (gcm_cmd_in[55], \gcm_cmd_in.iv [52]);
tran (gcm_cmd_in[54], \gcm_cmd_in.iv [51]);
tran (gcm_cmd_in[53], \gcm_cmd_in.iv [50]);
tran (gcm_cmd_in[52], \gcm_cmd_in.iv [49]);
tran (gcm_cmd_in[51], \gcm_cmd_in.iv [48]);
tran (gcm_cmd_in[50], \gcm_cmd_in.iv [47]);
tran (gcm_cmd_in[49], \gcm_cmd_in.iv [46]);
tran (gcm_cmd_in[48], \gcm_cmd_in.iv [45]);
tran (gcm_cmd_in[47], \gcm_cmd_in.iv [44]);
tran (gcm_cmd_in[46], \gcm_cmd_in.iv [43]);
tran (gcm_cmd_in[45], \gcm_cmd_in.iv [42]);
tran (gcm_cmd_in[44], \gcm_cmd_in.iv [41]);
tran (gcm_cmd_in[43], \gcm_cmd_in.iv [40]);
tran (gcm_cmd_in[42], \gcm_cmd_in.iv [39]);
tran (gcm_cmd_in[41], \gcm_cmd_in.iv [38]);
tran (gcm_cmd_in[40], \gcm_cmd_in.iv [37]);
tran (gcm_cmd_in[39], \gcm_cmd_in.iv [36]);
tran (gcm_cmd_in[38], \gcm_cmd_in.iv [35]);
tran (gcm_cmd_in[37], \gcm_cmd_in.iv [34]);
tran (gcm_cmd_in[36], \gcm_cmd_in.iv [33]);
tran (gcm_cmd_in[35], \gcm_cmd_in.iv [32]);
tran (gcm_cmd_in[34], \gcm_cmd_in.iv [31]);
tran (gcm_cmd_in[33], \gcm_cmd_in.iv [30]);
tran (gcm_cmd_in[32], \gcm_cmd_in.iv [29]);
tran (gcm_cmd_in[31], \gcm_cmd_in.iv [28]);
tran (gcm_cmd_in[30], \gcm_cmd_in.iv [27]);
tran (gcm_cmd_in[29], \gcm_cmd_in.iv [26]);
tran (gcm_cmd_in[28], \gcm_cmd_in.iv [25]);
tran (gcm_cmd_in[27], \gcm_cmd_in.iv [24]);
tran (gcm_cmd_in[26], \gcm_cmd_in.iv [23]);
tran (gcm_cmd_in[25], \gcm_cmd_in.iv [22]);
tran (gcm_cmd_in[24], \gcm_cmd_in.iv [21]);
tran (gcm_cmd_in[23], \gcm_cmd_in.iv [20]);
tran (gcm_cmd_in[22], \gcm_cmd_in.iv [19]);
tran (gcm_cmd_in[21], \gcm_cmd_in.iv [18]);
tran (gcm_cmd_in[20], \gcm_cmd_in.iv [17]);
tran (gcm_cmd_in[19], \gcm_cmd_in.iv [16]);
tran (gcm_cmd_in[18], \gcm_cmd_in.iv [15]);
tran (gcm_cmd_in[17], \gcm_cmd_in.iv [14]);
tran (gcm_cmd_in[16], \gcm_cmd_in.iv [13]);
tran (gcm_cmd_in[15], \gcm_cmd_in.iv [12]);
tran (gcm_cmd_in[14], \gcm_cmd_in.iv [11]);
tran (gcm_cmd_in[13], \gcm_cmd_in.iv [10]);
tran (gcm_cmd_in[12], \gcm_cmd_in.iv [9]);
tran (gcm_cmd_in[11], \gcm_cmd_in.iv [8]);
tran (gcm_cmd_in[10], \gcm_cmd_in.iv [7]);
tran (gcm_cmd_in[9], \gcm_cmd_in.iv [6]);
tran (gcm_cmd_in[8], \gcm_cmd_in.iv [5]);
tran (gcm_cmd_in[7], \gcm_cmd_in.iv [4]);
tran (gcm_cmd_in[6], \gcm_cmd_in.iv [3]);
tran (gcm_cmd_in[5], \gcm_cmd_in.iv [2]);
tran (gcm_cmd_in[4], \gcm_cmd_in.iv [1]);
tran (gcm_cmd_in[3], \gcm_cmd_in.iv [0]);
tran (gcm_cmd_in[2], \gcm_cmd_in.op [2]);
tran (gcm_cmd_in[1], \gcm_cmd_in.op [1]);
tran (gcm_cmd_in[0], \gcm_cmd_in.op [0]);
tran (keyfilter_cmd_in[0], \keyfilter_cmd_in.combo_mode [0]);
tran (kdfstream_cmd_in[262], \kdfstream_cmd_in.combo_mode [0]);
tran (kdfstream_cmd_in[261], \kdfstream_cmd_in.skip [0]);
tran (kdfstream_cmd_in[260], \kdfstream_cmd_in.guid [255]);
tran (kdfstream_cmd_in[259], \kdfstream_cmd_in.guid [254]);
tran (kdfstream_cmd_in[258], \kdfstream_cmd_in.guid [253]);
tran (kdfstream_cmd_in[257], \kdfstream_cmd_in.guid [252]);
tran (kdfstream_cmd_in[256], \kdfstream_cmd_in.guid [251]);
tran (kdfstream_cmd_in[255], \kdfstream_cmd_in.guid [250]);
tran (kdfstream_cmd_in[254], \kdfstream_cmd_in.guid [249]);
tran (kdfstream_cmd_in[253], \kdfstream_cmd_in.guid [248]);
tran (kdfstream_cmd_in[252], \kdfstream_cmd_in.guid [247]);
tran (kdfstream_cmd_in[251], \kdfstream_cmd_in.guid [246]);
tran (kdfstream_cmd_in[250], \kdfstream_cmd_in.guid [245]);
tran (kdfstream_cmd_in[249], \kdfstream_cmd_in.guid [244]);
tran (kdfstream_cmd_in[248], \kdfstream_cmd_in.guid [243]);
tran (kdfstream_cmd_in[247], \kdfstream_cmd_in.guid [242]);
tran (kdfstream_cmd_in[246], \kdfstream_cmd_in.guid [241]);
tran (kdfstream_cmd_in[245], \kdfstream_cmd_in.guid [240]);
tran (kdfstream_cmd_in[244], \kdfstream_cmd_in.guid [239]);
tran (kdfstream_cmd_in[243], \kdfstream_cmd_in.guid [238]);
tran (kdfstream_cmd_in[242], \kdfstream_cmd_in.guid [237]);
tran (kdfstream_cmd_in[241], \kdfstream_cmd_in.guid [236]);
tran (kdfstream_cmd_in[240], \kdfstream_cmd_in.guid [235]);
tran (kdfstream_cmd_in[239], \kdfstream_cmd_in.guid [234]);
tran (kdfstream_cmd_in[238], \kdfstream_cmd_in.guid [233]);
tran (kdfstream_cmd_in[237], \kdfstream_cmd_in.guid [232]);
tran (kdfstream_cmd_in[236], \kdfstream_cmd_in.guid [231]);
tran (kdfstream_cmd_in[235], \kdfstream_cmd_in.guid [230]);
tran (kdfstream_cmd_in[234], \kdfstream_cmd_in.guid [229]);
tran (kdfstream_cmd_in[233], \kdfstream_cmd_in.guid [228]);
tran (kdfstream_cmd_in[232], \kdfstream_cmd_in.guid [227]);
tran (kdfstream_cmd_in[231], \kdfstream_cmd_in.guid [226]);
tran (kdfstream_cmd_in[230], \kdfstream_cmd_in.guid [225]);
tran (kdfstream_cmd_in[229], \kdfstream_cmd_in.guid [224]);
tran (kdfstream_cmd_in[228], \kdfstream_cmd_in.guid [223]);
tran (kdfstream_cmd_in[227], \kdfstream_cmd_in.guid [222]);
tran (kdfstream_cmd_in[226], \kdfstream_cmd_in.guid [221]);
tran (kdfstream_cmd_in[225], \kdfstream_cmd_in.guid [220]);
tran (kdfstream_cmd_in[224], \kdfstream_cmd_in.guid [219]);
tran (kdfstream_cmd_in[223], \kdfstream_cmd_in.guid [218]);
tran (kdfstream_cmd_in[222], \kdfstream_cmd_in.guid [217]);
tran (kdfstream_cmd_in[221], \kdfstream_cmd_in.guid [216]);
tran (kdfstream_cmd_in[220], \kdfstream_cmd_in.guid [215]);
tran (kdfstream_cmd_in[219], \kdfstream_cmd_in.guid [214]);
tran (kdfstream_cmd_in[218], \kdfstream_cmd_in.guid [213]);
tran (kdfstream_cmd_in[217], \kdfstream_cmd_in.guid [212]);
tran (kdfstream_cmd_in[216], \kdfstream_cmd_in.guid [211]);
tran (kdfstream_cmd_in[215], \kdfstream_cmd_in.guid [210]);
tran (kdfstream_cmd_in[214], \kdfstream_cmd_in.guid [209]);
tran (kdfstream_cmd_in[213], \kdfstream_cmd_in.guid [208]);
tran (kdfstream_cmd_in[212], \kdfstream_cmd_in.guid [207]);
tran (kdfstream_cmd_in[211], \kdfstream_cmd_in.guid [206]);
tran (kdfstream_cmd_in[210], \kdfstream_cmd_in.guid [205]);
tran (kdfstream_cmd_in[209], \kdfstream_cmd_in.guid [204]);
tran (kdfstream_cmd_in[208], \kdfstream_cmd_in.guid [203]);
tran (kdfstream_cmd_in[207], \kdfstream_cmd_in.guid [202]);
tran (kdfstream_cmd_in[206], \kdfstream_cmd_in.guid [201]);
tran (kdfstream_cmd_in[205], \kdfstream_cmd_in.guid [200]);
tran (kdfstream_cmd_in[204], \kdfstream_cmd_in.guid [199]);
tran (kdfstream_cmd_in[203], \kdfstream_cmd_in.guid [198]);
tran (kdfstream_cmd_in[202], \kdfstream_cmd_in.guid [197]);
tran (kdfstream_cmd_in[201], \kdfstream_cmd_in.guid [196]);
tran (kdfstream_cmd_in[200], \kdfstream_cmd_in.guid [195]);
tran (kdfstream_cmd_in[199], \kdfstream_cmd_in.guid [194]);
tran (kdfstream_cmd_in[198], \kdfstream_cmd_in.guid [193]);
tran (kdfstream_cmd_in[197], \kdfstream_cmd_in.guid [192]);
tran (kdfstream_cmd_in[196], \kdfstream_cmd_in.guid [191]);
tran (kdfstream_cmd_in[195], \kdfstream_cmd_in.guid [190]);
tran (kdfstream_cmd_in[194], \kdfstream_cmd_in.guid [189]);
tran (kdfstream_cmd_in[193], \kdfstream_cmd_in.guid [188]);
tran (kdfstream_cmd_in[192], \kdfstream_cmd_in.guid [187]);
tran (kdfstream_cmd_in[191], \kdfstream_cmd_in.guid [186]);
tran (kdfstream_cmd_in[190], \kdfstream_cmd_in.guid [185]);
tran (kdfstream_cmd_in[189], \kdfstream_cmd_in.guid [184]);
tran (kdfstream_cmd_in[188], \kdfstream_cmd_in.guid [183]);
tran (kdfstream_cmd_in[187], \kdfstream_cmd_in.guid [182]);
tran (kdfstream_cmd_in[186], \kdfstream_cmd_in.guid [181]);
tran (kdfstream_cmd_in[185], \kdfstream_cmd_in.guid [180]);
tran (kdfstream_cmd_in[184], \kdfstream_cmd_in.guid [179]);
tran (kdfstream_cmd_in[183], \kdfstream_cmd_in.guid [178]);
tran (kdfstream_cmd_in[182], \kdfstream_cmd_in.guid [177]);
tran (kdfstream_cmd_in[181], \kdfstream_cmd_in.guid [176]);
tran (kdfstream_cmd_in[180], \kdfstream_cmd_in.guid [175]);
tran (kdfstream_cmd_in[179], \kdfstream_cmd_in.guid [174]);
tran (kdfstream_cmd_in[178], \kdfstream_cmd_in.guid [173]);
tran (kdfstream_cmd_in[177], \kdfstream_cmd_in.guid [172]);
tran (kdfstream_cmd_in[176], \kdfstream_cmd_in.guid [171]);
tran (kdfstream_cmd_in[175], \kdfstream_cmd_in.guid [170]);
tran (kdfstream_cmd_in[174], \kdfstream_cmd_in.guid [169]);
tran (kdfstream_cmd_in[173], \kdfstream_cmd_in.guid [168]);
tran (kdfstream_cmd_in[172], \kdfstream_cmd_in.guid [167]);
tran (kdfstream_cmd_in[171], \kdfstream_cmd_in.guid [166]);
tran (kdfstream_cmd_in[170], \kdfstream_cmd_in.guid [165]);
tran (kdfstream_cmd_in[169], \kdfstream_cmd_in.guid [164]);
tran (kdfstream_cmd_in[168], \kdfstream_cmd_in.guid [163]);
tran (kdfstream_cmd_in[167], \kdfstream_cmd_in.guid [162]);
tran (kdfstream_cmd_in[166], \kdfstream_cmd_in.guid [161]);
tran (kdfstream_cmd_in[165], \kdfstream_cmd_in.guid [160]);
tran (kdfstream_cmd_in[164], \kdfstream_cmd_in.guid [159]);
tran (kdfstream_cmd_in[163], \kdfstream_cmd_in.guid [158]);
tran (kdfstream_cmd_in[162], \kdfstream_cmd_in.guid [157]);
tran (kdfstream_cmd_in[161], \kdfstream_cmd_in.guid [156]);
tran (kdfstream_cmd_in[160], \kdfstream_cmd_in.guid [155]);
tran (kdfstream_cmd_in[159], \kdfstream_cmd_in.guid [154]);
tran (kdfstream_cmd_in[158], \kdfstream_cmd_in.guid [153]);
tran (kdfstream_cmd_in[157], \kdfstream_cmd_in.guid [152]);
tran (kdfstream_cmd_in[156], \kdfstream_cmd_in.guid [151]);
tran (kdfstream_cmd_in[155], \kdfstream_cmd_in.guid [150]);
tran (kdfstream_cmd_in[154], \kdfstream_cmd_in.guid [149]);
tran (kdfstream_cmd_in[153], \kdfstream_cmd_in.guid [148]);
tran (kdfstream_cmd_in[152], \kdfstream_cmd_in.guid [147]);
tran (kdfstream_cmd_in[151], \kdfstream_cmd_in.guid [146]);
tran (kdfstream_cmd_in[150], \kdfstream_cmd_in.guid [145]);
tran (kdfstream_cmd_in[149], \kdfstream_cmd_in.guid [144]);
tran (kdfstream_cmd_in[148], \kdfstream_cmd_in.guid [143]);
tran (kdfstream_cmd_in[147], \kdfstream_cmd_in.guid [142]);
tran (kdfstream_cmd_in[146], \kdfstream_cmd_in.guid [141]);
tran (kdfstream_cmd_in[145], \kdfstream_cmd_in.guid [140]);
tran (kdfstream_cmd_in[144], \kdfstream_cmd_in.guid [139]);
tran (kdfstream_cmd_in[143], \kdfstream_cmd_in.guid [138]);
tran (kdfstream_cmd_in[142], \kdfstream_cmd_in.guid [137]);
tran (kdfstream_cmd_in[141], \kdfstream_cmd_in.guid [136]);
tran (kdfstream_cmd_in[140], \kdfstream_cmd_in.guid [135]);
tran (kdfstream_cmd_in[139], \kdfstream_cmd_in.guid [134]);
tran (kdfstream_cmd_in[138], \kdfstream_cmd_in.guid [133]);
tran (kdfstream_cmd_in[137], \kdfstream_cmd_in.guid [132]);
tran (kdfstream_cmd_in[136], \kdfstream_cmd_in.guid [131]);
tran (kdfstream_cmd_in[135], \kdfstream_cmd_in.guid [130]);
tran (kdfstream_cmd_in[134], \kdfstream_cmd_in.guid [129]);
tran (kdfstream_cmd_in[133], \kdfstream_cmd_in.guid [128]);
tran (kdfstream_cmd_in[132], \kdfstream_cmd_in.guid [127]);
tran (kdfstream_cmd_in[131], \kdfstream_cmd_in.guid [126]);
tran (kdfstream_cmd_in[130], \kdfstream_cmd_in.guid [125]);
tran (kdfstream_cmd_in[129], \kdfstream_cmd_in.guid [124]);
tran (kdfstream_cmd_in[128], \kdfstream_cmd_in.guid [123]);
tran (kdfstream_cmd_in[127], \kdfstream_cmd_in.guid [122]);
tran (kdfstream_cmd_in[126], \kdfstream_cmd_in.guid [121]);
tran (kdfstream_cmd_in[125], \kdfstream_cmd_in.guid [120]);
tran (kdfstream_cmd_in[124], \kdfstream_cmd_in.guid [119]);
tran (kdfstream_cmd_in[123], \kdfstream_cmd_in.guid [118]);
tran (kdfstream_cmd_in[122], \kdfstream_cmd_in.guid [117]);
tran (kdfstream_cmd_in[121], \kdfstream_cmd_in.guid [116]);
tran (kdfstream_cmd_in[120], \kdfstream_cmd_in.guid [115]);
tran (kdfstream_cmd_in[119], \kdfstream_cmd_in.guid [114]);
tran (kdfstream_cmd_in[118], \kdfstream_cmd_in.guid [113]);
tran (kdfstream_cmd_in[117], \kdfstream_cmd_in.guid [112]);
tran (kdfstream_cmd_in[116], \kdfstream_cmd_in.guid [111]);
tran (kdfstream_cmd_in[115], \kdfstream_cmd_in.guid [110]);
tran (kdfstream_cmd_in[114], \kdfstream_cmd_in.guid [109]);
tran (kdfstream_cmd_in[113], \kdfstream_cmd_in.guid [108]);
tran (kdfstream_cmd_in[112], \kdfstream_cmd_in.guid [107]);
tran (kdfstream_cmd_in[111], \kdfstream_cmd_in.guid [106]);
tran (kdfstream_cmd_in[110], \kdfstream_cmd_in.guid [105]);
tran (kdfstream_cmd_in[109], \kdfstream_cmd_in.guid [104]);
tran (kdfstream_cmd_in[108], \kdfstream_cmd_in.guid [103]);
tran (kdfstream_cmd_in[107], \kdfstream_cmd_in.guid [102]);
tran (kdfstream_cmd_in[106], \kdfstream_cmd_in.guid [101]);
tran (kdfstream_cmd_in[105], \kdfstream_cmd_in.guid [100]);
tran (kdfstream_cmd_in[104], \kdfstream_cmd_in.guid [99]);
tran (kdfstream_cmd_in[103], \kdfstream_cmd_in.guid [98]);
tran (kdfstream_cmd_in[102], \kdfstream_cmd_in.guid [97]);
tran (kdfstream_cmd_in[101], \kdfstream_cmd_in.guid [96]);
tran (kdfstream_cmd_in[100], \kdfstream_cmd_in.guid [95]);
tran (kdfstream_cmd_in[99], \kdfstream_cmd_in.guid [94]);
tran (kdfstream_cmd_in[98], \kdfstream_cmd_in.guid [93]);
tran (kdfstream_cmd_in[97], \kdfstream_cmd_in.guid [92]);
tran (kdfstream_cmd_in[96], \kdfstream_cmd_in.guid [91]);
tran (kdfstream_cmd_in[95], \kdfstream_cmd_in.guid [90]);
tran (kdfstream_cmd_in[94], \kdfstream_cmd_in.guid [89]);
tran (kdfstream_cmd_in[93], \kdfstream_cmd_in.guid [88]);
tran (kdfstream_cmd_in[92], \kdfstream_cmd_in.guid [87]);
tran (kdfstream_cmd_in[91], \kdfstream_cmd_in.guid [86]);
tran (kdfstream_cmd_in[90], \kdfstream_cmd_in.guid [85]);
tran (kdfstream_cmd_in[89], \kdfstream_cmd_in.guid [84]);
tran (kdfstream_cmd_in[88], \kdfstream_cmd_in.guid [83]);
tran (kdfstream_cmd_in[87], \kdfstream_cmd_in.guid [82]);
tran (kdfstream_cmd_in[86], \kdfstream_cmd_in.guid [81]);
tran (kdfstream_cmd_in[85], \kdfstream_cmd_in.guid [80]);
tran (kdfstream_cmd_in[84], \kdfstream_cmd_in.guid [79]);
tran (kdfstream_cmd_in[83], \kdfstream_cmd_in.guid [78]);
tran (kdfstream_cmd_in[82], \kdfstream_cmd_in.guid [77]);
tran (kdfstream_cmd_in[81], \kdfstream_cmd_in.guid [76]);
tran (kdfstream_cmd_in[80], \kdfstream_cmd_in.guid [75]);
tran (kdfstream_cmd_in[79], \kdfstream_cmd_in.guid [74]);
tran (kdfstream_cmd_in[78], \kdfstream_cmd_in.guid [73]);
tran (kdfstream_cmd_in[77], \kdfstream_cmd_in.guid [72]);
tran (kdfstream_cmd_in[76], \kdfstream_cmd_in.guid [71]);
tran (kdfstream_cmd_in[75], \kdfstream_cmd_in.guid [70]);
tran (kdfstream_cmd_in[74], \kdfstream_cmd_in.guid [69]);
tran (kdfstream_cmd_in[73], \kdfstream_cmd_in.guid [68]);
tran (kdfstream_cmd_in[72], \kdfstream_cmd_in.guid [67]);
tran (kdfstream_cmd_in[71], \kdfstream_cmd_in.guid [66]);
tran (kdfstream_cmd_in[70], \kdfstream_cmd_in.guid [65]);
tran (kdfstream_cmd_in[69], \kdfstream_cmd_in.guid [64]);
tran (kdfstream_cmd_in[68], \kdfstream_cmd_in.guid [63]);
tran (kdfstream_cmd_in[67], \kdfstream_cmd_in.guid [62]);
tran (kdfstream_cmd_in[66], \kdfstream_cmd_in.guid [61]);
tran (kdfstream_cmd_in[65], \kdfstream_cmd_in.guid [60]);
tran (kdfstream_cmd_in[64], \kdfstream_cmd_in.guid [59]);
tran (kdfstream_cmd_in[63], \kdfstream_cmd_in.guid [58]);
tran (kdfstream_cmd_in[62], \kdfstream_cmd_in.guid [57]);
tran (kdfstream_cmd_in[61], \kdfstream_cmd_in.guid [56]);
tran (kdfstream_cmd_in[60], \kdfstream_cmd_in.guid [55]);
tran (kdfstream_cmd_in[59], \kdfstream_cmd_in.guid [54]);
tran (kdfstream_cmd_in[58], \kdfstream_cmd_in.guid [53]);
tran (kdfstream_cmd_in[57], \kdfstream_cmd_in.guid [52]);
tran (kdfstream_cmd_in[56], \kdfstream_cmd_in.guid [51]);
tran (kdfstream_cmd_in[55], \kdfstream_cmd_in.guid [50]);
tran (kdfstream_cmd_in[54], \kdfstream_cmd_in.guid [49]);
tran (kdfstream_cmd_in[53], \kdfstream_cmd_in.guid [48]);
tran (kdfstream_cmd_in[52], \kdfstream_cmd_in.guid [47]);
tran (kdfstream_cmd_in[51], \kdfstream_cmd_in.guid [46]);
tran (kdfstream_cmd_in[50], \kdfstream_cmd_in.guid [45]);
tran (kdfstream_cmd_in[49], \kdfstream_cmd_in.guid [44]);
tran (kdfstream_cmd_in[48], \kdfstream_cmd_in.guid [43]);
tran (kdfstream_cmd_in[47], \kdfstream_cmd_in.guid [42]);
tran (kdfstream_cmd_in[46], \kdfstream_cmd_in.guid [41]);
tran (kdfstream_cmd_in[45], \kdfstream_cmd_in.guid [40]);
tran (kdfstream_cmd_in[44], \kdfstream_cmd_in.guid [39]);
tran (kdfstream_cmd_in[43], \kdfstream_cmd_in.guid [38]);
tran (kdfstream_cmd_in[42], \kdfstream_cmd_in.guid [37]);
tran (kdfstream_cmd_in[41], \kdfstream_cmd_in.guid [36]);
tran (kdfstream_cmd_in[40], \kdfstream_cmd_in.guid [35]);
tran (kdfstream_cmd_in[39], \kdfstream_cmd_in.guid [34]);
tran (kdfstream_cmd_in[38], \kdfstream_cmd_in.guid [33]);
tran (kdfstream_cmd_in[37], \kdfstream_cmd_in.guid [32]);
tran (kdfstream_cmd_in[36], \kdfstream_cmd_in.guid [31]);
tran (kdfstream_cmd_in[35], \kdfstream_cmd_in.guid [30]);
tran (kdfstream_cmd_in[34], \kdfstream_cmd_in.guid [29]);
tran (kdfstream_cmd_in[33], \kdfstream_cmd_in.guid [28]);
tran (kdfstream_cmd_in[32], \kdfstream_cmd_in.guid [27]);
tran (kdfstream_cmd_in[31], \kdfstream_cmd_in.guid [26]);
tran (kdfstream_cmd_in[30], \kdfstream_cmd_in.guid [25]);
tran (kdfstream_cmd_in[29], \kdfstream_cmd_in.guid [24]);
tran (kdfstream_cmd_in[28], \kdfstream_cmd_in.guid [23]);
tran (kdfstream_cmd_in[27], \kdfstream_cmd_in.guid [22]);
tran (kdfstream_cmd_in[26], \kdfstream_cmd_in.guid [21]);
tran (kdfstream_cmd_in[25], \kdfstream_cmd_in.guid [20]);
tran (kdfstream_cmd_in[24], \kdfstream_cmd_in.guid [19]);
tran (kdfstream_cmd_in[23], \kdfstream_cmd_in.guid [18]);
tran (kdfstream_cmd_in[22], \kdfstream_cmd_in.guid [17]);
tran (kdfstream_cmd_in[21], \kdfstream_cmd_in.guid [16]);
tran (kdfstream_cmd_in[20], \kdfstream_cmd_in.guid [15]);
tran (kdfstream_cmd_in[19], \kdfstream_cmd_in.guid [14]);
tran (kdfstream_cmd_in[18], \kdfstream_cmd_in.guid [13]);
tran (kdfstream_cmd_in[17], \kdfstream_cmd_in.guid [12]);
tran (kdfstream_cmd_in[16], \kdfstream_cmd_in.guid [11]);
tran (kdfstream_cmd_in[15], \kdfstream_cmd_in.guid [10]);
tran (kdfstream_cmd_in[14], \kdfstream_cmd_in.guid [9]);
tran (kdfstream_cmd_in[13], \kdfstream_cmd_in.guid [8]);
tran (kdfstream_cmd_in[12], \kdfstream_cmd_in.guid [7]);
tran (kdfstream_cmd_in[11], \kdfstream_cmd_in.guid [6]);
tran (kdfstream_cmd_in[10], \kdfstream_cmd_in.guid [5]);
tran (kdfstream_cmd_in[9], \kdfstream_cmd_in.guid [4]);
tran (kdfstream_cmd_in[8], \kdfstream_cmd_in.guid [3]);
tran (kdfstream_cmd_in[7], \kdfstream_cmd_in.guid [2]);
tran (kdfstream_cmd_in[6], \kdfstream_cmd_in.guid [1]);
tran (kdfstream_cmd_in[5], \kdfstream_cmd_in.guid [0]);
tran (kdfstream_cmd_in[4], \kdfstream_cmd_in.label_index [2]);
tran (kdfstream_cmd_in[3], \kdfstream_cmd_in.label_index [1]);
tran (kdfstream_cmd_in[2], \kdfstream_cmd_in.label_index [0]);
tran (kdfstream_cmd_in[1], \kdfstream_cmd_in.num_iter [1]);
tran (kdfstream_cmd_in[0], \kdfstream_cmd_in.num_iter [0]);
tran (kdf_cmd_in[3], \kdf_cmd_in.kdf_dek_iter [0]);
tran (kdf_cmd_in[2], \kdf_cmd_in.combo_mode [0]);
tran (kdf_cmd_in[1], \kdf_cmd_in.dek_key_op [0]);
tran (kdf_cmd_in[0], \kdf_cmd_in.dak_key_op [0]);
tran (\labels[0][0] , \labels[0].delimiter[0] );
tran (\labels[0][1] , \labels[0].delimiter[1] );
tran (\labels[0][2] , \labels[0].delimiter[2] );
tran (\labels[0][3] , \labels[0].delimiter[3] );
tran (\labels[0][4] , \labels[0].delimiter[4] );
tran (\labels[0][5] , \labels[0].delimiter[5] );
tran (\labels[0][6] , \labels[0].delimiter[6] );
tran (\labels[0][7] , \labels[0].delimiter[7] );
tran (\labels[0][8] , \labels[0].delimiter_valid[0] );
tran (\labels[0][9] , \labels[0].label[0] );
tran (\labels[0][10] , \labels[0].label[1] );
tran (\labels[0][11] , \labels[0].label[2] );
tran (\labels[0][12] , \labels[0].label[3] );
tran (\labels[0][13] , \labels[0].label[4] );
tran (\labels[0][14] , \labels[0].label[5] );
tran (\labels[0][15] , \labels[0].label[6] );
tran (\labels[0][16] , \labels[0].label[7] );
tran (\labels[0][17] , \labels[0].label[8] );
tran (\labels[0][18] , \labels[0].label[9] );
tran (\labels[0][19] , \labels[0].label[10] );
tran (\labels[0][20] , \labels[0].label[11] );
tran (\labels[0][21] , \labels[0].label[12] );
tran (\labels[0][22] , \labels[0].label[13] );
tran (\labels[0][23] , \labels[0].label[14] );
tran (\labels[0][24] , \labels[0].label[15] );
tran (\labels[0][25] , \labels[0].label[16] );
tran (\labels[0][26] , \labels[0].label[17] );
tran (\labels[0][27] , \labels[0].label[18] );
tran (\labels[0][28] , \labels[0].label[19] );
tran (\labels[0][29] , \labels[0].label[20] );
tran (\labels[0][30] , \labels[0].label[21] );
tran (\labels[0][31] , \labels[0].label[22] );
tran (\labels[0][32] , \labels[0].label[23] );
tran (\labels[0][33] , \labels[0].label[24] );
tran (\labels[0][34] , \labels[0].label[25] );
tran (\labels[0][35] , \labels[0].label[26] );
tran (\labels[0][36] , \labels[0].label[27] );
tran (\labels[0][37] , \labels[0].label[28] );
tran (\labels[0][38] , \labels[0].label[29] );
tran (\labels[0][39] , \labels[0].label[30] );
tran (\labels[0][40] , \labels[0].label[31] );
tran (\labels[0][41] , \labels[0].label[32] );
tran (\labels[0][42] , \labels[0].label[33] );
tran (\labels[0][43] , \labels[0].label[34] );
tran (\labels[0][44] , \labels[0].label[35] );
tran (\labels[0][45] , \labels[0].label[36] );
tran (\labels[0][46] , \labels[0].label[37] );
tran (\labels[0][47] , \labels[0].label[38] );
tran (\labels[0][48] , \labels[0].label[39] );
tran (\labels[0][49] , \labels[0].label[40] );
tran (\labels[0][50] , \labels[0].label[41] );
tran (\labels[0][51] , \labels[0].label[42] );
tran (\labels[0][52] , \labels[0].label[43] );
tran (\labels[0][53] , \labels[0].label[44] );
tran (\labels[0][54] , \labels[0].label[45] );
tran (\labels[0][55] , \labels[0].label[46] );
tran (\labels[0][56] , \labels[0].label[47] );
tran (\labels[0][57] , \labels[0].label[48] );
tran (\labels[0][58] , \labels[0].label[49] );
tran (\labels[0][59] , \labels[0].label[50] );
tran (\labels[0][60] , \labels[0].label[51] );
tran (\labels[0][61] , \labels[0].label[52] );
tran (\labels[0][62] , \labels[0].label[53] );
tran (\labels[0][63] , \labels[0].label[54] );
tran (\labels[0][64] , \labels[0].label[55] );
tran (\labels[0][65] , \labels[0].label[56] );
tran (\labels[0][66] , \labels[0].label[57] );
tran (\labels[0][67] , \labels[0].label[58] );
tran (\labels[0][68] , \labels[0].label[59] );
tran (\labels[0][69] , \labels[0].label[60] );
tran (\labels[0][70] , \labels[0].label[61] );
tran (\labels[0][71] , \labels[0].label[62] );
tran (\labels[0][72] , \labels[0].label[63] );
tran (\labels[0][73] , \labels[0].label[64] );
tran (\labels[0][74] , \labels[0].label[65] );
tran (\labels[0][75] , \labels[0].label[66] );
tran (\labels[0][76] , \labels[0].label[67] );
tran (\labels[0][77] , \labels[0].label[68] );
tran (\labels[0][78] , \labels[0].label[69] );
tran (\labels[0][79] , \labels[0].label[70] );
tran (\labels[0][80] , \labels[0].label[71] );
tran (\labels[0][81] , \labels[0].label[72] );
tran (\labels[0][82] , \labels[0].label[73] );
tran (\labels[0][83] , \labels[0].label[74] );
tran (\labels[0][84] , \labels[0].label[75] );
tran (\labels[0][85] , \labels[0].label[76] );
tran (\labels[0][86] , \labels[0].label[77] );
tran (\labels[0][87] , \labels[0].label[78] );
tran (\labels[0][88] , \labels[0].label[79] );
tran (\labels[0][89] , \labels[0].label[80] );
tran (\labels[0][90] , \labels[0].label[81] );
tran (\labels[0][91] , \labels[0].label[82] );
tran (\labels[0][92] , \labels[0].label[83] );
tran (\labels[0][93] , \labels[0].label[84] );
tran (\labels[0][94] , \labels[0].label[85] );
tran (\labels[0][95] , \labels[0].label[86] );
tran (\labels[0][96] , \labels[0].label[87] );
tran (\labels[0][97] , \labels[0].label[88] );
tran (\labels[0][98] , \labels[0].label[89] );
tran (\labels[0][99] , \labels[0].label[90] );
tran (\labels[0][100] , \labels[0].label[91] );
tran (\labels[0][101] , \labels[0].label[92] );
tran (\labels[0][102] , \labels[0].label[93] );
tran (\labels[0][103] , \labels[0].label[94] );
tran (\labels[0][104] , \labels[0].label[95] );
tran (\labels[0][105] , \labels[0].label[96] );
tran (\labels[0][106] , \labels[0].label[97] );
tran (\labels[0][107] , \labels[0].label[98] );
tran (\labels[0][108] , \labels[0].label[99] );
tran (\labels[0][109] , \labels[0].label[100] );
tran (\labels[0][110] , \labels[0].label[101] );
tran (\labels[0][111] , \labels[0].label[102] );
tran (\labels[0][112] , \labels[0].label[103] );
tran (\labels[0][113] , \labels[0].label[104] );
tran (\labels[0][114] , \labels[0].label[105] );
tran (\labels[0][115] , \labels[0].label[106] );
tran (\labels[0][116] , \labels[0].label[107] );
tran (\labels[0][117] , \labels[0].label[108] );
tran (\labels[0][118] , \labels[0].label[109] );
tran (\labels[0][119] , \labels[0].label[110] );
tran (\labels[0][120] , \labels[0].label[111] );
tran (\labels[0][121] , \labels[0].label[112] );
tran (\labels[0][122] , \labels[0].label[113] );
tran (\labels[0][123] , \labels[0].label[114] );
tran (\labels[0][124] , \labels[0].label[115] );
tran (\labels[0][125] , \labels[0].label[116] );
tran (\labels[0][126] , \labels[0].label[117] );
tran (\labels[0][127] , \labels[0].label[118] );
tran (\labels[0][128] , \labels[0].label[119] );
tran (\labels[0][129] , \labels[0].label[120] );
tran (\labels[0][130] , \labels[0].label[121] );
tran (\labels[0][131] , \labels[0].label[122] );
tran (\labels[0][132] , \labels[0].label[123] );
tran (\labels[0][133] , \labels[0].label[124] );
tran (\labels[0][134] , \labels[0].label[125] );
tran (\labels[0][135] , \labels[0].label[126] );
tran (\labels[0][136] , \labels[0].label[127] );
tran (\labels[0][137] , \labels[0].label[128] );
tran (\labels[0][138] , \labels[0].label[129] );
tran (\labels[0][139] , \labels[0].label[130] );
tran (\labels[0][140] , \labels[0].label[131] );
tran (\labels[0][141] , \labels[0].label[132] );
tran (\labels[0][142] , \labels[0].label[133] );
tran (\labels[0][143] , \labels[0].label[134] );
tran (\labels[0][144] , \labels[0].label[135] );
tran (\labels[0][145] , \labels[0].label[136] );
tran (\labels[0][146] , \labels[0].label[137] );
tran (\labels[0][147] , \labels[0].label[138] );
tran (\labels[0][148] , \labels[0].label[139] );
tran (\labels[0][149] , \labels[0].label[140] );
tran (\labels[0][150] , \labels[0].label[141] );
tran (\labels[0][151] , \labels[0].label[142] );
tran (\labels[0][152] , \labels[0].label[143] );
tran (\labels[0][153] , \labels[0].label[144] );
tran (\labels[0][154] , \labels[0].label[145] );
tran (\labels[0][155] , \labels[0].label[146] );
tran (\labels[0][156] , \labels[0].label[147] );
tran (\labels[0][157] , \labels[0].label[148] );
tran (\labels[0][158] , \labels[0].label[149] );
tran (\labels[0][159] , \labels[0].label[150] );
tran (\labels[0][160] , \labels[0].label[151] );
tran (\labels[0][161] , \labels[0].label[152] );
tran (\labels[0][162] , \labels[0].label[153] );
tran (\labels[0][163] , \labels[0].label[154] );
tran (\labels[0][164] , \labels[0].label[155] );
tran (\labels[0][165] , \labels[0].label[156] );
tran (\labels[0][166] , \labels[0].label[157] );
tran (\labels[0][167] , \labels[0].label[158] );
tran (\labels[0][168] , \labels[0].label[159] );
tran (\labels[0][169] , \labels[0].label[160] );
tran (\labels[0][170] , \labels[0].label[161] );
tran (\labels[0][171] , \labels[0].label[162] );
tran (\labels[0][172] , \labels[0].label[163] );
tran (\labels[0][173] , \labels[0].label[164] );
tran (\labels[0][174] , \labels[0].label[165] );
tran (\labels[0][175] , \labels[0].label[166] );
tran (\labels[0][176] , \labels[0].label[167] );
tran (\labels[0][177] , \labels[0].label[168] );
tran (\labels[0][178] , \labels[0].label[169] );
tran (\labels[0][179] , \labels[0].label[170] );
tran (\labels[0][180] , \labels[0].label[171] );
tran (\labels[0][181] , \labels[0].label[172] );
tran (\labels[0][182] , \labels[0].label[173] );
tran (\labels[0][183] , \labels[0].label[174] );
tran (\labels[0][184] , \labels[0].label[175] );
tran (\labels[0][185] , \labels[0].label[176] );
tran (\labels[0][186] , \labels[0].label[177] );
tran (\labels[0][187] , \labels[0].label[178] );
tran (\labels[0][188] , \labels[0].label[179] );
tran (\labels[0][189] , \labels[0].label[180] );
tran (\labels[0][190] , \labels[0].label[181] );
tran (\labels[0][191] , \labels[0].label[182] );
tran (\labels[0][192] , \labels[0].label[183] );
tran (\labels[0][193] , \labels[0].label[184] );
tran (\labels[0][194] , \labels[0].label[185] );
tran (\labels[0][195] , \labels[0].label[186] );
tran (\labels[0][196] , \labels[0].label[187] );
tran (\labels[0][197] , \labels[0].label[188] );
tran (\labels[0][198] , \labels[0].label[189] );
tran (\labels[0][199] , \labels[0].label[190] );
tran (\labels[0][200] , \labels[0].label[191] );
tran (\labels[0][201] , \labels[0].label[192] );
tran (\labels[0][202] , \labels[0].label[193] );
tran (\labels[0][203] , \labels[0].label[194] );
tran (\labels[0][204] , \labels[0].label[195] );
tran (\labels[0][205] , \labels[0].label[196] );
tran (\labels[0][206] , \labels[0].label[197] );
tran (\labels[0][207] , \labels[0].label[198] );
tran (\labels[0][208] , \labels[0].label[199] );
tran (\labels[0][209] , \labels[0].label[200] );
tran (\labels[0][210] , \labels[0].label[201] );
tran (\labels[0][211] , \labels[0].label[202] );
tran (\labels[0][212] , \labels[0].label[203] );
tran (\labels[0][213] , \labels[0].label[204] );
tran (\labels[0][214] , \labels[0].label[205] );
tran (\labels[0][215] , \labels[0].label[206] );
tran (\labels[0][216] , \labels[0].label[207] );
tran (\labels[0][217] , \labels[0].label[208] );
tran (\labels[0][218] , \labels[0].label[209] );
tran (\labels[0][219] , \labels[0].label[210] );
tran (\labels[0][220] , \labels[0].label[211] );
tran (\labels[0][221] , \labels[0].label[212] );
tran (\labels[0][222] , \labels[0].label[213] );
tran (\labels[0][223] , \labels[0].label[214] );
tran (\labels[0][224] , \labels[0].label[215] );
tran (\labels[0][225] , \labels[0].label[216] );
tran (\labels[0][226] , \labels[0].label[217] );
tran (\labels[0][227] , \labels[0].label[218] );
tran (\labels[0][228] , \labels[0].label[219] );
tran (\labels[0][229] , \labels[0].label[220] );
tran (\labels[0][230] , \labels[0].label[221] );
tran (\labels[0][231] , \labels[0].label[222] );
tran (\labels[0][232] , \labels[0].label[223] );
tran (\labels[0][233] , \labels[0].label[224] );
tran (\labels[0][234] , \labels[0].label[225] );
tran (\labels[0][235] , \labels[0].label[226] );
tran (\labels[0][236] , \labels[0].label[227] );
tran (\labels[0][237] , \labels[0].label[228] );
tran (\labels[0][238] , \labels[0].label[229] );
tran (\labels[0][239] , \labels[0].label[230] );
tran (\labels[0][240] , \labels[0].label[231] );
tran (\labels[0][241] , \labels[0].label[232] );
tran (\labels[0][242] , \labels[0].label[233] );
tran (\labels[0][243] , \labels[0].label[234] );
tran (\labels[0][244] , \labels[0].label[235] );
tran (\labels[0][245] , \labels[0].label[236] );
tran (\labels[0][246] , \labels[0].label[237] );
tran (\labels[0][247] , \labels[0].label[238] );
tran (\labels[0][248] , \labels[0].label[239] );
tran (\labels[0][249] , \labels[0].label[240] );
tran (\labels[0][250] , \labels[0].label[241] );
tran (\labels[0][251] , \labels[0].label[242] );
tran (\labels[0][252] , \labels[0].label[243] );
tran (\labels[0][253] , \labels[0].label[244] );
tran (\labels[0][254] , \labels[0].label[245] );
tran (\labels[0][255] , \labels[0].label[246] );
tran (\labels[0][256] , \labels[0].label[247] );
tran (\labels[0][257] , \labels[0].label[248] );
tran (\labels[0][258] , \labels[0].label[249] );
tran (\labels[0][259] , \labels[0].label[250] );
tran (\labels[0][260] , \labels[0].label[251] );
tran (\labels[0][261] , \labels[0].label[252] );
tran (\labels[0][262] , \labels[0].label[253] );
tran (\labels[0][263] , \labels[0].label[254] );
tran (\labels[0][264] , \labels[0].label[255] );
tran (\labels[0][265] , \labels[0].label_size[0] );
tran (\labels[0][266] , \labels[0].label_size[1] );
tran (\labels[0][267] , \labels[0].label_size[2] );
tran (\labels[0][268] , \labels[0].label_size[3] );
tran (\labels[0][269] , \labels[0].label_size[4] );
tran (\labels[0][270] , \labels[0].label_size[5] );
tran (\labels[0][271] , \labels[0].guid_size[0] );
tran (\labels[1][0] , \labels[1].delimiter[0] );
tran (\labels[1][1] , \labels[1].delimiter[1] );
tran (\labels[1][2] , \labels[1].delimiter[2] );
tran (\labels[1][3] , \labels[1].delimiter[3] );
tran (\labels[1][4] , \labels[1].delimiter[4] );
tran (\labels[1][5] , \labels[1].delimiter[5] );
tran (\labels[1][6] , \labels[1].delimiter[6] );
tran (\labels[1][7] , \labels[1].delimiter[7] );
tran (\labels[1][8] , \labels[1].delimiter_valid[0] );
tran (\labels[1][9] , \labels[1].label[0] );
tran (\labels[1][10] , \labels[1].label[1] );
tran (\labels[1][11] , \labels[1].label[2] );
tran (\labels[1][12] , \labels[1].label[3] );
tran (\labels[1][13] , \labels[1].label[4] );
tran (\labels[1][14] , \labels[1].label[5] );
tran (\labels[1][15] , \labels[1].label[6] );
tran (\labels[1][16] , \labels[1].label[7] );
tran (\labels[1][17] , \labels[1].label[8] );
tran (\labels[1][18] , \labels[1].label[9] );
tran (\labels[1][19] , \labels[1].label[10] );
tran (\labels[1][20] , \labels[1].label[11] );
tran (\labels[1][21] , \labels[1].label[12] );
tran (\labels[1][22] , \labels[1].label[13] );
tran (\labels[1][23] , \labels[1].label[14] );
tran (\labels[1][24] , \labels[1].label[15] );
tran (\labels[1][25] , \labels[1].label[16] );
tran (\labels[1][26] , \labels[1].label[17] );
tran (\labels[1][27] , \labels[1].label[18] );
tran (\labels[1][28] , \labels[1].label[19] );
tran (\labels[1][29] , \labels[1].label[20] );
tran (\labels[1][30] , \labels[1].label[21] );
tran (\labels[1][31] , \labels[1].label[22] );
tran (\labels[1][32] , \labels[1].label[23] );
tran (\labels[1][33] , \labels[1].label[24] );
tran (\labels[1][34] , \labels[1].label[25] );
tran (\labels[1][35] , \labels[1].label[26] );
tran (\labels[1][36] , \labels[1].label[27] );
tran (\labels[1][37] , \labels[1].label[28] );
tran (\labels[1][38] , \labels[1].label[29] );
tran (\labels[1][39] , \labels[1].label[30] );
tran (\labels[1][40] , \labels[1].label[31] );
tran (\labels[1][41] , \labels[1].label[32] );
tran (\labels[1][42] , \labels[1].label[33] );
tran (\labels[1][43] , \labels[1].label[34] );
tran (\labels[1][44] , \labels[1].label[35] );
tran (\labels[1][45] , \labels[1].label[36] );
tran (\labels[1][46] , \labels[1].label[37] );
tran (\labels[1][47] , \labels[1].label[38] );
tran (\labels[1][48] , \labels[1].label[39] );
tran (\labels[1][49] , \labels[1].label[40] );
tran (\labels[1][50] , \labels[1].label[41] );
tran (\labels[1][51] , \labels[1].label[42] );
tran (\labels[1][52] , \labels[1].label[43] );
tran (\labels[1][53] , \labels[1].label[44] );
tran (\labels[1][54] , \labels[1].label[45] );
tran (\labels[1][55] , \labels[1].label[46] );
tran (\labels[1][56] , \labels[1].label[47] );
tran (\labels[1][57] , \labels[1].label[48] );
tran (\labels[1][58] , \labels[1].label[49] );
tran (\labels[1][59] , \labels[1].label[50] );
tran (\labels[1][60] , \labels[1].label[51] );
tran (\labels[1][61] , \labels[1].label[52] );
tran (\labels[1][62] , \labels[1].label[53] );
tran (\labels[1][63] , \labels[1].label[54] );
tran (\labels[1][64] , \labels[1].label[55] );
tran (\labels[1][65] , \labels[1].label[56] );
tran (\labels[1][66] , \labels[1].label[57] );
tran (\labels[1][67] , \labels[1].label[58] );
tran (\labels[1][68] , \labels[1].label[59] );
tran (\labels[1][69] , \labels[1].label[60] );
tran (\labels[1][70] , \labels[1].label[61] );
tran (\labels[1][71] , \labels[1].label[62] );
tran (\labels[1][72] , \labels[1].label[63] );
tran (\labels[1][73] , \labels[1].label[64] );
tran (\labels[1][74] , \labels[1].label[65] );
tran (\labels[1][75] , \labels[1].label[66] );
tran (\labels[1][76] , \labels[1].label[67] );
tran (\labels[1][77] , \labels[1].label[68] );
tran (\labels[1][78] , \labels[1].label[69] );
tran (\labels[1][79] , \labels[1].label[70] );
tran (\labels[1][80] , \labels[1].label[71] );
tran (\labels[1][81] , \labels[1].label[72] );
tran (\labels[1][82] , \labels[1].label[73] );
tran (\labels[1][83] , \labels[1].label[74] );
tran (\labels[1][84] , \labels[1].label[75] );
tran (\labels[1][85] , \labels[1].label[76] );
tran (\labels[1][86] , \labels[1].label[77] );
tran (\labels[1][87] , \labels[1].label[78] );
tran (\labels[1][88] , \labels[1].label[79] );
tran (\labels[1][89] , \labels[1].label[80] );
tran (\labels[1][90] , \labels[1].label[81] );
tran (\labels[1][91] , \labels[1].label[82] );
tran (\labels[1][92] , \labels[1].label[83] );
tran (\labels[1][93] , \labels[1].label[84] );
tran (\labels[1][94] , \labels[1].label[85] );
tran (\labels[1][95] , \labels[1].label[86] );
tran (\labels[1][96] , \labels[1].label[87] );
tran (\labels[1][97] , \labels[1].label[88] );
tran (\labels[1][98] , \labels[1].label[89] );
tran (\labels[1][99] , \labels[1].label[90] );
tran (\labels[1][100] , \labels[1].label[91] );
tran (\labels[1][101] , \labels[1].label[92] );
tran (\labels[1][102] , \labels[1].label[93] );
tran (\labels[1][103] , \labels[1].label[94] );
tran (\labels[1][104] , \labels[1].label[95] );
tran (\labels[1][105] , \labels[1].label[96] );
tran (\labels[1][106] , \labels[1].label[97] );
tran (\labels[1][107] , \labels[1].label[98] );
tran (\labels[1][108] , \labels[1].label[99] );
tran (\labels[1][109] , \labels[1].label[100] );
tran (\labels[1][110] , \labels[1].label[101] );
tran (\labels[1][111] , \labels[1].label[102] );
tran (\labels[1][112] , \labels[1].label[103] );
tran (\labels[1][113] , \labels[1].label[104] );
tran (\labels[1][114] , \labels[1].label[105] );
tran (\labels[1][115] , \labels[1].label[106] );
tran (\labels[1][116] , \labels[1].label[107] );
tran (\labels[1][117] , \labels[1].label[108] );
tran (\labels[1][118] , \labels[1].label[109] );
tran (\labels[1][119] , \labels[1].label[110] );
tran (\labels[1][120] , \labels[1].label[111] );
tran (\labels[1][121] , \labels[1].label[112] );
tran (\labels[1][122] , \labels[1].label[113] );
tran (\labels[1][123] , \labels[1].label[114] );
tran (\labels[1][124] , \labels[1].label[115] );
tran (\labels[1][125] , \labels[1].label[116] );
tran (\labels[1][126] , \labels[1].label[117] );
tran (\labels[1][127] , \labels[1].label[118] );
tran (\labels[1][128] , \labels[1].label[119] );
tran (\labels[1][129] , \labels[1].label[120] );
tran (\labels[1][130] , \labels[1].label[121] );
tran (\labels[1][131] , \labels[1].label[122] );
tran (\labels[1][132] , \labels[1].label[123] );
tran (\labels[1][133] , \labels[1].label[124] );
tran (\labels[1][134] , \labels[1].label[125] );
tran (\labels[1][135] , \labels[1].label[126] );
tran (\labels[1][136] , \labels[1].label[127] );
tran (\labels[1][137] , \labels[1].label[128] );
tran (\labels[1][138] , \labels[1].label[129] );
tran (\labels[1][139] , \labels[1].label[130] );
tran (\labels[1][140] , \labels[1].label[131] );
tran (\labels[1][141] , \labels[1].label[132] );
tran (\labels[1][142] , \labels[1].label[133] );
tran (\labels[1][143] , \labels[1].label[134] );
tran (\labels[1][144] , \labels[1].label[135] );
tran (\labels[1][145] , \labels[1].label[136] );
tran (\labels[1][146] , \labels[1].label[137] );
tran (\labels[1][147] , \labels[1].label[138] );
tran (\labels[1][148] , \labels[1].label[139] );
tran (\labels[1][149] , \labels[1].label[140] );
tran (\labels[1][150] , \labels[1].label[141] );
tran (\labels[1][151] , \labels[1].label[142] );
tran (\labels[1][152] , \labels[1].label[143] );
tran (\labels[1][153] , \labels[1].label[144] );
tran (\labels[1][154] , \labels[1].label[145] );
tran (\labels[1][155] , \labels[1].label[146] );
tran (\labels[1][156] , \labels[1].label[147] );
tran (\labels[1][157] , \labels[1].label[148] );
tran (\labels[1][158] , \labels[1].label[149] );
tran (\labels[1][159] , \labels[1].label[150] );
tran (\labels[1][160] , \labels[1].label[151] );
tran (\labels[1][161] , \labels[1].label[152] );
tran (\labels[1][162] , \labels[1].label[153] );
tran (\labels[1][163] , \labels[1].label[154] );
tran (\labels[1][164] , \labels[1].label[155] );
tran (\labels[1][165] , \labels[1].label[156] );
tran (\labels[1][166] , \labels[1].label[157] );
tran (\labels[1][167] , \labels[1].label[158] );
tran (\labels[1][168] , \labels[1].label[159] );
tran (\labels[1][169] , \labels[1].label[160] );
tran (\labels[1][170] , \labels[1].label[161] );
tran (\labels[1][171] , \labels[1].label[162] );
tran (\labels[1][172] , \labels[1].label[163] );
tran (\labels[1][173] , \labels[1].label[164] );
tran (\labels[1][174] , \labels[1].label[165] );
tran (\labels[1][175] , \labels[1].label[166] );
tran (\labels[1][176] , \labels[1].label[167] );
tran (\labels[1][177] , \labels[1].label[168] );
tran (\labels[1][178] , \labels[1].label[169] );
tran (\labels[1][179] , \labels[1].label[170] );
tran (\labels[1][180] , \labels[1].label[171] );
tran (\labels[1][181] , \labels[1].label[172] );
tran (\labels[1][182] , \labels[1].label[173] );
tran (\labels[1][183] , \labels[1].label[174] );
tran (\labels[1][184] , \labels[1].label[175] );
tran (\labels[1][185] , \labels[1].label[176] );
tran (\labels[1][186] , \labels[1].label[177] );
tran (\labels[1][187] , \labels[1].label[178] );
tran (\labels[1][188] , \labels[1].label[179] );
tran (\labels[1][189] , \labels[1].label[180] );
tran (\labels[1][190] , \labels[1].label[181] );
tran (\labels[1][191] , \labels[1].label[182] );
tran (\labels[1][192] , \labels[1].label[183] );
tran (\labels[1][193] , \labels[1].label[184] );
tran (\labels[1][194] , \labels[1].label[185] );
tran (\labels[1][195] , \labels[1].label[186] );
tran (\labels[1][196] , \labels[1].label[187] );
tran (\labels[1][197] , \labels[1].label[188] );
tran (\labels[1][198] , \labels[1].label[189] );
tran (\labels[1][199] , \labels[1].label[190] );
tran (\labels[1][200] , \labels[1].label[191] );
tran (\labels[1][201] , \labels[1].label[192] );
tran (\labels[1][202] , \labels[1].label[193] );
tran (\labels[1][203] , \labels[1].label[194] );
tran (\labels[1][204] , \labels[1].label[195] );
tran (\labels[1][205] , \labels[1].label[196] );
tran (\labels[1][206] , \labels[1].label[197] );
tran (\labels[1][207] , \labels[1].label[198] );
tran (\labels[1][208] , \labels[1].label[199] );
tran (\labels[1][209] , \labels[1].label[200] );
tran (\labels[1][210] , \labels[1].label[201] );
tran (\labels[1][211] , \labels[1].label[202] );
tran (\labels[1][212] , \labels[1].label[203] );
tran (\labels[1][213] , \labels[1].label[204] );
tran (\labels[1][214] , \labels[1].label[205] );
tran (\labels[1][215] , \labels[1].label[206] );
tran (\labels[1][216] , \labels[1].label[207] );
tran (\labels[1][217] , \labels[1].label[208] );
tran (\labels[1][218] , \labels[1].label[209] );
tran (\labels[1][219] , \labels[1].label[210] );
tran (\labels[1][220] , \labels[1].label[211] );
tran (\labels[1][221] , \labels[1].label[212] );
tran (\labels[1][222] , \labels[1].label[213] );
tran (\labels[1][223] , \labels[1].label[214] );
tran (\labels[1][224] , \labels[1].label[215] );
tran (\labels[1][225] , \labels[1].label[216] );
tran (\labels[1][226] , \labels[1].label[217] );
tran (\labels[1][227] , \labels[1].label[218] );
tran (\labels[1][228] , \labels[1].label[219] );
tran (\labels[1][229] , \labels[1].label[220] );
tran (\labels[1][230] , \labels[1].label[221] );
tran (\labels[1][231] , \labels[1].label[222] );
tran (\labels[1][232] , \labels[1].label[223] );
tran (\labels[1][233] , \labels[1].label[224] );
tran (\labels[1][234] , \labels[1].label[225] );
tran (\labels[1][235] , \labels[1].label[226] );
tran (\labels[1][236] , \labels[1].label[227] );
tran (\labels[1][237] , \labels[1].label[228] );
tran (\labels[1][238] , \labels[1].label[229] );
tran (\labels[1][239] , \labels[1].label[230] );
tran (\labels[1][240] , \labels[1].label[231] );
tran (\labels[1][241] , \labels[1].label[232] );
tran (\labels[1][242] , \labels[1].label[233] );
tran (\labels[1][243] , \labels[1].label[234] );
tran (\labels[1][244] , \labels[1].label[235] );
tran (\labels[1][245] , \labels[1].label[236] );
tran (\labels[1][246] , \labels[1].label[237] );
tran (\labels[1][247] , \labels[1].label[238] );
tran (\labels[1][248] , \labels[1].label[239] );
tran (\labels[1][249] , \labels[1].label[240] );
tran (\labels[1][250] , \labels[1].label[241] );
tran (\labels[1][251] , \labels[1].label[242] );
tran (\labels[1][252] , \labels[1].label[243] );
tran (\labels[1][253] , \labels[1].label[244] );
tran (\labels[1][254] , \labels[1].label[245] );
tran (\labels[1][255] , \labels[1].label[246] );
tran (\labels[1][256] , \labels[1].label[247] );
tran (\labels[1][257] , \labels[1].label[248] );
tran (\labels[1][258] , \labels[1].label[249] );
tran (\labels[1][259] , \labels[1].label[250] );
tran (\labels[1][260] , \labels[1].label[251] );
tran (\labels[1][261] , \labels[1].label[252] );
tran (\labels[1][262] , \labels[1].label[253] );
tran (\labels[1][263] , \labels[1].label[254] );
tran (\labels[1][264] , \labels[1].label[255] );
tran (\labels[1][265] , \labels[1].label_size[0] );
tran (\labels[1][266] , \labels[1].label_size[1] );
tran (\labels[1][267] , \labels[1].label_size[2] );
tran (\labels[1][268] , \labels[1].label_size[3] );
tran (\labels[1][269] , \labels[1].label_size[4] );
tran (\labels[1][270] , \labels[1].label_size[5] );
tran (\labels[1][271] , \labels[1].guid_size[0] );
tran (\labels[2][0] , \labels[2].delimiter[0] );
tran (\labels[2][1] , \labels[2].delimiter[1] );
tran (\labels[2][2] , \labels[2].delimiter[2] );
tran (\labels[2][3] , \labels[2].delimiter[3] );
tran (\labels[2][4] , \labels[2].delimiter[4] );
tran (\labels[2][5] , \labels[2].delimiter[5] );
tran (\labels[2][6] , \labels[2].delimiter[6] );
tran (\labels[2][7] , \labels[2].delimiter[7] );
tran (\labels[2][8] , \labels[2].delimiter_valid[0] );
tran (\labels[2][9] , \labels[2].label[0] );
tran (\labels[2][10] , \labels[2].label[1] );
tran (\labels[2][11] , \labels[2].label[2] );
tran (\labels[2][12] , \labels[2].label[3] );
tran (\labels[2][13] , \labels[2].label[4] );
tran (\labels[2][14] , \labels[2].label[5] );
tran (\labels[2][15] , \labels[2].label[6] );
tran (\labels[2][16] , \labels[2].label[7] );
tran (\labels[2][17] , \labels[2].label[8] );
tran (\labels[2][18] , \labels[2].label[9] );
tran (\labels[2][19] , \labels[2].label[10] );
tran (\labels[2][20] , \labels[2].label[11] );
tran (\labels[2][21] , \labels[2].label[12] );
tran (\labels[2][22] , \labels[2].label[13] );
tran (\labels[2][23] , \labels[2].label[14] );
tran (\labels[2][24] , \labels[2].label[15] );
tran (\labels[2][25] , \labels[2].label[16] );
tran (\labels[2][26] , \labels[2].label[17] );
tran (\labels[2][27] , \labels[2].label[18] );
tran (\labels[2][28] , \labels[2].label[19] );
tran (\labels[2][29] , \labels[2].label[20] );
tran (\labels[2][30] , \labels[2].label[21] );
tran (\labels[2][31] , \labels[2].label[22] );
tran (\labels[2][32] , \labels[2].label[23] );
tran (\labels[2][33] , \labels[2].label[24] );
tran (\labels[2][34] , \labels[2].label[25] );
tran (\labels[2][35] , \labels[2].label[26] );
tran (\labels[2][36] , \labels[2].label[27] );
tran (\labels[2][37] , \labels[2].label[28] );
tran (\labels[2][38] , \labels[2].label[29] );
tran (\labels[2][39] , \labels[2].label[30] );
tran (\labels[2][40] , \labels[2].label[31] );
tran (\labels[2][41] , \labels[2].label[32] );
tran (\labels[2][42] , \labels[2].label[33] );
tran (\labels[2][43] , \labels[2].label[34] );
tran (\labels[2][44] , \labels[2].label[35] );
tran (\labels[2][45] , \labels[2].label[36] );
tran (\labels[2][46] , \labels[2].label[37] );
tran (\labels[2][47] , \labels[2].label[38] );
tran (\labels[2][48] , \labels[2].label[39] );
tran (\labels[2][49] , \labels[2].label[40] );
tran (\labels[2][50] , \labels[2].label[41] );
tran (\labels[2][51] , \labels[2].label[42] );
tran (\labels[2][52] , \labels[2].label[43] );
tran (\labels[2][53] , \labels[2].label[44] );
tran (\labels[2][54] , \labels[2].label[45] );
tran (\labels[2][55] , \labels[2].label[46] );
tran (\labels[2][56] , \labels[2].label[47] );
tran (\labels[2][57] , \labels[2].label[48] );
tran (\labels[2][58] , \labels[2].label[49] );
tran (\labels[2][59] , \labels[2].label[50] );
tran (\labels[2][60] , \labels[2].label[51] );
tran (\labels[2][61] , \labels[2].label[52] );
tran (\labels[2][62] , \labels[2].label[53] );
tran (\labels[2][63] , \labels[2].label[54] );
tran (\labels[2][64] , \labels[2].label[55] );
tran (\labels[2][65] , \labels[2].label[56] );
tran (\labels[2][66] , \labels[2].label[57] );
tran (\labels[2][67] , \labels[2].label[58] );
tran (\labels[2][68] , \labels[2].label[59] );
tran (\labels[2][69] , \labels[2].label[60] );
tran (\labels[2][70] , \labels[2].label[61] );
tran (\labels[2][71] , \labels[2].label[62] );
tran (\labels[2][72] , \labels[2].label[63] );
tran (\labels[2][73] , \labels[2].label[64] );
tran (\labels[2][74] , \labels[2].label[65] );
tran (\labels[2][75] , \labels[2].label[66] );
tran (\labels[2][76] , \labels[2].label[67] );
tran (\labels[2][77] , \labels[2].label[68] );
tran (\labels[2][78] , \labels[2].label[69] );
tran (\labels[2][79] , \labels[2].label[70] );
tran (\labels[2][80] , \labels[2].label[71] );
tran (\labels[2][81] , \labels[2].label[72] );
tran (\labels[2][82] , \labels[2].label[73] );
tran (\labels[2][83] , \labels[2].label[74] );
tran (\labels[2][84] , \labels[2].label[75] );
tran (\labels[2][85] , \labels[2].label[76] );
tran (\labels[2][86] , \labels[2].label[77] );
tran (\labels[2][87] , \labels[2].label[78] );
tran (\labels[2][88] , \labels[2].label[79] );
tran (\labels[2][89] , \labels[2].label[80] );
tran (\labels[2][90] , \labels[2].label[81] );
tran (\labels[2][91] , \labels[2].label[82] );
tran (\labels[2][92] , \labels[2].label[83] );
tran (\labels[2][93] , \labels[2].label[84] );
tran (\labels[2][94] , \labels[2].label[85] );
tran (\labels[2][95] , \labels[2].label[86] );
tran (\labels[2][96] , \labels[2].label[87] );
tran (\labels[2][97] , \labels[2].label[88] );
tran (\labels[2][98] , \labels[2].label[89] );
tran (\labels[2][99] , \labels[2].label[90] );
tran (\labels[2][100] , \labels[2].label[91] );
tran (\labels[2][101] , \labels[2].label[92] );
tran (\labels[2][102] , \labels[2].label[93] );
tran (\labels[2][103] , \labels[2].label[94] );
tran (\labels[2][104] , \labels[2].label[95] );
tran (\labels[2][105] , \labels[2].label[96] );
tran (\labels[2][106] , \labels[2].label[97] );
tran (\labels[2][107] , \labels[2].label[98] );
tran (\labels[2][108] , \labels[2].label[99] );
tran (\labels[2][109] , \labels[2].label[100] );
tran (\labels[2][110] , \labels[2].label[101] );
tran (\labels[2][111] , \labels[2].label[102] );
tran (\labels[2][112] , \labels[2].label[103] );
tran (\labels[2][113] , \labels[2].label[104] );
tran (\labels[2][114] , \labels[2].label[105] );
tran (\labels[2][115] , \labels[2].label[106] );
tran (\labels[2][116] , \labels[2].label[107] );
tran (\labels[2][117] , \labels[2].label[108] );
tran (\labels[2][118] , \labels[2].label[109] );
tran (\labels[2][119] , \labels[2].label[110] );
tran (\labels[2][120] , \labels[2].label[111] );
tran (\labels[2][121] , \labels[2].label[112] );
tran (\labels[2][122] , \labels[2].label[113] );
tran (\labels[2][123] , \labels[2].label[114] );
tran (\labels[2][124] , \labels[2].label[115] );
tran (\labels[2][125] , \labels[2].label[116] );
tran (\labels[2][126] , \labels[2].label[117] );
tran (\labels[2][127] , \labels[2].label[118] );
tran (\labels[2][128] , \labels[2].label[119] );
tran (\labels[2][129] , \labels[2].label[120] );
tran (\labels[2][130] , \labels[2].label[121] );
tran (\labels[2][131] , \labels[2].label[122] );
tran (\labels[2][132] , \labels[2].label[123] );
tran (\labels[2][133] , \labels[2].label[124] );
tran (\labels[2][134] , \labels[2].label[125] );
tran (\labels[2][135] , \labels[2].label[126] );
tran (\labels[2][136] , \labels[2].label[127] );
tran (\labels[2][137] , \labels[2].label[128] );
tran (\labels[2][138] , \labels[2].label[129] );
tran (\labels[2][139] , \labels[2].label[130] );
tran (\labels[2][140] , \labels[2].label[131] );
tran (\labels[2][141] , \labels[2].label[132] );
tran (\labels[2][142] , \labels[2].label[133] );
tran (\labels[2][143] , \labels[2].label[134] );
tran (\labels[2][144] , \labels[2].label[135] );
tran (\labels[2][145] , \labels[2].label[136] );
tran (\labels[2][146] , \labels[2].label[137] );
tran (\labels[2][147] , \labels[2].label[138] );
tran (\labels[2][148] , \labels[2].label[139] );
tran (\labels[2][149] , \labels[2].label[140] );
tran (\labels[2][150] , \labels[2].label[141] );
tran (\labels[2][151] , \labels[2].label[142] );
tran (\labels[2][152] , \labels[2].label[143] );
tran (\labels[2][153] , \labels[2].label[144] );
tran (\labels[2][154] , \labels[2].label[145] );
tran (\labels[2][155] , \labels[2].label[146] );
tran (\labels[2][156] , \labels[2].label[147] );
tran (\labels[2][157] , \labels[2].label[148] );
tran (\labels[2][158] , \labels[2].label[149] );
tran (\labels[2][159] , \labels[2].label[150] );
tran (\labels[2][160] , \labels[2].label[151] );
tran (\labels[2][161] , \labels[2].label[152] );
tran (\labels[2][162] , \labels[2].label[153] );
tran (\labels[2][163] , \labels[2].label[154] );
tran (\labels[2][164] , \labels[2].label[155] );
tran (\labels[2][165] , \labels[2].label[156] );
tran (\labels[2][166] , \labels[2].label[157] );
tran (\labels[2][167] , \labels[2].label[158] );
tran (\labels[2][168] , \labels[2].label[159] );
tran (\labels[2][169] , \labels[2].label[160] );
tran (\labels[2][170] , \labels[2].label[161] );
tran (\labels[2][171] , \labels[2].label[162] );
tran (\labels[2][172] , \labels[2].label[163] );
tran (\labels[2][173] , \labels[2].label[164] );
tran (\labels[2][174] , \labels[2].label[165] );
tran (\labels[2][175] , \labels[2].label[166] );
tran (\labels[2][176] , \labels[2].label[167] );
tran (\labels[2][177] , \labels[2].label[168] );
tran (\labels[2][178] , \labels[2].label[169] );
tran (\labels[2][179] , \labels[2].label[170] );
tran (\labels[2][180] , \labels[2].label[171] );
tran (\labels[2][181] , \labels[2].label[172] );
tran (\labels[2][182] , \labels[2].label[173] );
tran (\labels[2][183] , \labels[2].label[174] );
tran (\labels[2][184] , \labels[2].label[175] );
tran (\labels[2][185] , \labels[2].label[176] );
tran (\labels[2][186] , \labels[2].label[177] );
tran (\labels[2][187] , \labels[2].label[178] );
tran (\labels[2][188] , \labels[2].label[179] );
tran (\labels[2][189] , \labels[2].label[180] );
tran (\labels[2][190] , \labels[2].label[181] );
tran (\labels[2][191] , \labels[2].label[182] );
tran (\labels[2][192] , \labels[2].label[183] );
tran (\labels[2][193] , \labels[2].label[184] );
tran (\labels[2][194] , \labels[2].label[185] );
tran (\labels[2][195] , \labels[2].label[186] );
tran (\labels[2][196] , \labels[2].label[187] );
tran (\labels[2][197] , \labels[2].label[188] );
tran (\labels[2][198] , \labels[2].label[189] );
tran (\labels[2][199] , \labels[2].label[190] );
tran (\labels[2][200] , \labels[2].label[191] );
tran (\labels[2][201] , \labels[2].label[192] );
tran (\labels[2][202] , \labels[2].label[193] );
tran (\labels[2][203] , \labels[2].label[194] );
tran (\labels[2][204] , \labels[2].label[195] );
tran (\labels[2][205] , \labels[2].label[196] );
tran (\labels[2][206] , \labels[2].label[197] );
tran (\labels[2][207] , \labels[2].label[198] );
tran (\labels[2][208] , \labels[2].label[199] );
tran (\labels[2][209] , \labels[2].label[200] );
tran (\labels[2][210] , \labels[2].label[201] );
tran (\labels[2][211] , \labels[2].label[202] );
tran (\labels[2][212] , \labels[2].label[203] );
tran (\labels[2][213] , \labels[2].label[204] );
tran (\labels[2][214] , \labels[2].label[205] );
tran (\labels[2][215] , \labels[2].label[206] );
tran (\labels[2][216] , \labels[2].label[207] );
tran (\labels[2][217] , \labels[2].label[208] );
tran (\labels[2][218] , \labels[2].label[209] );
tran (\labels[2][219] , \labels[2].label[210] );
tran (\labels[2][220] , \labels[2].label[211] );
tran (\labels[2][221] , \labels[2].label[212] );
tran (\labels[2][222] , \labels[2].label[213] );
tran (\labels[2][223] , \labels[2].label[214] );
tran (\labels[2][224] , \labels[2].label[215] );
tran (\labels[2][225] , \labels[2].label[216] );
tran (\labels[2][226] , \labels[2].label[217] );
tran (\labels[2][227] , \labels[2].label[218] );
tran (\labels[2][228] , \labels[2].label[219] );
tran (\labels[2][229] , \labels[2].label[220] );
tran (\labels[2][230] , \labels[2].label[221] );
tran (\labels[2][231] , \labels[2].label[222] );
tran (\labels[2][232] , \labels[2].label[223] );
tran (\labels[2][233] , \labels[2].label[224] );
tran (\labels[2][234] , \labels[2].label[225] );
tran (\labels[2][235] , \labels[2].label[226] );
tran (\labels[2][236] , \labels[2].label[227] );
tran (\labels[2][237] , \labels[2].label[228] );
tran (\labels[2][238] , \labels[2].label[229] );
tran (\labels[2][239] , \labels[2].label[230] );
tran (\labels[2][240] , \labels[2].label[231] );
tran (\labels[2][241] , \labels[2].label[232] );
tran (\labels[2][242] , \labels[2].label[233] );
tran (\labels[2][243] , \labels[2].label[234] );
tran (\labels[2][244] , \labels[2].label[235] );
tran (\labels[2][245] , \labels[2].label[236] );
tran (\labels[2][246] , \labels[2].label[237] );
tran (\labels[2][247] , \labels[2].label[238] );
tran (\labels[2][248] , \labels[2].label[239] );
tran (\labels[2][249] , \labels[2].label[240] );
tran (\labels[2][250] , \labels[2].label[241] );
tran (\labels[2][251] , \labels[2].label[242] );
tran (\labels[2][252] , \labels[2].label[243] );
tran (\labels[2][253] , \labels[2].label[244] );
tran (\labels[2][254] , \labels[2].label[245] );
tran (\labels[2][255] , \labels[2].label[246] );
tran (\labels[2][256] , \labels[2].label[247] );
tran (\labels[2][257] , \labels[2].label[248] );
tran (\labels[2][258] , \labels[2].label[249] );
tran (\labels[2][259] , \labels[2].label[250] );
tran (\labels[2][260] , \labels[2].label[251] );
tran (\labels[2][261] , \labels[2].label[252] );
tran (\labels[2][262] , \labels[2].label[253] );
tran (\labels[2][263] , \labels[2].label[254] );
tran (\labels[2][264] , \labels[2].label[255] );
tran (\labels[2][265] , \labels[2].label_size[0] );
tran (\labels[2][266] , \labels[2].label_size[1] );
tran (\labels[2][267] , \labels[2].label_size[2] );
tran (\labels[2][268] , \labels[2].label_size[3] );
tran (\labels[2][269] , \labels[2].label_size[4] );
tran (\labels[2][270] , \labels[2].label_size[5] );
tran (\labels[2][271] , \labels[2].guid_size[0] );
tran (\labels[3][0] , \labels[3].delimiter[0] );
tran (\labels[3][1] , \labels[3].delimiter[1] );
tran (\labels[3][2] , \labels[3].delimiter[2] );
tran (\labels[3][3] , \labels[3].delimiter[3] );
tran (\labels[3][4] , \labels[3].delimiter[4] );
tran (\labels[3][5] , \labels[3].delimiter[5] );
tran (\labels[3][6] , \labels[3].delimiter[6] );
tran (\labels[3][7] , \labels[3].delimiter[7] );
tran (\labels[3][8] , \labels[3].delimiter_valid[0] );
tran (\labels[3][9] , \labels[3].label[0] );
tran (\labels[3][10] , \labels[3].label[1] );
tran (\labels[3][11] , \labels[3].label[2] );
tran (\labels[3][12] , \labels[3].label[3] );
tran (\labels[3][13] , \labels[3].label[4] );
tran (\labels[3][14] , \labels[3].label[5] );
tran (\labels[3][15] , \labels[3].label[6] );
tran (\labels[3][16] , \labels[3].label[7] );
tran (\labels[3][17] , \labels[3].label[8] );
tran (\labels[3][18] , \labels[3].label[9] );
tran (\labels[3][19] , \labels[3].label[10] );
tran (\labels[3][20] , \labels[3].label[11] );
tran (\labels[3][21] , \labels[3].label[12] );
tran (\labels[3][22] , \labels[3].label[13] );
tran (\labels[3][23] , \labels[3].label[14] );
tran (\labels[3][24] , \labels[3].label[15] );
tran (\labels[3][25] , \labels[3].label[16] );
tran (\labels[3][26] , \labels[3].label[17] );
tran (\labels[3][27] , \labels[3].label[18] );
tran (\labels[3][28] , \labels[3].label[19] );
tran (\labels[3][29] , \labels[3].label[20] );
tran (\labels[3][30] , \labels[3].label[21] );
tran (\labels[3][31] , \labels[3].label[22] );
tran (\labels[3][32] , \labels[3].label[23] );
tran (\labels[3][33] , \labels[3].label[24] );
tran (\labels[3][34] , \labels[3].label[25] );
tran (\labels[3][35] , \labels[3].label[26] );
tran (\labels[3][36] , \labels[3].label[27] );
tran (\labels[3][37] , \labels[3].label[28] );
tran (\labels[3][38] , \labels[3].label[29] );
tran (\labels[3][39] , \labels[3].label[30] );
tran (\labels[3][40] , \labels[3].label[31] );
tran (\labels[3][41] , \labels[3].label[32] );
tran (\labels[3][42] , \labels[3].label[33] );
tran (\labels[3][43] , \labels[3].label[34] );
tran (\labels[3][44] , \labels[3].label[35] );
tran (\labels[3][45] , \labels[3].label[36] );
tran (\labels[3][46] , \labels[3].label[37] );
tran (\labels[3][47] , \labels[3].label[38] );
tran (\labels[3][48] , \labels[3].label[39] );
tran (\labels[3][49] , \labels[3].label[40] );
tran (\labels[3][50] , \labels[3].label[41] );
tran (\labels[3][51] , \labels[3].label[42] );
tran (\labels[3][52] , \labels[3].label[43] );
tran (\labels[3][53] , \labels[3].label[44] );
tran (\labels[3][54] , \labels[3].label[45] );
tran (\labels[3][55] , \labels[3].label[46] );
tran (\labels[3][56] , \labels[3].label[47] );
tran (\labels[3][57] , \labels[3].label[48] );
tran (\labels[3][58] , \labels[3].label[49] );
tran (\labels[3][59] , \labels[3].label[50] );
tran (\labels[3][60] , \labels[3].label[51] );
tran (\labels[3][61] , \labels[3].label[52] );
tran (\labels[3][62] , \labels[3].label[53] );
tran (\labels[3][63] , \labels[3].label[54] );
tran (\labels[3][64] , \labels[3].label[55] );
tran (\labels[3][65] , \labels[3].label[56] );
tran (\labels[3][66] , \labels[3].label[57] );
tran (\labels[3][67] , \labels[3].label[58] );
tran (\labels[3][68] , \labels[3].label[59] );
tran (\labels[3][69] , \labels[3].label[60] );
tran (\labels[3][70] , \labels[3].label[61] );
tran (\labels[3][71] , \labels[3].label[62] );
tran (\labels[3][72] , \labels[3].label[63] );
tran (\labels[3][73] , \labels[3].label[64] );
tran (\labels[3][74] , \labels[3].label[65] );
tran (\labels[3][75] , \labels[3].label[66] );
tran (\labels[3][76] , \labels[3].label[67] );
tran (\labels[3][77] , \labels[3].label[68] );
tran (\labels[3][78] , \labels[3].label[69] );
tran (\labels[3][79] , \labels[3].label[70] );
tran (\labels[3][80] , \labels[3].label[71] );
tran (\labels[3][81] , \labels[3].label[72] );
tran (\labels[3][82] , \labels[3].label[73] );
tran (\labels[3][83] , \labels[3].label[74] );
tran (\labels[3][84] , \labels[3].label[75] );
tran (\labels[3][85] , \labels[3].label[76] );
tran (\labels[3][86] , \labels[3].label[77] );
tran (\labels[3][87] , \labels[3].label[78] );
tran (\labels[3][88] , \labels[3].label[79] );
tran (\labels[3][89] , \labels[3].label[80] );
tran (\labels[3][90] , \labels[3].label[81] );
tran (\labels[3][91] , \labels[3].label[82] );
tran (\labels[3][92] , \labels[3].label[83] );
tran (\labels[3][93] , \labels[3].label[84] );
tran (\labels[3][94] , \labels[3].label[85] );
tran (\labels[3][95] , \labels[3].label[86] );
tran (\labels[3][96] , \labels[3].label[87] );
tran (\labels[3][97] , \labels[3].label[88] );
tran (\labels[3][98] , \labels[3].label[89] );
tran (\labels[3][99] , \labels[3].label[90] );
tran (\labels[3][100] , \labels[3].label[91] );
tran (\labels[3][101] , \labels[3].label[92] );
tran (\labels[3][102] , \labels[3].label[93] );
tran (\labels[3][103] , \labels[3].label[94] );
tran (\labels[3][104] , \labels[3].label[95] );
tran (\labels[3][105] , \labels[3].label[96] );
tran (\labels[3][106] , \labels[3].label[97] );
tran (\labels[3][107] , \labels[3].label[98] );
tran (\labels[3][108] , \labels[3].label[99] );
tran (\labels[3][109] , \labels[3].label[100] );
tran (\labels[3][110] , \labels[3].label[101] );
tran (\labels[3][111] , \labels[3].label[102] );
tran (\labels[3][112] , \labels[3].label[103] );
tran (\labels[3][113] , \labels[3].label[104] );
tran (\labels[3][114] , \labels[3].label[105] );
tran (\labels[3][115] , \labels[3].label[106] );
tran (\labels[3][116] , \labels[3].label[107] );
tran (\labels[3][117] , \labels[3].label[108] );
tran (\labels[3][118] , \labels[3].label[109] );
tran (\labels[3][119] , \labels[3].label[110] );
tran (\labels[3][120] , \labels[3].label[111] );
tran (\labels[3][121] , \labels[3].label[112] );
tran (\labels[3][122] , \labels[3].label[113] );
tran (\labels[3][123] , \labels[3].label[114] );
tran (\labels[3][124] , \labels[3].label[115] );
tran (\labels[3][125] , \labels[3].label[116] );
tran (\labels[3][126] , \labels[3].label[117] );
tran (\labels[3][127] , \labels[3].label[118] );
tran (\labels[3][128] , \labels[3].label[119] );
tran (\labels[3][129] , \labels[3].label[120] );
tran (\labels[3][130] , \labels[3].label[121] );
tran (\labels[3][131] , \labels[3].label[122] );
tran (\labels[3][132] , \labels[3].label[123] );
tran (\labels[3][133] , \labels[3].label[124] );
tran (\labels[3][134] , \labels[3].label[125] );
tran (\labels[3][135] , \labels[3].label[126] );
tran (\labels[3][136] , \labels[3].label[127] );
tran (\labels[3][137] , \labels[3].label[128] );
tran (\labels[3][138] , \labels[3].label[129] );
tran (\labels[3][139] , \labels[3].label[130] );
tran (\labels[3][140] , \labels[3].label[131] );
tran (\labels[3][141] , \labels[3].label[132] );
tran (\labels[3][142] , \labels[3].label[133] );
tran (\labels[3][143] , \labels[3].label[134] );
tran (\labels[3][144] , \labels[3].label[135] );
tran (\labels[3][145] , \labels[3].label[136] );
tran (\labels[3][146] , \labels[3].label[137] );
tran (\labels[3][147] , \labels[3].label[138] );
tran (\labels[3][148] , \labels[3].label[139] );
tran (\labels[3][149] , \labels[3].label[140] );
tran (\labels[3][150] , \labels[3].label[141] );
tran (\labels[3][151] , \labels[3].label[142] );
tran (\labels[3][152] , \labels[3].label[143] );
tran (\labels[3][153] , \labels[3].label[144] );
tran (\labels[3][154] , \labels[3].label[145] );
tran (\labels[3][155] , \labels[3].label[146] );
tran (\labels[3][156] , \labels[3].label[147] );
tran (\labels[3][157] , \labels[3].label[148] );
tran (\labels[3][158] , \labels[3].label[149] );
tran (\labels[3][159] , \labels[3].label[150] );
tran (\labels[3][160] , \labels[3].label[151] );
tran (\labels[3][161] , \labels[3].label[152] );
tran (\labels[3][162] , \labels[3].label[153] );
tran (\labels[3][163] , \labels[3].label[154] );
tran (\labels[3][164] , \labels[3].label[155] );
tran (\labels[3][165] , \labels[3].label[156] );
tran (\labels[3][166] , \labels[3].label[157] );
tran (\labels[3][167] , \labels[3].label[158] );
tran (\labels[3][168] , \labels[3].label[159] );
tran (\labels[3][169] , \labels[3].label[160] );
tran (\labels[3][170] , \labels[3].label[161] );
tran (\labels[3][171] , \labels[3].label[162] );
tran (\labels[3][172] , \labels[3].label[163] );
tran (\labels[3][173] , \labels[3].label[164] );
tran (\labels[3][174] , \labels[3].label[165] );
tran (\labels[3][175] , \labels[3].label[166] );
tran (\labels[3][176] , \labels[3].label[167] );
tran (\labels[3][177] , \labels[3].label[168] );
tran (\labels[3][178] , \labels[3].label[169] );
tran (\labels[3][179] , \labels[3].label[170] );
tran (\labels[3][180] , \labels[3].label[171] );
tran (\labels[3][181] , \labels[3].label[172] );
tran (\labels[3][182] , \labels[3].label[173] );
tran (\labels[3][183] , \labels[3].label[174] );
tran (\labels[3][184] , \labels[3].label[175] );
tran (\labels[3][185] , \labels[3].label[176] );
tran (\labels[3][186] , \labels[3].label[177] );
tran (\labels[3][187] , \labels[3].label[178] );
tran (\labels[3][188] , \labels[3].label[179] );
tran (\labels[3][189] , \labels[3].label[180] );
tran (\labels[3][190] , \labels[3].label[181] );
tran (\labels[3][191] , \labels[3].label[182] );
tran (\labels[3][192] , \labels[3].label[183] );
tran (\labels[3][193] , \labels[3].label[184] );
tran (\labels[3][194] , \labels[3].label[185] );
tran (\labels[3][195] , \labels[3].label[186] );
tran (\labels[3][196] , \labels[3].label[187] );
tran (\labels[3][197] , \labels[3].label[188] );
tran (\labels[3][198] , \labels[3].label[189] );
tran (\labels[3][199] , \labels[3].label[190] );
tran (\labels[3][200] , \labels[3].label[191] );
tran (\labels[3][201] , \labels[3].label[192] );
tran (\labels[3][202] , \labels[3].label[193] );
tran (\labels[3][203] , \labels[3].label[194] );
tran (\labels[3][204] , \labels[3].label[195] );
tran (\labels[3][205] , \labels[3].label[196] );
tran (\labels[3][206] , \labels[3].label[197] );
tran (\labels[3][207] , \labels[3].label[198] );
tran (\labels[3][208] , \labels[3].label[199] );
tran (\labels[3][209] , \labels[3].label[200] );
tran (\labels[3][210] , \labels[3].label[201] );
tran (\labels[3][211] , \labels[3].label[202] );
tran (\labels[3][212] , \labels[3].label[203] );
tran (\labels[3][213] , \labels[3].label[204] );
tran (\labels[3][214] , \labels[3].label[205] );
tran (\labels[3][215] , \labels[3].label[206] );
tran (\labels[3][216] , \labels[3].label[207] );
tran (\labels[3][217] , \labels[3].label[208] );
tran (\labels[3][218] , \labels[3].label[209] );
tran (\labels[3][219] , \labels[3].label[210] );
tran (\labels[3][220] , \labels[3].label[211] );
tran (\labels[3][221] , \labels[3].label[212] );
tran (\labels[3][222] , \labels[3].label[213] );
tran (\labels[3][223] , \labels[3].label[214] );
tran (\labels[3][224] , \labels[3].label[215] );
tran (\labels[3][225] , \labels[3].label[216] );
tran (\labels[3][226] , \labels[3].label[217] );
tran (\labels[3][227] , \labels[3].label[218] );
tran (\labels[3][228] , \labels[3].label[219] );
tran (\labels[3][229] , \labels[3].label[220] );
tran (\labels[3][230] , \labels[3].label[221] );
tran (\labels[3][231] , \labels[3].label[222] );
tran (\labels[3][232] , \labels[3].label[223] );
tran (\labels[3][233] , \labels[3].label[224] );
tran (\labels[3][234] , \labels[3].label[225] );
tran (\labels[3][235] , \labels[3].label[226] );
tran (\labels[3][236] , \labels[3].label[227] );
tran (\labels[3][237] , \labels[3].label[228] );
tran (\labels[3][238] , \labels[3].label[229] );
tran (\labels[3][239] , \labels[3].label[230] );
tran (\labels[3][240] , \labels[3].label[231] );
tran (\labels[3][241] , \labels[3].label[232] );
tran (\labels[3][242] , \labels[3].label[233] );
tran (\labels[3][243] , \labels[3].label[234] );
tran (\labels[3][244] , \labels[3].label[235] );
tran (\labels[3][245] , \labels[3].label[236] );
tran (\labels[3][246] , \labels[3].label[237] );
tran (\labels[3][247] , \labels[3].label[238] );
tran (\labels[3][248] , \labels[3].label[239] );
tran (\labels[3][249] , \labels[3].label[240] );
tran (\labels[3][250] , \labels[3].label[241] );
tran (\labels[3][251] , \labels[3].label[242] );
tran (\labels[3][252] , \labels[3].label[243] );
tran (\labels[3][253] , \labels[3].label[244] );
tran (\labels[3][254] , \labels[3].label[245] );
tran (\labels[3][255] , \labels[3].label[246] );
tran (\labels[3][256] , \labels[3].label[247] );
tran (\labels[3][257] , \labels[3].label[248] );
tran (\labels[3][258] , \labels[3].label[249] );
tran (\labels[3][259] , \labels[3].label[250] );
tran (\labels[3][260] , \labels[3].label[251] );
tran (\labels[3][261] , \labels[3].label[252] );
tran (\labels[3][262] , \labels[3].label[253] );
tran (\labels[3][263] , \labels[3].label[254] );
tran (\labels[3][264] , \labels[3].label[255] );
tran (\labels[3][265] , \labels[3].label_size[0] );
tran (\labels[3][266] , \labels[3].label_size[1] );
tran (\labels[3][267] , \labels[3].label_size[2] );
tran (\labels[3][268] , \labels[3].label_size[3] );
tran (\labels[3][269] , \labels[3].label_size[4] );
tran (\labels[3][270] , \labels[3].label_size[5] );
tran (\labels[3][271] , \labels[3].guid_size[0] );
tran (\labels[4][0] , \labels[4].delimiter[0] );
tran (\labels[4][1] , \labels[4].delimiter[1] );
tran (\labels[4][2] , \labels[4].delimiter[2] );
tran (\labels[4][3] , \labels[4].delimiter[3] );
tran (\labels[4][4] , \labels[4].delimiter[4] );
tran (\labels[4][5] , \labels[4].delimiter[5] );
tran (\labels[4][6] , \labels[4].delimiter[6] );
tran (\labels[4][7] , \labels[4].delimiter[7] );
tran (\labels[4][8] , \labels[4].delimiter_valid[0] );
tran (\labels[4][9] , \labels[4].label[0] );
tran (\labels[4][10] , \labels[4].label[1] );
tran (\labels[4][11] , \labels[4].label[2] );
tran (\labels[4][12] , \labels[4].label[3] );
tran (\labels[4][13] , \labels[4].label[4] );
tran (\labels[4][14] , \labels[4].label[5] );
tran (\labels[4][15] , \labels[4].label[6] );
tran (\labels[4][16] , \labels[4].label[7] );
tran (\labels[4][17] , \labels[4].label[8] );
tran (\labels[4][18] , \labels[4].label[9] );
tran (\labels[4][19] , \labels[4].label[10] );
tran (\labels[4][20] , \labels[4].label[11] );
tran (\labels[4][21] , \labels[4].label[12] );
tran (\labels[4][22] , \labels[4].label[13] );
tran (\labels[4][23] , \labels[4].label[14] );
tran (\labels[4][24] , \labels[4].label[15] );
tran (\labels[4][25] , \labels[4].label[16] );
tran (\labels[4][26] , \labels[4].label[17] );
tran (\labels[4][27] , \labels[4].label[18] );
tran (\labels[4][28] , \labels[4].label[19] );
tran (\labels[4][29] , \labels[4].label[20] );
tran (\labels[4][30] , \labels[4].label[21] );
tran (\labels[4][31] , \labels[4].label[22] );
tran (\labels[4][32] , \labels[4].label[23] );
tran (\labels[4][33] , \labels[4].label[24] );
tran (\labels[4][34] , \labels[4].label[25] );
tran (\labels[4][35] , \labels[4].label[26] );
tran (\labels[4][36] , \labels[4].label[27] );
tran (\labels[4][37] , \labels[4].label[28] );
tran (\labels[4][38] , \labels[4].label[29] );
tran (\labels[4][39] , \labels[4].label[30] );
tran (\labels[4][40] , \labels[4].label[31] );
tran (\labels[4][41] , \labels[4].label[32] );
tran (\labels[4][42] , \labels[4].label[33] );
tran (\labels[4][43] , \labels[4].label[34] );
tran (\labels[4][44] , \labels[4].label[35] );
tran (\labels[4][45] , \labels[4].label[36] );
tran (\labels[4][46] , \labels[4].label[37] );
tran (\labels[4][47] , \labels[4].label[38] );
tran (\labels[4][48] , \labels[4].label[39] );
tran (\labels[4][49] , \labels[4].label[40] );
tran (\labels[4][50] , \labels[4].label[41] );
tran (\labels[4][51] , \labels[4].label[42] );
tran (\labels[4][52] , \labels[4].label[43] );
tran (\labels[4][53] , \labels[4].label[44] );
tran (\labels[4][54] , \labels[4].label[45] );
tran (\labels[4][55] , \labels[4].label[46] );
tran (\labels[4][56] , \labels[4].label[47] );
tran (\labels[4][57] , \labels[4].label[48] );
tran (\labels[4][58] , \labels[4].label[49] );
tran (\labels[4][59] , \labels[4].label[50] );
tran (\labels[4][60] , \labels[4].label[51] );
tran (\labels[4][61] , \labels[4].label[52] );
tran (\labels[4][62] , \labels[4].label[53] );
tran (\labels[4][63] , \labels[4].label[54] );
tran (\labels[4][64] , \labels[4].label[55] );
tran (\labels[4][65] , \labels[4].label[56] );
tran (\labels[4][66] , \labels[4].label[57] );
tran (\labels[4][67] , \labels[4].label[58] );
tran (\labels[4][68] , \labels[4].label[59] );
tran (\labels[4][69] , \labels[4].label[60] );
tran (\labels[4][70] , \labels[4].label[61] );
tran (\labels[4][71] , \labels[4].label[62] );
tran (\labels[4][72] , \labels[4].label[63] );
tran (\labels[4][73] , \labels[4].label[64] );
tran (\labels[4][74] , \labels[4].label[65] );
tran (\labels[4][75] , \labels[4].label[66] );
tran (\labels[4][76] , \labels[4].label[67] );
tran (\labels[4][77] , \labels[4].label[68] );
tran (\labels[4][78] , \labels[4].label[69] );
tran (\labels[4][79] , \labels[4].label[70] );
tran (\labels[4][80] , \labels[4].label[71] );
tran (\labels[4][81] , \labels[4].label[72] );
tran (\labels[4][82] , \labels[4].label[73] );
tran (\labels[4][83] , \labels[4].label[74] );
tran (\labels[4][84] , \labels[4].label[75] );
tran (\labels[4][85] , \labels[4].label[76] );
tran (\labels[4][86] , \labels[4].label[77] );
tran (\labels[4][87] , \labels[4].label[78] );
tran (\labels[4][88] , \labels[4].label[79] );
tran (\labels[4][89] , \labels[4].label[80] );
tran (\labels[4][90] , \labels[4].label[81] );
tran (\labels[4][91] , \labels[4].label[82] );
tran (\labels[4][92] , \labels[4].label[83] );
tran (\labels[4][93] , \labels[4].label[84] );
tran (\labels[4][94] , \labels[4].label[85] );
tran (\labels[4][95] , \labels[4].label[86] );
tran (\labels[4][96] , \labels[4].label[87] );
tran (\labels[4][97] , \labels[4].label[88] );
tran (\labels[4][98] , \labels[4].label[89] );
tran (\labels[4][99] , \labels[4].label[90] );
tran (\labels[4][100] , \labels[4].label[91] );
tran (\labels[4][101] , \labels[4].label[92] );
tran (\labels[4][102] , \labels[4].label[93] );
tran (\labels[4][103] , \labels[4].label[94] );
tran (\labels[4][104] , \labels[4].label[95] );
tran (\labels[4][105] , \labels[4].label[96] );
tran (\labels[4][106] , \labels[4].label[97] );
tran (\labels[4][107] , \labels[4].label[98] );
tran (\labels[4][108] , \labels[4].label[99] );
tran (\labels[4][109] , \labels[4].label[100] );
tran (\labels[4][110] , \labels[4].label[101] );
tran (\labels[4][111] , \labels[4].label[102] );
tran (\labels[4][112] , \labels[4].label[103] );
tran (\labels[4][113] , \labels[4].label[104] );
tran (\labels[4][114] , \labels[4].label[105] );
tran (\labels[4][115] , \labels[4].label[106] );
tran (\labels[4][116] , \labels[4].label[107] );
tran (\labels[4][117] , \labels[4].label[108] );
tran (\labels[4][118] , \labels[4].label[109] );
tran (\labels[4][119] , \labels[4].label[110] );
tran (\labels[4][120] , \labels[4].label[111] );
tran (\labels[4][121] , \labels[4].label[112] );
tran (\labels[4][122] , \labels[4].label[113] );
tran (\labels[4][123] , \labels[4].label[114] );
tran (\labels[4][124] , \labels[4].label[115] );
tran (\labels[4][125] , \labels[4].label[116] );
tran (\labels[4][126] , \labels[4].label[117] );
tran (\labels[4][127] , \labels[4].label[118] );
tran (\labels[4][128] , \labels[4].label[119] );
tran (\labels[4][129] , \labels[4].label[120] );
tran (\labels[4][130] , \labels[4].label[121] );
tran (\labels[4][131] , \labels[4].label[122] );
tran (\labels[4][132] , \labels[4].label[123] );
tran (\labels[4][133] , \labels[4].label[124] );
tran (\labels[4][134] , \labels[4].label[125] );
tran (\labels[4][135] , \labels[4].label[126] );
tran (\labels[4][136] , \labels[4].label[127] );
tran (\labels[4][137] , \labels[4].label[128] );
tran (\labels[4][138] , \labels[4].label[129] );
tran (\labels[4][139] , \labels[4].label[130] );
tran (\labels[4][140] , \labels[4].label[131] );
tran (\labels[4][141] , \labels[4].label[132] );
tran (\labels[4][142] , \labels[4].label[133] );
tran (\labels[4][143] , \labels[4].label[134] );
tran (\labels[4][144] , \labels[4].label[135] );
tran (\labels[4][145] , \labels[4].label[136] );
tran (\labels[4][146] , \labels[4].label[137] );
tran (\labels[4][147] , \labels[4].label[138] );
tran (\labels[4][148] , \labels[4].label[139] );
tran (\labels[4][149] , \labels[4].label[140] );
tran (\labels[4][150] , \labels[4].label[141] );
tran (\labels[4][151] , \labels[4].label[142] );
tran (\labels[4][152] , \labels[4].label[143] );
tran (\labels[4][153] , \labels[4].label[144] );
tran (\labels[4][154] , \labels[4].label[145] );
tran (\labels[4][155] , \labels[4].label[146] );
tran (\labels[4][156] , \labels[4].label[147] );
tran (\labels[4][157] , \labels[4].label[148] );
tran (\labels[4][158] , \labels[4].label[149] );
tran (\labels[4][159] , \labels[4].label[150] );
tran (\labels[4][160] , \labels[4].label[151] );
tran (\labels[4][161] , \labels[4].label[152] );
tran (\labels[4][162] , \labels[4].label[153] );
tran (\labels[4][163] , \labels[4].label[154] );
tran (\labels[4][164] , \labels[4].label[155] );
tran (\labels[4][165] , \labels[4].label[156] );
tran (\labels[4][166] , \labels[4].label[157] );
tran (\labels[4][167] , \labels[4].label[158] );
tran (\labels[4][168] , \labels[4].label[159] );
tran (\labels[4][169] , \labels[4].label[160] );
tran (\labels[4][170] , \labels[4].label[161] );
tran (\labels[4][171] , \labels[4].label[162] );
tran (\labels[4][172] , \labels[4].label[163] );
tran (\labels[4][173] , \labels[4].label[164] );
tran (\labels[4][174] , \labels[4].label[165] );
tran (\labels[4][175] , \labels[4].label[166] );
tran (\labels[4][176] , \labels[4].label[167] );
tran (\labels[4][177] , \labels[4].label[168] );
tran (\labels[4][178] , \labels[4].label[169] );
tran (\labels[4][179] , \labels[4].label[170] );
tran (\labels[4][180] , \labels[4].label[171] );
tran (\labels[4][181] , \labels[4].label[172] );
tran (\labels[4][182] , \labels[4].label[173] );
tran (\labels[4][183] , \labels[4].label[174] );
tran (\labels[4][184] , \labels[4].label[175] );
tran (\labels[4][185] , \labels[4].label[176] );
tran (\labels[4][186] , \labels[4].label[177] );
tran (\labels[4][187] , \labels[4].label[178] );
tran (\labels[4][188] , \labels[4].label[179] );
tran (\labels[4][189] , \labels[4].label[180] );
tran (\labels[4][190] , \labels[4].label[181] );
tran (\labels[4][191] , \labels[4].label[182] );
tran (\labels[4][192] , \labels[4].label[183] );
tran (\labels[4][193] , \labels[4].label[184] );
tran (\labels[4][194] , \labels[4].label[185] );
tran (\labels[4][195] , \labels[4].label[186] );
tran (\labels[4][196] , \labels[4].label[187] );
tran (\labels[4][197] , \labels[4].label[188] );
tran (\labels[4][198] , \labels[4].label[189] );
tran (\labels[4][199] , \labels[4].label[190] );
tran (\labels[4][200] , \labels[4].label[191] );
tran (\labels[4][201] , \labels[4].label[192] );
tran (\labels[4][202] , \labels[4].label[193] );
tran (\labels[4][203] , \labels[4].label[194] );
tran (\labels[4][204] , \labels[4].label[195] );
tran (\labels[4][205] , \labels[4].label[196] );
tran (\labels[4][206] , \labels[4].label[197] );
tran (\labels[4][207] , \labels[4].label[198] );
tran (\labels[4][208] , \labels[4].label[199] );
tran (\labels[4][209] , \labels[4].label[200] );
tran (\labels[4][210] , \labels[4].label[201] );
tran (\labels[4][211] , \labels[4].label[202] );
tran (\labels[4][212] , \labels[4].label[203] );
tran (\labels[4][213] , \labels[4].label[204] );
tran (\labels[4][214] , \labels[4].label[205] );
tran (\labels[4][215] , \labels[4].label[206] );
tran (\labels[4][216] , \labels[4].label[207] );
tran (\labels[4][217] , \labels[4].label[208] );
tran (\labels[4][218] , \labels[4].label[209] );
tran (\labels[4][219] , \labels[4].label[210] );
tran (\labels[4][220] , \labels[4].label[211] );
tran (\labels[4][221] , \labels[4].label[212] );
tran (\labels[4][222] , \labels[4].label[213] );
tran (\labels[4][223] , \labels[4].label[214] );
tran (\labels[4][224] , \labels[4].label[215] );
tran (\labels[4][225] , \labels[4].label[216] );
tran (\labels[4][226] , \labels[4].label[217] );
tran (\labels[4][227] , \labels[4].label[218] );
tran (\labels[4][228] , \labels[4].label[219] );
tran (\labels[4][229] , \labels[4].label[220] );
tran (\labels[4][230] , \labels[4].label[221] );
tran (\labels[4][231] , \labels[4].label[222] );
tran (\labels[4][232] , \labels[4].label[223] );
tran (\labels[4][233] , \labels[4].label[224] );
tran (\labels[4][234] , \labels[4].label[225] );
tran (\labels[4][235] , \labels[4].label[226] );
tran (\labels[4][236] , \labels[4].label[227] );
tran (\labels[4][237] , \labels[4].label[228] );
tran (\labels[4][238] , \labels[4].label[229] );
tran (\labels[4][239] , \labels[4].label[230] );
tran (\labels[4][240] , \labels[4].label[231] );
tran (\labels[4][241] , \labels[4].label[232] );
tran (\labels[4][242] , \labels[4].label[233] );
tran (\labels[4][243] , \labels[4].label[234] );
tran (\labels[4][244] , \labels[4].label[235] );
tran (\labels[4][245] , \labels[4].label[236] );
tran (\labels[4][246] , \labels[4].label[237] );
tran (\labels[4][247] , \labels[4].label[238] );
tran (\labels[4][248] , \labels[4].label[239] );
tran (\labels[4][249] , \labels[4].label[240] );
tran (\labels[4][250] , \labels[4].label[241] );
tran (\labels[4][251] , \labels[4].label[242] );
tran (\labels[4][252] , \labels[4].label[243] );
tran (\labels[4][253] , \labels[4].label[244] );
tran (\labels[4][254] , \labels[4].label[245] );
tran (\labels[4][255] , \labels[4].label[246] );
tran (\labels[4][256] , \labels[4].label[247] );
tran (\labels[4][257] , \labels[4].label[248] );
tran (\labels[4][258] , \labels[4].label[249] );
tran (\labels[4][259] , \labels[4].label[250] );
tran (\labels[4][260] , \labels[4].label[251] );
tran (\labels[4][261] , \labels[4].label[252] );
tran (\labels[4][262] , \labels[4].label[253] );
tran (\labels[4][263] , \labels[4].label[254] );
tran (\labels[4][264] , \labels[4].label[255] );
tran (\labels[4][265] , \labels[4].label_size[0] );
tran (\labels[4][266] , \labels[4].label_size[1] );
tran (\labels[4][267] , \labels[4].label_size[2] );
tran (\labels[4][268] , \labels[4].label_size[3] );
tran (\labels[4][269] , \labels[4].label_size[4] );
tran (\labels[4][270] , \labels[4].label_size[5] );
tran (\labels[4][271] , \labels[4].guid_size[0] );
tran (\labels[5][0] , \labels[5].delimiter[0] );
tran (\labels[5][1] , \labels[5].delimiter[1] );
tran (\labels[5][2] , \labels[5].delimiter[2] );
tran (\labels[5][3] , \labels[5].delimiter[3] );
tran (\labels[5][4] , \labels[5].delimiter[4] );
tran (\labels[5][5] , \labels[5].delimiter[5] );
tran (\labels[5][6] , \labels[5].delimiter[6] );
tran (\labels[5][7] , \labels[5].delimiter[7] );
tran (\labels[5][8] , \labels[5].delimiter_valid[0] );
tran (\labels[5][9] , \labels[5].label[0] );
tran (\labels[5][10] , \labels[5].label[1] );
tran (\labels[5][11] , \labels[5].label[2] );
tran (\labels[5][12] , \labels[5].label[3] );
tran (\labels[5][13] , \labels[5].label[4] );
tran (\labels[5][14] , \labels[5].label[5] );
tran (\labels[5][15] , \labels[5].label[6] );
tran (\labels[5][16] , \labels[5].label[7] );
tran (\labels[5][17] , \labels[5].label[8] );
tran (\labels[5][18] , \labels[5].label[9] );
tran (\labels[5][19] , \labels[5].label[10] );
tran (\labels[5][20] , \labels[5].label[11] );
tran (\labels[5][21] , \labels[5].label[12] );
tran (\labels[5][22] , \labels[5].label[13] );
tran (\labels[5][23] , \labels[5].label[14] );
tran (\labels[5][24] , \labels[5].label[15] );
tran (\labels[5][25] , \labels[5].label[16] );
tran (\labels[5][26] , \labels[5].label[17] );
tran (\labels[5][27] , \labels[5].label[18] );
tran (\labels[5][28] , \labels[5].label[19] );
tran (\labels[5][29] , \labels[5].label[20] );
tran (\labels[5][30] , \labels[5].label[21] );
tran (\labels[5][31] , \labels[5].label[22] );
tran (\labels[5][32] , \labels[5].label[23] );
tran (\labels[5][33] , \labels[5].label[24] );
tran (\labels[5][34] , \labels[5].label[25] );
tran (\labels[5][35] , \labels[5].label[26] );
tran (\labels[5][36] , \labels[5].label[27] );
tran (\labels[5][37] , \labels[5].label[28] );
tran (\labels[5][38] , \labels[5].label[29] );
tran (\labels[5][39] , \labels[5].label[30] );
tran (\labels[5][40] , \labels[5].label[31] );
tran (\labels[5][41] , \labels[5].label[32] );
tran (\labels[5][42] , \labels[5].label[33] );
tran (\labels[5][43] , \labels[5].label[34] );
tran (\labels[5][44] , \labels[5].label[35] );
tran (\labels[5][45] , \labels[5].label[36] );
tran (\labels[5][46] , \labels[5].label[37] );
tran (\labels[5][47] , \labels[5].label[38] );
tran (\labels[5][48] , \labels[5].label[39] );
tran (\labels[5][49] , \labels[5].label[40] );
tran (\labels[5][50] , \labels[5].label[41] );
tran (\labels[5][51] , \labels[5].label[42] );
tran (\labels[5][52] , \labels[5].label[43] );
tran (\labels[5][53] , \labels[5].label[44] );
tran (\labels[5][54] , \labels[5].label[45] );
tran (\labels[5][55] , \labels[5].label[46] );
tran (\labels[5][56] , \labels[5].label[47] );
tran (\labels[5][57] , \labels[5].label[48] );
tran (\labels[5][58] , \labels[5].label[49] );
tran (\labels[5][59] , \labels[5].label[50] );
tran (\labels[5][60] , \labels[5].label[51] );
tran (\labels[5][61] , \labels[5].label[52] );
tran (\labels[5][62] , \labels[5].label[53] );
tran (\labels[5][63] , \labels[5].label[54] );
tran (\labels[5][64] , \labels[5].label[55] );
tran (\labels[5][65] , \labels[5].label[56] );
tran (\labels[5][66] , \labels[5].label[57] );
tran (\labels[5][67] , \labels[5].label[58] );
tran (\labels[5][68] , \labels[5].label[59] );
tran (\labels[5][69] , \labels[5].label[60] );
tran (\labels[5][70] , \labels[5].label[61] );
tran (\labels[5][71] , \labels[5].label[62] );
tran (\labels[5][72] , \labels[5].label[63] );
tran (\labels[5][73] , \labels[5].label[64] );
tran (\labels[5][74] , \labels[5].label[65] );
tran (\labels[5][75] , \labels[5].label[66] );
tran (\labels[5][76] , \labels[5].label[67] );
tran (\labels[5][77] , \labels[5].label[68] );
tran (\labels[5][78] , \labels[5].label[69] );
tran (\labels[5][79] , \labels[5].label[70] );
tran (\labels[5][80] , \labels[5].label[71] );
tran (\labels[5][81] , \labels[5].label[72] );
tran (\labels[5][82] , \labels[5].label[73] );
tran (\labels[5][83] , \labels[5].label[74] );
tran (\labels[5][84] , \labels[5].label[75] );
tran (\labels[5][85] , \labels[5].label[76] );
tran (\labels[5][86] , \labels[5].label[77] );
tran (\labels[5][87] , \labels[5].label[78] );
tran (\labels[5][88] , \labels[5].label[79] );
tran (\labels[5][89] , \labels[5].label[80] );
tran (\labels[5][90] , \labels[5].label[81] );
tran (\labels[5][91] , \labels[5].label[82] );
tran (\labels[5][92] , \labels[5].label[83] );
tran (\labels[5][93] , \labels[5].label[84] );
tran (\labels[5][94] , \labels[5].label[85] );
tran (\labels[5][95] , \labels[5].label[86] );
tran (\labels[5][96] , \labels[5].label[87] );
tran (\labels[5][97] , \labels[5].label[88] );
tran (\labels[5][98] , \labels[5].label[89] );
tran (\labels[5][99] , \labels[5].label[90] );
tran (\labels[5][100] , \labels[5].label[91] );
tran (\labels[5][101] , \labels[5].label[92] );
tran (\labels[5][102] , \labels[5].label[93] );
tran (\labels[5][103] , \labels[5].label[94] );
tran (\labels[5][104] , \labels[5].label[95] );
tran (\labels[5][105] , \labels[5].label[96] );
tran (\labels[5][106] , \labels[5].label[97] );
tran (\labels[5][107] , \labels[5].label[98] );
tran (\labels[5][108] , \labels[5].label[99] );
tran (\labels[5][109] , \labels[5].label[100] );
tran (\labels[5][110] , \labels[5].label[101] );
tran (\labels[5][111] , \labels[5].label[102] );
tran (\labels[5][112] , \labels[5].label[103] );
tran (\labels[5][113] , \labels[5].label[104] );
tran (\labels[5][114] , \labels[5].label[105] );
tran (\labels[5][115] , \labels[5].label[106] );
tran (\labels[5][116] , \labels[5].label[107] );
tran (\labels[5][117] , \labels[5].label[108] );
tran (\labels[5][118] , \labels[5].label[109] );
tran (\labels[5][119] , \labels[5].label[110] );
tran (\labels[5][120] , \labels[5].label[111] );
tran (\labels[5][121] , \labels[5].label[112] );
tran (\labels[5][122] , \labels[5].label[113] );
tran (\labels[5][123] , \labels[5].label[114] );
tran (\labels[5][124] , \labels[5].label[115] );
tran (\labels[5][125] , \labels[5].label[116] );
tran (\labels[5][126] , \labels[5].label[117] );
tran (\labels[5][127] , \labels[5].label[118] );
tran (\labels[5][128] , \labels[5].label[119] );
tran (\labels[5][129] , \labels[5].label[120] );
tran (\labels[5][130] , \labels[5].label[121] );
tran (\labels[5][131] , \labels[5].label[122] );
tran (\labels[5][132] , \labels[5].label[123] );
tran (\labels[5][133] , \labels[5].label[124] );
tran (\labels[5][134] , \labels[5].label[125] );
tran (\labels[5][135] , \labels[5].label[126] );
tran (\labels[5][136] , \labels[5].label[127] );
tran (\labels[5][137] , \labels[5].label[128] );
tran (\labels[5][138] , \labels[5].label[129] );
tran (\labels[5][139] , \labels[5].label[130] );
tran (\labels[5][140] , \labels[5].label[131] );
tran (\labels[5][141] , \labels[5].label[132] );
tran (\labels[5][142] , \labels[5].label[133] );
tran (\labels[5][143] , \labels[5].label[134] );
tran (\labels[5][144] , \labels[5].label[135] );
tran (\labels[5][145] , \labels[5].label[136] );
tran (\labels[5][146] , \labels[5].label[137] );
tran (\labels[5][147] , \labels[5].label[138] );
tran (\labels[5][148] , \labels[5].label[139] );
tran (\labels[5][149] , \labels[5].label[140] );
tran (\labels[5][150] , \labels[5].label[141] );
tran (\labels[5][151] , \labels[5].label[142] );
tran (\labels[5][152] , \labels[5].label[143] );
tran (\labels[5][153] , \labels[5].label[144] );
tran (\labels[5][154] , \labels[5].label[145] );
tran (\labels[5][155] , \labels[5].label[146] );
tran (\labels[5][156] , \labels[5].label[147] );
tran (\labels[5][157] , \labels[5].label[148] );
tran (\labels[5][158] , \labels[5].label[149] );
tran (\labels[5][159] , \labels[5].label[150] );
tran (\labels[5][160] , \labels[5].label[151] );
tran (\labels[5][161] , \labels[5].label[152] );
tran (\labels[5][162] , \labels[5].label[153] );
tran (\labels[5][163] , \labels[5].label[154] );
tran (\labels[5][164] , \labels[5].label[155] );
tran (\labels[5][165] , \labels[5].label[156] );
tran (\labels[5][166] , \labels[5].label[157] );
tran (\labels[5][167] , \labels[5].label[158] );
tran (\labels[5][168] , \labels[5].label[159] );
tran (\labels[5][169] , \labels[5].label[160] );
tran (\labels[5][170] , \labels[5].label[161] );
tran (\labels[5][171] , \labels[5].label[162] );
tran (\labels[5][172] , \labels[5].label[163] );
tran (\labels[5][173] , \labels[5].label[164] );
tran (\labels[5][174] , \labels[5].label[165] );
tran (\labels[5][175] , \labels[5].label[166] );
tran (\labels[5][176] , \labels[5].label[167] );
tran (\labels[5][177] , \labels[5].label[168] );
tran (\labels[5][178] , \labels[5].label[169] );
tran (\labels[5][179] , \labels[5].label[170] );
tran (\labels[5][180] , \labels[5].label[171] );
tran (\labels[5][181] , \labels[5].label[172] );
tran (\labels[5][182] , \labels[5].label[173] );
tran (\labels[5][183] , \labels[5].label[174] );
tran (\labels[5][184] , \labels[5].label[175] );
tran (\labels[5][185] , \labels[5].label[176] );
tran (\labels[5][186] , \labels[5].label[177] );
tran (\labels[5][187] , \labels[5].label[178] );
tran (\labels[5][188] , \labels[5].label[179] );
tran (\labels[5][189] , \labels[5].label[180] );
tran (\labels[5][190] , \labels[5].label[181] );
tran (\labels[5][191] , \labels[5].label[182] );
tran (\labels[5][192] , \labels[5].label[183] );
tran (\labels[5][193] , \labels[5].label[184] );
tran (\labels[5][194] , \labels[5].label[185] );
tran (\labels[5][195] , \labels[5].label[186] );
tran (\labels[5][196] , \labels[5].label[187] );
tran (\labels[5][197] , \labels[5].label[188] );
tran (\labels[5][198] , \labels[5].label[189] );
tran (\labels[5][199] , \labels[5].label[190] );
tran (\labels[5][200] , \labels[5].label[191] );
tran (\labels[5][201] , \labels[5].label[192] );
tran (\labels[5][202] , \labels[5].label[193] );
tran (\labels[5][203] , \labels[5].label[194] );
tran (\labels[5][204] , \labels[5].label[195] );
tran (\labels[5][205] , \labels[5].label[196] );
tran (\labels[5][206] , \labels[5].label[197] );
tran (\labels[5][207] , \labels[5].label[198] );
tran (\labels[5][208] , \labels[5].label[199] );
tran (\labels[5][209] , \labels[5].label[200] );
tran (\labels[5][210] , \labels[5].label[201] );
tran (\labels[5][211] , \labels[5].label[202] );
tran (\labels[5][212] , \labels[5].label[203] );
tran (\labels[5][213] , \labels[5].label[204] );
tran (\labels[5][214] , \labels[5].label[205] );
tran (\labels[5][215] , \labels[5].label[206] );
tran (\labels[5][216] , \labels[5].label[207] );
tran (\labels[5][217] , \labels[5].label[208] );
tran (\labels[5][218] , \labels[5].label[209] );
tran (\labels[5][219] , \labels[5].label[210] );
tran (\labels[5][220] , \labels[5].label[211] );
tran (\labels[5][221] , \labels[5].label[212] );
tran (\labels[5][222] , \labels[5].label[213] );
tran (\labels[5][223] , \labels[5].label[214] );
tran (\labels[5][224] , \labels[5].label[215] );
tran (\labels[5][225] , \labels[5].label[216] );
tran (\labels[5][226] , \labels[5].label[217] );
tran (\labels[5][227] , \labels[5].label[218] );
tran (\labels[5][228] , \labels[5].label[219] );
tran (\labels[5][229] , \labels[5].label[220] );
tran (\labels[5][230] , \labels[5].label[221] );
tran (\labels[5][231] , \labels[5].label[222] );
tran (\labels[5][232] , \labels[5].label[223] );
tran (\labels[5][233] , \labels[5].label[224] );
tran (\labels[5][234] , \labels[5].label[225] );
tran (\labels[5][235] , \labels[5].label[226] );
tran (\labels[5][236] , \labels[5].label[227] );
tran (\labels[5][237] , \labels[5].label[228] );
tran (\labels[5][238] , \labels[5].label[229] );
tran (\labels[5][239] , \labels[5].label[230] );
tran (\labels[5][240] , \labels[5].label[231] );
tran (\labels[5][241] , \labels[5].label[232] );
tran (\labels[5][242] , \labels[5].label[233] );
tran (\labels[5][243] , \labels[5].label[234] );
tran (\labels[5][244] , \labels[5].label[235] );
tran (\labels[5][245] , \labels[5].label[236] );
tran (\labels[5][246] , \labels[5].label[237] );
tran (\labels[5][247] , \labels[5].label[238] );
tran (\labels[5][248] , \labels[5].label[239] );
tran (\labels[5][249] , \labels[5].label[240] );
tran (\labels[5][250] , \labels[5].label[241] );
tran (\labels[5][251] , \labels[5].label[242] );
tran (\labels[5][252] , \labels[5].label[243] );
tran (\labels[5][253] , \labels[5].label[244] );
tran (\labels[5][254] , \labels[5].label[245] );
tran (\labels[5][255] , \labels[5].label[246] );
tran (\labels[5][256] , \labels[5].label[247] );
tran (\labels[5][257] , \labels[5].label[248] );
tran (\labels[5][258] , \labels[5].label[249] );
tran (\labels[5][259] , \labels[5].label[250] );
tran (\labels[5][260] , \labels[5].label[251] );
tran (\labels[5][261] , \labels[5].label[252] );
tran (\labels[5][262] , \labels[5].label[253] );
tran (\labels[5][263] , \labels[5].label[254] );
tran (\labels[5][264] , \labels[5].label[255] );
tran (\labels[5][265] , \labels[5].label_size[0] );
tran (\labels[5][266] , \labels[5].label_size[1] );
tran (\labels[5][267] , \labels[5].label_size[2] );
tran (\labels[5][268] , \labels[5].label_size[3] );
tran (\labels[5][269] , \labels[5].label_size[4] );
tran (\labels[5][270] , \labels[5].label_size[5] );
tran (\labels[5][271] , \labels[5].guid_size[0] );
tran (\labels[6][0] , \labels[6].delimiter[0] );
tran (\labels[6][1] , \labels[6].delimiter[1] );
tran (\labels[6][2] , \labels[6].delimiter[2] );
tran (\labels[6][3] , \labels[6].delimiter[3] );
tran (\labels[6][4] , \labels[6].delimiter[4] );
tran (\labels[6][5] , \labels[6].delimiter[5] );
tran (\labels[6][6] , \labels[6].delimiter[6] );
tran (\labels[6][7] , \labels[6].delimiter[7] );
tran (\labels[6][8] , \labels[6].delimiter_valid[0] );
tran (\labels[6][9] , \labels[6].label[0] );
tran (\labels[6][10] , \labels[6].label[1] );
tran (\labels[6][11] , \labels[6].label[2] );
tran (\labels[6][12] , \labels[6].label[3] );
tran (\labels[6][13] , \labels[6].label[4] );
tran (\labels[6][14] , \labels[6].label[5] );
tran (\labels[6][15] , \labels[6].label[6] );
tran (\labels[6][16] , \labels[6].label[7] );
tran (\labels[6][17] , \labels[6].label[8] );
tran (\labels[6][18] , \labels[6].label[9] );
tran (\labels[6][19] , \labels[6].label[10] );
tran (\labels[6][20] , \labels[6].label[11] );
tran (\labels[6][21] , \labels[6].label[12] );
tran (\labels[6][22] , \labels[6].label[13] );
tran (\labels[6][23] , \labels[6].label[14] );
tran (\labels[6][24] , \labels[6].label[15] );
tran (\labels[6][25] , \labels[6].label[16] );
tran (\labels[6][26] , \labels[6].label[17] );
tran (\labels[6][27] , \labels[6].label[18] );
tran (\labels[6][28] , \labels[6].label[19] );
tran (\labels[6][29] , \labels[6].label[20] );
tran (\labels[6][30] , \labels[6].label[21] );
tran (\labels[6][31] , \labels[6].label[22] );
tran (\labels[6][32] , \labels[6].label[23] );
tran (\labels[6][33] , \labels[6].label[24] );
tran (\labels[6][34] , \labels[6].label[25] );
tran (\labels[6][35] , \labels[6].label[26] );
tran (\labels[6][36] , \labels[6].label[27] );
tran (\labels[6][37] , \labels[6].label[28] );
tran (\labels[6][38] , \labels[6].label[29] );
tran (\labels[6][39] , \labels[6].label[30] );
tran (\labels[6][40] , \labels[6].label[31] );
tran (\labels[6][41] , \labels[6].label[32] );
tran (\labels[6][42] , \labels[6].label[33] );
tran (\labels[6][43] , \labels[6].label[34] );
tran (\labels[6][44] , \labels[6].label[35] );
tran (\labels[6][45] , \labels[6].label[36] );
tran (\labels[6][46] , \labels[6].label[37] );
tran (\labels[6][47] , \labels[6].label[38] );
tran (\labels[6][48] , \labels[6].label[39] );
tran (\labels[6][49] , \labels[6].label[40] );
tran (\labels[6][50] , \labels[6].label[41] );
tran (\labels[6][51] , \labels[6].label[42] );
tran (\labels[6][52] , \labels[6].label[43] );
tran (\labels[6][53] , \labels[6].label[44] );
tran (\labels[6][54] , \labels[6].label[45] );
tran (\labels[6][55] , \labels[6].label[46] );
tran (\labels[6][56] , \labels[6].label[47] );
tran (\labels[6][57] , \labels[6].label[48] );
tran (\labels[6][58] , \labels[6].label[49] );
tran (\labels[6][59] , \labels[6].label[50] );
tran (\labels[6][60] , \labels[6].label[51] );
tran (\labels[6][61] , \labels[6].label[52] );
tran (\labels[6][62] , \labels[6].label[53] );
tran (\labels[6][63] , \labels[6].label[54] );
tran (\labels[6][64] , \labels[6].label[55] );
tran (\labels[6][65] , \labels[6].label[56] );
tran (\labels[6][66] , \labels[6].label[57] );
tran (\labels[6][67] , \labels[6].label[58] );
tran (\labels[6][68] , \labels[6].label[59] );
tran (\labels[6][69] , \labels[6].label[60] );
tran (\labels[6][70] , \labels[6].label[61] );
tran (\labels[6][71] , \labels[6].label[62] );
tran (\labels[6][72] , \labels[6].label[63] );
tran (\labels[6][73] , \labels[6].label[64] );
tran (\labels[6][74] , \labels[6].label[65] );
tran (\labels[6][75] , \labels[6].label[66] );
tran (\labels[6][76] , \labels[6].label[67] );
tran (\labels[6][77] , \labels[6].label[68] );
tran (\labels[6][78] , \labels[6].label[69] );
tran (\labels[6][79] , \labels[6].label[70] );
tran (\labels[6][80] , \labels[6].label[71] );
tran (\labels[6][81] , \labels[6].label[72] );
tran (\labels[6][82] , \labels[6].label[73] );
tran (\labels[6][83] , \labels[6].label[74] );
tran (\labels[6][84] , \labels[6].label[75] );
tran (\labels[6][85] , \labels[6].label[76] );
tran (\labels[6][86] , \labels[6].label[77] );
tran (\labels[6][87] , \labels[6].label[78] );
tran (\labels[6][88] , \labels[6].label[79] );
tran (\labels[6][89] , \labels[6].label[80] );
tran (\labels[6][90] , \labels[6].label[81] );
tran (\labels[6][91] , \labels[6].label[82] );
tran (\labels[6][92] , \labels[6].label[83] );
tran (\labels[6][93] , \labels[6].label[84] );
tran (\labels[6][94] , \labels[6].label[85] );
tran (\labels[6][95] , \labels[6].label[86] );
tran (\labels[6][96] , \labels[6].label[87] );
tran (\labels[6][97] , \labels[6].label[88] );
tran (\labels[6][98] , \labels[6].label[89] );
tran (\labels[6][99] , \labels[6].label[90] );
tran (\labels[6][100] , \labels[6].label[91] );
tran (\labels[6][101] , \labels[6].label[92] );
tran (\labels[6][102] , \labels[6].label[93] );
tran (\labels[6][103] , \labels[6].label[94] );
tran (\labels[6][104] , \labels[6].label[95] );
tran (\labels[6][105] , \labels[6].label[96] );
tran (\labels[6][106] , \labels[6].label[97] );
tran (\labels[6][107] , \labels[6].label[98] );
tran (\labels[6][108] , \labels[6].label[99] );
tran (\labels[6][109] , \labels[6].label[100] );
tran (\labels[6][110] , \labels[6].label[101] );
tran (\labels[6][111] , \labels[6].label[102] );
tran (\labels[6][112] , \labels[6].label[103] );
tran (\labels[6][113] , \labels[6].label[104] );
tran (\labels[6][114] , \labels[6].label[105] );
tran (\labels[6][115] , \labels[6].label[106] );
tran (\labels[6][116] , \labels[6].label[107] );
tran (\labels[6][117] , \labels[6].label[108] );
tran (\labels[6][118] , \labels[6].label[109] );
tran (\labels[6][119] , \labels[6].label[110] );
tran (\labels[6][120] , \labels[6].label[111] );
tran (\labels[6][121] , \labels[6].label[112] );
tran (\labels[6][122] , \labels[6].label[113] );
tran (\labels[6][123] , \labels[6].label[114] );
tran (\labels[6][124] , \labels[6].label[115] );
tran (\labels[6][125] , \labels[6].label[116] );
tran (\labels[6][126] , \labels[6].label[117] );
tran (\labels[6][127] , \labels[6].label[118] );
tran (\labels[6][128] , \labels[6].label[119] );
tran (\labels[6][129] , \labels[6].label[120] );
tran (\labels[6][130] , \labels[6].label[121] );
tran (\labels[6][131] , \labels[6].label[122] );
tran (\labels[6][132] , \labels[6].label[123] );
tran (\labels[6][133] , \labels[6].label[124] );
tran (\labels[6][134] , \labels[6].label[125] );
tran (\labels[6][135] , \labels[6].label[126] );
tran (\labels[6][136] , \labels[6].label[127] );
tran (\labels[6][137] , \labels[6].label[128] );
tran (\labels[6][138] , \labels[6].label[129] );
tran (\labels[6][139] , \labels[6].label[130] );
tran (\labels[6][140] , \labels[6].label[131] );
tran (\labels[6][141] , \labels[6].label[132] );
tran (\labels[6][142] , \labels[6].label[133] );
tran (\labels[6][143] , \labels[6].label[134] );
tran (\labels[6][144] , \labels[6].label[135] );
tran (\labels[6][145] , \labels[6].label[136] );
tran (\labels[6][146] , \labels[6].label[137] );
tran (\labels[6][147] , \labels[6].label[138] );
tran (\labels[6][148] , \labels[6].label[139] );
tran (\labels[6][149] , \labels[6].label[140] );
tran (\labels[6][150] , \labels[6].label[141] );
tran (\labels[6][151] , \labels[6].label[142] );
tran (\labels[6][152] , \labels[6].label[143] );
tran (\labels[6][153] , \labels[6].label[144] );
tran (\labels[6][154] , \labels[6].label[145] );
tran (\labels[6][155] , \labels[6].label[146] );
tran (\labels[6][156] , \labels[6].label[147] );
tran (\labels[6][157] , \labels[6].label[148] );
tran (\labels[6][158] , \labels[6].label[149] );
tran (\labels[6][159] , \labels[6].label[150] );
tran (\labels[6][160] , \labels[6].label[151] );
tran (\labels[6][161] , \labels[6].label[152] );
tran (\labels[6][162] , \labels[6].label[153] );
tran (\labels[6][163] , \labels[6].label[154] );
tran (\labels[6][164] , \labels[6].label[155] );
tran (\labels[6][165] , \labels[6].label[156] );
tran (\labels[6][166] , \labels[6].label[157] );
tran (\labels[6][167] , \labels[6].label[158] );
tran (\labels[6][168] , \labels[6].label[159] );
tran (\labels[6][169] , \labels[6].label[160] );
tran (\labels[6][170] , \labels[6].label[161] );
tran (\labels[6][171] , \labels[6].label[162] );
tran (\labels[6][172] , \labels[6].label[163] );
tran (\labels[6][173] , \labels[6].label[164] );
tran (\labels[6][174] , \labels[6].label[165] );
tran (\labels[6][175] , \labels[6].label[166] );
tran (\labels[6][176] , \labels[6].label[167] );
tran (\labels[6][177] , \labels[6].label[168] );
tran (\labels[6][178] , \labels[6].label[169] );
tran (\labels[6][179] , \labels[6].label[170] );
tran (\labels[6][180] , \labels[6].label[171] );
tran (\labels[6][181] , \labels[6].label[172] );
tran (\labels[6][182] , \labels[6].label[173] );
tran (\labels[6][183] , \labels[6].label[174] );
tran (\labels[6][184] , \labels[6].label[175] );
tran (\labels[6][185] , \labels[6].label[176] );
tran (\labels[6][186] , \labels[6].label[177] );
tran (\labels[6][187] , \labels[6].label[178] );
tran (\labels[6][188] , \labels[6].label[179] );
tran (\labels[6][189] , \labels[6].label[180] );
tran (\labels[6][190] , \labels[6].label[181] );
tran (\labels[6][191] , \labels[6].label[182] );
tran (\labels[6][192] , \labels[6].label[183] );
tran (\labels[6][193] , \labels[6].label[184] );
tran (\labels[6][194] , \labels[6].label[185] );
tran (\labels[6][195] , \labels[6].label[186] );
tran (\labels[6][196] , \labels[6].label[187] );
tran (\labels[6][197] , \labels[6].label[188] );
tran (\labels[6][198] , \labels[6].label[189] );
tran (\labels[6][199] , \labels[6].label[190] );
tran (\labels[6][200] , \labels[6].label[191] );
tran (\labels[6][201] , \labels[6].label[192] );
tran (\labels[6][202] , \labels[6].label[193] );
tran (\labels[6][203] , \labels[6].label[194] );
tran (\labels[6][204] , \labels[6].label[195] );
tran (\labels[6][205] , \labels[6].label[196] );
tran (\labels[6][206] , \labels[6].label[197] );
tran (\labels[6][207] , \labels[6].label[198] );
tran (\labels[6][208] , \labels[6].label[199] );
tran (\labels[6][209] , \labels[6].label[200] );
tran (\labels[6][210] , \labels[6].label[201] );
tran (\labels[6][211] , \labels[6].label[202] );
tran (\labels[6][212] , \labels[6].label[203] );
tran (\labels[6][213] , \labels[6].label[204] );
tran (\labels[6][214] , \labels[6].label[205] );
tran (\labels[6][215] , \labels[6].label[206] );
tran (\labels[6][216] , \labels[6].label[207] );
tran (\labels[6][217] , \labels[6].label[208] );
tran (\labels[6][218] , \labels[6].label[209] );
tran (\labels[6][219] , \labels[6].label[210] );
tran (\labels[6][220] , \labels[6].label[211] );
tran (\labels[6][221] , \labels[6].label[212] );
tran (\labels[6][222] , \labels[6].label[213] );
tran (\labels[6][223] , \labels[6].label[214] );
tran (\labels[6][224] , \labels[6].label[215] );
tran (\labels[6][225] , \labels[6].label[216] );
tran (\labels[6][226] , \labels[6].label[217] );
tran (\labels[6][227] , \labels[6].label[218] );
tran (\labels[6][228] , \labels[6].label[219] );
tran (\labels[6][229] , \labels[6].label[220] );
tran (\labels[6][230] , \labels[6].label[221] );
tran (\labels[6][231] , \labels[6].label[222] );
tran (\labels[6][232] , \labels[6].label[223] );
tran (\labels[6][233] , \labels[6].label[224] );
tran (\labels[6][234] , \labels[6].label[225] );
tran (\labels[6][235] , \labels[6].label[226] );
tran (\labels[6][236] , \labels[6].label[227] );
tran (\labels[6][237] , \labels[6].label[228] );
tran (\labels[6][238] , \labels[6].label[229] );
tran (\labels[6][239] , \labels[6].label[230] );
tran (\labels[6][240] , \labels[6].label[231] );
tran (\labels[6][241] , \labels[6].label[232] );
tran (\labels[6][242] , \labels[6].label[233] );
tran (\labels[6][243] , \labels[6].label[234] );
tran (\labels[6][244] , \labels[6].label[235] );
tran (\labels[6][245] , \labels[6].label[236] );
tran (\labels[6][246] , \labels[6].label[237] );
tran (\labels[6][247] , \labels[6].label[238] );
tran (\labels[6][248] , \labels[6].label[239] );
tran (\labels[6][249] , \labels[6].label[240] );
tran (\labels[6][250] , \labels[6].label[241] );
tran (\labels[6][251] , \labels[6].label[242] );
tran (\labels[6][252] , \labels[6].label[243] );
tran (\labels[6][253] , \labels[6].label[244] );
tran (\labels[6][254] , \labels[6].label[245] );
tran (\labels[6][255] , \labels[6].label[246] );
tran (\labels[6][256] , \labels[6].label[247] );
tran (\labels[6][257] , \labels[6].label[248] );
tran (\labels[6][258] , \labels[6].label[249] );
tran (\labels[6][259] , \labels[6].label[250] );
tran (\labels[6][260] , \labels[6].label[251] );
tran (\labels[6][261] , \labels[6].label[252] );
tran (\labels[6][262] , \labels[6].label[253] );
tran (\labels[6][263] , \labels[6].label[254] );
tran (\labels[6][264] , \labels[6].label[255] );
tran (\labels[6][265] , \labels[6].label_size[0] );
tran (\labels[6][266] , \labels[6].label_size[1] );
tran (\labels[6][267] , \labels[6].label_size[2] );
tran (\labels[6][268] , \labels[6].label_size[3] );
tran (\labels[6][269] , \labels[6].label_size[4] );
tran (\labels[6][270] , \labels[6].label_size[5] );
tran (\labels[6][271] , \labels[6].guid_size[0] );
tran (\labels[7][0] , \labels[7].delimiter[0] );
tran (\labels[7][1] , \labels[7].delimiter[1] );
tran (\labels[7][2] , \labels[7].delimiter[2] );
tran (\labels[7][3] , \labels[7].delimiter[3] );
tran (\labels[7][4] , \labels[7].delimiter[4] );
tran (\labels[7][5] , \labels[7].delimiter[5] );
tran (\labels[7][6] , \labels[7].delimiter[6] );
tran (\labels[7][7] , \labels[7].delimiter[7] );
tran (\labels[7][8] , \labels[7].delimiter_valid[0] );
tran (\labels[7][9] , \labels[7].label[0] );
tran (\labels[7][10] , \labels[7].label[1] );
tran (\labels[7][11] , \labels[7].label[2] );
tran (\labels[7][12] , \labels[7].label[3] );
tran (\labels[7][13] , \labels[7].label[4] );
tran (\labels[7][14] , \labels[7].label[5] );
tran (\labels[7][15] , \labels[7].label[6] );
tran (\labels[7][16] , \labels[7].label[7] );
tran (\labels[7][17] , \labels[7].label[8] );
tran (\labels[7][18] , \labels[7].label[9] );
tran (\labels[7][19] , \labels[7].label[10] );
tran (\labels[7][20] , \labels[7].label[11] );
tran (\labels[7][21] , \labels[7].label[12] );
tran (\labels[7][22] , \labels[7].label[13] );
tran (\labels[7][23] , \labels[7].label[14] );
tran (\labels[7][24] , \labels[7].label[15] );
tran (\labels[7][25] , \labels[7].label[16] );
tran (\labels[7][26] , \labels[7].label[17] );
tran (\labels[7][27] , \labels[7].label[18] );
tran (\labels[7][28] , \labels[7].label[19] );
tran (\labels[7][29] , \labels[7].label[20] );
tran (\labels[7][30] , \labels[7].label[21] );
tran (\labels[7][31] , \labels[7].label[22] );
tran (\labels[7][32] , \labels[7].label[23] );
tran (\labels[7][33] , \labels[7].label[24] );
tran (\labels[7][34] , \labels[7].label[25] );
tran (\labels[7][35] , \labels[7].label[26] );
tran (\labels[7][36] , \labels[7].label[27] );
tran (\labels[7][37] , \labels[7].label[28] );
tran (\labels[7][38] , \labels[7].label[29] );
tran (\labels[7][39] , \labels[7].label[30] );
tran (\labels[7][40] , \labels[7].label[31] );
tran (\labels[7][41] , \labels[7].label[32] );
tran (\labels[7][42] , \labels[7].label[33] );
tran (\labels[7][43] , \labels[7].label[34] );
tran (\labels[7][44] , \labels[7].label[35] );
tran (\labels[7][45] , \labels[7].label[36] );
tran (\labels[7][46] , \labels[7].label[37] );
tran (\labels[7][47] , \labels[7].label[38] );
tran (\labels[7][48] , \labels[7].label[39] );
tran (\labels[7][49] , \labels[7].label[40] );
tran (\labels[7][50] , \labels[7].label[41] );
tran (\labels[7][51] , \labels[7].label[42] );
tran (\labels[7][52] , \labels[7].label[43] );
tran (\labels[7][53] , \labels[7].label[44] );
tran (\labels[7][54] , \labels[7].label[45] );
tran (\labels[7][55] , \labels[7].label[46] );
tran (\labels[7][56] , \labels[7].label[47] );
tran (\labels[7][57] , \labels[7].label[48] );
tran (\labels[7][58] , \labels[7].label[49] );
tran (\labels[7][59] , \labels[7].label[50] );
tran (\labels[7][60] , \labels[7].label[51] );
tran (\labels[7][61] , \labels[7].label[52] );
tran (\labels[7][62] , \labels[7].label[53] );
tran (\labels[7][63] , \labels[7].label[54] );
tran (\labels[7][64] , \labels[7].label[55] );
tran (\labels[7][65] , \labels[7].label[56] );
tran (\labels[7][66] , \labels[7].label[57] );
tran (\labels[7][67] , \labels[7].label[58] );
tran (\labels[7][68] , \labels[7].label[59] );
tran (\labels[7][69] , \labels[7].label[60] );
tran (\labels[7][70] , \labels[7].label[61] );
tran (\labels[7][71] , \labels[7].label[62] );
tran (\labels[7][72] , \labels[7].label[63] );
tran (\labels[7][73] , \labels[7].label[64] );
tran (\labels[7][74] , \labels[7].label[65] );
tran (\labels[7][75] , \labels[7].label[66] );
tran (\labels[7][76] , \labels[7].label[67] );
tran (\labels[7][77] , \labels[7].label[68] );
tran (\labels[7][78] , \labels[7].label[69] );
tran (\labels[7][79] , \labels[7].label[70] );
tran (\labels[7][80] , \labels[7].label[71] );
tran (\labels[7][81] , \labels[7].label[72] );
tran (\labels[7][82] , \labels[7].label[73] );
tran (\labels[7][83] , \labels[7].label[74] );
tran (\labels[7][84] , \labels[7].label[75] );
tran (\labels[7][85] , \labels[7].label[76] );
tran (\labels[7][86] , \labels[7].label[77] );
tran (\labels[7][87] , \labels[7].label[78] );
tran (\labels[7][88] , \labels[7].label[79] );
tran (\labels[7][89] , \labels[7].label[80] );
tran (\labels[7][90] , \labels[7].label[81] );
tran (\labels[7][91] , \labels[7].label[82] );
tran (\labels[7][92] , \labels[7].label[83] );
tran (\labels[7][93] , \labels[7].label[84] );
tran (\labels[7][94] , \labels[7].label[85] );
tran (\labels[7][95] , \labels[7].label[86] );
tran (\labels[7][96] , \labels[7].label[87] );
tran (\labels[7][97] , \labels[7].label[88] );
tran (\labels[7][98] , \labels[7].label[89] );
tran (\labels[7][99] , \labels[7].label[90] );
tran (\labels[7][100] , \labels[7].label[91] );
tran (\labels[7][101] , \labels[7].label[92] );
tran (\labels[7][102] , \labels[7].label[93] );
tran (\labels[7][103] , \labels[7].label[94] );
tran (\labels[7][104] , \labels[7].label[95] );
tran (\labels[7][105] , \labels[7].label[96] );
tran (\labels[7][106] , \labels[7].label[97] );
tran (\labels[7][107] , \labels[7].label[98] );
tran (\labels[7][108] , \labels[7].label[99] );
tran (\labels[7][109] , \labels[7].label[100] );
tran (\labels[7][110] , \labels[7].label[101] );
tran (\labels[7][111] , \labels[7].label[102] );
tran (\labels[7][112] , \labels[7].label[103] );
tran (\labels[7][113] , \labels[7].label[104] );
tran (\labels[7][114] , \labels[7].label[105] );
tran (\labels[7][115] , \labels[7].label[106] );
tran (\labels[7][116] , \labels[7].label[107] );
tran (\labels[7][117] , \labels[7].label[108] );
tran (\labels[7][118] , \labels[7].label[109] );
tran (\labels[7][119] , \labels[7].label[110] );
tran (\labels[7][120] , \labels[7].label[111] );
tran (\labels[7][121] , \labels[7].label[112] );
tran (\labels[7][122] , \labels[7].label[113] );
tran (\labels[7][123] , \labels[7].label[114] );
tran (\labels[7][124] , \labels[7].label[115] );
tran (\labels[7][125] , \labels[7].label[116] );
tran (\labels[7][126] , \labels[7].label[117] );
tran (\labels[7][127] , \labels[7].label[118] );
tran (\labels[7][128] , \labels[7].label[119] );
tran (\labels[7][129] , \labels[7].label[120] );
tran (\labels[7][130] , \labels[7].label[121] );
tran (\labels[7][131] , \labels[7].label[122] );
tran (\labels[7][132] , \labels[7].label[123] );
tran (\labels[7][133] , \labels[7].label[124] );
tran (\labels[7][134] , \labels[7].label[125] );
tran (\labels[7][135] , \labels[7].label[126] );
tran (\labels[7][136] , \labels[7].label[127] );
tran (\labels[7][137] , \labels[7].label[128] );
tran (\labels[7][138] , \labels[7].label[129] );
tran (\labels[7][139] , \labels[7].label[130] );
tran (\labels[7][140] , \labels[7].label[131] );
tran (\labels[7][141] , \labels[7].label[132] );
tran (\labels[7][142] , \labels[7].label[133] );
tran (\labels[7][143] , \labels[7].label[134] );
tran (\labels[7][144] , \labels[7].label[135] );
tran (\labels[7][145] , \labels[7].label[136] );
tran (\labels[7][146] , \labels[7].label[137] );
tran (\labels[7][147] , \labels[7].label[138] );
tran (\labels[7][148] , \labels[7].label[139] );
tran (\labels[7][149] , \labels[7].label[140] );
tran (\labels[7][150] , \labels[7].label[141] );
tran (\labels[7][151] , \labels[7].label[142] );
tran (\labels[7][152] , \labels[7].label[143] );
tran (\labels[7][153] , \labels[7].label[144] );
tran (\labels[7][154] , \labels[7].label[145] );
tran (\labels[7][155] , \labels[7].label[146] );
tran (\labels[7][156] , \labels[7].label[147] );
tran (\labels[7][157] , \labels[7].label[148] );
tran (\labels[7][158] , \labels[7].label[149] );
tran (\labels[7][159] , \labels[7].label[150] );
tran (\labels[7][160] , \labels[7].label[151] );
tran (\labels[7][161] , \labels[7].label[152] );
tran (\labels[7][162] , \labels[7].label[153] );
tran (\labels[7][163] , \labels[7].label[154] );
tran (\labels[7][164] , \labels[7].label[155] );
tran (\labels[7][165] , \labels[7].label[156] );
tran (\labels[7][166] , \labels[7].label[157] );
tran (\labels[7][167] , \labels[7].label[158] );
tran (\labels[7][168] , \labels[7].label[159] );
tran (\labels[7][169] , \labels[7].label[160] );
tran (\labels[7][170] , \labels[7].label[161] );
tran (\labels[7][171] , \labels[7].label[162] );
tran (\labels[7][172] , \labels[7].label[163] );
tran (\labels[7][173] , \labels[7].label[164] );
tran (\labels[7][174] , \labels[7].label[165] );
tran (\labels[7][175] , \labels[7].label[166] );
tran (\labels[7][176] , \labels[7].label[167] );
tran (\labels[7][177] , \labels[7].label[168] );
tran (\labels[7][178] , \labels[7].label[169] );
tran (\labels[7][179] , \labels[7].label[170] );
tran (\labels[7][180] , \labels[7].label[171] );
tran (\labels[7][181] , \labels[7].label[172] );
tran (\labels[7][182] , \labels[7].label[173] );
tran (\labels[7][183] , \labels[7].label[174] );
tran (\labels[7][184] , \labels[7].label[175] );
tran (\labels[7][185] , \labels[7].label[176] );
tran (\labels[7][186] , \labels[7].label[177] );
tran (\labels[7][187] , \labels[7].label[178] );
tran (\labels[7][188] , \labels[7].label[179] );
tran (\labels[7][189] , \labels[7].label[180] );
tran (\labels[7][190] , \labels[7].label[181] );
tran (\labels[7][191] , \labels[7].label[182] );
tran (\labels[7][192] , \labels[7].label[183] );
tran (\labels[7][193] , \labels[7].label[184] );
tran (\labels[7][194] , \labels[7].label[185] );
tran (\labels[7][195] , \labels[7].label[186] );
tran (\labels[7][196] , \labels[7].label[187] );
tran (\labels[7][197] , \labels[7].label[188] );
tran (\labels[7][198] , \labels[7].label[189] );
tran (\labels[7][199] , \labels[7].label[190] );
tran (\labels[7][200] , \labels[7].label[191] );
tran (\labels[7][201] , \labels[7].label[192] );
tran (\labels[7][202] , \labels[7].label[193] );
tran (\labels[7][203] , \labels[7].label[194] );
tran (\labels[7][204] , \labels[7].label[195] );
tran (\labels[7][205] , \labels[7].label[196] );
tran (\labels[7][206] , \labels[7].label[197] );
tran (\labels[7][207] , \labels[7].label[198] );
tran (\labels[7][208] , \labels[7].label[199] );
tran (\labels[7][209] , \labels[7].label[200] );
tran (\labels[7][210] , \labels[7].label[201] );
tran (\labels[7][211] , \labels[7].label[202] );
tran (\labels[7][212] , \labels[7].label[203] );
tran (\labels[7][213] , \labels[7].label[204] );
tran (\labels[7][214] , \labels[7].label[205] );
tran (\labels[7][215] , \labels[7].label[206] );
tran (\labels[7][216] , \labels[7].label[207] );
tran (\labels[7][217] , \labels[7].label[208] );
tran (\labels[7][218] , \labels[7].label[209] );
tran (\labels[7][219] , \labels[7].label[210] );
tran (\labels[7][220] , \labels[7].label[211] );
tran (\labels[7][221] , \labels[7].label[212] );
tran (\labels[7][222] , \labels[7].label[213] );
tran (\labels[7][223] , \labels[7].label[214] );
tran (\labels[7][224] , \labels[7].label[215] );
tran (\labels[7][225] , \labels[7].label[216] );
tran (\labels[7][226] , \labels[7].label[217] );
tran (\labels[7][227] , \labels[7].label[218] );
tran (\labels[7][228] , \labels[7].label[219] );
tran (\labels[7][229] , \labels[7].label[220] );
tran (\labels[7][230] , \labels[7].label[221] );
tran (\labels[7][231] , \labels[7].label[222] );
tran (\labels[7][232] , \labels[7].label[223] );
tran (\labels[7][233] , \labels[7].label[224] );
tran (\labels[7][234] , \labels[7].label[225] );
tran (\labels[7][235] , \labels[7].label[226] );
tran (\labels[7][236] , \labels[7].label[227] );
tran (\labels[7][237] , \labels[7].label[228] );
tran (\labels[7][238] , \labels[7].label[229] );
tran (\labels[7][239] , \labels[7].label[230] );
tran (\labels[7][240] , \labels[7].label[231] );
tran (\labels[7][241] , \labels[7].label[232] );
tran (\labels[7][242] , \labels[7].label[233] );
tran (\labels[7][243] , \labels[7].label[234] );
tran (\labels[7][244] , \labels[7].label[235] );
tran (\labels[7][245] , \labels[7].label[236] );
tran (\labels[7][246] , \labels[7].label[237] );
tran (\labels[7][247] , \labels[7].label[238] );
tran (\labels[7][248] , \labels[7].label[239] );
tran (\labels[7][249] , \labels[7].label[240] );
tran (\labels[7][250] , \labels[7].label[241] );
tran (\labels[7][251] , \labels[7].label[242] );
tran (\labels[7][252] , \labels[7].label[243] );
tran (\labels[7][253] , \labels[7].label[244] );
tran (\labels[7][254] , \labels[7].label[245] );
tran (\labels[7][255] , \labels[7].label[246] );
tran (\labels[7][256] , \labels[7].label[247] );
tran (\labels[7][257] , \labels[7].label[248] );
tran (\labels[7][258] , \labels[7].label[249] );
tran (\labels[7][259] , \labels[7].label[250] );
tran (\labels[7][260] , \labels[7].label[251] );
tran (\labels[7][261] , \labels[7].label[252] );
tran (\labels[7][262] , \labels[7].label[253] );
tran (\labels[7][263] , \labels[7].label[254] );
tran (\labels[7][264] , \labels[7].label[255] );
tran (\labels[7][265] , \labels[7].label_size[0] );
tran (\labels[7][266] , \labels[7].label_size[1] );
tran (\labels[7][267] , \labels[7].label_size[2] );
tran (\labels[7][268] , \labels[7].label_size[3] );
tran (\labels[7][269] , \labels[7].label_size[4] );
tran (\labels[7][270] , \labels[7].label_size[5] );
tran (\labels[7][271] , \labels[7].guid_size[0] );
tran (kme_internal_out[70], \kme_internal_out.sot [0]);
tran (kme_internal_out[69], \kme_internal_out.eoi [0]);
tran (kme_internal_out[68], \kme_internal_out.eot [0]);
tran (kme_internal_out[67], \kme_internal_out.id [3]);
tran (kme_internal_out[66], \kme_internal_out.id [2]);
tran (kme_internal_out[65], \kme_internal_out.id [1]);
tran (kme_internal_out[64], \kme_internal_out.id [0]);
tran (kme_internal_out[63], \kme_internal_out.tdata [63]);
tran (kme_internal_out[62], \kme_internal_out.tdata [62]);
tran (kme_internal_out[61], \kme_internal_out.tdata [61]);
tran (kme_internal_out[60], \kme_internal_out.tdata [60]);
tran (kme_internal_out[59], \kme_internal_out.tdata [59]);
tran (kme_internal_out[58], \kme_internal_out.tdata [58]);
tran (kme_internal_out[57], \kme_internal_out.tdata [57]);
tran (kme_internal_out[56], \kme_internal_out.tdata [56]);
tran (kme_internal_out[55], \kme_internal_out.tdata [55]);
tran (kme_internal_out[54], \kme_internal_out.tdata [54]);
tran (kme_internal_out[53], \kme_internal_out.tdata [53]);
tran (kme_internal_out[52], \kme_internal_out.tdata [52]);
tran (kme_internal_out[51], \kme_internal_out.tdata [51]);
tran (kme_internal_out[50], \kme_internal_out.tdata [50]);
tran (kme_internal_out[49], \kme_internal_out.tdata [49]);
tran (kme_internal_out[48], \kme_internal_out.tdata [48]);
tran (kme_internal_out[47], \kme_internal_out.tdata [47]);
tran (kme_internal_out[46], \kme_internal_out.tdata [46]);
tran (kme_internal_out[45], \kme_internal_out.tdata [45]);
tran (kme_internal_out[44], \kme_internal_out.tdata [44]);
tran (kme_internal_out[43], \kme_internal_out.tdata [43]);
tran (kme_internal_out[42], \kme_internal_out.tdata [42]);
tran (kme_internal_out[41], \kme_internal_out.tdata [41]);
tran (kme_internal_out[40], \kme_internal_out.tdata [40]);
tran (kme_internal_out[39], \kme_internal_out.tdata [39]);
tran (kme_internal_out[38], \kme_internal_out.tdata [38]);
tran (kme_internal_out[37], \kme_internal_out.tdata [37]);
tran (kme_internal_out[36], \kme_internal_out.tdata [36]);
tran (kme_internal_out[35], \kme_internal_out.tdata [35]);
tran (kme_internal_out[34], \kme_internal_out.tdata [34]);
tran (kme_internal_out[33], \kme_internal_out.tdata [33]);
tran (kme_internal_out[32], \kme_internal_out.tdata [32]);
tran (kme_internal_out[31], \kme_internal_out.tdata [31]);
tran (kme_internal_out[30], \kme_internal_out.tdata [30]);
tran (kme_internal_out[29], \kme_internal_out.tdata [29]);
tran (kme_internal_out[28], \kme_internal_out.tdata [28]);
tran (kme_internal_out[27], \kme_internal_out.tdata [27]);
tran (kme_internal_out[26], \kme_internal_out.tdata [26]);
tran (kme_internal_out[25], \kme_internal_out.tdata [25]);
tran (kme_internal_out[24], \kme_internal_out.tdata [24]);
tran (kme_internal_out[23], \kme_internal_out.tdata [23]);
tran (kme_internal_out[22], \kme_internal_out.tdata [22]);
tran (kme_internal_out[21], \kme_internal_out.tdata [21]);
tran (kme_internal_out[20], \kme_internal_out.tdata [20]);
tran (kme_internal_out[19], \kme_internal_out.tdata [19]);
tran (kme_internal_out[18], \kme_internal_out.tdata [18]);
tran (kme_internal_out[17], \kme_internal_out.tdata [17]);
tran (kme_internal_out[16], \kme_internal_out.tdata [16]);
tran (kme_internal_out[15], \kme_internal_out.tdata [15]);
tran (kme_internal_out[14], \kme_internal_out.tdata [14]);
tran (kme_internal_out[13], \kme_internal_out.tdata [13]);
tran (kme_internal_out[12], \kme_internal_out.tdata [12]);
tran (kme_internal_out[11], \kme_internal_out.tdata [11]);
tran (kme_internal_out[10], \kme_internal_out.tdata [10]);
tran (kme_internal_out[9], \kme_internal_out.tdata [9]);
tran (kme_internal_out[8], \kme_internal_out.tdata [8]);
tran (kme_internal_out[7], \kme_internal_out.tdata [7]);
tran (kme_internal_out[6], \kme_internal_out.tdata [6]);
tran (kme_internal_out[5], \kme_internal_out.tdata [5]);
tran (kme_internal_out[4], \kme_internal_out.tdata [4]);
tran (kme_internal_out[3], \kme_internal_out.tdata [3]);
tran (kme_internal_out[2], \kme_internal_out.tdata [2]);
tran (kme_internal_out[1], \kme_internal_out.tdata [1]);
tran (kme_internal_out[0], \kme_internal_out.tdata [0]);
tran (debug_cmd[31], \debug_cmd.tlvp_corrupt [0]);
tran (int_tlv_word0[63], \int_tlv_word0.tlv_bip2 [1]);
tran (int_tlv_word8[63], \int_tlv_word8.dek_kim_entry.valid [0]);
tran (int_tlv_word9[63], \int_tlv_word9.dak_kim_entry.valid [0]);
tran (debug_cmd[30], \debug_cmd.cmd_mode [1]);
tran (int_tlv_word0[62], \int_tlv_word0.tlv_bip2 [0]);
tran (int_tlv_word8[62], \int_tlv_word8.dek_kim_entry.label_index [2]);
tran (int_tlv_word9[62], \int_tlv_word9.dak_kim_entry.label_index [2]);
tran (debug_cmd[29], \debug_cmd.cmd_mode [0]);
tran (int_tlv_word0[61], \int_tlv_word0.resv0 [12]);
tran (int_tlv_word8[61], \int_tlv_word8.dek_kim_entry.label_index [1]);
tran (int_tlv_word9[61], \int_tlv_word9.dak_kim_entry.label_index [1]);
tran (debug_cmd[28], \debug_cmd.module_id [4]);
tran (int_tlv_word0[60], \int_tlv_word0.resv0 [11]);
tran (int_tlv_word8[60], \int_tlv_word8.dek_kim_entry.label_index [0]);
tran (int_tlv_word9[60], \int_tlv_word9.dak_kim_entry.label_index [0]);
tran (debug_cmd[27], \debug_cmd.module_id [3]);
tran (int_tlv_word0[59], \int_tlv_word0.resv0 [10]);
tran (int_tlv_word8[59], \int_tlv_word8.dek_kim_entry.ckv_length [1]);
tran (int_tlv_word9[59], \int_tlv_word9.dak_kim_entry.ckv_length [1]);
tran (debug_cmd[26], \debug_cmd.module_id [2]);
tran (int_tlv_word0[58], \int_tlv_word0.resv0 [9]);
tran (int_tlv_word8[58], \int_tlv_word8.dek_kim_entry.ckv_length [0]);
tran (int_tlv_word9[58], \int_tlv_word9.dak_kim_entry.ckv_length [0]);
tran (debug_cmd[25], \debug_cmd.module_id [1]);
tran (int_tlv_word0[57], \int_tlv_word0.resv0 [8]);
tran (int_tlv_word8[57], \int_tlv_word8.dek_kim_entry.ckv_pointer [14]);
tran (int_tlv_word9[57], \int_tlv_word9.dak_kim_entry.ckv_pointer [14]);
tran (debug_cmd[24], \debug_cmd.module_id [0]);
tran (int_tlv_word0[56], \int_tlv_word0.resv0 [7]);
tran (int_tlv_word8[56], \int_tlv_word8.dek_kim_entry.ckv_pointer [13]);
tran (int_tlv_word9[56], \int_tlv_word9.dak_kim_entry.ckv_pointer [13]);
tran (debug_cmd[23], \debug_cmd.cmd_type [0]);
tran (int_tlv_word0[55], \int_tlv_word0.resv0 [6]);
tran (int_tlv_word8[55], \int_tlv_word8.dek_kim_entry.ckv_pointer [12]);
tran (int_tlv_word9[55], \int_tlv_word9.dak_kim_entry.ckv_pointer [12]);
tran (int_tlv_word42[55], \int_tlv_word42.corrupt_crc32 [0]);
tran (debug_cmd[22], \debug_cmd.tlv_num [4]);
tran (int_tlv_word0[54], \int_tlv_word0.resv0 [5]);
tran (int_tlv_word8[54], \int_tlv_word8.dek_kim_entry.ckv_pointer [11]);
tran (int_tlv_word9[54], \int_tlv_word9.dak_kim_entry.ckv_pointer [11]);
tran (int_tlv_word42[54], \int_tlv_word42.unused [46]);
tran (debug_cmd[21], \debug_cmd.tlv_num [3]);
tran (int_tlv_word0[53], \int_tlv_word0.resv0 [4]);
tran (int_tlv_word8[53], \int_tlv_word8.dek_kim_entry.ckv_pointer [10]);
tran (int_tlv_word9[53], \int_tlv_word9.dak_kim_entry.ckv_pointer [10]);
tran (int_tlv_word42[53], \int_tlv_word42.unused [45]);
tran (debug_cmd[20], \debug_cmd.tlv_num [2]);
tran (int_tlv_word0[52], \int_tlv_word0.resv0 [3]);
tran (int_tlv_word8[52], \int_tlv_word8.dek_kim_entry.ckv_pointer [9]);
tran (int_tlv_word9[52], \int_tlv_word9.dak_kim_entry.ckv_pointer [9]);
tran (int_tlv_word42[52], \int_tlv_word42.unused [44]);
tran (debug_cmd[19], \debug_cmd.tlv_num [1]);
tran (int_tlv_word0[51], \int_tlv_word0.resv0 [2]);
tran (int_tlv_word8[51], \int_tlv_word8.dek_kim_entry.ckv_pointer [8]);
tran (int_tlv_word9[51], \int_tlv_word9.dak_kim_entry.ckv_pointer [8]);
tran (int_tlv_word42[51], \int_tlv_word42.unused [43]);
tran (debug_cmd[18], \debug_cmd.tlv_num [0]);
tran (int_tlv_word0[50], \int_tlv_word0.resv0 [1]);
tran (int_tlv_word8[50], \int_tlv_word8.dek_kim_entry.ckv_pointer [7]);
tran (int_tlv_word9[50], \int_tlv_word9.dak_kim_entry.ckv_pointer [7]);
tran (int_tlv_word42[50], \int_tlv_word42.unused [42]);
tran (debug_cmd[17], \debug_cmd.byte_num [9]);
tran (int_tlv_word0[49], \int_tlv_word0.resv0 [0]);
tran (int_tlv_word8[49], \int_tlv_word8.dek_kim_entry.ckv_pointer [6]);
tran (int_tlv_word9[49], \int_tlv_word9.dak_kim_entry.ckv_pointer [6]);
tran (int_tlv_word42[49], \int_tlv_word42.unused [41]);
tran (debug_cmd[16], \debug_cmd.byte_num [8]);
tran (int_tlv_word0[48], \int_tlv_word0.kdf_dek_iter [0]);
tran (int_tlv_word8[48], \int_tlv_word8.dek_kim_entry.ckv_pointer [5]);
tran (int_tlv_word9[48], \int_tlv_word9.dak_kim_entry.ckv_pointer [5]);
tran (int_tlv_word42[48], \int_tlv_word42.unused [40]);
tran (debug_cmd[15], \debug_cmd.byte_num [7]);
tran (int_tlv_word0[47], \int_tlv_word0.keyless_algos [0]);
tran (int_tlv_word8[47], \int_tlv_word8.dek_kim_entry.ckv_pointer [4]);
tran (int_tlv_word9[47], \int_tlv_word9.dak_kim_entry.ckv_pointer [4]);
tran (int_tlv_word42[47], \int_tlv_word42.unused [39]);
tran (debug_cmd[14], \debug_cmd.byte_num [6]);
tran (int_tlv_word0[46], \int_tlv_word0.needs_dek [0]);
tran (int_tlv_word8[46], \int_tlv_word8.dek_kim_entry.ckv_pointer [3]);
tran (int_tlv_word9[46], \int_tlv_word9.dak_kim_entry.ckv_pointer [3]);
tran (int_tlv_word42[46], \int_tlv_word42.unused [38]);
tran (debug_cmd[13], \debug_cmd.byte_num [5]);
tran (int_tlv_word0[45], \int_tlv_word0.needs_dak [0]);
tran (int_tlv_word8[45], \int_tlv_word8.dek_kim_entry.ckv_pointer [2]);
tran (int_tlv_word9[45], \int_tlv_word9.dak_kim_entry.ckv_pointer [2]);
tran (int_tlv_word42[45], \int_tlv_word42.unused [37]);
tran (debug_cmd[12], \debug_cmd.byte_num [4]);
tran (int_tlv_word0[44], \int_tlv_word0.key_type [5]);
tran (int_tlv_word8[44], \int_tlv_word8.dek_kim_entry.ckv_pointer [1]);
tran (int_tlv_word9[44], \int_tlv_word9.dak_kim_entry.ckv_pointer [1]);
tran (int_tlv_word42[44], \int_tlv_word42.unused [36]);
tran (debug_cmd[11], \debug_cmd.byte_num [3]);
tran (int_tlv_word0[43], \int_tlv_word0.key_type [4]);
tran (int_tlv_word8[43], \int_tlv_word8.dek_kim_entry.ckv_pointer [0]);
tran (int_tlv_word9[43], \int_tlv_word9.dak_kim_entry.ckv_pointer [0]);
tran (int_tlv_word42[43], \int_tlv_word42.unused [35]);
tran (debug_cmd[10], \debug_cmd.byte_num [2]);
tran (int_tlv_word0[42], \int_tlv_word0.key_type [3]);
tran (int_tlv_word8[42], \int_tlv_word8.dek_kim_entry.pf_num [3]);
tran (int_tlv_word9[42], \int_tlv_word9.dak_kim_entry.pf_num [3]);
tran (int_tlv_word42[42], \int_tlv_word42.unused [34]);
tran (debug_cmd[9], \debug_cmd.byte_num [1]);
tran (int_tlv_word0[41], \int_tlv_word0.key_type [2]);
tran (int_tlv_word8[41], \int_tlv_word8.dek_kim_entry.pf_num [2]);
tran (int_tlv_word9[41], \int_tlv_word9.dak_kim_entry.pf_num [2]);
tran (int_tlv_word42[41], \int_tlv_word42.unused [33]);
tran (debug_cmd[8], \debug_cmd.byte_num [0]);
tran (int_tlv_word0[40], \int_tlv_word0.key_type [1]);
tran (int_tlv_word8[40], \int_tlv_word8.dek_kim_entry.pf_num [1]);
tran (int_tlv_word9[40], \int_tlv_word9.dak_kim_entry.pf_num [1]);
tran (int_tlv_word42[40], \int_tlv_word42.unused [32]);
tran (debug_cmd[7], \debug_cmd.byte_msk [7]);
tran (int_tlv_word0[39], \int_tlv_word0.key_type [0]);
tran (int_tlv_word8[39], \int_tlv_word8.dek_kim_entry.pf_num [0]);
tran (int_tlv_word9[39], \int_tlv_word9.dak_kim_entry.pf_num [0]);
tran (int_tlv_word42[39], \int_tlv_word42.unused [31]);
tran (debug_cmd[6], \debug_cmd.byte_msk [6]);
tran (int_tlv_word0[38], \int_tlv_word0.tlv_frame_num [10]);
tran (int_tlv_word8[38], \int_tlv_word8.dek_kim_entry.vf_num [11]);
tran (int_tlv_word9[38], \int_tlv_word9.dak_kim_entry.vf_num [11]);
tran (int_tlv_word42[38], \int_tlv_word42.unused [30]);
tran (debug_cmd[5], \debug_cmd.byte_msk [5]);
tran (int_tlv_word0[37], \int_tlv_word0.tlv_frame_num [9]);
tran (int_tlv_word8[37], \int_tlv_word8.dek_kim_entry.vf_num [10]);
tran (int_tlv_word9[37], \int_tlv_word9.dak_kim_entry.vf_num [10]);
tran (int_tlv_word42[37], \int_tlv_word42.unused [29]);
tran (debug_cmd[4], \debug_cmd.byte_msk [4]);
tran (int_tlv_word0[36], \int_tlv_word0.tlv_frame_num [8]);
tran (int_tlv_word8[36], \int_tlv_word8.dek_kim_entry.vf_num [9]);
tran (int_tlv_word9[36], \int_tlv_word9.dak_kim_entry.vf_num [9]);
tran (int_tlv_word42[36], \int_tlv_word42.unused [28]);
tran (debug_cmd[3], \debug_cmd.byte_msk [3]);
tran (int_tlv_word0[35], \int_tlv_word0.tlv_frame_num [7]);
tran (int_tlv_word8[35], \int_tlv_word8.dek_kim_entry.vf_num [8]);
tran (int_tlv_word9[35], \int_tlv_word9.dak_kim_entry.vf_num [8]);
tran (int_tlv_word42[35], \int_tlv_word42.unused [27]);
tran (debug_cmd[2], \debug_cmd.byte_msk [2]);
tran (int_tlv_word0[34], \int_tlv_word0.tlv_frame_num [6]);
tran (int_tlv_word8[34], \int_tlv_word8.dek_kim_entry.vf_num [7]);
tran (int_tlv_word9[34], \int_tlv_word9.dak_kim_entry.vf_num [7]);
tran (int_tlv_word42[34], \int_tlv_word42.unused [26]);
tran (debug_cmd[1], \debug_cmd.byte_msk [1]);
tran (int_tlv_word0[33], \int_tlv_word0.tlv_frame_num [5]);
tran (int_tlv_word8[33], \int_tlv_word8.dek_kim_entry.vf_num [6]);
tran (int_tlv_word9[33], \int_tlv_word9.dak_kim_entry.vf_num [6]);
tran (int_tlv_word42[33], \int_tlv_word42.unused [25]);
tran (debug_cmd[0], \debug_cmd.byte_msk [0]);
tran (int_tlv_word0[32], \int_tlv_word0.tlv_frame_num [4]);
tran (int_tlv_word8[32], \int_tlv_word8.dek_kim_entry.vf_num [5]);
tran (int_tlv_word9[32], \int_tlv_word9.dak_kim_entry.vf_num [5]);
tran (int_tlv_word42[32], \int_tlv_word42.unused [24]);
tran (int_tlv_word0[31], \int_tlv_word0.tlv_frame_num [3]);
tran (int_tlv_word8[31], \int_tlv_word8.dek_kim_entry.vf_num [4]);
tran (int_tlv_word9[31], \int_tlv_word9.dak_kim_entry.vf_num [4]);
tran (int_tlv_word42[31], \int_tlv_word42.unused [23]);
tran (key_header[31], \key_header.dak_key_op [0]);
tran (int_tlv_word0[30], \int_tlv_word0.tlv_frame_num [2]);
tran (int_tlv_word8[30], \int_tlv_word8.dek_kim_entry.vf_num [3]);
tran (int_tlv_word9[30], \int_tlv_word9.dak_kim_entry.vf_num [3]);
tran (int_tlv_word42[30], \int_tlv_word42.unused [22]);
tran (key_header[30], \key_header.dak_key_ref [13]);
tran (int_tlv_word0[29], \int_tlv_word0.tlv_frame_num [1]);
tran (int_tlv_word8[29], \int_tlv_word8.dek_kim_entry.vf_num [2]);
tran (int_tlv_word9[29], \int_tlv_word9.dak_kim_entry.vf_num [2]);
tran (int_tlv_word42[29], \int_tlv_word42.unused [21]);
tran (key_header[29], \key_header.dak_key_ref [12]);
tran (int_tlv_word0[28], \int_tlv_word0.tlv_frame_num [0]);
tran (int_tlv_word8[28], \int_tlv_word8.dek_kim_entry.vf_num [1]);
tran (int_tlv_word9[28], \int_tlv_word9.dak_kim_entry.vf_num [1]);
tran (int_tlv_word42[28], \int_tlv_word42.unused [20]);
tran (key_header[28], \key_header.dak_key_ref [11]);
tran (int_tlv_word0[27], \int_tlv_word0.tlv_eng_id [3]);
tran (int_tlv_word8[27], \int_tlv_word8.dek_kim_entry.vf_num [0]);
tran (int_tlv_word9[27], \int_tlv_word9.dak_kim_entry.vf_num [0]);
tran (int_tlv_word42[27], \int_tlv_word42.unused [19]);
tran (key_header[27], \key_header.dak_key_ref [10]);
tran (int_tlv_word0[26], \int_tlv_word0.tlv_eng_id [2]);
tran (int_tlv_word8[26], \int_tlv_word8.dek_kim_entry.vf_valid [0]);
tran (int_tlv_word9[26], \int_tlv_word9.dak_kim_entry.vf_valid [0]);
tran (int_tlv_word42[26], \int_tlv_word42.unused [18]);
tran (key_header[26], \key_header.dak_key_ref [9]);
tran (int_tlv_word0[25], \int_tlv_word0.tlv_eng_id [1]);
tran (int_tlv_word8[25], \int_tlv_word8.unused [5]);
tran (int_tlv_word9[25], \int_tlv_word9.unused [7]);
tran (int_tlv_word42[25], \int_tlv_word42.unused [17]);
tran (key_header[25], \key_header.dak_key_ref [8]);
tran (int_tlv_word0[24], \int_tlv_word0.tlv_eng_id [0]);
tran (int_tlv_word8[24], \int_tlv_word8.unused [4]);
tran (int_tlv_word9[24], \int_tlv_word9.unused [6]);
tran (int_tlv_word42[24], \int_tlv_word42.unused [16]);
tran (key_header[24], \key_header.dak_key_ref [7]);
tran (int_tlv_word0[23], \int_tlv_word0.tlv_seq_num [7]);
tran (int_tlv_word8[23], \int_tlv_word8.unused [3]);
tran (int_tlv_word9[23], \int_tlv_word9.unused [5]);
tran (int_tlv_word42[23], \int_tlv_word42.unused [15]);
tran (key_header[23], \key_header.dak_key_ref [6]);
tran (int_tlv_word0[22], \int_tlv_word0.tlv_seq_num [6]);
tran (int_tlv_word8[22], \int_tlv_word8.unused [2]);
tran (int_tlv_word9[22], \int_tlv_word9.unused [4]);
tran (int_tlv_word42[22], \int_tlv_word42.unused [14]);
tran (key_header[22], \key_header.dak_key_ref [5]);
tran (int_tlv_word0[21], \int_tlv_word0.tlv_seq_num [5]);
tran (int_tlv_word8[21], \int_tlv_word8.unused [1]);
tran (int_tlv_word9[21], \int_tlv_word9.unused [3]);
tran (int_tlv_word42[21], \int_tlv_word42.unused [13]);
tran (key_header[21], \key_header.dak_key_ref [4]);
tran (int_tlv_word0[20], \int_tlv_word0.tlv_seq_num [4]);
tran (int_tlv_word8[20], \int_tlv_word8.unused [0]);
tran (int_tlv_word9[20], \int_tlv_word9.unused [2]);
tran (int_tlv_word42[20], \int_tlv_word42.unused [12]);
tran (key_header[20], \key_header.dak_key_ref [3]);
tran (int_tlv_word0[19], \int_tlv_word0.tlv_seq_num [3]);
tran (int_tlv_word8[19], \int_tlv_word8.missing_iv [0]);
tran (int_tlv_word9[19], \int_tlv_word9.unused [1]);
tran (int_tlv_word42[19], \int_tlv_word42.unused [11]);
tran (key_header[19], \key_header.dak_key_ref [2]);
tran (int_tlv_word0[18], \int_tlv_word0.tlv_seq_num [2]);
tran (int_tlv_word8[18], \int_tlv_word8.missing_guid [0]);
tran (int_tlv_word9[18], \int_tlv_word9.unused [0]);
tran (int_tlv_word42[18], \int_tlv_word42.unused [10]);
tran (key_header[18], \key_header.dak_key_ref [1]);
tran (int_tlv_word0[17], \int_tlv_word0.tlv_seq_num [1]);
tran (int_tlv_word8[17], \int_tlv_word8.validate_dek [0]);
tran (int_tlv_word9[17], \int_tlv_word9.validate_dak [0]);
tran (int_tlv_word42[17], \int_tlv_word42.unused [9]);
tran (key_header[17], \key_header.dak_key_ref [0]);
tran (int_tlv_word0[16], \int_tlv_word0.tlv_seq_num [0]);
tran (int_tlv_word8[16], \int_tlv_word8.vf_valid [0]);
tran (int_tlv_word9[16], \int_tlv_word9.vf_valid [0]);
tran (int_tlv_word42[16], \int_tlv_word42.unused [8]);
tran (key_header[16], \key_header.kdf_mode [1]);
tran (int_tlv_word0[15], \int_tlv_word0.tlv_len [7]);
tran (int_tlv_word8[15], \int_tlv_word8.pf_num [3]);
tran (int_tlv_word9[15], \int_tlv_word9.pf_num [3]);
tran (int_tlv_word42[15], \int_tlv_word42.unused [7]);
tran (key_header[15], \key_header.kdf_mode [0]);
tran (int_tlv_word0[14], \int_tlv_word0.tlv_len [6]);
tran (int_tlv_word8[14], \int_tlv_word8.pf_num [2]);
tran (int_tlv_word9[14], \int_tlv_word9.pf_num [2]);
tran (int_tlv_word42[14], \int_tlv_word42.unused [6]);
tran (key_header[14], \key_header.dek_key_op [0]);
tran (int_tlv_word0[13], \int_tlv_word0.tlv_len [5]);
tran (int_tlv_word8[13], \int_tlv_word8.pf_num [1]);
tran (int_tlv_word9[13], \int_tlv_word9.pf_num [1]);
tran (int_tlv_word42[13], \int_tlv_word42.unused [5]);
tran (key_header[13], \key_header.dek_key_ref [13]);
tran (int_tlv_word0[12], \int_tlv_word0.tlv_len [4]);
tran (int_tlv_word8[12], \int_tlv_word8.pf_num [0]);
tran (int_tlv_word9[12], \int_tlv_word9.pf_num [0]);
tran (int_tlv_word42[12], \int_tlv_word42.unused [4]);
tran (key_header[12], \key_header.dek_key_ref [12]);
tran (int_tlv_word0[11], \int_tlv_word0.tlv_len [3]);
tran (int_tlv_word8[11], \int_tlv_word8.vf_num [11]);
tran (int_tlv_word9[11], \int_tlv_word9.vf_num [11]);
tran (int_tlv_word42[11], \int_tlv_word42.unused [3]);
tran (key_header[11], \key_header.dek_key_ref [11]);
tran (int_tlv_word0[10], \int_tlv_word0.tlv_len [2]);
tran (int_tlv_word8[10], \int_tlv_word8.vf_num [10]);
tran (int_tlv_word9[10], \int_tlv_word9.vf_num [10]);
tran (int_tlv_word42[10], \int_tlv_word42.unused [2]);
tran (key_header[10], \key_header.dek_key_ref [10]);
tran (int_tlv_word0[9], \int_tlv_word0.tlv_len [1]);
tran (int_tlv_word8[9], \int_tlv_word8.vf_num [9]);
tran (int_tlv_word9[9], \int_tlv_word9.vf_num [9]);
tran (int_tlv_word42[9], \int_tlv_word42.unused [1]);
tran (key_header[9], \key_header.dek_key_ref [9]);
tran (int_tlv_word0[8], \int_tlv_word0.tlv_len [0]);
tran (int_tlv_word8[8], \int_tlv_word8.vf_num [8]);
tran (int_tlv_word9[8], \int_tlv_word9.vf_num [8]);
tran (int_tlv_word42[8], \int_tlv_word42.unused [0]);
tran (key_header[8], \key_header.dek_key_ref [8]);
tran (int_tlv_word0[7], \int_tlv_word0.tlv_type [7]);
tran (int_tlv_word8[7], \int_tlv_word8.vf_num [7]);
tran (int_tlv_word9[7], \int_tlv_word9.vf_num [7]);
tran (int_tlv_word42[7], \int_tlv_word42.error_code [7]);
tran (key_header[7], \key_header.dek_key_ref [7]);
tran (int_tlv_word0[6], \int_tlv_word0.tlv_type [6]);
tran (int_tlv_word8[6], \int_tlv_word8.vf_num [6]);
tran (int_tlv_word9[6], \int_tlv_word9.vf_num [6]);
tran (int_tlv_word42[6], \int_tlv_word42.error_code [6]);
tran (key_header[6], \key_header.dek_key_ref [6]);
tran (int_tlv_word0[5], \int_tlv_word0.tlv_type [5]);
tran (int_tlv_word8[5], \int_tlv_word8.vf_num [5]);
tran (int_tlv_word9[5], \int_tlv_word9.vf_num [5]);
tran (int_tlv_word42[5], \int_tlv_word42.error_code [5]);
tran (key_header[5], \key_header.dek_key_ref [5]);
tran (int_tlv_word0[4], \int_tlv_word0.tlv_type [4]);
tran (int_tlv_word8[4], \int_tlv_word8.vf_num [4]);
tran (int_tlv_word9[4], \int_tlv_word9.vf_num [4]);
tran (int_tlv_word42[4], \int_tlv_word42.error_code [4]);
tran (key_header[4], \key_header.dek_key_ref [4]);
tran (int_tlv_word0[3], \int_tlv_word0.tlv_type [3]);
tran (int_tlv_word8[3], \int_tlv_word8.vf_num [3]);
tran (int_tlv_word9[3], \int_tlv_word9.vf_num [3]);
tran (int_tlv_word42[3], \int_tlv_word42.error_code [3]);
tran (key_header[3], \key_header.dek_key_ref [3]);
tran (int_tlv_word0[2], \int_tlv_word0.tlv_type [2]);
tran (int_tlv_word8[2], \int_tlv_word8.vf_num [2]);
tran (int_tlv_word9[2], \int_tlv_word9.vf_num [2]);
tran (int_tlv_word42[2], \int_tlv_word42.error_code [2]);
tran (key_header[2], \key_header.dek_key_ref [2]);
tran (int_tlv_word0[1], \int_tlv_word0.tlv_type [1]);
tran (int_tlv_word8[1], \int_tlv_word8.vf_num [1]);
tran (int_tlv_word9[1], \int_tlv_word9.vf_num [1]);
tran (int_tlv_word42[1], \int_tlv_word42.error_code [1]);
tran (key_header[1], \key_header.dek_key_ref [1]);
tran (int_tlv_word0[0], \int_tlv_word0.tlv_type [0]);
tran (int_tlv_word8[0], \int_tlv_word8.vf_num [0]);
tran (int_tlv_word9[0], \int_tlv_word9.vf_num [0]);
tran (int_tlv_word42[0], \int_tlv_word42.error_code [0]);
tran (key_header[0], \key_header.dek_key_ref [0]);
tran (gcm_dak_cmd_in_nxt[0], \gcm_dak_cmd_in_nxt.op [0]);
tran (gcm_dak_cmd_in_nxt[1], \gcm_dak_cmd_in_nxt.op [1]);
tran (gcm_dak_cmd_in_nxt[2], \gcm_dak_cmd_in_nxt.op [2]);
tran (gcm_dak_cmd_in_nxt[3], \gcm_dak_cmd_in_nxt.iv [0]);
tran (gcm_dak_cmd_in_nxt[4], \gcm_dak_cmd_in_nxt.iv [1]);
tran (gcm_dak_cmd_in_nxt[5], \gcm_dak_cmd_in_nxt.iv [2]);
tran (gcm_dak_cmd_in_nxt[6], \gcm_dak_cmd_in_nxt.iv [3]);
tran (gcm_dak_cmd_in_nxt[7], \gcm_dak_cmd_in_nxt.iv [4]);
tran (gcm_dak_cmd_in_nxt[8], \gcm_dak_cmd_in_nxt.iv [5]);
tran (gcm_dak_cmd_in_nxt[9], \gcm_dak_cmd_in_nxt.iv [6]);
tran (gcm_dak_cmd_in_nxt[10], \gcm_dak_cmd_in_nxt.iv [7]);
tran (gcm_dak_cmd_in_nxt[11], \gcm_dak_cmd_in_nxt.iv [8]);
tran (gcm_dak_cmd_in_nxt[12], \gcm_dak_cmd_in_nxt.iv [9]);
tran (gcm_dak_cmd_in_nxt[13], \gcm_dak_cmd_in_nxt.iv [10]);
tran (gcm_dak_cmd_in_nxt[14], \gcm_dak_cmd_in_nxt.iv [11]);
tran (gcm_dak_cmd_in_nxt[15], \gcm_dak_cmd_in_nxt.iv [12]);
tran (gcm_dak_cmd_in_nxt[16], \gcm_dak_cmd_in_nxt.iv [13]);
tran (gcm_dak_cmd_in_nxt[17], \gcm_dak_cmd_in_nxt.iv [14]);
tran (gcm_dak_cmd_in_nxt[18], \gcm_dak_cmd_in_nxt.iv [15]);
tran (gcm_dak_cmd_in_nxt[19], \gcm_dak_cmd_in_nxt.iv [16]);
tran (gcm_dak_cmd_in_nxt[20], \gcm_dak_cmd_in_nxt.iv [17]);
tran (gcm_dak_cmd_in_nxt[21], \gcm_dak_cmd_in_nxt.iv [18]);
tran (gcm_dak_cmd_in_nxt[22], \gcm_dak_cmd_in_nxt.iv [19]);
tran (gcm_dak_cmd_in_nxt[23], \gcm_dak_cmd_in_nxt.iv [20]);
tran (gcm_dak_cmd_in_nxt[24], \gcm_dak_cmd_in_nxt.iv [21]);
tran (gcm_dak_cmd_in_nxt[25], \gcm_dak_cmd_in_nxt.iv [22]);
tran (gcm_dak_cmd_in_nxt[26], \gcm_dak_cmd_in_nxt.iv [23]);
tran (gcm_dak_cmd_in_nxt[27], \gcm_dak_cmd_in_nxt.iv [24]);
tran (gcm_dak_cmd_in_nxt[28], \gcm_dak_cmd_in_nxt.iv [25]);
tran (gcm_dak_cmd_in_nxt[29], \gcm_dak_cmd_in_nxt.iv [26]);
tran (gcm_dak_cmd_in_nxt[30], \gcm_dak_cmd_in_nxt.iv [27]);
tran (gcm_dak_cmd_in_nxt[31], \gcm_dak_cmd_in_nxt.iv [28]);
tran (gcm_dak_cmd_in_nxt[32], \gcm_dak_cmd_in_nxt.iv [29]);
tran (gcm_dak_cmd_in_nxt[33], \gcm_dak_cmd_in_nxt.iv [30]);
tran (gcm_dak_cmd_in_nxt[34], \gcm_dak_cmd_in_nxt.iv [31]);
tran (gcm_dak_cmd_in_nxt[35], \gcm_dak_cmd_in_nxt.iv [32]);
tran (gcm_dak_cmd_in_nxt[36], \gcm_dak_cmd_in_nxt.iv [33]);
tran (gcm_dak_cmd_in_nxt[37], \gcm_dak_cmd_in_nxt.iv [34]);
tran (gcm_dak_cmd_in_nxt[38], \gcm_dak_cmd_in_nxt.iv [35]);
tran (gcm_dak_cmd_in_nxt[39], \gcm_dak_cmd_in_nxt.iv [36]);
tran (gcm_dak_cmd_in_nxt[40], \gcm_dak_cmd_in_nxt.iv [37]);
tran (gcm_dak_cmd_in_nxt[41], \gcm_dak_cmd_in_nxt.iv [38]);
tran (gcm_dak_cmd_in_nxt[42], \gcm_dak_cmd_in_nxt.iv [39]);
tran (gcm_dak_cmd_in_nxt[43], \gcm_dak_cmd_in_nxt.iv [40]);
tran (gcm_dak_cmd_in_nxt[44], \gcm_dak_cmd_in_nxt.iv [41]);
tran (gcm_dak_cmd_in_nxt[45], \gcm_dak_cmd_in_nxt.iv [42]);
tran (gcm_dak_cmd_in_nxt[46], \gcm_dak_cmd_in_nxt.iv [43]);
tran (gcm_dak_cmd_in_nxt[47], \gcm_dak_cmd_in_nxt.iv [44]);
tran (gcm_dak_cmd_in_nxt[48], \gcm_dak_cmd_in_nxt.iv [45]);
tran (gcm_dak_cmd_in_nxt[49], \gcm_dak_cmd_in_nxt.iv [46]);
tran (gcm_dak_cmd_in_nxt[50], \gcm_dak_cmd_in_nxt.iv [47]);
tran (gcm_dak_cmd_in_nxt[51], \gcm_dak_cmd_in_nxt.iv [48]);
tran (gcm_dak_cmd_in_nxt[52], \gcm_dak_cmd_in_nxt.iv [49]);
tran (gcm_dak_cmd_in_nxt[53], \gcm_dak_cmd_in_nxt.iv [50]);
tran (gcm_dak_cmd_in_nxt[54], \gcm_dak_cmd_in_nxt.iv [51]);
tran (gcm_dak_cmd_in_nxt[55], \gcm_dak_cmd_in_nxt.iv [52]);
tran (gcm_dak_cmd_in_nxt[56], \gcm_dak_cmd_in_nxt.iv [53]);
tran (gcm_dak_cmd_in_nxt[57], \gcm_dak_cmd_in_nxt.iv [54]);
tran (gcm_dak_cmd_in_nxt[58], \gcm_dak_cmd_in_nxt.iv [55]);
tran (gcm_dak_cmd_in_nxt[59], \gcm_dak_cmd_in_nxt.iv [56]);
tran (gcm_dak_cmd_in_nxt[60], \gcm_dak_cmd_in_nxt.iv [57]);
tran (gcm_dak_cmd_in_nxt[61], \gcm_dak_cmd_in_nxt.iv [58]);
tran (gcm_dak_cmd_in_nxt[62], \gcm_dak_cmd_in_nxt.iv [59]);
tran (gcm_dak_cmd_in_nxt[63], \gcm_dak_cmd_in_nxt.iv [60]);
tran (gcm_dak_cmd_in_nxt[64], \gcm_dak_cmd_in_nxt.iv [61]);
tran (gcm_dak_cmd_in_nxt[65], \gcm_dak_cmd_in_nxt.iv [62]);
tran (gcm_dak_cmd_in_nxt[66], \gcm_dak_cmd_in_nxt.iv [63]);
tran (gcm_dak_cmd_in_nxt[67], \gcm_dak_cmd_in_nxt.iv [64]);
tran (gcm_dak_cmd_in_nxt[68], \gcm_dak_cmd_in_nxt.iv [65]);
tran (gcm_dak_cmd_in_nxt[69], \gcm_dak_cmd_in_nxt.iv [66]);
tran (gcm_dak_cmd_in_nxt[70], \gcm_dak_cmd_in_nxt.iv [67]);
tran (gcm_dak_cmd_in_nxt[71], \gcm_dak_cmd_in_nxt.iv [68]);
tran (gcm_dak_cmd_in_nxt[72], \gcm_dak_cmd_in_nxt.iv [69]);
tran (gcm_dak_cmd_in_nxt[73], \gcm_dak_cmd_in_nxt.iv [70]);
tran (gcm_dak_cmd_in_nxt[74], \gcm_dak_cmd_in_nxt.iv [71]);
tran (gcm_dak_cmd_in_nxt[75], \gcm_dak_cmd_in_nxt.iv [72]);
tran (gcm_dak_cmd_in_nxt[76], \gcm_dak_cmd_in_nxt.iv [73]);
tran (gcm_dak_cmd_in_nxt[77], \gcm_dak_cmd_in_nxt.iv [74]);
tran (gcm_dak_cmd_in_nxt[78], \gcm_dak_cmd_in_nxt.iv [75]);
tran (gcm_dak_cmd_in_nxt[79], \gcm_dak_cmd_in_nxt.iv [76]);
tran (gcm_dak_cmd_in_nxt[80], \gcm_dak_cmd_in_nxt.iv [77]);
tran (gcm_dak_cmd_in_nxt[81], \gcm_dak_cmd_in_nxt.iv [78]);
tran (gcm_dak_cmd_in_nxt[82], \gcm_dak_cmd_in_nxt.iv [79]);
tran (gcm_dak_cmd_in_nxt[83], \gcm_dak_cmd_in_nxt.iv [80]);
tran (gcm_dak_cmd_in_nxt[84], \gcm_dak_cmd_in_nxt.iv [81]);
tran (gcm_dak_cmd_in_nxt[85], \gcm_dak_cmd_in_nxt.iv [82]);
tran (gcm_dak_cmd_in_nxt[86], \gcm_dak_cmd_in_nxt.iv [83]);
tran (gcm_dak_cmd_in_nxt[87], \gcm_dak_cmd_in_nxt.iv [84]);
tran (gcm_dak_cmd_in_nxt[88], \gcm_dak_cmd_in_nxt.iv [85]);
tran (gcm_dak_cmd_in_nxt[89], \gcm_dak_cmd_in_nxt.iv [86]);
tran (gcm_dak_cmd_in_nxt[90], \gcm_dak_cmd_in_nxt.iv [87]);
tran (gcm_dak_cmd_in_nxt[91], \gcm_dak_cmd_in_nxt.iv [88]);
tran (gcm_dak_cmd_in_nxt[92], \gcm_dak_cmd_in_nxt.iv [89]);
tran (gcm_dak_cmd_in_nxt[93], \gcm_dak_cmd_in_nxt.iv [90]);
tran (gcm_dak_cmd_in_nxt[94], \gcm_dak_cmd_in_nxt.iv [91]);
tran (gcm_dak_cmd_in_nxt[95], \gcm_dak_cmd_in_nxt.iv [92]);
tran (gcm_dak_cmd_in_nxt[96], \gcm_dak_cmd_in_nxt.iv [93]);
tran (gcm_dak_cmd_in_nxt[97], \gcm_dak_cmd_in_nxt.iv [94]);
tran (gcm_dak_cmd_in_nxt[98], \gcm_dak_cmd_in_nxt.iv [95]);
tran (gcm_dak_cmd_in_nxt[99], \gcm_dak_cmd_in_nxt.key1 [0]);
tran (gcm_dak_cmd_in_nxt[100], \gcm_dak_cmd_in_nxt.key1 [1]);
tran (gcm_dak_cmd_in_nxt[101], \gcm_dak_cmd_in_nxt.key1 [2]);
tran (gcm_dak_cmd_in_nxt[102], \gcm_dak_cmd_in_nxt.key1 [3]);
tran (gcm_dak_cmd_in_nxt[103], \gcm_dak_cmd_in_nxt.key1 [4]);
tran (gcm_dak_cmd_in_nxt[104], \gcm_dak_cmd_in_nxt.key1 [5]);
tran (gcm_dak_cmd_in_nxt[105], \gcm_dak_cmd_in_nxt.key1 [6]);
tran (gcm_dak_cmd_in_nxt[106], \gcm_dak_cmd_in_nxt.key1 [7]);
tran (gcm_dak_cmd_in_nxt[107], \gcm_dak_cmd_in_nxt.key1 [8]);
tran (gcm_dak_cmd_in_nxt[108], \gcm_dak_cmd_in_nxt.key1 [9]);
tran (gcm_dak_cmd_in_nxt[109], \gcm_dak_cmd_in_nxt.key1 [10]);
tran (gcm_dak_cmd_in_nxt[110], \gcm_dak_cmd_in_nxt.key1 [11]);
tran (gcm_dak_cmd_in_nxt[111], \gcm_dak_cmd_in_nxt.key1 [12]);
tran (gcm_dak_cmd_in_nxt[112], \gcm_dak_cmd_in_nxt.key1 [13]);
tran (gcm_dak_cmd_in_nxt[113], \gcm_dak_cmd_in_nxt.key1 [14]);
tran (gcm_dak_cmd_in_nxt[114], \gcm_dak_cmd_in_nxt.key1 [15]);
tran (gcm_dak_cmd_in_nxt[115], \gcm_dak_cmd_in_nxt.key1 [16]);
tran (gcm_dak_cmd_in_nxt[116], \gcm_dak_cmd_in_nxt.key1 [17]);
tran (gcm_dak_cmd_in_nxt[117], \gcm_dak_cmd_in_nxt.key1 [18]);
tran (gcm_dak_cmd_in_nxt[118], \gcm_dak_cmd_in_nxt.key1 [19]);
tran (gcm_dak_cmd_in_nxt[119], \gcm_dak_cmd_in_nxt.key1 [20]);
tran (gcm_dak_cmd_in_nxt[120], \gcm_dak_cmd_in_nxt.key1 [21]);
tran (gcm_dak_cmd_in_nxt[121], \gcm_dak_cmd_in_nxt.key1 [22]);
tran (gcm_dak_cmd_in_nxt[122], \gcm_dak_cmd_in_nxt.key1 [23]);
tran (gcm_dak_cmd_in_nxt[123], \gcm_dak_cmd_in_nxt.key1 [24]);
tran (gcm_dak_cmd_in_nxt[124], \gcm_dak_cmd_in_nxt.key1 [25]);
tran (gcm_dak_cmd_in_nxt[125], \gcm_dak_cmd_in_nxt.key1 [26]);
tran (gcm_dak_cmd_in_nxt[126], \gcm_dak_cmd_in_nxt.key1 [27]);
tran (gcm_dak_cmd_in_nxt[127], \gcm_dak_cmd_in_nxt.key1 [28]);
tran (gcm_dak_cmd_in_nxt[128], \gcm_dak_cmd_in_nxt.key1 [29]);
tran (gcm_dak_cmd_in_nxt[129], \gcm_dak_cmd_in_nxt.key1 [30]);
tran (gcm_dak_cmd_in_nxt[130], \gcm_dak_cmd_in_nxt.key1 [31]);
tran (gcm_dak_cmd_in_nxt[131], \gcm_dak_cmd_in_nxt.key1 [32]);
tran (gcm_dak_cmd_in_nxt[132], \gcm_dak_cmd_in_nxt.key1 [33]);
tran (gcm_dak_cmd_in_nxt[133], \gcm_dak_cmd_in_nxt.key1 [34]);
tran (gcm_dak_cmd_in_nxt[134], \gcm_dak_cmd_in_nxt.key1 [35]);
tran (gcm_dak_cmd_in_nxt[135], \gcm_dak_cmd_in_nxt.key1 [36]);
tran (gcm_dak_cmd_in_nxt[136], \gcm_dak_cmd_in_nxt.key1 [37]);
tran (gcm_dak_cmd_in_nxt[137], \gcm_dak_cmd_in_nxt.key1 [38]);
tran (gcm_dak_cmd_in_nxt[138], \gcm_dak_cmd_in_nxt.key1 [39]);
tran (gcm_dak_cmd_in_nxt[139], \gcm_dak_cmd_in_nxt.key1 [40]);
tran (gcm_dak_cmd_in_nxt[140], \gcm_dak_cmd_in_nxt.key1 [41]);
tran (gcm_dak_cmd_in_nxt[141], \gcm_dak_cmd_in_nxt.key1 [42]);
tran (gcm_dak_cmd_in_nxt[142], \gcm_dak_cmd_in_nxt.key1 [43]);
tran (gcm_dak_cmd_in_nxt[143], \gcm_dak_cmd_in_nxt.key1 [44]);
tran (gcm_dak_cmd_in_nxt[144], \gcm_dak_cmd_in_nxt.key1 [45]);
tran (gcm_dak_cmd_in_nxt[145], \gcm_dak_cmd_in_nxt.key1 [46]);
tran (gcm_dak_cmd_in_nxt[146], \gcm_dak_cmd_in_nxt.key1 [47]);
tran (gcm_dak_cmd_in_nxt[147], \gcm_dak_cmd_in_nxt.key1 [48]);
tran (gcm_dak_cmd_in_nxt[148], \gcm_dak_cmd_in_nxt.key1 [49]);
tran (gcm_dak_cmd_in_nxt[149], \gcm_dak_cmd_in_nxt.key1 [50]);
tran (gcm_dak_cmd_in_nxt[150], \gcm_dak_cmd_in_nxt.key1 [51]);
tran (gcm_dak_cmd_in_nxt[151], \gcm_dak_cmd_in_nxt.key1 [52]);
tran (gcm_dak_cmd_in_nxt[152], \gcm_dak_cmd_in_nxt.key1 [53]);
tran (gcm_dak_cmd_in_nxt[153], \gcm_dak_cmd_in_nxt.key1 [54]);
tran (gcm_dak_cmd_in_nxt[154], \gcm_dak_cmd_in_nxt.key1 [55]);
tran (gcm_dak_cmd_in_nxt[155], \gcm_dak_cmd_in_nxt.key1 [56]);
tran (gcm_dak_cmd_in_nxt[156], \gcm_dak_cmd_in_nxt.key1 [57]);
tran (gcm_dak_cmd_in_nxt[157], \gcm_dak_cmd_in_nxt.key1 [58]);
tran (gcm_dak_cmd_in_nxt[158], \gcm_dak_cmd_in_nxt.key1 [59]);
tran (gcm_dak_cmd_in_nxt[159], \gcm_dak_cmd_in_nxt.key1 [60]);
tran (gcm_dak_cmd_in_nxt[160], \gcm_dak_cmd_in_nxt.key1 [61]);
tran (gcm_dak_cmd_in_nxt[161], \gcm_dak_cmd_in_nxt.key1 [62]);
tran (gcm_dak_cmd_in_nxt[162], \gcm_dak_cmd_in_nxt.key1 [63]);
tran (gcm_dak_cmd_in_nxt[163], \gcm_dak_cmd_in_nxt.key1 [64]);
tran (gcm_dak_cmd_in_nxt[164], \gcm_dak_cmd_in_nxt.key1 [65]);
tran (gcm_dak_cmd_in_nxt[165], \gcm_dak_cmd_in_nxt.key1 [66]);
tran (gcm_dak_cmd_in_nxt[166], \gcm_dak_cmd_in_nxt.key1 [67]);
tran (gcm_dak_cmd_in_nxt[167], \gcm_dak_cmd_in_nxt.key1 [68]);
tran (gcm_dak_cmd_in_nxt[168], \gcm_dak_cmd_in_nxt.key1 [69]);
tran (gcm_dak_cmd_in_nxt[169], \gcm_dak_cmd_in_nxt.key1 [70]);
tran (gcm_dak_cmd_in_nxt[170], \gcm_dak_cmd_in_nxt.key1 [71]);
tran (gcm_dak_cmd_in_nxt[171], \gcm_dak_cmd_in_nxt.key1 [72]);
tran (gcm_dak_cmd_in_nxt[172], \gcm_dak_cmd_in_nxt.key1 [73]);
tran (gcm_dak_cmd_in_nxt[173], \gcm_dak_cmd_in_nxt.key1 [74]);
tran (gcm_dak_cmd_in_nxt[174], \gcm_dak_cmd_in_nxt.key1 [75]);
tran (gcm_dak_cmd_in_nxt[175], \gcm_dak_cmd_in_nxt.key1 [76]);
tran (gcm_dak_cmd_in_nxt[176], \gcm_dak_cmd_in_nxt.key1 [77]);
tran (gcm_dak_cmd_in_nxt[177], \gcm_dak_cmd_in_nxt.key1 [78]);
tran (gcm_dak_cmd_in_nxt[178], \gcm_dak_cmd_in_nxt.key1 [79]);
tran (gcm_dak_cmd_in_nxt[179], \gcm_dak_cmd_in_nxt.key1 [80]);
tran (gcm_dak_cmd_in_nxt[180], \gcm_dak_cmd_in_nxt.key1 [81]);
tran (gcm_dak_cmd_in_nxt[181], \gcm_dak_cmd_in_nxt.key1 [82]);
tran (gcm_dak_cmd_in_nxt[182], \gcm_dak_cmd_in_nxt.key1 [83]);
tran (gcm_dak_cmd_in_nxt[183], \gcm_dak_cmd_in_nxt.key1 [84]);
tran (gcm_dak_cmd_in_nxt[184], \gcm_dak_cmd_in_nxt.key1 [85]);
tran (gcm_dak_cmd_in_nxt[185], \gcm_dak_cmd_in_nxt.key1 [86]);
tran (gcm_dak_cmd_in_nxt[186], \gcm_dak_cmd_in_nxt.key1 [87]);
tran (gcm_dak_cmd_in_nxt[187], \gcm_dak_cmd_in_nxt.key1 [88]);
tran (gcm_dak_cmd_in_nxt[188], \gcm_dak_cmd_in_nxt.key1 [89]);
tran (gcm_dak_cmd_in_nxt[189], \gcm_dak_cmd_in_nxt.key1 [90]);
tran (gcm_dak_cmd_in_nxt[190], \gcm_dak_cmd_in_nxt.key1 [91]);
tran (gcm_dak_cmd_in_nxt[191], \gcm_dak_cmd_in_nxt.key1 [92]);
tran (gcm_dak_cmd_in_nxt[192], \gcm_dak_cmd_in_nxt.key1 [93]);
tran (gcm_dak_cmd_in_nxt[193], \gcm_dak_cmd_in_nxt.key1 [94]);
tran (gcm_dak_cmd_in_nxt[194], \gcm_dak_cmd_in_nxt.key1 [95]);
tran (gcm_dak_cmd_in_nxt[195], \gcm_dak_cmd_in_nxt.key1 [96]);
tran (gcm_dak_cmd_in_nxt[196], \gcm_dak_cmd_in_nxt.key1 [97]);
tran (gcm_dak_cmd_in_nxt[197], \gcm_dak_cmd_in_nxt.key1 [98]);
tran (gcm_dak_cmd_in_nxt[198], \gcm_dak_cmd_in_nxt.key1 [99]);
tran (gcm_dak_cmd_in_nxt[199], \gcm_dak_cmd_in_nxt.key1 [100]);
tran (gcm_dak_cmd_in_nxt[200], \gcm_dak_cmd_in_nxt.key1 [101]);
tran (gcm_dak_cmd_in_nxt[201], \gcm_dak_cmd_in_nxt.key1 [102]);
tran (gcm_dak_cmd_in_nxt[202], \gcm_dak_cmd_in_nxt.key1 [103]);
tran (gcm_dak_cmd_in_nxt[203], \gcm_dak_cmd_in_nxt.key1 [104]);
tran (gcm_dak_cmd_in_nxt[204], \gcm_dak_cmd_in_nxt.key1 [105]);
tran (gcm_dak_cmd_in_nxt[205], \gcm_dak_cmd_in_nxt.key1 [106]);
tran (gcm_dak_cmd_in_nxt[206], \gcm_dak_cmd_in_nxt.key1 [107]);
tran (gcm_dak_cmd_in_nxt[207], \gcm_dak_cmd_in_nxt.key1 [108]);
tran (gcm_dak_cmd_in_nxt[208], \gcm_dak_cmd_in_nxt.key1 [109]);
tran (gcm_dak_cmd_in_nxt[209], \gcm_dak_cmd_in_nxt.key1 [110]);
tran (gcm_dak_cmd_in_nxt[210], \gcm_dak_cmd_in_nxt.key1 [111]);
tran (gcm_dak_cmd_in_nxt[211], \gcm_dak_cmd_in_nxt.key1 [112]);
tran (gcm_dak_cmd_in_nxt[212], \gcm_dak_cmd_in_nxt.key1 [113]);
tran (gcm_dak_cmd_in_nxt[213], \gcm_dak_cmd_in_nxt.key1 [114]);
tran (gcm_dak_cmd_in_nxt[214], \gcm_dak_cmd_in_nxt.key1 [115]);
tran (gcm_dak_cmd_in_nxt[215], \gcm_dak_cmd_in_nxt.key1 [116]);
tran (gcm_dak_cmd_in_nxt[216], \gcm_dak_cmd_in_nxt.key1 [117]);
tran (gcm_dak_cmd_in_nxt[217], \gcm_dak_cmd_in_nxt.key1 [118]);
tran (gcm_dak_cmd_in_nxt[218], \gcm_dak_cmd_in_nxt.key1 [119]);
tran (gcm_dak_cmd_in_nxt[219], \gcm_dak_cmd_in_nxt.key1 [120]);
tran (gcm_dak_cmd_in_nxt[220], \gcm_dak_cmd_in_nxt.key1 [121]);
tran (gcm_dak_cmd_in_nxt[221], \gcm_dak_cmd_in_nxt.key1 [122]);
tran (gcm_dak_cmd_in_nxt[222], \gcm_dak_cmd_in_nxt.key1 [123]);
tran (gcm_dak_cmd_in_nxt[223], \gcm_dak_cmd_in_nxt.key1 [124]);
tran (gcm_dak_cmd_in_nxt[224], \gcm_dak_cmd_in_nxt.key1 [125]);
tran (gcm_dak_cmd_in_nxt[225], \gcm_dak_cmd_in_nxt.key1 [126]);
tran (gcm_dak_cmd_in_nxt[226], \gcm_dak_cmd_in_nxt.key1 [127]);
tran (gcm_dak_cmd_in_nxt[227], \gcm_dak_cmd_in_nxt.key1 [128]);
tran (gcm_dak_cmd_in_nxt[228], \gcm_dak_cmd_in_nxt.key1 [129]);
tran (gcm_dak_cmd_in_nxt[229], \gcm_dak_cmd_in_nxt.key1 [130]);
tran (gcm_dak_cmd_in_nxt[230], \gcm_dak_cmd_in_nxt.key1 [131]);
tran (gcm_dak_cmd_in_nxt[231], \gcm_dak_cmd_in_nxt.key1 [132]);
tran (gcm_dak_cmd_in_nxt[232], \gcm_dak_cmd_in_nxt.key1 [133]);
tran (gcm_dak_cmd_in_nxt[233], \gcm_dak_cmd_in_nxt.key1 [134]);
tran (gcm_dak_cmd_in_nxt[234], \gcm_dak_cmd_in_nxt.key1 [135]);
tran (gcm_dak_cmd_in_nxt[235], \gcm_dak_cmd_in_nxt.key1 [136]);
tran (gcm_dak_cmd_in_nxt[236], \gcm_dak_cmd_in_nxt.key1 [137]);
tran (gcm_dak_cmd_in_nxt[237], \gcm_dak_cmd_in_nxt.key1 [138]);
tran (gcm_dak_cmd_in_nxt[238], \gcm_dak_cmd_in_nxt.key1 [139]);
tran (gcm_dak_cmd_in_nxt[239], \gcm_dak_cmd_in_nxt.key1 [140]);
tran (gcm_dak_cmd_in_nxt[240], \gcm_dak_cmd_in_nxt.key1 [141]);
tran (gcm_dak_cmd_in_nxt[241], \gcm_dak_cmd_in_nxt.key1 [142]);
tran (gcm_dak_cmd_in_nxt[242], \gcm_dak_cmd_in_nxt.key1 [143]);
tran (gcm_dak_cmd_in_nxt[243], \gcm_dak_cmd_in_nxt.key1 [144]);
tran (gcm_dak_cmd_in_nxt[244], \gcm_dak_cmd_in_nxt.key1 [145]);
tran (gcm_dak_cmd_in_nxt[245], \gcm_dak_cmd_in_nxt.key1 [146]);
tran (gcm_dak_cmd_in_nxt[246], \gcm_dak_cmd_in_nxt.key1 [147]);
tran (gcm_dak_cmd_in_nxt[247], \gcm_dak_cmd_in_nxt.key1 [148]);
tran (gcm_dak_cmd_in_nxt[248], \gcm_dak_cmd_in_nxt.key1 [149]);
tran (gcm_dak_cmd_in_nxt[249], \gcm_dak_cmd_in_nxt.key1 [150]);
tran (gcm_dak_cmd_in_nxt[250], \gcm_dak_cmd_in_nxt.key1 [151]);
tran (gcm_dak_cmd_in_nxt[251], \gcm_dak_cmd_in_nxt.key1 [152]);
tran (gcm_dak_cmd_in_nxt[252], \gcm_dak_cmd_in_nxt.key1 [153]);
tran (gcm_dak_cmd_in_nxt[253], \gcm_dak_cmd_in_nxt.key1 [154]);
tran (gcm_dak_cmd_in_nxt[254], \gcm_dak_cmd_in_nxt.key1 [155]);
tran (gcm_dak_cmd_in_nxt[255], \gcm_dak_cmd_in_nxt.key1 [156]);
tran (gcm_dak_cmd_in_nxt[256], \gcm_dak_cmd_in_nxt.key1 [157]);
tran (gcm_dak_cmd_in_nxt[257], \gcm_dak_cmd_in_nxt.key1 [158]);
tran (gcm_dak_cmd_in_nxt[258], \gcm_dak_cmd_in_nxt.key1 [159]);
tran (gcm_dak_cmd_in_nxt[259], \gcm_dak_cmd_in_nxt.key1 [160]);
tran (gcm_dak_cmd_in_nxt[260], \gcm_dak_cmd_in_nxt.key1 [161]);
tran (gcm_dak_cmd_in_nxt[261], \gcm_dak_cmd_in_nxt.key1 [162]);
tran (gcm_dak_cmd_in_nxt[262], \gcm_dak_cmd_in_nxt.key1 [163]);
tran (gcm_dak_cmd_in_nxt[263], \gcm_dak_cmd_in_nxt.key1 [164]);
tran (gcm_dak_cmd_in_nxt[264], \gcm_dak_cmd_in_nxt.key1 [165]);
tran (gcm_dak_cmd_in_nxt[265], \gcm_dak_cmd_in_nxt.key1 [166]);
tran (gcm_dak_cmd_in_nxt[266], \gcm_dak_cmd_in_nxt.key1 [167]);
tran (gcm_dak_cmd_in_nxt[267], \gcm_dak_cmd_in_nxt.key1 [168]);
tran (gcm_dak_cmd_in_nxt[268], \gcm_dak_cmd_in_nxt.key1 [169]);
tran (gcm_dak_cmd_in_nxt[269], \gcm_dak_cmd_in_nxt.key1 [170]);
tran (gcm_dak_cmd_in_nxt[270], \gcm_dak_cmd_in_nxt.key1 [171]);
tran (gcm_dak_cmd_in_nxt[271], \gcm_dak_cmd_in_nxt.key1 [172]);
tran (gcm_dak_cmd_in_nxt[272], \gcm_dak_cmd_in_nxt.key1 [173]);
tran (gcm_dak_cmd_in_nxt[273], \gcm_dak_cmd_in_nxt.key1 [174]);
tran (gcm_dak_cmd_in_nxt[274], \gcm_dak_cmd_in_nxt.key1 [175]);
tran (gcm_dak_cmd_in_nxt[275], \gcm_dak_cmd_in_nxt.key1 [176]);
tran (gcm_dak_cmd_in_nxt[276], \gcm_dak_cmd_in_nxt.key1 [177]);
tran (gcm_dak_cmd_in_nxt[277], \gcm_dak_cmd_in_nxt.key1 [178]);
tran (gcm_dak_cmd_in_nxt[278], \gcm_dak_cmd_in_nxt.key1 [179]);
tran (gcm_dak_cmd_in_nxt[279], \gcm_dak_cmd_in_nxt.key1 [180]);
tran (gcm_dak_cmd_in_nxt[280], \gcm_dak_cmd_in_nxt.key1 [181]);
tran (gcm_dak_cmd_in_nxt[281], \gcm_dak_cmd_in_nxt.key1 [182]);
tran (gcm_dak_cmd_in_nxt[282], \gcm_dak_cmd_in_nxt.key1 [183]);
tran (gcm_dak_cmd_in_nxt[283], \gcm_dak_cmd_in_nxt.key1 [184]);
tran (gcm_dak_cmd_in_nxt[284], \gcm_dak_cmd_in_nxt.key1 [185]);
tran (gcm_dak_cmd_in_nxt[285], \gcm_dak_cmd_in_nxt.key1 [186]);
tran (gcm_dak_cmd_in_nxt[286], \gcm_dak_cmd_in_nxt.key1 [187]);
tran (gcm_dak_cmd_in_nxt[287], \gcm_dak_cmd_in_nxt.key1 [188]);
tran (gcm_dak_cmd_in_nxt[288], \gcm_dak_cmd_in_nxt.key1 [189]);
tran (gcm_dak_cmd_in_nxt[289], \gcm_dak_cmd_in_nxt.key1 [190]);
tran (gcm_dak_cmd_in_nxt[290], \gcm_dak_cmd_in_nxt.key1 [191]);
tran (gcm_dak_cmd_in_nxt[291], \gcm_dak_cmd_in_nxt.key1 [192]);
tran (gcm_dak_cmd_in_nxt[292], \gcm_dak_cmd_in_nxt.key1 [193]);
tran (gcm_dak_cmd_in_nxt[293], \gcm_dak_cmd_in_nxt.key1 [194]);
tran (gcm_dak_cmd_in_nxt[294], \gcm_dak_cmd_in_nxt.key1 [195]);
tran (gcm_dak_cmd_in_nxt[295], \gcm_dak_cmd_in_nxt.key1 [196]);
tran (gcm_dak_cmd_in_nxt[296], \gcm_dak_cmd_in_nxt.key1 [197]);
tran (gcm_dak_cmd_in_nxt[297], \gcm_dak_cmd_in_nxt.key1 [198]);
tran (gcm_dak_cmd_in_nxt[298], \gcm_dak_cmd_in_nxt.key1 [199]);
tran (gcm_dak_cmd_in_nxt[299], \gcm_dak_cmd_in_nxt.key1 [200]);
tran (gcm_dak_cmd_in_nxt[300], \gcm_dak_cmd_in_nxt.key1 [201]);
tran (gcm_dak_cmd_in_nxt[301], \gcm_dak_cmd_in_nxt.key1 [202]);
tran (gcm_dak_cmd_in_nxt[302], \gcm_dak_cmd_in_nxt.key1 [203]);
tran (gcm_dak_cmd_in_nxt[303], \gcm_dak_cmd_in_nxt.key1 [204]);
tran (gcm_dak_cmd_in_nxt[304], \gcm_dak_cmd_in_nxt.key1 [205]);
tran (gcm_dak_cmd_in_nxt[305], \gcm_dak_cmd_in_nxt.key1 [206]);
tran (gcm_dak_cmd_in_nxt[306], \gcm_dak_cmd_in_nxt.key1 [207]);
tran (gcm_dak_cmd_in_nxt[307], \gcm_dak_cmd_in_nxt.key1 [208]);
tran (gcm_dak_cmd_in_nxt[308], \gcm_dak_cmd_in_nxt.key1 [209]);
tran (gcm_dak_cmd_in_nxt[309], \gcm_dak_cmd_in_nxt.key1 [210]);
tran (gcm_dak_cmd_in_nxt[310], \gcm_dak_cmd_in_nxt.key1 [211]);
tran (gcm_dak_cmd_in_nxt[311], \gcm_dak_cmd_in_nxt.key1 [212]);
tran (gcm_dak_cmd_in_nxt[312], \gcm_dak_cmd_in_nxt.key1 [213]);
tran (gcm_dak_cmd_in_nxt[313], \gcm_dak_cmd_in_nxt.key1 [214]);
tran (gcm_dak_cmd_in_nxt[314], \gcm_dak_cmd_in_nxt.key1 [215]);
tran (gcm_dak_cmd_in_nxt[315], \gcm_dak_cmd_in_nxt.key1 [216]);
tran (gcm_dak_cmd_in_nxt[316], \gcm_dak_cmd_in_nxt.key1 [217]);
tran (gcm_dak_cmd_in_nxt[317], \gcm_dak_cmd_in_nxt.key1 [218]);
tran (gcm_dak_cmd_in_nxt[318], \gcm_dak_cmd_in_nxt.key1 [219]);
tran (gcm_dak_cmd_in_nxt[319], \gcm_dak_cmd_in_nxt.key1 [220]);
tran (gcm_dak_cmd_in_nxt[320], \gcm_dak_cmd_in_nxt.key1 [221]);
tran (gcm_dak_cmd_in_nxt[321], \gcm_dak_cmd_in_nxt.key1 [222]);
tran (gcm_dak_cmd_in_nxt[322], \gcm_dak_cmd_in_nxt.key1 [223]);
tran (gcm_dak_cmd_in_nxt[323], \gcm_dak_cmd_in_nxt.key1 [224]);
tran (gcm_dak_cmd_in_nxt[324], \gcm_dak_cmd_in_nxt.key1 [225]);
tran (gcm_dak_cmd_in_nxt[325], \gcm_dak_cmd_in_nxt.key1 [226]);
tran (gcm_dak_cmd_in_nxt[326], \gcm_dak_cmd_in_nxt.key1 [227]);
tran (gcm_dak_cmd_in_nxt[327], \gcm_dak_cmd_in_nxt.key1 [228]);
tran (gcm_dak_cmd_in_nxt[328], \gcm_dak_cmd_in_nxt.key1 [229]);
tran (gcm_dak_cmd_in_nxt[329], \gcm_dak_cmd_in_nxt.key1 [230]);
tran (gcm_dak_cmd_in_nxt[330], \gcm_dak_cmd_in_nxt.key1 [231]);
tran (gcm_dak_cmd_in_nxt[331], \gcm_dak_cmd_in_nxt.key1 [232]);
tran (gcm_dak_cmd_in_nxt[332], \gcm_dak_cmd_in_nxt.key1 [233]);
tran (gcm_dak_cmd_in_nxt[333], \gcm_dak_cmd_in_nxt.key1 [234]);
tran (gcm_dak_cmd_in_nxt[334], \gcm_dak_cmd_in_nxt.key1 [235]);
tran (gcm_dak_cmd_in_nxt[335], \gcm_dak_cmd_in_nxt.key1 [236]);
tran (gcm_dak_cmd_in_nxt[336], \gcm_dak_cmd_in_nxt.key1 [237]);
tran (gcm_dak_cmd_in_nxt[337], \gcm_dak_cmd_in_nxt.key1 [238]);
tran (gcm_dak_cmd_in_nxt[338], \gcm_dak_cmd_in_nxt.key1 [239]);
tran (gcm_dak_cmd_in_nxt[339], \gcm_dak_cmd_in_nxt.key1 [240]);
tran (gcm_dak_cmd_in_nxt[340], \gcm_dak_cmd_in_nxt.key1 [241]);
tran (gcm_dak_cmd_in_nxt[341], \gcm_dak_cmd_in_nxt.key1 [242]);
tran (gcm_dak_cmd_in_nxt[342], \gcm_dak_cmd_in_nxt.key1 [243]);
tran (gcm_dak_cmd_in_nxt[343], \gcm_dak_cmd_in_nxt.key1 [244]);
tran (gcm_dak_cmd_in_nxt[344], \gcm_dak_cmd_in_nxt.key1 [245]);
tran (gcm_dak_cmd_in_nxt[345], \gcm_dak_cmd_in_nxt.key1 [246]);
tran (gcm_dak_cmd_in_nxt[346], \gcm_dak_cmd_in_nxt.key1 [247]);
tran (gcm_dak_cmd_in_nxt[347], \gcm_dak_cmd_in_nxt.key1 [248]);
tran (gcm_dak_cmd_in_nxt[348], \gcm_dak_cmd_in_nxt.key1 [249]);
tran (gcm_dak_cmd_in_nxt[349], \gcm_dak_cmd_in_nxt.key1 [250]);
tran (gcm_dak_cmd_in_nxt[350], \gcm_dak_cmd_in_nxt.key1 [251]);
tran (gcm_dak_cmd_in_nxt[351], \gcm_dak_cmd_in_nxt.key1 [252]);
tran (gcm_dak_cmd_in_nxt[352], \gcm_dak_cmd_in_nxt.key1 [253]);
tran (gcm_dak_cmd_in_nxt[353], \gcm_dak_cmd_in_nxt.key1 [254]);
tran (gcm_dak_cmd_in_nxt[354], \gcm_dak_cmd_in_nxt.key1 [255]);
tran (gcm_dak_cmd_in_nxt[355], \gcm_dak_cmd_in_nxt.key0 [0]);
tran (gcm_dak_cmd_in_nxt[356], \gcm_dak_cmd_in_nxt.key0 [1]);
tran (gcm_dak_cmd_in_nxt[357], \gcm_dak_cmd_in_nxt.key0 [2]);
tran (gcm_dak_cmd_in_nxt[358], \gcm_dak_cmd_in_nxt.key0 [3]);
tran (gcm_dak_cmd_in_nxt[359], \gcm_dak_cmd_in_nxt.key0 [4]);
tran (gcm_dak_cmd_in_nxt[360], \gcm_dak_cmd_in_nxt.key0 [5]);
tran (gcm_dak_cmd_in_nxt[361], \gcm_dak_cmd_in_nxt.key0 [6]);
tran (gcm_dak_cmd_in_nxt[362], \gcm_dak_cmd_in_nxt.key0 [7]);
tran (gcm_dak_cmd_in_nxt[363], \gcm_dak_cmd_in_nxt.key0 [8]);
tran (gcm_dak_cmd_in_nxt[364], \gcm_dak_cmd_in_nxt.key0 [9]);
tran (gcm_dak_cmd_in_nxt[365], \gcm_dak_cmd_in_nxt.key0 [10]);
tran (gcm_dak_cmd_in_nxt[366], \gcm_dak_cmd_in_nxt.key0 [11]);
tran (gcm_dak_cmd_in_nxt[367], \gcm_dak_cmd_in_nxt.key0 [12]);
tran (gcm_dak_cmd_in_nxt[368], \gcm_dak_cmd_in_nxt.key0 [13]);
tran (gcm_dak_cmd_in_nxt[369], \gcm_dak_cmd_in_nxt.key0 [14]);
tran (gcm_dak_cmd_in_nxt[370], \gcm_dak_cmd_in_nxt.key0 [15]);
tran (gcm_dak_cmd_in_nxt[371], \gcm_dak_cmd_in_nxt.key0 [16]);
tran (gcm_dak_cmd_in_nxt[372], \gcm_dak_cmd_in_nxt.key0 [17]);
tran (gcm_dak_cmd_in_nxt[373], \gcm_dak_cmd_in_nxt.key0 [18]);
tran (gcm_dak_cmd_in_nxt[374], \gcm_dak_cmd_in_nxt.key0 [19]);
tran (gcm_dak_cmd_in_nxt[375], \gcm_dak_cmd_in_nxt.key0 [20]);
tran (gcm_dak_cmd_in_nxt[376], \gcm_dak_cmd_in_nxt.key0 [21]);
tran (gcm_dak_cmd_in_nxt[377], \gcm_dak_cmd_in_nxt.key0 [22]);
tran (gcm_dak_cmd_in_nxt[378], \gcm_dak_cmd_in_nxt.key0 [23]);
tran (gcm_dak_cmd_in_nxt[379], \gcm_dak_cmd_in_nxt.key0 [24]);
tran (gcm_dak_cmd_in_nxt[380], \gcm_dak_cmd_in_nxt.key0 [25]);
tran (gcm_dak_cmd_in_nxt[381], \gcm_dak_cmd_in_nxt.key0 [26]);
tran (gcm_dak_cmd_in_nxt[382], \gcm_dak_cmd_in_nxt.key0 [27]);
tran (gcm_dak_cmd_in_nxt[383], \gcm_dak_cmd_in_nxt.key0 [28]);
tran (gcm_dak_cmd_in_nxt[384], \gcm_dak_cmd_in_nxt.key0 [29]);
tran (gcm_dak_cmd_in_nxt[385], \gcm_dak_cmd_in_nxt.key0 [30]);
tran (gcm_dak_cmd_in_nxt[386], \gcm_dak_cmd_in_nxt.key0 [31]);
tran (gcm_dak_cmd_in_nxt[387], \gcm_dak_cmd_in_nxt.key0 [32]);
tran (gcm_dak_cmd_in_nxt[388], \gcm_dak_cmd_in_nxt.key0 [33]);
tran (gcm_dak_cmd_in_nxt[389], \gcm_dak_cmd_in_nxt.key0 [34]);
tran (gcm_dak_cmd_in_nxt[390], \gcm_dak_cmd_in_nxt.key0 [35]);
tran (gcm_dak_cmd_in_nxt[391], \gcm_dak_cmd_in_nxt.key0 [36]);
tran (gcm_dak_cmd_in_nxt[392], \gcm_dak_cmd_in_nxt.key0 [37]);
tran (gcm_dak_cmd_in_nxt[393], \gcm_dak_cmd_in_nxt.key0 [38]);
tran (gcm_dak_cmd_in_nxt[394], \gcm_dak_cmd_in_nxt.key0 [39]);
tran (gcm_dak_cmd_in_nxt[395], \gcm_dak_cmd_in_nxt.key0 [40]);
tran (gcm_dak_cmd_in_nxt[396], \gcm_dak_cmd_in_nxt.key0 [41]);
tran (gcm_dak_cmd_in_nxt[397], \gcm_dak_cmd_in_nxt.key0 [42]);
tran (gcm_dak_cmd_in_nxt[398], \gcm_dak_cmd_in_nxt.key0 [43]);
tran (gcm_dak_cmd_in_nxt[399], \gcm_dak_cmd_in_nxt.key0 [44]);
tran (gcm_dak_cmd_in_nxt[400], \gcm_dak_cmd_in_nxt.key0 [45]);
tran (gcm_dak_cmd_in_nxt[401], \gcm_dak_cmd_in_nxt.key0 [46]);
tran (gcm_dak_cmd_in_nxt[402], \gcm_dak_cmd_in_nxt.key0 [47]);
tran (gcm_dak_cmd_in_nxt[403], \gcm_dak_cmd_in_nxt.key0 [48]);
tran (gcm_dak_cmd_in_nxt[404], \gcm_dak_cmd_in_nxt.key0 [49]);
tran (gcm_dak_cmd_in_nxt[405], \gcm_dak_cmd_in_nxt.key0 [50]);
tran (gcm_dak_cmd_in_nxt[406], \gcm_dak_cmd_in_nxt.key0 [51]);
tran (gcm_dak_cmd_in_nxt[407], \gcm_dak_cmd_in_nxt.key0 [52]);
tran (gcm_dak_cmd_in_nxt[408], \gcm_dak_cmd_in_nxt.key0 [53]);
tran (gcm_dak_cmd_in_nxt[409], \gcm_dak_cmd_in_nxt.key0 [54]);
tran (gcm_dak_cmd_in_nxt[410], \gcm_dak_cmd_in_nxt.key0 [55]);
tran (gcm_dak_cmd_in_nxt[411], \gcm_dak_cmd_in_nxt.key0 [56]);
tran (gcm_dak_cmd_in_nxt[412], \gcm_dak_cmd_in_nxt.key0 [57]);
tran (gcm_dak_cmd_in_nxt[413], \gcm_dak_cmd_in_nxt.key0 [58]);
tran (gcm_dak_cmd_in_nxt[414], \gcm_dak_cmd_in_nxt.key0 [59]);
tran (gcm_dak_cmd_in_nxt[415], \gcm_dak_cmd_in_nxt.key0 [60]);
tran (gcm_dak_cmd_in_nxt[416], \gcm_dak_cmd_in_nxt.key0 [61]);
tran (gcm_dak_cmd_in_nxt[417], \gcm_dak_cmd_in_nxt.key0 [62]);
tran (gcm_dak_cmd_in_nxt[418], \gcm_dak_cmd_in_nxt.key0 [63]);
tran (gcm_dak_cmd_in_nxt[419], \gcm_dak_cmd_in_nxt.key0 [64]);
tran (gcm_dak_cmd_in_nxt[420], \gcm_dak_cmd_in_nxt.key0 [65]);
tran (gcm_dak_cmd_in_nxt[421], \gcm_dak_cmd_in_nxt.key0 [66]);
tran (gcm_dak_cmd_in_nxt[422], \gcm_dak_cmd_in_nxt.key0 [67]);
tran (gcm_dak_cmd_in_nxt[423], \gcm_dak_cmd_in_nxt.key0 [68]);
tran (gcm_dak_cmd_in_nxt[424], \gcm_dak_cmd_in_nxt.key0 [69]);
tran (gcm_dak_cmd_in_nxt[425], \gcm_dak_cmd_in_nxt.key0 [70]);
tran (gcm_dak_cmd_in_nxt[426], \gcm_dak_cmd_in_nxt.key0 [71]);
tran (gcm_dak_cmd_in_nxt[427], \gcm_dak_cmd_in_nxt.key0 [72]);
tran (gcm_dak_cmd_in_nxt[428], \gcm_dak_cmd_in_nxt.key0 [73]);
tran (gcm_dak_cmd_in_nxt[429], \gcm_dak_cmd_in_nxt.key0 [74]);
tran (gcm_dak_cmd_in_nxt[430], \gcm_dak_cmd_in_nxt.key0 [75]);
tran (gcm_dak_cmd_in_nxt[431], \gcm_dak_cmd_in_nxt.key0 [76]);
tran (gcm_dak_cmd_in_nxt[432], \gcm_dak_cmd_in_nxt.key0 [77]);
tran (gcm_dak_cmd_in_nxt[433], \gcm_dak_cmd_in_nxt.key0 [78]);
tran (gcm_dak_cmd_in_nxt[434], \gcm_dak_cmd_in_nxt.key0 [79]);
tran (gcm_dak_cmd_in_nxt[435], \gcm_dak_cmd_in_nxt.key0 [80]);
tran (gcm_dak_cmd_in_nxt[436], \gcm_dak_cmd_in_nxt.key0 [81]);
tran (gcm_dak_cmd_in_nxt[437], \gcm_dak_cmd_in_nxt.key0 [82]);
tran (gcm_dak_cmd_in_nxt[438], \gcm_dak_cmd_in_nxt.key0 [83]);
tran (gcm_dak_cmd_in_nxt[439], \gcm_dak_cmd_in_nxt.key0 [84]);
tran (gcm_dak_cmd_in_nxt[440], \gcm_dak_cmd_in_nxt.key0 [85]);
tran (gcm_dak_cmd_in_nxt[441], \gcm_dak_cmd_in_nxt.key0 [86]);
tran (gcm_dak_cmd_in_nxt[442], \gcm_dak_cmd_in_nxt.key0 [87]);
tran (gcm_dak_cmd_in_nxt[443], \gcm_dak_cmd_in_nxt.key0 [88]);
tran (gcm_dak_cmd_in_nxt[444], \gcm_dak_cmd_in_nxt.key0 [89]);
tran (gcm_dak_cmd_in_nxt[445], \gcm_dak_cmd_in_nxt.key0 [90]);
tran (gcm_dak_cmd_in_nxt[446], \gcm_dak_cmd_in_nxt.key0 [91]);
tran (gcm_dak_cmd_in_nxt[447], \gcm_dak_cmd_in_nxt.key0 [92]);
tran (gcm_dak_cmd_in_nxt[448], \gcm_dak_cmd_in_nxt.key0 [93]);
tran (gcm_dak_cmd_in_nxt[449], \gcm_dak_cmd_in_nxt.key0 [94]);
tran (gcm_dak_cmd_in_nxt[450], \gcm_dak_cmd_in_nxt.key0 [95]);
tran (gcm_dak_cmd_in_nxt[451], \gcm_dak_cmd_in_nxt.key0 [96]);
tran (gcm_dak_cmd_in_nxt[452], \gcm_dak_cmd_in_nxt.key0 [97]);
tran (gcm_dak_cmd_in_nxt[453], \gcm_dak_cmd_in_nxt.key0 [98]);
tran (gcm_dak_cmd_in_nxt[454], \gcm_dak_cmd_in_nxt.key0 [99]);
tran (gcm_dak_cmd_in_nxt[455], \gcm_dak_cmd_in_nxt.key0 [100]);
tran (gcm_dak_cmd_in_nxt[456], \gcm_dak_cmd_in_nxt.key0 [101]);
tran (gcm_dak_cmd_in_nxt[457], \gcm_dak_cmd_in_nxt.key0 [102]);
tran (gcm_dak_cmd_in_nxt[458], \gcm_dak_cmd_in_nxt.key0 [103]);
tran (gcm_dak_cmd_in_nxt[459], \gcm_dak_cmd_in_nxt.key0 [104]);
tran (gcm_dak_cmd_in_nxt[460], \gcm_dak_cmd_in_nxt.key0 [105]);
tran (gcm_dak_cmd_in_nxt[461], \gcm_dak_cmd_in_nxt.key0 [106]);
tran (gcm_dak_cmd_in_nxt[462], \gcm_dak_cmd_in_nxt.key0 [107]);
tran (gcm_dak_cmd_in_nxt[463], \gcm_dak_cmd_in_nxt.key0 [108]);
tran (gcm_dak_cmd_in_nxt[464], \gcm_dak_cmd_in_nxt.key0 [109]);
tran (gcm_dak_cmd_in_nxt[465], \gcm_dak_cmd_in_nxt.key0 [110]);
tran (gcm_dak_cmd_in_nxt[466], \gcm_dak_cmd_in_nxt.key0 [111]);
tran (gcm_dak_cmd_in_nxt[467], \gcm_dak_cmd_in_nxt.key0 [112]);
tran (gcm_dak_cmd_in_nxt[468], \gcm_dak_cmd_in_nxt.key0 [113]);
tran (gcm_dak_cmd_in_nxt[469], \gcm_dak_cmd_in_nxt.key0 [114]);
tran (gcm_dak_cmd_in_nxt[470], \gcm_dak_cmd_in_nxt.key0 [115]);
tran (gcm_dak_cmd_in_nxt[471], \gcm_dak_cmd_in_nxt.key0 [116]);
tran (gcm_dak_cmd_in_nxt[472], \gcm_dak_cmd_in_nxt.key0 [117]);
tran (gcm_dak_cmd_in_nxt[473], \gcm_dak_cmd_in_nxt.key0 [118]);
tran (gcm_dak_cmd_in_nxt[474], \gcm_dak_cmd_in_nxt.key0 [119]);
tran (gcm_dak_cmd_in_nxt[475], \gcm_dak_cmd_in_nxt.key0 [120]);
tran (gcm_dak_cmd_in_nxt[476], \gcm_dak_cmd_in_nxt.key0 [121]);
tran (gcm_dak_cmd_in_nxt[477], \gcm_dak_cmd_in_nxt.key0 [122]);
tran (gcm_dak_cmd_in_nxt[478], \gcm_dak_cmd_in_nxt.key0 [123]);
tran (gcm_dak_cmd_in_nxt[479], \gcm_dak_cmd_in_nxt.key0 [124]);
tran (gcm_dak_cmd_in_nxt[480], \gcm_dak_cmd_in_nxt.key0 [125]);
tran (gcm_dak_cmd_in_nxt[481], \gcm_dak_cmd_in_nxt.key0 [126]);
tran (gcm_dak_cmd_in_nxt[482], \gcm_dak_cmd_in_nxt.key0 [127]);
tran (gcm_dak_cmd_in_nxt[483], \gcm_dak_cmd_in_nxt.key0 [128]);
tran (gcm_dak_cmd_in_nxt[484], \gcm_dak_cmd_in_nxt.key0 [129]);
tran (gcm_dak_cmd_in_nxt[485], \gcm_dak_cmd_in_nxt.key0 [130]);
tran (gcm_dak_cmd_in_nxt[486], \gcm_dak_cmd_in_nxt.key0 [131]);
tran (gcm_dak_cmd_in_nxt[487], \gcm_dak_cmd_in_nxt.key0 [132]);
tran (gcm_dak_cmd_in_nxt[488], \gcm_dak_cmd_in_nxt.key0 [133]);
tran (gcm_dak_cmd_in_nxt[489], \gcm_dak_cmd_in_nxt.key0 [134]);
tran (gcm_dak_cmd_in_nxt[490], \gcm_dak_cmd_in_nxt.key0 [135]);
tran (gcm_dak_cmd_in_nxt[491], \gcm_dak_cmd_in_nxt.key0 [136]);
tran (gcm_dak_cmd_in_nxt[492], \gcm_dak_cmd_in_nxt.key0 [137]);
tran (gcm_dak_cmd_in_nxt[493], \gcm_dak_cmd_in_nxt.key0 [138]);
tran (gcm_dak_cmd_in_nxt[494], \gcm_dak_cmd_in_nxt.key0 [139]);
tran (gcm_dak_cmd_in_nxt[495], \gcm_dak_cmd_in_nxt.key0 [140]);
tran (gcm_dak_cmd_in_nxt[496], \gcm_dak_cmd_in_nxt.key0 [141]);
tran (gcm_dak_cmd_in_nxt[497], \gcm_dak_cmd_in_nxt.key0 [142]);
tran (gcm_dak_cmd_in_nxt[498], \gcm_dak_cmd_in_nxt.key0 [143]);
tran (gcm_dak_cmd_in_nxt[499], \gcm_dak_cmd_in_nxt.key0 [144]);
tran (gcm_dak_cmd_in_nxt[500], \gcm_dak_cmd_in_nxt.key0 [145]);
tran (gcm_dak_cmd_in_nxt[501], \gcm_dak_cmd_in_nxt.key0 [146]);
tran (gcm_dak_cmd_in_nxt[502], \gcm_dak_cmd_in_nxt.key0 [147]);
tran (gcm_dak_cmd_in_nxt[503], \gcm_dak_cmd_in_nxt.key0 [148]);
tran (gcm_dak_cmd_in_nxt[504], \gcm_dak_cmd_in_nxt.key0 [149]);
tran (gcm_dak_cmd_in_nxt[505], \gcm_dak_cmd_in_nxt.key0 [150]);
tran (gcm_dak_cmd_in_nxt[506], \gcm_dak_cmd_in_nxt.key0 [151]);
tran (gcm_dak_cmd_in_nxt[507], \gcm_dak_cmd_in_nxt.key0 [152]);
tran (gcm_dak_cmd_in_nxt[508], \gcm_dak_cmd_in_nxt.key0 [153]);
tran (gcm_dak_cmd_in_nxt[509], \gcm_dak_cmd_in_nxt.key0 [154]);
tran (gcm_dak_cmd_in_nxt[510], \gcm_dak_cmd_in_nxt.key0 [155]);
tran (gcm_dak_cmd_in_nxt[511], \gcm_dak_cmd_in_nxt.key0 [156]);
tran (gcm_dak_cmd_in_nxt[512], \gcm_dak_cmd_in_nxt.key0 [157]);
tran (gcm_dak_cmd_in_nxt[513], \gcm_dak_cmd_in_nxt.key0 [158]);
tran (gcm_dak_cmd_in_nxt[514], \gcm_dak_cmd_in_nxt.key0 [159]);
tran (gcm_dak_cmd_in_nxt[515], \gcm_dak_cmd_in_nxt.key0 [160]);
tran (gcm_dak_cmd_in_nxt[516], \gcm_dak_cmd_in_nxt.key0 [161]);
tran (gcm_dak_cmd_in_nxt[517], \gcm_dak_cmd_in_nxt.key0 [162]);
tran (gcm_dak_cmd_in_nxt[518], \gcm_dak_cmd_in_nxt.key0 [163]);
tran (gcm_dak_cmd_in_nxt[519], \gcm_dak_cmd_in_nxt.key0 [164]);
tran (gcm_dak_cmd_in_nxt[520], \gcm_dak_cmd_in_nxt.key0 [165]);
tran (gcm_dak_cmd_in_nxt[521], \gcm_dak_cmd_in_nxt.key0 [166]);
tran (gcm_dak_cmd_in_nxt[522], \gcm_dak_cmd_in_nxt.key0 [167]);
tran (gcm_dak_cmd_in_nxt[523], \gcm_dak_cmd_in_nxt.key0 [168]);
tran (gcm_dak_cmd_in_nxt[524], \gcm_dak_cmd_in_nxt.key0 [169]);
tran (gcm_dak_cmd_in_nxt[525], \gcm_dak_cmd_in_nxt.key0 [170]);
tran (gcm_dak_cmd_in_nxt[526], \gcm_dak_cmd_in_nxt.key0 [171]);
tran (gcm_dak_cmd_in_nxt[527], \gcm_dak_cmd_in_nxt.key0 [172]);
tran (gcm_dak_cmd_in_nxt[528], \gcm_dak_cmd_in_nxt.key0 [173]);
tran (gcm_dak_cmd_in_nxt[529], \gcm_dak_cmd_in_nxt.key0 [174]);
tran (gcm_dak_cmd_in_nxt[530], \gcm_dak_cmd_in_nxt.key0 [175]);
tran (gcm_dak_cmd_in_nxt[531], \gcm_dak_cmd_in_nxt.key0 [176]);
tran (gcm_dak_cmd_in_nxt[532], \gcm_dak_cmd_in_nxt.key0 [177]);
tran (gcm_dak_cmd_in_nxt[533], \gcm_dak_cmd_in_nxt.key0 [178]);
tran (gcm_dak_cmd_in_nxt[534], \gcm_dak_cmd_in_nxt.key0 [179]);
tran (gcm_dak_cmd_in_nxt[535], \gcm_dak_cmd_in_nxt.key0 [180]);
tran (gcm_dak_cmd_in_nxt[536], \gcm_dak_cmd_in_nxt.key0 [181]);
tran (gcm_dak_cmd_in_nxt[537], \gcm_dak_cmd_in_nxt.key0 [182]);
tran (gcm_dak_cmd_in_nxt[538], \gcm_dak_cmd_in_nxt.key0 [183]);
tran (gcm_dak_cmd_in_nxt[539], \gcm_dak_cmd_in_nxt.key0 [184]);
tran (gcm_dak_cmd_in_nxt[540], \gcm_dak_cmd_in_nxt.key0 [185]);
tran (gcm_dak_cmd_in_nxt[541], \gcm_dak_cmd_in_nxt.key0 [186]);
tran (gcm_dak_cmd_in_nxt[542], \gcm_dak_cmd_in_nxt.key0 [187]);
tran (gcm_dak_cmd_in_nxt[543], \gcm_dak_cmd_in_nxt.key0 [188]);
tran (gcm_dak_cmd_in_nxt[544], \gcm_dak_cmd_in_nxt.key0 [189]);
tran (gcm_dak_cmd_in_nxt[545], \gcm_dak_cmd_in_nxt.key0 [190]);
tran (gcm_dak_cmd_in_nxt[546], \gcm_dak_cmd_in_nxt.key0 [191]);
tran (gcm_dak_cmd_in_nxt[547], \gcm_dak_cmd_in_nxt.key0 [192]);
tran (gcm_dak_cmd_in_nxt[548], \gcm_dak_cmd_in_nxt.key0 [193]);
tran (gcm_dak_cmd_in_nxt[549], \gcm_dak_cmd_in_nxt.key0 [194]);
tran (gcm_dak_cmd_in_nxt[550], \gcm_dak_cmd_in_nxt.key0 [195]);
tran (gcm_dak_cmd_in_nxt[551], \gcm_dak_cmd_in_nxt.key0 [196]);
tran (gcm_dak_cmd_in_nxt[552], \gcm_dak_cmd_in_nxt.key0 [197]);
tran (gcm_dak_cmd_in_nxt[553], \gcm_dak_cmd_in_nxt.key0 [198]);
tran (gcm_dak_cmd_in_nxt[554], \gcm_dak_cmd_in_nxt.key0 [199]);
tran (gcm_dak_cmd_in_nxt[555], \gcm_dak_cmd_in_nxt.key0 [200]);
tran (gcm_dak_cmd_in_nxt[556], \gcm_dak_cmd_in_nxt.key0 [201]);
tran (gcm_dak_cmd_in_nxt[557], \gcm_dak_cmd_in_nxt.key0 [202]);
tran (gcm_dak_cmd_in_nxt[558], \gcm_dak_cmd_in_nxt.key0 [203]);
tran (gcm_dak_cmd_in_nxt[559], \gcm_dak_cmd_in_nxt.key0 [204]);
tran (gcm_dak_cmd_in_nxt[560], \gcm_dak_cmd_in_nxt.key0 [205]);
tran (gcm_dak_cmd_in_nxt[561], \gcm_dak_cmd_in_nxt.key0 [206]);
tran (gcm_dak_cmd_in_nxt[562], \gcm_dak_cmd_in_nxt.key0 [207]);
tran (gcm_dak_cmd_in_nxt[563], \gcm_dak_cmd_in_nxt.key0 [208]);
tran (gcm_dak_cmd_in_nxt[564], \gcm_dak_cmd_in_nxt.key0 [209]);
tran (gcm_dak_cmd_in_nxt[565], \gcm_dak_cmd_in_nxt.key0 [210]);
tran (gcm_dak_cmd_in_nxt[566], \gcm_dak_cmd_in_nxt.key0 [211]);
tran (gcm_dak_cmd_in_nxt[567], \gcm_dak_cmd_in_nxt.key0 [212]);
tran (gcm_dak_cmd_in_nxt[568], \gcm_dak_cmd_in_nxt.key0 [213]);
tran (gcm_dak_cmd_in_nxt[569], \gcm_dak_cmd_in_nxt.key0 [214]);
tran (gcm_dak_cmd_in_nxt[570], \gcm_dak_cmd_in_nxt.key0 [215]);
tran (gcm_dak_cmd_in_nxt[571], \gcm_dak_cmd_in_nxt.key0 [216]);
tran (gcm_dak_cmd_in_nxt[572], \gcm_dak_cmd_in_nxt.key0 [217]);
tran (gcm_dak_cmd_in_nxt[573], \gcm_dak_cmd_in_nxt.key0 [218]);
tran (gcm_dak_cmd_in_nxt[574], \gcm_dak_cmd_in_nxt.key0 [219]);
tran (gcm_dak_cmd_in_nxt[575], \gcm_dak_cmd_in_nxt.key0 [220]);
tran (gcm_dak_cmd_in_nxt[576], \gcm_dak_cmd_in_nxt.key0 [221]);
tran (gcm_dak_cmd_in_nxt[577], \gcm_dak_cmd_in_nxt.key0 [222]);
tran (gcm_dak_cmd_in_nxt[578], \gcm_dak_cmd_in_nxt.key0 [223]);
tran (gcm_dak_cmd_in_nxt[579], \gcm_dak_cmd_in_nxt.key0 [224]);
tran (gcm_dak_cmd_in_nxt[580], \gcm_dak_cmd_in_nxt.key0 [225]);
tran (gcm_dak_cmd_in_nxt[581], \gcm_dak_cmd_in_nxt.key0 [226]);
tran (gcm_dak_cmd_in_nxt[582], \gcm_dak_cmd_in_nxt.key0 [227]);
tran (gcm_dak_cmd_in_nxt[583], \gcm_dak_cmd_in_nxt.key0 [228]);
tran (gcm_dak_cmd_in_nxt[584], \gcm_dak_cmd_in_nxt.key0 [229]);
tran (gcm_dak_cmd_in_nxt[585], \gcm_dak_cmd_in_nxt.key0 [230]);
tran (gcm_dak_cmd_in_nxt[586], \gcm_dak_cmd_in_nxt.key0 [231]);
tran (gcm_dak_cmd_in_nxt[587], \gcm_dak_cmd_in_nxt.key0 [232]);
tran (gcm_dak_cmd_in_nxt[588], \gcm_dak_cmd_in_nxt.key0 [233]);
tran (gcm_dak_cmd_in_nxt[589], \gcm_dak_cmd_in_nxt.key0 [234]);
tran (gcm_dak_cmd_in_nxt[590], \gcm_dak_cmd_in_nxt.key0 [235]);
tran (gcm_dak_cmd_in_nxt[591], \gcm_dak_cmd_in_nxt.key0 [236]);
tran (gcm_dak_cmd_in_nxt[592], \gcm_dak_cmd_in_nxt.key0 [237]);
tran (gcm_dak_cmd_in_nxt[593], \gcm_dak_cmd_in_nxt.key0 [238]);
tran (gcm_dak_cmd_in_nxt[594], \gcm_dak_cmd_in_nxt.key0 [239]);
tran (gcm_dak_cmd_in_nxt[595], \gcm_dak_cmd_in_nxt.key0 [240]);
tran (gcm_dak_cmd_in_nxt[596], \gcm_dak_cmd_in_nxt.key0 [241]);
tran (gcm_dak_cmd_in_nxt[597], \gcm_dak_cmd_in_nxt.key0 [242]);
tran (gcm_dak_cmd_in_nxt[598], \gcm_dak_cmd_in_nxt.key0 [243]);
tran (gcm_dak_cmd_in_nxt[599], \gcm_dak_cmd_in_nxt.key0 [244]);
tran (gcm_dak_cmd_in_nxt[600], \gcm_dak_cmd_in_nxt.key0 [245]);
tran (gcm_dak_cmd_in_nxt[601], \gcm_dak_cmd_in_nxt.key0 [246]);
tran (gcm_dak_cmd_in_nxt[602], \gcm_dak_cmd_in_nxt.key0 [247]);
tran (gcm_dak_cmd_in_nxt[603], \gcm_dak_cmd_in_nxt.key0 [248]);
tran (gcm_dak_cmd_in_nxt[604], \gcm_dak_cmd_in_nxt.key0 [249]);
tran (gcm_dak_cmd_in_nxt[605], \gcm_dak_cmd_in_nxt.key0 [250]);
tran (gcm_dak_cmd_in_nxt[606], \gcm_dak_cmd_in_nxt.key0 [251]);
tran (gcm_dak_cmd_in_nxt[607], \gcm_dak_cmd_in_nxt.key0 [252]);
tran (gcm_dak_cmd_in_nxt[608], \gcm_dak_cmd_in_nxt.key0 [253]);
tran (gcm_dak_cmd_in_nxt[609], \gcm_dak_cmd_in_nxt.key0 [254]);
tran (gcm_dak_cmd_in_nxt[610], \gcm_dak_cmd_in_nxt.key0 [255]);
tran (gcm_dek_cmd_in_nxt[0], \gcm_dek_cmd_in_nxt.op [0]);
tran (gcm_dek_cmd_in_nxt[1], \gcm_dek_cmd_in_nxt.op [1]);
tran (gcm_dek_cmd_in_nxt[2], \gcm_dek_cmd_in_nxt.op [2]);
tran (gcm_dek_cmd_in_nxt[3], \gcm_dek_cmd_in_nxt.iv [0]);
tran (gcm_dek_cmd_in_nxt[4], \gcm_dek_cmd_in_nxt.iv [1]);
tran (gcm_dek_cmd_in_nxt[5], \gcm_dek_cmd_in_nxt.iv [2]);
tran (gcm_dek_cmd_in_nxt[6], \gcm_dek_cmd_in_nxt.iv [3]);
tran (gcm_dek_cmd_in_nxt[7], \gcm_dek_cmd_in_nxt.iv [4]);
tran (gcm_dek_cmd_in_nxt[8], \gcm_dek_cmd_in_nxt.iv [5]);
tran (gcm_dek_cmd_in_nxt[9], \gcm_dek_cmd_in_nxt.iv [6]);
tran (gcm_dek_cmd_in_nxt[10], \gcm_dek_cmd_in_nxt.iv [7]);
tran (gcm_dek_cmd_in_nxt[11], \gcm_dek_cmd_in_nxt.iv [8]);
tran (gcm_dek_cmd_in_nxt[12], \gcm_dek_cmd_in_nxt.iv [9]);
tran (gcm_dek_cmd_in_nxt[13], \gcm_dek_cmd_in_nxt.iv [10]);
tran (gcm_dek_cmd_in_nxt[14], \gcm_dek_cmd_in_nxt.iv [11]);
tran (gcm_dek_cmd_in_nxt[15], \gcm_dek_cmd_in_nxt.iv [12]);
tran (gcm_dek_cmd_in_nxt[16], \gcm_dek_cmd_in_nxt.iv [13]);
tran (gcm_dek_cmd_in_nxt[17], \gcm_dek_cmd_in_nxt.iv [14]);
tran (gcm_dek_cmd_in_nxt[18], \gcm_dek_cmd_in_nxt.iv [15]);
tran (gcm_dek_cmd_in_nxt[19], \gcm_dek_cmd_in_nxt.iv [16]);
tran (gcm_dek_cmd_in_nxt[20], \gcm_dek_cmd_in_nxt.iv [17]);
tran (gcm_dek_cmd_in_nxt[21], \gcm_dek_cmd_in_nxt.iv [18]);
tran (gcm_dek_cmd_in_nxt[22], \gcm_dek_cmd_in_nxt.iv [19]);
tran (gcm_dek_cmd_in_nxt[23], \gcm_dek_cmd_in_nxt.iv [20]);
tran (gcm_dek_cmd_in_nxt[24], \gcm_dek_cmd_in_nxt.iv [21]);
tran (gcm_dek_cmd_in_nxt[25], \gcm_dek_cmd_in_nxt.iv [22]);
tran (gcm_dek_cmd_in_nxt[26], \gcm_dek_cmd_in_nxt.iv [23]);
tran (gcm_dek_cmd_in_nxt[27], \gcm_dek_cmd_in_nxt.iv [24]);
tran (gcm_dek_cmd_in_nxt[28], \gcm_dek_cmd_in_nxt.iv [25]);
tran (gcm_dek_cmd_in_nxt[29], \gcm_dek_cmd_in_nxt.iv [26]);
tran (gcm_dek_cmd_in_nxt[30], \gcm_dek_cmd_in_nxt.iv [27]);
tran (gcm_dek_cmd_in_nxt[31], \gcm_dek_cmd_in_nxt.iv [28]);
tran (gcm_dek_cmd_in_nxt[32], \gcm_dek_cmd_in_nxt.iv [29]);
tran (gcm_dek_cmd_in_nxt[33], \gcm_dek_cmd_in_nxt.iv [30]);
tran (gcm_dek_cmd_in_nxt[34], \gcm_dek_cmd_in_nxt.iv [31]);
tran (gcm_dek_cmd_in_nxt[35], \gcm_dek_cmd_in_nxt.iv [32]);
tran (gcm_dek_cmd_in_nxt[36], \gcm_dek_cmd_in_nxt.iv [33]);
tran (gcm_dek_cmd_in_nxt[37], \gcm_dek_cmd_in_nxt.iv [34]);
tran (gcm_dek_cmd_in_nxt[38], \gcm_dek_cmd_in_nxt.iv [35]);
tran (gcm_dek_cmd_in_nxt[39], \gcm_dek_cmd_in_nxt.iv [36]);
tran (gcm_dek_cmd_in_nxt[40], \gcm_dek_cmd_in_nxt.iv [37]);
tran (gcm_dek_cmd_in_nxt[41], \gcm_dek_cmd_in_nxt.iv [38]);
tran (gcm_dek_cmd_in_nxt[42], \gcm_dek_cmd_in_nxt.iv [39]);
tran (gcm_dek_cmd_in_nxt[43], \gcm_dek_cmd_in_nxt.iv [40]);
tran (gcm_dek_cmd_in_nxt[44], \gcm_dek_cmd_in_nxt.iv [41]);
tran (gcm_dek_cmd_in_nxt[45], \gcm_dek_cmd_in_nxt.iv [42]);
tran (gcm_dek_cmd_in_nxt[46], \gcm_dek_cmd_in_nxt.iv [43]);
tran (gcm_dek_cmd_in_nxt[47], \gcm_dek_cmd_in_nxt.iv [44]);
tran (gcm_dek_cmd_in_nxt[48], \gcm_dek_cmd_in_nxt.iv [45]);
tran (gcm_dek_cmd_in_nxt[49], \gcm_dek_cmd_in_nxt.iv [46]);
tran (gcm_dek_cmd_in_nxt[50], \gcm_dek_cmd_in_nxt.iv [47]);
tran (gcm_dek_cmd_in_nxt[51], \gcm_dek_cmd_in_nxt.iv [48]);
tran (gcm_dek_cmd_in_nxt[52], \gcm_dek_cmd_in_nxt.iv [49]);
tran (gcm_dek_cmd_in_nxt[53], \gcm_dek_cmd_in_nxt.iv [50]);
tran (gcm_dek_cmd_in_nxt[54], \gcm_dek_cmd_in_nxt.iv [51]);
tran (gcm_dek_cmd_in_nxt[55], \gcm_dek_cmd_in_nxt.iv [52]);
tran (gcm_dek_cmd_in_nxt[56], \gcm_dek_cmd_in_nxt.iv [53]);
tran (gcm_dek_cmd_in_nxt[57], \gcm_dek_cmd_in_nxt.iv [54]);
tran (gcm_dek_cmd_in_nxt[58], \gcm_dek_cmd_in_nxt.iv [55]);
tran (gcm_dek_cmd_in_nxt[59], \gcm_dek_cmd_in_nxt.iv [56]);
tran (gcm_dek_cmd_in_nxt[60], \gcm_dek_cmd_in_nxt.iv [57]);
tran (gcm_dek_cmd_in_nxt[61], \gcm_dek_cmd_in_nxt.iv [58]);
tran (gcm_dek_cmd_in_nxt[62], \gcm_dek_cmd_in_nxt.iv [59]);
tran (gcm_dek_cmd_in_nxt[63], \gcm_dek_cmd_in_nxt.iv [60]);
tran (gcm_dek_cmd_in_nxt[64], \gcm_dek_cmd_in_nxt.iv [61]);
tran (gcm_dek_cmd_in_nxt[65], \gcm_dek_cmd_in_nxt.iv [62]);
tran (gcm_dek_cmd_in_nxt[66], \gcm_dek_cmd_in_nxt.iv [63]);
tran (gcm_dek_cmd_in_nxt[67], \gcm_dek_cmd_in_nxt.iv [64]);
tran (gcm_dek_cmd_in_nxt[68], \gcm_dek_cmd_in_nxt.iv [65]);
tran (gcm_dek_cmd_in_nxt[69], \gcm_dek_cmd_in_nxt.iv [66]);
tran (gcm_dek_cmd_in_nxt[70], \gcm_dek_cmd_in_nxt.iv [67]);
tran (gcm_dek_cmd_in_nxt[71], \gcm_dek_cmd_in_nxt.iv [68]);
tran (gcm_dek_cmd_in_nxt[72], \gcm_dek_cmd_in_nxt.iv [69]);
tran (gcm_dek_cmd_in_nxt[73], \gcm_dek_cmd_in_nxt.iv [70]);
tran (gcm_dek_cmd_in_nxt[74], \gcm_dek_cmd_in_nxt.iv [71]);
tran (gcm_dek_cmd_in_nxt[75], \gcm_dek_cmd_in_nxt.iv [72]);
tran (gcm_dek_cmd_in_nxt[76], \gcm_dek_cmd_in_nxt.iv [73]);
tran (gcm_dek_cmd_in_nxt[77], \gcm_dek_cmd_in_nxt.iv [74]);
tran (gcm_dek_cmd_in_nxt[78], \gcm_dek_cmd_in_nxt.iv [75]);
tran (gcm_dek_cmd_in_nxt[79], \gcm_dek_cmd_in_nxt.iv [76]);
tran (gcm_dek_cmd_in_nxt[80], \gcm_dek_cmd_in_nxt.iv [77]);
tran (gcm_dek_cmd_in_nxt[81], \gcm_dek_cmd_in_nxt.iv [78]);
tran (gcm_dek_cmd_in_nxt[82], \gcm_dek_cmd_in_nxt.iv [79]);
tran (gcm_dek_cmd_in_nxt[83], \gcm_dek_cmd_in_nxt.iv [80]);
tran (gcm_dek_cmd_in_nxt[84], \gcm_dek_cmd_in_nxt.iv [81]);
tran (gcm_dek_cmd_in_nxt[85], \gcm_dek_cmd_in_nxt.iv [82]);
tran (gcm_dek_cmd_in_nxt[86], \gcm_dek_cmd_in_nxt.iv [83]);
tran (gcm_dek_cmd_in_nxt[87], \gcm_dek_cmd_in_nxt.iv [84]);
tran (gcm_dek_cmd_in_nxt[88], \gcm_dek_cmd_in_nxt.iv [85]);
tran (gcm_dek_cmd_in_nxt[89], \gcm_dek_cmd_in_nxt.iv [86]);
tran (gcm_dek_cmd_in_nxt[90], \gcm_dek_cmd_in_nxt.iv [87]);
tran (gcm_dek_cmd_in_nxt[91], \gcm_dek_cmd_in_nxt.iv [88]);
tran (gcm_dek_cmd_in_nxt[92], \gcm_dek_cmd_in_nxt.iv [89]);
tran (gcm_dek_cmd_in_nxt[93], \gcm_dek_cmd_in_nxt.iv [90]);
tran (gcm_dek_cmd_in_nxt[94], \gcm_dek_cmd_in_nxt.iv [91]);
tran (gcm_dek_cmd_in_nxt[95], \gcm_dek_cmd_in_nxt.iv [92]);
tran (gcm_dek_cmd_in_nxt[96], \gcm_dek_cmd_in_nxt.iv [93]);
tran (gcm_dek_cmd_in_nxt[97], \gcm_dek_cmd_in_nxt.iv [94]);
tran (gcm_dek_cmd_in_nxt[98], \gcm_dek_cmd_in_nxt.iv [95]);
tran (gcm_dek_cmd_in_nxt[99], \gcm_dek_cmd_in_nxt.key1 [0]);
tran (gcm_dek_cmd_in_nxt[100], \gcm_dek_cmd_in_nxt.key1 [1]);
tran (gcm_dek_cmd_in_nxt[101], \gcm_dek_cmd_in_nxt.key1 [2]);
tran (gcm_dek_cmd_in_nxt[102], \gcm_dek_cmd_in_nxt.key1 [3]);
tran (gcm_dek_cmd_in_nxt[103], \gcm_dek_cmd_in_nxt.key1 [4]);
tran (gcm_dek_cmd_in_nxt[104], \gcm_dek_cmd_in_nxt.key1 [5]);
tran (gcm_dek_cmd_in_nxt[105], \gcm_dek_cmd_in_nxt.key1 [6]);
tran (gcm_dek_cmd_in_nxt[106], \gcm_dek_cmd_in_nxt.key1 [7]);
tran (gcm_dek_cmd_in_nxt[107], \gcm_dek_cmd_in_nxt.key1 [8]);
tran (gcm_dek_cmd_in_nxt[108], \gcm_dek_cmd_in_nxt.key1 [9]);
tran (gcm_dek_cmd_in_nxt[109], \gcm_dek_cmd_in_nxt.key1 [10]);
tran (gcm_dek_cmd_in_nxt[110], \gcm_dek_cmd_in_nxt.key1 [11]);
tran (gcm_dek_cmd_in_nxt[111], \gcm_dek_cmd_in_nxt.key1 [12]);
tran (gcm_dek_cmd_in_nxt[112], \gcm_dek_cmd_in_nxt.key1 [13]);
tran (gcm_dek_cmd_in_nxt[113], \gcm_dek_cmd_in_nxt.key1 [14]);
tran (gcm_dek_cmd_in_nxt[114], \gcm_dek_cmd_in_nxt.key1 [15]);
tran (gcm_dek_cmd_in_nxt[115], \gcm_dek_cmd_in_nxt.key1 [16]);
tran (gcm_dek_cmd_in_nxt[116], \gcm_dek_cmd_in_nxt.key1 [17]);
tran (gcm_dek_cmd_in_nxt[117], \gcm_dek_cmd_in_nxt.key1 [18]);
tran (gcm_dek_cmd_in_nxt[118], \gcm_dek_cmd_in_nxt.key1 [19]);
tran (gcm_dek_cmd_in_nxt[119], \gcm_dek_cmd_in_nxt.key1 [20]);
tran (gcm_dek_cmd_in_nxt[120], \gcm_dek_cmd_in_nxt.key1 [21]);
tran (gcm_dek_cmd_in_nxt[121], \gcm_dek_cmd_in_nxt.key1 [22]);
tran (gcm_dek_cmd_in_nxt[122], \gcm_dek_cmd_in_nxt.key1 [23]);
tran (gcm_dek_cmd_in_nxt[123], \gcm_dek_cmd_in_nxt.key1 [24]);
tran (gcm_dek_cmd_in_nxt[124], \gcm_dek_cmd_in_nxt.key1 [25]);
tran (gcm_dek_cmd_in_nxt[125], \gcm_dek_cmd_in_nxt.key1 [26]);
tran (gcm_dek_cmd_in_nxt[126], \gcm_dek_cmd_in_nxt.key1 [27]);
tran (gcm_dek_cmd_in_nxt[127], \gcm_dek_cmd_in_nxt.key1 [28]);
tran (gcm_dek_cmd_in_nxt[128], \gcm_dek_cmd_in_nxt.key1 [29]);
tran (gcm_dek_cmd_in_nxt[129], \gcm_dek_cmd_in_nxt.key1 [30]);
tran (gcm_dek_cmd_in_nxt[130], \gcm_dek_cmd_in_nxt.key1 [31]);
tran (gcm_dek_cmd_in_nxt[131], \gcm_dek_cmd_in_nxt.key1 [32]);
tran (gcm_dek_cmd_in_nxt[132], \gcm_dek_cmd_in_nxt.key1 [33]);
tran (gcm_dek_cmd_in_nxt[133], \gcm_dek_cmd_in_nxt.key1 [34]);
tran (gcm_dek_cmd_in_nxt[134], \gcm_dek_cmd_in_nxt.key1 [35]);
tran (gcm_dek_cmd_in_nxt[135], \gcm_dek_cmd_in_nxt.key1 [36]);
tran (gcm_dek_cmd_in_nxt[136], \gcm_dek_cmd_in_nxt.key1 [37]);
tran (gcm_dek_cmd_in_nxt[137], \gcm_dek_cmd_in_nxt.key1 [38]);
tran (gcm_dek_cmd_in_nxt[138], \gcm_dek_cmd_in_nxt.key1 [39]);
tran (gcm_dek_cmd_in_nxt[139], \gcm_dek_cmd_in_nxt.key1 [40]);
tran (gcm_dek_cmd_in_nxt[140], \gcm_dek_cmd_in_nxt.key1 [41]);
tran (gcm_dek_cmd_in_nxt[141], \gcm_dek_cmd_in_nxt.key1 [42]);
tran (gcm_dek_cmd_in_nxt[142], \gcm_dek_cmd_in_nxt.key1 [43]);
tran (gcm_dek_cmd_in_nxt[143], \gcm_dek_cmd_in_nxt.key1 [44]);
tran (gcm_dek_cmd_in_nxt[144], \gcm_dek_cmd_in_nxt.key1 [45]);
tran (gcm_dek_cmd_in_nxt[145], \gcm_dek_cmd_in_nxt.key1 [46]);
tran (gcm_dek_cmd_in_nxt[146], \gcm_dek_cmd_in_nxt.key1 [47]);
tran (gcm_dek_cmd_in_nxt[147], \gcm_dek_cmd_in_nxt.key1 [48]);
tran (gcm_dek_cmd_in_nxt[148], \gcm_dek_cmd_in_nxt.key1 [49]);
tran (gcm_dek_cmd_in_nxt[149], \gcm_dek_cmd_in_nxt.key1 [50]);
tran (gcm_dek_cmd_in_nxt[150], \gcm_dek_cmd_in_nxt.key1 [51]);
tran (gcm_dek_cmd_in_nxt[151], \gcm_dek_cmd_in_nxt.key1 [52]);
tran (gcm_dek_cmd_in_nxt[152], \gcm_dek_cmd_in_nxt.key1 [53]);
tran (gcm_dek_cmd_in_nxt[153], \gcm_dek_cmd_in_nxt.key1 [54]);
tran (gcm_dek_cmd_in_nxt[154], \gcm_dek_cmd_in_nxt.key1 [55]);
tran (gcm_dek_cmd_in_nxt[155], \gcm_dek_cmd_in_nxt.key1 [56]);
tran (gcm_dek_cmd_in_nxt[156], \gcm_dek_cmd_in_nxt.key1 [57]);
tran (gcm_dek_cmd_in_nxt[157], \gcm_dek_cmd_in_nxt.key1 [58]);
tran (gcm_dek_cmd_in_nxt[158], \gcm_dek_cmd_in_nxt.key1 [59]);
tran (gcm_dek_cmd_in_nxt[159], \gcm_dek_cmd_in_nxt.key1 [60]);
tran (gcm_dek_cmd_in_nxt[160], \gcm_dek_cmd_in_nxt.key1 [61]);
tran (gcm_dek_cmd_in_nxt[161], \gcm_dek_cmd_in_nxt.key1 [62]);
tran (gcm_dek_cmd_in_nxt[162], \gcm_dek_cmd_in_nxt.key1 [63]);
tran (gcm_dek_cmd_in_nxt[163], \gcm_dek_cmd_in_nxt.key1 [64]);
tran (gcm_dek_cmd_in_nxt[164], \gcm_dek_cmd_in_nxt.key1 [65]);
tran (gcm_dek_cmd_in_nxt[165], \gcm_dek_cmd_in_nxt.key1 [66]);
tran (gcm_dek_cmd_in_nxt[166], \gcm_dek_cmd_in_nxt.key1 [67]);
tran (gcm_dek_cmd_in_nxt[167], \gcm_dek_cmd_in_nxt.key1 [68]);
tran (gcm_dek_cmd_in_nxt[168], \gcm_dek_cmd_in_nxt.key1 [69]);
tran (gcm_dek_cmd_in_nxt[169], \gcm_dek_cmd_in_nxt.key1 [70]);
tran (gcm_dek_cmd_in_nxt[170], \gcm_dek_cmd_in_nxt.key1 [71]);
tran (gcm_dek_cmd_in_nxt[171], \gcm_dek_cmd_in_nxt.key1 [72]);
tran (gcm_dek_cmd_in_nxt[172], \gcm_dek_cmd_in_nxt.key1 [73]);
tran (gcm_dek_cmd_in_nxt[173], \gcm_dek_cmd_in_nxt.key1 [74]);
tran (gcm_dek_cmd_in_nxt[174], \gcm_dek_cmd_in_nxt.key1 [75]);
tran (gcm_dek_cmd_in_nxt[175], \gcm_dek_cmd_in_nxt.key1 [76]);
tran (gcm_dek_cmd_in_nxt[176], \gcm_dek_cmd_in_nxt.key1 [77]);
tran (gcm_dek_cmd_in_nxt[177], \gcm_dek_cmd_in_nxt.key1 [78]);
tran (gcm_dek_cmd_in_nxt[178], \gcm_dek_cmd_in_nxt.key1 [79]);
tran (gcm_dek_cmd_in_nxt[179], \gcm_dek_cmd_in_nxt.key1 [80]);
tran (gcm_dek_cmd_in_nxt[180], \gcm_dek_cmd_in_nxt.key1 [81]);
tran (gcm_dek_cmd_in_nxt[181], \gcm_dek_cmd_in_nxt.key1 [82]);
tran (gcm_dek_cmd_in_nxt[182], \gcm_dek_cmd_in_nxt.key1 [83]);
tran (gcm_dek_cmd_in_nxt[183], \gcm_dek_cmd_in_nxt.key1 [84]);
tran (gcm_dek_cmd_in_nxt[184], \gcm_dek_cmd_in_nxt.key1 [85]);
tran (gcm_dek_cmd_in_nxt[185], \gcm_dek_cmd_in_nxt.key1 [86]);
tran (gcm_dek_cmd_in_nxt[186], \gcm_dek_cmd_in_nxt.key1 [87]);
tran (gcm_dek_cmd_in_nxt[187], \gcm_dek_cmd_in_nxt.key1 [88]);
tran (gcm_dek_cmd_in_nxt[188], \gcm_dek_cmd_in_nxt.key1 [89]);
tran (gcm_dek_cmd_in_nxt[189], \gcm_dek_cmd_in_nxt.key1 [90]);
tran (gcm_dek_cmd_in_nxt[190], \gcm_dek_cmd_in_nxt.key1 [91]);
tran (gcm_dek_cmd_in_nxt[191], \gcm_dek_cmd_in_nxt.key1 [92]);
tran (gcm_dek_cmd_in_nxt[192], \gcm_dek_cmd_in_nxt.key1 [93]);
tran (gcm_dek_cmd_in_nxt[193], \gcm_dek_cmd_in_nxt.key1 [94]);
tran (gcm_dek_cmd_in_nxt[194], \gcm_dek_cmd_in_nxt.key1 [95]);
tran (gcm_dek_cmd_in_nxt[195], \gcm_dek_cmd_in_nxt.key1 [96]);
tran (gcm_dek_cmd_in_nxt[196], \gcm_dek_cmd_in_nxt.key1 [97]);
tran (gcm_dek_cmd_in_nxt[197], \gcm_dek_cmd_in_nxt.key1 [98]);
tran (gcm_dek_cmd_in_nxt[198], \gcm_dek_cmd_in_nxt.key1 [99]);
tran (gcm_dek_cmd_in_nxt[199], \gcm_dek_cmd_in_nxt.key1 [100]);
tran (gcm_dek_cmd_in_nxt[200], \gcm_dek_cmd_in_nxt.key1 [101]);
tran (gcm_dek_cmd_in_nxt[201], \gcm_dek_cmd_in_nxt.key1 [102]);
tran (gcm_dek_cmd_in_nxt[202], \gcm_dek_cmd_in_nxt.key1 [103]);
tran (gcm_dek_cmd_in_nxt[203], \gcm_dek_cmd_in_nxt.key1 [104]);
tran (gcm_dek_cmd_in_nxt[204], \gcm_dek_cmd_in_nxt.key1 [105]);
tran (gcm_dek_cmd_in_nxt[205], \gcm_dek_cmd_in_nxt.key1 [106]);
tran (gcm_dek_cmd_in_nxt[206], \gcm_dek_cmd_in_nxt.key1 [107]);
tran (gcm_dek_cmd_in_nxt[207], \gcm_dek_cmd_in_nxt.key1 [108]);
tran (gcm_dek_cmd_in_nxt[208], \gcm_dek_cmd_in_nxt.key1 [109]);
tran (gcm_dek_cmd_in_nxt[209], \gcm_dek_cmd_in_nxt.key1 [110]);
tran (gcm_dek_cmd_in_nxt[210], \gcm_dek_cmd_in_nxt.key1 [111]);
tran (gcm_dek_cmd_in_nxt[211], \gcm_dek_cmd_in_nxt.key1 [112]);
tran (gcm_dek_cmd_in_nxt[212], \gcm_dek_cmd_in_nxt.key1 [113]);
tran (gcm_dek_cmd_in_nxt[213], \gcm_dek_cmd_in_nxt.key1 [114]);
tran (gcm_dek_cmd_in_nxt[214], \gcm_dek_cmd_in_nxt.key1 [115]);
tran (gcm_dek_cmd_in_nxt[215], \gcm_dek_cmd_in_nxt.key1 [116]);
tran (gcm_dek_cmd_in_nxt[216], \gcm_dek_cmd_in_nxt.key1 [117]);
tran (gcm_dek_cmd_in_nxt[217], \gcm_dek_cmd_in_nxt.key1 [118]);
tran (gcm_dek_cmd_in_nxt[218], \gcm_dek_cmd_in_nxt.key1 [119]);
tran (gcm_dek_cmd_in_nxt[219], \gcm_dek_cmd_in_nxt.key1 [120]);
tran (gcm_dek_cmd_in_nxt[220], \gcm_dek_cmd_in_nxt.key1 [121]);
tran (gcm_dek_cmd_in_nxt[221], \gcm_dek_cmd_in_nxt.key1 [122]);
tran (gcm_dek_cmd_in_nxt[222], \gcm_dek_cmd_in_nxt.key1 [123]);
tran (gcm_dek_cmd_in_nxt[223], \gcm_dek_cmd_in_nxt.key1 [124]);
tran (gcm_dek_cmd_in_nxt[224], \gcm_dek_cmd_in_nxt.key1 [125]);
tran (gcm_dek_cmd_in_nxt[225], \gcm_dek_cmd_in_nxt.key1 [126]);
tran (gcm_dek_cmd_in_nxt[226], \gcm_dek_cmd_in_nxt.key1 [127]);
tran (gcm_dek_cmd_in_nxt[227], \gcm_dek_cmd_in_nxt.key1 [128]);
tran (gcm_dek_cmd_in_nxt[228], \gcm_dek_cmd_in_nxt.key1 [129]);
tran (gcm_dek_cmd_in_nxt[229], \gcm_dek_cmd_in_nxt.key1 [130]);
tran (gcm_dek_cmd_in_nxt[230], \gcm_dek_cmd_in_nxt.key1 [131]);
tran (gcm_dek_cmd_in_nxt[231], \gcm_dek_cmd_in_nxt.key1 [132]);
tran (gcm_dek_cmd_in_nxt[232], \gcm_dek_cmd_in_nxt.key1 [133]);
tran (gcm_dek_cmd_in_nxt[233], \gcm_dek_cmd_in_nxt.key1 [134]);
tran (gcm_dek_cmd_in_nxt[234], \gcm_dek_cmd_in_nxt.key1 [135]);
tran (gcm_dek_cmd_in_nxt[235], \gcm_dek_cmd_in_nxt.key1 [136]);
tran (gcm_dek_cmd_in_nxt[236], \gcm_dek_cmd_in_nxt.key1 [137]);
tran (gcm_dek_cmd_in_nxt[237], \gcm_dek_cmd_in_nxt.key1 [138]);
tran (gcm_dek_cmd_in_nxt[238], \gcm_dek_cmd_in_nxt.key1 [139]);
tran (gcm_dek_cmd_in_nxt[239], \gcm_dek_cmd_in_nxt.key1 [140]);
tran (gcm_dek_cmd_in_nxt[240], \gcm_dek_cmd_in_nxt.key1 [141]);
tran (gcm_dek_cmd_in_nxt[241], \gcm_dek_cmd_in_nxt.key1 [142]);
tran (gcm_dek_cmd_in_nxt[242], \gcm_dek_cmd_in_nxt.key1 [143]);
tran (gcm_dek_cmd_in_nxt[243], \gcm_dek_cmd_in_nxt.key1 [144]);
tran (gcm_dek_cmd_in_nxt[244], \gcm_dek_cmd_in_nxt.key1 [145]);
tran (gcm_dek_cmd_in_nxt[245], \gcm_dek_cmd_in_nxt.key1 [146]);
tran (gcm_dek_cmd_in_nxt[246], \gcm_dek_cmd_in_nxt.key1 [147]);
tran (gcm_dek_cmd_in_nxt[247], \gcm_dek_cmd_in_nxt.key1 [148]);
tran (gcm_dek_cmd_in_nxt[248], \gcm_dek_cmd_in_nxt.key1 [149]);
tran (gcm_dek_cmd_in_nxt[249], \gcm_dek_cmd_in_nxt.key1 [150]);
tran (gcm_dek_cmd_in_nxt[250], \gcm_dek_cmd_in_nxt.key1 [151]);
tran (gcm_dek_cmd_in_nxt[251], \gcm_dek_cmd_in_nxt.key1 [152]);
tran (gcm_dek_cmd_in_nxt[252], \gcm_dek_cmd_in_nxt.key1 [153]);
tran (gcm_dek_cmd_in_nxt[253], \gcm_dek_cmd_in_nxt.key1 [154]);
tran (gcm_dek_cmd_in_nxt[254], \gcm_dek_cmd_in_nxt.key1 [155]);
tran (gcm_dek_cmd_in_nxt[255], \gcm_dek_cmd_in_nxt.key1 [156]);
tran (gcm_dek_cmd_in_nxt[256], \gcm_dek_cmd_in_nxt.key1 [157]);
tran (gcm_dek_cmd_in_nxt[257], \gcm_dek_cmd_in_nxt.key1 [158]);
tran (gcm_dek_cmd_in_nxt[258], \gcm_dek_cmd_in_nxt.key1 [159]);
tran (gcm_dek_cmd_in_nxt[259], \gcm_dek_cmd_in_nxt.key1 [160]);
tran (gcm_dek_cmd_in_nxt[260], \gcm_dek_cmd_in_nxt.key1 [161]);
tran (gcm_dek_cmd_in_nxt[261], \gcm_dek_cmd_in_nxt.key1 [162]);
tran (gcm_dek_cmd_in_nxt[262], \gcm_dek_cmd_in_nxt.key1 [163]);
tran (gcm_dek_cmd_in_nxt[263], \gcm_dek_cmd_in_nxt.key1 [164]);
tran (gcm_dek_cmd_in_nxt[264], \gcm_dek_cmd_in_nxt.key1 [165]);
tran (gcm_dek_cmd_in_nxt[265], \gcm_dek_cmd_in_nxt.key1 [166]);
tran (gcm_dek_cmd_in_nxt[266], \gcm_dek_cmd_in_nxt.key1 [167]);
tran (gcm_dek_cmd_in_nxt[267], \gcm_dek_cmd_in_nxt.key1 [168]);
tran (gcm_dek_cmd_in_nxt[268], \gcm_dek_cmd_in_nxt.key1 [169]);
tran (gcm_dek_cmd_in_nxt[269], \gcm_dek_cmd_in_nxt.key1 [170]);
tran (gcm_dek_cmd_in_nxt[270], \gcm_dek_cmd_in_nxt.key1 [171]);
tran (gcm_dek_cmd_in_nxt[271], \gcm_dek_cmd_in_nxt.key1 [172]);
tran (gcm_dek_cmd_in_nxt[272], \gcm_dek_cmd_in_nxt.key1 [173]);
tran (gcm_dek_cmd_in_nxt[273], \gcm_dek_cmd_in_nxt.key1 [174]);
tran (gcm_dek_cmd_in_nxt[274], \gcm_dek_cmd_in_nxt.key1 [175]);
tran (gcm_dek_cmd_in_nxt[275], \gcm_dek_cmd_in_nxt.key1 [176]);
tran (gcm_dek_cmd_in_nxt[276], \gcm_dek_cmd_in_nxt.key1 [177]);
tran (gcm_dek_cmd_in_nxt[277], \gcm_dek_cmd_in_nxt.key1 [178]);
tran (gcm_dek_cmd_in_nxt[278], \gcm_dek_cmd_in_nxt.key1 [179]);
tran (gcm_dek_cmd_in_nxt[279], \gcm_dek_cmd_in_nxt.key1 [180]);
tran (gcm_dek_cmd_in_nxt[280], \gcm_dek_cmd_in_nxt.key1 [181]);
tran (gcm_dek_cmd_in_nxt[281], \gcm_dek_cmd_in_nxt.key1 [182]);
tran (gcm_dek_cmd_in_nxt[282], \gcm_dek_cmd_in_nxt.key1 [183]);
tran (gcm_dek_cmd_in_nxt[283], \gcm_dek_cmd_in_nxt.key1 [184]);
tran (gcm_dek_cmd_in_nxt[284], \gcm_dek_cmd_in_nxt.key1 [185]);
tran (gcm_dek_cmd_in_nxt[285], \gcm_dek_cmd_in_nxt.key1 [186]);
tran (gcm_dek_cmd_in_nxt[286], \gcm_dek_cmd_in_nxt.key1 [187]);
tran (gcm_dek_cmd_in_nxt[287], \gcm_dek_cmd_in_nxt.key1 [188]);
tran (gcm_dek_cmd_in_nxt[288], \gcm_dek_cmd_in_nxt.key1 [189]);
tran (gcm_dek_cmd_in_nxt[289], \gcm_dek_cmd_in_nxt.key1 [190]);
tran (gcm_dek_cmd_in_nxt[290], \gcm_dek_cmd_in_nxt.key1 [191]);
tran (gcm_dek_cmd_in_nxt[291], \gcm_dek_cmd_in_nxt.key1 [192]);
tran (gcm_dek_cmd_in_nxt[292], \gcm_dek_cmd_in_nxt.key1 [193]);
tran (gcm_dek_cmd_in_nxt[293], \gcm_dek_cmd_in_nxt.key1 [194]);
tran (gcm_dek_cmd_in_nxt[294], \gcm_dek_cmd_in_nxt.key1 [195]);
tran (gcm_dek_cmd_in_nxt[295], \gcm_dek_cmd_in_nxt.key1 [196]);
tran (gcm_dek_cmd_in_nxt[296], \gcm_dek_cmd_in_nxt.key1 [197]);
tran (gcm_dek_cmd_in_nxt[297], \gcm_dek_cmd_in_nxt.key1 [198]);
tran (gcm_dek_cmd_in_nxt[298], \gcm_dek_cmd_in_nxt.key1 [199]);
tran (gcm_dek_cmd_in_nxt[299], \gcm_dek_cmd_in_nxt.key1 [200]);
tran (gcm_dek_cmd_in_nxt[300], \gcm_dek_cmd_in_nxt.key1 [201]);
tran (gcm_dek_cmd_in_nxt[301], \gcm_dek_cmd_in_nxt.key1 [202]);
tran (gcm_dek_cmd_in_nxt[302], \gcm_dek_cmd_in_nxt.key1 [203]);
tran (gcm_dek_cmd_in_nxt[303], \gcm_dek_cmd_in_nxt.key1 [204]);
tran (gcm_dek_cmd_in_nxt[304], \gcm_dek_cmd_in_nxt.key1 [205]);
tran (gcm_dek_cmd_in_nxt[305], \gcm_dek_cmd_in_nxt.key1 [206]);
tran (gcm_dek_cmd_in_nxt[306], \gcm_dek_cmd_in_nxt.key1 [207]);
tran (gcm_dek_cmd_in_nxt[307], \gcm_dek_cmd_in_nxt.key1 [208]);
tran (gcm_dek_cmd_in_nxt[308], \gcm_dek_cmd_in_nxt.key1 [209]);
tran (gcm_dek_cmd_in_nxt[309], \gcm_dek_cmd_in_nxt.key1 [210]);
tran (gcm_dek_cmd_in_nxt[310], \gcm_dek_cmd_in_nxt.key1 [211]);
tran (gcm_dek_cmd_in_nxt[311], \gcm_dek_cmd_in_nxt.key1 [212]);
tran (gcm_dek_cmd_in_nxt[312], \gcm_dek_cmd_in_nxt.key1 [213]);
tran (gcm_dek_cmd_in_nxt[313], \gcm_dek_cmd_in_nxt.key1 [214]);
tran (gcm_dek_cmd_in_nxt[314], \gcm_dek_cmd_in_nxt.key1 [215]);
tran (gcm_dek_cmd_in_nxt[315], \gcm_dek_cmd_in_nxt.key1 [216]);
tran (gcm_dek_cmd_in_nxt[316], \gcm_dek_cmd_in_nxt.key1 [217]);
tran (gcm_dek_cmd_in_nxt[317], \gcm_dek_cmd_in_nxt.key1 [218]);
tran (gcm_dek_cmd_in_nxt[318], \gcm_dek_cmd_in_nxt.key1 [219]);
tran (gcm_dek_cmd_in_nxt[319], \gcm_dek_cmd_in_nxt.key1 [220]);
tran (gcm_dek_cmd_in_nxt[320], \gcm_dek_cmd_in_nxt.key1 [221]);
tran (gcm_dek_cmd_in_nxt[321], \gcm_dek_cmd_in_nxt.key1 [222]);
tran (gcm_dek_cmd_in_nxt[322], \gcm_dek_cmd_in_nxt.key1 [223]);
tran (gcm_dek_cmd_in_nxt[323], \gcm_dek_cmd_in_nxt.key1 [224]);
tran (gcm_dek_cmd_in_nxt[324], \gcm_dek_cmd_in_nxt.key1 [225]);
tran (gcm_dek_cmd_in_nxt[325], \gcm_dek_cmd_in_nxt.key1 [226]);
tran (gcm_dek_cmd_in_nxt[326], \gcm_dek_cmd_in_nxt.key1 [227]);
tran (gcm_dek_cmd_in_nxt[327], \gcm_dek_cmd_in_nxt.key1 [228]);
tran (gcm_dek_cmd_in_nxt[328], \gcm_dek_cmd_in_nxt.key1 [229]);
tran (gcm_dek_cmd_in_nxt[329], \gcm_dek_cmd_in_nxt.key1 [230]);
tran (gcm_dek_cmd_in_nxt[330], \gcm_dek_cmd_in_nxt.key1 [231]);
tran (gcm_dek_cmd_in_nxt[331], \gcm_dek_cmd_in_nxt.key1 [232]);
tran (gcm_dek_cmd_in_nxt[332], \gcm_dek_cmd_in_nxt.key1 [233]);
tran (gcm_dek_cmd_in_nxt[333], \gcm_dek_cmd_in_nxt.key1 [234]);
tran (gcm_dek_cmd_in_nxt[334], \gcm_dek_cmd_in_nxt.key1 [235]);
tran (gcm_dek_cmd_in_nxt[335], \gcm_dek_cmd_in_nxt.key1 [236]);
tran (gcm_dek_cmd_in_nxt[336], \gcm_dek_cmd_in_nxt.key1 [237]);
tran (gcm_dek_cmd_in_nxt[337], \gcm_dek_cmd_in_nxt.key1 [238]);
tran (gcm_dek_cmd_in_nxt[338], \gcm_dek_cmd_in_nxt.key1 [239]);
tran (gcm_dek_cmd_in_nxt[339], \gcm_dek_cmd_in_nxt.key1 [240]);
tran (gcm_dek_cmd_in_nxt[340], \gcm_dek_cmd_in_nxt.key1 [241]);
tran (gcm_dek_cmd_in_nxt[341], \gcm_dek_cmd_in_nxt.key1 [242]);
tran (gcm_dek_cmd_in_nxt[342], \gcm_dek_cmd_in_nxt.key1 [243]);
tran (gcm_dek_cmd_in_nxt[343], \gcm_dek_cmd_in_nxt.key1 [244]);
tran (gcm_dek_cmd_in_nxt[344], \gcm_dek_cmd_in_nxt.key1 [245]);
tran (gcm_dek_cmd_in_nxt[345], \gcm_dek_cmd_in_nxt.key1 [246]);
tran (gcm_dek_cmd_in_nxt[346], \gcm_dek_cmd_in_nxt.key1 [247]);
tran (gcm_dek_cmd_in_nxt[347], \gcm_dek_cmd_in_nxt.key1 [248]);
tran (gcm_dek_cmd_in_nxt[348], \gcm_dek_cmd_in_nxt.key1 [249]);
tran (gcm_dek_cmd_in_nxt[349], \gcm_dek_cmd_in_nxt.key1 [250]);
tran (gcm_dek_cmd_in_nxt[350], \gcm_dek_cmd_in_nxt.key1 [251]);
tran (gcm_dek_cmd_in_nxt[351], \gcm_dek_cmd_in_nxt.key1 [252]);
tran (gcm_dek_cmd_in_nxt[352], \gcm_dek_cmd_in_nxt.key1 [253]);
tran (gcm_dek_cmd_in_nxt[353], \gcm_dek_cmd_in_nxt.key1 [254]);
tran (gcm_dek_cmd_in_nxt[354], \gcm_dek_cmd_in_nxt.key1 [255]);
tran (gcm_dek_cmd_in_nxt[355], \gcm_dek_cmd_in_nxt.key0 [0]);
tran (gcm_dek_cmd_in_nxt[356], \gcm_dek_cmd_in_nxt.key0 [1]);
tran (gcm_dek_cmd_in_nxt[357], \gcm_dek_cmd_in_nxt.key0 [2]);
tran (gcm_dek_cmd_in_nxt[358], \gcm_dek_cmd_in_nxt.key0 [3]);
tran (gcm_dek_cmd_in_nxt[359], \gcm_dek_cmd_in_nxt.key0 [4]);
tran (gcm_dek_cmd_in_nxt[360], \gcm_dek_cmd_in_nxt.key0 [5]);
tran (gcm_dek_cmd_in_nxt[361], \gcm_dek_cmd_in_nxt.key0 [6]);
tran (gcm_dek_cmd_in_nxt[362], \gcm_dek_cmd_in_nxt.key0 [7]);
tran (gcm_dek_cmd_in_nxt[363], \gcm_dek_cmd_in_nxt.key0 [8]);
tran (gcm_dek_cmd_in_nxt[364], \gcm_dek_cmd_in_nxt.key0 [9]);
tran (gcm_dek_cmd_in_nxt[365], \gcm_dek_cmd_in_nxt.key0 [10]);
tran (gcm_dek_cmd_in_nxt[366], \gcm_dek_cmd_in_nxt.key0 [11]);
tran (gcm_dek_cmd_in_nxt[367], \gcm_dek_cmd_in_nxt.key0 [12]);
tran (gcm_dek_cmd_in_nxt[368], \gcm_dek_cmd_in_nxt.key0 [13]);
tran (gcm_dek_cmd_in_nxt[369], \gcm_dek_cmd_in_nxt.key0 [14]);
tran (gcm_dek_cmd_in_nxt[370], \gcm_dek_cmd_in_nxt.key0 [15]);
tran (gcm_dek_cmd_in_nxt[371], \gcm_dek_cmd_in_nxt.key0 [16]);
tran (gcm_dek_cmd_in_nxt[372], \gcm_dek_cmd_in_nxt.key0 [17]);
tran (gcm_dek_cmd_in_nxt[373], \gcm_dek_cmd_in_nxt.key0 [18]);
tran (gcm_dek_cmd_in_nxt[374], \gcm_dek_cmd_in_nxt.key0 [19]);
tran (gcm_dek_cmd_in_nxt[375], \gcm_dek_cmd_in_nxt.key0 [20]);
tran (gcm_dek_cmd_in_nxt[376], \gcm_dek_cmd_in_nxt.key0 [21]);
tran (gcm_dek_cmd_in_nxt[377], \gcm_dek_cmd_in_nxt.key0 [22]);
tran (gcm_dek_cmd_in_nxt[378], \gcm_dek_cmd_in_nxt.key0 [23]);
tran (gcm_dek_cmd_in_nxt[379], \gcm_dek_cmd_in_nxt.key0 [24]);
tran (gcm_dek_cmd_in_nxt[380], \gcm_dek_cmd_in_nxt.key0 [25]);
tran (gcm_dek_cmd_in_nxt[381], \gcm_dek_cmd_in_nxt.key0 [26]);
tran (gcm_dek_cmd_in_nxt[382], \gcm_dek_cmd_in_nxt.key0 [27]);
tran (gcm_dek_cmd_in_nxt[383], \gcm_dek_cmd_in_nxt.key0 [28]);
tran (gcm_dek_cmd_in_nxt[384], \gcm_dek_cmd_in_nxt.key0 [29]);
tran (gcm_dek_cmd_in_nxt[385], \gcm_dek_cmd_in_nxt.key0 [30]);
tran (gcm_dek_cmd_in_nxt[386], \gcm_dek_cmd_in_nxt.key0 [31]);
tran (gcm_dek_cmd_in_nxt[387], \gcm_dek_cmd_in_nxt.key0 [32]);
tran (gcm_dek_cmd_in_nxt[388], \gcm_dek_cmd_in_nxt.key0 [33]);
tran (gcm_dek_cmd_in_nxt[389], \gcm_dek_cmd_in_nxt.key0 [34]);
tran (gcm_dek_cmd_in_nxt[390], \gcm_dek_cmd_in_nxt.key0 [35]);
tran (gcm_dek_cmd_in_nxt[391], \gcm_dek_cmd_in_nxt.key0 [36]);
tran (gcm_dek_cmd_in_nxt[392], \gcm_dek_cmd_in_nxt.key0 [37]);
tran (gcm_dek_cmd_in_nxt[393], \gcm_dek_cmd_in_nxt.key0 [38]);
tran (gcm_dek_cmd_in_nxt[394], \gcm_dek_cmd_in_nxt.key0 [39]);
tran (gcm_dek_cmd_in_nxt[395], \gcm_dek_cmd_in_nxt.key0 [40]);
tran (gcm_dek_cmd_in_nxt[396], \gcm_dek_cmd_in_nxt.key0 [41]);
tran (gcm_dek_cmd_in_nxt[397], \gcm_dek_cmd_in_nxt.key0 [42]);
tran (gcm_dek_cmd_in_nxt[398], \gcm_dek_cmd_in_nxt.key0 [43]);
tran (gcm_dek_cmd_in_nxt[399], \gcm_dek_cmd_in_nxt.key0 [44]);
tran (gcm_dek_cmd_in_nxt[400], \gcm_dek_cmd_in_nxt.key0 [45]);
tran (gcm_dek_cmd_in_nxt[401], \gcm_dek_cmd_in_nxt.key0 [46]);
tran (gcm_dek_cmd_in_nxt[402], \gcm_dek_cmd_in_nxt.key0 [47]);
tran (gcm_dek_cmd_in_nxt[403], \gcm_dek_cmd_in_nxt.key0 [48]);
tran (gcm_dek_cmd_in_nxt[404], \gcm_dek_cmd_in_nxt.key0 [49]);
tran (gcm_dek_cmd_in_nxt[405], \gcm_dek_cmd_in_nxt.key0 [50]);
tran (gcm_dek_cmd_in_nxt[406], \gcm_dek_cmd_in_nxt.key0 [51]);
tran (gcm_dek_cmd_in_nxt[407], \gcm_dek_cmd_in_nxt.key0 [52]);
tran (gcm_dek_cmd_in_nxt[408], \gcm_dek_cmd_in_nxt.key0 [53]);
tran (gcm_dek_cmd_in_nxt[409], \gcm_dek_cmd_in_nxt.key0 [54]);
tran (gcm_dek_cmd_in_nxt[410], \gcm_dek_cmd_in_nxt.key0 [55]);
tran (gcm_dek_cmd_in_nxt[411], \gcm_dek_cmd_in_nxt.key0 [56]);
tran (gcm_dek_cmd_in_nxt[412], \gcm_dek_cmd_in_nxt.key0 [57]);
tran (gcm_dek_cmd_in_nxt[413], \gcm_dek_cmd_in_nxt.key0 [58]);
tran (gcm_dek_cmd_in_nxt[414], \gcm_dek_cmd_in_nxt.key0 [59]);
tran (gcm_dek_cmd_in_nxt[415], \gcm_dek_cmd_in_nxt.key0 [60]);
tran (gcm_dek_cmd_in_nxt[416], \gcm_dek_cmd_in_nxt.key0 [61]);
tran (gcm_dek_cmd_in_nxt[417], \gcm_dek_cmd_in_nxt.key0 [62]);
tran (gcm_dek_cmd_in_nxt[418], \gcm_dek_cmd_in_nxt.key0 [63]);
tran (gcm_dek_cmd_in_nxt[419], \gcm_dek_cmd_in_nxt.key0 [64]);
tran (gcm_dek_cmd_in_nxt[420], \gcm_dek_cmd_in_nxt.key0 [65]);
tran (gcm_dek_cmd_in_nxt[421], \gcm_dek_cmd_in_nxt.key0 [66]);
tran (gcm_dek_cmd_in_nxt[422], \gcm_dek_cmd_in_nxt.key0 [67]);
tran (gcm_dek_cmd_in_nxt[423], \gcm_dek_cmd_in_nxt.key0 [68]);
tran (gcm_dek_cmd_in_nxt[424], \gcm_dek_cmd_in_nxt.key0 [69]);
tran (gcm_dek_cmd_in_nxt[425], \gcm_dek_cmd_in_nxt.key0 [70]);
tran (gcm_dek_cmd_in_nxt[426], \gcm_dek_cmd_in_nxt.key0 [71]);
tran (gcm_dek_cmd_in_nxt[427], \gcm_dek_cmd_in_nxt.key0 [72]);
tran (gcm_dek_cmd_in_nxt[428], \gcm_dek_cmd_in_nxt.key0 [73]);
tran (gcm_dek_cmd_in_nxt[429], \gcm_dek_cmd_in_nxt.key0 [74]);
tran (gcm_dek_cmd_in_nxt[430], \gcm_dek_cmd_in_nxt.key0 [75]);
tran (gcm_dek_cmd_in_nxt[431], \gcm_dek_cmd_in_nxt.key0 [76]);
tran (gcm_dek_cmd_in_nxt[432], \gcm_dek_cmd_in_nxt.key0 [77]);
tran (gcm_dek_cmd_in_nxt[433], \gcm_dek_cmd_in_nxt.key0 [78]);
tran (gcm_dek_cmd_in_nxt[434], \gcm_dek_cmd_in_nxt.key0 [79]);
tran (gcm_dek_cmd_in_nxt[435], \gcm_dek_cmd_in_nxt.key0 [80]);
tran (gcm_dek_cmd_in_nxt[436], \gcm_dek_cmd_in_nxt.key0 [81]);
tran (gcm_dek_cmd_in_nxt[437], \gcm_dek_cmd_in_nxt.key0 [82]);
tran (gcm_dek_cmd_in_nxt[438], \gcm_dek_cmd_in_nxt.key0 [83]);
tran (gcm_dek_cmd_in_nxt[439], \gcm_dek_cmd_in_nxt.key0 [84]);
tran (gcm_dek_cmd_in_nxt[440], \gcm_dek_cmd_in_nxt.key0 [85]);
tran (gcm_dek_cmd_in_nxt[441], \gcm_dek_cmd_in_nxt.key0 [86]);
tran (gcm_dek_cmd_in_nxt[442], \gcm_dek_cmd_in_nxt.key0 [87]);
tran (gcm_dek_cmd_in_nxt[443], \gcm_dek_cmd_in_nxt.key0 [88]);
tran (gcm_dek_cmd_in_nxt[444], \gcm_dek_cmd_in_nxt.key0 [89]);
tran (gcm_dek_cmd_in_nxt[445], \gcm_dek_cmd_in_nxt.key0 [90]);
tran (gcm_dek_cmd_in_nxt[446], \gcm_dek_cmd_in_nxt.key0 [91]);
tran (gcm_dek_cmd_in_nxt[447], \gcm_dek_cmd_in_nxt.key0 [92]);
tran (gcm_dek_cmd_in_nxt[448], \gcm_dek_cmd_in_nxt.key0 [93]);
tran (gcm_dek_cmd_in_nxt[449], \gcm_dek_cmd_in_nxt.key0 [94]);
tran (gcm_dek_cmd_in_nxt[450], \gcm_dek_cmd_in_nxt.key0 [95]);
tran (gcm_dek_cmd_in_nxt[451], \gcm_dek_cmd_in_nxt.key0 [96]);
tran (gcm_dek_cmd_in_nxt[452], \gcm_dek_cmd_in_nxt.key0 [97]);
tran (gcm_dek_cmd_in_nxt[453], \gcm_dek_cmd_in_nxt.key0 [98]);
tran (gcm_dek_cmd_in_nxt[454], \gcm_dek_cmd_in_nxt.key0 [99]);
tran (gcm_dek_cmd_in_nxt[455], \gcm_dek_cmd_in_nxt.key0 [100]);
tran (gcm_dek_cmd_in_nxt[456], \gcm_dek_cmd_in_nxt.key0 [101]);
tran (gcm_dek_cmd_in_nxt[457], \gcm_dek_cmd_in_nxt.key0 [102]);
tran (gcm_dek_cmd_in_nxt[458], \gcm_dek_cmd_in_nxt.key0 [103]);
tran (gcm_dek_cmd_in_nxt[459], \gcm_dek_cmd_in_nxt.key0 [104]);
tran (gcm_dek_cmd_in_nxt[460], \gcm_dek_cmd_in_nxt.key0 [105]);
tran (gcm_dek_cmd_in_nxt[461], \gcm_dek_cmd_in_nxt.key0 [106]);
tran (gcm_dek_cmd_in_nxt[462], \gcm_dek_cmd_in_nxt.key0 [107]);
tran (gcm_dek_cmd_in_nxt[463], \gcm_dek_cmd_in_nxt.key0 [108]);
tran (gcm_dek_cmd_in_nxt[464], \gcm_dek_cmd_in_nxt.key0 [109]);
tran (gcm_dek_cmd_in_nxt[465], \gcm_dek_cmd_in_nxt.key0 [110]);
tran (gcm_dek_cmd_in_nxt[466], \gcm_dek_cmd_in_nxt.key0 [111]);
tran (gcm_dek_cmd_in_nxt[467], \gcm_dek_cmd_in_nxt.key0 [112]);
tran (gcm_dek_cmd_in_nxt[468], \gcm_dek_cmd_in_nxt.key0 [113]);
tran (gcm_dek_cmd_in_nxt[469], \gcm_dek_cmd_in_nxt.key0 [114]);
tran (gcm_dek_cmd_in_nxt[470], \gcm_dek_cmd_in_nxt.key0 [115]);
tran (gcm_dek_cmd_in_nxt[471], \gcm_dek_cmd_in_nxt.key0 [116]);
tran (gcm_dek_cmd_in_nxt[472], \gcm_dek_cmd_in_nxt.key0 [117]);
tran (gcm_dek_cmd_in_nxt[473], \gcm_dek_cmd_in_nxt.key0 [118]);
tran (gcm_dek_cmd_in_nxt[474], \gcm_dek_cmd_in_nxt.key0 [119]);
tran (gcm_dek_cmd_in_nxt[475], \gcm_dek_cmd_in_nxt.key0 [120]);
tran (gcm_dek_cmd_in_nxt[476], \gcm_dek_cmd_in_nxt.key0 [121]);
tran (gcm_dek_cmd_in_nxt[477], \gcm_dek_cmd_in_nxt.key0 [122]);
tran (gcm_dek_cmd_in_nxt[478], \gcm_dek_cmd_in_nxt.key0 [123]);
tran (gcm_dek_cmd_in_nxt[479], \gcm_dek_cmd_in_nxt.key0 [124]);
tran (gcm_dek_cmd_in_nxt[480], \gcm_dek_cmd_in_nxt.key0 [125]);
tran (gcm_dek_cmd_in_nxt[481], \gcm_dek_cmd_in_nxt.key0 [126]);
tran (gcm_dek_cmd_in_nxt[482], \gcm_dek_cmd_in_nxt.key0 [127]);
tran (gcm_dek_cmd_in_nxt[483], \gcm_dek_cmd_in_nxt.key0 [128]);
tran (gcm_dek_cmd_in_nxt[484], \gcm_dek_cmd_in_nxt.key0 [129]);
tran (gcm_dek_cmd_in_nxt[485], \gcm_dek_cmd_in_nxt.key0 [130]);
tran (gcm_dek_cmd_in_nxt[486], \gcm_dek_cmd_in_nxt.key0 [131]);
tran (gcm_dek_cmd_in_nxt[487], \gcm_dek_cmd_in_nxt.key0 [132]);
tran (gcm_dek_cmd_in_nxt[488], \gcm_dek_cmd_in_nxt.key0 [133]);
tran (gcm_dek_cmd_in_nxt[489], \gcm_dek_cmd_in_nxt.key0 [134]);
tran (gcm_dek_cmd_in_nxt[490], \gcm_dek_cmd_in_nxt.key0 [135]);
tran (gcm_dek_cmd_in_nxt[491], \gcm_dek_cmd_in_nxt.key0 [136]);
tran (gcm_dek_cmd_in_nxt[492], \gcm_dek_cmd_in_nxt.key0 [137]);
tran (gcm_dek_cmd_in_nxt[493], \gcm_dek_cmd_in_nxt.key0 [138]);
tran (gcm_dek_cmd_in_nxt[494], \gcm_dek_cmd_in_nxt.key0 [139]);
tran (gcm_dek_cmd_in_nxt[495], \gcm_dek_cmd_in_nxt.key0 [140]);
tran (gcm_dek_cmd_in_nxt[496], \gcm_dek_cmd_in_nxt.key0 [141]);
tran (gcm_dek_cmd_in_nxt[497], \gcm_dek_cmd_in_nxt.key0 [142]);
tran (gcm_dek_cmd_in_nxt[498], \gcm_dek_cmd_in_nxt.key0 [143]);
tran (gcm_dek_cmd_in_nxt[499], \gcm_dek_cmd_in_nxt.key0 [144]);
tran (gcm_dek_cmd_in_nxt[500], \gcm_dek_cmd_in_nxt.key0 [145]);
tran (gcm_dek_cmd_in_nxt[501], \gcm_dek_cmd_in_nxt.key0 [146]);
tran (gcm_dek_cmd_in_nxt[502], \gcm_dek_cmd_in_nxt.key0 [147]);
tran (gcm_dek_cmd_in_nxt[503], \gcm_dek_cmd_in_nxt.key0 [148]);
tran (gcm_dek_cmd_in_nxt[504], \gcm_dek_cmd_in_nxt.key0 [149]);
tran (gcm_dek_cmd_in_nxt[505], \gcm_dek_cmd_in_nxt.key0 [150]);
tran (gcm_dek_cmd_in_nxt[506], \gcm_dek_cmd_in_nxt.key0 [151]);
tran (gcm_dek_cmd_in_nxt[507], \gcm_dek_cmd_in_nxt.key0 [152]);
tran (gcm_dek_cmd_in_nxt[508], \gcm_dek_cmd_in_nxt.key0 [153]);
tran (gcm_dek_cmd_in_nxt[509], \gcm_dek_cmd_in_nxt.key0 [154]);
tran (gcm_dek_cmd_in_nxt[510], \gcm_dek_cmd_in_nxt.key0 [155]);
tran (gcm_dek_cmd_in_nxt[511], \gcm_dek_cmd_in_nxt.key0 [156]);
tran (gcm_dek_cmd_in_nxt[512], \gcm_dek_cmd_in_nxt.key0 [157]);
tran (gcm_dek_cmd_in_nxt[513], \gcm_dek_cmd_in_nxt.key0 [158]);
tran (gcm_dek_cmd_in_nxt[514], \gcm_dek_cmd_in_nxt.key0 [159]);
tran (gcm_dek_cmd_in_nxt[515], \gcm_dek_cmd_in_nxt.key0 [160]);
tran (gcm_dek_cmd_in_nxt[516], \gcm_dek_cmd_in_nxt.key0 [161]);
tran (gcm_dek_cmd_in_nxt[517], \gcm_dek_cmd_in_nxt.key0 [162]);
tran (gcm_dek_cmd_in_nxt[518], \gcm_dek_cmd_in_nxt.key0 [163]);
tran (gcm_dek_cmd_in_nxt[519], \gcm_dek_cmd_in_nxt.key0 [164]);
tran (gcm_dek_cmd_in_nxt[520], \gcm_dek_cmd_in_nxt.key0 [165]);
tran (gcm_dek_cmd_in_nxt[521], \gcm_dek_cmd_in_nxt.key0 [166]);
tran (gcm_dek_cmd_in_nxt[522], \gcm_dek_cmd_in_nxt.key0 [167]);
tran (gcm_dek_cmd_in_nxt[523], \gcm_dek_cmd_in_nxt.key0 [168]);
tran (gcm_dek_cmd_in_nxt[524], \gcm_dek_cmd_in_nxt.key0 [169]);
tran (gcm_dek_cmd_in_nxt[525], \gcm_dek_cmd_in_nxt.key0 [170]);
tran (gcm_dek_cmd_in_nxt[526], \gcm_dek_cmd_in_nxt.key0 [171]);
tran (gcm_dek_cmd_in_nxt[527], \gcm_dek_cmd_in_nxt.key0 [172]);
tran (gcm_dek_cmd_in_nxt[528], \gcm_dek_cmd_in_nxt.key0 [173]);
tran (gcm_dek_cmd_in_nxt[529], \gcm_dek_cmd_in_nxt.key0 [174]);
tran (gcm_dek_cmd_in_nxt[530], \gcm_dek_cmd_in_nxt.key0 [175]);
tran (gcm_dek_cmd_in_nxt[531], \gcm_dek_cmd_in_nxt.key0 [176]);
tran (gcm_dek_cmd_in_nxt[532], \gcm_dek_cmd_in_nxt.key0 [177]);
tran (gcm_dek_cmd_in_nxt[533], \gcm_dek_cmd_in_nxt.key0 [178]);
tran (gcm_dek_cmd_in_nxt[534], \gcm_dek_cmd_in_nxt.key0 [179]);
tran (gcm_dek_cmd_in_nxt[535], \gcm_dek_cmd_in_nxt.key0 [180]);
tran (gcm_dek_cmd_in_nxt[536], \gcm_dek_cmd_in_nxt.key0 [181]);
tran (gcm_dek_cmd_in_nxt[537], \gcm_dek_cmd_in_nxt.key0 [182]);
tran (gcm_dek_cmd_in_nxt[538], \gcm_dek_cmd_in_nxt.key0 [183]);
tran (gcm_dek_cmd_in_nxt[539], \gcm_dek_cmd_in_nxt.key0 [184]);
tran (gcm_dek_cmd_in_nxt[540], \gcm_dek_cmd_in_nxt.key0 [185]);
tran (gcm_dek_cmd_in_nxt[541], \gcm_dek_cmd_in_nxt.key0 [186]);
tran (gcm_dek_cmd_in_nxt[542], \gcm_dek_cmd_in_nxt.key0 [187]);
tran (gcm_dek_cmd_in_nxt[543], \gcm_dek_cmd_in_nxt.key0 [188]);
tran (gcm_dek_cmd_in_nxt[544], \gcm_dek_cmd_in_nxt.key0 [189]);
tran (gcm_dek_cmd_in_nxt[545], \gcm_dek_cmd_in_nxt.key0 [190]);
tran (gcm_dek_cmd_in_nxt[546], \gcm_dek_cmd_in_nxt.key0 [191]);
tran (gcm_dek_cmd_in_nxt[547], \gcm_dek_cmd_in_nxt.key0 [192]);
tran (gcm_dek_cmd_in_nxt[548], \gcm_dek_cmd_in_nxt.key0 [193]);
tran (gcm_dek_cmd_in_nxt[549], \gcm_dek_cmd_in_nxt.key0 [194]);
tran (gcm_dek_cmd_in_nxt[550], \gcm_dek_cmd_in_nxt.key0 [195]);
tran (gcm_dek_cmd_in_nxt[551], \gcm_dek_cmd_in_nxt.key0 [196]);
tran (gcm_dek_cmd_in_nxt[552], \gcm_dek_cmd_in_nxt.key0 [197]);
tran (gcm_dek_cmd_in_nxt[553], \gcm_dek_cmd_in_nxt.key0 [198]);
tran (gcm_dek_cmd_in_nxt[554], \gcm_dek_cmd_in_nxt.key0 [199]);
tran (gcm_dek_cmd_in_nxt[555], \gcm_dek_cmd_in_nxt.key0 [200]);
tran (gcm_dek_cmd_in_nxt[556], \gcm_dek_cmd_in_nxt.key0 [201]);
tran (gcm_dek_cmd_in_nxt[557], \gcm_dek_cmd_in_nxt.key0 [202]);
tran (gcm_dek_cmd_in_nxt[558], \gcm_dek_cmd_in_nxt.key0 [203]);
tran (gcm_dek_cmd_in_nxt[559], \gcm_dek_cmd_in_nxt.key0 [204]);
tran (gcm_dek_cmd_in_nxt[560], \gcm_dek_cmd_in_nxt.key0 [205]);
tran (gcm_dek_cmd_in_nxt[561], \gcm_dek_cmd_in_nxt.key0 [206]);
tran (gcm_dek_cmd_in_nxt[562], \gcm_dek_cmd_in_nxt.key0 [207]);
tran (gcm_dek_cmd_in_nxt[563], \gcm_dek_cmd_in_nxt.key0 [208]);
tran (gcm_dek_cmd_in_nxt[564], \gcm_dek_cmd_in_nxt.key0 [209]);
tran (gcm_dek_cmd_in_nxt[565], \gcm_dek_cmd_in_nxt.key0 [210]);
tran (gcm_dek_cmd_in_nxt[566], \gcm_dek_cmd_in_nxt.key0 [211]);
tran (gcm_dek_cmd_in_nxt[567], \gcm_dek_cmd_in_nxt.key0 [212]);
tran (gcm_dek_cmd_in_nxt[568], \gcm_dek_cmd_in_nxt.key0 [213]);
tran (gcm_dek_cmd_in_nxt[569], \gcm_dek_cmd_in_nxt.key0 [214]);
tran (gcm_dek_cmd_in_nxt[570], \gcm_dek_cmd_in_nxt.key0 [215]);
tran (gcm_dek_cmd_in_nxt[571], \gcm_dek_cmd_in_nxt.key0 [216]);
tran (gcm_dek_cmd_in_nxt[572], \gcm_dek_cmd_in_nxt.key0 [217]);
tran (gcm_dek_cmd_in_nxt[573], \gcm_dek_cmd_in_nxt.key0 [218]);
tran (gcm_dek_cmd_in_nxt[574], \gcm_dek_cmd_in_nxt.key0 [219]);
tran (gcm_dek_cmd_in_nxt[575], \gcm_dek_cmd_in_nxt.key0 [220]);
tran (gcm_dek_cmd_in_nxt[576], \gcm_dek_cmd_in_nxt.key0 [221]);
tran (gcm_dek_cmd_in_nxt[577], \gcm_dek_cmd_in_nxt.key0 [222]);
tran (gcm_dek_cmd_in_nxt[578], \gcm_dek_cmd_in_nxt.key0 [223]);
tran (gcm_dek_cmd_in_nxt[579], \gcm_dek_cmd_in_nxt.key0 [224]);
tran (gcm_dek_cmd_in_nxt[580], \gcm_dek_cmd_in_nxt.key0 [225]);
tran (gcm_dek_cmd_in_nxt[581], \gcm_dek_cmd_in_nxt.key0 [226]);
tran (gcm_dek_cmd_in_nxt[582], \gcm_dek_cmd_in_nxt.key0 [227]);
tran (gcm_dek_cmd_in_nxt[583], \gcm_dek_cmd_in_nxt.key0 [228]);
tran (gcm_dek_cmd_in_nxt[584], \gcm_dek_cmd_in_nxt.key0 [229]);
tran (gcm_dek_cmd_in_nxt[585], \gcm_dek_cmd_in_nxt.key0 [230]);
tran (gcm_dek_cmd_in_nxt[586], \gcm_dek_cmd_in_nxt.key0 [231]);
tran (gcm_dek_cmd_in_nxt[587], \gcm_dek_cmd_in_nxt.key0 [232]);
tran (gcm_dek_cmd_in_nxt[588], \gcm_dek_cmd_in_nxt.key0 [233]);
tran (gcm_dek_cmd_in_nxt[589], \gcm_dek_cmd_in_nxt.key0 [234]);
tran (gcm_dek_cmd_in_nxt[590], \gcm_dek_cmd_in_nxt.key0 [235]);
tran (gcm_dek_cmd_in_nxt[591], \gcm_dek_cmd_in_nxt.key0 [236]);
tran (gcm_dek_cmd_in_nxt[592], \gcm_dek_cmd_in_nxt.key0 [237]);
tran (gcm_dek_cmd_in_nxt[593], \gcm_dek_cmd_in_nxt.key0 [238]);
tran (gcm_dek_cmd_in_nxt[594], \gcm_dek_cmd_in_nxt.key0 [239]);
tran (gcm_dek_cmd_in_nxt[595], \gcm_dek_cmd_in_nxt.key0 [240]);
tran (gcm_dek_cmd_in_nxt[596], \gcm_dek_cmd_in_nxt.key0 [241]);
tran (gcm_dek_cmd_in_nxt[597], \gcm_dek_cmd_in_nxt.key0 [242]);
tran (gcm_dek_cmd_in_nxt[598], \gcm_dek_cmd_in_nxt.key0 [243]);
tran (gcm_dek_cmd_in_nxt[599], \gcm_dek_cmd_in_nxt.key0 [244]);
tran (gcm_dek_cmd_in_nxt[600], \gcm_dek_cmd_in_nxt.key0 [245]);
tran (gcm_dek_cmd_in_nxt[601], \gcm_dek_cmd_in_nxt.key0 [246]);
tran (gcm_dek_cmd_in_nxt[602], \gcm_dek_cmd_in_nxt.key0 [247]);
tran (gcm_dek_cmd_in_nxt[603], \gcm_dek_cmd_in_nxt.key0 [248]);
tran (gcm_dek_cmd_in_nxt[604], \gcm_dek_cmd_in_nxt.key0 [249]);
tran (gcm_dek_cmd_in_nxt[605], \gcm_dek_cmd_in_nxt.key0 [250]);
tran (gcm_dek_cmd_in_nxt[606], \gcm_dek_cmd_in_nxt.key0 [251]);
tran (gcm_dek_cmd_in_nxt[607], \gcm_dek_cmd_in_nxt.key0 [252]);
tran (gcm_dek_cmd_in_nxt[608], \gcm_dek_cmd_in_nxt.key0 [253]);
tran (gcm_dek_cmd_in_nxt[609], \gcm_dek_cmd_in_nxt.key0 [254]);
tran (gcm_dek_cmd_in_nxt[610], \gcm_dek_cmd_in_nxt.key0 [255]);
tran (stream_cmd_in_nxt[0], \stream_cmd_in_nxt.num_iter [0]);
tran (stream_cmd_in_nxt[1], \stream_cmd_in_nxt.num_iter [1]);
tran (stream_cmd_in_nxt[2], \stream_cmd_in_nxt.label_index [0]);
tran (stream_cmd_in_nxt[3], \stream_cmd_in_nxt.label_index [1]);
tran (stream_cmd_in_nxt[4], \stream_cmd_in_nxt.label_index [2]);
tran (stream_cmd_in_nxt[5], \stream_cmd_in_nxt.guid [0]);
tran (stream_cmd_in_nxt[6], \stream_cmd_in_nxt.guid [1]);
tran (stream_cmd_in_nxt[7], \stream_cmd_in_nxt.guid [2]);
tran (stream_cmd_in_nxt[8], \stream_cmd_in_nxt.guid [3]);
tran (stream_cmd_in_nxt[9], \stream_cmd_in_nxt.guid [4]);
tran (stream_cmd_in_nxt[10], \stream_cmd_in_nxt.guid [5]);
tran (stream_cmd_in_nxt[11], \stream_cmd_in_nxt.guid [6]);
tran (stream_cmd_in_nxt[12], \stream_cmd_in_nxt.guid [7]);
tran (stream_cmd_in_nxt[13], \stream_cmd_in_nxt.guid [8]);
tran (stream_cmd_in_nxt[14], \stream_cmd_in_nxt.guid [9]);
tran (stream_cmd_in_nxt[15], \stream_cmd_in_nxt.guid [10]);
tran (stream_cmd_in_nxt[16], \stream_cmd_in_nxt.guid [11]);
tran (stream_cmd_in_nxt[17], \stream_cmd_in_nxt.guid [12]);
tran (stream_cmd_in_nxt[18], \stream_cmd_in_nxt.guid [13]);
tran (stream_cmd_in_nxt[19], \stream_cmd_in_nxt.guid [14]);
tran (stream_cmd_in_nxt[20], \stream_cmd_in_nxt.guid [15]);
tran (stream_cmd_in_nxt[21], \stream_cmd_in_nxt.guid [16]);
tran (stream_cmd_in_nxt[22], \stream_cmd_in_nxt.guid [17]);
tran (stream_cmd_in_nxt[23], \stream_cmd_in_nxt.guid [18]);
tran (stream_cmd_in_nxt[24], \stream_cmd_in_nxt.guid [19]);
tran (stream_cmd_in_nxt[25], \stream_cmd_in_nxt.guid [20]);
tran (stream_cmd_in_nxt[26], \stream_cmd_in_nxt.guid [21]);
tran (stream_cmd_in_nxt[27], \stream_cmd_in_nxt.guid [22]);
tran (stream_cmd_in_nxt[28], \stream_cmd_in_nxt.guid [23]);
tran (stream_cmd_in_nxt[29], \stream_cmd_in_nxt.guid [24]);
tran (stream_cmd_in_nxt[30], \stream_cmd_in_nxt.guid [25]);
tran (stream_cmd_in_nxt[31], \stream_cmd_in_nxt.guid [26]);
tran (stream_cmd_in_nxt[32], \stream_cmd_in_nxt.guid [27]);
tran (stream_cmd_in_nxt[33], \stream_cmd_in_nxt.guid [28]);
tran (stream_cmd_in_nxt[34], \stream_cmd_in_nxt.guid [29]);
tran (stream_cmd_in_nxt[35], \stream_cmd_in_nxt.guid [30]);
tran (stream_cmd_in_nxt[36], \stream_cmd_in_nxt.guid [31]);
tran (stream_cmd_in_nxt[37], \stream_cmd_in_nxt.guid [32]);
tran (stream_cmd_in_nxt[38], \stream_cmd_in_nxt.guid [33]);
tran (stream_cmd_in_nxt[39], \stream_cmd_in_nxt.guid [34]);
tran (stream_cmd_in_nxt[40], \stream_cmd_in_nxt.guid [35]);
tran (stream_cmd_in_nxt[41], \stream_cmd_in_nxt.guid [36]);
tran (stream_cmd_in_nxt[42], \stream_cmd_in_nxt.guid [37]);
tran (stream_cmd_in_nxt[43], \stream_cmd_in_nxt.guid [38]);
tran (stream_cmd_in_nxt[44], \stream_cmd_in_nxt.guid [39]);
tran (stream_cmd_in_nxt[45], \stream_cmd_in_nxt.guid [40]);
tran (stream_cmd_in_nxt[46], \stream_cmd_in_nxt.guid [41]);
tran (stream_cmd_in_nxt[47], \stream_cmd_in_nxt.guid [42]);
tran (stream_cmd_in_nxt[48], \stream_cmd_in_nxt.guid [43]);
tran (stream_cmd_in_nxt[49], \stream_cmd_in_nxt.guid [44]);
tran (stream_cmd_in_nxt[50], \stream_cmd_in_nxt.guid [45]);
tran (stream_cmd_in_nxt[51], \stream_cmd_in_nxt.guid [46]);
tran (stream_cmd_in_nxt[52], \stream_cmd_in_nxt.guid [47]);
tran (stream_cmd_in_nxt[53], \stream_cmd_in_nxt.guid [48]);
tran (stream_cmd_in_nxt[54], \stream_cmd_in_nxt.guid [49]);
tran (stream_cmd_in_nxt[55], \stream_cmd_in_nxt.guid [50]);
tran (stream_cmd_in_nxt[56], \stream_cmd_in_nxt.guid [51]);
tran (stream_cmd_in_nxt[57], \stream_cmd_in_nxt.guid [52]);
tran (stream_cmd_in_nxt[58], \stream_cmd_in_nxt.guid [53]);
tran (stream_cmd_in_nxt[59], \stream_cmd_in_nxt.guid [54]);
tran (stream_cmd_in_nxt[60], \stream_cmd_in_nxt.guid [55]);
tran (stream_cmd_in_nxt[61], \stream_cmd_in_nxt.guid [56]);
tran (stream_cmd_in_nxt[62], \stream_cmd_in_nxt.guid [57]);
tran (stream_cmd_in_nxt[63], \stream_cmd_in_nxt.guid [58]);
tran (stream_cmd_in_nxt[64], \stream_cmd_in_nxt.guid [59]);
tran (stream_cmd_in_nxt[65], \stream_cmd_in_nxt.guid [60]);
tran (stream_cmd_in_nxt[66], \stream_cmd_in_nxt.guid [61]);
tran (stream_cmd_in_nxt[67], \stream_cmd_in_nxt.guid [62]);
tran (stream_cmd_in_nxt[68], \stream_cmd_in_nxt.guid [63]);
tran (stream_cmd_in_nxt[69], \stream_cmd_in_nxt.guid [64]);
tran (stream_cmd_in_nxt[70], \stream_cmd_in_nxt.guid [65]);
tran (stream_cmd_in_nxt[71], \stream_cmd_in_nxt.guid [66]);
tran (stream_cmd_in_nxt[72], \stream_cmd_in_nxt.guid [67]);
tran (stream_cmd_in_nxt[73], \stream_cmd_in_nxt.guid [68]);
tran (stream_cmd_in_nxt[74], \stream_cmd_in_nxt.guid [69]);
tran (stream_cmd_in_nxt[75], \stream_cmd_in_nxt.guid [70]);
tran (stream_cmd_in_nxt[76], \stream_cmd_in_nxt.guid [71]);
tran (stream_cmd_in_nxt[77], \stream_cmd_in_nxt.guid [72]);
tran (stream_cmd_in_nxt[78], \stream_cmd_in_nxt.guid [73]);
tran (stream_cmd_in_nxt[79], \stream_cmd_in_nxt.guid [74]);
tran (stream_cmd_in_nxt[80], \stream_cmd_in_nxt.guid [75]);
tran (stream_cmd_in_nxt[81], \stream_cmd_in_nxt.guid [76]);
tran (stream_cmd_in_nxt[82], \stream_cmd_in_nxt.guid [77]);
tran (stream_cmd_in_nxt[83], \stream_cmd_in_nxt.guid [78]);
tran (stream_cmd_in_nxt[84], \stream_cmd_in_nxt.guid [79]);
tran (stream_cmd_in_nxt[85], \stream_cmd_in_nxt.guid [80]);
tran (stream_cmd_in_nxt[86], \stream_cmd_in_nxt.guid [81]);
tran (stream_cmd_in_nxt[87], \stream_cmd_in_nxt.guid [82]);
tran (stream_cmd_in_nxt[88], \stream_cmd_in_nxt.guid [83]);
tran (stream_cmd_in_nxt[89], \stream_cmd_in_nxt.guid [84]);
tran (stream_cmd_in_nxt[90], \stream_cmd_in_nxt.guid [85]);
tran (stream_cmd_in_nxt[91], \stream_cmd_in_nxt.guid [86]);
tran (stream_cmd_in_nxt[92], \stream_cmd_in_nxt.guid [87]);
tran (stream_cmd_in_nxt[93], \stream_cmd_in_nxt.guid [88]);
tran (stream_cmd_in_nxt[94], \stream_cmd_in_nxt.guid [89]);
tran (stream_cmd_in_nxt[95], \stream_cmd_in_nxt.guid [90]);
tran (stream_cmd_in_nxt[96], \stream_cmd_in_nxt.guid [91]);
tran (stream_cmd_in_nxt[97], \stream_cmd_in_nxt.guid [92]);
tran (stream_cmd_in_nxt[98], \stream_cmd_in_nxt.guid [93]);
tran (stream_cmd_in_nxt[99], \stream_cmd_in_nxt.guid [94]);
tran (stream_cmd_in_nxt[100], \stream_cmd_in_nxt.guid [95]);
tran (stream_cmd_in_nxt[101], \stream_cmd_in_nxt.guid [96]);
tran (stream_cmd_in_nxt[102], \stream_cmd_in_nxt.guid [97]);
tran (stream_cmd_in_nxt[103], \stream_cmd_in_nxt.guid [98]);
tran (stream_cmd_in_nxt[104], \stream_cmd_in_nxt.guid [99]);
tran (stream_cmd_in_nxt[105], \stream_cmd_in_nxt.guid [100]);
tran (stream_cmd_in_nxt[106], \stream_cmd_in_nxt.guid [101]);
tran (stream_cmd_in_nxt[107], \stream_cmd_in_nxt.guid [102]);
tran (stream_cmd_in_nxt[108], \stream_cmd_in_nxt.guid [103]);
tran (stream_cmd_in_nxt[109], \stream_cmd_in_nxt.guid [104]);
tran (stream_cmd_in_nxt[110], \stream_cmd_in_nxt.guid [105]);
tran (stream_cmd_in_nxt[111], \stream_cmd_in_nxt.guid [106]);
tran (stream_cmd_in_nxt[112], \stream_cmd_in_nxt.guid [107]);
tran (stream_cmd_in_nxt[113], \stream_cmd_in_nxt.guid [108]);
tran (stream_cmd_in_nxt[114], \stream_cmd_in_nxt.guid [109]);
tran (stream_cmd_in_nxt[115], \stream_cmd_in_nxt.guid [110]);
tran (stream_cmd_in_nxt[116], \stream_cmd_in_nxt.guid [111]);
tran (stream_cmd_in_nxt[117], \stream_cmd_in_nxt.guid [112]);
tran (stream_cmd_in_nxt[118], \stream_cmd_in_nxt.guid [113]);
tran (stream_cmd_in_nxt[119], \stream_cmd_in_nxt.guid [114]);
tran (stream_cmd_in_nxt[120], \stream_cmd_in_nxt.guid [115]);
tran (stream_cmd_in_nxt[121], \stream_cmd_in_nxt.guid [116]);
tran (stream_cmd_in_nxt[122], \stream_cmd_in_nxt.guid [117]);
tran (stream_cmd_in_nxt[123], \stream_cmd_in_nxt.guid [118]);
tran (stream_cmd_in_nxt[124], \stream_cmd_in_nxt.guid [119]);
tran (stream_cmd_in_nxt[125], \stream_cmd_in_nxt.guid [120]);
tran (stream_cmd_in_nxt[126], \stream_cmd_in_nxt.guid [121]);
tran (stream_cmd_in_nxt[127], \stream_cmd_in_nxt.guid [122]);
tran (stream_cmd_in_nxt[128], \stream_cmd_in_nxt.guid [123]);
tran (stream_cmd_in_nxt[129], \stream_cmd_in_nxt.guid [124]);
tran (stream_cmd_in_nxt[130], \stream_cmd_in_nxt.guid [125]);
tran (stream_cmd_in_nxt[131], \stream_cmd_in_nxt.guid [126]);
tran (stream_cmd_in_nxt[132], \stream_cmd_in_nxt.guid [127]);
tran (stream_cmd_in_nxt[133], \stream_cmd_in_nxt.guid [128]);
tran (stream_cmd_in_nxt[134], \stream_cmd_in_nxt.guid [129]);
tran (stream_cmd_in_nxt[135], \stream_cmd_in_nxt.guid [130]);
tran (stream_cmd_in_nxt[136], \stream_cmd_in_nxt.guid [131]);
tran (stream_cmd_in_nxt[137], \stream_cmd_in_nxt.guid [132]);
tran (stream_cmd_in_nxt[138], \stream_cmd_in_nxt.guid [133]);
tran (stream_cmd_in_nxt[139], \stream_cmd_in_nxt.guid [134]);
tran (stream_cmd_in_nxt[140], \stream_cmd_in_nxt.guid [135]);
tran (stream_cmd_in_nxt[141], \stream_cmd_in_nxt.guid [136]);
tran (stream_cmd_in_nxt[142], \stream_cmd_in_nxt.guid [137]);
tran (stream_cmd_in_nxt[143], \stream_cmd_in_nxt.guid [138]);
tran (stream_cmd_in_nxt[144], \stream_cmd_in_nxt.guid [139]);
tran (stream_cmd_in_nxt[145], \stream_cmd_in_nxt.guid [140]);
tran (stream_cmd_in_nxt[146], \stream_cmd_in_nxt.guid [141]);
tran (stream_cmd_in_nxt[147], \stream_cmd_in_nxt.guid [142]);
tran (stream_cmd_in_nxt[148], \stream_cmd_in_nxt.guid [143]);
tran (stream_cmd_in_nxt[149], \stream_cmd_in_nxt.guid [144]);
tran (stream_cmd_in_nxt[150], \stream_cmd_in_nxt.guid [145]);
tran (stream_cmd_in_nxt[151], \stream_cmd_in_nxt.guid [146]);
tran (stream_cmd_in_nxt[152], \stream_cmd_in_nxt.guid [147]);
tran (stream_cmd_in_nxt[153], \stream_cmd_in_nxt.guid [148]);
tran (stream_cmd_in_nxt[154], \stream_cmd_in_nxt.guid [149]);
tran (stream_cmd_in_nxt[155], \stream_cmd_in_nxt.guid [150]);
tran (stream_cmd_in_nxt[156], \stream_cmd_in_nxt.guid [151]);
tran (stream_cmd_in_nxt[157], \stream_cmd_in_nxt.guid [152]);
tran (stream_cmd_in_nxt[158], \stream_cmd_in_nxt.guid [153]);
tran (stream_cmd_in_nxt[159], \stream_cmd_in_nxt.guid [154]);
tran (stream_cmd_in_nxt[160], \stream_cmd_in_nxt.guid [155]);
tran (stream_cmd_in_nxt[161], \stream_cmd_in_nxt.guid [156]);
tran (stream_cmd_in_nxt[162], \stream_cmd_in_nxt.guid [157]);
tran (stream_cmd_in_nxt[163], \stream_cmd_in_nxt.guid [158]);
tran (stream_cmd_in_nxt[164], \stream_cmd_in_nxt.guid [159]);
tran (stream_cmd_in_nxt[165], \stream_cmd_in_nxt.guid [160]);
tran (stream_cmd_in_nxt[166], \stream_cmd_in_nxt.guid [161]);
tran (stream_cmd_in_nxt[167], \stream_cmd_in_nxt.guid [162]);
tran (stream_cmd_in_nxt[168], \stream_cmd_in_nxt.guid [163]);
tran (stream_cmd_in_nxt[169], \stream_cmd_in_nxt.guid [164]);
tran (stream_cmd_in_nxt[170], \stream_cmd_in_nxt.guid [165]);
tran (stream_cmd_in_nxt[171], \stream_cmd_in_nxt.guid [166]);
tran (stream_cmd_in_nxt[172], \stream_cmd_in_nxt.guid [167]);
tran (stream_cmd_in_nxt[173], \stream_cmd_in_nxt.guid [168]);
tran (stream_cmd_in_nxt[174], \stream_cmd_in_nxt.guid [169]);
tran (stream_cmd_in_nxt[175], \stream_cmd_in_nxt.guid [170]);
tran (stream_cmd_in_nxt[176], \stream_cmd_in_nxt.guid [171]);
tran (stream_cmd_in_nxt[177], \stream_cmd_in_nxt.guid [172]);
tran (stream_cmd_in_nxt[178], \stream_cmd_in_nxt.guid [173]);
tran (stream_cmd_in_nxt[179], \stream_cmd_in_nxt.guid [174]);
tran (stream_cmd_in_nxt[180], \stream_cmd_in_nxt.guid [175]);
tran (stream_cmd_in_nxt[181], \stream_cmd_in_nxt.guid [176]);
tran (stream_cmd_in_nxt[182], \stream_cmd_in_nxt.guid [177]);
tran (stream_cmd_in_nxt[183], \stream_cmd_in_nxt.guid [178]);
tran (stream_cmd_in_nxt[184], \stream_cmd_in_nxt.guid [179]);
tran (stream_cmd_in_nxt[185], \stream_cmd_in_nxt.guid [180]);
tran (stream_cmd_in_nxt[186], \stream_cmd_in_nxt.guid [181]);
tran (stream_cmd_in_nxt[187], \stream_cmd_in_nxt.guid [182]);
tran (stream_cmd_in_nxt[188], \stream_cmd_in_nxt.guid [183]);
tran (stream_cmd_in_nxt[189], \stream_cmd_in_nxt.guid [184]);
tran (stream_cmd_in_nxt[190], \stream_cmd_in_nxt.guid [185]);
tran (stream_cmd_in_nxt[191], \stream_cmd_in_nxt.guid [186]);
tran (stream_cmd_in_nxt[192], \stream_cmd_in_nxt.guid [187]);
tran (stream_cmd_in_nxt[193], \stream_cmd_in_nxt.guid [188]);
tran (stream_cmd_in_nxt[194], \stream_cmd_in_nxt.guid [189]);
tran (stream_cmd_in_nxt[195], \stream_cmd_in_nxt.guid [190]);
tran (stream_cmd_in_nxt[196], \stream_cmd_in_nxt.guid [191]);
tran (stream_cmd_in_nxt[197], \stream_cmd_in_nxt.guid [192]);
tran (stream_cmd_in_nxt[198], \stream_cmd_in_nxt.guid [193]);
tran (stream_cmd_in_nxt[199], \stream_cmd_in_nxt.guid [194]);
tran (stream_cmd_in_nxt[200], \stream_cmd_in_nxt.guid [195]);
tran (stream_cmd_in_nxt[201], \stream_cmd_in_nxt.guid [196]);
tran (stream_cmd_in_nxt[202], \stream_cmd_in_nxt.guid [197]);
tran (stream_cmd_in_nxt[203], \stream_cmd_in_nxt.guid [198]);
tran (stream_cmd_in_nxt[204], \stream_cmd_in_nxt.guid [199]);
tran (stream_cmd_in_nxt[205], \stream_cmd_in_nxt.guid [200]);
tran (stream_cmd_in_nxt[206], \stream_cmd_in_nxt.guid [201]);
tran (stream_cmd_in_nxt[207], \stream_cmd_in_nxt.guid [202]);
tran (stream_cmd_in_nxt[208], \stream_cmd_in_nxt.guid [203]);
tran (stream_cmd_in_nxt[209], \stream_cmd_in_nxt.guid [204]);
tran (stream_cmd_in_nxt[210], \stream_cmd_in_nxt.guid [205]);
tran (stream_cmd_in_nxt[211], \stream_cmd_in_nxt.guid [206]);
tran (stream_cmd_in_nxt[212], \stream_cmd_in_nxt.guid [207]);
tran (stream_cmd_in_nxt[213], \stream_cmd_in_nxt.guid [208]);
tran (stream_cmd_in_nxt[214], \stream_cmd_in_nxt.guid [209]);
tran (stream_cmd_in_nxt[215], \stream_cmd_in_nxt.guid [210]);
tran (stream_cmd_in_nxt[216], \stream_cmd_in_nxt.guid [211]);
tran (stream_cmd_in_nxt[217], \stream_cmd_in_nxt.guid [212]);
tran (stream_cmd_in_nxt[218], \stream_cmd_in_nxt.guid [213]);
tran (stream_cmd_in_nxt[219], \stream_cmd_in_nxt.guid [214]);
tran (stream_cmd_in_nxt[220], \stream_cmd_in_nxt.guid [215]);
tran (stream_cmd_in_nxt[221], \stream_cmd_in_nxt.guid [216]);
tran (stream_cmd_in_nxt[222], \stream_cmd_in_nxt.guid [217]);
tran (stream_cmd_in_nxt[223], \stream_cmd_in_nxt.guid [218]);
tran (stream_cmd_in_nxt[224], \stream_cmd_in_nxt.guid [219]);
tran (stream_cmd_in_nxt[225], \stream_cmd_in_nxt.guid [220]);
tran (stream_cmd_in_nxt[226], \stream_cmd_in_nxt.guid [221]);
tran (stream_cmd_in_nxt[227], \stream_cmd_in_nxt.guid [222]);
tran (stream_cmd_in_nxt[228], \stream_cmd_in_nxt.guid [223]);
tran (stream_cmd_in_nxt[229], \stream_cmd_in_nxt.guid [224]);
tran (stream_cmd_in_nxt[230], \stream_cmd_in_nxt.guid [225]);
tran (stream_cmd_in_nxt[231], \stream_cmd_in_nxt.guid [226]);
tran (stream_cmd_in_nxt[232], \stream_cmd_in_nxt.guid [227]);
tran (stream_cmd_in_nxt[233], \stream_cmd_in_nxt.guid [228]);
tran (stream_cmd_in_nxt[234], \stream_cmd_in_nxt.guid [229]);
tran (stream_cmd_in_nxt[235], \stream_cmd_in_nxt.guid [230]);
tran (stream_cmd_in_nxt[236], \stream_cmd_in_nxt.guid [231]);
tran (stream_cmd_in_nxt[237], \stream_cmd_in_nxt.guid [232]);
tran (stream_cmd_in_nxt[238], \stream_cmd_in_nxt.guid [233]);
tran (stream_cmd_in_nxt[239], \stream_cmd_in_nxt.guid [234]);
tran (stream_cmd_in_nxt[240], \stream_cmd_in_nxt.guid [235]);
tran (stream_cmd_in_nxt[241], \stream_cmd_in_nxt.guid [236]);
tran (stream_cmd_in_nxt[242], \stream_cmd_in_nxt.guid [237]);
tran (stream_cmd_in_nxt[243], \stream_cmd_in_nxt.guid [238]);
tran (stream_cmd_in_nxt[244], \stream_cmd_in_nxt.guid [239]);
tran (stream_cmd_in_nxt[245], \stream_cmd_in_nxt.guid [240]);
tran (stream_cmd_in_nxt[246], \stream_cmd_in_nxt.guid [241]);
tran (stream_cmd_in_nxt[247], \stream_cmd_in_nxt.guid [242]);
tran (stream_cmd_in_nxt[248], \stream_cmd_in_nxt.guid [243]);
tran (stream_cmd_in_nxt[249], \stream_cmd_in_nxt.guid [244]);
tran (stream_cmd_in_nxt[250], \stream_cmd_in_nxt.guid [245]);
tran (stream_cmd_in_nxt[251], \stream_cmd_in_nxt.guid [246]);
tran (stream_cmd_in_nxt[252], \stream_cmd_in_nxt.guid [247]);
tran (stream_cmd_in_nxt[253], \stream_cmd_in_nxt.guid [248]);
tran (stream_cmd_in_nxt[254], \stream_cmd_in_nxt.guid [249]);
tran (stream_cmd_in_nxt[255], \stream_cmd_in_nxt.guid [250]);
tran (stream_cmd_in_nxt[256], \stream_cmd_in_nxt.guid [251]);
tran (stream_cmd_in_nxt[257], \stream_cmd_in_nxt.guid [252]);
tran (stream_cmd_in_nxt[258], \stream_cmd_in_nxt.guid [253]);
tran (stream_cmd_in_nxt[259], \stream_cmd_in_nxt.guid [254]);
tran (stream_cmd_in_nxt[260], \stream_cmd_in_nxt.guid [255]);
tran (stream_cmd_in_nxt[261], \stream_cmd_in_nxt.skip [0]);
tran (stream_cmd_in_nxt[262], \stream_cmd_in_nxt.combo_mode [0]);
tran (gcm_dak_cmd_in[0], \gcm_dak_cmd_in.op [0]);
tran (gcm_dak_cmd_in[1], \gcm_dak_cmd_in.op [1]);
tran (gcm_dak_cmd_in[2], \gcm_dak_cmd_in.op [2]);
tran (gcm_dak_cmd_in[3], \gcm_dak_cmd_in.iv [0]);
tran (gcm_dak_cmd_in[4], \gcm_dak_cmd_in.iv [1]);
tran (gcm_dak_cmd_in[5], \gcm_dak_cmd_in.iv [2]);
tran (gcm_dak_cmd_in[6], \gcm_dak_cmd_in.iv [3]);
tran (gcm_dak_cmd_in[7], \gcm_dak_cmd_in.iv [4]);
tran (gcm_dak_cmd_in[8], \gcm_dak_cmd_in.iv [5]);
tran (gcm_dak_cmd_in[9], \gcm_dak_cmd_in.iv [6]);
tran (gcm_dak_cmd_in[10], \gcm_dak_cmd_in.iv [7]);
tran (gcm_dak_cmd_in[11], \gcm_dak_cmd_in.iv [8]);
tran (gcm_dak_cmd_in[12], \gcm_dak_cmd_in.iv [9]);
tran (gcm_dak_cmd_in[13], \gcm_dak_cmd_in.iv [10]);
tran (gcm_dak_cmd_in[14], \gcm_dak_cmd_in.iv [11]);
tran (gcm_dak_cmd_in[15], \gcm_dak_cmd_in.iv [12]);
tran (gcm_dak_cmd_in[16], \gcm_dak_cmd_in.iv [13]);
tran (gcm_dak_cmd_in[17], \gcm_dak_cmd_in.iv [14]);
tran (gcm_dak_cmd_in[18], \gcm_dak_cmd_in.iv [15]);
tran (gcm_dak_cmd_in[19], \gcm_dak_cmd_in.iv [16]);
tran (gcm_dak_cmd_in[20], \gcm_dak_cmd_in.iv [17]);
tran (gcm_dak_cmd_in[21], \gcm_dak_cmd_in.iv [18]);
tran (gcm_dak_cmd_in[22], \gcm_dak_cmd_in.iv [19]);
tran (gcm_dak_cmd_in[23], \gcm_dak_cmd_in.iv [20]);
tran (gcm_dak_cmd_in[24], \gcm_dak_cmd_in.iv [21]);
tran (gcm_dak_cmd_in[25], \gcm_dak_cmd_in.iv [22]);
tran (gcm_dak_cmd_in[26], \gcm_dak_cmd_in.iv [23]);
tran (gcm_dak_cmd_in[27], \gcm_dak_cmd_in.iv [24]);
tran (gcm_dak_cmd_in[28], \gcm_dak_cmd_in.iv [25]);
tran (gcm_dak_cmd_in[29], \gcm_dak_cmd_in.iv [26]);
tran (gcm_dak_cmd_in[30], \gcm_dak_cmd_in.iv [27]);
tran (gcm_dak_cmd_in[31], \gcm_dak_cmd_in.iv [28]);
tran (gcm_dak_cmd_in[32], \gcm_dak_cmd_in.iv [29]);
tran (gcm_dak_cmd_in[33], \gcm_dak_cmd_in.iv [30]);
tran (gcm_dak_cmd_in[34], \gcm_dak_cmd_in.iv [31]);
tran (gcm_dak_cmd_in[35], \gcm_dak_cmd_in.iv [32]);
tran (gcm_dak_cmd_in[36], \gcm_dak_cmd_in.iv [33]);
tran (gcm_dak_cmd_in[37], \gcm_dak_cmd_in.iv [34]);
tran (gcm_dak_cmd_in[38], \gcm_dak_cmd_in.iv [35]);
tran (gcm_dak_cmd_in[39], \gcm_dak_cmd_in.iv [36]);
tran (gcm_dak_cmd_in[40], \gcm_dak_cmd_in.iv [37]);
tran (gcm_dak_cmd_in[41], \gcm_dak_cmd_in.iv [38]);
tran (gcm_dak_cmd_in[42], \gcm_dak_cmd_in.iv [39]);
tran (gcm_dak_cmd_in[43], \gcm_dak_cmd_in.iv [40]);
tran (gcm_dak_cmd_in[44], \gcm_dak_cmd_in.iv [41]);
tran (gcm_dak_cmd_in[45], \gcm_dak_cmd_in.iv [42]);
tran (gcm_dak_cmd_in[46], \gcm_dak_cmd_in.iv [43]);
tran (gcm_dak_cmd_in[47], \gcm_dak_cmd_in.iv [44]);
tran (gcm_dak_cmd_in[48], \gcm_dak_cmd_in.iv [45]);
tran (gcm_dak_cmd_in[49], \gcm_dak_cmd_in.iv [46]);
tran (gcm_dak_cmd_in[50], \gcm_dak_cmd_in.iv [47]);
tran (gcm_dak_cmd_in[51], \gcm_dak_cmd_in.iv [48]);
tran (gcm_dak_cmd_in[52], \gcm_dak_cmd_in.iv [49]);
tran (gcm_dak_cmd_in[53], \gcm_dak_cmd_in.iv [50]);
tran (gcm_dak_cmd_in[54], \gcm_dak_cmd_in.iv [51]);
tran (gcm_dak_cmd_in[55], \gcm_dak_cmd_in.iv [52]);
tran (gcm_dak_cmd_in[56], \gcm_dak_cmd_in.iv [53]);
tran (gcm_dak_cmd_in[57], \gcm_dak_cmd_in.iv [54]);
tran (gcm_dak_cmd_in[58], \gcm_dak_cmd_in.iv [55]);
tran (gcm_dak_cmd_in[59], \gcm_dak_cmd_in.iv [56]);
tran (gcm_dak_cmd_in[60], \gcm_dak_cmd_in.iv [57]);
tran (gcm_dak_cmd_in[61], \gcm_dak_cmd_in.iv [58]);
tran (gcm_dak_cmd_in[62], \gcm_dak_cmd_in.iv [59]);
tran (gcm_dak_cmd_in[63], \gcm_dak_cmd_in.iv [60]);
tran (gcm_dak_cmd_in[64], \gcm_dak_cmd_in.iv [61]);
tran (gcm_dak_cmd_in[65], \gcm_dak_cmd_in.iv [62]);
tran (gcm_dak_cmd_in[66], \gcm_dak_cmd_in.iv [63]);
tran (gcm_dak_cmd_in[67], \gcm_dak_cmd_in.iv [64]);
tran (gcm_dak_cmd_in[68], \gcm_dak_cmd_in.iv [65]);
tran (gcm_dak_cmd_in[69], \gcm_dak_cmd_in.iv [66]);
tran (gcm_dak_cmd_in[70], \gcm_dak_cmd_in.iv [67]);
tran (gcm_dak_cmd_in[71], \gcm_dak_cmd_in.iv [68]);
tran (gcm_dak_cmd_in[72], \gcm_dak_cmd_in.iv [69]);
tran (gcm_dak_cmd_in[73], \gcm_dak_cmd_in.iv [70]);
tran (gcm_dak_cmd_in[74], \gcm_dak_cmd_in.iv [71]);
tran (gcm_dak_cmd_in[75], \gcm_dak_cmd_in.iv [72]);
tran (gcm_dak_cmd_in[76], \gcm_dak_cmd_in.iv [73]);
tran (gcm_dak_cmd_in[77], \gcm_dak_cmd_in.iv [74]);
tran (gcm_dak_cmd_in[78], \gcm_dak_cmd_in.iv [75]);
tran (gcm_dak_cmd_in[79], \gcm_dak_cmd_in.iv [76]);
tran (gcm_dak_cmd_in[80], \gcm_dak_cmd_in.iv [77]);
tran (gcm_dak_cmd_in[81], \gcm_dak_cmd_in.iv [78]);
tran (gcm_dak_cmd_in[82], \gcm_dak_cmd_in.iv [79]);
tran (gcm_dak_cmd_in[83], \gcm_dak_cmd_in.iv [80]);
tran (gcm_dak_cmd_in[84], \gcm_dak_cmd_in.iv [81]);
tran (gcm_dak_cmd_in[85], \gcm_dak_cmd_in.iv [82]);
tran (gcm_dak_cmd_in[86], \gcm_dak_cmd_in.iv [83]);
tran (gcm_dak_cmd_in[87], \gcm_dak_cmd_in.iv [84]);
tran (gcm_dak_cmd_in[88], \gcm_dak_cmd_in.iv [85]);
tran (gcm_dak_cmd_in[89], \gcm_dak_cmd_in.iv [86]);
tran (gcm_dak_cmd_in[90], \gcm_dak_cmd_in.iv [87]);
tran (gcm_dak_cmd_in[91], \gcm_dak_cmd_in.iv [88]);
tran (gcm_dak_cmd_in[92], \gcm_dak_cmd_in.iv [89]);
tran (gcm_dak_cmd_in[93], \gcm_dak_cmd_in.iv [90]);
tran (gcm_dak_cmd_in[94], \gcm_dak_cmd_in.iv [91]);
tran (gcm_dak_cmd_in[95], \gcm_dak_cmd_in.iv [92]);
tran (gcm_dak_cmd_in[96], \gcm_dak_cmd_in.iv [93]);
tran (gcm_dak_cmd_in[97], \gcm_dak_cmd_in.iv [94]);
tran (gcm_dak_cmd_in[98], \gcm_dak_cmd_in.iv [95]);
tran (gcm_dak_cmd_in[99], \gcm_dak_cmd_in.key1 [0]);
tran (gcm_dak_cmd_in[100], \gcm_dak_cmd_in.key1 [1]);
tran (gcm_dak_cmd_in[101], \gcm_dak_cmd_in.key1 [2]);
tran (gcm_dak_cmd_in[102], \gcm_dak_cmd_in.key1 [3]);
tran (gcm_dak_cmd_in[103], \gcm_dak_cmd_in.key1 [4]);
tran (gcm_dak_cmd_in[104], \gcm_dak_cmd_in.key1 [5]);
tran (gcm_dak_cmd_in[105], \gcm_dak_cmd_in.key1 [6]);
tran (gcm_dak_cmd_in[106], \gcm_dak_cmd_in.key1 [7]);
tran (gcm_dak_cmd_in[107], \gcm_dak_cmd_in.key1 [8]);
tran (gcm_dak_cmd_in[108], \gcm_dak_cmd_in.key1 [9]);
tran (gcm_dak_cmd_in[109], \gcm_dak_cmd_in.key1 [10]);
tran (gcm_dak_cmd_in[110], \gcm_dak_cmd_in.key1 [11]);
tran (gcm_dak_cmd_in[111], \gcm_dak_cmd_in.key1 [12]);
tran (gcm_dak_cmd_in[112], \gcm_dak_cmd_in.key1 [13]);
tran (gcm_dak_cmd_in[113], \gcm_dak_cmd_in.key1 [14]);
tran (gcm_dak_cmd_in[114], \gcm_dak_cmd_in.key1 [15]);
tran (gcm_dak_cmd_in[115], \gcm_dak_cmd_in.key1 [16]);
tran (gcm_dak_cmd_in[116], \gcm_dak_cmd_in.key1 [17]);
tran (gcm_dak_cmd_in[117], \gcm_dak_cmd_in.key1 [18]);
tran (gcm_dak_cmd_in[118], \gcm_dak_cmd_in.key1 [19]);
tran (gcm_dak_cmd_in[119], \gcm_dak_cmd_in.key1 [20]);
tran (gcm_dak_cmd_in[120], \gcm_dak_cmd_in.key1 [21]);
tran (gcm_dak_cmd_in[121], \gcm_dak_cmd_in.key1 [22]);
tran (gcm_dak_cmd_in[122], \gcm_dak_cmd_in.key1 [23]);
tran (gcm_dak_cmd_in[123], \gcm_dak_cmd_in.key1 [24]);
tran (gcm_dak_cmd_in[124], \gcm_dak_cmd_in.key1 [25]);
tran (gcm_dak_cmd_in[125], \gcm_dak_cmd_in.key1 [26]);
tran (gcm_dak_cmd_in[126], \gcm_dak_cmd_in.key1 [27]);
tran (gcm_dak_cmd_in[127], \gcm_dak_cmd_in.key1 [28]);
tran (gcm_dak_cmd_in[128], \gcm_dak_cmd_in.key1 [29]);
tran (gcm_dak_cmd_in[129], \gcm_dak_cmd_in.key1 [30]);
tran (gcm_dak_cmd_in[130], \gcm_dak_cmd_in.key1 [31]);
tran (gcm_dak_cmd_in[131], \gcm_dak_cmd_in.key1 [32]);
tran (gcm_dak_cmd_in[132], \gcm_dak_cmd_in.key1 [33]);
tran (gcm_dak_cmd_in[133], \gcm_dak_cmd_in.key1 [34]);
tran (gcm_dak_cmd_in[134], \gcm_dak_cmd_in.key1 [35]);
tran (gcm_dak_cmd_in[135], \gcm_dak_cmd_in.key1 [36]);
tran (gcm_dak_cmd_in[136], \gcm_dak_cmd_in.key1 [37]);
tran (gcm_dak_cmd_in[137], \gcm_dak_cmd_in.key1 [38]);
tran (gcm_dak_cmd_in[138], \gcm_dak_cmd_in.key1 [39]);
tran (gcm_dak_cmd_in[139], \gcm_dak_cmd_in.key1 [40]);
tran (gcm_dak_cmd_in[140], \gcm_dak_cmd_in.key1 [41]);
tran (gcm_dak_cmd_in[141], \gcm_dak_cmd_in.key1 [42]);
tran (gcm_dak_cmd_in[142], \gcm_dak_cmd_in.key1 [43]);
tran (gcm_dak_cmd_in[143], \gcm_dak_cmd_in.key1 [44]);
tran (gcm_dak_cmd_in[144], \gcm_dak_cmd_in.key1 [45]);
tran (gcm_dak_cmd_in[145], \gcm_dak_cmd_in.key1 [46]);
tran (gcm_dak_cmd_in[146], \gcm_dak_cmd_in.key1 [47]);
tran (gcm_dak_cmd_in[147], \gcm_dak_cmd_in.key1 [48]);
tran (gcm_dak_cmd_in[148], \gcm_dak_cmd_in.key1 [49]);
tran (gcm_dak_cmd_in[149], \gcm_dak_cmd_in.key1 [50]);
tran (gcm_dak_cmd_in[150], \gcm_dak_cmd_in.key1 [51]);
tran (gcm_dak_cmd_in[151], \gcm_dak_cmd_in.key1 [52]);
tran (gcm_dak_cmd_in[152], \gcm_dak_cmd_in.key1 [53]);
tran (gcm_dak_cmd_in[153], \gcm_dak_cmd_in.key1 [54]);
tran (gcm_dak_cmd_in[154], \gcm_dak_cmd_in.key1 [55]);
tran (gcm_dak_cmd_in[155], \gcm_dak_cmd_in.key1 [56]);
tran (gcm_dak_cmd_in[156], \gcm_dak_cmd_in.key1 [57]);
tran (gcm_dak_cmd_in[157], \gcm_dak_cmd_in.key1 [58]);
tran (gcm_dak_cmd_in[158], \gcm_dak_cmd_in.key1 [59]);
tran (gcm_dak_cmd_in[159], \gcm_dak_cmd_in.key1 [60]);
tran (gcm_dak_cmd_in[160], \gcm_dak_cmd_in.key1 [61]);
tran (gcm_dak_cmd_in[161], \gcm_dak_cmd_in.key1 [62]);
tran (gcm_dak_cmd_in[162], \gcm_dak_cmd_in.key1 [63]);
tran (gcm_dak_cmd_in[163], \gcm_dak_cmd_in.key1 [64]);
tran (gcm_dak_cmd_in[164], \gcm_dak_cmd_in.key1 [65]);
tran (gcm_dak_cmd_in[165], \gcm_dak_cmd_in.key1 [66]);
tran (gcm_dak_cmd_in[166], \gcm_dak_cmd_in.key1 [67]);
tran (gcm_dak_cmd_in[167], \gcm_dak_cmd_in.key1 [68]);
tran (gcm_dak_cmd_in[168], \gcm_dak_cmd_in.key1 [69]);
tran (gcm_dak_cmd_in[169], \gcm_dak_cmd_in.key1 [70]);
tran (gcm_dak_cmd_in[170], \gcm_dak_cmd_in.key1 [71]);
tran (gcm_dak_cmd_in[171], \gcm_dak_cmd_in.key1 [72]);
tran (gcm_dak_cmd_in[172], \gcm_dak_cmd_in.key1 [73]);
tran (gcm_dak_cmd_in[173], \gcm_dak_cmd_in.key1 [74]);
tran (gcm_dak_cmd_in[174], \gcm_dak_cmd_in.key1 [75]);
tran (gcm_dak_cmd_in[175], \gcm_dak_cmd_in.key1 [76]);
tran (gcm_dak_cmd_in[176], \gcm_dak_cmd_in.key1 [77]);
tran (gcm_dak_cmd_in[177], \gcm_dak_cmd_in.key1 [78]);
tran (gcm_dak_cmd_in[178], \gcm_dak_cmd_in.key1 [79]);
tran (gcm_dak_cmd_in[179], \gcm_dak_cmd_in.key1 [80]);
tran (gcm_dak_cmd_in[180], \gcm_dak_cmd_in.key1 [81]);
tran (gcm_dak_cmd_in[181], \gcm_dak_cmd_in.key1 [82]);
tran (gcm_dak_cmd_in[182], \gcm_dak_cmd_in.key1 [83]);
tran (gcm_dak_cmd_in[183], \gcm_dak_cmd_in.key1 [84]);
tran (gcm_dak_cmd_in[184], \gcm_dak_cmd_in.key1 [85]);
tran (gcm_dak_cmd_in[185], \gcm_dak_cmd_in.key1 [86]);
tran (gcm_dak_cmd_in[186], \gcm_dak_cmd_in.key1 [87]);
tran (gcm_dak_cmd_in[187], \gcm_dak_cmd_in.key1 [88]);
tran (gcm_dak_cmd_in[188], \gcm_dak_cmd_in.key1 [89]);
tran (gcm_dak_cmd_in[189], \gcm_dak_cmd_in.key1 [90]);
tran (gcm_dak_cmd_in[190], \gcm_dak_cmd_in.key1 [91]);
tran (gcm_dak_cmd_in[191], \gcm_dak_cmd_in.key1 [92]);
tran (gcm_dak_cmd_in[192], \gcm_dak_cmd_in.key1 [93]);
tran (gcm_dak_cmd_in[193], \gcm_dak_cmd_in.key1 [94]);
tran (gcm_dak_cmd_in[194], \gcm_dak_cmd_in.key1 [95]);
tran (gcm_dak_cmd_in[195], \gcm_dak_cmd_in.key1 [96]);
tran (gcm_dak_cmd_in[196], \gcm_dak_cmd_in.key1 [97]);
tran (gcm_dak_cmd_in[197], \gcm_dak_cmd_in.key1 [98]);
tran (gcm_dak_cmd_in[198], \gcm_dak_cmd_in.key1 [99]);
tran (gcm_dak_cmd_in[199], \gcm_dak_cmd_in.key1 [100]);
tran (gcm_dak_cmd_in[200], \gcm_dak_cmd_in.key1 [101]);
tran (gcm_dak_cmd_in[201], \gcm_dak_cmd_in.key1 [102]);
tran (gcm_dak_cmd_in[202], \gcm_dak_cmd_in.key1 [103]);
tran (gcm_dak_cmd_in[203], \gcm_dak_cmd_in.key1 [104]);
tran (gcm_dak_cmd_in[204], \gcm_dak_cmd_in.key1 [105]);
tran (gcm_dak_cmd_in[205], \gcm_dak_cmd_in.key1 [106]);
tran (gcm_dak_cmd_in[206], \gcm_dak_cmd_in.key1 [107]);
tran (gcm_dak_cmd_in[207], \gcm_dak_cmd_in.key1 [108]);
tran (gcm_dak_cmd_in[208], \gcm_dak_cmd_in.key1 [109]);
tran (gcm_dak_cmd_in[209], \gcm_dak_cmd_in.key1 [110]);
tran (gcm_dak_cmd_in[210], \gcm_dak_cmd_in.key1 [111]);
tran (gcm_dak_cmd_in[211], \gcm_dak_cmd_in.key1 [112]);
tran (gcm_dak_cmd_in[212], \gcm_dak_cmd_in.key1 [113]);
tran (gcm_dak_cmd_in[213], \gcm_dak_cmd_in.key1 [114]);
tran (gcm_dak_cmd_in[214], \gcm_dak_cmd_in.key1 [115]);
tran (gcm_dak_cmd_in[215], \gcm_dak_cmd_in.key1 [116]);
tran (gcm_dak_cmd_in[216], \gcm_dak_cmd_in.key1 [117]);
tran (gcm_dak_cmd_in[217], \gcm_dak_cmd_in.key1 [118]);
tran (gcm_dak_cmd_in[218], \gcm_dak_cmd_in.key1 [119]);
tran (gcm_dak_cmd_in[219], \gcm_dak_cmd_in.key1 [120]);
tran (gcm_dak_cmd_in[220], \gcm_dak_cmd_in.key1 [121]);
tran (gcm_dak_cmd_in[221], \gcm_dak_cmd_in.key1 [122]);
tran (gcm_dak_cmd_in[222], \gcm_dak_cmd_in.key1 [123]);
tran (gcm_dak_cmd_in[223], \gcm_dak_cmd_in.key1 [124]);
tran (gcm_dak_cmd_in[224], \gcm_dak_cmd_in.key1 [125]);
tran (gcm_dak_cmd_in[225], \gcm_dak_cmd_in.key1 [126]);
tran (gcm_dak_cmd_in[226], \gcm_dak_cmd_in.key1 [127]);
tran (gcm_dak_cmd_in[227], \gcm_dak_cmd_in.key1 [128]);
tran (gcm_dak_cmd_in[228], \gcm_dak_cmd_in.key1 [129]);
tran (gcm_dak_cmd_in[229], \gcm_dak_cmd_in.key1 [130]);
tran (gcm_dak_cmd_in[230], \gcm_dak_cmd_in.key1 [131]);
tran (gcm_dak_cmd_in[231], \gcm_dak_cmd_in.key1 [132]);
tran (gcm_dak_cmd_in[232], \gcm_dak_cmd_in.key1 [133]);
tran (gcm_dak_cmd_in[233], \gcm_dak_cmd_in.key1 [134]);
tran (gcm_dak_cmd_in[234], \gcm_dak_cmd_in.key1 [135]);
tran (gcm_dak_cmd_in[235], \gcm_dak_cmd_in.key1 [136]);
tran (gcm_dak_cmd_in[236], \gcm_dak_cmd_in.key1 [137]);
tran (gcm_dak_cmd_in[237], \gcm_dak_cmd_in.key1 [138]);
tran (gcm_dak_cmd_in[238], \gcm_dak_cmd_in.key1 [139]);
tran (gcm_dak_cmd_in[239], \gcm_dak_cmd_in.key1 [140]);
tran (gcm_dak_cmd_in[240], \gcm_dak_cmd_in.key1 [141]);
tran (gcm_dak_cmd_in[241], \gcm_dak_cmd_in.key1 [142]);
tran (gcm_dak_cmd_in[242], \gcm_dak_cmd_in.key1 [143]);
tran (gcm_dak_cmd_in[243], \gcm_dak_cmd_in.key1 [144]);
tran (gcm_dak_cmd_in[244], \gcm_dak_cmd_in.key1 [145]);
tran (gcm_dak_cmd_in[245], \gcm_dak_cmd_in.key1 [146]);
tran (gcm_dak_cmd_in[246], \gcm_dak_cmd_in.key1 [147]);
tran (gcm_dak_cmd_in[247], \gcm_dak_cmd_in.key1 [148]);
tran (gcm_dak_cmd_in[248], \gcm_dak_cmd_in.key1 [149]);
tran (gcm_dak_cmd_in[249], \gcm_dak_cmd_in.key1 [150]);
tran (gcm_dak_cmd_in[250], \gcm_dak_cmd_in.key1 [151]);
tran (gcm_dak_cmd_in[251], \gcm_dak_cmd_in.key1 [152]);
tran (gcm_dak_cmd_in[252], \gcm_dak_cmd_in.key1 [153]);
tran (gcm_dak_cmd_in[253], \gcm_dak_cmd_in.key1 [154]);
tran (gcm_dak_cmd_in[254], \gcm_dak_cmd_in.key1 [155]);
tran (gcm_dak_cmd_in[255], \gcm_dak_cmd_in.key1 [156]);
tran (gcm_dak_cmd_in[256], \gcm_dak_cmd_in.key1 [157]);
tran (gcm_dak_cmd_in[257], \gcm_dak_cmd_in.key1 [158]);
tran (gcm_dak_cmd_in[258], \gcm_dak_cmd_in.key1 [159]);
tran (gcm_dak_cmd_in[259], \gcm_dak_cmd_in.key1 [160]);
tran (gcm_dak_cmd_in[260], \gcm_dak_cmd_in.key1 [161]);
tran (gcm_dak_cmd_in[261], \gcm_dak_cmd_in.key1 [162]);
tran (gcm_dak_cmd_in[262], \gcm_dak_cmd_in.key1 [163]);
tran (gcm_dak_cmd_in[263], \gcm_dak_cmd_in.key1 [164]);
tran (gcm_dak_cmd_in[264], \gcm_dak_cmd_in.key1 [165]);
tran (gcm_dak_cmd_in[265], \gcm_dak_cmd_in.key1 [166]);
tran (gcm_dak_cmd_in[266], \gcm_dak_cmd_in.key1 [167]);
tran (gcm_dak_cmd_in[267], \gcm_dak_cmd_in.key1 [168]);
tran (gcm_dak_cmd_in[268], \gcm_dak_cmd_in.key1 [169]);
tran (gcm_dak_cmd_in[269], \gcm_dak_cmd_in.key1 [170]);
tran (gcm_dak_cmd_in[270], \gcm_dak_cmd_in.key1 [171]);
tran (gcm_dak_cmd_in[271], \gcm_dak_cmd_in.key1 [172]);
tran (gcm_dak_cmd_in[272], \gcm_dak_cmd_in.key1 [173]);
tran (gcm_dak_cmd_in[273], \gcm_dak_cmd_in.key1 [174]);
tran (gcm_dak_cmd_in[274], \gcm_dak_cmd_in.key1 [175]);
tran (gcm_dak_cmd_in[275], \gcm_dak_cmd_in.key1 [176]);
tran (gcm_dak_cmd_in[276], \gcm_dak_cmd_in.key1 [177]);
tran (gcm_dak_cmd_in[277], \gcm_dak_cmd_in.key1 [178]);
tran (gcm_dak_cmd_in[278], \gcm_dak_cmd_in.key1 [179]);
tran (gcm_dak_cmd_in[279], \gcm_dak_cmd_in.key1 [180]);
tran (gcm_dak_cmd_in[280], \gcm_dak_cmd_in.key1 [181]);
tran (gcm_dak_cmd_in[281], \gcm_dak_cmd_in.key1 [182]);
tran (gcm_dak_cmd_in[282], \gcm_dak_cmd_in.key1 [183]);
tran (gcm_dak_cmd_in[283], \gcm_dak_cmd_in.key1 [184]);
tran (gcm_dak_cmd_in[284], \gcm_dak_cmd_in.key1 [185]);
tran (gcm_dak_cmd_in[285], \gcm_dak_cmd_in.key1 [186]);
tran (gcm_dak_cmd_in[286], \gcm_dak_cmd_in.key1 [187]);
tran (gcm_dak_cmd_in[287], \gcm_dak_cmd_in.key1 [188]);
tran (gcm_dak_cmd_in[288], \gcm_dak_cmd_in.key1 [189]);
tran (gcm_dak_cmd_in[289], \gcm_dak_cmd_in.key1 [190]);
tran (gcm_dak_cmd_in[290], \gcm_dak_cmd_in.key1 [191]);
tran (gcm_dak_cmd_in[291], \gcm_dak_cmd_in.key1 [192]);
tran (gcm_dak_cmd_in[292], \gcm_dak_cmd_in.key1 [193]);
tran (gcm_dak_cmd_in[293], \gcm_dak_cmd_in.key1 [194]);
tran (gcm_dak_cmd_in[294], \gcm_dak_cmd_in.key1 [195]);
tran (gcm_dak_cmd_in[295], \gcm_dak_cmd_in.key1 [196]);
tran (gcm_dak_cmd_in[296], \gcm_dak_cmd_in.key1 [197]);
tran (gcm_dak_cmd_in[297], \gcm_dak_cmd_in.key1 [198]);
tran (gcm_dak_cmd_in[298], \gcm_dak_cmd_in.key1 [199]);
tran (gcm_dak_cmd_in[299], \gcm_dak_cmd_in.key1 [200]);
tran (gcm_dak_cmd_in[300], \gcm_dak_cmd_in.key1 [201]);
tran (gcm_dak_cmd_in[301], \gcm_dak_cmd_in.key1 [202]);
tran (gcm_dak_cmd_in[302], \gcm_dak_cmd_in.key1 [203]);
tran (gcm_dak_cmd_in[303], \gcm_dak_cmd_in.key1 [204]);
tran (gcm_dak_cmd_in[304], \gcm_dak_cmd_in.key1 [205]);
tran (gcm_dak_cmd_in[305], \gcm_dak_cmd_in.key1 [206]);
tran (gcm_dak_cmd_in[306], \gcm_dak_cmd_in.key1 [207]);
tran (gcm_dak_cmd_in[307], \gcm_dak_cmd_in.key1 [208]);
tran (gcm_dak_cmd_in[308], \gcm_dak_cmd_in.key1 [209]);
tran (gcm_dak_cmd_in[309], \gcm_dak_cmd_in.key1 [210]);
tran (gcm_dak_cmd_in[310], \gcm_dak_cmd_in.key1 [211]);
tran (gcm_dak_cmd_in[311], \gcm_dak_cmd_in.key1 [212]);
tran (gcm_dak_cmd_in[312], \gcm_dak_cmd_in.key1 [213]);
tran (gcm_dak_cmd_in[313], \gcm_dak_cmd_in.key1 [214]);
tran (gcm_dak_cmd_in[314], \gcm_dak_cmd_in.key1 [215]);
tran (gcm_dak_cmd_in[315], \gcm_dak_cmd_in.key1 [216]);
tran (gcm_dak_cmd_in[316], \gcm_dak_cmd_in.key1 [217]);
tran (gcm_dak_cmd_in[317], \gcm_dak_cmd_in.key1 [218]);
tran (gcm_dak_cmd_in[318], \gcm_dak_cmd_in.key1 [219]);
tran (gcm_dak_cmd_in[319], \gcm_dak_cmd_in.key1 [220]);
tran (gcm_dak_cmd_in[320], \gcm_dak_cmd_in.key1 [221]);
tran (gcm_dak_cmd_in[321], \gcm_dak_cmd_in.key1 [222]);
tran (gcm_dak_cmd_in[322], \gcm_dak_cmd_in.key1 [223]);
tran (gcm_dak_cmd_in[323], \gcm_dak_cmd_in.key1 [224]);
tran (gcm_dak_cmd_in[324], \gcm_dak_cmd_in.key1 [225]);
tran (gcm_dak_cmd_in[325], \gcm_dak_cmd_in.key1 [226]);
tran (gcm_dak_cmd_in[326], \gcm_dak_cmd_in.key1 [227]);
tran (gcm_dak_cmd_in[327], \gcm_dak_cmd_in.key1 [228]);
tran (gcm_dak_cmd_in[328], \gcm_dak_cmd_in.key1 [229]);
tran (gcm_dak_cmd_in[329], \gcm_dak_cmd_in.key1 [230]);
tran (gcm_dak_cmd_in[330], \gcm_dak_cmd_in.key1 [231]);
tran (gcm_dak_cmd_in[331], \gcm_dak_cmd_in.key1 [232]);
tran (gcm_dak_cmd_in[332], \gcm_dak_cmd_in.key1 [233]);
tran (gcm_dak_cmd_in[333], \gcm_dak_cmd_in.key1 [234]);
tran (gcm_dak_cmd_in[334], \gcm_dak_cmd_in.key1 [235]);
tran (gcm_dak_cmd_in[335], \gcm_dak_cmd_in.key1 [236]);
tran (gcm_dak_cmd_in[336], \gcm_dak_cmd_in.key1 [237]);
tran (gcm_dak_cmd_in[337], \gcm_dak_cmd_in.key1 [238]);
tran (gcm_dak_cmd_in[338], \gcm_dak_cmd_in.key1 [239]);
tran (gcm_dak_cmd_in[339], \gcm_dak_cmd_in.key1 [240]);
tran (gcm_dak_cmd_in[340], \gcm_dak_cmd_in.key1 [241]);
tran (gcm_dak_cmd_in[341], \gcm_dak_cmd_in.key1 [242]);
tran (gcm_dak_cmd_in[342], \gcm_dak_cmd_in.key1 [243]);
tran (gcm_dak_cmd_in[343], \gcm_dak_cmd_in.key1 [244]);
tran (gcm_dak_cmd_in[344], \gcm_dak_cmd_in.key1 [245]);
tran (gcm_dak_cmd_in[345], \gcm_dak_cmd_in.key1 [246]);
tran (gcm_dak_cmd_in[346], \gcm_dak_cmd_in.key1 [247]);
tran (gcm_dak_cmd_in[347], \gcm_dak_cmd_in.key1 [248]);
tran (gcm_dak_cmd_in[348], \gcm_dak_cmd_in.key1 [249]);
tran (gcm_dak_cmd_in[349], \gcm_dak_cmd_in.key1 [250]);
tran (gcm_dak_cmd_in[350], \gcm_dak_cmd_in.key1 [251]);
tran (gcm_dak_cmd_in[351], \gcm_dak_cmd_in.key1 [252]);
tran (gcm_dak_cmd_in[352], \gcm_dak_cmd_in.key1 [253]);
tran (gcm_dak_cmd_in[353], \gcm_dak_cmd_in.key1 [254]);
tran (gcm_dak_cmd_in[354], \gcm_dak_cmd_in.key1 [255]);
tran (gcm_dak_cmd_in[355], \gcm_dak_cmd_in.key0 [0]);
tran (gcm_dak_cmd_in[356], \gcm_dak_cmd_in.key0 [1]);
tran (gcm_dak_cmd_in[357], \gcm_dak_cmd_in.key0 [2]);
tran (gcm_dak_cmd_in[358], \gcm_dak_cmd_in.key0 [3]);
tran (gcm_dak_cmd_in[359], \gcm_dak_cmd_in.key0 [4]);
tran (gcm_dak_cmd_in[360], \gcm_dak_cmd_in.key0 [5]);
tran (gcm_dak_cmd_in[361], \gcm_dak_cmd_in.key0 [6]);
tran (gcm_dak_cmd_in[362], \gcm_dak_cmd_in.key0 [7]);
tran (gcm_dak_cmd_in[363], \gcm_dak_cmd_in.key0 [8]);
tran (gcm_dak_cmd_in[364], \gcm_dak_cmd_in.key0 [9]);
tran (gcm_dak_cmd_in[365], \gcm_dak_cmd_in.key0 [10]);
tran (gcm_dak_cmd_in[366], \gcm_dak_cmd_in.key0 [11]);
tran (gcm_dak_cmd_in[367], \gcm_dak_cmd_in.key0 [12]);
tran (gcm_dak_cmd_in[368], \gcm_dak_cmd_in.key0 [13]);
tran (gcm_dak_cmd_in[369], \gcm_dak_cmd_in.key0 [14]);
tran (gcm_dak_cmd_in[370], \gcm_dak_cmd_in.key0 [15]);
tran (gcm_dak_cmd_in[371], \gcm_dak_cmd_in.key0 [16]);
tran (gcm_dak_cmd_in[372], \gcm_dak_cmd_in.key0 [17]);
tran (gcm_dak_cmd_in[373], \gcm_dak_cmd_in.key0 [18]);
tran (gcm_dak_cmd_in[374], \gcm_dak_cmd_in.key0 [19]);
tran (gcm_dak_cmd_in[375], \gcm_dak_cmd_in.key0 [20]);
tran (gcm_dak_cmd_in[376], \gcm_dak_cmd_in.key0 [21]);
tran (gcm_dak_cmd_in[377], \gcm_dak_cmd_in.key0 [22]);
tran (gcm_dak_cmd_in[378], \gcm_dak_cmd_in.key0 [23]);
tran (gcm_dak_cmd_in[379], \gcm_dak_cmd_in.key0 [24]);
tran (gcm_dak_cmd_in[380], \gcm_dak_cmd_in.key0 [25]);
tran (gcm_dak_cmd_in[381], \gcm_dak_cmd_in.key0 [26]);
tran (gcm_dak_cmd_in[382], \gcm_dak_cmd_in.key0 [27]);
tran (gcm_dak_cmd_in[383], \gcm_dak_cmd_in.key0 [28]);
tran (gcm_dak_cmd_in[384], \gcm_dak_cmd_in.key0 [29]);
tran (gcm_dak_cmd_in[385], \gcm_dak_cmd_in.key0 [30]);
tran (gcm_dak_cmd_in[386], \gcm_dak_cmd_in.key0 [31]);
tran (gcm_dak_cmd_in[387], \gcm_dak_cmd_in.key0 [32]);
tran (gcm_dak_cmd_in[388], \gcm_dak_cmd_in.key0 [33]);
tran (gcm_dak_cmd_in[389], \gcm_dak_cmd_in.key0 [34]);
tran (gcm_dak_cmd_in[390], \gcm_dak_cmd_in.key0 [35]);
tran (gcm_dak_cmd_in[391], \gcm_dak_cmd_in.key0 [36]);
tran (gcm_dak_cmd_in[392], \gcm_dak_cmd_in.key0 [37]);
tran (gcm_dak_cmd_in[393], \gcm_dak_cmd_in.key0 [38]);
tran (gcm_dak_cmd_in[394], \gcm_dak_cmd_in.key0 [39]);
tran (gcm_dak_cmd_in[395], \gcm_dak_cmd_in.key0 [40]);
tran (gcm_dak_cmd_in[396], \gcm_dak_cmd_in.key0 [41]);
tran (gcm_dak_cmd_in[397], \gcm_dak_cmd_in.key0 [42]);
tran (gcm_dak_cmd_in[398], \gcm_dak_cmd_in.key0 [43]);
tran (gcm_dak_cmd_in[399], \gcm_dak_cmd_in.key0 [44]);
tran (gcm_dak_cmd_in[400], \gcm_dak_cmd_in.key0 [45]);
tran (gcm_dak_cmd_in[401], \gcm_dak_cmd_in.key0 [46]);
tran (gcm_dak_cmd_in[402], \gcm_dak_cmd_in.key0 [47]);
tran (gcm_dak_cmd_in[403], \gcm_dak_cmd_in.key0 [48]);
tran (gcm_dak_cmd_in[404], \gcm_dak_cmd_in.key0 [49]);
tran (gcm_dak_cmd_in[405], \gcm_dak_cmd_in.key0 [50]);
tran (gcm_dak_cmd_in[406], \gcm_dak_cmd_in.key0 [51]);
tran (gcm_dak_cmd_in[407], \gcm_dak_cmd_in.key0 [52]);
tran (gcm_dak_cmd_in[408], \gcm_dak_cmd_in.key0 [53]);
tran (gcm_dak_cmd_in[409], \gcm_dak_cmd_in.key0 [54]);
tran (gcm_dak_cmd_in[410], \gcm_dak_cmd_in.key0 [55]);
tran (gcm_dak_cmd_in[411], \gcm_dak_cmd_in.key0 [56]);
tran (gcm_dak_cmd_in[412], \gcm_dak_cmd_in.key0 [57]);
tran (gcm_dak_cmd_in[413], \gcm_dak_cmd_in.key0 [58]);
tran (gcm_dak_cmd_in[414], \gcm_dak_cmd_in.key0 [59]);
tran (gcm_dak_cmd_in[415], \gcm_dak_cmd_in.key0 [60]);
tran (gcm_dak_cmd_in[416], \gcm_dak_cmd_in.key0 [61]);
tran (gcm_dak_cmd_in[417], \gcm_dak_cmd_in.key0 [62]);
tran (gcm_dak_cmd_in[418], \gcm_dak_cmd_in.key0 [63]);
tran (gcm_dak_cmd_in[419], \gcm_dak_cmd_in.key0 [64]);
tran (gcm_dak_cmd_in[420], \gcm_dak_cmd_in.key0 [65]);
tran (gcm_dak_cmd_in[421], \gcm_dak_cmd_in.key0 [66]);
tran (gcm_dak_cmd_in[422], \gcm_dak_cmd_in.key0 [67]);
tran (gcm_dak_cmd_in[423], \gcm_dak_cmd_in.key0 [68]);
tran (gcm_dak_cmd_in[424], \gcm_dak_cmd_in.key0 [69]);
tran (gcm_dak_cmd_in[425], \gcm_dak_cmd_in.key0 [70]);
tran (gcm_dak_cmd_in[426], \gcm_dak_cmd_in.key0 [71]);
tran (gcm_dak_cmd_in[427], \gcm_dak_cmd_in.key0 [72]);
tran (gcm_dak_cmd_in[428], \gcm_dak_cmd_in.key0 [73]);
tran (gcm_dak_cmd_in[429], \gcm_dak_cmd_in.key0 [74]);
tran (gcm_dak_cmd_in[430], \gcm_dak_cmd_in.key0 [75]);
tran (gcm_dak_cmd_in[431], \gcm_dak_cmd_in.key0 [76]);
tran (gcm_dak_cmd_in[432], \gcm_dak_cmd_in.key0 [77]);
tran (gcm_dak_cmd_in[433], \gcm_dak_cmd_in.key0 [78]);
tran (gcm_dak_cmd_in[434], \gcm_dak_cmd_in.key0 [79]);
tran (gcm_dak_cmd_in[435], \gcm_dak_cmd_in.key0 [80]);
tran (gcm_dak_cmd_in[436], \gcm_dak_cmd_in.key0 [81]);
tran (gcm_dak_cmd_in[437], \gcm_dak_cmd_in.key0 [82]);
tran (gcm_dak_cmd_in[438], \gcm_dak_cmd_in.key0 [83]);
tran (gcm_dak_cmd_in[439], \gcm_dak_cmd_in.key0 [84]);
tran (gcm_dak_cmd_in[440], \gcm_dak_cmd_in.key0 [85]);
tran (gcm_dak_cmd_in[441], \gcm_dak_cmd_in.key0 [86]);
tran (gcm_dak_cmd_in[442], \gcm_dak_cmd_in.key0 [87]);
tran (gcm_dak_cmd_in[443], \gcm_dak_cmd_in.key0 [88]);
tran (gcm_dak_cmd_in[444], \gcm_dak_cmd_in.key0 [89]);
tran (gcm_dak_cmd_in[445], \gcm_dak_cmd_in.key0 [90]);
tran (gcm_dak_cmd_in[446], \gcm_dak_cmd_in.key0 [91]);
tran (gcm_dak_cmd_in[447], \gcm_dak_cmd_in.key0 [92]);
tran (gcm_dak_cmd_in[448], \gcm_dak_cmd_in.key0 [93]);
tran (gcm_dak_cmd_in[449], \gcm_dak_cmd_in.key0 [94]);
tran (gcm_dak_cmd_in[450], \gcm_dak_cmd_in.key0 [95]);
tran (gcm_dak_cmd_in[451], \gcm_dak_cmd_in.key0 [96]);
tran (gcm_dak_cmd_in[452], \gcm_dak_cmd_in.key0 [97]);
tran (gcm_dak_cmd_in[453], \gcm_dak_cmd_in.key0 [98]);
tran (gcm_dak_cmd_in[454], \gcm_dak_cmd_in.key0 [99]);
tran (gcm_dak_cmd_in[455], \gcm_dak_cmd_in.key0 [100]);
tran (gcm_dak_cmd_in[456], \gcm_dak_cmd_in.key0 [101]);
tran (gcm_dak_cmd_in[457], \gcm_dak_cmd_in.key0 [102]);
tran (gcm_dak_cmd_in[458], \gcm_dak_cmd_in.key0 [103]);
tran (gcm_dak_cmd_in[459], \gcm_dak_cmd_in.key0 [104]);
tran (gcm_dak_cmd_in[460], \gcm_dak_cmd_in.key0 [105]);
tran (gcm_dak_cmd_in[461], \gcm_dak_cmd_in.key0 [106]);
tran (gcm_dak_cmd_in[462], \gcm_dak_cmd_in.key0 [107]);
tran (gcm_dak_cmd_in[463], \gcm_dak_cmd_in.key0 [108]);
tran (gcm_dak_cmd_in[464], \gcm_dak_cmd_in.key0 [109]);
tran (gcm_dak_cmd_in[465], \gcm_dak_cmd_in.key0 [110]);
tran (gcm_dak_cmd_in[466], \gcm_dak_cmd_in.key0 [111]);
tran (gcm_dak_cmd_in[467], \gcm_dak_cmd_in.key0 [112]);
tran (gcm_dak_cmd_in[468], \gcm_dak_cmd_in.key0 [113]);
tran (gcm_dak_cmd_in[469], \gcm_dak_cmd_in.key0 [114]);
tran (gcm_dak_cmd_in[470], \gcm_dak_cmd_in.key0 [115]);
tran (gcm_dak_cmd_in[471], \gcm_dak_cmd_in.key0 [116]);
tran (gcm_dak_cmd_in[472], \gcm_dak_cmd_in.key0 [117]);
tran (gcm_dak_cmd_in[473], \gcm_dak_cmd_in.key0 [118]);
tran (gcm_dak_cmd_in[474], \gcm_dak_cmd_in.key0 [119]);
tran (gcm_dak_cmd_in[475], \gcm_dak_cmd_in.key0 [120]);
tran (gcm_dak_cmd_in[476], \gcm_dak_cmd_in.key0 [121]);
tran (gcm_dak_cmd_in[477], \gcm_dak_cmd_in.key0 [122]);
tran (gcm_dak_cmd_in[478], \gcm_dak_cmd_in.key0 [123]);
tran (gcm_dak_cmd_in[479], \gcm_dak_cmd_in.key0 [124]);
tran (gcm_dak_cmd_in[480], \gcm_dak_cmd_in.key0 [125]);
tran (gcm_dak_cmd_in[481], \gcm_dak_cmd_in.key0 [126]);
tran (gcm_dak_cmd_in[482], \gcm_dak_cmd_in.key0 [127]);
tran (gcm_dak_cmd_in[483], \gcm_dak_cmd_in.key0 [128]);
tran (gcm_dak_cmd_in[484], \gcm_dak_cmd_in.key0 [129]);
tran (gcm_dak_cmd_in[485], \gcm_dak_cmd_in.key0 [130]);
tran (gcm_dak_cmd_in[486], \gcm_dak_cmd_in.key0 [131]);
tran (gcm_dak_cmd_in[487], \gcm_dak_cmd_in.key0 [132]);
tran (gcm_dak_cmd_in[488], \gcm_dak_cmd_in.key0 [133]);
tran (gcm_dak_cmd_in[489], \gcm_dak_cmd_in.key0 [134]);
tran (gcm_dak_cmd_in[490], \gcm_dak_cmd_in.key0 [135]);
tran (gcm_dak_cmd_in[491], \gcm_dak_cmd_in.key0 [136]);
tran (gcm_dak_cmd_in[492], \gcm_dak_cmd_in.key0 [137]);
tran (gcm_dak_cmd_in[493], \gcm_dak_cmd_in.key0 [138]);
tran (gcm_dak_cmd_in[494], \gcm_dak_cmd_in.key0 [139]);
tran (gcm_dak_cmd_in[495], \gcm_dak_cmd_in.key0 [140]);
tran (gcm_dak_cmd_in[496], \gcm_dak_cmd_in.key0 [141]);
tran (gcm_dak_cmd_in[497], \gcm_dak_cmd_in.key0 [142]);
tran (gcm_dak_cmd_in[498], \gcm_dak_cmd_in.key0 [143]);
tran (gcm_dak_cmd_in[499], \gcm_dak_cmd_in.key0 [144]);
tran (gcm_dak_cmd_in[500], \gcm_dak_cmd_in.key0 [145]);
tran (gcm_dak_cmd_in[501], \gcm_dak_cmd_in.key0 [146]);
tran (gcm_dak_cmd_in[502], \gcm_dak_cmd_in.key0 [147]);
tran (gcm_dak_cmd_in[503], \gcm_dak_cmd_in.key0 [148]);
tran (gcm_dak_cmd_in[504], \gcm_dak_cmd_in.key0 [149]);
tran (gcm_dak_cmd_in[505], \gcm_dak_cmd_in.key0 [150]);
tran (gcm_dak_cmd_in[506], \gcm_dak_cmd_in.key0 [151]);
tran (gcm_dak_cmd_in[507], \gcm_dak_cmd_in.key0 [152]);
tran (gcm_dak_cmd_in[508], \gcm_dak_cmd_in.key0 [153]);
tran (gcm_dak_cmd_in[509], \gcm_dak_cmd_in.key0 [154]);
tran (gcm_dak_cmd_in[510], \gcm_dak_cmd_in.key0 [155]);
tran (gcm_dak_cmd_in[511], \gcm_dak_cmd_in.key0 [156]);
tran (gcm_dak_cmd_in[512], \gcm_dak_cmd_in.key0 [157]);
tran (gcm_dak_cmd_in[513], \gcm_dak_cmd_in.key0 [158]);
tran (gcm_dak_cmd_in[514], \gcm_dak_cmd_in.key0 [159]);
tran (gcm_dak_cmd_in[515], \gcm_dak_cmd_in.key0 [160]);
tran (gcm_dak_cmd_in[516], \gcm_dak_cmd_in.key0 [161]);
tran (gcm_dak_cmd_in[517], \gcm_dak_cmd_in.key0 [162]);
tran (gcm_dak_cmd_in[518], \gcm_dak_cmd_in.key0 [163]);
tran (gcm_dak_cmd_in[519], \gcm_dak_cmd_in.key0 [164]);
tran (gcm_dak_cmd_in[520], \gcm_dak_cmd_in.key0 [165]);
tran (gcm_dak_cmd_in[521], \gcm_dak_cmd_in.key0 [166]);
tran (gcm_dak_cmd_in[522], \gcm_dak_cmd_in.key0 [167]);
tran (gcm_dak_cmd_in[523], \gcm_dak_cmd_in.key0 [168]);
tran (gcm_dak_cmd_in[524], \gcm_dak_cmd_in.key0 [169]);
tran (gcm_dak_cmd_in[525], \gcm_dak_cmd_in.key0 [170]);
tran (gcm_dak_cmd_in[526], \gcm_dak_cmd_in.key0 [171]);
tran (gcm_dak_cmd_in[527], \gcm_dak_cmd_in.key0 [172]);
tran (gcm_dak_cmd_in[528], \gcm_dak_cmd_in.key0 [173]);
tran (gcm_dak_cmd_in[529], \gcm_dak_cmd_in.key0 [174]);
tran (gcm_dak_cmd_in[530], \gcm_dak_cmd_in.key0 [175]);
tran (gcm_dak_cmd_in[531], \gcm_dak_cmd_in.key0 [176]);
tran (gcm_dak_cmd_in[532], \gcm_dak_cmd_in.key0 [177]);
tran (gcm_dak_cmd_in[533], \gcm_dak_cmd_in.key0 [178]);
tran (gcm_dak_cmd_in[534], \gcm_dak_cmd_in.key0 [179]);
tran (gcm_dak_cmd_in[535], \gcm_dak_cmd_in.key0 [180]);
tran (gcm_dak_cmd_in[536], \gcm_dak_cmd_in.key0 [181]);
tran (gcm_dak_cmd_in[537], \gcm_dak_cmd_in.key0 [182]);
tran (gcm_dak_cmd_in[538], \gcm_dak_cmd_in.key0 [183]);
tran (gcm_dak_cmd_in[539], \gcm_dak_cmd_in.key0 [184]);
tran (gcm_dak_cmd_in[540], \gcm_dak_cmd_in.key0 [185]);
tran (gcm_dak_cmd_in[541], \gcm_dak_cmd_in.key0 [186]);
tran (gcm_dak_cmd_in[542], \gcm_dak_cmd_in.key0 [187]);
tran (gcm_dak_cmd_in[543], \gcm_dak_cmd_in.key0 [188]);
tran (gcm_dak_cmd_in[544], \gcm_dak_cmd_in.key0 [189]);
tran (gcm_dak_cmd_in[545], \gcm_dak_cmd_in.key0 [190]);
tran (gcm_dak_cmd_in[546], \gcm_dak_cmd_in.key0 [191]);
tran (gcm_dak_cmd_in[547], \gcm_dak_cmd_in.key0 [192]);
tran (gcm_dak_cmd_in[548], \gcm_dak_cmd_in.key0 [193]);
tran (gcm_dak_cmd_in[549], \gcm_dak_cmd_in.key0 [194]);
tran (gcm_dak_cmd_in[550], \gcm_dak_cmd_in.key0 [195]);
tran (gcm_dak_cmd_in[551], \gcm_dak_cmd_in.key0 [196]);
tran (gcm_dak_cmd_in[552], \gcm_dak_cmd_in.key0 [197]);
tran (gcm_dak_cmd_in[553], \gcm_dak_cmd_in.key0 [198]);
tran (gcm_dak_cmd_in[554], \gcm_dak_cmd_in.key0 [199]);
tran (gcm_dak_cmd_in[555], \gcm_dak_cmd_in.key0 [200]);
tran (gcm_dak_cmd_in[556], \gcm_dak_cmd_in.key0 [201]);
tran (gcm_dak_cmd_in[557], \gcm_dak_cmd_in.key0 [202]);
tran (gcm_dak_cmd_in[558], \gcm_dak_cmd_in.key0 [203]);
tran (gcm_dak_cmd_in[559], \gcm_dak_cmd_in.key0 [204]);
tran (gcm_dak_cmd_in[560], \gcm_dak_cmd_in.key0 [205]);
tran (gcm_dak_cmd_in[561], \gcm_dak_cmd_in.key0 [206]);
tran (gcm_dak_cmd_in[562], \gcm_dak_cmd_in.key0 [207]);
tran (gcm_dak_cmd_in[563], \gcm_dak_cmd_in.key0 [208]);
tran (gcm_dak_cmd_in[564], \gcm_dak_cmd_in.key0 [209]);
tran (gcm_dak_cmd_in[565], \gcm_dak_cmd_in.key0 [210]);
tran (gcm_dak_cmd_in[566], \gcm_dak_cmd_in.key0 [211]);
tran (gcm_dak_cmd_in[567], \gcm_dak_cmd_in.key0 [212]);
tran (gcm_dak_cmd_in[568], \gcm_dak_cmd_in.key0 [213]);
tran (gcm_dak_cmd_in[569], \gcm_dak_cmd_in.key0 [214]);
tran (gcm_dak_cmd_in[570], \gcm_dak_cmd_in.key0 [215]);
tran (gcm_dak_cmd_in[571], \gcm_dak_cmd_in.key0 [216]);
tran (gcm_dak_cmd_in[572], \gcm_dak_cmd_in.key0 [217]);
tran (gcm_dak_cmd_in[573], \gcm_dak_cmd_in.key0 [218]);
tran (gcm_dak_cmd_in[574], \gcm_dak_cmd_in.key0 [219]);
tran (gcm_dak_cmd_in[575], \gcm_dak_cmd_in.key0 [220]);
tran (gcm_dak_cmd_in[576], \gcm_dak_cmd_in.key0 [221]);
tran (gcm_dak_cmd_in[577], \gcm_dak_cmd_in.key0 [222]);
tran (gcm_dak_cmd_in[578], \gcm_dak_cmd_in.key0 [223]);
tran (gcm_dak_cmd_in[579], \gcm_dak_cmd_in.key0 [224]);
tran (gcm_dak_cmd_in[580], \gcm_dak_cmd_in.key0 [225]);
tran (gcm_dak_cmd_in[581], \gcm_dak_cmd_in.key0 [226]);
tran (gcm_dak_cmd_in[582], \gcm_dak_cmd_in.key0 [227]);
tran (gcm_dak_cmd_in[583], \gcm_dak_cmd_in.key0 [228]);
tran (gcm_dak_cmd_in[584], \gcm_dak_cmd_in.key0 [229]);
tran (gcm_dak_cmd_in[585], \gcm_dak_cmd_in.key0 [230]);
tran (gcm_dak_cmd_in[586], \gcm_dak_cmd_in.key0 [231]);
tran (gcm_dak_cmd_in[587], \gcm_dak_cmd_in.key0 [232]);
tran (gcm_dak_cmd_in[588], \gcm_dak_cmd_in.key0 [233]);
tran (gcm_dak_cmd_in[589], \gcm_dak_cmd_in.key0 [234]);
tran (gcm_dak_cmd_in[590], \gcm_dak_cmd_in.key0 [235]);
tran (gcm_dak_cmd_in[591], \gcm_dak_cmd_in.key0 [236]);
tran (gcm_dak_cmd_in[592], \gcm_dak_cmd_in.key0 [237]);
tran (gcm_dak_cmd_in[593], \gcm_dak_cmd_in.key0 [238]);
tran (gcm_dak_cmd_in[594], \gcm_dak_cmd_in.key0 [239]);
tran (gcm_dak_cmd_in[595], \gcm_dak_cmd_in.key0 [240]);
tran (gcm_dak_cmd_in[596], \gcm_dak_cmd_in.key0 [241]);
tran (gcm_dak_cmd_in[597], \gcm_dak_cmd_in.key0 [242]);
tran (gcm_dak_cmd_in[598], \gcm_dak_cmd_in.key0 [243]);
tran (gcm_dak_cmd_in[599], \gcm_dak_cmd_in.key0 [244]);
tran (gcm_dak_cmd_in[600], \gcm_dak_cmd_in.key0 [245]);
tran (gcm_dak_cmd_in[601], \gcm_dak_cmd_in.key0 [246]);
tran (gcm_dak_cmd_in[602], \gcm_dak_cmd_in.key0 [247]);
tran (gcm_dak_cmd_in[603], \gcm_dak_cmd_in.key0 [248]);
tran (gcm_dak_cmd_in[604], \gcm_dak_cmd_in.key0 [249]);
tran (gcm_dak_cmd_in[605], \gcm_dak_cmd_in.key0 [250]);
tran (gcm_dak_cmd_in[606], \gcm_dak_cmd_in.key0 [251]);
tran (gcm_dak_cmd_in[607], \gcm_dak_cmd_in.key0 [252]);
tran (gcm_dak_cmd_in[608], \gcm_dak_cmd_in.key0 [253]);
tran (gcm_dak_cmd_in[609], \gcm_dak_cmd_in.key0 [254]);
tran (gcm_dak_cmd_in[610], \gcm_dak_cmd_in.key0 [255]);
tran (gcm_dek_cmd_in[0], \gcm_dek_cmd_in.op [0]);
tran (gcm_dek_cmd_in[1], \gcm_dek_cmd_in.op [1]);
tran (gcm_dek_cmd_in[2], \gcm_dek_cmd_in.op [2]);
tran (gcm_dek_cmd_in[3], \gcm_dek_cmd_in.iv [0]);
tran (gcm_dek_cmd_in[4], \gcm_dek_cmd_in.iv [1]);
tran (gcm_dek_cmd_in[5], \gcm_dek_cmd_in.iv [2]);
tran (gcm_dek_cmd_in[6], \gcm_dek_cmd_in.iv [3]);
tran (gcm_dek_cmd_in[7], \gcm_dek_cmd_in.iv [4]);
tran (gcm_dek_cmd_in[8], \gcm_dek_cmd_in.iv [5]);
tran (gcm_dek_cmd_in[9], \gcm_dek_cmd_in.iv [6]);
tran (gcm_dek_cmd_in[10], \gcm_dek_cmd_in.iv [7]);
tran (gcm_dek_cmd_in[11], \gcm_dek_cmd_in.iv [8]);
tran (gcm_dek_cmd_in[12], \gcm_dek_cmd_in.iv [9]);
tran (gcm_dek_cmd_in[13], \gcm_dek_cmd_in.iv [10]);
tran (gcm_dek_cmd_in[14], \gcm_dek_cmd_in.iv [11]);
tran (gcm_dek_cmd_in[15], \gcm_dek_cmd_in.iv [12]);
tran (gcm_dek_cmd_in[16], \gcm_dek_cmd_in.iv [13]);
tran (gcm_dek_cmd_in[17], \gcm_dek_cmd_in.iv [14]);
tran (gcm_dek_cmd_in[18], \gcm_dek_cmd_in.iv [15]);
tran (gcm_dek_cmd_in[19], \gcm_dek_cmd_in.iv [16]);
tran (gcm_dek_cmd_in[20], \gcm_dek_cmd_in.iv [17]);
tran (gcm_dek_cmd_in[21], \gcm_dek_cmd_in.iv [18]);
tran (gcm_dek_cmd_in[22], \gcm_dek_cmd_in.iv [19]);
tran (gcm_dek_cmd_in[23], \gcm_dek_cmd_in.iv [20]);
tran (gcm_dek_cmd_in[24], \gcm_dek_cmd_in.iv [21]);
tran (gcm_dek_cmd_in[25], \gcm_dek_cmd_in.iv [22]);
tran (gcm_dek_cmd_in[26], \gcm_dek_cmd_in.iv [23]);
tran (gcm_dek_cmd_in[27], \gcm_dek_cmd_in.iv [24]);
tran (gcm_dek_cmd_in[28], \gcm_dek_cmd_in.iv [25]);
tran (gcm_dek_cmd_in[29], \gcm_dek_cmd_in.iv [26]);
tran (gcm_dek_cmd_in[30], \gcm_dek_cmd_in.iv [27]);
tran (gcm_dek_cmd_in[31], \gcm_dek_cmd_in.iv [28]);
tran (gcm_dek_cmd_in[32], \gcm_dek_cmd_in.iv [29]);
tran (gcm_dek_cmd_in[33], \gcm_dek_cmd_in.iv [30]);
tran (gcm_dek_cmd_in[34], \gcm_dek_cmd_in.iv [31]);
tran (gcm_dek_cmd_in[35], \gcm_dek_cmd_in.iv [32]);
tran (gcm_dek_cmd_in[36], \gcm_dek_cmd_in.iv [33]);
tran (gcm_dek_cmd_in[37], \gcm_dek_cmd_in.iv [34]);
tran (gcm_dek_cmd_in[38], \gcm_dek_cmd_in.iv [35]);
tran (gcm_dek_cmd_in[39], \gcm_dek_cmd_in.iv [36]);
tran (gcm_dek_cmd_in[40], \gcm_dek_cmd_in.iv [37]);
tran (gcm_dek_cmd_in[41], \gcm_dek_cmd_in.iv [38]);
tran (gcm_dek_cmd_in[42], \gcm_dek_cmd_in.iv [39]);
tran (gcm_dek_cmd_in[43], \gcm_dek_cmd_in.iv [40]);
tran (gcm_dek_cmd_in[44], \gcm_dek_cmd_in.iv [41]);
tran (gcm_dek_cmd_in[45], \gcm_dek_cmd_in.iv [42]);
tran (gcm_dek_cmd_in[46], \gcm_dek_cmd_in.iv [43]);
tran (gcm_dek_cmd_in[47], \gcm_dek_cmd_in.iv [44]);
tran (gcm_dek_cmd_in[48], \gcm_dek_cmd_in.iv [45]);
tran (gcm_dek_cmd_in[49], \gcm_dek_cmd_in.iv [46]);
tran (gcm_dek_cmd_in[50], \gcm_dek_cmd_in.iv [47]);
tran (gcm_dek_cmd_in[51], \gcm_dek_cmd_in.iv [48]);
tran (gcm_dek_cmd_in[52], \gcm_dek_cmd_in.iv [49]);
tran (gcm_dek_cmd_in[53], \gcm_dek_cmd_in.iv [50]);
tran (gcm_dek_cmd_in[54], \gcm_dek_cmd_in.iv [51]);
tran (gcm_dek_cmd_in[55], \gcm_dek_cmd_in.iv [52]);
tran (gcm_dek_cmd_in[56], \gcm_dek_cmd_in.iv [53]);
tran (gcm_dek_cmd_in[57], \gcm_dek_cmd_in.iv [54]);
tran (gcm_dek_cmd_in[58], \gcm_dek_cmd_in.iv [55]);
tran (gcm_dek_cmd_in[59], \gcm_dek_cmd_in.iv [56]);
tran (gcm_dek_cmd_in[60], \gcm_dek_cmd_in.iv [57]);
tran (gcm_dek_cmd_in[61], \gcm_dek_cmd_in.iv [58]);
tran (gcm_dek_cmd_in[62], \gcm_dek_cmd_in.iv [59]);
tran (gcm_dek_cmd_in[63], \gcm_dek_cmd_in.iv [60]);
tran (gcm_dek_cmd_in[64], \gcm_dek_cmd_in.iv [61]);
tran (gcm_dek_cmd_in[65], \gcm_dek_cmd_in.iv [62]);
tran (gcm_dek_cmd_in[66], \gcm_dek_cmd_in.iv [63]);
tran (gcm_dek_cmd_in[67], \gcm_dek_cmd_in.iv [64]);
tran (gcm_dek_cmd_in[68], \gcm_dek_cmd_in.iv [65]);
tran (gcm_dek_cmd_in[69], \gcm_dek_cmd_in.iv [66]);
tran (gcm_dek_cmd_in[70], \gcm_dek_cmd_in.iv [67]);
tran (gcm_dek_cmd_in[71], \gcm_dek_cmd_in.iv [68]);
tran (gcm_dek_cmd_in[72], \gcm_dek_cmd_in.iv [69]);
tran (gcm_dek_cmd_in[73], \gcm_dek_cmd_in.iv [70]);
tran (gcm_dek_cmd_in[74], \gcm_dek_cmd_in.iv [71]);
tran (gcm_dek_cmd_in[75], \gcm_dek_cmd_in.iv [72]);
tran (gcm_dek_cmd_in[76], \gcm_dek_cmd_in.iv [73]);
tran (gcm_dek_cmd_in[77], \gcm_dek_cmd_in.iv [74]);
tran (gcm_dek_cmd_in[78], \gcm_dek_cmd_in.iv [75]);
tran (gcm_dek_cmd_in[79], \gcm_dek_cmd_in.iv [76]);
tran (gcm_dek_cmd_in[80], \gcm_dek_cmd_in.iv [77]);
tran (gcm_dek_cmd_in[81], \gcm_dek_cmd_in.iv [78]);
tran (gcm_dek_cmd_in[82], \gcm_dek_cmd_in.iv [79]);
tran (gcm_dek_cmd_in[83], \gcm_dek_cmd_in.iv [80]);
tran (gcm_dek_cmd_in[84], \gcm_dek_cmd_in.iv [81]);
tran (gcm_dek_cmd_in[85], \gcm_dek_cmd_in.iv [82]);
tran (gcm_dek_cmd_in[86], \gcm_dek_cmd_in.iv [83]);
tran (gcm_dek_cmd_in[87], \gcm_dek_cmd_in.iv [84]);
tran (gcm_dek_cmd_in[88], \gcm_dek_cmd_in.iv [85]);
tran (gcm_dek_cmd_in[89], \gcm_dek_cmd_in.iv [86]);
tran (gcm_dek_cmd_in[90], \gcm_dek_cmd_in.iv [87]);
tran (gcm_dek_cmd_in[91], \gcm_dek_cmd_in.iv [88]);
tran (gcm_dek_cmd_in[92], \gcm_dek_cmd_in.iv [89]);
tran (gcm_dek_cmd_in[93], \gcm_dek_cmd_in.iv [90]);
tran (gcm_dek_cmd_in[94], \gcm_dek_cmd_in.iv [91]);
tran (gcm_dek_cmd_in[95], \gcm_dek_cmd_in.iv [92]);
tran (gcm_dek_cmd_in[96], \gcm_dek_cmd_in.iv [93]);
tran (gcm_dek_cmd_in[97], \gcm_dek_cmd_in.iv [94]);
tran (gcm_dek_cmd_in[98], \gcm_dek_cmd_in.iv [95]);
tran (gcm_dek_cmd_in[99], \gcm_dek_cmd_in.key1 [0]);
tran (gcm_dek_cmd_in[100], \gcm_dek_cmd_in.key1 [1]);
tran (gcm_dek_cmd_in[101], \gcm_dek_cmd_in.key1 [2]);
tran (gcm_dek_cmd_in[102], \gcm_dek_cmd_in.key1 [3]);
tran (gcm_dek_cmd_in[103], \gcm_dek_cmd_in.key1 [4]);
tran (gcm_dek_cmd_in[104], \gcm_dek_cmd_in.key1 [5]);
tran (gcm_dek_cmd_in[105], \gcm_dek_cmd_in.key1 [6]);
tran (gcm_dek_cmd_in[106], \gcm_dek_cmd_in.key1 [7]);
tran (gcm_dek_cmd_in[107], \gcm_dek_cmd_in.key1 [8]);
tran (gcm_dek_cmd_in[108], \gcm_dek_cmd_in.key1 [9]);
tran (gcm_dek_cmd_in[109], \gcm_dek_cmd_in.key1 [10]);
tran (gcm_dek_cmd_in[110], \gcm_dek_cmd_in.key1 [11]);
tran (gcm_dek_cmd_in[111], \gcm_dek_cmd_in.key1 [12]);
tran (gcm_dek_cmd_in[112], \gcm_dek_cmd_in.key1 [13]);
tran (gcm_dek_cmd_in[113], \gcm_dek_cmd_in.key1 [14]);
tran (gcm_dek_cmd_in[114], \gcm_dek_cmd_in.key1 [15]);
tran (gcm_dek_cmd_in[115], \gcm_dek_cmd_in.key1 [16]);
tran (gcm_dek_cmd_in[116], \gcm_dek_cmd_in.key1 [17]);
tran (gcm_dek_cmd_in[117], \gcm_dek_cmd_in.key1 [18]);
tran (gcm_dek_cmd_in[118], \gcm_dek_cmd_in.key1 [19]);
tran (gcm_dek_cmd_in[119], \gcm_dek_cmd_in.key1 [20]);
tran (gcm_dek_cmd_in[120], \gcm_dek_cmd_in.key1 [21]);
tran (gcm_dek_cmd_in[121], \gcm_dek_cmd_in.key1 [22]);
tran (gcm_dek_cmd_in[122], \gcm_dek_cmd_in.key1 [23]);
tran (gcm_dek_cmd_in[123], \gcm_dek_cmd_in.key1 [24]);
tran (gcm_dek_cmd_in[124], \gcm_dek_cmd_in.key1 [25]);
tran (gcm_dek_cmd_in[125], \gcm_dek_cmd_in.key1 [26]);
tran (gcm_dek_cmd_in[126], \gcm_dek_cmd_in.key1 [27]);
tran (gcm_dek_cmd_in[127], \gcm_dek_cmd_in.key1 [28]);
tran (gcm_dek_cmd_in[128], \gcm_dek_cmd_in.key1 [29]);
tran (gcm_dek_cmd_in[129], \gcm_dek_cmd_in.key1 [30]);
tran (gcm_dek_cmd_in[130], \gcm_dek_cmd_in.key1 [31]);
tran (gcm_dek_cmd_in[131], \gcm_dek_cmd_in.key1 [32]);
tran (gcm_dek_cmd_in[132], \gcm_dek_cmd_in.key1 [33]);
tran (gcm_dek_cmd_in[133], \gcm_dek_cmd_in.key1 [34]);
tran (gcm_dek_cmd_in[134], \gcm_dek_cmd_in.key1 [35]);
tran (gcm_dek_cmd_in[135], \gcm_dek_cmd_in.key1 [36]);
tran (gcm_dek_cmd_in[136], \gcm_dek_cmd_in.key1 [37]);
tran (gcm_dek_cmd_in[137], \gcm_dek_cmd_in.key1 [38]);
tran (gcm_dek_cmd_in[138], \gcm_dek_cmd_in.key1 [39]);
tran (gcm_dek_cmd_in[139], \gcm_dek_cmd_in.key1 [40]);
tran (gcm_dek_cmd_in[140], \gcm_dek_cmd_in.key1 [41]);
tran (gcm_dek_cmd_in[141], \gcm_dek_cmd_in.key1 [42]);
tran (gcm_dek_cmd_in[142], \gcm_dek_cmd_in.key1 [43]);
tran (gcm_dek_cmd_in[143], \gcm_dek_cmd_in.key1 [44]);
tran (gcm_dek_cmd_in[144], \gcm_dek_cmd_in.key1 [45]);
tran (gcm_dek_cmd_in[145], \gcm_dek_cmd_in.key1 [46]);
tran (gcm_dek_cmd_in[146], \gcm_dek_cmd_in.key1 [47]);
tran (gcm_dek_cmd_in[147], \gcm_dek_cmd_in.key1 [48]);
tran (gcm_dek_cmd_in[148], \gcm_dek_cmd_in.key1 [49]);
tran (gcm_dek_cmd_in[149], \gcm_dek_cmd_in.key1 [50]);
tran (gcm_dek_cmd_in[150], \gcm_dek_cmd_in.key1 [51]);
tran (gcm_dek_cmd_in[151], \gcm_dek_cmd_in.key1 [52]);
tran (gcm_dek_cmd_in[152], \gcm_dek_cmd_in.key1 [53]);
tran (gcm_dek_cmd_in[153], \gcm_dek_cmd_in.key1 [54]);
tran (gcm_dek_cmd_in[154], \gcm_dek_cmd_in.key1 [55]);
tran (gcm_dek_cmd_in[155], \gcm_dek_cmd_in.key1 [56]);
tran (gcm_dek_cmd_in[156], \gcm_dek_cmd_in.key1 [57]);
tran (gcm_dek_cmd_in[157], \gcm_dek_cmd_in.key1 [58]);
tran (gcm_dek_cmd_in[158], \gcm_dek_cmd_in.key1 [59]);
tran (gcm_dek_cmd_in[159], \gcm_dek_cmd_in.key1 [60]);
tran (gcm_dek_cmd_in[160], \gcm_dek_cmd_in.key1 [61]);
tran (gcm_dek_cmd_in[161], \gcm_dek_cmd_in.key1 [62]);
tran (gcm_dek_cmd_in[162], \gcm_dek_cmd_in.key1 [63]);
tran (gcm_dek_cmd_in[163], \gcm_dek_cmd_in.key1 [64]);
tran (gcm_dek_cmd_in[164], \gcm_dek_cmd_in.key1 [65]);
tran (gcm_dek_cmd_in[165], \gcm_dek_cmd_in.key1 [66]);
tran (gcm_dek_cmd_in[166], \gcm_dek_cmd_in.key1 [67]);
tran (gcm_dek_cmd_in[167], \gcm_dek_cmd_in.key1 [68]);
tran (gcm_dek_cmd_in[168], \gcm_dek_cmd_in.key1 [69]);
tran (gcm_dek_cmd_in[169], \gcm_dek_cmd_in.key1 [70]);
tran (gcm_dek_cmd_in[170], \gcm_dek_cmd_in.key1 [71]);
tran (gcm_dek_cmd_in[171], \gcm_dek_cmd_in.key1 [72]);
tran (gcm_dek_cmd_in[172], \gcm_dek_cmd_in.key1 [73]);
tran (gcm_dek_cmd_in[173], \gcm_dek_cmd_in.key1 [74]);
tran (gcm_dek_cmd_in[174], \gcm_dek_cmd_in.key1 [75]);
tran (gcm_dek_cmd_in[175], \gcm_dek_cmd_in.key1 [76]);
tran (gcm_dek_cmd_in[176], \gcm_dek_cmd_in.key1 [77]);
tran (gcm_dek_cmd_in[177], \gcm_dek_cmd_in.key1 [78]);
tran (gcm_dek_cmd_in[178], \gcm_dek_cmd_in.key1 [79]);
tran (gcm_dek_cmd_in[179], \gcm_dek_cmd_in.key1 [80]);
tran (gcm_dek_cmd_in[180], \gcm_dek_cmd_in.key1 [81]);
tran (gcm_dek_cmd_in[181], \gcm_dek_cmd_in.key1 [82]);
tran (gcm_dek_cmd_in[182], \gcm_dek_cmd_in.key1 [83]);
tran (gcm_dek_cmd_in[183], \gcm_dek_cmd_in.key1 [84]);
tran (gcm_dek_cmd_in[184], \gcm_dek_cmd_in.key1 [85]);
tran (gcm_dek_cmd_in[185], \gcm_dek_cmd_in.key1 [86]);
tran (gcm_dek_cmd_in[186], \gcm_dek_cmd_in.key1 [87]);
tran (gcm_dek_cmd_in[187], \gcm_dek_cmd_in.key1 [88]);
tran (gcm_dek_cmd_in[188], \gcm_dek_cmd_in.key1 [89]);
tran (gcm_dek_cmd_in[189], \gcm_dek_cmd_in.key1 [90]);
tran (gcm_dek_cmd_in[190], \gcm_dek_cmd_in.key1 [91]);
tran (gcm_dek_cmd_in[191], \gcm_dek_cmd_in.key1 [92]);
tran (gcm_dek_cmd_in[192], \gcm_dek_cmd_in.key1 [93]);
tran (gcm_dek_cmd_in[193], \gcm_dek_cmd_in.key1 [94]);
tran (gcm_dek_cmd_in[194], \gcm_dek_cmd_in.key1 [95]);
tran (gcm_dek_cmd_in[195], \gcm_dek_cmd_in.key1 [96]);
tran (gcm_dek_cmd_in[196], \gcm_dek_cmd_in.key1 [97]);
tran (gcm_dek_cmd_in[197], \gcm_dek_cmd_in.key1 [98]);
tran (gcm_dek_cmd_in[198], \gcm_dek_cmd_in.key1 [99]);
tran (gcm_dek_cmd_in[199], \gcm_dek_cmd_in.key1 [100]);
tran (gcm_dek_cmd_in[200], \gcm_dek_cmd_in.key1 [101]);
tran (gcm_dek_cmd_in[201], \gcm_dek_cmd_in.key1 [102]);
tran (gcm_dek_cmd_in[202], \gcm_dek_cmd_in.key1 [103]);
tran (gcm_dek_cmd_in[203], \gcm_dek_cmd_in.key1 [104]);
tran (gcm_dek_cmd_in[204], \gcm_dek_cmd_in.key1 [105]);
tran (gcm_dek_cmd_in[205], \gcm_dek_cmd_in.key1 [106]);
tran (gcm_dek_cmd_in[206], \gcm_dek_cmd_in.key1 [107]);
tran (gcm_dek_cmd_in[207], \gcm_dek_cmd_in.key1 [108]);
tran (gcm_dek_cmd_in[208], \gcm_dek_cmd_in.key1 [109]);
tran (gcm_dek_cmd_in[209], \gcm_dek_cmd_in.key1 [110]);
tran (gcm_dek_cmd_in[210], \gcm_dek_cmd_in.key1 [111]);
tran (gcm_dek_cmd_in[211], \gcm_dek_cmd_in.key1 [112]);
tran (gcm_dek_cmd_in[212], \gcm_dek_cmd_in.key1 [113]);
tran (gcm_dek_cmd_in[213], \gcm_dek_cmd_in.key1 [114]);
tran (gcm_dek_cmd_in[214], \gcm_dek_cmd_in.key1 [115]);
tran (gcm_dek_cmd_in[215], \gcm_dek_cmd_in.key1 [116]);
tran (gcm_dek_cmd_in[216], \gcm_dek_cmd_in.key1 [117]);
tran (gcm_dek_cmd_in[217], \gcm_dek_cmd_in.key1 [118]);
tran (gcm_dek_cmd_in[218], \gcm_dek_cmd_in.key1 [119]);
tran (gcm_dek_cmd_in[219], \gcm_dek_cmd_in.key1 [120]);
tran (gcm_dek_cmd_in[220], \gcm_dek_cmd_in.key1 [121]);
tran (gcm_dek_cmd_in[221], \gcm_dek_cmd_in.key1 [122]);
tran (gcm_dek_cmd_in[222], \gcm_dek_cmd_in.key1 [123]);
tran (gcm_dek_cmd_in[223], \gcm_dek_cmd_in.key1 [124]);
tran (gcm_dek_cmd_in[224], \gcm_dek_cmd_in.key1 [125]);
tran (gcm_dek_cmd_in[225], \gcm_dek_cmd_in.key1 [126]);
tran (gcm_dek_cmd_in[226], \gcm_dek_cmd_in.key1 [127]);
tran (gcm_dek_cmd_in[227], \gcm_dek_cmd_in.key1 [128]);
tran (gcm_dek_cmd_in[228], \gcm_dek_cmd_in.key1 [129]);
tran (gcm_dek_cmd_in[229], \gcm_dek_cmd_in.key1 [130]);
tran (gcm_dek_cmd_in[230], \gcm_dek_cmd_in.key1 [131]);
tran (gcm_dek_cmd_in[231], \gcm_dek_cmd_in.key1 [132]);
tran (gcm_dek_cmd_in[232], \gcm_dek_cmd_in.key1 [133]);
tran (gcm_dek_cmd_in[233], \gcm_dek_cmd_in.key1 [134]);
tran (gcm_dek_cmd_in[234], \gcm_dek_cmd_in.key1 [135]);
tran (gcm_dek_cmd_in[235], \gcm_dek_cmd_in.key1 [136]);
tran (gcm_dek_cmd_in[236], \gcm_dek_cmd_in.key1 [137]);
tran (gcm_dek_cmd_in[237], \gcm_dek_cmd_in.key1 [138]);
tran (gcm_dek_cmd_in[238], \gcm_dek_cmd_in.key1 [139]);
tran (gcm_dek_cmd_in[239], \gcm_dek_cmd_in.key1 [140]);
tran (gcm_dek_cmd_in[240], \gcm_dek_cmd_in.key1 [141]);
tran (gcm_dek_cmd_in[241], \gcm_dek_cmd_in.key1 [142]);
tran (gcm_dek_cmd_in[242], \gcm_dek_cmd_in.key1 [143]);
tran (gcm_dek_cmd_in[243], \gcm_dek_cmd_in.key1 [144]);
tran (gcm_dek_cmd_in[244], \gcm_dek_cmd_in.key1 [145]);
tran (gcm_dek_cmd_in[245], \gcm_dek_cmd_in.key1 [146]);
tran (gcm_dek_cmd_in[246], \gcm_dek_cmd_in.key1 [147]);
tran (gcm_dek_cmd_in[247], \gcm_dek_cmd_in.key1 [148]);
tran (gcm_dek_cmd_in[248], \gcm_dek_cmd_in.key1 [149]);
tran (gcm_dek_cmd_in[249], \gcm_dek_cmd_in.key1 [150]);
tran (gcm_dek_cmd_in[250], \gcm_dek_cmd_in.key1 [151]);
tran (gcm_dek_cmd_in[251], \gcm_dek_cmd_in.key1 [152]);
tran (gcm_dek_cmd_in[252], \gcm_dek_cmd_in.key1 [153]);
tran (gcm_dek_cmd_in[253], \gcm_dek_cmd_in.key1 [154]);
tran (gcm_dek_cmd_in[254], \gcm_dek_cmd_in.key1 [155]);
tran (gcm_dek_cmd_in[255], \gcm_dek_cmd_in.key1 [156]);
tran (gcm_dek_cmd_in[256], \gcm_dek_cmd_in.key1 [157]);
tran (gcm_dek_cmd_in[257], \gcm_dek_cmd_in.key1 [158]);
tran (gcm_dek_cmd_in[258], \gcm_dek_cmd_in.key1 [159]);
tran (gcm_dek_cmd_in[259], \gcm_dek_cmd_in.key1 [160]);
tran (gcm_dek_cmd_in[260], \gcm_dek_cmd_in.key1 [161]);
tran (gcm_dek_cmd_in[261], \gcm_dek_cmd_in.key1 [162]);
tran (gcm_dek_cmd_in[262], \gcm_dek_cmd_in.key1 [163]);
tran (gcm_dek_cmd_in[263], \gcm_dek_cmd_in.key1 [164]);
tran (gcm_dek_cmd_in[264], \gcm_dek_cmd_in.key1 [165]);
tran (gcm_dek_cmd_in[265], \gcm_dek_cmd_in.key1 [166]);
tran (gcm_dek_cmd_in[266], \gcm_dek_cmd_in.key1 [167]);
tran (gcm_dek_cmd_in[267], \gcm_dek_cmd_in.key1 [168]);
tran (gcm_dek_cmd_in[268], \gcm_dek_cmd_in.key1 [169]);
tran (gcm_dek_cmd_in[269], \gcm_dek_cmd_in.key1 [170]);
tran (gcm_dek_cmd_in[270], \gcm_dek_cmd_in.key1 [171]);
tran (gcm_dek_cmd_in[271], \gcm_dek_cmd_in.key1 [172]);
tran (gcm_dek_cmd_in[272], \gcm_dek_cmd_in.key1 [173]);
tran (gcm_dek_cmd_in[273], \gcm_dek_cmd_in.key1 [174]);
tran (gcm_dek_cmd_in[274], \gcm_dek_cmd_in.key1 [175]);
tran (gcm_dek_cmd_in[275], \gcm_dek_cmd_in.key1 [176]);
tran (gcm_dek_cmd_in[276], \gcm_dek_cmd_in.key1 [177]);
tran (gcm_dek_cmd_in[277], \gcm_dek_cmd_in.key1 [178]);
tran (gcm_dek_cmd_in[278], \gcm_dek_cmd_in.key1 [179]);
tran (gcm_dek_cmd_in[279], \gcm_dek_cmd_in.key1 [180]);
tran (gcm_dek_cmd_in[280], \gcm_dek_cmd_in.key1 [181]);
tran (gcm_dek_cmd_in[281], \gcm_dek_cmd_in.key1 [182]);
tran (gcm_dek_cmd_in[282], \gcm_dek_cmd_in.key1 [183]);
tran (gcm_dek_cmd_in[283], \gcm_dek_cmd_in.key1 [184]);
tran (gcm_dek_cmd_in[284], \gcm_dek_cmd_in.key1 [185]);
tran (gcm_dek_cmd_in[285], \gcm_dek_cmd_in.key1 [186]);
tran (gcm_dek_cmd_in[286], \gcm_dek_cmd_in.key1 [187]);
tran (gcm_dek_cmd_in[287], \gcm_dek_cmd_in.key1 [188]);
tran (gcm_dek_cmd_in[288], \gcm_dek_cmd_in.key1 [189]);
tran (gcm_dek_cmd_in[289], \gcm_dek_cmd_in.key1 [190]);
tran (gcm_dek_cmd_in[290], \gcm_dek_cmd_in.key1 [191]);
tran (gcm_dek_cmd_in[291], \gcm_dek_cmd_in.key1 [192]);
tran (gcm_dek_cmd_in[292], \gcm_dek_cmd_in.key1 [193]);
tran (gcm_dek_cmd_in[293], \gcm_dek_cmd_in.key1 [194]);
tran (gcm_dek_cmd_in[294], \gcm_dek_cmd_in.key1 [195]);
tran (gcm_dek_cmd_in[295], \gcm_dek_cmd_in.key1 [196]);
tran (gcm_dek_cmd_in[296], \gcm_dek_cmd_in.key1 [197]);
tran (gcm_dek_cmd_in[297], \gcm_dek_cmd_in.key1 [198]);
tran (gcm_dek_cmd_in[298], \gcm_dek_cmd_in.key1 [199]);
tran (gcm_dek_cmd_in[299], \gcm_dek_cmd_in.key1 [200]);
tran (gcm_dek_cmd_in[300], \gcm_dek_cmd_in.key1 [201]);
tran (gcm_dek_cmd_in[301], \gcm_dek_cmd_in.key1 [202]);
tran (gcm_dek_cmd_in[302], \gcm_dek_cmd_in.key1 [203]);
tran (gcm_dek_cmd_in[303], \gcm_dek_cmd_in.key1 [204]);
tran (gcm_dek_cmd_in[304], \gcm_dek_cmd_in.key1 [205]);
tran (gcm_dek_cmd_in[305], \gcm_dek_cmd_in.key1 [206]);
tran (gcm_dek_cmd_in[306], \gcm_dek_cmd_in.key1 [207]);
tran (gcm_dek_cmd_in[307], \gcm_dek_cmd_in.key1 [208]);
tran (gcm_dek_cmd_in[308], \gcm_dek_cmd_in.key1 [209]);
tran (gcm_dek_cmd_in[309], \gcm_dek_cmd_in.key1 [210]);
tran (gcm_dek_cmd_in[310], \gcm_dek_cmd_in.key1 [211]);
tran (gcm_dek_cmd_in[311], \gcm_dek_cmd_in.key1 [212]);
tran (gcm_dek_cmd_in[312], \gcm_dek_cmd_in.key1 [213]);
tran (gcm_dek_cmd_in[313], \gcm_dek_cmd_in.key1 [214]);
tran (gcm_dek_cmd_in[314], \gcm_dek_cmd_in.key1 [215]);
tran (gcm_dek_cmd_in[315], \gcm_dek_cmd_in.key1 [216]);
tran (gcm_dek_cmd_in[316], \gcm_dek_cmd_in.key1 [217]);
tran (gcm_dek_cmd_in[317], \gcm_dek_cmd_in.key1 [218]);
tran (gcm_dek_cmd_in[318], \gcm_dek_cmd_in.key1 [219]);
tran (gcm_dek_cmd_in[319], \gcm_dek_cmd_in.key1 [220]);
tran (gcm_dek_cmd_in[320], \gcm_dek_cmd_in.key1 [221]);
tran (gcm_dek_cmd_in[321], \gcm_dek_cmd_in.key1 [222]);
tran (gcm_dek_cmd_in[322], \gcm_dek_cmd_in.key1 [223]);
tran (gcm_dek_cmd_in[323], \gcm_dek_cmd_in.key1 [224]);
tran (gcm_dek_cmd_in[324], \gcm_dek_cmd_in.key1 [225]);
tran (gcm_dek_cmd_in[325], \gcm_dek_cmd_in.key1 [226]);
tran (gcm_dek_cmd_in[326], \gcm_dek_cmd_in.key1 [227]);
tran (gcm_dek_cmd_in[327], \gcm_dek_cmd_in.key1 [228]);
tran (gcm_dek_cmd_in[328], \gcm_dek_cmd_in.key1 [229]);
tran (gcm_dek_cmd_in[329], \gcm_dek_cmd_in.key1 [230]);
tran (gcm_dek_cmd_in[330], \gcm_dek_cmd_in.key1 [231]);
tran (gcm_dek_cmd_in[331], \gcm_dek_cmd_in.key1 [232]);
tran (gcm_dek_cmd_in[332], \gcm_dek_cmd_in.key1 [233]);
tran (gcm_dek_cmd_in[333], \gcm_dek_cmd_in.key1 [234]);
tran (gcm_dek_cmd_in[334], \gcm_dek_cmd_in.key1 [235]);
tran (gcm_dek_cmd_in[335], \gcm_dek_cmd_in.key1 [236]);
tran (gcm_dek_cmd_in[336], \gcm_dek_cmd_in.key1 [237]);
tran (gcm_dek_cmd_in[337], \gcm_dek_cmd_in.key1 [238]);
tran (gcm_dek_cmd_in[338], \gcm_dek_cmd_in.key1 [239]);
tran (gcm_dek_cmd_in[339], \gcm_dek_cmd_in.key1 [240]);
tran (gcm_dek_cmd_in[340], \gcm_dek_cmd_in.key1 [241]);
tran (gcm_dek_cmd_in[341], \gcm_dek_cmd_in.key1 [242]);
tran (gcm_dek_cmd_in[342], \gcm_dek_cmd_in.key1 [243]);
tran (gcm_dek_cmd_in[343], \gcm_dek_cmd_in.key1 [244]);
tran (gcm_dek_cmd_in[344], \gcm_dek_cmd_in.key1 [245]);
tran (gcm_dek_cmd_in[345], \gcm_dek_cmd_in.key1 [246]);
tran (gcm_dek_cmd_in[346], \gcm_dek_cmd_in.key1 [247]);
tran (gcm_dek_cmd_in[347], \gcm_dek_cmd_in.key1 [248]);
tran (gcm_dek_cmd_in[348], \gcm_dek_cmd_in.key1 [249]);
tran (gcm_dek_cmd_in[349], \gcm_dek_cmd_in.key1 [250]);
tran (gcm_dek_cmd_in[350], \gcm_dek_cmd_in.key1 [251]);
tran (gcm_dek_cmd_in[351], \gcm_dek_cmd_in.key1 [252]);
tran (gcm_dek_cmd_in[352], \gcm_dek_cmd_in.key1 [253]);
tran (gcm_dek_cmd_in[353], \gcm_dek_cmd_in.key1 [254]);
tran (gcm_dek_cmd_in[354], \gcm_dek_cmd_in.key1 [255]);
tran (gcm_dek_cmd_in[355], \gcm_dek_cmd_in.key0 [0]);
tran (gcm_dek_cmd_in[356], \gcm_dek_cmd_in.key0 [1]);
tran (gcm_dek_cmd_in[357], \gcm_dek_cmd_in.key0 [2]);
tran (gcm_dek_cmd_in[358], \gcm_dek_cmd_in.key0 [3]);
tran (gcm_dek_cmd_in[359], \gcm_dek_cmd_in.key0 [4]);
tran (gcm_dek_cmd_in[360], \gcm_dek_cmd_in.key0 [5]);
tran (gcm_dek_cmd_in[361], \gcm_dek_cmd_in.key0 [6]);
tran (gcm_dek_cmd_in[362], \gcm_dek_cmd_in.key0 [7]);
tran (gcm_dek_cmd_in[363], \gcm_dek_cmd_in.key0 [8]);
tran (gcm_dek_cmd_in[364], \gcm_dek_cmd_in.key0 [9]);
tran (gcm_dek_cmd_in[365], \gcm_dek_cmd_in.key0 [10]);
tran (gcm_dek_cmd_in[366], \gcm_dek_cmd_in.key0 [11]);
tran (gcm_dek_cmd_in[367], \gcm_dek_cmd_in.key0 [12]);
tran (gcm_dek_cmd_in[368], \gcm_dek_cmd_in.key0 [13]);
tran (gcm_dek_cmd_in[369], \gcm_dek_cmd_in.key0 [14]);
tran (gcm_dek_cmd_in[370], \gcm_dek_cmd_in.key0 [15]);
tran (gcm_dek_cmd_in[371], \gcm_dek_cmd_in.key0 [16]);
tran (gcm_dek_cmd_in[372], \gcm_dek_cmd_in.key0 [17]);
tran (gcm_dek_cmd_in[373], \gcm_dek_cmd_in.key0 [18]);
tran (gcm_dek_cmd_in[374], \gcm_dek_cmd_in.key0 [19]);
tran (gcm_dek_cmd_in[375], \gcm_dek_cmd_in.key0 [20]);
tran (gcm_dek_cmd_in[376], \gcm_dek_cmd_in.key0 [21]);
tran (gcm_dek_cmd_in[377], \gcm_dek_cmd_in.key0 [22]);
tran (gcm_dek_cmd_in[378], \gcm_dek_cmd_in.key0 [23]);
tran (gcm_dek_cmd_in[379], \gcm_dek_cmd_in.key0 [24]);
tran (gcm_dek_cmd_in[380], \gcm_dek_cmd_in.key0 [25]);
tran (gcm_dek_cmd_in[381], \gcm_dek_cmd_in.key0 [26]);
tran (gcm_dek_cmd_in[382], \gcm_dek_cmd_in.key0 [27]);
tran (gcm_dek_cmd_in[383], \gcm_dek_cmd_in.key0 [28]);
tran (gcm_dek_cmd_in[384], \gcm_dek_cmd_in.key0 [29]);
tran (gcm_dek_cmd_in[385], \gcm_dek_cmd_in.key0 [30]);
tran (gcm_dek_cmd_in[386], \gcm_dek_cmd_in.key0 [31]);
tran (gcm_dek_cmd_in[387], \gcm_dek_cmd_in.key0 [32]);
tran (gcm_dek_cmd_in[388], \gcm_dek_cmd_in.key0 [33]);
tran (gcm_dek_cmd_in[389], \gcm_dek_cmd_in.key0 [34]);
tran (gcm_dek_cmd_in[390], \gcm_dek_cmd_in.key0 [35]);
tran (gcm_dek_cmd_in[391], \gcm_dek_cmd_in.key0 [36]);
tran (gcm_dek_cmd_in[392], \gcm_dek_cmd_in.key0 [37]);
tran (gcm_dek_cmd_in[393], \gcm_dek_cmd_in.key0 [38]);
tran (gcm_dek_cmd_in[394], \gcm_dek_cmd_in.key0 [39]);
tran (gcm_dek_cmd_in[395], \gcm_dek_cmd_in.key0 [40]);
tran (gcm_dek_cmd_in[396], \gcm_dek_cmd_in.key0 [41]);
tran (gcm_dek_cmd_in[397], \gcm_dek_cmd_in.key0 [42]);
tran (gcm_dek_cmd_in[398], \gcm_dek_cmd_in.key0 [43]);
tran (gcm_dek_cmd_in[399], \gcm_dek_cmd_in.key0 [44]);
tran (gcm_dek_cmd_in[400], \gcm_dek_cmd_in.key0 [45]);
tran (gcm_dek_cmd_in[401], \gcm_dek_cmd_in.key0 [46]);
tran (gcm_dek_cmd_in[402], \gcm_dek_cmd_in.key0 [47]);
tran (gcm_dek_cmd_in[403], \gcm_dek_cmd_in.key0 [48]);
tran (gcm_dek_cmd_in[404], \gcm_dek_cmd_in.key0 [49]);
tran (gcm_dek_cmd_in[405], \gcm_dek_cmd_in.key0 [50]);
tran (gcm_dek_cmd_in[406], \gcm_dek_cmd_in.key0 [51]);
tran (gcm_dek_cmd_in[407], \gcm_dek_cmd_in.key0 [52]);
tran (gcm_dek_cmd_in[408], \gcm_dek_cmd_in.key0 [53]);
tran (gcm_dek_cmd_in[409], \gcm_dek_cmd_in.key0 [54]);
tran (gcm_dek_cmd_in[410], \gcm_dek_cmd_in.key0 [55]);
tran (gcm_dek_cmd_in[411], \gcm_dek_cmd_in.key0 [56]);
tran (gcm_dek_cmd_in[412], \gcm_dek_cmd_in.key0 [57]);
tran (gcm_dek_cmd_in[413], \gcm_dek_cmd_in.key0 [58]);
tran (gcm_dek_cmd_in[414], \gcm_dek_cmd_in.key0 [59]);
tran (gcm_dek_cmd_in[415], \gcm_dek_cmd_in.key0 [60]);
tran (gcm_dek_cmd_in[416], \gcm_dek_cmd_in.key0 [61]);
tran (gcm_dek_cmd_in[417], \gcm_dek_cmd_in.key0 [62]);
tran (gcm_dek_cmd_in[418], \gcm_dek_cmd_in.key0 [63]);
tran (gcm_dek_cmd_in[419], \gcm_dek_cmd_in.key0 [64]);
tran (gcm_dek_cmd_in[420], \gcm_dek_cmd_in.key0 [65]);
tran (gcm_dek_cmd_in[421], \gcm_dek_cmd_in.key0 [66]);
tran (gcm_dek_cmd_in[422], \gcm_dek_cmd_in.key0 [67]);
tran (gcm_dek_cmd_in[423], \gcm_dek_cmd_in.key0 [68]);
tran (gcm_dek_cmd_in[424], \gcm_dek_cmd_in.key0 [69]);
tran (gcm_dek_cmd_in[425], \gcm_dek_cmd_in.key0 [70]);
tran (gcm_dek_cmd_in[426], \gcm_dek_cmd_in.key0 [71]);
tran (gcm_dek_cmd_in[427], \gcm_dek_cmd_in.key0 [72]);
tran (gcm_dek_cmd_in[428], \gcm_dek_cmd_in.key0 [73]);
tran (gcm_dek_cmd_in[429], \gcm_dek_cmd_in.key0 [74]);
tran (gcm_dek_cmd_in[430], \gcm_dek_cmd_in.key0 [75]);
tran (gcm_dek_cmd_in[431], \gcm_dek_cmd_in.key0 [76]);
tran (gcm_dek_cmd_in[432], \gcm_dek_cmd_in.key0 [77]);
tran (gcm_dek_cmd_in[433], \gcm_dek_cmd_in.key0 [78]);
tran (gcm_dek_cmd_in[434], \gcm_dek_cmd_in.key0 [79]);
tran (gcm_dek_cmd_in[435], \gcm_dek_cmd_in.key0 [80]);
tran (gcm_dek_cmd_in[436], \gcm_dek_cmd_in.key0 [81]);
tran (gcm_dek_cmd_in[437], \gcm_dek_cmd_in.key0 [82]);
tran (gcm_dek_cmd_in[438], \gcm_dek_cmd_in.key0 [83]);
tran (gcm_dek_cmd_in[439], \gcm_dek_cmd_in.key0 [84]);
tran (gcm_dek_cmd_in[440], \gcm_dek_cmd_in.key0 [85]);
tran (gcm_dek_cmd_in[441], \gcm_dek_cmd_in.key0 [86]);
tran (gcm_dek_cmd_in[442], \gcm_dek_cmd_in.key0 [87]);
tran (gcm_dek_cmd_in[443], \gcm_dek_cmd_in.key0 [88]);
tran (gcm_dek_cmd_in[444], \gcm_dek_cmd_in.key0 [89]);
tran (gcm_dek_cmd_in[445], \gcm_dek_cmd_in.key0 [90]);
tran (gcm_dek_cmd_in[446], \gcm_dek_cmd_in.key0 [91]);
tran (gcm_dek_cmd_in[447], \gcm_dek_cmd_in.key0 [92]);
tran (gcm_dek_cmd_in[448], \gcm_dek_cmd_in.key0 [93]);
tran (gcm_dek_cmd_in[449], \gcm_dek_cmd_in.key0 [94]);
tran (gcm_dek_cmd_in[450], \gcm_dek_cmd_in.key0 [95]);
tran (gcm_dek_cmd_in[451], \gcm_dek_cmd_in.key0 [96]);
tran (gcm_dek_cmd_in[452], \gcm_dek_cmd_in.key0 [97]);
tran (gcm_dek_cmd_in[453], \gcm_dek_cmd_in.key0 [98]);
tran (gcm_dek_cmd_in[454], \gcm_dek_cmd_in.key0 [99]);
tran (gcm_dek_cmd_in[455], \gcm_dek_cmd_in.key0 [100]);
tran (gcm_dek_cmd_in[456], \gcm_dek_cmd_in.key0 [101]);
tran (gcm_dek_cmd_in[457], \gcm_dek_cmd_in.key0 [102]);
tran (gcm_dek_cmd_in[458], \gcm_dek_cmd_in.key0 [103]);
tran (gcm_dek_cmd_in[459], \gcm_dek_cmd_in.key0 [104]);
tran (gcm_dek_cmd_in[460], \gcm_dek_cmd_in.key0 [105]);
tran (gcm_dek_cmd_in[461], \gcm_dek_cmd_in.key0 [106]);
tran (gcm_dek_cmd_in[462], \gcm_dek_cmd_in.key0 [107]);
tran (gcm_dek_cmd_in[463], \gcm_dek_cmd_in.key0 [108]);
tran (gcm_dek_cmd_in[464], \gcm_dek_cmd_in.key0 [109]);
tran (gcm_dek_cmd_in[465], \gcm_dek_cmd_in.key0 [110]);
tran (gcm_dek_cmd_in[466], \gcm_dek_cmd_in.key0 [111]);
tran (gcm_dek_cmd_in[467], \gcm_dek_cmd_in.key0 [112]);
tran (gcm_dek_cmd_in[468], \gcm_dek_cmd_in.key0 [113]);
tran (gcm_dek_cmd_in[469], \gcm_dek_cmd_in.key0 [114]);
tran (gcm_dek_cmd_in[470], \gcm_dek_cmd_in.key0 [115]);
tran (gcm_dek_cmd_in[471], \gcm_dek_cmd_in.key0 [116]);
tran (gcm_dek_cmd_in[472], \gcm_dek_cmd_in.key0 [117]);
tran (gcm_dek_cmd_in[473], \gcm_dek_cmd_in.key0 [118]);
tran (gcm_dek_cmd_in[474], \gcm_dek_cmd_in.key0 [119]);
tran (gcm_dek_cmd_in[475], \gcm_dek_cmd_in.key0 [120]);
tran (gcm_dek_cmd_in[476], \gcm_dek_cmd_in.key0 [121]);
tran (gcm_dek_cmd_in[477], \gcm_dek_cmd_in.key0 [122]);
tran (gcm_dek_cmd_in[478], \gcm_dek_cmd_in.key0 [123]);
tran (gcm_dek_cmd_in[479], \gcm_dek_cmd_in.key0 [124]);
tran (gcm_dek_cmd_in[480], \gcm_dek_cmd_in.key0 [125]);
tran (gcm_dek_cmd_in[481], \gcm_dek_cmd_in.key0 [126]);
tran (gcm_dek_cmd_in[482], \gcm_dek_cmd_in.key0 [127]);
tran (gcm_dek_cmd_in[483], \gcm_dek_cmd_in.key0 [128]);
tran (gcm_dek_cmd_in[484], \gcm_dek_cmd_in.key0 [129]);
tran (gcm_dek_cmd_in[485], \gcm_dek_cmd_in.key0 [130]);
tran (gcm_dek_cmd_in[486], \gcm_dek_cmd_in.key0 [131]);
tran (gcm_dek_cmd_in[487], \gcm_dek_cmd_in.key0 [132]);
tran (gcm_dek_cmd_in[488], \gcm_dek_cmd_in.key0 [133]);
tran (gcm_dek_cmd_in[489], \gcm_dek_cmd_in.key0 [134]);
tran (gcm_dek_cmd_in[490], \gcm_dek_cmd_in.key0 [135]);
tran (gcm_dek_cmd_in[491], \gcm_dek_cmd_in.key0 [136]);
tran (gcm_dek_cmd_in[492], \gcm_dek_cmd_in.key0 [137]);
tran (gcm_dek_cmd_in[493], \gcm_dek_cmd_in.key0 [138]);
tran (gcm_dek_cmd_in[494], \gcm_dek_cmd_in.key0 [139]);
tran (gcm_dek_cmd_in[495], \gcm_dek_cmd_in.key0 [140]);
tran (gcm_dek_cmd_in[496], \gcm_dek_cmd_in.key0 [141]);
tran (gcm_dek_cmd_in[497], \gcm_dek_cmd_in.key0 [142]);
tran (gcm_dek_cmd_in[498], \gcm_dek_cmd_in.key0 [143]);
tran (gcm_dek_cmd_in[499], \gcm_dek_cmd_in.key0 [144]);
tran (gcm_dek_cmd_in[500], \gcm_dek_cmd_in.key0 [145]);
tran (gcm_dek_cmd_in[501], \gcm_dek_cmd_in.key0 [146]);
tran (gcm_dek_cmd_in[502], \gcm_dek_cmd_in.key0 [147]);
tran (gcm_dek_cmd_in[503], \gcm_dek_cmd_in.key0 [148]);
tran (gcm_dek_cmd_in[504], \gcm_dek_cmd_in.key0 [149]);
tran (gcm_dek_cmd_in[505], \gcm_dek_cmd_in.key0 [150]);
tran (gcm_dek_cmd_in[506], \gcm_dek_cmd_in.key0 [151]);
tran (gcm_dek_cmd_in[507], \gcm_dek_cmd_in.key0 [152]);
tran (gcm_dek_cmd_in[508], \gcm_dek_cmd_in.key0 [153]);
tran (gcm_dek_cmd_in[509], \gcm_dek_cmd_in.key0 [154]);
tran (gcm_dek_cmd_in[510], \gcm_dek_cmd_in.key0 [155]);
tran (gcm_dek_cmd_in[511], \gcm_dek_cmd_in.key0 [156]);
tran (gcm_dek_cmd_in[512], \gcm_dek_cmd_in.key0 [157]);
tran (gcm_dek_cmd_in[513], \gcm_dek_cmd_in.key0 [158]);
tran (gcm_dek_cmd_in[514], \gcm_dek_cmd_in.key0 [159]);
tran (gcm_dek_cmd_in[515], \gcm_dek_cmd_in.key0 [160]);
tran (gcm_dek_cmd_in[516], \gcm_dek_cmd_in.key0 [161]);
tran (gcm_dek_cmd_in[517], \gcm_dek_cmd_in.key0 [162]);
tran (gcm_dek_cmd_in[518], \gcm_dek_cmd_in.key0 [163]);
tran (gcm_dek_cmd_in[519], \gcm_dek_cmd_in.key0 [164]);
tran (gcm_dek_cmd_in[520], \gcm_dek_cmd_in.key0 [165]);
tran (gcm_dek_cmd_in[521], \gcm_dek_cmd_in.key0 [166]);
tran (gcm_dek_cmd_in[522], \gcm_dek_cmd_in.key0 [167]);
tran (gcm_dek_cmd_in[523], \gcm_dek_cmd_in.key0 [168]);
tran (gcm_dek_cmd_in[524], \gcm_dek_cmd_in.key0 [169]);
tran (gcm_dek_cmd_in[525], \gcm_dek_cmd_in.key0 [170]);
tran (gcm_dek_cmd_in[526], \gcm_dek_cmd_in.key0 [171]);
tran (gcm_dek_cmd_in[527], \gcm_dek_cmd_in.key0 [172]);
tran (gcm_dek_cmd_in[528], \gcm_dek_cmd_in.key0 [173]);
tran (gcm_dek_cmd_in[529], \gcm_dek_cmd_in.key0 [174]);
tran (gcm_dek_cmd_in[530], \gcm_dek_cmd_in.key0 [175]);
tran (gcm_dek_cmd_in[531], \gcm_dek_cmd_in.key0 [176]);
tran (gcm_dek_cmd_in[532], \gcm_dek_cmd_in.key0 [177]);
tran (gcm_dek_cmd_in[533], \gcm_dek_cmd_in.key0 [178]);
tran (gcm_dek_cmd_in[534], \gcm_dek_cmd_in.key0 [179]);
tran (gcm_dek_cmd_in[535], \gcm_dek_cmd_in.key0 [180]);
tran (gcm_dek_cmd_in[536], \gcm_dek_cmd_in.key0 [181]);
tran (gcm_dek_cmd_in[537], \gcm_dek_cmd_in.key0 [182]);
tran (gcm_dek_cmd_in[538], \gcm_dek_cmd_in.key0 [183]);
tran (gcm_dek_cmd_in[539], \gcm_dek_cmd_in.key0 [184]);
tran (gcm_dek_cmd_in[540], \gcm_dek_cmd_in.key0 [185]);
tran (gcm_dek_cmd_in[541], \gcm_dek_cmd_in.key0 [186]);
tran (gcm_dek_cmd_in[542], \gcm_dek_cmd_in.key0 [187]);
tran (gcm_dek_cmd_in[543], \gcm_dek_cmd_in.key0 [188]);
tran (gcm_dek_cmd_in[544], \gcm_dek_cmd_in.key0 [189]);
tran (gcm_dek_cmd_in[545], \gcm_dek_cmd_in.key0 [190]);
tran (gcm_dek_cmd_in[546], \gcm_dek_cmd_in.key0 [191]);
tran (gcm_dek_cmd_in[547], \gcm_dek_cmd_in.key0 [192]);
tran (gcm_dek_cmd_in[548], \gcm_dek_cmd_in.key0 [193]);
tran (gcm_dek_cmd_in[549], \gcm_dek_cmd_in.key0 [194]);
tran (gcm_dek_cmd_in[550], \gcm_dek_cmd_in.key0 [195]);
tran (gcm_dek_cmd_in[551], \gcm_dek_cmd_in.key0 [196]);
tran (gcm_dek_cmd_in[552], \gcm_dek_cmd_in.key0 [197]);
tran (gcm_dek_cmd_in[553], \gcm_dek_cmd_in.key0 [198]);
tran (gcm_dek_cmd_in[554], \gcm_dek_cmd_in.key0 [199]);
tran (gcm_dek_cmd_in[555], \gcm_dek_cmd_in.key0 [200]);
tran (gcm_dek_cmd_in[556], \gcm_dek_cmd_in.key0 [201]);
tran (gcm_dek_cmd_in[557], \gcm_dek_cmd_in.key0 [202]);
tran (gcm_dek_cmd_in[558], \gcm_dek_cmd_in.key0 [203]);
tran (gcm_dek_cmd_in[559], \gcm_dek_cmd_in.key0 [204]);
tran (gcm_dek_cmd_in[560], \gcm_dek_cmd_in.key0 [205]);
tran (gcm_dek_cmd_in[561], \gcm_dek_cmd_in.key0 [206]);
tran (gcm_dek_cmd_in[562], \gcm_dek_cmd_in.key0 [207]);
tran (gcm_dek_cmd_in[563], \gcm_dek_cmd_in.key0 [208]);
tran (gcm_dek_cmd_in[564], \gcm_dek_cmd_in.key0 [209]);
tran (gcm_dek_cmd_in[565], \gcm_dek_cmd_in.key0 [210]);
tran (gcm_dek_cmd_in[566], \gcm_dek_cmd_in.key0 [211]);
tran (gcm_dek_cmd_in[567], \gcm_dek_cmd_in.key0 [212]);
tran (gcm_dek_cmd_in[568], \gcm_dek_cmd_in.key0 [213]);
tran (gcm_dek_cmd_in[569], \gcm_dek_cmd_in.key0 [214]);
tran (gcm_dek_cmd_in[570], \gcm_dek_cmd_in.key0 [215]);
tran (gcm_dek_cmd_in[571], \gcm_dek_cmd_in.key0 [216]);
tran (gcm_dek_cmd_in[572], \gcm_dek_cmd_in.key0 [217]);
tran (gcm_dek_cmd_in[573], \gcm_dek_cmd_in.key0 [218]);
tran (gcm_dek_cmd_in[574], \gcm_dek_cmd_in.key0 [219]);
tran (gcm_dek_cmd_in[575], \gcm_dek_cmd_in.key0 [220]);
tran (gcm_dek_cmd_in[576], \gcm_dek_cmd_in.key0 [221]);
tran (gcm_dek_cmd_in[577], \gcm_dek_cmd_in.key0 [222]);
tran (gcm_dek_cmd_in[578], \gcm_dek_cmd_in.key0 [223]);
tran (gcm_dek_cmd_in[579], \gcm_dek_cmd_in.key0 [224]);
tran (gcm_dek_cmd_in[580], \gcm_dek_cmd_in.key0 [225]);
tran (gcm_dek_cmd_in[581], \gcm_dek_cmd_in.key0 [226]);
tran (gcm_dek_cmd_in[582], \gcm_dek_cmd_in.key0 [227]);
tran (gcm_dek_cmd_in[583], \gcm_dek_cmd_in.key0 [228]);
tran (gcm_dek_cmd_in[584], \gcm_dek_cmd_in.key0 [229]);
tran (gcm_dek_cmd_in[585], \gcm_dek_cmd_in.key0 [230]);
tran (gcm_dek_cmd_in[586], \gcm_dek_cmd_in.key0 [231]);
tran (gcm_dek_cmd_in[587], \gcm_dek_cmd_in.key0 [232]);
tran (gcm_dek_cmd_in[588], \gcm_dek_cmd_in.key0 [233]);
tran (gcm_dek_cmd_in[589], \gcm_dek_cmd_in.key0 [234]);
tran (gcm_dek_cmd_in[590], \gcm_dek_cmd_in.key0 [235]);
tran (gcm_dek_cmd_in[591], \gcm_dek_cmd_in.key0 [236]);
tran (gcm_dek_cmd_in[592], \gcm_dek_cmd_in.key0 [237]);
tran (gcm_dek_cmd_in[593], \gcm_dek_cmd_in.key0 [238]);
tran (gcm_dek_cmd_in[594], \gcm_dek_cmd_in.key0 [239]);
tran (gcm_dek_cmd_in[595], \gcm_dek_cmd_in.key0 [240]);
tran (gcm_dek_cmd_in[596], \gcm_dek_cmd_in.key0 [241]);
tran (gcm_dek_cmd_in[597], \gcm_dek_cmd_in.key0 [242]);
tran (gcm_dek_cmd_in[598], \gcm_dek_cmd_in.key0 [243]);
tran (gcm_dek_cmd_in[599], \gcm_dek_cmd_in.key0 [244]);
tran (gcm_dek_cmd_in[600], \gcm_dek_cmd_in.key0 [245]);
tran (gcm_dek_cmd_in[601], \gcm_dek_cmd_in.key0 [246]);
tran (gcm_dek_cmd_in[602], \gcm_dek_cmd_in.key0 [247]);
tran (gcm_dek_cmd_in[603], \gcm_dek_cmd_in.key0 [248]);
tran (gcm_dek_cmd_in[604], \gcm_dek_cmd_in.key0 [249]);
tran (gcm_dek_cmd_in[605], \gcm_dek_cmd_in.key0 [250]);
tran (gcm_dek_cmd_in[606], \gcm_dek_cmd_in.key0 [251]);
tran (gcm_dek_cmd_in[607], \gcm_dek_cmd_in.key0 [252]);
tran (gcm_dek_cmd_in[608], \gcm_dek_cmd_in.key0 [253]);
tran (gcm_dek_cmd_in[609], \gcm_dek_cmd_in.key0 [254]);
tran (gcm_dek_cmd_in[610], \gcm_dek_cmd_in.key0 [255]);
tran (stream_cmd_in[0], \stream_cmd_in.num_iter [0]);
tran (stream_cmd_in[1], \stream_cmd_in.num_iter [1]);
tran (stream_cmd_in[2], \stream_cmd_in.label_index [0]);
tran (stream_cmd_in[3], \stream_cmd_in.label_index [1]);
tran (stream_cmd_in[4], \stream_cmd_in.label_index [2]);
tran (stream_cmd_in[5], \stream_cmd_in.guid [0]);
tran (stream_cmd_in[6], \stream_cmd_in.guid [1]);
tran (stream_cmd_in[7], \stream_cmd_in.guid [2]);
tran (stream_cmd_in[8], \stream_cmd_in.guid [3]);
tran (stream_cmd_in[9], \stream_cmd_in.guid [4]);
tran (stream_cmd_in[10], \stream_cmd_in.guid [5]);
tran (stream_cmd_in[11], \stream_cmd_in.guid [6]);
tran (stream_cmd_in[12], \stream_cmd_in.guid [7]);
tran (stream_cmd_in[13], \stream_cmd_in.guid [8]);
tran (stream_cmd_in[14], \stream_cmd_in.guid [9]);
tran (stream_cmd_in[15], \stream_cmd_in.guid [10]);
tran (stream_cmd_in[16], \stream_cmd_in.guid [11]);
tran (stream_cmd_in[17], \stream_cmd_in.guid [12]);
tran (stream_cmd_in[18], \stream_cmd_in.guid [13]);
tran (stream_cmd_in[19], \stream_cmd_in.guid [14]);
tran (stream_cmd_in[20], \stream_cmd_in.guid [15]);
tran (stream_cmd_in[21], \stream_cmd_in.guid [16]);
tran (stream_cmd_in[22], \stream_cmd_in.guid [17]);
tran (stream_cmd_in[23], \stream_cmd_in.guid [18]);
tran (stream_cmd_in[24], \stream_cmd_in.guid [19]);
tran (stream_cmd_in[25], \stream_cmd_in.guid [20]);
tran (stream_cmd_in[26], \stream_cmd_in.guid [21]);
tran (stream_cmd_in[27], \stream_cmd_in.guid [22]);
tran (stream_cmd_in[28], \stream_cmd_in.guid [23]);
tran (stream_cmd_in[29], \stream_cmd_in.guid [24]);
tran (stream_cmd_in[30], \stream_cmd_in.guid [25]);
tran (stream_cmd_in[31], \stream_cmd_in.guid [26]);
tran (stream_cmd_in[32], \stream_cmd_in.guid [27]);
tran (stream_cmd_in[33], \stream_cmd_in.guid [28]);
tran (stream_cmd_in[34], \stream_cmd_in.guid [29]);
tran (stream_cmd_in[35], \stream_cmd_in.guid [30]);
tran (stream_cmd_in[36], \stream_cmd_in.guid [31]);
tran (stream_cmd_in[37], \stream_cmd_in.guid [32]);
tran (stream_cmd_in[38], \stream_cmd_in.guid [33]);
tran (stream_cmd_in[39], \stream_cmd_in.guid [34]);
tran (stream_cmd_in[40], \stream_cmd_in.guid [35]);
tran (stream_cmd_in[41], \stream_cmd_in.guid [36]);
tran (stream_cmd_in[42], \stream_cmd_in.guid [37]);
tran (stream_cmd_in[43], \stream_cmd_in.guid [38]);
tran (stream_cmd_in[44], \stream_cmd_in.guid [39]);
tran (stream_cmd_in[45], \stream_cmd_in.guid [40]);
tran (stream_cmd_in[46], \stream_cmd_in.guid [41]);
tran (stream_cmd_in[47], \stream_cmd_in.guid [42]);
tran (stream_cmd_in[48], \stream_cmd_in.guid [43]);
tran (stream_cmd_in[49], \stream_cmd_in.guid [44]);
tran (stream_cmd_in[50], \stream_cmd_in.guid [45]);
tran (stream_cmd_in[51], \stream_cmd_in.guid [46]);
tran (stream_cmd_in[52], \stream_cmd_in.guid [47]);
tran (stream_cmd_in[53], \stream_cmd_in.guid [48]);
tran (stream_cmd_in[54], \stream_cmd_in.guid [49]);
tran (stream_cmd_in[55], \stream_cmd_in.guid [50]);
tran (stream_cmd_in[56], \stream_cmd_in.guid [51]);
tran (stream_cmd_in[57], \stream_cmd_in.guid [52]);
tran (stream_cmd_in[58], \stream_cmd_in.guid [53]);
tran (stream_cmd_in[59], \stream_cmd_in.guid [54]);
tran (stream_cmd_in[60], \stream_cmd_in.guid [55]);
tran (stream_cmd_in[61], \stream_cmd_in.guid [56]);
tran (stream_cmd_in[62], \stream_cmd_in.guid [57]);
tran (stream_cmd_in[63], \stream_cmd_in.guid [58]);
tran (stream_cmd_in[64], \stream_cmd_in.guid [59]);
tran (stream_cmd_in[65], \stream_cmd_in.guid [60]);
tran (stream_cmd_in[66], \stream_cmd_in.guid [61]);
tran (stream_cmd_in[67], \stream_cmd_in.guid [62]);
tran (stream_cmd_in[68], \stream_cmd_in.guid [63]);
tran (stream_cmd_in[69], \stream_cmd_in.guid [64]);
tran (stream_cmd_in[70], \stream_cmd_in.guid [65]);
tran (stream_cmd_in[71], \stream_cmd_in.guid [66]);
tran (stream_cmd_in[72], \stream_cmd_in.guid [67]);
tran (stream_cmd_in[73], \stream_cmd_in.guid [68]);
tran (stream_cmd_in[74], \stream_cmd_in.guid [69]);
tran (stream_cmd_in[75], \stream_cmd_in.guid [70]);
tran (stream_cmd_in[76], \stream_cmd_in.guid [71]);
tran (stream_cmd_in[77], \stream_cmd_in.guid [72]);
tran (stream_cmd_in[78], \stream_cmd_in.guid [73]);
tran (stream_cmd_in[79], \stream_cmd_in.guid [74]);
tran (stream_cmd_in[80], \stream_cmd_in.guid [75]);
tran (stream_cmd_in[81], \stream_cmd_in.guid [76]);
tran (stream_cmd_in[82], \stream_cmd_in.guid [77]);
tran (stream_cmd_in[83], \stream_cmd_in.guid [78]);
tran (stream_cmd_in[84], \stream_cmd_in.guid [79]);
tran (stream_cmd_in[85], \stream_cmd_in.guid [80]);
tran (stream_cmd_in[86], \stream_cmd_in.guid [81]);
tran (stream_cmd_in[87], \stream_cmd_in.guid [82]);
tran (stream_cmd_in[88], \stream_cmd_in.guid [83]);
tran (stream_cmd_in[89], \stream_cmd_in.guid [84]);
tran (stream_cmd_in[90], \stream_cmd_in.guid [85]);
tran (stream_cmd_in[91], \stream_cmd_in.guid [86]);
tran (stream_cmd_in[92], \stream_cmd_in.guid [87]);
tran (stream_cmd_in[93], \stream_cmd_in.guid [88]);
tran (stream_cmd_in[94], \stream_cmd_in.guid [89]);
tran (stream_cmd_in[95], \stream_cmd_in.guid [90]);
tran (stream_cmd_in[96], \stream_cmd_in.guid [91]);
tran (stream_cmd_in[97], \stream_cmd_in.guid [92]);
tran (stream_cmd_in[98], \stream_cmd_in.guid [93]);
tran (stream_cmd_in[99], \stream_cmd_in.guid [94]);
tran (stream_cmd_in[100], \stream_cmd_in.guid [95]);
tran (stream_cmd_in[101], \stream_cmd_in.guid [96]);
tran (stream_cmd_in[102], \stream_cmd_in.guid [97]);
tran (stream_cmd_in[103], \stream_cmd_in.guid [98]);
tran (stream_cmd_in[104], \stream_cmd_in.guid [99]);
tran (stream_cmd_in[105], \stream_cmd_in.guid [100]);
tran (stream_cmd_in[106], \stream_cmd_in.guid [101]);
tran (stream_cmd_in[107], \stream_cmd_in.guid [102]);
tran (stream_cmd_in[108], \stream_cmd_in.guid [103]);
tran (stream_cmd_in[109], \stream_cmd_in.guid [104]);
tran (stream_cmd_in[110], \stream_cmd_in.guid [105]);
tran (stream_cmd_in[111], \stream_cmd_in.guid [106]);
tran (stream_cmd_in[112], \stream_cmd_in.guid [107]);
tran (stream_cmd_in[113], \stream_cmd_in.guid [108]);
tran (stream_cmd_in[114], \stream_cmd_in.guid [109]);
tran (stream_cmd_in[115], \stream_cmd_in.guid [110]);
tran (stream_cmd_in[116], \stream_cmd_in.guid [111]);
tran (stream_cmd_in[117], \stream_cmd_in.guid [112]);
tran (stream_cmd_in[118], \stream_cmd_in.guid [113]);
tran (stream_cmd_in[119], \stream_cmd_in.guid [114]);
tran (stream_cmd_in[120], \stream_cmd_in.guid [115]);
tran (stream_cmd_in[121], \stream_cmd_in.guid [116]);
tran (stream_cmd_in[122], \stream_cmd_in.guid [117]);
tran (stream_cmd_in[123], \stream_cmd_in.guid [118]);
tran (stream_cmd_in[124], \stream_cmd_in.guid [119]);
tran (stream_cmd_in[125], \stream_cmd_in.guid [120]);
tran (stream_cmd_in[126], \stream_cmd_in.guid [121]);
tran (stream_cmd_in[127], \stream_cmd_in.guid [122]);
tran (stream_cmd_in[128], \stream_cmd_in.guid [123]);
tran (stream_cmd_in[129], \stream_cmd_in.guid [124]);
tran (stream_cmd_in[130], \stream_cmd_in.guid [125]);
tran (stream_cmd_in[131], \stream_cmd_in.guid [126]);
tran (stream_cmd_in[132], \stream_cmd_in.guid [127]);
tran (stream_cmd_in[133], \stream_cmd_in.guid [128]);
tran (stream_cmd_in[134], \stream_cmd_in.guid [129]);
tran (stream_cmd_in[135], \stream_cmd_in.guid [130]);
tran (stream_cmd_in[136], \stream_cmd_in.guid [131]);
tran (stream_cmd_in[137], \stream_cmd_in.guid [132]);
tran (stream_cmd_in[138], \stream_cmd_in.guid [133]);
tran (stream_cmd_in[139], \stream_cmd_in.guid [134]);
tran (stream_cmd_in[140], \stream_cmd_in.guid [135]);
tran (stream_cmd_in[141], \stream_cmd_in.guid [136]);
tran (stream_cmd_in[142], \stream_cmd_in.guid [137]);
tran (stream_cmd_in[143], \stream_cmd_in.guid [138]);
tran (stream_cmd_in[144], \stream_cmd_in.guid [139]);
tran (stream_cmd_in[145], \stream_cmd_in.guid [140]);
tran (stream_cmd_in[146], \stream_cmd_in.guid [141]);
tran (stream_cmd_in[147], \stream_cmd_in.guid [142]);
tran (stream_cmd_in[148], \stream_cmd_in.guid [143]);
tran (stream_cmd_in[149], \stream_cmd_in.guid [144]);
tran (stream_cmd_in[150], \stream_cmd_in.guid [145]);
tran (stream_cmd_in[151], \stream_cmd_in.guid [146]);
tran (stream_cmd_in[152], \stream_cmd_in.guid [147]);
tran (stream_cmd_in[153], \stream_cmd_in.guid [148]);
tran (stream_cmd_in[154], \stream_cmd_in.guid [149]);
tran (stream_cmd_in[155], \stream_cmd_in.guid [150]);
tran (stream_cmd_in[156], \stream_cmd_in.guid [151]);
tran (stream_cmd_in[157], \stream_cmd_in.guid [152]);
tran (stream_cmd_in[158], \stream_cmd_in.guid [153]);
tran (stream_cmd_in[159], \stream_cmd_in.guid [154]);
tran (stream_cmd_in[160], \stream_cmd_in.guid [155]);
tran (stream_cmd_in[161], \stream_cmd_in.guid [156]);
tran (stream_cmd_in[162], \stream_cmd_in.guid [157]);
tran (stream_cmd_in[163], \stream_cmd_in.guid [158]);
tran (stream_cmd_in[164], \stream_cmd_in.guid [159]);
tran (stream_cmd_in[165], \stream_cmd_in.guid [160]);
tran (stream_cmd_in[166], \stream_cmd_in.guid [161]);
tran (stream_cmd_in[167], \stream_cmd_in.guid [162]);
tran (stream_cmd_in[168], \stream_cmd_in.guid [163]);
tran (stream_cmd_in[169], \stream_cmd_in.guid [164]);
tran (stream_cmd_in[170], \stream_cmd_in.guid [165]);
tran (stream_cmd_in[171], \stream_cmd_in.guid [166]);
tran (stream_cmd_in[172], \stream_cmd_in.guid [167]);
tran (stream_cmd_in[173], \stream_cmd_in.guid [168]);
tran (stream_cmd_in[174], \stream_cmd_in.guid [169]);
tran (stream_cmd_in[175], \stream_cmd_in.guid [170]);
tran (stream_cmd_in[176], \stream_cmd_in.guid [171]);
tran (stream_cmd_in[177], \stream_cmd_in.guid [172]);
tran (stream_cmd_in[178], \stream_cmd_in.guid [173]);
tran (stream_cmd_in[179], \stream_cmd_in.guid [174]);
tran (stream_cmd_in[180], \stream_cmd_in.guid [175]);
tran (stream_cmd_in[181], \stream_cmd_in.guid [176]);
tran (stream_cmd_in[182], \stream_cmd_in.guid [177]);
tran (stream_cmd_in[183], \stream_cmd_in.guid [178]);
tran (stream_cmd_in[184], \stream_cmd_in.guid [179]);
tran (stream_cmd_in[185], \stream_cmd_in.guid [180]);
tran (stream_cmd_in[186], \stream_cmd_in.guid [181]);
tran (stream_cmd_in[187], \stream_cmd_in.guid [182]);
tran (stream_cmd_in[188], \stream_cmd_in.guid [183]);
tran (stream_cmd_in[189], \stream_cmd_in.guid [184]);
tran (stream_cmd_in[190], \stream_cmd_in.guid [185]);
tran (stream_cmd_in[191], \stream_cmd_in.guid [186]);
tran (stream_cmd_in[192], \stream_cmd_in.guid [187]);
tran (stream_cmd_in[193], \stream_cmd_in.guid [188]);
tran (stream_cmd_in[194], \stream_cmd_in.guid [189]);
tran (stream_cmd_in[195], \stream_cmd_in.guid [190]);
tran (stream_cmd_in[196], \stream_cmd_in.guid [191]);
tran (stream_cmd_in[197], \stream_cmd_in.guid [192]);
tran (stream_cmd_in[198], \stream_cmd_in.guid [193]);
tran (stream_cmd_in[199], \stream_cmd_in.guid [194]);
tran (stream_cmd_in[200], \stream_cmd_in.guid [195]);
tran (stream_cmd_in[201], \stream_cmd_in.guid [196]);
tran (stream_cmd_in[202], \stream_cmd_in.guid [197]);
tran (stream_cmd_in[203], \stream_cmd_in.guid [198]);
tran (stream_cmd_in[204], \stream_cmd_in.guid [199]);
tran (stream_cmd_in[205], \stream_cmd_in.guid [200]);
tran (stream_cmd_in[206], \stream_cmd_in.guid [201]);
tran (stream_cmd_in[207], \stream_cmd_in.guid [202]);
tran (stream_cmd_in[208], \stream_cmd_in.guid [203]);
tran (stream_cmd_in[209], \stream_cmd_in.guid [204]);
tran (stream_cmd_in[210], \stream_cmd_in.guid [205]);
tran (stream_cmd_in[211], \stream_cmd_in.guid [206]);
tran (stream_cmd_in[212], \stream_cmd_in.guid [207]);
tran (stream_cmd_in[213], \stream_cmd_in.guid [208]);
tran (stream_cmd_in[214], \stream_cmd_in.guid [209]);
tran (stream_cmd_in[215], \stream_cmd_in.guid [210]);
tran (stream_cmd_in[216], \stream_cmd_in.guid [211]);
tran (stream_cmd_in[217], \stream_cmd_in.guid [212]);
tran (stream_cmd_in[218], \stream_cmd_in.guid [213]);
tran (stream_cmd_in[219], \stream_cmd_in.guid [214]);
tran (stream_cmd_in[220], \stream_cmd_in.guid [215]);
tran (stream_cmd_in[221], \stream_cmd_in.guid [216]);
tran (stream_cmd_in[222], \stream_cmd_in.guid [217]);
tran (stream_cmd_in[223], \stream_cmd_in.guid [218]);
tran (stream_cmd_in[224], \stream_cmd_in.guid [219]);
tran (stream_cmd_in[225], \stream_cmd_in.guid [220]);
tran (stream_cmd_in[226], \stream_cmd_in.guid [221]);
tran (stream_cmd_in[227], \stream_cmd_in.guid [222]);
tran (stream_cmd_in[228], \stream_cmd_in.guid [223]);
tran (stream_cmd_in[229], \stream_cmd_in.guid [224]);
tran (stream_cmd_in[230], \stream_cmd_in.guid [225]);
tran (stream_cmd_in[231], \stream_cmd_in.guid [226]);
tran (stream_cmd_in[232], \stream_cmd_in.guid [227]);
tran (stream_cmd_in[233], \stream_cmd_in.guid [228]);
tran (stream_cmd_in[234], \stream_cmd_in.guid [229]);
tran (stream_cmd_in[235], \stream_cmd_in.guid [230]);
tran (stream_cmd_in[236], \stream_cmd_in.guid [231]);
tran (stream_cmd_in[237], \stream_cmd_in.guid [232]);
tran (stream_cmd_in[238], \stream_cmd_in.guid [233]);
tran (stream_cmd_in[239], \stream_cmd_in.guid [234]);
tran (stream_cmd_in[240], \stream_cmd_in.guid [235]);
tran (stream_cmd_in[241], \stream_cmd_in.guid [236]);
tran (stream_cmd_in[242], \stream_cmd_in.guid [237]);
tran (stream_cmd_in[243], \stream_cmd_in.guid [238]);
tran (stream_cmd_in[244], \stream_cmd_in.guid [239]);
tran (stream_cmd_in[245], \stream_cmd_in.guid [240]);
tran (stream_cmd_in[246], \stream_cmd_in.guid [241]);
tran (stream_cmd_in[247], \stream_cmd_in.guid [242]);
tran (stream_cmd_in[248], \stream_cmd_in.guid [243]);
tran (stream_cmd_in[249], \stream_cmd_in.guid [244]);
tran (stream_cmd_in[250], \stream_cmd_in.guid [245]);
tran (stream_cmd_in[251], \stream_cmd_in.guid [246]);
tran (stream_cmd_in[252], \stream_cmd_in.guid [247]);
tran (stream_cmd_in[253], \stream_cmd_in.guid [248]);
tran (stream_cmd_in[254], \stream_cmd_in.guid [249]);
tran (stream_cmd_in[255], \stream_cmd_in.guid [250]);
tran (stream_cmd_in[256], \stream_cmd_in.guid [251]);
tran (stream_cmd_in[257], \stream_cmd_in.guid [252]);
tran (stream_cmd_in[258], \stream_cmd_in.guid [253]);
tran (stream_cmd_in[259], \stream_cmd_in.guid [254]);
tran (stream_cmd_in[260], \stream_cmd_in.guid [255]);
tran (stream_cmd_in[261], \stream_cmd_in.skip [0]);
tran (stream_cmd_in[262], \stream_cmd_in.combo_mode [0]);
Q_ASSIGN U0 ( .B(kme_internal_out[63]), .A(debug_cmd[31]));
Q_ASSIGN U1 ( .B(kme_internal_out[63]), .A(int_tlv_word0[63]));
Q_ASSIGN U2 ( .B(kme_internal_out[63]), .A(int_tlv_word8[63]));
Q_ASSIGN U3 ( .B(kme_internal_out[63]), .A(int_tlv_word9[63]));
Q_ASSIGN U4 ( .B(kme_internal_out[62]), .A(debug_cmd[30]));
Q_ASSIGN U5 ( .B(kme_internal_out[62]), .A(int_tlv_word0[62]));
Q_ASSIGN U6 ( .B(kme_internal_out[62]), .A(int_tlv_word8[62]));
Q_ASSIGN U7 ( .B(kme_internal_out[62]), .A(int_tlv_word9[62]));
Q_ASSIGN U8 ( .B(kme_internal_out[61]), .A(debug_cmd[29]));
Q_ASSIGN U9 ( .B(kme_internal_out[61]), .A(int_tlv_word0[61]));
Q_ASSIGN U10 ( .B(kme_internal_out[61]), .A(int_tlv_word8[61]));
Q_ASSIGN U11 ( .B(kme_internal_out[61]), .A(int_tlv_word9[61]));
Q_ASSIGN U12 ( .B(kme_internal_out[60]), .A(debug_cmd[28]));
Q_ASSIGN U13 ( .B(kme_internal_out[60]), .A(int_tlv_word0[60]));
Q_ASSIGN U14 ( .B(kme_internal_out[60]), .A(int_tlv_word8[60]));
Q_ASSIGN U15 ( .B(kme_internal_out[60]), .A(int_tlv_word9[60]));
Q_ASSIGN U16 ( .B(kme_internal_out[59]), .A(debug_cmd[27]));
Q_ASSIGN U17 ( .B(kme_internal_out[59]), .A(int_tlv_word0[59]));
Q_ASSIGN U18 ( .B(kme_internal_out[59]), .A(int_tlv_word8[59]));
Q_ASSIGN U19 ( .B(kme_internal_out[59]), .A(int_tlv_word9[59]));
Q_ASSIGN U20 ( .B(kme_internal_out[58]), .A(debug_cmd[26]));
Q_ASSIGN U21 ( .B(kme_internal_out[58]), .A(int_tlv_word0[58]));
Q_ASSIGN U22 ( .B(kme_internal_out[58]), .A(int_tlv_word8[58]));
Q_ASSIGN U23 ( .B(kme_internal_out[58]), .A(int_tlv_word9[58]));
Q_ASSIGN U24 ( .B(kme_internal_out[57]), .A(debug_cmd[25]));
Q_ASSIGN U25 ( .B(kme_internal_out[57]), .A(int_tlv_word0[57]));
Q_ASSIGN U26 ( .B(kme_internal_out[57]), .A(int_tlv_word8[57]));
Q_ASSIGN U27 ( .B(kme_internal_out[57]), .A(int_tlv_word9[57]));
Q_ASSIGN U28 ( .B(kme_internal_out[56]), .A(debug_cmd[24]));
Q_ASSIGN U29 ( .B(kme_internal_out[56]), .A(int_tlv_word0[56]));
Q_ASSIGN U30 ( .B(kme_internal_out[56]), .A(int_tlv_word8[56]));
Q_ASSIGN U31 ( .B(kme_internal_out[56]), .A(int_tlv_word9[56]));
Q_ASSIGN U32 ( .B(kme_internal_out[55]), .A(debug_cmd[23]));
Q_ASSIGN U33 ( .B(kme_internal_out[55]), .A(int_tlv_word0[55]));
Q_ASSIGN U34 ( .B(kme_internal_out[55]), .A(int_tlv_word8[55]));
Q_ASSIGN U35 ( .B(kme_internal_out[55]), .A(int_tlv_word9[55]));
Q_BUF U36 ( .A(corrupt_crc32), .Z(int_tlv_word42[55]));
Q_ASSIGN U37 ( .B(kme_internal_out[54]), .A(debug_cmd[22]));
Q_ASSIGN U38 ( .B(kme_internal_out[54]), .A(int_tlv_word0[54]));
Q_ASSIGN U39 ( .B(kme_internal_out[54]), .A(int_tlv_word8[54]));
Q_ASSIGN U40 ( .B(kme_internal_out[54]), .A(int_tlv_word9[54]));
Q_ASSIGN U41 ( .B(kme_internal_out[54]), .A(int_tlv_word42[54]));
Q_ASSIGN U42 ( .B(kme_internal_out[53]), .A(debug_cmd[21]));
Q_ASSIGN U43 ( .B(kme_internal_out[53]), .A(int_tlv_word0[53]));
Q_ASSIGN U44 ( .B(kme_internal_out[53]), .A(int_tlv_word8[53]));
Q_ASSIGN U45 ( .B(kme_internal_out[53]), .A(int_tlv_word9[53]));
Q_ASSIGN U46 ( .B(kme_internal_out[53]), .A(int_tlv_word42[53]));
Q_ASSIGN U47 ( .B(kme_internal_out[52]), .A(debug_cmd[20]));
Q_ASSIGN U48 ( .B(kme_internal_out[52]), .A(int_tlv_word0[52]));
Q_ASSIGN U49 ( .B(kme_internal_out[52]), .A(int_tlv_word8[52]));
Q_ASSIGN U50 ( .B(kme_internal_out[52]), .A(int_tlv_word9[52]));
Q_ASSIGN U51 ( .B(kme_internal_out[52]), .A(int_tlv_word42[52]));
Q_ASSIGN U52 ( .B(kme_internal_out[51]), .A(debug_cmd[19]));
Q_ASSIGN U53 ( .B(kme_internal_out[51]), .A(int_tlv_word0[51]));
Q_ASSIGN U54 ( .B(kme_internal_out[51]), .A(int_tlv_word8[51]));
Q_ASSIGN U55 ( .B(kme_internal_out[51]), .A(int_tlv_word9[51]));
Q_ASSIGN U56 ( .B(kme_internal_out[51]), .A(int_tlv_word42[51]));
Q_ASSIGN U57 ( .B(kme_internal_out[50]), .A(debug_cmd[18]));
Q_ASSIGN U58 ( .B(kme_internal_out[50]), .A(int_tlv_word0[50]));
Q_ASSIGN U59 ( .B(kme_internal_out[50]), .A(int_tlv_word8[50]));
Q_ASSIGN U60 ( .B(kme_internal_out[50]), .A(int_tlv_word9[50]));
Q_ASSIGN U61 ( .B(kme_internal_out[50]), .A(int_tlv_word42[50]));
Q_ASSIGN U62 ( .B(kme_internal_out[49]), .A(debug_cmd[17]));
Q_ASSIGN U63 ( .B(kme_internal_out[49]), .A(int_tlv_word0[49]));
Q_ASSIGN U64 ( .B(kme_internal_out[49]), .A(int_tlv_word8[49]));
Q_ASSIGN U65 ( .B(kme_internal_out[49]), .A(int_tlv_word9[49]));
Q_ASSIGN U66 ( .B(kme_internal_out[49]), .A(int_tlv_word42[49]));
Q_ASSIGN U67 ( .B(kme_internal_out[48]), .A(debug_cmd[16]));
Q_ASSIGN U68 ( .B(kme_internal_out[48]), .A(int_tlv_word0[48]));
Q_ASSIGN U69 ( .B(kme_internal_out[48]), .A(int_tlv_word8[48]));
Q_ASSIGN U70 ( .B(kme_internal_out[48]), .A(int_tlv_word9[48]));
Q_ASSIGN U71 ( .B(kme_internal_out[48]), .A(int_tlv_word42[48]));
Q_ASSIGN U72 ( .B(kme_internal_out[47]), .A(debug_cmd[15]));
Q_ASSIGN U73 ( .B(kme_internal_out[47]), .A(int_tlv_word0[47]));
Q_ASSIGN U74 ( .B(kme_internal_out[47]), .A(int_tlv_word8[47]));
Q_ASSIGN U75 ( .B(kme_internal_out[47]), .A(int_tlv_word9[47]));
Q_ASSIGN U76 ( .B(kme_internal_out[47]), .A(int_tlv_word42[47]));
Q_ASSIGN U77 ( .B(kme_internal_out[46]), .A(debug_cmd[14]));
Q_ASSIGN U78 ( .B(kme_internal_out[46]), .A(int_tlv_word0[46]));
Q_ASSIGN U79 ( .B(kme_internal_out[46]), .A(int_tlv_word8[46]));
Q_ASSIGN U80 ( .B(kme_internal_out[46]), .A(int_tlv_word9[46]));
Q_ASSIGN U81 ( .B(kme_internal_out[46]), .A(int_tlv_word42[46]));
Q_ASSIGN U82 ( .B(kme_internal_out[45]), .A(debug_cmd[13]));
Q_ASSIGN U83 ( .B(kme_internal_out[45]), .A(int_tlv_word0[45]));
Q_ASSIGN U84 ( .B(kme_internal_out[45]), .A(int_tlv_word8[45]));
Q_ASSIGN U85 ( .B(kme_internal_out[45]), .A(int_tlv_word9[45]));
Q_ASSIGN U86 ( .B(kme_internal_out[45]), .A(int_tlv_word42[45]));
Q_ASSIGN U87 ( .B(kme_internal_out[44]), .A(debug_cmd[12]));
Q_ASSIGN U88 ( .B(kme_internal_out[44]), .A(int_tlv_word0[44]));
Q_ASSIGN U89 ( .B(kme_internal_out[44]), .A(int_tlv_word8[44]));
Q_ASSIGN U90 ( .B(kme_internal_out[44]), .A(int_tlv_word9[44]));
Q_ASSIGN U91 ( .B(kme_internal_out[44]), .A(int_tlv_word42[44]));
Q_ASSIGN U92 ( .B(kme_internal_out[43]), .A(debug_cmd[11]));
Q_ASSIGN U93 ( .B(kme_internal_out[43]), .A(int_tlv_word0[43]));
Q_ASSIGN U94 ( .B(kme_internal_out[43]), .A(int_tlv_word8[43]));
Q_ASSIGN U95 ( .B(kme_internal_out[43]), .A(int_tlv_word9[43]));
Q_ASSIGN U96 ( .B(kme_internal_out[43]), .A(int_tlv_word42[43]));
Q_ASSIGN U97 ( .B(kme_internal_out[42]), .A(debug_cmd[10]));
Q_ASSIGN U98 ( .B(kme_internal_out[42]), .A(int_tlv_word0[42]));
Q_ASSIGN U99 ( .B(kme_internal_out[42]), .A(int_tlv_word8[42]));
Q_ASSIGN U100 ( .B(kme_internal_out[42]), .A(int_tlv_word9[42]));
Q_ASSIGN U101 ( .B(kme_internal_out[42]), .A(int_tlv_word42[42]));
Q_ASSIGN U102 ( .B(kme_internal_out[41]), .A(debug_cmd[9]));
Q_ASSIGN U103 ( .B(kme_internal_out[41]), .A(int_tlv_word0[41]));
Q_ASSIGN U104 ( .B(kme_internal_out[41]), .A(int_tlv_word8[41]));
Q_ASSIGN U105 ( .B(kme_internal_out[41]), .A(int_tlv_word9[41]));
Q_ASSIGN U106 ( .B(kme_internal_out[41]), .A(int_tlv_word42[41]));
Q_ASSIGN U107 ( .B(kme_internal_out[40]), .A(debug_cmd[8]));
Q_ASSIGN U108 ( .B(kme_internal_out[40]), .A(int_tlv_word0[40]));
Q_ASSIGN U109 ( .B(kme_internal_out[40]), .A(int_tlv_word8[40]));
Q_ASSIGN U110 ( .B(kme_internal_out[40]), .A(int_tlv_word9[40]));
Q_ASSIGN U111 ( .B(kme_internal_out[40]), .A(int_tlv_word42[40]));
Q_ASSIGN U112 ( .B(kme_internal_out[39]), .A(debug_cmd[7]));
Q_ASSIGN U113 ( .B(kme_internal_out[39]), .A(int_tlv_word0[39]));
Q_ASSIGN U114 ( .B(kme_internal_out[39]), .A(int_tlv_word8[39]));
Q_ASSIGN U115 ( .B(kme_internal_out[39]), .A(int_tlv_word9[39]));
Q_ASSIGN U116 ( .B(kme_internal_out[39]), .A(int_tlv_word42[39]));
Q_ASSIGN U117 ( .B(kme_internal_out[38]), .A(debug_cmd[6]));
Q_ASSIGN U118 ( .B(kme_internal_out[38]), .A(int_tlv_word0[38]));
Q_ASSIGN U119 ( .B(kme_internal_out[38]), .A(int_tlv_word8[38]));
Q_ASSIGN U120 ( .B(kme_internal_out[38]), .A(int_tlv_word9[38]));
Q_ASSIGN U121 ( .B(kme_internal_out[38]), .A(int_tlv_word42[38]));
Q_ASSIGN U122 ( .B(kme_internal_out[37]), .A(debug_cmd[5]));
Q_ASSIGN U123 ( .B(kme_internal_out[37]), .A(int_tlv_word0[37]));
Q_ASSIGN U124 ( .B(kme_internal_out[37]), .A(int_tlv_word8[37]));
Q_ASSIGN U125 ( .B(kme_internal_out[37]), .A(int_tlv_word9[37]));
Q_ASSIGN U126 ( .B(kme_internal_out[37]), .A(int_tlv_word42[37]));
Q_ASSIGN U127 ( .B(kme_internal_out[36]), .A(debug_cmd[4]));
Q_ASSIGN U128 ( .B(kme_internal_out[36]), .A(int_tlv_word0[36]));
Q_ASSIGN U129 ( .B(kme_internal_out[36]), .A(int_tlv_word8[36]));
Q_ASSIGN U130 ( .B(kme_internal_out[36]), .A(int_tlv_word9[36]));
Q_ASSIGN U131 ( .B(kme_internal_out[36]), .A(int_tlv_word42[36]));
Q_ASSIGN U132 ( .B(kme_internal_out[35]), .A(debug_cmd[3]));
Q_ASSIGN U133 ( .B(kme_internal_out[35]), .A(int_tlv_word0[35]));
Q_ASSIGN U134 ( .B(kme_internal_out[35]), .A(int_tlv_word8[35]));
Q_ASSIGN U135 ( .B(kme_internal_out[35]), .A(int_tlv_word9[35]));
Q_ASSIGN U136 ( .B(kme_internal_out[35]), .A(int_tlv_word42[35]));
Q_ASSIGN U137 ( .B(kme_internal_out[34]), .A(debug_cmd[2]));
Q_ASSIGN U138 ( .B(kme_internal_out[34]), .A(int_tlv_word0[34]));
Q_ASSIGN U139 ( .B(kme_internal_out[34]), .A(int_tlv_word8[34]));
Q_ASSIGN U140 ( .B(kme_internal_out[34]), .A(int_tlv_word9[34]));
Q_ASSIGN U141 ( .B(kme_internal_out[34]), .A(int_tlv_word42[34]));
Q_ASSIGN U142 ( .B(kme_internal_out[33]), .A(debug_cmd[1]));
Q_ASSIGN U143 ( .B(kme_internal_out[33]), .A(int_tlv_word0[33]));
Q_ASSIGN U144 ( .B(kme_internal_out[33]), .A(int_tlv_word8[33]));
Q_ASSIGN U145 ( .B(kme_internal_out[33]), .A(int_tlv_word9[33]));
Q_ASSIGN U146 ( .B(kme_internal_out[33]), .A(int_tlv_word42[33]));
Q_ASSIGN U147 ( .B(kme_internal_out[32]), .A(debug_cmd[0]));
Q_ASSIGN U148 ( .B(kme_internal_out[32]), .A(int_tlv_word0[32]));
Q_ASSIGN U149 ( .B(kme_internal_out[32]), .A(int_tlv_word8[32]));
Q_ASSIGN U150 ( .B(kme_internal_out[32]), .A(int_tlv_word9[32]));
Q_ASSIGN U151 ( .B(kme_internal_out[32]), .A(int_tlv_word42[32]));
Q_ASSIGN U152 ( .B(kme_internal_out[31]), .A(int_tlv_word0[31]));
Q_ASSIGN U153 ( .B(kme_internal_out[31]), .A(int_tlv_word8[31]));
Q_ASSIGN U154 ( .B(kme_internal_out[31]), .A(int_tlv_word9[31]));
Q_ASSIGN U155 ( .B(kme_internal_out[31]), .A(int_tlv_word42[31]));
Q_ASSIGN U156 ( .B(kme_internal_out[31]), .A(key_header[31]));
Q_ASSIGN U157 ( .B(kme_internal_out[30]), .A(int_tlv_word0[30]));
Q_ASSIGN U158 ( .B(kme_internal_out[30]), .A(int_tlv_word8[30]));
Q_ASSIGN U159 ( .B(kme_internal_out[30]), .A(int_tlv_word9[30]));
Q_ASSIGN U160 ( .B(kme_internal_out[30]), .A(int_tlv_word42[30]));
Q_ASSIGN U161 ( .B(kme_internal_out[30]), .A(key_header[30]));
Q_ASSIGN U162 ( .B(kme_internal_out[29]), .A(int_tlv_word0[29]));
Q_ASSIGN U163 ( .B(kme_internal_out[29]), .A(int_tlv_word8[29]));
Q_ASSIGN U164 ( .B(kme_internal_out[29]), .A(int_tlv_word9[29]));
Q_ASSIGN U165 ( .B(kme_internal_out[29]), .A(int_tlv_word42[29]));
Q_ASSIGN U166 ( .B(kme_internal_out[29]), .A(key_header[29]));
Q_ASSIGN U167 ( .B(kme_internal_out[28]), .A(int_tlv_word0[28]));
Q_ASSIGN U168 ( .B(kme_internal_out[28]), .A(int_tlv_word8[28]));
Q_ASSIGN U169 ( .B(kme_internal_out[28]), .A(int_tlv_word9[28]));
Q_ASSIGN U170 ( .B(kme_internal_out[28]), .A(int_tlv_word42[28]));
Q_ASSIGN U171 ( .B(kme_internal_out[28]), .A(key_header[28]));
Q_ASSIGN U172 ( .B(kme_internal_out[27]), .A(int_tlv_word0[27]));
Q_ASSIGN U173 ( .B(kme_internal_out[27]), .A(int_tlv_word8[27]));
Q_ASSIGN U174 ( .B(kme_internal_out[27]), .A(int_tlv_word9[27]));
Q_ASSIGN U175 ( .B(kme_internal_out[27]), .A(int_tlv_word42[27]));
Q_ASSIGN U176 ( .B(kme_internal_out[27]), .A(key_header[27]));
Q_ASSIGN U177 ( .B(kme_internal_out[26]), .A(int_tlv_word0[26]));
Q_ASSIGN U178 ( .B(kme_internal_out[26]), .A(int_tlv_word8[26]));
Q_ASSIGN U179 ( .B(kme_internal_out[26]), .A(int_tlv_word9[26]));
Q_ASSIGN U180 ( .B(kme_internal_out[26]), .A(int_tlv_word42[26]));
Q_ASSIGN U181 ( .B(kme_internal_out[26]), .A(key_header[26]));
Q_ASSIGN U182 ( .B(kme_internal_out[25]), .A(int_tlv_word0[25]));
Q_ASSIGN U183 ( .B(kme_internal_out[25]), .A(int_tlv_word8[25]));
Q_ASSIGN U184 ( .B(kme_internal_out[25]), .A(int_tlv_word9[25]));
Q_ASSIGN U185 ( .B(kme_internal_out[25]), .A(int_tlv_word42[25]));
Q_ASSIGN U186 ( .B(kme_internal_out[25]), .A(key_header[25]));
Q_ASSIGN U187 ( .B(kme_internal_out[24]), .A(int_tlv_word0[24]));
Q_ASSIGN U188 ( .B(kme_internal_out[24]), .A(int_tlv_word8[24]));
Q_ASSIGN U189 ( .B(kme_internal_out[24]), .A(int_tlv_word9[24]));
Q_ASSIGN U190 ( .B(kme_internal_out[24]), .A(int_tlv_word42[24]));
Q_ASSIGN U191 ( .B(kme_internal_out[24]), .A(key_header[24]));
Q_ASSIGN U192 ( .B(kme_internal_out[23]), .A(int_tlv_word0[23]));
Q_ASSIGN U193 ( .B(kme_internal_out[23]), .A(int_tlv_word8[23]));
Q_ASSIGN U194 ( .B(kme_internal_out[23]), .A(int_tlv_word9[23]));
Q_ASSIGN U195 ( .B(kme_internal_out[23]), .A(int_tlv_word42[23]));
Q_ASSIGN U196 ( .B(kme_internal_out[23]), .A(key_header[23]));
Q_ASSIGN U197 ( .B(kme_internal_out[22]), .A(int_tlv_word0[22]));
Q_ASSIGN U198 ( .B(kme_internal_out[22]), .A(int_tlv_word8[22]));
Q_ASSIGN U199 ( .B(kme_internal_out[22]), .A(int_tlv_word9[22]));
Q_ASSIGN U200 ( .B(kme_internal_out[22]), .A(int_tlv_word42[22]));
Q_ASSIGN U201 ( .B(kme_internal_out[22]), .A(key_header[22]));
Q_ASSIGN U202 ( .B(kme_internal_out[21]), .A(int_tlv_word0[21]));
Q_ASSIGN U203 ( .B(kme_internal_out[21]), .A(int_tlv_word8[21]));
Q_ASSIGN U204 ( .B(kme_internal_out[21]), .A(int_tlv_word9[21]));
Q_ASSIGN U205 ( .B(kme_internal_out[21]), .A(int_tlv_word42[21]));
Q_ASSIGN U206 ( .B(kme_internal_out[21]), .A(key_header[21]));
Q_ASSIGN U207 ( .B(kme_internal_out[20]), .A(int_tlv_word0[20]));
Q_ASSIGN U208 ( .B(kme_internal_out[20]), .A(int_tlv_word8[20]));
Q_ASSIGN U209 ( .B(kme_internal_out[20]), .A(int_tlv_word9[20]));
Q_ASSIGN U210 ( .B(kme_internal_out[20]), .A(int_tlv_word42[20]));
Q_ASSIGN U211 ( .B(kme_internal_out[20]), .A(key_header[20]));
Q_ASSIGN U212 ( .B(kme_internal_out[19]), .A(int_tlv_word0[19]));
Q_ASSIGN U213 ( .B(kme_internal_out[19]), .A(int_tlv_word8[19]));
Q_ASSIGN U214 ( .B(kme_internal_out[19]), .A(int_tlv_word9[19]));
Q_ASSIGN U215 ( .B(kme_internal_out[19]), .A(int_tlv_word42[19]));
Q_ASSIGN U216 ( .B(kme_internal_out[19]), .A(key_header[19]));
Q_ASSIGN U217 ( .B(kme_internal_out[18]), .A(int_tlv_word0[18]));
Q_ASSIGN U218 ( .B(kme_internal_out[18]), .A(int_tlv_word8[18]));
Q_ASSIGN U219 ( .B(kme_internal_out[18]), .A(int_tlv_word9[18]));
Q_ASSIGN U220 ( .B(kme_internal_out[18]), .A(int_tlv_word42[18]));
Q_ASSIGN U221 ( .B(kme_internal_out[18]), .A(key_header[18]));
Q_ASSIGN U222 ( .B(kme_internal_out[17]), .A(int_tlv_word0[17]));
Q_ASSIGN U223 ( .B(kme_internal_out[17]), .A(int_tlv_word8[17]));
Q_ASSIGN U224 ( .B(kme_internal_out[17]), .A(int_tlv_word9[17]));
Q_ASSIGN U225 ( .B(kme_internal_out[17]), .A(int_tlv_word42[17]));
Q_ASSIGN U226 ( .B(kme_internal_out[17]), .A(key_header[17]));
Q_ASSIGN U227 ( .B(kme_internal_out[16]), .A(int_tlv_word0[16]));
Q_ASSIGN U228 ( .B(kme_internal_out[16]), .A(int_tlv_word8[16]));
Q_ASSIGN U229 ( .B(kme_internal_out[16]), .A(int_tlv_word9[16]));
Q_ASSIGN U230 ( .B(kme_internal_out[16]), .A(int_tlv_word42[16]));
Q_ASSIGN U231 ( .B(kme_internal_out[16]), .A(key_header[16]));
Q_ASSIGN U232 ( .B(kme_internal_out[15]), .A(int_tlv_word0[15]));
Q_ASSIGN U233 ( .B(kme_internal_out[15]), .A(int_tlv_word8[15]));
Q_ASSIGN U234 ( .B(kme_internal_out[15]), .A(int_tlv_word9[15]));
Q_ASSIGN U235 ( .B(kme_internal_out[15]), .A(int_tlv_word42[15]));
Q_ASSIGN U236 ( .B(kme_internal_out[15]), .A(key_header[15]));
Q_ASSIGN U237 ( .B(kme_internal_out[14]), .A(int_tlv_word0[14]));
Q_ASSIGN U238 ( .B(kme_internal_out[14]), .A(int_tlv_word8[14]));
Q_ASSIGN U239 ( .B(kme_internal_out[14]), .A(int_tlv_word9[14]));
Q_ASSIGN U240 ( .B(kme_internal_out[14]), .A(int_tlv_word42[14]));
Q_ASSIGN U241 ( .B(kme_internal_out[14]), .A(key_header[14]));
Q_ASSIGN U242 ( .B(kme_internal_out[13]), .A(int_tlv_word0[13]));
Q_ASSIGN U243 ( .B(kme_internal_out[13]), .A(int_tlv_word8[13]));
Q_ASSIGN U244 ( .B(kme_internal_out[13]), .A(int_tlv_word9[13]));
Q_ASSIGN U245 ( .B(kme_internal_out[13]), .A(int_tlv_word42[13]));
Q_ASSIGN U246 ( .B(kme_internal_out[13]), .A(key_header[13]));
Q_ASSIGN U247 ( .B(kme_internal_out[12]), .A(int_tlv_word0[12]));
Q_ASSIGN U248 ( .B(kme_internal_out[12]), .A(int_tlv_word8[12]));
Q_ASSIGN U249 ( .B(kme_internal_out[12]), .A(int_tlv_word9[12]));
Q_ASSIGN U250 ( .B(kme_internal_out[12]), .A(int_tlv_word42[12]));
Q_ASSIGN U251 ( .B(kme_internal_out[12]), .A(key_header[12]));
Q_ASSIGN U252 ( .B(kme_internal_out[11]), .A(int_tlv_word0[11]));
Q_ASSIGN U253 ( .B(kme_internal_out[11]), .A(int_tlv_word8[11]));
Q_ASSIGN U254 ( .B(kme_internal_out[11]), .A(int_tlv_word9[11]));
Q_ASSIGN U255 ( .B(kme_internal_out[11]), .A(int_tlv_word42[11]));
Q_ASSIGN U256 ( .B(kme_internal_out[11]), .A(key_header[11]));
Q_ASSIGN U257 ( .B(kme_internal_out[10]), .A(int_tlv_word0[10]));
Q_ASSIGN U258 ( .B(kme_internal_out[10]), .A(int_tlv_word8[10]));
Q_ASSIGN U259 ( .B(kme_internal_out[10]), .A(int_tlv_word9[10]));
Q_ASSIGN U260 ( .B(kme_internal_out[10]), .A(int_tlv_word42[10]));
Q_ASSIGN U261 ( .B(kme_internal_out[10]), .A(key_header[10]));
Q_ASSIGN U262 ( .B(kme_internal_out[9]), .A(int_tlv_word0[9]));
Q_ASSIGN U263 ( .B(kme_internal_out[9]), .A(int_tlv_word8[9]));
Q_ASSIGN U264 ( .B(kme_internal_out[9]), .A(int_tlv_word9[9]));
Q_ASSIGN U265 ( .B(kme_internal_out[9]), .A(int_tlv_word42[9]));
Q_ASSIGN U266 ( .B(kme_internal_out[9]), .A(key_header[9]));
Q_ASSIGN U267 ( .B(kme_internal_out[8]), .A(int_tlv_word0[8]));
Q_ASSIGN U268 ( .B(kme_internal_out[8]), .A(int_tlv_word8[8]));
Q_ASSIGN U269 ( .B(kme_internal_out[8]), .A(int_tlv_word9[8]));
Q_ASSIGN U270 ( .B(kme_internal_out[8]), .A(int_tlv_word42[8]));
Q_ASSIGN U271 ( .B(kme_internal_out[8]), .A(key_header[8]));
Q_ASSIGN U272 ( .B(kme_internal_out[7]), .A(int_tlv_word0[7]));
Q_ASSIGN U273 ( .B(kme_internal_out[7]), .A(int_tlv_word8[7]));
Q_ASSIGN U274 ( .B(kme_internal_out[7]), .A(int_tlv_word9[7]));
Q_ASSIGN U275 ( .B(kme_internal_out[7]), .A(int_tlv_word42[7]));
Q_ASSIGN U276 ( .B(kme_internal_out[7]), .A(key_header[7]));
Q_ASSIGN U277 ( .B(kme_internal_out[6]), .A(int_tlv_word0[6]));
Q_ASSIGN U278 ( .B(kme_internal_out[6]), .A(int_tlv_word8[6]));
Q_ASSIGN U279 ( .B(kme_internal_out[6]), .A(int_tlv_word9[6]));
Q_ASSIGN U280 ( .B(kme_internal_out[6]), .A(int_tlv_word42[6]));
Q_ASSIGN U281 ( .B(kme_internal_out[6]), .A(key_header[6]));
Q_ASSIGN U282 ( .B(kme_internal_out[5]), .A(int_tlv_word0[5]));
Q_ASSIGN U283 ( .B(kme_internal_out[5]), .A(int_tlv_word8[5]));
Q_ASSIGN U284 ( .B(kme_internal_out[5]), .A(int_tlv_word9[5]));
Q_ASSIGN U285 ( .B(kme_internal_out[5]), .A(int_tlv_word42[5]));
Q_ASSIGN U286 ( .B(kme_internal_out[5]), .A(key_header[5]));
Q_ASSIGN U287 ( .B(kme_internal_out[4]), .A(int_tlv_word0[4]));
Q_ASSIGN U288 ( .B(kme_internal_out[4]), .A(int_tlv_word8[4]));
Q_ASSIGN U289 ( .B(kme_internal_out[4]), .A(int_tlv_word9[4]));
Q_ASSIGN U290 ( .B(kme_internal_out[4]), .A(int_tlv_word42[4]));
Q_ASSIGN U291 ( .B(kme_internal_out[4]), .A(key_header[4]));
Q_ASSIGN U292 ( .B(kme_internal_out[3]), .A(int_tlv_word0[3]));
Q_ASSIGN U293 ( .B(kme_internal_out[3]), .A(int_tlv_word8[3]));
Q_ASSIGN U294 ( .B(kme_internal_out[3]), .A(int_tlv_word9[3]));
Q_ASSIGN U295 ( .B(kme_internal_out[3]), .A(int_tlv_word42[3]));
Q_ASSIGN U296 ( .B(kme_internal_out[3]), .A(key_header[3]));
Q_ASSIGN U297 ( .B(kme_internal_out[2]), .A(int_tlv_word0[2]));
Q_ASSIGN U298 ( .B(kme_internal_out[2]), .A(int_tlv_word8[2]));
Q_ASSIGN U299 ( .B(kme_internal_out[2]), .A(int_tlv_word9[2]));
Q_ASSIGN U300 ( .B(kme_internal_out[2]), .A(int_tlv_word42[2]));
Q_ASSIGN U301 ( .B(kme_internal_out[2]), .A(key_header[2]));
Q_ASSIGN U302 ( .B(kme_internal_out[1]), .A(int_tlv_word0[1]));
Q_ASSIGN U303 ( .B(kme_internal_out[1]), .A(int_tlv_word8[1]));
Q_ASSIGN U304 ( .B(kme_internal_out[1]), .A(int_tlv_word9[1]));
Q_ASSIGN U305 ( .B(kme_internal_out[1]), .A(int_tlv_word42[1]));
Q_ASSIGN U306 ( .B(kme_internal_out[1]), .A(key_header[1]));
Q_ASSIGN U307 ( .B(kme_internal_out[0]), .A(int_tlv_word0[0]));
Q_ASSIGN U308 ( .B(kme_internal_out[0]), .A(int_tlv_word8[0]));
Q_ASSIGN U309 ( .B(kme_internal_out[0]), .A(int_tlv_word9[0]));
Q_ASSIGN U310 ( .B(kme_internal_out[0]), .A(int_tlv_word42[0]));
Q_ASSIGN U311 ( .B(kme_internal_out[0]), .A(key_header[0]));
Q_BUF U312 ( .A(_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_reset_or), .Z(_zy_sva_brcm_gcm_dek512_with_512bit_key_2_reset_or));
Q_BUF U313 ( .A(_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_reset_or), .Z(_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_reset_or));
Q_BUF U314 ( .A(_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_reset_or), .Z(_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_reset_or));
Q_BUF U315 ( .A(_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_reset_or), .Z(_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_reset_or));
Q_BUF U316 ( .A(_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_reset_or), .Z(_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_reset_or));
Q_BUF U317 ( .A(_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_reset_or), .Z(_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_reset_or));
Q_BUF U318 ( .A(_zy_sva_brcm_tlv_sb_stall_on_guid_9_reset_or), .Z(_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_reset_or));
Q_BUF U319 ( .A(_zy_sva_brcm_gcm_10_reset_or), .Z(_zy_sva_brcm_tlv_sb_stall_on_guid_9_reset_or));
Q_BUF U320 ( .A(_zy_sva_brcm_gcm_11_reset_or), .Z(_zy_sva_brcm_gcm_10_reset_or));
Q_BUF U321 ( .A(_zy_sva_brcm_gcm_12_reset_or), .Z(_zy_sva_brcm_gcm_11_reset_or));
Q_BUF U322 ( .A(_zy_sva_brcm_gcm_13_reset_or), .Z(_zy_sva_brcm_gcm_12_reset_or));
Q_BUF U323 ( .A(_zy_sva_brcm_gcm_14_reset_or), .Z(_zy_sva_brcm_gcm_13_reset_or));
Q_BUF U324 ( .A(_zy_sva_brcm_gcm_15_reset_or), .Z(_zy_sva_brcm_gcm_14_reset_or));
Q_BUF U325 ( .A(_zy_sva_brcm_gcm_16_reset_or), .Z(_zy_sva_brcm_gcm_15_reset_or));
Q_BUF U326 ( .A(_zy_sva_brcm_gcm_17_reset_or), .Z(_zy_sva_brcm_gcm_16_reset_or));
Q_BUF U327 ( .A(_zy_sva_brcm_kdf_label0_8_18_reset_or), .Z(_zy_sva_brcm_gcm_17_reset_or));
Q_BUF U328 ( .A(_zy_sva_brcm_kdf_label9_16_19_reset_or), .Z(_zy_sva_brcm_kdf_label0_8_18_reset_or));
Q_BUF U329 ( .A(_zy_sva_brcm_kdf_label17_24_20_reset_or), .Z(_zy_sva_brcm_kdf_label9_16_19_reset_or));
Q_BUF U330 ( .A(_zy_sva_brcm_kdf_label25_32_21_reset_or), .Z(_zy_sva_brcm_kdf_label17_24_20_reset_or));
Q_BUF U331 ( .A(_zy_sva_brcm_kdf_label0_8_22_reset_or), .Z(_zy_sva_brcm_kdf_label25_32_21_reset_or));
Q_BUF U332 ( .A(_zy_sva_brcm_kdf_label9_16_23_reset_or), .Z(_zy_sva_brcm_kdf_label0_8_22_reset_or));
Q_BUF U333 ( .A(_zy_sva_brcm_kdf_label17_24_24_reset_or), .Z(_zy_sva_brcm_kdf_label9_16_23_reset_or));
Q_BUF U334 ( .A(_zy_sva_brcm_kdf_label25_32_25_reset_or), .Z(_zy_sva_brcm_kdf_label17_24_24_reset_or));
Q_BUF U335 ( .A(_zy_sva_brcm_kdf_label0_8_26_reset_or), .Z(_zy_sva_brcm_kdf_label25_32_25_reset_or));
Q_BUF U336 ( .A(_zy_sva_brcm_kdf_label9_16_27_reset_or), .Z(_zy_sva_brcm_kdf_label0_8_26_reset_or));
Q_BUF U337 ( .A(_zy_sva_brcm_kdf_label17_24_28_reset_or), .Z(_zy_sva_brcm_kdf_label9_16_27_reset_or));
Q_BUF U338 ( .A(_zy_sva_brcm_kdf_label25_32_29_reset_or), .Z(_zy_sva_brcm_kdf_label17_24_28_reset_or));
Q_BUF U339 ( .A(_zy_sva_brcm_kdf_label0_8_30_reset_or), .Z(_zy_sva_brcm_kdf_label25_32_29_reset_or));
Q_BUF U340 ( .A(_zy_sva_brcm_kdf_label9_16_31_reset_or), .Z(_zy_sva_brcm_kdf_label0_8_30_reset_or));
Q_BUF U341 ( .A(_zy_sva_brcm_kdf_label17_24_32_reset_or), .Z(_zy_sva_brcm_kdf_label9_16_31_reset_or));
Q_BUF U342 ( .A(_zy_sva_brcm_kdf_label25_32_33_reset_or), .Z(_zy_sva_brcm_kdf_label17_24_32_reset_or));
Q_BUF U343 ( .A(_zy_sva_brcm_gcm_dek256_with_512bit_key_1_reset_or), .Z(_zy_sva_brcm_kdf_label25_32_33_reset_or));
Q_BUF U344 ( .A(keyfilter_cmd_in_valid), .Z(kdf_cmd_in_valid));
Q_BUF U345 ( .A(keyfilter_cmd_in[0]), .Z(kdf_cmd_in[2]));
Q_OR02 U346 ( .A0(n29), .A1(n28), .Z(n1));
Q_OR02 U347 ( .A0(n8), .A1(n7), .Z(n2801));
Q_MX08 U348 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][271] ), .A1(\labels[1][271] ), .A2(\labels[2][271] ), .A3(\labels[3][271] ), .A4(\labels[4][271] ), .A5(\labels[5][271] ), .A6(\labels[6][271] ), .A7(\labels[7][271] ), .Z(n2));
Q_MX08 U349 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][270] ), .A1(\labels[1][270] ), .A2(\labels[2][270] ), .A3(\labels[3][270] ), .A4(\labels[4][270] ), .A5(\labels[5][270] ), .A6(\labels[6][270] ), .A7(\labels[7][270] ), .Z(n3));
Q_MX08 U350 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][269] ), .A1(\labels[1][269] ), .A2(\labels[2][269] ), .A3(\labels[3][269] ), .A4(\labels[4][269] ), .A5(\labels[5][269] ), .A6(\labels[6][269] ), .A7(\labels[7][269] ), .Z(n4));
Q_MX08 U351 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][268] ), .A1(\labels[1][268] ), .A2(\labels[2][268] ), .A3(\labels[3][268] ), .A4(\labels[4][268] ), .A5(\labels[5][268] ), .A6(\labels[6][268] ), .A7(\labels[7][268] ), .Z(n5));
Q_MX08 U352 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][267] ), .A1(\labels[1][267] ), .A2(\labels[2][267] ), .A3(\labels[3][267] ), .A4(\labels[4][267] ), .A5(\labels[5][267] ), .A6(\labels[6][267] ), .A7(\labels[7][267] ), .Z(n6));
Q_MX08 U353 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][266] ), .A1(\labels[1][266] ), .A2(\labels[2][266] ), .A3(\labels[3][266] ), .A4(\labels[4][266] ), .A5(\labels[5][266] ), .A6(\labels[6][266] ), .A7(\labels[7][266] ), .Z(n7));
Q_MX08 U354 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][265] ), .A1(\labels[1][265] ), .A2(\labels[2][265] ), .A3(\labels[3][265] ), .A4(\labels[4][265] ), .A5(\labels[5][265] ), .A6(\labels[6][265] ), .A7(\labels[7][265] ), .Z(n8));
Q_MX08 U355 ( .S0(kdfstream_cmd_in[2]), .S1(kdfstream_cmd_in[3]), .S2(kdfstream_cmd_in[4]), .A0(\labels[0][8] ), .A1(\labels[1][8] ), .A2(\labels[2][8] ), .A3(\labels[3][8] ), .A4(\labels[4][8] ), .A5(\labels[5][8] ), .A6(\labels[6][8] ), .A7(\labels[7][8] ), .Z(n9));
Q_AN03 U356 ( .A0(kme_internal_out_ack), .A1(n12), .A2(n11), .Z(n10));
Q_INV U357 ( .A(kme_internal_out[69]), .Z(n11));
Q_NR02 U358 ( .A0(kme_internal_out[64]), .A1(n13), .Z(n12));
Q_OR03 U359 ( .A0(kme_internal_out[67]), .A1(n14), .A2(kme_internal_out[65]), .Z(n13));
Q_INV U360 ( .A(kme_internal_out[66]), .Z(n14));
Q_OR02 U361 ( .A0(n2735), .A1(n116), .Z(n83));
Q_INV U362 ( .A(kme_internal_out_ack), .Z(n128));
Q_OR03 U363 ( .A0(n11), .A1(n119), .A2(n83), .Z(n39));
Q_ND02 U364 ( .A0(kme_internal_out[69]), .A1(n63), .Z(n40));
Q_NR02 U365 ( .A0(n40), .A1(n83), .Z(n41));
Q_OR02 U366 ( .A0(n44), .A1(n83), .Z(n42));
Q_INV U367 ( .A(n42), .Z(gcm_cmd_in_valid));
Q_AN02 U368 ( .A0(kme_internal_out_ack), .A1(n16), .Z(n32));
Q_AN02 U369 ( .A0(kme_internal_out[69]), .A1(n32), .Z(n24));
Q_INV U370 ( .A(n15), .Z(n43));
Q_NR03 U371 ( .A0(n43), .A1(n16), .A2(n44), .Z(n45));
Q_INV U372 ( .A(n46), .Z(n44));
Q_OA21 U373 ( .A0(n15), .A1(n16), .B0(n46), .Z(gcm_tag_data_in_valid));
Q_AN02 U374 ( .A0(kme_internal_out[69]), .A1(kme_internal_out_ack), .Z(n46));
Q_OR02 U375 ( .A0(kme_internal_out[65]), .A1(n2731), .Z(n68));
Q_OA21 U376 ( .A0(n2735), .A1(n68), .B0(kme_internal_out[66]), .Z(n51));
Q_XOR2 U377 ( .A0(kme_internal_out[65]), .A1(n2731), .Z(n47));
Q_OA21 U378 ( .A0(n2735), .A1(n47), .B0(n14), .Z(n48));
Q_NR03 U379 ( .A0(n51), .A1(n48), .A2(n128), .Z(inspector_upsizer_valid));
Q_INV U380 ( .A(kme_internal_out[65]), .Z(n49));
Q_OR02 U381 ( .A0(n49), .A1(kme_internal_out[64]), .Z(n121));
Q_OA21 U382 ( .A0(n2735), .A1(n121), .B0(n14), .Z(n50));
Q_NR03 U383 ( .A0(n51), .A1(n50), .A2(n128), .Z(n52));
Q_OR03 U384 ( .A0(kme_internal_out[67]), .A1(n116), .A2(n53), .Z(n57));
Q_INV U385 ( .A(n63), .Z(n53));
Q_OR02 U386 ( .A0(kme_internal_out[69]), .A1(n57), .Z(n56));
Q_OA21 U387 ( .A0(n57), .A1(stream_cmd_in[262]), .B0(n58), .Z(n54));
Q_INV U388 ( .A(n54), .Z(kdfstream_cmd_in_valid));
Q_INV U389 ( .A(n56), .Z(n26));
Q_OR02 U390 ( .A0(n56), .A1(n55), .Z(n58));
Q_OR03 U391 ( .A0(n11), .A1(n57), .A2(stream_cmd_in[262]), .Z(n60));
Q_AN02 U392 ( .A0(n58), .A1(n60), .Z(n59));
Q_INV U393 ( .A(n59), .Z(n25));
Q_INV U394 ( .A(n60), .Z(n27));
Q_INV U395 ( .A(n68), .Z(n61));
Q_OR02 U396 ( .A0(kme_internal_out[67]), .A1(n61), .Z(n65));
Q_OR02 U397 ( .A0(n119), .A1(n65), .Z(n62));
Q_INV U398 ( .A(n62), .Z(n28));
Q_AN02 U399 ( .A0(kme_internal_out[65]), .A1(kme_internal_out[64]), .Z(n70));
Q_AN02 U400 ( .A0(kme_internal_out[67]), .A1(n70), .Z(n64));
Q_AN02 U401 ( .A0(kme_internal_out_ack), .A1(kme_internal_out[66]), .Z(n63));
Q_AN02 U402 ( .A0(n63), .A1(n64), .Z(n29));
Q_INV U403 ( .A(n65), .Z(n66));
Q_MX02 U404 ( .S(kme_internal_out[66]), .A0(n66), .A1(n64), .Z(n67));
Q_AN02 U405 ( .A0(kme_internal_out_ack), .A1(n67), .Z(tlv_sb_data_in_valid));
Q_OR02 U406 ( .A0(kme_internal_out[67]), .A1(n68), .Z(n125));
Q_OR02 U407 ( .A0(n119), .A1(n125), .Z(n31));
Q_NR02 U408 ( .A0(n143), .A1(n31), .Z(n69));
Q_INV U409 ( .A(n70), .Z(n71));
Q_OR02 U410 ( .A0(kme_internal_out[67]), .A1(n71), .Z(n87));
Q_OR02 U411 ( .A0(n119), .A1(n87), .Z(n72));
Q_OR03 U412 ( .A0(kme_internal_out[67]), .A1(n2731), .A2(n119), .Z(n30));
Q_AN02 U413 ( .A0(kme_internal_out_ack), .A1(n15), .Z(n33));
Q_OR02 U414 ( .A0(kme_internal_out[40]), .A1(kme_internal_out[39]), .Z(n98));
Q_INV U415 ( .A(n98), .Z(n73));
Q_OA21 U416 ( .A0(kme_internal_out[41]), .A1(n73), .B0(kme_internal_out[42]), .Z(n75));
Q_INV U417 ( .A(kme_internal_out[42]), .Z(n110));
Q_INV U418 ( .A(kme_internal_out[41]), .Z(n106));
Q_AN02 U419 ( .A0(kme_internal_out[40]), .A1(kme_internal_out[39]), .Z(n74));
Q_MX02 U420 ( .S(kme_internal_out[41]), .A0(n98), .A1(n74), .Z(n78));
Q_NR03 U421 ( .A0(n75), .A1(n79), .A2(n76), .Z(n77));
Q_OR03 U422 ( .A0(n128), .A1(n103), .A2(n114), .Z(n76));
Q_OA21 U423 ( .A0(n106), .A1(kme_internal_out[40]), .B0(kme_internal_out[42]), .Z(n80));
Q_AN02 U424 ( .A0(n78), .A1(n110), .Z(n79));
Q_OR03 U425 ( .A0(n80), .A1(n79), .A2(n81), .Z(n88));
Q_OR02 U426 ( .A0(kme_internal_out[67]), .A1(n114), .Z(n81));
Q_OR02 U427 ( .A0(n119), .A1(n88), .Z(n82));
Q_INV U428 ( .A(n82), .Z(n34));
Q_AO21 U429 ( .A0(n83), .A1(kme_internal_out[66]), .B0(n84), .Z(n85));
Q_AN02 U430 ( .A0(n88), .A1(n14), .Z(n84));
Q_OR02 U431 ( .A0(n128), .A1(n85), .Z(n86));
Q_AO21 U432 ( .A0(n87), .A1(kme_internal_out[66]), .B0(n84), .Z(n89));
Q_OR02 U433 ( .A0(n128), .A1(n89), .Z(n90));
Q_INV U434 ( .A(kme_internal_out[40]), .Z(n91));
Q_OR03 U435 ( .A0(n91), .A1(kme_internal_out[39]), .A2(kme_internal_out[41]), .Z(n92));
Q_AN02 U436 ( .A0(n98), .A1(kme_internal_out[41]), .Z(n93));
Q_INV U437 ( .A(kme_internal_out[39]), .Z(n99));
Q_OR02 U438 ( .A0(kme_internal_out[40]), .A1(n99), .Z(n108));
Q_AO21 U439 ( .A0(n108), .A1(n106), .B0(n93), .Z(n94));
Q_INV U440 ( .A(n94), .Z(n95));
Q_MX02 U441 ( .S(kme_internal_out[42]), .A0(n95), .A1(n92), .Z(n96));
Q_NR02 U442 ( .A0(n112), .A1(n96), .Z(n97));
Q_OR02 U443 ( .A0(n35), .A1(n97), .Z(n37));
Q_XOR2 U444 ( .A0(kme_internal_out[40]), .A1(n99), .Z(n107));
Q_INV U445 ( .A(n107), .Z(n104));
Q_NR02 U446 ( .A0(n107), .A1(kme_internal_out[41]), .Z(n100));
Q_NR03 U447 ( .A0(n93), .A1(n100), .A2(n101), .Z(n102));
Q_OR03 U448 ( .A0(kme_internal_out[43]), .A1(n110), .A2(kme_internal_out[44]), .Z(n101));
Q_OR03 U449 ( .A0(n103), .A1(n116), .A2(n128), .Z(n35));
Q_OR02 U450 ( .A0(kme_internal_out[66]), .A1(kme_internal_out[67]), .Z(n103));
Q_OR02 U451 ( .A0(n35), .A1(n102), .Z(n38));
Q_MX02 U452 ( .S(kme_internal_out[41]), .A0(n104), .A1(n108), .Z(n105));
Q_INV U453 ( .A(n108), .Z(n109));
Q_MX02 U454 ( .S(kme_internal_out[41]), .A0(n109), .A1(n107), .Z(n111));
Q_MX02 U455 ( .S(kme_internal_out[42]), .A0(n111), .A1(n105), .Z(n113));
Q_OR02 U456 ( .A0(kme_internal_out[44]), .A1(kme_internal_out[43]), .Z(n112));
Q_OR02 U457 ( .A0(n116), .A1(n112), .Z(n114));
Q_OR02 U458 ( .A0(kme_internal_out[65]), .A1(kme_internal_out[64]), .Z(n116));
Q_OR02 U459 ( .A0(n114), .A1(n113), .Z(n117));
Q_OR02 U460 ( .A0(kme_internal_out[67]), .A1(n117), .Z(n126));
Q_OR02 U461 ( .A0(n119), .A1(n126), .Z(n115));
Q_INV U462 ( .A(n115), .Z(n36));
Q_MX02 U463 ( .S(kme_internal_out[67]), .A0(n117), .A1(n116), .Z(n118));
Q_OR02 U464 ( .A0(n128), .A1(kme_internal_out[66]), .Z(n119));
Q_OR02 U465 ( .A0(n119), .A1(n118), .Z(n120));
Q_OA21 U466 ( .A0(kme_internal_out[67]), .A1(n121), .B0(kme_internal_out[66]), .Z(n123));
Q_AN02 U467 ( .A0(n126), .A1(n14), .Z(n122));
Q_OR03 U468 ( .A0(n123), .A1(n122), .A2(n128), .Z(n124));
Q_AO21 U469 ( .A0(n125), .A1(kme_internal_out[66]), .B0(n122), .Z(n127));
Q_OR02 U470 ( .A0(n128), .A1(n127), .Z(n129));
Q_OR03 U471 ( .A0(n131), .A1(n130), .A2(n133), .Z(n137));
Q_OR03 U472 ( .A0(n18), .A1(n17), .A2(n132), .Z(n133));
Q_OR03 U473 ( .A0(n135), .A1(n134), .A2(n136), .Z(n138));
Q_OR02 U474 ( .A0(n23), .A1(n22), .Z(n136));
Q_NR02 U475 ( .A0(n138), .A1(n137), .Z(n139));
Q_MX02 U476 ( .S(n31), .A0(n140), .A1(stream_cmd_in[1]), .Z(stream_cmd_in_nxt[1]));
Q_MX02 U477 ( .S(n31), .A0(n142), .A1(stream_cmd_in[0]), .Z(stream_cmd_in_nxt[0]));
Q_XOR2 U478 ( .A0(kme_internal_out[16]), .A1(n141), .Z(n140));
Q_AD01HF U479 ( .A0(kdf_dek_iter), .B0(n143), .S(n142), .CO(n141));
Q_INV U480 ( .A(kme_internal_out[16]), .Z(n143));
Q_MX02 U481 ( .S(n39), .A0(gcm_dek_cmd_in[610]), .A1(n144), .Z(gcm_cmd_in[610]));
Q_AN02 U482 ( .A0(n41), .A1(gcm_dak_cmd_in[610]), .Z(n144));
Q_MX02 U483 ( .S(n39), .A0(gcm_dek_cmd_in[609]), .A1(n145), .Z(gcm_cmd_in[609]));
Q_AN02 U484 ( .A0(n41), .A1(gcm_dak_cmd_in[609]), .Z(n145));
Q_MX02 U485 ( .S(n39), .A0(gcm_dek_cmd_in[608]), .A1(n146), .Z(gcm_cmd_in[608]));
Q_AN02 U486 ( .A0(n41), .A1(gcm_dak_cmd_in[608]), .Z(n146));
Q_MX02 U487 ( .S(n39), .A0(gcm_dek_cmd_in[607]), .A1(n147), .Z(gcm_cmd_in[607]));
Q_AN02 U488 ( .A0(n41), .A1(gcm_dak_cmd_in[607]), .Z(n147));
Q_MX02 U489 ( .S(n39), .A0(gcm_dek_cmd_in[606]), .A1(n148), .Z(gcm_cmd_in[606]));
Q_AN02 U490 ( .A0(n41), .A1(gcm_dak_cmd_in[606]), .Z(n148));
Q_MX02 U491 ( .S(n39), .A0(gcm_dek_cmd_in[605]), .A1(n149), .Z(gcm_cmd_in[605]));
Q_AN02 U492 ( .A0(n41), .A1(gcm_dak_cmd_in[605]), .Z(n149));
Q_MX02 U493 ( .S(n39), .A0(gcm_dek_cmd_in[604]), .A1(n150), .Z(gcm_cmd_in[604]));
Q_AN02 U494 ( .A0(n41), .A1(gcm_dak_cmd_in[604]), .Z(n150));
Q_MX02 U495 ( .S(n39), .A0(gcm_dek_cmd_in[603]), .A1(n151), .Z(gcm_cmd_in[603]));
Q_AN02 U496 ( .A0(n41), .A1(gcm_dak_cmd_in[603]), .Z(n151));
Q_MX02 U497 ( .S(n39), .A0(gcm_dek_cmd_in[602]), .A1(n152), .Z(gcm_cmd_in[602]));
Q_AN02 U498 ( .A0(n41), .A1(gcm_dak_cmd_in[602]), .Z(n152));
Q_MX02 U499 ( .S(n39), .A0(gcm_dek_cmd_in[601]), .A1(n153), .Z(gcm_cmd_in[601]));
Q_AN02 U500 ( .A0(n41), .A1(gcm_dak_cmd_in[601]), .Z(n153));
Q_MX02 U501 ( .S(n39), .A0(gcm_dek_cmd_in[600]), .A1(n154), .Z(gcm_cmd_in[600]));
Q_AN02 U502 ( .A0(n41), .A1(gcm_dak_cmd_in[600]), .Z(n154));
Q_MX02 U503 ( .S(n39), .A0(gcm_dek_cmd_in[599]), .A1(n155), .Z(gcm_cmd_in[599]));
Q_AN02 U504 ( .A0(n41), .A1(gcm_dak_cmd_in[599]), .Z(n155));
Q_MX02 U505 ( .S(n39), .A0(gcm_dek_cmd_in[598]), .A1(n156), .Z(gcm_cmd_in[598]));
Q_AN02 U506 ( .A0(n41), .A1(gcm_dak_cmd_in[598]), .Z(n156));
Q_MX02 U507 ( .S(n39), .A0(gcm_dek_cmd_in[597]), .A1(n157), .Z(gcm_cmd_in[597]));
Q_AN02 U508 ( .A0(n41), .A1(gcm_dak_cmd_in[597]), .Z(n157));
Q_MX02 U509 ( .S(n39), .A0(gcm_dek_cmd_in[596]), .A1(n158), .Z(gcm_cmd_in[596]));
Q_AN02 U510 ( .A0(n41), .A1(gcm_dak_cmd_in[596]), .Z(n158));
Q_MX02 U511 ( .S(n39), .A0(gcm_dek_cmd_in[595]), .A1(n159), .Z(gcm_cmd_in[595]));
Q_AN02 U512 ( .A0(n41), .A1(gcm_dak_cmd_in[595]), .Z(n159));
Q_MX02 U513 ( .S(n39), .A0(gcm_dek_cmd_in[594]), .A1(n160), .Z(gcm_cmd_in[594]));
Q_AN02 U514 ( .A0(n41), .A1(gcm_dak_cmd_in[594]), .Z(n160));
Q_MX02 U515 ( .S(n39), .A0(gcm_dek_cmd_in[593]), .A1(n161), .Z(gcm_cmd_in[593]));
Q_AN02 U516 ( .A0(n41), .A1(gcm_dak_cmd_in[593]), .Z(n161));
Q_MX02 U517 ( .S(n39), .A0(gcm_dek_cmd_in[592]), .A1(n162), .Z(gcm_cmd_in[592]));
Q_AN02 U518 ( .A0(n41), .A1(gcm_dak_cmd_in[592]), .Z(n162));
Q_MX02 U519 ( .S(n39), .A0(gcm_dek_cmd_in[591]), .A1(n163), .Z(gcm_cmd_in[591]));
Q_AN02 U520 ( .A0(n41), .A1(gcm_dak_cmd_in[591]), .Z(n163));
Q_MX02 U521 ( .S(n39), .A0(gcm_dek_cmd_in[590]), .A1(n164), .Z(gcm_cmd_in[590]));
Q_AN02 U522 ( .A0(n41), .A1(gcm_dak_cmd_in[590]), .Z(n164));
Q_MX02 U523 ( .S(n39), .A0(gcm_dek_cmd_in[589]), .A1(n165), .Z(gcm_cmd_in[589]));
Q_AN02 U524 ( .A0(n41), .A1(gcm_dak_cmd_in[589]), .Z(n165));
Q_MX02 U525 ( .S(n39), .A0(gcm_dek_cmd_in[588]), .A1(n166), .Z(gcm_cmd_in[588]));
Q_AN02 U526 ( .A0(n41), .A1(gcm_dak_cmd_in[588]), .Z(n166));
Q_MX02 U527 ( .S(n39), .A0(gcm_dek_cmd_in[587]), .A1(n167), .Z(gcm_cmd_in[587]));
Q_AN02 U528 ( .A0(n41), .A1(gcm_dak_cmd_in[587]), .Z(n167));
Q_MX02 U529 ( .S(n39), .A0(gcm_dek_cmd_in[586]), .A1(n168), .Z(gcm_cmd_in[586]));
Q_AN02 U530 ( .A0(n41), .A1(gcm_dak_cmd_in[586]), .Z(n168));
Q_MX02 U531 ( .S(n39), .A0(gcm_dek_cmd_in[585]), .A1(n169), .Z(gcm_cmd_in[585]));
Q_AN02 U532 ( .A0(n41), .A1(gcm_dak_cmd_in[585]), .Z(n169));
Q_MX02 U533 ( .S(n39), .A0(gcm_dek_cmd_in[584]), .A1(n170), .Z(gcm_cmd_in[584]));
Q_AN02 U534 ( .A0(n41), .A1(gcm_dak_cmd_in[584]), .Z(n170));
Q_MX02 U535 ( .S(n39), .A0(gcm_dek_cmd_in[583]), .A1(n171), .Z(gcm_cmd_in[583]));
Q_AN02 U536 ( .A0(n41), .A1(gcm_dak_cmd_in[583]), .Z(n171));
Q_MX02 U537 ( .S(n39), .A0(gcm_dek_cmd_in[582]), .A1(n172), .Z(gcm_cmd_in[582]));
Q_AN02 U538 ( .A0(n41), .A1(gcm_dak_cmd_in[582]), .Z(n172));
Q_MX02 U539 ( .S(n39), .A0(gcm_dek_cmd_in[581]), .A1(n173), .Z(gcm_cmd_in[581]));
Q_AN02 U540 ( .A0(n41), .A1(gcm_dak_cmd_in[581]), .Z(n173));
Q_MX02 U541 ( .S(n39), .A0(gcm_dek_cmd_in[580]), .A1(n174), .Z(gcm_cmd_in[580]));
Q_AN02 U542 ( .A0(n41), .A1(gcm_dak_cmd_in[580]), .Z(n174));
Q_MX02 U543 ( .S(n39), .A0(gcm_dek_cmd_in[579]), .A1(n175), .Z(gcm_cmd_in[579]));
Q_AN02 U544 ( .A0(n41), .A1(gcm_dak_cmd_in[579]), .Z(n175));
Q_MX02 U545 ( .S(n39), .A0(gcm_dek_cmd_in[578]), .A1(n176), .Z(gcm_cmd_in[578]));
Q_AN02 U546 ( .A0(n41), .A1(gcm_dak_cmd_in[578]), .Z(n176));
Q_MX02 U547 ( .S(n39), .A0(gcm_dek_cmd_in[577]), .A1(n177), .Z(gcm_cmd_in[577]));
Q_AN02 U548 ( .A0(n41), .A1(gcm_dak_cmd_in[577]), .Z(n177));
Q_MX02 U549 ( .S(n39), .A0(gcm_dek_cmd_in[576]), .A1(n178), .Z(gcm_cmd_in[576]));
Q_AN02 U550 ( .A0(n41), .A1(gcm_dak_cmd_in[576]), .Z(n178));
Q_MX02 U551 ( .S(n39), .A0(gcm_dek_cmd_in[575]), .A1(n179), .Z(gcm_cmd_in[575]));
Q_AN02 U552 ( .A0(n41), .A1(gcm_dak_cmd_in[575]), .Z(n179));
Q_MX02 U553 ( .S(n39), .A0(gcm_dek_cmd_in[574]), .A1(n180), .Z(gcm_cmd_in[574]));
Q_AN02 U554 ( .A0(n41), .A1(gcm_dak_cmd_in[574]), .Z(n180));
Q_MX02 U555 ( .S(n39), .A0(gcm_dek_cmd_in[573]), .A1(n181), .Z(gcm_cmd_in[573]));
Q_AN02 U556 ( .A0(n41), .A1(gcm_dak_cmd_in[573]), .Z(n181));
Q_MX02 U557 ( .S(n39), .A0(gcm_dek_cmd_in[572]), .A1(n182), .Z(gcm_cmd_in[572]));
Q_AN02 U558 ( .A0(n41), .A1(gcm_dak_cmd_in[572]), .Z(n182));
Q_MX02 U559 ( .S(n39), .A0(gcm_dek_cmd_in[571]), .A1(n183), .Z(gcm_cmd_in[571]));
Q_AN02 U560 ( .A0(n41), .A1(gcm_dak_cmd_in[571]), .Z(n183));
Q_MX02 U561 ( .S(n39), .A0(gcm_dek_cmd_in[570]), .A1(n184), .Z(gcm_cmd_in[570]));
Q_AN02 U562 ( .A0(n41), .A1(gcm_dak_cmd_in[570]), .Z(n184));
Q_MX02 U563 ( .S(n39), .A0(gcm_dek_cmd_in[569]), .A1(n185), .Z(gcm_cmd_in[569]));
Q_AN02 U564 ( .A0(n41), .A1(gcm_dak_cmd_in[569]), .Z(n185));
Q_MX02 U565 ( .S(n39), .A0(gcm_dek_cmd_in[568]), .A1(n186), .Z(gcm_cmd_in[568]));
Q_AN02 U566 ( .A0(n41), .A1(gcm_dak_cmd_in[568]), .Z(n186));
Q_MX02 U567 ( .S(n39), .A0(gcm_dek_cmd_in[567]), .A1(n187), .Z(gcm_cmd_in[567]));
Q_AN02 U568 ( .A0(n41), .A1(gcm_dak_cmd_in[567]), .Z(n187));
Q_MX02 U569 ( .S(n39), .A0(gcm_dek_cmd_in[566]), .A1(n188), .Z(gcm_cmd_in[566]));
Q_AN02 U570 ( .A0(n41), .A1(gcm_dak_cmd_in[566]), .Z(n188));
Q_MX02 U571 ( .S(n39), .A0(gcm_dek_cmd_in[565]), .A1(n189), .Z(gcm_cmd_in[565]));
Q_AN02 U572 ( .A0(n41), .A1(gcm_dak_cmd_in[565]), .Z(n189));
Q_MX02 U573 ( .S(n39), .A0(gcm_dek_cmd_in[564]), .A1(n190), .Z(gcm_cmd_in[564]));
Q_AN02 U574 ( .A0(n41), .A1(gcm_dak_cmd_in[564]), .Z(n190));
Q_MX02 U575 ( .S(n39), .A0(gcm_dek_cmd_in[563]), .A1(n191), .Z(gcm_cmd_in[563]));
Q_AN02 U576 ( .A0(n41), .A1(gcm_dak_cmd_in[563]), .Z(n191));
Q_MX02 U577 ( .S(n39), .A0(gcm_dek_cmd_in[562]), .A1(n192), .Z(gcm_cmd_in[562]));
Q_AN02 U578 ( .A0(n41), .A1(gcm_dak_cmd_in[562]), .Z(n192));
Q_MX02 U579 ( .S(n39), .A0(gcm_dek_cmd_in[561]), .A1(n193), .Z(gcm_cmd_in[561]));
Q_AN02 U580 ( .A0(n41), .A1(gcm_dak_cmd_in[561]), .Z(n193));
Q_MX02 U581 ( .S(n39), .A0(gcm_dek_cmd_in[560]), .A1(n194), .Z(gcm_cmd_in[560]));
Q_AN02 U582 ( .A0(n41), .A1(gcm_dak_cmd_in[560]), .Z(n194));
Q_MX02 U583 ( .S(n39), .A0(gcm_dek_cmd_in[559]), .A1(n195), .Z(gcm_cmd_in[559]));
Q_AN02 U584 ( .A0(n41), .A1(gcm_dak_cmd_in[559]), .Z(n195));
Q_MX02 U585 ( .S(n39), .A0(gcm_dek_cmd_in[558]), .A1(n196), .Z(gcm_cmd_in[558]));
Q_AN02 U586 ( .A0(n41), .A1(gcm_dak_cmd_in[558]), .Z(n196));
Q_MX02 U587 ( .S(n39), .A0(gcm_dek_cmd_in[557]), .A1(n197), .Z(gcm_cmd_in[557]));
Q_AN02 U588 ( .A0(n41), .A1(gcm_dak_cmd_in[557]), .Z(n197));
Q_MX02 U589 ( .S(n39), .A0(gcm_dek_cmd_in[556]), .A1(n198), .Z(gcm_cmd_in[556]));
Q_AN02 U590 ( .A0(n41), .A1(gcm_dak_cmd_in[556]), .Z(n198));
Q_MX02 U591 ( .S(n39), .A0(gcm_dek_cmd_in[555]), .A1(n199), .Z(gcm_cmd_in[555]));
Q_AN02 U592 ( .A0(n41), .A1(gcm_dak_cmd_in[555]), .Z(n199));
Q_MX02 U593 ( .S(n39), .A0(gcm_dek_cmd_in[554]), .A1(n200), .Z(gcm_cmd_in[554]));
Q_AN02 U594 ( .A0(n41), .A1(gcm_dak_cmd_in[554]), .Z(n200));
Q_MX02 U595 ( .S(n39), .A0(gcm_dek_cmd_in[553]), .A1(n201), .Z(gcm_cmd_in[553]));
Q_AN02 U596 ( .A0(n41), .A1(gcm_dak_cmd_in[553]), .Z(n201));
Q_MX02 U597 ( .S(n39), .A0(gcm_dek_cmd_in[552]), .A1(n202), .Z(gcm_cmd_in[552]));
Q_AN02 U598 ( .A0(n41), .A1(gcm_dak_cmd_in[552]), .Z(n202));
Q_MX02 U599 ( .S(n39), .A0(gcm_dek_cmd_in[551]), .A1(n203), .Z(gcm_cmd_in[551]));
Q_AN02 U600 ( .A0(n41), .A1(gcm_dak_cmd_in[551]), .Z(n203));
Q_MX02 U601 ( .S(n39), .A0(gcm_dek_cmd_in[550]), .A1(n204), .Z(gcm_cmd_in[550]));
Q_AN02 U602 ( .A0(n41), .A1(gcm_dak_cmd_in[550]), .Z(n204));
Q_MX02 U603 ( .S(n39), .A0(gcm_dek_cmd_in[549]), .A1(n205), .Z(gcm_cmd_in[549]));
Q_AN02 U604 ( .A0(n41), .A1(gcm_dak_cmd_in[549]), .Z(n205));
Q_MX02 U605 ( .S(n39), .A0(gcm_dek_cmd_in[548]), .A1(n206), .Z(gcm_cmd_in[548]));
Q_AN02 U606 ( .A0(n41), .A1(gcm_dak_cmd_in[548]), .Z(n206));
Q_MX02 U607 ( .S(n39), .A0(gcm_dek_cmd_in[547]), .A1(n207), .Z(gcm_cmd_in[547]));
Q_AN02 U608 ( .A0(n41), .A1(gcm_dak_cmd_in[547]), .Z(n207));
Q_MX02 U609 ( .S(n39), .A0(gcm_dek_cmd_in[546]), .A1(n208), .Z(gcm_cmd_in[546]));
Q_AN02 U610 ( .A0(n41), .A1(gcm_dak_cmd_in[546]), .Z(n208));
Q_MX02 U611 ( .S(n39), .A0(gcm_dek_cmd_in[545]), .A1(n209), .Z(gcm_cmd_in[545]));
Q_AN02 U612 ( .A0(n41), .A1(gcm_dak_cmd_in[545]), .Z(n209));
Q_MX02 U613 ( .S(n39), .A0(gcm_dek_cmd_in[544]), .A1(n210), .Z(gcm_cmd_in[544]));
Q_AN02 U614 ( .A0(n41), .A1(gcm_dak_cmd_in[544]), .Z(n210));
Q_MX02 U615 ( .S(n39), .A0(gcm_dek_cmd_in[543]), .A1(n211), .Z(gcm_cmd_in[543]));
Q_AN02 U616 ( .A0(n41), .A1(gcm_dak_cmd_in[543]), .Z(n211));
Q_MX02 U617 ( .S(n39), .A0(gcm_dek_cmd_in[542]), .A1(n212), .Z(gcm_cmd_in[542]));
Q_AN02 U618 ( .A0(n41), .A1(gcm_dak_cmd_in[542]), .Z(n212));
Q_MX02 U619 ( .S(n39), .A0(gcm_dek_cmd_in[541]), .A1(n213), .Z(gcm_cmd_in[541]));
Q_AN02 U620 ( .A0(n41), .A1(gcm_dak_cmd_in[541]), .Z(n213));
Q_MX02 U621 ( .S(n39), .A0(gcm_dek_cmd_in[540]), .A1(n214), .Z(gcm_cmd_in[540]));
Q_AN02 U622 ( .A0(n41), .A1(gcm_dak_cmd_in[540]), .Z(n214));
Q_MX02 U623 ( .S(n39), .A0(gcm_dek_cmd_in[539]), .A1(n215), .Z(gcm_cmd_in[539]));
Q_AN02 U624 ( .A0(n41), .A1(gcm_dak_cmd_in[539]), .Z(n215));
Q_MX02 U625 ( .S(n39), .A0(gcm_dek_cmd_in[538]), .A1(n216), .Z(gcm_cmd_in[538]));
Q_AN02 U626 ( .A0(n41), .A1(gcm_dak_cmd_in[538]), .Z(n216));
Q_MX02 U627 ( .S(n39), .A0(gcm_dek_cmd_in[537]), .A1(n217), .Z(gcm_cmd_in[537]));
Q_AN02 U628 ( .A0(n41), .A1(gcm_dak_cmd_in[537]), .Z(n217));
Q_MX02 U629 ( .S(n39), .A0(gcm_dek_cmd_in[536]), .A1(n218), .Z(gcm_cmd_in[536]));
Q_AN02 U630 ( .A0(n41), .A1(gcm_dak_cmd_in[536]), .Z(n218));
Q_MX02 U631 ( .S(n39), .A0(gcm_dek_cmd_in[535]), .A1(n219), .Z(gcm_cmd_in[535]));
Q_AN02 U632 ( .A0(n41), .A1(gcm_dak_cmd_in[535]), .Z(n219));
Q_MX02 U633 ( .S(n39), .A0(gcm_dek_cmd_in[534]), .A1(n220), .Z(gcm_cmd_in[534]));
Q_AN02 U634 ( .A0(n41), .A1(gcm_dak_cmd_in[534]), .Z(n220));
Q_MX02 U635 ( .S(n39), .A0(gcm_dek_cmd_in[533]), .A1(n221), .Z(gcm_cmd_in[533]));
Q_AN02 U636 ( .A0(n41), .A1(gcm_dak_cmd_in[533]), .Z(n221));
Q_MX02 U637 ( .S(n39), .A0(gcm_dek_cmd_in[532]), .A1(n222), .Z(gcm_cmd_in[532]));
Q_AN02 U638 ( .A0(n41), .A1(gcm_dak_cmd_in[532]), .Z(n222));
Q_MX02 U639 ( .S(n39), .A0(gcm_dek_cmd_in[531]), .A1(n223), .Z(gcm_cmd_in[531]));
Q_AN02 U640 ( .A0(n41), .A1(gcm_dak_cmd_in[531]), .Z(n223));
Q_MX02 U641 ( .S(n39), .A0(gcm_dek_cmd_in[530]), .A1(n224), .Z(gcm_cmd_in[530]));
Q_AN02 U642 ( .A0(n41), .A1(gcm_dak_cmd_in[530]), .Z(n224));
Q_MX02 U643 ( .S(n39), .A0(gcm_dek_cmd_in[529]), .A1(n225), .Z(gcm_cmd_in[529]));
Q_AN02 U644 ( .A0(n41), .A1(gcm_dak_cmd_in[529]), .Z(n225));
Q_MX02 U645 ( .S(n39), .A0(gcm_dek_cmd_in[528]), .A1(n226), .Z(gcm_cmd_in[528]));
Q_AN02 U646 ( .A0(n41), .A1(gcm_dak_cmd_in[528]), .Z(n226));
Q_MX02 U647 ( .S(n39), .A0(gcm_dek_cmd_in[527]), .A1(n227), .Z(gcm_cmd_in[527]));
Q_AN02 U648 ( .A0(n41), .A1(gcm_dak_cmd_in[527]), .Z(n227));
Q_MX02 U649 ( .S(n39), .A0(gcm_dek_cmd_in[526]), .A1(n228), .Z(gcm_cmd_in[526]));
Q_AN02 U650 ( .A0(n41), .A1(gcm_dak_cmd_in[526]), .Z(n228));
Q_MX02 U651 ( .S(n39), .A0(gcm_dek_cmd_in[525]), .A1(n229), .Z(gcm_cmd_in[525]));
Q_AN02 U652 ( .A0(n41), .A1(gcm_dak_cmd_in[525]), .Z(n229));
Q_MX02 U653 ( .S(n39), .A0(gcm_dek_cmd_in[524]), .A1(n230), .Z(gcm_cmd_in[524]));
Q_AN02 U654 ( .A0(n41), .A1(gcm_dak_cmd_in[524]), .Z(n230));
Q_MX02 U655 ( .S(n39), .A0(gcm_dek_cmd_in[523]), .A1(n231), .Z(gcm_cmd_in[523]));
Q_AN02 U656 ( .A0(n41), .A1(gcm_dak_cmd_in[523]), .Z(n231));
Q_MX02 U657 ( .S(n39), .A0(gcm_dek_cmd_in[522]), .A1(n232), .Z(gcm_cmd_in[522]));
Q_AN02 U658 ( .A0(n41), .A1(gcm_dak_cmd_in[522]), .Z(n232));
Q_MX02 U659 ( .S(n39), .A0(gcm_dek_cmd_in[521]), .A1(n233), .Z(gcm_cmd_in[521]));
Q_AN02 U660 ( .A0(n41), .A1(gcm_dak_cmd_in[521]), .Z(n233));
Q_MX02 U661 ( .S(n39), .A0(gcm_dek_cmd_in[520]), .A1(n234), .Z(gcm_cmd_in[520]));
Q_AN02 U662 ( .A0(n41), .A1(gcm_dak_cmd_in[520]), .Z(n234));
Q_MX02 U663 ( .S(n39), .A0(gcm_dek_cmd_in[519]), .A1(n235), .Z(gcm_cmd_in[519]));
Q_AN02 U664 ( .A0(n41), .A1(gcm_dak_cmd_in[519]), .Z(n235));
Q_MX02 U665 ( .S(n39), .A0(gcm_dek_cmd_in[518]), .A1(n236), .Z(gcm_cmd_in[518]));
Q_AN02 U666 ( .A0(n41), .A1(gcm_dak_cmd_in[518]), .Z(n236));
Q_MX02 U667 ( .S(n39), .A0(gcm_dek_cmd_in[517]), .A1(n237), .Z(gcm_cmd_in[517]));
Q_AN02 U668 ( .A0(n41), .A1(gcm_dak_cmd_in[517]), .Z(n237));
Q_MX02 U669 ( .S(n39), .A0(gcm_dek_cmd_in[516]), .A1(n238), .Z(gcm_cmd_in[516]));
Q_AN02 U670 ( .A0(n41), .A1(gcm_dak_cmd_in[516]), .Z(n238));
Q_MX02 U671 ( .S(n39), .A0(gcm_dek_cmd_in[515]), .A1(n239), .Z(gcm_cmd_in[515]));
Q_AN02 U672 ( .A0(n41), .A1(gcm_dak_cmd_in[515]), .Z(n239));
Q_MX02 U673 ( .S(n39), .A0(gcm_dek_cmd_in[514]), .A1(n240), .Z(gcm_cmd_in[514]));
Q_AN02 U674 ( .A0(n41), .A1(gcm_dak_cmd_in[514]), .Z(n240));
Q_MX02 U675 ( .S(n39), .A0(gcm_dek_cmd_in[513]), .A1(n241), .Z(gcm_cmd_in[513]));
Q_AN02 U676 ( .A0(n41), .A1(gcm_dak_cmd_in[513]), .Z(n241));
Q_MX02 U677 ( .S(n39), .A0(gcm_dek_cmd_in[512]), .A1(n242), .Z(gcm_cmd_in[512]));
Q_AN02 U678 ( .A0(n41), .A1(gcm_dak_cmd_in[512]), .Z(n242));
Q_MX02 U679 ( .S(n39), .A0(gcm_dek_cmd_in[511]), .A1(n243), .Z(gcm_cmd_in[511]));
Q_AN02 U680 ( .A0(n41), .A1(gcm_dak_cmd_in[511]), .Z(n243));
Q_MX02 U681 ( .S(n39), .A0(gcm_dek_cmd_in[510]), .A1(n244), .Z(gcm_cmd_in[510]));
Q_AN02 U682 ( .A0(n41), .A1(gcm_dak_cmd_in[510]), .Z(n244));
Q_MX02 U683 ( .S(n39), .A0(gcm_dek_cmd_in[509]), .A1(n245), .Z(gcm_cmd_in[509]));
Q_AN02 U684 ( .A0(n41), .A1(gcm_dak_cmd_in[509]), .Z(n245));
Q_MX02 U685 ( .S(n39), .A0(gcm_dek_cmd_in[508]), .A1(n246), .Z(gcm_cmd_in[508]));
Q_AN02 U686 ( .A0(n41), .A1(gcm_dak_cmd_in[508]), .Z(n246));
Q_MX02 U687 ( .S(n39), .A0(gcm_dek_cmd_in[507]), .A1(n247), .Z(gcm_cmd_in[507]));
Q_AN02 U688 ( .A0(n41), .A1(gcm_dak_cmd_in[507]), .Z(n247));
Q_MX02 U689 ( .S(n39), .A0(gcm_dek_cmd_in[506]), .A1(n248), .Z(gcm_cmd_in[506]));
Q_AN02 U690 ( .A0(n41), .A1(gcm_dak_cmd_in[506]), .Z(n248));
Q_MX02 U691 ( .S(n39), .A0(gcm_dek_cmd_in[505]), .A1(n249), .Z(gcm_cmd_in[505]));
Q_AN02 U692 ( .A0(n41), .A1(gcm_dak_cmd_in[505]), .Z(n249));
Q_MX02 U693 ( .S(n39), .A0(gcm_dek_cmd_in[504]), .A1(n250), .Z(gcm_cmd_in[504]));
Q_AN02 U694 ( .A0(n41), .A1(gcm_dak_cmd_in[504]), .Z(n250));
Q_MX02 U695 ( .S(n39), .A0(gcm_dek_cmd_in[503]), .A1(n251), .Z(gcm_cmd_in[503]));
Q_AN02 U696 ( .A0(n41), .A1(gcm_dak_cmd_in[503]), .Z(n251));
Q_MX02 U697 ( .S(n39), .A0(gcm_dek_cmd_in[502]), .A1(n252), .Z(gcm_cmd_in[502]));
Q_AN02 U698 ( .A0(n41), .A1(gcm_dak_cmd_in[502]), .Z(n252));
Q_MX02 U699 ( .S(n39), .A0(gcm_dek_cmd_in[501]), .A1(n253), .Z(gcm_cmd_in[501]));
Q_AN02 U700 ( .A0(n41), .A1(gcm_dak_cmd_in[501]), .Z(n253));
Q_MX02 U701 ( .S(n39), .A0(gcm_dek_cmd_in[500]), .A1(n254), .Z(gcm_cmd_in[500]));
Q_AN02 U702 ( .A0(n41), .A1(gcm_dak_cmd_in[500]), .Z(n254));
Q_MX02 U703 ( .S(n39), .A0(gcm_dek_cmd_in[499]), .A1(n255), .Z(gcm_cmd_in[499]));
Q_AN02 U704 ( .A0(n41), .A1(gcm_dak_cmd_in[499]), .Z(n255));
Q_MX02 U705 ( .S(n39), .A0(gcm_dek_cmd_in[498]), .A1(n256), .Z(gcm_cmd_in[498]));
Q_AN02 U706 ( .A0(n41), .A1(gcm_dak_cmd_in[498]), .Z(n256));
Q_MX02 U707 ( .S(n39), .A0(gcm_dek_cmd_in[497]), .A1(n257), .Z(gcm_cmd_in[497]));
Q_AN02 U708 ( .A0(n41), .A1(gcm_dak_cmd_in[497]), .Z(n257));
Q_MX02 U709 ( .S(n39), .A0(gcm_dek_cmd_in[496]), .A1(n258), .Z(gcm_cmd_in[496]));
Q_AN02 U710 ( .A0(n41), .A1(gcm_dak_cmd_in[496]), .Z(n258));
Q_MX02 U711 ( .S(n39), .A0(gcm_dek_cmd_in[495]), .A1(n259), .Z(gcm_cmd_in[495]));
Q_AN02 U712 ( .A0(n41), .A1(gcm_dak_cmd_in[495]), .Z(n259));
Q_MX02 U713 ( .S(n39), .A0(gcm_dek_cmd_in[494]), .A1(n260), .Z(gcm_cmd_in[494]));
Q_AN02 U714 ( .A0(n41), .A1(gcm_dak_cmd_in[494]), .Z(n260));
Q_MX02 U715 ( .S(n39), .A0(gcm_dek_cmd_in[493]), .A1(n261), .Z(gcm_cmd_in[493]));
Q_AN02 U716 ( .A0(n41), .A1(gcm_dak_cmd_in[493]), .Z(n261));
Q_MX02 U717 ( .S(n39), .A0(gcm_dek_cmd_in[492]), .A1(n262), .Z(gcm_cmd_in[492]));
Q_AN02 U718 ( .A0(n41), .A1(gcm_dak_cmd_in[492]), .Z(n262));
Q_MX02 U719 ( .S(n39), .A0(gcm_dek_cmd_in[491]), .A1(n263), .Z(gcm_cmd_in[491]));
Q_AN02 U720 ( .A0(n41), .A1(gcm_dak_cmd_in[491]), .Z(n263));
Q_MX02 U721 ( .S(n39), .A0(gcm_dek_cmd_in[490]), .A1(n264), .Z(gcm_cmd_in[490]));
Q_AN02 U722 ( .A0(n41), .A1(gcm_dak_cmd_in[490]), .Z(n264));
Q_MX02 U723 ( .S(n39), .A0(gcm_dek_cmd_in[489]), .A1(n265), .Z(gcm_cmd_in[489]));
Q_AN02 U724 ( .A0(n41), .A1(gcm_dak_cmd_in[489]), .Z(n265));
Q_MX02 U725 ( .S(n39), .A0(gcm_dek_cmd_in[488]), .A1(n266), .Z(gcm_cmd_in[488]));
Q_AN02 U726 ( .A0(n41), .A1(gcm_dak_cmd_in[488]), .Z(n266));
Q_MX02 U727 ( .S(n39), .A0(gcm_dek_cmd_in[487]), .A1(n267), .Z(gcm_cmd_in[487]));
Q_AN02 U728 ( .A0(n41), .A1(gcm_dak_cmd_in[487]), .Z(n267));
Q_MX02 U729 ( .S(n39), .A0(gcm_dek_cmd_in[486]), .A1(n268), .Z(gcm_cmd_in[486]));
Q_AN02 U730 ( .A0(n41), .A1(gcm_dak_cmd_in[486]), .Z(n268));
Q_MX02 U731 ( .S(n39), .A0(gcm_dek_cmd_in[485]), .A1(n269), .Z(gcm_cmd_in[485]));
Q_AN02 U732 ( .A0(n41), .A1(gcm_dak_cmd_in[485]), .Z(n269));
Q_MX02 U733 ( .S(n39), .A0(gcm_dek_cmd_in[484]), .A1(n270), .Z(gcm_cmd_in[484]));
Q_AN02 U734 ( .A0(n41), .A1(gcm_dak_cmd_in[484]), .Z(n270));
Q_MX02 U735 ( .S(n39), .A0(gcm_dek_cmd_in[483]), .A1(n271), .Z(gcm_cmd_in[483]));
Q_AN02 U736 ( .A0(n41), .A1(gcm_dak_cmd_in[483]), .Z(n271));
Q_MX02 U737 ( .S(n39), .A0(gcm_dek_cmd_in[482]), .A1(n272), .Z(gcm_cmd_in[482]));
Q_AN02 U738 ( .A0(n41), .A1(gcm_dak_cmd_in[482]), .Z(n272));
Q_MX02 U739 ( .S(n39), .A0(gcm_dek_cmd_in[481]), .A1(n273), .Z(gcm_cmd_in[481]));
Q_AN02 U740 ( .A0(n41), .A1(gcm_dak_cmd_in[481]), .Z(n273));
Q_MX02 U741 ( .S(n39), .A0(gcm_dek_cmd_in[480]), .A1(n274), .Z(gcm_cmd_in[480]));
Q_AN02 U742 ( .A0(n41), .A1(gcm_dak_cmd_in[480]), .Z(n274));
Q_MX02 U743 ( .S(n39), .A0(gcm_dek_cmd_in[479]), .A1(n275), .Z(gcm_cmd_in[479]));
Q_AN02 U744 ( .A0(n41), .A1(gcm_dak_cmd_in[479]), .Z(n275));
Q_MX02 U745 ( .S(n39), .A0(gcm_dek_cmd_in[478]), .A1(n276), .Z(gcm_cmd_in[478]));
Q_AN02 U746 ( .A0(n41), .A1(gcm_dak_cmd_in[478]), .Z(n276));
Q_MX02 U747 ( .S(n39), .A0(gcm_dek_cmd_in[477]), .A1(n277), .Z(gcm_cmd_in[477]));
Q_AN02 U748 ( .A0(n41), .A1(gcm_dak_cmd_in[477]), .Z(n277));
Q_MX02 U749 ( .S(n39), .A0(gcm_dek_cmd_in[476]), .A1(n278), .Z(gcm_cmd_in[476]));
Q_AN02 U750 ( .A0(n41), .A1(gcm_dak_cmd_in[476]), .Z(n278));
Q_MX02 U751 ( .S(n39), .A0(gcm_dek_cmd_in[475]), .A1(n279), .Z(gcm_cmd_in[475]));
Q_AN02 U752 ( .A0(n41), .A1(gcm_dak_cmd_in[475]), .Z(n279));
Q_MX02 U753 ( .S(n39), .A0(gcm_dek_cmd_in[474]), .A1(n280), .Z(gcm_cmd_in[474]));
Q_AN02 U754 ( .A0(n41), .A1(gcm_dak_cmd_in[474]), .Z(n280));
Q_MX02 U755 ( .S(n39), .A0(gcm_dek_cmd_in[473]), .A1(n281), .Z(gcm_cmd_in[473]));
Q_AN02 U756 ( .A0(n41), .A1(gcm_dak_cmd_in[473]), .Z(n281));
Q_MX02 U757 ( .S(n39), .A0(gcm_dek_cmd_in[472]), .A1(n282), .Z(gcm_cmd_in[472]));
Q_AN02 U758 ( .A0(n41), .A1(gcm_dak_cmd_in[472]), .Z(n282));
Q_MX02 U759 ( .S(n39), .A0(gcm_dek_cmd_in[471]), .A1(n283), .Z(gcm_cmd_in[471]));
Q_AN02 U760 ( .A0(n41), .A1(gcm_dak_cmd_in[471]), .Z(n283));
Q_MX02 U761 ( .S(n39), .A0(gcm_dek_cmd_in[470]), .A1(n284), .Z(gcm_cmd_in[470]));
Q_AN02 U762 ( .A0(n41), .A1(gcm_dak_cmd_in[470]), .Z(n284));
Q_MX02 U763 ( .S(n39), .A0(gcm_dek_cmd_in[469]), .A1(n285), .Z(gcm_cmd_in[469]));
Q_AN02 U764 ( .A0(n41), .A1(gcm_dak_cmd_in[469]), .Z(n285));
Q_MX02 U765 ( .S(n39), .A0(gcm_dek_cmd_in[468]), .A1(n286), .Z(gcm_cmd_in[468]));
Q_AN02 U766 ( .A0(n41), .A1(gcm_dak_cmd_in[468]), .Z(n286));
Q_MX02 U767 ( .S(n39), .A0(gcm_dek_cmd_in[467]), .A1(n287), .Z(gcm_cmd_in[467]));
Q_AN02 U768 ( .A0(n41), .A1(gcm_dak_cmd_in[467]), .Z(n287));
Q_MX02 U769 ( .S(n39), .A0(gcm_dek_cmd_in[466]), .A1(n288), .Z(gcm_cmd_in[466]));
Q_AN02 U770 ( .A0(n41), .A1(gcm_dak_cmd_in[466]), .Z(n288));
Q_MX02 U771 ( .S(n39), .A0(gcm_dek_cmd_in[465]), .A1(n289), .Z(gcm_cmd_in[465]));
Q_AN02 U772 ( .A0(n41), .A1(gcm_dak_cmd_in[465]), .Z(n289));
Q_MX02 U773 ( .S(n39), .A0(gcm_dek_cmd_in[464]), .A1(n290), .Z(gcm_cmd_in[464]));
Q_AN02 U774 ( .A0(n41), .A1(gcm_dak_cmd_in[464]), .Z(n290));
Q_MX02 U775 ( .S(n39), .A0(gcm_dek_cmd_in[463]), .A1(n291), .Z(gcm_cmd_in[463]));
Q_AN02 U776 ( .A0(n41), .A1(gcm_dak_cmd_in[463]), .Z(n291));
Q_MX02 U777 ( .S(n39), .A0(gcm_dek_cmd_in[462]), .A1(n292), .Z(gcm_cmd_in[462]));
Q_AN02 U778 ( .A0(n41), .A1(gcm_dak_cmd_in[462]), .Z(n292));
Q_MX02 U779 ( .S(n39), .A0(gcm_dek_cmd_in[461]), .A1(n293), .Z(gcm_cmd_in[461]));
Q_AN02 U780 ( .A0(n41), .A1(gcm_dak_cmd_in[461]), .Z(n293));
Q_MX02 U781 ( .S(n39), .A0(gcm_dek_cmd_in[460]), .A1(n294), .Z(gcm_cmd_in[460]));
Q_AN02 U782 ( .A0(n41), .A1(gcm_dak_cmd_in[460]), .Z(n294));
Q_MX02 U783 ( .S(n39), .A0(gcm_dek_cmd_in[459]), .A1(n295), .Z(gcm_cmd_in[459]));
Q_AN02 U784 ( .A0(n41), .A1(gcm_dak_cmd_in[459]), .Z(n295));
Q_MX02 U785 ( .S(n39), .A0(gcm_dek_cmd_in[458]), .A1(n296), .Z(gcm_cmd_in[458]));
Q_AN02 U786 ( .A0(n41), .A1(gcm_dak_cmd_in[458]), .Z(n296));
Q_MX02 U787 ( .S(n39), .A0(gcm_dek_cmd_in[457]), .A1(n297), .Z(gcm_cmd_in[457]));
Q_AN02 U788 ( .A0(n41), .A1(gcm_dak_cmd_in[457]), .Z(n297));
Q_MX02 U789 ( .S(n39), .A0(gcm_dek_cmd_in[456]), .A1(n298), .Z(gcm_cmd_in[456]));
Q_AN02 U790 ( .A0(n41), .A1(gcm_dak_cmd_in[456]), .Z(n298));
Q_MX02 U791 ( .S(n39), .A0(gcm_dek_cmd_in[455]), .A1(n299), .Z(gcm_cmd_in[455]));
Q_AN02 U792 ( .A0(n41), .A1(gcm_dak_cmd_in[455]), .Z(n299));
Q_MX02 U793 ( .S(n39), .A0(gcm_dek_cmd_in[454]), .A1(n300), .Z(gcm_cmd_in[454]));
Q_AN02 U794 ( .A0(n41), .A1(gcm_dak_cmd_in[454]), .Z(n300));
Q_MX02 U795 ( .S(n39), .A0(gcm_dek_cmd_in[453]), .A1(n301), .Z(gcm_cmd_in[453]));
Q_AN02 U796 ( .A0(n41), .A1(gcm_dak_cmd_in[453]), .Z(n301));
Q_MX02 U797 ( .S(n39), .A0(gcm_dek_cmd_in[452]), .A1(n302), .Z(gcm_cmd_in[452]));
Q_AN02 U798 ( .A0(n41), .A1(gcm_dak_cmd_in[452]), .Z(n302));
Q_MX02 U799 ( .S(n39), .A0(gcm_dek_cmd_in[451]), .A1(n303), .Z(gcm_cmd_in[451]));
Q_AN02 U800 ( .A0(n41), .A1(gcm_dak_cmd_in[451]), .Z(n303));
Q_MX02 U801 ( .S(n39), .A0(gcm_dek_cmd_in[450]), .A1(n304), .Z(gcm_cmd_in[450]));
Q_AN02 U802 ( .A0(n41), .A1(gcm_dak_cmd_in[450]), .Z(n304));
Q_MX02 U803 ( .S(n39), .A0(gcm_dek_cmd_in[449]), .A1(n305), .Z(gcm_cmd_in[449]));
Q_AN02 U804 ( .A0(n41), .A1(gcm_dak_cmd_in[449]), .Z(n305));
Q_MX02 U805 ( .S(n39), .A0(gcm_dek_cmd_in[448]), .A1(n306), .Z(gcm_cmd_in[448]));
Q_AN02 U806 ( .A0(n41), .A1(gcm_dak_cmd_in[448]), .Z(n306));
Q_MX02 U807 ( .S(n39), .A0(gcm_dek_cmd_in[447]), .A1(n307), .Z(gcm_cmd_in[447]));
Q_AN02 U808 ( .A0(n41), .A1(gcm_dak_cmd_in[447]), .Z(n307));
Q_MX02 U809 ( .S(n39), .A0(gcm_dek_cmd_in[446]), .A1(n308), .Z(gcm_cmd_in[446]));
Q_AN02 U810 ( .A0(n41), .A1(gcm_dak_cmd_in[446]), .Z(n308));
Q_MX02 U811 ( .S(n39), .A0(gcm_dek_cmd_in[445]), .A1(n309), .Z(gcm_cmd_in[445]));
Q_AN02 U812 ( .A0(n41), .A1(gcm_dak_cmd_in[445]), .Z(n309));
Q_MX02 U813 ( .S(n39), .A0(gcm_dek_cmd_in[444]), .A1(n310), .Z(gcm_cmd_in[444]));
Q_AN02 U814 ( .A0(n41), .A1(gcm_dak_cmd_in[444]), .Z(n310));
Q_MX02 U815 ( .S(n39), .A0(gcm_dek_cmd_in[443]), .A1(n311), .Z(gcm_cmd_in[443]));
Q_AN02 U816 ( .A0(n41), .A1(gcm_dak_cmd_in[443]), .Z(n311));
Q_MX02 U817 ( .S(n39), .A0(gcm_dek_cmd_in[442]), .A1(n312), .Z(gcm_cmd_in[442]));
Q_AN02 U818 ( .A0(n41), .A1(gcm_dak_cmd_in[442]), .Z(n312));
Q_MX02 U819 ( .S(n39), .A0(gcm_dek_cmd_in[441]), .A1(n313), .Z(gcm_cmd_in[441]));
Q_AN02 U820 ( .A0(n41), .A1(gcm_dak_cmd_in[441]), .Z(n313));
Q_MX02 U821 ( .S(n39), .A0(gcm_dek_cmd_in[440]), .A1(n314), .Z(gcm_cmd_in[440]));
Q_AN02 U822 ( .A0(n41), .A1(gcm_dak_cmd_in[440]), .Z(n314));
Q_MX02 U823 ( .S(n39), .A0(gcm_dek_cmd_in[439]), .A1(n315), .Z(gcm_cmd_in[439]));
Q_AN02 U824 ( .A0(n41), .A1(gcm_dak_cmd_in[439]), .Z(n315));
Q_MX02 U825 ( .S(n39), .A0(gcm_dek_cmd_in[438]), .A1(n316), .Z(gcm_cmd_in[438]));
Q_AN02 U826 ( .A0(n41), .A1(gcm_dak_cmd_in[438]), .Z(n316));
Q_MX02 U827 ( .S(n39), .A0(gcm_dek_cmd_in[437]), .A1(n317), .Z(gcm_cmd_in[437]));
Q_AN02 U828 ( .A0(n41), .A1(gcm_dak_cmd_in[437]), .Z(n317));
Q_MX02 U829 ( .S(n39), .A0(gcm_dek_cmd_in[436]), .A1(n318), .Z(gcm_cmd_in[436]));
Q_AN02 U830 ( .A0(n41), .A1(gcm_dak_cmd_in[436]), .Z(n318));
Q_MX02 U831 ( .S(n39), .A0(gcm_dek_cmd_in[435]), .A1(n319), .Z(gcm_cmd_in[435]));
Q_AN02 U832 ( .A0(n41), .A1(gcm_dak_cmd_in[435]), .Z(n319));
Q_MX02 U833 ( .S(n39), .A0(gcm_dek_cmd_in[434]), .A1(n320), .Z(gcm_cmd_in[434]));
Q_AN02 U834 ( .A0(n41), .A1(gcm_dak_cmd_in[434]), .Z(n320));
Q_MX02 U835 ( .S(n39), .A0(gcm_dek_cmd_in[433]), .A1(n321), .Z(gcm_cmd_in[433]));
Q_AN02 U836 ( .A0(n41), .A1(gcm_dak_cmd_in[433]), .Z(n321));
Q_MX02 U837 ( .S(n39), .A0(gcm_dek_cmd_in[432]), .A1(n322), .Z(gcm_cmd_in[432]));
Q_AN02 U838 ( .A0(n41), .A1(gcm_dak_cmd_in[432]), .Z(n322));
Q_MX02 U839 ( .S(n39), .A0(gcm_dek_cmd_in[431]), .A1(n323), .Z(gcm_cmd_in[431]));
Q_AN02 U840 ( .A0(n41), .A1(gcm_dak_cmd_in[431]), .Z(n323));
Q_MX02 U841 ( .S(n39), .A0(gcm_dek_cmd_in[430]), .A1(n324), .Z(gcm_cmd_in[430]));
Q_AN02 U842 ( .A0(n41), .A1(gcm_dak_cmd_in[430]), .Z(n324));
Q_MX02 U843 ( .S(n39), .A0(gcm_dek_cmd_in[429]), .A1(n325), .Z(gcm_cmd_in[429]));
Q_AN02 U844 ( .A0(n41), .A1(gcm_dak_cmd_in[429]), .Z(n325));
Q_MX02 U845 ( .S(n39), .A0(gcm_dek_cmd_in[428]), .A1(n326), .Z(gcm_cmd_in[428]));
Q_AN02 U846 ( .A0(n41), .A1(gcm_dak_cmd_in[428]), .Z(n326));
Q_MX02 U847 ( .S(n39), .A0(gcm_dek_cmd_in[427]), .A1(n327), .Z(gcm_cmd_in[427]));
Q_AN02 U848 ( .A0(n41), .A1(gcm_dak_cmd_in[427]), .Z(n327));
Q_MX02 U849 ( .S(n39), .A0(gcm_dek_cmd_in[426]), .A1(n328), .Z(gcm_cmd_in[426]));
Q_AN02 U850 ( .A0(n41), .A1(gcm_dak_cmd_in[426]), .Z(n328));
Q_MX02 U851 ( .S(n39), .A0(gcm_dek_cmd_in[425]), .A1(n329), .Z(gcm_cmd_in[425]));
Q_AN02 U852 ( .A0(n41), .A1(gcm_dak_cmd_in[425]), .Z(n329));
Q_MX02 U853 ( .S(n39), .A0(gcm_dek_cmd_in[424]), .A1(n330), .Z(gcm_cmd_in[424]));
Q_AN02 U854 ( .A0(n41), .A1(gcm_dak_cmd_in[424]), .Z(n330));
Q_MX02 U855 ( .S(n39), .A0(gcm_dek_cmd_in[423]), .A1(n331), .Z(gcm_cmd_in[423]));
Q_AN02 U856 ( .A0(n41), .A1(gcm_dak_cmd_in[423]), .Z(n331));
Q_MX02 U857 ( .S(n39), .A0(gcm_dek_cmd_in[422]), .A1(n332), .Z(gcm_cmd_in[422]));
Q_AN02 U858 ( .A0(n41), .A1(gcm_dak_cmd_in[422]), .Z(n332));
Q_MX02 U859 ( .S(n39), .A0(gcm_dek_cmd_in[421]), .A1(n333), .Z(gcm_cmd_in[421]));
Q_AN02 U860 ( .A0(n41), .A1(gcm_dak_cmd_in[421]), .Z(n333));
Q_MX02 U861 ( .S(n39), .A0(gcm_dek_cmd_in[420]), .A1(n334), .Z(gcm_cmd_in[420]));
Q_AN02 U862 ( .A0(n41), .A1(gcm_dak_cmd_in[420]), .Z(n334));
Q_MX02 U863 ( .S(n39), .A0(gcm_dek_cmd_in[419]), .A1(n335), .Z(gcm_cmd_in[419]));
Q_AN02 U864 ( .A0(n41), .A1(gcm_dak_cmd_in[419]), .Z(n335));
Q_MX02 U865 ( .S(n39), .A0(gcm_dek_cmd_in[418]), .A1(n336), .Z(gcm_cmd_in[418]));
Q_AN02 U866 ( .A0(n41), .A1(gcm_dak_cmd_in[418]), .Z(n336));
Q_MX02 U867 ( .S(n39), .A0(gcm_dek_cmd_in[417]), .A1(n337), .Z(gcm_cmd_in[417]));
Q_AN02 U868 ( .A0(n41), .A1(gcm_dak_cmd_in[417]), .Z(n337));
Q_MX02 U869 ( .S(n39), .A0(gcm_dek_cmd_in[416]), .A1(n338), .Z(gcm_cmd_in[416]));
Q_AN02 U870 ( .A0(n41), .A1(gcm_dak_cmd_in[416]), .Z(n338));
Q_MX02 U871 ( .S(n39), .A0(gcm_dek_cmd_in[415]), .A1(n339), .Z(gcm_cmd_in[415]));
Q_AN02 U872 ( .A0(n41), .A1(gcm_dak_cmd_in[415]), .Z(n339));
Q_MX02 U873 ( .S(n39), .A0(gcm_dek_cmd_in[414]), .A1(n340), .Z(gcm_cmd_in[414]));
Q_AN02 U874 ( .A0(n41), .A1(gcm_dak_cmd_in[414]), .Z(n340));
Q_MX02 U875 ( .S(n39), .A0(gcm_dek_cmd_in[413]), .A1(n341), .Z(gcm_cmd_in[413]));
Q_AN02 U876 ( .A0(n41), .A1(gcm_dak_cmd_in[413]), .Z(n341));
Q_MX02 U877 ( .S(n39), .A0(gcm_dek_cmd_in[412]), .A1(n342), .Z(gcm_cmd_in[412]));
Q_AN02 U878 ( .A0(n41), .A1(gcm_dak_cmd_in[412]), .Z(n342));
Q_MX02 U879 ( .S(n39), .A0(gcm_dek_cmd_in[411]), .A1(n343), .Z(gcm_cmd_in[411]));
Q_AN02 U880 ( .A0(n41), .A1(gcm_dak_cmd_in[411]), .Z(n343));
Q_MX02 U881 ( .S(n39), .A0(gcm_dek_cmd_in[410]), .A1(n344), .Z(gcm_cmd_in[410]));
Q_AN02 U882 ( .A0(n41), .A1(gcm_dak_cmd_in[410]), .Z(n344));
Q_MX02 U883 ( .S(n39), .A0(gcm_dek_cmd_in[409]), .A1(n345), .Z(gcm_cmd_in[409]));
Q_AN02 U884 ( .A0(n41), .A1(gcm_dak_cmd_in[409]), .Z(n345));
Q_MX02 U885 ( .S(n39), .A0(gcm_dek_cmd_in[408]), .A1(n346), .Z(gcm_cmd_in[408]));
Q_AN02 U886 ( .A0(n41), .A1(gcm_dak_cmd_in[408]), .Z(n346));
Q_MX02 U887 ( .S(n39), .A0(gcm_dek_cmd_in[407]), .A1(n347), .Z(gcm_cmd_in[407]));
Q_AN02 U888 ( .A0(n41), .A1(gcm_dak_cmd_in[407]), .Z(n347));
Q_MX02 U889 ( .S(n39), .A0(gcm_dek_cmd_in[406]), .A1(n348), .Z(gcm_cmd_in[406]));
Q_AN02 U890 ( .A0(n41), .A1(gcm_dak_cmd_in[406]), .Z(n348));
Q_MX02 U891 ( .S(n39), .A0(gcm_dek_cmd_in[405]), .A1(n349), .Z(gcm_cmd_in[405]));
Q_AN02 U892 ( .A0(n41), .A1(gcm_dak_cmd_in[405]), .Z(n349));
Q_MX02 U893 ( .S(n39), .A0(gcm_dek_cmd_in[404]), .A1(n350), .Z(gcm_cmd_in[404]));
Q_AN02 U894 ( .A0(n41), .A1(gcm_dak_cmd_in[404]), .Z(n350));
Q_MX02 U895 ( .S(n39), .A0(gcm_dek_cmd_in[403]), .A1(n351), .Z(gcm_cmd_in[403]));
Q_AN02 U896 ( .A0(n41), .A1(gcm_dak_cmd_in[403]), .Z(n351));
Q_MX02 U897 ( .S(n39), .A0(gcm_dek_cmd_in[402]), .A1(n352), .Z(gcm_cmd_in[402]));
Q_AN02 U898 ( .A0(n41), .A1(gcm_dak_cmd_in[402]), .Z(n352));
Q_MX02 U899 ( .S(n39), .A0(gcm_dek_cmd_in[401]), .A1(n353), .Z(gcm_cmd_in[401]));
Q_AN02 U900 ( .A0(n41), .A1(gcm_dak_cmd_in[401]), .Z(n353));
Q_MX02 U901 ( .S(n39), .A0(gcm_dek_cmd_in[400]), .A1(n354), .Z(gcm_cmd_in[400]));
Q_AN02 U902 ( .A0(n41), .A1(gcm_dak_cmd_in[400]), .Z(n354));
Q_MX02 U903 ( .S(n39), .A0(gcm_dek_cmd_in[399]), .A1(n355), .Z(gcm_cmd_in[399]));
Q_AN02 U904 ( .A0(n41), .A1(gcm_dak_cmd_in[399]), .Z(n355));
Q_MX02 U905 ( .S(n39), .A0(gcm_dek_cmd_in[398]), .A1(n356), .Z(gcm_cmd_in[398]));
Q_AN02 U906 ( .A0(n41), .A1(gcm_dak_cmd_in[398]), .Z(n356));
Q_MX02 U907 ( .S(n39), .A0(gcm_dek_cmd_in[397]), .A1(n357), .Z(gcm_cmd_in[397]));
Q_AN02 U908 ( .A0(n41), .A1(gcm_dak_cmd_in[397]), .Z(n357));
Q_MX02 U909 ( .S(n39), .A0(gcm_dek_cmd_in[396]), .A1(n358), .Z(gcm_cmd_in[396]));
Q_AN02 U910 ( .A0(n41), .A1(gcm_dak_cmd_in[396]), .Z(n358));
Q_MX02 U911 ( .S(n39), .A0(gcm_dek_cmd_in[395]), .A1(n359), .Z(gcm_cmd_in[395]));
Q_AN02 U912 ( .A0(n41), .A1(gcm_dak_cmd_in[395]), .Z(n359));
Q_MX02 U913 ( .S(n39), .A0(gcm_dek_cmd_in[394]), .A1(n360), .Z(gcm_cmd_in[394]));
Q_AN02 U914 ( .A0(n41), .A1(gcm_dak_cmd_in[394]), .Z(n360));
Q_MX02 U915 ( .S(n39), .A0(gcm_dek_cmd_in[393]), .A1(n361), .Z(gcm_cmd_in[393]));
Q_AN02 U916 ( .A0(n41), .A1(gcm_dak_cmd_in[393]), .Z(n361));
Q_MX02 U917 ( .S(n39), .A0(gcm_dek_cmd_in[392]), .A1(n362), .Z(gcm_cmd_in[392]));
Q_AN02 U918 ( .A0(n41), .A1(gcm_dak_cmd_in[392]), .Z(n362));
Q_MX02 U919 ( .S(n39), .A0(gcm_dek_cmd_in[391]), .A1(n363), .Z(gcm_cmd_in[391]));
Q_AN02 U920 ( .A0(n41), .A1(gcm_dak_cmd_in[391]), .Z(n363));
Q_MX02 U921 ( .S(n39), .A0(gcm_dek_cmd_in[390]), .A1(n364), .Z(gcm_cmd_in[390]));
Q_AN02 U922 ( .A0(n41), .A1(gcm_dak_cmd_in[390]), .Z(n364));
Q_MX02 U923 ( .S(n39), .A0(gcm_dek_cmd_in[389]), .A1(n365), .Z(gcm_cmd_in[389]));
Q_AN02 U924 ( .A0(n41), .A1(gcm_dak_cmd_in[389]), .Z(n365));
Q_MX02 U925 ( .S(n39), .A0(gcm_dek_cmd_in[388]), .A1(n366), .Z(gcm_cmd_in[388]));
Q_AN02 U926 ( .A0(n41), .A1(gcm_dak_cmd_in[388]), .Z(n366));
Q_MX02 U927 ( .S(n39), .A0(gcm_dek_cmd_in[387]), .A1(n367), .Z(gcm_cmd_in[387]));
Q_AN02 U928 ( .A0(n41), .A1(gcm_dak_cmd_in[387]), .Z(n367));
Q_MX02 U929 ( .S(n39), .A0(gcm_dek_cmd_in[386]), .A1(n368), .Z(gcm_cmd_in[386]));
Q_AN02 U930 ( .A0(n41), .A1(gcm_dak_cmd_in[386]), .Z(n368));
Q_MX02 U931 ( .S(n39), .A0(gcm_dek_cmd_in[385]), .A1(n369), .Z(gcm_cmd_in[385]));
Q_AN02 U932 ( .A0(n41), .A1(gcm_dak_cmd_in[385]), .Z(n369));
Q_MX02 U933 ( .S(n39), .A0(gcm_dek_cmd_in[384]), .A1(n370), .Z(gcm_cmd_in[384]));
Q_AN02 U934 ( .A0(n41), .A1(gcm_dak_cmd_in[384]), .Z(n370));
Q_MX02 U935 ( .S(n39), .A0(gcm_dek_cmd_in[383]), .A1(n371), .Z(gcm_cmd_in[383]));
Q_AN02 U936 ( .A0(n41), .A1(gcm_dak_cmd_in[383]), .Z(n371));
Q_MX02 U937 ( .S(n39), .A0(gcm_dek_cmd_in[382]), .A1(n372), .Z(gcm_cmd_in[382]));
Q_AN02 U938 ( .A0(n41), .A1(gcm_dak_cmd_in[382]), .Z(n372));
Q_MX02 U939 ( .S(n39), .A0(gcm_dek_cmd_in[381]), .A1(n373), .Z(gcm_cmd_in[381]));
Q_AN02 U940 ( .A0(n41), .A1(gcm_dak_cmd_in[381]), .Z(n373));
Q_MX02 U941 ( .S(n39), .A0(gcm_dek_cmd_in[380]), .A1(n374), .Z(gcm_cmd_in[380]));
Q_AN02 U942 ( .A0(n41), .A1(gcm_dak_cmd_in[380]), .Z(n374));
Q_MX02 U943 ( .S(n39), .A0(gcm_dek_cmd_in[379]), .A1(n375), .Z(gcm_cmd_in[379]));
Q_AN02 U944 ( .A0(n41), .A1(gcm_dak_cmd_in[379]), .Z(n375));
Q_MX02 U945 ( .S(n39), .A0(gcm_dek_cmd_in[378]), .A1(n376), .Z(gcm_cmd_in[378]));
Q_AN02 U946 ( .A0(n41), .A1(gcm_dak_cmd_in[378]), .Z(n376));
Q_MX02 U947 ( .S(n39), .A0(gcm_dek_cmd_in[377]), .A1(n377), .Z(gcm_cmd_in[377]));
Q_AN02 U948 ( .A0(n41), .A1(gcm_dak_cmd_in[377]), .Z(n377));
Q_MX02 U949 ( .S(n39), .A0(gcm_dek_cmd_in[376]), .A1(n378), .Z(gcm_cmd_in[376]));
Q_AN02 U950 ( .A0(n41), .A1(gcm_dak_cmd_in[376]), .Z(n378));
Q_MX02 U951 ( .S(n39), .A0(gcm_dek_cmd_in[375]), .A1(n379), .Z(gcm_cmd_in[375]));
Q_AN02 U952 ( .A0(n41), .A1(gcm_dak_cmd_in[375]), .Z(n379));
Q_MX02 U953 ( .S(n39), .A0(gcm_dek_cmd_in[374]), .A1(n380), .Z(gcm_cmd_in[374]));
Q_AN02 U954 ( .A0(n41), .A1(gcm_dak_cmd_in[374]), .Z(n380));
Q_MX02 U955 ( .S(n39), .A0(gcm_dek_cmd_in[373]), .A1(n381), .Z(gcm_cmd_in[373]));
Q_AN02 U956 ( .A0(n41), .A1(gcm_dak_cmd_in[373]), .Z(n381));
Q_MX02 U957 ( .S(n39), .A0(gcm_dek_cmd_in[372]), .A1(n382), .Z(gcm_cmd_in[372]));
Q_AN02 U958 ( .A0(n41), .A1(gcm_dak_cmd_in[372]), .Z(n382));
Q_MX02 U959 ( .S(n39), .A0(gcm_dek_cmd_in[371]), .A1(n383), .Z(gcm_cmd_in[371]));
Q_AN02 U960 ( .A0(n41), .A1(gcm_dak_cmd_in[371]), .Z(n383));
Q_MX02 U961 ( .S(n39), .A0(gcm_dek_cmd_in[370]), .A1(n384), .Z(gcm_cmd_in[370]));
Q_AN02 U962 ( .A0(n41), .A1(gcm_dak_cmd_in[370]), .Z(n384));
Q_MX02 U963 ( .S(n39), .A0(gcm_dek_cmd_in[369]), .A1(n385), .Z(gcm_cmd_in[369]));
Q_AN02 U964 ( .A0(n41), .A1(gcm_dak_cmd_in[369]), .Z(n385));
Q_MX02 U965 ( .S(n39), .A0(gcm_dek_cmd_in[368]), .A1(n386), .Z(gcm_cmd_in[368]));
Q_AN02 U966 ( .A0(n41), .A1(gcm_dak_cmd_in[368]), .Z(n386));
Q_MX02 U967 ( .S(n39), .A0(gcm_dek_cmd_in[367]), .A1(n387), .Z(gcm_cmd_in[367]));
Q_AN02 U968 ( .A0(n41), .A1(gcm_dak_cmd_in[367]), .Z(n387));
Q_MX02 U969 ( .S(n39), .A0(gcm_dek_cmd_in[366]), .A1(n388), .Z(gcm_cmd_in[366]));
Q_AN02 U970 ( .A0(n41), .A1(gcm_dak_cmd_in[366]), .Z(n388));
Q_MX02 U971 ( .S(n39), .A0(gcm_dek_cmd_in[365]), .A1(n389), .Z(gcm_cmd_in[365]));
Q_AN02 U972 ( .A0(n41), .A1(gcm_dak_cmd_in[365]), .Z(n389));
Q_MX02 U973 ( .S(n39), .A0(gcm_dek_cmd_in[364]), .A1(n390), .Z(gcm_cmd_in[364]));
Q_AN02 U974 ( .A0(n41), .A1(gcm_dak_cmd_in[364]), .Z(n390));
Q_MX02 U975 ( .S(n39), .A0(gcm_dek_cmd_in[363]), .A1(n391), .Z(gcm_cmd_in[363]));
Q_AN02 U976 ( .A0(n41), .A1(gcm_dak_cmd_in[363]), .Z(n391));
Q_MX02 U977 ( .S(n39), .A0(gcm_dek_cmd_in[362]), .A1(n392), .Z(gcm_cmd_in[362]));
Q_AN02 U978 ( .A0(n41), .A1(gcm_dak_cmd_in[362]), .Z(n392));
Q_MX02 U979 ( .S(n39), .A0(gcm_dek_cmd_in[361]), .A1(n393), .Z(gcm_cmd_in[361]));
Q_AN02 U980 ( .A0(n41), .A1(gcm_dak_cmd_in[361]), .Z(n393));
Q_MX02 U981 ( .S(n39), .A0(gcm_dek_cmd_in[360]), .A1(n394), .Z(gcm_cmd_in[360]));
Q_AN02 U982 ( .A0(n41), .A1(gcm_dak_cmd_in[360]), .Z(n394));
Q_MX02 U983 ( .S(n39), .A0(gcm_dek_cmd_in[359]), .A1(n395), .Z(gcm_cmd_in[359]));
Q_AN02 U984 ( .A0(n41), .A1(gcm_dak_cmd_in[359]), .Z(n395));
Q_MX02 U985 ( .S(n39), .A0(gcm_dek_cmd_in[358]), .A1(n396), .Z(gcm_cmd_in[358]));
Q_AN02 U986 ( .A0(n41), .A1(gcm_dak_cmd_in[358]), .Z(n396));
Q_MX02 U987 ( .S(n39), .A0(gcm_dek_cmd_in[357]), .A1(n397), .Z(gcm_cmd_in[357]));
Q_AN02 U988 ( .A0(n41), .A1(gcm_dak_cmd_in[357]), .Z(n397));
Q_MX02 U989 ( .S(n39), .A0(gcm_dek_cmd_in[356]), .A1(n398), .Z(gcm_cmd_in[356]));
Q_AN02 U990 ( .A0(n41), .A1(gcm_dak_cmd_in[356]), .Z(n398));
Q_MX02 U991 ( .S(n39), .A0(gcm_dek_cmd_in[355]), .A1(n399), .Z(gcm_cmd_in[355]));
Q_AN02 U992 ( .A0(n41), .A1(gcm_dak_cmd_in[355]), .Z(n399));
Q_MX02 U993 ( .S(n39), .A0(gcm_dek_cmd_in[354]), .A1(n400), .Z(gcm_cmd_in[354]));
Q_AN02 U994 ( .A0(n41), .A1(gcm_dak_cmd_in[354]), .Z(n400));
Q_MX02 U995 ( .S(n39), .A0(gcm_dek_cmd_in[353]), .A1(n401), .Z(gcm_cmd_in[353]));
Q_AN02 U996 ( .A0(n41), .A1(gcm_dak_cmd_in[353]), .Z(n401));
Q_MX02 U997 ( .S(n39), .A0(gcm_dek_cmd_in[352]), .A1(n402), .Z(gcm_cmd_in[352]));
Q_AN02 U998 ( .A0(n41), .A1(gcm_dak_cmd_in[352]), .Z(n402));
Q_MX02 U999 ( .S(n39), .A0(gcm_dek_cmd_in[351]), .A1(n403), .Z(gcm_cmd_in[351]));
Q_AN02 U1000 ( .A0(n41), .A1(gcm_dak_cmd_in[351]), .Z(n403));
Q_MX02 U1001 ( .S(n39), .A0(gcm_dek_cmd_in[350]), .A1(n404), .Z(gcm_cmd_in[350]));
Q_AN02 U1002 ( .A0(n41), .A1(gcm_dak_cmd_in[350]), .Z(n404));
Q_MX02 U1003 ( .S(n39), .A0(gcm_dek_cmd_in[349]), .A1(n405), .Z(gcm_cmd_in[349]));
Q_AN02 U1004 ( .A0(n41), .A1(gcm_dak_cmd_in[349]), .Z(n405));
Q_MX02 U1005 ( .S(n39), .A0(gcm_dek_cmd_in[348]), .A1(n406), .Z(gcm_cmd_in[348]));
Q_AN02 U1006 ( .A0(n41), .A1(gcm_dak_cmd_in[348]), .Z(n406));
Q_MX02 U1007 ( .S(n39), .A0(gcm_dek_cmd_in[347]), .A1(n407), .Z(gcm_cmd_in[347]));
Q_AN02 U1008 ( .A0(n41), .A1(gcm_dak_cmd_in[347]), .Z(n407));
Q_MX02 U1009 ( .S(n39), .A0(gcm_dek_cmd_in[346]), .A1(n408), .Z(gcm_cmd_in[346]));
Q_AN02 U1010 ( .A0(n41), .A1(gcm_dak_cmd_in[346]), .Z(n408));
Q_MX02 U1011 ( .S(n39), .A0(gcm_dek_cmd_in[345]), .A1(n409), .Z(gcm_cmd_in[345]));
Q_AN02 U1012 ( .A0(n41), .A1(gcm_dak_cmd_in[345]), .Z(n409));
Q_MX02 U1013 ( .S(n39), .A0(gcm_dek_cmd_in[344]), .A1(n410), .Z(gcm_cmd_in[344]));
Q_AN02 U1014 ( .A0(n41), .A1(gcm_dak_cmd_in[344]), .Z(n410));
Q_MX02 U1015 ( .S(n39), .A0(gcm_dek_cmd_in[343]), .A1(n411), .Z(gcm_cmd_in[343]));
Q_AN02 U1016 ( .A0(n41), .A1(gcm_dak_cmd_in[343]), .Z(n411));
Q_MX02 U1017 ( .S(n39), .A0(gcm_dek_cmd_in[342]), .A1(n412), .Z(gcm_cmd_in[342]));
Q_AN02 U1018 ( .A0(n41), .A1(gcm_dak_cmd_in[342]), .Z(n412));
Q_MX02 U1019 ( .S(n39), .A0(gcm_dek_cmd_in[341]), .A1(n413), .Z(gcm_cmd_in[341]));
Q_AN02 U1020 ( .A0(n41), .A1(gcm_dak_cmd_in[341]), .Z(n413));
Q_MX02 U1021 ( .S(n39), .A0(gcm_dek_cmd_in[340]), .A1(n414), .Z(gcm_cmd_in[340]));
Q_AN02 U1022 ( .A0(n41), .A1(gcm_dak_cmd_in[340]), .Z(n414));
Q_MX02 U1023 ( .S(n39), .A0(gcm_dek_cmd_in[339]), .A1(n415), .Z(gcm_cmd_in[339]));
Q_AN02 U1024 ( .A0(n41), .A1(gcm_dak_cmd_in[339]), .Z(n415));
Q_MX02 U1025 ( .S(n39), .A0(gcm_dek_cmd_in[338]), .A1(n416), .Z(gcm_cmd_in[338]));
Q_AN02 U1026 ( .A0(n41), .A1(gcm_dak_cmd_in[338]), .Z(n416));
Q_MX02 U1027 ( .S(n39), .A0(gcm_dek_cmd_in[337]), .A1(n417), .Z(gcm_cmd_in[337]));
Q_AN02 U1028 ( .A0(n41), .A1(gcm_dak_cmd_in[337]), .Z(n417));
Q_MX02 U1029 ( .S(n39), .A0(gcm_dek_cmd_in[336]), .A1(n418), .Z(gcm_cmd_in[336]));
Q_AN02 U1030 ( .A0(n41), .A1(gcm_dak_cmd_in[336]), .Z(n418));
Q_MX02 U1031 ( .S(n39), .A0(gcm_dek_cmd_in[335]), .A1(n419), .Z(gcm_cmd_in[335]));
Q_AN02 U1032 ( .A0(n41), .A1(gcm_dak_cmd_in[335]), .Z(n419));
Q_MX02 U1033 ( .S(n39), .A0(gcm_dek_cmd_in[334]), .A1(n420), .Z(gcm_cmd_in[334]));
Q_AN02 U1034 ( .A0(n41), .A1(gcm_dak_cmd_in[334]), .Z(n420));
Q_MX02 U1035 ( .S(n39), .A0(gcm_dek_cmd_in[333]), .A1(n421), .Z(gcm_cmd_in[333]));
Q_AN02 U1036 ( .A0(n41), .A1(gcm_dak_cmd_in[333]), .Z(n421));
Q_MX02 U1037 ( .S(n39), .A0(gcm_dek_cmd_in[332]), .A1(n422), .Z(gcm_cmd_in[332]));
Q_AN02 U1038 ( .A0(n41), .A1(gcm_dak_cmd_in[332]), .Z(n422));
Q_MX02 U1039 ( .S(n39), .A0(gcm_dek_cmd_in[331]), .A1(n423), .Z(gcm_cmd_in[331]));
Q_AN02 U1040 ( .A0(n41), .A1(gcm_dak_cmd_in[331]), .Z(n423));
Q_MX02 U1041 ( .S(n39), .A0(gcm_dek_cmd_in[330]), .A1(n424), .Z(gcm_cmd_in[330]));
Q_AN02 U1042 ( .A0(n41), .A1(gcm_dak_cmd_in[330]), .Z(n424));
Q_MX02 U1043 ( .S(n39), .A0(gcm_dek_cmd_in[329]), .A1(n425), .Z(gcm_cmd_in[329]));
Q_AN02 U1044 ( .A0(n41), .A1(gcm_dak_cmd_in[329]), .Z(n425));
Q_MX02 U1045 ( .S(n39), .A0(gcm_dek_cmd_in[328]), .A1(n426), .Z(gcm_cmd_in[328]));
Q_AN02 U1046 ( .A0(n41), .A1(gcm_dak_cmd_in[328]), .Z(n426));
Q_MX02 U1047 ( .S(n39), .A0(gcm_dek_cmd_in[327]), .A1(n427), .Z(gcm_cmd_in[327]));
Q_AN02 U1048 ( .A0(n41), .A1(gcm_dak_cmd_in[327]), .Z(n427));
Q_MX02 U1049 ( .S(n39), .A0(gcm_dek_cmd_in[326]), .A1(n428), .Z(gcm_cmd_in[326]));
Q_AN02 U1050 ( .A0(n41), .A1(gcm_dak_cmd_in[326]), .Z(n428));
Q_MX02 U1051 ( .S(n39), .A0(gcm_dek_cmd_in[325]), .A1(n429), .Z(gcm_cmd_in[325]));
Q_AN02 U1052 ( .A0(n41), .A1(gcm_dak_cmd_in[325]), .Z(n429));
Q_MX02 U1053 ( .S(n39), .A0(gcm_dek_cmd_in[324]), .A1(n430), .Z(gcm_cmd_in[324]));
Q_AN02 U1054 ( .A0(n41), .A1(gcm_dak_cmd_in[324]), .Z(n430));
Q_MX02 U1055 ( .S(n39), .A0(gcm_dek_cmd_in[323]), .A1(n431), .Z(gcm_cmd_in[323]));
Q_AN02 U1056 ( .A0(n41), .A1(gcm_dak_cmd_in[323]), .Z(n431));
Q_MX02 U1057 ( .S(n39), .A0(gcm_dek_cmd_in[322]), .A1(n432), .Z(gcm_cmd_in[322]));
Q_AN02 U1058 ( .A0(n41), .A1(gcm_dak_cmd_in[322]), .Z(n432));
Q_MX02 U1059 ( .S(n39), .A0(gcm_dek_cmd_in[321]), .A1(n433), .Z(gcm_cmd_in[321]));
Q_AN02 U1060 ( .A0(n41), .A1(gcm_dak_cmd_in[321]), .Z(n433));
Q_MX02 U1061 ( .S(n39), .A0(gcm_dek_cmd_in[320]), .A1(n434), .Z(gcm_cmd_in[320]));
Q_AN02 U1062 ( .A0(n41), .A1(gcm_dak_cmd_in[320]), .Z(n434));
Q_MX02 U1063 ( .S(n39), .A0(gcm_dek_cmd_in[319]), .A1(n435), .Z(gcm_cmd_in[319]));
Q_AN02 U1064 ( .A0(n41), .A1(gcm_dak_cmd_in[319]), .Z(n435));
Q_MX02 U1065 ( .S(n39), .A0(gcm_dek_cmd_in[318]), .A1(n436), .Z(gcm_cmd_in[318]));
Q_AN02 U1066 ( .A0(n41), .A1(gcm_dak_cmd_in[318]), .Z(n436));
Q_MX02 U1067 ( .S(n39), .A0(gcm_dek_cmd_in[317]), .A1(n437), .Z(gcm_cmd_in[317]));
Q_AN02 U1068 ( .A0(n41), .A1(gcm_dak_cmd_in[317]), .Z(n437));
Q_MX02 U1069 ( .S(n39), .A0(gcm_dek_cmd_in[316]), .A1(n438), .Z(gcm_cmd_in[316]));
Q_AN02 U1070 ( .A0(n41), .A1(gcm_dak_cmd_in[316]), .Z(n438));
Q_MX02 U1071 ( .S(n39), .A0(gcm_dek_cmd_in[315]), .A1(n439), .Z(gcm_cmd_in[315]));
Q_AN02 U1072 ( .A0(n41), .A1(gcm_dak_cmd_in[315]), .Z(n439));
Q_MX02 U1073 ( .S(n39), .A0(gcm_dek_cmd_in[314]), .A1(n440), .Z(gcm_cmd_in[314]));
Q_AN02 U1074 ( .A0(n41), .A1(gcm_dak_cmd_in[314]), .Z(n440));
Q_MX02 U1075 ( .S(n39), .A0(gcm_dek_cmd_in[313]), .A1(n441), .Z(gcm_cmd_in[313]));
Q_AN02 U1076 ( .A0(n41), .A1(gcm_dak_cmd_in[313]), .Z(n441));
Q_MX02 U1077 ( .S(n39), .A0(gcm_dek_cmd_in[312]), .A1(n442), .Z(gcm_cmd_in[312]));
Q_AN02 U1078 ( .A0(n41), .A1(gcm_dak_cmd_in[312]), .Z(n442));
Q_MX02 U1079 ( .S(n39), .A0(gcm_dek_cmd_in[311]), .A1(n443), .Z(gcm_cmd_in[311]));
Q_AN02 U1080 ( .A0(n41), .A1(gcm_dak_cmd_in[311]), .Z(n443));
Q_MX02 U1081 ( .S(n39), .A0(gcm_dek_cmd_in[310]), .A1(n444), .Z(gcm_cmd_in[310]));
Q_AN02 U1082 ( .A0(n41), .A1(gcm_dak_cmd_in[310]), .Z(n444));
Q_MX02 U1083 ( .S(n39), .A0(gcm_dek_cmd_in[309]), .A1(n445), .Z(gcm_cmd_in[309]));
Q_AN02 U1084 ( .A0(n41), .A1(gcm_dak_cmd_in[309]), .Z(n445));
Q_MX02 U1085 ( .S(n39), .A0(gcm_dek_cmd_in[308]), .A1(n446), .Z(gcm_cmd_in[308]));
Q_AN02 U1086 ( .A0(n41), .A1(gcm_dak_cmd_in[308]), .Z(n446));
Q_MX02 U1087 ( .S(n39), .A0(gcm_dek_cmd_in[307]), .A1(n447), .Z(gcm_cmd_in[307]));
Q_AN02 U1088 ( .A0(n41), .A1(gcm_dak_cmd_in[307]), .Z(n447));
Q_MX02 U1089 ( .S(n39), .A0(gcm_dek_cmd_in[306]), .A1(n448), .Z(gcm_cmd_in[306]));
Q_AN02 U1090 ( .A0(n41), .A1(gcm_dak_cmd_in[306]), .Z(n448));
Q_MX02 U1091 ( .S(n39), .A0(gcm_dek_cmd_in[305]), .A1(n449), .Z(gcm_cmd_in[305]));
Q_AN02 U1092 ( .A0(n41), .A1(gcm_dak_cmd_in[305]), .Z(n449));
Q_MX02 U1093 ( .S(n39), .A0(gcm_dek_cmd_in[304]), .A1(n450), .Z(gcm_cmd_in[304]));
Q_AN02 U1094 ( .A0(n41), .A1(gcm_dak_cmd_in[304]), .Z(n450));
Q_MX02 U1095 ( .S(n39), .A0(gcm_dek_cmd_in[303]), .A1(n451), .Z(gcm_cmd_in[303]));
Q_AN02 U1096 ( .A0(n41), .A1(gcm_dak_cmd_in[303]), .Z(n451));
Q_MX02 U1097 ( .S(n39), .A0(gcm_dek_cmd_in[302]), .A1(n452), .Z(gcm_cmd_in[302]));
Q_AN02 U1098 ( .A0(n41), .A1(gcm_dak_cmd_in[302]), .Z(n452));
Q_MX02 U1099 ( .S(n39), .A0(gcm_dek_cmd_in[301]), .A1(n453), .Z(gcm_cmd_in[301]));
Q_AN02 U1100 ( .A0(n41), .A1(gcm_dak_cmd_in[301]), .Z(n453));
Q_MX02 U1101 ( .S(n39), .A0(gcm_dek_cmd_in[300]), .A1(n454), .Z(gcm_cmd_in[300]));
Q_AN02 U1102 ( .A0(n41), .A1(gcm_dak_cmd_in[300]), .Z(n454));
Q_MX02 U1103 ( .S(n39), .A0(gcm_dek_cmd_in[299]), .A1(n455), .Z(gcm_cmd_in[299]));
Q_AN02 U1104 ( .A0(n41), .A1(gcm_dak_cmd_in[299]), .Z(n455));
Q_MX02 U1105 ( .S(n39), .A0(gcm_dek_cmd_in[298]), .A1(n456), .Z(gcm_cmd_in[298]));
Q_AN02 U1106 ( .A0(n41), .A1(gcm_dak_cmd_in[298]), .Z(n456));
Q_MX02 U1107 ( .S(n39), .A0(gcm_dek_cmd_in[297]), .A1(n457), .Z(gcm_cmd_in[297]));
Q_AN02 U1108 ( .A0(n41), .A1(gcm_dak_cmd_in[297]), .Z(n457));
Q_MX02 U1109 ( .S(n39), .A0(gcm_dek_cmd_in[296]), .A1(n458), .Z(gcm_cmd_in[296]));
Q_AN02 U1110 ( .A0(n41), .A1(gcm_dak_cmd_in[296]), .Z(n458));
Q_MX02 U1111 ( .S(n39), .A0(gcm_dek_cmd_in[295]), .A1(n459), .Z(gcm_cmd_in[295]));
Q_AN02 U1112 ( .A0(n41), .A1(gcm_dak_cmd_in[295]), .Z(n459));
Q_MX02 U1113 ( .S(n39), .A0(gcm_dek_cmd_in[294]), .A1(n460), .Z(gcm_cmd_in[294]));
Q_AN02 U1114 ( .A0(n41), .A1(gcm_dak_cmd_in[294]), .Z(n460));
Q_MX02 U1115 ( .S(n39), .A0(gcm_dek_cmd_in[293]), .A1(n461), .Z(gcm_cmd_in[293]));
Q_AN02 U1116 ( .A0(n41), .A1(gcm_dak_cmd_in[293]), .Z(n461));
Q_MX02 U1117 ( .S(n39), .A0(gcm_dek_cmd_in[292]), .A1(n462), .Z(gcm_cmd_in[292]));
Q_AN02 U1118 ( .A0(n41), .A1(gcm_dak_cmd_in[292]), .Z(n462));
Q_MX02 U1119 ( .S(n39), .A0(gcm_dek_cmd_in[291]), .A1(n463), .Z(gcm_cmd_in[291]));
Q_AN02 U1120 ( .A0(n41), .A1(gcm_dak_cmd_in[291]), .Z(n463));
Q_MX02 U1121 ( .S(n39), .A0(gcm_dek_cmd_in[290]), .A1(n464), .Z(gcm_cmd_in[290]));
Q_AN02 U1122 ( .A0(n41), .A1(gcm_dak_cmd_in[290]), .Z(n464));
Q_MX02 U1123 ( .S(n39), .A0(gcm_dek_cmd_in[289]), .A1(n465), .Z(gcm_cmd_in[289]));
Q_AN02 U1124 ( .A0(n41), .A1(gcm_dak_cmd_in[289]), .Z(n465));
Q_MX02 U1125 ( .S(n39), .A0(gcm_dek_cmd_in[288]), .A1(n466), .Z(gcm_cmd_in[288]));
Q_AN02 U1126 ( .A0(n41), .A1(gcm_dak_cmd_in[288]), .Z(n466));
Q_MX02 U1127 ( .S(n39), .A0(gcm_dek_cmd_in[287]), .A1(n467), .Z(gcm_cmd_in[287]));
Q_AN02 U1128 ( .A0(n41), .A1(gcm_dak_cmd_in[287]), .Z(n467));
Q_MX02 U1129 ( .S(n39), .A0(gcm_dek_cmd_in[286]), .A1(n468), .Z(gcm_cmd_in[286]));
Q_AN02 U1130 ( .A0(n41), .A1(gcm_dak_cmd_in[286]), .Z(n468));
Q_MX02 U1131 ( .S(n39), .A0(gcm_dek_cmd_in[285]), .A1(n469), .Z(gcm_cmd_in[285]));
Q_AN02 U1132 ( .A0(n41), .A1(gcm_dak_cmd_in[285]), .Z(n469));
Q_MX02 U1133 ( .S(n39), .A0(gcm_dek_cmd_in[284]), .A1(n470), .Z(gcm_cmd_in[284]));
Q_AN02 U1134 ( .A0(n41), .A1(gcm_dak_cmd_in[284]), .Z(n470));
Q_MX02 U1135 ( .S(n39), .A0(gcm_dek_cmd_in[283]), .A1(n471), .Z(gcm_cmd_in[283]));
Q_AN02 U1136 ( .A0(n41), .A1(gcm_dak_cmd_in[283]), .Z(n471));
Q_MX02 U1137 ( .S(n39), .A0(gcm_dek_cmd_in[282]), .A1(n472), .Z(gcm_cmd_in[282]));
Q_AN02 U1138 ( .A0(n41), .A1(gcm_dak_cmd_in[282]), .Z(n472));
Q_MX02 U1139 ( .S(n39), .A0(gcm_dek_cmd_in[281]), .A1(n473), .Z(gcm_cmd_in[281]));
Q_AN02 U1140 ( .A0(n41), .A1(gcm_dak_cmd_in[281]), .Z(n473));
Q_MX02 U1141 ( .S(n39), .A0(gcm_dek_cmd_in[280]), .A1(n474), .Z(gcm_cmd_in[280]));
Q_AN02 U1142 ( .A0(n41), .A1(gcm_dak_cmd_in[280]), .Z(n474));
Q_MX02 U1143 ( .S(n39), .A0(gcm_dek_cmd_in[279]), .A1(n475), .Z(gcm_cmd_in[279]));
Q_AN02 U1144 ( .A0(n41), .A1(gcm_dak_cmd_in[279]), .Z(n475));
Q_MX02 U1145 ( .S(n39), .A0(gcm_dek_cmd_in[278]), .A1(n476), .Z(gcm_cmd_in[278]));
Q_AN02 U1146 ( .A0(n41), .A1(gcm_dak_cmd_in[278]), .Z(n476));
Q_MX02 U1147 ( .S(n39), .A0(gcm_dek_cmd_in[277]), .A1(n477), .Z(gcm_cmd_in[277]));
Q_AN02 U1148 ( .A0(n41), .A1(gcm_dak_cmd_in[277]), .Z(n477));
Q_MX02 U1149 ( .S(n39), .A0(gcm_dek_cmd_in[276]), .A1(n478), .Z(gcm_cmd_in[276]));
Q_AN02 U1150 ( .A0(n41), .A1(gcm_dak_cmd_in[276]), .Z(n478));
Q_MX02 U1151 ( .S(n39), .A0(gcm_dek_cmd_in[275]), .A1(n479), .Z(gcm_cmd_in[275]));
Q_AN02 U1152 ( .A0(n41), .A1(gcm_dak_cmd_in[275]), .Z(n479));
Q_MX02 U1153 ( .S(n39), .A0(gcm_dek_cmd_in[274]), .A1(n480), .Z(gcm_cmd_in[274]));
Q_AN02 U1154 ( .A0(n41), .A1(gcm_dak_cmd_in[274]), .Z(n480));
Q_MX02 U1155 ( .S(n39), .A0(gcm_dek_cmd_in[273]), .A1(n481), .Z(gcm_cmd_in[273]));
Q_AN02 U1156 ( .A0(n41), .A1(gcm_dak_cmd_in[273]), .Z(n481));
Q_MX02 U1157 ( .S(n39), .A0(gcm_dek_cmd_in[272]), .A1(n482), .Z(gcm_cmd_in[272]));
Q_AN02 U1158 ( .A0(n41), .A1(gcm_dak_cmd_in[272]), .Z(n482));
Q_MX02 U1159 ( .S(n39), .A0(gcm_dek_cmd_in[271]), .A1(n483), .Z(gcm_cmd_in[271]));
Q_AN02 U1160 ( .A0(n41), .A1(gcm_dak_cmd_in[271]), .Z(n483));
Q_MX02 U1161 ( .S(n39), .A0(gcm_dek_cmd_in[270]), .A1(n484), .Z(gcm_cmd_in[270]));
Q_AN02 U1162 ( .A0(n41), .A1(gcm_dak_cmd_in[270]), .Z(n484));
Q_MX02 U1163 ( .S(n39), .A0(gcm_dek_cmd_in[269]), .A1(n485), .Z(gcm_cmd_in[269]));
Q_AN02 U1164 ( .A0(n41), .A1(gcm_dak_cmd_in[269]), .Z(n485));
Q_MX02 U1165 ( .S(n39), .A0(gcm_dek_cmd_in[268]), .A1(n486), .Z(gcm_cmd_in[268]));
Q_AN02 U1166 ( .A0(n41), .A1(gcm_dak_cmd_in[268]), .Z(n486));
Q_MX02 U1167 ( .S(n39), .A0(gcm_dek_cmd_in[267]), .A1(n487), .Z(gcm_cmd_in[267]));
Q_AN02 U1168 ( .A0(n41), .A1(gcm_dak_cmd_in[267]), .Z(n487));
Q_MX02 U1169 ( .S(n39), .A0(gcm_dek_cmd_in[266]), .A1(n488), .Z(gcm_cmd_in[266]));
Q_AN02 U1170 ( .A0(n41), .A1(gcm_dak_cmd_in[266]), .Z(n488));
Q_MX02 U1171 ( .S(n39), .A0(gcm_dek_cmd_in[265]), .A1(n489), .Z(gcm_cmd_in[265]));
Q_AN02 U1172 ( .A0(n41), .A1(gcm_dak_cmd_in[265]), .Z(n489));
Q_MX02 U1173 ( .S(n39), .A0(gcm_dek_cmd_in[264]), .A1(n490), .Z(gcm_cmd_in[264]));
Q_AN02 U1174 ( .A0(n41), .A1(gcm_dak_cmd_in[264]), .Z(n490));
Q_MX02 U1175 ( .S(n39), .A0(gcm_dek_cmd_in[263]), .A1(n491), .Z(gcm_cmd_in[263]));
Q_AN02 U1176 ( .A0(n41), .A1(gcm_dak_cmd_in[263]), .Z(n491));
Q_MX02 U1177 ( .S(n39), .A0(gcm_dek_cmd_in[262]), .A1(n492), .Z(gcm_cmd_in[262]));
Q_AN02 U1178 ( .A0(n41), .A1(gcm_dak_cmd_in[262]), .Z(n492));
Q_MX02 U1179 ( .S(n39), .A0(gcm_dek_cmd_in[261]), .A1(n493), .Z(gcm_cmd_in[261]));
Q_AN02 U1180 ( .A0(n41), .A1(gcm_dak_cmd_in[261]), .Z(n493));
Q_MX02 U1181 ( .S(n39), .A0(gcm_dek_cmd_in[260]), .A1(n494), .Z(gcm_cmd_in[260]));
Q_AN02 U1182 ( .A0(n41), .A1(gcm_dak_cmd_in[260]), .Z(n494));
Q_MX02 U1183 ( .S(n39), .A0(gcm_dek_cmd_in[259]), .A1(n495), .Z(gcm_cmd_in[259]));
Q_AN02 U1184 ( .A0(n41), .A1(gcm_dak_cmd_in[259]), .Z(n495));
Q_MX02 U1185 ( .S(n39), .A0(gcm_dek_cmd_in[258]), .A1(n496), .Z(gcm_cmd_in[258]));
Q_AN02 U1186 ( .A0(n41), .A1(gcm_dak_cmd_in[258]), .Z(n496));
Q_MX02 U1187 ( .S(n39), .A0(gcm_dek_cmd_in[257]), .A1(n497), .Z(gcm_cmd_in[257]));
Q_AN02 U1188 ( .A0(n41), .A1(gcm_dak_cmd_in[257]), .Z(n497));
Q_MX02 U1189 ( .S(n39), .A0(gcm_dek_cmd_in[256]), .A1(n498), .Z(gcm_cmd_in[256]));
Q_AN02 U1190 ( .A0(n41), .A1(gcm_dak_cmd_in[256]), .Z(n498));
Q_MX02 U1191 ( .S(n39), .A0(gcm_dek_cmd_in[255]), .A1(n499), .Z(gcm_cmd_in[255]));
Q_AN02 U1192 ( .A0(n41), .A1(gcm_dak_cmd_in[255]), .Z(n499));
Q_MX02 U1193 ( .S(n39), .A0(gcm_dek_cmd_in[254]), .A1(n500), .Z(gcm_cmd_in[254]));
Q_AN02 U1194 ( .A0(n41), .A1(gcm_dak_cmd_in[254]), .Z(n500));
Q_MX02 U1195 ( .S(n39), .A0(gcm_dek_cmd_in[253]), .A1(n501), .Z(gcm_cmd_in[253]));
Q_AN02 U1196 ( .A0(n41), .A1(gcm_dak_cmd_in[253]), .Z(n501));
Q_MX02 U1197 ( .S(n39), .A0(gcm_dek_cmd_in[252]), .A1(n502), .Z(gcm_cmd_in[252]));
Q_AN02 U1198 ( .A0(n41), .A1(gcm_dak_cmd_in[252]), .Z(n502));
Q_MX02 U1199 ( .S(n39), .A0(gcm_dek_cmd_in[251]), .A1(n503), .Z(gcm_cmd_in[251]));
Q_AN02 U1200 ( .A0(n41), .A1(gcm_dak_cmd_in[251]), .Z(n503));
Q_MX02 U1201 ( .S(n39), .A0(gcm_dek_cmd_in[250]), .A1(n504), .Z(gcm_cmd_in[250]));
Q_AN02 U1202 ( .A0(n41), .A1(gcm_dak_cmd_in[250]), .Z(n504));
Q_MX02 U1203 ( .S(n39), .A0(gcm_dek_cmd_in[249]), .A1(n505), .Z(gcm_cmd_in[249]));
Q_AN02 U1204 ( .A0(n41), .A1(gcm_dak_cmd_in[249]), .Z(n505));
Q_MX02 U1205 ( .S(n39), .A0(gcm_dek_cmd_in[248]), .A1(n506), .Z(gcm_cmd_in[248]));
Q_AN02 U1206 ( .A0(n41), .A1(gcm_dak_cmd_in[248]), .Z(n506));
Q_MX02 U1207 ( .S(n39), .A0(gcm_dek_cmd_in[247]), .A1(n507), .Z(gcm_cmd_in[247]));
Q_AN02 U1208 ( .A0(n41), .A1(gcm_dak_cmd_in[247]), .Z(n507));
Q_MX02 U1209 ( .S(n39), .A0(gcm_dek_cmd_in[246]), .A1(n508), .Z(gcm_cmd_in[246]));
Q_AN02 U1210 ( .A0(n41), .A1(gcm_dak_cmd_in[246]), .Z(n508));
Q_MX02 U1211 ( .S(n39), .A0(gcm_dek_cmd_in[245]), .A1(n509), .Z(gcm_cmd_in[245]));
Q_AN02 U1212 ( .A0(n41), .A1(gcm_dak_cmd_in[245]), .Z(n509));
Q_MX02 U1213 ( .S(n39), .A0(gcm_dek_cmd_in[244]), .A1(n510), .Z(gcm_cmd_in[244]));
Q_AN02 U1214 ( .A0(n41), .A1(gcm_dak_cmd_in[244]), .Z(n510));
Q_MX02 U1215 ( .S(n39), .A0(gcm_dek_cmd_in[243]), .A1(n511), .Z(gcm_cmd_in[243]));
Q_AN02 U1216 ( .A0(n41), .A1(gcm_dak_cmd_in[243]), .Z(n511));
Q_MX02 U1217 ( .S(n39), .A0(gcm_dek_cmd_in[242]), .A1(n512), .Z(gcm_cmd_in[242]));
Q_AN02 U1218 ( .A0(n41), .A1(gcm_dak_cmd_in[242]), .Z(n512));
Q_MX02 U1219 ( .S(n39), .A0(gcm_dek_cmd_in[241]), .A1(n513), .Z(gcm_cmd_in[241]));
Q_AN02 U1220 ( .A0(n41), .A1(gcm_dak_cmd_in[241]), .Z(n513));
Q_MX02 U1221 ( .S(n39), .A0(gcm_dek_cmd_in[240]), .A1(n514), .Z(gcm_cmd_in[240]));
Q_AN02 U1222 ( .A0(n41), .A1(gcm_dak_cmd_in[240]), .Z(n514));
Q_MX02 U1223 ( .S(n39), .A0(gcm_dek_cmd_in[239]), .A1(n515), .Z(gcm_cmd_in[239]));
Q_AN02 U1224 ( .A0(n41), .A1(gcm_dak_cmd_in[239]), .Z(n515));
Q_MX02 U1225 ( .S(n39), .A0(gcm_dek_cmd_in[238]), .A1(n516), .Z(gcm_cmd_in[238]));
Q_AN02 U1226 ( .A0(n41), .A1(gcm_dak_cmd_in[238]), .Z(n516));
Q_MX02 U1227 ( .S(n39), .A0(gcm_dek_cmd_in[237]), .A1(n517), .Z(gcm_cmd_in[237]));
Q_AN02 U1228 ( .A0(n41), .A1(gcm_dak_cmd_in[237]), .Z(n517));
Q_MX02 U1229 ( .S(n39), .A0(gcm_dek_cmd_in[236]), .A1(n518), .Z(gcm_cmd_in[236]));
Q_AN02 U1230 ( .A0(n41), .A1(gcm_dak_cmd_in[236]), .Z(n518));
Q_MX02 U1231 ( .S(n39), .A0(gcm_dek_cmd_in[235]), .A1(n519), .Z(gcm_cmd_in[235]));
Q_AN02 U1232 ( .A0(n41), .A1(gcm_dak_cmd_in[235]), .Z(n519));
Q_MX02 U1233 ( .S(n39), .A0(gcm_dek_cmd_in[234]), .A1(n520), .Z(gcm_cmd_in[234]));
Q_AN02 U1234 ( .A0(n41), .A1(gcm_dak_cmd_in[234]), .Z(n520));
Q_MX02 U1235 ( .S(n39), .A0(gcm_dek_cmd_in[233]), .A1(n521), .Z(gcm_cmd_in[233]));
Q_AN02 U1236 ( .A0(n41), .A1(gcm_dak_cmd_in[233]), .Z(n521));
Q_MX02 U1237 ( .S(n39), .A0(gcm_dek_cmd_in[232]), .A1(n522), .Z(gcm_cmd_in[232]));
Q_AN02 U1238 ( .A0(n41), .A1(gcm_dak_cmd_in[232]), .Z(n522));
Q_MX02 U1239 ( .S(n39), .A0(gcm_dek_cmd_in[231]), .A1(n523), .Z(gcm_cmd_in[231]));
Q_AN02 U1240 ( .A0(n41), .A1(gcm_dak_cmd_in[231]), .Z(n523));
Q_MX02 U1241 ( .S(n39), .A0(gcm_dek_cmd_in[230]), .A1(n524), .Z(gcm_cmd_in[230]));
Q_AN02 U1242 ( .A0(n41), .A1(gcm_dak_cmd_in[230]), .Z(n524));
Q_MX02 U1243 ( .S(n39), .A0(gcm_dek_cmd_in[229]), .A1(n525), .Z(gcm_cmd_in[229]));
Q_AN02 U1244 ( .A0(n41), .A1(gcm_dak_cmd_in[229]), .Z(n525));
Q_MX02 U1245 ( .S(n39), .A0(gcm_dek_cmd_in[228]), .A1(n526), .Z(gcm_cmd_in[228]));
Q_AN02 U1246 ( .A0(n41), .A1(gcm_dak_cmd_in[228]), .Z(n526));
Q_MX02 U1247 ( .S(n39), .A0(gcm_dek_cmd_in[227]), .A1(n527), .Z(gcm_cmd_in[227]));
Q_AN02 U1248 ( .A0(n41), .A1(gcm_dak_cmd_in[227]), .Z(n527));
Q_MX02 U1249 ( .S(n39), .A0(gcm_dek_cmd_in[226]), .A1(n528), .Z(gcm_cmd_in[226]));
Q_AN02 U1250 ( .A0(n41), .A1(gcm_dak_cmd_in[226]), .Z(n528));
Q_MX02 U1251 ( .S(n39), .A0(gcm_dek_cmd_in[225]), .A1(n529), .Z(gcm_cmd_in[225]));
Q_AN02 U1252 ( .A0(n41), .A1(gcm_dak_cmd_in[225]), .Z(n529));
Q_MX02 U1253 ( .S(n39), .A0(gcm_dek_cmd_in[224]), .A1(n530), .Z(gcm_cmd_in[224]));
Q_AN02 U1254 ( .A0(n41), .A1(gcm_dak_cmd_in[224]), .Z(n530));
Q_MX02 U1255 ( .S(n39), .A0(gcm_dek_cmd_in[223]), .A1(n531), .Z(gcm_cmd_in[223]));
Q_AN02 U1256 ( .A0(n41), .A1(gcm_dak_cmd_in[223]), .Z(n531));
Q_MX02 U1257 ( .S(n39), .A0(gcm_dek_cmd_in[222]), .A1(n532), .Z(gcm_cmd_in[222]));
Q_AN02 U1258 ( .A0(n41), .A1(gcm_dak_cmd_in[222]), .Z(n532));
Q_MX02 U1259 ( .S(n39), .A0(gcm_dek_cmd_in[221]), .A1(n533), .Z(gcm_cmd_in[221]));
Q_AN02 U1260 ( .A0(n41), .A1(gcm_dak_cmd_in[221]), .Z(n533));
Q_MX02 U1261 ( .S(n39), .A0(gcm_dek_cmd_in[220]), .A1(n534), .Z(gcm_cmd_in[220]));
Q_AN02 U1262 ( .A0(n41), .A1(gcm_dak_cmd_in[220]), .Z(n534));
Q_MX02 U1263 ( .S(n39), .A0(gcm_dek_cmd_in[219]), .A1(n535), .Z(gcm_cmd_in[219]));
Q_AN02 U1264 ( .A0(n41), .A1(gcm_dak_cmd_in[219]), .Z(n535));
Q_MX02 U1265 ( .S(n39), .A0(gcm_dek_cmd_in[218]), .A1(n536), .Z(gcm_cmd_in[218]));
Q_AN02 U1266 ( .A0(n41), .A1(gcm_dak_cmd_in[218]), .Z(n536));
Q_MX02 U1267 ( .S(n39), .A0(gcm_dek_cmd_in[217]), .A1(n537), .Z(gcm_cmd_in[217]));
Q_AN02 U1268 ( .A0(n41), .A1(gcm_dak_cmd_in[217]), .Z(n537));
Q_MX02 U1269 ( .S(n39), .A0(gcm_dek_cmd_in[216]), .A1(n538), .Z(gcm_cmd_in[216]));
Q_AN02 U1270 ( .A0(n41), .A1(gcm_dak_cmd_in[216]), .Z(n538));
Q_MX02 U1271 ( .S(n39), .A0(gcm_dek_cmd_in[215]), .A1(n539), .Z(gcm_cmd_in[215]));
Q_AN02 U1272 ( .A0(n41), .A1(gcm_dak_cmd_in[215]), .Z(n539));
Q_MX02 U1273 ( .S(n39), .A0(gcm_dek_cmd_in[214]), .A1(n540), .Z(gcm_cmd_in[214]));
Q_AN02 U1274 ( .A0(n41), .A1(gcm_dak_cmd_in[214]), .Z(n540));
Q_MX02 U1275 ( .S(n39), .A0(gcm_dek_cmd_in[213]), .A1(n541), .Z(gcm_cmd_in[213]));
Q_AN02 U1276 ( .A0(n41), .A1(gcm_dak_cmd_in[213]), .Z(n541));
Q_MX02 U1277 ( .S(n39), .A0(gcm_dek_cmd_in[212]), .A1(n542), .Z(gcm_cmd_in[212]));
Q_AN02 U1278 ( .A0(n41), .A1(gcm_dak_cmd_in[212]), .Z(n542));
Q_MX02 U1279 ( .S(n39), .A0(gcm_dek_cmd_in[211]), .A1(n543), .Z(gcm_cmd_in[211]));
Q_AN02 U1280 ( .A0(n41), .A1(gcm_dak_cmd_in[211]), .Z(n543));
Q_MX02 U1281 ( .S(n39), .A0(gcm_dek_cmd_in[210]), .A1(n544), .Z(gcm_cmd_in[210]));
Q_AN02 U1282 ( .A0(n41), .A1(gcm_dak_cmd_in[210]), .Z(n544));
Q_MX02 U1283 ( .S(n39), .A0(gcm_dek_cmd_in[209]), .A1(n545), .Z(gcm_cmd_in[209]));
Q_AN02 U1284 ( .A0(n41), .A1(gcm_dak_cmd_in[209]), .Z(n545));
Q_MX02 U1285 ( .S(n39), .A0(gcm_dek_cmd_in[208]), .A1(n546), .Z(gcm_cmd_in[208]));
Q_AN02 U1286 ( .A0(n41), .A1(gcm_dak_cmd_in[208]), .Z(n546));
Q_MX02 U1287 ( .S(n39), .A0(gcm_dek_cmd_in[207]), .A1(n547), .Z(gcm_cmd_in[207]));
Q_AN02 U1288 ( .A0(n41), .A1(gcm_dak_cmd_in[207]), .Z(n547));
Q_MX02 U1289 ( .S(n39), .A0(gcm_dek_cmd_in[206]), .A1(n548), .Z(gcm_cmd_in[206]));
Q_AN02 U1290 ( .A0(n41), .A1(gcm_dak_cmd_in[206]), .Z(n548));
Q_MX02 U1291 ( .S(n39), .A0(gcm_dek_cmd_in[205]), .A1(n549), .Z(gcm_cmd_in[205]));
Q_AN02 U1292 ( .A0(n41), .A1(gcm_dak_cmd_in[205]), .Z(n549));
Q_MX02 U1293 ( .S(n39), .A0(gcm_dek_cmd_in[204]), .A1(n550), .Z(gcm_cmd_in[204]));
Q_AN02 U1294 ( .A0(n41), .A1(gcm_dak_cmd_in[204]), .Z(n550));
Q_MX02 U1295 ( .S(n39), .A0(gcm_dek_cmd_in[203]), .A1(n551), .Z(gcm_cmd_in[203]));
Q_AN02 U1296 ( .A0(n41), .A1(gcm_dak_cmd_in[203]), .Z(n551));
Q_MX02 U1297 ( .S(n39), .A0(gcm_dek_cmd_in[202]), .A1(n552), .Z(gcm_cmd_in[202]));
Q_AN02 U1298 ( .A0(n41), .A1(gcm_dak_cmd_in[202]), .Z(n552));
Q_MX02 U1299 ( .S(n39), .A0(gcm_dek_cmd_in[201]), .A1(n553), .Z(gcm_cmd_in[201]));
Q_AN02 U1300 ( .A0(n41), .A1(gcm_dak_cmd_in[201]), .Z(n553));
Q_MX02 U1301 ( .S(n39), .A0(gcm_dek_cmd_in[200]), .A1(n554), .Z(gcm_cmd_in[200]));
Q_AN02 U1302 ( .A0(n41), .A1(gcm_dak_cmd_in[200]), .Z(n554));
Q_MX02 U1303 ( .S(n39), .A0(gcm_dek_cmd_in[199]), .A1(n555), .Z(gcm_cmd_in[199]));
Q_AN02 U1304 ( .A0(n41), .A1(gcm_dak_cmd_in[199]), .Z(n555));
Q_MX02 U1305 ( .S(n39), .A0(gcm_dek_cmd_in[198]), .A1(n556), .Z(gcm_cmd_in[198]));
Q_AN02 U1306 ( .A0(n41), .A1(gcm_dak_cmd_in[198]), .Z(n556));
Q_MX02 U1307 ( .S(n39), .A0(gcm_dek_cmd_in[197]), .A1(n557), .Z(gcm_cmd_in[197]));
Q_AN02 U1308 ( .A0(n41), .A1(gcm_dak_cmd_in[197]), .Z(n557));
Q_MX02 U1309 ( .S(n39), .A0(gcm_dek_cmd_in[196]), .A1(n558), .Z(gcm_cmd_in[196]));
Q_AN02 U1310 ( .A0(n41), .A1(gcm_dak_cmd_in[196]), .Z(n558));
Q_MX02 U1311 ( .S(n39), .A0(gcm_dek_cmd_in[195]), .A1(n559), .Z(gcm_cmd_in[195]));
Q_AN02 U1312 ( .A0(n41), .A1(gcm_dak_cmd_in[195]), .Z(n559));
Q_MX02 U1313 ( .S(n39), .A0(gcm_dek_cmd_in[194]), .A1(n560), .Z(gcm_cmd_in[194]));
Q_AN02 U1314 ( .A0(n41), .A1(gcm_dak_cmd_in[194]), .Z(n560));
Q_MX02 U1315 ( .S(n39), .A0(gcm_dek_cmd_in[193]), .A1(n561), .Z(gcm_cmd_in[193]));
Q_AN02 U1316 ( .A0(n41), .A1(gcm_dak_cmd_in[193]), .Z(n561));
Q_MX02 U1317 ( .S(n39), .A0(gcm_dek_cmd_in[192]), .A1(n562), .Z(gcm_cmd_in[192]));
Q_AN02 U1318 ( .A0(n41), .A1(gcm_dak_cmd_in[192]), .Z(n562));
Q_MX02 U1319 ( .S(n39), .A0(gcm_dek_cmd_in[191]), .A1(n563), .Z(gcm_cmd_in[191]));
Q_AN02 U1320 ( .A0(n41), .A1(gcm_dak_cmd_in[191]), .Z(n563));
Q_MX02 U1321 ( .S(n39), .A0(gcm_dek_cmd_in[190]), .A1(n564), .Z(gcm_cmd_in[190]));
Q_AN02 U1322 ( .A0(n41), .A1(gcm_dak_cmd_in[190]), .Z(n564));
Q_MX02 U1323 ( .S(n39), .A0(gcm_dek_cmd_in[189]), .A1(n565), .Z(gcm_cmd_in[189]));
Q_AN02 U1324 ( .A0(n41), .A1(gcm_dak_cmd_in[189]), .Z(n565));
Q_MX02 U1325 ( .S(n39), .A0(gcm_dek_cmd_in[188]), .A1(n566), .Z(gcm_cmd_in[188]));
Q_AN02 U1326 ( .A0(n41), .A1(gcm_dak_cmd_in[188]), .Z(n566));
Q_MX02 U1327 ( .S(n39), .A0(gcm_dek_cmd_in[187]), .A1(n567), .Z(gcm_cmd_in[187]));
Q_AN02 U1328 ( .A0(n41), .A1(gcm_dak_cmd_in[187]), .Z(n567));
Q_MX02 U1329 ( .S(n39), .A0(gcm_dek_cmd_in[186]), .A1(n568), .Z(gcm_cmd_in[186]));
Q_AN02 U1330 ( .A0(n41), .A1(gcm_dak_cmd_in[186]), .Z(n568));
Q_MX02 U1331 ( .S(n39), .A0(gcm_dek_cmd_in[185]), .A1(n569), .Z(gcm_cmd_in[185]));
Q_AN02 U1332 ( .A0(n41), .A1(gcm_dak_cmd_in[185]), .Z(n569));
Q_MX02 U1333 ( .S(n39), .A0(gcm_dek_cmd_in[184]), .A1(n570), .Z(gcm_cmd_in[184]));
Q_AN02 U1334 ( .A0(n41), .A1(gcm_dak_cmd_in[184]), .Z(n570));
Q_MX02 U1335 ( .S(n39), .A0(gcm_dek_cmd_in[183]), .A1(n571), .Z(gcm_cmd_in[183]));
Q_AN02 U1336 ( .A0(n41), .A1(gcm_dak_cmd_in[183]), .Z(n571));
Q_MX02 U1337 ( .S(n39), .A0(gcm_dek_cmd_in[182]), .A1(n572), .Z(gcm_cmd_in[182]));
Q_AN02 U1338 ( .A0(n41), .A1(gcm_dak_cmd_in[182]), .Z(n572));
Q_MX02 U1339 ( .S(n39), .A0(gcm_dek_cmd_in[181]), .A1(n573), .Z(gcm_cmd_in[181]));
Q_AN02 U1340 ( .A0(n41), .A1(gcm_dak_cmd_in[181]), .Z(n573));
Q_MX02 U1341 ( .S(n39), .A0(gcm_dek_cmd_in[180]), .A1(n574), .Z(gcm_cmd_in[180]));
Q_AN02 U1342 ( .A0(n41), .A1(gcm_dak_cmd_in[180]), .Z(n574));
Q_MX02 U1343 ( .S(n39), .A0(gcm_dek_cmd_in[179]), .A1(n575), .Z(gcm_cmd_in[179]));
Q_AN02 U1344 ( .A0(n41), .A1(gcm_dak_cmd_in[179]), .Z(n575));
Q_MX02 U1345 ( .S(n39), .A0(gcm_dek_cmd_in[178]), .A1(n576), .Z(gcm_cmd_in[178]));
Q_AN02 U1346 ( .A0(n41), .A1(gcm_dak_cmd_in[178]), .Z(n576));
Q_MX02 U1347 ( .S(n39), .A0(gcm_dek_cmd_in[177]), .A1(n577), .Z(gcm_cmd_in[177]));
Q_AN02 U1348 ( .A0(n41), .A1(gcm_dak_cmd_in[177]), .Z(n577));
Q_MX02 U1349 ( .S(n39), .A0(gcm_dek_cmd_in[176]), .A1(n578), .Z(gcm_cmd_in[176]));
Q_AN02 U1350 ( .A0(n41), .A1(gcm_dak_cmd_in[176]), .Z(n578));
Q_MX02 U1351 ( .S(n39), .A0(gcm_dek_cmd_in[175]), .A1(n579), .Z(gcm_cmd_in[175]));
Q_AN02 U1352 ( .A0(n41), .A1(gcm_dak_cmd_in[175]), .Z(n579));
Q_MX02 U1353 ( .S(n39), .A0(gcm_dek_cmd_in[174]), .A1(n580), .Z(gcm_cmd_in[174]));
Q_AN02 U1354 ( .A0(n41), .A1(gcm_dak_cmd_in[174]), .Z(n580));
Q_MX02 U1355 ( .S(n39), .A0(gcm_dek_cmd_in[173]), .A1(n581), .Z(gcm_cmd_in[173]));
Q_AN02 U1356 ( .A0(n41), .A1(gcm_dak_cmd_in[173]), .Z(n581));
Q_MX02 U1357 ( .S(n39), .A0(gcm_dek_cmd_in[172]), .A1(n582), .Z(gcm_cmd_in[172]));
Q_AN02 U1358 ( .A0(n41), .A1(gcm_dak_cmd_in[172]), .Z(n582));
Q_MX02 U1359 ( .S(n39), .A0(gcm_dek_cmd_in[171]), .A1(n583), .Z(gcm_cmd_in[171]));
Q_AN02 U1360 ( .A0(n41), .A1(gcm_dak_cmd_in[171]), .Z(n583));
Q_MX02 U1361 ( .S(n39), .A0(gcm_dek_cmd_in[170]), .A1(n584), .Z(gcm_cmd_in[170]));
Q_AN02 U1362 ( .A0(n41), .A1(gcm_dak_cmd_in[170]), .Z(n584));
Q_MX02 U1363 ( .S(n39), .A0(gcm_dek_cmd_in[169]), .A1(n585), .Z(gcm_cmd_in[169]));
Q_AN02 U1364 ( .A0(n41), .A1(gcm_dak_cmd_in[169]), .Z(n585));
Q_MX02 U1365 ( .S(n39), .A0(gcm_dek_cmd_in[168]), .A1(n586), .Z(gcm_cmd_in[168]));
Q_AN02 U1366 ( .A0(n41), .A1(gcm_dak_cmd_in[168]), .Z(n586));
Q_MX02 U1367 ( .S(n39), .A0(gcm_dek_cmd_in[167]), .A1(n587), .Z(gcm_cmd_in[167]));
Q_AN02 U1368 ( .A0(n41), .A1(gcm_dak_cmd_in[167]), .Z(n587));
Q_MX02 U1369 ( .S(n39), .A0(gcm_dek_cmd_in[166]), .A1(n588), .Z(gcm_cmd_in[166]));
Q_AN02 U1370 ( .A0(n41), .A1(gcm_dak_cmd_in[166]), .Z(n588));
Q_MX02 U1371 ( .S(n39), .A0(gcm_dek_cmd_in[165]), .A1(n589), .Z(gcm_cmd_in[165]));
Q_AN02 U1372 ( .A0(n41), .A1(gcm_dak_cmd_in[165]), .Z(n589));
Q_MX02 U1373 ( .S(n39), .A0(gcm_dek_cmd_in[164]), .A1(n590), .Z(gcm_cmd_in[164]));
Q_AN02 U1374 ( .A0(n41), .A1(gcm_dak_cmd_in[164]), .Z(n590));
Q_MX02 U1375 ( .S(n39), .A0(gcm_dek_cmd_in[163]), .A1(n591), .Z(gcm_cmd_in[163]));
Q_AN02 U1376 ( .A0(n41), .A1(gcm_dak_cmd_in[163]), .Z(n591));
Q_MX02 U1377 ( .S(n39), .A0(gcm_dek_cmd_in[162]), .A1(n592), .Z(gcm_cmd_in[162]));
Q_AN02 U1378 ( .A0(n41), .A1(gcm_dak_cmd_in[162]), .Z(n592));
Q_MX02 U1379 ( .S(n39), .A0(gcm_dek_cmd_in[161]), .A1(n593), .Z(gcm_cmd_in[161]));
Q_AN02 U1380 ( .A0(n41), .A1(gcm_dak_cmd_in[161]), .Z(n593));
Q_MX02 U1381 ( .S(n39), .A0(gcm_dek_cmd_in[160]), .A1(n594), .Z(gcm_cmd_in[160]));
Q_AN02 U1382 ( .A0(n41), .A1(gcm_dak_cmd_in[160]), .Z(n594));
Q_MX02 U1383 ( .S(n39), .A0(gcm_dek_cmd_in[159]), .A1(n595), .Z(gcm_cmd_in[159]));
Q_AN02 U1384 ( .A0(n41), .A1(gcm_dak_cmd_in[159]), .Z(n595));
Q_MX02 U1385 ( .S(n39), .A0(gcm_dek_cmd_in[158]), .A1(n596), .Z(gcm_cmd_in[158]));
Q_AN02 U1386 ( .A0(n41), .A1(gcm_dak_cmd_in[158]), .Z(n596));
Q_MX02 U1387 ( .S(n39), .A0(gcm_dek_cmd_in[157]), .A1(n597), .Z(gcm_cmd_in[157]));
Q_AN02 U1388 ( .A0(n41), .A1(gcm_dak_cmd_in[157]), .Z(n597));
Q_MX02 U1389 ( .S(n39), .A0(gcm_dek_cmd_in[156]), .A1(n598), .Z(gcm_cmd_in[156]));
Q_AN02 U1390 ( .A0(n41), .A1(gcm_dak_cmd_in[156]), .Z(n598));
Q_MX02 U1391 ( .S(n39), .A0(gcm_dek_cmd_in[155]), .A1(n599), .Z(gcm_cmd_in[155]));
Q_AN02 U1392 ( .A0(n41), .A1(gcm_dak_cmd_in[155]), .Z(n599));
Q_MX02 U1393 ( .S(n39), .A0(gcm_dek_cmd_in[154]), .A1(n600), .Z(gcm_cmd_in[154]));
Q_AN02 U1394 ( .A0(n41), .A1(gcm_dak_cmd_in[154]), .Z(n600));
Q_MX02 U1395 ( .S(n39), .A0(gcm_dek_cmd_in[153]), .A1(n601), .Z(gcm_cmd_in[153]));
Q_AN02 U1396 ( .A0(n41), .A1(gcm_dak_cmd_in[153]), .Z(n601));
Q_MX02 U1397 ( .S(n39), .A0(gcm_dek_cmd_in[152]), .A1(n602), .Z(gcm_cmd_in[152]));
Q_AN02 U1398 ( .A0(n41), .A1(gcm_dak_cmd_in[152]), .Z(n602));
Q_MX02 U1399 ( .S(n39), .A0(gcm_dek_cmd_in[151]), .A1(n603), .Z(gcm_cmd_in[151]));
Q_AN02 U1400 ( .A0(n41), .A1(gcm_dak_cmd_in[151]), .Z(n603));
Q_MX02 U1401 ( .S(n39), .A0(gcm_dek_cmd_in[150]), .A1(n604), .Z(gcm_cmd_in[150]));
Q_AN02 U1402 ( .A0(n41), .A1(gcm_dak_cmd_in[150]), .Z(n604));
Q_MX02 U1403 ( .S(n39), .A0(gcm_dek_cmd_in[149]), .A1(n605), .Z(gcm_cmd_in[149]));
Q_AN02 U1404 ( .A0(n41), .A1(gcm_dak_cmd_in[149]), .Z(n605));
Q_MX02 U1405 ( .S(n39), .A0(gcm_dek_cmd_in[148]), .A1(n606), .Z(gcm_cmd_in[148]));
Q_AN02 U1406 ( .A0(n41), .A1(gcm_dak_cmd_in[148]), .Z(n606));
Q_MX02 U1407 ( .S(n39), .A0(gcm_dek_cmd_in[147]), .A1(n607), .Z(gcm_cmd_in[147]));
Q_AN02 U1408 ( .A0(n41), .A1(gcm_dak_cmd_in[147]), .Z(n607));
Q_MX02 U1409 ( .S(n39), .A0(gcm_dek_cmd_in[146]), .A1(n608), .Z(gcm_cmd_in[146]));
Q_AN02 U1410 ( .A0(n41), .A1(gcm_dak_cmd_in[146]), .Z(n608));
Q_MX02 U1411 ( .S(n39), .A0(gcm_dek_cmd_in[145]), .A1(n609), .Z(gcm_cmd_in[145]));
Q_AN02 U1412 ( .A0(n41), .A1(gcm_dak_cmd_in[145]), .Z(n609));
Q_MX02 U1413 ( .S(n39), .A0(gcm_dek_cmd_in[144]), .A1(n610), .Z(gcm_cmd_in[144]));
Q_AN02 U1414 ( .A0(n41), .A1(gcm_dak_cmd_in[144]), .Z(n610));
Q_MX02 U1415 ( .S(n39), .A0(gcm_dek_cmd_in[143]), .A1(n611), .Z(gcm_cmd_in[143]));
Q_AN02 U1416 ( .A0(n41), .A1(gcm_dak_cmd_in[143]), .Z(n611));
Q_MX02 U1417 ( .S(n39), .A0(gcm_dek_cmd_in[142]), .A1(n612), .Z(gcm_cmd_in[142]));
Q_AN02 U1418 ( .A0(n41), .A1(gcm_dak_cmd_in[142]), .Z(n612));
Q_MX02 U1419 ( .S(n39), .A0(gcm_dek_cmd_in[141]), .A1(n613), .Z(gcm_cmd_in[141]));
Q_AN02 U1420 ( .A0(n41), .A1(gcm_dak_cmd_in[141]), .Z(n613));
Q_MX02 U1421 ( .S(n39), .A0(gcm_dek_cmd_in[140]), .A1(n614), .Z(gcm_cmd_in[140]));
Q_AN02 U1422 ( .A0(n41), .A1(gcm_dak_cmd_in[140]), .Z(n614));
Q_MX02 U1423 ( .S(n39), .A0(gcm_dek_cmd_in[139]), .A1(n615), .Z(gcm_cmd_in[139]));
Q_AN02 U1424 ( .A0(n41), .A1(gcm_dak_cmd_in[139]), .Z(n615));
Q_MX02 U1425 ( .S(n39), .A0(gcm_dek_cmd_in[138]), .A1(n616), .Z(gcm_cmd_in[138]));
Q_AN02 U1426 ( .A0(n41), .A1(gcm_dak_cmd_in[138]), .Z(n616));
Q_MX02 U1427 ( .S(n39), .A0(gcm_dek_cmd_in[137]), .A1(n617), .Z(gcm_cmd_in[137]));
Q_AN02 U1428 ( .A0(n41), .A1(gcm_dak_cmd_in[137]), .Z(n617));
Q_MX02 U1429 ( .S(n39), .A0(gcm_dek_cmd_in[136]), .A1(n618), .Z(gcm_cmd_in[136]));
Q_AN02 U1430 ( .A0(n41), .A1(gcm_dak_cmd_in[136]), .Z(n618));
Q_MX02 U1431 ( .S(n39), .A0(gcm_dek_cmd_in[135]), .A1(n619), .Z(gcm_cmd_in[135]));
Q_AN02 U1432 ( .A0(n41), .A1(gcm_dak_cmd_in[135]), .Z(n619));
Q_MX02 U1433 ( .S(n39), .A0(gcm_dek_cmd_in[134]), .A1(n620), .Z(gcm_cmd_in[134]));
Q_AN02 U1434 ( .A0(n41), .A1(gcm_dak_cmd_in[134]), .Z(n620));
Q_MX02 U1435 ( .S(n39), .A0(gcm_dek_cmd_in[133]), .A1(n621), .Z(gcm_cmd_in[133]));
Q_AN02 U1436 ( .A0(n41), .A1(gcm_dak_cmd_in[133]), .Z(n621));
Q_MX02 U1437 ( .S(n39), .A0(gcm_dek_cmd_in[132]), .A1(n622), .Z(gcm_cmd_in[132]));
Q_AN02 U1438 ( .A0(n41), .A1(gcm_dak_cmd_in[132]), .Z(n622));
Q_MX02 U1439 ( .S(n39), .A0(gcm_dek_cmd_in[131]), .A1(n623), .Z(gcm_cmd_in[131]));
Q_AN02 U1440 ( .A0(n41), .A1(gcm_dak_cmd_in[131]), .Z(n623));
Q_MX02 U1441 ( .S(n39), .A0(gcm_dek_cmd_in[130]), .A1(n624), .Z(gcm_cmd_in[130]));
Q_AN02 U1442 ( .A0(n41), .A1(gcm_dak_cmd_in[130]), .Z(n624));
Q_MX02 U1443 ( .S(n39), .A0(gcm_dek_cmd_in[129]), .A1(n625), .Z(gcm_cmd_in[129]));
Q_AN02 U1444 ( .A0(n41), .A1(gcm_dak_cmd_in[129]), .Z(n625));
Q_MX02 U1445 ( .S(n39), .A0(gcm_dek_cmd_in[128]), .A1(n626), .Z(gcm_cmd_in[128]));
Q_AN02 U1446 ( .A0(n41), .A1(gcm_dak_cmd_in[128]), .Z(n626));
Q_MX02 U1447 ( .S(n39), .A0(gcm_dek_cmd_in[127]), .A1(n627), .Z(gcm_cmd_in[127]));
Q_AN02 U1448 ( .A0(n41), .A1(gcm_dak_cmd_in[127]), .Z(n627));
Q_MX02 U1449 ( .S(n39), .A0(gcm_dek_cmd_in[126]), .A1(n628), .Z(gcm_cmd_in[126]));
Q_AN02 U1450 ( .A0(n41), .A1(gcm_dak_cmd_in[126]), .Z(n628));
Q_MX02 U1451 ( .S(n39), .A0(gcm_dek_cmd_in[125]), .A1(n629), .Z(gcm_cmd_in[125]));
Q_AN02 U1452 ( .A0(n41), .A1(gcm_dak_cmd_in[125]), .Z(n629));
Q_MX02 U1453 ( .S(n39), .A0(gcm_dek_cmd_in[124]), .A1(n630), .Z(gcm_cmd_in[124]));
Q_AN02 U1454 ( .A0(n41), .A1(gcm_dak_cmd_in[124]), .Z(n630));
Q_MX02 U1455 ( .S(n39), .A0(gcm_dek_cmd_in[123]), .A1(n631), .Z(gcm_cmd_in[123]));
Q_AN02 U1456 ( .A0(n41), .A1(gcm_dak_cmd_in[123]), .Z(n631));
Q_MX02 U1457 ( .S(n39), .A0(gcm_dek_cmd_in[122]), .A1(n632), .Z(gcm_cmd_in[122]));
Q_AN02 U1458 ( .A0(n41), .A1(gcm_dak_cmd_in[122]), .Z(n632));
Q_MX02 U1459 ( .S(n39), .A0(gcm_dek_cmd_in[121]), .A1(n633), .Z(gcm_cmd_in[121]));
Q_AN02 U1460 ( .A0(n41), .A1(gcm_dak_cmd_in[121]), .Z(n633));
Q_MX02 U1461 ( .S(n39), .A0(gcm_dek_cmd_in[120]), .A1(n634), .Z(gcm_cmd_in[120]));
Q_AN02 U1462 ( .A0(n41), .A1(gcm_dak_cmd_in[120]), .Z(n634));
Q_MX02 U1463 ( .S(n39), .A0(gcm_dek_cmd_in[119]), .A1(n635), .Z(gcm_cmd_in[119]));
Q_AN02 U1464 ( .A0(n41), .A1(gcm_dak_cmd_in[119]), .Z(n635));
Q_MX02 U1465 ( .S(n39), .A0(gcm_dek_cmd_in[118]), .A1(n636), .Z(gcm_cmd_in[118]));
Q_AN02 U1466 ( .A0(n41), .A1(gcm_dak_cmd_in[118]), .Z(n636));
Q_MX02 U1467 ( .S(n39), .A0(gcm_dek_cmd_in[117]), .A1(n637), .Z(gcm_cmd_in[117]));
Q_AN02 U1468 ( .A0(n41), .A1(gcm_dak_cmd_in[117]), .Z(n637));
Q_MX02 U1469 ( .S(n39), .A0(gcm_dek_cmd_in[116]), .A1(n638), .Z(gcm_cmd_in[116]));
Q_AN02 U1470 ( .A0(n41), .A1(gcm_dak_cmd_in[116]), .Z(n638));
Q_MX02 U1471 ( .S(n39), .A0(gcm_dek_cmd_in[115]), .A1(n639), .Z(gcm_cmd_in[115]));
Q_AN02 U1472 ( .A0(n41), .A1(gcm_dak_cmd_in[115]), .Z(n639));
Q_MX02 U1473 ( .S(n39), .A0(gcm_dek_cmd_in[114]), .A1(n640), .Z(gcm_cmd_in[114]));
Q_AN02 U1474 ( .A0(n41), .A1(gcm_dak_cmd_in[114]), .Z(n640));
Q_MX02 U1475 ( .S(n39), .A0(gcm_dek_cmd_in[113]), .A1(n641), .Z(gcm_cmd_in[113]));
Q_AN02 U1476 ( .A0(n41), .A1(gcm_dak_cmd_in[113]), .Z(n641));
Q_MX02 U1477 ( .S(n39), .A0(gcm_dek_cmd_in[112]), .A1(n642), .Z(gcm_cmd_in[112]));
Q_AN02 U1478 ( .A0(n41), .A1(gcm_dak_cmd_in[112]), .Z(n642));
Q_MX02 U1479 ( .S(n39), .A0(gcm_dek_cmd_in[111]), .A1(n643), .Z(gcm_cmd_in[111]));
Q_AN02 U1480 ( .A0(n41), .A1(gcm_dak_cmd_in[111]), .Z(n643));
Q_MX02 U1481 ( .S(n39), .A0(gcm_dek_cmd_in[110]), .A1(n644), .Z(gcm_cmd_in[110]));
Q_AN02 U1482 ( .A0(n41), .A1(gcm_dak_cmd_in[110]), .Z(n644));
Q_MX02 U1483 ( .S(n39), .A0(gcm_dek_cmd_in[109]), .A1(n645), .Z(gcm_cmd_in[109]));
Q_AN02 U1484 ( .A0(n41), .A1(gcm_dak_cmd_in[109]), .Z(n645));
Q_MX02 U1485 ( .S(n39), .A0(gcm_dek_cmd_in[108]), .A1(n646), .Z(gcm_cmd_in[108]));
Q_AN02 U1486 ( .A0(n41), .A1(gcm_dak_cmd_in[108]), .Z(n646));
Q_MX02 U1487 ( .S(n39), .A0(gcm_dek_cmd_in[107]), .A1(n647), .Z(gcm_cmd_in[107]));
Q_AN02 U1488 ( .A0(n41), .A1(gcm_dak_cmd_in[107]), .Z(n647));
Q_MX02 U1489 ( .S(n39), .A0(gcm_dek_cmd_in[106]), .A1(n648), .Z(gcm_cmd_in[106]));
Q_AN02 U1490 ( .A0(n41), .A1(gcm_dak_cmd_in[106]), .Z(n648));
Q_MX02 U1491 ( .S(n39), .A0(gcm_dek_cmd_in[105]), .A1(n649), .Z(gcm_cmd_in[105]));
Q_AN02 U1492 ( .A0(n41), .A1(gcm_dak_cmd_in[105]), .Z(n649));
Q_MX02 U1493 ( .S(n39), .A0(gcm_dek_cmd_in[104]), .A1(n650), .Z(gcm_cmd_in[104]));
Q_AN02 U1494 ( .A0(n41), .A1(gcm_dak_cmd_in[104]), .Z(n650));
Q_MX02 U1495 ( .S(n39), .A0(gcm_dek_cmd_in[103]), .A1(n651), .Z(gcm_cmd_in[103]));
Q_AN02 U1496 ( .A0(n41), .A1(gcm_dak_cmd_in[103]), .Z(n651));
Q_MX02 U1497 ( .S(n39), .A0(gcm_dek_cmd_in[102]), .A1(n652), .Z(gcm_cmd_in[102]));
Q_AN02 U1498 ( .A0(n41), .A1(gcm_dak_cmd_in[102]), .Z(n652));
Q_MX02 U1499 ( .S(n39), .A0(gcm_dek_cmd_in[101]), .A1(n653), .Z(gcm_cmd_in[101]));
Q_AN02 U1500 ( .A0(n41), .A1(gcm_dak_cmd_in[101]), .Z(n653));
Q_MX02 U1501 ( .S(n39), .A0(gcm_dek_cmd_in[100]), .A1(n654), .Z(gcm_cmd_in[100]));
Q_AN02 U1502 ( .A0(n41), .A1(gcm_dak_cmd_in[100]), .Z(n654));
Q_MX02 U1503 ( .S(n39), .A0(gcm_dek_cmd_in[99]), .A1(n655), .Z(gcm_cmd_in[99]));
Q_AN02 U1504 ( .A0(n41), .A1(gcm_dak_cmd_in[99]), .Z(n655));
Q_MX02 U1505 ( .S(n39), .A0(n2653), .A1(n656), .Z(gcm_cmd_in[98]));
Q_AN02 U1506 ( .A0(n41), .A1(n2557), .Z(n656));
Q_MX02 U1507 ( .S(n39), .A0(n2654), .A1(n657), .Z(gcm_cmd_in[97]));
Q_AN02 U1508 ( .A0(n41), .A1(n2558), .Z(n657));
Q_MX02 U1509 ( .S(n39), .A0(n2655), .A1(n658), .Z(gcm_cmd_in[96]));
Q_AN02 U1510 ( .A0(n41), .A1(n2559), .Z(n658));
Q_MX02 U1511 ( .S(n39), .A0(n2656), .A1(n659), .Z(gcm_cmd_in[95]));
Q_AN02 U1512 ( .A0(n41), .A1(n2560), .Z(n659));
Q_MX02 U1513 ( .S(n39), .A0(n2657), .A1(n660), .Z(gcm_cmd_in[94]));
Q_AN02 U1514 ( .A0(n41), .A1(n2561), .Z(n660));
Q_MX02 U1515 ( .S(n39), .A0(n2658), .A1(n661), .Z(gcm_cmd_in[93]));
Q_AN02 U1516 ( .A0(n41), .A1(n2562), .Z(n661));
Q_MX02 U1517 ( .S(n39), .A0(n2659), .A1(n662), .Z(gcm_cmd_in[92]));
Q_AN02 U1518 ( .A0(n41), .A1(n2563), .Z(n662));
Q_MX02 U1519 ( .S(n39), .A0(n2660), .A1(n663), .Z(gcm_cmd_in[91]));
Q_AN02 U1520 ( .A0(n41), .A1(n2564), .Z(n663));
Q_MX02 U1521 ( .S(n39), .A0(n2661), .A1(n664), .Z(gcm_cmd_in[90]));
Q_AN02 U1522 ( .A0(n41), .A1(n2565), .Z(n664));
Q_MX02 U1523 ( .S(n39), .A0(n2662), .A1(n665), .Z(gcm_cmd_in[89]));
Q_AN02 U1524 ( .A0(n41), .A1(n2566), .Z(n665));
Q_MX02 U1525 ( .S(n39), .A0(n2663), .A1(n666), .Z(gcm_cmd_in[88]));
Q_AN02 U1526 ( .A0(n41), .A1(n2567), .Z(n666));
Q_MX02 U1527 ( .S(n39), .A0(n2664), .A1(n667), .Z(gcm_cmd_in[87]));
Q_AN02 U1528 ( .A0(n41), .A1(n2568), .Z(n667));
Q_MX02 U1529 ( .S(n39), .A0(n2665), .A1(n668), .Z(gcm_cmd_in[86]));
Q_AN02 U1530 ( .A0(n41), .A1(n2569), .Z(n668));
Q_MX02 U1531 ( .S(n39), .A0(n2666), .A1(n669), .Z(gcm_cmd_in[85]));
Q_AN02 U1532 ( .A0(n41), .A1(n2570), .Z(n669));
Q_MX02 U1533 ( .S(n39), .A0(n2667), .A1(n670), .Z(gcm_cmd_in[84]));
Q_AN02 U1534 ( .A0(n41), .A1(n2571), .Z(n670));
Q_MX02 U1535 ( .S(n39), .A0(n2668), .A1(n671), .Z(gcm_cmd_in[83]));
Q_AN02 U1536 ( .A0(n41), .A1(n2572), .Z(n671));
Q_MX02 U1537 ( .S(n39), .A0(n2669), .A1(n672), .Z(gcm_cmd_in[82]));
Q_AN02 U1538 ( .A0(n41), .A1(n2573), .Z(n672));
Q_MX02 U1539 ( .S(n39), .A0(n2670), .A1(n673), .Z(gcm_cmd_in[81]));
Q_AN02 U1540 ( .A0(n41), .A1(n2574), .Z(n673));
Q_MX02 U1541 ( .S(n39), .A0(n2671), .A1(n674), .Z(gcm_cmd_in[80]));
Q_AN02 U1542 ( .A0(n41), .A1(n2575), .Z(n674));
Q_MX02 U1543 ( .S(n39), .A0(n2672), .A1(n675), .Z(gcm_cmd_in[79]));
Q_AN02 U1544 ( .A0(n41), .A1(n2576), .Z(n675));
Q_MX02 U1545 ( .S(n39), .A0(n2673), .A1(n676), .Z(gcm_cmd_in[78]));
Q_AN02 U1546 ( .A0(n41), .A1(n2577), .Z(n676));
Q_MX02 U1547 ( .S(n39), .A0(n2674), .A1(n677), .Z(gcm_cmd_in[77]));
Q_AN02 U1548 ( .A0(n41), .A1(n2578), .Z(n677));
Q_MX02 U1549 ( .S(n39), .A0(n2675), .A1(n678), .Z(gcm_cmd_in[76]));
Q_AN02 U1550 ( .A0(n41), .A1(n2579), .Z(n678));
Q_MX02 U1551 ( .S(n39), .A0(n2676), .A1(n679), .Z(gcm_cmd_in[75]));
Q_AN02 U1552 ( .A0(n41), .A1(n2580), .Z(n679));
Q_MX02 U1553 ( .S(n39), .A0(n2677), .A1(n680), .Z(gcm_cmd_in[74]));
Q_AN02 U1554 ( .A0(n41), .A1(n2581), .Z(n680));
Q_MX02 U1555 ( .S(n39), .A0(n2678), .A1(n681), .Z(gcm_cmd_in[73]));
Q_AN02 U1556 ( .A0(n41), .A1(n2582), .Z(n681));
Q_MX02 U1557 ( .S(n39), .A0(n2679), .A1(n682), .Z(gcm_cmd_in[72]));
Q_AN02 U1558 ( .A0(n41), .A1(n2583), .Z(n682));
Q_MX02 U1559 ( .S(n39), .A0(n2680), .A1(n683), .Z(gcm_cmd_in[71]));
Q_AN02 U1560 ( .A0(n41), .A1(n2584), .Z(n683));
Q_MX02 U1561 ( .S(n39), .A0(n2681), .A1(n684), .Z(gcm_cmd_in[70]));
Q_AN02 U1562 ( .A0(n41), .A1(n2585), .Z(n684));
Q_MX02 U1563 ( .S(n39), .A0(n2682), .A1(n685), .Z(gcm_cmd_in[69]));
Q_AN02 U1564 ( .A0(n41), .A1(n2586), .Z(n685));
Q_MX02 U1565 ( .S(n39), .A0(n2683), .A1(n686), .Z(gcm_cmd_in[68]));
Q_AN02 U1566 ( .A0(n41), .A1(n2587), .Z(n686));
Q_MX02 U1567 ( .S(n39), .A0(n2684), .A1(n687), .Z(gcm_cmd_in[67]));
Q_AN02 U1568 ( .A0(n41), .A1(n2588), .Z(n687));
Q_MX02 U1569 ( .S(n39), .A0(n2685), .A1(n688), .Z(gcm_cmd_in[66]));
Q_AN02 U1570 ( .A0(n41), .A1(n2589), .Z(n688));
Q_MX02 U1571 ( .S(n39), .A0(n2686), .A1(n689), .Z(gcm_cmd_in[65]));
Q_AN02 U1572 ( .A0(n41), .A1(n2590), .Z(n689));
Q_MX02 U1573 ( .S(n39), .A0(n2687), .A1(n690), .Z(gcm_cmd_in[64]));
Q_AN02 U1574 ( .A0(n41), .A1(n2591), .Z(n690));
Q_MX02 U1575 ( .S(n39), .A0(n2688), .A1(n691), .Z(gcm_cmd_in[63]));
Q_AN02 U1576 ( .A0(n41), .A1(n2592), .Z(n691));
Q_MX02 U1577 ( .S(n39), .A0(n2689), .A1(n692), .Z(gcm_cmd_in[62]));
Q_AN02 U1578 ( .A0(n41), .A1(n2593), .Z(n692));
Q_MX02 U1579 ( .S(n39), .A0(n2690), .A1(n693), .Z(gcm_cmd_in[61]));
Q_AN02 U1580 ( .A0(n41), .A1(n2594), .Z(n693));
Q_MX02 U1581 ( .S(n39), .A0(n2691), .A1(n694), .Z(gcm_cmd_in[60]));
Q_AN02 U1582 ( .A0(n41), .A1(n2595), .Z(n694));
Q_MX02 U1583 ( .S(n39), .A0(n2692), .A1(n695), .Z(gcm_cmd_in[59]));
Q_AN02 U1584 ( .A0(n41), .A1(n2596), .Z(n695));
Q_MX02 U1585 ( .S(n39), .A0(n2693), .A1(n696), .Z(gcm_cmd_in[58]));
Q_AN02 U1586 ( .A0(n41), .A1(n2597), .Z(n696));
Q_MX02 U1587 ( .S(n39), .A0(n2694), .A1(n697), .Z(gcm_cmd_in[57]));
Q_AN02 U1588 ( .A0(n41), .A1(n2598), .Z(n697));
Q_MX02 U1589 ( .S(n39), .A0(n2695), .A1(n698), .Z(gcm_cmd_in[56]));
Q_AN02 U1590 ( .A0(n41), .A1(n2599), .Z(n698));
Q_MX02 U1591 ( .S(n39), .A0(n2696), .A1(n699), .Z(gcm_cmd_in[55]));
Q_AN02 U1592 ( .A0(n41), .A1(n2600), .Z(n699));
Q_MX02 U1593 ( .S(n39), .A0(n2697), .A1(n700), .Z(gcm_cmd_in[54]));
Q_AN02 U1594 ( .A0(n41), .A1(n2601), .Z(n700));
Q_MX02 U1595 ( .S(n39), .A0(n2698), .A1(n701), .Z(gcm_cmd_in[53]));
Q_AN02 U1596 ( .A0(n41), .A1(n2602), .Z(n701));
Q_MX02 U1597 ( .S(n39), .A0(n2699), .A1(n702), .Z(gcm_cmd_in[52]));
Q_AN02 U1598 ( .A0(n41), .A1(n2603), .Z(n702));
Q_MX02 U1599 ( .S(n39), .A0(n2700), .A1(n703), .Z(gcm_cmd_in[51]));
Q_AN02 U1600 ( .A0(n41), .A1(n2604), .Z(n703));
Q_MX02 U1601 ( .S(n39), .A0(n2701), .A1(n704), .Z(gcm_cmd_in[50]));
Q_AN02 U1602 ( .A0(n41), .A1(n2605), .Z(n704));
Q_MX02 U1603 ( .S(n39), .A0(n2702), .A1(n705), .Z(gcm_cmd_in[49]));
Q_AN02 U1604 ( .A0(n41), .A1(n2606), .Z(n705));
Q_MX02 U1605 ( .S(n39), .A0(n2703), .A1(n706), .Z(gcm_cmd_in[48]));
Q_AN02 U1606 ( .A0(n41), .A1(n2607), .Z(n706));
Q_MX02 U1607 ( .S(n39), .A0(n2704), .A1(n707), .Z(gcm_cmd_in[47]));
Q_AN02 U1608 ( .A0(n41), .A1(n2608), .Z(n707));
Q_MX02 U1609 ( .S(n39), .A0(n2705), .A1(n708), .Z(gcm_cmd_in[46]));
Q_AN02 U1610 ( .A0(n41), .A1(n2609), .Z(n708));
Q_MX02 U1611 ( .S(n39), .A0(n2706), .A1(n709), .Z(gcm_cmd_in[45]));
Q_AN02 U1612 ( .A0(n41), .A1(n2610), .Z(n709));
Q_MX02 U1613 ( .S(n39), .A0(n2707), .A1(n710), .Z(gcm_cmd_in[44]));
Q_AN02 U1614 ( .A0(n41), .A1(n2611), .Z(n710));
Q_MX02 U1615 ( .S(n39), .A0(n2708), .A1(n711), .Z(gcm_cmd_in[43]));
Q_AN02 U1616 ( .A0(n41), .A1(n2612), .Z(n711));
Q_MX02 U1617 ( .S(n39), .A0(n2709), .A1(n712), .Z(gcm_cmd_in[42]));
Q_AN02 U1618 ( .A0(n41), .A1(n2613), .Z(n712));
Q_MX02 U1619 ( .S(n39), .A0(n2710), .A1(n713), .Z(gcm_cmd_in[41]));
Q_AN02 U1620 ( .A0(n41), .A1(n2614), .Z(n713));
Q_MX02 U1621 ( .S(n39), .A0(n2711), .A1(n714), .Z(gcm_cmd_in[40]));
Q_AN02 U1622 ( .A0(n41), .A1(n2615), .Z(n714));
Q_MX02 U1623 ( .S(n39), .A0(n2712), .A1(n715), .Z(gcm_cmd_in[39]));
Q_AN02 U1624 ( .A0(n41), .A1(n2616), .Z(n715));
Q_MX02 U1625 ( .S(n39), .A0(n2713), .A1(n716), .Z(gcm_cmd_in[38]));
Q_AN02 U1626 ( .A0(n41), .A1(n2617), .Z(n716));
Q_MX02 U1627 ( .S(n39), .A0(n2714), .A1(n717), .Z(gcm_cmd_in[37]));
Q_AN02 U1628 ( .A0(n41), .A1(n2618), .Z(n717));
Q_MX02 U1629 ( .S(n39), .A0(n2715), .A1(n718), .Z(gcm_cmd_in[36]));
Q_AN02 U1630 ( .A0(n41), .A1(n2619), .Z(n718));
Q_MX02 U1631 ( .S(n39), .A0(n2716), .A1(n719), .Z(gcm_cmd_in[35]));
Q_AN02 U1632 ( .A0(n41), .A1(n2620), .Z(n719));
Q_MX02 U1633 ( .S(n39), .A0(n2621), .A1(n720), .Z(gcm_cmd_in[34]));
Q_AN02 U1634 ( .A0(n41), .A1(n2525), .Z(n720));
Q_MX02 U1635 ( .S(n39), .A0(n2622), .A1(n721), .Z(gcm_cmd_in[33]));
Q_AN02 U1636 ( .A0(n41), .A1(n2526), .Z(n721));
Q_MX02 U1637 ( .S(n39), .A0(n2623), .A1(n722), .Z(gcm_cmd_in[32]));
Q_AN02 U1638 ( .A0(n41), .A1(n2527), .Z(n722));
Q_MX02 U1639 ( .S(n39), .A0(n2624), .A1(n723), .Z(gcm_cmd_in[31]));
Q_AN02 U1640 ( .A0(n41), .A1(n2528), .Z(n723));
Q_MX02 U1641 ( .S(n39), .A0(n2625), .A1(n724), .Z(gcm_cmd_in[30]));
Q_AN02 U1642 ( .A0(n41), .A1(n2529), .Z(n724));
Q_MX02 U1643 ( .S(n39), .A0(n2626), .A1(n725), .Z(gcm_cmd_in[29]));
Q_AN02 U1644 ( .A0(n41), .A1(n2530), .Z(n725));
Q_MX02 U1645 ( .S(n39), .A0(n2627), .A1(n726), .Z(gcm_cmd_in[28]));
Q_AN02 U1646 ( .A0(n41), .A1(n2531), .Z(n726));
Q_MX02 U1647 ( .S(n39), .A0(n2628), .A1(n727), .Z(gcm_cmd_in[27]));
Q_AN02 U1648 ( .A0(n41), .A1(n2532), .Z(n727));
Q_MX02 U1649 ( .S(n39), .A0(n2629), .A1(n728), .Z(gcm_cmd_in[26]));
Q_AN02 U1650 ( .A0(n41), .A1(n2533), .Z(n728));
Q_MX02 U1651 ( .S(n39), .A0(n2630), .A1(n729), .Z(gcm_cmd_in[25]));
Q_AN02 U1652 ( .A0(n41), .A1(n2534), .Z(n729));
Q_MX02 U1653 ( .S(n39), .A0(n2631), .A1(n730), .Z(gcm_cmd_in[24]));
Q_AN02 U1654 ( .A0(n41), .A1(n2535), .Z(n730));
Q_MX02 U1655 ( .S(n39), .A0(n2632), .A1(n731), .Z(gcm_cmd_in[23]));
Q_AN02 U1656 ( .A0(n41), .A1(n2536), .Z(n731));
Q_MX02 U1657 ( .S(n39), .A0(n2633), .A1(n732), .Z(gcm_cmd_in[22]));
Q_AN02 U1658 ( .A0(n41), .A1(n2537), .Z(n732));
Q_MX02 U1659 ( .S(n39), .A0(n2634), .A1(n733), .Z(gcm_cmd_in[21]));
Q_AN02 U1660 ( .A0(n41), .A1(n2538), .Z(n733));
Q_MX02 U1661 ( .S(n39), .A0(n2635), .A1(n734), .Z(gcm_cmd_in[20]));
Q_AN02 U1662 ( .A0(n41), .A1(n2539), .Z(n734));
Q_MX02 U1663 ( .S(n39), .A0(n2636), .A1(n735), .Z(gcm_cmd_in[19]));
Q_AN02 U1664 ( .A0(n41), .A1(n2540), .Z(n735));
Q_MX02 U1665 ( .S(n39), .A0(n2637), .A1(n736), .Z(gcm_cmd_in[18]));
Q_AN02 U1666 ( .A0(n41), .A1(n2541), .Z(n736));
Q_MX02 U1667 ( .S(n39), .A0(n2638), .A1(n737), .Z(gcm_cmd_in[17]));
Q_AN02 U1668 ( .A0(n41), .A1(n2542), .Z(n737));
Q_MX02 U1669 ( .S(n39), .A0(n2639), .A1(n738), .Z(gcm_cmd_in[16]));
Q_AN02 U1670 ( .A0(n41), .A1(n2543), .Z(n738));
Q_MX02 U1671 ( .S(n39), .A0(n2640), .A1(n739), .Z(gcm_cmd_in[15]));
Q_AN02 U1672 ( .A0(n41), .A1(n2544), .Z(n739));
Q_MX02 U1673 ( .S(n39), .A0(n2641), .A1(n740), .Z(gcm_cmd_in[14]));
Q_AN02 U1674 ( .A0(n41), .A1(n2545), .Z(n740));
Q_MX02 U1675 ( .S(n39), .A0(n2642), .A1(n741), .Z(gcm_cmd_in[13]));
Q_AN02 U1676 ( .A0(n41), .A1(n2546), .Z(n741));
Q_MX02 U1677 ( .S(n39), .A0(n2643), .A1(n742), .Z(gcm_cmd_in[12]));
Q_AN02 U1678 ( .A0(n41), .A1(n2547), .Z(n742));
Q_MX02 U1679 ( .S(n39), .A0(n2644), .A1(n743), .Z(gcm_cmd_in[11]));
Q_AN02 U1680 ( .A0(n41), .A1(n2548), .Z(n743));
Q_MX02 U1681 ( .S(n39), .A0(n2645), .A1(n744), .Z(gcm_cmd_in[10]));
Q_AN02 U1682 ( .A0(n41), .A1(n2549), .Z(n744));
Q_MX02 U1683 ( .S(n39), .A0(n2646), .A1(n745), .Z(gcm_cmd_in[9]));
Q_AN02 U1684 ( .A0(n41), .A1(n2550), .Z(n745));
Q_MX02 U1685 ( .S(n39), .A0(n2647), .A1(n746), .Z(gcm_cmd_in[8]));
Q_AN02 U1686 ( .A0(n41), .A1(n2551), .Z(n746));
Q_MX02 U1687 ( .S(n39), .A0(n2648), .A1(n747), .Z(gcm_cmd_in[7]));
Q_AN02 U1688 ( .A0(n41), .A1(n2552), .Z(n747));
Q_MX02 U1689 ( .S(n39), .A0(n2649), .A1(n748), .Z(gcm_cmd_in[6]));
Q_AN02 U1690 ( .A0(n41), .A1(n2553), .Z(n748));
Q_MX02 U1691 ( .S(n39), .A0(n2650), .A1(n749), .Z(gcm_cmd_in[5]));
Q_AN02 U1692 ( .A0(n41), .A1(n2554), .Z(n749));
Q_MX02 U1693 ( .S(n39), .A0(n2651), .A1(n750), .Z(gcm_cmd_in[4]));
Q_AN02 U1694 ( .A0(n41), .A1(n2555), .Z(n750));
Q_MX02 U1695 ( .S(n39), .A0(n2652), .A1(n751), .Z(gcm_cmd_in[3]));
Q_AN02 U1696 ( .A0(n41), .A1(n2556), .Z(n751));
Q_MX02 U1697 ( .S(n39), .A0(gcm_dek_cmd_in[2]), .A1(n752), .Z(gcm_cmd_in[2]));
Q_AN02 U1698 ( .A0(n41), .A1(gcm_dak_cmd_in[2]), .Z(n752));
Q_MX02 U1699 ( .S(n39), .A0(gcm_dek_cmd_in[1]), .A1(n753), .Z(gcm_cmd_in[1]));
Q_AN02 U1700 ( .A0(n41), .A1(gcm_dak_cmd_in[1]), .Z(n753));
Q_MX02 U1701 ( .S(n39), .A0(gcm_dek_cmd_in[0]), .A1(n754), .Z(gcm_cmd_in[0]));
Q_AN02 U1702 ( .A0(n41), .A1(gcm_dak_cmd_in[0]), .Z(n754));
Q_MX02 U1703 ( .S(n24), .A0(n755), .A1(n2365), .Z(gcm_tag_data_in[95]));
Q_AN02 U1704 ( .A0(n45), .A1(n2461), .Z(n755));
Q_MX02 U1705 ( .S(n24), .A0(n756), .A1(n2366), .Z(gcm_tag_data_in[94]));
Q_AN02 U1706 ( .A0(n45), .A1(n2462), .Z(n756));
Q_MX02 U1707 ( .S(n24), .A0(n757), .A1(n2367), .Z(gcm_tag_data_in[93]));
Q_AN02 U1708 ( .A0(n45), .A1(n2463), .Z(n757));
Q_MX02 U1709 ( .S(n24), .A0(n758), .A1(n2368), .Z(gcm_tag_data_in[92]));
Q_AN02 U1710 ( .A0(n45), .A1(n2464), .Z(n758));
Q_MX02 U1711 ( .S(n24), .A0(n759), .A1(n2369), .Z(gcm_tag_data_in[91]));
Q_AN02 U1712 ( .A0(n45), .A1(n2465), .Z(n759));
Q_MX02 U1713 ( .S(n24), .A0(n760), .A1(n2370), .Z(gcm_tag_data_in[90]));
Q_AN02 U1714 ( .A0(n45), .A1(n2466), .Z(n760));
Q_MX02 U1715 ( .S(n24), .A0(n761), .A1(n2371), .Z(gcm_tag_data_in[89]));
Q_AN02 U1716 ( .A0(n45), .A1(n2467), .Z(n761));
Q_MX02 U1717 ( .S(n24), .A0(n762), .A1(n2372), .Z(gcm_tag_data_in[88]));
Q_AN02 U1718 ( .A0(n45), .A1(n2468), .Z(n762));
Q_MX02 U1719 ( .S(n24), .A0(n763), .A1(n2373), .Z(gcm_tag_data_in[87]));
Q_AN02 U1720 ( .A0(n45), .A1(n2469), .Z(n763));
Q_MX02 U1721 ( .S(n24), .A0(n764), .A1(n2374), .Z(gcm_tag_data_in[86]));
Q_AN02 U1722 ( .A0(n45), .A1(n2470), .Z(n764));
Q_MX02 U1723 ( .S(n24), .A0(n765), .A1(n2375), .Z(gcm_tag_data_in[85]));
Q_AN02 U1724 ( .A0(n45), .A1(n2471), .Z(n765));
Q_MX02 U1725 ( .S(n24), .A0(n766), .A1(n2376), .Z(gcm_tag_data_in[84]));
Q_AN02 U1726 ( .A0(n45), .A1(n2472), .Z(n766));
Q_MX02 U1727 ( .S(n24), .A0(n767), .A1(n2377), .Z(gcm_tag_data_in[83]));
Q_AN02 U1728 ( .A0(n45), .A1(n2473), .Z(n767));
Q_MX02 U1729 ( .S(n24), .A0(n768), .A1(n2378), .Z(gcm_tag_data_in[82]));
Q_AN02 U1730 ( .A0(n45), .A1(n2474), .Z(n768));
Q_MX02 U1731 ( .S(n24), .A0(n769), .A1(n2379), .Z(gcm_tag_data_in[81]));
Q_AN02 U1732 ( .A0(n45), .A1(n2475), .Z(n769));
Q_MX02 U1733 ( .S(n24), .A0(n770), .A1(n2380), .Z(gcm_tag_data_in[80]));
Q_AN02 U1734 ( .A0(n45), .A1(n2476), .Z(n770));
Q_MX02 U1735 ( .S(n24), .A0(n771), .A1(n2381), .Z(gcm_tag_data_in[79]));
Q_AN02 U1736 ( .A0(n45), .A1(n2477), .Z(n771));
Q_MX02 U1737 ( .S(n24), .A0(n772), .A1(n2382), .Z(gcm_tag_data_in[78]));
Q_AN02 U1738 ( .A0(n45), .A1(n2478), .Z(n772));
Q_MX02 U1739 ( .S(n24), .A0(n773), .A1(n2383), .Z(gcm_tag_data_in[77]));
Q_AN02 U1740 ( .A0(n45), .A1(n2479), .Z(n773));
Q_MX02 U1741 ( .S(n24), .A0(n774), .A1(n2384), .Z(gcm_tag_data_in[76]));
Q_AN02 U1742 ( .A0(n45), .A1(n2480), .Z(n774));
Q_MX02 U1743 ( .S(n24), .A0(n775), .A1(n2385), .Z(gcm_tag_data_in[75]));
Q_AN02 U1744 ( .A0(n45), .A1(n2481), .Z(n775));
Q_MX02 U1745 ( .S(n24), .A0(n776), .A1(n2386), .Z(gcm_tag_data_in[74]));
Q_AN02 U1746 ( .A0(n45), .A1(n2482), .Z(n776));
Q_MX02 U1747 ( .S(n24), .A0(n777), .A1(n2387), .Z(gcm_tag_data_in[73]));
Q_AN02 U1748 ( .A0(n45), .A1(n2483), .Z(n777));
Q_MX02 U1749 ( .S(n24), .A0(n778), .A1(n2388), .Z(gcm_tag_data_in[72]));
Q_AN02 U1750 ( .A0(n45), .A1(n2484), .Z(n778));
Q_MX02 U1751 ( .S(n24), .A0(n779), .A1(n2389), .Z(gcm_tag_data_in[71]));
Q_AN02 U1752 ( .A0(n45), .A1(n2485), .Z(n779));
Q_MX02 U1753 ( .S(n24), .A0(n780), .A1(n2390), .Z(gcm_tag_data_in[70]));
Q_AN02 U1754 ( .A0(n45), .A1(n2486), .Z(n780));
Q_MX02 U1755 ( .S(n24), .A0(n781), .A1(n2391), .Z(gcm_tag_data_in[69]));
Q_AN02 U1756 ( .A0(n45), .A1(n2487), .Z(n781));
Q_MX02 U1757 ( .S(n24), .A0(n782), .A1(n2392), .Z(gcm_tag_data_in[68]));
Q_AN02 U1758 ( .A0(n45), .A1(n2488), .Z(n782));
Q_MX02 U1759 ( .S(n24), .A0(n783), .A1(n2393), .Z(gcm_tag_data_in[67]));
Q_AN02 U1760 ( .A0(n45), .A1(n2489), .Z(n783));
Q_MX02 U1761 ( .S(n24), .A0(n784), .A1(n2394), .Z(gcm_tag_data_in[66]));
Q_AN02 U1762 ( .A0(n45), .A1(n2490), .Z(n784));
Q_MX02 U1763 ( .S(n24), .A0(n785), .A1(n2395), .Z(gcm_tag_data_in[65]));
Q_AN02 U1764 ( .A0(n45), .A1(n2491), .Z(n785));
Q_MX02 U1765 ( .S(n24), .A0(n786), .A1(n2396), .Z(gcm_tag_data_in[64]));
Q_AN02 U1766 ( .A0(n45), .A1(n2492), .Z(n786));
Q_MX02 U1767 ( .S(n24), .A0(n787), .A1(n2397), .Z(gcm_tag_data_in[63]));
Q_AN02 U1768 ( .A0(n45), .A1(n2493), .Z(n787));
Q_MX02 U1769 ( .S(n24), .A0(n788), .A1(n2398), .Z(gcm_tag_data_in[62]));
Q_AN02 U1770 ( .A0(n45), .A1(n2494), .Z(n788));
Q_MX02 U1771 ( .S(n24), .A0(n789), .A1(n2399), .Z(gcm_tag_data_in[61]));
Q_AN02 U1772 ( .A0(n45), .A1(n2495), .Z(n789));
Q_MX02 U1773 ( .S(n24), .A0(n790), .A1(n2400), .Z(gcm_tag_data_in[60]));
Q_AN02 U1774 ( .A0(n45), .A1(n2496), .Z(n790));
Q_MX02 U1775 ( .S(n24), .A0(n791), .A1(n2401), .Z(gcm_tag_data_in[59]));
Q_AN02 U1776 ( .A0(n45), .A1(n2497), .Z(n791));
Q_MX02 U1777 ( .S(n24), .A0(n792), .A1(n2402), .Z(gcm_tag_data_in[58]));
Q_AN02 U1778 ( .A0(n45), .A1(n2498), .Z(n792));
Q_MX02 U1779 ( .S(n24), .A0(n793), .A1(n2403), .Z(gcm_tag_data_in[57]));
Q_AN02 U1780 ( .A0(n45), .A1(n2499), .Z(n793));
Q_MX02 U1781 ( .S(n24), .A0(n794), .A1(n2404), .Z(gcm_tag_data_in[56]));
Q_AN02 U1782 ( .A0(n45), .A1(n2500), .Z(n794));
Q_MX02 U1783 ( .S(n24), .A0(n795), .A1(n2405), .Z(gcm_tag_data_in[55]));
Q_AN02 U1784 ( .A0(n45), .A1(n2501), .Z(n795));
Q_MX02 U1785 ( .S(n24), .A0(n796), .A1(n2406), .Z(gcm_tag_data_in[54]));
Q_AN02 U1786 ( .A0(n45), .A1(n2502), .Z(n796));
Q_MX02 U1787 ( .S(n24), .A0(n797), .A1(n2407), .Z(gcm_tag_data_in[53]));
Q_AN02 U1788 ( .A0(n45), .A1(n2503), .Z(n797));
Q_MX02 U1789 ( .S(n24), .A0(n798), .A1(n2408), .Z(gcm_tag_data_in[52]));
Q_AN02 U1790 ( .A0(n45), .A1(n2504), .Z(n798));
Q_MX02 U1791 ( .S(n24), .A0(n799), .A1(n2409), .Z(gcm_tag_data_in[51]));
Q_AN02 U1792 ( .A0(n45), .A1(n2505), .Z(n799));
Q_MX02 U1793 ( .S(n24), .A0(n800), .A1(n2410), .Z(gcm_tag_data_in[50]));
Q_AN02 U1794 ( .A0(n45), .A1(n2506), .Z(n800));
Q_MX02 U1795 ( .S(n24), .A0(n801), .A1(n2411), .Z(gcm_tag_data_in[49]));
Q_AN02 U1796 ( .A0(n45), .A1(n2507), .Z(n801));
Q_MX02 U1797 ( .S(n24), .A0(n802), .A1(n2412), .Z(gcm_tag_data_in[48]));
Q_AN02 U1798 ( .A0(n45), .A1(n2508), .Z(n802));
Q_MX02 U1799 ( .S(n24), .A0(n803), .A1(n2413), .Z(gcm_tag_data_in[47]));
Q_AN02 U1800 ( .A0(n45), .A1(n2509), .Z(n803));
Q_MX02 U1801 ( .S(n24), .A0(n804), .A1(n2414), .Z(gcm_tag_data_in[46]));
Q_AN02 U1802 ( .A0(n45), .A1(n2510), .Z(n804));
Q_MX02 U1803 ( .S(n24), .A0(n805), .A1(n2415), .Z(gcm_tag_data_in[45]));
Q_AN02 U1804 ( .A0(n45), .A1(n2511), .Z(n805));
Q_MX02 U1805 ( .S(n24), .A0(n806), .A1(n2416), .Z(gcm_tag_data_in[44]));
Q_AN02 U1806 ( .A0(n45), .A1(n2512), .Z(n806));
Q_MX02 U1807 ( .S(n24), .A0(n807), .A1(n2417), .Z(gcm_tag_data_in[43]));
Q_AN02 U1808 ( .A0(n45), .A1(n2513), .Z(n807));
Q_MX02 U1809 ( .S(n24), .A0(n808), .A1(n2418), .Z(gcm_tag_data_in[42]));
Q_AN02 U1810 ( .A0(n45), .A1(n2514), .Z(n808));
Q_MX02 U1811 ( .S(n24), .A0(n809), .A1(n2419), .Z(gcm_tag_data_in[41]));
Q_AN02 U1812 ( .A0(n45), .A1(n2515), .Z(n809));
Q_MX02 U1813 ( .S(n24), .A0(n810), .A1(n2420), .Z(gcm_tag_data_in[40]));
Q_AN02 U1814 ( .A0(n45), .A1(n2516), .Z(n810));
Q_MX02 U1815 ( .S(n24), .A0(n811), .A1(n2421), .Z(gcm_tag_data_in[39]));
Q_AN02 U1816 ( .A0(n45), .A1(n2517), .Z(n811));
Q_MX02 U1817 ( .S(n24), .A0(n812), .A1(n2422), .Z(gcm_tag_data_in[38]));
Q_AN02 U1818 ( .A0(n45), .A1(n2518), .Z(n812));
Q_MX02 U1819 ( .S(n24), .A0(n813), .A1(n2423), .Z(gcm_tag_data_in[37]));
Q_AN02 U1820 ( .A0(n45), .A1(n2519), .Z(n813));
Q_MX02 U1821 ( .S(n24), .A0(n814), .A1(n2424), .Z(gcm_tag_data_in[36]));
Q_AN02 U1822 ( .A0(n45), .A1(n2520), .Z(n814));
Q_MX02 U1823 ( .S(n24), .A0(n815), .A1(n2425), .Z(gcm_tag_data_in[35]));
Q_AN02 U1824 ( .A0(n45), .A1(n2521), .Z(n815));
Q_MX02 U1825 ( .S(n24), .A0(n816), .A1(n2426), .Z(gcm_tag_data_in[34]));
Q_AN02 U1826 ( .A0(n45), .A1(n2522), .Z(n816));
Q_MX02 U1827 ( .S(n24), .A0(n817), .A1(n2427), .Z(gcm_tag_data_in[33]));
Q_AN02 U1828 ( .A0(n45), .A1(n2523), .Z(n817));
Q_MX02 U1829 ( .S(n24), .A0(n818), .A1(n2428), .Z(gcm_tag_data_in[32]));
Q_AN02 U1830 ( .A0(n45), .A1(n2524), .Z(n818));
Q_MX02 U1831 ( .S(n24), .A0(n819), .A1(n2333), .Z(gcm_tag_data_in[31]));
Q_AN02 U1832 ( .A0(n45), .A1(n2429), .Z(n819));
Q_MX02 U1833 ( .S(n24), .A0(n820), .A1(n2334), .Z(gcm_tag_data_in[30]));
Q_AN02 U1834 ( .A0(n45), .A1(n2430), .Z(n820));
Q_MX02 U1835 ( .S(n24), .A0(n821), .A1(n2335), .Z(gcm_tag_data_in[29]));
Q_AN02 U1836 ( .A0(n45), .A1(n2431), .Z(n821));
Q_MX02 U1837 ( .S(n24), .A0(n822), .A1(n2336), .Z(gcm_tag_data_in[28]));
Q_AN02 U1838 ( .A0(n45), .A1(n2432), .Z(n822));
Q_MX02 U1839 ( .S(n24), .A0(n823), .A1(n2337), .Z(gcm_tag_data_in[27]));
Q_AN02 U1840 ( .A0(n45), .A1(n2433), .Z(n823));
Q_MX02 U1841 ( .S(n24), .A0(n824), .A1(n2338), .Z(gcm_tag_data_in[26]));
Q_AN02 U1842 ( .A0(n45), .A1(n2434), .Z(n824));
Q_MX02 U1843 ( .S(n24), .A0(n825), .A1(n2339), .Z(gcm_tag_data_in[25]));
Q_AN02 U1844 ( .A0(n45), .A1(n2435), .Z(n825));
Q_MX02 U1845 ( .S(n24), .A0(n826), .A1(n2340), .Z(gcm_tag_data_in[24]));
Q_AN02 U1846 ( .A0(n45), .A1(n2436), .Z(n826));
Q_MX02 U1847 ( .S(n24), .A0(n827), .A1(n2341), .Z(gcm_tag_data_in[23]));
Q_AN02 U1848 ( .A0(n45), .A1(n2437), .Z(n827));
Q_MX02 U1849 ( .S(n24), .A0(n828), .A1(n2342), .Z(gcm_tag_data_in[22]));
Q_AN02 U1850 ( .A0(n45), .A1(n2438), .Z(n828));
Q_MX02 U1851 ( .S(n24), .A0(n829), .A1(n2343), .Z(gcm_tag_data_in[21]));
Q_AN02 U1852 ( .A0(n45), .A1(n2439), .Z(n829));
Q_MX02 U1853 ( .S(n24), .A0(n830), .A1(n2344), .Z(gcm_tag_data_in[20]));
Q_AN02 U1854 ( .A0(n45), .A1(n2440), .Z(n830));
Q_MX02 U1855 ( .S(n24), .A0(n831), .A1(n2345), .Z(gcm_tag_data_in[19]));
Q_AN02 U1856 ( .A0(n45), .A1(n2441), .Z(n831));
Q_MX02 U1857 ( .S(n24), .A0(n832), .A1(n2346), .Z(gcm_tag_data_in[18]));
Q_AN02 U1858 ( .A0(n45), .A1(n2442), .Z(n832));
Q_MX02 U1859 ( .S(n24), .A0(n833), .A1(n2347), .Z(gcm_tag_data_in[17]));
Q_AN02 U1860 ( .A0(n45), .A1(n2443), .Z(n833));
Q_MX02 U1861 ( .S(n24), .A0(n834), .A1(n2348), .Z(gcm_tag_data_in[16]));
Q_AN02 U1862 ( .A0(n45), .A1(n2444), .Z(n834));
Q_MX02 U1863 ( .S(n24), .A0(n835), .A1(n2349), .Z(gcm_tag_data_in[15]));
Q_AN02 U1864 ( .A0(n45), .A1(n2445), .Z(n835));
Q_MX02 U1865 ( .S(n24), .A0(n836), .A1(n2350), .Z(gcm_tag_data_in[14]));
Q_AN02 U1866 ( .A0(n45), .A1(n2446), .Z(n836));
Q_MX02 U1867 ( .S(n24), .A0(n837), .A1(n2351), .Z(gcm_tag_data_in[13]));
Q_AN02 U1868 ( .A0(n45), .A1(n2447), .Z(n837));
Q_MX02 U1869 ( .S(n24), .A0(n838), .A1(n2352), .Z(gcm_tag_data_in[12]));
Q_AN02 U1870 ( .A0(n45), .A1(n2448), .Z(n838));
Q_MX02 U1871 ( .S(n24), .A0(n839), .A1(n2353), .Z(gcm_tag_data_in[11]));
Q_AN02 U1872 ( .A0(n45), .A1(n2449), .Z(n839));
Q_MX02 U1873 ( .S(n24), .A0(n840), .A1(n2354), .Z(gcm_tag_data_in[10]));
Q_AN02 U1874 ( .A0(n45), .A1(n2450), .Z(n840));
Q_MX02 U1875 ( .S(n24), .A0(n841), .A1(n2355), .Z(gcm_tag_data_in[9]));
Q_AN02 U1876 ( .A0(n45), .A1(n2451), .Z(n841));
Q_MX02 U1877 ( .S(n24), .A0(n842), .A1(n2356), .Z(gcm_tag_data_in[8]));
Q_AN02 U1878 ( .A0(n45), .A1(n2452), .Z(n842));
Q_MX02 U1879 ( .S(n24), .A0(n843), .A1(n2357), .Z(gcm_tag_data_in[7]));
Q_AN02 U1880 ( .A0(n45), .A1(n2453), .Z(n843));
Q_MX02 U1881 ( .S(n24), .A0(n844), .A1(n2358), .Z(gcm_tag_data_in[6]));
Q_AN02 U1882 ( .A0(n45), .A1(n2454), .Z(n844));
Q_MX02 U1883 ( .S(n24), .A0(n845), .A1(n2359), .Z(gcm_tag_data_in[5]));
Q_AN02 U1884 ( .A0(n45), .A1(n2455), .Z(n845));
Q_MX02 U1885 ( .S(n24), .A0(n846), .A1(n2360), .Z(gcm_tag_data_in[4]));
Q_AN02 U1886 ( .A0(n45), .A1(n2456), .Z(n846));
Q_MX02 U1887 ( .S(n24), .A0(n847), .A1(n2361), .Z(gcm_tag_data_in[3]));
Q_AN02 U1888 ( .A0(n45), .A1(n2457), .Z(n847));
Q_MX02 U1889 ( .S(n24), .A0(n848), .A1(n2362), .Z(gcm_tag_data_in[2]));
Q_AN02 U1890 ( .A0(n45), .A1(n2458), .Z(n848));
Q_MX02 U1891 ( .S(n24), .A0(n849), .A1(n2363), .Z(gcm_tag_data_in[1]));
Q_AN02 U1892 ( .A0(n45), .A1(n2459), .Z(n849));
Q_MX02 U1893 ( .S(n24), .A0(n850), .A1(n2364), .Z(gcm_tag_data_in[0]));
Q_AN02 U1894 ( .A0(n45), .A1(n2460), .Z(n850));
Q_AN02 U1895 ( .A0(n52), .A1(kme_internal_out[69]), .Z(inspector_upsizer_eof));
Q_AN02 U1896 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[63]), .Z(inspector_upsizer_data[63]));
Q_AN02 U1897 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[62]), .Z(inspector_upsizer_data[62]));
Q_AN02 U1898 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[61]), .Z(inspector_upsizer_data[61]));
Q_AN02 U1899 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[60]), .Z(inspector_upsizer_data[60]));
Q_AN02 U1900 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[59]), .Z(inspector_upsizer_data[59]));
Q_AN02 U1901 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[58]), .Z(inspector_upsizer_data[58]));
Q_AN02 U1902 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[57]), .Z(inspector_upsizer_data[57]));
Q_AN02 U1903 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[56]), .Z(inspector_upsizer_data[56]));
Q_AN02 U1904 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[55]), .Z(inspector_upsizer_data[55]));
Q_AN02 U1905 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[54]), .Z(inspector_upsizer_data[54]));
Q_AN02 U1906 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[53]), .Z(inspector_upsizer_data[53]));
Q_AN02 U1907 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[52]), .Z(inspector_upsizer_data[52]));
Q_AN02 U1908 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[51]), .Z(inspector_upsizer_data[51]));
Q_AN02 U1909 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[50]), .Z(inspector_upsizer_data[50]));
Q_AN02 U1910 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[49]), .Z(inspector_upsizer_data[49]));
Q_AN02 U1911 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[48]), .Z(inspector_upsizer_data[48]));
Q_AN02 U1912 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[47]), .Z(inspector_upsizer_data[47]));
Q_AN02 U1913 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[46]), .Z(inspector_upsizer_data[46]));
Q_AN02 U1914 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[45]), .Z(inspector_upsizer_data[45]));
Q_AN02 U1915 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[44]), .Z(inspector_upsizer_data[44]));
Q_AN02 U1916 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[43]), .Z(inspector_upsizer_data[43]));
Q_AN02 U1917 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[42]), .Z(inspector_upsizer_data[42]));
Q_AN02 U1918 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[41]), .Z(inspector_upsizer_data[41]));
Q_AN02 U1919 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[40]), .Z(inspector_upsizer_data[40]));
Q_AN02 U1920 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[39]), .Z(inspector_upsizer_data[39]));
Q_AN02 U1921 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[38]), .Z(inspector_upsizer_data[38]));
Q_AN02 U1922 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[37]), .Z(inspector_upsizer_data[37]));
Q_AN02 U1923 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[36]), .Z(inspector_upsizer_data[36]));
Q_AN02 U1924 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[35]), .Z(inspector_upsizer_data[35]));
Q_AN02 U1925 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[34]), .Z(inspector_upsizer_data[34]));
Q_AN02 U1926 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[33]), .Z(inspector_upsizer_data[33]));
Q_AN02 U1927 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[32]), .Z(inspector_upsizer_data[32]));
Q_AN02 U1928 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[31]), .Z(inspector_upsizer_data[31]));
Q_AN02 U1929 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[30]), .Z(inspector_upsizer_data[30]));
Q_AN02 U1930 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[29]), .Z(inspector_upsizer_data[29]));
Q_AN02 U1931 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[28]), .Z(inspector_upsizer_data[28]));
Q_AN02 U1932 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[27]), .Z(inspector_upsizer_data[27]));
Q_AN02 U1933 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[26]), .Z(inspector_upsizer_data[26]));
Q_AN02 U1934 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[25]), .Z(inspector_upsizer_data[25]));
Q_AN02 U1935 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[24]), .Z(inspector_upsizer_data[24]));
Q_AN02 U1936 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[23]), .Z(inspector_upsizer_data[23]));
Q_AN02 U1937 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[22]), .Z(inspector_upsizer_data[22]));
Q_AN02 U1938 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[21]), .Z(inspector_upsizer_data[21]));
Q_AN02 U1939 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[20]), .Z(inspector_upsizer_data[20]));
Q_AN02 U1940 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[19]), .Z(inspector_upsizer_data[19]));
Q_AN02 U1941 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[18]), .Z(inspector_upsizer_data[18]));
Q_AN02 U1942 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[17]), .Z(inspector_upsizer_data[17]));
Q_AN02 U1943 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[16]), .Z(inspector_upsizer_data[16]));
Q_AN02 U1944 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[15]), .Z(inspector_upsizer_data[15]));
Q_AN02 U1945 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[14]), .Z(inspector_upsizer_data[14]));
Q_AN02 U1946 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[13]), .Z(inspector_upsizer_data[13]));
Q_AN02 U1947 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[12]), .Z(inspector_upsizer_data[12]));
Q_AN02 U1948 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[11]), .Z(inspector_upsizer_data[11]));
Q_AN02 U1949 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[10]), .Z(inspector_upsizer_data[10]));
Q_AN02 U1950 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[9]), .Z(inspector_upsizer_data[9]));
Q_AN02 U1951 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[8]), .Z(inspector_upsizer_data[8]));
Q_AN02 U1952 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[7]), .Z(inspector_upsizer_data[7]));
Q_AN02 U1953 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[6]), .Z(inspector_upsizer_data[6]));
Q_AN02 U1954 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[5]), .Z(inspector_upsizer_data[5]));
Q_AN02 U1955 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[4]), .Z(inspector_upsizer_data[4]));
Q_AN02 U1956 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[3]), .Z(inspector_upsizer_data[3]));
Q_AN02 U1957 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[2]), .Z(inspector_upsizer_data[2]));
Q_AN02 U1958 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[1]), .Z(inspector_upsizer_data[1]));
Q_AN02 U1959 ( .A0(inspector_upsizer_valid), .A1(kme_internal_out[0]), .Z(inspector_upsizer_data[0]));
Q_AN02 U1960 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[262]), .Z(kdfstream_cmd_in[262]));
Q_MX02 U1961 ( .S(n56), .A0(n852), .A1(n851), .Z(kdfstream_cmd_in[261]));
Q_AN02 U1962 ( .A0(n25), .A1(skip_dak_kdf), .Z(n851));
Q_MX02 U1963 ( .S(n59), .A0(stream_cmd_in[261]), .A1(skip_dek_kdf), .Z(n852));
Q_AN02 U1964 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[260]), .Z(kdfstream_cmd_in[260]));
Q_AN02 U1965 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[259]), .Z(kdfstream_cmd_in[259]));
Q_AN02 U1966 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[258]), .Z(kdfstream_cmd_in[258]));
Q_AN02 U1967 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[257]), .Z(kdfstream_cmd_in[257]));
Q_AN02 U1968 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[256]), .Z(kdfstream_cmd_in[256]));
Q_AN02 U1969 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[255]), .Z(kdfstream_cmd_in[255]));
Q_AN02 U1970 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[254]), .Z(kdfstream_cmd_in[254]));
Q_AN02 U1971 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[253]), .Z(kdfstream_cmd_in[253]));
Q_AN02 U1972 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[252]), .Z(kdfstream_cmd_in[252]));
Q_AN02 U1973 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[251]), .Z(kdfstream_cmd_in[251]));
Q_AN02 U1974 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[250]), .Z(kdfstream_cmd_in[250]));
Q_AN02 U1975 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[249]), .Z(kdfstream_cmd_in[249]));
Q_AN02 U1976 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[248]), .Z(kdfstream_cmd_in[248]));
Q_AN02 U1977 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[247]), .Z(kdfstream_cmd_in[247]));
Q_AN02 U1978 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[246]), .Z(kdfstream_cmd_in[246]));
Q_AN02 U1979 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[245]), .Z(kdfstream_cmd_in[245]));
Q_AN02 U1980 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[244]), .Z(kdfstream_cmd_in[244]));
Q_AN02 U1981 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[243]), .Z(kdfstream_cmd_in[243]));
Q_AN02 U1982 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[242]), .Z(kdfstream_cmd_in[242]));
Q_AN02 U1983 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[241]), .Z(kdfstream_cmd_in[241]));
Q_AN02 U1984 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[240]), .Z(kdfstream_cmd_in[240]));
Q_AN02 U1985 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[239]), .Z(kdfstream_cmd_in[239]));
Q_AN02 U1986 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[238]), .Z(kdfstream_cmd_in[238]));
Q_AN02 U1987 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[237]), .Z(kdfstream_cmd_in[237]));
Q_AN02 U1988 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[236]), .Z(kdfstream_cmd_in[236]));
Q_AN02 U1989 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[235]), .Z(kdfstream_cmd_in[235]));
Q_AN02 U1990 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[234]), .Z(kdfstream_cmd_in[234]));
Q_AN02 U1991 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[233]), .Z(kdfstream_cmd_in[233]));
Q_AN02 U1992 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[232]), .Z(kdfstream_cmd_in[232]));
Q_AN02 U1993 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[231]), .Z(kdfstream_cmd_in[231]));
Q_AN02 U1994 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[230]), .Z(kdfstream_cmd_in[230]));
Q_AN02 U1995 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[229]), .Z(kdfstream_cmd_in[229]));
Q_AN02 U1996 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[228]), .Z(kdfstream_cmd_in[228]));
Q_AN02 U1997 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[227]), .Z(kdfstream_cmd_in[227]));
Q_AN02 U1998 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[226]), .Z(kdfstream_cmd_in[226]));
Q_AN02 U1999 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[225]), .Z(kdfstream_cmd_in[225]));
Q_AN02 U2000 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[224]), .Z(kdfstream_cmd_in[224]));
Q_AN02 U2001 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[223]), .Z(kdfstream_cmd_in[223]));
Q_AN02 U2002 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[222]), .Z(kdfstream_cmd_in[222]));
Q_AN02 U2003 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[221]), .Z(kdfstream_cmd_in[221]));
Q_AN02 U2004 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[220]), .Z(kdfstream_cmd_in[220]));
Q_AN02 U2005 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[219]), .Z(kdfstream_cmd_in[219]));
Q_AN02 U2006 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[218]), .Z(kdfstream_cmd_in[218]));
Q_AN02 U2007 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[217]), .Z(kdfstream_cmd_in[217]));
Q_AN02 U2008 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[216]), .Z(kdfstream_cmd_in[216]));
Q_AN02 U2009 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[215]), .Z(kdfstream_cmd_in[215]));
Q_AN02 U2010 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[214]), .Z(kdfstream_cmd_in[214]));
Q_AN02 U2011 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[213]), .Z(kdfstream_cmd_in[213]));
Q_AN02 U2012 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[212]), .Z(kdfstream_cmd_in[212]));
Q_AN02 U2013 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[211]), .Z(kdfstream_cmd_in[211]));
Q_AN02 U2014 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[210]), .Z(kdfstream_cmd_in[210]));
Q_AN02 U2015 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[209]), .Z(kdfstream_cmd_in[209]));
Q_AN02 U2016 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[208]), .Z(kdfstream_cmd_in[208]));
Q_AN02 U2017 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[207]), .Z(kdfstream_cmd_in[207]));
Q_AN02 U2018 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[206]), .Z(kdfstream_cmd_in[206]));
Q_AN02 U2019 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[205]), .Z(kdfstream_cmd_in[205]));
Q_AN02 U2020 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[204]), .Z(kdfstream_cmd_in[204]));
Q_AN02 U2021 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[203]), .Z(kdfstream_cmd_in[203]));
Q_AN02 U2022 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[202]), .Z(kdfstream_cmd_in[202]));
Q_AN02 U2023 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[201]), .Z(kdfstream_cmd_in[201]));
Q_AN02 U2024 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[200]), .Z(kdfstream_cmd_in[200]));
Q_AN02 U2025 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[199]), .Z(kdfstream_cmd_in[199]));
Q_AN02 U2026 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[198]), .Z(kdfstream_cmd_in[198]));
Q_AN02 U2027 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[197]), .Z(kdfstream_cmd_in[197]));
Q_AN02 U2028 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[196]), .Z(kdfstream_cmd_in[196]));
Q_AN02 U2029 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[195]), .Z(kdfstream_cmd_in[195]));
Q_AN02 U2030 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[194]), .Z(kdfstream_cmd_in[194]));
Q_AN02 U2031 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[193]), .Z(kdfstream_cmd_in[193]));
Q_AN02 U2032 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[192]), .Z(kdfstream_cmd_in[192]));
Q_AN02 U2033 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[191]), .Z(kdfstream_cmd_in[191]));
Q_AN02 U2034 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[190]), .Z(kdfstream_cmd_in[190]));
Q_AN02 U2035 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[189]), .Z(kdfstream_cmd_in[189]));
Q_AN02 U2036 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[188]), .Z(kdfstream_cmd_in[188]));
Q_AN02 U2037 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[187]), .Z(kdfstream_cmd_in[187]));
Q_AN02 U2038 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[186]), .Z(kdfstream_cmd_in[186]));
Q_AN02 U2039 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[185]), .Z(kdfstream_cmd_in[185]));
Q_AN02 U2040 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[184]), .Z(kdfstream_cmd_in[184]));
Q_AN02 U2041 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[183]), .Z(kdfstream_cmd_in[183]));
Q_AN02 U2042 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[182]), .Z(kdfstream_cmd_in[182]));
Q_AN02 U2043 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[181]), .Z(kdfstream_cmd_in[181]));
Q_AN02 U2044 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[180]), .Z(kdfstream_cmd_in[180]));
Q_AN02 U2045 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[179]), .Z(kdfstream_cmd_in[179]));
Q_AN02 U2046 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[178]), .Z(kdfstream_cmd_in[178]));
Q_AN02 U2047 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[177]), .Z(kdfstream_cmd_in[177]));
Q_AN02 U2048 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[176]), .Z(kdfstream_cmd_in[176]));
Q_AN02 U2049 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[175]), .Z(kdfstream_cmd_in[175]));
Q_AN02 U2050 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[174]), .Z(kdfstream_cmd_in[174]));
Q_AN02 U2051 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[173]), .Z(kdfstream_cmd_in[173]));
Q_AN02 U2052 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[172]), .Z(kdfstream_cmd_in[172]));
Q_AN02 U2053 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[171]), .Z(kdfstream_cmd_in[171]));
Q_AN02 U2054 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[170]), .Z(kdfstream_cmd_in[170]));
Q_AN02 U2055 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[169]), .Z(kdfstream_cmd_in[169]));
Q_AN02 U2056 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[168]), .Z(kdfstream_cmd_in[168]));
Q_AN02 U2057 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[167]), .Z(kdfstream_cmd_in[167]));
Q_AN02 U2058 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[166]), .Z(kdfstream_cmd_in[166]));
Q_AN02 U2059 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[165]), .Z(kdfstream_cmd_in[165]));
Q_AN02 U2060 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[164]), .Z(kdfstream_cmd_in[164]));
Q_AN02 U2061 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[163]), .Z(kdfstream_cmd_in[163]));
Q_AN02 U2062 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[162]), .Z(kdfstream_cmd_in[162]));
Q_AN02 U2063 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[161]), .Z(kdfstream_cmd_in[161]));
Q_AN02 U2064 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[160]), .Z(kdfstream_cmd_in[160]));
Q_AN02 U2065 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[159]), .Z(kdfstream_cmd_in[159]));
Q_AN02 U2066 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[158]), .Z(kdfstream_cmd_in[158]));
Q_AN02 U2067 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[157]), .Z(kdfstream_cmd_in[157]));
Q_AN02 U2068 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[156]), .Z(kdfstream_cmd_in[156]));
Q_AN02 U2069 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[155]), .Z(kdfstream_cmd_in[155]));
Q_AN02 U2070 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[154]), .Z(kdfstream_cmd_in[154]));
Q_AN02 U2071 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[153]), .Z(kdfstream_cmd_in[153]));
Q_AN02 U2072 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[152]), .Z(kdfstream_cmd_in[152]));
Q_AN02 U2073 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[151]), .Z(kdfstream_cmd_in[151]));
Q_AN02 U2074 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[150]), .Z(kdfstream_cmd_in[150]));
Q_AN02 U2075 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[149]), .Z(kdfstream_cmd_in[149]));
Q_AN02 U2076 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[148]), .Z(kdfstream_cmd_in[148]));
Q_AN02 U2077 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[147]), .Z(kdfstream_cmd_in[147]));
Q_AN02 U2078 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[146]), .Z(kdfstream_cmd_in[146]));
Q_AN02 U2079 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[145]), .Z(kdfstream_cmd_in[145]));
Q_AN02 U2080 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[144]), .Z(kdfstream_cmd_in[144]));
Q_AN02 U2081 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[143]), .Z(kdfstream_cmd_in[143]));
Q_AN02 U2082 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[142]), .Z(kdfstream_cmd_in[142]));
Q_AN02 U2083 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[141]), .Z(kdfstream_cmd_in[141]));
Q_AN02 U2084 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[140]), .Z(kdfstream_cmd_in[140]));
Q_AN02 U2085 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[139]), .Z(kdfstream_cmd_in[139]));
Q_AN02 U2086 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[138]), .Z(kdfstream_cmd_in[138]));
Q_AN02 U2087 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[137]), .Z(kdfstream_cmd_in[137]));
Q_AN02 U2088 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[136]), .Z(kdfstream_cmd_in[136]));
Q_AN02 U2089 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[135]), .Z(kdfstream_cmd_in[135]));
Q_AN02 U2090 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[134]), .Z(kdfstream_cmd_in[134]));
Q_AN02 U2091 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[133]), .Z(kdfstream_cmd_in[133]));
Q_AN02 U2092 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[132]), .Z(kdfstream_cmd_in[132]));
Q_AN02 U2093 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[131]), .Z(kdfstream_cmd_in[131]));
Q_AN02 U2094 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[130]), .Z(kdfstream_cmd_in[130]));
Q_AN02 U2095 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[129]), .Z(kdfstream_cmd_in[129]));
Q_AN02 U2096 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[128]), .Z(kdfstream_cmd_in[128]));
Q_AN02 U2097 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[127]), .Z(kdfstream_cmd_in[127]));
Q_AN02 U2098 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[126]), .Z(kdfstream_cmd_in[126]));
Q_AN02 U2099 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[125]), .Z(kdfstream_cmd_in[125]));
Q_AN02 U2100 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[124]), .Z(kdfstream_cmd_in[124]));
Q_AN02 U2101 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[123]), .Z(kdfstream_cmd_in[123]));
Q_AN02 U2102 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[122]), .Z(kdfstream_cmd_in[122]));
Q_AN02 U2103 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[121]), .Z(kdfstream_cmd_in[121]));
Q_AN02 U2104 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[120]), .Z(kdfstream_cmd_in[120]));
Q_AN02 U2105 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[119]), .Z(kdfstream_cmd_in[119]));
Q_AN02 U2106 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[118]), .Z(kdfstream_cmd_in[118]));
Q_AN02 U2107 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[117]), .Z(kdfstream_cmd_in[117]));
Q_AN02 U2108 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[116]), .Z(kdfstream_cmd_in[116]));
Q_AN02 U2109 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[115]), .Z(kdfstream_cmd_in[115]));
Q_AN02 U2110 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[114]), .Z(kdfstream_cmd_in[114]));
Q_AN02 U2111 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[113]), .Z(kdfstream_cmd_in[113]));
Q_AN02 U2112 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[112]), .Z(kdfstream_cmd_in[112]));
Q_AN02 U2113 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[111]), .Z(kdfstream_cmd_in[111]));
Q_AN02 U2114 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[110]), .Z(kdfstream_cmd_in[110]));
Q_AN02 U2115 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[109]), .Z(kdfstream_cmd_in[109]));
Q_AN02 U2116 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[108]), .Z(kdfstream_cmd_in[108]));
Q_AN02 U2117 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[107]), .Z(kdfstream_cmd_in[107]));
Q_AN02 U2118 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[106]), .Z(kdfstream_cmd_in[106]));
Q_AN02 U2119 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[105]), .Z(kdfstream_cmd_in[105]));
Q_AN02 U2120 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[104]), .Z(kdfstream_cmd_in[104]));
Q_AN02 U2121 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[103]), .Z(kdfstream_cmd_in[103]));
Q_AN02 U2122 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[102]), .Z(kdfstream_cmd_in[102]));
Q_AN02 U2123 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[101]), .Z(kdfstream_cmd_in[101]));
Q_AN02 U2124 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[100]), .Z(kdfstream_cmd_in[100]));
Q_AN02 U2125 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[99]), .Z(kdfstream_cmd_in[99]));
Q_AN02 U2126 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[98]), .Z(kdfstream_cmd_in[98]));
Q_AN02 U2127 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[97]), .Z(kdfstream_cmd_in[97]));
Q_AN02 U2128 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[96]), .Z(kdfstream_cmd_in[96]));
Q_AN02 U2129 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[95]), .Z(kdfstream_cmd_in[95]));
Q_AN02 U2130 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[94]), .Z(kdfstream_cmd_in[94]));
Q_AN02 U2131 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[93]), .Z(kdfstream_cmd_in[93]));
Q_AN02 U2132 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[92]), .Z(kdfstream_cmd_in[92]));
Q_AN02 U2133 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[91]), .Z(kdfstream_cmd_in[91]));
Q_AN02 U2134 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[90]), .Z(kdfstream_cmd_in[90]));
Q_AN02 U2135 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[89]), .Z(kdfstream_cmd_in[89]));
Q_AN02 U2136 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[88]), .Z(kdfstream_cmd_in[88]));
Q_AN02 U2137 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[87]), .Z(kdfstream_cmd_in[87]));
Q_AN02 U2138 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[86]), .Z(kdfstream_cmd_in[86]));
Q_AN02 U2139 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[85]), .Z(kdfstream_cmd_in[85]));
Q_AN02 U2140 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[84]), .Z(kdfstream_cmd_in[84]));
Q_AN02 U2141 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[83]), .Z(kdfstream_cmd_in[83]));
Q_AN02 U2142 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[82]), .Z(kdfstream_cmd_in[82]));
Q_AN02 U2143 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[81]), .Z(kdfstream_cmd_in[81]));
Q_AN02 U2144 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[80]), .Z(kdfstream_cmd_in[80]));
Q_AN02 U2145 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[79]), .Z(kdfstream_cmd_in[79]));
Q_AN02 U2146 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[78]), .Z(kdfstream_cmd_in[78]));
Q_AN02 U2147 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[77]), .Z(kdfstream_cmd_in[77]));
Q_AN02 U2148 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[76]), .Z(kdfstream_cmd_in[76]));
Q_AN02 U2149 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[75]), .Z(kdfstream_cmd_in[75]));
Q_AN02 U2150 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[74]), .Z(kdfstream_cmd_in[74]));
Q_AN02 U2151 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[73]), .Z(kdfstream_cmd_in[73]));
Q_AN02 U2152 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[72]), .Z(kdfstream_cmd_in[72]));
Q_AN02 U2153 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[71]), .Z(kdfstream_cmd_in[71]));
Q_AN02 U2154 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[70]), .Z(kdfstream_cmd_in[70]));
Q_AN02 U2155 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[69]), .Z(kdfstream_cmd_in[69]));
Q_AN02 U2156 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[68]), .Z(kdfstream_cmd_in[68]));
Q_AN02 U2157 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[67]), .Z(kdfstream_cmd_in[67]));
Q_AN02 U2158 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[66]), .Z(kdfstream_cmd_in[66]));
Q_AN02 U2159 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[65]), .Z(kdfstream_cmd_in[65]));
Q_AN02 U2160 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[64]), .Z(kdfstream_cmd_in[64]));
Q_AN02 U2161 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[63]), .Z(kdfstream_cmd_in[63]));
Q_AN02 U2162 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[62]), .Z(kdfstream_cmd_in[62]));
Q_AN02 U2163 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[61]), .Z(kdfstream_cmd_in[61]));
Q_AN02 U2164 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[60]), .Z(kdfstream_cmd_in[60]));
Q_AN02 U2165 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[59]), .Z(kdfstream_cmd_in[59]));
Q_AN02 U2166 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[58]), .Z(kdfstream_cmd_in[58]));
Q_AN02 U2167 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[57]), .Z(kdfstream_cmd_in[57]));
Q_AN02 U2168 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[56]), .Z(kdfstream_cmd_in[56]));
Q_AN02 U2169 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[55]), .Z(kdfstream_cmd_in[55]));
Q_AN02 U2170 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[54]), .Z(kdfstream_cmd_in[54]));
Q_AN02 U2171 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[53]), .Z(kdfstream_cmd_in[53]));
Q_AN02 U2172 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[52]), .Z(kdfstream_cmd_in[52]));
Q_AN02 U2173 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[51]), .Z(kdfstream_cmd_in[51]));
Q_AN02 U2174 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[50]), .Z(kdfstream_cmd_in[50]));
Q_AN02 U2175 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[49]), .Z(kdfstream_cmd_in[49]));
Q_AN02 U2176 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[48]), .Z(kdfstream_cmd_in[48]));
Q_AN02 U2177 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[47]), .Z(kdfstream_cmd_in[47]));
Q_AN02 U2178 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[46]), .Z(kdfstream_cmd_in[46]));
Q_AN02 U2179 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[45]), .Z(kdfstream_cmd_in[45]));
Q_AN02 U2180 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[44]), .Z(kdfstream_cmd_in[44]));
Q_AN02 U2181 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[43]), .Z(kdfstream_cmd_in[43]));
Q_AN02 U2182 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[42]), .Z(kdfstream_cmd_in[42]));
Q_AN02 U2183 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[41]), .Z(kdfstream_cmd_in[41]));
Q_AN02 U2184 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[40]), .Z(kdfstream_cmd_in[40]));
Q_AN02 U2185 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[39]), .Z(kdfstream_cmd_in[39]));
Q_AN02 U2186 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[38]), .Z(kdfstream_cmd_in[38]));
Q_AN02 U2187 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[37]), .Z(kdfstream_cmd_in[37]));
Q_AN02 U2188 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[36]), .Z(kdfstream_cmd_in[36]));
Q_AN02 U2189 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[35]), .Z(kdfstream_cmd_in[35]));
Q_AN02 U2190 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[34]), .Z(kdfstream_cmd_in[34]));
Q_AN02 U2191 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[33]), .Z(kdfstream_cmd_in[33]));
Q_AN02 U2192 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[32]), .Z(kdfstream_cmd_in[32]));
Q_AN02 U2193 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[31]), .Z(kdfstream_cmd_in[31]));
Q_AN02 U2194 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[30]), .Z(kdfstream_cmd_in[30]));
Q_AN02 U2195 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[29]), .Z(kdfstream_cmd_in[29]));
Q_AN02 U2196 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[28]), .Z(kdfstream_cmd_in[28]));
Q_AN02 U2197 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[27]), .Z(kdfstream_cmd_in[27]));
Q_AN02 U2198 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[26]), .Z(kdfstream_cmd_in[26]));
Q_AN02 U2199 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[25]), .Z(kdfstream_cmd_in[25]));
Q_AN02 U2200 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[24]), .Z(kdfstream_cmd_in[24]));
Q_AN02 U2201 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[23]), .Z(kdfstream_cmd_in[23]));
Q_AN02 U2202 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[22]), .Z(kdfstream_cmd_in[22]));
Q_AN02 U2203 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[21]), .Z(kdfstream_cmd_in[21]));
Q_AN02 U2204 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[20]), .Z(kdfstream_cmd_in[20]));
Q_AN02 U2205 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[19]), .Z(kdfstream_cmd_in[19]));
Q_AN02 U2206 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[18]), .Z(kdfstream_cmd_in[18]));
Q_AN02 U2207 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[17]), .Z(kdfstream_cmd_in[17]));
Q_AN02 U2208 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[16]), .Z(kdfstream_cmd_in[16]));
Q_AN02 U2209 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[15]), .Z(kdfstream_cmd_in[15]));
Q_AN02 U2210 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[14]), .Z(kdfstream_cmd_in[14]));
Q_AN02 U2211 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[13]), .Z(kdfstream_cmd_in[13]));
Q_AN02 U2212 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[12]), .Z(kdfstream_cmd_in[12]));
Q_AN02 U2213 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[11]), .Z(kdfstream_cmd_in[11]));
Q_AN02 U2214 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[10]), .Z(kdfstream_cmd_in[10]));
Q_AN02 U2215 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[9]), .Z(kdfstream_cmd_in[9]));
Q_AN02 U2216 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[8]), .Z(kdfstream_cmd_in[8]));
Q_AN02 U2217 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[7]), .Z(kdfstream_cmd_in[7]));
Q_AN02 U2218 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[6]), .Z(kdfstream_cmd_in[6]));
Q_AN02 U2219 ( .A0(kdfstream_cmd_in_valid), .A1(stream_cmd_in[5]), .Z(kdfstream_cmd_in[5]));
Q_AN02 U2220 ( .A0(kdfstream_cmd_in_valid), .A1(kme_internal_out[62]), .Z(kdfstream_cmd_in[4]));
Q_AN02 U2221 ( .A0(kdfstream_cmd_in_valid), .A1(kme_internal_out[61]), .Z(kdfstream_cmd_in[3]));
Q_AN02 U2222 ( .A0(kdfstream_cmd_in_valid), .A1(kme_internal_out[60]), .Z(kdfstream_cmd_in[2]));
Q_AN02 U2223 ( .A0(n26), .A1(stream_cmd_in[1]), .Z(kdfstream_cmd_in[1]));
Q_MX02 U2224 ( .S(n56), .A0(stream_cmd_in[0]), .A1(n27), .Z(kdfstream_cmd_in[0]));
Q_AN02 U2225 ( .A0(keyfilter_cmd_in_valid), .A1(kdf_dek_iter), .Z(kdf_cmd_in[3]));
Q_AN02 U2226 ( .A0(keyfilter_cmd_in_valid), .A1(kme_internal_out[16]), .Z(keyfilter_cmd_in[0]));
Q_AN02 U2227 ( .A0(keyfilter_cmd_in_valid), .A1(kme_internal_out[14]), .Z(kdf_cmd_in[1]));
Q_AN02 U2228 ( .A0(keyfilter_cmd_in_valid), .A1(kme_internal_out[31]), .Z(kdf_cmd_in[0]));
Q_AN02 U2229 ( .A0(n28), .A1(kme_internal_out[63]), .Z(tlv_sb_data_in[63]));
Q_AN02 U2230 ( .A0(n28), .A1(kme_internal_out[62]), .Z(tlv_sb_data_in[62]));
Q_AN02 U2231 ( .A0(n28), .A1(kme_internal_out[61]), .Z(tlv_sb_data_in[61]));
Q_AN02 U2232 ( .A0(n28), .A1(kme_internal_out[60]), .Z(tlv_sb_data_in[60]));
Q_AN02 U2233 ( .A0(n28), .A1(kme_internal_out[59]), .Z(tlv_sb_data_in[59]));
Q_AN02 U2234 ( .A0(n28), .A1(kme_internal_out[58]), .Z(tlv_sb_data_in[58]));
Q_AN02 U2235 ( .A0(n28), .A1(kme_internal_out[57]), .Z(tlv_sb_data_in[57]));
Q_AN02 U2236 ( .A0(n28), .A1(kme_internal_out[56]), .Z(tlv_sb_data_in[56]));
Q_MX02 U2237 ( .S(n62), .A0(kme_internal_out[55]), .A1(n853), .Z(tlv_sb_data_in[55]));
Q_AN02 U2238 ( .A0(n29), .A1(int_tlv_word42[55]), .Z(n853));
Q_AN02 U2239 ( .A0(n1), .A1(kme_internal_out[54]), .Z(tlv_sb_data_in[54]));
Q_AN02 U2240 ( .A0(n1), .A1(kme_internal_out[53]), .Z(tlv_sb_data_in[53]));
Q_AN02 U2241 ( .A0(n1), .A1(kme_internal_out[52]), .Z(tlv_sb_data_in[52]));
Q_AN02 U2242 ( .A0(n1), .A1(kme_internal_out[51]), .Z(tlv_sb_data_in[51]));
Q_AN02 U2243 ( .A0(n1), .A1(kme_internal_out[50]), .Z(tlv_sb_data_in[50]));
Q_AN02 U2244 ( .A0(n1), .A1(kme_internal_out[49]), .Z(tlv_sb_data_in[49]));
Q_AN02 U2245 ( .A0(n1), .A1(kme_internal_out[48]), .Z(tlv_sb_data_in[48]));
Q_AN02 U2246 ( .A0(n1), .A1(kme_internal_out[47]), .Z(tlv_sb_data_in[47]));
Q_AN02 U2247 ( .A0(n1), .A1(kme_internal_out[46]), .Z(tlv_sb_data_in[46]));
Q_AN02 U2248 ( .A0(n1), .A1(kme_internal_out[45]), .Z(tlv_sb_data_in[45]));
Q_AN02 U2249 ( .A0(n1), .A1(kme_internal_out[44]), .Z(tlv_sb_data_in[44]));
Q_AN02 U2250 ( .A0(n1), .A1(kme_internal_out[43]), .Z(tlv_sb_data_in[43]));
Q_AN02 U2251 ( .A0(n1), .A1(kme_internal_out[42]), .Z(tlv_sb_data_in[42]));
Q_AN02 U2252 ( .A0(n1), .A1(kme_internal_out[41]), .Z(tlv_sb_data_in[41]));
Q_AN02 U2253 ( .A0(n1), .A1(kme_internal_out[40]), .Z(tlv_sb_data_in[40]));
Q_AN02 U2254 ( .A0(n1), .A1(kme_internal_out[39]), .Z(tlv_sb_data_in[39]));
Q_AN02 U2255 ( .A0(n1), .A1(kme_internal_out[38]), .Z(tlv_sb_data_in[38]));
Q_AN02 U2256 ( .A0(n1), .A1(kme_internal_out[37]), .Z(tlv_sb_data_in[37]));
Q_AN02 U2257 ( .A0(n1), .A1(kme_internal_out[36]), .Z(tlv_sb_data_in[36]));
Q_AN02 U2258 ( .A0(n1), .A1(kme_internal_out[35]), .Z(tlv_sb_data_in[35]));
Q_AN02 U2259 ( .A0(n1), .A1(kme_internal_out[34]), .Z(tlv_sb_data_in[34]));
Q_AN02 U2260 ( .A0(n1), .A1(kme_internal_out[33]), .Z(tlv_sb_data_in[33]));
Q_AN02 U2261 ( .A0(n1), .A1(kme_internal_out[32]), .Z(tlv_sb_data_in[32]));
Q_AN02 U2262 ( .A0(n1), .A1(kme_internal_out[31]), .Z(tlv_sb_data_in[31]));
Q_AN02 U2263 ( .A0(n1), .A1(kme_internal_out[30]), .Z(tlv_sb_data_in[30]));
Q_AN02 U2264 ( .A0(n1), .A1(kme_internal_out[29]), .Z(tlv_sb_data_in[29]));
Q_AN02 U2265 ( .A0(n1), .A1(kme_internal_out[28]), .Z(tlv_sb_data_in[28]));
Q_AN02 U2266 ( .A0(n1), .A1(kme_internal_out[27]), .Z(tlv_sb_data_in[27]));
Q_AN02 U2267 ( .A0(n1), .A1(kme_internal_out[26]), .Z(tlv_sb_data_in[26]));
Q_AN02 U2268 ( .A0(n1), .A1(kme_internal_out[25]), .Z(tlv_sb_data_in[25]));
Q_AN02 U2269 ( .A0(n1), .A1(kme_internal_out[24]), .Z(tlv_sb_data_in[24]));
Q_AN02 U2270 ( .A0(n1), .A1(kme_internal_out[23]), .Z(tlv_sb_data_in[23]));
Q_AN02 U2271 ( .A0(n1), .A1(kme_internal_out[22]), .Z(tlv_sb_data_in[22]));
Q_AN02 U2272 ( .A0(n1), .A1(kme_internal_out[21]), .Z(tlv_sb_data_in[21]));
Q_AN02 U2273 ( .A0(n1), .A1(kme_internal_out[20]), .Z(tlv_sb_data_in[20]));
Q_AN02 U2274 ( .A0(n1), .A1(kme_internal_out[19]), .Z(tlv_sb_data_in[19]));
Q_AN02 U2275 ( .A0(n1), .A1(kme_internal_out[18]), .Z(tlv_sb_data_in[18]));
Q_AN02 U2276 ( .A0(n1), .A1(kme_internal_out[17]), .Z(tlv_sb_data_in[17]));
Q_AN02 U2277 ( .A0(n1), .A1(kme_internal_out[16]), .Z(tlv_sb_data_in[16]));
Q_AN02 U2278 ( .A0(n1), .A1(kme_internal_out[15]), .Z(tlv_sb_data_in[15]));
Q_AN02 U2279 ( .A0(n1), .A1(kme_internal_out[14]), .Z(tlv_sb_data_in[14]));
Q_AN02 U2280 ( .A0(n1), .A1(kme_internal_out[13]), .Z(tlv_sb_data_in[13]));
Q_AN02 U2281 ( .A0(n1), .A1(kme_internal_out[12]), .Z(tlv_sb_data_in[12]));
Q_AN02 U2282 ( .A0(n1), .A1(kme_internal_out[11]), .Z(tlv_sb_data_in[11]));
Q_AN02 U2283 ( .A0(n1), .A1(kme_internal_out[10]), .Z(tlv_sb_data_in[10]));
Q_AN02 U2284 ( .A0(n1), .A1(kme_internal_out[9]), .Z(tlv_sb_data_in[9]));
Q_AN02 U2285 ( .A0(n1), .A1(kme_internal_out[8]), .Z(tlv_sb_data_in[8]));
Q_AN02 U2286 ( .A0(n1), .A1(kme_internal_out[7]), .Z(tlv_sb_data_in[7]));
Q_AN02 U2287 ( .A0(n1), .A1(kme_internal_out[6]), .Z(tlv_sb_data_in[6]));
Q_AN02 U2288 ( .A0(n1), .A1(kme_internal_out[5]), .Z(tlv_sb_data_in[5]));
Q_AN02 U2289 ( .A0(n1), .A1(kme_internal_out[4]), .Z(tlv_sb_data_in[4]));
Q_AN02 U2290 ( .A0(n1), .A1(kme_internal_out[3]), .Z(tlv_sb_data_in[3]));
Q_AN02 U2291 ( .A0(n1), .A1(kme_internal_out[2]), .Z(tlv_sb_data_in[2]));
Q_AN02 U2292 ( .A0(n1), .A1(kme_internal_out[1]), .Z(tlv_sb_data_in[1]));
Q_AN02 U2293 ( .A0(n1), .A1(kme_internal_out[0]), .Z(tlv_sb_data_in[0]));
Q_MX02 U2294 ( .S(n31), .A0(n69), .A1(stream_cmd_in[262]), .Z(stream_cmd_in_nxt[262]));
Q_AN02 U2295 ( .A0(n31), .A1(stream_cmd_in[261]), .Z(stream_cmd_in_nxt[261]));
Q_MX02 U2296 ( .S(n72), .A0(stream_cmd_in[196]), .A1(n854), .Z(stream_cmd_in_nxt[260]));
Q_AN02 U2297 ( .A0(n30), .A1(stream_cmd_in[260]), .Z(n854));
Q_MX02 U2298 ( .S(n72), .A0(stream_cmd_in[195]), .A1(n855), .Z(stream_cmd_in_nxt[259]));
Q_AN02 U2299 ( .A0(n30), .A1(stream_cmd_in[259]), .Z(n855));
Q_MX02 U2300 ( .S(n72), .A0(stream_cmd_in[194]), .A1(n856), .Z(stream_cmd_in_nxt[258]));
Q_AN02 U2301 ( .A0(n30), .A1(stream_cmd_in[258]), .Z(n856));
Q_MX02 U2302 ( .S(n72), .A0(stream_cmd_in[193]), .A1(n857), .Z(stream_cmd_in_nxt[257]));
Q_AN02 U2303 ( .A0(n30), .A1(stream_cmd_in[257]), .Z(n857));
Q_MX02 U2304 ( .S(n72), .A0(stream_cmd_in[192]), .A1(n858), .Z(stream_cmd_in_nxt[256]));
Q_AN02 U2305 ( .A0(n30), .A1(stream_cmd_in[256]), .Z(n858));
Q_MX02 U2306 ( .S(n72), .A0(stream_cmd_in[191]), .A1(n859), .Z(stream_cmd_in_nxt[255]));
Q_AN02 U2307 ( .A0(n30), .A1(stream_cmd_in[255]), .Z(n859));
Q_MX02 U2308 ( .S(n72), .A0(stream_cmd_in[190]), .A1(n860), .Z(stream_cmd_in_nxt[254]));
Q_AN02 U2309 ( .A0(n30), .A1(stream_cmd_in[254]), .Z(n860));
Q_MX02 U2310 ( .S(n72), .A0(stream_cmd_in[189]), .A1(n861), .Z(stream_cmd_in_nxt[253]));
Q_AN02 U2311 ( .A0(n30), .A1(stream_cmd_in[253]), .Z(n861));
Q_MX02 U2312 ( .S(n72), .A0(stream_cmd_in[188]), .A1(n862), .Z(stream_cmd_in_nxt[252]));
Q_AN02 U2313 ( .A0(n30), .A1(stream_cmd_in[252]), .Z(n862));
Q_MX02 U2314 ( .S(n72), .A0(stream_cmd_in[187]), .A1(n863), .Z(stream_cmd_in_nxt[251]));
Q_AN02 U2315 ( .A0(n30), .A1(stream_cmd_in[251]), .Z(n863));
Q_MX02 U2316 ( .S(n72), .A0(stream_cmd_in[186]), .A1(n864), .Z(stream_cmd_in_nxt[250]));
Q_AN02 U2317 ( .A0(n30), .A1(stream_cmd_in[250]), .Z(n864));
Q_MX02 U2318 ( .S(n72), .A0(stream_cmd_in[185]), .A1(n865), .Z(stream_cmd_in_nxt[249]));
Q_AN02 U2319 ( .A0(n30), .A1(stream_cmd_in[249]), .Z(n865));
Q_MX02 U2320 ( .S(n72), .A0(stream_cmd_in[184]), .A1(n866), .Z(stream_cmd_in_nxt[248]));
Q_AN02 U2321 ( .A0(n30), .A1(stream_cmd_in[248]), .Z(n866));
Q_MX02 U2322 ( .S(n72), .A0(stream_cmd_in[183]), .A1(n867), .Z(stream_cmd_in_nxt[247]));
Q_AN02 U2323 ( .A0(n30), .A1(stream_cmd_in[247]), .Z(n867));
Q_MX02 U2324 ( .S(n72), .A0(stream_cmd_in[182]), .A1(n868), .Z(stream_cmd_in_nxt[246]));
Q_AN02 U2325 ( .A0(n30), .A1(stream_cmd_in[246]), .Z(n868));
Q_MX02 U2326 ( .S(n72), .A0(stream_cmd_in[181]), .A1(n869), .Z(stream_cmd_in_nxt[245]));
Q_AN02 U2327 ( .A0(n30), .A1(stream_cmd_in[245]), .Z(n869));
Q_MX02 U2328 ( .S(n72), .A0(stream_cmd_in[180]), .A1(n870), .Z(stream_cmd_in_nxt[244]));
Q_AN02 U2329 ( .A0(n30), .A1(stream_cmd_in[244]), .Z(n870));
Q_MX02 U2330 ( .S(n72), .A0(stream_cmd_in[179]), .A1(n871), .Z(stream_cmd_in_nxt[243]));
Q_AN02 U2331 ( .A0(n30), .A1(stream_cmd_in[243]), .Z(n871));
Q_MX02 U2332 ( .S(n72), .A0(stream_cmd_in[178]), .A1(n872), .Z(stream_cmd_in_nxt[242]));
Q_AN02 U2333 ( .A0(n30), .A1(stream_cmd_in[242]), .Z(n872));
Q_MX02 U2334 ( .S(n72), .A0(stream_cmd_in[177]), .A1(n873), .Z(stream_cmd_in_nxt[241]));
Q_AN02 U2335 ( .A0(n30), .A1(stream_cmd_in[241]), .Z(n873));
Q_MX02 U2336 ( .S(n72), .A0(stream_cmd_in[176]), .A1(n874), .Z(stream_cmd_in_nxt[240]));
Q_AN02 U2337 ( .A0(n30), .A1(stream_cmd_in[240]), .Z(n874));
Q_MX02 U2338 ( .S(n72), .A0(stream_cmd_in[175]), .A1(n875), .Z(stream_cmd_in_nxt[239]));
Q_AN02 U2339 ( .A0(n30), .A1(stream_cmd_in[239]), .Z(n875));
Q_MX02 U2340 ( .S(n72), .A0(stream_cmd_in[174]), .A1(n876), .Z(stream_cmd_in_nxt[238]));
Q_AN02 U2341 ( .A0(n30), .A1(stream_cmd_in[238]), .Z(n876));
Q_MX02 U2342 ( .S(n72), .A0(stream_cmd_in[173]), .A1(n877), .Z(stream_cmd_in_nxt[237]));
Q_AN02 U2343 ( .A0(n30), .A1(stream_cmd_in[237]), .Z(n877));
Q_MX02 U2344 ( .S(n72), .A0(stream_cmd_in[172]), .A1(n878), .Z(stream_cmd_in_nxt[236]));
Q_AN02 U2345 ( .A0(n30), .A1(stream_cmd_in[236]), .Z(n878));
Q_MX02 U2346 ( .S(n72), .A0(stream_cmd_in[171]), .A1(n879), .Z(stream_cmd_in_nxt[235]));
Q_AN02 U2347 ( .A0(n30), .A1(stream_cmd_in[235]), .Z(n879));
Q_MX02 U2348 ( .S(n72), .A0(stream_cmd_in[170]), .A1(n880), .Z(stream_cmd_in_nxt[234]));
Q_AN02 U2349 ( .A0(n30), .A1(stream_cmd_in[234]), .Z(n880));
Q_MX02 U2350 ( .S(n72), .A0(stream_cmd_in[169]), .A1(n881), .Z(stream_cmd_in_nxt[233]));
Q_AN02 U2351 ( .A0(n30), .A1(stream_cmd_in[233]), .Z(n881));
Q_MX02 U2352 ( .S(n72), .A0(stream_cmd_in[168]), .A1(n882), .Z(stream_cmd_in_nxt[232]));
Q_AN02 U2353 ( .A0(n30), .A1(stream_cmd_in[232]), .Z(n882));
Q_MX02 U2354 ( .S(n72), .A0(stream_cmd_in[167]), .A1(n883), .Z(stream_cmd_in_nxt[231]));
Q_AN02 U2355 ( .A0(n30), .A1(stream_cmd_in[231]), .Z(n883));
Q_MX02 U2356 ( .S(n72), .A0(stream_cmd_in[166]), .A1(n884), .Z(stream_cmd_in_nxt[230]));
Q_AN02 U2357 ( .A0(n30), .A1(stream_cmd_in[230]), .Z(n884));
Q_MX02 U2358 ( .S(n72), .A0(stream_cmd_in[165]), .A1(n885), .Z(stream_cmd_in_nxt[229]));
Q_AN02 U2359 ( .A0(n30), .A1(stream_cmd_in[229]), .Z(n885));
Q_MX02 U2360 ( .S(n72), .A0(stream_cmd_in[164]), .A1(n886), .Z(stream_cmd_in_nxt[228]));
Q_AN02 U2361 ( .A0(n30), .A1(stream_cmd_in[228]), .Z(n886));
Q_MX02 U2362 ( .S(n72), .A0(stream_cmd_in[163]), .A1(n887), .Z(stream_cmd_in_nxt[227]));
Q_AN02 U2363 ( .A0(n30), .A1(stream_cmd_in[227]), .Z(n887));
Q_MX02 U2364 ( .S(n72), .A0(stream_cmd_in[162]), .A1(n888), .Z(stream_cmd_in_nxt[226]));
Q_AN02 U2365 ( .A0(n30), .A1(stream_cmd_in[226]), .Z(n888));
Q_MX02 U2366 ( .S(n72), .A0(stream_cmd_in[161]), .A1(n889), .Z(stream_cmd_in_nxt[225]));
Q_AN02 U2367 ( .A0(n30), .A1(stream_cmd_in[225]), .Z(n889));
Q_MX02 U2368 ( .S(n72), .A0(stream_cmd_in[160]), .A1(n890), .Z(stream_cmd_in_nxt[224]));
Q_AN02 U2369 ( .A0(n30), .A1(stream_cmd_in[224]), .Z(n890));
Q_MX02 U2370 ( .S(n72), .A0(stream_cmd_in[159]), .A1(n891), .Z(stream_cmd_in_nxt[223]));
Q_AN02 U2371 ( .A0(n30), .A1(stream_cmd_in[223]), .Z(n891));
Q_MX02 U2372 ( .S(n72), .A0(stream_cmd_in[158]), .A1(n892), .Z(stream_cmd_in_nxt[222]));
Q_AN02 U2373 ( .A0(n30), .A1(stream_cmd_in[222]), .Z(n892));
Q_MX02 U2374 ( .S(n72), .A0(stream_cmd_in[157]), .A1(n893), .Z(stream_cmd_in_nxt[221]));
Q_AN02 U2375 ( .A0(n30), .A1(stream_cmd_in[221]), .Z(n893));
Q_MX02 U2376 ( .S(n72), .A0(stream_cmd_in[156]), .A1(n894), .Z(stream_cmd_in_nxt[220]));
Q_AN02 U2377 ( .A0(n30), .A1(stream_cmd_in[220]), .Z(n894));
Q_MX02 U2378 ( .S(n72), .A0(stream_cmd_in[155]), .A1(n895), .Z(stream_cmd_in_nxt[219]));
Q_AN02 U2379 ( .A0(n30), .A1(stream_cmd_in[219]), .Z(n895));
Q_MX02 U2380 ( .S(n72), .A0(stream_cmd_in[154]), .A1(n896), .Z(stream_cmd_in_nxt[218]));
Q_AN02 U2381 ( .A0(n30), .A1(stream_cmd_in[218]), .Z(n896));
Q_MX02 U2382 ( .S(n72), .A0(stream_cmd_in[153]), .A1(n897), .Z(stream_cmd_in_nxt[217]));
Q_AN02 U2383 ( .A0(n30), .A1(stream_cmd_in[217]), .Z(n897));
Q_MX02 U2384 ( .S(n72), .A0(stream_cmd_in[152]), .A1(n898), .Z(stream_cmd_in_nxt[216]));
Q_AN02 U2385 ( .A0(n30), .A1(stream_cmd_in[216]), .Z(n898));
Q_MX02 U2386 ( .S(n72), .A0(stream_cmd_in[151]), .A1(n899), .Z(stream_cmd_in_nxt[215]));
Q_AN02 U2387 ( .A0(n30), .A1(stream_cmd_in[215]), .Z(n899));
Q_MX02 U2388 ( .S(n72), .A0(stream_cmd_in[150]), .A1(n900), .Z(stream_cmd_in_nxt[214]));
Q_AN02 U2389 ( .A0(n30), .A1(stream_cmd_in[214]), .Z(n900));
Q_MX02 U2390 ( .S(n72), .A0(stream_cmd_in[149]), .A1(n901), .Z(stream_cmd_in_nxt[213]));
Q_AN02 U2391 ( .A0(n30), .A1(stream_cmd_in[213]), .Z(n901));
Q_MX02 U2392 ( .S(n72), .A0(stream_cmd_in[148]), .A1(n902), .Z(stream_cmd_in_nxt[212]));
Q_AN02 U2393 ( .A0(n30), .A1(stream_cmd_in[212]), .Z(n902));
Q_MX02 U2394 ( .S(n72), .A0(stream_cmd_in[147]), .A1(n903), .Z(stream_cmd_in_nxt[211]));
Q_AN02 U2395 ( .A0(n30), .A1(stream_cmd_in[211]), .Z(n903));
Q_MX02 U2396 ( .S(n72), .A0(stream_cmd_in[146]), .A1(n904), .Z(stream_cmd_in_nxt[210]));
Q_AN02 U2397 ( .A0(n30), .A1(stream_cmd_in[210]), .Z(n904));
Q_MX02 U2398 ( .S(n72), .A0(stream_cmd_in[145]), .A1(n905), .Z(stream_cmd_in_nxt[209]));
Q_AN02 U2399 ( .A0(n30), .A1(stream_cmd_in[209]), .Z(n905));
Q_MX02 U2400 ( .S(n72), .A0(stream_cmd_in[144]), .A1(n906), .Z(stream_cmd_in_nxt[208]));
Q_AN02 U2401 ( .A0(n30), .A1(stream_cmd_in[208]), .Z(n906));
Q_MX02 U2402 ( .S(n72), .A0(stream_cmd_in[143]), .A1(n907), .Z(stream_cmd_in_nxt[207]));
Q_AN02 U2403 ( .A0(n30), .A1(stream_cmd_in[207]), .Z(n907));
Q_MX02 U2404 ( .S(n72), .A0(stream_cmd_in[142]), .A1(n908), .Z(stream_cmd_in_nxt[206]));
Q_AN02 U2405 ( .A0(n30), .A1(stream_cmd_in[206]), .Z(n908));
Q_MX02 U2406 ( .S(n72), .A0(stream_cmd_in[141]), .A1(n909), .Z(stream_cmd_in_nxt[205]));
Q_AN02 U2407 ( .A0(n30), .A1(stream_cmd_in[205]), .Z(n909));
Q_MX02 U2408 ( .S(n72), .A0(stream_cmd_in[140]), .A1(n910), .Z(stream_cmd_in_nxt[204]));
Q_AN02 U2409 ( .A0(n30), .A1(stream_cmd_in[204]), .Z(n910));
Q_MX02 U2410 ( .S(n72), .A0(stream_cmd_in[139]), .A1(n911), .Z(stream_cmd_in_nxt[203]));
Q_AN02 U2411 ( .A0(n30), .A1(stream_cmd_in[203]), .Z(n911));
Q_MX02 U2412 ( .S(n72), .A0(stream_cmd_in[138]), .A1(n912), .Z(stream_cmd_in_nxt[202]));
Q_AN02 U2413 ( .A0(n30), .A1(stream_cmd_in[202]), .Z(n912));
Q_MX02 U2414 ( .S(n72), .A0(stream_cmd_in[137]), .A1(n913), .Z(stream_cmd_in_nxt[201]));
Q_AN02 U2415 ( .A0(n30), .A1(stream_cmd_in[201]), .Z(n913));
Q_MX02 U2416 ( .S(n72), .A0(stream_cmd_in[136]), .A1(n914), .Z(stream_cmd_in_nxt[200]));
Q_AN02 U2417 ( .A0(n30), .A1(stream_cmd_in[200]), .Z(n914));
Q_MX02 U2418 ( .S(n72), .A0(stream_cmd_in[135]), .A1(n915), .Z(stream_cmd_in_nxt[199]));
Q_AN02 U2419 ( .A0(n30), .A1(stream_cmd_in[199]), .Z(n915));
Q_MX02 U2420 ( .S(n72), .A0(stream_cmd_in[134]), .A1(n916), .Z(stream_cmd_in_nxt[198]));
Q_AN02 U2421 ( .A0(n30), .A1(stream_cmd_in[198]), .Z(n916));
Q_MX02 U2422 ( .S(n72), .A0(stream_cmd_in[133]), .A1(n917), .Z(stream_cmd_in_nxt[197]));
Q_AN02 U2423 ( .A0(n30), .A1(stream_cmd_in[197]), .Z(n917));
Q_MX02 U2424 ( .S(n72), .A0(stream_cmd_in[132]), .A1(n918), .Z(stream_cmd_in_nxt[196]));
Q_AN02 U2425 ( .A0(n30), .A1(stream_cmd_in[196]), .Z(n918));
Q_MX02 U2426 ( .S(n72), .A0(stream_cmd_in[131]), .A1(n919), .Z(stream_cmd_in_nxt[195]));
Q_AN02 U2427 ( .A0(n30), .A1(stream_cmd_in[195]), .Z(n919));
Q_MX02 U2428 ( .S(n72), .A0(stream_cmd_in[130]), .A1(n920), .Z(stream_cmd_in_nxt[194]));
Q_AN02 U2429 ( .A0(n30), .A1(stream_cmd_in[194]), .Z(n920));
Q_MX02 U2430 ( .S(n72), .A0(stream_cmd_in[129]), .A1(n921), .Z(stream_cmd_in_nxt[193]));
Q_AN02 U2431 ( .A0(n30), .A1(stream_cmd_in[193]), .Z(n921));
Q_MX02 U2432 ( .S(n72), .A0(stream_cmd_in[128]), .A1(n922), .Z(stream_cmd_in_nxt[192]));
Q_AN02 U2433 ( .A0(n30), .A1(stream_cmd_in[192]), .Z(n922));
Q_MX02 U2434 ( .S(n72), .A0(stream_cmd_in[127]), .A1(n923), .Z(stream_cmd_in_nxt[191]));
Q_AN02 U2435 ( .A0(n30), .A1(stream_cmd_in[191]), .Z(n923));
Q_MX02 U2436 ( .S(n72), .A0(stream_cmd_in[126]), .A1(n924), .Z(stream_cmd_in_nxt[190]));
Q_AN02 U2437 ( .A0(n30), .A1(stream_cmd_in[190]), .Z(n924));
Q_MX02 U2438 ( .S(n72), .A0(stream_cmd_in[125]), .A1(n925), .Z(stream_cmd_in_nxt[189]));
Q_AN02 U2439 ( .A0(n30), .A1(stream_cmd_in[189]), .Z(n925));
Q_MX02 U2440 ( .S(n72), .A0(stream_cmd_in[124]), .A1(n926), .Z(stream_cmd_in_nxt[188]));
Q_AN02 U2441 ( .A0(n30), .A1(stream_cmd_in[188]), .Z(n926));
Q_MX02 U2442 ( .S(n72), .A0(stream_cmd_in[123]), .A1(n927), .Z(stream_cmd_in_nxt[187]));
Q_AN02 U2443 ( .A0(n30), .A1(stream_cmd_in[187]), .Z(n927));
Q_MX02 U2444 ( .S(n72), .A0(stream_cmd_in[122]), .A1(n928), .Z(stream_cmd_in_nxt[186]));
Q_AN02 U2445 ( .A0(n30), .A1(stream_cmd_in[186]), .Z(n928));
Q_MX02 U2446 ( .S(n72), .A0(stream_cmd_in[121]), .A1(n929), .Z(stream_cmd_in_nxt[185]));
Q_AN02 U2447 ( .A0(n30), .A1(stream_cmd_in[185]), .Z(n929));
Q_MX02 U2448 ( .S(n72), .A0(stream_cmd_in[120]), .A1(n930), .Z(stream_cmd_in_nxt[184]));
Q_AN02 U2449 ( .A0(n30), .A1(stream_cmd_in[184]), .Z(n930));
Q_MX02 U2450 ( .S(n72), .A0(stream_cmd_in[119]), .A1(n931), .Z(stream_cmd_in_nxt[183]));
Q_AN02 U2451 ( .A0(n30), .A1(stream_cmd_in[183]), .Z(n931));
Q_MX02 U2452 ( .S(n72), .A0(stream_cmd_in[118]), .A1(n932), .Z(stream_cmd_in_nxt[182]));
Q_AN02 U2453 ( .A0(n30), .A1(stream_cmd_in[182]), .Z(n932));
Q_MX02 U2454 ( .S(n72), .A0(stream_cmd_in[117]), .A1(n933), .Z(stream_cmd_in_nxt[181]));
Q_AN02 U2455 ( .A0(n30), .A1(stream_cmd_in[181]), .Z(n933));
Q_MX02 U2456 ( .S(n72), .A0(stream_cmd_in[116]), .A1(n934), .Z(stream_cmd_in_nxt[180]));
Q_AN02 U2457 ( .A0(n30), .A1(stream_cmd_in[180]), .Z(n934));
Q_MX02 U2458 ( .S(n72), .A0(stream_cmd_in[115]), .A1(n935), .Z(stream_cmd_in_nxt[179]));
Q_AN02 U2459 ( .A0(n30), .A1(stream_cmd_in[179]), .Z(n935));
Q_MX02 U2460 ( .S(n72), .A0(stream_cmd_in[114]), .A1(n936), .Z(stream_cmd_in_nxt[178]));
Q_AN02 U2461 ( .A0(n30), .A1(stream_cmd_in[178]), .Z(n936));
Q_MX02 U2462 ( .S(n72), .A0(stream_cmd_in[113]), .A1(n937), .Z(stream_cmd_in_nxt[177]));
Q_AN02 U2463 ( .A0(n30), .A1(stream_cmd_in[177]), .Z(n937));
Q_MX02 U2464 ( .S(n72), .A0(stream_cmd_in[112]), .A1(n938), .Z(stream_cmd_in_nxt[176]));
Q_AN02 U2465 ( .A0(n30), .A1(stream_cmd_in[176]), .Z(n938));
Q_MX02 U2466 ( .S(n72), .A0(stream_cmd_in[111]), .A1(n939), .Z(stream_cmd_in_nxt[175]));
Q_AN02 U2467 ( .A0(n30), .A1(stream_cmd_in[175]), .Z(n939));
Q_MX02 U2468 ( .S(n72), .A0(stream_cmd_in[110]), .A1(n940), .Z(stream_cmd_in_nxt[174]));
Q_AN02 U2469 ( .A0(n30), .A1(stream_cmd_in[174]), .Z(n940));
Q_MX02 U2470 ( .S(n72), .A0(stream_cmd_in[109]), .A1(n941), .Z(stream_cmd_in_nxt[173]));
Q_AN02 U2471 ( .A0(n30), .A1(stream_cmd_in[173]), .Z(n941));
Q_MX02 U2472 ( .S(n72), .A0(stream_cmd_in[108]), .A1(n942), .Z(stream_cmd_in_nxt[172]));
Q_AN02 U2473 ( .A0(n30), .A1(stream_cmd_in[172]), .Z(n942));
Q_MX02 U2474 ( .S(n72), .A0(stream_cmd_in[107]), .A1(n943), .Z(stream_cmd_in_nxt[171]));
Q_AN02 U2475 ( .A0(n30), .A1(stream_cmd_in[171]), .Z(n943));
Q_MX02 U2476 ( .S(n72), .A0(stream_cmd_in[106]), .A1(n944), .Z(stream_cmd_in_nxt[170]));
Q_AN02 U2477 ( .A0(n30), .A1(stream_cmd_in[170]), .Z(n944));
Q_MX02 U2478 ( .S(n72), .A0(stream_cmd_in[105]), .A1(n945), .Z(stream_cmd_in_nxt[169]));
Q_AN02 U2479 ( .A0(n30), .A1(stream_cmd_in[169]), .Z(n945));
Q_MX02 U2480 ( .S(n72), .A0(stream_cmd_in[104]), .A1(n946), .Z(stream_cmd_in_nxt[168]));
Q_AN02 U2481 ( .A0(n30), .A1(stream_cmd_in[168]), .Z(n946));
Q_MX02 U2482 ( .S(n72), .A0(stream_cmd_in[103]), .A1(n947), .Z(stream_cmd_in_nxt[167]));
Q_AN02 U2483 ( .A0(n30), .A1(stream_cmd_in[167]), .Z(n947));
Q_MX02 U2484 ( .S(n72), .A0(stream_cmd_in[102]), .A1(n948), .Z(stream_cmd_in_nxt[166]));
Q_AN02 U2485 ( .A0(n30), .A1(stream_cmd_in[166]), .Z(n948));
Q_MX02 U2486 ( .S(n72), .A0(stream_cmd_in[101]), .A1(n949), .Z(stream_cmd_in_nxt[165]));
Q_AN02 U2487 ( .A0(n30), .A1(stream_cmd_in[165]), .Z(n949));
Q_MX02 U2488 ( .S(n72), .A0(stream_cmd_in[100]), .A1(n950), .Z(stream_cmd_in_nxt[164]));
Q_AN02 U2489 ( .A0(n30), .A1(stream_cmd_in[164]), .Z(n950));
Q_MX02 U2490 ( .S(n72), .A0(stream_cmd_in[99]), .A1(n951), .Z(stream_cmd_in_nxt[163]));
Q_AN02 U2491 ( .A0(n30), .A1(stream_cmd_in[163]), .Z(n951));
Q_MX02 U2492 ( .S(n72), .A0(stream_cmd_in[98]), .A1(n952), .Z(stream_cmd_in_nxt[162]));
Q_AN02 U2493 ( .A0(n30), .A1(stream_cmd_in[162]), .Z(n952));
Q_MX02 U2494 ( .S(n72), .A0(stream_cmd_in[97]), .A1(n953), .Z(stream_cmd_in_nxt[161]));
Q_AN02 U2495 ( .A0(n30), .A1(stream_cmd_in[161]), .Z(n953));
Q_MX02 U2496 ( .S(n72), .A0(stream_cmd_in[96]), .A1(n954), .Z(stream_cmd_in_nxt[160]));
Q_AN02 U2497 ( .A0(n30), .A1(stream_cmd_in[160]), .Z(n954));
Q_MX02 U2498 ( .S(n72), .A0(stream_cmd_in[95]), .A1(n955), .Z(stream_cmd_in_nxt[159]));
Q_AN02 U2499 ( .A0(n30), .A1(stream_cmd_in[159]), .Z(n955));
Q_MX02 U2500 ( .S(n72), .A0(stream_cmd_in[94]), .A1(n956), .Z(stream_cmd_in_nxt[158]));
Q_AN02 U2501 ( .A0(n30), .A1(stream_cmd_in[158]), .Z(n956));
Q_MX02 U2502 ( .S(n72), .A0(stream_cmd_in[93]), .A1(n957), .Z(stream_cmd_in_nxt[157]));
Q_AN02 U2503 ( .A0(n30), .A1(stream_cmd_in[157]), .Z(n957));
Q_MX02 U2504 ( .S(n72), .A0(stream_cmd_in[92]), .A1(n958), .Z(stream_cmd_in_nxt[156]));
Q_AN02 U2505 ( .A0(n30), .A1(stream_cmd_in[156]), .Z(n958));
Q_MX02 U2506 ( .S(n72), .A0(stream_cmd_in[91]), .A1(n959), .Z(stream_cmd_in_nxt[155]));
Q_AN02 U2507 ( .A0(n30), .A1(stream_cmd_in[155]), .Z(n959));
Q_MX02 U2508 ( .S(n72), .A0(stream_cmd_in[90]), .A1(n960), .Z(stream_cmd_in_nxt[154]));
Q_AN02 U2509 ( .A0(n30), .A1(stream_cmd_in[154]), .Z(n960));
Q_MX02 U2510 ( .S(n72), .A0(stream_cmd_in[89]), .A1(n961), .Z(stream_cmd_in_nxt[153]));
Q_AN02 U2511 ( .A0(n30), .A1(stream_cmd_in[153]), .Z(n961));
Q_MX02 U2512 ( .S(n72), .A0(stream_cmd_in[88]), .A1(n962), .Z(stream_cmd_in_nxt[152]));
Q_AN02 U2513 ( .A0(n30), .A1(stream_cmd_in[152]), .Z(n962));
Q_MX02 U2514 ( .S(n72), .A0(stream_cmd_in[87]), .A1(n963), .Z(stream_cmd_in_nxt[151]));
Q_AN02 U2515 ( .A0(n30), .A1(stream_cmd_in[151]), .Z(n963));
Q_MX02 U2516 ( .S(n72), .A0(stream_cmd_in[86]), .A1(n964), .Z(stream_cmd_in_nxt[150]));
Q_AN02 U2517 ( .A0(n30), .A1(stream_cmd_in[150]), .Z(n964));
Q_MX02 U2518 ( .S(n72), .A0(stream_cmd_in[85]), .A1(n965), .Z(stream_cmd_in_nxt[149]));
Q_AN02 U2519 ( .A0(n30), .A1(stream_cmd_in[149]), .Z(n965));
Q_MX02 U2520 ( .S(n72), .A0(stream_cmd_in[84]), .A1(n966), .Z(stream_cmd_in_nxt[148]));
Q_AN02 U2521 ( .A0(n30), .A1(stream_cmd_in[148]), .Z(n966));
Q_MX02 U2522 ( .S(n72), .A0(stream_cmd_in[83]), .A1(n967), .Z(stream_cmd_in_nxt[147]));
Q_AN02 U2523 ( .A0(n30), .A1(stream_cmd_in[147]), .Z(n967));
Q_MX02 U2524 ( .S(n72), .A0(stream_cmd_in[82]), .A1(n968), .Z(stream_cmd_in_nxt[146]));
Q_AN02 U2525 ( .A0(n30), .A1(stream_cmd_in[146]), .Z(n968));
Q_MX02 U2526 ( .S(n72), .A0(stream_cmd_in[81]), .A1(n969), .Z(stream_cmd_in_nxt[145]));
Q_AN02 U2527 ( .A0(n30), .A1(stream_cmd_in[145]), .Z(n969));
Q_MX02 U2528 ( .S(n72), .A0(stream_cmd_in[80]), .A1(n970), .Z(stream_cmd_in_nxt[144]));
Q_AN02 U2529 ( .A0(n30), .A1(stream_cmd_in[144]), .Z(n970));
Q_MX02 U2530 ( .S(n72), .A0(stream_cmd_in[79]), .A1(n971), .Z(stream_cmd_in_nxt[143]));
Q_AN02 U2531 ( .A0(n30), .A1(stream_cmd_in[143]), .Z(n971));
Q_MX02 U2532 ( .S(n72), .A0(stream_cmd_in[78]), .A1(n972), .Z(stream_cmd_in_nxt[142]));
Q_AN02 U2533 ( .A0(n30), .A1(stream_cmd_in[142]), .Z(n972));
Q_MX02 U2534 ( .S(n72), .A0(stream_cmd_in[77]), .A1(n973), .Z(stream_cmd_in_nxt[141]));
Q_AN02 U2535 ( .A0(n30), .A1(stream_cmd_in[141]), .Z(n973));
Q_MX02 U2536 ( .S(n72), .A0(stream_cmd_in[76]), .A1(n974), .Z(stream_cmd_in_nxt[140]));
Q_AN02 U2537 ( .A0(n30), .A1(stream_cmd_in[140]), .Z(n974));
Q_MX02 U2538 ( .S(n72), .A0(stream_cmd_in[75]), .A1(n975), .Z(stream_cmd_in_nxt[139]));
Q_AN02 U2539 ( .A0(n30), .A1(stream_cmd_in[139]), .Z(n975));
Q_MX02 U2540 ( .S(n72), .A0(stream_cmd_in[74]), .A1(n976), .Z(stream_cmd_in_nxt[138]));
Q_AN02 U2541 ( .A0(n30), .A1(stream_cmd_in[138]), .Z(n976));
Q_MX02 U2542 ( .S(n72), .A0(stream_cmd_in[73]), .A1(n977), .Z(stream_cmd_in_nxt[137]));
Q_AN02 U2543 ( .A0(n30), .A1(stream_cmd_in[137]), .Z(n977));
Q_MX02 U2544 ( .S(n72), .A0(stream_cmd_in[72]), .A1(n978), .Z(stream_cmd_in_nxt[136]));
Q_AN02 U2545 ( .A0(n30), .A1(stream_cmd_in[136]), .Z(n978));
Q_MX02 U2546 ( .S(n72), .A0(stream_cmd_in[71]), .A1(n979), .Z(stream_cmd_in_nxt[135]));
Q_AN02 U2547 ( .A0(n30), .A1(stream_cmd_in[135]), .Z(n979));
Q_MX02 U2548 ( .S(n72), .A0(stream_cmd_in[70]), .A1(n980), .Z(stream_cmd_in_nxt[134]));
Q_AN02 U2549 ( .A0(n30), .A1(stream_cmd_in[134]), .Z(n980));
Q_MX02 U2550 ( .S(n72), .A0(stream_cmd_in[69]), .A1(n981), .Z(stream_cmd_in_nxt[133]));
Q_AN02 U2551 ( .A0(n30), .A1(stream_cmd_in[133]), .Z(n981));
Q_MX02 U2552 ( .S(n72), .A0(stream_cmd_in[68]), .A1(n982), .Z(stream_cmd_in_nxt[132]));
Q_AN02 U2553 ( .A0(n30), .A1(stream_cmd_in[132]), .Z(n982));
Q_MX02 U2554 ( .S(n72), .A0(stream_cmd_in[67]), .A1(n983), .Z(stream_cmd_in_nxt[131]));
Q_AN02 U2555 ( .A0(n30), .A1(stream_cmd_in[131]), .Z(n983));
Q_MX02 U2556 ( .S(n72), .A0(stream_cmd_in[66]), .A1(n984), .Z(stream_cmd_in_nxt[130]));
Q_AN02 U2557 ( .A0(n30), .A1(stream_cmd_in[130]), .Z(n984));
Q_MX02 U2558 ( .S(n72), .A0(stream_cmd_in[65]), .A1(n985), .Z(stream_cmd_in_nxt[129]));
Q_AN02 U2559 ( .A0(n30), .A1(stream_cmd_in[129]), .Z(n985));
Q_MX02 U2560 ( .S(n72), .A0(stream_cmd_in[64]), .A1(n986), .Z(stream_cmd_in_nxt[128]));
Q_AN02 U2561 ( .A0(n30), .A1(stream_cmd_in[128]), .Z(n986));
Q_MX02 U2562 ( .S(n72), .A0(stream_cmd_in[63]), .A1(n987), .Z(stream_cmd_in_nxt[127]));
Q_AN02 U2563 ( .A0(n30), .A1(stream_cmd_in[127]), .Z(n987));
Q_MX02 U2564 ( .S(n72), .A0(stream_cmd_in[62]), .A1(n988), .Z(stream_cmd_in_nxt[126]));
Q_AN02 U2565 ( .A0(n30), .A1(stream_cmd_in[126]), .Z(n988));
Q_MX02 U2566 ( .S(n72), .A0(stream_cmd_in[61]), .A1(n989), .Z(stream_cmd_in_nxt[125]));
Q_AN02 U2567 ( .A0(n30), .A1(stream_cmd_in[125]), .Z(n989));
Q_MX02 U2568 ( .S(n72), .A0(stream_cmd_in[60]), .A1(n990), .Z(stream_cmd_in_nxt[124]));
Q_AN02 U2569 ( .A0(n30), .A1(stream_cmd_in[124]), .Z(n990));
Q_MX02 U2570 ( .S(n72), .A0(stream_cmd_in[59]), .A1(n991), .Z(stream_cmd_in_nxt[123]));
Q_AN02 U2571 ( .A0(n30), .A1(stream_cmd_in[123]), .Z(n991));
Q_MX02 U2572 ( .S(n72), .A0(stream_cmd_in[58]), .A1(n992), .Z(stream_cmd_in_nxt[122]));
Q_AN02 U2573 ( .A0(n30), .A1(stream_cmd_in[122]), .Z(n992));
Q_MX02 U2574 ( .S(n72), .A0(stream_cmd_in[57]), .A1(n993), .Z(stream_cmd_in_nxt[121]));
Q_AN02 U2575 ( .A0(n30), .A1(stream_cmd_in[121]), .Z(n993));
Q_MX02 U2576 ( .S(n72), .A0(stream_cmd_in[56]), .A1(n994), .Z(stream_cmd_in_nxt[120]));
Q_AN02 U2577 ( .A0(n30), .A1(stream_cmd_in[120]), .Z(n994));
Q_MX02 U2578 ( .S(n72), .A0(stream_cmd_in[55]), .A1(n995), .Z(stream_cmd_in_nxt[119]));
Q_AN02 U2579 ( .A0(n30), .A1(stream_cmd_in[119]), .Z(n995));
Q_MX02 U2580 ( .S(n72), .A0(stream_cmd_in[54]), .A1(n996), .Z(stream_cmd_in_nxt[118]));
Q_AN02 U2581 ( .A0(n30), .A1(stream_cmd_in[118]), .Z(n996));
Q_MX02 U2582 ( .S(n72), .A0(stream_cmd_in[53]), .A1(n997), .Z(stream_cmd_in_nxt[117]));
Q_AN02 U2583 ( .A0(n30), .A1(stream_cmd_in[117]), .Z(n997));
Q_MX02 U2584 ( .S(n72), .A0(stream_cmd_in[52]), .A1(n998), .Z(stream_cmd_in_nxt[116]));
Q_AN02 U2585 ( .A0(n30), .A1(stream_cmd_in[116]), .Z(n998));
Q_MX02 U2586 ( .S(n72), .A0(stream_cmd_in[51]), .A1(n999), .Z(stream_cmd_in_nxt[115]));
Q_AN02 U2587 ( .A0(n30), .A1(stream_cmd_in[115]), .Z(n999));
Q_MX02 U2588 ( .S(n72), .A0(stream_cmd_in[50]), .A1(n1000), .Z(stream_cmd_in_nxt[114]));
Q_AN02 U2589 ( .A0(n30), .A1(stream_cmd_in[114]), .Z(n1000));
Q_MX02 U2590 ( .S(n72), .A0(stream_cmd_in[49]), .A1(n1001), .Z(stream_cmd_in_nxt[113]));
Q_AN02 U2591 ( .A0(n30), .A1(stream_cmd_in[113]), .Z(n1001));
Q_MX02 U2592 ( .S(n72), .A0(stream_cmd_in[48]), .A1(n1002), .Z(stream_cmd_in_nxt[112]));
Q_AN02 U2593 ( .A0(n30), .A1(stream_cmd_in[112]), .Z(n1002));
Q_MX02 U2594 ( .S(n72), .A0(stream_cmd_in[47]), .A1(n1003), .Z(stream_cmd_in_nxt[111]));
Q_AN02 U2595 ( .A0(n30), .A1(stream_cmd_in[111]), .Z(n1003));
Q_MX02 U2596 ( .S(n72), .A0(stream_cmd_in[46]), .A1(n1004), .Z(stream_cmd_in_nxt[110]));
Q_AN02 U2597 ( .A0(n30), .A1(stream_cmd_in[110]), .Z(n1004));
Q_MX02 U2598 ( .S(n72), .A0(stream_cmd_in[45]), .A1(n1005), .Z(stream_cmd_in_nxt[109]));
Q_AN02 U2599 ( .A0(n30), .A1(stream_cmd_in[109]), .Z(n1005));
Q_MX02 U2600 ( .S(n72), .A0(stream_cmd_in[44]), .A1(n1006), .Z(stream_cmd_in_nxt[108]));
Q_AN02 U2601 ( .A0(n30), .A1(stream_cmd_in[108]), .Z(n1006));
Q_MX02 U2602 ( .S(n72), .A0(stream_cmd_in[43]), .A1(n1007), .Z(stream_cmd_in_nxt[107]));
Q_AN02 U2603 ( .A0(n30), .A1(stream_cmd_in[107]), .Z(n1007));
Q_MX02 U2604 ( .S(n72), .A0(stream_cmd_in[42]), .A1(n1008), .Z(stream_cmd_in_nxt[106]));
Q_AN02 U2605 ( .A0(n30), .A1(stream_cmd_in[106]), .Z(n1008));
Q_MX02 U2606 ( .S(n72), .A0(stream_cmd_in[41]), .A1(n1009), .Z(stream_cmd_in_nxt[105]));
Q_AN02 U2607 ( .A0(n30), .A1(stream_cmd_in[105]), .Z(n1009));
Q_MX02 U2608 ( .S(n72), .A0(stream_cmd_in[40]), .A1(n1010), .Z(stream_cmd_in_nxt[104]));
Q_AN02 U2609 ( .A0(n30), .A1(stream_cmd_in[104]), .Z(n1010));
Q_MX02 U2610 ( .S(n72), .A0(stream_cmd_in[39]), .A1(n1011), .Z(stream_cmd_in_nxt[103]));
Q_AN02 U2611 ( .A0(n30), .A1(stream_cmd_in[103]), .Z(n1011));
Q_MX02 U2612 ( .S(n72), .A0(stream_cmd_in[38]), .A1(n1012), .Z(stream_cmd_in_nxt[102]));
Q_AN02 U2613 ( .A0(n30), .A1(stream_cmd_in[102]), .Z(n1012));
Q_MX02 U2614 ( .S(n72), .A0(stream_cmd_in[37]), .A1(n1013), .Z(stream_cmd_in_nxt[101]));
Q_AN02 U2615 ( .A0(n30), .A1(stream_cmd_in[101]), .Z(n1013));
Q_MX02 U2616 ( .S(n72), .A0(stream_cmd_in[36]), .A1(n1014), .Z(stream_cmd_in_nxt[100]));
Q_AN02 U2617 ( .A0(n30), .A1(stream_cmd_in[100]), .Z(n1014));
Q_MX02 U2618 ( .S(n72), .A0(stream_cmd_in[35]), .A1(n1015), .Z(stream_cmd_in_nxt[99]));
Q_AN02 U2619 ( .A0(n30), .A1(stream_cmd_in[99]), .Z(n1015));
Q_MX02 U2620 ( .S(n72), .A0(stream_cmd_in[34]), .A1(n1016), .Z(stream_cmd_in_nxt[98]));
Q_AN02 U2621 ( .A0(n30), .A1(stream_cmd_in[98]), .Z(n1016));
Q_MX02 U2622 ( .S(n72), .A0(stream_cmd_in[33]), .A1(n1017), .Z(stream_cmd_in_nxt[97]));
Q_AN02 U2623 ( .A0(n30), .A1(stream_cmd_in[97]), .Z(n1017));
Q_MX02 U2624 ( .S(n72), .A0(stream_cmd_in[32]), .A1(n1018), .Z(stream_cmd_in_nxt[96]));
Q_AN02 U2625 ( .A0(n30), .A1(stream_cmd_in[96]), .Z(n1018));
Q_MX02 U2626 ( .S(n72), .A0(stream_cmd_in[31]), .A1(n1019), .Z(stream_cmd_in_nxt[95]));
Q_AN02 U2627 ( .A0(n30), .A1(stream_cmd_in[95]), .Z(n1019));
Q_MX02 U2628 ( .S(n72), .A0(stream_cmd_in[30]), .A1(n1020), .Z(stream_cmd_in_nxt[94]));
Q_AN02 U2629 ( .A0(n30), .A1(stream_cmd_in[94]), .Z(n1020));
Q_MX02 U2630 ( .S(n72), .A0(stream_cmd_in[29]), .A1(n1021), .Z(stream_cmd_in_nxt[93]));
Q_AN02 U2631 ( .A0(n30), .A1(stream_cmd_in[93]), .Z(n1021));
Q_MX02 U2632 ( .S(n72), .A0(stream_cmd_in[28]), .A1(n1022), .Z(stream_cmd_in_nxt[92]));
Q_AN02 U2633 ( .A0(n30), .A1(stream_cmd_in[92]), .Z(n1022));
Q_MX02 U2634 ( .S(n72), .A0(stream_cmd_in[27]), .A1(n1023), .Z(stream_cmd_in_nxt[91]));
Q_AN02 U2635 ( .A0(n30), .A1(stream_cmd_in[91]), .Z(n1023));
Q_MX02 U2636 ( .S(n72), .A0(stream_cmd_in[26]), .A1(n1024), .Z(stream_cmd_in_nxt[90]));
Q_AN02 U2637 ( .A0(n30), .A1(stream_cmd_in[90]), .Z(n1024));
Q_MX02 U2638 ( .S(n72), .A0(stream_cmd_in[25]), .A1(n1025), .Z(stream_cmd_in_nxt[89]));
Q_AN02 U2639 ( .A0(n30), .A1(stream_cmd_in[89]), .Z(n1025));
Q_MX02 U2640 ( .S(n72), .A0(stream_cmd_in[24]), .A1(n1026), .Z(stream_cmd_in_nxt[88]));
Q_AN02 U2641 ( .A0(n30), .A1(stream_cmd_in[88]), .Z(n1026));
Q_MX02 U2642 ( .S(n72), .A0(stream_cmd_in[23]), .A1(n1027), .Z(stream_cmd_in_nxt[87]));
Q_AN02 U2643 ( .A0(n30), .A1(stream_cmd_in[87]), .Z(n1027));
Q_MX02 U2644 ( .S(n72), .A0(stream_cmd_in[22]), .A1(n1028), .Z(stream_cmd_in_nxt[86]));
Q_AN02 U2645 ( .A0(n30), .A1(stream_cmd_in[86]), .Z(n1028));
Q_MX02 U2646 ( .S(n72), .A0(stream_cmd_in[21]), .A1(n1029), .Z(stream_cmd_in_nxt[85]));
Q_AN02 U2647 ( .A0(n30), .A1(stream_cmd_in[85]), .Z(n1029));
Q_MX02 U2648 ( .S(n72), .A0(stream_cmd_in[20]), .A1(n1030), .Z(stream_cmd_in_nxt[84]));
Q_AN02 U2649 ( .A0(n30), .A1(stream_cmd_in[84]), .Z(n1030));
Q_MX02 U2650 ( .S(n72), .A0(stream_cmd_in[19]), .A1(n1031), .Z(stream_cmd_in_nxt[83]));
Q_AN02 U2651 ( .A0(n30), .A1(stream_cmd_in[83]), .Z(n1031));
Q_MX02 U2652 ( .S(n72), .A0(stream_cmd_in[18]), .A1(n1032), .Z(stream_cmd_in_nxt[82]));
Q_AN02 U2653 ( .A0(n30), .A1(stream_cmd_in[82]), .Z(n1032));
Q_MX02 U2654 ( .S(n72), .A0(stream_cmd_in[17]), .A1(n1033), .Z(stream_cmd_in_nxt[81]));
Q_AN02 U2655 ( .A0(n30), .A1(stream_cmd_in[81]), .Z(n1033));
Q_MX02 U2656 ( .S(n72), .A0(stream_cmd_in[16]), .A1(n1034), .Z(stream_cmd_in_nxt[80]));
Q_AN02 U2657 ( .A0(n30), .A1(stream_cmd_in[80]), .Z(n1034));
Q_MX02 U2658 ( .S(n72), .A0(stream_cmd_in[15]), .A1(n1035), .Z(stream_cmd_in_nxt[79]));
Q_AN02 U2659 ( .A0(n30), .A1(stream_cmd_in[79]), .Z(n1035));
Q_MX02 U2660 ( .S(n72), .A0(stream_cmd_in[14]), .A1(n1036), .Z(stream_cmd_in_nxt[78]));
Q_AN02 U2661 ( .A0(n30), .A1(stream_cmd_in[78]), .Z(n1036));
Q_MX02 U2662 ( .S(n72), .A0(stream_cmd_in[13]), .A1(n1037), .Z(stream_cmd_in_nxt[77]));
Q_AN02 U2663 ( .A0(n30), .A1(stream_cmd_in[77]), .Z(n1037));
Q_MX02 U2664 ( .S(n72), .A0(stream_cmd_in[12]), .A1(n1038), .Z(stream_cmd_in_nxt[76]));
Q_AN02 U2665 ( .A0(n30), .A1(stream_cmd_in[76]), .Z(n1038));
Q_MX02 U2666 ( .S(n72), .A0(stream_cmd_in[11]), .A1(n1039), .Z(stream_cmd_in_nxt[75]));
Q_AN02 U2667 ( .A0(n30), .A1(stream_cmd_in[75]), .Z(n1039));
Q_MX02 U2668 ( .S(n72), .A0(stream_cmd_in[10]), .A1(n1040), .Z(stream_cmd_in_nxt[74]));
Q_AN02 U2669 ( .A0(n30), .A1(stream_cmd_in[74]), .Z(n1040));
Q_MX02 U2670 ( .S(n72), .A0(stream_cmd_in[9]), .A1(n1041), .Z(stream_cmd_in_nxt[73]));
Q_AN02 U2671 ( .A0(n30), .A1(stream_cmd_in[73]), .Z(n1041));
Q_MX02 U2672 ( .S(n72), .A0(stream_cmd_in[8]), .A1(n1042), .Z(stream_cmd_in_nxt[72]));
Q_AN02 U2673 ( .A0(n30), .A1(stream_cmd_in[72]), .Z(n1042));
Q_MX02 U2674 ( .S(n72), .A0(stream_cmd_in[7]), .A1(n1043), .Z(stream_cmd_in_nxt[71]));
Q_AN02 U2675 ( .A0(n30), .A1(stream_cmd_in[71]), .Z(n1043));
Q_MX02 U2676 ( .S(n72), .A0(stream_cmd_in[6]), .A1(n1044), .Z(stream_cmd_in_nxt[70]));
Q_AN02 U2677 ( .A0(n30), .A1(stream_cmd_in[70]), .Z(n1044));
Q_MX02 U2678 ( .S(n72), .A0(stream_cmd_in[5]), .A1(n1045), .Z(stream_cmd_in_nxt[69]));
Q_AN02 U2679 ( .A0(n30), .A1(stream_cmd_in[69]), .Z(n1045));
Q_MX02 U2680 ( .S(n72), .A0(kme_internal_out[63]), .A1(n1046), .Z(stream_cmd_in_nxt[68]));
Q_AN02 U2681 ( .A0(n30), .A1(stream_cmd_in[68]), .Z(n1046));
Q_MX02 U2682 ( .S(n72), .A0(kme_internal_out[62]), .A1(n1047), .Z(stream_cmd_in_nxt[67]));
Q_AN02 U2683 ( .A0(n30), .A1(stream_cmd_in[67]), .Z(n1047));
Q_MX02 U2684 ( .S(n72), .A0(kme_internal_out[61]), .A1(n1048), .Z(stream_cmd_in_nxt[66]));
Q_AN02 U2685 ( .A0(n30), .A1(stream_cmd_in[66]), .Z(n1048));
Q_MX02 U2686 ( .S(n72), .A0(kme_internal_out[60]), .A1(n1049), .Z(stream_cmd_in_nxt[65]));
Q_AN02 U2687 ( .A0(n30), .A1(stream_cmd_in[65]), .Z(n1049));
Q_MX02 U2688 ( .S(n72), .A0(kme_internal_out[59]), .A1(n1050), .Z(stream_cmd_in_nxt[64]));
Q_AN02 U2689 ( .A0(n30), .A1(stream_cmd_in[64]), .Z(n1050));
Q_MX02 U2690 ( .S(n72), .A0(kme_internal_out[58]), .A1(n1051), .Z(stream_cmd_in_nxt[63]));
Q_AN02 U2691 ( .A0(n30), .A1(stream_cmd_in[63]), .Z(n1051));
Q_MX02 U2692 ( .S(n72), .A0(kme_internal_out[57]), .A1(n1052), .Z(stream_cmd_in_nxt[62]));
Q_AN02 U2693 ( .A0(n30), .A1(stream_cmd_in[62]), .Z(n1052));
Q_MX02 U2694 ( .S(n72), .A0(kme_internal_out[56]), .A1(n1053), .Z(stream_cmd_in_nxt[61]));
Q_AN02 U2695 ( .A0(n30), .A1(stream_cmd_in[61]), .Z(n1053));
Q_MX02 U2696 ( .S(n72), .A0(kme_internal_out[55]), .A1(n1054), .Z(stream_cmd_in_nxt[60]));
Q_AN02 U2697 ( .A0(n30), .A1(stream_cmd_in[60]), .Z(n1054));
Q_MX02 U2698 ( .S(n72), .A0(kme_internal_out[54]), .A1(n1055), .Z(stream_cmd_in_nxt[59]));
Q_AN02 U2699 ( .A0(n30), .A1(stream_cmd_in[59]), .Z(n1055));
Q_MX02 U2700 ( .S(n72), .A0(kme_internal_out[53]), .A1(n1056), .Z(stream_cmd_in_nxt[58]));
Q_AN02 U2701 ( .A0(n30), .A1(stream_cmd_in[58]), .Z(n1056));
Q_MX02 U2702 ( .S(n72), .A0(kme_internal_out[52]), .A1(n1057), .Z(stream_cmd_in_nxt[57]));
Q_AN02 U2703 ( .A0(n30), .A1(stream_cmd_in[57]), .Z(n1057));
Q_MX02 U2704 ( .S(n72), .A0(kme_internal_out[51]), .A1(n1058), .Z(stream_cmd_in_nxt[56]));
Q_AN02 U2705 ( .A0(n30), .A1(stream_cmd_in[56]), .Z(n1058));
Q_MX02 U2706 ( .S(n72), .A0(kme_internal_out[50]), .A1(n1059), .Z(stream_cmd_in_nxt[55]));
Q_AN02 U2707 ( .A0(n30), .A1(stream_cmd_in[55]), .Z(n1059));
Q_MX02 U2708 ( .S(n72), .A0(kme_internal_out[49]), .A1(n1060), .Z(stream_cmd_in_nxt[54]));
Q_AN02 U2709 ( .A0(n30), .A1(stream_cmd_in[54]), .Z(n1060));
Q_MX02 U2710 ( .S(n72), .A0(kme_internal_out[48]), .A1(n1061), .Z(stream_cmd_in_nxt[53]));
Q_AN02 U2711 ( .A0(n30), .A1(stream_cmd_in[53]), .Z(n1061));
Q_MX02 U2712 ( .S(n72), .A0(kme_internal_out[47]), .A1(n1062), .Z(stream_cmd_in_nxt[52]));
Q_AN02 U2713 ( .A0(n30), .A1(stream_cmd_in[52]), .Z(n1062));
Q_MX02 U2714 ( .S(n72), .A0(kme_internal_out[46]), .A1(n1063), .Z(stream_cmd_in_nxt[51]));
Q_AN02 U2715 ( .A0(n30), .A1(stream_cmd_in[51]), .Z(n1063));
Q_MX02 U2716 ( .S(n72), .A0(kme_internal_out[45]), .A1(n1064), .Z(stream_cmd_in_nxt[50]));
Q_AN02 U2717 ( .A0(n30), .A1(stream_cmd_in[50]), .Z(n1064));
Q_MX02 U2718 ( .S(n72), .A0(kme_internal_out[44]), .A1(n1065), .Z(stream_cmd_in_nxt[49]));
Q_AN02 U2719 ( .A0(n30), .A1(stream_cmd_in[49]), .Z(n1065));
Q_MX02 U2720 ( .S(n72), .A0(kme_internal_out[43]), .A1(n1066), .Z(stream_cmd_in_nxt[48]));
Q_AN02 U2721 ( .A0(n30), .A1(stream_cmd_in[48]), .Z(n1066));
Q_MX02 U2722 ( .S(n72), .A0(kme_internal_out[42]), .A1(n1067), .Z(stream_cmd_in_nxt[47]));
Q_AN02 U2723 ( .A0(n30), .A1(stream_cmd_in[47]), .Z(n1067));
Q_MX02 U2724 ( .S(n72), .A0(kme_internal_out[41]), .A1(n1068), .Z(stream_cmd_in_nxt[46]));
Q_AN02 U2725 ( .A0(n30), .A1(stream_cmd_in[46]), .Z(n1068));
Q_MX02 U2726 ( .S(n72), .A0(kme_internal_out[40]), .A1(n1069), .Z(stream_cmd_in_nxt[45]));
Q_AN02 U2727 ( .A0(n30), .A1(stream_cmd_in[45]), .Z(n1069));
Q_MX02 U2728 ( .S(n72), .A0(kme_internal_out[39]), .A1(n1070), .Z(stream_cmd_in_nxt[44]));
Q_AN02 U2729 ( .A0(n30), .A1(stream_cmd_in[44]), .Z(n1070));
Q_MX02 U2730 ( .S(n72), .A0(kme_internal_out[38]), .A1(n1071), .Z(stream_cmd_in_nxt[43]));
Q_AN02 U2731 ( .A0(n30), .A1(stream_cmd_in[43]), .Z(n1071));
Q_MX02 U2732 ( .S(n72), .A0(kme_internal_out[37]), .A1(n1072), .Z(stream_cmd_in_nxt[42]));
Q_AN02 U2733 ( .A0(n30), .A1(stream_cmd_in[42]), .Z(n1072));
Q_MX02 U2734 ( .S(n72), .A0(kme_internal_out[36]), .A1(n1073), .Z(stream_cmd_in_nxt[41]));
Q_AN02 U2735 ( .A0(n30), .A1(stream_cmd_in[41]), .Z(n1073));
Q_MX02 U2736 ( .S(n72), .A0(kme_internal_out[35]), .A1(n1074), .Z(stream_cmd_in_nxt[40]));
Q_AN02 U2737 ( .A0(n30), .A1(stream_cmd_in[40]), .Z(n1074));
Q_MX02 U2738 ( .S(n72), .A0(kme_internal_out[34]), .A1(n1075), .Z(stream_cmd_in_nxt[39]));
Q_AN02 U2739 ( .A0(n30), .A1(stream_cmd_in[39]), .Z(n1075));
Q_MX02 U2740 ( .S(n72), .A0(kme_internal_out[33]), .A1(n1076), .Z(stream_cmd_in_nxt[38]));
Q_AN02 U2741 ( .A0(n30), .A1(stream_cmd_in[38]), .Z(n1076));
Q_MX02 U2742 ( .S(n72), .A0(kme_internal_out[32]), .A1(n1077), .Z(stream_cmd_in_nxt[37]));
Q_AN02 U2743 ( .A0(n30), .A1(stream_cmd_in[37]), .Z(n1077));
Q_MX02 U2744 ( .S(n72), .A0(kme_internal_out[31]), .A1(n1078), .Z(stream_cmd_in_nxt[36]));
Q_AN02 U2745 ( .A0(n30), .A1(stream_cmd_in[36]), .Z(n1078));
Q_MX02 U2746 ( .S(n72), .A0(kme_internal_out[30]), .A1(n1079), .Z(stream_cmd_in_nxt[35]));
Q_AN02 U2747 ( .A0(n30), .A1(stream_cmd_in[35]), .Z(n1079));
Q_MX02 U2748 ( .S(n72), .A0(kme_internal_out[29]), .A1(n1080), .Z(stream_cmd_in_nxt[34]));
Q_AN02 U2749 ( .A0(n30), .A1(stream_cmd_in[34]), .Z(n1080));
Q_MX02 U2750 ( .S(n72), .A0(kme_internal_out[28]), .A1(n1081), .Z(stream_cmd_in_nxt[33]));
Q_AN02 U2751 ( .A0(n30), .A1(stream_cmd_in[33]), .Z(n1081));
Q_MX02 U2752 ( .S(n72), .A0(kme_internal_out[27]), .A1(n1082), .Z(stream_cmd_in_nxt[32]));
Q_AN02 U2753 ( .A0(n30), .A1(stream_cmd_in[32]), .Z(n1082));
Q_MX02 U2754 ( .S(n72), .A0(kme_internal_out[26]), .A1(n1083), .Z(stream_cmd_in_nxt[31]));
Q_AN02 U2755 ( .A0(n30), .A1(stream_cmd_in[31]), .Z(n1083));
Q_MX02 U2756 ( .S(n72), .A0(kme_internal_out[25]), .A1(n1084), .Z(stream_cmd_in_nxt[30]));
Q_AN02 U2757 ( .A0(n30), .A1(stream_cmd_in[30]), .Z(n1084));
Q_MX02 U2758 ( .S(n72), .A0(kme_internal_out[24]), .A1(n1085), .Z(stream_cmd_in_nxt[29]));
Q_AN02 U2759 ( .A0(n30), .A1(stream_cmd_in[29]), .Z(n1085));
Q_MX02 U2760 ( .S(n72), .A0(kme_internal_out[23]), .A1(n1086), .Z(stream_cmd_in_nxt[28]));
Q_AN02 U2761 ( .A0(n30), .A1(stream_cmd_in[28]), .Z(n1086));
Q_MX02 U2762 ( .S(n72), .A0(kme_internal_out[22]), .A1(n1087), .Z(stream_cmd_in_nxt[27]));
Q_AN02 U2763 ( .A0(n30), .A1(stream_cmd_in[27]), .Z(n1087));
Q_MX02 U2764 ( .S(n72), .A0(kme_internal_out[21]), .A1(n1088), .Z(stream_cmd_in_nxt[26]));
Q_AN02 U2765 ( .A0(n30), .A1(stream_cmd_in[26]), .Z(n1088));
Q_MX02 U2766 ( .S(n72), .A0(kme_internal_out[20]), .A1(n1089), .Z(stream_cmd_in_nxt[25]));
Q_AN02 U2767 ( .A0(n30), .A1(stream_cmd_in[25]), .Z(n1089));
Q_MX02 U2768 ( .S(n72), .A0(kme_internal_out[19]), .A1(n1090), .Z(stream_cmd_in_nxt[24]));
Q_AN02 U2769 ( .A0(n30), .A1(stream_cmd_in[24]), .Z(n1090));
Q_MX02 U2770 ( .S(n72), .A0(kme_internal_out[18]), .A1(n1091), .Z(stream_cmd_in_nxt[23]));
Q_AN02 U2771 ( .A0(n30), .A1(stream_cmd_in[23]), .Z(n1091));
Q_MX02 U2772 ( .S(n72), .A0(kme_internal_out[17]), .A1(n1092), .Z(stream_cmd_in_nxt[22]));
Q_AN02 U2773 ( .A0(n30), .A1(stream_cmd_in[22]), .Z(n1092));
Q_MX02 U2774 ( .S(n72), .A0(kme_internal_out[16]), .A1(n1093), .Z(stream_cmd_in_nxt[21]));
Q_AN02 U2775 ( .A0(n30), .A1(stream_cmd_in[21]), .Z(n1093));
Q_MX02 U2776 ( .S(n72), .A0(kme_internal_out[15]), .A1(n1094), .Z(stream_cmd_in_nxt[20]));
Q_AN02 U2777 ( .A0(n30), .A1(stream_cmd_in[20]), .Z(n1094));
Q_MX02 U2778 ( .S(n72), .A0(kme_internal_out[14]), .A1(n1095), .Z(stream_cmd_in_nxt[19]));
Q_AN02 U2779 ( .A0(n30), .A1(stream_cmd_in[19]), .Z(n1095));
Q_MX02 U2780 ( .S(n72), .A0(kme_internal_out[13]), .A1(n1096), .Z(stream_cmd_in_nxt[18]));
Q_AN02 U2781 ( .A0(n30), .A1(stream_cmd_in[18]), .Z(n1096));
Q_MX02 U2782 ( .S(n72), .A0(kme_internal_out[12]), .A1(n1097), .Z(stream_cmd_in_nxt[17]));
Q_AN02 U2783 ( .A0(n30), .A1(stream_cmd_in[17]), .Z(n1097));
Q_MX02 U2784 ( .S(n72), .A0(kme_internal_out[11]), .A1(n1098), .Z(stream_cmd_in_nxt[16]));
Q_AN02 U2785 ( .A0(n30), .A1(stream_cmd_in[16]), .Z(n1098));
Q_MX02 U2786 ( .S(n72), .A0(kme_internal_out[10]), .A1(n1099), .Z(stream_cmd_in_nxt[15]));
Q_AN02 U2787 ( .A0(n30), .A1(stream_cmd_in[15]), .Z(n1099));
Q_MX02 U2788 ( .S(n72), .A0(kme_internal_out[9]), .A1(n1100), .Z(stream_cmd_in_nxt[14]));
Q_AN02 U2789 ( .A0(n30), .A1(stream_cmd_in[14]), .Z(n1100));
Q_MX02 U2790 ( .S(n72), .A0(kme_internal_out[8]), .A1(n1101), .Z(stream_cmd_in_nxt[13]));
Q_AN02 U2791 ( .A0(n30), .A1(stream_cmd_in[13]), .Z(n1101));
Q_MX02 U2792 ( .S(n72), .A0(kme_internal_out[7]), .A1(n1102), .Z(stream_cmd_in_nxt[12]));
Q_AN02 U2793 ( .A0(n30), .A1(stream_cmd_in[12]), .Z(n1102));
Q_MX02 U2794 ( .S(n72), .A0(kme_internal_out[6]), .A1(n1103), .Z(stream_cmd_in_nxt[11]));
Q_AN02 U2795 ( .A0(n30), .A1(stream_cmd_in[11]), .Z(n1103));
Q_MX02 U2796 ( .S(n72), .A0(kme_internal_out[5]), .A1(n1104), .Z(stream_cmd_in_nxt[10]));
Q_AN02 U2797 ( .A0(n30), .A1(stream_cmd_in[10]), .Z(n1104));
Q_MX02 U2798 ( .S(n72), .A0(kme_internal_out[4]), .A1(n1105), .Z(stream_cmd_in_nxt[9]));
Q_AN02 U2799 ( .A0(n30), .A1(stream_cmd_in[9]), .Z(n1105));
Q_MX02 U2800 ( .S(n72), .A0(kme_internal_out[3]), .A1(n1106), .Z(stream_cmd_in_nxt[8]));
Q_AN02 U2801 ( .A0(n30), .A1(stream_cmd_in[8]), .Z(n1106));
Q_MX02 U2802 ( .S(n72), .A0(kme_internal_out[2]), .A1(n1107), .Z(stream_cmd_in_nxt[7]));
Q_AN02 U2803 ( .A0(n30), .A1(stream_cmd_in[7]), .Z(n1107));
Q_MX02 U2804 ( .S(n72), .A0(kme_internal_out[1]), .A1(n1108), .Z(stream_cmd_in_nxt[6]));
Q_AN02 U2805 ( .A0(n30), .A1(stream_cmd_in[6]), .Z(n1108));
Q_MX02 U2806 ( .S(n72), .A0(kme_internal_out[0]), .A1(n1109), .Z(stream_cmd_in_nxt[5]));
Q_AN02 U2807 ( .A0(n30), .A1(stream_cmd_in[5]), .Z(n1109));
Q_AN02 U2808 ( .A0(n31), .A1(stream_cmd_in[4]), .Z(stream_cmd_in_nxt[4]));
Q_AN02 U2809 ( .A0(n31), .A1(stream_cmd_in[3]), .Z(stream_cmd_in_nxt[3]));
Q_AN02 U2810 ( .A0(n31), .A1(stream_cmd_in[2]), .Z(stream_cmd_in_nxt[2]));
Q_MX02 U2811 ( .S(keyfilter_cmd_in_valid), .A0(skip_dek_kdf), .A1(n2718), .Z(skip_dek_kdf_nxt));
Q_MX02 U2812 ( .S(keyfilter_cmd_in_valid), .A0(skip_dak_kdf), .A1(n2717), .Z(skip_dak_kdf_nxt));
Q_MX02 U2813 ( .S(n35), .A0(kme_internal_out[48]), .A1(kdf_dek_iter), .Z(kdf_dek_iter_nxt));
Q_MX02 U2814 ( .S(n32), .A0(gcm_dak_tag[31]), .A1(n2333), .Z(gcm_dak_tag_nxt[31]));
Q_MX02 U2815 ( .S(n32), .A0(gcm_dak_tag[30]), .A1(n2334), .Z(gcm_dak_tag_nxt[30]));
Q_MX02 U2816 ( .S(n32), .A0(gcm_dak_tag[29]), .A1(n2335), .Z(gcm_dak_tag_nxt[29]));
Q_MX02 U2817 ( .S(n32), .A0(gcm_dak_tag[28]), .A1(n2336), .Z(gcm_dak_tag_nxt[28]));
Q_MX02 U2818 ( .S(n32), .A0(gcm_dak_tag[27]), .A1(n2337), .Z(gcm_dak_tag_nxt[27]));
Q_MX02 U2819 ( .S(n32), .A0(gcm_dak_tag[26]), .A1(n2338), .Z(gcm_dak_tag_nxt[26]));
Q_MX02 U2820 ( .S(n32), .A0(gcm_dak_tag[25]), .A1(n2339), .Z(gcm_dak_tag_nxt[25]));
Q_MX02 U2821 ( .S(n32), .A0(gcm_dak_tag[24]), .A1(n2340), .Z(gcm_dak_tag_nxt[24]));
Q_MX02 U2822 ( .S(n32), .A0(gcm_dak_tag[23]), .A1(n2341), .Z(gcm_dak_tag_nxt[23]));
Q_MX02 U2823 ( .S(n32), .A0(gcm_dak_tag[22]), .A1(n2342), .Z(gcm_dak_tag_nxt[22]));
Q_MX02 U2824 ( .S(n32), .A0(gcm_dak_tag[21]), .A1(n2343), .Z(gcm_dak_tag_nxt[21]));
Q_MX02 U2825 ( .S(n32), .A0(gcm_dak_tag[20]), .A1(n2344), .Z(gcm_dak_tag_nxt[20]));
Q_MX02 U2826 ( .S(n32), .A0(gcm_dak_tag[19]), .A1(n2345), .Z(gcm_dak_tag_nxt[19]));
Q_MX02 U2827 ( .S(n32), .A0(gcm_dak_tag[18]), .A1(n2346), .Z(gcm_dak_tag_nxt[18]));
Q_MX02 U2828 ( .S(n32), .A0(gcm_dak_tag[17]), .A1(n2347), .Z(gcm_dak_tag_nxt[17]));
Q_MX02 U2829 ( .S(n32), .A0(gcm_dak_tag[16]), .A1(n2348), .Z(gcm_dak_tag_nxt[16]));
Q_MX02 U2830 ( .S(n32), .A0(gcm_dak_tag[15]), .A1(n2349), .Z(gcm_dak_tag_nxt[15]));
Q_MX02 U2831 ( .S(n32), .A0(gcm_dak_tag[14]), .A1(n2350), .Z(gcm_dak_tag_nxt[14]));
Q_MX02 U2832 ( .S(n32), .A0(gcm_dak_tag[13]), .A1(n2351), .Z(gcm_dak_tag_nxt[13]));
Q_MX02 U2833 ( .S(n32), .A0(gcm_dak_tag[12]), .A1(n2352), .Z(gcm_dak_tag_nxt[12]));
Q_MX02 U2834 ( .S(n32), .A0(gcm_dak_tag[11]), .A1(n2353), .Z(gcm_dak_tag_nxt[11]));
Q_MX02 U2835 ( .S(n32), .A0(gcm_dak_tag[10]), .A1(n2354), .Z(gcm_dak_tag_nxt[10]));
Q_MX02 U2836 ( .S(n32), .A0(gcm_dak_tag[9]), .A1(n2355), .Z(gcm_dak_tag_nxt[9]));
Q_MX02 U2837 ( .S(n32), .A0(gcm_dak_tag[8]), .A1(n2356), .Z(gcm_dak_tag_nxt[8]));
Q_MX02 U2838 ( .S(n32), .A0(gcm_dak_tag[7]), .A1(n2357), .Z(gcm_dak_tag_nxt[7]));
Q_MX02 U2839 ( .S(n32), .A0(gcm_dak_tag[6]), .A1(n2358), .Z(gcm_dak_tag_nxt[6]));
Q_MX02 U2840 ( .S(n32), .A0(gcm_dak_tag[5]), .A1(n2359), .Z(gcm_dak_tag_nxt[5]));
Q_MX02 U2841 ( .S(n32), .A0(gcm_dak_tag[4]), .A1(n2360), .Z(gcm_dak_tag_nxt[4]));
Q_MX02 U2842 ( .S(n32), .A0(gcm_dak_tag[3]), .A1(n2361), .Z(gcm_dak_tag_nxt[3]));
Q_MX02 U2843 ( .S(n32), .A0(gcm_dak_tag[2]), .A1(n2362), .Z(gcm_dak_tag_nxt[2]));
Q_MX02 U2844 ( .S(n32), .A0(gcm_dak_tag[1]), .A1(n2363), .Z(gcm_dak_tag_nxt[1]));
Q_MX02 U2845 ( .S(n32), .A0(gcm_dak_tag[0]), .A1(n2364), .Z(gcm_dak_tag_nxt[0]));
Q_MX02 U2846 ( .S(n32), .A0(gcm_dak_tag[95]), .A1(n2365), .Z(gcm_dak_tag_nxt[95]));
Q_MX02 U2847 ( .S(n32), .A0(gcm_dak_tag[94]), .A1(n2366), .Z(gcm_dak_tag_nxt[94]));
Q_MX02 U2848 ( .S(n32), .A0(gcm_dak_tag[93]), .A1(n2367), .Z(gcm_dak_tag_nxt[93]));
Q_MX02 U2849 ( .S(n32), .A0(gcm_dak_tag[92]), .A1(n2368), .Z(gcm_dak_tag_nxt[92]));
Q_MX02 U2850 ( .S(n32), .A0(gcm_dak_tag[91]), .A1(n2369), .Z(gcm_dak_tag_nxt[91]));
Q_MX02 U2851 ( .S(n32), .A0(gcm_dak_tag[90]), .A1(n2370), .Z(gcm_dak_tag_nxt[90]));
Q_MX02 U2852 ( .S(n32), .A0(gcm_dak_tag[89]), .A1(n2371), .Z(gcm_dak_tag_nxt[89]));
Q_MX02 U2853 ( .S(n32), .A0(gcm_dak_tag[88]), .A1(n2372), .Z(gcm_dak_tag_nxt[88]));
Q_MX02 U2854 ( .S(n32), .A0(gcm_dak_tag[87]), .A1(n2373), .Z(gcm_dak_tag_nxt[87]));
Q_MX02 U2855 ( .S(n32), .A0(gcm_dak_tag[86]), .A1(n2374), .Z(gcm_dak_tag_nxt[86]));
Q_MX02 U2856 ( .S(n32), .A0(gcm_dak_tag[85]), .A1(n2375), .Z(gcm_dak_tag_nxt[85]));
Q_MX02 U2857 ( .S(n32), .A0(gcm_dak_tag[84]), .A1(n2376), .Z(gcm_dak_tag_nxt[84]));
Q_MX02 U2858 ( .S(n32), .A0(gcm_dak_tag[83]), .A1(n2377), .Z(gcm_dak_tag_nxt[83]));
Q_MX02 U2859 ( .S(n32), .A0(gcm_dak_tag[82]), .A1(n2378), .Z(gcm_dak_tag_nxt[82]));
Q_MX02 U2860 ( .S(n32), .A0(gcm_dak_tag[81]), .A1(n2379), .Z(gcm_dak_tag_nxt[81]));
Q_MX02 U2861 ( .S(n32), .A0(gcm_dak_tag[80]), .A1(n2380), .Z(gcm_dak_tag_nxt[80]));
Q_MX02 U2862 ( .S(n32), .A0(gcm_dak_tag[79]), .A1(n2381), .Z(gcm_dak_tag_nxt[79]));
Q_MX02 U2863 ( .S(n32), .A0(gcm_dak_tag[78]), .A1(n2382), .Z(gcm_dak_tag_nxt[78]));
Q_MX02 U2864 ( .S(n32), .A0(gcm_dak_tag[77]), .A1(n2383), .Z(gcm_dak_tag_nxt[77]));
Q_MX02 U2865 ( .S(n32), .A0(gcm_dak_tag[76]), .A1(n2384), .Z(gcm_dak_tag_nxt[76]));
Q_MX02 U2866 ( .S(n32), .A0(gcm_dak_tag[75]), .A1(n2385), .Z(gcm_dak_tag_nxt[75]));
Q_MX02 U2867 ( .S(n32), .A0(gcm_dak_tag[74]), .A1(n2386), .Z(gcm_dak_tag_nxt[74]));
Q_MX02 U2868 ( .S(n32), .A0(gcm_dak_tag[73]), .A1(n2387), .Z(gcm_dak_tag_nxt[73]));
Q_MX02 U2869 ( .S(n32), .A0(gcm_dak_tag[72]), .A1(n2388), .Z(gcm_dak_tag_nxt[72]));
Q_MX02 U2870 ( .S(n32), .A0(gcm_dak_tag[71]), .A1(n2389), .Z(gcm_dak_tag_nxt[71]));
Q_MX02 U2871 ( .S(n32), .A0(gcm_dak_tag[70]), .A1(n2390), .Z(gcm_dak_tag_nxt[70]));
Q_MX02 U2872 ( .S(n32), .A0(gcm_dak_tag[69]), .A1(n2391), .Z(gcm_dak_tag_nxt[69]));
Q_MX02 U2873 ( .S(n32), .A0(gcm_dak_tag[68]), .A1(n2392), .Z(gcm_dak_tag_nxt[68]));
Q_MX02 U2874 ( .S(n32), .A0(gcm_dak_tag[67]), .A1(n2393), .Z(gcm_dak_tag_nxt[67]));
Q_MX02 U2875 ( .S(n32), .A0(gcm_dak_tag[66]), .A1(n2394), .Z(gcm_dak_tag_nxt[66]));
Q_MX02 U2876 ( .S(n32), .A0(gcm_dak_tag[65]), .A1(n2395), .Z(gcm_dak_tag_nxt[65]));
Q_MX02 U2877 ( .S(n32), .A0(gcm_dak_tag[64]), .A1(n2396), .Z(gcm_dak_tag_nxt[64]));
Q_MX02 U2878 ( .S(n32), .A0(gcm_dak_tag[63]), .A1(n2397), .Z(gcm_dak_tag_nxt[63]));
Q_MX02 U2879 ( .S(n32), .A0(gcm_dak_tag[62]), .A1(n2398), .Z(gcm_dak_tag_nxt[62]));
Q_MX02 U2880 ( .S(n32), .A0(gcm_dak_tag[61]), .A1(n2399), .Z(gcm_dak_tag_nxt[61]));
Q_MX02 U2881 ( .S(n32), .A0(gcm_dak_tag[60]), .A1(n2400), .Z(gcm_dak_tag_nxt[60]));
Q_MX02 U2882 ( .S(n32), .A0(gcm_dak_tag[59]), .A1(n2401), .Z(gcm_dak_tag_nxt[59]));
Q_MX02 U2883 ( .S(n32), .A0(gcm_dak_tag[58]), .A1(n2402), .Z(gcm_dak_tag_nxt[58]));
Q_MX02 U2884 ( .S(n32), .A0(gcm_dak_tag[57]), .A1(n2403), .Z(gcm_dak_tag_nxt[57]));
Q_MX02 U2885 ( .S(n32), .A0(gcm_dak_tag[56]), .A1(n2404), .Z(gcm_dak_tag_nxt[56]));
Q_MX02 U2886 ( .S(n32), .A0(gcm_dak_tag[55]), .A1(n2405), .Z(gcm_dak_tag_nxt[55]));
Q_MX02 U2887 ( .S(n32), .A0(gcm_dak_tag[54]), .A1(n2406), .Z(gcm_dak_tag_nxt[54]));
Q_MX02 U2888 ( .S(n32), .A0(gcm_dak_tag[53]), .A1(n2407), .Z(gcm_dak_tag_nxt[53]));
Q_MX02 U2889 ( .S(n32), .A0(gcm_dak_tag[52]), .A1(n2408), .Z(gcm_dak_tag_nxt[52]));
Q_MX02 U2890 ( .S(n32), .A0(gcm_dak_tag[51]), .A1(n2409), .Z(gcm_dak_tag_nxt[51]));
Q_MX02 U2891 ( .S(n32), .A0(gcm_dak_tag[50]), .A1(n2410), .Z(gcm_dak_tag_nxt[50]));
Q_MX02 U2892 ( .S(n32), .A0(gcm_dak_tag[49]), .A1(n2411), .Z(gcm_dak_tag_nxt[49]));
Q_MX02 U2893 ( .S(n32), .A0(gcm_dak_tag[48]), .A1(n2412), .Z(gcm_dak_tag_nxt[48]));
Q_MX02 U2894 ( .S(n32), .A0(gcm_dak_tag[47]), .A1(n2413), .Z(gcm_dak_tag_nxt[47]));
Q_MX02 U2895 ( .S(n32), .A0(gcm_dak_tag[46]), .A1(n2414), .Z(gcm_dak_tag_nxt[46]));
Q_MX02 U2896 ( .S(n32), .A0(gcm_dak_tag[45]), .A1(n2415), .Z(gcm_dak_tag_nxt[45]));
Q_MX02 U2897 ( .S(n32), .A0(gcm_dak_tag[44]), .A1(n2416), .Z(gcm_dak_tag_nxt[44]));
Q_MX02 U2898 ( .S(n32), .A0(gcm_dak_tag[43]), .A1(n2417), .Z(gcm_dak_tag_nxt[43]));
Q_MX02 U2899 ( .S(n32), .A0(gcm_dak_tag[42]), .A1(n2418), .Z(gcm_dak_tag_nxt[42]));
Q_MX02 U2900 ( .S(n32), .A0(gcm_dak_tag[41]), .A1(n2419), .Z(gcm_dak_tag_nxt[41]));
Q_MX02 U2901 ( .S(n32), .A0(gcm_dak_tag[40]), .A1(n2420), .Z(gcm_dak_tag_nxt[40]));
Q_MX02 U2902 ( .S(n32), .A0(gcm_dak_tag[39]), .A1(n2421), .Z(gcm_dak_tag_nxt[39]));
Q_MX02 U2903 ( .S(n32), .A0(gcm_dak_tag[38]), .A1(n2422), .Z(gcm_dak_tag_nxt[38]));
Q_MX02 U2904 ( .S(n32), .A0(gcm_dak_tag[37]), .A1(n2423), .Z(gcm_dak_tag_nxt[37]));
Q_MX02 U2905 ( .S(n32), .A0(gcm_dak_tag[36]), .A1(n2424), .Z(gcm_dak_tag_nxt[36]));
Q_MX02 U2906 ( .S(n32), .A0(gcm_dak_tag[35]), .A1(n2425), .Z(gcm_dak_tag_nxt[35]));
Q_MX02 U2907 ( .S(n32), .A0(gcm_dak_tag[34]), .A1(n2426), .Z(gcm_dak_tag_nxt[34]));
Q_MX02 U2908 ( .S(n32), .A0(gcm_dak_tag[33]), .A1(n2427), .Z(gcm_dak_tag_nxt[33]));
Q_MX02 U2909 ( .S(n32), .A0(gcm_dak_tag[32]), .A1(n2428), .Z(gcm_dak_tag_nxt[32]));
Q_MX02 U2910 ( .S(n33), .A0(gcm_dek_tag[31]), .A1(n2429), .Z(gcm_dek_tag_nxt[31]));
Q_MX02 U2911 ( .S(n33), .A0(gcm_dek_tag[30]), .A1(n2430), .Z(gcm_dek_tag_nxt[30]));
Q_MX02 U2912 ( .S(n33), .A0(gcm_dek_tag[29]), .A1(n2431), .Z(gcm_dek_tag_nxt[29]));
Q_MX02 U2913 ( .S(n33), .A0(gcm_dek_tag[28]), .A1(n2432), .Z(gcm_dek_tag_nxt[28]));
Q_MX02 U2914 ( .S(n33), .A0(gcm_dek_tag[27]), .A1(n2433), .Z(gcm_dek_tag_nxt[27]));
Q_MX02 U2915 ( .S(n33), .A0(gcm_dek_tag[26]), .A1(n2434), .Z(gcm_dek_tag_nxt[26]));
Q_MX02 U2916 ( .S(n33), .A0(gcm_dek_tag[25]), .A1(n2435), .Z(gcm_dek_tag_nxt[25]));
Q_MX02 U2917 ( .S(n33), .A0(gcm_dek_tag[24]), .A1(n2436), .Z(gcm_dek_tag_nxt[24]));
Q_MX02 U2918 ( .S(n33), .A0(gcm_dek_tag[23]), .A1(n2437), .Z(gcm_dek_tag_nxt[23]));
Q_MX02 U2919 ( .S(n33), .A0(gcm_dek_tag[22]), .A1(n2438), .Z(gcm_dek_tag_nxt[22]));
Q_MX02 U2920 ( .S(n33), .A0(gcm_dek_tag[21]), .A1(n2439), .Z(gcm_dek_tag_nxt[21]));
Q_MX02 U2921 ( .S(n33), .A0(gcm_dek_tag[20]), .A1(n2440), .Z(gcm_dek_tag_nxt[20]));
Q_MX02 U2922 ( .S(n33), .A0(gcm_dek_tag[19]), .A1(n2441), .Z(gcm_dek_tag_nxt[19]));
Q_MX02 U2923 ( .S(n33), .A0(gcm_dek_tag[18]), .A1(n2442), .Z(gcm_dek_tag_nxt[18]));
Q_MX02 U2924 ( .S(n33), .A0(gcm_dek_tag[17]), .A1(n2443), .Z(gcm_dek_tag_nxt[17]));
Q_MX02 U2925 ( .S(n33), .A0(gcm_dek_tag[16]), .A1(n2444), .Z(gcm_dek_tag_nxt[16]));
Q_MX02 U2926 ( .S(n33), .A0(gcm_dek_tag[15]), .A1(n2445), .Z(gcm_dek_tag_nxt[15]));
Q_MX02 U2927 ( .S(n33), .A0(gcm_dek_tag[14]), .A1(n2446), .Z(gcm_dek_tag_nxt[14]));
Q_MX02 U2928 ( .S(n33), .A0(gcm_dek_tag[13]), .A1(n2447), .Z(gcm_dek_tag_nxt[13]));
Q_MX02 U2929 ( .S(n33), .A0(gcm_dek_tag[12]), .A1(n2448), .Z(gcm_dek_tag_nxt[12]));
Q_MX02 U2930 ( .S(n33), .A0(gcm_dek_tag[11]), .A1(n2449), .Z(gcm_dek_tag_nxt[11]));
Q_MX02 U2931 ( .S(n33), .A0(gcm_dek_tag[10]), .A1(n2450), .Z(gcm_dek_tag_nxt[10]));
Q_MX02 U2932 ( .S(n33), .A0(gcm_dek_tag[9]), .A1(n2451), .Z(gcm_dek_tag_nxt[9]));
Q_MX02 U2933 ( .S(n33), .A0(gcm_dek_tag[8]), .A1(n2452), .Z(gcm_dek_tag_nxt[8]));
Q_MX02 U2934 ( .S(n33), .A0(gcm_dek_tag[7]), .A1(n2453), .Z(gcm_dek_tag_nxt[7]));
Q_MX02 U2935 ( .S(n33), .A0(gcm_dek_tag[6]), .A1(n2454), .Z(gcm_dek_tag_nxt[6]));
Q_MX02 U2936 ( .S(n33), .A0(gcm_dek_tag[5]), .A1(n2455), .Z(gcm_dek_tag_nxt[5]));
Q_MX02 U2937 ( .S(n33), .A0(gcm_dek_tag[4]), .A1(n2456), .Z(gcm_dek_tag_nxt[4]));
Q_MX02 U2938 ( .S(n33), .A0(gcm_dek_tag[3]), .A1(n2457), .Z(gcm_dek_tag_nxt[3]));
Q_MX02 U2939 ( .S(n33), .A0(gcm_dek_tag[2]), .A1(n2458), .Z(gcm_dek_tag_nxt[2]));
Q_MX02 U2940 ( .S(n33), .A0(gcm_dek_tag[1]), .A1(n2459), .Z(gcm_dek_tag_nxt[1]));
Q_MX02 U2941 ( .S(n33), .A0(gcm_dek_tag[0]), .A1(n2460), .Z(gcm_dek_tag_nxt[0]));
Q_MX02 U2942 ( .S(n33), .A0(gcm_dek_tag[95]), .A1(n2461), .Z(gcm_dek_tag_nxt[95]));
Q_MX02 U2943 ( .S(n33), .A0(gcm_dek_tag[94]), .A1(n2462), .Z(gcm_dek_tag_nxt[94]));
Q_MX02 U2944 ( .S(n33), .A0(gcm_dek_tag[93]), .A1(n2463), .Z(gcm_dek_tag_nxt[93]));
Q_MX02 U2945 ( .S(n33), .A0(gcm_dek_tag[92]), .A1(n2464), .Z(gcm_dek_tag_nxt[92]));
Q_MX02 U2946 ( .S(n33), .A0(gcm_dek_tag[91]), .A1(n2465), .Z(gcm_dek_tag_nxt[91]));
Q_MX02 U2947 ( .S(n33), .A0(gcm_dek_tag[90]), .A1(n2466), .Z(gcm_dek_tag_nxt[90]));
Q_MX02 U2948 ( .S(n33), .A0(gcm_dek_tag[89]), .A1(n2467), .Z(gcm_dek_tag_nxt[89]));
Q_MX02 U2949 ( .S(n33), .A0(gcm_dek_tag[88]), .A1(n2468), .Z(gcm_dek_tag_nxt[88]));
Q_MX02 U2950 ( .S(n33), .A0(gcm_dek_tag[87]), .A1(n2469), .Z(gcm_dek_tag_nxt[87]));
Q_MX02 U2951 ( .S(n33), .A0(gcm_dek_tag[86]), .A1(n2470), .Z(gcm_dek_tag_nxt[86]));
Q_MX02 U2952 ( .S(n33), .A0(gcm_dek_tag[85]), .A1(n2471), .Z(gcm_dek_tag_nxt[85]));
Q_MX02 U2953 ( .S(n33), .A0(gcm_dek_tag[84]), .A1(n2472), .Z(gcm_dek_tag_nxt[84]));
Q_MX02 U2954 ( .S(n33), .A0(gcm_dek_tag[83]), .A1(n2473), .Z(gcm_dek_tag_nxt[83]));
Q_MX02 U2955 ( .S(n33), .A0(gcm_dek_tag[82]), .A1(n2474), .Z(gcm_dek_tag_nxt[82]));
Q_MX02 U2956 ( .S(n33), .A0(gcm_dek_tag[81]), .A1(n2475), .Z(gcm_dek_tag_nxt[81]));
Q_MX02 U2957 ( .S(n33), .A0(gcm_dek_tag[80]), .A1(n2476), .Z(gcm_dek_tag_nxt[80]));
Q_MX02 U2958 ( .S(n33), .A0(gcm_dek_tag[79]), .A1(n2477), .Z(gcm_dek_tag_nxt[79]));
Q_MX02 U2959 ( .S(n33), .A0(gcm_dek_tag[78]), .A1(n2478), .Z(gcm_dek_tag_nxt[78]));
Q_MX02 U2960 ( .S(n33), .A0(gcm_dek_tag[77]), .A1(n2479), .Z(gcm_dek_tag_nxt[77]));
Q_MX02 U2961 ( .S(n33), .A0(gcm_dek_tag[76]), .A1(n2480), .Z(gcm_dek_tag_nxt[76]));
Q_MX02 U2962 ( .S(n33), .A0(gcm_dek_tag[75]), .A1(n2481), .Z(gcm_dek_tag_nxt[75]));
Q_MX02 U2963 ( .S(n33), .A0(gcm_dek_tag[74]), .A1(n2482), .Z(gcm_dek_tag_nxt[74]));
Q_MX02 U2964 ( .S(n33), .A0(gcm_dek_tag[73]), .A1(n2483), .Z(gcm_dek_tag_nxt[73]));
Q_MX02 U2965 ( .S(n33), .A0(gcm_dek_tag[72]), .A1(n2484), .Z(gcm_dek_tag_nxt[72]));
Q_MX02 U2966 ( .S(n33), .A0(gcm_dek_tag[71]), .A1(n2485), .Z(gcm_dek_tag_nxt[71]));
Q_MX02 U2967 ( .S(n33), .A0(gcm_dek_tag[70]), .A1(n2486), .Z(gcm_dek_tag_nxt[70]));
Q_MX02 U2968 ( .S(n33), .A0(gcm_dek_tag[69]), .A1(n2487), .Z(gcm_dek_tag_nxt[69]));
Q_MX02 U2969 ( .S(n33), .A0(gcm_dek_tag[68]), .A1(n2488), .Z(gcm_dek_tag_nxt[68]));
Q_MX02 U2970 ( .S(n33), .A0(gcm_dek_tag[67]), .A1(n2489), .Z(gcm_dek_tag_nxt[67]));
Q_MX02 U2971 ( .S(n33), .A0(gcm_dek_tag[66]), .A1(n2490), .Z(gcm_dek_tag_nxt[66]));
Q_MX02 U2972 ( .S(n33), .A0(gcm_dek_tag[65]), .A1(n2491), .Z(gcm_dek_tag_nxt[65]));
Q_MX02 U2973 ( .S(n33), .A0(gcm_dek_tag[64]), .A1(n2492), .Z(gcm_dek_tag_nxt[64]));
Q_MX02 U2974 ( .S(n33), .A0(gcm_dek_tag[63]), .A1(n2493), .Z(gcm_dek_tag_nxt[63]));
Q_MX02 U2975 ( .S(n33), .A0(gcm_dek_tag[62]), .A1(n2494), .Z(gcm_dek_tag_nxt[62]));
Q_MX02 U2976 ( .S(n33), .A0(gcm_dek_tag[61]), .A1(n2495), .Z(gcm_dek_tag_nxt[61]));
Q_MX02 U2977 ( .S(n33), .A0(gcm_dek_tag[60]), .A1(n2496), .Z(gcm_dek_tag_nxt[60]));
Q_MX02 U2978 ( .S(n33), .A0(gcm_dek_tag[59]), .A1(n2497), .Z(gcm_dek_tag_nxt[59]));
Q_MX02 U2979 ( .S(n33), .A0(gcm_dek_tag[58]), .A1(n2498), .Z(gcm_dek_tag_nxt[58]));
Q_MX02 U2980 ( .S(n33), .A0(gcm_dek_tag[57]), .A1(n2499), .Z(gcm_dek_tag_nxt[57]));
Q_MX02 U2981 ( .S(n33), .A0(gcm_dek_tag[56]), .A1(n2500), .Z(gcm_dek_tag_nxt[56]));
Q_MX02 U2982 ( .S(n33), .A0(gcm_dek_tag[55]), .A1(n2501), .Z(gcm_dek_tag_nxt[55]));
Q_MX02 U2983 ( .S(n33), .A0(gcm_dek_tag[54]), .A1(n2502), .Z(gcm_dek_tag_nxt[54]));
Q_MX02 U2984 ( .S(n33), .A0(gcm_dek_tag[53]), .A1(n2503), .Z(gcm_dek_tag_nxt[53]));
Q_MX02 U2985 ( .S(n33), .A0(gcm_dek_tag[52]), .A1(n2504), .Z(gcm_dek_tag_nxt[52]));
Q_MX02 U2986 ( .S(n33), .A0(gcm_dek_tag[51]), .A1(n2505), .Z(gcm_dek_tag_nxt[51]));
Q_MX02 U2987 ( .S(n33), .A0(gcm_dek_tag[50]), .A1(n2506), .Z(gcm_dek_tag_nxt[50]));
Q_MX02 U2988 ( .S(n33), .A0(gcm_dek_tag[49]), .A1(n2507), .Z(gcm_dek_tag_nxt[49]));
Q_MX02 U2989 ( .S(n33), .A0(gcm_dek_tag[48]), .A1(n2508), .Z(gcm_dek_tag_nxt[48]));
Q_MX02 U2990 ( .S(n33), .A0(gcm_dek_tag[47]), .A1(n2509), .Z(gcm_dek_tag_nxt[47]));
Q_MX02 U2991 ( .S(n33), .A0(gcm_dek_tag[46]), .A1(n2510), .Z(gcm_dek_tag_nxt[46]));
Q_MX02 U2992 ( .S(n33), .A0(gcm_dek_tag[45]), .A1(n2511), .Z(gcm_dek_tag_nxt[45]));
Q_MX02 U2993 ( .S(n33), .A0(gcm_dek_tag[44]), .A1(n2512), .Z(gcm_dek_tag_nxt[44]));
Q_MX02 U2994 ( .S(n33), .A0(gcm_dek_tag[43]), .A1(n2513), .Z(gcm_dek_tag_nxt[43]));
Q_MX02 U2995 ( .S(n33), .A0(gcm_dek_tag[42]), .A1(n2514), .Z(gcm_dek_tag_nxt[42]));
Q_MX02 U2996 ( .S(n33), .A0(gcm_dek_tag[41]), .A1(n2515), .Z(gcm_dek_tag_nxt[41]));
Q_MX02 U2997 ( .S(n33), .A0(gcm_dek_tag[40]), .A1(n2516), .Z(gcm_dek_tag_nxt[40]));
Q_MX02 U2998 ( .S(n33), .A0(gcm_dek_tag[39]), .A1(n2517), .Z(gcm_dek_tag_nxt[39]));
Q_MX02 U2999 ( .S(n33), .A0(gcm_dek_tag[38]), .A1(n2518), .Z(gcm_dek_tag_nxt[38]));
Q_MX02 U3000 ( .S(n33), .A0(gcm_dek_tag[37]), .A1(n2519), .Z(gcm_dek_tag_nxt[37]));
Q_MX02 U3001 ( .S(n33), .A0(gcm_dek_tag[36]), .A1(n2520), .Z(gcm_dek_tag_nxt[36]));
Q_MX02 U3002 ( .S(n33), .A0(gcm_dek_tag[35]), .A1(n2521), .Z(gcm_dek_tag_nxt[35]));
Q_MX02 U3003 ( .S(n33), .A0(gcm_dek_tag[34]), .A1(n2522), .Z(gcm_dek_tag_nxt[34]));
Q_MX02 U3004 ( .S(n33), .A0(gcm_dek_tag[33]), .A1(n2523), .Z(gcm_dek_tag_nxt[33]));
Q_MX02 U3005 ( .S(n33), .A0(gcm_dek_tag[32]), .A1(n2524), .Z(gcm_dek_tag_nxt[32]));
Q_AO21 U3006 ( .A0(n35), .A1(gcm_dak_cmd_in[0]), .B0(n34), .Z(gcm_dak_cmd_in_nxt[0]));
Q_AO21 U3007 ( .A0(n35), .A1(gcm_dak_cmd_in[1]), .B0(n1111), .Z(gcm_dak_cmd_in_nxt[1]));
Q_AO21 U3008 ( .A0(n35), .A1(gcm_dak_cmd_in[2]), .B0(n1110), .Z(gcm_dak_cmd_in_nxt[2]));
Q_XNR2 U3009 ( .A0(n77), .A1(n82), .Z(n1110));
Q_NR02 U3010 ( .A0(n77), .A1(n82), .Z(n1111));
Q_AN02 U3011 ( .A0(n35), .A1(n1112), .Z(gcm_dak_cmd_in_nxt[34]));
Q_MX02 U3012 ( .S(n86), .A0(n2525), .A1(gcm_dak_cmd_in[34]), .Z(n1112));
Q_AN02 U3013 ( .A0(n35), .A1(n1113), .Z(gcm_dak_cmd_in_nxt[33]));
Q_MX02 U3014 ( .S(n86), .A0(n2526), .A1(gcm_dak_cmd_in[33]), .Z(n1113));
Q_AN02 U3015 ( .A0(n35), .A1(n1114), .Z(gcm_dak_cmd_in_nxt[32]));
Q_MX02 U3016 ( .S(n86), .A0(n2527), .A1(gcm_dak_cmd_in[32]), .Z(n1114));
Q_AN02 U3017 ( .A0(n35), .A1(n1115), .Z(gcm_dak_cmd_in_nxt[31]));
Q_MX02 U3018 ( .S(n86), .A0(n2528), .A1(gcm_dak_cmd_in[31]), .Z(n1115));
Q_AN02 U3019 ( .A0(n35), .A1(n1116), .Z(gcm_dak_cmd_in_nxt[30]));
Q_MX02 U3020 ( .S(n86), .A0(n2529), .A1(gcm_dak_cmd_in[30]), .Z(n1116));
Q_AN02 U3021 ( .A0(n35), .A1(n1117), .Z(gcm_dak_cmd_in_nxt[29]));
Q_MX02 U3022 ( .S(n86), .A0(n2530), .A1(gcm_dak_cmd_in[29]), .Z(n1117));
Q_AN02 U3023 ( .A0(n35), .A1(n1118), .Z(gcm_dak_cmd_in_nxt[28]));
Q_MX02 U3024 ( .S(n86), .A0(n2531), .A1(gcm_dak_cmd_in[28]), .Z(n1118));
Q_AN02 U3025 ( .A0(n35), .A1(n1119), .Z(gcm_dak_cmd_in_nxt[27]));
Q_MX02 U3026 ( .S(n86), .A0(n2532), .A1(gcm_dak_cmd_in[27]), .Z(n1119));
Q_AN02 U3027 ( .A0(n35), .A1(n1120), .Z(gcm_dak_cmd_in_nxt[26]));
Q_MX02 U3028 ( .S(n86), .A0(n2533), .A1(gcm_dak_cmd_in[26]), .Z(n1120));
Q_AN02 U3029 ( .A0(n35), .A1(n1121), .Z(gcm_dak_cmd_in_nxt[25]));
Q_MX02 U3030 ( .S(n86), .A0(n2534), .A1(gcm_dak_cmd_in[25]), .Z(n1121));
Q_AN02 U3031 ( .A0(n35), .A1(n1122), .Z(gcm_dak_cmd_in_nxt[24]));
Q_MX02 U3032 ( .S(n86), .A0(n2535), .A1(gcm_dak_cmd_in[24]), .Z(n1122));
Q_AN02 U3033 ( .A0(n35), .A1(n1123), .Z(gcm_dak_cmd_in_nxt[23]));
Q_MX02 U3034 ( .S(n86), .A0(n2536), .A1(gcm_dak_cmd_in[23]), .Z(n1123));
Q_AN02 U3035 ( .A0(n35), .A1(n1124), .Z(gcm_dak_cmd_in_nxt[22]));
Q_MX02 U3036 ( .S(n86), .A0(n2537), .A1(gcm_dak_cmd_in[22]), .Z(n1124));
Q_AN02 U3037 ( .A0(n35), .A1(n1125), .Z(gcm_dak_cmd_in_nxt[21]));
Q_MX02 U3038 ( .S(n86), .A0(n2538), .A1(gcm_dak_cmd_in[21]), .Z(n1125));
Q_AN02 U3039 ( .A0(n35), .A1(n1126), .Z(gcm_dak_cmd_in_nxt[20]));
Q_MX02 U3040 ( .S(n86), .A0(n2539), .A1(gcm_dak_cmd_in[20]), .Z(n1126));
Q_AN02 U3041 ( .A0(n35), .A1(n1127), .Z(gcm_dak_cmd_in_nxt[19]));
Q_MX02 U3042 ( .S(n86), .A0(n2540), .A1(gcm_dak_cmd_in[19]), .Z(n1127));
Q_AN02 U3043 ( .A0(n35), .A1(n1128), .Z(gcm_dak_cmd_in_nxt[18]));
Q_MX02 U3044 ( .S(n86), .A0(n2541), .A1(gcm_dak_cmd_in[18]), .Z(n1128));
Q_AN02 U3045 ( .A0(n35), .A1(n1129), .Z(gcm_dak_cmd_in_nxt[17]));
Q_MX02 U3046 ( .S(n86), .A0(n2542), .A1(gcm_dak_cmd_in[17]), .Z(n1129));
Q_AN02 U3047 ( .A0(n35), .A1(n1130), .Z(gcm_dak_cmd_in_nxt[16]));
Q_MX02 U3048 ( .S(n86), .A0(n2543), .A1(gcm_dak_cmd_in[16]), .Z(n1130));
Q_AN02 U3049 ( .A0(n35), .A1(n1131), .Z(gcm_dak_cmd_in_nxt[15]));
Q_MX02 U3050 ( .S(n86), .A0(n2544), .A1(gcm_dak_cmd_in[15]), .Z(n1131));
Q_AN02 U3051 ( .A0(n35), .A1(n1132), .Z(gcm_dak_cmd_in_nxt[14]));
Q_MX02 U3052 ( .S(n86), .A0(n2545), .A1(gcm_dak_cmd_in[14]), .Z(n1132));
Q_AN02 U3053 ( .A0(n35), .A1(n1133), .Z(gcm_dak_cmd_in_nxt[13]));
Q_MX02 U3054 ( .S(n86), .A0(n2546), .A1(gcm_dak_cmd_in[13]), .Z(n1133));
Q_AN02 U3055 ( .A0(n35), .A1(n1134), .Z(gcm_dak_cmd_in_nxt[12]));
Q_MX02 U3056 ( .S(n86), .A0(n2547), .A1(gcm_dak_cmd_in[12]), .Z(n1134));
Q_AN02 U3057 ( .A0(n35), .A1(n1135), .Z(gcm_dak_cmd_in_nxt[11]));
Q_MX02 U3058 ( .S(n86), .A0(n2548), .A1(gcm_dak_cmd_in[11]), .Z(n1135));
Q_AN02 U3059 ( .A0(n35), .A1(n1136), .Z(gcm_dak_cmd_in_nxt[10]));
Q_MX02 U3060 ( .S(n86), .A0(n2549), .A1(gcm_dak_cmd_in[10]), .Z(n1136));
Q_AN02 U3061 ( .A0(n35), .A1(n1137), .Z(gcm_dak_cmd_in_nxt[9]));
Q_MX02 U3062 ( .S(n86), .A0(n2550), .A1(gcm_dak_cmd_in[9]), .Z(n1137));
Q_AN02 U3063 ( .A0(n35), .A1(n1138), .Z(gcm_dak_cmd_in_nxt[8]));
Q_MX02 U3064 ( .S(n86), .A0(n2551), .A1(gcm_dak_cmd_in[8]), .Z(n1138));
Q_AN02 U3065 ( .A0(n35), .A1(n1139), .Z(gcm_dak_cmd_in_nxt[7]));
Q_MX02 U3066 ( .S(n86), .A0(n2552), .A1(gcm_dak_cmd_in[7]), .Z(n1139));
Q_AN02 U3067 ( .A0(n35), .A1(n1140), .Z(gcm_dak_cmd_in_nxt[6]));
Q_MX02 U3068 ( .S(n86), .A0(n2553), .A1(gcm_dak_cmd_in[6]), .Z(n1140));
Q_AN02 U3069 ( .A0(n35), .A1(n1141), .Z(gcm_dak_cmd_in_nxt[5]));
Q_MX02 U3070 ( .S(n86), .A0(n2554), .A1(gcm_dak_cmd_in[5]), .Z(n1141));
Q_AN02 U3071 ( .A0(n35), .A1(n1142), .Z(gcm_dak_cmd_in_nxt[4]));
Q_MX02 U3072 ( .S(n86), .A0(n2555), .A1(gcm_dak_cmd_in[4]), .Z(n1142));
Q_AN02 U3073 ( .A0(n35), .A1(n1143), .Z(gcm_dak_cmd_in_nxt[3]));
Q_MX02 U3074 ( .S(n86), .A0(n2556), .A1(gcm_dak_cmd_in[3]), .Z(n1143));
Q_AN02 U3075 ( .A0(n35), .A1(n1144), .Z(gcm_dak_cmd_in_nxt[98]));
Q_MX02 U3076 ( .S(n86), .A0(n2557), .A1(gcm_dak_cmd_in[98]), .Z(n1144));
Q_AN02 U3077 ( .A0(n35), .A1(n1145), .Z(gcm_dak_cmd_in_nxt[97]));
Q_MX02 U3078 ( .S(n86), .A0(n2558), .A1(gcm_dak_cmd_in[97]), .Z(n1145));
Q_AN02 U3079 ( .A0(n35), .A1(n1146), .Z(gcm_dak_cmd_in_nxt[96]));
Q_MX02 U3080 ( .S(n86), .A0(n2559), .A1(gcm_dak_cmd_in[96]), .Z(n1146));
Q_AN02 U3081 ( .A0(n35), .A1(n1147), .Z(gcm_dak_cmd_in_nxt[95]));
Q_MX02 U3082 ( .S(n86), .A0(n2560), .A1(gcm_dak_cmd_in[95]), .Z(n1147));
Q_AN02 U3083 ( .A0(n35), .A1(n1148), .Z(gcm_dak_cmd_in_nxt[94]));
Q_MX02 U3084 ( .S(n86), .A0(n2561), .A1(gcm_dak_cmd_in[94]), .Z(n1148));
Q_AN02 U3085 ( .A0(n35), .A1(n1149), .Z(gcm_dak_cmd_in_nxt[93]));
Q_MX02 U3086 ( .S(n86), .A0(n2562), .A1(gcm_dak_cmd_in[93]), .Z(n1149));
Q_AN02 U3087 ( .A0(n35), .A1(n1150), .Z(gcm_dak_cmd_in_nxt[92]));
Q_MX02 U3088 ( .S(n86), .A0(n2563), .A1(gcm_dak_cmd_in[92]), .Z(n1150));
Q_AN02 U3089 ( .A0(n35), .A1(n1151), .Z(gcm_dak_cmd_in_nxt[91]));
Q_MX02 U3090 ( .S(n86), .A0(n2564), .A1(gcm_dak_cmd_in[91]), .Z(n1151));
Q_AN02 U3091 ( .A0(n35), .A1(n1152), .Z(gcm_dak_cmd_in_nxt[90]));
Q_MX02 U3092 ( .S(n86), .A0(n2565), .A1(gcm_dak_cmd_in[90]), .Z(n1152));
Q_AN02 U3093 ( .A0(n35), .A1(n1153), .Z(gcm_dak_cmd_in_nxt[89]));
Q_MX02 U3094 ( .S(n86), .A0(n2566), .A1(gcm_dak_cmd_in[89]), .Z(n1153));
Q_AN02 U3095 ( .A0(n35), .A1(n1154), .Z(gcm_dak_cmd_in_nxt[88]));
Q_MX02 U3096 ( .S(n86), .A0(n2567), .A1(gcm_dak_cmd_in[88]), .Z(n1154));
Q_AN02 U3097 ( .A0(n35), .A1(n1155), .Z(gcm_dak_cmd_in_nxt[87]));
Q_MX02 U3098 ( .S(n86), .A0(n2568), .A1(gcm_dak_cmd_in[87]), .Z(n1155));
Q_AN02 U3099 ( .A0(n35), .A1(n1156), .Z(gcm_dak_cmd_in_nxt[86]));
Q_MX02 U3100 ( .S(n86), .A0(n2569), .A1(gcm_dak_cmd_in[86]), .Z(n1156));
Q_AN02 U3101 ( .A0(n35), .A1(n1157), .Z(gcm_dak_cmd_in_nxt[85]));
Q_MX02 U3102 ( .S(n86), .A0(n2570), .A1(gcm_dak_cmd_in[85]), .Z(n1157));
Q_AN02 U3103 ( .A0(n35), .A1(n1158), .Z(gcm_dak_cmd_in_nxt[84]));
Q_MX02 U3104 ( .S(n86), .A0(n2571), .A1(gcm_dak_cmd_in[84]), .Z(n1158));
Q_AN02 U3105 ( .A0(n35), .A1(n1159), .Z(gcm_dak_cmd_in_nxt[83]));
Q_MX02 U3106 ( .S(n86), .A0(n2572), .A1(gcm_dak_cmd_in[83]), .Z(n1159));
Q_AN02 U3107 ( .A0(n35), .A1(n1160), .Z(gcm_dak_cmd_in_nxt[82]));
Q_MX02 U3108 ( .S(n86), .A0(n2573), .A1(gcm_dak_cmd_in[82]), .Z(n1160));
Q_AN02 U3109 ( .A0(n35), .A1(n1161), .Z(gcm_dak_cmd_in_nxt[81]));
Q_MX02 U3110 ( .S(n86), .A0(n2574), .A1(gcm_dak_cmd_in[81]), .Z(n1161));
Q_AN02 U3111 ( .A0(n35), .A1(n1162), .Z(gcm_dak_cmd_in_nxt[80]));
Q_MX02 U3112 ( .S(n86), .A0(n2575), .A1(gcm_dak_cmd_in[80]), .Z(n1162));
Q_AN02 U3113 ( .A0(n35), .A1(n1163), .Z(gcm_dak_cmd_in_nxt[79]));
Q_MX02 U3114 ( .S(n86), .A0(n2576), .A1(gcm_dak_cmd_in[79]), .Z(n1163));
Q_AN02 U3115 ( .A0(n35), .A1(n1164), .Z(gcm_dak_cmd_in_nxt[78]));
Q_MX02 U3116 ( .S(n86), .A0(n2577), .A1(gcm_dak_cmd_in[78]), .Z(n1164));
Q_AN02 U3117 ( .A0(n35), .A1(n1165), .Z(gcm_dak_cmd_in_nxt[77]));
Q_MX02 U3118 ( .S(n86), .A0(n2578), .A1(gcm_dak_cmd_in[77]), .Z(n1165));
Q_AN02 U3119 ( .A0(n35), .A1(n1166), .Z(gcm_dak_cmd_in_nxt[76]));
Q_MX02 U3120 ( .S(n86), .A0(n2579), .A1(gcm_dak_cmd_in[76]), .Z(n1166));
Q_AN02 U3121 ( .A0(n35), .A1(n1167), .Z(gcm_dak_cmd_in_nxt[75]));
Q_MX02 U3122 ( .S(n86), .A0(n2580), .A1(gcm_dak_cmd_in[75]), .Z(n1167));
Q_AN02 U3123 ( .A0(n35), .A1(n1168), .Z(gcm_dak_cmd_in_nxt[74]));
Q_MX02 U3124 ( .S(n86), .A0(n2581), .A1(gcm_dak_cmd_in[74]), .Z(n1168));
Q_AN02 U3125 ( .A0(n35), .A1(n1169), .Z(gcm_dak_cmd_in_nxt[73]));
Q_MX02 U3126 ( .S(n86), .A0(n2582), .A1(gcm_dak_cmd_in[73]), .Z(n1169));
Q_AN02 U3127 ( .A0(n35), .A1(n1170), .Z(gcm_dak_cmd_in_nxt[72]));
Q_MX02 U3128 ( .S(n86), .A0(n2583), .A1(gcm_dak_cmd_in[72]), .Z(n1170));
Q_AN02 U3129 ( .A0(n35), .A1(n1171), .Z(gcm_dak_cmd_in_nxt[71]));
Q_MX02 U3130 ( .S(n86), .A0(n2584), .A1(gcm_dak_cmd_in[71]), .Z(n1171));
Q_AN02 U3131 ( .A0(n35), .A1(n1172), .Z(gcm_dak_cmd_in_nxt[70]));
Q_MX02 U3132 ( .S(n86), .A0(n2585), .A1(gcm_dak_cmd_in[70]), .Z(n1172));
Q_AN02 U3133 ( .A0(n35), .A1(n1173), .Z(gcm_dak_cmd_in_nxt[69]));
Q_MX02 U3134 ( .S(n86), .A0(n2586), .A1(gcm_dak_cmd_in[69]), .Z(n1173));
Q_AN02 U3135 ( .A0(n35), .A1(n1174), .Z(gcm_dak_cmd_in_nxt[68]));
Q_MX02 U3136 ( .S(n86), .A0(n2587), .A1(gcm_dak_cmd_in[68]), .Z(n1174));
Q_AN02 U3137 ( .A0(n35), .A1(n1175), .Z(gcm_dak_cmd_in_nxt[67]));
Q_MX02 U3138 ( .S(n86), .A0(n2588), .A1(gcm_dak_cmd_in[67]), .Z(n1175));
Q_AN02 U3139 ( .A0(n35), .A1(n1176), .Z(gcm_dak_cmd_in_nxt[66]));
Q_MX02 U3140 ( .S(n86), .A0(n2589), .A1(gcm_dak_cmd_in[66]), .Z(n1176));
Q_AN02 U3141 ( .A0(n35), .A1(n1177), .Z(gcm_dak_cmd_in_nxt[65]));
Q_MX02 U3142 ( .S(n86), .A0(n2590), .A1(gcm_dak_cmd_in[65]), .Z(n1177));
Q_AN02 U3143 ( .A0(n35), .A1(n1178), .Z(gcm_dak_cmd_in_nxt[64]));
Q_MX02 U3144 ( .S(n86), .A0(n2591), .A1(gcm_dak_cmd_in[64]), .Z(n1178));
Q_AN02 U3145 ( .A0(n35), .A1(n1179), .Z(gcm_dak_cmd_in_nxt[63]));
Q_MX02 U3146 ( .S(n86), .A0(n2592), .A1(gcm_dak_cmd_in[63]), .Z(n1179));
Q_AN02 U3147 ( .A0(n35), .A1(n1180), .Z(gcm_dak_cmd_in_nxt[62]));
Q_MX02 U3148 ( .S(n86), .A0(n2593), .A1(gcm_dak_cmd_in[62]), .Z(n1180));
Q_AN02 U3149 ( .A0(n35), .A1(n1181), .Z(gcm_dak_cmd_in_nxt[61]));
Q_MX02 U3150 ( .S(n86), .A0(n2594), .A1(gcm_dak_cmd_in[61]), .Z(n1181));
Q_AN02 U3151 ( .A0(n35), .A1(n1182), .Z(gcm_dak_cmd_in_nxt[60]));
Q_MX02 U3152 ( .S(n86), .A0(n2595), .A1(gcm_dak_cmd_in[60]), .Z(n1182));
Q_AN02 U3153 ( .A0(n35), .A1(n1183), .Z(gcm_dak_cmd_in_nxt[59]));
Q_MX02 U3154 ( .S(n86), .A0(n2596), .A1(gcm_dak_cmd_in[59]), .Z(n1183));
Q_AN02 U3155 ( .A0(n35), .A1(n1184), .Z(gcm_dak_cmd_in_nxt[58]));
Q_MX02 U3156 ( .S(n86), .A0(n2597), .A1(gcm_dak_cmd_in[58]), .Z(n1184));
Q_AN02 U3157 ( .A0(n35), .A1(n1185), .Z(gcm_dak_cmd_in_nxt[57]));
Q_MX02 U3158 ( .S(n86), .A0(n2598), .A1(gcm_dak_cmd_in[57]), .Z(n1185));
Q_AN02 U3159 ( .A0(n35), .A1(n1186), .Z(gcm_dak_cmd_in_nxt[56]));
Q_MX02 U3160 ( .S(n86), .A0(n2599), .A1(gcm_dak_cmd_in[56]), .Z(n1186));
Q_AN02 U3161 ( .A0(n35), .A1(n1187), .Z(gcm_dak_cmd_in_nxt[55]));
Q_MX02 U3162 ( .S(n86), .A0(n2600), .A1(gcm_dak_cmd_in[55]), .Z(n1187));
Q_AN02 U3163 ( .A0(n35), .A1(n1188), .Z(gcm_dak_cmd_in_nxt[54]));
Q_MX02 U3164 ( .S(n86), .A0(n2601), .A1(gcm_dak_cmd_in[54]), .Z(n1188));
Q_AN02 U3165 ( .A0(n35), .A1(n1189), .Z(gcm_dak_cmd_in_nxt[53]));
Q_MX02 U3166 ( .S(n86), .A0(n2602), .A1(gcm_dak_cmd_in[53]), .Z(n1189));
Q_AN02 U3167 ( .A0(n35), .A1(n1190), .Z(gcm_dak_cmd_in_nxt[52]));
Q_MX02 U3168 ( .S(n86), .A0(n2603), .A1(gcm_dak_cmd_in[52]), .Z(n1190));
Q_AN02 U3169 ( .A0(n35), .A1(n1191), .Z(gcm_dak_cmd_in_nxt[51]));
Q_MX02 U3170 ( .S(n86), .A0(n2604), .A1(gcm_dak_cmd_in[51]), .Z(n1191));
Q_AN02 U3171 ( .A0(n35), .A1(n1192), .Z(gcm_dak_cmd_in_nxt[50]));
Q_MX02 U3172 ( .S(n86), .A0(n2605), .A1(gcm_dak_cmd_in[50]), .Z(n1192));
Q_AN02 U3173 ( .A0(n35), .A1(n1193), .Z(gcm_dak_cmd_in_nxt[49]));
Q_MX02 U3174 ( .S(n86), .A0(n2606), .A1(gcm_dak_cmd_in[49]), .Z(n1193));
Q_AN02 U3175 ( .A0(n35), .A1(n1194), .Z(gcm_dak_cmd_in_nxt[48]));
Q_MX02 U3176 ( .S(n86), .A0(n2607), .A1(gcm_dak_cmd_in[48]), .Z(n1194));
Q_AN02 U3177 ( .A0(n35), .A1(n1195), .Z(gcm_dak_cmd_in_nxt[47]));
Q_MX02 U3178 ( .S(n86), .A0(n2608), .A1(gcm_dak_cmd_in[47]), .Z(n1195));
Q_AN02 U3179 ( .A0(n35), .A1(n1196), .Z(gcm_dak_cmd_in_nxt[46]));
Q_MX02 U3180 ( .S(n86), .A0(n2609), .A1(gcm_dak_cmd_in[46]), .Z(n1196));
Q_AN02 U3181 ( .A0(n35), .A1(n1197), .Z(gcm_dak_cmd_in_nxt[45]));
Q_MX02 U3182 ( .S(n86), .A0(n2610), .A1(gcm_dak_cmd_in[45]), .Z(n1197));
Q_AN02 U3183 ( .A0(n35), .A1(n1198), .Z(gcm_dak_cmd_in_nxt[44]));
Q_MX02 U3184 ( .S(n86), .A0(n2611), .A1(gcm_dak_cmd_in[44]), .Z(n1198));
Q_AN02 U3185 ( .A0(n35), .A1(n1199), .Z(gcm_dak_cmd_in_nxt[43]));
Q_MX02 U3186 ( .S(n86), .A0(n2612), .A1(gcm_dak_cmd_in[43]), .Z(n1199));
Q_AN02 U3187 ( .A0(n35), .A1(n1200), .Z(gcm_dak_cmd_in_nxt[42]));
Q_MX02 U3188 ( .S(n86), .A0(n2613), .A1(gcm_dak_cmd_in[42]), .Z(n1200));
Q_AN02 U3189 ( .A0(n35), .A1(n1201), .Z(gcm_dak_cmd_in_nxt[41]));
Q_MX02 U3190 ( .S(n86), .A0(n2614), .A1(gcm_dak_cmd_in[41]), .Z(n1201));
Q_AN02 U3191 ( .A0(n35), .A1(n1202), .Z(gcm_dak_cmd_in_nxt[40]));
Q_MX02 U3192 ( .S(n86), .A0(n2615), .A1(gcm_dak_cmd_in[40]), .Z(n1202));
Q_AN02 U3193 ( .A0(n35), .A1(n1203), .Z(gcm_dak_cmd_in_nxt[39]));
Q_MX02 U3194 ( .S(n86), .A0(n2616), .A1(gcm_dak_cmd_in[39]), .Z(n1203));
Q_AN02 U3195 ( .A0(n35), .A1(n1204), .Z(gcm_dak_cmd_in_nxt[38]));
Q_MX02 U3196 ( .S(n86), .A0(n2617), .A1(gcm_dak_cmd_in[38]), .Z(n1204));
Q_AN02 U3197 ( .A0(n35), .A1(n1205), .Z(gcm_dak_cmd_in_nxt[37]));
Q_MX02 U3198 ( .S(n86), .A0(n2618), .A1(gcm_dak_cmd_in[37]), .Z(n1205));
Q_AN02 U3199 ( .A0(n35), .A1(n1206), .Z(gcm_dak_cmd_in_nxt[36]));
Q_MX02 U3200 ( .S(n86), .A0(n2619), .A1(gcm_dak_cmd_in[36]), .Z(n1206));
Q_AN02 U3201 ( .A0(n35), .A1(n1207), .Z(gcm_dak_cmd_in_nxt[35]));
Q_MX02 U3202 ( .S(n86), .A0(n2620), .A1(gcm_dak_cmd_in[35]), .Z(n1207));
Q_AN02 U3203 ( .A0(n35), .A1(n1208), .Z(gcm_dak_cmd_in_nxt[354]));
Q_MX02 U3204 ( .S(n90), .A0(gcm_dak_cmd_in[290]), .A1(gcm_dak_cmd_in[354]), .Z(n1208));
Q_AN02 U3205 ( .A0(n35), .A1(n1209), .Z(gcm_dak_cmd_in_nxt[353]));
Q_MX02 U3206 ( .S(n90), .A0(gcm_dak_cmd_in[289]), .A1(gcm_dak_cmd_in[353]), .Z(n1209));
Q_AN02 U3207 ( .A0(n35), .A1(n1210), .Z(gcm_dak_cmd_in_nxt[352]));
Q_MX02 U3208 ( .S(n90), .A0(gcm_dak_cmd_in[288]), .A1(gcm_dak_cmd_in[352]), .Z(n1210));
Q_AN02 U3209 ( .A0(n35), .A1(n1211), .Z(gcm_dak_cmd_in_nxt[351]));
Q_MX02 U3210 ( .S(n90), .A0(gcm_dak_cmd_in[287]), .A1(gcm_dak_cmd_in[351]), .Z(n1211));
Q_AN02 U3211 ( .A0(n35), .A1(n1212), .Z(gcm_dak_cmd_in_nxt[350]));
Q_MX02 U3212 ( .S(n90), .A0(gcm_dak_cmd_in[286]), .A1(gcm_dak_cmd_in[350]), .Z(n1212));
Q_AN02 U3213 ( .A0(n35), .A1(n1213), .Z(gcm_dak_cmd_in_nxt[349]));
Q_MX02 U3214 ( .S(n90), .A0(gcm_dak_cmd_in[285]), .A1(gcm_dak_cmd_in[349]), .Z(n1213));
Q_AN02 U3215 ( .A0(n35), .A1(n1214), .Z(gcm_dak_cmd_in_nxt[348]));
Q_MX02 U3216 ( .S(n90), .A0(gcm_dak_cmd_in[284]), .A1(gcm_dak_cmd_in[348]), .Z(n1214));
Q_AN02 U3217 ( .A0(n35), .A1(n1215), .Z(gcm_dak_cmd_in_nxt[347]));
Q_MX02 U3218 ( .S(n90), .A0(gcm_dak_cmd_in[283]), .A1(gcm_dak_cmd_in[347]), .Z(n1215));
Q_AN02 U3219 ( .A0(n35), .A1(n1216), .Z(gcm_dak_cmd_in_nxt[346]));
Q_MX02 U3220 ( .S(n90), .A0(gcm_dak_cmd_in[282]), .A1(gcm_dak_cmd_in[346]), .Z(n1216));
Q_AN02 U3221 ( .A0(n35), .A1(n1217), .Z(gcm_dak_cmd_in_nxt[345]));
Q_MX02 U3222 ( .S(n90), .A0(gcm_dak_cmd_in[281]), .A1(gcm_dak_cmd_in[345]), .Z(n1217));
Q_AN02 U3223 ( .A0(n35), .A1(n1218), .Z(gcm_dak_cmd_in_nxt[344]));
Q_MX02 U3224 ( .S(n90), .A0(gcm_dak_cmd_in[280]), .A1(gcm_dak_cmd_in[344]), .Z(n1218));
Q_AN02 U3225 ( .A0(n35), .A1(n1219), .Z(gcm_dak_cmd_in_nxt[343]));
Q_MX02 U3226 ( .S(n90), .A0(gcm_dak_cmd_in[279]), .A1(gcm_dak_cmd_in[343]), .Z(n1219));
Q_AN02 U3227 ( .A0(n35), .A1(n1220), .Z(gcm_dak_cmd_in_nxt[342]));
Q_MX02 U3228 ( .S(n90), .A0(gcm_dak_cmd_in[278]), .A1(gcm_dak_cmd_in[342]), .Z(n1220));
Q_AN02 U3229 ( .A0(n35), .A1(n1221), .Z(gcm_dak_cmd_in_nxt[341]));
Q_MX02 U3230 ( .S(n90), .A0(gcm_dak_cmd_in[277]), .A1(gcm_dak_cmd_in[341]), .Z(n1221));
Q_AN02 U3231 ( .A0(n35), .A1(n1222), .Z(gcm_dak_cmd_in_nxt[340]));
Q_MX02 U3232 ( .S(n90), .A0(gcm_dak_cmd_in[276]), .A1(gcm_dak_cmd_in[340]), .Z(n1222));
Q_AN02 U3233 ( .A0(n35), .A1(n1223), .Z(gcm_dak_cmd_in_nxt[339]));
Q_MX02 U3234 ( .S(n90), .A0(gcm_dak_cmd_in[275]), .A1(gcm_dak_cmd_in[339]), .Z(n1223));
Q_AN02 U3235 ( .A0(n35), .A1(n1224), .Z(gcm_dak_cmd_in_nxt[338]));
Q_MX02 U3236 ( .S(n90), .A0(gcm_dak_cmd_in[274]), .A1(gcm_dak_cmd_in[338]), .Z(n1224));
Q_AN02 U3237 ( .A0(n35), .A1(n1225), .Z(gcm_dak_cmd_in_nxt[337]));
Q_MX02 U3238 ( .S(n90), .A0(gcm_dak_cmd_in[273]), .A1(gcm_dak_cmd_in[337]), .Z(n1225));
Q_AN02 U3239 ( .A0(n35), .A1(n1226), .Z(gcm_dak_cmd_in_nxt[336]));
Q_MX02 U3240 ( .S(n90), .A0(gcm_dak_cmd_in[272]), .A1(gcm_dak_cmd_in[336]), .Z(n1226));
Q_AN02 U3241 ( .A0(n35), .A1(n1227), .Z(gcm_dak_cmd_in_nxt[335]));
Q_MX02 U3242 ( .S(n90), .A0(gcm_dak_cmd_in[271]), .A1(gcm_dak_cmd_in[335]), .Z(n1227));
Q_AN02 U3243 ( .A0(n35), .A1(n1228), .Z(gcm_dak_cmd_in_nxt[334]));
Q_MX02 U3244 ( .S(n90), .A0(gcm_dak_cmd_in[270]), .A1(gcm_dak_cmd_in[334]), .Z(n1228));
Q_AN02 U3245 ( .A0(n35), .A1(n1229), .Z(gcm_dak_cmd_in_nxt[333]));
Q_MX02 U3246 ( .S(n90), .A0(gcm_dak_cmd_in[269]), .A1(gcm_dak_cmd_in[333]), .Z(n1229));
Q_AN02 U3247 ( .A0(n35), .A1(n1230), .Z(gcm_dak_cmd_in_nxt[332]));
Q_MX02 U3248 ( .S(n90), .A0(gcm_dak_cmd_in[268]), .A1(gcm_dak_cmd_in[332]), .Z(n1230));
Q_AN02 U3249 ( .A0(n35), .A1(n1231), .Z(gcm_dak_cmd_in_nxt[331]));
Q_MX02 U3250 ( .S(n90), .A0(gcm_dak_cmd_in[267]), .A1(gcm_dak_cmd_in[331]), .Z(n1231));
Q_AN02 U3251 ( .A0(n35), .A1(n1232), .Z(gcm_dak_cmd_in_nxt[330]));
Q_MX02 U3252 ( .S(n90), .A0(gcm_dak_cmd_in[266]), .A1(gcm_dak_cmd_in[330]), .Z(n1232));
Q_AN02 U3253 ( .A0(n35), .A1(n1233), .Z(gcm_dak_cmd_in_nxt[329]));
Q_MX02 U3254 ( .S(n90), .A0(gcm_dak_cmd_in[265]), .A1(gcm_dak_cmd_in[329]), .Z(n1233));
Q_AN02 U3255 ( .A0(n35), .A1(n1234), .Z(gcm_dak_cmd_in_nxt[328]));
Q_MX02 U3256 ( .S(n90), .A0(gcm_dak_cmd_in[264]), .A1(gcm_dak_cmd_in[328]), .Z(n1234));
Q_AN02 U3257 ( .A0(n35), .A1(n1235), .Z(gcm_dak_cmd_in_nxt[327]));
Q_MX02 U3258 ( .S(n90), .A0(gcm_dak_cmd_in[263]), .A1(gcm_dak_cmd_in[327]), .Z(n1235));
Q_AN02 U3259 ( .A0(n35), .A1(n1236), .Z(gcm_dak_cmd_in_nxt[326]));
Q_MX02 U3260 ( .S(n90), .A0(gcm_dak_cmd_in[262]), .A1(gcm_dak_cmd_in[326]), .Z(n1236));
Q_AN02 U3261 ( .A0(n35), .A1(n1237), .Z(gcm_dak_cmd_in_nxt[325]));
Q_MX02 U3262 ( .S(n90), .A0(gcm_dak_cmd_in[261]), .A1(gcm_dak_cmd_in[325]), .Z(n1237));
Q_AN02 U3263 ( .A0(n35), .A1(n1238), .Z(gcm_dak_cmd_in_nxt[324]));
Q_MX02 U3264 ( .S(n90), .A0(gcm_dak_cmd_in[260]), .A1(gcm_dak_cmd_in[324]), .Z(n1238));
Q_AN02 U3265 ( .A0(n35), .A1(n1239), .Z(gcm_dak_cmd_in_nxt[323]));
Q_MX02 U3266 ( .S(n90), .A0(gcm_dak_cmd_in[259]), .A1(gcm_dak_cmd_in[323]), .Z(n1239));
Q_AN02 U3267 ( .A0(n35), .A1(n1240), .Z(gcm_dak_cmd_in_nxt[322]));
Q_MX02 U3268 ( .S(n90), .A0(gcm_dak_cmd_in[258]), .A1(gcm_dak_cmd_in[322]), .Z(n1240));
Q_AN02 U3269 ( .A0(n35), .A1(n1241), .Z(gcm_dak_cmd_in_nxt[321]));
Q_MX02 U3270 ( .S(n90), .A0(gcm_dak_cmd_in[257]), .A1(gcm_dak_cmd_in[321]), .Z(n1241));
Q_AN02 U3271 ( .A0(n35), .A1(n1242), .Z(gcm_dak_cmd_in_nxt[320]));
Q_MX02 U3272 ( .S(n90), .A0(gcm_dak_cmd_in[256]), .A1(gcm_dak_cmd_in[320]), .Z(n1242));
Q_AN02 U3273 ( .A0(n35), .A1(n1243), .Z(gcm_dak_cmd_in_nxt[319]));
Q_MX02 U3274 ( .S(n90), .A0(gcm_dak_cmd_in[255]), .A1(gcm_dak_cmd_in[319]), .Z(n1243));
Q_AN02 U3275 ( .A0(n35), .A1(n1244), .Z(gcm_dak_cmd_in_nxt[318]));
Q_MX02 U3276 ( .S(n90), .A0(gcm_dak_cmd_in[254]), .A1(gcm_dak_cmd_in[318]), .Z(n1244));
Q_AN02 U3277 ( .A0(n35), .A1(n1245), .Z(gcm_dak_cmd_in_nxt[317]));
Q_MX02 U3278 ( .S(n90), .A0(gcm_dak_cmd_in[253]), .A1(gcm_dak_cmd_in[317]), .Z(n1245));
Q_AN02 U3279 ( .A0(n35), .A1(n1246), .Z(gcm_dak_cmd_in_nxt[316]));
Q_MX02 U3280 ( .S(n90), .A0(gcm_dak_cmd_in[252]), .A1(gcm_dak_cmd_in[316]), .Z(n1246));
Q_AN02 U3281 ( .A0(n35), .A1(n1247), .Z(gcm_dak_cmd_in_nxt[315]));
Q_MX02 U3282 ( .S(n90), .A0(gcm_dak_cmd_in[251]), .A1(gcm_dak_cmd_in[315]), .Z(n1247));
Q_AN02 U3283 ( .A0(n35), .A1(n1248), .Z(gcm_dak_cmd_in_nxt[314]));
Q_MX02 U3284 ( .S(n90), .A0(gcm_dak_cmd_in[250]), .A1(gcm_dak_cmd_in[314]), .Z(n1248));
Q_AN02 U3285 ( .A0(n35), .A1(n1249), .Z(gcm_dak_cmd_in_nxt[313]));
Q_MX02 U3286 ( .S(n90), .A0(gcm_dak_cmd_in[249]), .A1(gcm_dak_cmd_in[313]), .Z(n1249));
Q_AN02 U3287 ( .A0(n35), .A1(n1250), .Z(gcm_dak_cmd_in_nxt[312]));
Q_MX02 U3288 ( .S(n90), .A0(gcm_dak_cmd_in[248]), .A1(gcm_dak_cmd_in[312]), .Z(n1250));
Q_AN02 U3289 ( .A0(n35), .A1(n1251), .Z(gcm_dak_cmd_in_nxt[311]));
Q_MX02 U3290 ( .S(n90), .A0(gcm_dak_cmd_in[247]), .A1(gcm_dak_cmd_in[311]), .Z(n1251));
Q_AN02 U3291 ( .A0(n35), .A1(n1252), .Z(gcm_dak_cmd_in_nxt[310]));
Q_MX02 U3292 ( .S(n90), .A0(gcm_dak_cmd_in[246]), .A1(gcm_dak_cmd_in[310]), .Z(n1252));
Q_AN02 U3293 ( .A0(n35), .A1(n1253), .Z(gcm_dak_cmd_in_nxt[309]));
Q_MX02 U3294 ( .S(n90), .A0(gcm_dak_cmd_in[245]), .A1(gcm_dak_cmd_in[309]), .Z(n1253));
Q_AN02 U3295 ( .A0(n35), .A1(n1254), .Z(gcm_dak_cmd_in_nxt[308]));
Q_MX02 U3296 ( .S(n90), .A0(gcm_dak_cmd_in[244]), .A1(gcm_dak_cmd_in[308]), .Z(n1254));
Q_AN02 U3297 ( .A0(n35), .A1(n1255), .Z(gcm_dak_cmd_in_nxt[307]));
Q_MX02 U3298 ( .S(n90), .A0(gcm_dak_cmd_in[243]), .A1(gcm_dak_cmd_in[307]), .Z(n1255));
Q_AN02 U3299 ( .A0(n35), .A1(n1256), .Z(gcm_dak_cmd_in_nxt[306]));
Q_MX02 U3300 ( .S(n90), .A0(gcm_dak_cmd_in[242]), .A1(gcm_dak_cmd_in[306]), .Z(n1256));
Q_AN02 U3301 ( .A0(n35), .A1(n1257), .Z(gcm_dak_cmd_in_nxt[305]));
Q_MX02 U3302 ( .S(n90), .A0(gcm_dak_cmd_in[241]), .A1(gcm_dak_cmd_in[305]), .Z(n1257));
Q_AN02 U3303 ( .A0(n35), .A1(n1258), .Z(gcm_dak_cmd_in_nxt[304]));
Q_MX02 U3304 ( .S(n90), .A0(gcm_dak_cmd_in[240]), .A1(gcm_dak_cmd_in[304]), .Z(n1258));
Q_AN02 U3305 ( .A0(n35), .A1(n1259), .Z(gcm_dak_cmd_in_nxt[303]));
Q_MX02 U3306 ( .S(n90), .A0(gcm_dak_cmd_in[239]), .A1(gcm_dak_cmd_in[303]), .Z(n1259));
Q_AN02 U3307 ( .A0(n35), .A1(n1260), .Z(gcm_dak_cmd_in_nxt[302]));
Q_MX02 U3308 ( .S(n90), .A0(gcm_dak_cmd_in[238]), .A1(gcm_dak_cmd_in[302]), .Z(n1260));
Q_AN02 U3309 ( .A0(n35), .A1(n1261), .Z(gcm_dak_cmd_in_nxt[301]));
Q_MX02 U3310 ( .S(n90), .A0(gcm_dak_cmd_in[237]), .A1(gcm_dak_cmd_in[301]), .Z(n1261));
Q_AN02 U3311 ( .A0(n35), .A1(n1262), .Z(gcm_dak_cmd_in_nxt[300]));
Q_MX02 U3312 ( .S(n90), .A0(gcm_dak_cmd_in[236]), .A1(gcm_dak_cmd_in[300]), .Z(n1262));
Q_AN02 U3313 ( .A0(n35), .A1(n1263), .Z(gcm_dak_cmd_in_nxt[299]));
Q_MX02 U3314 ( .S(n90), .A0(gcm_dak_cmd_in[235]), .A1(gcm_dak_cmd_in[299]), .Z(n1263));
Q_AN02 U3315 ( .A0(n35), .A1(n1264), .Z(gcm_dak_cmd_in_nxt[298]));
Q_MX02 U3316 ( .S(n90), .A0(gcm_dak_cmd_in[234]), .A1(gcm_dak_cmd_in[298]), .Z(n1264));
Q_AN02 U3317 ( .A0(n35), .A1(n1265), .Z(gcm_dak_cmd_in_nxt[297]));
Q_MX02 U3318 ( .S(n90), .A0(gcm_dak_cmd_in[233]), .A1(gcm_dak_cmd_in[297]), .Z(n1265));
Q_AN02 U3319 ( .A0(n35), .A1(n1266), .Z(gcm_dak_cmd_in_nxt[296]));
Q_MX02 U3320 ( .S(n90), .A0(gcm_dak_cmd_in[232]), .A1(gcm_dak_cmd_in[296]), .Z(n1266));
Q_AN02 U3321 ( .A0(n35), .A1(n1267), .Z(gcm_dak_cmd_in_nxt[295]));
Q_MX02 U3322 ( .S(n90), .A0(gcm_dak_cmd_in[231]), .A1(gcm_dak_cmd_in[295]), .Z(n1267));
Q_AN02 U3323 ( .A0(n35), .A1(n1268), .Z(gcm_dak_cmd_in_nxt[294]));
Q_MX02 U3324 ( .S(n90), .A0(gcm_dak_cmd_in[230]), .A1(gcm_dak_cmd_in[294]), .Z(n1268));
Q_AN02 U3325 ( .A0(n35), .A1(n1269), .Z(gcm_dak_cmd_in_nxt[293]));
Q_MX02 U3326 ( .S(n90), .A0(gcm_dak_cmd_in[229]), .A1(gcm_dak_cmd_in[293]), .Z(n1269));
Q_AN02 U3327 ( .A0(n35), .A1(n1270), .Z(gcm_dak_cmd_in_nxt[292]));
Q_MX02 U3328 ( .S(n90), .A0(gcm_dak_cmd_in[228]), .A1(gcm_dak_cmd_in[292]), .Z(n1270));
Q_AN02 U3329 ( .A0(n35), .A1(n1271), .Z(gcm_dak_cmd_in_nxt[291]));
Q_MX02 U3330 ( .S(n90), .A0(gcm_dak_cmd_in[227]), .A1(gcm_dak_cmd_in[291]), .Z(n1271));
Q_AN02 U3331 ( .A0(n35), .A1(n1272), .Z(gcm_dak_cmd_in_nxt[290]));
Q_MX02 U3332 ( .S(n90), .A0(gcm_dak_cmd_in[226]), .A1(gcm_dak_cmd_in[290]), .Z(n1272));
Q_AN02 U3333 ( .A0(n35), .A1(n1273), .Z(gcm_dak_cmd_in_nxt[289]));
Q_MX02 U3334 ( .S(n90), .A0(gcm_dak_cmd_in[225]), .A1(gcm_dak_cmd_in[289]), .Z(n1273));
Q_AN02 U3335 ( .A0(n35), .A1(n1274), .Z(gcm_dak_cmd_in_nxt[288]));
Q_MX02 U3336 ( .S(n90), .A0(gcm_dak_cmd_in[224]), .A1(gcm_dak_cmd_in[288]), .Z(n1274));
Q_AN02 U3337 ( .A0(n35), .A1(n1275), .Z(gcm_dak_cmd_in_nxt[287]));
Q_MX02 U3338 ( .S(n90), .A0(gcm_dak_cmd_in[223]), .A1(gcm_dak_cmd_in[287]), .Z(n1275));
Q_AN02 U3339 ( .A0(n35), .A1(n1276), .Z(gcm_dak_cmd_in_nxt[286]));
Q_MX02 U3340 ( .S(n90), .A0(gcm_dak_cmd_in[222]), .A1(gcm_dak_cmd_in[286]), .Z(n1276));
Q_AN02 U3341 ( .A0(n35), .A1(n1277), .Z(gcm_dak_cmd_in_nxt[285]));
Q_MX02 U3342 ( .S(n90), .A0(gcm_dak_cmd_in[221]), .A1(gcm_dak_cmd_in[285]), .Z(n1277));
Q_AN02 U3343 ( .A0(n35), .A1(n1278), .Z(gcm_dak_cmd_in_nxt[284]));
Q_MX02 U3344 ( .S(n90), .A0(gcm_dak_cmd_in[220]), .A1(gcm_dak_cmd_in[284]), .Z(n1278));
Q_AN02 U3345 ( .A0(n35), .A1(n1279), .Z(gcm_dak_cmd_in_nxt[283]));
Q_MX02 U3346 ( .S(n90), .A0(gcm_dak_cmd_in[219]), .A1(gcm_dak_cmd_in[283]), .Z(n1279));
Q_AN02 U3347 ( .A0(n35), .A1(n1280), .Z(gcm_dak_cmd_in_nxt[282]));
Q_MX02 U3348 ( .S(n90), .A0(gcm_dak_cmd_in[218]), .A1(gcm_dak_cmd_in[282]), .Z(n1280));
Q_AN02 U3349 ( .A0(n35), .A1(n1281), .Z(gcm_dak_cmd_in_nxt[281]));
Q_MX02 U3350 ( .S(n90), .A0(gcm_dak_cmd_in[217]), .A1(gcm_dak_cmd_in[281]), .Z(n1281));
Q_AN02 U3351 ( .A0(n35), .A1(n1282), .Z(gcm_dak_cmd_in_nxt[280]));
Q_MX02 U3352 ( .S(n90), .A0(gcm_dak_cmd_in[216]), .A1(gcm_dak_cmd_in[280]), .Z(n1282));
Q_AN02 U3353 ( .A0(n35), .A1(n1283), .Z(gcm_dak_cmd_in_nxt[279]));
Q_MX02 U3354 ( .S(n90), .A0(gcm_dak_cmd_in[215]), .A1(gcm_dak_cmd_in[279]), .Z(n1283));
Q_AN02 U3355 ( .A0(n35), .A1(n1284), .Z(gcm_dak_cmd_in_nxt[278]));
Q_MX02 U3356 ( .S(n90), .A0(gcm_dak_cmd_in[214]), .A1(gcm_dak_cmd_in[278]), .Z(n1284));
Q_AN02 U3357 ( .A0(n35), .A1(n1285), .Z(gcm_dak_cmd_in_nxt[277]));
Q_MX02 U3358 ( .S(n90), .A0(gcm_dak_cmd_in[213]), .A1(gcm_dak_cmd_in[277]), .Z(n1285));
Q_AN02 U3359 ( .A0(n35), .A1(n1286), .Z(gcm_dak_cmd_in_nxt[276]));
Q_MX02 U3360 ( .S(n90), .A0(gcm_dak_cmd_in[212]), .A1(gcm_dak_cmd_in[276]), .Z(n1286));
Q_AN02 U3361 ( .A0(n35), .A1(n1287), .Z(gcm_dak_cmd_in_nxt[275]));
Q_MX02 U3362 ( .S(n90), .A0(gcm_dak_cmd_in[211]), .A1(gcm_dak_cmd_in[275]), .Z(n1287));
Q_AN02 U3363 ( .A0(n35), .A1(n1288), .Z(gcm_dak_cmd_in_nxt[274]));
Q_MX02 U3364 ( .S(n90), .A0(gcm_dak_cmd_in[210]), .A1(gcm_dak_cmd_in[274]), .Z(n1288));
Q_AN02 U3365 ( .A0(n35), .A1(n1289), .Z(gcm_dak_cmd_in_nxt[273]));
Q_MX02 U3366 ( .S(n90), .A0(gcm_dak_cmd_in[209]), .A1(gcm_dak_cmd_in[273]), .Z(n1289));
Q_AN02 U3367 ( .A0(n35), .A1(n1290), .Z(gcm_dak_cmd_in_nxt[272]));
Q_MX02 U3368 ( .S(n90), .A0(gcm_dak_cmd_in[208]), .A1(gcm_dak_cmd_in[272]), .Z(n1290));
Q_AN02 U3369 ( .A0(n35), .A1(n1291), .Z(gcm_dak_cmd_in_nxt[271]));
Q_MX02 U3370 ( .S(n90), .A0(gcm_dak_cmd_in[207]), .A1(gcm_dak_cmd_in[271]), .Z(n1291));
Q_AN02 U3371 ( .A0(n35), .A1(n1292), .Z(gcm_dak_cmd_in_nxt[270]));
Q_MX02 U3372 ( .S(n90), .A0(gcm_dak_cmd_in[206]), .A1(gcm_dak_cmd_in[270]), .Z(n1292));
Q_AN02 U3373 ( .A0(n35), .A1(n1293), .Z(gcm_dak_cmd_in_nxt[269]));
Q_MX02 U3374 ( .S(n90), .A0(gcm_dak_cmd_in[205]), .A1(gcm_dak_cmd_in[269]), .Z(n1293));
Q_AN02 U3375 ( .A0(n35), .A1(n1294), .Z(gcm_dak_cmd_in_nxt[268]));
Q_MX02 U3376 ( .S(n90), .A0(gcm_dak_cmd_in[204]), .A1(gcm_dak_cmd_in[268]), .Z(n1294));
Q_AN02 U3377 ( .A0(n35), .A1(n1295), .Z(gcm_dak_cmd_in_nxt[267]));
Q_MX02 U3378 ( .S(n90), .A0(gcm_dak_cmd_in[203]), .A1(gcm_dak_cmd_in[267]), .Z(n1295));
Q_AN02 U3379 ( .A0(n35), .A1(n1296), .Z(gcm_dak_cmd_in_nxt[266]));
Q_MX02 U3380 ( .S(n90), .A0(gcm_dak_cmd_in[202]), .A1(gcm_dak_cmd_in[266]), .Z(n1296));
Q_AN02 U3381 ( .A0(n35), .A1(n1297), .Z(gcm_dak_cmd_in_nxt[265]));
Q_MX02 U3382 ( .S(n90), .A0(gcm_dak_cmd_in[201]), .A1(gcm_dak_cmd_in[265]), .Z(n1297));
Q_AN02 U3383 ( .A0(n35), .A1(n1298), .Z(gcm_dak_cmd_in_nxt[264]));
Q_MX02 U3384 ( .S(n90), .A0(gcm_dak_cmd_in[200]), .A1(gcm_dak_cmd_in[264]), .Z(n1298));
Q_AN02 U3385 ( .A0(n35), .A1(n1299), .Z(gcm_dak_cmd_in_nxt[263]));
Q_MX02 U3386 ( .S(n90), .A0(gcm_dak_cmd_in[199]), .A1(gcm_dak_cmd_in[263]), .Z(n1299));
Q_AN02 U3387 ( .A0(n35), .A1(n1300), .Z(gcm_dak_cmd_in_nxt[262]));
Q_MX02 U3388 ( .S(n90), .A0(gcm_dak_cmd_in[198]), .A1(gcm_dak_cmd_in[262]), .Z(n1300));
Q_AN02 U3389 ( .A0(n35), .A1(n1301), .Z(gcm_dak_cmd_in_nxt[261]));
Q_MX02 U3390 ( .S(n90), .A0(gcm_dak_cmd_in[197]), .A1(gcm_dak_cmd_in[261]), .Z(n1301));
Q_AN02 U3391 ( .A0(n35), .A1(n1302), .Z(gcm_dak_cmd_in_nxt[260]));
Q_MX02 U3392 ( .S(n90), .A0(gcm_dak_cmd_in[196]), .A1(gcm_dak_cmd_in[260]), .Z(n1302));
Q_AN02 U3393 ( .A0(n35), .A1(n1303), .Z(gcm_dak_cmd_in_nxt[259]));
Q_MX02 U3394 ( .S(n90), .A0(gcm_dak_cmd_in[195]), .A1(gcm_dak_cmd_in[259]), .Z(n1303));
Q_AN02 U3395 ( .A0(n35), .A1(n1304), .Z(gcm_dak_cmd_in_nxt[258]));
Q_MX02 U3396 ( .S(n90), .A0(gcm_dak_cmd_in[194]), .A1(gcm_dak_cmd_in[258]), .Z(n1304));
Q_AN02 U3397 ( .A0(n35), .A1(n1305), .Z(gcm_dak_cmd_in_nxt[257]));
Q_MX02 U3398 ( .S(n90), .A0(gcm_dak_cmd_in[193]), .A1(gcm_dak_cmd_in[257]), .Z(n1305));
Q_AN02 U3399 ( .A0(n35), .A1(n1306), .Z(gcm_dak_cmd_in_nxt[256]));
Q_MX02 U3400 ( .S(n90), .A0(gcm_dak_cmd_in[192]), .A1(gcm_dak_cmd_in[256]), .Z(n1306));
Q_AN02 U3401 ( .A0(n35), .A1(n1307), .Z(gcm_dak_cmd_in_nxt[255]));
Q_MX02 U3402 ( .S(n90), .A0(gcm_dak_cmd_in[191]), .A1(gcm_dak_cmd_in[255]), .Z(n1307));
Q_AN02 U3403 ( .A0(n35), .A1(n1308), .Z(gcm_dak_cmd_in_nxt[254]));
Q_MX02 U3404 ( .S(n90), .A0(gcm_dak_cmd_in[190]), .A1(gcm_dak_cmd_in[254]), .Z(n1308));
Q_AN02 U3405 ( .A0(n35), .A1(n1309), .Z(gcm_dak_cmd_in_nxt[253]));
Q_MX02 U3406 ( .S(n90), .A0(gcm_dak_cmd_in[189]), .A1(gcm_dak_cmd_in[253]), .Z(n1309));
Q_AN02 U3407 ( .A0(n35), .A1(n1310), .Z(gcm_dak_cmd_in_nxt[252]));
Q_MX02 U3408 ( .S(n90), .A0(gcm_dak_cmd_in[188]), .A1(gcm_dak_cmd_in[252]), .Z(n1310));
Q_AN02 U3409 ( .A0(n35), .A1(n1311), .Z(gcm_dak_cmd_in_nxt[251]));
Q_MX02 U3410 ( .S(n90), .A0(gcm_dak_cmd_in[187]), .A1(gcm_dak_cmd_in[251]), .Z(n1311));
Q_AN02 U3411 ( .A0(n35), .A1(n1312), .Z(gcm_dak_cmd_in_nxt[250]));
Q_MX02 U3412 ( .S(n90), .A0(gcm_dak_cmd_in[186]), .A1(gcm_dak_cmd_in[250]), .Z(n1312));
Q_AN02 U3413 ( .A0(n35), .A1(n1313), .Z(gcm_dak_cmd_in_nxt[249]));
Q_MX02 U3414 ( .S(n90), .A0(gcm_dak_cmd_in[185]), .A1(gcm_dak_cmd_in[249]), .Z(n1313));
Q_AN02 U3415 ( .A0(n35), .A1(n1314), .Z(gcm_dak_cmd_in_nxt[248]));
Q_MX02 U3416 ( .S(n90), .A0(gcm_dak_cmd_in[184]), .A1(gcm_dak_cmd_in[248]), .Z(n1314));
Q_AN02 U3417 ( .A0(n35), .A1(n1315), .Z(gcm_dak_cmd_in_nxt[247]));
Q_MX02 U3418 ( .S(n90), .A0(gcm_dak_cmd_in[183]), .A1(gcm_dak_cmd_in[247]), .Z(n1315));
Q_AN02 U3419 ( .A0(n35), .A1(n1316), .Z(gcm_dak_cmd_in_nxt[246]));
Q_MX02 U3420 ( .S(n90), .A0(gcm_dak_cmd_in[182]), .A1(gcm_dak_cmd_in[246]), .Z(n1316));
Q_AN02 U3421 ( .A0(n35), .A1(n1317), .Z(gcm_dak_cmd_in_nxt[245]));
Q_MX02 U3422 ( .S(n90), .A0(gcm_dak_cmd_in[181]), .A1(gcm_dak_cmd_in[245]), .Z(n1317));
Q_AN02 U3423 ( .A0(n35), .A1(n1318), .Z(gcm_dak_cmd_in_nxt[244]));
Q_MX02 U3424 ( .S(n90), .A0(gcm_dak_cmd_in[180]), .A1(gcm_dak_cmd_in[244]), .Z(n1318));
Q_AN02 U3425 ( .A0(n35), .A1(n1319), .Z(gcm_dak_cmd_in_nxt[243]));
Q_MX02 U3426 ( .S(n90), .A0(gcm_dak_cmd_in[179]), .A1(gcm_dak_cmd_in[243]), .Z(n1319));
Q_AN02 U3427 ( .A0(n35), .A1(n1320), .Z(gcm_dak_cmd_in_nxt[242]));
Q_MX02 U3428 ( .S(n90), .A0(gcm_dak_cmd_in[178]), .A1(gcm_dak_cmd_in[242]), .Z(n1320));
Q_AN02 U3429 ( .A0(n35), .A1(n1321), .Z(gcm_dak_cmd_in_nxt[241]));
Q_MX02 U3430 ( .S(n90), .A0(gcm_dak_cmd_in[177]), .A1(gcm_dak_cmd_in[241]), .Z(n1321));
Q_AN02 U3431 ( .A0(n35), .A1(n1322), .Z(gcm_dak_cmd_in_nxt[240]));
Q_MX02 U3432 ( .S(n90), .A0(gcm_dak_cmd_in[176]), .A1(gcm_dak_cmd_in[240]), .Z(n1322));
Q_AN02 U3433 ( .A0(n35), .A1(n1323), .Z(gcm_dak_cmd_in_nxt[239]));
Q_MX02 U3434 ( .S(n90), .A0(gcm_dak_cmd_in[175]), .A1(gcm_dak_cmd_in[239]), .Z(n1323));
Q_AN02 U3435 ( .A0(n35), .A1(n1324), .Z(gcm_dak_cmd_in_nxt[238]));
Q_MX02 U3436 ( .S(n90), .A0(gcm_dak_cmd_in[174]), .A1(gcm_dak_cmd_in[238]), .Z(n1324));
Q_AN02 U3437 ( .A0(n35), .A1(n1325), .Z(gcm_dak_cmd_in_nxt[237]));
Q_MX02 U3438 ( .S(n90), .A0(gcm_dak_cmd_in[173]), .A1(gcm_dak_cmd_in[237]), .Z(n1325));
Q_AN02 U3439 ( .A0(n35), .A1(n1326), .Z(gcm_dak_cmd_in_nxt[236]));
Q_MX02 U3440 ( .S(n90), .A0(gcm_dak_cmd_in[172]), .A1(gcm_dak_cmd_in[236]), .Z(n1326));
Q_AN02 U3441 ( .A0(n35), .A1(n1327), .Z(gcm_dak_cmd_in_nxt[235]));
Q_MX02 U3442 ( .S(n90), .A0(gcm_dak_cmd_in[171]), .A1(gcm_dak_cmd_in[235]), .Z(n1327));
Q_AN02 U3443 ( .A0(n35), .A1(n1328), .Z(gcm_dak_cmd_in_nxt[234]));
Q_MX02 U3444 ( .S(n90), .A0(gcm_dak_cmd_in[170]), .A1(gcm_dak_cmd_in[234]), .Z(n1328));
Q_AN02 U3445 ( .A0(n35), .A1(n1329), .Z(gcm_dak_cmd_in_nxt[233]));
Q_MX02 U3446 ( .S(n90), .A0(gcm_dak_cmd_in[169]), .A1(gcm_dak_cmd_in[233]), .Z(n1329));
Q_AN02 U3447 ( .A0(n35), .A1(n1330), .Z(gcm_dak_cmd_in_nxt[232]));
Q_MX02 U3448 ( .S(n90), .A0(gcm_dak_cmd_in[168]), .A1(gcm_dak_cmd_in[232]), .Z(n1330));
Q_AN02 U3449 ( .A0(n35), .A1(n1331), .Z(gcm_dak_cmd_in_nxt[231]));
Q_MX02 U3450 ( .S(n90), .A0(gcm_dak_cmd_in[167]), .A1(gcm_dak_cmd_in[231]), .Z(n1331));
Q_AN02 U3451 ( .A0(n35), .A1(n1332), .Z(gcm_dak_cmd_in_nxt[230]));
Q_MX02 U3452 ( .S(n90), .A0(gcm_dak_cmd_in[166]), .A1(gcm_dak_cmd_in[230]), .Z(n1332));
Q_AN02 U3453 ( .A0(n35), .A1(n1333), .Z(gcm_dak_cmd_in_nxt[229]));
Q_MX02 U3454 ( .S(n90), .A0(gcm_dak_cmd_in[165]), .A1(gcm_dak_cmd_in[229]), .Z(n1333));
Q_AN02 U3455 ( .A0(n35), .A1(n1334), .Z(gcm_dak_cmd_in_nxt[228]));
Q_MX02 U3456 ( .S(n90), .A0(gcm_dak_cmd_in[164]), .A1(gcm_dak_cmd_in[228]), .Z(n1334));
Q_AN02 U3457 ( .A0(n35), .A1(n1335), .Z(gcm_dak_cmd_in_nxt[227]));
Q_MX02 U3458 ( .S(n90), .A0(gcm_dak_cmd_in[163]), .A1(gcm_dak_cmd_in[227]), .Z(n1335));
Q_AN02 U3459 ( .A0(n35), .A1(n1336), .Z(gcm_dak_cmd_in_nxt[226]));
Q_MX02 U3460 ( .S(n90), .A0(gcm_dak_cmd_in[162]), .A1(gcm_dak_cmd_in[226]), .Z(n1336));
Q_AN02 U3461 ( .A0(n35), .A1(n1337), .Z(gcm_dak_cmd_in_nxt[225]));
Q_MX02 U3462 ( .S(n90), .A0(gcm_dak_cmd_in[161]), .A1(gcm_dak_cmd_in[225]), .Z(n1337));
Q_AN02 U3463 ( .A0(n35), .A1(n1338), .Z(gcm_dak_cmd_in_nxt[224]));
Q_MX02 U3464 ( .S(n90), .A0(gcm_dak_cmd_in[160]), .A1(gcm_dak_cmd_in[224]), .Z(n1338));
Q_AN02 U3465 ( .A0(n35), .A1(n1339), .Z(gcm_dak_cmd_in_nxt[223]));
Q_MX02 U3466 ( .S(n90), .A0(gcm_dak_cmd_in[159]), .A1(gcm_dak_cmd_in[223]), .Z(n1339));
Q_AN02 U3467 ( .A0(n35), .A1(n1340), .Z(gcm_dak_cmd_in_nxt[222]));
Q_MX02 U3468 ( .S(n90), .A0(gcm_dak_cmd_in[158]), .A1(gcm_dak_cmd_in[222]), .Z(n1340));
Q_AN02 U3469 ( .A0(n35), .A1(n1341), .Z(gcm_dak_cmd_in_nxt[221]));
Q_MX02 U3470 ( .S(n90), .A0(gcm_dak_cmd_in[157]), .A1(gcm_dak_cmd_in[221]), .Z(n1341));
Q_AN02 U3471 ( .A0(n35), .A1(n1342), .Z(gcm_dak_cmd_in_nxt[220]));
Q_MX02 U3472 ( .S(n90), .A0(gcm_dak_cmd_in[156]), .A1(gcm_dak_cmd_in[220]), .Z(n1342));
Q_AN02 U3473 ( .A0(n35), .A1(n1343), .Z(gcm_dak_cmd_in_nxt[219]));
Q_MX02 U3474 ( .S(n90), .A0(gcm_dak_cmd_in[155]), .A1(gcm_dak_cmd_in[219]), .Z(n1343));
Q_AN02 U3475 ( .A0(n35), .A1(n1344), .Z(gcm_dak_cmd_in_nxt[218]));
Q_MX02 U3476 ( .S(n90), .A0(gcm_dak_cmd_in[154]), .A1(gcm_dak_cmd_in[218]), .Z(n1344));
Q_AN02 U3477 ( .A0(n35), .A1(n1345), .Z(gcm_dak_cmd_in_nxt[217]));
Q_MX02 U3478 ( .S(n90), .A0(gcm_dak_cmd_in[153]), .A1(gcm_dak_cmd_in[217]), .Z(n1345));
Q_AN02 U3479 ( .A0(n35), .A1(n1346), .Z(gcm_dak_cmd_in_nxt[216]));
Q_MX02 U3480 ( .S(n90), .A0(gcm_dak_cmd_in[152]), .A1(gcm_dak_cmd_in[216]), .Z(n1346));
Q_AN02 U3481 ( .A0(n35), .A1(n1347), .Z(gcm_dak_cmd_in_nxt[215]));
Q_MX02 U3482 ( .S(n90), .A0(gcm_dak_cmd_in[151]), .A1(gcm_dak_cmd_in[215]), .Z(n1347));
Q_AN02 U3483 ( .A0(n35), .A1(n1348), .Z(gcm_dak_cmd_in_nxt[214]));
Q_MX02 U3484 ( .S(n90), .A0(gcm_dak_cmd_in[150]), .A1(gcm_dak_cmd_in[214]), .Z(n1348));
Q_AN02 U3485 ( .A0(n35), .A1(n1349), .Z(gcm_dak_cmd_in_nxt[213]));
Q_MX02 U3486 ( .S(n90), .A0(gcm_dak_cmd_in[149]), .A1(gcm_dak_cmd_in[213]), .Z(n1349));
Q_AN02 U3487 ( .A0(n35), .A1(n1350), .Z(gcm_dak_cmd_in_nxt[212]));
Q_MX02 U3488 ( .S(n90), .A0(gcm_dak_cmd_in[148]), .A1(gcm_dak_cmd_in[212]), .Z(n1350));
Q_AN02 U3489 ( .A0(n35), .A1(n1351), .Z(gcm_dak_cmd_in_nxt[211]));
Q_MX02 U3490 ( .S(n90), .A0(gcm_dak_cmd_in[147]), .A1(gcm_dak_cmd_in[211]), .Z(n1351));
Q_AN02 U3491 ( .A0(n35), .A1(n1352), .Z(gcm_dak_cmd_in_nxt[210]));
Q_MX02 U3492 ( .S(n90), .A0(gcm_dak_cmd_in[146]), .A1(gcm_dak_cmd_in[210]), .Z(n1352));
Q_AN02 U3493 ( .A0(n35), .A1(n1353), .Z(gcm_dak_cmd_in_nxt[209]));
Q_MX02 U3494 ( .S(n90), .A0(gcm_dak_cmd_in[145]), .A1(gcm_dak_cmd_in[209]), .Z(n1353));
Q_AN02 U3495 ( .A0(n35), .A1(n1354), .Z(gcm_dak_cmd_in_nxt[208]));
Q_MX02 U3496 ( .S(n90), .A0(gcm_dak_cmd_in[144]), .A1(gcm_dak_cmd_in[208]), .Z(n1354));
Q_AN02 U3497 ( .A0(n35), .A1(n1355), .Z(gcm_dak_cmd_in_nxt[207]));
Q_MX02 U3498 ( .S(n90), .A0(gcm_dak_cmd_in[143]), .A1(gcm_dak_cmd_in[207]), .Z(n1355));
Q_AN02 U3499 ( .A0(n35), .A1(n1356), .Z(gcm_dak_cmd_in_nxt[206]));
Q_MX02 U3500 ( .S(n90), .A0(gcm_dak_cmd_in[142]), .A1(gcm_dak_cmd_in[206]), .Z(n1356));
Q_AN02 U3501 ( .A0(n35), .A1(n1357), .Z(gcm_dak_cmd_in_nxt[205]));
Q_MX02 U3502 ( .S(n90), .A0(gcm_dak_cmd_in[141]), .A1(gcm_dak_cmd_in[205]), .Z(n1357));
Q_AN02 U3503 ( .A0(n35), .A1(n1358), .Z(gcm_dak_cmd_in_nxt[204]));
Q_MX02 U3504 ( .S(n90), .A0(gcm_dak_cmd_in[140]), .A1(gcm_dak_cmd_in[204]), .Z(n1358));
Q_AN02 U3505 ( .A0(n35), .A1(n1359), .Z(gcm_dak_cmd_in_nxt[203]));
Q_MX02 U3506 ( .S(n90), .A0(gcm_dak_cmd_in[139]), .A1(gcm_dak_cmd_in[203]), .Z(n1359));
Q_AN02 U3507 ( .A0(n35), .A1(n1360), .Z(gcm_dak_cmd_in_nxt[202]));
Q_MX02 U3508 ( .S(n90), .A0(gcm_dak_cmd_in[138]), .A1(gcm_dak_cmd_in[202]), .Z(n1360));
Q_AN02 U3509 ( .A0(n35), .A1(n1361), .Z(gcm_dak_cmd_in_nxt[201]));
Q_MX02 U3510 ( .S(n90), .A0(gcm_dak_cmd_in[137]), .A1(gcm_dak_cmd_in[201]), .Z(n1361));
Q_AN02 U3511 ( .A0(n35), .A1(n1362), .Z(gcm_dak_cmd_in_nxt[200]));
Q_MX02 U3512 ( .S(n90), .A0(gcm_dak_cmd_in[136]), .A1(gcm_dak_cmd_in[200]), .Z(n1362));
Q_AN02 U3513 ( .A0(n35), .A1(n1363), .Z(gcm_dak_cmd_in_nxt[199]));
Q_MX02 U3514 ( .S(n90), .A0(gcm_dak_cmd_in[135]), .A1(gcm_dak_cmd_in[199]), .Z(n1363));
Q_AN02 U3515 ( .A0(n35), .A1(n1364), .Z(gcm_dak_cmd_in_nxt[198]));
Q_MX02 U3516 ( .S(n90), .A0(gcm_dak_cmd_in[134]), .A1(gcm_dak_cmd_in[198]), .Z(n1364));
Q_AN02 U3517 ( .A0(n35), .A1(n1365), .Z(gcm_dak_cmd_in_nxt[197]));
Q_MX02 U3518 ( .S(n90), .A0(gcm_dak_cmd_in[133]), .A1(gcm_dak_cmd_in[197]), .Z(n1365));
Q_AN02 U3519 ( .A0(n35), .A1(n1366), .Z(gcm_dak_cmd_in_nxt[196]));
Q_MX02 U3520 ( .S(n90), .A0(gcm_dak_cmd_in[132]), .A1(gcm_dak_cmd_in[196]), .Z(n1366));
Q_AN02 U3521 ( .A0(n35), .A1(n1367), .Z(gcm_dak_cmd_in_nxt[195]));
Q_MX02 U3522 ( .S(n90), .A0(gcm_dak_cmd_in[131]), .A1(gcm_dak_cmd_in[195]), .Z(n1367));
Q_AN02 U3523 ( .A0(n35), .A1(n1368), .Z(gcm_dak_cmd_in_nxt[194]));
Q_MX02 U3524 ( .S(n90), .A0(gcm_dak_cmd_in[130]), .A1(gcm_dak_cmd_in[194]), .Z(n1368));
Q_AN02 U3525 ( .A0(n35), .A1(n1369), .Z(gcm_dak_cmd_in_nxt[193]));
Q_MX02 U3526 ( .S(n90), .A0(gcm_dak_cmd_in[129]), .A1(gcm_dak_cmd_in[193]), .Z(n1369));
Q_AN02 U3527 ( .A0(n35), .A1(n1370), .Z(gcm_dak_cmd_in_nxt[192]));
Q_MX02 U3528 ( .S(n90), .A0(gcm_dak_cmd_in[128]), .A1(gcm_dak_cmd_in[192]), .Z(n1370));
Q_AN02 U3529 ( .A0(n35), .A1(n1371), .Z(gcm_dak_cmd_in_nxt[191]));
Q_MX02 U3530 ( .S(n90), .A0(gcm_dak_cmd_in[127]), .A1(gcm_dak_cmd_in[191]), .Z(n1371));
Q_AN02 U3531 ( .A0(n35), .A1(n1372), .Z(gcm_dak_cmd_in_nxt[190]));
Q_MX02 U3532 ( .S(n90), .A0(gcm_dak_cmd_in[126]), .A1(gcm_dak_cmd_in[190]), .Z(n1372));
Q_AN02 U3533 ( .A0(n35), .A1(n1373), .Z(gcm_dak_cmd_in_nxt[189]));
Q_MX02 U3534 ( .S(n90), .A0(gcm_dak_cmd_in[125]), .A1(gcm_dak_cmd_in[189]), .Z(n1373));
Q_AN02 U3535 ( .A0(n35), .A1(n1374), .Z(gcm_dak_cmd_in_nxt[188]));
Q_MX02 U3536 ( .S(n90), .A0(gcm_dak_cmd_in[124]), .A1(gcm_dak_cmd_in[188]), .Z(n1374));
Q_AN02 U3537 ( .A0(n35), .A1(n1375), .Z(gcm_dak_cmd_in_nxt[187]));
Q_MX02 U3538 ( .S(n90), .A0(gcm_dak_cmd_in[123]), .A1(gcm_dak_cmd_in[187]), .Z(n1375));
Q_AN02 U3539 ( .A0(n35), .A1(n1376), .Z(gcm_dak_cmd_in_nxt[186]));
Q_MX02 U3540 ( .S(n90), .A0(gcm_dak_cmd_in[122]), .A1(gcm_dak_cmd_in[186]), .Z(n1376));
Q_AN02 U3541 ( .A0(n35), .A1(n1377), .Z(gcm_dak_cmd_in_nxt[185]));
Q_MX02 U3542 ( .S(n90), .A0(gcm_dak_cmd_in[121]), .A1(gcm_dak_cmd_in[185]), .Z(n1377));
Q_AN02 U3543 ( .A0(n35), .A1(n1378), .Z(gcm_dak_cmd_in_nxt[184]));
Q_MX02 U3544 ( .S(n90), .A0(gcm_dak_cmd_in[120]), .A1(gcm_dak_cmd_in[184]), .Z(n1378));
Q_AN02 U3545 ( .A0(n35), .A1(n1379), .Z(gcm_dak_cmd_in_nxt[183]));
Q_MX02 U3546 ( .S(n90), .A0(gcm_dak_cmd_in[119]), .A1(gcm_dak_cmd_in[183]), .Z(n1379));
Q_AN02 U3547 ( .A0(n35), .A1(n1380), .Z(gcm_dak_cmd_in_nxt[182]));
Q_MX02 U3548 ( .S(n90), .A0(gcm_dak_cmd_in[118]), .A1(gcm_dak_cmd_in[182]), .Z(n1380));
Q_AN02 U3549 ( .A0(n35), .A1(n1381), .Z(gcm_dak_cmd_in_nxt[181]));
Q_MX02 U3550 ( .S(n90), .A0(gcm_dak_cmd_in[117]), .A1(gcm_dak_cmd_in[181]), .Z(n1381));
Q_AN02 U3551 ( .A0(n35), .A1(n1382), .Z(gcm_dak_cmd_in_nxt[180]));
Q_MX02 U3552 ( .S(n90), .A0(gcm_dak_cmd_in[116]), .A1(gcm_dak_cmd_in[180]), .Z(n1382));
Q_AN02 U3553 ( .A0(n35), .A1(n1383), .Z(gcm_dak_cmd_in_nxt[179]));
Q_MX02 U3554 ( .S(n90), .A0(gcm_dak_cmd_in[115]), .A1(gcm_dak_cmd_in[179]), .Z(n1383));
Q_AN02 U3555 ( .A0(n35), .A1(n1384), .Z(gcm_dak_cmd_in_nxt[178]));
Q_MX02 U3556 ( .S(n90), .A0(gcm_dak_cmd_in[114]), .A1(gcm_dak_cmd_in[178]), .Z(n1384));
Q_AN02 U3557 ( .A0(n35), .A1(n1385), .Z(gcm_dak_cmd_in_nxt[177]));
Q_MX02 U3558 ( .S(n90), .A0(gcm_dak_cmd_in[113]), .A1(gcm_dak_cmd_in[177]), .Z(n1385));
Q_AN02 U3559 ( .A0(n35), .A1(n1386), .Z(gcm_dak_cmd_in_nxt[176]));
Q_MX02 U3560 ( .S(n90), .A0(gcm_dak_cmd_in[112]), .A1(gcm_dak_cmd_in[176]), .Z(n1386));
Q_AN02 U3561 ( .A0(n35), .A1(n1387), .Z(gcm_dak_cmd_in_nxt[175]));
Q_MX02 U3562 ( .S(n90), .A0(gcm_dak_cmd_in[111]), .A1(gcm_dak_cmd_in[175]), .Z(n1387));
Q_AN02 U3563 ( .A0(n35), .A1(n1388), .Z(gcm_dak_cmd_in_nxt[174]));
Q_MX02 U3564 ( .S(n90), .A0(gcm_dak_cmd_in[110]), .A1(gcm_dak_cmd_in[174]), .Z(n1388));
Q_AN02 U3565 ( .A0(n35), .A1(n1389), .Z(gcm_dak_cmd_in_nxt[173]));
Q_MX02 U3566 ( .S(n90), .A0(gcm_dak_cmd_in[109]), .A1(gcm_dak_cmd_in[173]), .Z(n1389));
Q_AN02 U3567 ( .A0(n35), .A1(n1390), .Z(gcm_dak_cmd_in_nxt[172]));
Q_MX02 U3568 ( .S(n90), .A0(gcm_dak_cmd_in[108]), .A1(gcm_dak_cmd_in[172]), .Z(n1390));
Q_AN02 U3569 ( .A0(n35), .A1(n1391), .Z(gcm_dak_cmd_in_nxt[171]));
Q_MX02 U3570 ( .S(n90), .A0(gcm_dak_cmd_in[107]), .A1(gcm_dak_cmd_in[171]), .Z(n1391));
Q_AN02 U3571 ( .A0(n35), .A1(n1392), .Z(gcm_dak_cmd_in_nxt[170]));
Q_MX02 U3572 ( .S(n90), .A0(gcm_dak_cmd_in[106]), .A1(gcm_dak_cmd_in[170]), .Z(n1392));
Q_AN02 U3573 ( .A0(n35), .A1(n1393), .Z(gcm_dak_cmd_in_nxt[169]));
Q_MX02 U3574 ( .S(n90), .A0(gcm_dak_cmd_in[105]), .A1(gcm_dak_cmd_in[169]), .Z(n1393));
Q_AN02 U3575 ( .A0(n35), .A1(n1394), .Z(gcm_dak_cmd_in_nxt[168]));
Q_MX02 U3576 ( .S(n90), .A0(gcm_dak_cmd_in[104]), .A1(gcm_dak_cmd_in[168]), .Z(n1394));
Q_AN02 U3577 ( .A0(n35), .A1(n1395), .Z(gcm_dak_cmd_in_nxt[167]));
Q_MX02 U3578 ( .S(n90), .A0(gcm_dak_cmd_in[103]), .A1(gcm_dak_cmd_in[167]), .Z(n1395));
Q_AN02 U3579 ( .A0(n35), .A1(n1396), .Z(gcm_dak_cmd_in_nxt[166]));
Q_MX02 U3580 ( .S(n90), .A0(gcm_dak_cmd_in[102]), .A1(gcm_dak_cmd_in[166]), .Z(n1396));
Q_AN02 U3581 ( .A0(n35), .A1(n1397), .Z(gcm_dak_cmd_in_nxt[165]));
Q_MX02 U3582 ( .S(n90), .A0(gcm_dak_cmd_in[101]), .A1(gcm_dak_cmd_in[165]), .Z(n1397));
Q_AN02 U3583 ( .A0(n35), .A1(n1398), .Z(gcm_dak_cmd_in_nxt[164]));
Q_MX02 U3584 ( .S(n90), .A0(gcm_dak_cmd_in[100]), .A1(gcm_dak_cmd_in[164]), .Z(n1398));
Q_AN02 U3585 ( .A0(n35), .A1(n1399), .Z(gcm_dak_cmd_in_nxt[163]));
Q_MX02 U3586 ( .S(n90), .A0(gcm_dak_cmd_in[99]), .A1(gcm_dak_cmd_in[163]), .Z(n1399));
Q_AN02 U3587 ( .A0(n35), .A1(n1400), .Z(gcm_dak_cmd_in_nxt[162]));
Q_MX02 U3588 ( .S(n90), .A0(kme_internal_out[63]), .A1(gcm_dak_cmd_in[162]), .Z(n1400));
Q_AN02 U3589 ( .A0(n35), .A1(n1401), .Z(gcm_dak_cmd_in_nxt[161]));
Q_MX02 U3590 ( .S(n90), .A0(kme_internal_out[62]), .A1(gcm_dak_cmd_in[161]), .Z(n1401));
Q_AN02 U3591 ( .A0(n35), .A1(n1402), .Z(gcm_dak_cmd_in_nxt[160]));
Q_MX02 U3592 ( .S(n90), .A0(kme_internal_out[61]), .A1(gcm_dak_cmd_in[160]), .Z(n1402));
Q_AN02 U3593 ( .A0(n35), .A1(n1403), .Z(gcm_dak_cmd_in_nxt[159]));
Q_MX02 U3594 ( .S(n90), .A0(kme_internal_out[60]), .A1(gcm_dak_cmd_in[159]), .Z(n1403));
Q_AN02 U3595 ( .A0(n35), .A1(n1404), .Z(gcm_dak_cmd_in_nxt[158]));
Q_MX02 U3596 ( .S(n90), .A0(kme_internal_out[59]), .A1(gcm_dak_cmd_in[158]), .Z(n1404));
Q_AN02 U3597 ( .A0(n35), .A1(n1405), .Z(gcm_dak_cmd_in_nxt[157]));
Q_MX02 U3598 ( .S(n90), .A0(kme_internal_out[58]), .A1(gcm_dak_cmd_in[157]), .Z(n1405));
Q_AN02 U3599 ( .A0(n35), .A1(n1406), .Z(gcm_dak_cmd_in_nxt[156]));
Q_MX02 U3600 ( .S(n90), .A0(kme_internal_out[57]), .A1(gcm_dak_cmd_in[156]), .Z(n1406));
Q_AN02 U3601 ( .A0(n35), .A1(n1407), .Z(gcm_dak_cmd_in_nxt[155]));
Q_MX02 U3602 ( .S(n90), .A0(kme_internal_out[56]), .A1(gcm_dak_cmd_in[155]), .Z(n1407));
Q_AN02 U3603 ( .A0(n35), .A1(n1408), .Z(gcm_dak_cmd_in_nxt[154]));
Q_MX02 U3604 ( .S(n90), .A0(kme_internal_out[55]), .A1(gcm_dak_cmd_in[154]), .Z(n1408));
Q_AN02 U3605 ( .A0(n35), .A1(n1409), .Z(gcm_dak_cmd_in_nxt[153]));
Q_MX02 U3606 ( .S(n90), .A0(kme_internal_out[54]), .A1(gcm_dak_cmd_in[153]), .Z(n1409));
Q_AN02 U3607 ( .A0(n35), .A1(n1410), .Z(gcm_dak_cmd_in_nxt[152]));
Q_MX02 U3608 ( .S(n90), .A0(kme_internal_out[53]), .A1(gcm_dak_cmd_in[152]), .Z(n1410));
Q_AN02 U3609 ( .A0(n35), .A1(n1411), .Z(gcm_dak_cmd_in_nxt[151]));
Q_MX02 U3610 ( .S(n90), .A0(kme_internal_out[52]), .A1(gcm_dak_cmd_in[151]), .Z(n1411));
Q_AN02 U3611 ( .A0(n35), .A1(n1412), .Z(gcm_dak_cmd_in_nxt[150]));
Q_MX02 U3612 ( .S(n90), .A0(kme_internal_out[51]), .A1(gcm_dak_cmd_in[150]), .Z(n1412));
Q_AN02 U3613 ( .A0(n35), .A1(n1413), .Z(gcm_dak_cmd_in_nxt[149]));
Q_MX02 U3614 ( .S(n90), .A0(kme_internal_out[50]), .A1(gcm_dak_cmd_in[149]), .Z(n1413));
Q_AN02 U3615 ( .A0(n35), .A1(n1414), .Z(gcm_dak_cmd_in_nxt[148]));
Q_MX02 U3616 ( .S(n90), .A0(kme_internal_out[49]), .A1(gcm_dak_cmd_in[148]), .Z(n1414));
Q_AN02 U3617 ( .A0(n35), .A1(n1415), .Z(gcm_dak_cmd_in_nxt[147]));
Q_MX02 U3618 ( .S(n90), .A0(kme_internal_out[48]), .A1(gcm_dak_cmd_in[147]), .Z(n1415));
Q_AN02 U3619 ( .A0(n35), .A1(n1416), .Z(gcm_dak_cmd_in_nxt[146]));
Q_MX02 U3620 ( .S(n90), .A0(kme_internal_out[47]), .A1(gcm_dak_cmd_in[146]), .Z(n1416));
Q_AN02 U3621 ( .A0(n35), .A1(n1417), .Z(gcm_dak_cmd_in_nxt[145]));
Q_MX02 U3622 ( .S(n90), .A0(kme_internal_out[46]), .A1(gcm_dak_cmd_in[145]), .Z(n1417));
Q_AN02 U3623 ( .A0(n35), .A1(n1418), .Z(gcm_dak_cmd_in_nxt[144]));
Q_MX02 U3624 ( .S(n90), .A0(kme_internal_out[45]), .A1(gcm_dak_cmd_in[144]), .Z(n1418));
Q_AN02 U3625 ( .A0(n35), .A1(n1419), .Z(gcm_dak_cmd_in_nxt[143]));
Q_MX02 U3626 ( .S(n90), .A0(kme_internal_out[44]), .A1(gcm_dak_cmd_in[143]), .Z(n1419));
Q_AN02 U3627 ( .A0(n35), .A1(n1420), .Z(gcm_dak_cmd_in_nxt[142]));
Q_MX02 U3628 ( .S(n90), .A0(kme_internal_out[43]), .A1(gcm_dak_cmd_in[142]), .Z(n1420));
Q_AN02 U3629 ( .A0(n35), .A1(n1421), .Z(gcm_dak_cmd_in_nxt[141]));
Q_MX02 U3630 ( .S(n90), .A0(kme_internal_out[42]), .A1(gcm_dak_cmd_in[141]), .Z(n1421));
Q_AN02 U3631 ( .A0(n35), .A1(n1422), .Z(gcm_dak_cmd_in_nxt[140]));
Q_MX02 U3632 ( .S(n90), .A0(kme_internal_out[41]), .A1(gcm_dak_cmd_in[140]), .Z(n1422));
Q_AN02 U3633 ( .A0(n35), .A1(n1423), .Z(gcm_dak_cmd_in_nxt[139]));
Q_MX02 U3634 ( .S(n90), .A0(kme_internal_out[40]), .A1(gcm_dak_cmd_in[139]), .Z(n1423));
Q_AN02 U3635 ( .A0(n35), .A1(n1424), .Z(gcm_dak_cmd_in_nxt[138]));
Q_MX02 U3636 ( .S(n90), .A0(kme_internal_out[39]), .A1(gcm_dak_cmd_in[138]), .Z(n1424));
Q_AN02 U3637 ( .A0(n35), .A1(n1425), .Z(gcm_dak_cmd_in_nxt[137]));
Q_MX02 U3638 ( .S(n90), .A0(kme_internal_out[38]), .A1(gcm_dak_cmd_in[137]), .Z(n1425));
Q_AN02 U3639 ( .A0(n35), .A1(n1426), .Z(gcm_dak_cmd_in_nxt[136]));
Q_MX02 U3640 ( .S(n90), .A0(kme_internal_out[37]), .A1(gcm_dak_cmd_in[136]), .Z(n1426));
Q_AN02 U3641 ( .A0(n35), .A1(n1427), .Z(gcm_dak_cmd_in_nxt[135]));
Q_MX02 U3642 ( .S(n90), .A0(kme_internal_out[36]), .A1(gcm_dak_cmd_in[135]), .Z(n1427));
Q_AN02 U3643 ( .A0(n35), .A1(n1428), .Z(gcm_dak_cmd_in_nxt[134]));
Q_MX02 U3644 ( .S(n90), .A0(kme_internal_out[35]), .A1(gcm_dak_cmd_in[134]), .Z(n1428));
Q_AN02 U3645 ( .A0(n35), .A1(n1429), .Z(gcm_dak_cmd_in_nxt[133]));
Q_MX02 U3646 ( .S(n90), .A0(kme_internal_out[34]), .A1(gcm_dak_cmd_in[133]), .Z(n1429));
Q_AN02 U3647 ( .A0(n35), .A1(n1430), .Z(gcm_dak_cmd_in_nxt[132]));
Q_MX02 U3648 ( .S(n90), .A0(kme_internal_out[33]), .A1(gcm_dak_cmd_in[132]), .Z(n1430));
Q_AN02 U3649 ( .A0(n35), .A1(n1431), .Z(gcm_dak_cmd_in_nxt[131]));
Q_MX02 U3650 ( .S(n90), .A0(kme_internal_out[32]), .A1(gcm_dak_cmd_in[131]), .Z(n1431));
Q_AN02 U3651 ( .A0(n35), .A1(n1432), .Z(gcm_dak_cmd_in_nxt[130]));
Q_MX02 U3652 ( .S(n90), .A0(kme_internal_out[31]), .A1(gcm_dak_cmd_in[130]), .Z(n1432));
Q_AN02 U3653 ( .A0(n35), .A1(n1433), .Z(gcm_dak_cmd_in_nxt[129]));
Q_MX02 U3654 ( .S(n90), .A0(kme_internal_out[30]), .A1(gcm_dak_cmd_in[129]), .Z(n1433));
Q_AN02 U3655 ( .A0(n35), .A1(n1434), .Z(gcm_dak_cmd_in_nxt[128]));
Q_MX02 U3656 ( .S(n90), .A0(kme_internal_out[29]), .A1(gcm_dak_cmd_in[128]), .Z(n1434));
Q_AN02 U3657 ( .A0(n35), .A1(n1435), .Z(gcm_dak_cmd_in_nxt[127]));
Q_MX02 U3658 ( .S(n90), .A0(kme_internal_out[28]), .A1(gcm_dak_cmd_in[127]), .Z(n1435));
Q_AN02 U3659 ( .A0(n35), .A1(n1436), .Z(gcm_dak_cmd_in_nxt[126]));
Q_MX02 U3660 ( .S(n90), .A0(kme_internal_out[27]), .A1(gcm_dak_cmd_in[126]), .Z(n1436));
Q_AN02 U3661 ( .A0(n35), .A1(n1437), .Z(gcm_dak_cmd_in_nxt[125]));
Q_MX02 U3662 ( .S(n90), .A0(kme_internal_out[26]), .A1(gcm_dak_cmd_in[125]), .Z(n1437));
Q_AN02 U3663 ( .A0(n35), .A1(n1438), .Z(gcm_dak_cmd_in_nxt[124]));
Q_MX02 U3664 ( .S(n90), .A0(kme_internal_out[25]), .A1(gcm_dak_cmd_in[124]), .Z(n1438));
Q_AN02 U3665 ( .A0(n35), .A1(n1439), .Z(gcm_dak_cmd_in_nxt[123]));
Q_MX02 U3666 ( .S(n90), .A0(kme_internal_out[24]), .A1(gcm_dak_cmd_in[123]), .Z(n1439));
Q_AN02 U3667 ( .A0(n35), .A1(n1440), .Z(gcm_dak_cmd_in_nxt[122]));
Q_MX02 U3668 ( .S(n90), .A0(kme_internal_out[23]), .A1(gcm_dak_cmd_in[122]), .Z(n1440));
Q_AN02 U3669 ( .A0(n35), .A1(n1441), .Z(gcm_dak_cmd_in_nxt[121]));
Q_MX02 U3670 ( .S(n90), .A0(kme_internal_out[22]), .A1(gcm_dak_cmd_in[121]), .Z(n1441));
Q_AN02 U3671 ( .A0(n35), .A1(n1442), .Z(gcm_dak_cmd_in_nxt[120]));
Q_MX02 U3672 ( .S(n90), .A0(kme_internal_out[21]), .A1(gcm_dak_cmd_in[120]), .Z(n1442));
Q_AN02 U3673 ( .A0(n35), .A1(n1443), .Z(gcm_dak_cmd_in_nxt[119]));
Q_MX02 U3674 ( .S(n90), .A0(kme_internal_out[20]), .A1(gcm_dak_cmd_in[119]), .Z(n1443));
Q_AN02 U3675 ( .A0(n35), .A1(n1444), .Z(gcm_dak_cmd_in_nxt[118]));
Q_MX02 U3676 ( .S(n90), .A0(kme_internal_out[19]), .A1(gcm_dak_cmd_in[118]), .Z(n1444));
Q_AN02 U3677 ( .A0(n35), .A1(n1445), .Z(gcm_dak_cmd_in_nxt[117]));
Q_MX02 U3678 ( .S(n90), .A0(kme_internal_out[18]), .A1(gcm_dak_cmd_in[117]), .Z(n1445));
Q_AN02 U3679 ( .A0(n35), .A1(n1446), .Z(gcm_dak_cmd_in_nxt[116]));
Q_MX02 U3680 ( .S(n90), .A0(kme_internal_out[17]), .A1(gcm_dak_cmd_in[116]), .Z(n1446));
Q_AN02 U3681 ( .A0(n35), .A1(n1447), .Z(gcm_dak_cmd_in_nxt[115]));
Q_MX02 U3682 ( .S(n90), .A0(kme_internal_out[16]), .A1(gcm_dak_cmd_in[115]), .Z(n1447));
Q_AN02 U3683 ( .A0(n35), .A1(n1448), .Z(gcm_dak_cmd_in_nxt[114]));
Q_MX02 U3684 ( .S(n90), .A0(kme_internal_out[15]), .A1(gcm_dak_cmd_in[114]), .Z(n1448));
Q_AN02 U3685 ( .A0(n35), .A1(n1449), .Z(gcm_dak_cmd_in_nxt[113]));
Q_MX02 U3686 ( .S(n90), .A0(kme_internal_out[14]), .A1(gcm_dak_cmd_in[113]), .Z(n1449));
Q_AN02 U3687 ( .A0(n35), .A1(n1450), .Z(gcm_dak_cmd_in_nxt[112]));
Q_MX02 U3688 ( .S(n90), .A0(kme_internal_out[13]), .A1(gcm_dak_cmd_in[112]), .Z(n1450));
Q_AN02 U3689 ( .A0(n35), .A1(n1451), .Z(gcm_dak_cmd_in_nxt[111]));
Q_MX02 U3690 ( .S(n90), .A0(kme_internal_out[12]), .A1(gcm_dak_cmd_in[111]), .Z(n1451));
Q_AN02 U3691 ( .A0(n35), .A1(n1452), .Z(gcm_dak_cmd_in_nxt[110]));
Q_MX02 U3692 ( .S(n90), .A0(kme_internal_out[11]), .A1(gcm_dak_cmd_in[110]), .Z(n1452));
Q_AN02 U3693 ( .A0(n35), .A1(n1453), .Z(gcm_dak_cmd_in_nxt[109]));
Q_MX02 U3694 ( .S(n90), .A0(kme_internal_out[10]), .A1(gcm_dak_cmd_in[109]), .Z(n1453));
Q_AN02 U3695 ( .A0(n35), .A1(n1454), .Z(gcm_dak_cmd_in_nxt[108]));
Q_MX02 U3696 ( .S(n90), .A0(kme_internal_out[9]), .A1(gcm_dak_cmd_in[108]), .Z(n1454));
Q_AN02 U3697 ( .A0(n35), .A1(n1455), .Z(gcm_dak_cmd_in_nxt[107]));
Q_MX02 U3698 ( .S(n90), .A0(kme_internal_out[8]), .A1(gcm_dak_cmd_in[107]), .Z(n1455));
Q_AN02 U3699 ( .A0(n35), .A1(n1456), .Z(gcm_dak_cmd_in_nxt[106]));
Q_MX02 U3700 ( .S(n90), .A0(kme_internal_out[7]), .A1(gcm_dak_cmd_in[106]), .Z(n1456));
Q_AN02 U3701 ( .A0(n35), .A1(n1457), .Z(gcm_dak_cmd_in_nxt[105]));
Q_MX02 U3702 ( .S(n90), .A0(kme_internal_out[6]), .A1(gcm_dak_cmd_in[105]), .Z(n1457));
Q_AN02 U3703 ( .A0(n35), .A1(n1458), .Z(gcm_dak_cmd_in_nxt[104]));
Q_MX02 U3704 ( .S(n90), .A0(kme_internal_out[5]), .A1(gcm_dak_cmd_in[104]), .Z(n1458));
Q_AN02 U3705 ( .A0(n35), .A1(n1459), .Z(gcm_dak_cmd_in_nxt[103]));
Q_MX02 U3706 ( .S(n90), .A0(kme_internal_out[4]), .A1(gcm_dak_cmd_in[103]), .Z(n1459));
Q_AN02 U3707 ( .A0(n35), .A1(n1460), .Z(gcm_dak_cmd_in_nxt[102]));
Q_MX02 U3708 ( .S(n90), .A0(kme_internal_out[3]), .A1(gcm_dak_cmd_in[102]), .Z(n1460));
Q_AN02 U3709 ( .A0(n35), .A1(n1461), .Z(gcm_dak_cmd_in_nxt[101]));
Q_MX02 U3710 ( .S(n90), .A0(kme_internal_out[2]), .A1(gcm_dak_cmd_in[101]), .Z(n1461));
Q_AN02 U3711 ( .A0(n35), .A1(n1462), .Z(gcm_dak_cmd_in_nxt[100]));
Q_MX02 U3712 ( .S(n90), .A0(kme_internal_out[1]), .A1(gcm_dak_cmd_in[100]), .Z(n1462));
Q_AN02 U3713 ( .A0(n35), .A1(n1463), .Z(gcm_dak_cmd_in_nxt[99]));
Q_MX02 U3714 ( .S(n90), .A0(kme_internal_out[0]), .A1(gcm_dak_cmd_in[99]), .Z(n1463));
Q_AN02 U3715 ( .A0(n35), .A1(n1464), .Z(gcm_dak_cmd_in_nxt[610]));
Q_MX02 U3716 ( .S(n90), .A0(gcm_dak_cmd_in[546]), .A1(gcm_dak_cmd_in[610]), .Z(n1464));
Q_AN02 U3717 ( .A0(n35), .A1(n1465), .Z(gcm_dak_cmd_in_nxt[609]));
Q_MX02 U3718 ( .S(n90), .A0(gcm_dak_cmd_in[545]), .A1(gcm_dak_cmd_in[609]), .Z(n1465));
Q_AN02 U3719 ( .A0(n35), .A1(n1466), .Z(gcm_dak_cmd_in_nxt[608]));
Q_MX02 U3720 ( .S(n90), .A0(gcm_dak_cmd_in[544]), .A1(gcm_dak_cmd_in[608]), .Z(n1466));
Q_AN02 U3721 ( .A0(n35), .A1(n1467), .Z(gcm_dak_cmd_in_nxt[607]));
Q_MX02 U3722 ( .S(n90), .A0(gcm_dak_cmd_in[543]), .A1(gcm_dak_cmd_in[607]), .Z(n1467));
Q_AN02 U3723 ( .A0(n35), .A1(n1468), .Z(gcm_dak_cmd_in_nxt[606]));
Q_MX02 U3724 ( .S(n90), .A0(gcm_dak_cmd_in[542]), .A1(gcm_dak_cmd_in[606]), .Z(n1468));
Q_AN02 U3725 ( .A0(n35), .A1(n1469), .Z(gcm_dak_cmd_in_nxt[605]));
Q_MX02 U3726 ( .S(n90), .A0(gcm_dak_cmd_in[541]), .A1(gcm_dak_cmd_in[605]), .Z(n1469));
Q_AN02 U3727 ( .A0(n35), .A1(n1470), .Z(gcm_dak_cmd_in_nxt[604]));
Q_MX02 U3728 ( .S(n90), .A0(gcm_dak_cmd_in[540]), .A1(gcm_dak_cmd_in[604]), .Z(n1470));
Q_AN02 U3729 ( .A0(n35), .A1(n1471), .Z(gcm_dak_cmd_in_nxt[603]));
Q_MX02 U3730 ( .S(n90), .A0(gcm_dak_cmd_in[539]), .A1(gcm_dak_cmd_in[603]), .Z(n1471));
Q_AN02 U3731 ( .A0(n35), .A1(n1472), .Z(gcm_dak_cmd_in_nxt[602]));
Q_MX02 U3732 ( .S(n90), .A0(gcm_dak_cmd_in[538]), .A1(gcm_dak_cmd_in[602]), .Z(n1472));
Q_AN02 U3733 ( .A0(n35), .A1(n1473), .Z(gcm_dak_cmd_in_nxt[601]));
Q_MX02 U3734 ( .S(n90), .A0(gcm_dak_cmd_in[537]), .A1(gcm_dak_cmd_in[601]), .Z(n1473));
Q_AN02 U3735 ( .A0(n35), .A1(n1474), .Z(gcm_dak_cmd_in_nxt[600]));
Q_MX02 U3736 ( .S(n90), .A0(gcm_dak_cmd_in[536]), .A1(gcm_dak_cmd_in[600]), .Z(n1474));
Q_AN02 U3737 ( .A0(n35), .A1(n1475), .Z(gcm_dak_cmd_in_nxt[599]));
Q_MX02 U3738 ( .S(n90), .A0(gcm_dak_cmd_in[535]), .A1(gcm_dak_cmd_in[599]), .Z(n1475));
Q_AN02 U3739 ( .A0(n35), .A1(n1476), .Z(gcm_dak_cmd_in_nxt[598]));
Q_MX02 U3740 ( .S(n90), .A0(gcm_dak_cmd_in[534]), .A1(gcm_dak_cmd_in[598]), .Z(n1476));
Q_AN02 U3741 ( .A0(n35), .A1(n1477), .Z(gcm_dak_cmd_in_nxt[597]));
Q_MX02 U3742 ( .S(n90), .A0(gcm_dak_cmd_in[533]), .A1(gcm_dak_cmd_in[597]), .Z(n1477));
Q_AN02 U3743 ( .A0(n35), .A1(n1478), .Z(gcm_dak_cmd_in_nxt[596]));
Q_MX02 U3744 ( .S(n90), .A0(gcm_dak_cmd_in[532]), .A1(gcm_dak_cmd_in[596]), .Z(n1478));
Q_AN02 U3745 ( .A0(n35), .A1(n1479), .Z(gcm_dak_cmd_in_nxt[595]));
Q_MX02 U3746 ( .S(n90), .A0(gcm_dak_cmd_in[531]), .A1(gcm_dak_cmd_in[595]), .Z(n1479));
Q_AN02 U3747 ( .A0(n35), .A1(n1480), .Z(gcm_dak_cmd_in_nxt[594]));
Q_MX02 U3748 ( .S(n90), .A0(gcm_dak_cmd_in[530]), .A1(gcm_dak_cmd_in[594]), .Z(n1480));
Q_AN02 U3749 ( .A0(n35), .A1(n1481), .Z(gcm_dak_cmd_in_nxt[593]));
Q_MX02 U3750 ( .S(n90), .A0(gcm_dak_cmd_in[529]), .A1(gcm_dak_cmd_in[593]), .Z(n1481));
Q_AN02 U3751 ( .A0(n35), .A1(n1482), .Z(gcm_dak_cmd_in_nxt[592]));
Q_MX02 U3752 ( .S(n90), .A0(gcm_dak_cmd_in[528]), .A1(gcm_dak_cmd_in[592]), .Z(n1482));
Q_AN02 U3753 ( .A0(n35), .A1(n1483), .Z(gcm_dak_cmd_in_nxt[591]));
Q_MX02 U3754 ( .S(n90), .A0(gcm_dak_cmd_in[527]), .A1(gcm_dak_cmd_in[591]), .Z(n1483));
Q_AN02 U3755 ( .A0(n35), .A1(n1484), .Z(gcm_dak_cmd_in_nxt[590]));
Q_MX02 U3756 ( .S(n90), .A0(gcm_dak_cmd_in[526]), .A1(gcm_dak_cmd_in[590]), .Z(n1484));
Q_AN02 U3757 ( .A0(n35), .A1(n1485), .Z(gcm_dak_cmd_in_nxt[589]));
Q_MX02 U3758 ( .S(n90), .A0(gcm_dak_cmd_in[525]), .A1(gcm_dak_cmd_in[589]), .Z(n1485));
Q_AN02 U3759 ( .A0(n35), .A1(n1486), .Z(gcm_dak_cmd_in_nxt[588]));
Q_MX02 U3760 ( .S(n90), .A0(gcm_dak_cmd_in[524]), .A1(gcm_dak_cmd_in[588]), .Z(n1486));
Q_AN02 U3761 ( .A0(n35), .A1(n1487), .Z(gcm_dak_cmd_in_nxt[587]));
Q_MX02 U3762 ( .S(n90), .A0(gcm_dak_cmd_in[523]), .A1(gcm_dak_cmd_in[587]), .Z(n1487));
Q_AN02 U3763 ( .A0(n35), .A1(n1488), .Z(gcm_dak_cmd_in_nxt[586]));
Q_MX02 U3764 ( .S(n90), .A0(gcm_dak_cmd_in[522]), .A1(gcm_dak_cmd_in[586]), .Z(n1488));
Q_AN02 U3765 ( .A0(n35), .A1(n1489), .Z(gcm_dak_cmd_in_nxt[585]));
Q_MX02 U3766 ( .S(n90), .A0(gcm_dak_cmd_in[521]), .A1(gcm_dak_cmd_in[585]), .Z(n1489));
Q_AN02 U3767 ( .A0(n35), .A1(n1490), .Z(gcm_dak_cmd_in_nxt[584]));
Q_MX02 U3768 ( .S(n90), .A0(gcm_dak_cmd_in[520]), .A1(gcm_dak_cmd_in[584]), .Z(n1490));
Q_AN02 U3769 ( .A0(n35), .A1(n1491), .Z(gcm_dak_cmd_in_nxt[583]));
Q_MX02 U3770 ( .S(n90), .A0(gcm_dak_cmd_in[519]), .A1(gcm_dak_cmd_in[583]), .Z(n1491));
Q_AN02 U3771 ( .A0(n35), .A1(n1492), .Z(gcm_dak_cmd_in_nxt[582]));
Q_MX02 U3772 ( .S(n90), .A0(gcm_dak_cmd_in[518]), .A1(gcm_dak_cmd_in[582]), .Z(n1492));
Q_AN02 U3773 ( .A0(n35), .A1(n1493), .Z(gcm_dak_cmd_in_nxt[581]));
Q_MX02 U3774 ( .S(n90), .A0(gcm_dak_cmd_in[517]), .A1(gcm_dak_cmd_in[581]), .Z(n1493));
Q_AN02 U3775 ( .A0(n35), .A1(n1494), .Z(gcm_dak_cmd_in_nxt[580]));
Q_MX02 U3776 ( .S(n90), .A0(gcm_dak_cmd_in[516]), .A1(gcm_dak_cmd_in[580]), .Z(n1494));
Q_AN02 U3777 ( .A0(n35), .A1(n1495), .Z(gcm_dak_cmd_in_nxt[579]));
Q_MX02 U3778 ( .S(n90), .A0(gcm_dak_cmd_in[515]), .A1(gcm_dak_cmd_in[579]), .Z(n1495));
Q_AN02 U3779 ( .A0(n35), .A1(n1496), .Z(gcm_dak_cmd_in_nxt[578]));
Q_MX02 U3780 ( .S(n90), .A0(gcm_dak_cmd_in[514]), .A1(gcm_dak_cmd_in[578]), .Z(n1496));
Q_AN02 U3781 ( .A0(n35), .A1(n1497), .Z(gcm_dak_cmd_in_nxt[577]));
Q_MX02 U3782 ( .S(n90), .A0(gcm_dak_cmd_in[513]), .A1(gcm_dak_cmd_in[577]), .Z(n1497));
Q_AN02 U3783 ( .A0(n35), .A1(n1498), .Z(gcm_dak_cmd_in_nxt[576]));
Q_MX02 U3784 ( .S(n90), .A0(gcm_dak_cmd_in[512]), .A1(gcm_dak_cmd_in[576]), .Z(n1498));
Q_AN02 U3785 ( .A0(n35), .A1(n1499), .Z(gcm_dak_cmd_in_nxt[575]));
Q_MX02 U3786 ( .S(n90), .A0(gcm_dak_cmd_in[511]), .A1(gcm_dak_cmd_in[575]), .Z(n1499));
Q_AN02 U3787 ( .A0(n35), .A1(n1500), .Z(gcm_dak_cmd_in_nxt[574]));
Q_MX02 U3788 ( .S(n90), .A0(gcm_dak_cmd_in[510]), .A1(gcm_dak_cmd_in[574]), .Z(n1500));
Q_AN02 U3789 ( .A0(n35), .A1(n1501), .Z(gcm_dak_cmd_in_nxt[573]));
Q_MX02 U3790 ( .S(n90), .A0(gcm_dak_cmd_in[509]), .A1(gcm_dak_cmd_in[573]), .Z(n1501));
Q_AN02 U3791 ( .A0(n35), .A1(n1502), .Z(gcm_dak_cmd_in_nxt[572]));
Q_MX02 U3792 ( .S(n90), .A0(gcm_dak_cmd_in[508]), .A1(gcm_dak_cmd_in[572]), .Z(n1502));
Q_AN02 U3793 ( .A0(n35), .A1(n1503), .Z(gcm_dak_cmd_in_nxt[571]));
Q_MX02 U3794 ( .S(n90), .A0(gcm_dak_cmd_in[507]), .A1(gcm_dak_cmd_in[571]), .Z(n1503));
Q_AN02 U3795 ( .A0(n35), .A1(n1504), .Z(gcm_dak_cmd_in_nxt[570]));
Q_MX02 U3796 ( .S(n90), .A0(gcm_dak_cmd_in[506]), .A1(gcm_dak_cmd_in[570]), .Z(n1504));
Q_AN02 U3797 ( .A0(n35), .A1(n1505), .Z(gcm_dak_cmd_in_nxt[569]));
Q_MX02 U3798 ( .S(n90), .A0(gcm_dak_cmd_in[505]), .A1(gcm_dak_cmd_in[569]), .Z(n1505));
Q_AN02 U3799 ( .A0(n35), .A1(n1506), .Z(gcm_dak_cmd_in_nxt[568]));
Q_MX02 U3800 ( .S(n90), .A0(gcm_dak_cmd_in[504]), .A1(gcm_dak_cmd_in[568]), .Z(n1506));
Q_AN02 U3801 ( .A0(n35), .A1(n1507), .Z(gcm_dak_cmd_in_nxt[567]));
Q_MX02 U3802 ( .S(n90), .A0(gcm_dak_cmd_in[503]), .A1(gcm_dak_cmd_in[567]), .Z(n1507));
Q_AN02 U3803 ( .A0(n35), .A1(n1508), .Z(gcm_dak_cmd_in_nxt[566]));
Q_MX02 U3804 ( .S(n90), .A0(gcm_dak_cmd_in[502]), .A1(gcm_dak_cmd_in[566]), .Z(n1508));
Q_AN02 U3805 ( .A0(n35), .A1(n1509), .Z(gcm_dak_cmd_in_nxt[565]));
Q_MX02 U3806 ( .S(n90), .A0(gcm_dak_cmd_in[501]), .A1(gcm_dak_cmd_in[565]), .Z(n1509));
Q_AN02 U3807 ( .A0(n35), .A1(n1510), .Z(gcm_dak_cmd_in_nxt[564]));
Q_MX02 U3808 ( .S(n90), .A0(gcm_dak_cmd_in[500]), .A1(gcm_dak_cmd_in[564]), .Z(n1510));
Q_AN02 U3809 ( .A0(n35), .A1(n1511), .Z(gcm_dak_cmd_in_nxt[563]));
Q_MX02 U3810 ( .S(n90), .A0(gcm_dak_cmd_in[499]), .A1(gcm_dak_cmd_in[563]), .Z(n1511));
Q_AN02 U3811 ( .A0(n35), .A1(n1512), .Z(gcm_dak_cmd_in_nxt[562]));
Q_MX02 U3812 ( .S(n90), .A0(gcm_dak_cmd_in[498]), .A1(gcm_dak_cmd_in[562]), .Z(n1512));
Q_AN02 U3813 ( .A0(n35), .A1(n1513), .Z(gcm_dak_cmd_in_nxt[561]));
Q_MX02 U3814 ( .S(n90), .A0(gcm_dak_cmd_in[497]), .A1(gcm_dak_cmd_in[561]), .Z(n1513));
Q_AN02 U3815 ( .A0(n35), .A1(n1514), .Z(gcm_dak_cmd_in_nxt[560]));
Q_MX02 U3816 ( .S(n90), .A0(gcm_dak_cmd_in[496]), .A1(gcm_dak_cmd_in[560]), .Z(n1514));
Q_AN02 U3817 ( .A0(n35), .A1(n1515), .Z(gcm_dak_cmd_in_nxt[559]));
Q_MX02 U3818 ( .S(n90), .A0(gcm_dak_cmd_in[495]), .A1(gcm_dak_cmd_in[559]), .Z(n1515));
Q_AN02 U3819 ( .A0(n35), .A1(n1516), .Z(gcm_dak_cmd_in_nxt[558]));
Q_MX02 U3820 ( .S(n90), .A0(gcm_dak_cmd_in[494]), .A1(gcm_dak_cmd_in[558]), .Z(n1516));
Q_AN02 U3821 ( .A0(n35), .A1(n1517), .Z(gcm_dak_cmd_in_nxt[557]));
Q_MX02 U3822 ( .S(n90), .A0(gcm_dak_cmd_in[493]), .A1(gcm_dak_cmd_in[557]), .Z(n1517));
Q_AN02 U3823 ( .A0(n35), .A1(n1518), .Z(gcm_dak_cmd_in_nxt[556]));
Q_MX02 U3824 ( .S(n90), .A0(gcm_dak_cmd_in[492]), .A1(gcm_dak_cmd_in[556]), .Z(n1518));
Q_AN02 U3825 ( .A0(n35), .A1(n1519), .Z(gcm_dak_cmd_in_nxt[555]));
Q_MX02 U3826 ( .S(n90), .A0(gcm_dak_cmd_in[491]), .A1(gcm_dak_cmd_in[555]), .Z(n1519));
Q_AN02 U3827 ( .A0(n35), .A1(n1520), .Z(gcm_dak_cmd_in_nxt[554]));
Q_MX02 U3828 ( .S(n90), .A0(gcm_dak_cmd_in[490]), .A1(gcm_dak_cmd_in[554]), .Z(n1520));
Q_AN02 U3829 ( .A0(n35), .A1(n1521), .Z(gcm_dak_cmd_in_nxt[553]));
Q_MX02 U3830 ( .S(n90), .A0(gcm_dak_cmd_in[489]), .A1(gcm_dak_cmd_in[553]), .Z(n1521));
Q_AN02 U3831 ( .A0(n35), .A1(n1522), .Z(gcm_dak_cmd_in_nxt[552]));
Q_MX02 U3832 ( .S(n90), .A0(gcm_dak_cmd_in[488]), .A1(gcm_dak_cmd_in[552]), .Z(n1522));
Q_AN02 U3833 ( .A0(n35), .A1(n1523), .Z(gcm_dak_cmd_in_nxt[551]));
Q_MX02 U3834 ( .S(n90), .A0(gcm_dak_cmd_in[487]), .A1(gcm_dak_cmd_in[551]), .Z(n1523));
Q_AN02 U3835 ( .A0(n35), .A1(n1524), .Z(gcm_dak_cmd_in_nxt[550]));
Q_MX02 U3836 ( .S(n90), .A0(gcm_dak_cmd_in[486]), .A1(gcm_dak_cmd_in[550]), .Z(n1524));
Q_AN02 U3837 ( .A0(n35), .A1(n1525), .Z(gcm_dak_cmd_in_nxt[549]));
Q_MX02 U3838 ( .S(n90), .A0(gcm_dak_cmd_in[485]), .A1(gcm_dak_cmd_in[549]), .Z(n1525));
Q_AN02 U3839 ( .A0(n35), .A1(n1526), .Z(gcm_dak_cmd_in_nxt[548]));
Q_MX02 U3840 ( .S(n90), .A0(gcm_dak_cmd_in[484]), .A1(gcm_dak_cmd_in[548]), .Z(n1526));
Q_AN02 U3841 ( .A0(n35), .A1(n1527), .Z(gcm_dak_cmd_in_nxt[547]));
Q_MX02 U3842 ( .S(n90), .A0(gcm_dak_cmd_in[483]), .A1(gcm_dak_cmd_in[547]), .Z(n1527));
Q_AN02 U3843 ( .A0(n35), .A1(n1528), .Z(gcm_dak_cmd_in_nxt[546]));
Q_MX02 U3844 ( .S(n90), .A0(gcm_dak_cmd_in[482]), .A1(gcm_dak_cmd_in[546]), .Z(n1528));
Q_AN02 U3845 ( .A0(n35), .A1(n1529), .Z(gcm_dak_cmd_in_nxt[545]));
Q_MX02 U3846 ( .S(n90), .A0(gcm_dak_cmd_in[481]), .A1(gcm_dak_cmd_in[545]), .Z(n1529));
Q_AN02 U3847 ( .A0(n35), .A1(n1530), .Z(gcm_dak_cmd_in_nxt[544]));
Q_MX02 U3848 ( .S(n90), .A0(gcm_dak_cmd_in[480]), .A1(gcm_dak_cmd_in[544]), .Z(n1530));
Q_AN02 U3849 ( .A0(n35), .A1(n1531), .Z(gcm_dak_cmd_in_nxt[543]));
Q_MX02 U3850 ( .S(n90), .A0(gcm_dak_cmd_in[479]), .A1(gcm_dak_cmd_in[543]), .Z(n1531));
Q_AN02 U3851 ( .A0(n35), .A1(n1532), .Z(gcm_dak_cmd_in_nxt[542]));
Q_MX02 U3852 ( .S(n90), .A0(gcm_dak_cmd_in[478]), .A1(gcm_dak_cmd_in[542]), .Z(n1532));
Q_AN02 U3853 ( .A0(n35), .A1(n1533), .Z(gcm_dak_cmd_in_nxt[541]));
Q_MX02 U3854 ( .S(n90), .A0(gcm_dak_cmd_in[477]), .A1(gcm_dak_cmd_in[541]), .Z(n1533));
Q_AN02 U3855 ( .A0(n35), .A1(n1534), .Z(gcm_dak_cmd_in_nxt[540]));
Q_MX02 U3856 ( .S(n90), .A0(gcm_dak_cmd_in[476]), .A1(gcm_dak_cmd_in[540]), .Z(n1534));
Q_AN02 U3857 ( .A0(n35), .A1(n1535), .Z(gcm_dak_cmd_in_nxt[539]));
Q_MX02 U3858 ( .S(n90), .A0(gcm_dak_cmd_in[475]), .A1(gcm_dak_cmd_in[539]), .Z(n1535));
Q_AN02 U3859 ( .A0(n35), .A1(n1536), .Z(gcm_dak_cmd_in_nxt[538]));
Q_MX02 U3860 ( .S(n90), .A0(gcm_dak_cmd_in[474]), .A1(gcm_dak_cmd_in[538]), .Z(n1536));
Q_AN02 U3861 ( .A0(n35), .A1(n1537), .Z(gcm_dak_cmd_in_nxt[537]));
Q_MX02 U3862 ( .S(n90), .A0(gcm_dak_cmd_in[473]), .A1(gcm_dak_cmd_in[537]), .Z(n1537));
Q_AN02 U3863 ( .A0(n35), .A1(n1538), .Z(gcm_dak_cmd_in_nxt[536]));
Q_MX02 U3864 ( .S(n90), .A0(gcm_dak_cmd_in[472]), .A1(gcm_dak_cmd_in[536]), .Z(n1538));
Q_AN02 U3865 ( .A0(n35), .A1(n1539), .Z(gcm_dak_cmd_in_nxt[535]));
Q_MX02 U3866 ( .S(n90), .A0(gcm_dak_cmd_in[471]), .A1(gcm_dak_cmd_in[535]), .Z(n1539));
Q_AN02 U3867 ( .A0(n35), .A1(n1540), .Z(gcm_dak_cmd_in_nxt[534]));
Q_MX02 U3868 ( .S(n90), .A0(gcm_dak_cmd_in[470]), .A1(gcm_dak_cmd_in[534]), .Z(n1540));
Q_AN02 U3869 ( .A0(n35), .A1(n1541), .Z(gcm_dak_cmd_in_nxt[533]));
Q_MX02 U3870 ( .S(n90), .A0(gcm_dak_cmd_in[469]), .A1(gcm_dak_cmd_in[533]), .Z(n1541));
Q_AN02 U3871 ( .A0(n35), .A1(n1542), .Z(gcm_dak_cmd_in_nxt[532]));
Q_MX02 U3872 ( .S(n90), .A0(gcm_dak_cmd_in[468]), .A1(gcm_dak_cmd_in[532]), .Z(n1542));
Q_AN02 U3873 ( .A0(n35), .A1(n1543), .Z(gcm_dak_cmd_in_nxt[531]));
Q_MX02 U3874 ( .S(n90), .A0(gcm_dak_cmd_in[467]), .A1(gcm_dak_cmd_in[531]), .Z(n1543));
Q_AN02 U3875 ( .A0(n35), .A1(n1544), .Z(gcm_dak_cmd_in_nxt[530]));
Q_MX02 U3876 ( .S(n90), .A0(gcm_dak_cmd_in[466]), .A1(gcm_dak_cmd_in[530]), .Z(n1544));
Q_AN02 U3877 ( .A0(n35), .A1(n1545), .Z(gcm_dak_cmd_in_nxt[529]));
Q_MX02 U3878 ( .S(n90), .A0(gcm_dak_cmd_in[465]), .A1(gcm_dak_cmd_in[529]), .Z(n1545));
Q_AN02 U3879 ( .A0(n35), .A1(n1546), .Z(gcm_dak_cmd_in_nxt[528]));
Q_MX02 U3880 ( .S(n90), .A0(gcm_dak_cmd_in[464]), .A1(gcm_dak_cmd_in[528]), .Z(n1546));
Q_AN02 U3881 ( .A0(n35), .A1(n1547), .Z(gcm_dak_cmd_in_nxt[527]));
Q_MX02 U3882 ( .S(n90), .A0(gcm_dak_cmd_in[463]), .A1(gcm_dak_cmd_in[527]), .Z(n1547));
Q_AN02 U3883 ( .A0(n35), .A1(n1548), .Z(gcm_dak_cmd_in_nxt[526]));
Q_MX02 U3884 ( .S(n90), .A0(gcm_dak_cmd_in[462]), .A1(gcm_dak_cmd_in[526]), .Z(n1548));
Q_AN02 U3885 ( .A0(n35), .A1(n1549), .Z(gcm_dak_cmd_in_nxt[525]));
Q_MX02 U3886 ( .S(n90), .A0(gcm_dak_cmd_in[461]), .A1(gcm_dak_cmd_in[525]), .Z(n1549));
Q_AN02 U3887 ( .A0(n35), .A1(n1550), .Z(gcm_dak_cmd_in_nxt[524]));
Q_MX02 U3888 ( .S(n90), .A0(gcm_dak_cmd_in[460]), .A1(gcm_dak_cmd_in[524]), .Z(n1550));
Q_AN02 U3889 ( .A0(n35), .A1(n1551), .Z(gcm_dak_cmd_in_nxt[523]));
Q_MX02 U3890 ( .S(n90), .A0(gcm_dak_cmd_in[459]), .A1(gcm_dak_cmd_in[523]), .Z(n1551));
Q_AN02 U3891 ( .A0(n35), .A1(n1552), .Z(gcm_dak_cmd_in_nxt[522]));
Q_MX02 U3892 ( .S(n90), .A0(gcm_dak_cmd_in[458]), .A1(gcm_dak_cmd_in[522]), .Z(n1552));
Q_AN02 U3893 ( .A0(n35), .A1(n1553), .Z(gcm_dak_cmd_in_nxt[521]));
Q_MX02 U3894 ( .S(n90), .A0(gcm_dak_cmd_in[457]), .A1(gcm_dak_cmd_in[521]), .Z(n1553));
Q_AN02 U3895 ( .A0(n35), .A1(n1554), .Z(gcm_dak_cmd_in_nxt[520]));
Q_MX02 U3896 ( .S(n90), .A0(gcm_dak_cmd_in[456]), .A1(gcm_dak_cmd_in[520]), .Z(n1554));
Q_AN02 U3897 ( .A0(n35), .A1(n1555), .Z(gcm_dak_cmd_in_nxt[519]));
Q_MX02 U3898 ( .S(n90), .A0(gcm_dak_cmd_in[455]), .A1(gcm_dak_cmd_in[519]), .Z(n1555));
Q_AN02 U3899 ( .A0(n35), .A1(n1556), .Z(gcm_dak_cmd_in_nxt[518]));
Q_MX02 U3900 ( .S(n90), .A0(gcm_dak_cmd_in[454]), .A1(gcm_dak_cmd_in[518]), .Z(n1556));
Q_AN02 U3901 ( .A0(n35), .A1(n1557), .Z(gcm_dak_cmd_in_nxt[517]));
Q_MX02 U3902 ( .S(n90), .A0(gcm_dak_cmd_in[453]), .A1(gcm_dak_cmd_in[517]), .Z(n1557));
Q_AN02 U3903 ( .A0(n35), .A1(n1558), .Z(gcm_dak_cmd_in_nxt[516]));
Q_MX02 U3904 ( .S(n90), .A0(gcm_dak_cmd_in[452]), .A1(gcm_dak_cmd_in[516]), .Z(n1558));
Q_AN02 U3905 ( .A0(n35), .A1(n1559), .Z(gcm_dak_cmd_in_nxt[515]));
Q_MX02 U3906 ( .S(n90), .A0(gcm_dak_cmd_in[451]), .A1(gcm_dak_cmd_in[515]), .Z(n1559));
Q_AN02 U3907 ( .A0(n35), .A1(n1560), .Z(gcm_dak_cmd_in_nxt[514]));
Q_MX02 U3908 ( .S(n90), .A0(gcm_dak_cmd_in[450]), .A1(gcm_dak_cmd_in[514]), .Z(n1560));
Q_AN02 U3909 ( .A0(n35), .A1(n1561), .Z(gcm_dak_cmd_in_nxt[513]));
Q_MX02 U3910 ( .S(n90), .A0(gcm_dak_cmd_in[449]), .A1(gcm_dak_cmd_in[513]), .Z(n1561));
Q_AN02 U3911 ( .A0(n35), .A1(n1562), .Z(gcm_dak_cmd_in_nxt[512]));
Q_MX02 U3912 ( .S(n90), .A0(gcm_dak_cmd_in[448]), .A1(gcm_dak_cmd_in[512]), .Z(n1562));
Q_AN02 U3913 ( .A0(n35), .A1(n1563), .Z(gcm_dak_cmd_in_nxt[511]));
Q_MX02 U3914 ( .S(n90), .A0(gcm_dak_cmd_in[447]), .A1(gcm_dak_cmd_in[511]), .Z(n1563));
Q_AN02 U3915 ( .A0(n35), .A1(n1564), .Z(gcm_dak_cmd_in_nxt[510]));
Q_MX02 U3916 ( .S(n90), .A0(gcm_dak_cmd_in[446]), .A1(gcm_dak_cmd_in[510]), .Z(n1564));
Q_AN02 U3917 ( .A0(n35), .A1(n1565), .Z(gcm_dak_cmd_in_nxt[509]));
Q_MX02 U3918 ( .S(n90), .A0(gcm_dak_cmd_in[445]), .A1(gcm_dak_cmd_in[509]), .Z(n1565));
Q_AN02 U3919 ( .A0(n35), .A1(n1566), .Z(gcm_dak_cmd_in_nxt[508]));
Q_MX02 U3920 ( .S(n90), .A0(gcm_dak_cmd_in[444]), .A1(gcm_dak_cmd_in[508]), .Z(n1566));
Q_AN02 U3921 ( .A0(n35), .A1(n1567), .Z(gcm_dak_cmd_in_nxt[507]));
Q_MX02 U3922 ( .S(n90), .A0(gcm_dak_cmd_in[443]), .A1(gcm_dak_cmd_in[507]), .Z(n1567));
Q_AN02 U3923 ( .A0(n35), .A1(n1568), .Z(gcm_dak_cmd_in_nxt[506]));
Q_MX02 U3924 ( .S(n90), .A0(gcm_dak_cmd_in[442]), .A1(gcm_dak_cmd_in[506]), .Z(n1568));
Q_AN02 U3925 ( .A0(n35), .A1(n1569), .Z(gcm_dak_cmd_in_nxt[505]));
Q_MX02 U3926 ( .S(n90), .A0(gcm_dak_cmd_in[441]), .A1(gcm_dak_cmd_in[505]), .Z(n1569));
Q_AN02 U3927 ( .A0(n35), .A1(n1570), .Z(gcm_dak_cmd_in_nxt[504]));
Q_MX02 U3928 ( .S(n90), .A0(gcm_dak_cmd_in[440]), .A1(gcm_dak_cmd_in[504]), .Z(n1570));
Q_AN02 U3929 ( .A0(n35), .A1(n1571), .Z(gcm_dak_cmd_in_nxt[503]));
Q_MX02 U3930 ( .S(n90), .A0(gcm_dak_cmd_in[439]), .A1(gcm_dak_cmd_in[503]), .Z(n1571));
Q_AN02 U3931 ( .A0(n35), .A1(n1572), .Z(gcm_dak_cmd_in_nxt[502]));
Q_MX02 U3932 ( .S(n90), .A0(gcm_dak_cmd_in[438]), .A1(gcm_dak_cmd_in[502]), .Z(n1572));
Q_AN02 U3933 ( .A0(n35), .A1(n1573), .Z(gcm_dak_cmd_in_nxt[501]));
Q_MX02 U3934 ( .S(n90), .A0(gcm_dak_cmd_in[437]), .A1(gcm_dak_cmd_in[501]), .Z(n1573));
Q_AN02 U3935 ( .A0(n35), .A1(n1574), .Z(gcm_dak_cmd_in_nxt[500]));
Q_MX02 U3936 ( .S(n90), .A0(gcm_dak_cmd_in[436]), .A1(gcm_dak_cmd_in[500]), .Z(n1574));
Q_AN02 U3937 ( .A0(n35), .A1(n1575), .Z(gcm_dak_cmd_in_nxt[499]));
Q_MX02 U3938 ( .S(n90), .A0(gcm_dak_cmd_in[435]), .A1(gcm_dak_cmd_in[499]), .Z(n1575));
Q_AN02 U3939 ( .A0(n35), .A1(n1576), .Z(gcm_dak_cmd_in_nxt[498]));
Q_MX02 U3940 ( .S(n90), .A0(gcm_dak_cmd_in[434]), .A1(gcm_dak_cmd_in[498]), .Z(n1576));
Q_AN02 U3941 ( .A0(n35), .A1(n1577), .Z(gcm_dak_cmd_in_nxt[497]));
Q_MX02 U3942 ( .S(n90), .A0(gcm_dak_cmd_in[433]), .A1(gcm_dak_cmd_in[497]), .Z(n1577));
Q_AN02 U3943 ( .A0(n35), .A1(n1578), .Z(gcm_dak_cmd_in_nxt[496]));
Q_MX02 U3944 ( .S(n90), .A0(gcm_dak_cmd_in[432]), .A1(gcm_dak_cmd_in[496]), .Z(n1578));
Q_AN02 U3945 ( .A0(n35), .A1(n1579), .Z(gcm_dak_cmd_in_nxt[495]));
Q_MX02 U3946 ( .S(n90), .A0(gcm_dak_cmd_in[431]), .A1(gcm_dak_cmd_in[495]), .Z(n1579));
Q_AN02 U3947 ( .A0(n35), .A1(n1580), .Z(gcm_dak_cmd_in_nxt[494]));
Q_MX02 U3948 ( .S(n90), .A0(gcm_dak_cmd_in[430]), .A1(gcm_dak_cmd_in[494]), .Z(n1580));
Q_AN02 U3949 ( .A0(n35), .A1(n1581), .Z(gcm_dak_cmd_in_nxt[493]));
Q_MX02 U3950 ( .S(n90), .A0(gcm_dak_cmd_in[429]), .A1(gcm_dak_cmd_in[493]), .Z(n1581));
Q_AN02 U3951 ( .A0(n35), .A1(n1582), .Z(gcm_dak_cmd_in_nxt[492]));
Q_MX02 U3952 ( .S(n90), .A0(gcm_dak_cmd_in[428]), .A1(gcm_dak_cmd_in[492]), .Z(n1582));
Q_AN02 U3953 ( .A0(n35), .A1(n1583), .Z(gcm_dak_cmd_in_nxt[491]));
Q_MX02 U3954 ( .S(n90), .A0(gcm_dak_cmd_in[427]), .A1(gcm_dak_cmd_in[491]), .Z(n1583));
Q_AN02 U3955 ( .A0(n35), .A1(n1584), .Z(gcm_dak_cmd_in_nxt[490]));
Q_MX02 U3956 ( .S(n90), .A0(gcm_dak_cmd_in[426]), .A1(gcm_dak_cmd_in[490]), .Z(n1584));
Q_AN02 U3957 ( .A0(n35), .A1(n1585), .Z(gcm_dak_cmd_in_nxt[489]));
Q_MX02 U3958 ( .S(n90), .A0(gcm_dak_cmd_in[425]), .A1(gcm_dak_cmd_in[489]), .Z(n1585));
Q_AN02 U3959 ( .A0(n35), .A1(n1586), .Z(gcm_dak_cmd_in_nxt[488]));
Q_MX02 U3960 ( .S(n90), .A0(gcm_dak_cmd_in[424]), .A1(gcm_dak_cmd_in[488]), .Z(n1586));
Q_AN02 U3961 ( .A0(n35), .A1(n1587), .Z(gcm_dak_cmd_in_nxt[487]));
Q_MX02 U3962 ( .S(n90), .A0(gcm_dak_cmd_in[423]), .A1(gcm_dak_cmd_in[487]), .Z(n1587));
Q_AN02 U3963 ( .A0(n35), .A1(n1588), .Z(gcm_dak_cmd_in_nxt[486]));
Q_MX02 U3964 ( .S(n90), .A0(gcm_dak_cmd_in[422]), .A1(gcm_dak_cmd_in[486]), .Z(n1588));
Q_AN02 U3965 ( .A0(n35), .A1(n1589), .Z(gcm_dak_cmd_in_nxt[485]));
Q_MX02 U3966 ( .S(n90), .A0(gcm_dak_cmd_in[421]), .A1(gcm_dak_cmd_in[485]), .Z(n1589));
Q_AN02 U3967 ( .A0(n35), .A1(n1590), .Z(gcm_dak_cmd_in_nxt[484]));
Q_MX02 U3968 ( .S(n90), .A0(gcm_dak_cmd_in[420]), .A1(gcm_dak_cmd_in[484]), .Z(n1590));
Q_AN02 U3969 ( .A0(n35), .A1(n1591), .Z(gcm_dak_cmd_in_nxt[483]));
Q_MX02 U3970 ( .S(n90), .A0(gcm_dak_cmd_in[419]), .A1(gcm_dak_cmd_in[483]), .Z(n1591));
Q_AN02 U3971 ( .A0(n35), .A1(n1592), .Z(gcm_dak_cmd_in_nxt[482]));
Q_MX02 U3972 ( .S(n90), .A0(gcm_dak_cmd_in[418]), .A1(gcm_dak_cmd_in[482]), .Z(n1592));
Q_AN02 U3973 ( .A0(n35), .A1(n1593), .Z(gcm_dak_cmd_in_nxt[481]));
Q_MX02 U3974 ( .S(n90), .A0(gcm_dak_cmd_in[417]), .A1(gcm_dak_cmd_in[481]), .Z(n1593));
Q_AN02 U3975 ( .A0(n35), .A1(n1594), .Z(gcm_dak_cmd_in_nxt[480]));
Q_MX02 U3976 ( .S(n90), .A0(gcm_dak_cmd_in[416]), .A1(gcm_dak_cmd_in[480]), .Z(n1594));
Q_AN02 U3977 ( .A0(n35), .A1(n1595), .Z(gcm_dak_cmd_in_nxt[479]));
Q_MX02 U3978 ( .S(n90), .A0(gcm_dak_cmd_in[415]), .A1(gcm_dak_cmd_in[479]), .Z(n1595));
Q_AN02 U3979 ( .A0(n35), .A1(n1596), .Z(gcm_dak_cmd_in_nxt[478]));
Q_MX02 U3980 ( .S(n90), .A0(gcm_dak_cmd_in[414]), .A1(gcm_dak_cmd_in[478]), .Z(n1596));
Q_AN02 U3981 ( .A0(n35), .A1(n1597), .Z(gcm_dak_cmd_in_nxt[477]));
Q_MX02 U3982 ( .S(n90), .A0(gcm_dak_cmd_in[413]), .A1(gcm_dak_cmd_in[477]), .Z(n1597));
Q_AN02 U3983 ( .A0(n35), .A1(n1598), .Z(gcm_dak_cmd_in_nxt[476]));
Q_MX02 U3984 ( .S(n90), .A0(gcm_dak_cmd_in[412]), .A1(gcm_dak_cmd_in[476]), .Z(n1598));
Q_AN02 U3985 ( .A0(n35), .A1(n1599), .Z(gcm_dak_cmd_in_nxt[475]));
Q_MX02 U3986 ( .S(n90), .A0(gcm_dak_cmd_in[411]), .A1(gcm_dak_cmd_in[475]), .Z(n1599));
Q_AN02 U3987 ( .A0(n35), .A1(n1600), .Z(gcm_dak_cmd_in_nxt[474]));
Q_MX02 U3988 ( .S(n90), .A0(gcm_dak_cmd_in[410]), .A1(gcm_dak_cmd_in[474]), .Z(n1600));
Q_AN02 U3989 ( .A0(n35), .A1(n1601), .Z(gcm_dak_cmd_in_nxt[473]));
Q_MX02 U3990 ( .S(n90), .A0(gcm_dak_cmd_in[409]), .A1(gcm_dak_cmd_in[473]), .Z(n1601));
Q_AN02 U3991 ( .A0(n35), .A1(n1602), .Z(gcm_dak_cmd_in_nxt[472]));
Q_MX02 U3992 ( .S(n90), .A0(gcm_dak_cmd_in[408]), .A1(gcm_dak_cmd_in[472]), .Z(n1602));
Q_AN02 U3993 ( .A0(n35), .A1(n1603), .Z(gcm_dak_cmd_in_nxt[471]));
Q_MX02 U3994 ( .S(n90), .A0(gcm_dak_cmd_in[407]), .A1(gcm_dak_cmd_in[471]), .Z(n1603));
Q_AN02 U3995 ( .A0(n35), .A1(n1604), .Z(gcm_dak_cmd_in_nxt[470]));
Q_MX02 U3996 ( .S(n90), .A0(gcm_dak_cmd_in[406]), .A1(gcm_dak_cmd_in[470]), .Z(n1604));
Q_AN02 U3997 ( .A0(n35), .A1(n1605), .Z(gcm_dak_cmd_in_nxt[469]));
Q_MX02 U3998 ( .S(n90), .A0(gcm_dak_cmd_in[405]), .A1(gcm_dak_cmd_in[469]), .Z(n1605));
Q_AN02 U3999 ( .A0(n35), .A1(n1606), .Z(gcm_dak_cmd_in_nxt[468]));
Q_MX02 U4000 ( .S(n90), .A0(gcm_dak_cmd_in[404]), .A1(gcm_dak_cmd_in[468]), .Z(n1606));
Q_AN02 U4001 ( .A0(n35), .A1(n1607), .Z(gcm_dak_cmd_in_nxt[467]));
Q_MX02 U4002 ( .S(n90), .A0(gcm_dak_cmd_in[403]), .A1(gcm_dak_cmd_in[467]), .Z(n1607));
Q_AN02 U4003 ( .A0(n35), .A1(n1608), .Z(gcm_dak_cmd_in_nxt[466]));
Q_MX02 U4004 ( .S(n90), .A0(gcm_dak_cmd_in[402]), .A1(gcm_dak_cmd_in[466]), .Z(n1608));
Q_AN02 U4005 ( .A0(n35), .A1(n1609), .Z(gcm_dak_cmd_in_nxt[465]));
Q_MX02 U4006 ( .S(n90), .A0(gcm_dak_cmd_in[401]), .A1(gcm_dak_cmd_in[465]), .Z(n1609));
Q_AN02 U4007 ( .A0(n35), .A1(n1610), .Z(gcm_dak_cmd_in_nxt[464]));
Q_MX02 U4008 ( .S(n90), .A0(gcm_dak_cmd_in[400]), .A1(gcm_dak_cmd_in[464]), .Z(n1610));
Q_AN02 U4009 ( .A0(n35), .A1(n1611), .Z(gcm_dak_cmd_in_nxt[463]));
Q_MX02 U4010 ( .S(n90), .A0(gcm_dak_cmd_in[399]), .A1(gcm_dak_cmd_in[463]), .Z(n1611));
Q_AN02 U4011 ( .A0(n35), .A1(n1612), .Z(gcm_dak_cmd_in_nxt[462]));
Q_MX02 U4012 ( .S(n90), .A0(gcm_dak_cmd_in[398]), .A1(gcm_dak_cmd_in[462]), .Z(n1612));
Q_AN02 U4013 ( .A0(n35), .A1(n1613), .Z(gcm_dak_cmd_in_nxt[461]));
Q_MX02 U4014 ( .S(n90), .A0(gcm_dak_cmd_in[397]), .A1(gcm_dak_cmd_in[461]), .Z(n1613));
Q_AN02 U4015 ( .A0(n35), .A1(n1614), .Z(gcm_dak_cmd_in_nxt[460]));
Q_MX02 U4016 ( .S(n90), .A0(gcm_dak_cmd_in[396]), .A1(gcm_dak_cmd_in[460]), .Z(n1614));
Q_AN02 U4017 ( .A0(n35), .A1(n1615), .Z(gcm_dak_cmd_in_nxt[459]));
Q_MX02 U4018 ( .S(n90), .A0(gcm_dak_cmd_in[395]), .A1(gcm_dak_cmd_in[459]), .Z(n1615));
Q_AN02 U4019 ( .A0(n35), .A1(n1616), .Z(gcm_dak_cmd_in_nxt[458]));
Q_MX02 U4020 ( .S(n90), .A0(gcm_dak_cmd_in[394]), .A1(gcm_dak_cmd_in[458]), .Z(n1616));
Q_AN02 U4021 ( .A0(n35), .A1(n1617), .Z(gcm_dak_cmd_in_nxt[457]));
Q_MX02 U4022 ( .S(n90), .A0(gcm_dak_cmd_in[393]), .A1(gcm_dak_cmd_in[457]), .Z(n1617));
Q_AN02 U4023 ( .A0(n35), .A1(n1618), .Z(gcm_dak_cmd_in_nxt[456]));
Q_MX02 U4024 ( .S(n90), .A0(gcm_dak_cmd_in[392]), .A1(gcm_dak_cmd_in[456]), .Z(n1618));
Q_AN02 U4025 ( .A0(n35), .A1(n1619), .Z(gcm_dak_cmd_in_nxt[455]));
Q_MX02 U4026 ( .S(n90), .A0(gcm_dak_cmd_in[391]), .A1(gcm_dak_cmd_in[455]), .Z(n1619));
Q_AN02 U4027 ( .A0(n35), .A1(n1620), .Z(gcm_dak_cmd_in_nxt[454]));
Q_MX02 U4028 ( .S(n90), .A0(gcm_dak_cmd_in[390]), .A1(gcm_dak_cmd_in[454]), .Z(n1620));
Q_AN02 U4029 ( .A0(n35), .A1(n1621), .Z(gcm_dak_cmd_in_nxt[453]));
Q_MX02 U4030 ( .S(n90), .A0(gcm_dak_cmd_in[389]), .A1(gcm_dak_cmd_in[453]), .Z(n1621));
Q_AN02 U4031 ( .A0(n35), .A1(n1622), .Z(gcm_dak_cmd_in_nxt[452]));
Q_MX02 U4032 ( .S(n90), .A0(gcm_dak_cmd_in[388]), .A1(gcm_dak_cmd_in[452]), .Z(n1622));
Q_AN02 U4033 ( .A0(n35), .A1(n1623), .Z(gcm_dak_cmd_in_nxt[451]));
Q_MX02 U4034 ( .S(n90), .A0(gcm_dak_cmd_in[387]), .A1(gcm_dak_cmd_in[451]), .Z(n1623));
Q_AN02 U4035 ( .A0(n35), .A1(n1624), .Z(gcm_dak_cmd_in_nxt[450]));
Q_MX02 U4036 ( .S(n90), .A0(gcm_dak_cmd_in[386]), .A1(gcm_dak_cmd_in[450]), .Z(n1624));
Q_AN02 U4037 ( .A0(n35), .A1(n1625), .Z(gcm_dak_cmd_in_nxt[449]));
Q_MX02 U4038 ( .S(n90), .A0(gcm_dak_cmd_in[385]), .A1(gcm_dak_cmd_in[449]), .Z(n1625));
Q_AN02 U4039 ( .A0(n35), .A1(n1626), .Z(gcm_dak_cmd_in_nxt[448]));
Q_MX02 U4040 ( .S(n90), .A0(gcm_dak_cmd_in[384]), .A1(gcm_dak_cmd_in[448]), .Z(n1626));
Q_AN02 U4041 ( .A0(n35), .A1(n1627), .Z(gcm_dak_cmd_in_nxt[447]));
Q_MX02 U4042 ( .S(n90), .A0(gcm_dak_cmd_in[383]), .A1(gcm_dak_cmd_in[447]), .Z(n1627));
Q_AN02 U4043 ( .A0(n35), .A1(n1628), .Z(gcm_dak_cmd_in_nxt[446]));
Q_MX02 U4044 ( .S(n90), .A0(gcm_dak_cmd_in[382]), .A1(gcm_dak_cmd_in[446]), .Z(n1628));
Q_AN02 U4045 ( .A0(n35), .A1(n1629), .Z(gcm_dak_cmd_in_nxt[445]));
Q_MX02 U4046 ( .S(n90), .A0(gcm_dak_cmd_in[381]), .A1(gcm_dak_cmd_in[445]), .Z(n1629));
Q_AN02 U4047 ( .A0(n35), .A1(n1630), .Z(gcm_dak_cmd_in_nxt[444]));
Q_MX02 U4048 ( .S(n90), .A0(gcm_dak_cmd_in[380]), .A1(gcm_dak_cmd_in[444]), .Z(n1630));
Q_AN02 U4049 ( .A0(n35), .A1(n1631), .Z(gcm_dak_cmd_in_nxt[443]));
Q_MX02 U4050 ( .S(n90), .A0(gcm_dak_cmd_in[379]), .A1(gcm_dak_cmd_in[443]), .Z(n1631));
Q_AN02 U4051 ( .A0(n35), .A1(n1632), .Z(gcm_dak_cmd_in_nxt[442]));
Q_MX02 U4052 ( .S(n90), .A0(gcm_dak_cmd_in[378]), .A1(gcm_dak_cmd_in[442]), .Z(n1632));
Q_AN02 U4053 ( .A0(n35), .A1(n1633), .Z(gcm_dak_cmd_in_nxt[441]));
Q_MX02 U4054 ( .S(n90), .A0(gcm_dak_cmd_in[377]), .A1(gcm_dak_cmd_in[441]), .Z(n1633));
Q_AN02 U4055 ( .A0(n35), .A1(n1634), .Z(gcm_dak_cmd_in_nxt[440]));
Q_MX02 U4056 ( .S(n90), .A0(gcm_dak_cmd_in[376]), .A1(gcm_dak_cmd_in[440]), .Z(n1634));
Q_AN02 U4057 ( .A0(n35), .A1(n1635), .Z(gcm_dak_cmd_in_nxt[439]));
Q_MX02 U4058 ( .S(n90), .A0(gcm_dak_cmd_in[375]), .A1(gcm_dak_cmd_in[439]), .Z(n1635));
Q_AN02 U4059 ( .A0(n35), .A1(n1636), .Z(gcm_dak_cmd_in_nxt[438]));
Q_MX02 U4060 ( .S(n90), .A0(gcm_dak_cmd_in[374]), .A1(gcm_dak_cmd_in[438]), .Z(n1636));
Q_AN02 U4061 ( .A0(n35), .A1(n1637), .Z(gcm_dak_cmd_in_nxt[437]));
Q_MX02 U4062 ( .S(n90), .A0(gcm_dak_cmd_in[373]), .A1(gcm_dak_cmd_in[437]), .Z(n1637));
Q_AN02 U4063 ( .A0(n35), .A1(n1638), .Z(gcm_dak_cmd_in_nxt[436]));
Q_MX02 U4064 ( .S(n90), .A0(gcm_dak_cmd_in[372]), .A1(gcm_dak_cmd_in[436]), .Z(n1638));
Q_AN02 U4065 ( .A0(n35), .A1(n1639), .Z(gcm_dak_cmd_in_nxt[435]));
Q_MX02 U4066 ( .S(n90), .A0(gcm_dak_cmd_in[371]), .A1(gcm_dak_cmd_in[435]), .Z(n1639));
Q_AN02 U4067 ( .A0(n35), .A1(n1640), .Z(gcm_dak_cmd_in_nxt[434]));
Q_MX02 U4068 ( .S(n90), .A0(gcm_dak_cmd_in[370]), .A1(gcm_dak_cmd_in[434]), .Z(n1640));
Q_AN02 U4069 ( .A0(n35), .A1(n1641), .Z(gcm_dak_cmd_in_nxt[433]));
Q_MX02 U4070 ( .S(n90), .A0(gcm_dak_cmd_in[369]), .A1(gcm_dak_cmd_in[433]), .Z(n1641));
Q_AN02 U4071 ( .A0(n35), .A1(n1642), .Z(gcm_dak_cmd_in_nxt[432]));
Q_MX02 U4072 ( .S(n90), .A0(gcm_dak_cmd_in[368]), .A1(gcm_dak_cmd_in[432]), .Z(n1642));
Q_AN02 U4073 ( .A0(n35), .A1(n1643), .Z(gcm_dak_cmd_in_nxt[431]));
Q_MX02 U4074 ( .S(n90), .A0(gcm_dak_cmd_in[367]), .A1(gcm_dak_cmd_in[431]), .Z(n1643));
Q_AN02 U4075 ( .A0(n35), .A1(n1644), .Z(gcm_dak_cmd_in_nxt[430]));
Q_MX02 U4076 ( .S(n90), .A0(gcm_dak_cmd_in[366]), .A1(gcm_dak_cmd_in[430]), .Z(n1644));
Q_AN02 U4077 ( .A0(n35), .A1(n1645), .Z(gcm_dak_cmd_in_nxt[429]));
Q_MX02 U4078 ( .S(n90), .A0(gcm_dak_cmd_in[365]), .A1(gcm_dak_cmd_in[429]), .Z(n1645));
Q_AN02 U4079 ( .A0(n35), .A1(n1646), .Z(gcm_dak_cmd_in_nxt[428]));
Q_MX02 U4080 ( .S(n90), .A0(gcm_dak_cmd_in[364]), .A1(gcm_dak_cmd_in[428]), .Z(n1646));
Q_AN02 U4081 ( .A0(n35), .A1(n1647), .Z(gcm_dak_cmd_in_nxt[427]));
Q_MX02 U4082 ( .S(n90), .A0(gcm_dak_cmd_in[363]), .A1(gcm_dak_cmd_in[427]), .Z(n1647));
Q_AN02 U4083 ( .A0(n35), .A1(n1648), .Z(gcm_dak_cmd_in_nxt[426]));
Q_MX02 U4084 ( .S(n90), .A0(gcm_dak_cmd_in[362]), .A1(gcm_dak_cmd_in[426]), .Z(n1648));
Q_AN02 U4085 ( .A0(n35), .A1(n1649), .Z(gcm_dak_cmd_in_nxt[425]));
Q_MX02 U4086 ( .S(n90), .A0(gcm_dak_cmd_in[361]), .A1(gcm_dak_cmd_in[425]), .Z(n1649));
Q_AN02 U4087 ( .A0(n35), .A1(n1650), .Z(gcm_dak_cmd_in_nxt[424]));
Q_MX02 U4088 ( .S(n90), .A0(gcm_dak_cmd_in[360]), .A1(gcm_dak_cmd_in[424]), .Z(n1650));
Q_AN02 U4089 ( .A0(n35), .A1(n1651), .Z(gcm_dak_cmd_in_nxt[423]));
Q_MX02 U4090 ( .S(n90), .A0(gcm_dak_cmd_in[359]), .A1(gcm_dak_cmd_in[423]), .Z(n1651));
Q_AN02 U4091 ( .A0(n35), .A1(n1652), .Z(gcm_dak_cmd_in_nxt[422]));
Q_MX02 U4092 ( .S(n90), .A0(gcm_dak_cmd_in[358]), .A1(gcm_dak_cmd_in[422]), .Z(n1652));
Q_AN02 U4093 ( .A0(n35), .A1(n1653), .Z(gcm_dak_cmd_in_nxt[421]));
Q_MX02 U4094 ( .S(n90), .A0(gcm_dak_cmd_in[357]), .A1(gcm_dak_cmd_in[421]), .Z(n1653));
Q_AN02 U4095 ( .A0(n35), .A1(n1654), .Z(gcm_dak_cmd_in_nxt[420]));
Q_MX02 U4096 ( .S(n90), .A0(gcm_dak_cmd_in[356]), .A1(gcm_dak_cmd_in[420]), .Z(n1654));
Q_AN02 U4097 ( .A0(n35), .A1(n1655), .Z(gcm_dak_cmd_in_nxt[419]));
Q_MX02 U4098 ( .S(n90), .A0(gcm_dak_cmd_in[355]), .A1(gcm_dak_cmd_in[419]), .Z(n1655));
Q_AN02 U4099 ( .A0(n35), .A1(n1656), .Z(gcm_dak_cmd_in_nxt[418]));
Q_MX02 U4100 ( .S(n90), .A0(kme_internal_out[63]), .A1(gcm_dak_cmd_in[418]), .Z(n1656));
Q_AN02 U4101 ( .A0(n35), .A1(n1657), .Z(gcm_dak_cmd_in_nxt[417]));
Q_MX02 U4102 ( .S(n90), .A0(kme_internal_out[62]), .A1(gcm_dak_cmd_in[417]), .Z(n1657));
Q_AN02 U4103 ( .A0(n35), .A1(n1658), .Z(gcm_dak_cmd_in_nxt[416]));
Q_MX02 U4104 ( .S(n90), .A0(kme_internal_out[61]), .A1(gcm_dak_cmd_in[416]), .Z(n1658));
Q_AN02 U4105 ( .A0(n35), .A1(n1659), .Z(gcm_dak_cmd_in_nxt[415]));
Q_MX02 U4106 ( .S(n90), .A0(kme_internal_out[60]), .A1(gcm_dak_cmd_in[415]), .Z(n1659));
Q_AN02 U4107 ( .A0(n35), .A1(n1660), .Z(gcm_dak_cmd_in_nxt[414]));
Q_MX02 U4108 ( .S(n90), .A0(kme_internal_out[59]), .A1(gcm_dak_cmd_in[414]), .Z(n1660));
Q_AN02 U4109 ( .A0(n35), .A1(n1661), .Z(gcm_dak_cmd_in_nxt[413]));
Q_MX02 U4110 ( .S(n90), .A0(kme_internal_out[58]), .A1(gcm_dak_cmd_in[413]), .Z(n1661));
Q_AN02 U4111 ( .A0(n35), .A1(n1662), .Z(gcm_dak_cmd_in_nxt[412]));
Q_MX02 U4112 ( .S(n90), .A0(kme_internal_out[57]), .A1(gcm_dak_cmd_in[412]), .Z(n1662));
Q_AN02 U4113 ( .A0(n35), .A1(n1663), .Z(gcm_dak_cmd_in_nxt[411]));
Q_MX02 U4114 ( .S(n90), .A0(kme_internal_out[56]), .A1(gcm_dak_cmd_in[411]), .Z(n1663));
Q_AN02 U4115 ( .A0(n35), .A1(n1664), .Z(gcm_dak_cmd_in_nxt[410]));
Q_MX02 U4116 ( .S(n90), .A0(kme_internal_out[55]), .A1(gcm_dak_cmd_in[410]), .Z(n1664));
Q_AN02 U4117 ( .A0(n35), .A1(n1665), .Z(gcm_dak_cmd_in_nxt[409]));
Q_MX02 U4118 ( .S(n90), .A0(kme_internal_out[54]), .A1(gcm_dak_cmd_in[409]), .Z(n1665));
Q_AN02 U4119 ( .A0(n35), .A1(n1666), .Z(gcm_dak_cmd_in_nxt[408]));
Q_MX02 U4120 ( .S(n90), .A0(kme_internal_out[53]), .A1(gcm_dak_cmd_in[408]), .Z(n1666));
Q_AN02 U4121 ( .A0(n35), .A1(n1667), .Z(gcm_dak_cmd_in_nxt[407]));
Q_MX02 U4122 ( .S(n90), .A0(kme_internal_out[52]), .A1(gcm_dak_cmd_in[407]), .Z(n1667));
Q_AN02 U4123 ( .A0(n35), .A1(n1668), .Z(gcm_dak_cmd_in_nxt[406]));
Q_MX02 U4124 ( .S(n90), .A0(kme_internal_out[51]), .A1(gcm_dak_cmd_in[406]), .Z(n1668));
Q_AN02 U4125 ( .A0(n35), .A1(n1669), .Z(gcm_dak_cmd_in_nxt[405]));
Q_MX02 U4126 ( .S(n90), .A0(kme_internal_out[50]), .A1(gcm_dak_cmd_in[405]), .Z(n1669));
Q_AN02 U4127 ( .A0(n35), .A1(n1670), .Z(gcm_dak_cmd_in_nxt[404]));
Q_MX02 U4128 ( .S(n90), .A0(kme_internal_out[49]), .A1(gcm_dak_cmd_in[404]), .Z(n1670));
Q_AN02 U4129 ( .A0(n35), .A1(n1671), .Z(gcm_dak_cmd_in_nxt[403]));
Q_MX02 U4130 ( .S(n90), .A0(kme_internal_out[48]), .A1(gcm_dak_cmd_in[403]), .Z(n1671));
Q_AN02 U4131 ( .A0(n35), .A1(n1672), .Z(gcm_dak_cmd_in_nxt[402]));
Q_MX02 U4132 ( .S(n90), .A0(kme_internal_out[47]), .A1(gcm_dak_cmd_in[402]), .Z(n1672));
Q_AN02 U4133 ( .A0(n35), .A1(n1673), .Z(gcm_dak_cmd_in_nxt[401]));
Q_MX02 U4134 ( .S(n90), .A0(kme_internal_out[46]), .A1(gcm_dak_cmd_in[401]), .Z(n1673));
Q_AN02 U4135 ( .A0(n35), .A1(n1674), .Z(gcm_dak_cmd_in_nxt[400]));
Q_MX02 U4136 ( .S(n90), .A0(kme_internal_out[45]), .A1(gcm_dak_cmd_in[400]), .Z(n1674));
Q_AN02 U4137 ( .A0(n35), .A1(n1675), .Z(gcm_dak_cmd_in_nxt[399]));
Q_MX02 U4138 ( .S(n90), .A0(kme_internal_out[44]), .A1(gcm_dak_cmd_in[399]), .Z(n1675));
Q_AN02 U4139 ( .A0(n35), .A1(n1676), .Z(gcm_dak_cmd_in_nxt[398]));
Q_MX02 U4140 ( .S(n90), .A0(kme_internal_out[43]), .A1(gcm_dak_cmd_in[398]), .Z(n1676));
Q_AN02 U4141 ( .A0(n35), .A1(n1677), .Z(gcm_dak_cmd_in_nxt[397]));
Q_MX02 U4142 ( .S(n90), .A0(kme_internal_out[42]), .A1(gcm_dak_cmd_in[397]), .Z(n1677));
Q_AN02 U4143 ( .A0(n35), .A1(n1678), .Z(gcm_dak_cmd_in_nxt[396]));
Q_MX02 U4144 ( .S(n90), .A0(kme_internal_out[41]), .A1(gcm_dak_cmd_in[396]), .Z(n1678));
Q_AN02 U4145 ( .A0(n35), .A1(n1679), .Z(gcm_dak_cmd_in_nxt[395]));
Q_MX02 U4146 ( .S(n90), .A0(kme_internal_out[40]), .A1(gcm_dak_cmd_in[395]), .Z(n1679));
Q_AN02 U4147 ( .A0(n35), .A1(n1680), .Z(gcm_dak_cmd_in_nxt[394]));
Q_MX02 U4148 ( .S(n90), .A0(kme_internal_out[39]), .A1(gcm_dak_cmd_in[394]), .Z(n1680));
Q_AN02 U4149 ( .A0(n35), .A1(n1681), .Z(gcm_dak_cmd_in_nxt[393]));
Q_MX02 U4150 ( .S(n90), .A0(kme_internal_out[38]), .A1(gcm_dak_cmd_in[393]), .Z(n1681));
Q_AN02 U4151 ( .A0(n35), .A1(n1682), .Z(gcm_dak_cmd_in_nxt[392]));
Q_MX02 U4152 ( .S(n90), .A0(kme_internal_out[37]), .A1(gcm_dak_cmd_in[392]), .Z(n1682));
Q_AN02 U4153 ( .A0(n35), .A1(n1683), .Z(gcm_dak_cmd_in_nxt[391]));
Q_MX02 U4154 ( .S(n90), .A0(kme_internal_out[36]), .A1(gcm_dak_cmd_in[391]), .Z(n1683));
Q_AN02 U4155 ( .A0(n35), .A1(n1684), .Z(gcm_dak_cmd_in_nxt[390]));
Q_MX02 U4156 ( .S(n90), .A0(kme_internal_out[35]), .A1(gcm_dak_cmd_in[390]), .Z(n1684));
Q_AN02 U4157 ( .A0(n35), .A1(n1685), .Z(gcm_dak_cmd_in_nxt[389]));
Q_MX02 U4158 ( .S(n90), .A0(kme_internal_out[34]), .A1(gcm_dak_cmd_in[389]), .Z(n1685));
Q_AN02 U4159 ( .A0(n35), .A1(n1686), .Z(gcm_dak_cmd_in_nxt[388]));
Q_MX02 U4160 ( .S(n90), .A0(kme_internal_out[33]), .A1(gcm_dak_cmd_in[388]), .Z(n1686));
Q_AN02 U4161 ( .A0(n35), .A1(n1687), .Z(gcm_dak_cmd_in_nxt[387]));
Q_MX02 U4162 ( .S(n90), .A0(kme_internal_out[32]), .A1(gcm_dak_cmd_in[387]), .Z(n1687));
Q_AN02 U4163 ( .A0(n35), .A1(n1688), .Z(gcm_dak_cmd_in_nxt[386]));
Q_MX02 U4164 ( .S(n90), .A0(kme_internal_out[31]), .A1(gcm_dak_cmd_in[386]), .Z(n1688));
Q_AN02 U4165 ( .A0(n35), .A1(n1689), .Z(gcm_dak_cmd_in_nxt[385]));
Q_MX02 U4166 ( .S(n90), .A0(kme_internal_out[30]), .A1(gcm_dak_cmd_in[385]), .Z(n1689));
Q_AN02 U4167 ( .A0(n35), .A1(n1690), .Z(gcm_dak_cmd_in_nxt[384]));
Q_MX02 U4168 ( .S(n90), .A0(kme_internal_out[29]), .A1(gcm_dak_cmd_in[384]), .Z(n1690));
Q_AN02 U4169 ( .A0(n35), .A1(n1691), .Z(gcm_dak_cmd_in_nxt[383]));
Q_MX02 U4170 ( .S(n90), .A0(kme_internal_out[28]), .A1(gcm_dak_cmd_in[383]), .Z(n1691));
Q_AN02 U4171 ( .A0(n35), .A1(n1692), .Z(gcm_dak_cmd_in_nxt[382]));
Q_MX02 U4172 ( .S(n90), .A0(kme_internal_out[27]), .A1(gcm_dak_cmd_in[382]), .Z(n1692));
Q_AN02 U4173 ( .A0(n35), .A1(n1693), .Z(gcm_dak_cmd_in_nxt[381]));
Q_MX02 U4174 ( .S(n90), .A0(kme_internal_out[26]), .A1(gcm_dak_cmd_in[381]), .Z(n1693));
Q_AN02 U4175 ( .A0(n35), .A1(n1694), .Z(gcm_dak_cmd_in_nxt[380]));
Q_MX02 U4176 ( .S(n90), .A0(kme_internal_out[25]), .A1(gcm_dak_cmd_in[380]), .Z(n1694));
Q_AN02 U4177 ( .A0(n35), .A1(n1695), .Z(gcm_dak_cmd_in_nxt[379]));
Q_MX02 U4178 ( .S(n90), .A0(kme_internal_out[24]), .A1(gcm_dak_cmd_in[379]), .Z(n1695));
Q_AN02 U4179 ( .A0(n35), .A1(n1696), .Z(gcm_dak_cmd_in_nxt[378]));
Q_MX02 U4180 ( .S(n90), .A0(kme_internal_out[23]), .A1(gcm_dak_cmd_in[378]), .Z(n1696));
Q_AN02 U4181 ( .A0(n35), .A1(n1697), .Z(gcm_dak_cmd_in_nxt[377]));
Q_MX02 U4182 ( .S(n90), .A0(kme_internal_out[22]), .A1(gcm_dak_cmd_in[377]), .Z(n1697));
Q_AN02 U4183 ( .A0(n35), .A1(n1698), .Z(gcm_dak_cmd_in_nxt[376]));
Q_MX02 U4184 ( .S(n90), .A0(kme_internal_out[21]), .A1(gcm_dak_cmd_in[376]), .Z(n1698));
Q_AN02 U4185 ( .A0(n35), .A1(n1699), .Z(gcm_dak_cmd_in_nxt[375]));
Q_MX02 U4186 ( .S(n90), .A0(kme_internal_out[20]), .A1(gcm_dak_cmd_in[375]), .Z(n1699));
Q_AN02 U4187 ( .A0(n35), .A1(n1700), .Z(gcm_dak_cmd_in_nxt[374]));
Q_MX02 U4188 ( .S(n90), .A0(kme_internal_out[19]), .A1(gcm_dak_cmd_in[374]), .Z(n1700));
Q_AN02 U4189 ( .A0(n35), .A1(n1701), .Z(gcm_dak_cmd_in_nxt[373]));
Q_MX02 U4190 ( .S(n90), .A0(kme_internal_out[18]), .A1(gcm_dak_cmd_in[373]), .Z(n1701));
Q_AN02 U4191 ( .A0(n35), .A1(n1702), .Z(gcm_dak_cmd_in_nxt[372]));
Q_MX02 U4192 ( .S(n90), .A0(kme_internal_out[17]), .A1(gcm_dak_cmd_in[372]), .Z(n1702));
Q_AN02 U4193 ( .A0(n35), .A1(n1703), .Z(gcm_dak_cmd_in_nxt[371]));
Q_MX02 U4194 ( .S(n90), .A0(kme_internal_out[16]), .A1(gcm_dak_cmd_in[371]), .Z(n1703));
Q_AN02 U4195 ( .A0(n35), .A1(n1704), .Z(gcm_dak_cmd_in_nxt[370]));
Q_MX02 U4196 ( .S(n90), .A0(kme_internal_out[15]), .A1(gcm_dak_cmd_in[370]), .Z(n1704));
Q_AN02 U4197 ( .A0(n35), .A1(n1705), .Z(gcm_dak_cmd_in_nxt[369]));
Q_MX02 U4198 ( .S(n90), .A0(kme_internal_out[14]), .A1(gcm_dak_cmd_in[369]), .Z(n1705));
Q_AN02 U4199 ( .A0(n35), .A1(n1706), .Z(gcm_dak_cmd_in_nxt[368]));
Q_MX02 U4200 ( .S(n90), .A0(kme_internal_out[13]), .A1(gcm_dak_cmd_in[368]), .Z(n1706));
Q_AN02 U4201 ( .A0(n35), .A1(n1707), .Z(gcm_dak_cmd_in_nxt[367]));
Q_MX02 U4202 ( .S(n90), .A0(kme_internal_out[12]), .A1(gcm_dak_cmd_in[367]), .Z(n1707));
Q_AN02 U4203 ( .A0(n35), .A1(n1708), .Z(gcm_dak_cmd_in_nxt[366]));
Q_MX02 U4204 ( .S(n90), .A0(kme_internal_out[11]), .A1(gcm_dak_cmd_in[366]), .Z(n1708));
Q_AN02 U4205 ( .A0(n35), .A1(n1709), .Z(gcm_dak_cmd_in_nxt[365]));
Q_MX02 U4206 ( .S(n90), .A0(kme_internal_out[10]), .A1(gcm_dak_cmd_in[365]), .Z(n1709));
Q_AN02 U4207 ( .A0(n35), .A1(n1710), .Z(gcm_dak_cmd_in_nxt[364]));
Q_MX02 U4208 ( .S(n90), .A0(kme_internal_out[9]), .A1(gcm_dak_cmd_in[364]), .Z(n1710));
Q_AN02 U4209 ( .A0(n35), .A1(n1711), .Z(gcm_dak_cmd_in_nxt[363]));
Q_MX02 U4210 ( .S(n90), .A0(kme_internal_out[8]), .A1(gcm_dak_cmd_in[363]), .Z(n1711));
Q_AN02 U4211 ( .A0(n35), .A1(n1712), .Z(gcm_dak_cmd_in_nxt[362]));
Q_MX02 U4212 ( .S(n90), .A0(kme_internal_out[7]), .A1(gcm_dak_cmd_in[362]), .Z(n1712));
Q_AN02 U4213 ( .A0(n35), .A1(n1713), .Z(gcm_dak_cmd_in_nxt[361]));
Q_MX02 U4214 ( .S(n90), .A0(kme_internal_out[6]), .A1(gcm_dak_cmd_in[361]), .Z(n1713));
Q_AN02 U4215 ( .A0(n35), .A1(n1714), .Z(gcm_dak_cmd_in_nxt[360]));
Q_MX02 U4216 ( .S(n90), .A0(kme_internal_out[5]), .A1(gcm_dak_cmd_in[360]), .Z(n1714));
Q_AN02 U4217 ( .A0(n35), .A1(n1715), .Z(gcm_dak_cmd_in_nxt[359]));
Q_MX02 U4218 ( .S(n90), .A0(kme_internal_out[4]), .A1(gcm_dak_cmd_in[359]), .Z(n1715));
Q_AN02 U4219 ( .A0(n35), .A1(n1716), .Z(gcm_dak_cmd_in_nxt[358]));
Q_MX02 U4220 ( .S(n90), .A0(kme_internal_out[3]), .A1(gcm_dak_cmd_in[358]), .Z(n1716));
Q_AN02 U4221 ( .A0(n35), .A1(n1717), .Z(gcm_dak_cmd_in_nxt[357]));
Q_MX02 U4222 ( .S(n90), .A0(kme_internal_out[2]), .A1(gcm_dak_cmd_in[357]), .Z(n1717));
Q_AN02 U4223 ( .A0(n35), .A1(n1718), .Z(gcm_dak_cmd_in_nxt[356]));
Q_MX02 U4224 ( .S(n90), .A0(kme_internal_out[1]), .A1(gcm_dak_cmd_in[356]), .Z(n1718));
Q_AN02 U4225 ( .A0(n35), .A1(n1719), .Z(gcm_dak_cmd_in_nxt[355]));
Q_MX02 U4226 ( .S(n90), .A0(kme_internal_out[0]), .A1(gcm_dak_cmd_in[355]), .Z(n1719));
Q_AO21 U4227 ( .A0(n1720), .A1(gcm_dek_cmd_in[0]), .B0(n1724), .Z(gcm_dek_cmd_in_nxt[0]));
Q_AO21 U4228 ( .A0(n1720), .A1(gcm_dek_cmd_in[1]), .B0(n1723), .Z(gcm_dek_cmd_in_nxt[1]));
Q_AO21 U4229 ( .A0(n1720), .A1(gcm_dek_cmd_in[2]), .B0(n1721), .Z(gcm_dek_cmd_in_nxt[2]));
Q_AN02 U4230 ( .A0(n37), .A1(n38), .Z(n1720));
Q_XOR2 U4231 ( .A0(n38), .A1(n115), .Z(n1722));
Q_NR02 U4232 ( .A0(n37), .A1(n1722), .Z(n1721));
Q_MX02 U4233 ( .S(n37), .A0(n36), .A1(n1722), .Z(n1723));
Q_MX02 U4234 ( .S(n37), .A0(n38), .A1(n36), .Z(n1724));
Q_AN03 U4235 ( .A0(n38), .A1(n1725), .A2(n37), .Z(gcm_dek_cmd_in_nxt[34]));
Q_MX02 U4236 ( .S(n120), .A0(n2621), .A1(gcm_dek_cmd_in[34]), .Z(n1725));
Q_AN03 U4237 ( .A0(n38), .A1(n1726), .A2(n37), .Z(gcm_dek_cmd_in_nxt[33]));
Q_MX02 U4238 ( .S(n120), .A0(n2622), .A1(gcm_dek_cmd_in[33]), .Z(n1726));
Q_AN03 U4239 ( .A0(n38), .A1(n1727), .A2(n37), .Z(gcm_dek_cmd_in_nxt[32]));
Q_MX02 U4240 ( .S(n120), .A0(n2623), .A1(gcm_dek_cmd_in[32]), .Z(n1727));
Q_AN03 U4241 ( .A0(n38), .A1(n1728), .A2(n37), .Z(gcm_dek_cmd_in_nxt[31]));
Q_MX02 U4242 ( .S(n120), .A0(n2624), .A1(gcm_dek_cmd_in[31]), .Z(n1728));
Q_AN03 U4243 ( .A0(n38), .A1(n1729), .A2(n37), .Z(gcm_dek_cmd_in_nxt[30]));
Q_MX02 U4244 ( .S(n120), .A0(n2625), .A1(gcm_dek_cmd_in[30]), .Z(n1729));
Q_AN03 U4245 ( .A0(n38), .A1(n1730), .A2(n37), .Z(gcm_dek_cmd_in_nxt[29]));
Q_MX02 U4246 ( .S(n120), .A0(n2626), .A1(gcm_dek_cmd_in[29]), .Z(n1730));
Q_AN03 U4247 ( .A0(n38), .A1(n1731), .A2(n37), .Z(gcm_dek_cmd_in_nxt[28]));
Q_MX02 U4248 ( .S(n120), .A0(n2627), .A1(gcm_dek_cmd_in[28]), .Z(n1731));
Q_AN03 U4249 ( .A0(n38), .A1(n1732), .A2(n37), .Z(gcm_dek_cmd_in_nxt[27]));
Q_MX02 U4250 ( .S(n120), .A0(n2628), .A1(gcm_dek_cmd_in[27]), .Z(n1732));
Q_AN03 U4251 ( .A0(n38), .A1(n1733), .A2(n37), .Z(gcm_dek_cmd_in_nxt[26]));
Q_MX02 U4252 ( .S(n120), .A0(n2629), .A1(gcm_dek_cmd_in[26]), .Z(n1733));
Q_AN03 U4253 ( .A0(n38), .A1(n1734), .A2(n37), .Z(gcm_dek_cmd_in_nxt[25]));
Q_MX02 U4254 ( .S(n120), .A0(n2630), .A1(gcm_dek_cmd_in[25]), .Z(n1734));
Q_AN03 U4255 ( .A0(n38), .A1(n1735), .A2(n37), .Z(gcm_dek_cmd_in_nxt[24]));
Q_MX02 U4256 ( .S(n120), .A0(n2631), .A1(gcm_dek_cmd_in[24]), .Z(n1735));
Q_AN03 U4257 ( .A0(n38), .A1(n1736), .A2(n37), .Z(gcm_dek_cmd_in_nxt[23]));
Q_MX02 U4258 ( .S(n120), .A0(n2632), .A1(gcm_dek_cmd_in[23]), .Z(n1736));
Q_AN03 U4259 ( .A0(n38), .A1(n1737), .A2(n37), .Z(gcm_dek_cmd_in_nxt[22]));
Q_MX02 U4260 ( .S(n120), .A0(n2633), .A1(gcm_dek_cmd_in[22]), .Z(n1737));
Q_AN03 U4261 ( .A0(n38), .A1(n1738), .A2(n37), .Z(gcm_dek_cmd_in_nxt[21]));
Q_MX02 U4262 ( .S(n120), .A0(n2634), .A1(gcm_dek_cmd_in[21]), .Z(n1738));
Q_AN03 U4263 ( .A0(n38), .A1(n1739), .A2(n37), .Z(gcm_dek_cmd_in_nxt[20]));
Q_MX02 U4264 ( .S(n120), .A0(n2635), .A1(gcm_dek_cmd_in[20]), .Z(n1739));
Q_AN03 U4265 ( .A0(n38), .A1(n1740), .A2(n37), .Z(gcm_dek_cmd_in_nxt[19]));
Q_MX02 U4266 ( .S(n120), .A0(n2636), .A1(gcm_dek_cmd_in[19]), .Z(n1740));
Q_AN03 U4267 ( .A0(n38), .A1(n1741), .A2(n37), .Z(gcm_dek_cmd_in_nxt[18]));
Q_MX02 U4268 ( .S(n120), .A0(n2637), .A1(gcm_dek_cmd_in[18]), .Z(n1741));
Q_AN03 U4269 ( .A0(n38), .A1(n1742), .A2(n37), .Z(gcm_dek_cmd_in_nxt[17]));
Q_MX02 U4270 ( .S(n120), .A0(n2638), .A1(gcm_dek_cmd_in[17]), .Z(n1742));
Q_AN03 U4271 ( .A0(n38), .A1(n1743), .A2(n37), .Z(gcm_dek_cmd_in_nxt[16]));
Q_MX02 U4272 ( .S(n120), .A0(n2639), .A1(gcm_dek_cmd_in[16]), .Z(n1743));
Q_AN03 U4273 ( .A0(n38), .A1(n1744), .A2(n37), .Z(gcm_dek_cmd_in_nxt[15]));
Q_MX02 U4274 ( .S(n120), .A0(n2640), .A1(gcm_dek_cmd_in[15]), .Z(n1744));
Q_AN03 U4275 ( .A0(n38), .A1(n1745), .A2(n37), .Z(gcm_dek_cmd_in_nxt[14]));
Q_MX02 U4276 ( .S(n120), .A0(n2641), .A1(gcm_dek_cmd_in[14]), .Z(n1745));
Q_AN03 U4277 ( .A0(n38), .A1(n1746), .A2(n37), .Z(gcm_dek_cmd_in_nxt[13]));
Q_MX02 U4278 ( .S(n120), .A0(n2642), .A1(gcm_dek_cmd_in[13]), .Z(n1746));
Q_AN03 U4279 ( .A0(n38), .A1(n1747), .A2(n37), .Z(gcm_dek_cmd_in_nxt[12]));
Q_MX02 U4280 ( .S(n120), .A0(n2643), .A1(gcm_dek_cmd_in[12]), .Z(n1747));
Q_AN03 U4281 ( .A0(n38), .A1(n1748), .A2(n37), .Z(gcm_dek_cmd_in_nxt[11]));
Q_MX02 U4282 ( .S(n120), .A0(n2644), .A1(gcm_dek_cmd_in[11]), .Z(n1748));
Q_AN03 U4283 ( .A0(n38), .A1(n1749), .A2(n37), .Z(gcm_dek_cmd_in_nxt[10]));
Q_MX02 U4284 ( .S(n120), .A0(n2645), .A1(gcm_dek_cmd_in[10]), .Z(n1749));
Q_AN03 U4285 ( .A0(n38), .A1(n1750), .A2(n37), .Z(gcm_dek_cmd_in_nxt[9]));
Q_MX02 U4286 ( .S(n120), .A0(n2646), .A1(gcm_dek_cmd_in[9]), .Z(n1750));
Q_AN03 U4287 ( .A0(n38), .A1(n1751), .A2(n37), .Z(gcm_dek_cmd_in_nxt[8]));
Q_MX02 U4288 ( .S(n120), .A0(n2647), .A1(gcm_dek_cmd_in[8]), .Z(n1751));
Q_AN03 U4289 ( .A0(n38), .A1(n1752), .A2(n37), .Z(gcm_dek_cmd_in_nxt[7]));
Q_MX02 U4290 ( .S(n120), .A0(n2648), .A1(gcm_dek_cmd_in[7]), .Z(n1752));
Q_AN03 U4291 ( .A0(n38), .A1(n1753), .A2(n37), .Z(gcm_dek_cmd_in_nxt[6]));
Q_MX02 U4292 ( .S(n120), .A0(n2649), .A1(gcm_dek_cmd_in[6]), .Z(n1753));
Q_AN03 U4293 ( .A0(n38), .A1(n1754), .A2(n37), .Z(gcm_dek_cmd_in_nxt[5]));
Q_MX02 U4294 ( .S(n120), .A0(n2650), .A1(gcm_dek_cmd_in[5]), .Z(n1754));
Q_AN03 U4295 ( .A0(n38), .A1(n1755), .A2(n37), .Z(gcm_dek_cmd_in_nxt[4]));
Q_MX02 U4296 ( .S(n120), .A0(n2651), .A1(gcm_dek_cmd_in[4]), .Z(n1755));
Q_AN03 U4297 ( .A0(n38), .A1(n1756), .A2(n37), .Z(gcm_dek_cmd_in_nxt[3]));
Q_MX02 U4298 ( .S(n120), .A0(n2652), .A1(gcm_dek_cmd_in[3]), .Z(n1756));
Q_AN03 U4299 ( .A0(n38), .A1(n1757), .A2(n37), .Z(gcm_dek_cmd_in_nxt[98]));
Q_MX02 U4300 ( .S(n120), .A0(n2653), .A1(gcm_dek_cmd_in[98]), .Z(n1757));
Q_AN03 U4301 ( .A0(n38), .A1(n1758), .A2(n37), .Z(gcm_dek_cmd_in_nxt[97]));
Q_MX02 U4302 ( .S(n120), .A0(n2654), .A1(gcm_dek_cmd_in[97]), .Z(n1758));
Q_AN03 U4303 ( .A0(n38), .A1(n1759), .A2(n37), .Z(gcm_dek_cmd_in_nxt[96]));
Q_MX02 U4304 ( .S(n120), .A0(n2655), .A1(gcm_dek_cmd_in[96]), .Z(n1759));
Q_AN03 U4305 ( .A0(n38), .A1(n1760), .A2(n37), .Z(gcm_dek_cmd_in_nxt[95]));
Q_MX02 U4306 ( .S(n120), .A0(n2656), .A1(gcm_dek_cmd_in[95]), .Z(n1760));
Q_AN03 U4307 ( .A0(n38), .A1(n1761), .A2(n37), .Z(gcm_dek_cmd_in_nxt[94]));
Q_MX02 U4308 ( .S(n120), .A0(n2657), .A1(gcm_dek_cmd_in[94]), .Z(n1761));
Q_AN03 U4309 ( .A0(n38), .A1(n1762), .A2(n37), .Z(gcm_dek_cmd_in_nxt[93]));
Q_MX02 U4310 ( .S(n120), .A0(n2658), .A1(gcm_dek_cmd_in[93]), .Z(n1762));
Q_AN03 U4311 ( .A0(n38), .A1(n1763), .A2(n37), .Z(gcm_dek_cmd_in_nxt[92]));
Q_MX02 U4312 ( .S(n120), .A0(n2659), .A1(gcm_dek_cmd_in[92]), .Z(n1763));
Q_AN03 U4313 ( .A0(n38), .A1(n1764), .A2(n37), .Z(gcm_dek_cmd_in_nxt[91]));
Q_MX02 U4314 ( .S(n120), .A0(n2660), .A1(gcm_dek_cmd_in[91]), .Z(n1764));
Q_AN03 U4315 ( .A0(n38), .A1(n1765), .A2(n37), .Z(gcm_dek_cmd_in_nxt[90]));
Q_MX02 U4316 ( .S(n120), .A0(n2661), .A1(gcm_dek_cmd_in[90]), .Z(n1765));
Q_AN03 U4317 ( .A0(n38), .A1(n1766), .A2(n37), .Z(gcm_dek_cmd_in_nxt[89]));
Q_MX02 U4318 ( .S(n120), .A0(n2662), .A1(gcm_dek_cmd_in[89]), .Z(n1766));
Q_AN03 U4319 ( .A0(n38), .A1(n1767), .A2(n37), .Z(gcm_dek_cmd_in_nxt[88]));
Q_MX02 U4320 ( .S(n120), .A0(n2663), .A1(gcm_dek_cmd_in[88]), .Z(n1767));
Q_AN03 U4321 ( .A0(n38), .A1(n1768), .A2(n37), .Z(gcm_dek_cmd_in_nxt[87]));
Q_MX02 U4322 ( .S(n120), .A0(n2664), .A1(gcm_dek_cmd_in[87]), .Z(n1768));
Q_AN03 U4323 ( .A0(n38), .A1(n1769), .A2(n37), .Z(gcm_dek_cmd_in_nxt[86]));
Q_MX02 U4324 ( .S(n120), .A0(n2665), .A1(gcm_dek_cmd_in[86]), .Z(n1769));
Q_AN03 U4325 ( .A0(n38), .A1(n1770), .A2(n37), .Z(gcm_dek_cmd_in_nxt[85]));
Q_MX02 U4326 ( .S(n120), .A0(n2666), .A1(gcm_dek_cmd_in[85]), .Z(n1770));
Q_AN03 U4327 ( .A0(n38), .A1(n1771), .A2(n37), .Z(gcm_dek_cmd_in_nxt[84]));
Q_MX02 U4328 ( .S(n120), .A0(n2667), .A1(gcm_dek_cmd_in[84]), .Z(n1771));
Q_AN03 U4329 ( .A0(n38), .A1(n1772), .A2(n37), .Z(gcm_dek_cmd_in_nxt[83]));
Q_MX02 U4330 ( .S(n120), .A0(n2668), .A1(gcm_dek_cmd_in[83]), .Z(n1772));
Q_AN03 U4331 ( .A0(n38), .A1(n1773), .A2(n37), .Z(gcm_dek_cmd_in_nxt[82]));
Q_MX02 U4332 ( .S(n120), .A0(n2669), .A1(gcm_dek_cmd_in[82]), .Z(n1773));
Q_AN03 U4333 ( .A0(n38), .A1(n1774), .A2(n37), .Z(gcm_dek_cmd_in_nxt[81]));
Q_MX02 U4334 ( .S(n120), .A0(n2670), .A1(gcm_dek_cmd_in[81]), .Z(n1774));
Q_AN03 U4335 ( .A0(n38), .A1(n1775), .A2(n37), .Z(gcm_dek_cmd_in_nxt[80]));
Q_MX02 U4336 ( .S(n120), .A0(n2671), .A1(gcm_dek_cmd_in[80]), .Z(n1775));
Q_AN03 U4337 ( .A0(n38), .A1(n1776), .A2(n37), .Z(gcm_dek_cmd_in_nxt[79]));
Q_MX02 U4338 ( .S(n120), .A0(n2672), .A1(gcm_dek_cmd_in[79]), .Z(n1776));
Q_AN03 U4339 ( .A0(n38), .A1(n1777), .A2(n37), .Z(gcm_dek_cmd_in_nxt[78]));
Q_MX02 U4340 ( .S(n120), .A0(n2673), .A1(gcm_dek_cmd_in[78]), .Z(n1777));
Q_AN03 U4341 ( .A0(n38), .A1(n1778), .A2(n37), .Z(gcm_dek_cmd_in_nxt[77]));
Q_MX02 U4342 ( .S(n120), .A0(n2674), .A1(gcm_dek_cmd_in[77]), .Z(n1778));
Q_AN03 U4343 ( .A0(n38), .A1(n1779), .A2(n37), .Z(gcm_dek_cmd_in_nxt[76]));
Q_MX02 U4344 ( .S(n120), .A0(n2675), .A1(gcm_dek_cmd_in[76]), .Z(n1779));
Q_AN03 U4345 ( .A0(n38), .A1(n1780), .A2(n37), .Z(gcm_dek_cmd_in_nxt[75]));
Q_MX02 U4346 ( .S(n120), .A0(n2676), .A1(gcm_dek_cmd_in[75]), .Z(n1780));
Q_AN03 U4347 ( .A0(n38), .A1(n1781), .A2(n37), .Z(gcm_dek_cmd_in_nxt[74]));
Q_MX02 U4348 ( .S(n120), .A0(n2677), .A1(gcm_dek_cmd_in[74]), .Z(n1781));
Q_AN03 U4349 ( .A0(n38), .A1(n1782), .A2(n37), .Z(gcm_dek_cmd_in_nxt[73]));
Q_MX02 U4350 ( .S(n120), .A0(n2678), .A1(gcm_dek_cmd_in[73]), .Z(n1782));
Q_AN03 U4351 ( .A0(n38), .A1(n1783), .A2(n37), .Z(gcm_dek_cmd_in_nxt[72]));
Q_MX02 U4352 ( .S(n120), .A0(n2679), .A1(gcm_dek_cmd_in[72]), .Z(n1783));
Q_AN03 U4353 ( .A0(n38), .A1(n1784), .A2(n37), .Z(gcm_dek_cmd_in_nxt[71]));
Q_MX02 U4354 ( .S(n120), .A0(n2680), .A1(gcm_dek_cmd_in[71]), .Z(n1784));
Q_AN03 U4355 ( .A0(n38), .A1(n1785), .A2(n37), .Z(gcm_dek_cmd_in_nxt[70]));
Q_MX02 U4356 ( .S(n120), .A0(n2681), .A1(gcm_dek_cmd_in[70]), .Z(n1785));
Q_AN03 U4357 ( .A0(n38), .A1(n1786), .A2(n37), .Z(gcm_dek_cmd_in_nxt[69]));
Q_MX02 U4358 ( .S(n120), .A0(n2682), .A1(gcm_dek_cmd_in[69]), .Z(n1786));
Q_AN03 U4359 ( .A0(n38), .A1(n1787), .A2(n37), .Z(gcm_dek_cmd_in_nxt[68]));
Q_MX02 U4360 ( .S(n120), .A0(n2683), .A1(gcm_dek_cmd_in[68]), .Z(n1787));
Q_AN03 U4361 ( .A0(n38), .A1(n1788), .A2(n37), .Z(gcm_dek_cmd_in_nxt[67]));
Q_MX02 U4362 ( .S(n120), .A0(n2684), .A1(gcm_dek_cmd_in[67]), .Z(n1788));
Q_AN03 U4363 ( .A0(n38), .A1(n1789), .A2(n37), .Z(gcm_dek_cmd_in_nxt[66]));
Q_MX02 U4364 ( .S(n120), .A0(n2685), .A1(gcm_dek_cmd_in[66]), .Z(n1789));
Q_AN03 U4365 ( .A0(n38), .A1(n1790), .A2(n37), .Z(gcm_dek_cmd_in_nxt[65]));
Q_MX02 U4366 ( .S(n120), .A0(n2686), .A1(gcm_dek_cmd_in[65]), .Z(n1790));
Q_AN03 U4367 ( .A0(n38), .A1(n1791), .A2(n37), .Z(gcm_dek_cmd_in_nxt[64]));
Q_MX02 U4368 ( .S(n120), .A0(n2687), .A1(gcm_dek_cmd_in[64]), .Z(n1791));
Q_AN03 U4369 ( .A0(n38), .A1(n1792), .A2(n37), .Z(gcm_dek_cmd_in_nxt[63]));
Q_MX02 U4370 ( .S(n120), .A0(n2688), .A1(gcm_dek_cmd_in[63]), .Z(n1792));
Q_AN03 U4371 ( .A0(n38), .A1(n1793), .A2(n37), .Z(gcm_dek_cmd_in_nxt[62]));
Q_MX02 U4372 ( .S(n120), .A0(n2689), .A1(gcm_dek_cmd_in[62]), .Z(n1793));
Q_AN03 U4373 ( .A0(n38), .A1(n1794), .A2(n37), .Z(gcm_dek_cmd_in_nxt[61]));
Q_MX02 U4374 ( .S(n120), .A0(n2690), .A1(gcm_dek_cmd_in[61]), .Z(n1794));
Q_AN03 U4375 ( .A0(n38), .A1(n1795), .A2(n37), .Z(gcm_dek_cmd_in_nxt[60]));
Q_MX02 U4376 ( .S(n120), .A0(n2691), .A1(gcm_dek_cmd_in[60]), .Z(n1795));
Q_AN03 U4377 ( .A0(n38), .A1(n1796), .A2(n37), .Z(gcm_dek_cmd_in_nxt[59]));
Q_MX02 U4378 ( .S(n120), .A0(n2692), .A1(gcm_dek_cmd_in[59]), .Z(n1796));
Q_AN03 U4379 ( .A0(n38), .A1(n1797), .A2(n37), .Z(gcm_dek_cmd_in_nxt[58]));
Q_MX02 U4380 ( .S(n120), .A0(n2693), .A1(gcm_dek_cmd_in[58]), .Z(n1797));
Q_AN03 U4381 ( .A0(n38), .A1(n1798), .A2(n37), .Z(gcm_dek_cmd_in_nxt[57]));
Q_MX02 U4382 ( .S(n120), .A0(n2694), .A1(gcm_dek_cmd_in[57]), .Z(n1798));
Q_AN03 U4383 ( .A0(n38), .A1(n1799), .A2(n37), .Z(gcm_dek_cmd_in_nxt[56]));
Q_MX02 U4384 ( .S(n120), .A0(n2695), .A1(gcm_dek_cmd_in[56]), .Z(n1799));
Q_AN03 U4385 ( .A0(n38), .A1(n1800), .A2(n37), .Z(gcm_dek_cmd_in_nxt[55]));
Q_MX02 U4386 ( .S(n120), .A0(n2696), .A1(gcm_dek_cmd_in[55]), .Z(n1800));
Q_AN03 U4387 ( .A0(n38), .A1(n1801), .A2(n37), .Z(gcm_dek_cmd_in_nxt[54]));
Q_MX02 U4388 ( .S(n120), .A0(n2697), .A1(gcm_dek_cmd_in[54]), .Z(n1801));
Q_AN03 U4389 ( .A0(n38), .A1(n1802), .A2(n37), .Z(gcm_dek_cmd_in_nxt[53]));
Q_MX02 U4390 ( .S(n120), .A0(n2698), .A1(gcm_dek_cmd_in[53]), .Z(n1802));
Q_AN03 U4391 ( .A0(n38), .A1(n1803), .A2(n37), .Z(gcm_dek_cmd_in_nxt[52]));
Q_MX02 U4392 ( .S(n120), .A0(n2699), .A1(gcm_dek_cmd_in[52]), .Z(n1803));
Q_AN03 U4393 ( .A0(n38), .A1(n1804), .A2(n37), .Z(gcm_dek_cmd_in_nxt[51]));
Q_MX02 U4394 ( .S(n120), .A0(n2700), .A1(gcm_dek_cmd_in[51]), .Z(n1804));
Q_AN03 U4395 ( .A0(n38), .A1(n1805), .A2(n37), .Z(gcm_dek_cmd_in_nxt[50]));
Q_MX02 U4396 ( .S(n120), .A0(n2701), .A1(gcm_dek_cmd_in[50]), .Z(n1805));
Q_AN03 U4397 ( .A0(n38), .A1(n1806), .A2(n37), .Z(gcm_dek_cmd_in_nxt[49]));
Q_MX02 U4398 ( .S(n120), .A0(n2702), .A1(gcm_dek_cmd_in[49]), .Z(n1806));
Q_AN03 U4399 ( .A0(n38), .A1(n1807), .A2(n37), .Z(gcm_dek_cmd_in_nxt[48]));
Q_MX02 U4400 ( .S(n120), .A0(n2703), .A1(gcm_dek_cmd_in[48]), .Z(n1807));
Q_AN03 U4401 ( .A0(n38), .A1(n1808), .A2(n37), .Z(gcm_dek_cmd_in_nxt[47]));
Q_MX02 U4402 ( .S(n120), .A0(n2704), .A1(gcm_dek_cmd_in[47]), .Z(n1808));
Q_AN03 U4403 ( .A0(n38), .A1(n1809), .A2(n37), .Z(gcm_dek_cmd_in_nxt[46]));
Q_MX02 U4404 ( .S(n120), .A0(n2705), .A1(gcm_dek_cmd_in[46]), .Z(n1809));
Q_AN03 U4405 ( .A0(n38), .A1(n1810), .A2(n37), .Z(gcm_dek_cmd_in_nxt[45]));
Q_MX02 U4406 ( .S(n120), .A0(n2706), .A1(gcm_dek_cmd_in[45]), .Z(n1810));
Q_AN03 U4407 ( .A0(n38), .A1(n1811), .A2(n37), .Z(gcm_dek_cmd_in_nxt[44]));
Q_MX02 U4408 ( .S(n120), .A0(n2707), .A1(gcm_dek_cmd_in[44]), .Z(n1811));
Q_AN03 U4409 ( .A0(n38), .A1(n1812), .A2(n37), .Z(gcm_dek_cmd_in_nxt[43]));
Q_MX02 U4410 ( .S(n120), .A0(n2708), .A1(gcm_dek_cmd_in[43]), .Z(n1812));
Q_AN03 U4411 ( .A0(n38), .A1(n1813), .A2(n37), .Z(gcm_dek_cmd_in_nxt[42]));
Q_MX02 U4412 ( .S(n120), .A0(n2709), .A1(gcm_dek_cmd_in[42]), .Z(n1813));
Q_AN03 U4413 ( .A0(n38), .A1(n1814), .A2(n37), .Z(gcm_dek_cmd_in_nxt[41]));
Q_MX02 U4414 ( .S(n120), .A0(n2710), .A1(gcm_dek_cmd_in[41]), .Z(n1814));
Q_AN03 U4415 ( .A0(n38), .A1(n1815), .A2(n37), .Z(gcm_dek_cmd_in_nxt[40]));
Q_MX02 U4416 ( .S(n120), .A0(n2711), .A1(gcm_dek_cmd_in[40]), .Z(n1815));
Q_AN03 U4417 ( .A0(n38), .A1(n1816), .A2(n37), .Z(gcm_dek_cmd_in_nxt[39]));
Q_MX02 U4418 ( .S(n120), .A0(n2712), .A1(gcm_dek_cmd_in[39]), .Z(n1816));
Q_AN03 U4419 ( .A0(n38), .A1(n1817), .A2(n37), .Z(gcm_dek_cmd_in_nxt[38]));
Q_MX02 U4420 ( .S(n120), .A0(n2713), .A1(gcm_dek_cmd_in[38]), .Z(n1817));
Q_AN03 U4421 ( .A0(n38), .A1(n1818), .A2(n37), .Z(gcm_dek_cmd_in_nxt[37]));
Q_MX02 U4422 ( .S(n120), .A0(n2714), .A1(gcm_dek_cmd_in[37]), .Z(n1818));
Q_AN03 U4423 ( .A0(n38), .A1(n1819), .A2(n37), .Z(gcm_dek_cmd_in_nxt[36]));
Q_MX02 U4424 ( .S(n120), .A0(n2715), .A1(gcm_dek_cmd_in[36]), .Z(n1819));
Q_AN03 U4425 ( .A0(n38), .A1(n1820), .A2(n37), .Z(gcm_dek_cmd_in_nxt[35]));
Q_MX02 U4426 ( .S(n120), .A0(n2716), .A1(gcm_dek_cmd_in[35]), .Z(n1820));
Q_AN03 U4427 ( .A0(n38), .A1(n1821), .A2(n37), .Z(gcm_dek_cmd_in_nxt[354]));
Q_MX02 U4428 ( .S(n124), .A0(gcm_dek_cmd_in[290]), .A1(gcm_dek_cmd_in[354]), .Z(n1821));
Q_AN03 U4429 ( .A0(n38), .A1(n1822), .A2(n37), .Z(gcm_dek_cmd_in_nxt[353]));
Q_MX02 U4430 ( .S(n124), .A0(gcm_dek_cmd_in[289]), .A1(gcm_dek_cmd_in[353]), .Z(n1822));
Q_AN03 U4431 ( .A0(n38), .A1(n1823), .A2(n37), .Z(gcm_dek_cmd_in_nxt[352]));
Q_MX02 U4432 ( .S(n124), .A0(gcm_dek_cmd_in[288]), .A1(gcm_dek_cmd_in[352]), .Z(n1823));
Q_AN03 U4433 ( .A0(n38), .A1(n1824), .A2(n37), .Z(gcm_dek_cmd_in_nxt[351]));
Q_MX02 U4434 ( .S(n124), .A0(gcm_dek_cmd_in[287]), .A1(gcm_dek_cmd_in[351]), .Z(n1824));
Q_AN03 U4435 ( .A0(n38), .A1(n1825), .A2(n37), .Z(gcm_dek_cmd_in_nxt[350]));
Q_MX02 U4436 ( .S(n124), .A0(gcm_dek_cmd_in[286]), .A1(gcm_dek_cmd_in[350]), .Z(n1825));
Q_AN03 U4437 ( .A0(n38), .A1(n1826), .A2(n37), .Z(gcm_dek_cmd_in_nxt[349]));
Q_MX02 U4438 ( .S(n124), .A0(gcm_dek_cmd_in[285]), .A1(gcm_dek_cmd_in[349]), .Z(n1826));
Q_AN03 U4439 ( .A0(n38), .A1(n1827), .A2(n37), .Z(gcm_dek_cmd_in_nxt[348]));
Q_MX02 U4440 ( .S(n124), .A0(gcm_dek_cmd_in[284]), .A1(gcm_dek_cmd_in[348]), .Z(n1827));
Q_AN03 U4441 ( .A0(n38), .A1(n1828), .A2(n37), .Z(gcm_dek_cmd_in_nxt[347]));
Q_MX02 U4442 ( .S(n124), .A0(gcm_dek_cmd_in[283]), .A1(gcm_dek_cmd_in[347]), .Z(n1828));
Q_AN03 U4443 ( .A0(n38), .A1(n1829), .A2(n37), .Z(gcm_dek_cmd_in_nxt[346]));
Q_MX02 U4444 ( .S(n124), .A0(gcm_dek_cmd_in[282]), .A1(gcm_dek_cmd_in[346]), .Z(n1829));
Q_AN03 U4445 ( .A0(n38), .A1(n1830), .A2(n37), .Z(gcm_dek_cmd_in_nxt[345]));
Q_MX02 U4446 ( .S(n124), .A0(gcm_dek_cmd_in[281]), .A1(gcm_dek_cmd_in[345]), .Z(n1830));
Q_AN03 U4447 ( .A0(n38), .A1(n1831), .A2(n37), .Z(gcm_dek_cmd_in_nxt[344]));
Q_MX02 U4448 ( .S(n124), .A0(gcm_dek_cmd_in[280]), .A1(gcm_dek_cmd_in[344]), .Z(n1831));
Q_AN03 U4449 ( .A0(n38), .A1(n1832), .A2(n37), .Z(gcm_dek_cmd_in_nxt[343]));
Q_MX02 U4450 ( .S(n124), .A0(gcm_dek_cmd_in[279]), .A1(gcm_dek_cmd_in[343]), .Z(n1832));
Q_AN03 U4451 ( .A0(n38), .A1(n1833), .A2(n37), .Z(gcm_dek_cmd_in_nxt[342]));
Q_MX02 U4452 ( .S(n124), .A0(gcm_dek_cmd_in[278]), .A1(gcm_dek_cmd_in[342]), .Z(n1833));
Q_AN03 U4453 ( .A0(n38), .A1(n1834), .A2(n37), .Z(gcm_dek_cmd_in_nxt[341]));
Q_MX02 U4454 ( .S(n124), .A0(gcm_dek_cmd_in[277]), .A1(gcm_dek_cmd_in[341]), .Z(n1834));
Q_AN03 U4455 ( .A0(n38), .A1(n1835), .A2(n37), .Z(gcm_dek_cmd_in_nxt[340]));
Q_MX02 U4456 ( .S(n124), .A0(gcm_dek_cmd_in[276]), .A1(gcm_dek_cmd_in[340]), .Z(n1835));
Q_AN03 U4457 ( .A0(n38), .A1(n1836), .A2(n37), .Z(gcm_dek_cmd_in_nxt[339]));
Q_MX02 U4458 ( .S(n124), .A0(gcm_dek_cmd_in[275]), .A1(gcm_dek_cmd_in[339]), .Z(n1836));
Q_AN03 U4459 ( .A0(n38), .A1(n1837), .A2(n37), .Z(gcm_dek_cmd_in_nxt[338]));
Q_MX02 U4460 ( .S(n124), .A0(gcm_dek_cmd_in[274]), .A1(gcm_dek_cmd_in[338]), .Z(n1837));
Q_AN03 U4461 ( .A0(n38), .A1(n1838), .A2(n37), .Z(gcm_dek_cmd_in_nxt[337]));
Q_MX02 U4462 ( .S(n124), .A0(gcm_dek_cmd_in[273]), .A1(gcm_dek_cmd_in[337]), .Z(n1838));
Q_AN03 U4463 ( .A0(n38), .A1(n1839), .A2(n37), .Z(gcm_dek_cmd_in_nxt[336]));
Q_MX02 U4464 ( .S(n124), .A0(gcm_dek_cmd_in[272]), .A1(gcm_dek_cmd_in[336]), .Z(n1839));
Q_AN03 U4465 ( .A0(n38), .A1(n1840), .A2(n37), .Z(gcm_dek_cmd_in_nxt[335]));
Q_MX02 U4466 ( .S(n124), .A0(gcm_dek_cmd_in[271]), .A1(gcm_dek_cmd_in[335]), .Z(n1840));
Q_AN03 U4467 ( .A0(n38), .A1(n1841), .A2(n37), .Z(gcm_dek_cmd_in_nxt[334]));
Q_MX02 U4468 ( .S(n124), .A0(gcm_dek_cmd_in[270]), .A1(gcm_dek_cmd_in[334]), .Z(n1841));
Q_AN03 U4469 ( .A0(n38), .A1(n1842), .A2(n37), .Z(gcm_dek_cmd_in_nxt[333]));
Q_MX02 U4470 ( .S(n124), .A0(gcm_dek_cmd_in[269]), .A1(gcm_dek_cmd_in[333]), .Z(n1842));
Q_AN03 U4471 ( .A0(n38), .A1(n1843), .A2(n37), .Z(gcm_dek_cmd_in_nxt[332]));
Q_MX02 U4472 ( .S(n124), .A0(gcm_dek_cmd_in[268]), .A1(gcm_dek_cmd_in[332]), .Z(n1843));
Q_AN03 U4473 ( .A0(n38), .A1(n1844), .A2(n37), .Z(gcm_dek_cmd_in_nxt[331]));
Q_MX02 U4474 ( .S(n124), .A0(gcm_dek_cmd_in[267]), .A1(gcm_dek_cmd_in[331]), .Z(n1844));
Q_AN03 U4475 ( .A0(n38), .A1(n1845), .A2(n37), .Z(gcm_dek_cmd_in_nxt[330]));
Q_MX02 U4476 ( .S(n124), .A0(gcm_dek_cmd_in[266]), .A1(gcm_dek_cmd_in[330]), .Z(n1845));
Q_AN03 U4477 ( .A0(n38), .A1(n1846), .A2(n37), .Z(gcm_dek_cmd_in_nxt[329]));
Q_MX02 U4478 ( .S(n124), .A0(gcm_dek_cmd_in[265]), .A1(gcm_dek_cmd_in[329]), .Z(n1846));
Q_AN03 U4479 ( .A0(n38), .A1(n1847), .A2(n37), .Z(gcm_dek_cmd_in_nxt[328]));
Q_MX02 U4480 ( .S(n124), .A0(gcm_dek_cmd_in[264]), .A1(gcm_dek_cmd_in[328]), .Z(n1847));
Q_AN03 U4481 ( .A0(n38), .A1(n1848), .A2(n37), .Z(gcm_dek_cmd_in_nxt[327]));
Q_MX02 U4482 ( .S(n124), .A0(gcm_dek_cmd_in[263]), .A1(gcm_dek_cmd_in[327]), .Z(n1848));
Q_AN03 U4483 ( .A0(n38), .A1(n1849), .A2(n37), .Z(gcm_dek_cmd_in_nxt[326]));
Q_MX02 U4484 ( .S(n124), .A0(gcm_dek_cmd_in[262]), .A1(gcm_dek_cmd_in[326]), .Z(n1849));
Q_AN03 U4485 ( .A0(n38), .A1(n1850), .A2(n37), .Z(gcm_dek_cmd_in_nxt[325]));
Q_MX02 U4486 ( .S(n124), .A0(gcm_dek_cmd_in[261]), .A1(gcm_dek_cmd_in[325]), .Z(n1850));
Q_AN03 U4487 ( .A0(n38), .A1(n1851), .A2(n37), .Z(gcm_dek_cmd_in_nxt[324]));
Q_MX02 U4488 ( .S(n124), .A0(gcm_dek_cmd_in[260]), .A1(gcm_dek_cmd_in[324]), .Z(n1851));
Q_AN03 U4489 ( .A0(n38), .A1(n1852), .A2(n37), .Z(gcm_dek_cmd_in_nxt[323]));
Q_MX02 U4490 ( .S(n124), .A0(gcm_dek_cmd_in[259]), .A1(gcm_dek_cmd_in[323]), .Z(n1852));
Q_AN03 U4491 ( .A0(n38), .A1(n1853), .A2(n37), .Z(gcm_dek_cmd_in_nxt[322]));
Q_MX02 U4492 ( .S(n124), .A0(gcm_dek_cmd_in[258]), .A1(gcm_dek_cmd_in[322]), .Z(n1853));
Q_AN03 U4493 ( .A0(n38), .A1(n1854), .A2(n37), .Z(gcm_dek_cmd_in_nxt[321]));
Q_MX02 U4494 ( .S(n124), .A0(gcm_dek_cmd_in[257]), .A1(gcm_dek_cmd_in[321]), .Z(n1854));
Q_AN03 U4495 ( .A0(n38), .A1(n1855), .A2(n37), .Z(gcm_dek_cmd_in_nxt[320]));
Q_MX02 U4496 ( .S(n124), .A0(gcm_dek_cmd_in[256]), .A1(gcm_dek_cmd_in[320]), .Z(n1855));
Q_AN03 U4497 ( .A0(n38), .A1(n1856), .A2(n37), .Z(gcm_dek_cmd_in_nxt[319]));
Q_MX02 U4498 ( .S(n124), .A0(gcm_dek_cmd_in[255]), .A1(gcm_dek_cmd_in[319]), .Z(n1856));
Q_AN03 U4499 ( .A0(n38), .A1(n1857), .A2(n37), .Z(gcm_dek_cmd_in_nxt[318]));
Q_MX02 U4500 ( .S(n124), .A0(gcm_dek_cmd_in[254]), .A1(gcm_dek_cmd_in[318]), .Z(n1857));
Q_AN03 U4501 ( .A0(n38), .A1(n1858), .A2(n37), .Z(gcm_dek_cmd_in_nxt[317]));
Q_MX02 U4502 ( .S(n124), .A0(gcm_dek_cmd_in[253]), .A1(gcm_dek_cmd_in[317]), .Z(n1858));
Q_AN03 U4503 ( .A0(n38), .A1(n1859), .A2(n37), .Z(gcm_dek_cmd_in_nxt[316]));
Q_MX02 U4504 ( .S(n124), .A0(gcm_dek_cmd_in[252]), .A1(gcm_dek_cmd_in[316]), .Z(n1859));
Q_AN03 U4505 ( .A0(n38), .A1(n1860), .A2(n37), .Z(gcm_dek_cmd_in_nxt[315]));
Q_MX02 U4506 ( .S(n124), .A0(gcm_dek_cmd_in[251]), .A1(gcm_dek_cmd_in[315]), .Z(n1860));
Q_AN03 U4507 ( .A0(n38), .A1(n1861), .A2(n37), .Z(gcm_dek_cmd_in_nxt[314]));
Q_MX02 U4508 ( .S(n124), .A0(gcm_dek_cmd_in[250]), .A1(gcm_dek_cmd_in[314]), .Z(n1861));
Q_AN03 U4509 ( .A0(n38), .A1(n1862), .A2(n37), .Z(gcm_dek_cmd_in_nxt[313]));
Q_MX02 U4510 ( .S(n124), .A0(gcm_dek_cmd_in[249]), .A1(gcm_dek_cmd_in[313]), .Z(n1862));
Q_AN03 U4511 ( .A0(n38), .A1(n1863), .A2(n37), .Z(gcm_dek_cmd_in_nxt[312]));
Q_MX02 U4512 ( .S(n124), .A0(gcm_dek_cmd_in[248]), .A1(gcm_dek_cmd_in[312]), .Z(n1863));
Q_AN03 U4513 ( .A0(n38), .A1(n1864), .A2(n37), .Z(gcm_dek_cmd_in_nxt[311]));
Q_MX02 U4514 ( .S(n124), .A0(gcm_dek_cmd_in[247]), .A1(gcm_dek_cmd_in[311]), .Z(n1864));
Q_AN03 U4515 ( .A0(n38), .A1(n1865), .A2(n37), .Z(gcm_dek_cmd_in_nxt[310]));
Q_MX02 U4516 ( .S(n124), .A0(gcm_dek_cmd_in[246]), .A1(gcm_dek_cmd_in[310]), .Z(n1865));
Q_AN03 U4517 ( .A0(n38), .A1(n1866), .A2(n37), .Z(gcm_dek_cmd_in_nxt[309]));
Q_MX02 U4518 ( .S(n124), .A0(gcm_dek_cmd_in[245]), .A1(gcm_dek_cmd_in[309]), .Z(n1866));
Q_AN03 U4519 ( .A0(n38), .A1(n1867), .A2(n37), .Z(gcm_dek_cmd_in_nxt[308]));
Q_MX02 U4520 ( .S(n124), .A0(gcm_dek_cmd_in[244]), .A1(gcm_dek_cmd_in[308]), .Z(n1867));
Q_AN03 U4521 ( .A0(n38), .A1(n1868), .A2(n37), .Z(gcm_dek_cmd_in_nxt[307]));
Q_MX02 U4522 ( .S(n124), .A0(gcm_dek_cmd_in[243]), .A1(gcm_dek_cmd_in[307]), .Z(n1868));
Q_AN03 U4523 ( .A0(n38), .A1(n1869), .A2(n37), .Z(gcm_dek_cmd_in_nxt[306]));
Q_MX02 U4524 ( .S(n124), .A0(gcm_dek_cmd_in[242]), .A1(gcm_dek_cmd_in[306]), .Z(n1869));
Q_AN03 U4525 ( .A0(n38), .A1(n1870), .A2(n37), .Z(gcm_dek_cmd_in_nxt[305]));
Q_MX02 U4526 ( .S(n124), .A0(gcm_dek_cmd_in[241]), .A1(gcm_dek_cmd_in[305]), .Z(n1870));
Q_AN03 U4527 ( .A0(n38), .A1(n1871), .A2(n37), .Z(gcm_dek_cmd_in_nxt[304]));
Q_MX02 U4528 ( .S(n124), .A0(gcm_dek_cmd_in[240]), .A1(gcm_dek_cmd_in[304]), .Z(n1871));
Q_AN03 U4529 ( .A0(n38), .A1(n1872), .A2(n37), .Z(gcm_dek_cmd_in_nxt[303]));
Q_MX02 U4530 ( .S(n124), .A0(gcm_dek_cmd_in[239]), .A1(gcm_dek_cmd_in[303]), .Z(n1872));
Q_AN03 U4531 ( .A0(n38), .A1(n1873), .A2(n37), .Z(gcm_dek_cmd_in_nxt[302]));
Q_MX02 U4532 ( .S(n124), .A0(gcm_dek_cmd_in[238]), .A1(gcm_dek_cmd_in[302]), .Z(n1873));
Q_AN03 U4533 ( .A0(n38), .A1(n1874), .A2(n37), .Z(gcm_dek_cmd_in_nxt[301]));
Q_MX02 U4534 ( .S(n124), .A0(gcm_dek_cmd_in[237]), .A1(gcm_dek_cmd_in[301]), .Z(n1874));
Q_AN03 U4535 ( .A0(n38), .A1(n1875), .A2(n37), .Z(gcm_dek_cmd_in_nxt[300]));
Q_MX02 U4536 ( .S(n124), .A0(gcm_dek_cmd_in[236]), .A1(gcm_dek_cmd_in[300]), .Z(n1875));
Q_AN03 U4537 ( .A0(n38), .A1(n1876), .A2(n37), .Z(gcm_dek_cmd_in_nxt[299]));
Q_MX02 U4538 ( .S(n124), .A0(gcm_dek_cmd_in[235]), .A1(gcm_dek_cmd_in[299]), .Z(n1876));
Q_AN03 U4539 ( .A0(n38), .A1(n1877), .A2(n37), .Z(gcm_dek_cmd_in_nxt[298]));
Q_MX02 U4540 ( .S(n124), .A0(gcm_dek_cmd_in[234]), .A1(gcm_dek_cmd_in[298]), .Z(n1877));
Q_AN03 U4541 ( .A0(n38), .A1(n1878), .A2(n37), .Z(gcm_dek_cmd_in_nxt[297]));
Q_MX02 U4542 ( .S(n124), .A0(gcm_dek_cmd_in[233]), .A1(gcm_dek_cmd_in[297]), .Z(n1878));
Q_AN03 U4543 ( .A0(n38), .A1(n1879), .A2(n37), .Z(gcm_dek_cmd_in_nxt[296]));
Q_MX02 U4544 ( .S(n124), .A0(gcm_dek_cmd_in[232]), .A1(gcm_dek_cmd_in[296]), .Z(n1879));
Q_AN03 U4545 ( .A0(n38), .A1(n1880), .A2(n37), .Z(gcm_dek_cmd_in_nxt[295]));
Q_MX02 U4546 ( .S(n124), .A0(gcm_dek_cmd_in[231]), .A1(gcm_dek_cmd_in[295]), .Z(n1880));
Q_AN03 U4547 ( .A0(n38), .A1(n1881), .A2(n37), .Z(gcm_dek_cmd_in_nxt[294]));
Q_MX02 U4548 ( .S(n124), .A0(gcm_dek_cmd_in[230]), .A1(gcm_dek_cmd_in[294]), .Z(n1881));
Q_AN03 U4549 ( .A0(n38), .A1(n1882), .A2(n37), .Z(gcm_dek_cmd_in_nxt[293]));
Q_MX02 U4550 ( .S(n124), .A0(gcm_dek_cmd_in[229]), .A1(gcm_dek_cmd_in[293]), .Z(n1882));
Q_AN03 U4551 ( .A0(n38), .A1(n1883), .A2(n37), .Z(gcm_dek_cmd_in_nxt[292]));
Q_MX02 U4552 ( .S(n124), .A0(gcm_dek_cmd_in[228]), .A1(gcm_dek_cmd_in[292]), .Z(n1883));
Q_AN03 U4553 ( .A0(n38), .A1(n1884), .A2(n37), .Z(gcm_dek_cmd_in_nxt[291]));
Q_MX02 U4554 ( .S(n124), .A0(gcm_dek_cmd_in[227]), .A1(gcm_dek_cmd_in[291]), .Z(n1884));
Q_AN03 U4555 ( .A0(n38), .A1(n1885), .A2(n37), .Z(gcm_dek_cmd_in_nxt[290]));
Q_MX02 U4556 ( .S(n124), .A0(gcm_dek_cmd_in[226]), .A1(gcm_dek_cmd_in[290]), .Z(n1885));
Q_AN03 U4557 ( .A0(n38), .A1(n1886), .A2(n37), .Z(gcm_dek_cmd_in_nxt[289]));
Q_MX02 U4558 ( .S(n124), .A0(gcm_dek_cmd_in[225]), .A1(gcm_dek_cmd_in[289]), .Z(n1886));
Q_AN03 U4559 ( .A0(n38), .A1(n1887), .A2(n37), .Z(gcm_dek_cmd_in_nxt[288]));
Q_MX02 U4560 ( .S(n124), .A0(gcm_dek_cmd_in[224]), .A1(gcm_dek_cmd_in[288]), .Z(n1887));
Q_AN03 U4561 ( .A0(n38), .A1(n1888), .A2(n37), .Z(gcm_dek_cmd_in_nxt[287]));
Q_MX02 U4562 ( .S(n124), .A0(gcm_dek_cmd_in[223]), .A1(gcm_dek_cmd_in[287]), .Z(n1888));
Q_AN03 U4563 ( .A0(n38), .A1(n1889), .A2(n37), .Z(gcm_dek_cmd_in_nxt[286]));
Q_MX02 U4564 ( .S(n124), .A0(gcm_dek_cmd_in[222]), .A1(gcm_dek_cmd_in[286]), .Z(n1889));
Q_AN03 U4565 ( .A0(n38), .A1(n1890), .A2(n37), .Z(gcm_dek_cmd_in_nxt[285]));
Q_MX02 U4566 ( .S(n124), .A0(gcm_dek_cmd_in[221]), .A1(gcm_dek_cmd_in[285]), .Z(n1890));
Q_AN03 U4567 ( .A0(n38), .A1(n1891), .A2(n37), .Z(gcm_dek_cmd_in_nxt[284]));
Q_MX02 U4568 ( .S(n124), .A0(gcm_dek_cmd_in[220]), .A1(gcm_dek_cmd_in[284]), .Z(n1891));
Q_AN03 U4569 ( .A0(n38), .A1(n1892), .A2(n37), .Z(gcm_dek_cmd_in_nxt[283]));
Q_MX02 U4570 ( .S(n124), .A0(gcm_dek_cmd_in[219]), .A1(gcm_dek_cmd_in[283]), .Z(n1892));
Q_AN03 U4571 ( .A0(n38), .A1(n1893), .A2(n37), .Z(gcm_dek_cmd_in_nxt[282]));
Q_MX02 U4572 ( .S(n124), .A0(gcm_dek_cmd_in[218]), .A1(gcm_dek_cmd_in[282]), .Z(n1893));
Q_AN03 U4573 ( .A0(n38), .A1(n1894), .A2(n37), .Z(gcm_dek_cmd_in_nxt[281]));
Q_MX02 U4574 ( .S(n124), .A0(gcm_dek_cmd_in[217]), .A1(gcm_dek_cmd_in[281]), .Z(n1894));
Q_AN03 U4575 ( .A0(n38), .A1(n1895), .A2(n37), .Z(gcm_dek_cmd_in_nxt[280]));
Q_MX02 U4576 ( .S(n124), .A0(gcm_dek_cmd_in[216]), .A1(gcm_dek_cmd_in[280]), .Z(n1895));
Q_AN03 U4577 ( .A0(n38), .A1(n1896), .A2(n37), .Z(gcm_dek_cmd_in_nxt[279]));
Q_MX02 U4578 ( .S(n124), .A0(gcm_dek_cmd_in[215]), .A1(gcm_dek_cmd_in[279]), .Z(n1896));
Q_AN03 U4579 ( .A0(n38), .A1(n1897), .A2(n37), .Z(gcm_dek_cmd_in_nxt[278]));
Q_MX02 U4580 ( .S(n124), .A0(gcm_dek_cmd_in[214]), .A1(gcm_dek_cmd_in[278]), .Z(n1897));
Q_AN03 U4581 ( .A0(n38), .A1(n1898), .A2(n37), .Z(gcm_dek_cmd_in_nxt[277]));
Q_MX02 U4582 ( .S(n124), .A0(gcm_dek_cmd_in[213]), .A1(gcm_dek_cmd_in[277]), .Z(n1898));
Q_AN03 U4583 ( .A0(n38), .A1(n1899), .A2(n37), .Z(gcm_dek_cmd_in_nxt[276]));
Q_MX02 U4584 ( .S(n124), .A0(gcm_dek_cmd_in[212]), .A1(gcm_dek_cmd_in[276]), .Z(n1899));
Q_AN03 U4585 ( .A0(n38), .A1(n1900), .A2(n37), .Z(gcm_dek_cmd_in_nxt[275]));
Q_MX02 U4586 ( .S(n124), .A0(gcm_dek_cmd_in[211]), .A1(gcm_dek_cmd_in[275]), .Z(n1900));
Q_AN03 U4587 ( .A0(n38), .A1(n1901), .A2(n37), .Z(gcm_dek_cmd_in_nxt[274]));
Q_MX02 U4588 ( .S(n124), .A0(gcm_dek_cmd_in[210]), .A1(gcm_dek_cmd_in[274]), .Z(n1901));
Q_AN03 U4589 ( .A0(n38), .A1(n1902), .A2(n37), .Z(gcm_dek_cmd_in_nxt[273]));
Q_MX02 U4590 ( .S(n124), .A0(gcm_dek_cmd_in[209]), .A1(gcm_dek_cmd_in[273]), .Z(n1902));
Q_AN03 U4591 ( .A0(n38), .A1(n1903), .A2(n37), .Z(gcm_dek_cmd_in_nxt[272]));
Q_MX02 U4592 ( .S(n124), .A0(gcm_dek_cmd_in[208]), .A1(gcm_dek_cmd_in[272]), .Z(n1903));
Q_AN03 U4593 ( .A0(n38), .A1(n1904), .A2(n37), .Z(gcm_dek_cmd_in_nxt[271]));
Q_MX02 U4594 ( .S(n124), .A0(gcm_dek_cmd_in[207]), .A1(gcm_dek_cmd_in[271]), .Z(n1904));
Q_AN03 U4595 ( .A0(n38), .A1(n1905), .A2(n37), .Z(gcm_dek_cmd_in_nxt[270]));
Q_MX02 U4596 ( .S(n124), .A0(gcm_dek_cmd_in[206]), .A1(gcm_dek_cmd_in[270]), .Z(n1905));
Q_AN03 U4597 ( .A0(n38), .A1(n1906), .A2(n37), .Z(gcm_dek_cmd_in_nxt[269]));
Q_MX02 U4598 ( .S(n124), .A0(gcm_dek_cmd_in[205]), .A1(gcm_dek_cmd_in[269]), .Z(n1906));
Q_AN03 U4599 ( .A0(n38), .A1(n1907), .A2(n37), .Z(gcm_dek_cmd_in_nxt[268]));
Q_MX02 U4600 ( .S(n124), .A0(gcm_dek_cmd_in[204]), .A1(gcm_dek_cmd_in[268]), .Z(n1907));
Q_AN03 U4601 ( .A0(n38), .A1(n1908), .A2(n37), .Z(gcm_dek_cmd_in_nxt[267]));
Q_MX02 U4602 ( .S(n124), .A0(gcm_dek_cmd_in[203]), .A1(gcm_dek_cmd_in[267]), .Z(n1908));
Q_AN03 U4603 ( .A0(n38), .A1(n1909), .A2(n37), .Z(gcm_dek_cmd_in_nxt[266]));
Q_MX02 U4604 ( .S(n124), .A0(gcm_dek_cmd_in[202]), .A1(gcm_dek_cmd_in[266]), .Z(n1909));
Q_AN03 U4605 ( .A0(n38), .A1(n1910), .A2(n37), .Z(gcm_dek_cmd_in_nxt[265]));
Q_MX02 U4606 ( .S(n124), .A0(gcm_dek_cmd_in[201]), .A1(gcm_dek_cmd_in[265]), .Z(n1910));
Q_AN03 U4607 ( .A0(n38), .A1(n1911), .A2(n37), .Z(gcm_dek_cmd_in_nxt[264]));
Q_MX02 U4608 ( .S(n124), .A0(gcm_dek_cmd_in[200]), .A1(gcm_dek_cmd_in[264]), .Z(n1911));
Q_AN03 U4609 ( .A0(n38), .A1(n1912), .A2(n37), .Z(gcm_dek_cmd_in_nxt[263]));
Q_MX02 U4610 ( .S(n124), .A0(gcm_dek_cmd_in[199]), .A1(gcm_dek_cmd_in[263]), .Z(n1912));
Q_AN03 U4611 ( .A0(n38), .A1(n1913), .A2(n37), .Z(gcm_dek_cmd_in_nxt[262]));
Q_MX02 U4612 ( .S(n124), .A0(gcm_dek_cmd_in[198]), .A1(gcm_dek_cmd_in[262]), .Z(n1913));
Q_AN03 U4613 ( .A0(n38), .A1(n1914), .A2(n37), .Z(gcm_dek_cmd_in_nxt[261]));
Q_MX02 U4614 ( .S(n124), .A0(gcm_dek_cmd_in[197]), .A1(gcm_dek_cmd_in[261]), .Z(n1914));
Q_AN03 U4615 ( .A0(n38), .A1(n1915), .A2(n37), .Z(gcm_dek_cmd_in_nxt[260]));
Q_MX02 U4616 ( .S(n124), .A0(gcm_dek_cmd_in[196]), .A1(gcm_dek_cmd_in[260]), .Z(n1915));
Q_AN03 U4617 ( .A0(n38), .A1(n1916), .A2(n37), .Z(gcm_dek_cmd_in_nxt[259]));
Q_MX02 U4618 ( .S(n124), .A0(gcm_dek_cmd_in[195]), .A1(gcm_dek_cmd_in[259]), .Z(n1916));
Q_AN03 U4619 ( .A0(n38), .A1(n1917), .A2(n37), .Z(gcm_dek_cmd_in_nxt[258]));
Q_MX02 U4620 ( .S(n124), .A0(gcm_dek_cmd_in[194]), .A1(gcm_dek_cmd_in[258]), .Z(n1917));
Q_AN03 U4621 ( .A0(n38), .A1(n1918), .A2(n37), .Z(gcm_dek_cmd_in_nxt[257]));
Q_MX02 U4622 ( .S(n124), .A0(gcm_dek_cmd_in[193]), .A1(gcm_dek_cmd_in[257]), .Z(n1918));
Q_AN03 U4623 ( .A0(n38), .A1(n1919), .A2(n37), .Z(gcm_dek_cmd_in_nxt[256]));
Q_MX02 U4624 ( .S(n124), .A0(gcm_dek_cmd_in[192]), .A1(gcm_dek_cmd_in[256]), .Z(n1919));
Q_AN03 U4625 ( .A0(n38), .A1(n1920), .A2(n37), .Z(gcm_dek_cmd_in_nxt[255]));
Q_MX02 U4626 ( .S(n124), .A0(gcm_dek_cmd_in[191]), .A1(gcm_dek_cmd_in[255]), .Z(n1920));
Q_AN03 U4627 ( .A0(n38), .A1(n1921), .A2(n37), .Z(gcm_dek_cmd_in_nxt[254]));
Q_MX02 U4628 ( .S(n124), .A0(gcm_dek_cmd_in[190]), .A1(gcm_dek_cmd_in[254]), .Z(n1921));
Q_AN03 U4629 ( .A0(n38), .A1(n1922), .A2(n37), .Z(gcm_dek_cmd_in_nxt[253]));
Q_MX02 U4630 ( .S(n124), .A0(gcm_dek_cmd_in[189]), .A1(gcm_dek_cmd_in[253]), .Z(n1922));
Q_AN03 U4631 ( .A0(n38), .A1(n1923), .A2(n37), .Z(gcm_dek_cmd_in_nxt[252]));
Q_MX02 U4632 ( .S(n124), .A0(gcm_dek_cmd_in[188]), .A1(gcm_dek_cmd_in[252]), .Z(n1923));
Q_AN03 U4633 ( .A0(n38), .A1(n1924), .A2(n37), .Z(gcm_dek_cmd_in_nxt[251]));
Q_MX02 U4634 ( .S(n124), .A0(gcm_dek_cmd_in[187]), .A1(gcm_dek_cmd_in[251]), .Z(n1924));
Q_AN03 U4635 ( .A0(n38), .A1(n1925), .A2(n37), .Z(gcm_dek_cmd_in_nxt[250]));
Q_MX02 U4636 ( .S(n124), .A0(gcm_dek_cmd_in[186]), .A1(gcm_dek_cmd_in[250]), .Z(n1925));
Q_AN03 U4637 ( .A0(n38), .A1(n1926), .A2(n37), .Z(gcm_dek_cmd_in_nxt[249]));
Q_MX02 U4638 ( .S(n124), .A0(gcm_dek_cmd_in[185]), .A1(gcm_dek_cmd_in[249]), .Z(n1926));
Q_AN03 U4639 ( .A0(n38), .A1(n1927), .A2(n37), .Z(gcm_dek_cmd_in_nxt[248]));
Q_MX02 U4640 ( .S(n124), .A0(gcm_dek_cmd_in[184]), .A1(gcm_dek_cmd_in[248]), .Z(n1927));
Q_AN03 U4641 ( .A0(n38), .A1(n1928), .A2(n37), .Z(gcm_dek_cmd_in_nxt[247]));
Q_MX02 U4642 ( .S(n124), .A0(gcm_dek_cmd_in[183]), .A1(gcm_dek_cmd_in[247]), .Z(n1928));
Q_AN03 U4643 ( .A0(n38), .A1(n1929), .A2(n37), .Z(gcm_dek_cmd_in_nxt[246]));
Q_MX02 U4644 ( .S(n124), .A0(gcm_dek_cmd_in[182]), .A1(gcm_dek_cmd_in[246]), .Z(n1929));
Q_AN03 U4645 ( .A0(n38), .A1(n1930), .A2(n37), .Z(gcm_dek_cmd_in_nxt[245]));
Q_MX02 U4646 ( .S(n124), .A0(gcm_dek_cmd_in[181]), .A1(gcm_dek_cmd_in[245]), .Z(n1930));
Q_AN03 U4647 ( .A0(n38), .A1(n1931), .A2(n37), .Z(gcm_dek_cmd_in_nxt[244]));
Q_MX02 U4648 ( .S(n124), .A0(gcm_dek_cmd_in[180]), .A1(gcm_dek_cmd_in[244]), .Z(n1931));
Q_AN03 U4649 ( .A0(n38), .A1(n1932), .A2(n37), .Z(gcm_dek_cmd_in_nxt[243]));
Q_MX02 U4650 ( .S(n124), .A0(gcm_dek_cmd_in[179]), .A1(gcm_dek_cmd_in[243]), .Z(n1932));
Q_AN03 U4651 ( .A0(n38), .A1(n1933), .A2(n37), .Z(gcm_dek_cmd_in_nxt[242]));
Q_MX02 U4652 ( .S(n124), .A0(gcm_dek_cmd_in[178]), .A1(gcm_dek_cmd_in[242]), .Z(n1933));
Q_AN03 U4653 ( .A0(n38), .A1(n1934), .A2(n37), .Z(gcm_dek_cmd_in_nxt[241]));
Q_MX02 U4654 ( .S(n124), .A0(gcm_dek_cmd_in[177]), .A1(gcm_dek_cmd_in[241]), .Z(n1934));
Q_AN03 U4655 ( .A0(n38), .A1(n1935), .A2(n37), .Z(gcm_dek_cmd_in_nxt[240]));
Q_MX02 U4656 ( .S(n124), .A0(gcm_dek_cmd_in[176]), .A1(gcm_dek_cmd_in[240]), .Z(n1935));
Q_AN03 U4657 ( .A0(n38), .A1(n1936), .A2(n37), .Z(gcm_dek_cmd_in_nxt[239]));
Q_MX02 U4658 ( .S(n124), .A0(gcm_dek_cmd_in[175]), .A1(gcm_dek_cmd_in[239]), .Z(n1936));
Q_AN03 U4659 ( .A0(n38), .A1(n1937), .A2(n37), .Z(gcm_dek_cmd_in_nxt[238]));
Q_MX02 U4660 ( .S(n124), .A0(gcm_dek_cmd_in[174]), .A1(gcm_dek_cmd_in[238]), .Z(n1937));
Q_AN03 U4661 ( .A0(n38), .A1(n1938), .A2(n37), .Z(gcm_dek_cmd_in_nxt[237]));
Q_MX02 U4662 ( .S(n124), .A0(gcm_dek_cmd_in[173]), .A1(gcm_dek_cmd_in[237]), .Z(n1938));
Q_AN03 U4663 ( .A0(n38), .A1(n1939), .A2(n37), .Z(gcm_dek_cmd_in_nxt[236]));
Q_MX02 U4664 ( .S(n124), .A0(gcm_dek_cmd_in[172]), .A1(gcm_dek_cmd_in[236]), .Z(n1939));
Q_AN03 U4665 ( .A0(n38), .A1(n1940), .A2(n37), .Z(gcm_dek_cmd_in_nxt[235]));
Q_MX02 U4666 ( .S(n124), .A0(gcm_dek_cmd_in[171]), .A1(gcm_dek_cmd_in[235]), .Z(n1940));
Q_AN03 U4667 ( .A0(n38), .A1(n1941), .A2(n37), .Z(gcm_dek_cmd_in_nxt[234]));
Q_MX02 U4668 ( .S(n124), .A0(gcm_dek_cmd_in[170]), .A1(gcm_dek_cmd_in[234]), .Z(n1941));
Q_AN03 U4669 ( .A0(n38), .A1(n1942), .A2(n37), .Z(gcm_dek_cmd_in_nxt[233]));
Q_MX02 U4670 ( .S(n124), .A0(gcm_dek_cmd_in[169]), .A1(gcm_dek_cmd_in[233]), .Z(n1942));
Q_AN03 U4671 ( .A0(n38), .A1(n1943), .A2(n37), .Z(gcm_dek_cmd_in_nxt[232]));
Q_MX02 U4672 ( .S(n124), .A0(gcm_dek_cmd_in[168]), .A1(gcm_dek_cmd_in[232]), .Z(n1943));
Q_AN03 U4673 ( .A0(n38), .A1(n1944), .A2(n37), .Z(gcm_dek_cmd_in_nxt[231]));
Q_MX02 U4674 ( .S(n124), .A0(gcm_dek_cmd_in[167]), .A1(gcm_dek_cmd_in[231]), .Z(n1944));
Q_AN03 U4675 ( .A0(n38), .A1(n1945), .A2(n37), .Z(gcm_dek_cmd_in_nxt[230]));
Q_MX02 U4676 ( .S(n124), .A0(gcm_dek_cmd_in[166]), .A1(gcm_dek_cmd_in[230]), .Z(n1945));
Q_AN03 U4677 ( .A0(n38), .A1(n1946), .A2(n37), .Z(gcm_dek_cmd_in_nxt[229]));
Q_MX02 U4678 ( .S(n124), .A0(gcm_dek_cmd_in[165]), .A1(gcm_dek_cmd_in[229]), .Z(n1946));
Q_AN03 U4679 ( .A0(n38), .A1(n1947), .A2(n37), .Z(gcm_dek_cmd_in_nxt[228]));
Q_MX02 U4680 ( .S(n124), .A0(gcm_dek_cmd_in[164]), .A1(gcm_dek_cmd_in[228]), .Z(n1947));
Q_AN03 U4681 ( .A0(n38), .A1(n1948), .A2(n37), .Z(gcm_dek_cmd_in_nxt[227]));
Q_MX02 U4682 ( .S(n124), .A0(gcm_dek_cmd_in[163]), .A1(gcm_dek_cmd_in[227]), .Z(n1948));
Q_AN03 U4683 ( .A0(n38), .A1(n1949), .A2(n37), .Z(gcm_dek_cmd_in_nxt[226]));
Q_MX02 U4684 ( .S(n124), .A0(gcm_dek_cmd_in[162]), .A1(gcm_dek_cmd_in[226]), .Z(n1949));
Q_AN03 U4685 ( .A0(n38), .A1(n1950), .A2(n37), .Z(gcm_dek_cmd_in_nxt[225]));
Q_MX02 U4686 ( .S(n124), .A0(gcm_dek_cmd_in[161]), .A1(gcm_dek_cmd_in[225]), .Z(n1950));
Q_AN03 U4687 ( .A0(n38), .A1(n1951), .A2(n37), .Z(gcm_dek_cmd_in_nxt[224]));
Q_MX02 U4688 ( .S(n124), .A0(gcm_dek_cmd_in[160]), .A1(gcm_dek_cmd_in[224]), .Z(n1951));
Q_AN03 U4689 ( .A0(n38), .A1(n1952), .A2(n37), .Z(gcm_dek_cmd_in_nxt[223]));
Q_MX02 U4690 ( .S(n124), .A0(gcm_dek_cmd_in[159]), .A1(gcm_dek_cmd_in[223]), .Z(n1952));
Q_AN03 U4691 ( .A0(n38), .A1(n1953), .A2(n37), .Z(gcm_dek_cmd_in_nxt[222]));
Q_MX02 U4692 ( .S(n124), .A0(gcm_dek_cmd_in[158]), .A1(gcm_dek_cmd_in[222]), .Z(n1953));
Q_AN03 U4693 ( .A0(n38), .A1(n1954), .A2(n37), .Z(gcm_dek_cmd_in_nxt[221]));
Q_MX02 U4694 ( .S(n124), .A0(gcm_dek_cmd_in[157]), .A1(gcm_dek_cmd_in[221]), .Z(n1954));
Q_AN03 U4695 ( .A0(n38), .A1(n1955), .A2(n37), .Z(gcm_dek_cmd_in_nxt[220]));
Q_MX02 U4696 ( .S(n124), .A0(gcm_dek_cmd_in[156]), .A1(gcm_dek_cmd_in[220]), .Z(n1955));
Q_AN03 U4697 ( .A0(n38), .A1(n1956), .A2(n37), .Z(gcm_dek_cmd_in_nxt[219]));
Q_MX02 U4698 ( .S(n124), .A0(gcm_dek_cmd_in[155]), .A1(gcm_dek_cmd_in[219]), .Z(n1956));
Q_AN03 U4699 ( .A0(n38), .A1(n1957), .A2(n37), .Z(gcm_dek_cmd_in_nxt[218]));
Q_MX02 U4700 ( .S(n124), .A0(gcm_dek_cmd_in[154]), .A1(gcm_dek_cmd_in[218]), .Z(n1957));
Q_AN03 U4701 ( .A0(n38), .A1(n1958), .A2(n37), .Z(gcm_dek_cmd_in_nxt[217]));
Q_MX02 U4702 ( .S(n124), .A0(gcm_dek_cmd_in[153]), .A1(gcm_dek_cmd_in[217]), .Z(n1958));
Q_AN03 U4703 ( .A0(n38), .A1(n1959), .A2(n37), .Z(gcm_dek_cmd_in_nxt[216]));
Q_MX02 U4704 ( .S(n124), .A0(gcm_dek_cmd_in[152]), .A1(gcm_dek_cmd_in[216]), .Z(n1959));
Q_AN03 U4705 ( .A0(n38), .A1(n1960), .A2(n37), .Z(gcm_dek_cmd_in_nxt[215]));
Q_MX02 U4706 ( .S(n124), .A0(gcm_dek_cmd_in[151]), .A1(gcm_dek_cmd_in[215]), .Z(n1960));
Q_AN03 U4707 ( .A0(n38), .A1(n1961), .A2(n37), .Z(gcm_dek_cmd_in_nxt[214]));
Q_MX02 U4708 ( .S(n124), .A0(gcm_dek_cmd_in[150]), .A1(gcm_dek_cmd_in[214]), .Z(n1961));
Q_AN03 U4709 ( .A0(n38), .A1(n1962), .A2(n37), .Z(gcm_dek_cmd_in_nxt[213]));
Q_MX02 U4710 ( .S(n124), .A0(gcm_dek_cmd_in[149]), .A1(gcm_dek_cmd_in[213]), .Z(n1962));
Q_AN03 U4711 ( .A0(n38), .A1(n1963), .A2(n37), .Z(gcm_dek_cmd_in_nxt[212]));
Q_MX02 U4712 ( .S(n124), .A0(gcm_dek_cmd_in[148]), .A1(gcm_dek_cmd_in[212]), .Z(n1963));
Q_AN03 U4713 ( .A0(n38), .A1(n1964), .A2(n37), .Z(gcm_dek_cmd_in_nxt[211]));
Q_MX02 U4714 ( .S(n124), .A0(gcm_dek_cmd_in[147]), .A1(gcm_dek_cmd_in[211]), .Z(n1964));
Q_AN03 U4715 ( .A0(n38), .A1(n1965), .A2(n37), .Z(gcm_dek_cmd_in_nxt[210]));
Q_MX02 U4716 ( .S(n124), .A0(gcm_dek_cmd_in[146]), .A1(gcm_dek_cmd_in[210]), .Z(n1965));
Q_AN03 U4717 ( .A0(n38), .A1(n1966), .A2(n37), .Z(gcm_dek_cmd_in_nxt[209]));
Q_MX02 U4718 ( .S(n124), .A0(gcm_dek_cmd_in[145]), .A1(gcm_dek_cmd_in[209]), .Z(n1966));
Q_AN03 U4719 ( .A0(n38), .A1(n1967), .A2(n37), .Z(gcm_dek_cmd_in_nxt[208]));
Q_MX02 U4720 ( .S(n124), .A0(gcm_dek_cmd_in[144]), .A1(gcm_dek_cmd_in[208]), .Z(n1967));
Q_AN03 U4721 ( .A0(n38), .A1(n1968), .A2(n37), .Z(gcm_dek_cmd_in_nxt[207]));
Q_MX02 U4722 ( .S(n124), .A0(gcm_dek_cmd_in[143]), .A1(gcm_dek_cmd_in[207]), .Z(n1968));
Q_AN03 U4723 ( .A0(n38), .A1(n1969), .A2(n37), .Z(gcm_dek_cmd_in_nxt[206]));
Q_MX02 U4724 ( .S(n124), .A0(gcm_dek_cmd_in[142]), .A1(gcm_dek_cmd_in[206]), .Z(n1969));
Q_AN03 U4725 ( .A0(n38), .A1(n1970), .A2(n37), .Z(gcm_dek_cmd_in_nxt[205]));
Q_MX02 U4726 ( .S(n124), .A0(gcm_dek_cmd_in[141]), .A1(gcm_dek_cmd_in[205]), .Z(n1970));
Q_AN03 U4727 ( .A0(n38), .A1(n1971), .A2(n37), .Z(gcm_dek_cmd_in_nxt[204]));
Q_MX02 U4728 ( .S(n124), .A0(gcm_dek_cmd_in[140]), .A1(gcm_dek_cmd_in[204]), .Z(n1971));
Q_AN03 U4729 ( .A0(n38), .A1(n1972), .A2(n37), .Z(gcm_dek_cmd_in_nxt[203]));
Q_MX02 U4730 ( .S(n124), .A0(gcm_dek_cmd_in[139]), .A1(gcm_dek_cmd_in[203]), .Z(n1972));
Q_AN03 U4731 ( .A0(n38), .A1(n1973), .A2(n37), .Z(gcm_dek_cmd_in_nxt[202]));
Q_MX02 U4732 ( .S(n124), .A0(gcm_dek_cmd_in[138]), .A1(gcm_dek_cmd_in[202]), .Z(n1973));
Q_AN03 U4733 ( .A0(n38), .A1(n1974), .A2(n37), .Z(gcm_dek_cmd_in_nxt[201]));
Q_MX02 U4734 ( .S(n124), .A0(gcm_dek_cmd_in[137]), .A1(gcm_dek_cmd_in[201]), .Z(n1974));
Q_AN03 U4735 ( .A0(n38), .A1(n1975), .A2(n37), .Z(gcm_dek_cmd_in_nxt[200]));
Q_MX02 U4736 ( .S(n124), .A0(gcm_dek_cmd_in[136]), .A1(gcm_dek_cmd_in[200]), .Z(n1975));
Q_AN03 U4737 ( .A0(n38), .A1(n1976), .A2(n37), .Z(gcm_dek_cmd_in_nxt[199]));
Q_MX02 U4738 ( .S(n124), .A0(gcm_dek_cmd_in[135]), .A1(gcm_dek_cmd_in[199]), .Z(n1976));
Q_AN03 U4739 ( .A0(n38), .A1(n1977), .A2(n37), .Z(gcm_dek_cmd_in_nxt[198]));
Q_MX02 U4740 ( .S(n124), .A0(gcm_dek_cmd_in[134]), .A1(gcm_dek_cmd_in[198]), .Z(n1977));
Q_AN03 U4741 ( .A0(n38), .A1(n1978), .A2(n37), .Z(gcm_dek_cmd_in_nxt[197]));
Q_MX02 U4742 ( .S(n124), .A0(gcm_dek_cmd_in[133]), .A1(gcm_dek_cmd_in[197]), .Z(n1978));
Q_AN03 U4743 ( .A0(n38), .A1(n1979), .A2(n37), .Z(gcm_dek_cmd_in_nxt[196]));
Q_MX02 U4744 ( .S(n124), .A0(gcm_dek_cmd_in[132]), .A1(gcm_dek_cmd_in[196]), .Z(n1979));
Q_AN03 U4745 ( .A0(n38), .A1(n1980), .A2(n37), .Z(gcm_dek_cmd_in_nxt[195]));
Q_MX02 U4746 ( .S(n124), .A0(gcm_dek_cmd_in[131]), .A1(gcm_dek_cmd_in[195]), .Z(n1980));
Q_AN03 U4747 ( .A0(n38), .A1(n1981), .A2(n37), .Z(gcm_dek_cmd_in_nxt[194]));
Q_MX02 U4748 ( .S(n124), .A0(gcm_dek_cmd_in[130]), .A1(gcm_dek_cmd_in[194]), .Z(n1981));
Q_AN03 U4749 ( .A0(n38), .A1(n1982), .A2(n37), .Z(gcm_dek_cmd_in_nxt[193]));
Q_MX02 U4750 ( .S(n124), .A0(gcm_dek_cmd_in[129]), .A1(gcm_dek_cmd_in[193]), .Z(n1982));
Q_AN03 U4751 ( .A0(n38), .A1(n1983), .A2(n37), .Z(gcm_dek_cmd_in_nxt[192]));
Q_MX02 U4752 ( .S(n124), .A0(gcm_dek_cmd_in[128]), .A1(gcm_dek_cmd_in[192]), .Z(n1983));
Q_AN03 U4753 ( .A0(n38), .A1(n1984), .A2(n37), .Z(gcm_dek_cmd_in_nxt[191]));
Q_MX02 U4754 ( .S(n124), .A0(gcm_dek_cmd_in[127]), .A1(gcm_dek_cmd_in[191]), .Z(n1984));
Q_AN03 U4755 ( .A0(n38), .A1(n1985), .A2(n37), .Z(gcm_dek_cmd_in_nxt[190]));
Q_MX02 U4756 ( .S(n124), .A0(gcm_dek_cmd_in[126]), .A1(gcm_dek_cmd_in[190]), .Z(n1985));
Q_AN03 U4757 ( .A0(n38), .A1(n1986), .A2(n37), .Z(gcm_dek_cmd_in_nxt[189]));
Q_MX02 U4758 ( .S(n124), .A0(gcm_dek_cmd_in[125]), .A1(gcm_dek_cmd_in[189]), .Z(n1986));
Q_AN03 U4759 ( .A0(n38), .A1(n1987), .A2(n37), .Z(gcm_dek_cmd_in_nxt[188]));
Q_MX02 U4760 ( .S(n124), .A0(gcm_dek_cmd_in[124]), .A1(gcm_dek_cmd_in[188]), .Z(n1987));
Q_AN03 U4761 ( .A0(n38), .A1(n1988), .A2(n37), .Z(gcm_dek_cmd_in_nxt[187]));
Q_MX02 U4762 ( .S(n124), .A0(gcm_dek_cmd_in[123]), .A1(gcm_dek_cmd_in[187]), .Z(n1988));
Q_AN03 U4763 ( .A0(n38), .A1(n1989), .A2(n37), .Z(gcm_dek_cmd_in_nxt[186]));
Q_MX02 U4764 ( .S(n124), .A0(gcm_dek_cmd_in[122]), .A1(gcm_dek_cmd_in[186]), .Z(n1989));
Q_AN03 U4765 ( .A0(n38), .A1(n1990), .A2(n37), .Z(gcm_dek_cmd_in_nxt[185]));
Q_MX02 U4766 ( .S(n124), .A0(gcm_dek_cmd_in[121]), .A1(gcm_dek_cmd_in[185]), .Z(n1990));
Q_AN03 U4767 ( .A0(n38), .A1(n1991), .A2(n37), .Z(gcm_dek_cmd_in_nxt[184]));
Q_MX02 U4768 ( .S(n124), .A0(gcm_dek_cmd_in[120]), .A1(gcm_dek_cmd_in[184]), .Z(n1991));
Q_AN03 U4769 ( .A0(n38), .A1(n1992), .A2(n37), .Z(gcm_dek_cmd_in_nxt[183]));
Q_MX02 U4770 ( .S(n124), .A0(gcm_dek_cmd_in[119]), .A1(gcm_dek_cmd_in[183]), .Z(n1992));
Q_AN03 U4771 ( .A0(n38), .A1(n1993), .A2(n37), .Z(gcm_dek_cmd_in_nxt[182]));
Q_MX02 U4772 ( .S(n124), .A0(gcm_dek_cmd_in[118]), .A1(gcm_dek_cmd_in[182]), .Z(n1993));
Q_AN03 U4773 ( .A0(n38), .A1(n1994), .A2(n37), .Z(gcm_dek_cmd_in_nxt[181]));
Q_MX02 U4774 ( .S(n124), .A0(gcm_dek_cmd_in[117]), .A1(gcm_dek_cmd_in[181]), .Z(n1994));
Q_AN03 U4775 ( .A0(n38), .A1(n1995), .A2(n37), .Z(gcm_dek_cmd_in_nxt[180]));
Q_MX02 U4776 ( .S(n124), .A0(gcm_dek_cmd_in[116]), .A1(gcm_dek_cmd_in[180]), .Z(n1995));
Q_AN03 U4777 ( .A0(n38), .A1(n1996), .A2(n37), .Z(gcm_dek_cmd_in_nxt[179]));
Q_MX02 U4778 ( .S(n124), .A0(gcm_dek_cmd_in[115]), .A1(gcm_dek_cmd_in[179]), .Z(n1996));
Q_AN03 U4779 ( .A0(n38), .A1(n1997), .A2(n37), .Z(gcm_dek_cmd_in_nxt[178]));
Q_MX02 U4780 ( .S(n124), .A0(gcm_dek_cmd_in[114]), .A1(gcm_dek_cmd_in[178]), .Z(n1997));
Q_AN03 U4781 ( .A0(n38), .A1(n1998), .A2(n37), .Z(gcm_dek_cmd_in_nxt[177]));
Q_MX02 U4782 ( .S(n124), .A0(gcm_dek_cmd_in[113]), .A1(gcm_dek_cmd_in[177]), .Z(n1998));
Q_AN03 U4783 ( .A0(n38), .A1(n1999), .A2(n37), .Z(gcm_dek_cmd_in_nxt[176]));
Q_MX02 U4784 ( .S(n124), .A0(gcm_dek_cmd_in[112]), .A1(gcm_dek_cmd_in[176]), .Z(n1999));
Q_AN03 U4785 ( .A0(n38), .A1(n2000), .A2(n37), .Z(gcm_dek_cmd_in_nxt[175]));
Q_MX02 U4786 ( .S(n124), .A0(gcm_dek_cmd_in[111]), .A1(gcm_dek_cmd_in[175]), .Z(n2000));
Q_AN03 U4787 ( .A0(n38), .A1(n2001), .A2(n37), .Z(gcm_dek_cmd_in_nxt[174]));
Q_MX02 U4788 ( .S(n124), .A0(gcm_dek_cmd_in[110]), .A1(gcm_dek_cmd_in[174]), .Z(n2001));
Q_AN03 U4789 ( .A0(n38), .A1(n2002), .A2(n37), .Z(gcm_dek_cmd_in_nxt[173]));
Q_MX02 U4790 ( .S(n124), .A0(gcm_dek_cmd_in[109]), .A1(gcm_dek_cmd_in[173]), .Z(n2002));
Q_AN03 U4791 ( .A0(n38), .A1(n2003), .A2(n37), .Z(gcm_dek_cmd_in_nxt[172]));
Q_MX02 U4792 ( .S(n124), .A0(gcm_dek_cmd_in[108]), .A1(gcm_dek_cmd_in[172]), .Z(n2003));
Q_AN03 U4793 ( .A0(n38), .A1(n2004), .A2(n37), .Z(gcm_dek_cmd_in_nxt[171]));
Q_MX02 U4794 ( .S(n124), .A0(gcm_dek_cmd_in[107]), .A1(gcm_dek_cmd_in[171]), .Z(n2004));
Q_AN03 U4795 ( .A0(n38), .A1(n2005), .A2(n37), .Z(gcm_dek_cmd_in_nxt[170]));
Q_MX02 U4796 ( .S(n124), .A0(gcm_dek_cmd_in[106]), .A1(gcm_dek_cmd_in[170]), .Z(n2005));
Q_AN03 U4797 ( .A0(n38), .A1(n2006), .A2(n37), .Z(gcm_dek_cmd_in_nxt[169]));
Q_MX02 U4798 ( .S(n124), .A0(gcm_dek_cmd_in[105]), .A1(gcm_dek_cmd_in[169]), .Z(n2006));
Q_AN03 U4799 ( .A0(n38), .A1(n2007), .A2(n37), .Z(gcm_dek_cmd_in_nxt[168]));
Q_MX02 U4800 ( .S(n124), .A0(gcm_dek_cmd_in[104]), .A1(gcm_dek_cmd_in[168]), .Z(n2007));
Q_AN03 U4801 ( .A0(n38), .A1(n2008), .A2(n37), .Z(gcm_dek_cmd_in_nxt[167]));
Q_MX02 U4802 ( .S(n124), .A0(gcm_dek_cmd_in[103]), .A1(gcm_dek_cmd_in[167]), .Z(n2008));
Q_AN03 U4803 ( .A0(n38), .A1(n2009), .A2(n37), .Z(gcm_dek_cmd_in_nxt[166]));
Q_MX02 U4804 ( .S(n124), .A0(gcm_dek_cmd_in[102]), .A1(gcm_dek_cmd_in[166]), .Z(n2009));
Q_AN03 U4805 ( .A0(n38), .A1(n2010), .A2(n37), .Z(gcm_dek_cmd_in_nxt[165]));
Q_MX02 U4806 ( .S(n124), .A0(gcm_dek_cmd_in[101]), .A1(gcm_dek_cmd_in[165]), .Z(n2010));
Q_AN03 U4807 ( .A0(n38), .A1(n2011), .A2(n37), .Z(gcm_dek_cmd_in_nxt[164]));
Q_MX02 U4808 ( .S(n124), .A0(gcm_dek_cmd_in[100]), .A1(gcm_dek_cmd_in[164]), .Z(n2011));
Q_AN03 U4809 ( .A0(n38), .A1(n2012), .A2(n37), .Z(gcm_dek_cmd_in_nxt[163]));
Q_MX02 U4810 ( .S(n124), .A0(gcm_dek_cmd_in[99]), .A1(gcm_dek_cmd_in[163]), .Z(n2012));
Q_AN03 U4811 ( .A0(n38), .A1(n2013), .A2(n37), .Z(gcm_dek_cmd_in_nxt[162]));
Q_MX02 U4812 ( .S(n124), .A0(kme_internal_out[63]), .A1(gcm_dek_cmd_in[162]), .Z(n2013));
Q_AN03 U4813 ( .A0(n38), .A1(n2014), .A2(n37), .Z(gcm_dek_cmd_in_nxt[161]));
Q_MX02 U4814 ( .S(n124), .A0(kme_internal_out[62]), .A1(gcm_dek_cmd_in[161]), .Z(n2014));
Q_AN03 U4815 ( .A0(n38), .A1(n2015), .A2(n37), .Z(gcm_dek_cmd_in_nxt[160]));
Q_MX02 U4816 ( .S(n124), .A0(kme_internal_out[61]), .A1(gcm_dek_cmd_in[160]), .Z(n2015));
Q_AN03 U4817 ( .A0(n38), .A1(n2016), .A2(n37), .Z(gcm_dek_cmd_in_nxt[159]));
Q_MX02 U4818 ( .S(n124), .A0(kme_internal_out[60]), .A1(gcm_dek_cmd_in[159]), .Z(n2016));
Q_AN03 U4819 ( .A0(n38), .A1(n2017), .A2(n37), .Z(gcm_dek_cmd_in_nxt[158]));
Q_MX02 U4820 ( .S(n124), .A0(kme_internal_out[59]), .A1(gcm_dek_cmd_in[158]), .Z(n2017));
Q_AN03 U4821 ( .A0(n38), .A1(n2018), .A2(n37), .Z(gcm_dek_cmd_in_nxt[157]));
Q_MX02 U4822 ( .S(n124), .A0(kme_internal_out[58]), .A1(gcm_dek_cmd_in[157]), .Z(n2018));
Q_AN03 U4823 ( .A0(n38), .A1(n2019), .A2(n37), .Z(gcm_dek_cmd_in_nxt[156]));
Q_MX02 U4824 ( .S(n124), .A0(kme_internal_out[57]), .A1(gcm_dek_cmd_in[156]), .Z(n2019));
Q_AN03 U4825 ( .A0(n38), .A1(n2020), .A2(n37), .Z(gcm_dek_cmd_in_nxt[155]));
Q_MX02 U4826 ( .S(n124), .A0(kme_internal_out[56]), .A1(gcm_dek_cmd_in[155]), .Z(n2020));
Q_AN03 U4827 ( .A0(n38), .A1(n2021), .A2(n37), .Z(gcm_dek_cmd_in_nxt[154]));
Q_MX02 U4828 ( .S(n124), .A0(kme_internal_out[55]), .A1(gcm_dek_cmd_in[154]), .Z(n2021));
Q_AN03 U4829 ( .A0(n38), .A1(n2022), .A2(n37), .Z(gcm_dek_cmd_in_nxt[153]));
Q_MX02 U4830 ( .S(n124), .A0(kme_internal_out[54]), .A1(gcm_dek_cmd_in[153]), .Z(n2022));
Q_AN03 U4831 ( .A0(n38), .A1(n2023), .A2(n37), .Z(gcm_dek_cmd_in_nxt[152]));
Q_MX02 U4832 ( .S(n124), .A0(kme_internal_out[53]), .A1(gcm_dek_cmd_in[152]), .Z(n2023));
Q_AN03 U4833 ( .A0(n38), .A1(n2024), .A2(n37), .Z(gcm_dek_cmd_in_nxt[151]));
Q_MX02 U4834 ( .S(n124), .A0(kme_internal_out[52]), .A1(gcm_dek_cmd_in[151]), .Z(n2024));
Q_AN03 U4835 ( .A0(n38), .A1(n2025), .A2(n37), .Z(gcm_dek_cmd_in_nxt[150]));
Q_MX02 U4836 ( .S(n124), .A0(kme_internal_out[51]), .A1(gcm_dek_cmd_in[150]), .Z(n2025));
Q_AN03 U4837 ( .A0(n38), .A1(n2026), .A2(n37), .Z(gcm_dek_cmd_in_nxt[149]));
Q_MX02 U4838 ( .S(n124), .A0(kme_internal_out[50]), .A1(gcm_dek_cmd_in[149]), .Z(n2026));
Q_AN03 U4839 ( .A0(n38), .A1(n2027), .A2(n37), .Z(gcm_dek_cmd_in_nxt[148]));
Q_MX02 U4840 ( .S(n124), .A0(kme_internal_out[49]), .A1(gcm_dek_cmd_in[148]), .Z(n2027));
Q_AN03 U4841 ( .A0(n38), .A1(n2028), .A2(n37), .Z(gcm_dek_cmd_in_nxt[147]));
Q_MX02 U4842 ( .S(n124), .A0(kme_internal_out[48]), .A1(gcm_dek_cmd_in[147]), .Z(n2028));
Q_AN03 U4843 ( .A0(n38), .A1(n2029), .A2(n37), .Z(gcm_dek_cmd_in_nxt[146]));
Q_MX02 U4844 ( .S(n124), .A0(kme_internal_out[47]), .A1(gcm_dek_cmd_in[146]), .Z(n2029));
Q_AN03 U4845 ( .A0(n38), .A1(n2030), .A2(n37), .Z(gcm_dek_cmd_in_nxt[145]));
Q_MX02 U4846 ( .S(n124), .A0(kme_internal_out[46]), .A1(gcm_dek_cmd_in[145]), .Z(n2030));
Q_AN03 U4847 ( .A0(n38), .A1(n2031), .A2(n37), .Z(gcm_dek_cmd_in_nxt[144]));
Q_MX02 U4848 ( .S(n124), .A0(kme_internal_out[45]), .A1(gcm_dek_cmd_in[144]), .Z(n2031));
Q_AN03 U4849 ( .A0(n38), .A1(n2032), .A2(n37), .Z(gcm_dek_cmd_in_nxt[143]));
Q_MX02 U4850 ( .S(n124), .A0(kme_internal_out[44]), .A1(gcm_dek_cmd_in[143]), .Z(n2032));
Q_AN03 U4851 ( .A0(n38), .A1(n2033), .A2(n37), .Z(gcm_dek_cmd_in_nxt[142]));
Q_MX02 U4852 ( .S(n124), .A0(kme_internal_out[43]), .A1(gcm_dek_cmd_in[142]), .Z(n2033));
Q_AN03 U4853 ( .A0(n38), .A1(n2034), .A2(n37), .Z(gcm_dek_cmd_in_nxt[141]));
Q_MX02 U4854 ( .S(n124), .A0(kme_internal_out[42]), .A1(gcm_dek_cmd_in[141]), .Z(n2034));
Q_AN03 U4855 ( .A0(n38), .A1(n2035), .A2(n37), .Z(gcm_dek_cmd_in_nxt[140]));
Q_MX02 U4856 ( .S(n124), .A0(kme_internal_out[41]), .A1(gcm_dek_cmd_in[140]), .Z(n2035));
Q_AN03 U4857 ( .A0(n38), .A1(n2036), .A2(n37), .Z(gcm_dek_cmd_in_nxt[139]));
Q_MX02 U4858 ( .S(n124), .A0(kme_internal_out[40]), .A1(gcm_dek_cmd_in[139]), .Z(n2036));
Q_AN03 U4859 ( .A0(n38), .A1(n2037), .A2(n37), .Z(gcm_dek_cmd_in_nxt[138]));
Q_MX02 U4860 ( .S(n124), .A0(kme_internal_out[39]), .A1(gcm_dek_cmd_in[138]), .Z(n2037));
Q_AN03 U4861 ( .A0(n38), .A1(n2038), .A2(n37), .Z(gcm_dek_cmd_in_nxt[137]));
Q_MX02 U4862 ( .S(n124), .A0(kme_internal_out[38]), .A1(gcm_dek_cmd_in[137]), .Z(n2038));
Q_AN03 U4863 ( .A0(n38), .A1(n2039), .A2(n37), .Z(gcm_dek_cmd_in_nxt[136]));
Q_MX02 U4864 ( .S(n124), .A0(kme_internal_out[37]), .A1(gcm_dek_cmd_in[136]), .Z(n2039));
Q_AN03 U4865 ( .A0(n38), .A1(n2040), .A2(n37), .Z(gcm_dek_cmd_in_nxt[135]));
Q_MX02 U4866 ( .S(n124), .A0(kme_internal_out[36]), .A1(gcm_dek_cmd_in[135]), .Z(n2040));
Q_AN03 U4867 ( .A0(n38), .A1(n2041), .A2(n37), .Z(gcm_dek_cmd_in_nxt[134]));
Q_MX02 U4868 ( .S(n124), .A0(kme_internal_out[35]), .A1(gcm_dek_cmd_in[134]), .Z(n2041));
Q_AN03 U4869 ( .A0(n38), .A1(n2042), .A2(n37), .Z(gcm_dek_cmd_in_nxt[133]));
Q_MX02 U4870 ( .S(n124), .A0(kme_internal_out[34]), .A1(gcm_dek_cmd_in[133]), .Z(n2042));
Q_AN03 U4871 ( .A0(n38), .A1(n2043), .A2(n37), .Z(gcm_dek_cmd_in_nxt[132]));
Q_MX02 U4872 ( .S(n124), .A0(kme_internal_out[33]), .A1(gcm_dek_cmd_in[132]), .Z(n2043));
Q_AN03 U4873 ( .A0(n38), .A1(n2044), .A2(n37), .Z(gcm_dek_cmd_in_nxt[131]));
Q_MX02 U4874 ( .S(n124), .A0(kme_internal_out[32]), .A1(gcm_dek_cmd_in[131]), .Z(n2044));
Q_AN03 U4875 ( .A0(n38), .A1(n2045), .A2(n37), .Z(gcm_dek_cmd_in_nxt[130]));
Q_MX02 U4876 ( .S(n124), .A0(kme_internal_out[31]), .A1(gcm_dek_cmd_in[130]), .Z(n2045));
Q_AN03 U4877 ( .A0(n38), .A1(n2046), .A2(n37), .Z(gcm_dek_cmd_in_nxt[129]));
Q_MX02 U4878 ( .S(n124), .A0(kme_internal_out[30]), .A1(gcm_dek_cmd_in[129]), .Z(n2046));
Q_AN03 U4879 ( .A0(n38), .A1(n2047), .A2(n37), .Z(gcm_dek_cmd_in_nxt[128]));
Q_MX02 U4880 ( .S(n124), .A0(kme_internal_out[29]), .A1(gcm_dek_cmd_in[128]), .Z(n2047));
Q_AN03 U4881 ( .A0(n38), .A1(n2048), .A2(n37), .Z(gcm_dek_cmd_in_nxt[127]));
Q_MX02 U4882 ( .S(n124), .A0(kme_internal_out[28]), .A1(gcm_dek_cmd_in[127]), .Z(n2048));
Q_AN03 U4883 ( .A0(n38), .A1(n2049), .A2(n37), .Z(gcm_dek_cmd_in_nxt[126]));
Q_MX02 U4884 ( .S(n124), .A0(kme_internal_out[27]), .A1(gcm_dek_cmd_in[126]), .Z(n2049));
Q_AN03 U4885 ( .A0(n38), .A1(n2050), .A2(n37), .Z(gcm_dek_cmd_in_nxt[125]));
Q_MX02 U4886 ( .S(n124), .A0(kme_internal_out[26]), .A1(gcm_dek_cmd_in[125]), .Z(n2050));
Q_AN03 U4887 ( .A0(n38), .A1(n2051), .A2(n37), .Z(gcm_dek_cmd_in_nxt[124]));
Q_MX02 U4888 ( .S(n124), .A0(kme_internal_out[25]), .A1(gcm_dek_cmd_in[124]), .Z(n2051));
Q_AN03 U4889 ( .A0(n38), .A1(n2052), .A2(n37), .Z(gcm_dek_cmd_in_nxt[123]));
Q_MX02 U4890 ( .S(n124), .A0(kme_internal_out[24]), .A1(gcm_dek_cmd_in[123]), .Z(n2052));
Q_AN03 U4891 ( .A0(n38), .A1(n2053), .A2(n37), .Z(gcm_dek_cmd_in_nxt[122]));
Q_MX02 U4892 ( .S(n124), .A0(kme_internal_out[23]), .A1(gcm_dek_cmd_in[122]), .Z(n2053));
Q_AN03 U4893 ( .A0(n38), .A1(n2054), .A2(n37), .Z(gcm_dek_cmd_in_nxt[121]));
Q_MX02 U4894 ( .S(n124), .A0(kme_internal_out[22]), .A1(gcm_dek_cmd_in[121]), .Z(n2054));
Q_AN03 U4895 ( .A0(n38), .A1(n2055), .A2(n37), .Z(gcm_dek_cmd_in_nxt[120]));
Q_MX02 U4896 ( .S(n124), .A0(kme_internal_out[21]), .A1(gcm_dek_cmd_in[120]), .Z(n2055));
Q_AN03 U4897 ( .A0(n38), .A1(n2056), .A2(n37), .Z(gcm_dek_cmd_in_nxt[119]));
Q_MX02 U4898 ( .S(n124), .A0(kme_internal_out[20]), .A1(gcm_dek_cmd_in[119]), .Z(n2056));
Q_AN03 U4899 ( .A0(n38), .A1(n2057), .A2(n37), .Z(gcm_dek_cmd_in_nxt[118]));
Q_MX02 U4900 ( .S(n124), .A0(kme_internal_out[19]), .A1(gcm_dek_cmd_in[118]), .Z(n2057));
Q_AN03 U4901 ( .A0(n38), .A1(n2058), .A2(n37), .Z(gcm_dek_cmd_in_nxt[117]));
Q_MX02 U4902 ( .S(n124), .A0(kme_internal_out[18]), .A1(gcm_dek_cmd_in[117]), .Z(n2058));
Q_AN03 U4903 ( .A0(n38), .A1(n2059), .A2(n37), .Z(gcm_dek_cmd_in_nxt[116]));
Q_MX02 U4904 ( .S(n124), .A0(kme_internal_out[17]), .A1(gcm_dek_cmd_in[116]), .Z(n2059));
Q_AN03 U4905 ( .A0(n38), .A1(n2060), .A2(n37), .Z(gcm_dek_cmd_in_nxt[115]));
Q_MX02 U4906 ( .S(n124), .A0(kme_internal_out[16]), .A1(gcm_dek_cmd_in[115]), .Z(n2060));
Q_AN03 U4907 ( .A0(n38), .A1(n2061), .A2(n37), .Z(gcm_dek_cmd_in_nxt[114]));
Q_MX02 U4908 ( .S(n124), .A0(kme_internal_out[15]), .A1(gcm_dek_cmd_in[114]), .Z(n2061));
Q_AN03 U4909 ( .A0(n38), .A1(n2062), .A2(n37), .Z(gcm_dek_cmd_in_nxt[113]));
Q_MX02 U4910 ( .S(n124), .A0(kme_internal_out[14]), .A1(gcm_dek_cmd_in[113]), .Z(n2062));
Q_AN03 U4911 ( .A0(n38), .A1(n2063), .A2(n37), .Z(gcm_dek_cmd_in_nxt[112]));
Q_MX02 U4912 ( .S(n124), .A0(kme_internal_out[13]), .A1(gcm_dek_cmd_in[112]), .Z(n2063));
Q_AN03 U4913 ( .A0(n38), .A1(n2064), .A2(n37), .Z(gcm_dek_cmd_in_nxt[111]));
Q_MX02 U4914 ( .S(n124), .A0(kme_internal_out[12]), .A1(gcm_dek_cmd_in[111]), .Z(n2064));
Q_AN03 U4915 ( .A0(n38), .A1(n2065), .A2(n37), .Z(gcm_dek_cmd_in_nxt[110]));
Q_MX02 U4916 ( .S(n124), .A0(kme_internal_out[11]), .A1(gcm_dek_cmd_in[110]), .Z(n2065));
Q_AN03 U4917 ( .A0(n38), .A1(n2066), .A2(n37), .Z(gcm_dek_cmd_in_nxt[109]));
Q_MX02 U4918 ( .S(n124), .A0(kme_internal_out[10]), .A1(gcm_dek_cmd_in[109]), .Z(n2066));
Q_AN03 U4919 ( .A0(n38), .A1(n2067), .A2(n37), .Z(gcm_dek_cmd_in_nxt[108]));
Q_MX02 U4920 ( .S(n124), .A0(kme_internal_out[9]), .A1(gcm_dek_cmd_in[108]), .Z(n2067));
Q_AN03 U4921 ( .A0(n38), .A1(n2068), .A2(n37), .Z(gcm_dek_cmd_in_nxt[107]));
Q_MX02 U4922 ( .S(n124), .A0(kme_internal_out[8]), .A1(gcm_dek_cmd_in[107]), .Z(n2068));
Q_AN03 U4923 ( .A0(n38), .A1(n2069), .A2(n37), .Z(gcm_dek_cmd_in_nxt[106]));
Q_MX02 U4924 ( .S(n124), .A0(kme_internal_out[7]), .A1(gcm_dek_cmd_in[106]), .Z(n2069));
Q_AN03 U4925 ( .A0(n38), .A1(n2070), .A2(n37), .Z(gcm_dek_cmd_in_nxt[105]));
Q_MX02 U4926 ( .S(n124), .A0(kme_internal_out[6]), .A1(gcm_dek_cmd_in[105]), .Z(n2070));
Q_AN03 U4927 ( .A0(n38), .A1(n2071), .A2(n37), .Z(gcm_dek_cmd_in_nxt[104]));
Q_MX02 U4928 ( .S(n124), .A0(kme_internal_out[5]), .A1(gcm_dek_cmd_in[104]), .Z(n2071));
Q_AN03 U4929 ( .A0(n38), .A1(n2072), .A2(n37), .Z(gcm_dek_cmd_in_nxt[103]));
Q_MX02 U4930 ( .S(n124), .A0(kme_internal_out[4]), .A1(gcm_dek_cmd_in[103]), .Z(n2072));
Q_AN03 U4931 ( .A0(n38), .A1(n2073), .A2(n37), .Z(gcm_dek_cmd_in_nxt[102]));
Q_MX02 U4932 ( .S(n124), .A0(kme_internal_out[3]), .A1(gcm_dek_cmd_in[102]), .Z(n2073));
Q_AN03 U4933 ( .A0(n38), .A1(n2074), .A2(n37), .Z(gcm_dek_cmd_in_nxt[101]));
Q_MX02 U4934 ( .S(n124), .A0(kme_internal_out[2]), .A1(gcm_dek_cmd_in[101]), .Z(n2074));
Q_AN03 U4935 ( .A0(n38), .A1(n2075), .A2(n37), .Z(gcm_dek_cmd_in_nxt[100]));
Q_MX02 U4936 ( .S(n124), .A0(kme_internal_out[1]), .A1(gcm_dek_cmd_in[100]), .Z(n2075));
Q_AN03 U4937 ( .A0(n38), .A1(n2076), .A2(n37), .Z(gcm_dek_cmd_in_nxt[99]));
Q_MX02 U4938 ( .S(n124), .A0(kme_internal_out[0]), .A1(gcm_dek_cmd_in[99]), .Z(n2076));
Q_AN03 U4939 ( .A0(n38), .A1(n2077), .A2(n37), .Z(gcm_dek_cmd_in_nxt[610]));
Q_MX02 U4940 ( .S(n129), .A0(gcm_dek_cmd_in[546]), .A1(gcm_dek_cmd_in[610]), .Z(n2077));
Q_AN03 U4941 ( .A0(n38), .A1(n2078), .A2(n37), .Z(gcm_dek_cmd_in_nxt[609]));
Q_MX02 U4942 ( .S(n129), .A0(gcm_dek_cmd_in[545]), .A1(gcm_dek_cmd_in[609]), .Z(n2078));
Q_AN03 U4943 ( .A0(n38), .A1(n2079), .A2(n37), .Z(gcm_dek_cmd_in_nxt[608]));
Q_MX02 U4944 ( .S(n129), .A0(gcm_dek_cmd_in[544]), .A1(gcm_dek_cmd_in[608]), .Z(n2079));
Q_AN03 U4945 ( .A0(n38), .A1(n2080), .A2(n37), .Z(gcm_dek_cmd_in_nxt[607]));
Q_MX02 U4946 ( .S(n129), .A0(gcm_dek_cmd_in[543]), .A1(gcm_dek_cmd_in[607]), .Z(n2080));
Q_AN03 U4947 ( .A0(n38), .A1(n2081), .A2(n37), .Z(gcm_dek_cmd_in_nxt[606]));
Q_MX02 U4948 ( .S(n129), .A0(gcm_dek_cmd_in[542]), .A1(gcm_dek_cmd_in[606]), .Z(n2081));
Q_AN03 U4949 ( .A0(n38), .A1(n2082), .A2(n37), .Z(gcm_dek_cmd_in_nxt[605]));
Q_MX02 U4950 ( .S(n129), .A0(gcm_dek_cmd_in[541]), .A1(gcm_dek_cmd_in[605]), .Z(n2082));
Q_AN03 U4951 ( .A0(n38), .A1(n2083), .A2(n37), .Z(gcm_dek_cmd_in_nxt[604]));
Q_MX02 U4952 ( .S(n129), .A0(gcm_dek_cmd_in[540]), .A1(gcm_dek_cmd_in[604]), .Z(n2083));
Q_AN03 U4953 ( .A0(n38), .A1(n2084), .A2(n37), .Z(gcm_dek_cmd_in_nxt[603]));
Q_MX02 U4954 ( .S(n129), .A0(gcm_dek_cmd_in[539]), .A1(gcm_dek_cmd_in[603]), .Z(n2084));
Q_AN03 U4955 ( .A0(n38), .A1(n2085), .A2(n37), .Z(gcm_dek_cmd_in_nxt[602]));
Q_MX02 U4956 ( .S(n129), .A0(gcm_dek_cmd_in[538]), .A1(gcm_dek_cmd_in[602]), .Z(n2085));
Q_AN03 U4957 ( .A0(n38), .A1(n2086), .A2(n37), .Z(gcm_dek_cmd_in_nxt[601]));
Q_MX02 U4958 ( .S(n129), .A0(gcm_dek_cmd_in[537]), .A1(gcm_dek_cmd_in[601]), .Z(n2086));
Q_AN03 U4959 ( .A0(n38), .A1(n2087), .A2(n37), .Z(gcm_dek_cmd_in_nxt[600]));
Q_MX02 U4960 ( .S(n129), .A0(gcm_dek_cmd_in[536]), .A1(gcm_dek_cmd_in[600]), .Z(n2087));
Q_AN03 U4961 ( .A0(n38), .A1(n2088), .A2(n37), .Z(gcm_dek_cmd_in_nxt[599]));
Q_MX02 U4962 ( .S(n129), .A0(gcm_dek_cmd_in[535]), .A1(gcm_dek_cmd_in[599]), .Z(n2088));
Q_AN03 U4963 ( .A0(n38), .A1(n2089), .A2(n37), .Z(gcm_dek_cmd_in_nxt[598]));
Q_MX02 U4964 ( .S(n129), .A0(gcm_dek_cmd_in[534]), .A1(gcm_dek_cmd_in[598]), .Z(n2089));
Q_AN03 U4965 ( .A0(n38), .A1(n2090), .A2(n37), .Z(gcm_dek_cmd_in_nxt[597]));
Q_MX02 U4966 ( .S(n129), .A0(gcm_dek_cmd_in[533]), .A1(gcm_dek_cmd_in[597]), .Z(n2090));
Q_AN03 U4967 ( .A0(n38), .A1(n2091), .A2(n37), .Z(gcm_dek_cmd_in_nxt[596]));
Q_MX02 U4968 ( .S(n129), .A0(gcm_dek_cmd_in[532]), .A1(gcm_dek_cmd_in[596]), .Z(n2091));
Q_AN03 U4969 ( .A0(n38), .A1(n2092), .A2(n37), .Z(gcm_dek_cmd_in_nxt[595]));
Q_MX02 U4970 ( .S(n129), .A0(gcm_dek_cmd_in[531]), .A1(gcm_dek_cmd_in[595]), .Z(n2092));
Q_AN03 U4971 ( .A0(n38), .A1(n2093), .A2(n37), .Z(gcm_dek_cmd_in_nxt[594]));
Q_MX02 U4972 ( .S(n129), .A0(gcm_dek_cmd_in[530]), .A1(gcm_dek_cmd_in[594]), .Z(n2093));
Q_AN03 U4973 ( .A0(n38), .A1(n2094), .A2(n37), .Z(gcm_dek_cmd_in_nxt[593]));
Q_MX02 U4974 ( .S(n129), .A0(gcm_dek_cmd_in[529]), .A1(gcm_dek_cmd_in[593]), .Z(n2094));
Q_AN03 U4975 ( .A0(n38), .A1(n2095), .A2(n37), .Z(gcm_dek_cmd_in_nxt[592]));
Q_MX02 U4976 ( .S(n129), .A0(gcm_dek_cmd_in[528]), .A1(gcm_dek_cmd_in[592]), .Z(n2095));
Q_AN03 U4977 ( .A0(n38), .A1(n2096), .A2(n37), .Z(gcm_dek_cmd_in_nxt[591]));
Q_MX02 U4978 ( .S(n129), .A0(gcm_dek_cmd_in[527]), .A1(gcm_dek_cmd_in[591]), .Z(n2096));
Q_AN03 U4979 ( .A0(n38), .A1(n2097), .A2(n37), .Z(gcm_dek_cmd_in_nxt[590]));
Q_MX02 U4980 ( .S(n129), .A0(gcm_dek_cmd_in[526]), .A1(gcm_dek_cmd_in[590]), .Z(n2097));
Q_AN03 U4981 ( .A0(n38), .A1(n2098), .A2(n37), .Z(gcm_dek_cmd_in_nxt[589]));
Q_MX02 U4982 ( .S(n129), .A0(gcm_dek_cmd_in[525]), .A1(gcm_dek_cmd_in[589]), .Z(n2098));
Q_AN03 U4983 ( .A0(n38), .A1(n2099), .A2(n37), .Z(gcm_dek_cmd_in_nxt[588]));
Q_MX02 U4984 ( .S(n129), .A0(gcm_dek_cmd_in[524]), .A1(gcm_dek_cmd_in[588]), .Z(n2099));
Q_AN03 U4985 ( .A0(n38), .A1(n2100), .A2(n37), .Z(gcm_dek_cmd_in_nxt[587]));
Q_MX02 U4986 ( .S(n129), .A0(gcm_dek_cmd_in[523]), .A1(gcm_dek_cmd_in[587]), .Z(n2100));
Q_AN03 U4987 ( .A0(n38), .A1(n2101), .A2(n37), .Z(gcm_dek_cmd_in_nxt[586]));
Q_MX02 U4988 ( .S(n129), .A0(gcm_dek_cmd_in[522]), .A1(gcm_dek_cmd_in[586]), .Z(n2101));
Q_AN03 U4989 ( .A0(n38), .A1(n2102), .A2(n37), .Z(gcm_dek_cmd_in_nxt[585]));
Q_MX02 U4990 ( .S(n129), .A0(gcm_dek_cmd_in[521]), .A1(gcm_dek_cmd_in[585]), .Z(n2102));
Q_AN03 U4991 ( .A0(n38), .A1(n2103), .A2(n37), .Z(gcm_dek_cmd_in_nxt[584]));
Q_MX02 U4992 ( .S(n129), .A0(gcm_dek_cmd_in[520]), .A1(gcm_dek_cmd_in[584]), .Z(n2103));
Q_AN03 U4993 ( .A0(n38), .A1(n2104), .A2(n37), .Z(gcm_dek_cmd_in_nxt[583]));
Q_MX02 U4994 ( .S(n129), .A0(gcm_dek_cmd_in[519]), .A1(gcm_dek_cmd_in[583]), .Z(n2104));
Q_AN03 U4995 ( .A0(n38), .A1(n2105), .A2(n37), .Z(gcm_dek_cmd_in_nxt[582]));
Q_MX02 U4996 ( .S(n129), .A0(gcm_dek_cmd_in[518]), .A1(gcm_dek_cmd_in[582]), .Z(n2105));
Q_AN03 U4997 ( .A0(n38), .A1(n2106), .A2(n37), .Z(gcm_dek_cmd_in_nxt[581]));
Q_MX02 U4998 ( .S(n129), .A0(gcm_dek_cmd_in[517]), .A1(gcm_dek_cmd_in[581]), .Z(n2106));
Q_AN03 U4999 ( .A0(n38), .A1(n2107), .A2(n37), .Z(gcm_dek_cmd_in_nxt[580]));
Q_MX02 U5000 ( .S(n129), .A0(gcm_dek_cmd_in[516]), .A1(gcm_dek_cmd_in[580]), .Z(n2107));
Q_AN03 U5001 ( .A0(n38), .A1(n2108), .A2(n37), .Z(gcm_dek_cmd_in_nxt[579]));
Q_MX02 U5002 ( .S(n129), .A0(gcm_dek_cmd_in[515]), .A1(gcm_dek_cmd_in[579]), .Z(n2108));
Q_AN03 U5003 ( .A0(n38), .A1(n2109), .A2(n37), .Z(gcm_dek_cmd_in_nxt[578]));
Q_MX02 U5004 ( .S(n129), .A0(gcm_dek_cmd_in[514]), .A1(gcm_dek_cmd_in[578]), .Z(n2109));
Q_AN03 U5005 ( .A0(n38), .A1(n2110), .A2(n37), .Z(gcm_dek_cmd_in_nxt[577]));
Q_MX02 U5006 ( .S(n129), .A0(gcm_dek_cmd_in[513]), .A1(gcm_dek_cmd_in[577]), .Z(n2110));
Q_AN03 U5007 ( .A0(n38), .A1(n2111), .A2(n37), .Z(gcm_dek_cmd_in_nxt[576]));
Q_MX02 U5008 ( .S(n129), .A0(gcm_dek_cmd_in[512]), .A1(gcm_dek_cmd_in[576]), .Z(n2111));
Q_AN03 U5009 ( .A0(n38), .A1(n2112), .A2(n37), .Z(gcm_dek_cmd_in_nxt[575]));
Q_MX02 U5010 ( .S(n129), .A0(gcm_dek_cmd_in[511]), .A1(gcm_dek_cmd_in[575]), .Z(n2112));
Q_AN03 U5011 ( .A0(n38), .A1(n2113), .A2(n37), .Z(gcm_dek_cmd_in_nxt[574]));
Q_MX02 U5012 ( .S(n129), .A0(gcm_dek_cmd_in[510]), .A1(gcm_dek_cmd_in[574]), .Z(n2113));
Q_AN03 U5013 ( .A0(n38), .A1(n2114), .A2(n37), .Z(gcm_dek_cmd_in_nxt[573]));
Q_MX02 U5014 ( .S(n129), .A0(gcm_dek_cmd_in[509]), .A1(gcm_dek_cmd_in[573]), .Z(n2114));
Q_AN03 U5015 ( .A0(n38), .A1(n2115), .A2(n37), .Z(gcm_dek_cmd_in_nxt[572]));
Q_MX02 U5016 ( .S(n129), .A0(gcm_dek_cmd_in[508]), .A1(gcm_dek_cmd_in[572]), .Z(n2115));
Q_AN03 U5017 ( .A0(n38), .A1(n2116), .A2(n37), .Z(gcm_dek_cmd_in_nxt[571]));
Q_MX02 U5018 ( .S(n129), .A0(gcm_dek_cmd_in[507]), .A1(gcm_dek_cmd_in[571]), .Z(n2116));
Q_AN03 U5019 ( .A0(n38), .A1(n2117), .A2(n37), .Z(gcm_dek_cmd_in_nxt[570]));
Q_MX02 U5020 ( .S(n129), .A0(gcm_dek_cmd_in[506]), .A1(gcm_dek_cmd_in[570]), .Z(n2117));
Q_AN03 U5021 ( .A0(n38), .A1(n2118), .A2(n37), .Z(gcm_dek_cmd_in_nxt[569]));
Q_MX02 U5022 ( .S(n129), .A0(gcm_dek_cmd_in[505]), .A1(gcm_dek_cmd_in[569]), .Z(n2118));
Q_AN03 U5023 ( .A0(n38), .A1(n2119), .A2(n37), .Z(gcm_dek_cmd_in_nxt[568]));
Q_MX02 U5024 ( .S(n129), .A0(gcm_dek_cmd_in[504]), .A1(gcm_dek_cmd_in[568]), .Z(n2119));
Q_AN03 U5025 ( .A0(n38), .A1(n2120), .A2(n37), .Z(gcm_dek_cmd_in_nxt[567]));
Q_MX02 U5026 ( .S(n129), .A0(gcm_dek_cmd_in[503]), .A1(gcm_dek_cmd_in[567]), .Z(n2120));
Q_AN03 U5027 ( .A0(n38), .A1(n2121), .A2(n37), .Z(gcm_dek_cmd_in_nxt[566]));
Q_MX02 U5028 ( .S(n129), .A0(gcm_dek_cmd_in[502]), .A1(gcm_dek_cmd_in[566]), .Z(n2121));
Q_AN03 U5029 ( .A0(n38), .A1(n2122), .A2(n37), .Z(gcm_dek_cmd_in_nxt[565]));
Q_MX02 U5030 ( .S(n129), .A0(gcm_dek_cmd_in[501]), .A1(gcm_dek_cmd_in[565]), .Z(n2122));
Q_AN03 U5031 ( .A0(n38), .A1(n2123), .A2(n37), .Z(gcm_dek_cmd_in_nxt[564]));
Q_MX02 U5032 ( .S(n129), .A0(gcm_dek_cmd_in[500]), .A1(gcm_dek_cmd_in[564]), .Z(n2123));
Q_AN03 U5033 ( .A0(n38), .A1(n2124), .A2(n37), .Z(gcm_dek_cmd_in_nxt[563]));
Q_MX02 U5034 ( .S(n129), .A0(gcm_dek_cmd_in[499]), .A1(gcm_dek_cmd_in[563]), .Z(n2124));
Q_AN03 U5035 ( .A0(n38), .A1(n2125), .A2(n37), .Z(gcm_dek_cmd_in_nxt[562]));
Q_MX02 U5036 ( .S(n129), .A0(gcm_dek_cmd_in[498]), .A1(gcm_dek_cmd_in[562]), .Z(n2125));
Q_AN03 U5037 ( .A0(n38), .A1(n2126), .A2(n37), .Z(gcm_dek_cmd_in_nxt[561]));
Q_MX02 U5038 ( .S(n129), .A0(gcm_dek_cmd_in[497]), .A1(gcm_dek_cmd_in[561]), .Z(n2126));
Q_AN03 U5039 ( .A0(n38), .A1(n2127), .A2(n37), .Z(gcm_dek_cmd_in_nxt[560]));
Q_MX02 U5040 ( .S(n129), .A0(gcm_dek_cmd_in[496]), .A1(gcm_dek_cmd_in[560]), .Z(n2127));
Q_AN03 U5041 ( .A0(n38), .A1(n2128), .A2(n37), .Z(gcm_dek_cmd_in_nxt[559]));
Q_MX02 U5042 ( .S(n129), .A0(gcm_dek_cmd_in[495]), .A1(gcm_dek_cmd_in[559]), .Z(n2128));
Q_AN03 U5043 ( .A0(n38), .A1(n2129), .A2(n37), .Z(gcm_dek_cmd_in_nxt[558]));
Q_MX02 U5044 ( .S(n129), .A0(gcm_dek_cmd_in[494]), .A1(gcm_dek_cmd_in[558]), .Z(n2129));
Q_AN03 U5045 ( .A0(n38), .A1(n2130), .A2(n37), .Z(gcm_dek_cmd_in_nxt[557]));
Q_MX02 U5046 ( .S(n129), .A0(gcm_dek_cmd_in[493]), .A1(gcm_dek_cmd_in[557]), .Z(n2130));
Q_AN03 U5047 ( .A0(n38), .A1(n2131), .A2(n37), .Z(gcm_dek_cmd_in_nxt[556]));
Q_MX02 U5048 ( .S(n129), .A0(gcm_dek_cmd_in[492]), .A1(gcm_dek_cmd_in[556]), .Z(n2131));
Q_AN03 U5049 ( .A0(n38), .A1(n2132), .A2(n37), .Z(gcm_dek_cmd_in_nxt[555]));
Q_MX02 U5050 ( .S(n129), .A0(gcm_dek_cmd_in[491]), .A1(gcm_dek_cmd_in[555]), .Z(n2132));
Q_AN03 U5051 ( .A0(n38), .A1(n2133), .A2(n37), .Z(gcm_dek_cmd_in_nxt[554]));
Q_MX02 U5052 ( .S(n129), .A0(gcm_dek_cmd_in[490]), .A1(gcm_dek_cmd_in[554]), .Z(n2133));
Q_AN03 U5053 ( .A0(n38), .A1(n2134), .A2(n37), .Z(gcm_dek_cmd_in_nxt[553]));
Q_MX02 U5054 ( .S(n129), .A0(gcm_dek_cmd_in[489]), .A1(gcm_dek_cmd_in[553]), .Z(n2134));
Q_AN03 U5055 ( .A0(n38), .A1(n2135), .A2(n37), .Z(gcm_dek_cmd_in_nxt[552]));
Q_MX02 U5056 ( .S(n129), .A0(gcm_dek_cmd_in[488]), .A1(gcm_dek_cmd_in[552]), .Z(n2135));
Q_AN03 U5057 ( .A0(n38), .A1(n2136), .A2(n37), .Z(gcm_dek_cmd_in_nxt[551]));
Q_MX02 U5058 ( .S(n129), .A0(gcm_dek_cmd_in[487]), .A1(gcm_dek_cmd_in[551]), .Z(n2136));
Q_AN03 U5059 ( .A0(n38), .A1(n2137), .A2(n37), .Z(gcm_dek_cmd_in_nxt[550]));
Q_MX02 U5060 ( .S(n129), .A0(gcm_dek_cmd_in[486]), .A1(gcm_dek_cmd_in[550]), .Z(n2137));
Q_AN03 U5061 ( .A0(n38), .A1(n2138), .A2(n37), .Z(gcm_dek_cmd_in_nxt[549]));
Q_MX02 U5062 ( .S(n129), .A0(gcm_dek_cmd_in[485]), .A1(gcm_dek_cmd_in[549]), .Z(n2138));
Q_AN03 U5063 ( .A0(n38), .A1(n2139), .A2(n37), .Z(gcm_dek_cmd_in_nxt[548]));
Q_MX02 U5064 ( .S(n129), .A0(gcm_dek_cmd_in[484]), .A1(gcm_dek_cmd_in[548]), .Z(n2139));
Q_AN03 U5065 ( .A0(n38), .A1(n2140), .A2(n37), .Z(gcm_dek_cmd_in_nxt[547]));
Q_MX02 U5066 ( .S(n129), .A0(gcm_dek_cmd_in[483]), .A1(gcm_dek_cmd_in[547]), .Z(n2140));
Q_AN03 U5067 ( .A0(n38), .A1(n2141), .A2(n37), .Z(gcm_dek_cmd_in_nxt[546]));
Q_MX02 U5068 ( .S(n129), .A0(gcm_dek_cmd_in[482]), .A1(gcm_dek_cmd_in[546]), .Z(n2141));
Q_AN03 U5069 ( .A0(n38), .A1(n2142), .A2(n37), .Z(gcm_dek_cmd_in_nxt[545]));
Q_MX02 U5070 ( .S(n129), .A0(gcm_dek_cmd_in[481]), .A1(gcm_dek_cmd_in[545]), .Z(n2142));
Q_AN03 U5071 ( .A0(n38), .A1(n2143), .A2(n37), .Z(gcm_dek_cmd_in_nxt[544]));
Q_MX02 U5072 ( .S(n129), .A0(gcm_dek_cmd_in[480]), .A1(gcm_dek_cmd_in[544]), .Z(n2143));
Q_AN03 U5073 ( .A0(n38), .A1(n2144), .A2(n37), .Z(gcm_dek_cmd_in_nxt[543]));
Q_MX02 U5074 ( .S(n129), .A0(gcm_dek_cmd_in[479]), .A1(gcm_dek_cmd_in[543]), .Z(n2144));
Q_AN03 U5075 ( .A0(n38), .A1(n2145), .A2(n37), .Z(gcm_dek_cmd_in_nxt[542]));
Q_MX02 U5076 ( .S(n129), .A0(gcm_dek_cmd_in[478]), .A1(gcm_dek_cmd_in[542]), .Z(n2145));
Q_AN03 U5077 ( .A0(n38), .A1(n2146), .A2(n37), .Z(gcm_dek_cmd_in_nxt[541]));
Q_MX02 U5078 ( .S(n129), .A0(gcm_dek_cmd_in[477]), .A1(gcm_dek_cmd_in[541]), .Z(n2146));
Q_AN03 U5079 ( .A0(n38), .A1(n2147), .A2(n37), .Z(gcm_dek_cmd_in_nxt[540]));
Q_MX02 U5080 ( .S(n129), .A0(gcm_dek_cmd_in[476]), .A1(gcm_dek_cmd_in[540]), .Z(n2147));
Q_AN03 U5081 ( .A0(n38), .A1(n2148), .A2(n37), .Z(gcm_dek_cmd_in_nxt[539]));
Q_MX02 U5082 ( .S(n129), .A0(gcm_dek_cmd_in[475]), .A1(gcm_dek_cmd_in[539]), .Z(n2148));
Q_AN03 U5083 ( .A0(n38), .A1(n2149), .A2(n37), .Z(gcm_dek_cmd_in_nxt[538]));
Q_MX02 U5084 ( .S(n129), .A0(gcm_dek_cmd_in[474]), .A1(gcm_dek_cmd_in[538]), .Z(n2149));
Q_AN03 U5085 ( .A0(n38), .A1(n2150), .A2(n37), .Z(gcm_dek_cmd_in_nxt[537]));
Q_MX02 U5086 ( .S(n129), .A0(gcm_dek_cmd_in[473]), .A1(gcm_dek_cmd_in[537]), .Z(n2150));
Q_AN03 U5087 ( .A0(n38), .A1(n2151), .A2(n37), .Z(gcm_dek_cmd_in_nxt[536]));
Q_MX02 U5088 ( .S(n129), .A0(gcm_dek_cmd_in[472]), .A1(gcm_dek_cmd_in[536]), .Z(n2151));
Q_AN03 U5089 ( .A0(n38), .A1(n2152), .A2(n37), .Z(gcm_dek_cmd_in_nxt[535]));
Q_MX02 U5090 ( .S(n129), .A0(gcm_dek_cmd_in[471]), .A1(gcm_dek_cmd_in[535]), .Z(n2152));
Q_AN03 U5091 ( .A0(n38), .A1(n2153), .A2(n37), .Z(gcm_dek_cmd_in_nxt[534]));
Q_MX02 U5092 ( .S(n129), .A0(gcm_dek_cmd_in[470]), .A1(gcm_dek_cmd_in[534]), .Z(n2153));
Q_AN03 U5093 ( .A0(n38), .A1(n2154), .A2(n37), .Z(gcm_dek_cmd_in_nxt[533]));
Q_MX02 U5094 ( .S(n129), .A0(gcm_dek_cmd_in[469]), .A1(gcm_dek_cmd_in[533]), .Z(n2154));
Q_AN03 U5095 ( .A0(n38), .A1(n2155), .A2(n37), .Z(gcm_dek_cmd_in_nxt[532]));
Q_MX02 U5096 ( .S(n129), .A0(gcm_dek_cmd_in[468]), .A1(gcm_dek_cmd_in[532]), .Z(n2155));
Q_AN03 U5097 ( .A0(n38), .A1(n2156), .A2(n37), .Z(gcm_dek_cmd_in_nxt[531]));
Q_MX02 U5098 ( .S(n129), .A0(gcm_dek_cmd_in[467]), .A1(gcm_dek_cmd_in[531]), .Z(n2156));
Q_AN03 U5099 ( .A0(n38), .A1(n2157), .A2(n37), .Z(gcm_dek_cmd_in_nxt[530]));
Q_MX02 U5100 ( .S(n129), .A0(gcm_dek_cmd_in[466]), .A1(gcm_dek_cmd_in[530]), .Z(n2157));
Q_AN03 U5101 ( .A0(n38), .A1(n2158), .A2(n37), .Z(gcm_dek_cmd_in_nxt[529]));
Q_MX02 U5102 ( .S(n129), .A0(gcm_dek_cmd_in[465]), .A1(gcm_dek_cmd_in[529]), .Z(n2158));
Q_AN03 U5103 ( .A0(n38), .A1(n2159), .A2(n37), .Z(gcm_dek_cmd_in_nxt[528]));
Q_MX02 U5104 ( .S(n129), .A0(gcm_dek_cmd_in[464]), .A1(gcm_dek_cmd_in[528]), .Z(n2159));
Q_AN03 U5105 ( .A0(n38), .A1(n2160), .A2(n37), .Z(gcm_dek_cmd_in_nxt[527]));
Q_MX02 U5106 ( .S(n129), .A0(gcm_dek_cmd_in[463]), .A1(gcm_dek_cmd_in[527]), .Z(n2160));
Q_AN03 U5107 ( .A0(n38), .A1(n2161), .A2(n37), .Z(gcm_dek_cmd_in_nxt[526]));
Q_MX02 U5108 ( .S(n129), .A0(gcm_dek_cmd_in[462]), .A1(gcm_dek_cmd_in[526]), .Z(n2161));
Q_AN03 U5109 ( .A0(n38), .A1(n2162), .A2(n37), .Z(gcm_dek_cmd_in_nxt[525]));
Q_MX02 U5110 ( .S(n129), .A0(gcm_dek_cmd_in[461]), .A1(gcm_dek_cmd_in[525]), .Z(n2162));
Q_AN03 U5111 ( .A0(n38), .A1(n2163), .A2(n37), .Z(gcm_dek_cmd_in_nxt[524]));
Q_MX02 U5112 ( .S(n129), .A0(gcm_dek_cmd_in[460]), .A1(gcm_dek_cmd_in[524]), .Z(n2163));
Q_AN03 U5113 ( .A0(n38), .A1(n2164), .A2(n37), .Z(gcm_dek_cmd_in_nxt[523]));
Q_MX02 U5114 ( .S(n129), .A0(gcm_dek_cmd_in[459]), .A1(gcm_dek_cmd_in[523]), .Z(n2164));
Q_AN03 U5115 ( .A0(n38), .A1(n2165), .A2(n37), .Z(gcm_dek_cmd_in_nxt[522]));
Q_MX02 U5116 ( .S(n129), .A0(gcm_dek_cmd_in[458]), .A1(gcm_dek_cmd_in[522]), .Z(n2165));
Q_AN03 U5117 ( .A0(n38), .A1(n2166), .A2(n37), .Z(gcm_dek_cmd_in_nxt[521]));
Q_MX02 U5118 ( .S(n129), .A0(gcm_dek_cmd_in[457]), .A1(gcm_dek_cmd_in[521]), .Z(n2166));
Q_AN03 U5119 ( .A0(n38), .A1(n2167), .A2(n37), .Z(gcm_dek_cmd_in_nxt[520]));
Q_MX02 U5120 ( .S(n129), .A0(gcm_dek_cmd_in[456]), .A1(gcm_dek_cmd_in[520]), .Z(n2167));
Q_AN03 U5121 ( .A0(n38), .A1(n2168), .A2(n37), .Z(gcm_dek_cmd_in_nxt[519]));
Q_MX02 U5122 ( .S(n129), .A0(gcm_dek_cmd_in[455]), .A1(gcm_dek_cmd_in[519]), .Z(n2168));
Q_AN03 U5123 ( .A0(n38), .A1(n2169), .A2(n37), .Z(gcm_dek_cmd_in_nxt[518]));
Q_MX02 U5124 ( .S(n129), .A0(gcm_dek_cmd_in[454]), .A1(gcm_dek_cmd_in[518]), .Z(n2169));
Q_AN03 U5125 ( .A0(n38), .A1(n2170), .A2(n37), .Z(gcm_dek_cmd_in_nxt[517]));
Q_MX02 U5126 ( .S(n129), .A0(gcm_dek_cmd_in[453]), .A1(gcm_dek_cmd_in[517]), .Z(n2170));
Q_AN03 U5127 ( .A0(n38), .A1(n2171), .A2(n37), .Z(gcm_dek_cmd_in_nxt[516]));
Q_MX02 U5128 ( .S(n129), .A0(gcm_dek_cmd_in[452]), .A1(gcm_dek_cmd_in[516]), .Z(n2171));
Q_AN03 U5129 ( .A0(n38), .A1(n2172), .A2(n37), .Z(gcm_dek_cmd_in_nxt[515]));
Q_MX02 U5130 ( .S(n129), .A0(gcm_dek_cmd_in[451]), .A1(gcm_dek_cmd_in[515]), .Z(n2172));
Q_AN03 U5131 ( .A0(n38), .A1(n2173), .A2(n37), .Z(gcm_dek_cmd_in_nxt[514]));
Q_MX02 U5132 ( .S(n129), .A0(gcm_dek_cmd_in[450]), .A1(gcm_dek_cmd_in[514]), .Z(n2173));
Q_AN03 U5133 ( .A0(n38), .A1(n2174), .A2(n37), .Z(gcm_dek_cmd_in_nxt[513]));
Q_MX02 U5134 ( .S(n129), .A0(gcm_dek_cmd_in[449]), .A1(gcm_dek_cmd_in[513]), .Z(n2174));
Q_AN03 U5135 ( .A0(n38), .A1(n2175), .A2(n37), .Z(gcm_dek_cmd_in_nxt[512]));
Q_MX02 U5136 ( .S(n129), .A0(gcm_dek_cmd_in[448]), .A1(gcm_dek_cmd_in[512]), .Z(n2175));
Q_AN03 U5137 ( .A0(n38), .A1(n2176), .A2(n37), .Z(gcm_dek_cmd_in_nxt[511]));
Q_MX02 U5138 ( .S(n129), .A0(gcm_dek_cmd_in[447]), .A1(gcm_dek_cmd_in[511]), .Z(n2176));
Q_AN03 U5139 ( .A0(n38), .A1(n2177), .A2(n37), .Z(gcm_dek_cmd_in_nxt[510]));
Q_MX02 U5140 ( .S(n129), .A0(gcm_dek_cmd_in[446]), .A1(gcm_dek_cmd_in[510]), .Z(n2177));
Q_AN03 U5141 ( .A0(n38), .A1(n2178), .A2(n37), .Z(gcm_dek_cmd_in_nxt[509]));
Q_MX02 U5142 ( .S(n129), .A0(gcm_dek_cmd_in[445]), .A1(gcm_dek_cmd_in[509]), .Z(n2178));
Q_AN03 U5143 ( .A0(n38), .A1(n2179), .A2(n37), .Z(gcm_dek_cmd_in_nxt[508]));
Q_MX02 U5144 ( .S(n129), .A0(gcm_dek_cmd_in[444]), .A1(gcm_dek_cmd_in[508]), .Z(n2179));
Q_AN03 U5145 ( .A0(n38), .A1(n2180), .A2(n37), .Z(gcm_dek_cmd_in_nxt[507]));
Q_MX02 U5146 ( .S(n129), .A0(gcm_dek_cmd_in[443]), .A1(gcm_dek_cmd_in[507]), .Z(n2180));
Q_AN03 U5147 ( .A0(n38), .A1(n2181), .A2(n37), .Z(gcm_dek_cmd_in_nxt[506]));
Q_MX02 U5148 ( .S(n129), .A0(gcm_dek_cmd_in[442]), .A1(gcm_dek_cmd_in[506]), .Z(n2181));
Q_AN03 U5149 ( .A0(n38), .A1(n2182), .A2(n37), .Z(gcm_dek_cmd_in_nxt[505]));
Q_MX02 U5150 ( .S(n129), .A0(gcm_dek_cmd_in[441]), .A1(gcm_dek_cmd_in[505]), .Z(n2182));
Q_AN03 U5151 ( .A0(n38), .A1(n2183), .A2(n37), .Z(gcm_dek_cmd_in_nxt[504]));
Q_MX02 U5152 ( .S(n129), .A0(gcm_dek_cmd_in[440]), .A1(gcm_dek_cmd_in[504]), .Z(n2183));
Q_AN03 U5153 ( .A0(n38), .A1(n2184), .A2(n37), .Z(gcm_dek_cmd_in_nxt[503]));
Q_MX02 U5154 ( .S(n129), .A0(gcm_dek_cmd_in[439]), .A1(gcm_dek_cmd_in[503]), .Z(n2184));
Q_AN03 U5155 ( .A0(n38), .A1(n2185), .A2(n37), .Z(gcm_dek_cmd_in_nxt[502]));
Q_MX02 U5156 ( .S(n129), .A0(gcm_dek_cmd_in[438]), .A1(gcm_dek_cmd_in[502]), .Z(n2185));
Q_AN03 U5157 ( .A0(n38), .A1(n2186), .A2(n37), .Z(gcm_dek_cmd_in_nxt[501]));
Q_MX02 U5158 ( .S(n129), .A0(gcm_dek_cmd_in[437]), .A1(gcm_dek_cmd_in[501]), .Z(n2186));
Q_AN03 U5159 ( .A0(n38), .A1(n2187), .A2(n37), .Z(gcm_dek_cmd_in_nxt[500]));
Q_MX02 U5160 ( .S(n129), .A0(gcm_dek_cmd_in[436]), .A1(gcm_dek_cmd_in[500]), .Z(n2187));
Q_AN03 U5161 ( .A0(n38), .A1(n2188), .A2(n37), .Z(gcm_dek_cmd_in_nxt[499]));
Q_MX02 U5162 ( .S(n129), .A0(gcm_dek_cmd_in[435]), .A1(gcm_dek_cmd_in[499]), .Z(n2188));
Q_AN03 U5163 ( .A0(n38), .A1(n2189), .A2(n37), .Z(gcm_dek_cmd_in_nxt[498]));
Q_MX02 U5164 ( .S(n129), .A0(gcm_dek_cmd_in[434]), .A1(gcm_dek_cmd_in[498]), .Z(n2189));
Q_AN03 U5165 ( .A0(n38), .A1(n2190), .A2(n37), .Z(gcm_dek_cmd_in_nxt[497]));
Q_MX02 U5166 ( .S(n129), .A0(gcm_dek_cmd_in[433]), .A1(gcm_dek_cmd_in[497]), .Z(n2190));
Q_AN03 U5167 ( .A0(n38), .A1(n2191), .A2(n37), .Z(gcm_dek_cmd_in_nxt[496]));
Q_MX02 U5168 ( .S(n129), .A0(gcm_dek_cmd_in[432]), .A1(gcm_dek_cmd_in[496]), .Z(n2191));
Q_AN03 U5169 ( .A0(n38), .A1(n2192), .A2(n37), .Z(gcm_dek_cmd_in_nxt[495]));
Q_MX02 U5170 ( .S(n129), .A0(gcm_dek_cmd_in[431]), .A1(gcm_dek_cmd_in[495]), .Z(n2192));
Q_AN03 U5171 ( .A0(n38), .A1(n2193), .A2(n37), .Z(gcm_dek_cmd_in_nxt[494]));
Q_MX02 U5172 ( .S(n129), .A0(gcm_dek_cmd_in[430]), .A1(gcm_dek_cmd_in[494]), .Z(n2193));
Q_AN03 U5173 ( .A0(n38), .A1(n2194), .A2(n37), .Z(gcm_dek_cmd_in_nxt[493]));
Q_MX02 U5174 ( .S(n129), .A0(gcm_dek_cmd_in[429]), .A1(gcm_dek_cmd_in[493]), .Z(n2194));
Q_AN03 U5175 ( .A0(n38), .A1(n2195), .A2(n37), .Z(gcm_dek_cmd_in_nxt[492]));
Q_MX02 U5176 ( .S(n129), .A0(gcm_dek_cmd_in[428]), .A1(gcm_dek_cmd_in[492]), .Z(n2195));
Q_AN03 U5177 ( .A0(n38), .A1(n2196), .A2(n37), .Z(gcm_dek_cmd_in_nxt[491]));
Q_MX02 U5178 ( .S(n129), .A0(gcm_dek_cmd_in[427]), .A1(gcm_dek_cmd_in[491]), .Z(n2196));
Q_AN03 U5179 ( .A0(n38), .A1(n2197), .A2(n37), .Z(gcm_dek_cmd_in_nxt[490]));
Q_MX02 U5180 ( .S(n129), .A0(gcm_dek_cmd_in[426]), .A1(gcm_dek_cmd_in[490]), .Z(n2197));
Q_AN03 U5181 ( .A0(n38), .A1(n2198), .A2(n37), .Z(gcm_dek_cmd_in_nxt[489]));
Q_MX02 U5182 ( .S(n129), .A0(gcm_dek_cmd_in[425]), .A1(gcm_dek_cmd_in[489]), .Z(n2198));
Q_AN03 U5183 ( .A0(n38), .A1(n2199), .A2(n37), .Z(gcm_dek_cmd_in_nxt[488]));
Q_MX02 U5184 ( .S(n129), .A0(gcm_dek_cmd_in[424]), .A1(gcm_dek_cmd_in[488]), .Z(n2199));
Q_AN03 U5185 ( .A0(n38), .A1(n2200), .A2(n37), .Z(gcm_dek_cmd_in_nxt[487]));
Q_MX02 U5186 ( .S(n129), .A0(gcm_dek_cmd_in[423]), .A1(gcm_dek_cmd_in[487]), .Z(n2200));
Q_AN03 U5187 ( .A0(n38), .A1(n2201), .A2(n37), .Z(gcm_dek_cmd_in_nxt[486]));
Q_MX02 U5188 ( .S(n129), .A0(gcm_dek_cmd_in[422]), .A1(gcm_dek_cmd_in[486]), .Z(n2201));
Q_AN03 U5189 ( .A0(n38), .A1(n2202), .A2(n37), .Z(gcm_dek_cmd_in_nxt[485]));
Q_MX02 U5190 ( .S(n129), .A0(gcm_dek_cmd_in[421]), .A1(gcm_dek_cmd_in[485]), .Z(n2202));
Q_AN03 U5191 ( .A0(n38), .A1(n2203), .A2(n37), .Z(gcm_dek_cmd_in_nxt[484]));
Q_MX02 U5192 ( .S(n129), .A0(gcm_dek_cmd_in[420]), .A1(gcm_dek_cmd_in[484]), .Z(n2203));
Q_AN03 U5193 ( .A0(n38), .A1(n2204), .A2(n37), .Z(gcm_dek_cmd_in_nxt[483]));
Q_MX02 U5194 ( .S(n129), .A0(gcm_dek_cmd_in[419]), .A1(gcm_dek_cmd_in[483]), .Z(n2204));
Q_AN03 U5195 ( .A0(n38), .A1(n2205), .A2(n37), .Z(gcm_dek_cmd_in_nxt[482]));
Q_MX02 U5196 ( .S(n129), .A0(gcm_dek_cmd_in[418]), .A1(gcm_dek_cmd_in[482]), .Z(n2205));
Q_AN03 U5197 ( .A0(n38), .A1(n2206), .A2(n37), .Z(gcm_dek_cmd_in_nxt[481]));
Q_MX02 U5198 ( .S(n129), .A0(gcm_dek_cmd_in[417]), .A1(gcm_dek_cmd_in[481]), .Z(n2206));
Q_AN03 U5199 ( .A0(n38), .A1(n2207), .A2(n37), .Z(gcm_dek_cmd_in_nxt[480]));
Q_MX02 U5200 ( .S(n129), .A0(gcm_dek_cmd_in[416]), .A1(gcm_dek_cmd_in[480]), .Z(n2207));
Q_AN03 U5201 ( .A0(n38), .A1(n2208), .A2(n37), .Z(gcm_dek_cmd_in_nxt[479]));
Q_MX02 U5202 ( .S(n129), .A0(gcm_dek_cmd_in[415]), .A1(gcm_dek_cmd_in[479]), .Z(n2208));
Q_AN03 U5203 ( .A0(n38), .A1(n2209), .A2(n37), .Z(gcm_dek_cmd_in_nxt[478]));
Q_MX02 U5204 ( .S(n129), .A0(gcm_dek_cmd_in[414]), .A1(gcm_dek_cmd_in[478]), .Z(n2209));
Q_AN03 U5205 ( .A0(n38), .A1(n2210), .A2(n37), .Z(gcm_dek_cmd_in_nxt[477]));
Q_MX02 U5206 ( .S(n129), .A0(gcm_dek_cmd_in[413]), .A1(gcm_dek_cmd_in[477]), .Z(n2210));
Q_AN03 U5207 ( .A0(n38), .A1(n2211), .A2(n37), .Z(gcm_dek_cmd_in_nxt[476]));
Q_MX02 U5208 ( .S(n129), .A0(gcm_dek_cmd_in[412]), .A1(gcm_dek_cmd_in[476]), .Z(n2211));
Q_AN03 U5209 ( .A0(n38), .A1(n2212), .A2(n37), .Z(gcm_dek_cmd_in_nxt[475]));
Q_MX02 U5210 ( .S(n129), .A0(gcm_dek_cmd_in[411]), .A1(gcm_dek_cmd_in[475]), .Z(n2212));
Q_AN03 U5211 ( .A0(n38), .A1(n2213), .A2(n37), .Z(gcm_dek_cmd_in_nxt[474]));
Q_MX02 U5212 ( .S(n129), .A0(gcm_dek_cmd_in[410]), .A1(gcm_dek_cmd_in[474]), .Z(n2213));
Q_AN03 U5213 ( .A0(n38), .A1(n2214), .A2(n37), .Z(gcm_dek_cmd_in_nxt[473]));
Q_MX02 U5214 ( .S(n129), .A0(gcm_dek_cmd_in[409]), .A1(gcm_dek_cmd_in[473]), .Z(n2214));
Q_AN03 U5215 ( .A0(n38), .A1(n2215), .A2(n37), .Z(gcm_dek_cmd_in_nxt[472]));
Q_MX02 U5216 ( .S(n129), .A0(gcm_dek_cmd_in[408]), .A1(gcm_dek_cmd_in[472]), .Z(n2215));
Q_AN03 U5217 ( .A0(n38), .A1(n2216), .A2(n37), .Z(gcm_dek_cmd_in_nxt[471]));
Q_MX02 U5218 ( .S(n129), .A0(gcm_dek_cmd_in[407]), .A1(gcm_dek_cmd_in[471]), .Z(n2216));
Q_AN03 U5219 ( .A0(n38), .A1(n2217), .A2(n37), .Z(gcm_dek_cmd_in_nxt[470]));
Q_MX02 U5220 ( .S(n129), .A0(gcm_dek_cmd_in[406]), .A1(gcm_dek_cmd_in[470]), .Z(n2217));
Q_AN03 U5221 ( .A0(n38), .A1(n2218), .A2(n37), .Z(gcm_dek_cmd_in_nxt[469]));
Q_MX02 U5222 ( .S(n129), .A0(gcm_dek_cmd_in[405]), .A1(gcm_dek_cmd_in[469]), .Z(n2218));
Q_AN03 U5223 ( .A0(n38), .A1(n2219), .A2(n37), .Z(gcm_dek_cmd_in_nxt[468]));
Q_MX02 U5224 ( .S(n129), .A0(gcm_dek_cmd_in[404]), .A1(gcm_dek_cmd_in[468]), .Z(n2219));
Q_AN03 U5225 ( .A0(n38), .A1(n2220), .A2(n37), .Z(gcm_dek_cmd_in_nxt[467]));
Q_MX02 U5226 ( .S(n129), .A0(gcm_dek_cmd_in[403]), .A1(gcm_dek_cmd_in[467]), .Z(n2220));
Q_AN03 U5227 ( .A0(n38), .A1(n2221), .A2(n37), .Z(gcm_dek_cmd_in_nxt[466]));
Q_MX02 U5228 ( .S(n129), .A0(gcm_dek_cmd_in[402]), .A1(gcm_dek_cmd_in[466]), .Z(n2221));
Q_AN03 U5229 ( .A0(n38), .A1(n2222), .A2(n37), .Z(gcm_dek_cmd_in_nxt[465]));
Q_MX02 U5230 ( .S(n129), .A0(gcm_dek_cmd_in[401]), .A1(gcm_dek_cmd_in[465]), .Z(n2222));
Q_AN03 U5231 ( .A0(n38), .A1(n2223), .A2(n37), .Z(gcm_dek_cmd_in_nxt[464]));
Q_MX02 U5232 ( .S(n129), .A0(gcm_dek_cmd_in[400]), .A1(gcm_dek_cmd_in[464]), .Z(n2223));
Q_AN03 U5233 ( .A0(n38), .A1(n2224), .A2(n37), .Z(gcm_dek_cmd_in_nxt[463]));
Q_MX02 U5234 ( .S(n129), .A0(gcm_dek_cmd_in[399]), .A1(gcm_dek_cmd_in[463]), .Z(n2224));
Q_AN03 U5235 ( .A0(n38), .A1(n2225), .A2(n37), .Z(gcm_dek_cmd_in_nxt[462]));
Q_MX02 U5236 ( .S(n129), .A0(gcm_dek_cmd_in[398]), .A1(gcm_dek_cmd_in[462]), .Z(n2225));
Q_AN03 U5237 ( .A0(n38), .A1(n2226), .A2(n37), .Z(gcm_dek_cmd_in_nxt[461]));
Q_MX02 U5238 ( .S(n129), .A0(gcm_dek_cmd_in[397]), .A1(gcm_dek_cmd_in[461]), .Z(n2226));
Q_AN03 U5239 ( .A0(n38), .A1(n2227), .A2(n37), .Z(gcm_dek_cmd_in_nxt[460]));
Q_MX02 U5240 ( .S(n129), .A0(gcm_dek_cmd_in[396]), .A1(gcm_dek_cmd_in[460]), .Z(n2227));
Q_AN03 U5241 ( .A0(n38), .A1(n2228), .A2(n37), .Z(gcm_dek_cmd_in_nxt[459]));
Q_MX02 U5242 ( .S(n129), .A0(gcm_dek_cmd_in[395]), .A1(gcm_dek_cmd_in[459]), .Z(n2228));
Q_AN03 U5243 ( .A0(n38), .A1(n2229), .A2(n37), .Z(gcm_dek_cmd_in_nxt[458]));
Q_MX02 U5244 ( .S(n129), .A0(gcm_dek_cmd_in[394]), .A1(gcm_dek_cmd_in[458]), .Z(n2229));
Q_AN03 U5245 ( .A0(n38), .A1(n2230), .A2(n37), .Z(gcm_dek_cmd_in_nxt[457]));
Q_MX02 U5246 ( .S(n129), .A0(gcm_dek_cmd_in[393]), .A1(gcm_dek_cmd_in[457]), .Z(n2230));
Q_AN03 U5247 ( .A0(n38), .A1(n2231), .A2(n37), .Z(gcm_dek_cmd_in_nxt[456]));
Q_MX02 U5248 ( .S(n129), .A0(gcm_dek_cmd_in[392]), .A1(gcm_dek_cmd_in[456]), .Z(n2231));
Q_AN03 U5249 ( .A0(n38), .A1(n2232), .A2(n37), .Z(gcm_dek_cmd_in_nxt[455]));
Q_MX02 U5250 ( .S(n129), .A0(gcm_dek_cmd_in[391]), .A1(gcm_dek_cmd_in[455]), .Z(n2232));
Q_AN03 U5251 ( .A0(n38), .A1(n2233), .A2(n37), .Z(gcm_dek_cmd_in_nxt[454]));
Q_MX02 U5252 ( .S(n129), .A0(gcm_dek_cmd_in[390]), .A1(gcm_dek_cmd_in[454]), .Z(n2233));
Q_AN03 U5253 ( .A0(n38), .A1(n2234), .A2(n37), .Z(gcm_dek_cmd_in_nxt[453]));
Q_MX02 U5254 ( .S(n129), .A0(gcm_dek_cmd_in[389]), .A1(gcm_dek_cmd_in[453]), .Z(n2234));
Q_AN03 U5255 ( .A0(n38), .A1(n2235), .A2(n37), .Z(gcm_dek_cmd_in_nxt[452]));
Q_MX02 U5256 ( .S(n129), .A0(gcm_dek_cmd_in[388]), .A1(gcm_dek_cmd_in[452]), .Z(n2235));
Q_AN03 U5257 ( .A0(n38), .A1(n2236), .A2(n37), .Z(gcm_dek_cmd_in_nxt[451]));
Q_MX02 U5258 ( .S(n129), .A0(gcm_dek_cmd_in[387]), .A1(gcm_dek_cmd_in[451]), .Z(n2236));
Q_AN03 U5259 ( .A0(n38), .A1(n2237), .A2(n37), .Z(gcm_dek_cmd_in_nxt[450]));
Q_MX02 U5260 ( .S(n129), .A0(gcm_dek_cmd_in[386]), .A1(gcm_dek_cmd_in[450]), .Z(n2237));
Q_AN03 U5261 ( .A0(n38), .A1(n2238), .A2(n37), .Z(gcm_dek_cmd_in_nxt[449]));
Q_MX02 U5262 ( .S(n129), .A0(gcm_dek_cmd_in[385]), .A1(gcm_dek_cmd_in[449]), .Z(n2238));
Q_AN03 U5263 ( .A0(n38), .A1(n2239), .A2(n37), .Z(gcm_dek_cmd_in_nxt[448]));
Q_MX02 U5264 ( .S(n129), .A0(gcm_dek_cmd_in[384]), .A1(gcm_dek_cmd_in[448]), .Z(n2239));
Q_AN03 U5265 ( .A0(n38), .A1(n2240), .A2(n37), .Z(gcm_dek_cmd_in_nxt[447]));
Q_MX02 U5266 ( .S(n129), .A0(gcm_dek_cmd_in[383]), .A1(gcm_dek_cmd_in[447]), .Z(n2240));
Q_AN03 U5267 ( .A0(n38), .A1(n2241), .A2(n37), .Z(gcm_dek_cmd_in_nxt[446]));
Q_MX02 U5268 ( .S(n129), .A0(gcm_dek_cmd_in[382]), .A1(gcm_dek_cmd_in[446]), .Z(n2241));
Q_AN03 U5269 ( .A0(n38), .A1(n2242), .A2(n37), .Z(gcm_dek_cmd_in_nxt[445]));
Q_MX02 U5270 ( .S(n129), .A0(gcm_dek_cmd_in[381]), .A1(gcm_dek_cmd_in[445]), .Z(n2242));
Q_AN03 U5271 ( .A0(n38), .A1(n2243), .A2(n37), .Z(gcm_dek_cmd_in_nxt[444]));
Q_MX02 U5272 ( .S(n129), .A0(gcm_dek_cmd_in[380]), .A1(gcm_dek_cmd_in[444]), .Z(n2243));
Q_AN03 U5273 ( .A0(n38), .A1(n2244), .A2(n37), .Z(gcm_dek_cmd_in_nxt[443]));
Q_MX02 U5274 ( .S(n129), .A0(gcm_dek_cmd_in[379]), .A1(gcm_dek_cmd_in[443]), .Z(n2244));
Q_AN03 U5275 ( .A0(n38), .A1(n2245), .A2(n37), .Z(gcm_dek_cmd_in_nxt[442]));
Q_MX02 U5276 ( .S(n129), .A0(gcm_dek_cmd_in[378]), .A1(gcm_dek_cmd_in[442]), .Z(n2245));
Q_AN03 U5277 ( .A0(n38), .A1(n2246), .A2(n37), .Z(gcm_dek_cmd_in_nxt[441]));
Q_MX02 U5278 ( .S(n129), .A0(gcm_dek_cmd_in[377]), .A1(gcm_dek_cmd_in[441]), .Z(n2246));
Q_AN03 U5279 ( .A0(n38), .A1(n2247), .A2(n37), .Z(gcm_dek_cmd_in_nxt[440]));
Q_MX02 U5280 ( .S(n129), .A0(gcm_dek_cmd_in[376]), .A1(gcm_dek_cmd_in[440]), .Z(n2247));
Q_AN03 U5281 ( .A0(n38), .A1(n2248), .A2(n37), .Z(gcm_dek_cmd_in_nxt[439]));
Q_MX02 U5282 ( .S(n129), .A0(gcm_dek_cmd_in[375]), .A1(gcm_dek_cmd_in[439]), .Z(n2248));
Q_AN03 U5283 ( .A0(n38), .A1(n2249), .A2(n37), .Z(gcm_dek_cmd_in_nxt[438]));
Q_MX02 U5284 ( .S(n129), .A0(gcm_dek_cmd_in[374]), .A1(gcm_dek_cmd_in[438]), .Z(n2249));
Q_AN03 U5285 ( .A0(n38), .A1(n2250), .A2(n37), .Z(gcm_dek_cmd_in_nxt[437]));
Q_MX02 U5286 ( .S(n129), .A0(gcm_dek_cmd_in[373]), .A1(gcm_dek_cmd_in[437]), .Z(n2250));
Q_AN03 U5287 ( .A0(n38), .A1(n2251), .A2(n37), .Z(gcm_dek_cmd_in_nxt[436]));
Q_MX02 U5288 ( .S(n129), .A0(gcm_dek_cmd_in[372]), .A1(gcm_dek_cmd_in[436]), .Z(n2251));
Q_AN03 U5289 ( .A0(n38), .A1(n2252), .A2(n37), .Z(gcm_dek_cmd_in_nxt[435]));
Q_MX02 U5290 ( .S(n129), .A0(gcm_dek_cmd_in[371]), .A1(gcm_dek_cmd_in[435]), .Z(n2252));
Q_AN03 U5291 ( .A0(n38), .A1(n2253), .A2(n37), .Z(gcm_dek_cmd_in_nxt[434]));
Q_MX02 U5292 ( .S(n129), .A0(gcm_dek_cmd_in[370]), .A1(gcm_dek_cmd_in[434]), .Z(n2253));
Q_AN03 U5293 ( .A0(n38), .A1(n2254), .A2(n37), .Z(gcm_dek_cmd_in_nxt[433]));
Q_MX02 U5294 ( .S(n129), .A0(gcm_dek_cmd_in[369]), .A1(gcm_dek_cmd_in[433]), .Z(n2254));
Q_AN03 U5295 ( .A0(n38), .A1(n2255), .A2(n37), .Z(gcm_dek_cmd_in_nxt[432]));
Q_MX02 U5296 ( .S(n129), .A0(gcm_dek_cmd_in[368]), .A1(gcm_dek_cmd_in[432]), .Z(n2255));
Q_AN03 U5297 ( .A0(n38), .A1(n2256), .A2(n37), .Z(gcm_dek_cmd_in_nxt[431]));
Q_MX02 U5298 ( .S(n129), .A0(gcm_dek_cmd_in[367]), .A1(gcm_dek_cmd_in[431]), .Z(n2256));
Q_AN03 U5299 ( .A0(n38), .A1(n2257), .A2(n37), .Z(gcm_dek_cmd_in_nxt[430]));
Q_MX02 U5300 ( .S(n129), .A0(gcm_dek_cmd_in[366]), .A1(gcm_dek_cmd_in[430]), .Z(n2257));
Q_AN03 U5301 ( .A0(n38), .A1(n2258), .A2(n37), .Z(gcm_dek_cmd_in_nxt[429]));
Q_MX02 U5302 ( .S(n129), .A0(gcm_dek_cmd_in[365]), .A1(gcm_dek_cmd_in[429]), .Z(n2258));
Q_AN03 U5303 ( .A0(n38), .A1(n2259), .A2(n37), .Z(gcm_dek_cmd_in_nxt[428]));
Q_MX02 U5304 ( .S(n129), .A0(gcm_dek_cmd_in[364]), .A1(gcm_dek_cmd_in[428]), .Z(n2259));
Q_AN03 U5305 ( .A0(n38), .A1(n2260), .A2(n37), .Z(gcm_dek_cmd_in_nxt[427]));
Q_MX02 U5306 ( .S(n129), .A0(gcm_dek_cmd_in[363]), .A1(gcm_dek_cmd_in[427]), .Z(n2260));
Q_AN03 U5307 ( .A0(n38), .A1(n2261), .A2(n37), .Z(gcm_dek_cmd_in_nxt[426]));
Q_MX02 U5308 ( .S(n129), .A0(gcm_dek_cmd_in[362]), .A1(gcm_dek_cmd_in[426]), .Z(n2261));
Q_AN03 U5309 ( .A0(n38), .A1(n2262), .A2(n37), .Z(gcm_dek_cmd_in_nxt[425]));
Q_MX02 U5310 ( .S(n129), .A0(gcm_dek_cmd_in[361]), .A1(gcm_dek_cmd_in[425]), .Z(n2262));
Q_AN03 U5311 ( .A0(n38), .A1(n2263), .A2(n37), .Z(gcm_dek_cmd_in_nxt[424]));
Q_MX02 U5312 ( .S(n129), .A0(gcm_dek_cmd_in[360]), .A1(gcm_dek_cmd_in[424]), .Z(n2263));
Q_AN03 U5313 ( .A0(n38), .A1(n2264), .A2(n37), .Z(gcm_dek_cmd_in_nxt[423]));
Q_MX02 U5314 ( .S(n129), .A0(gcm_dek_cmd_in[359]), .A1(gcm_dek_cmd_in[423]), .Z(n2264));
Q_AN03 U5315 ( .A0(n38), .A1(n2265), .A2(n37), .Z(gcm_dek_cmd_in_nxt[422]));
Q_MX02 U5316 ( .S(n129), .A0(gcm_dek_cmd_in[358]), .A1(gcm_dek_cmd_in[422]), .Z(n2265));
Q_AN03 U5317 ( .A0(n38), .A1(n2266), .A2(n37), .Z(gcm_dek_cmd_in_nxt[421]));
Q_MX02 U5318 ( .S(n129), .A0(gcm_dek_cmd_in[357]), .A1(gcm_dek_cmd_in[421]), .Z(n2266));
Q_AN03 U5319 ( .A0(n38), .A1(n2267), .A2(n37), .Z(gcm_dek_cmd_in_nxt[420]));
Q_MX02 U5320 ( .S(n129), .A0(gcm_dek_cmd_in[356]), .A1(gcm_dek_cmd_in[420]), .Z(n2267));
Q_AN03 U5321 ( .A0(n38), .A1(n2268), .A2(n37), .Z(gcm_dek_cmd_in_nxt[419]));
Q_MX02 U5322 ( .S(n129), .A0(gcm_dek_cmd_in[355]), .A1(gcm_dek_cmd_in[419]), .Z(n2268));
Q_AN03 U5323 ( .A0(n38), .A1(n2269), .A2(n37), .Z(gcm_dek_cmd_in_nxt[418]));
Q_MX02 U5324 ( .S(n129), .A0(kme_internal_out[63]), .A1(gcm_dek_cmd_in[418]), .Z(n2269));
Q_AN03 U5325 ( .A0(n38), .A1(n2270), .A2(n37), .Z(gcm_dek_cmd_in_nxt[417]));
Q_MX02 U5326 ( .S(n129), .A0(kme_internal_out[62]), .A1(gcm_dek_cmd_in[417]), .Z(n2270));
Q_AN03 U5327 ( .A0(n38), .A1(n2271), .A2(n37), .Z(gcm_dek_cmd_in_nxt[416]));
Q_MX02 U5328 ( .S(n129), .A0(kme_internal_out[61]), .A1(gcm_dek_cmd_in[416]), .Z(n2271));
Q_AN03 U5329 ( .A0(n38), .A1(n2272), .A2(n37), .Z(gcm_dek_cmd_in_nxt[415]));
Q_MX02 U5330 ( .S(n129), .A0(kme_internal_out[60]), .A1(gcm_dek_cmd_in[415]), .Z(n2272));
Q_AN03 U5331 ( .A0(n38), .A1(n2273), .A2(n37), .Z(gcm_dek_cmd_in_nxt[414]));
Q_MX02 U5332 ( .S(n129), .A0(kme_internal_out[59]), .A1(gcm_dek_cmd_in[414]), .Z(n2273));
Q_AN03 U5333 ( .A0(n38), .A1(n2274), .A2(n37), .Z(gcm_dek_cmd_in_nxt[413]));
Q_MX02 U5334 ( .S(n129), .A0(kme_internal_out[58]), .A1(gcm_dek_cmd_in[413]), .Z(n2274));
Q_AN03 U5335 ( .A0(n38), .A1(n2275), .A2(n37), .Z(gcm_dek_cmd_in_nxt[412]));
Q_MX02 U5336 ( .S(n129), .A0(kme_internal_out[57]), .A1(gcm_dek_cmd_in[412]), .Z(n2275));
Q_AN03 U5337 ( .A0(n38), .A1(n2276), .A2(n37), .Z(gcm_dek_cmd_in_nxt[411]));
Q_MX02 U5338 ( .S(n129), .A0(kme_internal_out[56]), .A1(gcm_dek_cmd_in[411]), .Z(n2276));
Q_AN03 U5339 ( .A0(n38), .A1(n2277), .A2(n37), .Z(gcm_dek_cmd_in_nxt[410]));
Q_MX02 U5340 ( .S(n129), .A0(kme_internal_out[55]), .A1(gcm_dek_cmd_in[410]), .Z(n2277));
Q_AN03 U5341 ( .A0(n38), .A1(n2278), .A2(n37), .Z(gcm_dek_cmd_in_nxt[409]));
Q_MX02 U5342 ( .S(n129), .A0(kme_internal_out[54]), .A1(gcm_dek_cmd_in[409]), .Z(n2278));
Q_AN03 U5343 ( .A0(n38), .A1(n2279), .A2(n37), .Z(gcm_dek_cmd_in_nxt[408]));
Q_MX02 U5344 ( .S(n129), .A0(kme_internal_out[53]), .A1(gcm_dek_cmd_in[408]), .Z(n2279));
Q_AN03 U5345 ( .A0(n38), .A1(n2280), .A2(n37), .Z(gcm_dek_cmd_in_nxt[407]));
Q_MX02 U5346 ( .S(n129), .A0(kme_internal_out[52]), .A1(gcm_dek_cmd_in[407]), .Z(n2280));
Q_AN03 U5347 ( .A0(n38), .A1(n2281), .A2(n37), .Z(gcm_dek_cmd_in_nxt[406]));
Q_MX02 U5348 ( .S(n129), .A0(kme_internal_out[51]), .A1(gcm_dek_cmd_in[406]), .Z(n2281));
Q_AN03 U5349 ( .A0(n38), .A1(n2282), .A2(n37), .Z(gcm_dek_cmd_in_nxt[405]));
Q_MX02 U5350 ( .S(n129), .A0(kme_internal_out[50]), .A1(gcm_dek_cmd_in[405]), .Z(n2282));
Q_AN03 U5351 ( .A0(n38), .A1(n2283), .A2(n37), .Z(gcm_dek_cmd_in_nxt[404]));
Q_MX02 U5352 ( .S(n129), .A0(kme_internal_out[49]), .A1(gcm_dek_cmd_in[404]), .Z(n2283));
Q_AN03 U5353 ( .A0(n38), .A1(n2284), .A2(n37), .Z(gcm_dek_cmd_in_nxt[403]));
Q_MX02 U5354 ( .S(n129), .A0(kme_internal_out[48]), .A1(gcm_dek_cmd_in[403]), .Z(n2284));
Q_AN03 U5355 ( .A0(n38), .A1(n2285), .A2(n37), .Z(gcm_dek_cmd_in_nxt[402]));
Q_MX02 U5356 ( .S(n129), .A0(kme_internal_out[47]), .A1(gcm_dek_cmd_in[402]), .Z(n2285));
Q_AN03 U5357 ( .A0(n38), .A1(n2286), .A2(n37), .Z(gcm_dek_cmd_in_nxt[401]));
Q_MX02 U5358 ( .S(n129), .A0(kme_internal_out[46]), .A1(gcm_dek_cmd_in[401]), .Z(n2286));
Q_AN03 U5359 ( .A0(n38), .A1(n2287), .A2(n37), .Z(gcm_dek_cmd_in_nxt[400]));
Q_MX02 U5360 ( .S(n129), .A0(kme_internal_out[45]), .A1(gcm_dek_cmd_in[400]), .Z(n2287));
Q_AN03 U5361 ( .A0(n38), .A1(n2288), .A2(n37), .Z(gcm_dek_cmd_in_nxt[399]));
Q_MX02 U5362 ( .S(n129), .A0(kme_internal_out[44]), .A1(gcm_dek_cmd_in[399]), .Z(n2288));
Q_AN03 U5363 ( .A0(n38), .A1(n2289), .A2(n37), .Z(gcm_dek_cmd_in_nxt[398]));
Q_MX02 U5364 ( .S(n129), .A0(kme_internal_out[43]), .A1(gcm_dek_cmd_in[398]), .Z(n2289));
Q_AN03 U5365 ( .A0(n38), .A1(n2290), .A2(n37), .Z(gcm_dek_cmd_in_nxt[397]));
Q_MX02 U5366 ( .S(n129), .A0(kme_internal_out[42]), .A1(gcm_dek_cmd_in[397]), .Z(n2290));
Q_AN03 U5367 ( .A0(n38), .A1(n2291), .A2(n37), .Z(gcm_dek_cmd_in_nxt[396]));
Q_MX02 U5368 ( .S(n129), .A0(kme_internal_out[41]), .A1(gcm_dek_cmd_in[396]), .Z(n2291));
Q_AN03 U5369 ( .A0(n38), .A1(n2292), .A2(n37), .Z(gcm_dek_cmd_in_nxt[395]));
Q_MX02 U5370 ( .S(n129), .A0(kme_internal_out[40]), .A1(gcm_dek_cmd_in[395]), .Z(n2292));
Q_AN03 U5371 ( .A0(n38), .A1(n2293), .A2(n37), .Z(gcm_dek_cmd_in_nxt[394]));
Q_MX02 U5372 ( .S(n129), .A0(kme_internal_out[39]), .A1(gcm_dek_cmd_in[394]), .Z(n2293));
Q_AN03 U5373 ( .A0(n38), .A1(n2294), .A2(n37), .Z(gcm_dek_cmd_in_nxt[393]));
Q_MX02 U5374 ( .S(n129), .A0(kme_internal_out[38]), .A1(gcm_dek_cmd_in[393]), .Z(n2294));
Q_AN03 U5375 ( .A0(n38), .A1(n2295), .A2(n37), .Z(gcm_dek_cmd_in_nxt[392]));
Q_MX02 U5376 ( .S(n129), .A0(kme_internal_out[37]), .A1(gcm_dek_cmd_in[392]), .Z(n2295));
Q_AN03 U5377 ( .A0(n38), .A1(n2296), .A2(n37), .Z(gcm_dek_cmd_in_nxt[391]));
Q_MX02 U5378 ( .S(n129), .A0(kme_internal_out[36]), .A1(gcm_dek_cmd_in[391]), .Z(n2296));
Q_AN03 U5379 ( .A0(n38), .A1(n2297), .A2(n37), .Z(gcm_dek_cmd_in_nxt[390]));
Q_MX02 U5380 ( .S(n129), .A0(kme_internal_out[35]), .A1(gcm_dek_cmd_in[390]), .Z(n2297));
Q_AN03 U5381 ( .A0(n38), .A1(n2298), .A2(n37), .Z(gcm_dek_cmd_in_nxt[389]));
Q_MX02 U5382 ( .S(n129), .A0(kme_internal_out[34]), .A1(gcm_dek_cmd_in[389]), .Z(n2298));
Q_AN03 U5383 ( .A0(n38), .A1(n2299), .A2(n37), .Z(gcm_dek_cmd_in_nxt[388]));
Q_MX02 U5384 ( .S(n129), .A0(kme_internal_out[33]), .A1(gcm_dek_cmd_in[388]), .Z(n2299));
Q_AN03 U5385 ( .A0(n38), .A1(n2300), .A2(n37), .Z(gcm_dek_cmd_in_nxt[387]));
Q_MX02 U5386 ( .S(n129), .A0(kme_internal_out[32]), .A1(gcm_dek_cmd_in[387]), .Z(n2300));
Q_AN03 U5387 ( .A0(n38), .A1(n2301), .A2(n37), .Z(gcm_dek_cmd_in_nxt[386]));
Q_MX02 U5388 ( .S(n129), .A0(kme_internal_out[31]), .A1(gcm_dek_cmd_in[386]), .Z(n2301));
Q_AN03 U5389 ( .A0(n38), .A1(n2302), .A2(n37), .Z(gcm_dek_cmd_in_nxt[385]));
Q_MX02 U5390 ( .S(n129), .A0(kme_internal_out[30]), .A1(gcm_dek_cmd_in[385]), .Z(n2302));
Q_AN03 U5391 ( .A0(n38), .A1(n2303), .A2(n37), .Z(gcm_dek_cmd_in_nxt[384]));
Q_MX02 U5392 ( .S(n129), .A0(kme_internal_out[29]), .A1(gcm_dek_cmd_in[384]), .Z(n2303));
Q_AN03 U5393 ( .A0(n38), .A1(n2304), .A2(n37), .Z(gcm_dek_cmd_in_nxt[383]));
Q_MX02 U5394 ( .S(n129), .A0(kme_internal_out[28]), .A1(gcm_dek_cmd_in[383]), .Z(n2304));
Q_AN03 U5395 ( .A0(n38), .A1(n2305), .A2(n37), .Z(gcm_dek_cmd_in_nxt[382]));
Q_MX02 U5396 ( .S(n129), .A0(kme_internal_out[27]), .A1(gcm_dek_cmd_in[382]), .Z(n2305));
Q_AN03 U5397 ( .A0(n38), .A1(n2306), .A2(n37), .Z(gcm_dek_cmd_in_nxt[381]));
Q_MX02 U5398 ( .S(n129), .A0(kme_internal_out[26]), .A1(gcm_dek_cmd_in[381]), .Z(n2306));
Q_AN03 U5399 ( .A0(n38), .A1(n2307), .A2(n37), .Z(gcm_dek_cmd_in_nxt[380]));
Q_MX02 U5400 ( .S(n129), .A0(kme_internal_out[25]), .A1(gcm_dek_cmd_in[380]), .Z(n2307));
Q_AN03 U5401 ( .A0(n38), .A1(n2308), .A2(n37), .Z(gcm_dek_cmd_in_nxt[379]));
Q_MX02 U5402 ( .S(n129), .A0(kme_internal_out[24]), .A1(gcm_dek_cmd_in[379]), .Z(n2308));
Q_AN03 U5403 ( .A0(n38), .A1(n2309), .A2(n37), .Z(gcm_dek_cmd_in_nxt[378]));
Q_MX02 U5404 ( .S(n129), .A0(kme_internal_out[23]), .A1(gcm_dek_cmd_in[378]), .Z(n2309));
Q_AN03 U5405 ( .A0(n38), .A1(n2310), .A2(n37), .Z(gcm_dek_cmd_in_nxt[377]));
Q_MX02 U5406 ( .S(n129), .A0(kme_internal_out[22]), .A1(gcm_dek_cmd_in[377]), .Z(n2310));
Q_AN03 U5407 ( .A0(n38), .A1(n2311), .A2(n37), .Z(gcm_dek_cmd_in_nxt[376]));
Q_MX02 U5408 ( .S(n129), .A0(kme_internal_out[21]), .A1(gcm_dek_cmd_in[376]), .Z(n2311));
Q_AN03 U5409 ( .A0(n38), .A1(n2312), .A2(n37), .Z(gcm_dek_cmd_in_nxt[375]));
Q_MX02 U5410 ( .S(n129), .A0(kme_internal_out[20]), .A1(gcm_dek_cmd_in[375]), .Z(n2312));
Q_AN03 U5411 ( .A0(n38), .A1(n2313), .A2(n37), .Z(gcm_dek_cmd_in_nxt[374]));
Q_MX02 U5412 ( .S(n129), .A0(kme_internal_out[19]), .A1(gcm_dek_cmd_in[374]), .Z(n2313));
Q_AN03 U5413 ( .A0(n38), .A1(n2314), .A2(n37), .Z(gcm_dek_cmd_in_nxt[373]));
Q_MX02 U5414 ( .S(n129), .A0(kme_internal_out[18]), .A1(gcm_dek_cmd_in[373]), .Z(n2314));
Q_AN03 U5415 ( .A0(n38), .A1(n2315), .A2(n37), .Z(gcm_dek_cmd_in_nxt[372]));
Q_MX02 U5416 ( .S(n129), .A0(kme_internal_out[17]), .A1(gcm_dek_cmd_in[372]), .Z(n2315));
Q_AN03 U5417 ( .A0(n38), .A1(n2316), .A2(n37), .Z(gcm_dek_cmd_in_nxt[371]));
Q_MX02 U5418 ( .S(n129), .A0(kme_internal_out[16]), .A1(gcm_dek_cmd_in[371]), .Z(n2316));
Q_AN03 U5419 ( .A0(n38), .A1(n2317), .A2(n37), .Z(gcm_dek_cmd_in_nxt[370]));
Q_MX02 U5420 ( .S(n129), .A0(kme_internal_out[15]), .A1(gcm_dek_cmd_in[370]), .Z(n2317));
Q_AN03 U5421 ( .A0(n38), .A1(n2318), .A2(n37), .Z(gcm_dek_cmd_in_nxt[369]));
Q_MX02 U5422 ( .S(n129), .A0(kme_internal_out[14]), .A1(gcm_dek_cmd_in[369]), .Z(n2318));
Q_AN03 U5423 ( .A0(n38), .A1(n2319), .A2(n37), .Z(gcm_dek_cmd_in_nxt[368]));
Q_MX02 U5424 ( .S(n129), .A0(kme_internal_out[13]), .A1(gcm_dek_cmd_in[368]), .Z(n2319));
Q_AN03 U5425 ( .A0(n38), .A1(n2320), .A2(n37), .Z(gcm_dek_cmd_in_nxt[367]));
Q_MX02 U5426 ( .S(n129), .A0(kme_internal_out[12]), .A1(gcm_dek_cmd_in[367]), .Z(n2320));
Q_AN03 U5427 ( .A0(n38), .A1(n2321), .A2(n37), .Z(gcm_dek_cmd_in_nxt[366]));
Q_MX02 U5428 ( .S(n129), .A0(kme_internal_out[11]), .A1(gcm_dek_cmd_in[366]), .Z(n2321));
Q_AN03 U5429 ( .A0(n38), .A1(n2322), .A2(n37), .Z(gcm_dek_cmd_in_nxt[365]));
Q_MX02 U5430 ( .S(n129), .A0(kme_internal_out[10]), .A1(gcm_dek_cmd_in[365]), .Z(n2322));
Q_AN03 U5431 ( .A0(n38), .A1(n2323), .A2(n37), .Z(gcm_dek_cmd_in_nxt[364]));
Q_MX02 U5432 ( .S(n129), .A0(kme_internal_out[9]), .A1(gcm_dek_cmd_in[364]), .Z(n2323));
Q_AN03 U5433 ( .A0(n38), .A1(n2324), .A2(n37), .Z(gcm_dek_cmd_in_nxt[363]));
Q_MX02 U5434 ( .S(n129), .A0(kme_internal_out[8]), .A1(gcm_dek_cmd_in[363]), .Z(n2324));
Q_AN03 U5435 ( .A0(n38), .A1(n2325), .A2(n37), .Z(gcm_dek_cmd_in_nxt[362]));
Q_MX02 U5436 ( .S(n129), .A0(kme_internal_out[7]), .A1(gcm_dek_cmd_in[362]), .Z(n2325));
Q_AN03 U5437 ( .A0(n38), .A1(n2326), .A2(n37), .Z(gcm_dek_cmd_in_nxt[361]));
Q_MX02 U5438 ( .S(n129), .A0(kme_internal_out[6]), .A1(gcm_dek_cmd_in[361]), .Z(n2326));
Q_AN03 U5439 ( .A0(n38), .A1(n2327), .A2(n37), .Z(gcm_dek_cmd_in_nxt[360]));
Q_MX02 U5440 ( .S(n129), .A0(kme_internal_out[5]), .A1(gcm_dek_cmd_in[360]), .Z(n2327));
Q_AN03 U5441 ( .A0(n38), .A1(n2328), .A2(n37), .Z(gcm_dek_cmd_in_nxt[359]));
Q_MX02 U5442 ( .S(n129), .A0(kme_internal_out[4]), .A1(gcm_dek_cmd_in[359]), .Z(n2328));
Q_AN03 U5443 ( .A0(n38), .A1(n2329), .A2(n37), .Z(gcm_dek_cmd_in_nxt[358]));
Q_MX02 U5444 ( .S(n129), .A0(kme_internal_out[3]), .A1(gcm_dek_cmd_in[358]), .Z(n2329));
Q_AN03 U5445 ( .A0(n38), .A1(n2330), .A2(n37), .Z(gcm_dek_cmd_in_nxt[357]));
Q_MX02 U5446 ( .S(n129), .A0(kme_internal_out[2]), .A1(gcm_dek_cmd_in[357]), .Z(n2330));
Q_AN03 U5447 ( .A0(n38), .A1(n2331), .A2(n37), .Z(gcm_dek_cmd_in_nxt[356]));
Q_MX02 U5448 ( .S(n129), .A0(kme_internal_out[1]), .A1(gcm_dek_cmd_in[356]), .Z(n2331));
Q_AN03 U5449 ( .A0(n38), .A1(n2332), .A2(n37), .Z(gcm_dek_cmd_in_nxt[355]));
Q_MX02 U5450 ( .S(n129), .A0(kme_internal_out[0]), .A1(gcm_dek_cmd_in[355]), .Z(n2332));
Q_MX02 U5451 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[31]), .A1(kme_internal_out[63]), .Z(n2333));
Q_MX02 U5452 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[30]), .A1(kme_internal_out[62]), .Z(n2334));
Q_MX02 U5453 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[29]), .A1(kme_internal_out[61]), .Z(n2335));
Q_MX02 U5454 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[28]), .A1(kme_internal_out[60]), .Z(n2336));
Q_MX02 U5455 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[27]), .A1(kme_internal_out[59]), .Z(n2337));
Q_MX02 U5456 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[26]), .A1(kme_internal_out[58]), .Z(n2338));
Q_MX02 U5457 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[25]), .A1(kme_internal_out[57]), .Z(n2339));
Q_MX02 U5458 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[24]), .A1(kme_internal_out[56]), .Z(n2340));
Q_MX02 U5459 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[23]), .A1(kme_internal_out[55]), .Z(n2341));
Q_MX02 U5460 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[22]), .A1(kme_internal_out[54]), .Z(n2342));
Q_MX02 U5461 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[21]), .A1(kme_internal_out[53]), .Z(n2343));
Q_MX02 U5462 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[20]), .A1(kme_internal_out[52]), .Z(n2344));
Q_MX02 U5463 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[19]), .A1(kme_internal_out[51]), .Z(n2345));
Q_MX02 U5464 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[18]), .A1(kme_internal_out[50]), .Z(n2346));
Q_MX02 U5465 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[17]), .A1(kme_internal_out[49]), .Z(n2347));
Q_MX02 U5466 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[16]), .A1(kme_internal_out[48]), .Z(n2348));
Q_MX02 U5467 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[15]), .A1(kme_internal_out[47]), .Z(n2349));
Q_MX02 U5468 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[14]), .A1(kme_internal_out[46]), .Z(n2350));
Q_MX02 U5469 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[13]), .A1(kme_internal_out[45]), .Z(n2351));
Q_MX02 U5470 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[12]), .A1(kme_internal_out[44]), .Z(n2352));
Q_MX02 U5471 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[11]), .A1(kme_internal_out[43]), .Z(n2353));
Q_MX02 U5472 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[10]), .A1(kme_internal_out[42]), .Z(n2354));
Q_MX02 U5473 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[9]), .A1(kme_internal_out[41]), .Z(n2355));
Q_MX02 U5474 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[8]), .A1(kme_internal_out[40]), .Z(n2356));
Q_MX02 U5475 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[7]), .A1(kme_internal_out[39]), .Z(n2357));
Q_MX02 U5476 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[6]), .A1(kme_internal_out[38]), .Z(n2358));
Q_MX02 U5477 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[5]), .A1(kme_internal_out[37]), .Z(n2359));
Q_MX02 U5478 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[4]), .A1(kme_internal_out[36]), .Z(n2360));
Q_MX02 U5479 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[3]), .A1(kme_internal_out[35]), .Z(n2361));
Q_MX02 U5480 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[2]), .A1(kme_internal_out[34]), .Z(n2362));
Q_MX02 U5481 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[1]), .A1(kme_internal_out[33]), .Z(n2363));
Q_MX02 U5482 ( .S(kme_internal_out[69]), .A0(gcm_dak_tag[0]), .A1(kme_internal_out[32]), .Z(n2364));
Q_MX02 U5483 ( .S(kme_internal_out[69]), .A0(kme_internal_out[63]), .A1(gcm_dak_tag[95]), .Z(n2365));
Q_MX02 U5484 ( .S(kme_internal_out[69]), .A0(kme_internal_out[62]), .A1(gcm_dak_tag[94]), .Z(n2366));
Q_MX02 U5485 ( .S(kme_internal_out[69]), .A0(kme_internal_out[61]), .A1(gcm_dak_tag[93]), .Z(n2367));
Q_MX02 U5486 ( .S(kme_internal_out[69]), .A0(kme_internal_out[60]), .A1(gcm_dak_tag[92]), .Z(n2368));
Q_MX02 U5487 ( .S(kme_internal_out[69]), .A0(kme_internal_out[59]), .A1(gcm_dak_tag[91]), .Z(n2369));
Q_MX02 U5488 ( .S(kme_internal_out[69]), .A0(kme_internal_out[58]), .A1(gcm_dak_tag[90]), .Z(n2370));
Q_MX02 U5489 ( .S(kme_internal_out[69]), .A0(kme_internal_out[57]), .A1(gcm_dak_tag[89]), .Z(n2371));
Q_MX02 U5490 ( .S(kme_internal_out[69]), .A0(kme_internal_out[56]), .A1(gcm_dak_tag[88]), .Z(n2372));
Q_MX02 U5491 ( .S(kme_internal_out[69]), .A0(kme_internal_out[55]), .A1(gcm_dak_tag[87]), .Z(n2373));
Q_MX02 U5492 ( .S(kme_internal_out[69]), .A0(kme_internal_out[54]), .A1(gcm_dak_tag[86]), .Z(n2374));
Q_MX02 U5493 ( .S(kme_internal_out[69]), .A0(kme_internal_out[53]), .A1(gcm_dak_tag[85]), .Z(n2375));
Q_MX02 U5494 ( .S(kme_internal_out[69]), .A0(kme_internal_out[52]), .A1(gcm_dak_tag[84]), .Z(n2376));
Q_MX02 U5495 ( .S(kme_internal_out[69]), .A0(kme_internal_out[51]), .A1(gcm_dak_tag[83]), .Z(n2377));
Q_MX02 U5496 ( .S(kme_internal_out[69]), .A0(kme_internal_out[50]), .A1(gcm_dak_tag[82]), .Z(n2378));
Q_MX02 U5497 ( .S(kme_internal_out[69]), .A0(kme_internal_out[49]), .A1(gcm_dak_tag[81]), .Z(n2379));
Q_MX02 U5498 ( .S(kme_internal_out[69]), .A0(kme_internal_out[48]), .A1(gcm_dak_tag[80]), .Z(n2380));
Q_MX02 U5499 ( .S(kme_internal_out[69]), .A0(kme_internal_out[47]), .A1(gcm_dak_tag[79]), .Z(n2381));
Q_MX02 U5500 ( .S(kme_internal_out[69]), .A0(kme_internal_out[46]), .A1(gcm_dak_tag[78]), .Z(n2382));
Q_MX02 U5501 ( .S(kme_internal_out[69]), .A0(kme_internal_out[45]), .A1(gcm_dak_tag[77]), .Z(n2383));
Q_MX02 U5502 ( .S(kme_internal_out[69]), .A0(kme_internal_out[44]), .A1(gcm_dak_tag[76]), .Z(n2384));
Q_MX02 U5503 ( .S(kme_internal_out[69]), .A0(kme_internal_out[43]), .A1(gcm_dak_tag[75]), .Z(n2385));
Q_MX02 U5504 ( .S(kme_internal_out[69]), .A0(kme_internal_out[42]), .A1(gcm_dak_tag[74]), .Z(n2386));
Q_MX02 U5505 ( .S(kme_internal_out[69]), .A0(kme_internal_out[41]), .A1(gcm_dak_tag[73]), .Z(n2387));
Q_MX02 U5506 ( .S(kme_internal_out[69]), .A0(kme_internal_out[40]), .A1(gcm_dak_tag[72]), .Z(n2388));
Q_MX02 U5507 ( .S(kme_internal_out[69]), .A0(kme_internal_out[39]), .A1(gcm_dak_tag[71]), .Z(n2389));
Q_MX02 U5508 ( .S(kme_internal_out[69]), .A0(kme_internal_out[38]), .A1(gcm_dak_tag[70]), .Z(n2390));
Q_MX02 U5509 ( .S(kme_internal_out[69]), .A0(kme_internal_out[37]), .A1(gcm_dak_tag[69]), .Z(n2391));
Q_MX02 U5510 ( .S(kme_internal_out[69]), .A0(kme_internal_out[36]), .A1(gcm_dak_tag[68]), .Z(n2392));
Q_MX02 U5511 ( .S(kme_internal_out[69]), .A0(kme_internal_out[35]), .A1(gcm_dak_tag[67]), .Z(n2393));
Q_MX02 U5512 ( .S(kme_internal_out[69]), .A0(kme_internal_out[34]), .A1(gcm_dak_tag[66]), .Z(n2394));
Q_MX02 U5513 ( .S(kme_internal_out[69]), .A0(kme_internal_out[33]), .A1(gcm_dak_tag[65]), .Z(n2395));
Q_MX02 U5514 ( .S(kme_internal_out[69]), .A0(kme_internal_out[32]), .A1(gcm_dak_tag[64]), .Z(n2396));
Q_MX02 U5515 ( .S(kme_internal_out[69]), .A0(kme_internal_out[31]), .A1(gcm_dak_tag[63]), .Z(n2397));
Q_MX02 U5516 ( .S(kme_internal_out[69]), .A0(kme_internal_out[30]), .A1(gcm_dak_tag[62]), .Z(n2398));
Q_MX02 U5517 ( .S(kme_internal_out[69]), .A0(kme_internal_out[29]), .A1(gcm_dak_tag[61]), .Z(n2399));
Q_MX02 U5518 ( .S(kme_internal_out[69]), .A0(kme_internal_out[28]), .A1(gcm_dak_tag[60]), .Z(n2400));
Q_MX02 U5519 ( .S(kme_internal_out[69]), .A0(kme_internal_out[27]), .A1(gcm_dak_tag[59]), .Z(n2401));
Q_MX02 U5520 ( .S(kme_internal_out[69]), .A0(kme_internal_out[26]), .A1(gcm_dak_tag[58]), .Z(n2402));
Q_MX02 U5521 ( .S(kme_internal_out[69]), .A0(kme_internal_out[25]), .A1(gcm_dak_tag[57]), .Z(n2403));
Q_MX02 U5522 ( .S(kme_internal_out[69]), .A0(kme_internal_out[24]), .A1(gcm_dak_tag[56]), .Z(n2404));
Q_MX02 U5523 ( .S(kme_internal_out[69]), .A0(kme_internal_out[23]), .A1(gcm_dak_tag[55]), .Z(n2405));
Q_MX02 U5524 ( .S(kme_internal_out[69]), .A0(kme_internal_out[22]), .A1(gcm_dak_tag[54]), .Z(n2406));
Q_MX02 U5525 ( .S(kme_internal_out[69]), .A0(kme_internal_out[21]), .A1(gcm_dak_tag[53]), .Z(n2407));
Q_MX02 U5526 ( .S(kme_internal_out[69]), .A0(kme_internal_out[20]), .A1(gcm_dak_tag[52]), .Z(n2408));
Q_MX02 U5527 ( .S(kme_internal_out[69]), .A0(kme_internal_out[19]), .A1(gcm_dak_tag[51]), .Z(n2409));
Q_MX02 U5528 ( .S(kme_internal_out[69]), .A0(kme_internal_out[18]), .A1(gcm_dak_tag[50]), .Z(n2410));
Q_MX02 U5529 ( .S(kme_internal_out[69]), .A0(kme_internal_out[17]), .A1(gcm_dak_tag[49]), .Z(n2411));
Q_MX02 U5530 ( .S(kme_internal_out[69]), .A0(kme_internal_out[16]), .A1(gcm_dak_tag[48]), .Z(n2412));
Q_MX02 U5531 ( .S(kme_internal_out[69]), .A0(kme_internal_out[15]), .A1(gcm_dak_tag[47]), .Z(n2413));
Q_MX02 U5532 ( .S(kme_internal_out[69]), .A0(kme_internal_out[14]), .A1(gcm_dak_tag[46]), .Z(n2414));
Q_MX02 U5533 ( .S(kme_internal_out[69]), .A0(kme_internal_out[13]), .A1(gcm_dak_tag[45]), .Z(n2415));
Q_MX02 U5534 ( .S(kme_internal_out[69]), .A0(kme_internal_out[12]), .A1(gcm_dak_tag[44]), .Z(n2416));
Q_MX02 U5535 ( .S(kme_internal_out[69]), .A0(kme_internal_out[11]), .A1(gcm_dak_tag[43]), .Z(n2417));
Q_MX02 U5536 ( .S(kme_internal_out[69]), .A0(kme_internal_out[10]), .A1(gcm_dak_tag[42]), .Z(n2418));
Q_MX02 U5537 ( .S(kme_internal_out[69]), .A0(kme_internal_out[9]), .A1(gcm_dak_tag[41]), .Z(n2419));
Q_MX02 U5538 ( .S(kme_internal_out[69]), .A0(kme_internal_out[8]), .A1(gcm_dak_tag[40]), .Z(n2420));
Q_MX02 U5539 ( .S(kme_internal_out[69]), .A0(kme_internal_out[7]), .A1(gcm_dak_tag[39]), .Z(n2421));
Q_MX02 U5540 ( .S(kme_internal_out[69]), .A0(kme_internal_out[6]), .A1(gcm_dak_tag[38]), .Z(n2422));
Q_MX02 U5541 ( .S(kme_internal_out[69]), .A0(kme_internal_out[5]), .A1(gcm_dak_tag[37]), .Z(n2423));
Q_MX02 U5542 ( .S(kme_internal_out[69]), .A0(kme_internal_out[4]), .A1(gcm_dak_tag[36]), .Z(n2424));
Q_MX02 U5543 ( .S(kme_internal_out[69]), .A0(kme_internal_out[3]), .A1(gcm_dak_tag[35]), .Z(n2425));
Q_MX02 U5544 ( .S(kme_internal_out[69]), .A0(kme_internal_out[2]), .A1(gcm_dak_tag[34]), .Z(n2426));
Q_MX02 U5545 ( .S(kme_internal_out[69]), .A0(kme_internal_out[1]), .A1(gcm_dak_tag[33]), .Z(n2427));
Q_MX02 U5546 ( .S(kme_internal_out[69]), .A0(kme_internal_out[0]), .A1(gcm_dak_tag[32]), .Z(n2428));
Q_MX02 U5547 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[31]), .A1(kme_internal_out[63]), .Z(n2429));
Q_MX02 U5548 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[30]), .A1(kme_internal_out[62]), .Z(n2430));
Q_MX02 U5549 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[29]), .A1(kme_internal_out[61]), .Z(n2431));
Q_MX02 U5550 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[28]), .A1(kme_internal_out[60]), .Z(n2432));
Q_MX02 U5551 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[27]), .A1(kme_internal_out[59]), .Z(n2433));
Q_MX02 U5552 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[26]), .A1(kme_internal_out[58]), .Z(n2434));
Q_MX02 U5553 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[25]), .A1(kme_internal_out[57]), .Z(n2435));
Q_MX02 U5554 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[24]), .A1(kme_internal_out[56]), .Z(n2436));
Q_MX02 U5555 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[23]), .A1(kme_internal_out[55]), .Z(n2437));
Q_MX02 U5556 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[22]), .A1(kme_internal_out[54]), .Z(n2438));
Q_MX02 U5557 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[21]), .A1(kme_internal_out[53]), .Z(n2439));
Q_MX02 U5558 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[20]), .A1(kme_internal_out[52]), .Z(n2440));
Q_MX02 U5559 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[19]), .A1(kme_internal_out[51]), .Z(n2441));
Q_MX02 U5560 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[18]), .A1(kme_internal_out[50]), .Z(n2442));
Q_MX02 U5561 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[17]), .A1(kme_internal_out[49]), .Z(n2443));
Q_MX02 U5562 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[16]), .A1(kme_internal_out[48]), .Z(n2444));
Q_MX02 U5563 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[15]), .A1(kme_internal_out[47]), .Z(n2445));
Q_MX02 U5564 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[14]), .A1(kme_internal_out[46]), .Z(n2446));
Q_MX02 U5565 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[13]), .A1(kme_internal_out[45]), .Z(n2447));
Q_MX02 U5566 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[12]), .A1(kme_internal_out[44]), .Z(n2448));
Q_MX02 U5567 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[11]), .A1(kme_internal_out[43]), .Z(n2449));
Q_MX02 U5568 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[10]), .A1(kme_internal_out[42]), .Z(n2450));
Q_MX02 U5569 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[9]), .A1(kme_internal_out[41]), .Z(n2451));
Q_MX02 U5570 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[8]), .A1(kme_internal_out[40]), .Z(n2452));
Q_MX02 U5571 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[7]), .A1(kme_internal_out[39]), .Z(n2453));
Q_MX02 U5572 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[6]), .A1(kme_internal_out[38]), .Z(n2454));
Q_MX02 U5573 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[5]), .A1(kme_internal_out[37]), .Z(n2455));
Q_MX02 U5574 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[4]), .A1(kme_internal_out[36]), .Z(n2456));
Q_MX02 U5575 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[3]), .A1(kme_internal_out[35]), .Z(n2457));
Q_MX02 U5576 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[2]), .A1(kme_internal_out[34]), .Z(n2458));
Q_MX02 U5577 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[1]), .A1(kme_internal_out[33]), .Z(n2459));
Q_MX02 U5578 ( .S(kme_internal_out[69]), .A0(gcm_dek_tag[0]), .A1(kme_internal_out[32]), .Z(n2460));
Q_MX02 U5579 ( .S(kme_internal_out[69]), .A0(kme_internal_out[63]), .A1(gcm_dek_tag[95]), .Z(n2461));
Q_MX02 U5580 ( .S(kme_internal_out[69]), .A0(kme_internal_out[62]), .A1(gcm_dek_tag[94]), .Z(n2462));
Q_MX02 U5581 ( .S(kme_internal_out[69]), .A0(kme_internal_out[61]), .A1(gcm_dek_tag[93]), .Z(n2463));
Q_MX02 U5582 ( .S(kme_internal_out[69]), .A0(kme_internal_out[60]), .A1(gcm_dek_tag[92]), .Z(n2464));
Q_MX02 U5583 ( .S(kme_internal_out[69]), .A0(kme_internal_out[59]), .A1(gcm_dek_tag[91]), .Z(n2465));
Q_MX02 U5584 ( .S(kme_internal_out[69]), .A0(kme_internal_out[58]), .A1(gcm_dek_tag[90]), .Z(n2466));
Q_MX02 U5585 ( .S(kme_internal_out[69]), .A0(kme_internal_out[57]), .A1(gcm_dek_tag[89]), .Z(n2467));
Q_MX02 U5586 ( .S(kme_internal_out[69]), .A0(kme_internal_out[56]), .A1(gcm_dek_tag[88]), .Z(n2468));
Q_MX02 U5587 ( .S(kme_internal_out[69]), .A0(kme_internal_out[55]), .A1(gcm_dek_tag[87]), .Z(n2469));
Q_MX02 U5588 ( .S(kme_internal_out[69]), .A0(kme_internal_out[54]), .A1(gcm_dek_tag[86]), .Z(n2470));
Q_MX02 U5589 ( .S(kme_internal_out[69]), .A0(kme_internal_out[53]), .A1(gcm_dek_tag[85]), .Z(n2471));
Q_MX02 U5590 ( .S(kme_internal_out[69]), .A0(kme_internal_out[52]), .A1(gcm_dek_tag[84]), .Z(n2472));
Q_MX02 U5591 ( .S(kme_internal_out[69]), .A0(kme_internal_out[51]), .A1(gcm_dek_tag[83]), .Z(n2473));
Q_MX02 U5592 ( .S(kme_internal_out[69]), .A0(kme_internal_out[50]), .A1(gcm_dek_tag[82]), .Z(n2474));
Q_MX02 U5593 ( .S(kme_internal_out[69]), .A0(kme_internal_out[49]), .A1(gcm_dek_tag[81]), .Z(n2475));
Q_MX02 U5594 ( .S(kme_internal_out[69]), .A0(kme_internal_out[48]), .A1(gcm_dek_tag[80]), .Z(n2476));
Q_MX02 U5595 ( .S(kme_internal_out[69]), .A0(kme_internal_out[47]), .A1(gcm_dek_tag[79]), .Z(n2477));
Q_MX02 U5596 ( .S(kme_internal_out[69]), .A0(kme_internal_out[46]), .A1(gcm_dek_tag[78]), .Z(n2478));
Q_MX02 U5597 ( .S(kme_internal_out[69]), .A0(kme_internal_out[45]), .A1(gcm_dek_tag[77]), .Z(n2479));
Q_MX02 U5598 ( .S(kme_internal_out[69]), .A0(kme_internal_out[44]), .A1(gcm_dek_tag[76]), .Z(n2480));
Q_MX02 U5599 ( .S(kme_internal_out[69]), .A0(kme_internal_out[43]), .A1(gcm_dek_tag[75]), .Z(n2481));
Q_MX02 U5600 ( .S(kme_internal_out[69]), .A0(kme_internal_out[42]), .A1(gcm_dek_tag[74]), .Z(n2482));
Q_MX02 U5601 ( .S(kme_internal_out[69]), .A0(kme_internal_out[41]), .A1(gcm_dek_tag[73]), .Z(n2483));
Q_MX02 U5602 ( .S(kme_internal_out[69]), .A0(kme_internal_out[40]), .A1(gcm_dek_tag[72]), .Z(n2484));
Q_MX02 U5603 ( .S(kme_internal_out[69]), .A0(kme_internal_out[39]), .A1(gcm_dek_tag[71]), .Z(n2485));
Q_MX02 U5604 ( .S(kme_internal_out[69]), .A0(kme_internal_out[38]), .A1(gcm_dek_tag[70]), .Z(n2486));
Q_MX02 U5605 ( .S(kme_internal_out[69]), .A0(kme_internal_out[37]), .A1(gcm_dek_tag[69]), .Z(n2487));
Q_MX02 U5606 ( .S(kme_internal_out[69]), .A0(kme_internal_out[36]), .A1(gcm_dek_tag[68]), .Z(n2488));
Q_MX02 U5607 ( .S(kme_internal_out[69]), .A0(kme_internal_out[35]), .A1(gcm_dek_tag[67]), .Z(n2489));
Q_MX02 U5608 ( .S(kme_internal_out[69]), .A0(kme_internal_out[34]), .A1(gcm_dek_tag[66]), .Z(n2490));
Q_MX02 U5609 ( .S(kme_internal_out[69]), .A0(kme_internal_out[33]), .A1(gcm_dek_tag[65]), .Z(n2491));
Q_MX02 U5610 ( .S(kme_internal_out[69]), .A0(kme_internal_out[32]), .A1(gcm_dek_tag[64]), .Z(n2492));
Q_MX02 U5611 ( .S(kme_internal_out[69]), .A0(kme_internal_out[31]), .A1(gcm_dek_tag[63]), .Z(n2493));
Q_MX02 U5612 ( .S(kme_internal_out[69]), .A0(kme_internal_out[30]), .A1(gcm_dek_tag[62]), .Z(n2494));
Q_MX02 U5613 ( .S(kme_internal_out[69]), .A0(kme_internal_out[29]), .A1(gcm_dek_tag[61]), .Z(n2495));
Q_MX02 U5614 ( .S(kme_internal_out[69]), .A0(kme_internal_out[28]), .A1(gcm_dek_tag[60]), .Z(n2496));
Q_MX02 U5615 ( .S(kme_internal_out[69]), .A0(kme_internal_out[27]), .A1(gcm_dek_tag[59]), .Z(n2497));
Q_MX02 U5616 ( .S(kme_internal_out[69]), .A0(kme_internal_out[26]), .A1(gcm_dek_tag[58]), .Z(n2498));
Q_MX02 U5617 ( .S(kme_internal_out[69]), .A0(kme_internal_out[25]), .A1(gcm_dek_tag[57]), .Z(n2499));
Q_MX02 U5618 ( .S(kme_internal_out[69]), .A0(kme_internal_out[24]), .A1(gcm_dek_tag[56]), .Z(n2500));
Q_MX02 U5619 ( .S(kme_internal_out[69]), .A0(kme_internal_out[23]), .A1(gcm_dek_tag[55]), .Z(n2501));
Q_MX02 U5620 ( .S(kme_internal_out[69]), .A0(kme_internal_out[22]), .A1(gcm_dek_tag[54]), .Z(n2502));
Q_MX02 U5621 ( .S(kme_internal_out[69]), .A0(kme_internal_out[21]), .A1(gcm_dek_tag[53]), .Z(n2503));
Q_MX02 U5622 ( .S(kme_internal_out[69]), .A0(kme_internal_out[20]), .A1(gcm_dek_tag[52]), .Z(n2504));
Q_MX02 U5623 ( .S(kme_internal_out[69]), .A0(kme_internal_out[19]), .A1(gcm_dek_tag[51]), .Z(n2505));
Q_MX02 U5624 ( .S(kme_internal_out[69]), .A0(kme_internal_out[18]), .A1(gcm_dek_tag[50]), .Z(n2506));
Q_MX02 U5625 ( .S(kme_internal_out[69]), .A0(kme_internal_out[17]), .A1(gcm_dek_tag[49]), .Z(n2507));
Q_MX02 U5626 ( .S(kme_internal_out[69]), .A0(kme_internal_out[16]), .A1(gcm_dek_tag[48]), .Z(n2508));
Q_MX02 U5627 ( .S(kme_internal_out[69]), .A0(kme_internal_out[15]), .A1(gcm_dek_tag[47]), .Z(n2509));
Q_MX02 U5628 ( .S(kme_internal_out[69]), .A0(kme_internal_out[14]), .A1(gcm_dek_tag[46]), .Z(n2510));
Q_MX02 U5629 ( .S(kme_internal_out[69]), .A0(kme_internal_out[13]), .A1(gcm_dek_tag[45]), .Z(n2511));
Q_MX02 U5630 ( .S(kme_internal_out[69]), .A0(kme_internal_out[12]), .A1(gcm_dek_tag[44]), .Z(n2512));
Q_MX02 U5631 ( .S(kme_internal_out[69]), .A0(kme_internal_out[11]), .A1(gcm_dek_tag[43]), .Z(n2513));
Q_MX02 U5632 ( .S(kme_internal_out[69]), .A0(kme_internal_out[10]), .A1(gcm_dek_tag[42]), .Z(n2514));
Q_MX02 U5633 ( .S(kme_internal_out[69]), .A0(kme_internal_out[9]), .A1(gcm_dek_tag[41]), .Z(n2515));
Q_MX02 U5634 ( .S(kme_internal_out[69]), .A0(kme_internal_out[8]), .A1(gcm_dek_tag[40]), .Z(n2516));
Q_MX02 U5635 ( .S(kme_internal_out[69]), .A0(kme_internal_out[7]), .A1(gcm_dek_tag[39]), .Z(n2517));
Q_MX02 U5636 ( .S(kme_internal_out[69]), .A0(kme_internal_out[6]), .A1(gcm_dek_tag[38]), .Z(n2518));
Q_MX02 U5637 ( .S(kme_internal_out[69]), .A0(kme_internal_out[5]), .A1(gcm_dek_tag[37]), .Z(n2519));
Q_MX02 U5638 ( .S(kme_internal_out[69]), .A0(kme_internal_out[4]), .A1(gcm_dek_tag[36]), .Z(n2520));
Q_MX02 U5639 ( .S(kme_internal_out[69]), .A0(kme_internal_out[3]), .A1(gcm_dek_tag[35]), .Z(n2521));
Q_MX02 U5640 ( .S(kme_internal_out[69]), .A0(kme_internal_out[2]), .A1(gcm_dek_tag[34]), .Z(n2522));
Q_MX02 U5641 ( .S(kme_internal_out[69]), .A0(kme_internal_out[1]), .A1(gcm_dek_tag[33]), .Z(n2523));
Q_MX02 U5642 ( .S(kme_internal_out[69]), .A0(kme_internal_out[0]), .A1(gcm_dek_tag[32]), .Z(n2524));
Q_MX02 U5643 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[34]), .A1(kme_internal_out[63]), .Z(n2525));
Q_MX02 U5644 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[33]), .A1(kme_internal_out[62]), .Z(n2526));
Q_MX02 U5645 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[32]), .A1(kme_internal_out[61]), .Z(n2527));
Q_MX02 U5646 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[31]), .A1(kme_internal_out[60]), .Z(n2528));
Q_MX02 U5647 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[30]), .A1(kme_internal_out[59]), .Z(n2529));
Q_MX02 U5648 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[29]), .A1(kme_internal_out[58]), .Z(n2530));
Q_MX02 U5649 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[28]), .A1(kme_internal_out[57]), .Z(n2531));
Q_MX02 U5650 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[27]), .A1(kme_internal_out[56]), .Z(n2532));
Q_MX02 U5651 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[26]), .A1(kme_internal_out[55]), .Z(n2533));
Q_MX02 U5652 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[25]), .A1(kme_internal_out[54]), .Z(n2534));
Q_MX02 U5653 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[24]), .A1(kme_internal_out[53]), .Z(n2535));
Q_MX02 U5654 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[23]), .A1(kme_internal_out[52]), .Z(n2536));
Q_MX02 U5655 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[22]), .A1(kme_internal_out[51]), .Z(n2537));
Q_MX02 U5656 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[21]), .A1(kme_internal_out[50]), .Z(n2538));
Q_MX02 U5657 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[20]), .A1(kme_internal_out[49]), .Z(n2539));
Q_MX02 U5658 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[19]), .A1(kme_internal_out[48]), .Z(n2540));
Q_MX02 U5659 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[18]), .A1(kme_internal_out[47]), .Z(n2541));
Q_MX02 U5660 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[17]), .A1(kme_internal_out[46]), .Z(n2542));
Q_MX02 U5661 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[16]), .A1(kme_internal_out[45]), .Z(n2543));
Q_MX02 U5662 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[15]), .A1(kme_internal_out[44]), .Z(n2544));
Q_MX02 U5663 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[14]), .A1(kme_internal_out[43]), .Z(n2545));
Q_MX02 U5664 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[13]), .A1(kme_internal_out[42]), .Z(n2546));
Q_MX02 U5665 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[12]), .A1(kme_internal_out[41]), .Z(n2547));
Q_MX02 U5666 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[11]), .A1(kme_internal_out[40]), .Z(n2548));
Q_MX02 U5667 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[10]), .A1(kme_internal_out[39]), .Z(n2549));
Q_MX02 U5668 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[9]), .A1(kme_internal_out[38]), .Z(n2550));
Q_MX02 U5669 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[8]), .A1(kme_internal_out[37]), .Z(n2551));
Q_MX02 U5670 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[7]), .A1(kme_internal_out[36]), .Z(n2552));
Q_MX02 U5671 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[6]), .A1(kme_internal_out[35]), .Z(n2553));
Q_MX02 U5672 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[5]), .A1(kme_internal_out[34]), .Z(n2554));
Q_MX02 U5673 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[4]), .A1(kme_internal_out[33]), .Z(n2555));
Q_MX02 U5674 ( .S(kme_internal_out[69]), .A0(gcm_dak_cmd_in[3]), .A1(kme_internal_out[32]), .Z(n2556));
Q_MX02 U5675 ( .S(kme_internal_out[69]), .A0(kme_internal_out[63]), .A1(gcm_dak_cmd_in[98]), .Z(n2557));
Q_MX02 U5676 ( .S(kme_internal_out[69]), .A0(kme_internal_out[62]), .A1(gcm_dak_cmd_in[97]), .Z(n2558));
Q_MX02 U5677 ( .S(kme_internal_out[69]), .A0(kme_internal_out[61]), .A1(gcm_dak_cmd_in[96]), .Z(n2559));
Q_MX02 U5678 ( .S(kme_internal_out[69]), .A0(kme_internal_out[60]), .A1(gcm_dak_cmd_in[95]), .Z(n2560));
Q_MX02 U5679 ( .S(kme_internal_out[69]), .A0(kme_internal_out[59]), .A1(gcm_dak_cmd_in[94]), .Z(n2561));
Q_MX02 U5680 ( .S(kme_internal_out[69]), .A0(kme_internal_out[58]), .A1(gcm_dak_cmd_in[93]), .Z(n2562));
Q_MX02 U5681 ( .S(kme_internal_out[69]), .A0(kme_internal_out[57]), .A1(gcm_dak_cmd_in[92]), .Z(n2563));
Q_MX02 U5682 ( .S(kme_internal_out[69]), .A0(kme_internal_out[56]), .A1(gcm_dak_cmd_in[91]), .Z(n2564));
Q_MX02 U5683 ( .S(kme_internal_out[69]), .A0(kme_internal_out[55]), .A1(gcm_dak_cmd_in[90]), .Z(n2565));
Q_MX02 U5684 ( .S(kme_internal_out[69]), .A0(kme_internal_out[54]), .A1(gcm_dak_cmd_in[89]), .Z(n2566));
Q_MX02 U5685 ( .S(kme_internal_out[69]), .A0(kme_internal_out[53]), .A1(gcm_dak_cmd_in[88]), .Z(n2567));
Q_MX02 U5686 ( .S(kme_internal_out[69]), .A0(kme_internal_out[52]), .A1(gcm_dak_cmd_in[87]), .Z(n2568));
Q_MX02 U5687 ( .S(kme_internal_out[69]), .A0(kme_internal_out[51]), .A1(gcm_dak_cmd_in[86]), .Z(n2569));
Q_MX02 U5688 ( .S(kme_internal_out[69]), .A0(kme_internal_out[50]), .A1(gcm_dak_cmd_in[85]), .Z(n2570));
Q_MX02 U5689 ( .S(kme_internal_out[69]), .A0(kme_internal_out[49]), .A1(gcm_dak_cmd_in[84]), .Z(n2571));
Q_MX02 U5690 ( .S(kme_internal_out[69]), .A0(kme_internal_out[48]), .A1(gcm_dak_cmd_in[83]), .Z(n2572));
Q_MX02 U5691 ( .S(kme_internal_out[69]), .A0(kme_internal_out[47]), .A1(gcm_dak_cmd_in[82]), .Z(n2573));
Q_MX02 U5692 ( .S(kme_internal_out[69]), .A0(kme_internal_out[46]), .A1(gcm_dak_cmd_in[81]), .Z(n2574));
Q_MX02 U5693 ( .S(kme_internal_out[69]), .A0(kme_internal_out[45]), .A1(gcm_dak_cmd_in[80]), .Z(n2575));
Q_MX02 U5694 ( .S(kme_internal_out[69]), .A0(kme_internal_out[44]), .A1(gcm_dak_cmd_in[79]), .Z(n2576));
Q_MX02 U5695 ( .S(kme_internal_out[69]), .A0(kme_internal_out[43]), .A1(gcm_dak_cmd_in[78]), .Z(n2577));
Q_MX02 U5696 ( .S(kme_internal_out[69]), .A0(kme_internal_out[42]), .A1(gcm_dak_cmd_in[77]), .Z(n2578));
Q_MX02 U5697 ( .S(kme_internal_out[69]), .A0(kme_internal_out[41]), .A1(gcm_dak_cmd_in[76]), .Z(n2579));
Q_MX02 U5698 ( .S(kme_internal_out[69]), .A0(kme_internal_out[40]), .A1(gcm_dak_cmd_in[75]), .Z(n2580));
Q_MX02 U5699 ( .S(kme_internal_out[69]), .A0(kme_internal_out[39]), .A1(gcm_dak_cmd_in[74]), .Z(n2581));
Q_MX02 U5700 ( .S(kme_internal_out[69]), .A0(kme_internal_out[38]), .A1(gcm_dak_cmd_in[73]), .Z(n2582));
Q_MX02 U5701 ( .S(kme_internal_out[69]), .A0(kme_internal_out[37]), .A1(gcm_dak_cmd_in[72]), .Z(n2583));
Q_MX02 U5702 ( .S(kme_internal_out[69]), .A0(kme_internal_out[36]), .A1(gcm_dak_cmd_in[71]), .Z(n2584));
Q_MX02 U5703 ( .S(kme_internal_out[69]), .A0(kme_internal_out[35]), .A1(gcm_dak_cmd_in[70]), .Z(n2585));
Q_MX02 U5704 ( .S(kme_internal_out[69]), .A0(kme_internal_out[34]), .A1(gcm_dak_cmd_in[69]), .Z(n2586));
Q_MX02 U5705 ( .S(kme_internal_out[69]), .A0(kme_internal_out[33]), .A1(gcm_dak_cmd_in[68]), .Z(n2587));
Q_MX02 U5706 ( .S(kme_internal_out[69]), .A0(kme_internal_out[32]), .A1(gcm_dak_cmd_in[67]), .Z(n2588));
Q_MX02 U5707 ( .S(kme_internal_out[69]), .A0(kme_internal_out[31]), .A1(gcm_dak_cmd_in[66]), .Z(n2589));
Q_MX02 U5708 ( .S(kme_internal_out[69]), .A0(kme_internal_out[30]), .A1(gcm_dak_cmd_in[65]), .Z(n2590));
Q_MX02 U5709 ( .S(kme_internal_out[69]), .A0(kme_internal_out[29]), .A1(gcm_dak_cmd_in[64]), .Z(n2591));
Q_MX02 U5710 ( .S(kme_internal_out[69]), .A0(kme_internal_out[28]), .A1(gcm_dak_cmd_in[63]), .Z(n2592));
Q_MX02 U5711 ( .S(kme_internal_out[69]), .A0(kme_internal_out[27]), .A1(gcm_dak_cmd_in[62]), .Z(n2593));
Q_MX02 U5712 ( .S(kme_internal_out[69]), .A0(kme_internal_out[26]), .A1(gcm_dak_cmd_in[61]), .Z(n2594));
Q_MX02 U5713 ( .S(kme_internal_out[69]), .A0(kme_internal_out[25]), .A1(gcm_dak_cmd_in[60]), .Z(n2595));
Q_MX02 U5714 ( .S(kme_internal_out[69]), .A0(kme_internal_out[24]), .A1(gcm_dak_cmd_in[59]), .Z(n2596));
Q_MX02 U5715 ( .S(kme_internal_out[69]), .A0(kme_internal_out[23]), .A1(gcm_dak_cmd_in[58]), .Z(n2597));
Q_MX02 U5716 ( .S(kme_internal_out[69]), .A0(kme_internal_out[22]), .A1(gcm_dak_cmd_in[57]), .Z(n2598));
Q_MX02 U5717 ( .S(kme_internal_out[69]), .A0(kme_internal_out[21]), .A1(gcm_dak_cmd_in[56]), .Z(n2599));
Q_MX02 U5718 ( .S(kme_internal_out[69]), .A0(kme_internal_out[20]), .A1(gcm_dak_cmd_in[55]), .Z(n2600));
Q_MX02 U5719 ( .S(kme_internal_out[69]), .A0(kme_internal_out[19]), .A1(gcm_dak_cmd_in[54]), .Z(n2601));
Q_MX02 U5720 ( .S(kme_internal_out[69]), .A0(kme_internal_out[18]), .A1(gcm_dak_cmd_in[53]), .Z(n2602));
Q_MX02 U5721 ( .S(kme_internal_out[69]), .A0(kme_internal_out[17]), .A1(gcm_dak_cmd_in[52]), .Z(n2603));
Q_MX02 U5722 ( .S(kme_internal_out[69]), .A0(kme_internal_out[16]), .A1(gcm_dak_cmd_in[51]), .Z(n2604));
Q_MX02 U5723 ( .S(kme_internal_out[69]), .A0(kme_internal_out[15]), .A1(gcm_dak_cmd_in[50]), .Z(n2605));
Q_MX02 U5724 ( .S(kme_internal_out[69]), .A0(kme_internal_out[14]), .A1(gcm_dak_cmd_in[49]), .Z(n2606));
Q_MX02 U5725 ( .S(kme_internal_out[69]), .A0(kme_internal_out[13]), .A1(gcm_dak_cmd_in[48]), .Z(n2607));
Q_MX02 U5726 ( .S(kme_internal_out[69]), .A0(kme_internal_out[12]), .A1(gcm_dak_cmd_in[47]), .Z(n2608));
Q_MX02 U5727 ( .S(kme_internal_out[69]), .A0(kme_internal_out[11]), .A1(gcm_dak_cmd_in[46]), .Z(n2609));
Q_MX02 U5728 ( .S(kme_internal_out[69]), .A0(kme_internal_out[10]), .A1(gcm_dak_cmd_in[45]), .Z(n2610));
Q_MX02 U5729 ( .S(kme_internal_out[69]), .A0(kme_internal_out[9]), .A1(gcm_dak_cmd_in[44]), .Z(n2611));
Q_MX02 U5730 ( .S(kme_internal_out[69]), .A0(kme_internal_out[8]), .A1(gcm_dak_cmd_in[43]), .Z(n2612));
Q_MX02 U5731 ( .S(kme_internal_out[69]), .A0(kme_internal_out[7]), .A1(gcm_dak_cmd_in[42]), .Z(n2613));
Q_MX02 U5732 ( .S(kme_internal_out[69]), .A0(kme_internal_out[6]), .A1(gcm_dak_cmd_in[41]), .Z(n2614));
Q_MX02 U5733 ( .S(kme_internal_out[69]), .A0(kme_internal_out[5]), .A1(gcm_dak_cmd_in[40]), .Z(n2615));
Q_MX02 U5734 ( .S(kme_internal_out[69]), .A0(kme_internal_out[4]), .A1(gcm_dak_cmd_in[39]), .Z(n2616));
Q_MX02 U5735 ( .S(kme_internal_out[69]), .A0(kme_internal_out[3]), .A1(gcm_dak_cmd_in[38]), .Z(n2617));
Q_MX02 U5736 ( .S(kme_internal_out[69]), .A0(kme_internal_out[2]), .A1(gcm_dak_cmd_in[37]), .Z(n2618));
Q_MX02 U5737 ( .S(kme_internal_out[69]), .A0(kme_internal_out[1]), .A1(gcm_dak_cmd_in[36]), .Z(n2619));
Q_MX02 U5738 ( .S(kme_internal_out[69]), .A0(kme_internal_out[0]), .A1(gcm_dak_cmd_in[35]), .Z(n2620));
Q_MX02 U5739 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[34]), .A1(kme_internal_out[63]), .Z(n2621));
Q_MX02 U5740 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[33]), .A1(kme_internal_out[62]), .Z(n2622));
Q_MX02 U5741 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[32]), .A1(kme_internal_out[61]), .Z(n2623));
Q_MX02 U5742 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[31]), .A1(kme_internal_out[60]), .Z(n2624));
Q_MX02 U5743 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[30]), .A1(kme_internal_out[59]), .Z(n2625));
Q_MX02 U5744 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[29]), .A1(kme_internal_out[58]), .Z(n2626));
Q_MX02 U5745 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[28]), .A1(kme_internal_out[57]), .Z(n2627));
Q_MX02 U5746 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[27]), .A1(kme_internal_out[56]), .Z(n2628));
Q_MX02 U5747 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[26]), .A1(kme_internal_out[55]), .Z(n2629));
Q_MX02 U5748 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[25]), .A1(kme_internal_out[54]), .Z(n2630));
Q_MX02 U5749 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[24]), .A1(kme_internal_out[53]), .Z(n2631));
Q_MX02 U5750 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[23]), .A1(kme_internal_out[52]), .Z(n2632));
Q_MX02 U5751 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[22]), .A1(kme_internal_out[51]), .Z(n2633));
Q_MX02 U5752 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[21]), .A1(kme_internal_out[50]), .Z(n2634));
Q_MX02 U5753 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[20]), .A1(kme_internal_out[49]), .Z(n2635));
Q_MX02 U5754 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[19]), .A1(kme_internal_out[48]), .Z(n2636));
Q_MX02 U5755 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[18]), .A1(kme_internal_out[47]), .Z(n2637));
Q_MX02 U5756 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[17]), .A1(kme_internal_out[46]), .Z(n2638));
Q_MX02 U5757 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[16]), .A1(kme_internal_out[45]), .Z(n2639));
Q_MX02 U5758 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[15]), .A1(kme_internal_out[44]), .Z(n2640));
Q_MX02 U5759 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[14]), .A1(kme_internal_out[43]), .Z(n2641));
Q_MX02 U5760 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[13]), .A1(kme_internal_out[42]), .Z(n2642));
Q_MX02 U5761 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[12]), .A1(kme_internal_out[41]), .Z(n2643));
Q_MX02 U5762 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[11]), .A1(kme_internal_out[40]), .Z(n2644));
Q_MX02 U5763 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[10]), .A1(kme_internal_out[39]), .Z(n2645));
Q_MX02 U5764 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[9]), .A1(kme_internal_out[38]), .Z(n2646));
Q_MX02 U5765 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[8]), .A1(kme_internal_out[37]), .Z(n2647));
Q_MX02 U5766 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[7]), .A1(kme_internal_out[36]), .Z(n2648));
Q_MX02 U5767 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[6]), .A1(kme_internal_out[35]), .Z(n2649));
Q_MX02 U5768 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[5]), .A1(kme_internal_out[34]), .Z(n2650));
Q_MX02 U5769 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[4]), .A1(kme_internal_out[33]), .Z(n2651));
Q_MX02 U5770 ( .S(kme_internal_out[69]), .A0(gcm_dek_cmd_in[3]), .A1(kme_internal_out[32]), .Z(n2652));
Q_MX02 U5771 ( .S(kme_internal_out[69]), .A0(kme_internal_out[63]), .A1(gcm_dek_cmd_in[98]), .Z(n2653));
Q_MX02 U5772 ( .S(kme_internal_out[69]), .A0(kme_internal_out[62]), .A1(gcm_dek_cmd_in[97]), .Z(n2654));
Q_MX02 U5773 ( .S(kme_internal_out[69]), .A0(kme_internal_out[61]), .A1(gcm_dek_cmd_in[96]), .Z(n2655));
Q_MX02 U5774 ( .S(kme_internal_out[69]), .A0(kme_internal_out[60]), .A1(gcm_dek_cmd_in[95]), .Z(n2656));
Q_MX02 U5775 ( .S(kme_internal_out[69]), .A0(kme_internal_out[59]), .A1(gcm_dek_cmd_in[94]), .Z(n2657));
Q_MX02 U5776 ( .S(kme_internal_out[69]), .A0(kme_internal_out[58]), .A1(gcm_dek_cmd_in[93]), .Z(n2658));
Q_MX02 U5777 ( .S(kme_internal_out[69]), .A0(kme_internal_out[57]), .A1(gcm_dek_cmd_in[92]), .Z(n2659));
Q_MX02 U5778 ( .S(kme_internal_out[69]), .A0(kme_internal_out[56]), .A1(gcm_dek_cmd_in[91]), .Z(n2660));
Q_MX02 U5779 ( .S(kme_internal_out[69]), .A0(kme_internal_out[55]), .A1(gcm_dek_cmd_in[90]), .Z(n2661));
Q_MX02 U5780 ( .S(kme_internal_out[69]), .A0(kme_internal_out[54]), .A1(gcm_dek_cmd_in[89]), .Z(n2662));
Q_MX02 U5781 ( .S(kme_internal_out[69]), .A0(kme_internal_out[53]), .A1(gcm_dek_cmd_in[88]), .Z(n2663));
Q_MX02 U5782 ( .S(kme_internal_out[69]), .A0(kme_internal_out[52]), .A1(gcm_dek_cmd_in[87]), .Z(n2664));
Q_MX02 U5783 ( .S(kme_internal_out[69]), .A0(kme_internal_out[51]), .A1(gcm_dek_cmd_in[86]), .Z(n2665));
Q_MX02 U5784 ( .S(kme_internal_out[69]), .A0(kme_internal_out[50]), .A1(gcm_dek_cmd_in[85]), .Z(n2666));
Q_MX02 U5785 ( .S(kme_internal_out[69]), .A0(kme_internal_out[49]), .A1(gcm_dek_cmd_in[84]), .Z(n2667));
Q_MX02 U5786 ( .S(kme_internal_out[69]), .A0(kme_internal_out[48]), .A1(gcm_dek_cmd_in[83]), .Z(n2668));
Q_MX02 U5787 ( .S(kme_internal_out[69]), .A0(kme_internal_out[47]), .A1(gcm_dek_cmd_in[82]), .Z(n2669));
Q_MX02 U5788 ( .S(kme_internal_out[69]), .A0(kme_internal_out[46]), .A1(gcm_dek_cmd_in[81]), .Z(n2670));
Q_MX02 U5789 ( .S(kme_internal_out[69]), .A0(kme_internal_out[45]), .A1(gcm_dek_cmd_in[80]), .Z(n2671));
Q_MX02 U5790 ( .S(kme_internal_out[69]), .A0(kme_internal_out[44]), .A1(gcm_dek_cmd_in[79]), .Z(n2672));
Q_MX02 U5791 ( .S(kme_internal_out[69]), .A0(kme_internal_out[43]), .A1(gcm_dek_cmd_in[78]), .Z(n2673));
Q_MX02 U5792 ( .S(kme_internal_out[69]), .A0(kme_internal_out[42]), .A1(gcm_dek_cmd_in[77]), .Z(n2674));
Q_MX02 U5793 ( .S(kme_internal_out[69]), .A0(kme_internal_out[41]), .A1(gcm_dek_cmd_in[76]), .Z(n2675));
Q_MX02 U5794 ( .S(kme_internal_out[69]), .A0(kme_internal_out[40]), .A1(gcm_dek_cmd_in[75]), .Z(n2676));
Q_MX02 U5795 ( .S(kme_internal_out[69]), .A0(kme_internal_out[39]), .A1(gcm_dek_cmd_in[74]), .Z(n2677));
Q_MX02 U5796 ( .S(kme_internal_out[69]), .A0(kme_internal_out[38]), .A1(gcm_dek_cmd_in[73]), .Z(n2678));
Q_MX02 U5797 ( .S(kme_internal_out[69]), .A0(kme_internal_out[37]), .A1(gcm_dek_cmd_in[72]), .Z(n2679));
Q_MX02 U5798 ( .S(kme_internal_out[69]), .A0(kme_internal_out[36]), .A1(gcm_dek_cmd_in[71]), .Z(n2680));
Q_MX02 U5799 ( .S(kme_internal_out[69]), .A0(kme_internal_out[35]), .A1(gcm_dek_cmd_in[70]), .Z(n2681));
Q_MX02 U5800 ( .S(kme_internal_out[69]), .A0(kme_internal_out[34]), .A1(gcm_dek_cmd_in[69]), .Z(n2682));
Q_MX02 U5801 ( .S(kme_internal_out[69]), .A0(kme_internal_out[33]), .A1(gcm_dek_cmd_in[68]), .Z(n2683));
Q_MX02 U5802 ( .S(kme_internal_out[69]), .A0(kme_internal_out[32]), .A1(gcm_dek_cmd_in[67]), .Z(n2684));
Q_MX02 U5803 ( .S(kme_internal_out[69]), .A0(kme_internal_out[31]), .A1(gcm_dek_cmd_in[66]), .Z(n2685));
Q_MX02 U5804 ( .S(kme_internal_out[69]), .A0(kme_internal_out[30]), .A1(gcm_dek_cmd_in[65]), .Z(n2686));
Q_MX02 U5805 ( .S(kme_internal_out[69]), .A0(kme_internal_out[29]), .A1(gcm_dek_cmd_in[64]), .Z(n2687));
Q_MX02 U5806 ( .S(kme_internal_out[69]), .A0(kme_internal_out[28]), .A1(gcm_dek_cmd_in[63]), .Z(n2688));
Q_MX02 U5807 ( .S(kme_internal_out[69]), .A0(kme_internal_out[27]), .A1(gcm_dek_cmd_in[62]), .Z(n2689));
Q_MX02 U5808 ( .S(kme_internal_out[69]), .A0(kme_internal_out[26]), .A1(gcm_dek_cmd_in[61]), .Z(n2690));
Q_MX02 U5809 ( .S(kme_internal_out[69]), .A0(kme_internal_out[25]), .A1(gcm_dek_cmd_in[60]), .Z(n2691));
Q_MX02 U5810 ( .S(kme_internal_out[69]), .A0(kme_internal_out[24]), .A1(gcm_dek_cmd_in[59]), .Z(n2692));
Q_MX02 U5811 ( .S(kme_internal_out[69]), .A0(kme_internal_out[23]), .A1(gcm_dek_cmd_in[58]), .Z(n2693));
Q_MX02 U5812 ( .S(kme_internal_out[69]), .A0(kme_internal_out[22]), .A1(gcm_dek_cmd_in[57]), .Z(n2694));
Q_MX02 U5813 ( .S(kme_internal_out[69]), .A0(kme_internal_out[21]), .A1(gcm_dek_cmd_in[56]), .Z(n2695));
Q_MX02 U5814 ( .S(kme_internal_out[69]), .A0(kme_internal_out[20]), .A1(gcm_dek_cmd_in[55]), .Z(n2696));
Q_MX02 U5815 ( .S(kme_internal_out[69]), .A0(kme_internal_out[19]), .A1(gcm_dek_cmd_in[54]), .Z(n2697));
Q_MX02 U5816 ( .S(kme_internal_out[69]), .A0(kme_internal_out[18]), .A1(gcm_dek_cmd_in[53]), .Z(n2698));
Q_MX02 U5817 ( .S(kme_internal_out[69]), .A0(kme_internal_out[17]), .A1(gcm_dek_cmd_in[52]), .Z(n2699));
Q_MX02 U5818 ( .S(kme_internal_out[69]), .A0(kme_internal_out[16]), .A1(gcm_dek_cmd_in[51]), .Z(n2700));
Q_MX02 U5819 ( .S(kme_internal_out[69]), .A0(kme_internal_out[15]), .A1(gcm_dek_cmd_in[50]), .Z(n2701));
Q_MX02 U5820 ( .S(kme_internal_out[69]), .A0(kme_internal_out[14]), .A1(gcm_dek_cmd_in[49]), .Z(n2702));
Q_MX02 U5821 ( .S(kme_internal_out[69]), .A0(kme_internal_out[13]), .A1(gcm_dek_cmd_in[48]), .Z(n2703));
Q_MX02 U5822 ( .S(kme_internal_out[69]), .A0(kme_internal_out[12]), .A1(gcm_dek_cmd_in[47]), .Z(n2704));
Q_MX02 U5823 ( .S(kme_internal_out[69]), .A0(kme_internal_out[11]), .A1(gcm_dek_cmd_in[46]), .Z(n2705));
Q_MX02 U5824 ( .S(kme_internal_out[69]), .A0(kme_internal_out[10]), .A1(gcm_dek_cmd_in[45]), .Z(n2706));
Q_MX02 U5825 ( .S(kme_internal_out[69]), .A0(kme_internal_out[9]), .A1(gcm_dek_cmd_in[44]), .Z(n2707));
Q_MX02 U5826 ( .S(kme_internal_out[69]), .A0(kme_internal_out[8]), .A1(gcm_dek_cmd_in[43]), .Z(n2708));
Q_MX02 U5827 ( .S(kme_internal_out[69]), .A0(kme_internal_out[7]), .A1(gcm_dek_cmd_in[42]), .Z(n2709));
Q_MX02 U5828 ( .S(kme_internal_out[69]), .A0(kme_internal_out[6]), .A1(gcm_dek_cmd_in[41]), .Z(n2710));
Q_MX02 U5829 ( .S(kme_internal_out[69]), .A0(kme_internal_out[5]), .A1(gcm_dek_cmd_in[40]), .Z(n2711));
Q_MX02 U5830 ( .S(kme_internal_out[69]), .A0(kme_internal_out[4]), .A1(gcm_dek_cmd_in[39]), .Z(n2712));
Q_MX02 U5831 ( .S(kme_internal_out[69]), .A0(kme_internal_out[3]), .A1(gcm_dek_cmd_in[38]), .Z(n2713));
Q_MX02 U5832 ( .S(kme_internal_out[69]), .A0(kme_internal_out[2]), .A1(gcm_dek_cmd_in[37]), .Z(n2714));
Q_MX02 U5833 ( .S(kme_internal_out[69]), .A0(kme_internal_out[1]), .A1(gcm_dek_cmd_in[36]), .Z(n2715));
Q_MX02 U5834 ( .S(kme_internal_out[69]), .A0(kme_internal_out[0]), .A1(gcm_dek_cmd_in[35]), .Z(n2716));
Q_AN02 U5835 ( .A0(kme_internal_out_ack), .A1(n2729), .Z(keyfilter_cmd_in_valid));
Q_AN02 U5836 ( .A0(n139), .A1(kme_internal_out_valid), .Z(kme_internal_out_ack));
Q_INV U5837 ( .A(kme_internal_out[31]), .Z(n2717));
Q_INV U5838 ( .A(kme_internal_out[14]), .Z(n2718));
Q_AO21 U5839 ( .A0(n2719), .A1(upsizer_inspector_stall), .B0(n19), .Z(n131));
Q_AN02 U5840 ( .A0(kme_internal_out[64]), .A1(n2720), .Z(n2719));
Q_AN03 U5841 ( .A0(kme_internal_out[67]), .A1(n14), .A2(n49), .Z(n2720));
Q_OA21 U5842 ( .A0(n2721), .A1(n2723), .B0(upsizer_inspector_stall), .Z(n132));
Q_AN02 U5843 ( .A0(n2731), .A1(n2722), .Z(n2721));
Q_AN03 U5844 ( .A0(kme_internal_out[67]), .A1(n14), .A2(kme_internal_out[65]), .Z(n2722));
Q_AN02 U5845 ( .A0(kme_internal_out[64]), .A1(n2724), .Z(n2723));
Q_AN03 U5846 ( .A0(kme_internal_out[67]), .A1(kme_internal_out[66]), .A2(n49), .Z(n2724));
Q_AN03 U5847 ( .A0(n2725), .A1(kme_internal_out[69]), .A2(gcm_cmd_in_stall), .Z(n17));
Q_NR02 U5848 ( .A0(kme_internal_out[64]), .A1(n2853), .Z(n2725));
Q_AN03 U5849 ( .A0(n2726), .A1(kme_internal_out[69]), .A2(gcm_cmd_in_stall), .Z(n18));
Q_AN02 U5850 ( .A0(n2731), .A1(n2724), .Z(n2726));
Q_AN03 U5851 ( .A0(n15), .A1(kme_internal_out[69]), .A2(gcm_tag_data_in_stall), .Z(n19));
Q_AN02 U5852 ( .A0(kme_internal_out[64]), .A1(n2722), .Z(n15));
Q_AN03 U5853 ( .A0(n16), .A1(kme_internal_out[69]), .A2(gcm_tag_data_in_stall), .Z(n20));
Q_AN02 U5854 ( .A0(n2731), .A1(n2727), .Z(n16));
Q_AN03 U5855 ( .A0(kme_internal_out[67]), .A1(kme_internal_out[66]), .A2(kme_internal_out[65]), .Z(n2727));
Q_AO21 U5856 ( .A0(n2728), .A1(kdf_cmd_in_stall), .B0(n20), .Z(n134));
Q_AO21 U5857 ( .A0(n2728), .A1(keyfilter_cmd_in_stall), .B0(n21), .Z(n130));
Q_AN02 U5858 ( .A0(n2729), .A1(kme_internal_out[69]), .Z(n2728));
Q_NR02 U5859 ( .A0(n2731), .A1(n2730), .Z(n2729));
Q_OR03 U5860 ( .A0(kme_internal_out[67]), .A1(kme_internal_out[66]), .A2(kme_internal_out[65]), .Z(n2730));
Q_INV U5861 ( .A(kme_internal_out[64]), .Z(n2731));
Q_AO21 U5862 ( .A0(n12), .A1(kdfstream_cmd_in_stall), .B0(_zy_sva_b8_t), .Z(n135));
Q_AN03 U5863 ( .A0(n2732), .A1(kme_internal_out[69]), .A2(tlv_sb_data_in_stall), .Z(n21));
Q_NR02 U5864 ( .A0(kme_internal_out[64]), .A1(n2730), .Z(n2732));
Q_AN03 U5865 ( .A0(n2733), .A1(kme_internal_out_valid), .A2(tlv_sb_data_in_stall), .Z(_zy_sva_b8_t));
Q_AN02 U5866 ( .A0(kme_internal_out[64]), .A1(n2734), .Z(n2733));
Q_AN03 U5867 ( .A0(n2735), .A1(n14), .A2(kme_internal_out[65]), .Z(n2734));
Q_INV U5868 ( .A(kme_internal_out[67]), .Z(n2735));
Q_AN03 U5869 ( .A0(n2736), .A1(kme_internal_out_valid), .A2(tlv_sb_data_in_stall), .Z(n22));
Q_NR02 U5870 ( .A0(kme_internal_out[64]), .A1(n2852), .Z(n2736));
Q_AN03 U5871 ( .A0(n2737), .A1(kme_internal_out_valid), .A2(tlv_sb_data_in_stall), .Z(n23));
Q_AN02 U5872 ( .A0(kme_internal_out[64]), .A1(n2727), .Z(n2737));
Q_INV U5873 ( .A(kme_internal_out[62]), .Z(n2753));
Q_INV U5874 ( .A(kme_internal_out[61]), .Z(n2752));
Q_NR02 U5875 ( .A0(kme_internal_out[62]), .A1(kme_internal_out[61]), .Z(n2745));
Q_AN02 U5876 ( .A0(n2738), .A1(n2745), .Z(n2750));
Q_AO21 U5877 ( .A0(n2750), .A1(kme_internal_out[32]), .B0(n2760), .Z(n2746));
Q_AN02 U5878 ( .A0(n2737), .A1(rst_corrupt_crc32), .Z(n2760));
Q_AN02 U5879 ( .A0(kme_internal_out_ack), .A1(n2746), .Z(n2739));
Q_AN03 U5880 ( .A0(n2738), .A1(n2752), .A2(kme_internal_out[32]), .Z(n2748));
Q_AN02 U5881 ( .A0(n2738), .A1(n2753), .Z(n2747));
Q_AO21 U5882 ( .A0(n2747), .A1(kme_internal_out[32]), .B0(n2760), .Z(n2749));
Q_OA21 U5883 ( .A0(n2749), .A1(n2748), .B0(kme_internal_out_ack), .Z(n2740));
Q_INV U5884 ( .A(kme_internal_out[32]), .Z(n2754));
Q_AO21 U5885 ( .A0(n2750), .A1(n2754), .B0(n2758), .Z(n2751));
Q_AN02 U5886 ( .A0(n2737), .A1(rst_corrupt_kme_error_bit_0), .Z(n2758));
Q_AN02 U5887 ( .A0(kme_internal_out_ack), .A1(n2751), .Z(n2741));
Q_ND02 U5888 ( .A0(kme_internal_out[62]), .A1(kme_internal_out[61]), .Z(n2755));
Q_AN03 U5889 ( .A0(n2738), .A1(n2754), .A2(n2755), .Z(n2756));
Q_OA21 U5890 ( .A0(n2756), .A1(n2758), .B0(kme_internal_out_ack), .Z(n2742));
Q_NR02 U5891 ( .A0(kme_internal_out[62]), .A1(n2758), .Z(n2757));
Q_INV U5892 ( .A(n2758), .Z(n2743));
Q_NR02 U5893 ( .A0(n2760), .A1(kme_internal_out[62]), .Z(n2759));
Q_INV U5894 ( .A(n2760), .Z(n2744));
Q_AN02 U5895 ( .A0(n2762), .A1(n2761), .Z(n2738));
Q_AN03 U5896 ( .A0(kme_internal_out[55]), .A1(n2764), .A2(n2729), .Z(n2761));
Q_AN03 U5897 ( .A0(kme_internal_out[57]), .A1(kme_internal_out[56]), .A2(n2763), .Z(n2762));
Q_AN03 U5898 ( .A0(kme_internal_out[60]), .A1(kme_internal_out[59]), .A2(kme_internal_out[58]), .Z(n2763));
Q_INV U5899 ( .A(kme_internal_out[63]), .Z(n2764));
Q_FDP1 \stream_cmd_in_REG[262] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[262]), .Q(stream_cmd_in[262]), .QN(n55));
Q_FDP1 \stream_cmd_in_REG[261] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[261]), .Q(stream_cmd_in[261]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[260] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[260]), .Q(stream_cmd_in[260]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[259] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[259]), .Q(stream_cmd_in[259]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[258] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[258]), .Q(stream_cmd_in[258]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[257] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[257]), .Q(stream_cmd_in[257]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[256] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[256]), .Q(stream_cmd_in[256]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[255] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[255]), .Q(stream_cmd_in[255]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[254] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[254]), .Q(stream_cmd_in[254]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[253] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[253]), .Q(stream_cmd_in[253]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[252] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[252]), .Q(stream_cmd_in[252]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[251] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[251]), .Q(stream_cmd_in[251]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[250] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[250]), .Q(stream_cmd_in[250]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[249] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[249]), .Q(stream_cmd_in[249]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[248] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[248]), .Q(stream_cmd_in[248]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[247] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[247]), .Q(stream_cmd_in[247]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[246] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[246]), .Q(stream_cmd_in[246]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[245] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[245]), .Q(stream_cmd_in[245]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[244] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[244]), .Q(stream_cmd_in[244]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[243] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[243]), .Q(stream_cmd_in[243]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[242] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[242]), .Q(stream_cmd_in[242]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[241] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[241]), .Q(stream_cmd_in[241]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[240] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[240]), .Q(stream_cmd_in[240]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[239] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[239]), .Q(stream_cmd_in[239]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[238] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[238]), .Q(stream_cmd_in[238]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[237] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[237]), .Q(stream_cmd_in[237]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[236] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[236]), .Q(stream_cmd_in[236]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[235] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[235]), .Q(stream_cmd_in[235]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[234] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[234]), .Q(stream_cmd_in[234]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[233] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[233]), .Q(stream_cmd_in[233]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[232] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[232]), .Q(stream_cmd_in[232]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[231] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[231]), .Q(stream_cmd_in[231]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[230] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[230]), .Q(stream_cmd_in[230]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[229] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[229]), .Q(stream_cmd_in[229]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[228] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[228]), .Q(stream_cmd_in[228]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[227] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[227]), .Q(stream_cmd_in[227]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[226] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[226]), .Q(stream_cmd_in[226]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[225] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[225]), .Q(stream_cmd_in[225]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[224] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[224]), .Q(stream_cmd_in[224]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[223] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[223]), .Q(stream_cmd_in[223]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[222] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[222]), .Q(stream_cmd_in[222]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[221] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[221]), .Q(stream_cmd_in[221]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[220] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[220]), .Q(stream_cmd_in[220]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[219] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[219]), .Q(stream_cmd_in[219]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[218] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[218]), .Q(stream_cmd_in[218]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[217] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[217]), .Q(stream_cmd_in[217]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[216] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[216]), .Q(stream_cmd_in[216]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[215] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[215]), .Q(stream_cmd_in[215]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[214] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[214]), .Q(stream_cmd_in[214]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[213] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[213]), .Q(stream_cmd_in[213]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[212] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[212]), .Q(stream_cmd_in[212]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[211] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[211]), .Q(stream_cmd_in[211]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[210] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[210]), .Q(stream_cmd_in[210]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[209] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[209]), .Q(stream_cmd_in[209]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[208] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[208]), .Q(stream_cmd_in[208]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[207] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[207]), .Q(stream_cmd_in[207]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[206] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[206]), .Q(stream_cmd_in[206]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[205] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[205]), .Q(stream_cmd_in[205]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[204] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[204]), .Q(stream_cmd_in[204]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[203] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[203]), .Q(stream_cmd_in[203]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[202] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[202]), .Q(stream_cmd_in[202]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[201] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[201]), .Q(stream_cmd_in[201]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[200] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[200]), .Q(stream_cmd_in[200]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[199] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[199]), .Q(stream_cmd_in[199]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[198] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[198]), .Q(stream_cmd_in[198]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[197] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[197]), .Q(stream_cmd_in[197]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[196] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[196]), .Q(stream_cmd_in[196]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[195] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[195]), .Q(stream_cmd_in[195]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[194] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[194]), .Q(stream_cmd_in[194]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[193] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[193]), .Q(stream_cmd_in[193]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[192] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[192]), .Q(stream_cmd_in[192]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[191] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[191]), .Q(stream_cmd_in[191]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[190] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[190]), .Q(stream_cmd_in[190]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[189] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[189]), .Q(stream_cmd_in[189]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[188] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[188]), .Q(stream_cmd_in[188]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[187] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[187]), .Q(stream_cmd_in[187]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[186] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[186]), .Q(stream_cmd_in[186]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[185] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[185]), .Q(stream_cmd_in[185]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[184] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[184]), .Q(stream_cmd_in[184]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[183] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[183]), .Q(stream_cmd_in[183]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[182] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[182]), .Q(stream_cmd_in[182]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[181] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[181]), .Q(stream_cmd_in[181]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[180] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[180]), .Q(stream_cmd_in[180]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[179] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[179]), .Q(stream_cmd_in[179]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[178] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[178]), .Q(stream_cmd_in[178]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[177] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[177]), .Q(stream_cmd_in[177]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[176] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[176]), .Q(stream_cmd_in[176]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[175] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[175]), .Q(stream_cmd_in[175]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[174] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[174]), .Q(stream_cmd_in[174]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[173] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[173]), .Q(stream_cmd_in[173]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[172] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[172]), .Q(stream_cmd_in[172]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[171] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[171]), .Q(stream_cmd_in[171]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[170] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[170]), .Q(stream_cmd_in[170]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[169] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[169]), .Q(stream_cmd_in[169]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[168] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[168]), .Q(stream_cmd_in[168]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[167] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[167]), .Q(stream_cmd_in[167]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[166] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[166]), .Q(stream_cmd_in[166]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[165] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[165]), .Q(stream_cmd_in[165]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[164] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[164]), .Q(stream_cmd_in[164]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[163] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[163]), .Q(stream_cmd_in[163]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[162] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[162]), .Q(stream_cmd_in[162]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[161] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[161]), .Q(stream_cmd_in[161]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[160] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[160]), .Q(stream_cmd_in[160]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[159] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[159]), .Q(stream_cmd_in[159]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[158] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[158]), .Q(stream_cmd_in[158]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[157] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[157]), .Q(stream_cmd_in[157]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[156] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[156]), .Q(stream_cmd_in[156]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[155] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[155]), .Q(stream_cmd_in[155]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[154] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[154]), .Q(stream_cmd_in[154]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[153] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[153]), .Q(stream_cmd_in[153]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[152] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[152]), .Q(stream_cmd_in[152]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[151] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[151]), .Q(stream_cmd_in[151]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[150] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[150]), .Q(stream_cmd_in[150]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[149] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[149]), .Q(stream_cmd_in[149]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[148] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[148]), .Q(stream_cmd_in[148]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[147] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[147]), .Q(stream_cmd_in[147]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[146] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[146]), .Q(stream_cmd_in[146]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[145] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[145]), .Q(stream_cmd_in[145]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[144] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[144]), .Q(stream_cmd_in[144]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[143] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[143]), .Q(stream_cmd_in[143]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[142] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[142]), .Q(stream_cmd_in[142]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[141] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[141]), .Q(stream_cmd_in[141]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[140] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[140]), .Q(stream_cmd_in[140]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[139] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[139]), .Q(stream_cmd_in[139]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[138] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[138]), .Q(stream_cmd_in[138]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[137] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[137]), .Q(stream_cmd_in[137]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[136] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[136]), .Q(stream_cmd_in[136]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[135] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[135]), .Q(stream_cmd_in[135]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[134] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[134]), .Q(stream_cmd_in[134]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[133] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[133]), .Q(stream_cmd_in[133]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[132] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[132]), .Q(stream_cmd_in[132]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[131] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[131]), .Q(stream_cmd_in[131]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[130] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[130]), .Q(stream_cmd_in[130]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[129] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[129]), .Q(stream_cmd_in[129]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[128] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[128]), .Q(stream_cmd_in[128]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[127] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[127]), .Q(stream_cmd_in[127]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[126] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[126]), .Q(stream_cmd_in[126]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[125] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[125]), .Q(stream_cmd_in[125]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[124] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[124]), .Q(stream_cmd_in[124]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[123] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[123]), .Q(stream_cmd_in[123]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[122] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[122]), .Q(stream_cmd_in[122]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[121] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[121]), .Q(stream_cmd_in[121]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[120] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[120]), .Q(stream_cmd_in[120]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[119] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[119]), .Q(stream_cmd_in[119]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[118] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[118]), .Q(stream_cmd_in[118]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[117] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[117]), .Q(stream_cmd_in[117]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[116] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[116]), .Q(stream_cmd_in[116]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[115] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[115]), .Q(stream_cmd_in[115]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[114] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[114]), .Q(stream_cmd_in[114]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[113] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[113]), .Q(stream_cmd_in[113]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[112] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[112]), .Q(stream_cmd_in[112]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[111] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[111]), .Q(stream_cmd_in[111]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[110] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[110]), .Q(stream_cmd_in[110]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[109] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[109]), .Q(stream_cmd_in[109]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[108] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[108]), .Q(stream_cmd_in[108]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[107] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[107]), .Q(stream_cmd_in[107]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[106] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[106]), .Q(stream_cmd_in[106]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[105] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[105]), .Q(stream_cmd_in[105]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[104] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[104]), .Q(stream_cmd_in[104]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[103] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[103]), .Q(stream_cmd_in[103]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[102] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[102]), .Q(stream_cmd_in[102]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[101] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[101]), .Q(stream_cmd_in[101]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[100] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[100]), .Q(stream_cmd_in[100]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[99] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[99]), .Q(stream_cmd_in[99]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[98] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[98]), .Q(stream_cmd_in[98]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[97] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[97]), .Q(stream_cmd_in[97]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[96] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[96]), .Q(stream_cmd_in[96]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[95] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[95]), .Q(stream_cmd_in[95]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[94] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[94]), .Q(stream_cmd_in[94]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[93] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[93]), .Q(stream_cmd_in[93]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[92] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[92]), .Q(stream_cmd_in[92]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[91] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[91]), .Q(stream_cmd_in[91]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[90] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[90]), .Q(stream_cmd_in[90]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[89] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[89]), .Q(stream_cmd_in[89]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[88] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[88]), .Q(stream_cmd_in[88]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[87] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[87]), .Q(stream_cmd_in[87]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[86] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[86]), .Q(stream_cmd_in[86]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[85] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[85]), .Q(stream_cmd_in[85]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[84] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[84]), .Q(stream_cmd_in[84]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[83] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[83]), .Q(stream_cmd_in[83]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[82] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[82]), .Q(stream_cmd_in[82]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[81] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[81]), .Q(stream_cmd_in[81]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[80] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[80]), .Q(stream_cmd_in[80]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[79] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[79]), .Q(stream_cmd_in[79]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[78] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[78]), .Q(stream_cmd_in[78]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[77] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[77]), .Q(stream_cmd_in[77]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[76] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[76]), .Q(stream_cmd_in[76]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[75] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[75]), .Q(stream_cmd_in[75]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[74] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[74]), .Q(stream_cmd_in[74]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[73] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[73]), .Q(stream_cmd_in[73]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[72] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[72]), .Q(stream_cmd_in[72]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[71] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[71]), .Q(stream_cmd_in[71]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[70] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[70]), .Q(stream_cmd_in[70]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[69] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[69]), .Q(stream_cmd_in[69]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[68] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[68]), .Q(stream_cmd_in[68]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[67] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[67]), .Q(stream_cmd_in[67]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[66] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[66]), .Q(stream_cmd_in[66]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[65] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[65]), .Q(stream_cmd_in[65]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[64] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[64]), .Q(stream_cmd_in[64]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[63] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[63]), .Q(stream_cmd_in[63]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[62] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[62]), .Q(stream_cmd_in[62]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[61] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[61]), .Q(stream_cmd_in[61]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[60] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[60]), .Q(stream_cmd_in[60]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[59] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[59]), .Q(stream_cmd_in[59]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[58] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[58]), .Q(stream_cmd_in[58]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[57] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[57]), .Q(stream_cmd_in[57]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[56] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[56]), .Q(stream_cmd_in[56]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[55] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[55]), .Q(stream_cmd_in[55]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[54] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[54]), .Q(stream_cmd_in[54]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[53] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[53]), .Q(stream_cmd_in[53]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[52] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[52]), .Q(stream_cmd_in[52]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[51] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[51]), .Q(stream_cmd_in[51]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[50] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[50]), .Q(stream_cmd_in[50]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[49] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[49]), .Q(stream_cmd_in[49]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[48] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[48]), .Q(stream_cmd_in[48]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[47] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[47]), .Q(stream_cmd_in[47]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[46] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[46]), .Q(stream_cmd_in[46]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[45] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[45]), .Q(stream_cmd_in[45]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[44] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[44]), .Q(stream_cmd_in[44]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[43] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[43]), .Q(stream_cmd_in[43]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[42] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[42]), .Q(stream_cmd_in[42]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[41] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[41]), .Q(stream_cmd_in[41]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[40] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[40]), .Q(stream_cmd_in[40]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[39] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[39]), .Q(stream_cmd_in[39]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[38] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[38]), .Q(stream_cmd_in[38]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[37] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[37]), .Q(stream_cmd_in[37]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[36] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[36]), .Q(stream_cmd_in[36]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[35] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[35]), .Q(stream_cmd_in[35]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[34] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[34]), .Q(stream_cmd_in[34]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[33] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[33]), .Q(stream_cmd_in[33]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[32] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[32]), .Q(stream_cmd_in[32]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[31] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[31]), .Q(stream_cmd_in[31]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[30] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[30]), .Q(stream_cmd_in[30]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[29] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[29]), .Q(stream_cmd_in[29]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[28] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[28]), .Q(stream_cmd_in[28]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[27] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[27]), .Q(stream_cmd_in[27]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[26] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[26]), .Q(stream_cmd_in[26]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[25] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[25]), .Q(stream_cmd_in[25]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[24] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[24]), .Q(stream_cmd_in[24]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[23] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[23]), .Q(stream_cmd_in[23]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[22] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[22]), .Q(stream_cmd_in[22]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[21] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[21]), .Q(stream_cmd_in[21]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[20] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[20]), .Q(stream_cmd_in[20]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[19] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[19]), .Q(stream_cmd_in[19]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[18] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[18]), .Q(stream_cmd_in[18]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[17] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[17]), .Q(stream_cmd_in[17]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[16] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[16]), .Q(stream_cmd_in[16]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[15] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[15]), .Q(stream_cmd_in[15]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[14] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[14]), .Q(stream_cmd_in[14]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[13] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[13]), .Q(stream_cmd_in[13]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[12] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[12]), .Q(stream_cmd_in[12]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[11] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[11]), .Q(stream_cmd_in[11]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[10] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[10]), .Q(stream_cmd_in[10]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[9] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[9]), .Q(stream_cmd_in[9]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[8] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[8]), .Q(stream_cmd_in[8]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[7] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[7]), .Q(stream_cmd_in[7]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[6] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[6]), .Q(stream_cmd_in[6]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[5] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[5]), .Q(stream_cmd_in[5]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[4] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[4]), .Q(stream_cmd_in[4]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[3] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[3]), .Q(stream_cmd_in[3]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[2] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[2]), .Q(stream_cmd_in[2]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[1] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[1]), .Q(stream_cmd_in[1]), .QN( ));
Q_FDP1 \stream_cmd_in_REG[0] ( .CK(clk), .R(rst_n), .D(stream_cmd_in_nxt[0]), .Q(stream_cmd_in[0]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[610] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[610]), .Q(gcm_dek_cmd_in[610]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[609] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[609]), .Q(gcm_dek_cmd_in[609]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[608] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[608]), .Q(gcm_dek_cmd_in[608]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[607] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[607]), .Q(gcm_dek_cmd_in[607]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[606] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[606]), .Q(gcm_dek_cmd_in[606]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[605] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[605]), .Q(gcm_dek_cmd_in[605]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[604] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[604]), .Q(gcm_dek_cmd_in[604]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[603] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[603]), .Q(gcm_dek_cmd_in[603]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[602] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[602]), .Q(gcm_dek_cmd_in[602]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[601] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[601]), .Q(gcm_dek_cmd_in[601]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[600] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[600]), .Q(gcm_dek_cmd_in[600]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[599] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[599]), .Q(gcm_dek_cmd_in[599]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[598] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[598]), .Q(gcm_dek_cmd_in[598]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[597] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[597]), .Q(gcm_dek_cmd_in[597]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[596] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[596]), .Q(gcm_dek_cmd_in[596]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[595] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[595]), .Q(gcm_dek_cmd_in[595]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[594] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[594]), .Q(gcm_dek_cmd_in[594]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[593] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[593]), .Q(gcm_dek_cmd_in[593]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[592] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[592]), .Q(gcm_dek_cmd_in[592]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[591] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[591]), .Q(gcm_dek_cmd_in[591]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[590] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[590]), .Q(gcm_dek_cmd_in[590]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[589] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[589]), .Q(gcm_dek_cmd_in[589]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[588] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[588]), .Q(gcm_dek_cmd_in[588]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[587] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[587]), .Q(gcm_dek_cmd_in[587]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[586] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[586]), .Q(gcm_dek_cmd_in[586]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[585] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[585]), .Q(gcm_dek_cmd_in[585]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[584] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[584]), .Q(gcm_dek_cmd_in[584]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[583] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[583]), .Q(gcm_dek_cmd_in[583]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[582] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[582]), .Q(gcm_dek_cmd_in[582]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[581] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[581]), .Q(gcm_dek_cmd_in[581]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[580] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[580]), .Q(gcm_dek_cmd_in[580]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[579] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[579]), .Q(gcm_dek_cmd_in[579]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[578] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[578]), .Q(gcm_dek_cmd_in[578]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[577] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[577]), .Q(gcm_dek_cmd_in[577]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[576] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[576]), .Q(gcm_dek_cmd_in[576]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[575] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[575]), .Q(gcm_dek_cmd_in[575]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[574] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[574]), .Q(gcm_dek_cmd_in[574]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[573] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[573]), .Q(gcm_dek_cmd_in[573]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[572] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[572]), .Q(gcm_dek_cmd_in[572]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[571] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[571]), .Q(gcm_dek_cmd_in[571]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[570] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[570]), .Q(gcm_dek_cmd_in[570]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[569] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[569]), .Q(gcm_dek_cmd_in[569]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[568] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[568]), .Q(gcm_dek_cmd_in[568]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[567] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[567]), .Q(gcm_dek_cmd_in[567]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[566] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[566]), .Q(gcm_dek_cmd_in[566]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[565] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[565]), .Q(gcm_dek_cmd_in[565]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[564] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[564]), .Q(gcm_dek_cmd_in[564]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[563] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[563]), .Q(gcm_dek_cmd_in[563]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[562] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[562]), .Q(gcm_dek_cmd_in[562]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[561] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[561]), .Q(gcm_dek_cmd_in[561]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[560] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[560]), .Q(gcm_dek_cmd_in[560]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[559] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[559]), .Q(gcm_dek_cmd_in[559]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[558] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[558]), .Q(gcm_dek_cmd_in[558]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[557] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[557]), .Q(gcm_dek_cmd_in[557]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[556] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[556]), .Q(gcm_dek_cmd_in[556]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[555] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[555]), .Q(gcm_dek_cmd_in[555]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[554] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[554]), .Q(gcm_dek_cmd_in[554]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[553] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[553]), .Q(gcm_dek_cmd_in[553]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[552] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[552]), .Q(gcm_dek_cmd_in[552]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[551] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[551]), .Q(gcm_dek_cmd_in[551]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[550] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[550]), .Q(gcm_dek_cmd_in[550]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[549] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[549]), .Q(gcm_dek_cmd_in[549]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[548] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[548]), .Q(gcm_dek_cmd_in[548]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[547] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[547]), .Q(gcm_dek_cmd_in[547]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[546] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[546]), .Q(gcm_dek_cmd_in[546]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[545] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[545]), .Q(gcm_dek_cmd_in[545]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[544] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[544]), .Q(gcm_dek_cmd_in[544]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[543] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[543]), .Q(gcm_dek_cmd_in[543]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[542] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[542]), .Q(gcm_dek_cmd_in[542]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[541] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[541]), .Q(gcm_dek_cmd_in[541]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[540] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[540]), .Q(gcm_dek_cmd_in[540]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[539] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[539]), .Q(gcm_dek_cmd_in[539]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[538] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[538]), .Q(gcm_dek_cmd_in[538]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[537] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[537]), .Q(gcm_dek_cmd_in[537]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[536] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[536]), .Q(gcm_dek_cmd_in[536]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[535] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[535]), .Q(gcm_dek_cmd_in[535]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[534] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[534]), .Q(gcm_dek_cmd_in[534]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[533] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[533]), .Q(gcm_dek_cmd_in[533]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[532] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[532]), .Q(gcm_dek_cmd_in[532]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[531] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[531]), .Q(gcm_dek_cmd_in[531]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[530] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[530]), .Q(gcm_dek_cmd_in[530]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[529] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[529]), .Q(gcm_dek_cmd_in[529]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[528] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[528]), .Q(gcm_dek_cmd_in[528]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[527] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[527]), .Q(gcm_dek_cmd_in[527]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[526] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[526]), .Q(gcm_dek_cmd_in[526]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[525] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[525]), .Q(gcm_dek_cmd_in[525]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[524] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[524]), .Q(gcm_dek_cmd_in[524]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[523] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[523]), .Q(gcm_dek_cmd_in[523]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[522] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[522]), .Q(gcm_dek_cmd_in[522]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[521] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[521]), .Q(gcm_dek_cmd_in[521]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[520] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[520]), .Q(gcm_dek_cmd_in[520]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[519] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[519]), .Q(gcm_dek_cmd_in[519]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[518] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[518]), .Q(gcm_dek_cmd_in[518]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[517] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[517]), .Q(gcm_dek_cmd_in[517]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[516] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[516]), .Q(gcm_dek_cmd_in[516]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[515] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[515]), .Q(gcm_dek_cmd_in[515]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[514] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[514]), .Q(gcm_dek_cmd_in[514]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[513] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[513]), .Q(gcm_dek_cmd_in[513]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[512] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[512]), .Q(gcm_dek_cmd_in[512]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[511] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[511]), .Q(gcm_dek_cmd_in[511]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[510] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[510]), .Q(gcm_dek_cmd_in[510]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[509] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[509]), .Q(gcm_dek_cmd_in[509]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[508] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[508]), .Q(gcm_dek_cmd_in[508]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[507] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[507]), .Q(gcm_dek_cmd_in[507]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[506] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[506]), .Q(gcm_dek_cmd_in[506]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[505] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[505]), .Q(gcm_dek_cmd_in[505]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[504] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[504]), .Q(gcm_dek_cmd_in[504]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[503] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[503]), .Q(gcm_dek_cmd_in[503]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[502] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[502]), .Q(gcm_dek_cmd_in[502]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[501] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[501]), .Q(gcm_dek_cmd_in[501]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[500] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[500]), .Q(gcm_dek_cmd_in[500]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[499] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[499]), .Q(gcm_dek_cmd_in[499]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[498] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[498]), .Q(gcm_dek_cmd_in[498]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[497] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[497]), .Q(gcm_dek_cmd_in[497]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[496] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[496]), .Q(gcm_dek_cmd_in[496]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[495] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[495]), .Q(gcm_dek_cmd_in[495]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[494] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[494]), .Q(gcm_dek_cmd_in[494]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[493] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[493]), .Q(gcm_dek_cmd_in[493]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[492] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[492]), .Q(gcm_dek_cmd_in[492]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[491] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[491]), .Q(gcm_dek_cmd_in[491]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[490] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[490]), .Q(gcm_dek_cmd_in[490]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[489] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[489]), .Q(gcm_dek_cmd_in[489]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[488] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[488]), .Q(gcm_dek_cmd_in[488]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[487] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[487]), .Q(gcm_dek_cmd_in[487]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[486] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[486]), .Q(gcm_dek_cmd_in[486]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[485] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[485]), .Q(gcm_dek_cmd_in[485]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[484] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[484]), .Q(gcm_dek_cmd_in[484]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[483] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[483]), .Q(gcm_dek_cmd_in[483]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[482] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[482]), .Q(gcm_dek_cmd_in[482]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[481] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[481]), .Q(gcm_dek_cmd_in[481]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[480] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[480]), .Q(gcm_dek_cmd_in[480]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[479] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[479]), .Q(gcm_dek_cmd_in[479]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[478] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[478]), .Q(gcm_dek_cmd_in[478]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[477] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[477]), .Q(gcm_dek_cmd_in[477]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[476] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[476]), .Q(gcm_dek_cmd_in[476]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[475] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[475]), .Q(gcm_dek_cmd_in[475]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[474] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[474]), .Q(gcm_dek_cmd_in[474]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[473] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[473]), .Q(gcm_dek_cmd_in[473]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[472] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[472]), .Q(gcm_dek_cmd_in[472]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[471] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[471]), .Q(gcm_dek_cmd_in[471]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[470] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[470]), .Q(gcm_dek_cmd_in[470]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[469] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[469]), .Q(gcm_dek_cmd_in[469]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[468] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[468]), .Q(gcm_dek_cmd_in[468]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[467] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[467]), .Q(gcm_dek_cmd_in[467]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[466] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[466]), .Q(gcm_dek_cmd_in[466]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[465] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[465]), .Q(gcm_dek_cmd_in[465]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[464] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[464]), .Q(gcm_dek_cmd_in[464]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[463] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[463]), .Q(gcm_dek_cmd_in[463]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[462] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[462]), .Q(gcm_dek_cmd_in[462]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[461] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[461]), .Q(gcm_dek_cmd_in[461]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[460] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[460]), .Q(gcm_dek_cmd_in[460]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[459] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[459]), .Q(gcm_dek_cmd_in[459]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[458] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[458]), .Q(gcm_dek_cmd_in[458]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[457] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[457]), .Q(gcm_dek_cmd_in[457]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[456] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[456]), .Q(gcm_dek_cmd_in[456]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[455] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[455]), .Q(gcm_dek_cmd_in[455]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[454] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[454]), .Q(gcm_dek_cmd_in[454]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[453] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[453]), .Q(gcm_dek_cmd_in[453]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[452] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[452]), .Q(gcm_dek_cmd_in[452]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[451] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[451]), .Q(gcm_dek_cmd_in[451]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[450] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[450]), .Q(gcm_dek_cmd_in[450]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[449] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[449]), .Q(gcm_dek_cmd_in[449]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[448] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[448]), .Q(gcm_dek_cmd_in[448]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[447] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[447]), .Q(gcm_dek_cmd_in[447]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[446] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[446]), .Q(gcm_dek_cmd_in[446]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[445] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[445]), .Q(gcm_dek_cmd_in[445]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[444] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[444]), .Q(gcm_dek_cmd_in[444]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[443] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[443]), .Q(gcm_dek_cmd_in[443]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[442] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[442]), .Q(gcm_dek_cmd_in[442]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[441] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[441]), .Q(gcm_dek_cmd_in[441]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[440] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[440]), .Q(gcm_dek_cmd_in[440]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[439] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[439]), .Q(gcm_dek_cmd_in[439]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[438] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[438]), .Q(gcm_dek_cmd_in[438]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[437] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[437]), .Q(gcm_dek_cmd_in[437]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[436] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[436]), .Q(gcm_dek_cmd_in[436]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[435] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[435]), .Q(gcm_dek_cmd_in[435]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[434] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[434]), .Q(gcm_dek_cmd_in[434]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[433] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[433]), .Q(gcm_dek_cmd_in[433]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[432] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[432]), .Q(gcm_dek_cmd_in[432]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[431] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[431]), .Q(gcm_dek_cmd_in[431]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[430] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[430]), .Q(gcm_dek_cmd_in[430]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[429] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[429]), .Q(gcm_dek_cmd_in[429]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[428] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[428]), .Q(gcm_dek_cmd_in[428]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[427] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[427]), .Q(gcm_dek_cmd_in[427]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[426] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[426]), .Q(gcm_dek_cmd_in[426]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[425] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[425]), .Q(gcm_dek_cmd_in[425]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[424] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[424]), .Q(gcm_dek_cmd_in[424]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[423] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[423]), .Q(gcm_dek_cmd_in[423]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[422] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[422]), .Q(gcm_dek_cmd_in[422]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[421] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[421]), .Q(gcm_dek_cmd_in[421]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[420] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[420]), .Q(gcm_dek_cmd_in[420]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[419] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[419]), .Q(gcm_dek_cmd_in[419]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[418] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[418]), .Q(gcm_dek_cmd_in[418]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[417] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[417]), .Q(gcm_dek_cmd_in[417]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[416] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[416]), .Q(gcm_dek_cmd_in[416]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[415] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[415]), .Q(gcm_dek_cmd_in[415]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[414] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[414]), .Q(gcm_dek_cmd_in[414]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[413] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[413]), .Q(gcm_dek_cmd_in[413]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[412] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[412]), .Q(gcm_dek_cmd_in[412]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[411] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[411]), .Q(gcm_dek_cmd_in[411]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[410] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[410]), .Q(gcm_dek_cmd_in[410]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[409] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[409]), .Q(gcm_dek_cmd_in[409]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[408] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[408]), .Q(gcm_dek_cmd_in[408]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[407] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[407]), .Q(gcm_dek_cmd_in[407]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[406] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[406]), .Q(gcm_dek_cmd_in[406]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[405] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[405]), .Q(gcm_dek_cmd_in[405]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[404] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[404]), .Q(gcm_dek_cmd_in[404]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[403] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[403]), .Q(gcm_dek_cmd_in[403]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[402] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[402]), .Q(gcm_dek_cmd_in[402]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[401] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[401]), .Q(gcm_dek_cmd_in[401]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[400] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[400]), .Q(gcm_dek_cmd_in[400]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[399] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[399]), .Q(gcm_dek_cmd_in[399]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[398] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[398]), .Q(gcm_dek_cmd_in[398]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[397] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[397]), .Q(gcm_dek_cmd_in[397]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[396] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[396]), .Q(gcm_dek_cmd_in[396]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[395] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[395]), .Q(gcm_dek_cmd_in[395]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[394] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[394]), .Q(gcm_dek_cmd_in[394]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[393] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[393]), .Q(gcm_dek_cmd_in[393]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[392] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[392]), .Q(gcm_dek_cmd_in[392]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[391] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[391]), .Q(gcm_dek_cmd_in[391]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[390] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[390]), .Q(gcm_dek_cmd_in[390]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[389] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[389]), .Q(gcm_dek_cmd_in[389]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[388] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[388]), .Q(gcm_dek_cmd_in[388]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[387] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[387]), .Q(gcm_dek_cmd_in[387]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[386] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[386]), .Q(gcm_dek_cmd_in[386]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[385] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[385]), .Q(gcm_dek_cmd_in[385]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[384] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[384]), .Q(gcm_dek_cmd_in[384]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[383] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[383]), .Q(gcm_dek_cmd_in[383]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[382] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[382]), .Q(gcm_dek_cmd_in[382]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[381] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[381]), .Q(gcm_dek_cmd_in[381]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[380] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[380]), .Q(gcm_dek_cmd_in[380]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[379] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[379]), .Q(gcm_dek_cmd_in[379]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[378] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[378]), .Q(gcm_dek_cmd_in[378]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[377] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[377]), .Q(gcm_dek_cmd_in[377]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[376] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[376]), .Q(gcm_dek_cmd_in[376]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[375] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[375]), .Q(gcm_dek_cmd_in[375]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[374] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[374]), .Q(gcm_dek_cmd_in[374]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[373] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[373]), .Q(gcm_dek_cmd_in[373]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[372] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[372]), .Q(gcm_dek_cmd_in[372]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[371] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[371]), .Q(gcm_dek_cmd_in[371]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[370] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[370]), .Q(gcm_dek_cmd_in[370]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[369] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[369]), .Q(gcm_dek_cmd_in[369]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[368] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[368]), .Q(gcm_dek_cmd_in[368]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[367] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[367]), .Q(gcm_dek_cmd_in[367]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[366] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[366]), .Q(gcm_dek_cmd_in[366]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[365] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[365]), .Q(gcm_dek_cmd_in[365]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[364] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[364]), .Q(gcm_dek_cmd_in[364]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[363] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[363]), .Q(gcm_dek_cmd_in[363]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[362] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[362]), .Q(gcm_dek_cmd_in[362]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[361] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[361]), .Q(gcm_dek_cmd_in[361]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[360] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[360]), .Q(gcm_dek_cmd_in[360]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[359] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[359]), .Q(gcm_dek_cmd_in[359]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[358] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[358]), .Q(gcm_dek_cmd_in[358]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[357] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[357]), .Q(gcm_dek_cmd_in[357]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[356] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[356]), .Q(gcm_dek_cmd_in[356]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[355] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[355]), .Q(gcm_dek_cmd_in[355]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[354] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[354]), .Q(gcm_dek_cmd_in[354]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[353] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[353]), .Q(gcm_dek_cmd_in[353]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[352] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[352]), .Q(gcm_dek_cmd_in[352]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[351] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[351]), .Q(gcm_dek_cmd_in[351]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[350] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[350]), .Q(gcm_dek_cmd_in[350]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[349] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[349]), .Q(gcm_dek_cmd_in[349]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[348] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[348]), .Q(gcm_dek_cmd_in[348]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[347] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[347]), .Q(gcm_dek_cmd_in[347]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[346] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[346]), .Q(gcm_dek_cmd_in[346]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[345] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[345]), .Q(gcm_dek_cmd_in[345]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[344] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[344]), .Q(gcm_dek_cmd_in[344]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[343] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[343]), .Q(gcm_dek_cmd_in[343]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[342] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[342]), .Q(gcm_dek_cmd_in[342]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[341] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[341]), .Q(gcm_dek_cmd_in[341]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[340] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[340]), .Q(gcm_dek_cmd_in[340]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[339] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[339]), .Q(gcm_dek_cmd_in[339]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[338] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[338]), .Q(gcm_dek_cmd_in[338]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[337] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[337]), .Q(gcm_dek_cmd_in[337]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[336] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[336]), .Q(gcm_dek_cmd_in[336]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[335] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[335]), .Q(gcm_dek_cmd_in[335]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[334] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[334]), .Q(gcm_dek_cmd_in[334]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[333] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[333]), .Q(gcm_dek_cmd_in[333]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[332] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[332]), .Q(gcm_dek_cmd_in[332]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[331] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[331]), .Q(gcm_dek_cmd_in[331]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[330] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[330]), .Q(gcm_dek_cmd_in[330]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[329] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[329]), .Q(gcm_dek_cmd_in[329]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[328] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[328]), .Q(gcm_dek_cmd_in[328]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[327] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[327]), .Q(gcm_dek_cmd_in[327]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[326] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[326]), .Q(gcm_dek_cmd_in[326]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[325] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[325]), .Q(gcm_dek_cmd_in[325]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[324] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[324]), .Q(gcm_dek_cmd_in[324]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[323] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[323]), .Q(gcm_dek_cmd_in[323]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[322] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[322]), .Q(gcm_dek_cmd_in[322]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[321] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[321]), .Q(gcm_dek_cmd_in[321]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[320] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[320]), .Q(gcm_dek_cmd_in[320]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[319] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[319]), .Q(gcm_dek_cmd_in[319]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[318] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[318]), .Q(gcm_dek_cmd_in[318]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[317] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[317]), .Q(gcm_dek_cmd_in[317]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[316] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[316]), .Q(gcm_dek_cmd_in[316]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[315] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[315]), .Q(gcm_dek_cmd_in[315]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[314] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[314]), .Q(gcm_dek_cmd_in[314]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[313] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[313]), .Q(gcm_dek_cmd_in[313]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[312] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[312]), .Q(gcm_dek_cmd_in[312]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[311] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[311]), .Q(gcm_dek_cmd_in[311]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[310] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[310]), .Q(gcm_dek_cmd_in[310]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[309] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[309]), .Q(gcm_dek_cmd_in[309]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[308] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[308]), .Q(gcm_dek_cmd_in[308]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[307] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[307]), .Q(gcm_dek_cmd_in[307]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[306] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[306]), .Q(gcm_dek_cmd_in[306]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[305] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[305]), .Q(gcm_dek_cmd_in[305]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[304] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[304]), .Q(gcm_dek_cmd_in[304]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[303] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[303]), .Q(gcm_dek_cmd_in[303]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[302] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[302]), .Q(gcm_dek_cmd_in[302]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[301] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[301]), .Q(gcm_dek_cmd_in[301]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[300] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[300]), .Q(gcm_dek_cmd_in[300]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[299] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[299]), .Q(gcm_dek_cmd_in[299]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[298] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[298]), .Q(gcm_dek_cmd_in[298]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[297] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[297]), .Q(gcm_dek_cmd_in[297]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[296] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[296]), .Q(gcm_dek_cmd_in[296]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[295] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[295]), .Q(gcm_dek_cmd_in[295]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[294] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[294]), .Q(gcm_dek_cmd_in[294]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[293] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[293]), .Q(gcm_dek_cmd_in[293]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[292] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[292]), .Q(gcm_dek_cmd_in[292]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[291] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[291]), .Q(gcm_dek_cmd_in[291]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[290] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[290]), .Q(gcm_dek_cmd_in[290]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[289] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[289]), .Q(gcm_dek_cmd_in[289]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[288] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[288]), .Q(gcm_dek_cmd_in[288]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[287] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[287]), .Q(gcm_dek_cmd_in[287]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[286] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[286]), .Q(gcm_dek_cmd_in[286]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[285] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[285]), .Q(gcm_dek_cmd_in[285]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[284] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[284]), .Q(gcm_dek_cmd_in[284]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[283] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[283]), .Q(gcm_dek_cmd_in[283]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[282] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[282]), .Q(gcm_dek_cmd_in[282]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[281] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[281]), .Q(gcm_dek_cmd_in[281]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[280] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[280]), .Q(gcm_dek_cmd_in[280]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[279] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[279]), .Q(gcm_dek_cmd_in[279]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[278] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[278]), .Q(gcm_dek_cmd_in[278]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[277] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[277]), .Q(gcm_dek_cmd_in[277]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[276] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[276]), .Q(gcm_dek_cmd_in[276]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[275] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[275]), .Q(gcm_dek_cmd_in[275]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[274] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[274]), .Q(gcm_dek_cmd_in[274]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[273] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[273]), .Q(gcm_dek_cmd_in[273]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[272] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[272]), .Q(gcm_dek_cmd_in[272]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[271] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[271]), .Q(gcm_dek_cmd_in[271]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[270] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[270]), .Q(gcm_dek_cmd_in[270]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[269] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[269]), .Q(gcm_dek_cmd_in[269]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[268] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[268]), .Q(gcm_dek_cmd_in[268]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[267] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[267]), .Q(gcm_dek_cmd_in[267]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[266] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[266]), .Q(gcm_dek_cmd_in[266]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[265] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[265]), .Q(gcm_dek_cmd_in[265]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[264] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[264]), .Q(gcm_dek_cmd_in[264]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[263] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[263]), .Q(gcm_dek_cmd_in[263]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[262] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[262]), .Q(gcm_dek_cmd_in[262]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[261] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[261]), .Q(gcm_dek_cmd_in[261]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[260] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[260]), .Q(gcm_dek_cmd_in[260]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[259] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[259]), .Q(gcm_dek_cmd_in[259]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[258] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[258]), .Q(gcm_dek_cmd_in[258]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[257] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[257]), .Q(gcm_dek_cmd_in[257]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[256] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[256]), .Q(gcm_dek_cmd_in[256]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[255] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[255]), .Q(gcm_dek_cmd_in[255]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[254] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[254]), .Q(gcm_dek_cmd_in[254]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[253] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[253]), .Q(gcm_dek_cmd_in[253]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[252] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[252]), .Q(gcm_dek_cmd_in[252]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[251] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[251]), .Q(gcm_dek_cmd_in[251]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[250] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[250]), .Q(gcm_dek_cmd_in[250]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[249] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[249]), .Q(gcm_dek_cmd_in[249]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[248] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[248]), .Q(gcm_dek_cmd_in[248]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[247] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[247]), .Q(gcm_dek_cmd_in[247]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[246] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[246]), .Q(gcm_dek_cmd_in[246]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[245] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[245]), .Q(gcm_dek_cmd_in[245]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[244] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[244]), .Q(gcm_dek_cmd_in[244]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[243] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[243]), .Q(gcm_dek_cmd_in[243]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[242] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[242]), .Q(gcm_dek_cmd_in[242]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[241] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[241]), .Q(gcm_dek_cmd_in[241]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[240] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[240]), .Q(gcm_dek_cmd_in[240]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[239] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[239]), .Q(gcm_dek_cmd_in[239]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[238] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[238]), .Q(gcm_dek_cmd_in[238]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[237] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[237]), .Q(gcm_dek_cmd_in[237]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[236] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[236]), .Q(gcm_dek_cmd_in[236]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[235] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[235]), .Q(gcm_dek_cmd_in[235]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[234] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[234]), .Q(gcm_dek_cmd_in[234]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[233] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[233]), .Q(gcm_dek_cmd_in[233]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[232] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[232]), .Q(gcm_dek_cmd_in[232]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[231] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[231]), .Q(gcm_dek_cmd_in[231]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[230] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[230]), .Q(gcm_dek_cmd_in[230]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[229] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[229]), .Q(gcm_dek_cmd_in[229]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[228] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[228]), .Q(gcm_dek_cmd_in[228]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[227] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[227]), .Q(gcm_dek_cmd_in[227]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[226] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[226]), .Q(gcm_dek_cmd_in[226]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[225] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[225]), .Q(gcm_dek_cmd_in[225]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[224] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[224]), .Q(gcm_dek_cmd_in[224]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[223] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[223]), .Q(gcm_dek_cmd_in[223]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[222] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[222]), .Q(gcm_dek_cmd_in[222]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[221] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[221]), .Q(gcm_dek_cmd_in[221]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[220] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[220]), .Q(gcm_dek_cmd_in[220]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[219] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[219]), .Q(gcm_dek_cmd_in[219]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[218] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[218]), .Q(gcm_dek_cmd_in[218]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[217] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[217]), .Q(gcm_dek_cmd_in[217]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[216] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[216]), .Q(gcm_dek_cmd_in[216]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[215] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[215]), .Q(gcm_dek_cmd_in[215]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[214] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[214]), .Q(gcm_dek_cmd_in[214]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[213] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[213]), .Q(gcm_dek_cmd_in[213]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[212] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[212]), .Q(gcm_dek_cmd_in[212]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[211] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[211]), .Q(gcm_dek_cmd_in[211]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[210] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[210]), .Q(gcm_dek_cmd_in[210]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[209] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[209]), .Q(gcm_dek_cmd_in[209]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[208] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[208]), .Q(gcm_dek_cmd_in[208]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[207] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[207]), .Q(gcm_dek_cmd_in[207]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[206] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[206]), .Q(gcm_dek_cmd_in[206]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[205] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[205]), .Q(gcm_dek_cmd_in[205]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[204] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[204]), .Q(gcm_dek_cmd_in[204]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[203] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[203]), .Q(gcm_dek_cmd_in[203]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[202] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[202]), .Q(gcm_dek_cmd_in[202]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[201] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[201]), .Q(gcm_dek_cmd_in[201]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[200] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[200]), .Q(gcm_dek_cmd_in[200]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[199] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[199]), .Q(gcm_dek_cmd_in[199]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[198] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[198]), .Q(gcm_dek_cmd_in[198]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[197] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[197]), .Q(gcm_dek_cmd_in[197]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[196] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[196]), .Q(gcm_dek_cmd_in[196]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[195] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[195]), .Q(gcm_dek_cmd_in[195]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[194] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[194]), .Q(gcm_dek_cmd_in[194]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[193] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[193]), .Q(gcm_dek_cmd_in[193]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[192] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[192]), .Q(gcm_dek_cmd_in[192]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[191] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[191]), .Q(gcm_dek_cmd_in[191]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[190] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[190]), .Q(gcm_dek_cmd_in[190]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[189] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[189]), .Q(gcm_dek_cmd_in[189]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[188] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[188]), .Q(gcm_dek_cmd_in[188]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[187] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[187]), .Q(gcm_dek_cmd_in[187]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[186] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[186]), .Q(gcm_dek_cmd_in[186]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[185] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[185]), .Q(gcm_dek_cmd_in[185]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[184] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[184]), .Q(gcm_dek_cmd_in[184]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[183] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[183]), .Q(gcm_dek_cmd_in[183]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[182] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[182]), .Q(gcm_dek_cmd_in[182]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[181] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[181]), .Q(gcm_dek_cmd_in[181]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[180] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[180]), .Q(gcm_dek_cmd_in[180]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[179] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[179]), .Q(gcm_dek_cmd_in[179]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[178] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[178]), .Q(gcm_dek_cmd_in[178]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[177] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[177]), .Q(gcm_dek_cmd_in[177]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[176] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[176]), .Q(gcm_dek_cmd_in[176]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[175] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[175]), .Q(gcm_dek_cmd_in[175]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[174] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[174]), .Q(gcm_dek_cmd_in[174]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[173] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[173]), .Q(gcm_dek_cmd_in[173]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[172] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[172]), .Q(gcm_dek_cmd_in[172]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[171] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[171]), .Q(gcm_dek_cmd_in[171]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[170] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[170]), .Q(gcm_dek_cmd_in[170]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[169] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[169]), .Q(gcm_dek_cmd_in[169]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[168] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[168]), .Q(gcm_dek_cmd_in[168]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[167] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[167]), .Q(gcm_dek_cmd_in[167]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[166] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[166]), .Q(gcm_dek_cmd_in[166]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[165] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[165]), .Q(gcm_dek_cmd_in[165]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[164] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[164]), .Q(gcm_dek_cmd_in[164]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[163] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[163]), .Q(gcm_dek_cmd_in[163]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[162] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[162]), .Q(gcm_dek_cmd_in[162]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[161] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[161]), .Q(gcm_dek_cmd_in[161]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[160] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[160]), .Q(gcm_dek_cmd_in[160]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[159] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[159]), .Q(gcm_dek_cmd_in[159]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[158] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[158]), .Q(gcm_dek_cmd_in[158]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[157] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[157]), .Q(gcm_dek_cmd_in[157]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[156] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[156]), .Q(gcm_dek_cmd_in[156]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[155] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[155]), .Q(gcm_dek_cmd_in[155]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[154] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[154]), .Q(gcm_dek_cmd_in[154]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[153] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[153]), .Q(gcm_dek_cmd_in[153]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[152] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[152]), .Q(gcm_dek_cmd_in[152]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[151] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[151]), .Q(gcm_dek_cmd_in[151]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[150] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[150]), .Q(gcm_dek_cmd_in[150]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[149] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[149]), .Q(gcm_dek_cmd_in[149]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[148] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[148]), .Q(gcm_dek_cmd_in[148]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[147] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[147]), .Q(gcm_dek_cmd_in[147]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[146] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[146]), .Q(gcm_dek_cmd_in[146]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[145] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[145]), .Q(gcm_dek_cmd_in[145]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[144] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[144]), .Q(gcm_dek_cmd_in[144]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[143] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[143]), .Q(gcm_dek_cmd_in[143]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[142] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[142]), .Q(gcm_dek_cmd_in[142]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[141] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[141]), .Q(gcm_dek_cmd_in[141]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[140] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[140]), .Q(gcm_dek_cmd_in[140]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[139] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[139]), .Q(gcm_dek_cmd_in[139]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[138] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[138]), .Q(gcm_dek_cmd_in[138]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[137] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[137]), .Q(gcm_dek_cmd_in[137]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[136] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[136]), .Q(gcm_dek_cmd_in[136]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[135] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[135]), .Q(gcm_dek_cmd_in[135]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[134] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[134]), .Q(gcm_dek_cmd_in[134]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[133] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[133]), .Q(gcm_dek_cmd_in[133]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[132] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[132]), .Q(gcm_dek_cmd_in[132]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[131] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[131]), .Q(gcm_dek_cmd_in[131]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[130] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[130]), .Q(gcm_dek_cmd_in[130]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[129] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[129]), .Q(gcm_dek_cmd_in[129]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[128] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[128]), .Q(gcm_dek_cmd_in[128]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[127] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[127]), .Q(gcm_dek_cmd_in[127]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[126] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[126]), .Q(gcm_dek_cmd_in[126]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[125] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[125]), .Q(gcm_dek_cmd_in[125]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[124] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[124]), .Q(gcm_dek_cmd_in[124]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[123] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[123]), .Q(gcm_dek_cmd_in[123]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[122] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[122]), .Q(gcm_dek_cmd_in[122]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[121] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[121]), .Q(gcm_dek_cmd_in[121]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[120] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[120]), .Q(gcm_dek_cmd_in[120]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[119] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[119]), .Q(gcm_dek_cmd_in[119]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[118] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[118]), .Q(gcm_dek_cmd_in[118]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[117] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[117]), .Q(gcm_dek_cmd_in[117]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[116] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[116]), .Q(gcm_dek_cmd_in[116]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[115] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[115]), .Q(gcm_dek_cmd_in[115]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[114] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[114]), .Q(gcm_dek_cmd_in[114]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[113] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[113]), .Q(gcm_dek_cmd_in[113]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[112] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[112]), .Q(gcm_dek_cmd_in[112]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[111] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[111]), .Q(gcm_dek_cmd_in[111]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[110] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[110]), .Q(gcm_dek_cmd_in[110]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[109] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[109]), .Q(gcm_dek_cmd_in[109]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[108] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[108]), .Q(gcm_dek_cmd_in[108]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[107] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[107]), .Q(gcm_dek_cmd_in[107]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[106] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[106]), .Q(gcm_dek_cmd_in[106]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[105] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[105]), .Q(gcm_dek_cmd_in[105]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[104] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[104]), .Q(gcm_dek_cmd_in[104]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[103] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[103]), .Q(gcm_dek_cmd_in[103]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[102] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[102]), .Q(gcm_dek_cmd_in[102]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[101] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[101]), .Q(gcm_dek_cmd_in[101]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[100] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[100]), .Q(gcm_dek_cmd_in[100]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[99] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[99]), .Q(gcm_dek_cmd_in[99]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[98] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[98]), .Q(gcm_dek_cmd_in[98]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[97] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[97]), .Q(gcm_dek_cmd_in[97]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[96] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[96]), .Q(gcm_dek_cmd_in[96]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[95] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[95]), .Q(gcm_dek_cmd_in[95]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[94] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[94]), .Q(gcm_dek_cmd_in[94]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[93] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[93]), .Q(gcm_dek_cmd_in[93]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[92] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[92]), .Q(gcm_dek_cmd_in[92]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[91] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[91]), .Q(gcm_dek_cmd_in[91]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[90] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[90]), .Q(gcm_dek_cmd_in[90]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[89] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[89]), .Q(gcm_dek_cmd_in[89]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[88] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[88]), .Q(gcm_dek_cmd_in[88]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[87] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[87]), .Q(gcm_dek_cmd_in[87]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[86] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[86]), .Q(gcm_dek_cmd_in[86]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[85] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[85]), .Q(gcm_dek_cmd_in[85]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[84] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[84]), .Q(gcm_dek_cmd_in[84]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[83] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[83]), .Q(gcm_dek_cmd_in[83]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[82] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[82]), .Q(gcm_dek_cmd_in[82]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[81] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[81]), .Q(gcm_dek_cmd_in[81]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[80] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[80]), .Q(gcm_dek_cmd_in[80]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[79] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[79]), .Q(gcm_dek_cmd_in[79]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[78] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[78]), .Q(gcm_dek_cmd_in[78]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[77] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[77]), .Q(gcm_dek_cmd_in[77]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[76] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[76]), .Q(gcm_dek_cmd_in[76]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[75] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[75]), .Q(gcm_dek_cmd_in[75]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[74] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[74]), .Q(gcm_dek_cmd_in[74]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[73] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[73]), .Q(gcm_dek_cmd_in[73]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[72] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[72]), .Q(gcm_dek_cmd_in[72]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[71] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[71]), .Q(gcm_dek_cmd_in[71]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[70] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[70]), .Q(gcm_dek_cmd_in[70]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[69] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[69]), .Q(gcm_dek_cmd_in[69]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[68] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[68]), .Q(gcm_dek_cmd_in[68]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[67] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[67]), .Q(gcm_dek_cmd_in[67]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[66] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[66]), .Q(gcm_dek_cmd_in[66]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[65] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[65]), .Q(gcm_dek_cmd_in[65]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[64] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[64]), .Q(gcm_dek_cmd_in[64]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[63] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[63]), .Q(gcm_dek_cmd_in[63]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[62] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[62]), .Q(gcm_dek_cmd_in[62]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[61] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[61]), .Q(gcm_dek_cmd_in[61]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[60] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[60]), .Q(gcm_dek_cmd_in[60]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[59] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[59]), .Q(gcm_dek_cmd_in[59]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[58] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[58]), .Q(gcm_dek_cmd_in[58]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[57] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[57]), .Q(gcm_dek_cmd_in[57]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[56] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[56]), .Q(gcm_dek_cmd_in[56]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[55] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[55]), .Q(gcm_dek_cmd_in[55]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[54] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[54]), .Q(gcm_dek_cmd_in[54]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[53] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[53]), .Q(gcm_dek_cmd_in[53]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[52] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[52]), .Q(gcm_dek_cmd_in[52]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[51] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[51]), .Q(gcm_dek_cmd_in[51]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[50] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[50]), .Q(gcm_dek_cmd_in[50]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[49] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[49]), .Q(gcm_dek_cmd_in[49]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[48] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[48]), .Q(gcm_dek_cmd_in[48]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[47] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[47]), .Q(gcm_dek_cmd_in[47]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[46] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[46]), .Q(gcm_dek_cmd_in[46]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[45] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[45]), .Q(gcm_dek_cmd_in[45]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[44] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[44]), .Q(gcm_dek_cmd_in[44]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[43] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[43]), .Q(gcm_dek_cmd_in[43]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[42] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[42]), .Q(gcm_dek_cmd_in[42]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[41] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[41]), .Q(gcm_dek_cmd_in[41]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[40] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[40]), .Q(gcm_dek_cmd_in[40]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[39] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[39]), .Q(gcm_dek_cmd_in[39]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[38] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[38]), .Q(gcm_dek_cmd_in[38]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[37] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[37]), .Q(gcm_dek_cmd_in[37]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[36] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[36]), .Q(gcm_dek_cmd_in[36]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[35] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[35]), .Q(gcm_dek_cmd_in[35]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[34] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[34]), .Q(gcm_dek_cmd_in[34]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[33] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[33]), .Q(gcm_dek_cmd_in[33]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[32] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[32]), .Q(gcm_dek_cmd_in[32]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[31] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[31]), .Q(gcm_dek_cmd_in[31]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[30] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[30]), .Q(gcm_dek_cmd_in[30]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[29] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[29]), .Q(gcm_dek_cmd_in[29]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[28] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[28]), .Q(gcm_dek_cmd_in[28]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[27] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[27]), .Q(gcm_dek_cmd_in[27]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[26] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[26]), .Q(gcm_dek_cmd_in[26]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[25] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[25]), .Q(gcm_dek_cmd_in[25]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[24] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[24]), .Q(gcm_dek_cmd_in[24]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[23] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[23]), .Q(gcm_dek_cmd_in[23]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[22] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[22]), .Q(gcm_dek_cmd_in[22]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[21] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[21]), .Q(gcm_dek_cmd_in[21]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[20] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[20]), .Q(gcm_dek_cmd_in[20]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[19] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[19]), .Q(gcm_dek_cmd_in[19]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[18] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[18]), .Q(gcm_dek_cmd_in[18]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[17] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[17]), .Q(gcm_dek_cmd_in[17]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[16] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[16]), .Q(gcm_dek_cmd_in[16]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[15] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[15]), .Q(gcm_dek_cmd_in[15]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[14] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[14]), .Q(gcm_dek_cmd_in[14]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[13] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[13]), .Q(gcm_dek_cmd_in[13]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[12] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[12]), .Q(gcm_dek_cmd_in[12]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[11] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[11]), .Q(gcm_dek_cmd_in[11]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[10] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[10]), .Q(gcm_dek_cmd_in[10]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[9] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[9]), .Q(gcm_dek_cmd_in[9]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[8] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[8]), .Q(gcm_dek_cmd_in[8]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[7] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[7]), .Q(gcm_dek_cmd_in[7]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[6] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[6]), .Q(gcm_dek_cmd_in[6]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[5] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[5]), .Q(gcm_dek_cmd_in[5]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[4] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[4]), .Q(gcm_dek_cmd_in[4]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[3] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[3]), .Q(gcm_dek_cmd_in[3]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[2] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[2]), .Q(gcm_dek_cmd_in[2]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[1] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[1]), .Q(gcm_dek_cmd_in[1]), .QN( ));
Q_FDP1 \gcm_dek_cmd_in_REG[0] ( .CK(clk), .R(rst_n), .D(gcm_dek_cmd_in_nxt[0]), .Q(gcm_dek_cmd_in[0]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[610] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[610]), .Q(gcm_dak_cmd_in[610]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[609] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[609]), .Q(gcm_dak_cmd_in[609]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[608] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[608]), .Q(gcm_dak_cmd_in[608]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[607] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[607]), .Q(gcm_dak_cmd_in[607]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[606] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[606]), .Q(gcm_dak_cmd_in[606]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[605] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[605]), .Q(gcm_dak_cmd_in[605]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[604] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[604]), .Q(gcm_dak_cmd_in[604]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[603] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[603]), .Q(gcm_dak_cmd_in[603]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[602] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[602]), .Q(gcm_dak_cmd_in[602]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[601] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[601]), .Q(gcm_dak_cmd_in[601]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[600] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[600]), .Q(gcm_dak_cmd_in[600]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[599] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[599]), .Q(gcm_dak_cmd_in[599]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[598] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[598]), .Q(gcm_dak_cmd_in[598]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[597] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[597]), .Q(gcm_dak_cmd_in[597]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[596] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[596]), .Q(gcm_dak_cmd_in[596]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[595] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[595]), .Q(gcm_dak_cmd_in[595]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[594] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[594]), .Q(gcm_dak_cmd_in[594]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[593] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[593]), .Q(gcm_dak_cmd_in[593]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[592] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[592]), .Q(gcm_dak_cmd_in[592]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[591] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[591]), .Q(gcm_dak_cmd_in[591]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[590] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[590]), .Q(gcm_dak_cmd_in[590]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[589] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[589]), .Q(gcm_dak_cmd_in[589]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[588] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[588]), .Q(gcm_dak_cmd_in[588]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[587] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[587]), .Q(gcm_dak_cmd_in[587]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[586] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[586]), .Q(gcm_dak_cmd_in[586]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[585] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[585]), .Q(gcm_dak_cmd_in[585]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[584] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[584]), .Q(gcm_dak_cmd_in[584]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[583] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[583]), .Q(gcm_dak_cmd_in[583]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[582] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[582]), .Q(gcm_dak_cmd_in[582]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[581] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[581]), .Q(gcm_dak_cmd_in[581]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[580] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[580]), .Q(gcm_dak_cmd_in[580]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[579] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[579]), .Q(gcm_dak_cmd_in[579]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[578] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[578]), .Q(gcm_dak_cmd_in[578]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[577] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[577]), .Q(gcm_dak_cmd_in[577]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[576] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[576]), .Q(gcm_dak_cmd_in[576]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[575] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[575]), .Q(gcm_dak_cmd_in[575]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[574] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[574]), .Q(gcm_dak_cmd_in[574]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[573] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[573]), .Q(gcm_dak_cmd_in[573]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[572] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[572]), .Q(gcm_dak_cmd_in[572]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[571] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[571]), .Q(gcm_dak_cmd_in[571]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[570] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[570]), .Q(gcm_dak_cmd_in[570]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[569] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[569]), .Q(gcm_dak_cmd_in[569]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[568] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[568]), .Q(gcm_dak_cmd_in[568]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[567] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[567]), .Q(gcm_dak_cmd_in[567]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[566] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[566]), .Q(gcm_dak_cmd_in[566]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[565] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[565]), .Q(gcm_dak_cmd_in[565]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[564] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[564]), .Q(gcm_dak_cmd_in[564]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[563] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[563]), .Q(gcm_dak_cmd_in[563]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[562] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[562]), .Q(gcm_dak_cmd_in[562]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[561] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[561]), .Q(gcm_dak_cmd_in[561]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[560] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[560]), .Q(gcm_dak_cmd_in[560]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[559] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[559]), .Q(gcm_dak_cmd_in[559]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[558] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[558]), .Q(gcm_dak_cmd_in[558]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[557] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[557]), .Q(gcm_dak_cmd_in[557]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[556] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[556]), .Q(gcm_dak_cmd_in[556]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[555] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[555]), .Q(gcm_dak_cmd_in[555]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[554] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[554]), .Q(gcm_dak_cmd_in[554]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[553] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[553]), .Q(gcm_dak_cmd_in[553]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[552] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[552]), .Q(gcm_dak_cmd_in[552]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[551] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[551]), .Q(gcm_dak_cmd_in[551]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[550] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[550]), .Q(gcm_dak_cmd_in[550]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[549] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[549]), .Q(gcm_dak_cmd_in[549]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[548] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[548]), .Q(gcm_dak_cmd_in[548]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[547] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[547]), .Q(gcm_dak_cmd_in[547]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[546] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[546]), .Q(gcm_dak_cmd_in[546]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[545] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[545]), .Q(gcm_dak_cmd_in[545]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[544] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[544]), .Q(gcm_dak_cmd_in[544]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[543] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[543]), .Q(gcm_dak_cmd_in[543]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[542] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[542]), .Q(gcm_dak_cmd_in[542]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[541] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[541]), .Q(gcm_dak_cmd_in[541]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[540] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[540]), .Q(gcm_dak_cmd_in[540]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[539] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[539]), .Q(gcm_dak_cmd_in[539]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[538] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[538]), .Q(gcm_dak_cmd_in[538]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[537] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[537]), .Q(gcm_dak_cmd_in[537]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[536] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[536]), .Q(gcm_dak_cmd_in[536]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[535] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[535]), .Q(gcm_dak_cmd_in[535]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[534] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[534]), .Q(gcm_dak_cmd_in[534]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[533] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[533]), .Q(gcm_dak_cmd_in[533]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[532] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[532]), .Q(gcm_dak_cmd_in[532]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[531] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[531]), .Q(gcm_dak_cmd_in[531]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[530] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[530]), .Q(gcm_dak_cmd_in[530]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[529] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[529]), .Q(gcm_dak_cmd_in[529]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[528] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[528]), .Q(gcm_dak_cmd_in[528]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[527] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[527]), .Q(gcm_dak_cmd_in[527]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[526] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[526]), .Q(gcm_dak_cmd_in[526]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[525] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[525]), .Q(gcm_dak_cmd_in[525]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[524] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[524]), .Q(gcm_dak_cmd_in[524]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[523] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[523]), .Q(gcm_dak_cmd_in[523]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[522] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[522]), .Q(gcm_dak_cmd_in[522]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[521] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[521]), .Q(gcm_dak_cmd_in[521]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[520] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[520]), .Q(gcm_dak_cmd_in[520]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[519] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[519]), .Q(gcm_dak_cmd_in[519]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[518] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[518]), .Q(gcm_dak_cmd_in[518]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[517] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[517]), .Q(gcm_dak_cmd_in[517]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[516] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[516]), .Q(gcm_dak_cmd_in[516]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[515] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[515]), .Q(gcm_dak_cmd_in[515]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[514] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[514]), .Q(gcm_dak_cmd_in[514]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[513] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[513]), .Q(gcm_dak_cmd_in[513]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[512] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[512]), .Q(gcm_dak_cmd_in[512]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[511] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[511]), .Q(gcm_dak_cmd_in[511]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[510] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[510]), .Q(gcm_dak_cmd_in[510]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[509] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[509]), .Q(gcm_dak_cmd_in[509]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[508] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[508]), .Q(gcm_dak_cmd_in[508]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[507] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[507]), .Q(gcm_dak_cmd_in[507]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[506] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[506]), .Q(gcm_dak_cmd_in[506]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[505] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[505]), .Q(gcm_dak_cmd_in[505]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[504] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[504]), .Q(gcm_dak_cmd_in[504]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[503] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[503]), .Q(gcm_dak_cmd_in[503]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[502] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[502]), .Q(gcm_dak_cmd_in[502]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[501] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[501]), .Q(gcm_dak_cmd_in[501]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[500] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[500]), .Q(gcm_dak_cmd_in[500]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[499] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[499]), .Q(gcm_dak_cmd_in[499]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[498] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[498]), .Q(gcm_dak_cmd_in[498]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[497] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[497]), .Q(gcm_dak_cmd_in[497]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[496] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[496]), .Q(gcm_dak_cmd_in[496]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[495] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[495]), .Q(gcm_dak_cmd_in[495]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[494] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[494]), .Q(gcm_dak_cmd_in[494]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[493] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[493]), .Q(gcm_dak_cmd_in[493]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[492] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[492]), .Q(gcm_dak_cmd_in[492]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[491] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[491]), .Q(gcm_dak_cmd_in[491]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[490] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[490]), .Q(gcm_dak_cmd_in[490]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[489] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[489]), .Q(gcm_dak_cmd_in[489]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[488] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[488]), .Q(gcm_dak_cmd_in[488]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[487] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[487]), .Q(gcm_dak_cmd_in[487]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[486] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[486]), .Q(gcm_dak_cmd_in[486]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[485] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[485]), .Q(gcm_dak_cmd_in[485]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[484] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[484]), .Q(gcm_dak_cmd_in[484]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[483] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[483]), .Q(gcm_dak_cmd_in[483]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[482] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[482]), .Q(gcm_dak_cmd_in[482]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[481] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[481]), .Q(gcm_dak_cmd_in[481]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[480] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[480]), .Q(gcm_dak_cmd_in[480]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[479] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[479]), .Q(gcm_dak_cmd_in[479]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[478] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[478]), .Q(gcm_dak_cmd_in[478]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[477] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[477]), .Q(gcm_dak_cmd_in[477]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[476] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[476]), .Q(gcm_dak_cmd_in[476]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[475] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[475]), .Q(gcm_dak_cmd_in[475]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[474] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[474]), .Q(gcm_dak_cmd_in[474]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[473] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[473]), .Q(gcm_dak_cmd_in[473]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[472] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[472]), .Q(gcm_dak_cmd_in[472]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[471] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[471]), .Q(gcm_dak_cmd_in[471]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[470] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[470]), .Q(gcm_dak_cmd_in[470]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[469] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[469]), .Q(gcm_dak_cmd_in[469]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[468] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[468]), .Q(gcm_dak_cmd_in[468]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[467] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[467]), .Q(gcm_dak_cmd_in[467]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[466] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[466]), .Q(gcm_dak_cmd_in[466]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[465] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[465]), .Q(gcm_dak_cmd_in[465]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[464] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[464]), .Q(gcm_dak_cmd_in[464]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[463] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[463]), .Q(gcm_dak_cmd_in[463]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[462] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[462]), .Q(gcm_dak_cmd_in[462]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[461] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[461]), .Q(gcm_dak_cmd_in[461]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[460] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[460]), .Q(gcm_dak_cmd_in[460]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[459] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[459]), .Q(gcm_dak_cmd_in[459]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[458] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[458]), .Q(gcm_dak_cmd_in[458]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[457] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[457]), .Q(gcm_dak_cmd_in[457]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[456] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[456]), .Q(gcm_dak_cmd_in[456]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[455] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[455]), .Q(gcm_dak_cmd_in[455]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[454] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[454]), .Q(gcm_dak_cmd_in[454]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[453] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[453]), .Q(gcm_dak_cmd_in[453]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[452] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[452]), .Q(gcm_dak_cmd_in[452]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[451] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[451]), .Q(gcm_dak_cmd_in[451]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[450] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[450]), .Q(gcm_dak_cmd_in[450]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[449] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[449]), .Q(gcm_dak_cmd_in[449]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[448] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[448]), .Q(gcm_dak_cmd_in[448]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[447] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[447]), .Q(gcm_dak_cmd_in[447]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[446] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[446]), .Q(gcm_dak_cmd_in[446]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[445] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[445]), .Q(gcm_dak_cmd_in[445]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[444] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[444]), .Q(gcm_dak_cmd_in[444]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[443] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[443]), .Q(gcm_dak_cmd_in[443]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[442] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[442]), .Q(gcm_dak_cmd_in[442]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[441] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[441]), .Q(gcm_dak_cmd_in[441]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[440] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[440]), .Q(gcm_dak_cmd_in[440]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[439] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[439]), .Q(gcm_dak_cmd_in[439]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[438] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[438]), .Q(gcm_dak_cmd_in[438]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[437] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[437]), .Q(gcm_dak_cmd_in[437]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[436] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[436]), .Q(gcm_dak_cmd_in[436]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[435] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[435]), .Q(gcm_dak_cmd_in[435]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[434] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[434]), .Q(gcm_dak_cmd_in[434]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[433] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[433]), .Q(gcm_dak_cmd_in[433]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[432] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[432]), .Q(gcm_dak_cmd_in[432]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[431] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[431]), .Q(gcm_dak_cmd_in[431]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[430] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[430]), .Q(gcm_dak_cmd_in[430]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[429] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[429]), .Q(gcm_dak_cmd_in[429]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[428] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[428]), .Q(gcm_dak_cmd_in[428]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[427] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[427]), .Q(gcm_dak_cmd_in[427]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[426] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[426]), .Q(gcm_dak_cmd_in[426]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[425] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[425]), .Q(gcm_dak_cmd_in[425]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[424] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[424]), .Q(gcm_dak_cmd_in[424]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[423] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[423]), .Q(gcm_dak_cmd_in[423]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[422] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[422]), .Q(gcm_dak_cmd_in[422]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[421] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[421]), .Q(gcm_dak_cmd_in[421]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[420] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[420]), .Q(gcm_dak_cmd_in[420]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[419] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[419]), .Q(gcm_dak_cmd_in[419]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[418] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[418]), .Q(gcm_dak_cmd_in[418]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[417] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[417]), .Q(gcm_dak_cmd_in[417]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[416] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[416]), .Q(gcm_dak_cmd_in[416]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[415] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[415]), .Q(gcm_dak_cmd_in[415]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[414] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[414]), .Q(gcm_dak_cmd_in[414]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[413] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[413]), .Q(gcm_dak_cmd_in[413]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[412] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[412]), .Q(gcm_dak_cmd_in[412]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[411] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[411]), .Q(gcm_dak_cmd_in[411]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[410] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[410]), .Q(gcm_dak_cmd_in[410]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[409] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[409]), .Q(gcm_dak_cmd_in[409]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[408] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[408]), .Q(gcm_dak_cmd_in[408]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[407] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[407]), .Q(gcm_dak_cmd_in[407]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[406] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[406]), .Q(gcm_dak_cmd_in[406]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[405] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[405]), .Q(gcm_dak_cmd_in[405]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[404] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[404]), .Q(gcm_dak_cmd_in[404]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[403] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[403]), .Q(gcm_dak_cmd_in[403]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[402] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[402]), .Q(gcm_dak_cmd_in[402]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[401] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[401]), .Q(gcm_dak_cmd_in[401]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[400] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[400]), .Q(gcm_dak_cmd_in[400]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[399] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[399]), .Q(gcm_dak_cmd_in[399]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[398] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[398]), .Q(gcm_dak_cmd_in[398]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[397] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[397]), .Q(gcm_dak_cmd_in[397]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[396] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[396]), .Q(gcm_dak_cmd_in[396]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[395] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[395]), .Q(gcm_dak_cmd_in[395]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[394] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[394]), .Q(gcm_dak_cmd_in[394]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[393] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[393]), .Q(gcm_dak_cmd_in[393]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[392] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[392]), .Q(gcm_dak_cmd_in[392]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[391] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[391]), .Q(gcm_dak_cmd_in[391]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[390] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[390]), .Q(gcm_dak_cmd_in[390]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[389] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[389]), .Q(gcm_dak_cmd_in[389]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[388] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[388]), .Q(gcm_dak_cmd_in[388]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[387] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[387]), .Q(gcm_dak_cmd_in[387]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[386] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[386]), .Q(gcm_dak_cmd_in[386]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[385] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[385]), .Q(gcm_dak_cmd_in[385]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[384] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[384]), .Q(gcm_dak_cmd_in[384]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[383] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[383]), .Q(gcm_dak_cmd_in[383]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[382] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[382]), .Q(gcm_dak_cmd_in[382]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[381] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[381]), .Q(gcm_dak_cmd_in[381]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[380] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[380]), .Q(gcm_dak_cmd_in[380]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[379] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[379]), .Q(gcm_dak_cmd_in[379]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[378] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[378]), .Q(gcm_dak_cmd_in[378]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[377] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[377]), .Q(gcm_dak_cmd_in[377]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[376] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[376]), .Q(gcm_dak_cmd_in[376]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[375] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[375]), .Q(gcm_dak_cmd_in[375]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[374] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[374]), .Q(gcm_dak_cmd_in[374]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[373] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[373]), .Q(gcm_dak_cmd_in[373]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[372] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[372]), .Q(gcm_dak_cmd_in[372]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[371] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[371]), .Q(gcm_dak_cmd_in[371]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[370] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[370]), .Q(gcm_dak_cmd_in[370]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[369] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[369]), .Q(gcm_dak_cmd_in[369]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[368] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[368]), .Q(gcm_dak_cmd_in[368]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[367] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[367]), .Q(gcm_dak_cmd_in[367]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[366] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[366]), .Q(gcm_dak_cmd_in[366]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[365] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[365]), .Q(gcm_dak_cmd_in[365]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[364] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[364]), .Q(gcm_dak_cmd_in[364]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[363] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[363]), .Q(gcm_dak_cmd_in[363]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[362] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[362]), .Q(gcm_dak_cmd_in[362]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[361] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[361]), .Q(gcm_dak_cmd_in[361]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[360] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[360]), .Q(gcm_dak_cmd_in[360]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[359] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[359]), .Q(gcm_dak_cmd_in[359]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[358] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[358]), .Q(gcm_dak_cmd_in[358]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[357] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[357]), .Q(gcm_dak_cmd_in[357]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[356] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[356]), .Q(gcm_dak_cmd_in[356]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[355] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[355]), .Q(gcm_dak_cmd_in[355]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[354] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[354]), .Q(gcm_dak_cmd_in[354]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[353] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[353]), .Q(gcm_dak_cmd_in[353]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[352] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[352]), .Q(gcm_dak_cmd_in[352]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[351] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[351]), .Q(gcm_dak_cmd_in[351]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[350] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[350]), .Q(gcm_dak_cmd_in[350]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[349] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[349]), .Q(gcm_dak_cmd_in[349]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[348] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[348]), .Q(gcm_dak_cmd_in[348]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[347] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[347]), .Q(gcm_dak_cmd_in[347]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[346] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[346]), .Q(gcm_dak_cmd_in[346]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[345] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[345]), .Q(gcm_dak_cmd_in[345]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[344] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[344]), .Q(gcm_dak_cmd_in[344]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[343] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[343]), .Q(gcm_dak_cmd_in[343]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[342] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[342]), .Q(gcm_dak_cmd_in[342]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[341] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[341]), .Q(gcm_dak_cmd_in[341]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[340] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[340]), .Q(gcm_dak_cmd_in[340]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[339] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[339]), .Q(gcm_dak_cmd_in[339]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[338] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[338]), .Q(gcm_dak_cmd_in[338]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[337] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[337]), .Q(gcm_dak_cmd_in[337]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[336] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[336]), .Q(gcm_dak_cmd_in[336]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[335] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[335]), .Q(gcm_dak_cmd_in[335]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[334] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[334]), .Q(gcm_dak_cmd_in[334]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[333] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[333]), .Q(gcm_dak_cmd_in[333]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[332] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[332]), .Q(gcm_dak_cmd_in[332]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[331] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[331]), .Q(gcm_dak_cmd_in[331]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[330] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[330]), .Q(gcm_dak_cmd_in[330]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[329] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[329]), .Q(gcm_dak_cmd_in[329]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[328] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[328]), .Q(gcm_dak_cmd_in[328]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[327] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[327]), .Q(gcm_dak_cmd_in[327]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[326] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[326]), .Q(gcm_dak_cmd_in[326]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[325] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[325]), .Q(gcm_dak_cmd_in[325]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[324] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[324]), .Q(gcm_dak_cmd_in[324]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[323] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[323]), .Q(gcm_dak_cmd_in[323]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[322] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[322]), .Q(gcm_dak_cmd_in[322]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[321] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[321]), .Q(gcm_dak_cmd_in[321]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[320] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[320]), .Q(gcm_dak_cmd_in[320]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[319] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[319]), .Q(gcm_dak_cmd_in[319]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[318] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[318]), .Q(gcm_dak_cmd_in[318]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[317] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[317]), .Q(gcm_dak_cmd_in[317]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[316] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[316]), .Q(gcm_dak_cmd_in[316]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[315] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[315]), .Q(gcm_dak_cmd_in[315]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[314] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[314]), .Q(gcm_dak_cmd_in[314]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[313] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[313]), .Q(gcm_dak_cmd_in[313]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[312] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[312]), .Q(gcm_dak_cmd_in[312]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[311] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[311]), .Q(gcm_dak_cmd_in[311]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[310] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[310]), .Q(gcm_dak_cmd_in[310]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[309] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[309]), .Q(gcm_dak_cmd_in[309]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[308] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[308]), .Q(gcm_dak_cmd_in[308]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[307] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[307]), .Q(gcm_dak_cmd_in[307]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[306] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[306]), .Q(gcm_dak_cmd_in[306]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[305] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[305]), .Q(gcm_dak_cmd_in[305]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[304] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[304]), .Q(gcm_dak_cmd_in[304]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[303] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[303]), .Q(gcm_dak_cmd_in[303]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[302] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[302]), .Q(gcm_dak_cmd_in[302]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[301] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[301]), .Q(gcm_dak_cmd_in[301]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[300] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[300]), .Q(gcm_dak_cmd_in[300]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[299] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[299]), .Q(gcm_dak_cmd_in[299]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[298] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[298]), .Q(gcm_dak_cmd_in[298]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[297] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[297]), .Q(gcm_dak_cmd_in[297]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[296] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[296]), .Q(gcm_dak_cmd_in[296]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[295] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[295]), .Q(gcm_dak_cmd_in[295]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[294] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[294]), .Q(gcm_dak_cmd_in[294]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[293] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[293]), .Q(gcm_dak_cmd_in[293]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[292] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[292]), .Q(gcm_dak_cmd_in[292]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[291] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[291]), .Q(gcm_dak_cmd_in[291]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[290] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[290]), .Q(gcm_dak_cmd_in[290]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[289] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[289]), .Q(gcm_dak_cmd_in[289]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[288] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[288]), .Q(gcm_dak_cmd_in[288]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[287] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[287]), .Q(gcm_dak_cmd_in[287]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[286] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[286]), .Q(gcm_dak_cmd_in[286]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[285] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[285]), .Q(gcm_dak_cmd_in[285]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[284] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[284]), .Q(gcm_dak_cmd_in[284]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[283] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[283]), .Q(gcm_dak_cmd_in[283]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[282] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[282]), .Q(gcm_dak_cmd_in[282]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[281] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[281]), .Q(gcm_dak_cmd_in[281]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[280] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[280]), .Q(gcm_dak_cmd_in[280]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[279] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[279]), .Q(gcm_dak_cmd_in[279]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[278] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[278]), .Q(gcm_dak_cmd_in[278]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[277] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[277]), .Q(gcm_dak_cmd_in[277]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[276] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[276]), .Q(gcm_dak_cmd_in[276]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[275] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[275]), .Q(gcm_dak_cmd_in[275]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[274] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[274]), .Q(gcm_dak_cmd_in[274]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[273] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[273]), .Q(gcm_dak_cmd_in[273]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[272] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[272]), .Q(gcm_dak_cmd_in[272]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[271] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[271]), .Q(gcm_dak_cmd_in[271]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[270] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[270]), .Q(gcm_dak_cmd_in[270]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[269] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[269]), .Q(gcm_dak_cmd_in[269]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[268] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[268]), .Q(gcm_dak_cmd_in[268]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[267] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[267]), .Q(gcm_dak_cmd_in[267]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[266] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[266]), .Q(gcm_dak_cmd_in[266]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[265] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[265]), .Q(gcm_dak_cmd_in[265]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[264] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[264]), .Q(gcm_dak_cmd_in[264]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[263] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[263]), .Q(gcm_dak_cmd_in[263]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[262] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[262]), .Q(gcm_dak_cmd_in[262]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[261] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[261]), .Q(gcm_dak_cmd_in[261]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[260] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[260]), .Q(gcm_dak_cmd_in[260]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[259] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[259]), .Q(gcm_dak_cmd_in[259]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[258] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[258]), .Q(gcm_dak_cmd_in[258]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[257] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[257]), .Q(gcm_dak_cmd_in[257]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[256] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[256]), .Q(gcm_dak_cmd_in[256]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[255] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[255]), .Q(gcm_dak_cmd_in[255]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[254] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[254]), .Q(gcm_dak_cmd_in[254]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[253] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[253]), .Q(gcm_dak_cmd_in[253]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[252] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[252]), .Q(gcm_dak_cmd_in[252]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[251] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[251]), .Q(gcm_dak_cmd_in[251]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[250] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[250]), .Q(gcm_dak_cmd_in[250]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[249] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[249]), .Q(gcm_dak_cmd_in[249]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[248] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[248]), .Q(gcm_dak_cmd_in[248]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[247] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[247]), .Q(gcm_dak_cmd_in[247]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[246] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[246]), .Q(gcm_dak_cmd_in[246]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[245] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[245]), .Q(gcm_dak_cmd_in[245]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[244] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[244]), .Q(gcm_dak_cmd_in[244]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[243] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[243]), .Q(gcm_dak_cmd_in[243]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[242] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[242]), .Q(gcm_dak_cmd_in[242]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[241] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[241]), .Q(gcm_dak_cmd_in[241]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[240] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[240]), .Q(gcm_dak_cmd_in[240]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[239] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[239]), .Q(gcm_dak_cmd_in[239]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[238] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[238]), .Q(gcm_dak_cmd_in[238]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[237] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[237]), .Q(gcm_dak_cmd_in[237]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[236] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[236]), .Q(gcm_dak_cmd_in[236]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[235] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[235]), .Q(gcm_dak_cmd_in[235]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[234] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[234]), .Q(gcm_dak_cmd_in[234]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[233] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[233]), .Q(gcm_dak_cmd_in[233]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[232] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[232]), .Q(gcm_dak_cmd_in[232]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[231] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[231]), .Q(gcm_dak_cmd_in[231]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[230] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[230]), .Q(gcm_dak_cmd_in[230]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[229] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[229]), .Q(gcm_dak_cmd_in[229]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[228] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[228]), .Q(gcm_dak_cmd_in[228]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[227] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[227]), .Q(gcm_dak_cmd_in[227]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[226] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[226]), .Q(gcm_dak_cmd_in[226]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[225] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[225]), .Q(gcm_dak_cmd_in[225]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[224] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[224]), .Q(gcm_dak_cmd_in[224]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[223] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[223]), .Q(gcm_dak_cmd_in[223]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[222] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[222]), .Q(gcm_dak_cmd_in[222]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[221] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[221]), .Q(gcm_dak_cmd_in[221]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[220] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[220]), .Q(gcm_dak_cmd_in[220]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[219] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[219]), .Q(gcm_dak_cmd_in[219]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[218] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[218]), .Q(gcm_dak_cmd_in[218]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[217] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[217]), .Q(gcm_dak_cmd_in[217]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[216] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[216]), .Q(gcm_dak_cmd_in[216]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[215] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[215]), .Q(gcm_dak_cmd_in[215]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[214] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[214]), .Q(gcm_dak_cmd_in[214]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[213] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[213]), .Q(gcm_dak_cmd_in[213]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[212] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[212]), .Q(gcm_dak_cmd_in[212]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[211] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[211]), .Q(gcm_dak_cmd_in[211]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[210] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[210]), .Q(gcm_dak_cmd_in[210]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[209] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[209]), .Q(gcm_dak_cmd_in[209]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[208] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[208]), .Q(gcm_dak_cmd_in[208]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[207] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[207]), .Q(gcm_dak_cmd_in[207]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[206] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[206]), .Q(gcm_dak_cmd_in[206]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[205] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[205]), .Q(gcm_dak_cmd_in[205]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[204] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[204]), .Q(gcm_dak_cmd_in[204]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[203] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[203]), .Q(gcm_dak_cmd_in[203]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[202] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[202]), .Q(gcm_dak_cmd_in[202]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[201] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[201]), .Q(gcm_dak_cmd_in[201]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[200] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[200]), .Q(gcm_dak_cmd_in[200]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[199] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[199]), .Q(gcm_dak_cmd_in[199]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[198] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[198]), .Q(gcm_dak_cmd_in[198]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[197] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[197]), .Q(gcm_dak_cmd_in[197]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[196] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[196]), .Q(gcm_dak_cmd_in[196]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[195] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[195]), .Q(gcm_dak_cmd_in[195]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[194] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[194]), .Q(gcm_dak_cmd_in[194]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[193] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[193]), .Q(gcm_dak_cmd_in[193]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[192] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[192]), .Q(gcm_dak_cmd_in[192]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[191] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[191]), .Q(gcm_dak_cmd_in[191]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[190] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[190]), .Q(gcm_dak_cmd_in[190]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[189] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[189]), .Q(gcm_dak_cmd_in[189]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[188] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[188]), .Q(gcm_dak_cmd_in[188]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[187] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[187]), .Q(gcm_dak_cmd_in[187]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[186] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[186]), .Q(gcm_dak_cmd_in[186]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[185] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[185]), .Q(gcm_dak_cmd_in[185]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[184] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[184]), .Q(gcm_dak_cmd_in[184]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[183] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[183]), .Q(gcm_dak_cmd_in[183]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[182] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[182]), .Q(gcm_dak_cmd_in[182]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[181] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[181]), .Q(gcm_dak_cmd_in[181]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[180] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[180]), .Q(gcm_dak_cmd_in[180]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[179] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[179]), .Q(gcm_dak_cmd_in[179]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[178] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[178]), .Q(gcm_dak_cmd_in[178]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[177] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[177]), .Q(gcm_dak_cmd_in[177]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[176] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[176]), .Q(gcm_dak_cmd_in[176]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[175] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[175]), .Q(gcm_dak_cmd_in[175]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[174] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[174]), .Q(gcm_dak_cmd_in[174]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[173] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[173]), .Q(gcm_dak_cmd_in[173]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[172] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[172]), .Q(gcm_dak_cmd_in[172]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[171] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[171]), .Q(gcm_dak_cmd_in[171]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[170] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[170]), .Q(gcm_dak_cmd_in[170]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[169] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[169]), .Q(gcm_dak_cmd_in[169]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[168] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[168]), .Q(gcm_dak_cmd_in[168]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[167] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[167]), .Q(gcm_dak_cmd_in[167]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[166] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[166]), .Q(gcm_dak_cmd_in[166]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[165] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[165]), .Q(gcm_dak_cmd_in[165]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[164] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[164]), .Q(gcm_dak_cmd_in[164]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[163] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[163]), .Q(gcm_dak_cmd_in[163]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[162] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[162]), .Q(gcm_dak_cmd_in[162]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[161] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[161]), .Q(gcm_dak_cmd_in[161]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[160] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[160]), .Q(gcm_dak_cmd_in[160]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[159] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[159]), .Q(gcm_dak_cmd_in[159]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[158] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[158]), .Q(gcm_dak_cmd_in[158]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[157] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[157]), .Q(gcm_dak_cmd_in[157]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[156] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[156]), .Q(gcm_dak_cmd_in[156]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[155] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[155]), .Q(gcm_dak_cmd_in[155]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[154] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[154]), .Q(gcm_dak_cmd_in[154]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[153] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[153]), .Q(gcm_dak_cmd_in[153]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[152] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[152]), .Q(gcm_dak_cmd_in[152]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[151] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[151]), .Q(gcm_dak_cmd_in[151]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[150] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[150]), .Q(gcm_dak_cmd_in[150]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[149] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[149]), .Q(gcm_dak_cmd_in[149]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[148] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[148]), .Q(gcm_dak_cmd_in[148]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[147] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[147]), .Q(gcm_dak_cmd_in[147]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[146] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[146]), .Q(gcm_dak_cmd_in[146]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[145] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[145]), .Q(gcm_dak_cmd_in[145]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[144] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[144]), .Q(gcm_dak_cmd_in[144]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[143] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[143]), .Q(gcm_dak_cmd_in[143]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[142] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[142]), .Q(gcm_dak_cmd_in[142]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[141] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[141]), .Q(gcm_dak_cmd_in[141]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[140] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[140]), .Q(gcm_dak_cmd_in[140]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[139] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[139]), .Q(gcm_dak_cmd_in[139]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[138] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[138]), .Q(gcm_dak_cmd_in[138]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[137] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[137]), .Q(gcm_dak_cmd_in[137]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[136] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[136]), .Q(gcm_dak_cmd_in[136]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[135] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[135]), .Q(gcm_dak_cmd_in[135]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[134] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[134]), .Q(gcm_dak_cmd_in[134]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[133] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[133]), .Q(gcm_dak_cmd_in[133]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[132] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[132]), .Q(gcm_dak_cmd_in[132]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[131] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[131]), .Q(gcm_dak_cmd_in[131]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[130] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[130]), .Q(gcm_dak_cmd_in[130]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[129] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[129]), .Q(gcm_dak_cmd_in[129]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[128] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[128]), .Q(gcm_dak_cmd_in[128]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[127] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[127]), .Q(gcm_dak_cmd_in[127]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[126] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[126]), .Q(gcm_dak_cmd_in[126]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[125] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[125]), .Q(gcm_dak_cmd_in[125]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[124] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[124]), .Q(gcm_dak_cmd_in[124]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[123] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[123]), .Q(gcm_dak_cmd_in[123]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[122] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[122]), .Q(gcm_dak_cmd_in[122]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[121] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[121]), .Q(gcm_dak_cmd_in[121]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[120] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[120]), .Q(gcm_dak_cmd_in[120]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[119] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[119]), .Q(gcm_dak_cmd_in[119]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[118] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[118]), .Q(gcm_dak_cmd_in[118]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[117] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[117]), .Q(gcm_dak_cmd_in[117]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[116] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[116]), .Q(gcm_dak_cmd_in[116]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[115] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[115]), .Q(gcm_dak_cmd_in[115]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[114] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[114]), .Q(gcm_dak_cmd_in[114]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[113] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[113]), .Q(gcm_dak_cmd_in[113]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[112] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[112]), .Q(gcm_dak_cmd_in[112]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[111] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[111]), .Q(gcm_dak_cmd_in[111]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[110] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[110]), .Q(gcm_dak_cmd_in[110]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[109] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[109]), .Q(gcm_dak_cmd_in[109]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[108] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[108]), .Q(gcm_dak_cmd_in[108]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[107] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[107]), .Q(gcm_dak_cmd_in[107]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[106] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[106]), .Q(gcm_dak_cmd_in[106]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[105] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[105]), .Q(gcm_dak_cmd_in[105]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[104] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[104]), .Q(gcm_dak_cmd_in[104]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[103] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[103]), .Q(gcm_dak_cmd_in[103]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[102] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[102]), .Q(gcm_dak_cmd_in[102]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[101] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[101]), .Q(gcm_dak_cmd_in[101]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[100] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[100]), .Q(gcm_dak_cmd_in[100]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[99] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[99]), .Q(gcm_dak_cmd_in[99]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[98] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[98]), .Q(gcm_dak_cmd_in[98]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[97] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[97]), .Q(gcm_dak_cmd_in[97]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[96] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[96]), .Q(gcm_dak_cmd_in[96]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[95] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[95]), .Q(gcm_dak_cmd_in[95]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[94] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[94]), .Q(gcm_dak_cmd_in[94]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[93] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[93]), .Q(gcm_dak_cmd_in[93]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[92] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[92]), .Q(gcm_dak_cmd_in[92]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[91] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[91]), .Q(gcm_dak_cmd_in[91]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[90] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[90]), .Q(gcm_dak_cmd_in[90]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[89] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[89]), .Q(gcm_dak_cmd_in[89]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[88] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[88]), .Q(gcm_dak_cmd_in[88]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[87] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[87]), .Q(gcm_dak_cmd_in[87]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[86] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[86]), .Q(gcm_dak_cmd_in[86]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[85] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[85]), .Q(gcm_dak_cmd_in[85]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[84] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[84]), .Q(gcm_dak_cmd_in[84]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[83] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[83]), .Q(gcm_dak_cmd_in[83]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[82] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[82]), .Q(gcm_dak_cmd_in[82]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[81] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[81]), .Q(gcm_dak_cmd_in[81]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[80] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[80]), .Q(gcm_dak_cmd_in[80]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[79] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[79]), .Q(gcm_dak_cmd_in[79]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[78] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[78]), .Q(gcm_dak_cmd_in[78]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[77] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[77]), .Q(gcm_dak_cmd_in[77]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[76] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[76]), .Q(gcm_dak_cmd_in[76]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[75] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[75]), .Q(gcm_dak_cmd_in[75]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[74] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[74]), .Q(gcm_dak_cmd_in[74]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[73] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[73]), .Q(gcm_dak_cmd_in[73]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[72] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[72]), .Q(gcm_dak_cmd_in[72]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[71] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[71]), .Q(gcm_dak_cmd_in[71]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[70] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[70]), .Q(gcm_dak_cmd_in[70]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[69] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[69]), .Q(gcm_dak_cmd_in[69]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[68] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[68]), .Q(gcm_dak_cmd_in[68]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[67] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[67]), .Q(gcm_dak_cmd_in[67]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[66] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[66]), .Q(gcm_dak_cmd_in[66]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[65] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[65]), .Q(gcm_dak_cmd_in[65]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[64] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[64]), .Q(gcm_dak_cmd_in[64]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[63] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[63]), .Q(gcm_dak_cmd_in[63]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[62] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[62]), .Q(gcm_dak_cmd_in[62]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[61] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[61]), .Q(gcm_dak_cmd_in[61]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[60] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[60]), .Q(gcm_dak_cmd_in[60]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[59] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[59]), .Q(gcm_dak_cmd_in[59]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[58] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[58]), .Q(gcm_dak_cmd_in[58]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[57] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[57]), .Q(gcm_dak_cmd_in[57]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[56] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[56]), .Q(gcm_dak_cmd_in[56]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[55] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[55]), .Q(gcm_dak_cmd_in[55]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[54] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[54]), .Q(gcm_dak_cmd_in[54]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[53] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[53]), .Q(gcm_dak_cmd_in[53]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[52] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[52]), .Q(gcm_dak_cmd_in[52]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[51] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[51]), .Q(gcm_dak_cmd_in[51]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[50] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[50]), .Q(gcm_dak_cmd_in[50]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[49] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[49]), .Q(gcm_dak_cmd_in[49]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[48] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[48]), .Q(gcm_dak_cmd_in[48]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[47] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[47]), .Q(gcm_dak_cmd_in[47]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[46] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[46]), .Q(gcm_dak_cmd_in[46]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[45] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[45]), .Q(gcm_dak_cmd_in[45]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[44] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[44]), .Q(gcm_dak_cmd_in[44]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[43] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[43]), .Q(gcm_dak_cmd_in[43]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[42] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[42]), .Q(gcm_dak_cmd_in[42]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[41] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[41]), .Q(gcm_dak_cmd_in[41]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[40] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[40]), .Q(gcm_dak_cmd_in[40]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[39] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[39]), .Q(gcm_dak_cmd_in[39]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[38] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[38]), .Q(gcm_dak_cmd_in[38]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[37] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[37]), .Q(gcm_dak_cmd_in[37]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[36] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[36]), .Q(gcm_dak_cmd_in[36]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[35] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[35]), .Q(gcm_dak_cmd_in[35]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[34] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[34]), .Q(gcm_dak_cmd_in[34]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[33] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[33]), .Q(gcm_dak_cmd_in[33]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[32] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[32]), .Q(gcm_dak_cmd_in[32]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[31] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[31]), .Q(gcm_dak_cmd_in[31]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[30] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[30]), .Q(gcm_dak_cmd_in[30]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[29] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[29]), .Q(gcm_dak_cmd_in[29]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[28] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[28]), .Q(gcm_dak_cmd_in[28]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[27] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[27]), .Q(gcm_dak_cmd_in[27]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[26] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[26]), .Q(gcm_dak_cmd_in[26]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[25] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[25]), .Q(gcm_dak_cmd_in[25]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[24] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[24]), .Q(gcm_dak_cmd_in[24]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[23] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[23]), .Q(gcm_dak_cmd_in[23]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[22] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[22]), .Q(gcm_dak_cmd_in[22]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[21] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[21]), .Q(gcm_dak_cmd_in[21]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[20] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[20]), .Q(gcm_dak_cmd_in[20]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[19] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[19]), .Q(gcm_dak_cmd_in[19]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[18] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[18]), .Q(gcm_dak_cmd_in[18]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[17] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[17]), .Q(gcm_dak_cmd_in[17]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[16] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[16]), .Q(gcm_dak_cmd_in[16]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[15] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[15]), .Q(gcm_dak_cmd_in[15]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[14] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[14]), .Q(gcm_dak_cmd_in[14]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[13] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[13]), .Q(gcm_dak_cmd_in[13]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[12] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[12]), .Q(gcm_dak_cmd_in[12]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[11] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[11]), .Q(gcm_dak_cmd_in[11]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[10] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[10]), .Q(gcm_dak_cmd_in[10]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[9] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[9]), .Q(gcm_dak_cmd_in[9]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[8] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[8]), .Q(gcm_dak_cmd_in[8]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[7] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[7]), .Q(gcm_dak_cmd_in[7]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[6] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[6]), .Q(gcm_dak_cmd_in[6]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[5] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[5]), .Q(gcm_dak_cmd_in[5]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[4] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[4]), .Q(gcm_dak_cmd_in[4]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[3] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[3]), .Q(gcm_dak_cmd_in[3]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[2] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[2]), .Q(gcm_dak_cmd_in[2]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[1] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[1]), .Q(gcm_dak_cmd_in[1]), .QN( ));
Q_FDP1 \gcm_dak_cmd_in_REG[0] ( .CK(clk), .R(rst_n), .D(gcm_dak_cmd_in_nxt[0]), .Q(gcm_dak_cmd_in[0]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[95] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[95]), .Q(gcm_dek_tag[95]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[94] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[94]), .Q(gcm_dek_tag[94]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[93] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[93]), .Q(gcm_dek_tag[93]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[92] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[92]), .Q(gcm_dek_tag[92]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[91] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[91]), .Q(gcm_dek_tag[91]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[90] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[90]), .Q(gcm_dek_tag[90]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[89] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[89]), .Q(gcm_dek_tag[89]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[88] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[88]), .Q(gcm_dek_tag[88]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[87] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[87]), .Q(gcm_dek_tag[87]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[86] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[86]), .Q(gcm_dek_tag[86]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[85] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[85]), .Q(gcm_dek_tag[85]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[84] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[84]), .Q(gcm_dek_tag[84]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[83] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[83]), .Q(gcm_dek_tag[83]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[82] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[82]), .Q(gcm_dek_tag[82]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[81] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[81]), .Q(gcm_dek_tag[81]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[80] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[80]), .Q(gcm_dek_tag[80]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[79] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[79]), .Q(gcm_dek_tag[79]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[78] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[78]), .Q(gcm_dek_tag[78]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[77] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[77]), .Q(gcm_dek_tag[77]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[76] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[76]), .Q(gcm_dek_tag[76]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[75] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[75]), .Q(gcm_dek_tag[75]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[74] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[74]), .Q(gcm_dek_tag[74]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[73] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[73]), .Q(gcm_dek_tag[73]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[72] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[72]), .Q(gcm_dek_tag[72]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[71] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[71]), .Q(gcm_dek_tag[71]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[70] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[70]), .Q(gcm_dek_tag[70]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[69] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[69]), .Q(gcm_dek_tag[69]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[68] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[68]), .Q(gcm_dek_tag[68]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[67] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[67]), .Q(gcm_dek_tag[67]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[66] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[66]), .Q(gcm_dek_tag[66]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[65] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[65]), .Q(gcm_dek_tag[65]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[64] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[64]), .Q(gcm_dek_tag[64]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[63] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[63]), .Q(gcm_dek_tag[63]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[62] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[62]), .Q(gcm_dek_tag[62]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[61] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[61]), .Q(gcm_dek_tag[61]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[60] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[60]), .Q(gcm_dek_tag[60]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[59] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[59]), .Q(gcm_dek_tag[59]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[58] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[58]), .Q(gcm_dek_tag[58]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[57] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[57]), .Q(gcm_dek_tag[57]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[56] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[56]), .Q(gcm_dek_tag[56]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[55] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[55]), .Q(gcm_dek_tag[55]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[54] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[54]), .Q(gcm_dek_tag[54]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[53] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[53]), .Q(gcm_dek_tag[53]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[52] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[52]), .Q(gcm_dek_tag[52]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[51] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[51]), .Q(gcm_dek_tag[51]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[50] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[50]), .Q(gcm_dek_tag[50]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[49] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[49]), .Q(gcm_dek_tag[49]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[48] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[48]), .Q(gcm_dek_tag[48]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[47] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[47]), .Q(gcm_dek_tag[47]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[46] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[46]), .Q(gcm_dek_tag[46]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[45] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[45]), .Q(gcm_dek_tag[45]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[44] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[44]), .Q(gcm_dek_tag[44]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[43] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[43]), .Q(gcm_dek_tag[43]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[42] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[42]), .Q(gcm_dek_tag[42]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[41] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[41]), .Q(gcm_dek_tag[41]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[40] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[40]), .Q(gcm_dek_tag[40]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[39] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[39]), .Q(gcm_dek_tag[39]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[38] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[38]), .Q(gcm_dek_tag[38]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[37] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[37]), .Q(gcm_dek_tag[37]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[36] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[36]), .Q(gcm_dek_tag[36]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[35] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[35]), .Q(gcm_dek_tag[35]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[34] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[34]), .Q(gcm_dek_tag[34]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[33] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[33]), .Q(gcm_dek_tag[33]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[32] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[32]), .Q(gcm_dek_tag[32]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[31] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[31]), .Q(gcm_dek_tag[31]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[30] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[30]), .Q(gcm_dek_tag[30]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[29] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[29]), .Q(gcm_dek_tag[29]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[28] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[28]), .Q(gcm_dek_tag[28]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[27] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[27]), .Q(gcm_dek_tag[27]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[26] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[26]), .Q(gcm_dek_tag[26]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[25] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[25]), .Q(gcm_dek_tag[25]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[24] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[24]), .Q(gcm_dek_tag[24]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[23] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[23]), .Q(gcm_dek_tag[23]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[22] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[22]), .Q(gcm_dek_tag[22]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[21] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[21]), .Q(gcm_dek_tag[21]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[20] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[20]), .Q(gcm_dek_tag[20]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[19] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[19]), .Q(gcm_dek_tag[19]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[18] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[18]), .Q(gcm_dek_tag[18]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[17] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[17]), .Q(gcm_dek_tag[17]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[16] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[16]), .Q(gcm_dek_tag[16]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[15] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[15]), .Q(gcm_dek_tag[15]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[14] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[14]), .Q(gcm_dek_tag[14]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[13] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[13]), .Q(gcm_dek_tag[13]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[12] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[12]), .Q(gcm_dek_tag[12]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[11] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[11]), .Q(gcm_dek_tag[11]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[10] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[10]), .Q(gcm_dek_tag[10]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[9] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[9]), .Q(gcm_dek_tag[9]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[8] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[8]), .Q(gcm_dek_tag[8]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[7] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[7]), .Q(gcm_dek_tag[7]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[6] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[6]), .Q(gcm_dek_tag[6]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[5] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[5]), .Q(gcm_dek_tag[5]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[4] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[4]), .Q(gcm_dek_tag[4]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[3] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[3]), .Q(gcm_dek_tag[3]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[2] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[2]), .Q(gcm_dek_tag[2]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[1] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[1]), .Q(gcm_dek_tag[1]), .QN( ));
Q_FDP1 \gcm_dek_tag_REG[0] ( .CK(clk), .R(rst_n), .D(gcm_dek_tag_nxt[0]), .Q(gcm_dek_tag[0]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[95] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[95]), .Q(gcm_dak_tag[95]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[94] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[94]), .Q(gcm_dak_tag[94]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[93] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[93]), .Q(gcm_dak_tag[93]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[92] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[92]), .Q(gcm_dak_tag[92]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[91] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[91]), .Q(gcm_dak_tag[91]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[90] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[90]), .Q(gcm_dak_tag[90]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[89] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[89]), .Q(gcm_dak_tag[89]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[88] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[88]), .Q(gcm_dak_tag[88]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[87] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[87]), .Q(gcm_dak_tag[87]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[86] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[86]), .Q(gcm_dak_tag[86]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[85] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[85]), .Q(gcm_dak_tag[85]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[84] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[84]), .Q(gcm_dak_tag[84]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[83] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[83]), .Q(gcm_dak_tag[83]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[82] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[82]), .Q(gcm_dak_tag[82]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[81] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[81]), .Q(gcm_dak_tag[81]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[80] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[80]), .Q(gcm_dak_tag[80]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[79] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[79]), .Q(gcm_dak_tag[79]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[78] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[78]), .Q(gcm_dak_tag[78]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[77] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[77]), .Q(gcm_dak_tag[77]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[76] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[76]), .Q(gcm_dak_tag[76]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[75] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[75]), .Q(gcm_dak_tag[75]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[74] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[74]), .Q(gcm_dak_tag[74]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[73] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[73]), .Q(gcm_dak_tag[73]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[72] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[72]), .Q(gcm_dak_tag[72]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[71] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[71]), .Q(gcm_dak_tag[71]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[70] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[70]), .Q(gcm_dak_tag[70]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[69] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[69]), .Q(gcm_dak_tag[69]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[68] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[68]), .Q(gcm_dak_tag[68]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[67] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[67]), .Q(gcm_dak_tag[67]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[66] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[66]), .Q(gcm_dak_tag[66]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[65] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[65]), .Q(gcm_dak_tag[65]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[64] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[64]), .Q(gcm_dak_tag[64]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[63] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[63]), .Q(gcm_dak_tag[63]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[62] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[62]), .Q(gcm_dak_tag[62]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[61] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[61]), .Q(gcm_dak_tag[61]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[60] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[60]), .Q(gcm_dak_tag[60]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[59] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[59]), .Q(gcm_dak_tag[59]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[58] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[58]), .Q(gcm_dak_tag[58]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[57] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[57]), .Q(gcm_dak_tag[57]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[56] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[56]), .Q(gcm_dak_tag[56]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[55] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[55]), .Q(gcm_dak_tag[55]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[54] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[54]), .Q(gcm_dak_tag[54]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[53] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[53]), .Q(gcm_dak_tag[53]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[52] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[52]), .Q(gcm_dak_tag[52]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[51] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[51]), .Q(gcm_dak_tag[51]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[50] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[50]), .Q(gcm_dak_tag[50]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[49] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[49]), .Q(gcm_dak_tag[49]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[48] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[48]), .Q(gcm_dak_tag[48]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[47] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[47]), .Q(gcm_dak_tag[47]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[46] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[46]), .Q(gcm_dak_tag[46]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[45] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[45]), .Q(gcm_dak_tag[45]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[44] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[44]), .Q(gcm_dak_tag[44]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[43] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[43]), .Q(gcm_dak_tag[43]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[42] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[42]), .Q(gcm_dak_tag[42]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[41] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[41]), .Q(gcm_dak_tag[41]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[40] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[40]), .Q(gcm_dak_tag[40]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[39] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[39]), .Q(gcm_dak_tag[39]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[38] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[38]), .Q(gcm_dak_tag[38]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[37] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[37]), .Q(gcm_dak_tag[37]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[36] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[36]), .Q(gcm_dak_tag[36]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[35] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[35]), .Q(gcm_dak_tag[35]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[34] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[34]), .Q(gcm_dak_tag[34]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[33] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[33]), .Q(gcm_dak_tag[33]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[32] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[32]), .Q(gcm_dak_tag[32]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[31] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[31]), .Q(gcm_dak_tag[31]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[30] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[30]), .Q(gcm_dak_tag[30]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[29] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[29]), .Q(gcm_dak_tag[29]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[28] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[28]), .Q(gcm_dak_tag[28]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[27] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[27]), .Q(gcm_dak_tag[27]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[26] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[26]), .Q(gcm_dak_tag[26]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[25] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[25]), .Q(gcm_dak_tag[25]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[24] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[24]), .Q(gcm_dak_tag[24]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[23] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[23]), .Q(gcm_dak_tag[23]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[22] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[22]), .Q(gcm_dak_tag[22]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[21] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[21]), .Q(gcm_dak_tag[21]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[20] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[20]), .Q(gcm_dak_tag[20]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[19] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[19]), .Q(gcm_dak_tag[19]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[18] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[18]), .Q(gcm_dak_tag[18]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[17] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[17]), .Q(gcm_dak_tag[17]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[16] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[16]), .Q(gcm_dak_tag[16]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[15] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[15]), .Q(gcm_dak_tag[15]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[14] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[14]), .Q(gcm_dak_tag[14]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[13] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[13]), .Q(gcm_dak_tag[13]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[12] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[12]), .Q(gcm_dak_tag[12]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[11] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[11]), .Q(gcm_dak_tag[11]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[10] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[10]), .Q(gcm_dak_tag[10]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[9] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[9]), .Q(gcm_dak_tag[9]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[8] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[8]), .Q(gcm_dak_tag[8]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[7] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[7]), .Q(gcm_dak_tag[7]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[6] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[6]), .Q(gcm_dak_tag[6]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[5] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[5]), .Q(gcm_dak_tag[5]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[4] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[4]), .Q(gcm_dak_tag[4]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[3] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[3]), .Q(gcm_dak_tag[3]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[2] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[2]), .Q(gcm_dak_tag[2]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[1] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[1]), .Q(gcm_dak_tag[1]), .QN( ));
Q_FDP1 \gcm_dak_tag_REG[0] ( .CK(clk), .R(rst_n), .D(gcm_dak_tag_nxt[0]), .Q(gcm_dak_tag[0]), .QN( ));
Q_FDP1 skip_dek_kdf_REG  ( .CK(clk), .R(rst_n), .D(skip_dek_kdf_nxt), .Q(skip_dek_kdf), .QN( ));
Q_FDP1 skip_dak_kdf_REG  ( .CK(clk), .R(rst_n), .D(skip_dak_kdf_nxt), .Q(skip_dak_kdf), .QN( ));
Q_FDP1 kdf_dek_iter_REG  ( .CK(clk), .R(rst_n), .D(kdf_dek_iter_nxt), .Q(kdf_dek_iter), .QN( ));
Q_AN02 U7580 ( .A0(rst_n), .A1(_zy_sva_b32), .Z(n2765));
Q_AN02 U7581 ( .A0(rst_n), .A1(_zy_sva_b31), .Z(n2766));
Q_AN02 U7582 ( .A0(rst_n), .A1(_zy_sva_b30), .Z(n2767));
Q_AN02 U7583 ( .A0(rst_n), .A1(_zy_sva_b29), .Z(n2768));
Q_AN02 U7584 ( .A0(rst_n), .A1(_zy_sva_b28), .Z(n2769));
Q_AN02 U7585 ( .A0(rst_n), .A1(_zy_sva_b27), .Z(n2770));
Q_AN02 U7586 ( .A0(rst_n), .A1(_zy_sva_b26), .Z(n2771));
Q_AN02 U7587 ( .A0(rst_n), .A1(_zy_sva_b25), .Z(n2772));
Q_AN02 U7588 ( .A0(rst_n), .A1(_zy_sva_b24), .Z(n2773));
Q_AN02 U7589 ( .A0(rst_n), .A1(_zy_sva_b23), .Z(n2774));
Q_AN02 U7590 ( .A0(rst_n), .A1(_zy_sva_b22), .Z(n2775));
Q_AN02 U7591 ( .A0(rst_n), .A1(_zy_sva_b21), .Z(n2776));
Q_AN02 U7592 ( .A0(rst_n), .A1(_zy_sva_b20), .Z(n2777));
Q_AN02 U7593 ( .A0(rst_n), .A1(_zy_sva_b19), .Z(n2778));
Q_AN02 U7594 ( .A0(rst_n), .A1(_zy_sva_b18), .Z(n2779));
Q_AN02 U7595 ( .A0(rst_n), .A1(_zy_sva_b17), .Z(n2780));
Q_AN02 U7596 ( .A0(rst_n), .A1(_zy_sva_b16), .Z(n2781));
Q_AN02 U7597 ( .A0(rst_n), .A1(_zy_sva_b15), .Z(n2782));
Q_AN02 U7598 ( .A0(rst_n), .A1(_zy_sva_b14), .Z(n2783));
Q_AN02 U7599 ( .A0(rst_n), .A1(_zy_sva_b13), .Z(n2784));
Q_AN02 U7600 ( .A0(rst_n), .A1(_zy_sva_b12), .Z(n2785));
Q_AN02 U7601 ( .A0(rst_n), .A1(_zy_sva_b11), .Z(n2786));
Q_AN02 U7602 ( .A0(rst_n), .A1(_zy_sva_b10), .Z(n2787));
Q_AN02 U7603 ( .A0(rst_n), .A1(_zy_sva_b9), .Z(n2788));
Q_AN02 U7604 ( .A0(rst_n), .A1(_zy_sva_b8), .Z(n2789));
Q_AN02 U7605 ( .A0(rst_n), .A1(_zy_sva_b7), .Z(n2790));
Q_AN02 U7606 ( .A0(rst_n), .A1(_zy_sva_b6), .Z(n2791));
Q_AN02 U7607 ( .A0(rst_n), .A1(_zy_sva_b5), .Z(n2792));
Q_AN02 U7608 ( .A0(rst_n), .A1(_zy_sva_b4), .Z(n2793));
Q_AN02 U7609 ( .A0(rst_n), .A1(_zy_sva_b3), .Z(n2794));
Q_AN02 U7610 ( .A0(rst_n), .A1(_zy_sva_b2), .Z(n2795));
Q_AN02 U7611 ( .A0(rst_n), .A1(_zy_sva_b1), .Z(n2796));
Q_AN02 U7612 ( .A0(rst_n), .A1(_zy_sva_b0), .Z(n2797));
ixc_assign _zz_strnp_0 ( _zy_simnet_kme_internal_out_ack_0_w$, 
	kme_internal_out_ack);
ixc_assign_611 _zz_strnp_1 ( _zy_simnet_gcm_cmd_in_1_w$[0:610], 
	gcm_cmd_in[610:0]);
ixc_assign _zz_strnp_2 ( _zy_simnet_gcm_cmd_in_valid_2_w$, gcm_cmd_in_valid);
ixc_assign_96 _zz_strnp_3 ( _zy_simnet_gcm_tag_data_in_3_w$[0:95], 
	gcm_tag_data_in[95:0]);
ixc_assign _zz_strnp_4 ( _zy_simnet_gcm_tag_data_in_valid_4_w$, 
	gcm_tag_data_in_valid);
ixc_assign _zz_strnp_5 ( _zy_simnet_inspector_upsizer_valid_5_w$, 
	inspector_upsizer_valid);
ixc_assign _zz_strnp_6 ( _zy_simnet_inspector_upsizer_eof_6_w$, 
	inspector_upsizer_eof);
ixc_assign_64 _zz_strnp_7 ( _zy_simnet_inspector_upsizer_data_7_w$[0:63], 
	inspector_upsizer_data[63:0]);
ixc_assign _zz_strnp_8 ( _zy_simnet_keyfilter_cmd_in_8_w$, 
	keyfilter_cmd_in[0]);
ixc_assign _zz_strnp_9 ( _zy_simnet_keyfilter_cmd_in_valid_9_w$, 
	keyfilter_cmd_in_valid);
ixc_assign_263 _zz_strnp_10 ( _zy_simnet_kdfstream_cmd_in_10_w$[0:262], 
	kdfstream_cmd_in[262:0]);
ixc_assign _zz_strnp_11 ( _zy_simnet_kdfstream_cmd_in_valid_11_w$, 
	kdfstream_cmd_in_valid);
ixc_assign_4 _zz_strnp_12 ( _zy_simnet_kdf_cmd_in_12_w$[0:3], { kdf_cmd_in[3], 
	keyfilter_cmd_in[0], kdf_cmd_in[1], kdf_cmd_in[0]});
ixc_assign _zz_strnp_13 ( _zy_simnet_kdf_cmd_in_valid_13_w$, 
	keyfilter_cmd_in_valid);
ixc_assign_64 _zz_strnp_14 ( _zy_simnet_tlv_sb_data_in_14_w$[0:63], 
	tlv_sb_data_in[63:0]);
ixc_assign _zz_strnp_15 ( _zy_simnet_tlv_sb_data_in_valid_15_w$, 
	tlv_sb_data_in_valid);
Q_INV U7629 ( .A(rst_n), .Z(_zy_sva_brcm_gcm_dek256_with_512bit_key_1_reset_or));
Q_INV U7630 ( .A(gcm_cmd_in[1]), .Z(n2848));
Q_AN03 U7631 ( .A0(gcm_cmd_in_valid), .A1(n2846), .A2(n2840), .Z(_zy_sva_b0_t));
Q_INV U7632 ( .A(gcm_cmd_in[2]), .Z(n2847));
Q_AN03 U7633 ( .A0(gcm_cmd_in_valid), .A1(n2846), .A2(n2839), .Z(_zy_sva_b1_t));
Q_AN03 U7634 ( .A0(gcm_cmd_in_valid), .A1(n2846), .A2(n2837), .Z(_zy_sva_b2_t));
Q_AN02 U7635 ( .A0(n2849), .A1(dek_ckv_length_q[1]), .Z(n2846));
Q_INV U7636 ( .A(gcm_cmd_in[0]), .Z(n2845));
Q_AN03 U7637 ( .A0(gcm_cmd_in_valid), .A1(n2846), .A2(n2836), .Z(_zy_sva_b3_t));
Q_NR03 U7638 ( .A0(n42), .A1(kek_tag_q), .A2(n2841), .Z(_zy_sva_b4_t));
Q_AN03 U7639 ( .A0(gcm_cmd_in_valid), .A1(n2844), .A2(n2839), .Z(_zy_sva_b5_t));
Q_AN03 U7640 ( .A0(gcm_cmd_in_valid), .A1(n2844), .A2(n2837), .Z(_zy_sva_b6_t));
Q_AN03 U7641 ( .A0(gcm_cmd_in_valid), .A1(n2844), .A2(n2836), .Z(_zy_sva_b7_t));
Q_OR03 U7642 ( .A0(gcm_cmd_in[0]), .A1(gcm_cmd_in[1]), .A2(gcm_cmd_in[2]), .Z(n2843));
Q_NR02 U7643 ( .A0(n42), .A1(n2843), .Z(_zy_sva_b9_t));
Q_OR03 U7644 ( .A0(n2845), .A1(gcm_cmd_in[1]), .A2(gcm_cmd_in[2]), .Z(n2842));
Q_NR02 U7645 ( .A0(n42), .A1(n2842), .Z(_zy_sva_b10_t));
Q_OR03 U7646 ( .A0(gcm_cmd_in[0]), .A1(n2848), .A2(gcm_cmd_in[2]), .Z(n2841));
Q_INV U7647 ( .A(n2841), .Z(n2840));
Q_NR02 U7648 ( .A0(n42), .A1(n2841), .Z(_zy_sva_b11_t));
Q_AN03 U7649 ( .A0(gcm_cmd_in[0]), .A1(gcm_cmd_in[1]), .A2(n2847), .Z(n2839));
Q_AN02 U7650 ( .A0(gcm_cmd_in_valid), .A1(n2839), .Z(_zy_sva_b12_t));
Q_OR03 U7651 ( .A0(gcm_cmd_in[0]), .A1(gcm_cmd_in[1]), .A2(n2847), .Z(n2838));
Q_NR02 U7652 ( .A0(n42), .A1(n2838), .Z(_zy_sva_b13_t));
Q_AN03 U7653 ( .A0(gcm_cmd_in[0]), .A1(n2848), .A2(gcm_cmd_in[2]), .Z(n2837));
Q_AN02 U7654 ( .A0(gcm_cmd_in_valid), .A1(n2837), .Z(_zy_sva_b14_t));
Q_AN03 U7655 ( .A0(n2845), .A1(gcm_cmd_in[1]), .A2(gcm_cmd_in[2]), .Z(n2836));
Q_AN02 U7656 ( .A0(gcm_cmd_in_valid), .A1(n2836), .Z(_zy_sva_b15_t));
Q_AN03 U7657 ( .A0(gcm_cmd_in[0]), .A1(gcm_cmd_in[1]), .A2(gcm_cmd_in[2]), .Z(n2835));
Q_AN02 U7658 ( .A0(gcm_cmd_in_valid), .A1(n2835), .Z(_zy_sva_b16_t));
Q_AN02 U7659 ( .A0(n2834), .A1(n2827), .Z(_zy_sva_b17_t));
Q_AN03 U7660 ( .A0(n2834), .A1(n2823), .A2(n2819), .Z(_zy_sva_b18_t));
Q_AN03 U7661 ( .A0(n2834), .A1(n2816), .A2(n2812), .Z(_zy_sva_b19_t));
Q_NR03 U7662 ( .A0(n9), .A1(n2), .A2(n54), .Z(n2834));
Q_AN03 U7663 ( .A0(n2834), .A1(n2804), .A2(n2799), .Z(_zy_sva_b20_t));
Q_AN02 U7664 ( .A0(n2832), .A1(n2827), .Z(_zy_sva_b21_t));
Q_AN03 U7665 ( .A0(n2832), .A1(n2823), .A2(n2819), .Z(_zy_sva_b22_t));
Q_AN03 U7666 ( .A0(n2832), .A1(n2816), .A2(n2812), .Z(_zy_sva_b23_t));
Q_INV U7667 ( .A(n2), .Z(n2833));
Q_AN03 U7668 ( .A0(n9), .A1(n2833), .A2(kdfstream_cmd_in_valid), .Z(n2832));
Q_AN03 U7669 ( .A0(n2832), .A1(n2804), .A2(n2799), .Z(_zy_sva_b24_t));
Q_AN02 U7670 ( .A0(n2830), .A1(n2827), .Z(_zy_sva_b25_t));
Q_AN03 U7671 ( .A0(n2830), .A1(n2823), .A2(n2819), .Z(_zy_sva_b26_t));
Q_AN03 U7672 ( .A0(n2830), .A1(n2816), .A2(n2812), .Z(_zy_sva_b27_t));
Q_INV U7673 ( .A(n9), .Z(n2831));
Q_AN03 U7674 ( .A0(n2831), .A1(n2), .A2(kdfstream_cmd_in_valid), .Z(n2830));
Q_AN03 U7675 ( .A0(n2830), .A1(n2804), .A2(n2799), .Z(_zy_sva_b28_t));
Q_AO21 U7676 ( .A0(n5), .A1(n6), .B0(n2854), .Z(n2829));
Q_AO21 U7677 ( .A0(n5), .A1(n2801), .B0(n2829), .Z(n2828));
Q_INV U7678 ( .A(n2828), .Z(n2827));
Q_AN02 U7679 ( .A0(n2798), .A1(n2827), .Z(_zy_sva_b29_t));
Q_AN02 U7680 ( .A0(n2808), .A1(n2811), .Z(n2826));
Q_AN02 U7681 ( .A0(n2808), .A1(n2810), .Z(n2825));
Q_AO21 U7682 ( .A0(n2825), .A1(n2855), .B0(n2826), .Z(n2824));
Q_INV U7683 ( .A(n2824), .Z(n2823));
Q_AN02 U7684 ( .A0(n4), .A1(n6), .Z(n2822));
Q_OR03 U7685 ( .A0(n2815), .A1(n2822), .A2(n3), .Z(n2821));
Q_AO21 U7686 ( .A0(n4), .A1(n2801), .B0(n2821), .Z(n2820));
Q_INV U7687 ( .A(n2820), .Z(n2819));
Q_AN03 U7688 ( .A0(n2798), .A1(n2823), .A2(n2819), .Z(_zy_sva_b30_t));
Q_AN02 U7689 ( .A0(n2809), .A1(n2810), .Z(n2818));
Q_AO21 U7690 ( .A0(n2818), .A1(n2855), .B0(n2808), .Z(n2817));
Q_INV U7691 ( .A(n2817), .Z(n2816));
Q_AN02 U7692 ( .A0(n4), .A1(n5), .Z(n2815));
Q_AO21 U7693 ( .A0(n2815), .A1(n6), .B0(n3), .Z(n2814));
Q_AO21 U7694 ( .A0(n2815), .A1(n2801), .B0(n2814), .Z(n2813));
Q_INV U7695 ( .A(n2813), .Z(n2812));
Q_AN03 U7696 ( .A0(n2798), .A1(n2816), .A2(n2812), .Z(_zy_sva_b31_t));
Q_INV U7697 ( .A(n5), .Z(n2811));
Q_INV U7698 ( .A(n6), .Z(n2810));
Q_NR02 U7699 ( .A0(n3), .A1(n5), .Z(n2809));
Q_NR02 U7700 ( .A0(n3), .A1(n4), .Z(n2808));
Q_OR02 U7701 ( .A0(n2808), .A1(n2809), .Z(n2807));
Q_NR02 U7702 ( .A0(n3), .A1(n6), .Z(n2806));
Q_AO21 U7703 ( .A0(n2806), .A1(n2855), .B0(n2807), .Z(n2805));
Q_INV U7704 ( .A(n2805), .Z(n2804));
Q_OR02 U7705 ( .A0(n5), .A1(n6), .Z(n2803));
Q_OA21 U7706 ( .A0(n4), .A1(n2803), .B0(n3), .Z(n2802));
Q_AO21 U7707 ( .A0(n3), .A1(n2801), .B0(n2802), .Z(n2800));
Q_INV U7708 ( .A(n2800), .Z(n2799));
Q_AN03 U7709 ( .A0(n9), .A1(n2), .A2(kdfstream_cmd_in_valid), .Z(n2798));
Q_AN03 U7710 ( .A0(n2798), .A1(n2804), .A2(n2799), .Z(_zy_sva_b32_t));
ixc_sample_logic_1_3 _zz_zy_sva_b0 ( _zy_sva_b0, _zy_sva_b0_t);
ixc_sample_logic_1_3 _zz_zy_sva_b1 ( _zy_sva_b1, _zy_sva_b1_t);
ixc_sample_logic_1_3 _zz_zy_sva_b2 ( _zy_sva_b2, _zy_sva_b2_t);
ixc_sample_logic_1_3 _zz_zy_sva_b3 ( _zy_sva_b3, _zy_sva_b3_t);
ixc_sample_logic_1_3 _zz_zy_sva_b4 ( _zy_sva_b4, _zy_sva_b4_t);
ixc_sample_logic_1_3 _zz_zy_sva_b5 ( _zy_sva_b5, _zy_sva_b5_t);
ixc_sample_logic_1_3 _zz_zy_sva_b6 ( _zy_sva_b6, _zy_sva_b6_t);
ixc_sample_logic_1_3 _zz_zy_sva_b7 ( _zy_sva_b7, _zy_sva_b7_t);
ixc_sample_logic_1_3 _zz_zy_sva_b8 ( _zy_sva_b8, _zy_sva_b8_t);
ixc_sample_logic_1_3 _zz_zy_sva_b9 ( _zy_sva_b9, _zy_sva_b9_t);
ixc_sample_logic_1_3 _zz_zy_sva_b10 ( _zy_sva_b10, _zy_sva_b10_t);
ixc_sample_logic_1_3 _zz_zy_sva_b11 ( _zy_sva_b11, _zy_sva_b11_t);
ixc_sample_logic_1_3 _zz_zy_sva_b12 ( _zy_sva_b12, _zy_sva_b12_t);
ixc_sample_logic_1_3 _zz_zy_sva_b13 ( _zy_sva_b13, _zy_sva_b13_t);
ixc_sample_logic_1_3 _zz_zy_sva_b14 ( _zy_sva_b14, _zy_sva_b14_t);
ixc_sample_logic_1_3 _zz_zy_sva_b15 ( _zy_sva_b15, _zy_sva_b15_t);
ixc_sample_logic_1_3 _zz_zy_sva_b16 ( _zy_sva_b16, _zy_sva_b16_t);
ixc_sample_logic_1_3 _zz_zy_sva_b17 ( _zy_sva_b17, _zy_sva_b17_t);
ixc_sample_logic_1_3 _zz_zy_sva_b18 ( _zy_sva_b18, _zy_sva_b18_t);
ixc_sample_logic_1_3 _zz_zy_sva_b19 ( _zy_sva_b19, _zy_sva_b19_t);
ixc_sample_logic_1_3 _zz_zy_sva_b20 ( _zy_sva_b20, _zy_sva_b20_t);
ixc_sample_logic_1_3 _zz_zy_sva_b21 ( _zy_sva_b21, _zy_sva_b21_t);
ixc_sample_logic_1_3 _zz_zy_sva_b22 ( _zy_sva_b22, _zy_sva_b22_t);
ixc_sample_logic_1_3 _zz_zy_sva_b23 ( _zy_sva_b23, _zy_sva_b23_t);
ixc_sample_logic_1_3 _zz_zy_sva_b24 ( _zy_sva_b24, _zy_sva_b24_t);
ixc_sample_logic_1_3 _zz_zy_sva_b25 ( _zy_sva_b25, _zy_sva_b25_t);
ixc_sample_logic_1_3 _zz_zy_sva_b26 ( _zy_sva_b26, _zy_sva_b26_t);
ixc_sample_logic_1_3 _zz_zy_sva_b27 ( _zy_sva_b27, _zy_sva_b27_t);
ixc_sample_logic_1_3 _zz_zy_sva_b28 ( _zy_sva_b28, _zy_sva_b28_t);
ixc_sample_logic_1_3 _zz_zy_sva_b29 ( _zy_sva_b29, _zy_sva_b29_t);
ixc_sample_logic_1_3 _zz_zy_sva_b30 ( _zy_sva_b30, _zy_sva_b30_t);
ixc_sample_logic_1_3 _zz_zy_sva_b31 ( _zy_sva_b31, _zy_sva_b31_t);
ixc_sample_logic_1_3 _zz_zy_sva_b32 ( _zy_sva_b32, _zy_sva_b32_t);
wire [2:0] n2857 = 3'b000;
Q_ASSERT \op_0_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_10_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_10_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2857[0]));
// pragma CVASTRPROP INSTANCE "\op_0_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_0_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_0_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2858 = 3'b000;
Q_ASSERT \op_1_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_11_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_11_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2858[0]));
// pragma CVASTRPROP INSTANCE "\op_1_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_1_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_1_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2859 = 3'b000;
Q_ASSERT \op_2_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_12_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_12_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2859[0]));
// pragma CVASTRPROP INSTANCE "\op_2_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_2_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_2_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2860 = 3'b000;
Q_ASSERT \op_3_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_13_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_13_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2860[0]));
// pragma CVASTRPROP INSTANCE "\op_3_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_3_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_3_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2861 = 3'b000;
Q_ASSERT \op_4_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_14_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_14_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2861[0]));
// pragma CVASTRPROP INSTANCE "\op_4_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_4_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_4_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2862 = 3'b000;
Q_ASSERT \op_5_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_15_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_15_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2862[0]));
// pragma CVASTRPROP INSTANCE "\op_5_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_5_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_5_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2863 = 3'b000;
Q_ASSERT \op_6_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_16_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_16_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2863[0]));
// pragma CVASTRPROP INSTANCE "\op_6_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_6_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_6_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2864 = 3'b000;
Q_ASSERT \op_7_.brcm_gcm  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_17_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_17_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2864[0]));
// pragma CVASTRPROP INSTANCE "\op_7_.brcm_gcm " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\op_7_.brcm_gcm " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\op_7_.brcm_gcm " ASSERT_LINE 573
wire [2:0] n2865 = 3'b000;
Q_ASSERT \guid_0_.delimiter_0_.brcm_kdf_label0_8  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label0_8_18_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label0_8_18_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2865[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label0_8 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label0_8 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label0_8 " ASSERT_LINE 595
wire [2:0] n2866 = 3'b000;
Q_ASSERT \guid_0_.delimiter_0_.brcm_kdf_label9_16  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label9_16_19_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label9_16_19_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2866[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label9_16 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label9_16 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label9_16 " ASSERT_LINE 600
wire [2:0] n2867 = 3'b000;
Q_ASSERT \guid_0_.delimiter_0_.brcm_kdf_label17_24  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label17_24_20_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label17_24_20_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2867[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label17_24 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label17_24 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label17_24 " ASSERT_LINE 605
wire [2:0] n2868 = 3'b000;
Q_ASSERT \guid_0_.delimiter_0_.brcm_kdf_label25_32  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label25_32_21_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label25_32_21_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2868[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label25_32 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label25_32 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_0_.brcm_kdf_label25_32 " ASSERT_LINE 610
wire [2:0] n2869 = 3'b000;
Q_ASSERT \guid_0_.delimiter_1_.brcm_kdf_label0_8  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label0_8_22_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label0_8_22_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2869[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label0_8 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label0_8 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label0_8 " ASSERT_LINE 595
wire [2:0] n2870 = 3'b000;
Q_ASSERT \guid_0_.delimiter_1_.brcm_kdf_label9_16  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label9_16_23_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label9_16_23_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2870[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label9_16 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label9_16 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label9_16 " ASSERT_LINE 600
wire [2:0] n2871 = 3'b000;
Q_ASSERT \guid_0_.delimiter_1_.brcm_kdf_label17_24  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label17_24_24_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label17_24_24_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2871[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label17_24 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label17_24 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label17_24 " ASSERT_LINE 605
wire [2:0] n2872 = 3'b000;
Q_ASSERT \guid_0_.delimiter_1_.brcm_kdf_label25_32  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label25_32_25_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label25_32_25_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2872[0]));
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label25_32 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label25_32 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_0_.delimiter_1_.brcm_kdf_label25_32 " ASSERT_LINE 610
wire [2:0] n2873 = 3'b000;
Q_ASSERT \guid_1_.delimiter_0_.brcm_kdf_label0_8  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label0_8_26_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label0_8_26_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2873[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label0_8 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label0_8 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label0_8 " ASSERT_LINE 595
wire [2:0] n2874 = 3'b000;
Q_ASSERT \guid_1_.delimiter_0_.brcm_kdf_label9_16  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label9_16_27_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label9_16_27_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2874[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label9_16 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label9_16 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label9_16 " ASSERT_LINE 600
wire [2:0] n2875 = 3'b000;
Q_ASSERT \guid_1_.delimiter_0_.brcm_kdf_label17_24  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label17_24_28_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label17_24_28_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2875[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label17_24 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label17_24 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label17_24 " ASSERT_LINE 605
wire [2:0] n2876 = 3'b000;
Q_ASSERT \guid_1_.delimiter_0_.brcm_kdf_label25_32  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label25_32_29_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label25_32_29_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2876[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label25_32 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label25_32 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_0_.brcm_kdf_label25_32 " ASSERT_LINE 610
wire [2:0] n2877 = 3'b000;
Q_ASSERT \guid_1_.delimiter_1_.brcm_kdf_label0_8  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label0_8_30_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label0_8_30_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2877[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label0_8 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label0_8 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label0_8 " ASSERT_LINE 595
wire [2:0] n2878 = 3'b000;
Q_ASSERT \guid_1_.delimiter_1_.brcm_kdf_label9_16  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label9_16_31_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label9_16_31_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2878[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label9_16 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label9_16 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label9_16 " ASSERT_LINE 600
wire [2:0] n2879 = 3'b000;
Q_ASSERT \guid_1_.delimiter_1_.brcm_kdf_label17_24  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label17_24_32_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label17_24_32_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2879[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label17_24 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label17_24 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label17_24 " ASSERT_LINE 605
wire [2:0] n2880 = 3'b000;
Q_ASSERT \guid_1_.delimiter_1_.brcm_kdf_label25_32  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_kdf_label25_32_33_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_kdf_label25_32_33_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2880[0]));
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label25_32 " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label25_32 " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "\guid_1_.delimiter_1_.brcm_kdf_label25_32 " ASSERT_LINE 610
wire [2:0] n2881 = 3'b000;
Q_ASSERT brcm_gcm_dek256_with_512bit_key ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_dek256_with_512bit_key_1_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_dek256_with_512bit_key_1_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2881[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek256_with_512bit_key" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek256_with_512bit_key" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_dek256_with_512bit_key" ASSERT_LINE 577
wire [2:0] n2882 = 3'b000;
Q_ASSERT brcm_gcm_dek512_with_512bit_key ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_dek512_with_512bit_key_2_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_dek512_with_512bit_key_2_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2882[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek512_with_512bit_key" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek512_with_512bit_key" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_dek512_with_512bit_key" ASSERT_LINE 578
wire [2:0] n2883 = 3'b000;
Q_ASSERT brcm_gcm_dek256dak_with_512bit_key ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2883[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek256dak_with_512bit_key" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek256dak_with_512bit_key" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_dek256dak_with_512bit_key" ASSERT_LINE 579
wire [2:0] n2884 = 3'b000;
Q_ASSERT brcm_gcm_dek512dak_with_512bit_key ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2884[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek512dak_with_512bit_key" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_dek512dak_with_512bit_key" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_dek512dak_with_512bit_key" ASSERT_LINE 580
wire [2:0] n2885 = 3'b000;
Q_ASSERT brcm_gcm_enc_dek256_no_kbk ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2885[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek256_no_kbk" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek256_no_kbk" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_enc_dek256_no_kbk" ASSERT_LINE 583
wire [2:0] n2886 = 3'b000;
Q_ASSERT brcm_gcm_enc_dek512_no_kbk ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2886[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek512_no_kbk" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek512_no_kbk" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_enc_dek512_no_kbk" ASSERT_LINE 584
wire [2:0] n2887 = 3'b000;
Q_ASSERT brcm_gcm_enc_dek256_comb_no_kbk ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2887[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek256_comb_no_kbk" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek256_comb_no_kbk" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_enc_dek256_comb_no_kbk" ASSERT_LINE 585
wire [2:0] n2888 = 3'b000;
Q_ASSERT brcm_gcm_enc_dek512_comb_no_kbk ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2888[0]));
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek512_comb_no_kbk" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_gcm_enc_dek512_comb_no_kbk" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_gcm_enc_dek512_comb_no_kbk" ASSERT_LINE 586
wire [2:0] n2889 = 3'b000;
Q_ASSERT brcm_tlv_sb_stall_on_guid ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_tlv_sb_stall_on_guid_9_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_tlv_sb_stall_on_guid_9_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n2889[0]));
// pragma CVASTRPROP INSTANCE "brcm_tlv_sb_stall_on_guid" HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "brcm_tlv_sb_stall_on_guid" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_kop_tlv_inspector.v"
//pragma CVAINTPROP INSTANCE "brcm_tlv_sb_stall_on_guid" ASSERT_LINE 615
Q_INV U7777 ( .A(n2734), .Z(n2852));
Q_INV U7778 ( .A(n2720), .Z(n2853));
Q_INV U7779 ( .A(n2808), .Z(n2854));
Q_INV U7780 ( .A(n2801), .Z(n2855));
Q_FDP4EP \_zy_sva_brcm_gcm_dek256_with_512bit_key_1_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek256_with_512bit_key_1_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek256_with_512bit_key_1_cpass_REG[0] ( .CK(clk), .CE(n2797), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek256_with_512bit_key_1_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek512_with_512bit_key_2_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek512_with_512bit_key_2_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek512_with_512bit_key_2_cpass_REG[0] ( .CK(clk), .CE(n2796), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek512_with_512bit_key_2_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_cpass_REG[0] ( .CK(clk), .CE(n2795), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek256dak_with_512bit_key_3_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_cpass_REG[0] ( .CK(clk), .CE(n2794), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_dek512dak_with_512bit_key_4_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_cpass_REG[0] ( .CK(clk), .CE(n2793), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek256_no_kbk_5_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_cpass_REG[0] ( .CK(clk), .CE(n2792), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek512_no_kbk_6_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_cpass_REG[0] ( .CK(clk), .CE(n2791), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek256_comb_no_kbk_7_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_cpass_REG[0] ( .CK(clk), .CE(n2790), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_enc_dek512_comb_no_kbk_8_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_tlv_sb_stall_on_guid_9_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_tlv_sb_stall_on_guid_9_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_tlv_sb_stall_on_guid_9_cpass_REG[0] ( .CK(clk), .CE(n2789), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_tlv_sb_stall_on_guid_9_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_10_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_10_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_10_cpass_REG[0] ( .CK(clk), .CE(n2788), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_10_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_11_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_11_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_11_cpass_REG[0] ( .CK(clk), .CE(n2787), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_11_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_12_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_12_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_12_cpass_REG[0] ( .CK(clk), .CE(n2786), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_12_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_13_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_13_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_13_cpass_REG[0] ( .CK(clk), .CE(n2785), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_13_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_14_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_14_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_14_cpass_REG[0] ( .CK(clk), .CE(n2784), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_14_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_15_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_15_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_15_cpass_REG[0] ( .CK(clk), .CE(n2783), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_15_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_16_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_16_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_16_cpass_REG[0] ( .CK(clk), .CE(n2782), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_16_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_17_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_17_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_gcm_17_cpass_REG[0] ( .CK(clk), .CE(n2781), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_gcm_17_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_18_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_18_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_18_cpass_REG[0] ( .CK(clk), .CE(n2780), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_18_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_19_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_19_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_19_cpass_REG[0] ( .CK(clk), .CE(n2779), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_19_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_20_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_20_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_20_cpass_REG[0] ( .CK(clk), .CE(n2778), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_20_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_21_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_21_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_21_cpass_REG[0] ( .CK(clk), .CE(n2777), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_21_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_22_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_22_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_22_cpass_REG[0] ( .CK(clk), .CE(n2776), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_22_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_23_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_23_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_23_cpass_REG[0] ( .CK(clk), .CE(n2775), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_23_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_24_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_24_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_24_cpass_REG[0] ( .CK(clk), .CE(n2774), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_24_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_25_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_25_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_25_cpass_REG[0] ( .CK(clk), .CE(n2773), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_25_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_26_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_26_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_26_cpass_REG[0] ( .CK(clk), .CE(n2772), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_26_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_27_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_27_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_27_cpass_REG[0] ( .CK(clk), .CE(n2771), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_27_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_28_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_28_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_28_cpass_REG[0] ( .CK(clk), .CE(n2770), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_28_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_29_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_29_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_29_cpass_REG[0] ( .CK(clk), .CE(n2769), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_29_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_30_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_30_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label0_8_30_cpass_REG[0] ( .CK(clk), .CE(n2768), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label0_8_30_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_31_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_31_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label9_16_31_cpass_REG[0] ( .CK(clk), .CE(n2767), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label9_16_31_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_32_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_32_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label17_24_32_cpass_REG[0] ( .CK(clk), .CE(n2766), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label17_24_32_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_33_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_33_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_kdf_label25_32_33_cpass_REG[0] ( .CK(clk), .CE(n2765), .R(n2851), .D(n2850), .Q(_zy_sva_brcm_kdf_label25_32_33_cpass[0]));
Q_FDP4EP corrupt_kme_error_bit_0_REG  ( .CK(clk), .CE(n2742), .R(n2856), .D(n2757), .Q(corrupt_kme_error_bit_0));
Q_INV U7848 ( .A(rst_n), .Z(n2856));
Q_FDP4EP rst_corrupt_kme_error_bit_0_REG  ( .CK(clk), .CE(n2741), .R(n2856), .D(n2743), .Q(rst_corrupt_kme_error_bit_0));
Q_FDP4EP corrupt_crc32_REG  ( .CK(clk), .CE(n2740), .R(n2856), .D(n2759), .Q(corrupt_crc32));
Q_FDP4EP rst_corrupt_crc32_REG  ( .CK(clk), .CE(n2739), .R(n2856), .D(n2744), .Q(rst_corrupt_crc32));
Q_FDP4EP \dek_ckv_length_q_REG[1] ( .CK(clk), .CE(n10), .R(n2856), .D(kme_internal_out[59]), .Q(dek_ckv_length_q[1]));
Q_FDP4EP \dek_ckv_length_q_REG[0] ( .CK(clk), .CE(n10), .R(n2856), .D(kme_internal_out[58]), .Q(dek_ckv_length_q[0]));
Q_INV U7854 ( .A(dek_ckv_length_q[0]), .Z(n2849));
Q_FDP4EP kek_tag_q_REG  ( .CK(clk), .CE(n10), .R(n2856), .D(kme_internal_out[15]), .Q(kek_tag_q));
Q_INV U7856 ( .A(kek_tag_q), .Z(n2844));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\gcm_cmd_in.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\gcm_cmd_in.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\gcm_cmd_in.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\gcm_cmd_in.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\keyfilter_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\kdfstream_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\kdfstream_cmd_in.skip  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\kdfstream_cmd_in.guid  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\kdfstream_cmd_in.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\kdfstream_cmd_in.num_iter  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\kdf_cmd_in.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\kdf_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\kdf_cmd_in.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\kdf_cmd_in.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\labels%s.guid_size  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\labels%s.label_size  1 5 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\labels%s.label  1 255 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\labels%s.delimiter_valid  1 0 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\labels%s.delimiter  1 7 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "labels (2,0) 1 271 0 7 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\kme_internal_out.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\kme_internal_out.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\kme_internal_out.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\kme_internal_out.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\kme_internal_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\debug_cmd.tlvp_corrupt  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\debug_cmd.cmd_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\debug_cmd.module_id  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\debug_cmd.cmd_type  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\debug_cmd.tlv_num  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\debug_cmd.byte_num  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\debug_cmd.byte_msk  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\int_tlv_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\int_tlv_word0.resv0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\int_tlv_word0.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\int_tlv_word0.keyless_algos  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\int_tlv_word0.needs_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\int_tlv_word0.needs_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\int_tlv_word0.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\int_tlv_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\int_tlv_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\int_tlv_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\int_tlv_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\int_tlv_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\int_tlv_word8.dek_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\int_tlv_word8.dek_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\int_tlv_word8.dek_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\int_tlv_word8.dek_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\int_tlv_word8.dek_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\int_tlv_word8.dek_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\int_tlv_word8.dek_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\int_tlv_word8.unused  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\int_tlv_word8.missing_iv  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\int_tlv_word8.missing_guid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\int_tlv_word8.validate_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\int_tlv_word8.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\int_tlv_word8.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\int_tlv_word8.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\int_tlv_word9.dak_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\int_tlv_word9.dak_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\int_tlv_word9.dak_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\int_tlv_word9.dak_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\int_tlv_word9.dak_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\int_tlv_word9.dak_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\int_tlv_word9.dak_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\int_tlv_word9.unused  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\int_tlv_word9.validate_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\int_tlv_word9.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\int_tlv_word9.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\int_tlv_word9.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\int_tlv_word42.corrupt_crc32  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\int_tlv_word42.unused  (1,0) 1 46 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\int_tlv_word42.error_code  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\key_header.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\key_header.dak_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\key_header.kdf_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\key_header.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m78 "\key_header.dek_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m79 "\stream_cmd_in.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m80 "\stream_cmd_in.skip  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m81 "\stream_cmd_in.guid  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m82 "\stream_cmd_in.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m83 "\stream_cmd_in.num_iter  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m84 "\stream_cmd_in_nxt.combo_mode  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m85 "\stream_cmd_in_nxt.skip  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m86 "\stream_cmd_in_nxt.guid  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m87 "\stream_cmd_in_nxt.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m88 "\stream_cmd_in_nxt.num_iter  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m89 "\gcm_dek_cmd_in.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m90 "\gcm_dek_cmd_in.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m91 "\gcm_dek_cmd_in.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m92 "\gcm_dek_cmd_in.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m93 "\gcm_dek_cmd_in_nxt.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m94 "\gcm_dek_cmd_in_nxt.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m95 "\gcm_dek_cmd_in_nxt.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m96 "\gcm_dek_cmd_in_nxt.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m97 "\gcm_dak_cmd_in.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m98 "\gcm_dak_cmd_in.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m99 "\gcm_dak_cmd_in.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m100 "\gcm_dak_cmd_in.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m101 "\gcm_dak_cmd_in_nxt.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m102 "\gcm_dak_cmd_in_nxt.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m103 "\gcm_dak_cmd_in_nxt.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m104 "\gcm_dak_cmd_in_nxt.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "104"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "gcm_cmd_in 4 \gcm_cmd_in.key0  \gcm_cmd_in.key1  \gcm_cmd_in.iv  \gcm_cmd_in.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "keyfilter_cmd_in 1 \keyfilter_cmd_in.combo_mode "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "kdfstream_cmd_in 5 \kdfstream_cmd_in.combo_mode  \kdfstream_cmd_in.skip  \kdfstream_cmd_in.guid  \kdfstream_cmd_in.label_index  \kdfstream_cmd_in.num_iter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "kdf_cmd_in 4 \kdf_cmd_in.kdf_dek_iter  \kdf_cmd_in.combo_mode  \kdf_cmd_in.dek_key_op  \kdf_cmd_in.dak_key_op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "labels%s 5 \labels%s.guid_size  \labels%s.label_size  \labels%s.label  \labels%s.delimiter_valid  \labels%s.delimiter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "kme_internal_out 5 \kme_internal_out.sot  \kme_internal_out.eoi  \kme_internal_out.eot  \kme_internal_out.id  \kme_internal_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "debug_cmd 7 \debug_cmd.tlvp_corrupt  \debug_cmd.cmd_mode  \debug_cmd.module_id  \debug_cmd.cmd_type  \debug_cmd.tlv_num  \debug_cmd.byte_num  \debug_cmd.byte_msk "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "int_tlv_word0 12 \int_tlv_word0.tlv_bip2  \int_tlv_word0.resv0  \int_tlv_word0.kdf_dek_iter  \int_tlv_word0.keyless_algos  \int_tlv_word0.needs_dek  \int_tlv_word0.needs_dak  \int_tlv_word0.key_type  \int_tlv_word0.tlv_frame_num  \int_tlv_word0.tlv_eng_id  \int_tlv_word0.tlv_seq_num  \int_tlv_word0.tlv_len  \int_tlv_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "int_tlv_word8 8 \int_tlv_word8.dek_kim_entry  { \int_tlv_word8.dek_kim_entry.valid  \int_tlv_word8.dek_kim_entry.label_index  \int_tlv_word8.dek_kim_entry.ckv_length  \int_tlv_word8.dek_kim_entry.ckv_pointer  \int_tlv_word8.dek_kim_entry.pf_num  \int_tlv_word8.dek_kim_entry.vf_num  \int_tlv_word8.dek_kim_entry.vf_valid  } \int_tlv_word8.unused  \int_tlv_word8.missing_iv  \int_tlv_word8.missing_guid  \int_tlv_word8.validate_dek  \int_tlv_word8.vf_valid  \int_tlv_word8.pf_num  \int_tlv_word8.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r10 "int_tlv_word9 6 \int_tlv_word9.dak_kim_entry  { \int_tlv_word9.dak_kim_entry.valid  \int_tlv_word9.dak_kim_entry.label_index  \int_tlv_word9.dak_kim_entry.ckv_length  \int_tlv_word9.dak_kim_entry.ckv_pointer  \int_tlv_word9.dak_kim_entry.pf_num  \int_tlv_word9.dak_kim_entry.vf_num  \int_tlv_word9.dak_kim_entry.vf_valid  } \int_tlv_word9.unused  \int_tlv_word9.validate_dak  \int_tlv_word9.vf_valid  \int_tlv_word9.pf_num  \int_tlv_word9.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r11 "int_tlv_word42 3 \int_tlv_word42.corrupt_crc32  \int_tlv_word42.unused  \int_tlv_word42.error_code "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r12 "key_header 5 \key_header.dak_key_op  \key_header.dak_key_ref  \key_header.kdf_mode  \key_header.dek_key_op  \key_header.dek_key_ref "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r13 "stream_cmd_in 5 \stream_cmd_in.combo_mode  \stream_cmd_in.skip  \stream_cmd_in.guid  \stream_cmd_in.label_index  \stream_cmd_in.num_iter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r14 "stream_cmd_in_nxt 5 \stream_cmd_in_nxt.combo_mode  \stream_cmd_in_nxt.skip  \stream_cmd_in_nxt.guid  \stream_cmd_in_nxt.label_index  \stream_cmd_in_nxt.num_iter "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r15 "gcm_dek_cmd_in 4 \gcm_dek_cmd_in.key0  \gcm_dek_cmd_in.key1  \gcm_dek_cmd_in.iv  \gcm_dek_cmd_in.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r16 "gcm_dek_cmd_in_nxt 4 \gcm_dek_cmd_in_nxt.key0  \gcm_dek_cmd_in_nxt.key1  \gcm_dek_cmd_in_nxt.iv  \gcm_dek_cmd_in_nxt.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r17 "gcm_dak_cmd_in 4 \gcm_dak_cmd_in.key0  \gcm_dak_cmd_in.key1  \gcm_dak_cmd_in.iv  \gcm_dak_cmd_in.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r18 "gcm_dak_cmd_in_nxt 4 \gcm_dak_cmd_in_nxt.key0  \gcm_dak_cmd_in_nxt.key1  \gcm_dak_cmd_in_nxt.iv  \gcm_dak_cmd_in_nxt.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "18"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_2 "1 delimiter 0 1 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 guid 0 1 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 op 0 7 "
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "guid[1].delimiter[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "guid[1].delimiter[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "guid[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "guid[0].delimiter[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "guid[0].delimiter[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "guid[0]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[7]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[6]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[5]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[4]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "op[0]"
endmodule
