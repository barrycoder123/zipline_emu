
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module IXC_SV_GFIFO_VXE_256 ( rdCnt);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input [63:0] rdCnt;
wire hasMultiLevelGFIFO;
wire fclk;
wire GFreq;
wire [19:0] GFcbid;
wire [11:0] GFlen;
wire [511:0] GFidata;
wire GFtsReq;
wire GFfull;
wire LBreq;
wire LBempty;
wire LBfull;
wire flushTbc;
wire [63:0] timeStampPkt;
wire flushTbc_x$tbc;
wire svGFbusy1;
wire svGFbusy2;
`_2_ wire GFtsAdd;
wire [3:0] LBrd;
wire [3:0] LBwr;
wire [3:0] LBwrI;
wire [3:0] LBfill;
`_2_ wire [11:0] argLen;
`_2_ wire [18:0] wLen;
`_2_ wire [17:0] rLen;
`_2_ wire wSync;
`_2_ wire rSync;
`_2_ wire [543:0] xdata;
`_2_ wire [63:0] wrtCnt;
`_2_ wire [63:0] wrtCntD;
wire [7:0] ackId;
wire [7:0] ackIdNew;
wire ackClk;
wire [17:0] ackLen;
`_2_ wire [14:0] ofifoAddr0;
`_2_ wire [14:0] ofifoAddr0N;
`_2_ wire [14:0] ofifoAddr1;
`_2_ wire [14:0] ofifoAddr1N;
`_2_ wire [14:0] ofifoAddr2;
`_2_ wire [14:0] ofifoAddr2N;
`_2_ wire [767:0] ofifoData;
`_2_ wire [767:0] ofifoDataN;
`_2_ wire [5:0] writeLen;
`_2_ wire reqD;
`_2_ wire GFfullD;
`_2_ wire [4:0] oFill;
`_2_ wire [4:0] oFillN;
`_2_ wire [14:0] ofifoWptr;
`_2_ wire [14:0] ofifoWptrN;
`_2_ wire [7:0] shiftCount;
`_2_ wire [767:0] shiftedXdata;
wire gfTsReqO;
wire [63:0] gfTsValO;
wire gfTsEn;
supply1 n1572;
supply0 n1584;
supply0 n1585;
supply0 n1611;
Q_BUF U0 ( .A(n1572), .Z(timeStampPkt[31]));
Q_BUF U1 ( .A(n1572), .Z(xc_top.hasGFIFO1));
Q_BUF U2 ( .A(n1611), .Z(shiftCount[0]));
Q_BUF U3 ( .A(n1611), .Z(shiftCount[1]));
Q_BUF U4 ( .A(n1611), .Z(shiftCount[2]));
Q_BUF U5 ( .A(n1611), .Z(shiftCount[3]));
Q_BUF U6 ( .A(n1611), .Z(shiftCount[4]));
Q_BUF U7 ( .A(gfTsValO[55]), .Z(timeStampPkt[63]));
Q_BUF U8 ( .A(gfTsValO[54]), .Z(timeStampPkt[62]));
Q_BUF U9 ( .A(gfTsValO[53]), .Z(timeStampPkt[61]));
Q_BUF U10 ( .A(gfTsValO[52]), .Z(timeStampPkt[60]));
Q_BUF U11 ( .A(gfTsValO[51]), .Z(timeStampPkt[59]));
Q_BUF U12 ( .A(gfTsValO[50]), .Z(timeStampPkt[58]));
Q_BUF U13 ( .A(gfTsValO[49]), .Z(timeStampPkt[57]));
Q_BUF U14 ( .A(gfTsValO[48]), .Z(timeStampPkt[56]));
Q_BUF U15 ( .A(gfTsValO[47]), .Z(timeStampPkt[55]));
Q_BUF U16 ( .A(gfTsValO[46]), .Z(timeStampPkt[54]));
Q_BUF U17 ( .A(gfTsValO[45]), .Z(timeStampPkt[53]));
Q_BUF U18 ( .A(gfTsValO[44]), .Z(timeStampPkt[52]));
Q_BUF U19 ( .A(gfTsValO[43]), .Z(timeStampPkt[51]));
Q_BUF U20 ( .A(gfTsValO[42]), .Z(timeStampPkt[50]));
Q_BUF U21 ( .A(gfTsValO[41]), .Z(timeStampPkt[49]));
Q_BUF U22 ( .A(gfTsValO[40]), .Z(timeStampPkt[48]));
Q_BUF U23 ( .A(gfTsValO[39]), .Z(timeStampPkt[47]));
Q_BUF U24 ( .A(gfTsValO[38]), .Z(timeStampPkt[46]));
Q_BUF U25 ( .A(gfTsValO[37]), .Z(timeStampPkt[45]));
Q_BUF U26 ( .A(gfTsValO[36]), .Z(timeStampPkt[44]));
Q_BUF U27 ( .A(gfTsValO[35]), .Z(timeStampPkt[43]));
Q_BUF U28 ( .A(gfTsValO[34]), .Z(timeStampPkt[42]));
Q_BUF U29 ( .A(gfTsValO[33]), .Z(timeStampPkt[41]));
Q_BUF U30 ( .A(gfTsValO[32]), .Z(timeStampPkt[40]));
Q_BUF U31 ( .A(gfTsValO[31]), .Z(timeStampPkt[39]));
Q_BUF U32 ( .A(gfTsValO[30]), .Z(timeStampPkt[38]));
Q_BUF U33 ( .A(gfTsValO[29]), .Z(timeStampPkt[37]));
Q_BUF U34 ( .A(gfTsValO[28]), .Z(timeStampPkt[36]));
Q_BUF U35 ( .A(gfTsValO[27]), .Z(timeStampPkt[35]));
Q_BUF U36 ( .A(gfTsValO[26]), .Z(timeStampPkt[34]));
Q_BUF U37 ( .A(gfTsValO[25]), .Z(timeStampPkt[33]));
Q_BUF U38 ( .A(gfTsValO[24]), .Z(timeStampPkt[32]));
Q_BUF U39 ( .A(gfTsValO[23]), .Z(timeStampPkt[23]));
Q_BUF U40 ( .A(gfTsValO[22]), .Z(timeStampPkt[22]));
Q_BUF U41 ( .A(gfTsValO[21]), .Z(timeStampPkt[21]));
Q_BUF U42 ( .A(gfTsValO[20]), .Z(timeStampPkt[20]));
Q_BUF U43 ( .A(gfTsValO[19]), .Z(timeStampPkt[19]));
Q_BUF U44 ( .A(gfTsValO[18]), .Z(timeStampPkt[18]));
Q_BUF U45 ( .A(gfTsValO[17]), .Z(timeStampPkt[17]));
Q_BUF U46 ( .A(gfTsValO[16]), .Z(timeStampPkt[16]));
Q_BUF U47 ( .A(gfTsValO[15]), .Z(timeStampPkt[15]));
Q_BUF U48 ( .A(gfTsValO[14]), .Z(timeStampPkt[14]));
Q_BUF U49 ( .A(gfTsValO[13]), .Z(timeStampPkt[13]));
Q_BUF U50 ( .A(gfTsValO[12]), .Z(timeStampPkt[12]));
Q_BUF U51 ( .A(gfTsValO[11]), .Z(timeStampPkt[11]));
Q_BUF U52 ( .A(gfTsValO[10]), .Z(timeStampPkt[10]));
Q_BUF U53 ( .A(gfTsValO[9]), .Z(timeStampPkt[9]));
Q_BUF U54 ( .A(gfTsValO[8]), .Z(timeStampPkt[8]));
Q_BUF U55 ( .A(gfTsValO[7]), .Z(timeStampPkt[7]));
Q_BUF U56 ( .A(gfTsValO[6]), .Z(timeStampPkt[6]));
Q_BUF U57 ( .A(gfTsValO[5]), .Z(timeStampPkt[5]));
Q_BUF U58 ( .A(gfTsValO[4]), .Z(timeStampPkt[4]));
Q_BUF U59 ( .A(gfTsValO[3]), .Z(timeStampPkt[3]));
Q_BUF U60 ( .A(gfTsValO[2]), .Z(timeStampPkt[2]));
Q_BUF U61 ( .A(gfTsValO[1]), .Z(timeStampPkt[1]));
Q_BUF U62 ( .A(gfTsValO[0]), .Z(timeStampPkt[0]));
Q_BUF U63 ( .A(oFill[0]), .Z(shiftCount[5]));
Q_BUF U64 ( .A(oFill[1]), .Z(shiftCount[6]));
Q_BUF U65 ( .A(oFill[2]), .Z(shiftCount[7]));
Q_BUF U66 ( .A(ofifoAddr2N[0]), .Z(ofifoAddr0N[0]));
Q_BUF U67 ( .A(ofifoWptr[0]), .Z(ofifoAddr2N[0]));
Q_BUF U68 ( .A(ofifoWptr[1]), .Z(ofifoAddr0N[1]));
Q_BUF U69 ( .A(ofifoWptr[2]), .Z(ofifoAddr0N[2]));
Q_BUF U70 ( .A(ofifoWptr[3]), .Z(ofifoAddr0N[3]));
Q_BUF U71 ( .A(ofifoWptr[4]), .Z(ofifoAddr0N[4]));
Q_BUF U72 ( .A(ofifoWptr[5]), .Z(ofifoAddr0N[5]));
Q_BUF U73 ( .A(ofifoWptr[6]), .Z(ofifoAddr0N[6]));
Q_BUF U74 ( .A(ofifoWptr[7]), .Z(ofifoAddr0N[7]));
Q_BUF U75 ( .A(ofifoWptr[8]), .Z(ofifoAddr0N[8]));
Q_BUF U76 ( .A(ofifoWptr[9]), .Z(ofifoAddr0N[9]));
Q_BUF U77 ( .A(ofifoWptr[10]), .Z(ofifoAddr0N[10]));
Q_BUF U78 ( .A(ofifoWptr[11]), .Z(ofifoAddr0N[11]));
Q_BUF U79 ( .A(ofifoWptr[12]), .Z(ofifoAddr0N[12]));
Q_BUF U80 ( .A(ofifoWptr[13]), .Z(ofifoAddr0N[13]));
Q_BUF U81 ( .A(ofifoWptr[14]), .Z(ofifoAddr0N[14]));
Q_AN02 U82 ( .A0(n6677), .A1(n6718), .Z(n6741));
Q_XOR2 U83 ( .A0(writeLen[4]), .A1(n1628), .Z(oFillN[4]));
Q_XOR2 U84 ( .A0(n3893), .A1(n3862), .Z(n3894));
Q_OR02 U85 ( .A0(n5814), .A1(GFlen[11]), .Z(n3926));
Q_XOR2 U86 ( .A0(n4416), .A1(n4423), .Z(n4417));
Q_MX08 U87 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][64] ), .A1(\TsBuf[1][64] ), .A2(\TsBuf[2][64] ), .A3(\TsBuf[3][64] ), .A4(\TsBuf[4][64] ), .A5(\TsBuf[5][64] ), .A6(\TsBuf[6][64] ), .A7(\TsBuf[7][64] ), .Z(gfTsReqO));
Q_MX08 U88 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][63] ), .A1(\TsBuf[1][63] ), .A2(\TsBuf[2][63] ), .A3(\TsBuf[3][63] ), .A4(\TsBuf[4][63] ), .A5(\TsBuf[5][63] ), .A6(\TsBuf[6][63] ), .A7(\TsBuf[7][63] ), .Z(gfTsValO[63]));
Q_MX08 U89 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][62] ), .A1(\TsBuf[1][62] ), .A2(\TsBuf[2][62] ), .A3(\TsBuf[3][62] ), .A4(\TsBuf[4][62] ), .A5(\TsBuf[5][62] ), .A6(\TsBuf[6][62] ), .A7(\TsBuf[7][62] ), .Z(gfTsValO[62]));
Q_MX08 U90 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][61] ), .A1(\TsBuf[1][61] ), .A2(\TsBuf[2][61] ), .A3(\TsBuf[3][61] ), .A4(\TsBuf[4][61] ), .A5(\TsBuf[5][61] ), .A6(\TsBuf[6][61] ), .A7(\TsBuf[7][61] ), .Z(gfTsValO[61]));
Q_MX08 U91 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][60] ), .A1(\TsBuf[1][60] ), .A2(\TsBuf[2][60] ), .A3(\TsBuf[3][60] ), .A4(\TsBuf[4][60] ), .A5(\TsBuf[5][60] ), .A6(\TsBuf[6][60] ), .A7(\TsBuf[7][60] ), .Z(gfTsValO[60]));
Q_MX08 U92 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][59] ), .A1(\TsBuf[1][59] ), .A2(\TsBuf[2][59] ), .A3(\TsBuf[3][59] ), .A4(\TsBuf[4][59] ), .A5(\TsBuf[5][59] ), .A6(\TsBuf[6][59] ), .A7(\TsBuf[7][59] ), .Z(gfTsValO[59]));
Q_MX08 U93 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][58] ), .A1(\TsBuf[1][58] ), .A2(\TsBuf[2][58] ), .A3(\TsBuf[3][58] ), .A4(\TsBuf[4][58] ), .A5(\TsBuf[5][58] ), .A6(\TsBuf[6][58] ), .A7(\TsBuf[7][58] ), .Z(gfTsValO[58]));
Q_MX08 U94 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][57] ), .A1(\TsBuf[1][57] ), .A2(\TsBuf[2][57] ), .A3(\TsBuf[3][57] ), .A4(\TsBuf[4][57] ), .A5(\TsBuf[5][57] ), .A6(\TsBuf[6][57] ), .A7(\TsBuf[7][57] ), .Z(gfTsValO[57]));
Q_MX08 U95 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][56] ), .A1(\TsBuf[1][56] ), .A2(\TsBuf[2][56] ), .A3(\TsBuf[3][56] ), .A4(\TsBuf[4][56] ), .A5(\TsBuf[5][56] ), .A6(\TsBuf[6][56] ), .A7(\TsBuf[7][56] ), .Z(gfTsValO[56]));
Q_MX08 U96 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][55] ), .A1(\TsBuf[1][55] ), .A2(\TsBuf[2][55] ), .A3(\TsBuf[3][55] ), .A4(\TsBuf[4][55] ), .A5(\TsBuf[5][55] ), .A6(\TsBuf[6][55] ), .A7(\TsBuf[7][55] ), .Z(gfTsValO[55]));
Q_MX08 U97 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][54] ), .A1(\TsBuf[1][54] ), .A2(\TsBuf[2][54] ), .A3(\TsBuf[3][54] ), .A4(\TsBuf[4][54] ), .A5(\TsBuf[5][54] ), .A6(\TsBuf[6][54] ), .A7(\TsBuf[7][54] ), .Z(gfTsValO[54]));
Q_MX08 U98 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][53] ), .A1(\TsBuf[1][53] ), .A2(\TsBuf[2][53] ), .A3(\TsBuf[3][53] ), .A4(\TsBuf[4][53] ), .A5(\TsBuf[5][53] ), .A6(\TsBuf[6][53] ), .A7(\TsBuf[7][53] ), .Z(gfTsValO[53]));
Q_MX08 U99 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][52] ), .A1(\TsBuf[1][52] ), .A2(\TsBuf[2][52] ), .A3(\TsBuf[3][52] ), .A4(\TsBuf[4][52] ), .A5(\TsBuf[5][52] ), .A6(\TsBuf[6][52] ), .A7(\TsBuf[7][52] ), .Z(gfTsValO[52]));
Q_MX08 U100 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][51] ), .A1(\TsBuf[1][51] ), .A2(\TsBuf[2][51] ), .A3(\TsBuf[3][51] ), .A4(\TsBuf[4][51] ), .A5(\TsBuf[5][51] ), .A6(\TsBuf[6][51] ), .A7(\TsBuf[7][51] ), .Z(gfTsValO[51]));
Q_MX08 U101 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][50] ), .A1(\TsBuf[1][50] ), .A2(\TsBuf[2][50] ), .A3(\TsBuf[3][50] ), .A4(\TsBuf[4][50] ), .A5(\TsBuf[5][50] ), .A6(\TsBuf[6][50] ), .A7(\TsBuf[7][50] ), .Z(gfTsValO[50]));
Q_MX08 U102 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][49] ), .A1(\TsBuf[1][49] ), .A2(\TsBuf[2][49] ), .A3(\TsBuf[3][49] ), .A4(\TsBuf[4][49] ), .A5(\TsBuf[5][49] ), .A6(\TsBuf[6][49] ), .A7(\TsBuf[7][49] ), .Z(gfTsValO[49]));
Q_MX08 U103 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][48] ), .A1(\TsBuf[1][48] ), .A2(\TsBuf[2][48] ), .A3(\TsBuf[3][48] ), .A4(\TsBuf[4][48] ), .A5(\TsBuf[5][48] ), .A6(\TsBuf[6][48] ), .A7(\TsBuf[7][48] ), .Z(gfTsValO[48]));
Q_MX08 U104 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][47] ), .A1(\TsBuf[1][47] ), .A2(\TsBuf[2][47] ), .A3(\TsBuf[3][47] ), .A4(\TsBuf[4][47] ), .A5(\TsBuf[5][47] ), .A6(\TsBuf[6][47] ), .A7(\TsBuf[7][47] ), .Z(gfTsValO[47]));
Q_MX08 U105 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][46] ), .A1(\TsBuf[1][46] ), .A2(\TsBuf[2][46] ), .A3(\TsBuf[3][46] ), .A4(\TsBuf[4][46] ), .A5(\TsBuf[5][46] ), .A6(\TsBuf[6][46] ), .A7(\TsBuf[7][46] ), .Z(gfTsValO[46]));
Q_MX08 U106 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][45] ), .A1(\TsBuf[1][45] ), .A2(\TsBuf[2][45] ), .A3(\TsBuf[3][45] ), .A4(\TsBuf[4][45] ), .A5(\TsBuf[5][45] ), .A6(\TsBuf[6][45] ), .A7(\TsBuf[7][45] ), .Z(gfTsValO[45]));
Q_MX08 U107 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][44] ), .A1(\TsBuf[1][44] ), .A2(\TsBuf[2][44] ), .A3(\TsBuf[3][44] ), .A4(\TsBuf[4][44] ), .A5(\TsBuf[5][44] ), .A6(\TsBuf[6][44] ), .A7(\TsBuf[7][44] ), .Z(gfTsValO[44]));
Q_MX08 U108 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][43] ), .A1(\TsBuf[1][43] ), .A2(\TsBuf[2][43] ), .A3(\TsBuf[3][43] ), .A4(\TsBuf[4][43] ), .A5(\TsBuf[5][43] ), .A6(\TsBuf[6][43] ), .A7(\TsBuf[7][43] ), .Z(gfTsValO[43]));
Q_MX08 U109 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][42] ), .A1(\TsBuf[1][42] ), .A2(\TsBuf[2][42] ), .A3(\TsBuf[3][42] ), .A4(\TsBuf[4][42] ), .A5(\TsBuf[5][42] ), .A6(\TsBuf[6][42] ), .A7(\TsBuf[7][42] ), .Z(gfTsValO[42]));
Q_MX08 U110 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][41] ), .A1(\TsBuf[1][41] ), .A2(\TsBuf[2][41] ), .A3(\TsBuf[3][41] ), .A4(\TsBuf[4][41] ), .A5(\TsBuf[5][41] ), .A6(\TsBuf[6][41] ), .A7(\TsBuf[7][41] ), .Z(gfTsValO[41]));
Q_MX08 U111 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][40] ), .A1(\TsBuf[1][40] ), .A2(\TsBuf[2][40] ), .A3(\TsBuf[3][40] ), .A4(\TsBuf[4][40] ), .A5(\TsBuf[5][40] ), .A6(\TsBuf[6][40] ), .A7(\TsBuf[7][40] ), .Z(gfTsValO[40]));
Q_MX08 U112 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][39] ), .A1(\TsBuf[1][39] ), .A2(\TsBuf[2][39] ), .A3(\TsBuf[3][39] ), .A4(\TsBuf[4][39] ), .A5(\TsBuf[5][39] ), .A6(\TsBuf[6][39] ), .A7(\TsBuf[7][39] ), .Z(gfTsValO[39]));
Q_MX08 U113 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][38] ), .A1(\TsBuf[1][38] ), .A2(\TsBuf[2][38] ), .A3(\TsBuf[3][38] ), .A4(\TsBuf[4][38] ), .A5(\TsBuf[5][38] ), .A6(\TsBuf[6][38] ), .A7(\TsBuf[7][38] ), .Z(gfTsValO[38]));
Q_MX08 U114 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][37] ), .A1(\TsBuf[1][37] ), .A2(\TsBuf[2][37] ), .A3(\TsBuf[3][37] ), .A4(\TsBuf[4][37] ), .A5(\TsBuf[5][37] ), .A6(\TsBuf[6][37] ), .A7(\TsBuf[7][37] ), .Z(gfTsValO[37]));
Q_MX08 U115 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][36] ), .A1(\TsBuf[1][36] ), .A2(\TsBuf[2][36] ), .A3(\TsBuf[3][36] ), .A4(\TsBuf[4][36] ), .A5(\TsBuf[5][36] ), .A6(\TsBuf[6][36] ), .A7(\TsBuf[7][36] ), .Z(gfTsValO[36]));
Q_MX08 U116 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][35] ), .A1(\TsBuf[1][35] ), .A2(\TsBuf[2][35] ), .A3(\TsBuf[3][35] ), .A4(\TsBuf[4][35] ), .A5(\TsBuf[5][35] ), .A6(\TsBuf[6][35] ), .A7(\TsBuf[7][35] ), .Z(gfTsValO[35]));
Q_MX08 U117 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][34] ), .A1(\TsBuf[1][34] ), .A2(\TsBuf[2][34] ), .A3(\TsBuf[3][34] ), .A4(\TsBuf[4][34] ), .A5(\TsBuf[5][34] ), .A6(\TsBuf[6][34] ), .A7(\TsBuf[7][34] ), .Z(gfTsValO[34]));
Q_MX08 U118 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][33] ), .A1(\TsBuf[1][33] ), .A2(\TsBuf[2][33] ), .A3(\TsBuf[3][33] ), .A4(\TsBuf[4][33] ), .A5(\TsBuf[5][33] ), .A6(\TsBuf[6][33] ), .A7(\TsBuf[7][33] ), .Z(gfTsValO[33]));
Q_MX08 U119 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][32] ), .A1(\TsBuf[1][32] ), .A2(\TsBuf[2][32] ), .A3(\TsBuf[3][32] ), .A4(\TsBuf[4][32] ), .A5(\TsBuf[5][32] ), .A6(\TsBuf[6][32] ), .A7(\TsBuf[7][32] ), .Z(gfTsValO[32]));
Q_MX08 U120 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][31] ), .A1(\TsBuf[1][31] ), .A2(\TsBuf[2][31] ), .A3(\TsBuf[3][31] ), .A4(\TsBuf[4][31] ), .A5(\TsBuf[5][31] ), .A6(\TsBuf[6][31] ), .A7(\TsBuf[7][31] ), .Z(gfTsValO[31]));
Q_MX08 U121 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][30] ), .A1(\TsBuf[1][30] ), .A2(\TsBuf[2][30] ), .A3(\TsBuf[3][30] ), .A4(\TsBuf[4][30] ), .A5(\TsBuf[5][30] ), .A6(\TsBuf[6][30] ), .A7(\TsBuf[7][30] ), .Z(gfTsValO[30]));
Q_MX08 U122 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][29] ), .A1(\TsBuf[1][29] ), .A2(\TsBuf[2][29] ), .A3(\TsBuf[3][29] ), .A4(\TsBuf[4][29] ), .A5(\TsBuf[5][29] ), .A6(\TsBuf[6][29] ), .A7(\TsBuf[7][29] ), .Z(gfTsValO[29]));
Q_MX08 U123 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][28] ), .A1(\TsBuf[1][28] ), .A2(\TsBuf[2][28] ), .A3(\TsBuf[3][28] ), .A4(\TsBuf[4][28] ), .A5(\TsBuf[5][28] ), .A6(\TsBuf[6][28] ), .A7(\TsBuf[7][28] ), .Z(gfTsValO[28]));
Q_MX08 U124 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][27] ), .A1(\TsBuf[1][27] ), .A2(\TsBuf[2][27] ), .A3(\TsBuf[3][27] ), .A4(\TsBuf[4][27] ), .A5(\TsBuf[5][27] ), .A6(\TsBuf[6][27] ), .A7(\TsBuf[7][27] ), .Z(gfTsValO[27]));
Q_MX08 U125 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][26] ), .A1(\TsBuf[1][26] ), .A2(\TsBuf[2][26] ), .A3(\TsBuf[3][26] ), .A4(\TsBuf[4][26] ), .A5(\TsBuf[5][26] ), .A6(\TsBuf[6][26] ), .A7(\TsBuf[7][26] ), .Z(gfTsValO[26]));
Q_MX08 U126 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][25] ), .A1(\TsBuf[1][25] ), .A2(\TsBuf[2][25] ), .A3(\TsBuf[3][25] ), .A4(\TsBuf[4][25] ), .A5(\TsBuf[5][25] ), .A6(\TsBuf[6][25] ), .A7(\TsBuf[7][25] ), .Z(gfTsValO[25]));
Q_MX08 U127 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][24] ), .A1(\TsBuf[1][24] ), .A2(\TsBuf[2][24] ), .A3(\TsBuf[3][24] ), .A4(\TsBuf[4][24] ), .A5(\TsBuf[5][24] ), .A6(\TsBuf[6][24] ), .A7(\TsBuf[7][24] ), .Z(gfTsValO[24]));
Q_MX08 U128 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][23] ), .A1(\TsBuf[1][23] ), .A2(\TsBuf[2][23] ), .A3(\TsBuf[3][23] ), .A4(\TsBuf[4][23] ), .A5(\TsBuf[5][23] ), .A6(\TsBuf[6][23] ), .A7(\TsBuf[7][23] ), .Z(gfTsValO[23]));
Q_MX08 U129 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][22] ), .A1(\TsBuf[1][22] ), .A2(\TsBuf[2][22] ), .A3(\TsBuf[3][22] ), .A4(\TsBuf[4][22] ), .A5(\TsBuf[5][22] ), .A6(\TsBuf[6][22] ), .A7(\TsBuf[7][22] ), .Z(gfTsValO[22]));
Q_MX08 U130 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][21] ), .A1(\TsBuf[1][21] ), .A2(\TsBuf[2][21] ), .A3(\TsBuf[3][21] ), .A4(\TsBuf[4][21] ), .A5(\TsBuf[5][21] ), .A6(\TsBuf[6][21] ), .A7(\TsBuf[7][21] ), .Z(gfTsValO[21]));
Q_MX08 U131 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][20] ), .A1(\TsBuf[1][20] ), .A2(\TsBuf[2][20] ), .A3(\TsBuf[3][20] ), .A4(\TsBuf[4][20] ), .A5(\TsBuf[5][20] ), .A6(\TsBuf[6][20] ), .A7(\TsBuf[7][20] ), .Z(gfTsValO[20]));
Q_MX08 U132 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][19] ), .A1(\TsBuf[1][19] ), .A2(\TsBuf[2][19] ), .A3(\TsBuf[3][19] ), .A4(\TsBuf[4][19] ), .A5(\TsBuf[5][19] ), .A6(\TsBuf[6][19] ), .A7(\TsBuf[7][19] ), .Z(gfTsValO[19]));
Q_MX08 U133 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][18] ), .A1(\TsBuf[1][18] ), .A2(\TsBuf[2][18] ), .A3(\TsBuf[3][18] ), .A4(\TsBuf[4][18] ), .A5(\TsBuf[5][18] ), .A6(\TsBuf[6][18] ), .A7(\TsBuf[7][18] ), .Z(gfTsValO[18]));
Q_MX08 U134 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][17] ), .A1(\TsBuf[1][17] ), .A2(\TsBuf[2][17] ), .A3(\TsBuf[3][17] ), .A4(\TsBuf[4][17] ), .A5(\TsBuf[5][17] ), .A6(\TsBuf[6][17] ), .A7(\TsBuf[7][17] ), .Z(gfTsValO[17]));
Q_MX08 U135 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][16] ), .A1(\TsBuf[1][16] ), .A2(\TsBuf[2][16] ), .A3(\TsBuf[3][16] ), .A4(\TsBuf[4][16] ), .A5(\TsBuf[5][16] ), .A6(\TsBuf[6][16] ), .A7(\TsBuf[7][16] ), .Z(gfTsValO[16]));
Q_MX08 U136 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][15] ), .A1(\TsBuf[1][15] ), .A2(\TsBuf[2][15] ), .A3(\TsBuf[3][15] ), .A4(\TsBuf[4][15] ), .A5(\TsBuf[5][15] ), .A6(\TsBuf[6][15] ), .A7(\TsBuf[7][15] ), .Z(gfTsValO[15]));
Q_MX08 U137 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][14] ), .A1(\TsBuf[1][14] ), .A2(\TsBuf[2][14] ), .A3(\TsBuf[3][14] ), .A4(\TsBuf[4][14] ), .A5(\TsBuf[5][14] ), .A6(\TsBuf[6][14] ), .A7(\TsBuf[7][14] ), .Z(gfTsValO[14]));
Q_MX08 U138 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][13] ), .A1(\TsBuf[1][13] ), .A2(\TsBuf[2][13] ), .A3(\TsBuf[3][13] ), .A4(\TsBuf[4][13] ), .A5(\TsBuf[5][13] ), .A6(\TsBuf[6][13] ), .A7(\TsBuf[7][13] ), .Z(gfTsValO[13]));
Q_MX08 U139 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][12] ), .A1(\TsBuf[1][12] ), .A2(\TsBuf[2][12] ), .A3(\TsBuf[3][12] ), .A4(\TsBuf[4][12] ), .A5(\TsBuf[5][12] ), .A6(\TsBuf[6][12] ), .A7(\TsBuf[7][12] ), .Z(gfTsValO[12]));
Q_MX08 U140 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][11] ), .A1(\TsBuf[1][11] ), .A2(\TsBuf[2][11] ), .A3(\TsBuf[3][11] ), .A4(\TsBuf[4][11] ), .A5(\TsBuf[5][11] ), .A6(\TsBuf[6][11] ), .A7(\TsBuf[7][11] ), .Z(gfTsValO[11]));
Q_MX08 U141 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][10] ), .A1(\TsBuf[1][10] ), .A2(\TsBuf[2][10] ), .A3(\TsBuf[3][10] ), .A4(\TsBuf[4][10] ), .A5(\TsBuf[5][10] ), .A6(\TsBuf[6][10] ), .A7(\TsBuf[7][10] ), .Z(gfTsValO[10]));
Q_MX08 U142 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][9] ), .A1(\TsBuf[1][9] ), .A2(\TsBuf[2][9] ), .A3(\TsBuf[3][9] ), .A4(\TsBuf[4][9] ), .A5(\TsBuf[5][9] ), .A6(\TsBuf[6][9] ), .A7(\TsBuf[7][9] ), .Z(gfTsValO[9]));
Q_MX08 U143 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][8] ), .A1(\TsBuf[1][8] ), .A2(\TsBuf[2][8] ), .A3(\TsBuf[3][8] ), .A4(\TsBuf[4][8] ), .A5(\TsBuf[5][8] ), .A6(\TsBuf[6][8] ), .A7(\TsBuf[7][8] ), .Z(gfTsValO[8]));
Q_MX08 U144 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][7] ), .A1(\TsBuf[1][7] ), .A2(\TsBuf[2][7] ), .A3(\TsBuf[3][7] ), .A4(\TsBuf[4][7] ), .A5(\TsBuf[5][7] ), .A6(\TsBuf[6][7] ), .A7(\TsBuf[7][7] ), .Z(gfTsValO[7]));
Q_MX08 U145 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][6] ), .A1(\TsBuf[1][6] ), .A2(\TsBuf[2][6] ), .A3(\TsBuf[3][6] ), .A4(\TsBuf[4][6] ), .A5(\TsBuf[5][6] ), .A6(\TsBuf[6][6] ), .A7(\TsBuf[7][6] ), .Z(gfTsValO[6]));
Q_MX08 U146 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][5] ), .A1(\TsBuf[1][5] ), .A2(\TsBuf[2][5] ), .A3(\TsBuf[3][5] ), .A4(\TsBuf[4][5] ), .A5(\TsBuf[5][5] ), .A6(\TsBuf[6][5] ), .A7(\TsBuf[7][5] ), .Z(gfTsValO[5]));
Q_MX08 U147 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][4] ), .A1(\TsBuf[1][4] ), .A2(\TsBuf[2][4] ), .A3(\TsBuf[3][4] ), .A4(\TsBuf[4][4] ), .A5(\TsBuf[5][4] ), .A6(\TsBuf[6][4] ), .A7(\TsBuf[7][4] ), .Z(gfTsValO[4]));
Q_MX08 U148 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][3] ), .A1(\TsBuf[1][3] ), .A2(\TsBuf[2][3] ), .A3(\TsBuf[3][3] ), .A4(\TsBuf[4][3] ), .A5(\TsBuf[5][3] ), .A6(\TsBuf[6][3] ), .A7(\TsBuf[7][3] ), .Z(gfTsValO[3]));
Q_MX08 U149 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][2] ), .A1(\TsBuf[1][2] ), .A2(\TsBuf[2][2] ), .A3(\TsBuf[3][2] ), .A4(\TsBuf[4][2] ), .A5(\TsBuf[5][2] ), .A6(\TsBuf[6][2] ), .A7(\TsBuf[7][2] ), .Z(gfTsValO[2]));
Q_MX08 U150 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][1] ), .A1(\TsBuf[1][1] ), .A2(\TsBuf[2][1] ), .A3(\TsBuf[3][1] ), .A4(\TsBuf[4][1] ), .A5(\TsBuf[5][1] ), .A6(\TsBuf[6][1] ), .A7(\TsBuf[7][1] ), .Z(gfTsValO[1]));
Q_MX08 U151 ( .S0(LBrd[0]), .S1(LBrd[1]), .S2(LBrd[2]), .A0(\TsBuf[0][0] ), .A1(\TsBuf[1][0] ), .A2(\TsBuf[2][0] ), .A3(\TsBuf[3][0] ), .A4(\TsBuf[4][0] ), .A5(\TsBuf[5][0] ), .A6(\TsBuf[6][0] ), .A7(\TsBuf[7][0] ), .Z(gfTsValO[0]));
Q_LDP0 \TsBuf_REG[7][64] ( .G(n6739), .D(GFtsReq), .Q(\TsBuf[7][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][63] ( .G(n6739), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[7][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][62] ( .G(n6739), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[7][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][61] ( .G(n6739), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[7][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][60] ( .G(n6739), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[7][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][59] ( .G(n6739), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[7][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][58] ( .G(n6739), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[7][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][57] ( .G(n6739), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[7][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][56] ( .G(n6739), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[7][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][55] ( .G(n6739), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[7][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][54] ( .G(n6739), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[7][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][53] ( .G(n6739), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[7][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][52] ( .G(n6739), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[7][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][51] ( .G(n6739), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[7][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][50] ( .G(n6739), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[7][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][49] ( .G(n6739), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[7][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][48] ( .G(n6739), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[7][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][47] ( .G(n6739), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[7][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][46] ( .G(n6739), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[7][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][45] ( .G(n6739), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[7][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][44] ( .G(n6739), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[7][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][43] ( .G(n6739), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[7][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][42] ( .G(n6739), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[7][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][41] ( .G(n6739), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[7][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][40] ( .G(n6739), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[7][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][39] ( .G(n6739), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[7][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][38] ( .G(n6739), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[7][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][37] ( .G(n6739), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[7][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][36] ( .G(n6739), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[7][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][35] ( .G(n6739), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[7][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][34] ( .G(n6739), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[7][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][33] ( .G(n6739), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[7][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][32] ( .G(n6739), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[7][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][31] ( .G(n6739), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[7][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][30] ( .G(n6739), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[7][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][29] ( .G(n6739), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[7][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][28] ( .G(n6739), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[7][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][27] ( .G(n6739), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[7][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][26] ( .G(n6739), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[7][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][25] ( .G(n6739), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[7][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][24] ( .G(n6739), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[7][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][23] ( .G(n6739), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[7][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][22] ( .G(n6739), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[7][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][21] ( .G(n6739), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[7][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][20] ( .G(n6739), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[7][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][19] ( .G(n6739), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[7][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][18] ( .G(n6739), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[7][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][17] ( .G(n6739), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[7][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][16] ( .G(n6739), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[7][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][15] ( .G(n6739), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[7][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][14] ( .G(n6739), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[7][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][13] ( .G(n6739), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[7][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][12] ( .G(n6739), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[7][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][11] ( .G(n6739), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[7][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][10] ( .G(n6739), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[7][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][9] ( .G(n6739), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[7][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][8] ( .G(n6739), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[7][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][7] ( .G(n6739), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[7][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][6] ( .G(n6739), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[7][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][5] ( .G(n6739), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[7][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][4] ( .G(n6739), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[7][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][3] ( .G(n6739), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[7][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][2] ( .G(n6739), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[7][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][1] ( .G(n6739), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[7][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[7][0] ( .G(n6739), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[7][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][64] ( .G(n6738), .D(GFtsReq), .Q(\TsBuf[6][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][63] ( .G(n6738), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[6][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][62] ( .G(n6738), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[6][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][61] ( .G(n6738), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[6][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][60] ( .G(n6738), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[6][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][59] ( .G(n6738), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[6][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][58] ( .G(n6738), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[6][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][57] ( .G(n6738), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[6][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][56] ( .G(n6738), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[6][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][55] ( .G(n6738), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[6][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][54] ( .G(n6738), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[6][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][53] ( .G(n6738), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[6][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][52] ( .G(n6738), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[6][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][51] ( .G(n6738), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[6][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][50] ( .G(n6738), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[6][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][49] ( .G(n6738), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[6][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][48] ( .G(n6738), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[6][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][47] ( .G(n6738), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[6][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][46] ( .G(n6738), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[6][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][45] ( .G(n6738), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[6][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][44] ( .G(n6738), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[6][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][43] ( .G(n6738), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[6][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][42] ( .G(n6738), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[6][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][41] ( .G(n6738), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[6][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][40] ( .G(n6738), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[6][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][39] ( .G(n6738), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[6][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][38] ( .G(n6738), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[6][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][37] ( .G(n6738), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[6][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][36] ( .G(n6738), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[6][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][35] ( .G(n6738), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[6][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][34] ( .G(n6738), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[6][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][33] ( .G(n6738), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[6][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][32] ( .G(n6738), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[6][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][31] ( .G(n6738), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[6][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][30] ( .G(n6738), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[6][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][29] ( .G(n6738), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[6][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][28] ( .G(n6738), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[6][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][27] ( .G(n6738), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[6][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][26] ( .G(n6738), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[6][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][25] ( .G(n6738), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[6][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][24] ( .G(n6738), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[6][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][23] ( .G(n6738), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[6][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][22] ( .G(n6738), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[6][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][21] ( .G(n6738), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[6][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][20] ( .G(n6738), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[6][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][19] ( .G(n6738), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[6][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][18] ( .G(n6738), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[6][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][17] ( .G(n6738), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[6][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][16] ( .G(n6738), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[6][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][15] ( .G(n6738), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[6][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][14] ( .G(n6738), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[6][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][13] ( .G(n6738), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[6][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][12] ( .G(n6738), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[6][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][11] ( .G(n6738), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[6][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][10] ( .G(n6738), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[6][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][9] ( .G(n6738), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[6][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][8] ( .G(n6738), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[6][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][7] ( .G(n6738), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[6][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][6] ( .G(n6738), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[6][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][5] ( .G(n6738), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[6][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][4] ( .G(n6738), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[6][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][3] ( .G(n6738), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[6][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][2] ( .G(n6738), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[6][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][1] ( .G(n6738), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[6][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[6][0] ( .G(n6738), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[6][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][64] ( .G(n6737), .D(GFtsReq), .Q(\TsBuf[5][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][63] ( .G(n6737), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[5][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][62] ( .G(n6737), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[5][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][61] ( .G(n6737), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[5][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][60] ( .G(n6737), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[5][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][59] ( .G(n6737), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[5][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][58] ( .G(n6737), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[5][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][57] ( .G(n6737), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[5][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][56] ( .G(n6737), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[5][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][55] ( .G(n6737), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[5][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][54] ( .G(n6737), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[5][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][53] ( .G(n6737), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[5][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][52] ( .G(n6737), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[5][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][51] ( .G(n6737), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[5][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][50] ( .G(n6737), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[5][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][49] ( .G(n6737), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[5][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][48] ( .G(n6737), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[5][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][47] ( .G(n6737), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[5][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][46] ( .G(n6737), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[5][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][45] ( .G(n6737), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[5][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][44] ( .G(n6737), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[5][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][43] ( .G(n6737), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[5][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][42] ( .G(n6737), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[5][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][41] ( .G(n6737), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[5][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][40] ( .G(n6737), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[5][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][39] ( .G(n6737), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[5][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][38] ( .G(n6737), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[5][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][37] ( .G(n6737), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[5][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][36] ( .G(n6737), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[5][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][35] ( .G(n6737), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[5][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][34] ( .G(n6737), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[5][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][33] ( .G(n6737), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[5][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][32] ( .G(n6737), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[5][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][31] ( .G(n6737), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[5][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][30] ( .G(n6737), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[5][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][29] ( .G(n6737), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[5][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][28] ( .G(n6737), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[5][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][27] ( .G(n6737), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[5][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][26] ( .G(n6737), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[5][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][25] ( .G(n6737), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[5][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][24] ( .G(n6737), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[5][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][23] ( .G(n6737), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[5][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][22] ( .G(n6737), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[5][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][21] ( .G(n6737), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[5][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][20] ( .G(n6737), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[5][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][19] ( .G(n6737), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[5][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][18] ( .G(n6737), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[5][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][17] ( .G(n6737), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[5][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][16] ( .G(n6737), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[5][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][15] ( .G(n6737), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[5][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][14] ( .G(n6737), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[5][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][13] ( .G(n6737), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[5][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][12] ( .G(n6737), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[5][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][11] ( .G(n6737), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[5][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][10] ( .G(n6737), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[5][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][9] ( .G(n6737), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[5][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][8] ( .G(n6737), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[5][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][7] ( .G(n6737), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[5][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][6] ( .G(n6737), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[5][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][5] ( .G(n6737), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[5][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][4] ( .G(n6737), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[5][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][3] ( .G(n6737), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[5][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][2] ( .G(n6737), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[5][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][1] ( .G(n6737), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[5][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[5][0] ( .G(n6737), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[5][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][64] ( .G(n6736), .D(GFtsReq), .Q(\TsBuf[4][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][63] ( .G(n6736), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[4][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][62] ( .G(n6736), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[4][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][61] ( .G(n6736), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[4][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][60] ( .G(n6736), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[4][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][59] ( .G(n6736), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[4][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][58] ( .G(n6736), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[4][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][57] ( .G(n6736), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[4][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][56] ( .G(n6736), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[4][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][55] ( .G(n6736), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[4][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][54] ( .G(n6736), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[4][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][53] ( .G(n6736), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[4][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][52] ( .G(n6736), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[4][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][51] ( .G(n6736), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[4][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][50] ( .G(n6736), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[4][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][49] ( .G(n6736), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[4][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][48] ( .G(n6736), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[4][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][47] ( .G(n6736), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[4][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][46] ( .G(n6736), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[4][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][45] ( .G(n6736), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[4][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][44] ( .G(n6736), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[4][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][43] ( .G(n6736), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[4][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][42] ( .G(n6736), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[4][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][41] ( .G(n6736), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[4][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][40] ( .G(n6736), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[4][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][39] ( .G(n6736), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[4][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][38] ( .G(n6736), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[4][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][37] ( .G(n6736), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[4][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][36] ( .G(n6736), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[4][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][35] ( .G(n6736), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[4][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][34] ( .G(n6736), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[4][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][33] ( .G(n6736), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[4][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][32] ( .G(n6736), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[4][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][31] ( .G(n6736), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[4][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][30] ( .G(n6736), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[4][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][29] ( .G(n6736), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[4][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][28] ( .G(n6736), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[4][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][27] ( .G(n6736), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[4][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][26] ( .G(n6736), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[4][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][25] ( .G(n6736), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[4][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][24] ( .G(n6736), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[4][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][23] ( .G(n6736), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[4][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][22] ( .G(n6736), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[4][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][21] ( .G(n6736), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[4][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][20] ( .G(n6736), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[4][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][19] ( .G(n6736), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[4][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][18] ( .G(n6736), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[4][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][17] ( .G(n6736), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[4][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][16] ( .G(n6736), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[4][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][15] ( .G(n6736), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[4][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][14] ( .G(n6736), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[4][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][13] ( .G(n6736), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[4][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][12] ( .G(n6736), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[4][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][11] ( .G(n6736), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[4][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][10] ( .G(n6736), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[4][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][9] ( .G(n6736), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[4][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][8] ( .G(n6736), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[4][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][7] ( .G(n6736), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[4][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][6] ( .G(n6736), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[4][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][5] ( .G(n6736), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[4][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][4] ( .G(n6736), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[4][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][3] ( .G(n6736), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[4][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][2] ( .G(n6736), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[4][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][1] ( .G(n6736), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[4][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[4][0] ( .G(n6736), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[4][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][64] ( .G(n6735), .D(GFtsReq), .Q(\TsBuf[3][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][63] ( .G(n6735), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[3][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][62] ( .G(n6735), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[3][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][61] ( .G(n6735), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[3][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][60] ( .G(n6735), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[3][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][59] ( .G(n6735), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[3][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][58] ( .G(n6735), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[3][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][57] ( .G(n6735), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[3][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][56] ( .G(n6735), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[3][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][55] ( .G(n6735), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[3][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][54] ( .G(n6735), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[3][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][53] ( .G(n6735), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[3][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][52] ( .G(n6735), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[3][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][51] ( .G(n6735), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[3][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][50] ( .G(n6735), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[3][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][49] ( .G(n6735), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[3][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][48] ( .G(n6735), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[3][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][47] ( .G(n6735), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[3][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][46] ( .G(n6735), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[3][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][45] ( .G(n6735), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[3][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][44] ( .G(n6735), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[3][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][43] ( .G(n6735), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[3][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][42] ( .G(n6735), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[3][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][41] ( .G(n6735), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[3][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][40] ( .G(n6735), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[3][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][39] ( .G(n6735), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[3][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][38] ( .G(n6735), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[3][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][37] ( .G(n6735), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[3][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][36] ( .G(n6735), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[3][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][35] ( .G(n6735), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[3][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][34] ( .G(n6735), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[3][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][33] ( .G(n6735), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[3][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][32] ( .G(n6735), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[3][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][31] ( .G(n6735), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[3][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][30] ( .G(n6735), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[3][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][29] ( .G(n6735), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[3][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][28] ( .G(n6735), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[3][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][27] ( .G(n6735), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[3][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][26] ( .G(n6735), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[3][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][25] ( .G(n6735), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[3][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][24] ( .G(n6735), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[3][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][23] ( .G(n6735), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[3][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][22] ( .G(n6735), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[3][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][21] ( .G(n6735), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[3][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][20] ( .G(n6735), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[3][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][19] ( .G(n6735), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[3][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][18] ( .G(n6735), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[3][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][17] ( .G(n6735), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[3][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][16] ( .G(n6735), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[3][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][15] ( .G(n6735), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[3][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][14] ( .G(n6735), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[3][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][13] ( .G(n6735), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[3][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][12] ( .G(n6735), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[3][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][11] ( .G(n6735), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[3][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][10] ( .G(n6735), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[3][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][9] ( .G(n6735), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[3][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][8] ( .G(n6735), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[3][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][7] ( .G(n6735), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[3][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][6] ( .G(n6735), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[3][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][5] ( .G(n6735), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[3][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][4] ( .G(n6735), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[3][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][3] ( .G(n6735), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[3][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][2] ( .G(n6735), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[3][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][1] ( .G(n6735), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[3][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[3][0] ( .G(n6735), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[3][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][64] ( .G(n6734), .D(GFtsReq), .Q(\TsBuf[2][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][63] ( .G(n6734), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[2][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][62] ( .G(n6734), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[2][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][61] ( .G(n6734), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[2][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][60] ( .G(n6734), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[2][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][59] ( .G(n6734), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[2][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][58] ( .G(n6734), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[2][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][57] ( .G(n6734), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[2][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][56] ( .G(n6734), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[2][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][55] ( .G(n6734), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[2][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][54] ( .G(n6734), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[2][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][53] ( .G(n6734), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[2][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][52] ( .G(n6734), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[2][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][51] ( .G(n6734), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[2][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][50] ( .G(n6734), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[2][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][49] ( .G(n6734), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[2][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][48] ( .G(n6734), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[2][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][47] ( .G(n6734), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[2][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][46] ( .G(n6734), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[2][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][45] ( .G(n6734), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[2][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][44] ( .G(n6734), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[2][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][43] ( .G(n6734), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[2][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][42] ( .G(n6734), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[2][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][41] ( .G(n6734), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[2][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][40] ( .G(n6734), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[2][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][39] ( .G(n6734), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[2][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][38] ( .G(n6734), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[2][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][37] ( .G(n6734), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[2][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][36] ( .G(n6734), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[2][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][35] ( .G(n6734), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[2][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][34] ( .G(n6734), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[2][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][33] ( .G(n6734), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[2][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][32] ( .G(n6734), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[2][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][31] ( .G(n6734), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[2][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][30] ( .G(n6734), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[2][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][29] ( .G(n6734), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[2][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][28] ( .G(n6734), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[2][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][27] ( .G(n6734), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[2][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][26] ( .G(n6734), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[2][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][25] ( .G(n6734), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[2][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][24] ( .G(n6734), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[2][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][23] ( .G(n6734), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[2][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][22] ( .G(n6734), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[2][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][21] ( .G(n6734), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[2][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][20] ( .G(n6734), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[2][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][19] ( .G(n6734), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[2][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][18] ( .G(n6734), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[2][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][17] ( .G(n6734), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[2][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][16] ( .G(n6734), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[2][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][15] ( .G(n6734), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[2][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][14] ( .G(n6734), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[2][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][13] ( .G(n6734), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[2][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][12] ( .G(n6734), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[2][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][11] ( .G(n6734), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[2][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][10] ( .G(n6734), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[2][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][9] ( .G(n6734), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[2][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][8] ( .G(n6734), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[2][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][7] ( .G(n6734), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[2][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][6] ( .G(n6734), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[2][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][5] ( .G(n6734), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[2][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][4] ( .G(n6734), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[2][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][3] ( .G(n6734), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[2][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][2] ( .G(n6734), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[2][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][1] ( .G(n6734), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[2][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[2][0] ( .G(n6734), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[2][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][64] ( .G(n6733), .D(GFtsReq), .Q(\TsBuf[1][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][63] ( .G(n6733), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[1][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][62] ( .G(n6733), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[1][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][61] ( .G(n6733), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[1][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][60] ( .G(n6733), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[1][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][59] ( .G(n6733), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[1][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][58] ( .G(n6733), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[1][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][57] ( .G(n6733), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[1][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][56] ( .G(n6733), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[1][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][55] ( .G(n6733), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[1][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][54] ( .G(n6733), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[1][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][53] ( .G(n6733), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[1][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][52] ( .G(n6733), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[1][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][51] ( .G(n6733), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[1][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][50] ( .G(n6733), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[1][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][49] ( .G(n6733), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[1][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][48] ( .G(n6733), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[1][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][47] ( .G(n6733), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[1][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][46] ( .G(n6733), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[1][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][45] ( .G(n6733), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[1][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][44] ( .G(n6733), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[1][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][43] ( .G(n6733), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[1][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][42] ( .G(n6733), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[1][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][41] ( .G(n6733), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[1][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][40] ( .G(n6733), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[1][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][39] ( .G(n6733), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[1][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][38] ( .G(n6733), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[1][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][37] ( .G(n6733), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[1][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][36] ( .G(n6733), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[1][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][35] ( .G(n6733), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[1][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][34] ( .G(n6733), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[1][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][33] ( .G(n6733), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[1][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][32] ( .G(n6733), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[1][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][31] ( .G(n6733), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[1][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][30] ( .G(n6733), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[1][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][29] ( .G(n6733), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[1][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][28] ( .G(n6733), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[1][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][27] ( .G(n6733), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[1][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][26] ( .G(n6733), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[1][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][25] ( .G(n6733), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[1][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][24] ( .G(n6733), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[1][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][23] ( .G(n6733), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[1][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][22] ( .G(n6733), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[1][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][21] ( .G(n6733), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[1][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][20] ( .G(n6733), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[1][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][19] ( .G(n6733), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[1][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][18] ( .G(n6733), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[1][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][17] ( .G(n6733), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[1][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][16] ( .G(n6733), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[1][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][15] ( .G(n6733), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[1][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][14] ( .G(n6733), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[1][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][13] ( .G(n6733), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[1][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][12] ( .G(n6733), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[1][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][11] ( .G(n6733), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[1][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][10] ( .G(n6733), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[1][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][9] ( .G(n6733), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[1][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][8] ( .G(n6733), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[1][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][7] ( .G(n6733), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[1][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][6] ( .G(n6733), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[1][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][5] ( .G(n6733), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[1][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][4] ( .G(n6733), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[1][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][3] ( .G(n6733), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[1][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][2] ( .G(n6733), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[1][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][1] ( .G(n6733), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[1][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[1][0] ( .G(n6733), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[1][0] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][64] ( .G(n6740), .D(GFtsReq), .Q(\TsBuf[0][64] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][63] ( .G(n6740), .D(xc_top.ixcSimTime[63]), .Q(\TsBuf[0][63] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][62] ( .G(n6740), .D(xc_top.ixcSimTime[62]), .Q(\TsBuf[0][62] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][61] ( .G(n6740), .D(xc_top.ixcSimTime[61]), .Q(\TsBuf[0][61] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][60] ( .G(n6740), .D(xc_top.ixcSimTime[60]), .Q(\TsBuf[0][60] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][59] ( .G(n6740), .D(xc_top.ixcSimTime[59]), .Q(\TsBuf[0][59] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][58] ( .G(n6740), .D(xc_top.ixcSimTime[58]), .Q(\TsBuf[0][58] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][57] ( .G(n6740), .D(xc_top.ixcSimTime[57]), .Q(\TsBuf[0][57] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][56] ( .G(n6740), .D(xc_top.ixcSimTime[56]), .Q(\TsBuf[0][56] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][55] ( .G(n6740), .D(xc_top.ixcSimTime[55]), .Q(\TsBuf[0][55] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][54] ( .G(n6740), .D(xc_top.ixcSimTime[54]), .Q(\TsBuf[0][54] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][53] ( .G(n6740), .D(xc_top.ixcSimTime[53]), .Q(\TsBuf[0][53] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][52] ( .G(n6740), .D(xc_top.ixcSimTime[52]), .Q(\TsBuf[0][52] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][51] ( .G(n6740), .D(xc_top.ixcSimTime[51]), .Q(\TsBuf[0][51] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][50] ( .G(n6740), .D(xc_top.ixcSimTime[50]), .Q(\TsBuf[0][50] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][49] ( .G(n6740), .D(xc_top.ixcSimTime[49]), .Q(\TsBuf[0][49] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][48] ( .G(n6740), .D(xc_top.ixcSimTime[48]), .Q(\TsBuf[0][48] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][47] ( .G(n6740), .D(xc_top.ixcSimTime[47]), .Q(\TsBuf[0][47] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][46] ( .G(n6740), .D(xc_top.ixcSimTime[46]), .Q(\TsBuf[0][46] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][45] ( .G(n6740), .D(xc_top.ixcSimTime[45]), .Q(\TsBuf[0][45] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][44] ( .G(n6740), .D(xc_top.ixcSimTime[44]), .Q(\TsBuf[0][44] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][43] ( .G(n6740), .D(xc_top.ixcSimTime[43]), .Q(\TsBuf[0][43] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][42] ( .G(n6740), .D(xc_top.ixcSimTime[42]), .Q(\TsBuf[0][42] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][41] ( .G(n6740), .D(xc_top.ixcSimTime[41]), .Q(\TsBuf[0][41] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][40] ( .G(n6740), .D(xc_top.ixcSimTime[40]), .Q(\TsBuf[0][40] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][39] ( .G(n6740), .D(xc_top.ixcSimTime[39]), .Q(\TsBuf[0][39] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][38] ( .G(n6740), .D(xc_top.ixcSimTime[38]), .Q(\TsBuf[0][38] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][37] ( .G(n6740), .D(xc_top.ixcSimTime[37]), .Q(\TsBuf[0][37] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][36] ( .G(n6740), .D(xc_top.ixcSimTime[36]), .Q(\TsBuf[0][36] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][35] ( .G(n6740), .D(xc_top.ixcSimTime[35]), .Q(\TsBuf[0][35] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][34] ( .G(n6740), .D(xc_top.ixcSimTime[34]), .Q(\TsBuf[0][34] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][33] ( .G(n6740), .D(xc_top.ixcSimTime[33]), .Q(\TsBuf[0][33] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][32] ( .G(n6740), .D(xc_top.ixcSimTime[32]), .Q(\TsBuf[0][32] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][31] ( .G(n6740), .D(xc_top.ixcSimTime[31]), .Q(\TsBuf[0][31] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][30] ( .G(n6740), .D(xc_top.ixcSimTime[30]), .Q(\TsBuf[0][30] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][29] ( .G(n6740), .D(xc_top.ixcSimTime[29]), .Q(\TsBuf[0][29] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][28] ( .G(n6740), .D(xc_top.ixcSimTime[28]), .Q(\TsBuf[0][28] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][27] ( .G(n6740), .D(xc_top.ixcSimTime[27]), .Q(\TsBuf[0][27] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][26] ( .G(n6740), .D(xc_top.ixcSimTime[26]), .Q(\TsBuf[0][26] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][25] ( .G(n6740), .D(xc_top.ixcSimTime[25]), .Q(\TsBuf[0][25] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][24] ( .G(n6740), .D(xc_top.ixcSimTime[24]), .Q(\TsBuf[0][24] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][23] ( .G(n6740), .D(xc_top.ixcSimTime[23]), .Q(\TsBuf[0][23] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][22] ( .G(n6740), .D(xc_top.ixcSimTime[22]), .Q(\TsBuf[0][22] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][21] ( .G(n6740), .D(xc_top.ixcSimTime[21]), .Q(\TsBuf[0][21] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][20] ( .G(n6740), .D(xc_top.ixcSimTime[20]), .Q(\TsBuf[0][20] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][19] ( .G(n6740), .D(xc_top.ixcSimTime[19]), .Q(\TsBuf[0][19] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][18] ( .G(n6740), .D(xc_top.ixcSimTime[18]), .Q(\TsBuf[0][18] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][17] ( .G(n6740), .D(xc_top.ixcSimTime[17]), .Q(\TsBuf[0][17] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][16] ( .G(n6740), .D(xc_top.ixcSimTime[16]), .Q(\TsBuf[0][16] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][15] ( .G(n6740), .D(xc_top.ixcSimTime[15]), .Q(\TsBuf[0][15] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][14] ( .G(n6740), .D(xc_top.ixcSimTime[14]), .Q(\TsBuf[0][14] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][13] ( .G(n6740), .D(xc_top.ixcSimTime[13]), .Q(\TsBuf[0][13] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][12] ( .G(n6740), .D(xc_top.ixcSimTime[12]), .Q(\TsBuf[0][12] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][11] ( .G(n6740), .D(xc_top.ixcSimTime[11]), .Q(\TsBuf[0][11] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][10] ( .G(n6740), .D(xc_top.ixcSimTime[10]), .Q(\TsBuf[0][10] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][9] ( .G(n6740), .D(xc_top.ixcSimTime[9]), .Q(\TsBuf[0][9] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][8] ( .G(n6740), .D(xc_top.ixcSimTime[8]), .Q(\TsBuf[0][8] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][7] ( .G(n6740), .D(xc_top.ixcSimTime[7]), .Q(\TsBuf[0][7] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][6] ( .G(n6740), .D(xc_top.ixcSimTime[6]), .Q(\TsBuf[0][6] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][5] ( .G(n6740), .D(xc_top.ixcSimTime[5]), .Q(\TsBuf[0][5] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][4] ( .G(n6740), .D(xc_top.ixcSimTime[4]), .Q(\TsBuf[0][4] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][3] ( .G(n6740), .D(xc_top.ixcSimTime[3]), .Q(\TsBuf[0][3] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][2] ( .G(n6740), .D(xc_top.ixcSimTime[2]), .Q(\TsBuf[0][2] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][1] ( .G(n6740), .D(xc_top.ixcSimTime[1]), .Q(\TsBuf[0][1] ), .QN( ));
Q_LDP0 \TsBuf_REG[0][0] ( .G(n6740), .D(xc_top.ixcSimTime[0]), .Q(\TsBuf[0][0] ), .QN( ));
Q_AN02 U672 ( .A0(n6732), .A1(n6723), .Z(n6739));
Q_AN02 U673 ( .A0(n6732), .A1(n6726), .Z(n6738));
Q_AN02 U674 ( .A0(n6731), .A1(n6723), .Z(n6737));
Q_AN02 U675 ( .A0(n6731), .A1(n6726), .Z(n6736));
Q_AN02 U676 ( .A0(n6730), .A1(n6723), .Z(n6735));
Q_AN02 U677 ( .A0(n6730), .A1(n6726), .Z(n6734));
Q_AN02 U678 ( .A0(n6729), .A1(n6723), .Z(n6733));
Q_AN03 U679 ( .A0(n6729), .A1(n6726), .A2(n3648), .Z(n6740));
Q_AN02 U680 ( .A0(n6725), .A1(n6724), .Z(n6732));
Q_AN02 U681 ( .A0(n6725), .A1(n6727), .Z(n6731));
Q_AN02 U682 ( .A0(n6728), .A1(n6724), .Z(n6730));
Q_NR02 U683 ( .A0(n6725), .A1(n6724), .Z(n6729));
Q_INV U684 ( .A(n6725), .Z(n6728));
Q_INV U685 ( .A(n6724), .Z(n6727));
Q_INV U686 ( .A(n6723), .Z(n6726));
Q_AN02 U687 ( .A0(LBwr[2]), .A1(n3648), .Z(n6725));
Q_AN02 U688 ( .A0(LBwr[1]), .A1(n3648), .Z(n6724));
Q_AN02 U689 ( .A0(LBwr[0]), .A1(n3648), .Z(n6723));
Q_FDP0UA U690 ( .D(svGFbusy1), .QTFCLK( ), .Q(svGFbusy2));
Q_INV U691 ( .A(LBreq), .Z(n6717));
Q_ND02 U692 ( .A0(LBreq), .A1(n1610), .Z(n6712));
Q_INV U693 ( .A(xc_top.GFReset), .Z(n6720));
Q_AN02 U694 ( .A0(n6720), .A1(n6712), .Z(n6716));
Q_INV U695 ( .A(GFreq), .Z(n6715));
Q_AN03 U696 ( .A0(n6715), .A1(svGFbusy1), .A2(n6714), .Z(n6713));
Q_INV U697 ( .A(gfTsEn), .Z(n6714));
Q_OR02 U698 ( .A0(n6713), .A1(xc_top.GFReset), .Z(n6722));
Q_AN02 U699 ( .A0(n6720), .A1(n6713), .Z(n6719));
Q_INV U700 ( .A(n6722), .Z(n6721));
Q_INV U701 ( .A(n6712), .Z(n6718));
Q_FDP0UA U702 ( .D(n6719), .QTFCLK( ), .Q(gfTsEn));
Q_FDP0UA U703 ( .D(n6697), .QTFCLK( ), .Q(LBfill[0]));
Q_FDP0UA U704 ( .D(n6699), .QTFCLK( ), .Q(LBfill[1]));
Q_FDP0UA U705 ( .D(n6701), .QTFCLK( ), .Q(LBfill[2]));
Q_FDP0UA U706 ( .D(n6703), .QTFCLK( ), .Q(LBfill[3]));
Q_MX02 U707 ( .S(n6716), .A0(n6688), .A1(LBwrI[0]), .Z(n6711));
Q_FDP0UA U708 ( .D(n6711), .QTFCLK( ), .Q(LBwrI[0]));
Q_MX02 U709 ( .S(n6716), .A0(n6689), .A1(LBwrI[1]), .Z(n6710));
Q_FDP0UA U710 ( .D(n6710), .QTFCLK( ), .Q(LBwrI[1]));
Q_MX02 U711 ( .S(n6716), .A0(n6690), .A1(LBwrI[2]), .Z(n6709));
Q_FDP0UA U712 ( .D(n6709), .QTFCLK( ), .Q(LBwrI[2]));
Q_MX02 U713 ( .S(n6716), .A0(n6691), .A1(LBwrI[3]), .Z(n6708));
Q_FDP0UA U714 ( .D(n6708), .QTFCLK( ), .Q(LBwrI[3]));
Q_MX02 U715 ( .S(n6722), .A0(LBrd[0]), .A1(n6692), .Z(n6707));
Q_FDP0UA U716 ( .D(n6707), .QTFCLK( ), .Q(LBrd[0]));
Q_MX02 U717 ( .S(n6722), .A0(LBrd[1]), .A1(n6693), .Z(n6706));
Q_FDP0UA U718 ( .D(n6706), .QTFCLK( ), .Q(LBrd[1]));
Q_MX02 U719 ( .S(n6722), .A0(LBrd[2]), .A1(n6694), .Z(n6705));
Q_FDP0UA U720 ( .D(n6705), .QTFCLK( ), .Q(LBrd[2]));
Q_MX02 U721 ( .S(n6722), .A0(LBrd[3]), .A1(n6695), .Z(n6704));
Q_FDP0UA U722 ( .D(n6704), .QTFCLK( ), .Q(LBrd[3]));
Q_MX02 U723 ( .S(n6719), .A0(n6702), .A1(n6687), .Z(n6703));
Q_AN02 U724 ( .A0(n6721), .A1(n6681), .Z(n6702));
Q_MX02 U725 ( .S(n6719), .A0(n6700), .A1(n6685), .Z(n6701));
Q_AN02 U726 ( .A0(n6721), .A1(n6680), .Z(n6700));
Q_MX02 U727 ( .S(n6719), .A0(n6698), .A1(n6683), .Z(n6699));
Q_AN02 U728 ( .A0(n6721), .A1(n6679), .Z(n6698));
Q_MX02 U729 ( .S(n6719), .A0(n6696), .A1(n6682), .Z(n6697));
Q_AN02 U730 ( .A0(n6721), .A1(n6678), .Z(n6696));
Q_XNR2 U731 ( .A0(n6681), .A1(n6686), .Z(n6687));
Q_OR02 U732 ( .A0(n6680), .A1(n6684), .Z(n6686));
Q_XNR2 U733 ( .A0(n6680), .A1(n6684), .Z(n6685));
Q_OR02 U734 ( .A0(n6678), .A1(n6679), .Z(n6684));
Q_XNR2 U735 ( .A0(n6678), .A1(n6679), .Z(n6683));
Q_INV U736 ( .A(n6678), .Z(n6682));
Q_MX02 U737 ( .S(n6712), .A0(n6676), .A1(LBfill[2]), .Z(n6680));
Q_MX02 U738 ( .S(n6712), .A0(n6674), .A1(LBfill[1]), .Z(n6679));
Q_XOR2 U739 ( .A0(n6718), .A1(LBfill[0]), .Z(n6678));
Q_XOR2 U740 ( .A0(LBfill[3]), .A1(n6741), .Z(n6681));
Q_AD01HF U741 ( .A0(LBfill[2]), .B0(n6675), .S(n6676), .CO(n6677));
Q_AD01HF U742 ( .A0(LBfill[1]), .B0(LBfill[0]), .S(n6674), .CO(n6675));
Q_AN03 U743 ( .A0(n6673), .A1(n6669), .A2(n6720), .Z(n6691));
Q_AN03 U744 ( .A0(n6673), .A1(n6667), .A2(n6720), .Z(n6690));
Q_AN03 U745 ( .A0(n6673), .A1(n6665), .A2(n6720), .Z(n6689));
Q_AN03 U746 ( .A0(n6673), .A1(n6664), .A2(n6720), .Z(n6688));
Q_OR03 U747 ( .A0(n6671), .A1(n6669), .A2(n6672), .Z(n6673));
Q_OR03 U748 ( .A0(n6670), .A1(n6664), .A2(n6665), .Z(n6672));
Q_INV U749 ( .A(n6667), .Z(n6671));
Q_AD01HF U750 ( .A0(LBwrI[3]), .B0(n6668), .S(n6669), .CO(n6670));
Q_AD01HF U751 ( .A0(LBwrI[2]), .B0(n6666), .S(n6667), .CO(n6668));
Q_AD01HF U752 ( .A0(LBwrI[1]), .B0(LBwrI[0]), .S(n6665), .CO(n6666));
Q_INV U753 ( .A(LBwrI[0]), .Z(n6664));
Q_AN03 U754 ( .A0(n6663), .A1(n6659), .A2(n6720), .Z(n6695));
Q_AN03 U755 ( .A0(n6663), .A1(n6657), .A2(n6720), .Z(n6694));
Q_AN03 U756 ( .A0(n6663), .A1(n6655), .A2(n6720), .Z(n6693));
Q_AN03 U757 ( .A0(n6663), .A1(n6654), .A2(n6720), .Z(n6692));
Q_OR03 U758 ( .A0(n6661), .A1(n6659), .A2(n6662), .Z(n6663));
Q_OR03 U759 ( .A0(n6660), .A1(n6654), .A2(n6655), .Z(n6662));
Q_INV U760 ( .A(n6657), .Z(n6661));
Q_AD01HF U761 ( .A0(LBrd[3]), .B0(n6658), .S(n6659), .CO(n6660));
Q_AD01HF U762 ( .A0(LBrd[2]), .B0(n6656), .S(n6657), .CO(n6658));
Q_AD01HF U763 ( .A0(LBrd[1]), .B0(LBrd[0]), .S(n6655), .CO(n6656));
Q_INV U764 ( .A(LBrd[0]), .Z(n6654));
Q_FDP0UA U765 ( .D(n5824), .QTFCLK( ), .Q(ofifoWptr[0]));
Q_FDP0UA U766 ( .D(n5825), .QTFCLK( ), .Q(ofifoWptr[1]));
Q_FDP0UA U767 ( .D(n5826), .QTFCLK( ), .Q(ofifoWptr[2]));
Q_FDP0UA U768 ( .D(n5827), .QTFCLK( ), .Q(ofifoWptr[3]));
Q_FDP0UA U769 ( .D(n5828), .QTFCLK( ), .Q(ofifoWptr[4]));
Q_FDP0UA U770 ( .D(n5829), .QTFCLK( ), .Q(ofifoWptr[5]));
Q_FDP0UA U771 ( .D(n5830), .QTFCLK( ), .Q(ofifoWptr[6]));
Q_FDP0UA U772 ( .D(n5831), .QTFCLK( ), .Q(ofifoWptr[7]));
Q_FDP0UA U773 ( .D(n5832), .QTFCLK( ), .Q(ofifoWptr[8]));
Q_FDP0UA U774 ( .D(n5833), .QTFCLK( ), .Q(ofifoWptr[9]));
Q_FDP0UA U775 ( .D(n5834), .QTFCLK( ), .Q(ofifoWptr[10]));
Q_FDP0UA U776 ( .D(n5835), .QTFCLK( ), .Q(ofifoWptr[11]));
Q_FDP0UA U777 ( .D(n5836), .QTFCLK( ), .Q(ofifoWptr[12]));
Q_FDP0UA U778 ( .D(n5837), .QTFCLK( ), .Q(ofifoWptr[13]));
Q_FDP0UA U779 ( .D(n5838), .QTFCLK( ), .Q(ofifoWptr[14]));
Q_FDP0UA U780 ( .D(n5839), .QTFCLK( ), .Q(oFill[0]));
Q_FDP0UA U781 ( .D(n5840), .QTFCLK( ), .Q(oFill[1]));
Q_FDP0UA U782 ( .D(n5841), .QTFCLK( ), .Q(oFill[2]));
Q_FDP0UA U783 ( .D(n5842), .QTFCLK( ), .Q(oFill[3]));
Q_FDP0UA U784 ( .D(n5843), .QTFCLK( ), .Q(oFill[4]));
Q_FDP0UA U785 ( .D(n5844), .QTFCLK( ), .Q(ofifoData[0]));
Q_FDP0UA U786 ( .D(n5845), .QTFCLK( ), .Q(ofifoData[1]));
Q_FDP0UA U787 ( .D(n5846), .QTFCLK( ), .Q(ofifoData[2]));
Q_FDP0UA U788 ( .D(n5847), .QTFCLK( ), .Q(ofifoData[3]));
Q_FDP0UA U789 ( .D(n5848), .QTFCLK( ), .Q(ofifoData[4]));
Q_FDP0UA U790 ( .D(n5849), .QTFCLK( ), .Q(ofifoData[5]));
Q_FDP0UA U791 ( .D(n5850), .QTFCLK( ), .Q(ofifoData[6]));
Q_FDP0UA U792 ( .D(n5851), .QTFCLK( ), .Q(ofifoData[7]));
Q_FDP0UA U793 ( .D(n5852), .QTFCLK( ), .Q(ofifoData[8]));
Q_FDP0UA U794 ( .D(n5853), .QTFCLK( ), .Q(ofifoData[9]));
Q_FDP0UA U795 ( .D(n5854), .QTFCLK( ), .Q(ofifoData[10]));
Q_FDP0UA U796 ( .D(n5855), .QTFCLK( ), .Q(ofifoData[11]));
Q_FDP0UA U797 ( .D(n5856), .QTFCLK( ), .Q(ofifoData[12]));
Q_FDP0UA U798 ( .D(n5857), .QTFCLK( ), .Q(ofifoData[13]));
Q_FDP0UA U799 ( .D(n5858), .QTFCLK( ), .Q(ofifoData[14]));
Q_FDP0UA U800 ( .D(n5859), .QTFCLK( ), .Q(ofifoData[15]));
Q_FDP0UA U801 ( .D(n5860), .QTFCLK( ), .Q(ofifoData[16]));
Q_FDP0UA U802 ( .D(n5861), .QTFCLK( ), .Q(ofifoData[17]));
Q_FDP0UA U803 ( .D(n5862), .QTFCLK( ), .Q(ofifoData[18]));
Q_FDP0UA U804 ( .D(n5863), .QTFCLK( ), .Q(ofifoData[19]));
Q_FDP0UA U805 ( .D(n5864), .QTFCLK( ), .Q(ofifoData[20]));
Q_FDP0UA U806 ( .D(n5865), .QTFCLK( ), .Q(ofifoData[21]));
Q_FDP0UA U807 ( .D(n5866), .QTFCLK( ), .Q(ofifoData[22]));
Q_FDP0UA U808 ( .D(n5867), .QTFCLK( ), .Q(ofifoData[23]));
Q_FDP0UA U809 ( .D(n5868), .QTFCLK( ), .Q(ofifoData[24]));
Q_FDP0UA U810 ( .D(n5869), .QTFCLK( ), .Q(ofifoData[25]));
Q_FDP0UA U811 ( .D(n5870), .QTFCLK( ), .Q(ofifoData[26]));
Q_FDP0UA U812 ( .D(n5871), .QTFCLK( ), .Q(ofifoData[27]));
Q_FDP0UA U813 ( .D(n5872), .QTFCLK( ), .Q(ofifoData[28]));
Q_FDP0UA U814 ( .D(n5873), .QTFCLK( ), .Q(ofifoData[29]));
Q_FDP0UA U815 ( .D(n5874), .QTFCLK( ), .Q(ofifoData[30]));
Q_FDP0UA U816 ( .D(n5875), .QTFCLK( ), .Q(ofifoData[31]));
Q_FDP0UA U817 ( .D(n5876), .QTFCLK( ), .Q(ofifoData[32]));
Q_FDP0UA U818 ( .D(n5877), .QTFCLK( ), .Q(ofifoData[33]));
Q_FDP0UA U819 ( .D(n5878), .QTFCLK( ), .Q(ofifoData[34]));
Q_FDP0UA U820 ( .D(n5879), .QTFCLK( ), .Q(ofifoData[35]));
Q_FDP0UA U821 ( .D(n5880), .QTFCLK( ), .Q(ofifoData[36]));
Q_FDP0UA U822 ( .D(n5881), .QTFCLK( ), .Q(ofifoData[37]));
Q_FDP0UA U823 ( .D(n5882), .QTFCLK( ), .Q(ofifoData[38]));
Q_FDP0UA U824 ( .D(n5883), .QTFCLK( ), .Q(ofifoData[39]));
Q_FDP0UA U825 ( .D(n5884), .QTFCLK( ), .Q(ofifoData[40]));
Q_FDP0UA U826 ( .D(n5885), .QTFCLK( ), .Q(ofifoData[41]));
Q_FDP0UA U827 ( .D(n5886), .QTFCLK( ), .Q(ofifoData[42]));
Q_FDP0UA U828 ( .D(n5887), .QTFCLK( ), .Q(ofifoData[43]));
Q_FDP0UA U829 ( .D(n5888), .QTFCLK( ), .Q(ofifoData[44]));
Q_FDP0UA U830 ( .D(n5889), .QTFCLK( ), .Q(ofifoData[45]));
Q_FDP0UA U831 ( .D(n5890), .QTFCLK( ), .Q(ofifoData[46]));
Q_FDP0UA U832 ( .D(n5891), .QTFCLK( ), .Q(ofifoData[47]));
Q_FDP0UA U833 ( .D(n5892), .QTFCLK( ), .Q(ofifoData[48]));
Q_FDP0UA U834 ( .D(n5893), .QTFCLK( ), .Q(ofifoData[49]));
Q_FDP0UA U835 ( .D(n5894), .QTFCLK( ), .Q(ofifoData[50]));
Q_FDP0UA U836 ( .D(n5895), .QTFCLK( ), .Q(ofifoData[51]));
Q_FDP0UA U837 ( .D(n5896), .QTFCLK( ), .Q(ofifoData[52]));
Q_FDP0UA U838 ( .D(n5897), .QTFCLK( ), .Q(ofifoData[53]));
Q_FDP0UA U839 ( .D(n5898), .QTFCLK( ), .Q(ofifoData[54]));
Q_FDP0UA U840 ( .D(n5899), .QTFCLK( ), .Q(ofifoData[55]));
Q_FDP0UA U841 ( .D(n5900), .QTFCLK( ), .Q(ofifoData[56]));
Q_FDP0UA U842 ( .D(n5901), .QTFCLK( ), .Q(ofifoData[57]));
Q_FDP0UA U843 ( .D(n5902), .QTFCLK( ), .Q(ofifoData[58]));
Q_FDP0UA U844 ( .D(n5903), .QTFCLK( ), .Q(ofifoData[59]));
Q_FDP0UA U845 ( .D(n5904), .QTFCLK( ), .Q(ofifoData[60]));
Q_FDP0UA U846 ( .D(n5905), .QTFCLK( ), .Q(ofifoData[61]));
Q_FDP0UA U847 ( .D(n5906), .QTFCLK( ), .Q(ofifoData[62]));
Q_FDP0UA U848 ( .D(n5907), .QTFCLK( ), .Q(ofifoData[63]));
Q_FDP0UA U849 ( .D(n5908), .QTFCLK( ), .Q(ofifoData[64]));
Q_FDP0UA U850 ( .D(n5909), .QTFCLK( ), .Q(ofifoData[65]));
Q_FDP0UA U851 ( .D(n5910), .QTFCLK( ), .Q(ofifoData[66]));
Q_FDP0UA U852 ( .D(n5911), .QTFCLK( ), .Q(ofifoData[67]));
Q_FDP0UA U853 ( .D(n5912), .QTFCLK( ), .Q(ofifoData[68]));
Q_FDP0UA U854 ( .D(n5913), .QTFCLK( ), .Q(ofifoData[69]));
Q_FDP0UA U855 ( .D(n5914), .QTFCLK( ), .Q(ofifoData[70]));
Q_FDP0UA U856 ( .D(n5915), .QTFCLK( ), .Q(ofifoData[71]));
Q_FDP0UA U857 ( .D(n5916), .QTFCLK( ), .Q(ofifoData[72]));
Q_FDP0UA U858 ( .D(n5917), .QTFCLK( ), .Q(ofifoData[73]));
Q_FDP0UA U859 ( .D(n5918), .QTFCLK( ), .Q(ofifoData[74]));
Q_FDP0UA U860 ( .D(n5919), .QTFCLK( ), .Q(ofifoData[75]));
Q_FDP0UA U861 ( .D(n5920), .QTFCLK( ), .Q(ofifoData[76]));
Q_FDP0UA U862 ( .D(n5921), .QTFCLK( ), .Q(ofifoData[77]));
Q_FDP0UA U863 ( .D(n5922), .QTFCLK( ), .Q(ofifoData[78]));
Q_FDP0UA U864 ( .D(n5923), .QTFCLK( ), .Q(ofifoData[79]));
Q_FDP0UA U865 ( .D(n5924), .QTFCLK( ), .Q(ofifoData[80]));
Q_FDP0UA U866 ( .D(n5925), .QTFCLK( ), .Q(ofifoData[81]));
Q_FDP0UA U867 ( .D(n5926), .QTFCLK( ), .Q(ofifoData[82]));
Q_FDP0UA U868 ( .D(n5927), .QTFCLK( ), .Q(ofifoData[83]));
Q_FDP0UA U869 ( .D(n5928), .QTFCLK( ), .Q(ofifoData[84]));
Q_FDP0UA U870 ( .D(n5929), .QTFCLK( ), .Q(ofifoData[85]));
Q_FDP0UA U871 ( .D(n5930), .QTFCLK( ), .Q(ofifoData[86]));
Q_FDP0UA U872 ( .D(n5931), .QTFCLK( ), .Q(ofifoData[87]));
Q_FDP0UA U873 ( .D(n5932), .QTFCLK( ), .Q(ofifoData[88]));
Q_FDP0UA U874 ( .D(n5933), .QTFCLK( ), .Q(ofifoData[89]));
Q_FDP0UA U875 ( .D(n5934), .QTFCLK( ), .Q(ofifoData[90]));
Q_FDP0UA U876 ( .D(n5935), .QTFCLK( ), .Q(ofifoData[91]));
Q_FDP0UA U877 ( .D(n5936), .QTFCLK( ), .Q(ofifoData[92]));
Q_FDP0UA U878 ( .D(n5937), .QTFCLK( ), .Q(ofifoData[93]));
Q_FDP0UA U879 ( .D(n5938), .QTFCLK( ), .Q(ofifoData[94]));
Q_FDP0UA U880 ( .D(n5939), .QTFCLK( ), .Q(ofifoData[95]));
Q_FDP0UA U881 ( .D(n5940), .QTFCLK( ), .Q(ofifoData[96]));
Q_FDP0UA U882 ( .D(n5941), .QTFCLK( ), .Q(ofifoData[97]));
Q_FDP0UA U883 ( .D(n5942), .QTFCLK( ), .Q(ofifoData[98]));
Q_FDP0UA U884 ( .D(n5943), .QTFCLK( ), .Q(ofifoData[99]));
Q_FDP0UA U885 ( .D(n5944), .QTFCLK( ), .Q(ofifoData[100]));
Q_FDP0UA U886 ( .D(n5945), .QTFCLK( ), .Q(ofifoData[101]));
Q_FDP0UA U887 ( .D(n5946), .QTFCLK( ), .Q(ofifoData[102]));
Q_FDP0UA U888 ( .D(n5947), .QTFCLK( ), .Q(ofifoData[103]));
Q_FDP0UA U889 ( .D(n5948), .QTFCLK( ), .Q(ofifoData[104]));
Q_FDP0UA U890 ( .D(n5949), .QTFCLK( ), .Q(ofifoData[105]));
Q_FDP0UA U891 ( .D(n5950), .QTFCLK( ), .Q(ofifoData[106]));
Q_FDP0UA U892 ( .D(n5951), .QTFCLK( ), .Q(ofifoData[107]));
Q_FDP0UA U893 ( .D(n5952), .QTFCLK( ), .Q(ofifoData[108]));
Q_FDP0UA U894 ( .D(n5953), .QTFCLK( ), .Q(ofifoData[109]));
Q_FDP0UA U895 ( .D(n5954), .QTFCLK( ), .Q(ofifoData[110]));
Q_FDP0UA U896 ( .D(n5955), .QTFCLK( ), .Q(ofifoData[111]));
Q_FDP0UA U897 ( .D(n5956), .QTFCLK( ), .Q(ofifoData[112]));
Q_FDP0UA U898 ( .D(n5957), .QTFCLK( ), .Q(ofifoData[113]));
Q_FDP0UA U899 ( .D(n5958), .QTFCLK( ), .Q(ofifoData[114]));
Q_FDP0UA U900 ( .D(n5959), .QTFCLK( ), .Q(ofifoData[115]));
Q_FDP0UA U901 ( .D(n5960), .QTFCLK( ), .Q(ofifoData[116]));
Q_FDP0UA U902 ( .D(n5961), .QTFCLK( ), .Q(ofifoData[117]));
Q_FDP0UA U903 ( .D(n5962), .QTFCLK( ), .Q(ofifoData[118]));
Q_FDP0UA U904 ( .D(n5963), .QTFCLK( ), .Q(ofifoData[119]));
Q_FDP0UA U905 ( .D(n5964), .QTFCLK( ), .Q(ofifoData[120]));
Q_FDP0UA U906 ( .D(n5965), .QTFCLK( ), .Q(ofifoData[121]));
Q_FDP0UA U907 ( .D(n5966), .QTFCLK( ), .Q(ofifoData[122]));
Q_FDP0UA U908 ( .D(n5967), .QTFCLK( ), .Q(ofifoData[123]));
Q_FDP0UA U909 ( .D(n5968), .QTFCLK( ), .Q(ofifoData[124]));
Q_FDP0UA U910 ( .D(n5969), .QTFCLK( ), .Q(ofifoData[125]));
Q_FDP0UA U911 ( .D(n5970), .QTFCLK( ), .Q(ofifoData[126]));
Q_FDP0UA U912 ( .D(n5971), .QTFCLK( ), .Q(ofifoData[127]));
Q_FDP0UA U913 ( .D(n5972), .QTFCLK( ), .Q(ofifoData[128]));
Q_FDP0UA U914 ( .D(n5973), .QTFCLK( ), .Q(ofifoData[129]));
Q_FDP0UA U915 ( .D(n5974), .QTFCLK( ), .Q(ofifoData[130]));
Q_FDP0UA U916 ( .D(n5975), .QTFCLK( ), .Q(ofifoData[131]));
Q_FDP0UA U917 ( .D(n5976), .QTFCLK( ), .Q(ofifoData[132]));
Q_FDP0UA U918 ( .D(n5977), .QTFCLK( ), .Q(ofifoData[133]));
Q_FDP0UA U919 ( .D(n5978), .QTFCLK( ), .Q(ofifoData[134]));
Q_FDP0UA U920 ( .D(n5979), .QTFCLK( ), .Q(ofifoData[135]));
Q_FDP0UA U921 ( .D(n5980), .QTFCLK( ), .Q(ofifoData[136]));
Q_FDP0UA U922 ( .D(n5981), .QTFCLK( ), .Q(ofifoData[137]));
Q_FDP0UA U923 ( .D(n5982), .QTFCLK( ), .Q(ofifoData[138]));
Q_FDP0UA U924 ( .D(n5983), .QTFCLK( ), .Q(ofifoData[139]));
Q_FDP0UA U925 ( .D(n5984), .QTFCLK( ), .Q(ofifoData[140]));
Q_FDP0UA U926 ( .D(n5985), .QTFCLK( ), .Q(ofifoData[141]));
Q_FDP0UA U927 ( .D(n5986), .QTFCLK( ), .Q(ofifoData[142]));
Q_FDP0UA U928 ( .D(n5987), .QTFCLK( ), .Q(ofifoData[143]));
Q_FDP0UA U929 ( .D(n5988), .QTFCLK( ), .Q(ofifoData[144]));
Q_FDP0UA U930 ( .D(n5989), .QTFCLK( ), .Q(ofifoData[145]));
Q_FDP0UA U931 ( .D(n5990), .QTFCLK( ), .Q(ofifoData[146]));
Q_FDP0UA U932 ( .D(n5991), .QTFCLK( ), .Q(ofifoData[147]));
Q_FDP0UA U933 ( .D(n5992), .QTFCLK( ), .Q(ofifoData[148]));
Q_FDP0UA U934 ( .D(n5993), .QTFCLK( ), .Q(ofifoData[149]));
Q_FDP0UA U935 ( .D(n5994), .QTFCLK( ), .Q(ofifoData[150]));
Q_FDP0UA U936 ( .D(n5995), .QTFCLK( ), .Q(ofifoData[151]));
Q_FDP0UA U937 ( .D(n5996), .QTFCLK( ), .Q(ofifoData[152]));
Q_FDP0UA U938 ( .D(n5997), .QTFCLK( ), .Q(ofifoData[153]));
Q_FDP0UA U939 ( .D(n5998), .QTFCLK( ), .Q(ofifoData[154]));
Q_FDP0UA U940 ( .D(n5999), .QTFCLK( ), .Q(ofifoData[155]));
Q_FDP0UA U941 ( .D(n6000), .QTFCLK( ), .Q(ofifoData[156]));
Q_FDP0UA U942 ( .D(n6001), .QTFCLK( ), .Q(ofifoData[157]));
Q_FDP0UA U943 ( .D(n6002), .QTFCLK( ), .Q(ofifoData[158]));
Q_FDP0UA U944 ( .D(n6003), .QTFCLK( ), .Q(ofifoData[159]));
Q_FDP0UA U945 ( .D(n6004), .QTFCLK( ), .Q(ofifoData[160]));
Q_FDP0UA U946 ( .D(n6005), .QTFCLK( ), .Q(ofifoData[161]));
Q_FDP0UA U947 ( .D(n6006), .QTFCLK( ), .Q(ofifoData[162]));
Q_FDP0UA U948 ( .D(n6007), .QTFCLK( ), .Q(ofifoData[163]));
Q_FDP0UA U949 ( .D(n6008), .QTFCLK( ), .Q(ofifoData[164]));
Q_FDP0UA U950 ( .D(n6009), .QTFCLK( ), .Q(ofifoData[165]));
Q_FDP0UA U951 ( .D(n6010), .QTFCLK( ), .Q(ofifoData[166]));
Q_FDP0UA U952 ( .D(n6011), .QTFCLK( ), .Q(ofifoData[167]));
Q_FDP0UA U953 ( .D(n6012), .QTFCLK( ), .Q(ofifoData[168]));
Q_FDP0UA U954 ( .D(n6013), .QTFCLK( ), .Q(ofifoData[169]));
Q_FDP0UA U955 ( .D(n6014), .QTFCLK( ), .Q(ofifoData[170]));
Q_FDP0UA U956 ( .D(n6015), .QTFCLK( ), .Q(ofifoData[171]));
Q_FDP0UA U957 ( .D(n6016), .QTFCLK( ), .Q(ofifoData[172]));
Q_FDP0UA U958 ( .D(n6017), .QTFCLK( ), .Q(ofifoData[173]));
Q_FDP0UA U959 ( .D(n6018), .QTFCLK( ), .Q(ofifoData[174]));
Q_FDP0UA U960 ( .D(n6019), .QTFCLK( ), .Q(ofifoData[175]));
Q_FDP0UA U961 ( .D(n6020), .QTFCLK( ), .Q(ofifoData[176]));
Q_FDP0UA U962 ( .D(n6021), .QTFCLK( ), .Q(ofifoData[177]));
Q_FDP0UA U963 ( .D(n6022), .QTFCLK( ), .Q(ofifoData[178]));
Q_FDP0UA U964 ( .D(n6023), .QTFCLK( ), .Q(ofifoData[179]));
Q_FDP0UA U965 ( .D(n6024), .QTFCLK( ), .Q(ofifoData[180]));
Q_FDP0UA U966 ( .D(n6025), .QTFCLK( ), .Q(ofifoData[181]));
Q_FDP0UA U967 ( .D(n6026), .QTFCLK( ), .Q(ofifoData[182]));
Q_FDP0UA U968 ( .D(n6027), .QTFCLK( ), .Q(ofifoData[183]));
Q_FDP0UA U969 ( .D(n6028), .QTFCLK( ), .Q(ofifoData[184]));
Q_FDP0UA U970 ( .D(n6029), .QTFCLK( ), .Q(ofifoData[185]));
Q_FDP0UA U971 ( .D(n6030), .QTFCLK( ), .Q(ofifoData[186]));
Q_FDP0UA U972 ( .D(n6031), .QTFCLK( ), .Q(ofifoData[187]));
Q_FDP0UA U973 ( .D(n6032), .QTFCLK( ), .Q(ofifoData[188]));
Q_FDP0UA U974 ( .D(n6033), .QTFCLK( ), .Q(ofifoData[189]));
Q_FDP0UA U975 ( .D(n6034), .QTFCLK( ), .Q(ofifoData[190]));
Q_FDP0UA U976 ( .D(n6035), .QTFCLK( ), .Q(ofifoData[191]));
Q_FDP0UA U977 ( .D(n6036), .QTFCLK( ), .Q(ofifoData[192]));
Q_FDP0UA U978 ( .D(n6037), .QTFCLK( ), .Q(ofifoData[193]));
Q_FDP0UA U979 ( .D(n6038), .QTFCLK( ), .Q(ofifoData[194]));
Q_FDP0UA U980 ( .D(n6039), .QTFCLK( ), .Q(ofifoData[195]));
Q_FDP0UA U981 ( .D(n6040), .QTFCLK( ), .Q(ofifoData[196]));
Q_FDP0UA U982 ( .D(n6041), .QTFCLK( ), .Q(ofifoData[197]));
Q_FDP0UA U983 ( .D(n6042), .QTFCLK( ), .Q(ofifoData[198]));
Q_FDP0UA U984 ( .D(n6043), .QTFCLK( ), .Q(ofifoData[199]));
Q_FDP0UA U985 ( .D(n6044), .QTFCLK( ), .Q(ofifoData[200]));
Q_FDP0UA U986 ( .D(n6045), .QTFCLK( ), .Q(ofifoData[201]));
Q_FDP0UA U987 ( .D(n6046), .QTFCLK( ), .Q(ofifoData[202]));
Q_FDP0UA U988 ( .D(n6047), .QTFCLK( ), .Q(ofifoData[203]));
Q_FDP0UA U989 ( .D(n6048), .QTFCLK( ), .Q(ofifoData[204]));
Q_FDP0UA U990 ( .D(n6049), .QTFCLK( ), .Q(ofifoData[205]));
Q_FDP0UA U991 ( .D(n6050), .QTFCLK( ), .Q(ofifoData[206]));
Q_FDP0UA U992 ( .D(n6051), .QTFCLK( ), .Q(ofifoData[207]));
Q_FDP0UA U993 ( .D(n6052), .QTFCLK( ), .Q(ofifoData[208]));
Q_FDP0UA U994 ( .D(n6053), .QTFCLK( ), .Q(ofifoData[209]));
Q_FDP0UA U995 ( .D(n6054), .QTFCLK( ), .Q(ofifoData[210]));
Q_FDP0UA U996 ( .D(n6055), .QTFCLK( ), .Q(ofifoData[211]));
Q_FDP0UA U997 ( .D(n6056), .QTFCLK( ), .Q(ofifoData[212]));
Q_FDP0UA U998 ( .D(n6057), .QTFCLK( ), .Q(ofifoData[213]));
Q_FDP0UA U999 ( .D(n6058), .QTFCLK( ), .Q(ofifoData[214]));
Q_FDP0UA U1000 ( .D(n6059), .QTFCLK( ), .Q(ofifoData[215]));
Q_FDP0UA U1001 ( .D(n6060), .QTFCLK( ), .Q(ofifoData[216]));
Q_FDP0UA U1002 ( .D(n6061), .QTFCLK( ), .Q(ofifoData[217]));
Q_FDP0UA U1003 ( .D(n6062), .QTFCLK( ), .Q(ofifoData[218]));
Q_FDP0UA U1004 ( .D(n6063), .QTFCLK( ), .Q(ofifoData[219]));
Q_FDP0UA U1005 ( .D(n6064), .QTFCLK( ), .Q(ofifoData[220]));
Q_FDP0UA U1006 ( .D(n6065), .QTFCLK( ), .Q(ofifoData[221]));
Q_FDP0UA U1007 ( .D(n6066), .QTFCLK( ), .Q(ofifoData[222]));
Q_FDP0UA U1008 ( .D(n6067), .QTFCLK( ), .Q(ofifoData[223]));
Q_FDP0UA U1009 ( .D(n6068), .QTFCLK( ), .Q(ofifoData[224]));
Q_FDP0UA U1010 ( .D(n6069), .QTFCLK( ), .Q(ofifoData[225]));
Q_FDP0UA U1011 ( .D(n6070), .QTFCLK( ), .Q(ofifoData[226]));
Q_FDP0UA U1012 ( .D(n6071), .QTFCLK( ), .Q(ofifoData[227]));
Q_FDP0UA U1013 ( .D(n6072), .QTFCLK( ), .Q(ofifoData[228]));
Q_FDP0UA U1014 ( .D(n6073), .QTFCLK( ), .Q(ofifoData[229]));
Q_FDP0UA U1015 ( .D(n6074), .QTFCLK( ), .Q(ofifoData[230]));
Q_FDP0UA U1016 ( .D(n6075), .QTFCLK( ), .Q(ofifoData[231]));
Q_FDP0UA U1017 ( .D(n6076), .QTFCLK( ), .Q(ofifoData[232]));
Q_FDP0UA U1018 ( .D(n6077), .QTFCLK( ), .Q(ofifoData[233]));
Q_FDP0UA U1019 ( .D(n6078), .QTFCLK( ), .Q(ofifoData[234]));
Q_FDP0UA U1020 ( .D(n6079), .QTFCLK( ), .Q(ofifoData[235]));
Q_FDP0UA U1021 ( .D(n6080), .QTFCLK( ), .Q(ofifoData[236]));
Q_FDP0UA U1022 ( .D(n6081), .QTFCLK( ), .Q(ofifoData[237]));
Q_FDP0UA U1023 ( .D(n6082), .QTFCLK( ), .Q(ofifoData[238]));
Q_FDP0UA U1024 ( .D(n6083), .QTFCLK( ), .Q(ofifoData[239]));
Q_FDP0UA U1025 ( .D(n6084), .QTFCLK( ), .Q(ofifoData[240]));
Q_FDP0UA U1026 ( .D(n6085), .QTFCLK( ), .Q(ofifoData[241]));
Q_FDP0UA U1027 ( .D(n6086), .QTFCLK( ), .Q(ofifoData[242]));
Q_FDP0UA U1028 ( .D(n6087), .QTFCLK( ), .Q(ofifoData[243]));
Q_FDP0UA U1029 ( .D(n6088), .QTFCLK( ), .Q(ofifoData[244]));
Q_FDP0UA U1030 ( .D(n6089), .QTFCLK( ), .Q(ofifoData[245]));
Q_FDP0UA U1031 ( .D(n6090), .QTFCLK( ), .Q(ofifoData[246]));
Q_FDP0UA U1032 ( .D(n6091), .QTFCLK( ), .Q(ofifoData[247]));
Q_FDP0UA U1033 ( .D(n6092), .QTFCLK( ), .Q(ofifoData[248]));
Q_FDP0UA U1034 ( .D(n6093), .QTFCLK( ), .Q(ofifoData[249]));
Q_FDP0UA U1035 ( .D(n6094), .QTFCLK( ), .Q(ofifoData[250]));
Q_FDP0UA U1036 ( .D(n6095), .QTFCLK( ), .Q(ofifoData[251]));
Q_FDP0UA U1037 ( .D(n6096), .QTFCLK( ), .Q(ofifoData[252]));
Q_FDP0UA U1038 ( .D(n6097), .QTFCLK( ), .Q(ofifoData[253]));
Q_FDP0UA U1039 ( .D(n6098), .QTFCLK( ), .Q(ofifoData[254]));
Q_FDP0UA U1040 ( .D(n6099), .QTFCLK( ), .Q(ofifoData[255]));
Q_FDP0UA U1041 ( .D(n6100), .QTFCLK( ), .Q(ofifoData[256]));
Q_FDP0UA U1042 ( .D(n6101), .QTFCLK( ), .Q(ofifoData[257]));
Q_FDP0UA U1043 ( .D(n6102), .QTFCLK( ), .Q(ofifoData[258]));
Q_FDP0UA U1044 ( .D(n6103), .QTFCLK( ), .Q(ofifoData[259]));
Q_FDP0UA U1045 ( .D(n6104), .QTFCLK( ), .Q(ofifoData[260]));
Q_FDP0UA U1046 ( .D(n6105), .QTFCLK( ), .Q(ofifoData[261]));
Q_FDP0UA U1047 ( .D(n6106), .QTFCLK( ), .Q(ofifoData[262]));
Q_FDP0UA U1048 ( .D(n6107), .QTFCLK( ), .Q(ofifoData[263]));
Q_FDP0UA U1049 ( .D(n6108), .QTFCLK( ), .Q(ofifoData[264]));
Q_FDP0UA U1050 ( .D(n6109), .QTFCLK( ), .Q(ofifoData[265]));
Q_FDP0UA U1051 ( .D(n6110), .QTFCLK( ), .Q(ofifoData[266]));
Q_FDP0UA U1052 ( .D(n6111), .QTFCLK( ), .Q(ofifoData[267]));
Q_FDP0UA U1053 ( .D(n6112), .QTFCLK( ), .Q(ofifoData[268]));
Q_FDP0UA U1054 ( .D(n6113), .QTFCLK( ), .Q(ofifoData[269]));
Q_FDP0UA U1055 ( .D(n6114), .QTFCLK( ), .Q(ofifoData[270]));
Q_FDP0UA U1056 ( .D(n6115), .QTFCLK( ), .Q(ofifoData[271]));
Q_FDP0UA U1057 ( .D(n6116), .QTFCLK( ), .Q(ofifoData[272]));
Q_FDP0UA U1058 ( .D(n6117), .QTFCLK( ), .Q(ofifoData[273]));
Q_FDP0UA U1059 ( .D(n6118), .QTFCLK( ), .Q(ofifoData[274]));
Q_FDP0UA U1060 ( .D(n6119), .QTFCLK( ), .Q(ofifoData[275]));
Q_FDP0UA U1061 ( .D(n6120), .QTFCLK( ), .Q(ofifoData[276]));
Q_FDP0UA U1062 ( .D(n6121), .QTFCLK( ), .Q(ofifoData[277]));
Q_FDP0UA U1063 ( .D(n6122), .QTFCLK( ), .Q(ofifoData[278]));
Q_FDP0UA U1064 ( .D(n6123), .QTFCLK( ), .Q(ofifoData[279]));
Q_FDP0UA U1065 ( .D(n6124), .QTFCLK( ), .Q(ofifoData[280]));
Q_FDP0UA U1066 ( .D(n6125), .QTFCLK( ), .Q(ofifoData[281]));
Q_FDP0UA U1067 ( .D(n6126), .QTFCLK( ), .Q(ofifoData[282]));
Q_FDP0UA U1068 ( .D(n6127), .QTFCLK( ), .Q(ofifoData[283]));
Q_FDP0UA U1069 ( .D(n6128), .QTFCLK( ), .Q(ofifoData[284]));
Q_FDP0UA U1070 ( .D(n6129), .QTFCLK( ), .Q(ofifoData[285]));
Q_FDP0UA U1071 ( .D(n6130), .QTFCLK( ), .Q(ofifoData[286]));
Q_FDP0UA U1072 ( .D(n6131), .QTFCLK( ), .Q(ofifoData[287]));
Q_FDP0UA U1073 ( .D(n6132), .QTFCLK( ), .Q(ofifoData[288]));
Q_FDP0UA U1074 ( .D(n6133), .QTFCLK( ), .Q(ofifoData[289]));
Q_FDP0UA U1075 ( .D(n6134), .QTFCLK( ), .Q(ofifoData[290]));
Q_FDP0UA U1076 ( .D(n6135), .QTFCLK( ), .Q(ofifoData[291]));
Q_FDP0UA U1077 ( .D(n6136), .QTFCLK( ), .Q(ofifoData[292]));
Q_FDP0UA U1078 ( .D(n6137), .QTFCLK( ), .Q(ofifoData[293]));
Q_FDP0UA U1079 ( .D(n6138), .QTFCLK( ), .Q(ofifoData[294]));
Q_FDP0UA U1080 ( .D(n6139), .QTFCLK( ), .Q(ofifoData[295]));
Q_FDP0UA U1081 ( .D(n6140), .QTFCLK( ), .Q(ofifoData[296]));
Q_FDP0UA U1082 ( .D(n6141), .QTFCLK( ), .Q(ofifoData[297]));
Q_FDP0UA U1083 ( .D(n6142), .QTFCLK( ), .Q(ofifoData[298]));
Q_FDP0UA U1084 ( .D(n6143), .QTFCLK( ), .Q(ofifoData[299]));
Q_FDP0UA U1085 ( .D(n6144), .QTFCLK( ), .Q(ofifoData[300]));
Q_FDP0UA U1086 ( .D(n6145), .QTFCLK( ), .Q(ofifoData[301]));
Q_FDP0UA U1087 ( .D(n6146), .QTFCLK( ), .Q(ofifoData[302]));
Q_FDP0UA U1088 ( .D(n6147), .QTFCLK( ), .Q(ofifoData[303]));
Q_FDP0UA U1089 ( .D(n6148), .QTFCLK( ), .Q(ofifoData[304]));
Q_FDP0UA U1090 ( .D(n6149), .QTFCLK( ), .Q(ofifoData[305]));
Q_FDP0UA U1091 ( .D(n6150), .QTFCLK( ), .Q(ofifoData[306]));
Q_FDP0UA U1092 ( .D(n6151), .QTFCLK( ), .Q(ofifoData[307]));
Q_FDP0UA U1093 ( .D(n6152), .QTFCLK( ), .Q(ofifoData[308]));
Q_FDP0UA U1094 ( .D(n6153), .QTFCLK( ), .Q(ofifoData[309]));
Q_FDP0UA U1095 ( .D(n6154), .QTFCLK( ), .Q(ofifoData[310]));
Q_FDP0UA U1096 ( .D(n6155), .QTFCLK( ), .Q(ofifoData[311]));
Q_FDP0UA U1097 ( .D(n6156), .QTFCLK( ), .Q(ofifoData[312]));
Q_FDP0UA U1098 ( .D(n6157), .QTFCLK( ), .Q(ofifoData[313]));
Q_FDP0UA U1099 ( .D(n6158), .QTFCLK( ), .Q(ofifoData[314]));
Q_FDP0UA U1100 ( .D(n6159), .QTFCLK( ), .Q(ofifoData[315]));
Q_FDP0UA U1101 ( .D(n6160), .QTFCLK( ), .Q(ofifoData[316]));
Q_FDP0UA U1102 ( .D(n6161), .QTFCLK( ), .Q(ofifoData[317]));
Q_FDP0UA U1103 ( .D(n6162), .QTFCLK( ), .Q(ofifoData[318]));
Q_FDP0UA U1104 ( .D(n6163), .QTFCLK( ), .Q(ofifoData[319]));
Q_FDP0UA U1105 ( .D(n6164), .QTFCLK( ), .Q(ofifoData[320]));
Q_FDP0UA U1106 ( .D(n6165), .QTFCLK( ), .Q(ofifoData[321]));
Q_FDP0UA U1107 ( .D(n6166), .QTFCLK( ), .Q(ofifoData[322]));
Q_FDP0UA U1108 ( .D(n6167), .QTFCLK( ), .Q(ofifoData[323]));
Q_FDP0UA U1109 ( .D(n6168), .QTFCLK( ), .Q(ofifoData[324]));
Q_FDP0UA U1110 ( .D(n6169), .QTFCLK( ), .Q(ofifoData[325]));
Q_FDP0UA U1111 ( .D(n6170), .QTFCLK( ), .Q(ofifoData[326]));
Q_FDP0UA U1112 ( .D(n6171), .QTFCLK( ), .Q(ofifoData[327]));
Q_FDP0UA U1113 ( .D(n6172), .QTFCLK( ), .Q(ofifoData[328]));
Q_FDP0UA U1114 ( .D(n6173), .QTFCLK( ), .Q(ofifoData[329]));
Q_FDP0UA U1115 ( .D(n6174), .QTFCLK( ), .Q(ofifoData[330]));
Q_FDP0UA U1116 ( .D(n6175), .QTFCLK( ), .Q(ofifoData[331]));
Q_FDP0UA U1117 ( .D(n6176), .QTFCLK( ), .Q(ofifoData[332]));
Q_FDP0UA U1118 ( .D(n6177), .QTFCLK( ), .Q(ofifoData[333]));
Q_FDP0UA U1119 ( .D(n6178), .QTFCLK( ), .Q(ofifoData[334]));
Q_FDP0UA U1120 ( .D(n6179), .QTFCLK( ), .Q(ofifoData[335]));
Q_FDP0UA U1121 ( .D(n6180), .QTFCLK( ), .Q(ofifoData[336]));
Q_FDP0UA U1122 ( .D(n6181), .QTFCLK( ), .Q(ofifoData[337]));
Q_FDP0UA U1123 ( .D(n6182), .QTFCLK( ), .Q(ofifoData[338]));
Q_FDP0UA U1124 ( .D(n6183), .QTFCLK( ), .Q(ofifoData[339]));
Q_FDP0UA U1125 ( .D(n6184), .QTFCLK( ), .Q(ofifoData[340]));
Q_FDP0UA U1126 ( .D(n6185), .QTFCLK( ), .Q(ofifoData[341]));
Q_FDP0UA U1127 ( .D(n6186), .QTFCLK( ), .Q(ofifoData[342]));
Q_FDP0UA U1128 ( .D(n6187), .QTFCLK( ), .Q(ofifoData[343]));
Q_FDP0UA U1129 ( .D(n6188), .QTFCLK( ), .Q(ofifoData[344]));
Q_FDP0UA U1130 ( .D(n6189), .QTFCLK( ), .Q(ofifoData[345]));
Q_FDP0UA U1131 ( .D(n6190), .QTFCLK( ), .Q(ofifoData[346]));
Q_FDP0UA U1132 ( .D(n6191), .QTFCLK( ), .Q(ofifoData[347]));
Q_FDP0UA U1133 ( .D(n6192), .QTFCLK( ), .Q(ofifoData[348]));
Q_FDP0UA U1134 ( .D(n6193), .QTFCLK( ), .Q(ofifoData[349]));
Q_FDP0UA U1135 ( .D(n6194), .QTFCLK( ), .Q(ofifoData[350]));
Q_FDP0UA U1136 ( .D(n6195), .QTFCLK( ), .Q(ofifoData[351]));
Q_FDP0UA U1137 ( .D(n6196), .QTFCLK( ), .Q(ofifoData[352]));
Q_FDP0UA U1138 ( .D(n6197), .QTFCLK( ), .Q(ofifoData[353]));
Q_FDP0UA U1139 ( .D(n6198), .QTFCLK( ), .Q(ofifoData[354]));
Q_FDP0UA U1140 ( .D(n6199), .QTFCLK( ), .Q(ofifoData[355]));
Q_FDP0UA U1141 ( .D(n6200), .QTFCLK( ), .Q(ofifoData[356]));
Q_FDP0UA U1142 ( .D(n6201), .QTFCLK( ), .Q(ofifoData[357]));
Q_FDP0UA U1143 ( .D(n6202), .QTFCLK( ), .Q(ofifoData[358]));
Q_FDP0UA U1144 ( .D(n6203), .QTFCLK( ), .Q(ofifoData[359]));
Q_FDP0UA U1145 ( .D(n6204), .QTFCLK( ), .Q(ofifoData[360]));
Q_FDP0UA U1146 ( .D(n6205), .QTFCLK( ), .Q(ofifoData[361]));
Q_FDP0UA U1147 ( .D(n6206), .QTFCLK( ), .Q(ofifoData[362]));
Q_FDP0UA U1148 ( .D(n6207), .QTFCLK( ), .Q(ofifoData[363]));
Q_FDP0UA U1149 ( .D(n6208), .QTFCLK( ), .Q(ofifoData[364]));
Q_FDP0UA U1150 ( .D(n6209), .QTFCLK( ), .Q(ofifoData[365]));
Q_FDP0UA U1151 ( .D(n6210), .QTFCLK( ), .Q(ofifoData[366]));
Q_FDP0UA U1152 ( .D(n6211), .QTFCLK( ), .Q(ofifoData[367]));
Q_FDP0UA U1153 ( .D(n6212), .QTFCLK( ), .Q(ofifoData[368]));
Q_FDP0UA U1154 ( .D(n6213), .QTFCLK( ), .Q(ofifoData[369]));
Q_FDP0UA U1155 ( .D(n6214), .QTFCLK( ), .Q(ofifoData[370]));
Q_FDP0UA U1156 ( .D(n6215), .QTFCLK( ), .Q(ofifoData[371]));
Q_FDP0UA U1157 ( .D(n6216), .QTFCLK( ), .Q(ofifoData[372]));
Q_FDP0UA U1158 ( .D(n6217), .QTFCLK( ), .Q(ofifoData[373]));
Q_FDP0UA U1159 ( .D(n6218), .QTFCLK( ), .Q(ofifoData[374]));
Q_FDP0UA U1160 ( .D(n6219), .QTFCLK( ), .Q(ofifoData[375]));
Q_FDP0UA U1161 ( .D(n6220), .QTFCLK( ), .Q(ofifoData[376]));
Q_FDP0UA U1162 ( .D(n6221), .QTFCLK( ), .Q(ofifoData[377]));
Q_FDP0UA U1163 ( .D(n6222), .QTFCLK( ), .Q(ofifoData[378]));
Q_FDP0UA U1164 ( .D(n6223), .QTFCLK( ), .Q(ofifoData[379]));
Q_FDP0UA U1165 ( .D(n6224), .QTFCLK( ), .Q(ofifoData[380]));
Q_FDP0UA U1166 ( .D(n6225), .QTFCLK( ), .Q(ofifoData[381]));
Q_FDP0UA U1167 ( .D(n6226), .QTFCLK( ), .Q(ofifoData[382]));
Q_FDP0UA U1168 ( .D(n6227), .QTFCLK( ), .Q(ofifoData[383]));
Q_FDP0UA U1169 ( .D(n6228), .QTFCLK( ), .Q(ofifoData[384]));
Q_FDP0UA U1170 ( .D(n6229), .QTFCLK( ), .Q(ofifoData[385]));
Q_FDP0UA U1171 ( .D(n6230), .QTFCLK( ), .Q(ofifoData[386]));
Q_FDP0UA U1172 ( .D(n6231), .QTFCLK( ), .Q(ofifoData[387]));
Q_FDP0UA U1173 ( .D(n6232), .QTFCLK( ), .Q(ofifoData[388]));
Q_FDP0UA U1174 ( .D(n6233), .QTFCLK( ), .Q(ofifoData[389]));
Q_FDP0UA U1175 ( .D(n6234), .QTFCLK( ), .Q(ofifoData[390]));
Q_FDP0UA U1176 ( .D(n6235), .QTFCLK( ), .Q(ofifoData[391]));
Q_FDP0UA U1177 ( .D(n6236), .QTFCLK( ), .Q(ofifoData[392]));
Q_FDP0UA U1178 ( .D(n6237), .QTFCLK( ), .Q(ofifoData[393]));
Q_FDP0UA U1179 ( .D(n6238), .QTFCLK( ), .Q(ofifoData[394]));
Q_FDP0UA U1180 ( .D(n6239), .QTFCLK( ), .Q(ofifoData[395]));
Q_FDP0UA U1181 ( .D(n6240), .QTFCLK( ), .Q(ofifoData[396]));
Q_FDP0UA U1182 ( .D(n6241), .QTFCLK( ), .Q(ofifoData[397]));
Q_FDP0UA U1183 ( .D(n6242), .QTFCLK( ), .Q(ofifoData[398]));
Q_FDP0UA U1184 ( .D(n6243), .QTFCLK( ), .Q(ofifoData[399]));
Q_FDP0UA U1185 ( .D(n6244), .QTFCLK( ), .Q(ofifoData[400]));
Q_FDP0UA U1186 ( .D(n6245), .QTFCLK( ), .Q(ofifoData[401]));
Q_FDP0UA U1187 ( .D(n6246), .QTFCLK( ), .Q(ofifoData[402]));
Q_FDP0UA U1188 ( .D(n6247), .QTFCLK( ), .Q(ofifoData[403]));
Q_FDP0UA U1189 ( .D(n6248), .QTFCLK( ), .Q(ofifoData[404]));
Q_FDP0UA U1190 ( .D(n6249), .QTFCLK( ), .Q(ofifoData[405]));
Q_FDP0UA U1191 ( .D(n6250), .QTFCLK( ), .Q(ofifoData[406]));
Q_FDP0UA U1192 ( .D(n6251), .QTFCLK( ), .Q(ofifoData[407]));
Q_FDP0UA U1193 ( .D(n6252), .QTFCLK( ), .Q(ofifoData[408]));
Q_FDP0UA U1194 ( .D(n6253), .QTFCLK( ), .Q(ofifoData[409]));
Q_FDP0UA U1195 ( .D(n6254), .QTFCLK( ), .Q(ofifoData[410]));
Q_FDP0UA U1196 ( .D(n6255), .QTFCLK( ), .Q(ofifoData[411]));
Q_FDP0UA U1197 ( .D(n6256), .QTFCLK( ), .Q(ofifoData[412]));
Q_FDP0UA U1198 ( .D(n6257), .QTFCLK( ), .Q(ofifoData[413]));
Q_FDP0UA U1199 ( .D(n6258), .QTFCLK( ), .Q(ofifoData[414]));
Q_FDP0UA U1200 ( .D(n6259), .QTFCLK( ), .Q(ofifoData[415]));
Q_FDP0UA U1201 ( .D(n6260), .QTFCLK( ), .Q(ofifoData[416]));
Q_FDP0UA U1202 ( .D(n6261), .QTFCLK( ), .Q(ofifoData[417]));
Q_FDP0UA U1203 ( .D(n6262), .QTFCLK( ), .Q(ofifoData[418]));
Q_FDP0UA U1204 ( .D(n6263), .QTFCLK( ), .Q(ofifoData[419]));
Q_FDP0UA U1205 ( .D(n6264), .QTFCLK( ), .Q(ofifoData[420]));
Q_FDP0UA U1206 ( .D(n6265), .QTFCLK( ), .Q(ofifoData[421]));
Q_FDP0UA U1207 ( .D(n6266), .QTFCLK( ), .Q(ofifoData[422]));
Q_FDP0UA U1208 ( .D(n6267), .QTFCLK( ), .Q(ofifoData[423]));
Q_FDP0UA U1209 ( .D(n6268), .QTFCLK( ), .Q(ofifoData[424]));
Q_FDP0UA U1210 ( .D(n6269), .QTFCLK( ), .Q(ofifoData[425]));
Q_FDP0UA U1211 ( .D(n6270), .QTFCLK( ), .Q(ofifoData[426]));
Q_FDP0UA U1212 ( .D(n6271), .QTFCLK( ), .Q(ofifoData[427]));
Q_FDP0UA U1213 ( .D(n6272), .QTFCLK( ), .Q(ofifoData[428]));
Q_FDP0UA U1214 ( .D(n6273), .QTFCLK( ), .Q(ofifoData[429]));
Q_FDP0UA U1215 ( .D(n6274), .QTFCLK( ), .Q(ofifoData[430]));
Q_FDP0UA U1216 ( .D(n6275), .QTFCLK( ), .Q(ofifoData[431]));
Q_FDP0UA U1217 ( .D(n6276), .QTFCLK( ), .Q(ofifoData[432]));
Q_FDP0UA U1218 ( .D(n6277), .QTFCLK( ), .Q(ofifoData[433]));
Q_FDP0UA U1219 ( .D(n6278), .QTFCLK( ), .Q(ofifoData[434]));
Q_FDP0UA U1220 ( .D(n6279), .QTFCLK( ), .Q(ofifoData[435]));
Q_FDP0UA U1221 ( .D(n6280), .QTFCLK( ), .Q(ofifoData[436]));
Q_FDP0UA U1222 ( .D(n6281), .QTFCLK( ), .Q(ofifoData[437]));
Q_FDP0UA U1223 ( .D(n6282), .QTFCLK( ), .Q(ofifoData[438]));
Q_FDP0UA U1224 ( .D(n6283), .QTFCLK( ), .Q(ofifoData[439]));
Q_FDP0UA U1225 ( .D(n6284), .QTFCLK( ), .Q(ofifoData[440]));
Q_FDP0UA U1226 ( .D(n6285), .QTFCLK( ), .Q(ofifoData[441]));
Q_FDP0UA U1227 ( .D(n6286), .QTFCLK( ), .Q(ofifoData[442]));
Q_FDP0UA U1228 ( .D(n6287), .QTFCLK( ), .Q(ofifoData[443]));
Q_FDP0UA U1229 ( .D(n6288), .QTFCLK( ), .Q(ofifoData[444]));
Q_FDP0UA U1230 ( .D(n6289), .QTFCLK( ), .Q(ofifoData[445]));
Q_FDP0UA U1231 ( .D(n6290), .QTFCLK( ), .Q(ofifoData[446]));
Q_FDP0UA U1232 ( .D(n6291), .QTFCLK( ), .Q(ofifoData[447]));
Q_FDP0UA U1233 ( .D(n6292), .QTFCLK( ), .Q(ofifoData[448]));
Q_FDP0UA U1234 ( .D(n6293), .QTFCLK( ), .Q(ofifoData[449]));
Q_FDP0UA U1235 ( .D(n6294), .QTFCLK( ), .Q(ofifoData[450]));
Q_FDP0UA U1236 ( .D(n6295), .QTFCLK( ), .Q(ofifoData[451]));
Q_FDP0UA U1237 ( .D(n6296), .QTFCLK( ), .Q(ofifoData[452]));
Q_FDP0UA U1238 ( .D(n6297), .QTFCLK( ), .Q(ofifoData[453]));
Q_FDP0UA U1239 ( .D(n6298), .QTFCLK( ), .Q(ofifoData[454]));
Q_FDP0UA U1240 ( .D(n6299), .QTFCLK( ), .Q(ofifoData[455]));
Q_FDP0UA U1241 ( .D(n6300), .QTFCLK( ), .Q(ofifoData[456]));
Q_FDP0UA U1242 ( .D(n6301), .QTFCLK( ), .Q(ofifoData[457]));
Q_FDP0UA U1243 ( .D(n6302), .QTFCLK( ), .Q(ofifoData[458]));
Q_FDP0UA U1244 ( .D(n6303), .QTFCLK( ), .Q(ofifoData[459]));
Q_FDP0UA U1245 ( .D(n6304), .QTFCLK( ), .Q(ofifoData[460]));
Q_FDP0UA U1246 ( .D(n6305), .QTFCLK( ), .Q(ofifoData[461]));
Q_FDP0UA U1247 ( .D(n6306), .QTFCLK( ), .Q(ofifoData[462]));
Q_FDP0UA U1248 ( .D(n6307), .QTFCLK( ), .Q(ofifoData[463]));
Q_FDP0UA U1249 ( .D(n6308), .QTFCLK( ), .Q(ofifoData[464]));
Q_FDP0UA U1250 ( .D(n6309), .QTFCLK( ), .Q(ofifoData[465]));
Q_FDP0UA U1251 ( .D(n6310), .QTFCLK( ), .Q(ofifoData[466]));
Q_FDP0UA U1252 ( .D(n6311), .QTFCLK( ), .Q(ofifoData[467]));
Q_FDP0UA U1253 ( .D(n6312), .QTFCLK( ), .Q(ofifoData[468]));
Q_FDP0UA U1254 ( .D(n6313), .QTFCLK( ), .Q(ofifoData[469]));
Q_FDP0UA U1255 ( .D(n6314), .QTFCLK( ), .Q(ofifoData[470]));
Q_FDP0UA U1256 ( .D(n6315), .QTFCLK( ), .Q(ofifoData[471]));
Q_FDP0UA U1257 ( .D(n6316), .QTFCLK( ), .Q(ofifoData[472]));
Q_FDP0UA U1258 ( .D(n6317), .QTFCLK( ), .Q(ofifoData[473]));
Q_FDP0UA U1259 ( .D(n6318), .QTFCLK( ), .Q(ofifoData[474]));
Q_FDP0UA U1260 ( .D(n6319), .QTFCLK( ), .Q(ofifoData[475]));
Q_FDP0UA U1261 ( .D(n6320), .QTFCLK( ), .Q(ofifoData[476]));
Q_FDP0UA U1262 ( .D(n6321), .QTFCLK( ), .Q(ofifoData[477]));
Q_FDP0UA U1263 ( .D(n6322), .QTFCLK( ), .Q(ofifoData[478]));
Q_FDP0UA U1264 ( .D(n6323), .QTFCLK( ), .Q(ofifoData[479]));
Q_FDP0UA U1265 ( .D(n6324), .QTFCLK( ), .Q(ofifoData[480]));
Q_FDP0UA U1266 ( .D(n6325), .QTFCLK( ), .Q(ofifoData[481]));
Q_FDP0UA U1267 ( .D(n6326), .QTFCLK( ), .Q(ofifoData[482]));
Q_FDP0UA U1268 ( .D(n6327), .QTFCLK( ), .Q(ofifoData[483]));
Q_FDP0UA U1269 ( .D(n6328), .QTFCLK( ), .Q(ofifoData[484]));
Q_FDP0UA U1270 ( .D(n6329), .QTFCLK( ), .Q(ofifoData[485]));
Q_FDP0UA U1271 ( .D(n6330), .QTFCLK( ), .Q(ofifoData[486]));
Q_FDP0UA U1272 ( .D(n6331), .QTFCLK( ), .Q(ofifoData[487]));
Q_FDP0UA U1273 ( .D(n6332), .QTFCLK( ), .Q(ofifoData[488]));
Q_FDP0UA U1274 ( .D(n6333), .QTFCLK( ), .Q(ofifoData[489]));
Q_FDP0UA U1275 ( .D(n6334), .QTFCLK( ), .Q(ofifoData[490]));
Q_FDP0UA U1276 ( .D(n6335), .QTFCLK( ), .Q(ofifoData[491]));
Q_FDP0UA U1277 ( .D(n6336), .QTFCLK( ), .Q(ofifoData[492]));
Q_FDP0UA U1278 ( .D(n6337), .QTFCLK( ), .Q(ofifoData[493]));
Q_FDP0UA U1279 ( .D(n6338), .QTFCLK( ), .Q(ofifoData[494]));
Q_FDP0UA U1280 ( .D(n6339), .QTFCLK( ), .Q(ofifoData[495]));
Q_FDP0UA U1281 ( .D(n6340), .QTFCLK( ), .Q(ofifoData[496]));
Q_FDP0UA U1282 ( .D(n6341), .QTFCLK( ), .Q(ofifoData[497]));
Q_FDP0UA U1283 ( .D(n6342), .QTFCLK( ), .Q(ofifoData[498]));
Q_FDP0UA U1284 ( .D(n6343), .QTFCLK( ), .Q(ofifoData[499]));
Q_FDP0UA U1285 ( .D(n6344), .QTFCLK( ), .Q(ofifoData[500]));
Q_FDP0UA U1286 ( .D(n6345), .QTFCLK( ), .Q(ofifoData[501]));
Q_FDP0UA U1287 ( .D(n6346), .QTFCLK( ), .Q(ofifoData[502]));
Q_FDP0UA U1288 ( .D(n6347), .QTFCLK( ), .Q(ofifoData[503]));
Q_FDP0UA U1289 ( .D(n6348), .QTFCLK( ), .Q(ofifoData[504]));
Q_FDP0UA U1290 ( .D(n6349), .QTFCLK( ), .Q(ofifoData[505]));
Q_FDP0UA U1291 ( .D(n6350), .QTFCLK( ), .Q(ofifoData[506]));
Q_FDP0UA U1292 ( .D(n6351), .QTFCLK( ), .Q(ofifoData[507]));
Q_FDP0UA U1293 ( .D(n6352), .QTFCLK( ), .Q(ofifoData[508]));
Q_FDP0UA U1294 ( .D(n6353), .QTFCLK( ), .Q(ofifoData[509]));
Q_FDP0UA U1295 ( .D(n6354), .QTFCLK( ), .Q(ofifoData[510]));
Q_FDP0UA U1296 ( .D(n6355), .QTFCLK( ), .Q(ofifoData[511]));
Q_FDP0UA U1297 ( .D(n6356), .QTFCLK( ), .Q(ofifoData[512]));
Q_FDP0UA U1298 ( .D(n6357), .QTFCLK( ), .Q(ofifoData[513]));
Q_FDP0UA U1299 ( .D(n6358), .QTFCLK( ), .Q(ofifoData[514]));
Q_FDP0UA U1300 ( .D(n6359), .QTFCLK( ), .Q(ofifoData[515]));
Q_FDP0UA U1301 ( .D(n6360), .QTFCLK( ), .Q(ofifoData[516]));
Q_FDP0UA U1302 ( .D(n6361), .QTFCLK( ), .Q(ofifoData[517]));
Q_FDP0UA U1303 ( .D(n6362), .QTFCLK( ), .Q(ofifoData[518]));
Q_FDP0UA U1304 ( .D(n6363), .QTFCLK( ), .Q(ofifoData[519]));
Q_FDP0UA U1305 ( .D(n6364), .QTFCLK( ), .Q(ofifoData[520]));
Q_FDP0UA U1306 ( .D(n6365), .QTFCLK( ), .Q(ofifoData[521]));
Q_FDP0UA U1307 ( .D(n6366), .QTFCLK( ), .Q(ofifoData[522]));
Q_FDP0UA U1308 ( .D(n6367), .QTFCLK( ), .Q(ofifoData[523]));
Q_FDP0UA U1309 ( .D(n6368), .QTFCLK( ), .Q(ofifoData[524]));
Q_FDP0UA U1310 ( .D(n6369), .QTFCLK( ), .Q(ofifoData[525]));
Q_FDP0UA U1311 ( .D(n6370), .QTFCLK( ), .Q(ofifoData[526]));
Q_FDP0UA U1312 ( .D(n6371), .QTFCLK( ), .Q(ofifoData[527]));
Q_FDP0UA U1313 ( .D(n6372), .QTFCLK( ), .Q(ofifoData[528]));
Q_FDP0UA U1314 ( .D(n6373), .QTFCLK( ), .Q(ofifoData[529]));
Q_FDP0UA U1315 ( .D(n6374), .QTFCLK( ), .Q(ofifoData[530]));
Q_FDP0UA U1316 ( .D(n6375), .QTFCLK( ), .Q(ofifoData[531]));
Q_FDP0UA U1317 ( .D(n6376), .QTFCLK( ), .Q(ofifoData[532]));
Q_FDP0UA U1318 ( .D(n6377), .QTFCLK( ), .Q(ofifoData[533]));
Q_FDP0UA U1319 ( .D(n6378), .QTFCLK( ), .Q(ofifoData[534]));
Q_FDP0UA U1320 ( .D(n6379), .QTFCLK( ), .Q(ofifoData[535]));
Q_FDP0UA U1321 ( .D(n6380), .QTFCLK( ), .Q(ofifoData[536]));
Q_FDP0UA U1322 ( .D(n6381), .QTFCLK( ), .Q(ofifoData[537]));
Q_FDP0UA U1323 ( .D(n6382), .QTFCLK( ), .Q(ofifoData[538]));
Q_FDP0UA U1324 ( .D(n6383), .QTFCLK( ), .Q(ofifoData[539]));
Q_FDP0UA U1325 ( .D(n6384), .QTFCLK( ), .Q(ofifoData[540]));
Q_FDP0UA U1326 ( .D(n6385), .QTFCLK( ), .Q(ofifoData[541]));
Q_FDP0UA U1327 ( .D(n6386), .QTFCLK( ), .Q(ofifoData[542]));
Q_FDP0UA U1328 ( .D(n6387), .QTFCLK( ), .Q(ofifoData[543]));
Q_FDP0UA U1329 ( .D(n6388), .QTFCLK( ), .Q(ofifoData[544]));
Q_FDP0UA U1330 ( .D(n6389), .QTFCLK( ), .Q(ofifoData[545]));
Q_FDP0UA U1331 ( .D(n6390), .QTFCLK( ), .Q(ofifoData[546]));
Q_FDP0UA U1332 ( .D(n6391), .QTFCLK( ), .Q(ofifoData[547]));
Q_FDP0UA U1333 ( .D(n6392), .QTFCLK( ), .Q(ofifoData[548]));
Q_FDP0UA U1334 ( .D(n6393), .QTFCLK( ), .Q(ofifoData[549]));
Q_FDP0UA U1335 ( .D(n6394), .QTFCLK( ), .Q(ofifoData[550]));
Q_FDP0UA U1336 ( .D(n6395), .QTFCLK( ), .Q(ofifoData[551]));
Q_FDP0UA U1337 ( .D(n6396), .QTFCLK( ), .Q(ofifoData[552]));
Q_FDP0UA U1338 ( .D(n6397), .QTFCLK( ), .Q(ofifoData[553]));
Q_FDP0UA U1339 ( .D(n6398), .QTFCLK( ), .Q(ofifoData[554]));
Q_FDP0UA U1340 ( .D(n6399), .QTFCLK( ), .Q(ofifoData[555]));
Q_FDP0UA U1341 ( .D(n6400), .QTFCLK( ), .Q(ofifoData[556]));
Q_FDP0UA U1342 ( .D(n6401), .QTFCLK( ), .Q(ofifoData[557]));
Q_FDP0UA U1343 ( .D(n6402), .QTFCLK( ), .Q(ofifoData[558]));
Q_FDP0UA U1344 ( .D(n6403), .QTFCLK( ), .Q(ofifoData[559]));
Q_FDP0UA U1345 ( .D(n6404), .QTFCLK( ), .Q(ofifoData[560]));
Q_FDP0UA U1346 ( .D(n6405), .QTFCLK( ), .Q(ofifoData[561]));
Q_FDP0UA U1347 ( .D(n6406), .QTFCLK( ), .Q(ofifoData[562]));
Q_FDP0UA U1348 ( .D(n6407), .QTFCLK( ), .Q(ofifoData[563]));
Q_FDP0UA U1349 ( .D(n6408), .QTFCLK( ), .Q(ofifoData[564]));
Q_FDP0UA U1350 ( .D(n6409), .QTFCLK( ), .Q(ofifoData[565]));
Q_FDP0UA U1351 ( .D(n6410), .QTFCLK( ), .Q(ofifoData[566]));
Q_FDP0UA U1352 ( .D(n6411), .QTFCLK( ), .Q(ofifoData[567]));
Q_FDP0UA U1353 ( .D(n6412), .QTFCLK( ), .Q(ofifoData[568]));
Q_FDP0UA U1354 ( .D(n6413), .QTFCLK( ), .Q(ofifoData[569]));
Q_FDP0UA U1355 ( .D(n6414), .QTFCLK( ), .Q(ofifoData[570]));
Q_FDP0UA U1356 ( .D(n6415), .QTFCLK( ), .Q(ofifoData[571]));
Q_FDP0UA U1357 ( .D(n6416), .QTFCLK( ), .Q(ofifoData[572]));
Q_FDP0UA U1358 ( .D(n6417), .QTFCLK( ), .Q(ofifoData[573]));
Q_FDP0UA U1359 ( .D(n6418), .QTFCLK( ), .Q(ofifoData[574]));
Q_FDP0UA U1360 ( .D(n6419), .QTFCLK( ), .Q(ofifoData[575]));
Q_FDP0UA U1361 ( .D(n6420), .QTFCLK( ), .Q(ofifoData[576]));
Q_FDP0UA U1362 ( .D(n6421), .QTFCLK( ), .Q(ofifoData[577]));
Q_FDP0UA U1363 ( .D(n6422), .QTFCLK( ), .Q(ofifoData[578]));
Q_FDP0UA U1364 ( .D(n6423), .QTFCLK( ), .Q(ofifoData[579]));
Q_FDP0UA U1365 ( .D(n6424), .QTFCLK( ), .Q(ofifoData[580]));
Q_FDP0UA U1366 ( .D(n6425), .QTFCLK( ), .Q(ofifoData[581]));
Q_FDP0UA U1367 ( .D(n6426), .QTFCLK( ), .Q(ofifoData[582]));
Q_FDP0UA U1368 ( .D(n6427), .QTFCLK( ), .Q(ofifoData[583]));
Q_FDP0UA U1369 ( .D(n6428), .QTFCLK( ), .Q(ofifoData[584]));
Q_FDP0UA U1370 ( .D(n6429), .QTFCLK( ), .Q(ofifoData[585]));
Q_FDP0UA U1371 ( .D(n6430), .QTFCLK( ), .Q(ofifoData[586]));
Q_FDP0UA U1372 ( .D(n6431), .QTFCLK( ), .Q(ofifoData[587]));
Q_FDP0UA U1373 ( .D(n6432), .QTFCLK( ), .Q(ofifoData[588]));
Q_FDP0UA U1374 ( .D(n6433), .QTFCLK( ), .Q(ofifoData[589]));
Q_FDP0UA U1375 ( .D(n6434), .QTFCLK( ), .Q(ofifoData[590]));
Q_FDP0UA U1376 ( .D(n6435), .QTFCLK( ), .Q(ofifoData[591]));
Q_FDP0UA U1377 ( .D(n6436), .QTFCLK( ), .Q(ofifoData[592]));
Q_FDP0UA U1378 ( .D(n6437), .QTFCLK( ), .Q(ofifoData[593]));
Q_FDP0UA U1379 ( .D(n6438), .QTFCLK( ), .Q(ofifoData[594]));
Q_FDP0UA U1380 ( .D(n6439), .QTFCLK( ), .Q(ofifoData[595]));
Q_FDP0UA U1381 ( .D(n6440), .QTFCLK( ), .Q(ofifoData[596]));
Q_FDP0UA U1382 ( .D(n6441), .QTFCLK( ), .Q(ofifoData[597]));
Q_FDP0UA U1383 ( .D(n6442), .QTFCLK( ), .Q(ofifoData[598]));
Q_FDP0UA U1384 ( .D(n6443), .QTFCLK( ), .Q(ofifoData[599]));
Q_FDP0UA U1385 ( .D(n6444), .QTFCLK( ), .Q(ofifoData[600]));
Q_FDP0UA U1386 ( .D(n6445), .QTFCLK( ), .Q(ofifoData[601]));
Q_FDP0UA U1387 ( .D(n6446), .QTFCLK( ), .Q(ofifoData[602]));
Q_FDP0UA U1388 ( .D(n6447), .QTFCLK( ), .Q(ofifoData[603]));
Q_FDP0UA U1389 ( .D(n6448), .QTFCLK( ), .Q(ofifoData[604]));
Q_FDP0UA U1390 ( .D(n6449), .QTFCLK( ), .Q(ofifoData[605]));
Q_FDP0UA U1391 ( .D(n6450), .QTFCLK( ), .Q(ofifoData[606]));
Q_FDP0UA U1392 ( .D(n6451), .QTFCLK( ), .Q(ofifoData[607]));
Q_FDP0UA U1393 ( .D(n6452), .QTFCLK( ), .Q(ofifoData[608]));
Q_FDP0UA U1394 ( .D(n6453), .QTFCLK( ), .Q(ofifoData[609]));
Q_FDP0UA U1395 ( .D(n6454), .QTFCLK( ), .Q(ofifoData[610]));
Q_FDP0UA U1396 ( .D(n6455), .QTFCLK( ), .Q(ofifoData[611]));
Q_FDP0UA U1397 ( .D(n6456), .QTFCLK( ), .Q(ofifoData[612]));
Q_FDP0UA U1398 ( .D(n6457), .QTFCLK( ), .Q(ofifoData[613]));
Q_FDP0UA U1399 ( .D(n6458), .QTFCLK( ), .Q(ofifoData[614]));
Q_FDP0UA U1400 ( .D(n6459), .QTFCLK( ), .Q(ofifoData[615]));
Q_FDP0UA U1401 ( .D(n6460), .QTFCLK( ), .Q(ofifoData[616]));
Q_FDP0UA U1402 ( .D(n6461), .QTFCLK( ), .Q(ofifoData[617]));
Q_FDP0UA U1403 ( .D(n6462), .QTFCLK( ), .Q(ofifoData[618]));
Q_FDP0UA U1404 ( .D(n6463), .QTFCLK( ), .Q(ofifoData[619]));
Q_FDP0UA U1405 ( .D(n6464), .QTFCLK( ), .Q(ofifoData[620]));
Q_FDP0UA U1406 ( .D(n6465), .QTFCLK( ), .Q(ofifoData[621]));
Q_FDP0UA U1407 ( .D(n6466), .QTFCLK( ), .Q(ofifoData[622]));
Q_FDP0UA U1408 ( .D(n6467), .QTFCLK( ), .Q(ofifoData[623]));
Q_FDP0UA U1409 ( .D(n6468), .QTFCLK( ), .Q(ofifoData[624]));
Q_FDP0UA U1410 ( .D(n6469), .QTFCLK( ), .Q(ofifoData[625]));
Q_FDP0UA U1411 ( .D(n6470), .QTFCLK( ), .Q(ofifoData[626]));
Q_FDP0UA U1412 ( .D(n6471), .QTFCLK( ), .Q(ofifoData[627]));
Q_FDP0UA U1413 ( .D(n6472), .QTFCLK( ), .Q(ofifoData[628]));
Q_FDP0UA U1414 ( .D(n6473), .QTFCLK( ), .Q(ofifoData[629]));
Q_FDP0UA U1415 ( .D(n6474), .QTFCLK( ), .Q(ofifoData[630]));
Q_FDP0UA U1416 ( .D(n6475), .QTFCLK( ), .Q(ofifoData[631]));
Q_FDP0UA U1417 ( .D(n6476), .QTFCLK( ), .Q(ofifoData[632]));
Q_FDP0UA U1418 ( .D(n6477), .QTFCLK( ), .Q(ofifoData[633]));
Q_FDP0UA U1419 ( .D(n6478), .QTFCLK( ), .Q(ofifoData[634]));
Q_FDP0UA U1420 ( .D(n6479), .QTFCLK( ), .Q(ofifoData[635]));
Q_FDP0UA U1421 ( .D(n6480), .QTFCLK( ), .Q(ofifoData[636]));
Q_FDP0UA U1422 ( .D(n6481), .QTFCLK( ), .Q(ofifoData[637]));
Q_FDP0UA U1423 ( .D(n6482), .QTFCLK( ), .Q(ofifoData[638]));
Q_FDP0UA U1424 ( .D(n6483), .QTFCLK( ), .Q(ofifoData[639]));
Q_FDP0UA U1425 ( .D(n6484), .QTFCLK( ), .Q(ofifoData[640]));
Q_FDP0UA U1426 ( .D(n6485), .QTFCLK( ), .Q(ofifoData[641]));
Q_FDP0UA U1427 ( .D(n6486), .QTFCLK( ), .Q(ofifoData[642]));
Q_FDP0UA U1428 ( .D(n6487), .QTFCLK( ), .Q(ofifoData[643]));
Q_FDP0UA U1429 ( .D(n6488), .QTFCLK( ), .Q(ofifoData[644]));
Q_FDP0UA U1430 ( .D(n6489), .QTFCLK( ), .Q(ofifoData[645]));
Q_FDP0UA U1431 ( .D(n6490), .QTFCLK( ), .Q(ofifoData[646]));
Q_FDP0UA U1432 ( .D(n6491), .QTFCLK( ), .Q(ofifoData[647]));
Q_FDP0UA U1433 ( .D(n6492), .QTFCLK( ), .Q(ofifoData[648]));
Q_FDP0UA U1434 ( .D(n6493), .QTFCLK( ), .Q(ofifoData[649]));
Q_FDP0UA U1435 ( .D(n6494), .QTFCLK( ), .Q(ofifoData[650]));
Q_FDP0UA U1436 ( .D(n6495), .QTFCLK( ), .Q(ofifoData[651]));
Q_FDP0UA U1437 ( .D(n6496), .QTFCLK( ), .Q(ofifoData[652]));
Q_FDP0UA U1438 ( .D(n6497), .QTFCLK( ), .Q(ofifoData[653]));
Q_FDP0UA U1439 ( .D(n6498), .QTFCLK( ), .Q(ofifoData[654]));
Q_FDP0UA U1440 ( .D(n6499), .QTFCLK( ), .Q(ofifoData[655]));
Q_FDP0UA U1441 ( .D(n6500), .QTFCLK( ), .Q(ofifoData[656]));
Q_FDP0UA U1442 ( .D(n6501), .QTFCLK( ), .Q(ofifoData[657]));
Q_FDP0UA U1443 ( .D(n6502), .QTFCLK( ), .Q(ofifoData[658]));
Q_FDP0UA U1444 ( .D(n6503), .QTFCLK( ), .Q(ofifoData[659]));
Q_FDP0UA U1445 ( .D(n6504), .QTFCLK( ), .Q(ofifoData[660]));
Q_FDP0UA U1446 ( .D(n6505), .QTFCLK( ), .Q(ofifoData[661]));
Q_FDP0UA U1447 ( .D(n6506), .QTFCLK( ), .Q(ofifoData[662]));
Q_FDP0UA U1448 ( .D(n6507), .QTFCLK( ), .Q(ofifoData[663]));
Q_FDP0UA U1449 ( .D(n6508), .QTFCLK( ), .Q(ofifoData[664]));
Q_FDP0UA U1450 ( .D(n6509), .QTFCLK( ), .Q(ofifoData[665]));
Q_FDP0UA U1451 ( .D(n6510), .QTFCLK( ), .Q(ofifoData[666]));
Q_FDP0UA U1452 ( .D(n6511), .QTFCLK( ), .Q(ofifoData[667]));
Q_FDP0UA U1453 ( .D(n6512), .QTFCLK( ), .Q(ofifoData[668]));
Q_FDP0UA U1454 ( .D(n6513), .QTFCLK( ), .Q(ofifoData[669]));
Q_FDP0UA U1455 ( .D(n6514), .QTFCLK( ), .Q(ofifoData[670]));
Q_FDP0UA U1456 ( .D(n6515), .QTFCLK( ), .Q(ofifoData[671]));
Q_FDP0UA U1457 ( .D(n6516), .QTFCLK( ), .Q(ofifoData[672]));
Q_FDP0UA U1458 ( .D(n6517), .QTFCLK( ), .Q(ofifoData[673]));
Q_FDP0UA U1459 ( .D(n6518), .QTFCLK( ), .Q(ofifoData[674]));
Q_FDP0UA U1460 ( .D(n6519), .QTFCLK( ), .Q(ofifoData[675]));
Q_FDP0UA U1461 ( .D(n6520), .QTFCLK( ), .Q(ofifoData[676]));
Q_FDP0UA U1462 ( .D(n6521), .QTFCLK( ), .Q(ofifoData[677]));
Q_FDP0UA U1463 ( .D(n6522), .QTFCLK( ), .Q(ofifoData[678]));
Q_FDP0UA U1464 ( .D(n6523), .QTFCLK( ), .Q(ofifoData[679]));
Q_FDP0UA U1465 ( .D(n6524), .QTFCLK( ), .Q(ofifoData[680]));
Q_FDP0UA U1466 ( .D(n6525), .QTFCLK( ), .Q(ofifoData[681]));
Q_FDP0UA U1467 ( .D(n6526), .QTFCLK( ), .Q(ofifoData[682]));
Q_FDP0UA U1468 ( .D(n6527), .QTFCLK( ), .Q(ofifoData[683]));
Q_FDP0UA U1469 ( .D(n6528), .QTFCLK( ), .Q(ofifoData[684]));
Q_FDP0UA U1470 ( .D(n6529), .QTFCLK( ), .Q(ofifoData[685]));
Q_FDP0UA U1471 ( .D(n6530), .QTFCLK( ), .Q(ofifoData[686]));
Q_FDP0UA U1472 ( .D(n6531), .QTFCLK( ), .Q(ofifoData[687]));
Q_FDP0UA U1473 ( .D(n6532), .QTFCLK( ), .Q(ofifoData[688]));
Q_FDP0UA U1474 ( .D(n6533), .QTFCLK( ), .Q(ofifoData[689]));
Q_FDP0UA U1475 ( .D(n6534), .QTFCLK( ), .Q(ofifoData[690]));
Q_FDP0UA U1476 ( .D(n6535), .QTFCLK( ), .Q(ofifoData[691]));
Q_FDP0UA U1477 ( .D(n6536), .QTFCLK( ), .Q(ofifoData[692]));
Q_FDP0UA U1478 ( .D(n6537), .QTFCLK( ), .Q(ofifoData[693]));
Q_FDP0UA U1479 ( .D(n6538), .QTFCLK( ), .Q(ofifoData[694]));
Q_FDP0UA U1480 ( .D(n6539), .QTFCLK( ), .Q(ofifoData[695]));
Q_FDP0UA U1481 ( .D(n6540), .QTFCLK( ), .Q(ofifoData[696]));
Q_FDP0UA U1482 ( .D(n6541), .QTFCLK( ), .Q(ofifoData[697]));
Q_FDP0UA U1483 ( .D(n6542), .QTFCLK( ), .Q(ofifoData[698]));
Q_FDP0UA U1484 ( .D(n6543), .QTFCLK( ), .Q(ofifoData[699]));
Q_FDP0UA U1485 ( .D(n6544), .QTFCLK( ), .Q(ofifoData[700]));
Q_FDP0UA U1486 ( .D(n6545), .QTFCLK( ), .Q(ofifoData[701]));
Q_FDP0UA U1487 ( .D(n6546), .QTFCLK( ), .Q(ofifoData[702]));
Q_FDP0UA U1488 ( .D(n6547), .QTFCLK( ), .Q(ofifoData[703]));
Q_FDP0UA U1489 ( .D(n6548), .QTFCLK( ), .Q(ofifoData[704]));
Q_FDP0UA U1490 ( .D(n6549), .QTFCLK( ), .Q(ofifoData[705]));
Q_FDP0UA U1491 ( .D(n6550), .QTFCLK( ), .Q(ofifoData[706]));
Q_FDP0UA U1492 ( .D(n6551), .QTFCLK( ), .Q(ofifoData[707]));
Q_FDP0UA U1493 ( .D(n6552), .QTFCLK( ), .Q(ofifoData[708]));
Q_FDP0UA U1494 ( .D(n6553), .QTFCLK( ), .Q(ofifoData[709]));
Q_FDP0UA U1495 ( .D(n6554), .QTFCLK( ), .Q(ofifoData[710]));
Q_FDP0UA U1496 ( .D(n6555), .QTFCLK( ), .Q(ofifoData[711]));
Q_FDP0UA U1497 ( .D(n6556), .QTFCLK( ), .Q(ofifoData[712]));
Q_FDP0UA U1498 ( .D(n6557), .QTFCLK( ), .Q(ofifoData[713]));
Q_FDP0UA U1499 ( .D(n6558), .QTFCLK( ), .Q(ofifoData[714]));
Q_FDP0UA U1500 ( .D(n6559), .QTFCLK( ), .Q(ofifoData[715]));
Q_FDP0UA U1501 ( .D(n6560), .QTFCLK( ), .Q(ofifoData[716]));
Q_FDP0UA U1502 ( .D(n6561), .QTFCLK( ), .Q(ofifoData[717]));
Q_FDP0UA U1503 ( .D(n6562), .QTFCLK( ), .Q(ofifoData[718]));
Q_FDP0UA U1504 ( .D(n6563), .QTFCLK( ), .Q(ofifoData[719]));
Q_FDP0UA U1505 ( .D(n6564), .QTFCLK( ), .Q(ofifoData[720]));
Q_FDP0UA U1506 ( .D(n6565), .QTFCLK( ), .Q(ofifoData[721]));
Q_FDP0UA U1507 ( .D(n6566), .QTFCLK( ), .Q(ofifoData[722]));
Q_FDP0UA U1508 ( .D(n6567), .QTFCLK( ), .Q(ofifoData[723]));
Q_FDP0UA U1509 ( .D(n6568), .QTFCLK( ), .Q(ofifoData[724]));
Q_FDP0UA U1510 ( .D(n6569), .QTFCLK( ), .Q(ofifoData[725]));
Q_FDP0UA U1511 ( .D(n6570), .QTFCLK( ), .Q(ofifoData[726]));
Q_FDP0UA U1512 ( .D(n6571), .QTFCLK( ), .Q(ofifoData[727]));
Q_FDP0UA U1513 ( .D(n6572), .QTFCLK( ), .Q(ofifoData[728]));
Q_FDP0UA U1514 ( .D(n6573), .QTFCLK( ), .Q(ofifoData[729]));
Q_FDP0UA U1515 ( .D(n6574), .QTFCLK( ), .Q(ofifoData[730]));
Q_FDP0UA U1516 ( .D(n6575), .QTFCLK( ), .Q(ofifoData[731]));
Q_FDP0UA U1517 ( .D(n6576), .QTFCLK( ), .Q(ofifoData[732]));
Q_FDP0UA U1518 ( .D(n6577), .QTFCLK( ), .Q(ofifoData[733]));
Q_FDP0UA U1519 ( .D(n6578), .QTFCLK( ), .Q(ofifoData[734]));
Q_FDP0UA U1520 ( .D(n6579), .QTFCLK( ), .Q(ofifoData[735]));
Q_FDP0UA U1521 ( .D(n6580), .QTFCLK( ), .Q(ofifoData[736]));
Q_FDP0UA U1522 ( .D(n6581), .QTFCLK( ), .Q(ofifoData[737]));
Q_FDP0UA U1523 ( .D(n6582), .QTFCLK( ), .Q(ofifoData[738]));
Q_FDP0UA U1524 ( .D(n6583), .QTFCLK( ), .Q(ofifoData[739]));
Q_FDP0UA U1525 ( .D(n6584), .QTFCLK( ), .Q(ofifoData[740]));
Q_FDP0UA U1526 ( .D(n6585), .QTFCLK( ), .Q(ofifoData[741]));
Q_FDP0UA U1527 ( .D(n6586), .QTFCLK( ), .Q(ofifoData[742]));
Q_FDP0UA U1528 ( .D(n6587), .QTFCLK( ), .Q(ofifoData[743]));
Q_FDP0UA U1529 ( .D(n6588), .QTFCLK( ), .Q(ofifoData[744]));
Q_FDP0UA U1530 ( .D(n6589), .QTFCLK( ), .Q(ofifoData[745]));
Q_FDP0UA U1531 ( .D(n6590), .QTFCLK( ), .Q(ofifoData[746]));
Q_FDP0UA U1532 ( .D(n6591), .QTFCLK( ), .Q(ofifoData[747]));
Q_FDP0UA U1533 ( .D(n6592), .QTFCLK( ), .Q(ofifoData[748]));
Q_FDP0UA U1534 ( .D(n6593), .QTFCLK( ), .Q(ofifoData[749]));
Q_FDP0UA U1535 ( .D(n6594), .QTFCLK( ), .Q(ofifoData[750]));
Q_FDP0UA U1536 ( .D(n6595), .QTFCLK( ), .Q(ofifoData[751]));
Q_FDP0UA U1537 ( .D(n6596), .QTFCLK( ), .Q(ofifoData[752]));
Q_FDP0UA U1538 ( .D(n6597), .QTFCLK( ), .Q(ofifoData[753]));
Q_FDP0UA U1539 ( .D(n6598), .QTFCLK( ), .Q(ofifoData[754]));
Q_FDP0UA U1540 ( .D(n6599), .QTFCLK( ), .Q(ofifoData[755]));
Q_FDP0UA U1541 ( .D(n6600), .QTFCLK( ), .Q(ofifoData[756]));
Q_FDP0UA U1542 ( .D(n6601), .QTFCLK( ), .Q(ofifoData[757]));
Q_FDP0UA U1543 ( .D(n6602), .QTFCLK( ), .Q(ofifoData[758]));
Q_FDP0UA U1544 ( .D(n6603), .QTFCLK( ), .Q(ofifoData[759]));
Q_FDP0UA U1545 ( .D(n6604), .QTFCLK( ), .Q(ofifoData[760]));
Q_FDP0UA U1546 ( .D(n6605), .QTFCLK( ), .Q(ofifoData[761]));
Q_FDP0UA U1547 ( .D(n6606), .QTFCLK( ), .Q(ofifoData[762]));
Q_FDP0UA U1548 ( .D(n6607), .QTFCLK( ), .Q(ofifoData[763]));
Q_FDP0UA U1549 ( .D(n6608), .QTFCLK( ), .Q(ofifoData[764]));
Q_FDP0UA U1550 ( .D(n6609), .QTFCLK( ), .Q(ofifoData[765]));
Q_FDP0UA U1551 ( .D(n6610), .QTFCLK( ), .Q(ofifoData[766]));
Q_FDP0UA U1552 ( .D(n6611), .QTFCLK( ), .Q(ofifoData[767]));
Q_FDP0UA U1553 ( .D(n6639), .QTFCLK( ), .Q(ofifoAddr2[0]));
Q_FDP0UA U1554 ( .D(n1569), .QTFCLK( ), .Q(ofifoAddr2[1]));
Q_FDP0UA U1555 ( .D(n6612), .QTFCLK( ), .Q(ofifoAddr2[2]));
Q_FDP0UA U1556 ( .D(n6613), .QTFCLK( ), .Q(ofifoAddr2[3]));
Q_FDP0UA U1557 ( .D(n6614), .QTFCLK( ), .Q(ofifoAddr2[4]));
Q_FDP0UA U1558 ( .D(n6615), .QTFCLK( ), .Q(ofifoAddr2[5]));
Q_FDP0UA U1559 ( .D(n6616), .QTFCLK( ), .Q(ofifoAddr2[6]));
Q_FDP0UA U1560 ( .D(n6617), .QTFCLK( ), .Q(ofifoAddr2[7]));
Q_FDP0UA U1561 ( .D(n6618), .QTFCLK( ), .Q(ofifoAddr2[8]));
Q_FDP0UA U1562 ( .D(n6619), .QTFCLK( ), .Q(ofifoAddr2[9]));
Q_FDP0UA U1563 ( .D(n6620), .QTFCLK( ), .Q(ofifoAddr2[10]));
Q_FDP0UA U1564 ( .D(n6621), .QTFCLK( ), .Q(ofifoAddr2[11]));
Q_FDP0UA U1565 ( .D(n6622), .QTFCLK( ), .Q(ofifoAddr2[12]));
Q_FDP0UA U1566 ( .D(n6623), .QTFCLK( ), .Q(ofifoAddr2[13]));
Q_FDP0UA U1567 ( .D(n6624), .QTFCLK( ), .Q(ofifoAddr2[14]));
Q_FDP0UA U1568 ( .D(n1570), .QTFCLK( ), .Q(ofifoAddr1[0]));
Q_FDP0UA U1569 ( .D(n6625), .QTFCLK( ), .Q(ofifoAddr1[1]));
Q_FDP0UA U1570 ( .D(n6626), .QTFCLK( ), .Q(ofifoAddr1[2]));
Q_FDP0UA U1571 ( .D(n6627), .QTFCLK( ), .Q(ofifoAddr1[3]));
Q_FDP0UA U1572 ( .D(n6628), .QTFCLK( ), .Q(ofifoAddr1[4]));
Q_FDP0UA U1573 ( .D(n6629), .QTFCLK( ), .Q(ofifoAddr1[5]));
Q_FDP0UA U1574 ( .D(n6630), .QTFCLK( ), .Q(ofifoAddr1[6]));
Q_FDP0UA U1575 ( .D(n6631), .QTFCLK( ), .Q(ofifoAddr1[7]));
Q_FDP0UA U1576 ( .D(n6632), .QTFCLK( ), .Q(ofifoAddr1[8]));
Q_FDP0UA U1577 ( .D(n6633), .QTFCLK( ), .Q(ofifoAddr1[9]));
Q_FDP0UA U1578 ( .D(n6634), .QTFCLK( ), .Q(ofifoAddr1[10]));
Q_FDP0UA U1579 ( .D(n6635), .QTFCLK( ), .Q(ofifoAddr1[11]));
Q_FDP0UA U1580 ( .D(n6636), .QTFCLK( ), .Q(ofifoAddr1[12]));
Q_FDP0UA U1581 ( .D(n6637), .QTFCLK( ), .Q(ofifoAddr1[13]));
Q_FDP0UA U1582 ( .D(n6638), .QTFCLK( ), .Q(ofifoAddr1[14]));
Q_FDP0UA U1583 ( .D(n6639), .QTFCLK( ), .Q(ofifoAddr0[0]));
Q_FDP0UA U1584 ( .D(n6640), .QTFCLK( ), .Q(ofifoAddr0[1]));
Q_FDP0UA U1585 ( .D(n6641), .QTFCLK( ), .Q(ofifoAddr0[2]));
Q_FDP0UA U1586 ( .D(n6642), .QTFCLK( ), .Q(ofifoAddr0[3]));
Q_FDP0UA U1587 ( .D(n6643), .QTFCLK( ), .Q(ofifoAddr0[4]));
Q_FDP0UA U1588 ( .D(n6644), .QTFCLK( ), .Q(ofifoAddr0[5]));
Q_FDP0UA U1589 ( .D(n6645), .QTFCLK( ), .Q(ofifoAddr0[6]));
Q_FDP0UA U1590 ( .D(n6646), .QTFCLK( ), .Q(ofifoAddr0[7]));
Q_FDP0UA U1591 ( .D(n6647), .QTFCLK( ), .Q(ofifoAddr0[8]));
Q_FDP0UA U1592 ( .D(n6648), .QTFCLK( ), .Q(ofifoAddr0[9]));
Q_FDP0UA U1593 ( .D(n6649), .QTFCLK( ), .Q(ofifoAddr0[10]));
Q_FDP0UA U1594 ( .D(n6650), .QTFCLK( ), .Q(ofifoAddr0[11]));
Q_FDP0UA U1595 ( .D(n6651), .QTFCLK( ), .Q(ofifoAddr0[12]));
Q_FDP0UA U1596 ( .D(n6652), .QTFCLK( ), .Q(ofifoAddr0[13]));
Q_FDP0UA U1597 ( .D(n6653), .QTFCLK( ), .Q(ofifoAddr0[14]));
Q_AN02 U1598 ( .A0(n6720), .A1(ofifoAddr0N[14]), .Z(n6653));
Q_AN02 U1599 ( .A0(n6720), .A1(ofifoAddr0N[13]), .Z(n6652));
Q_AN02 U1600 ( .A0(n6720), .A1(ofifoAddr0N[12]), .Z(n6651));
Q_AN02 U1601 ( .A0(n6720), .A1(ofifoAddr0N[11]), .Z(n6650));
Q_AN02 U1602 ( .A0(n6720), .A1(ofifoAddr0N[10]), .Z(n6649));
Q_AN02 U1603 ( .A0(n6720), .A1(ofifoAddr0N[9]), .Z(n6648));
Q_AN02 U1604 ( .A0(n6720), .A1(ofifoAddr0N[8]), .Z(n6647));
Q_AN02 U1605 ( .A0(n6720), .A1(ofifoAddr0N[7]), .Z(n6646));
Q_AN02 U1606 ( .A0(n6720), .A1(ofifoAddr0N[6]), .Z(n6645));
Q_AN02 U1607 ( .A0(n6720), .A1(ofifoAddr0N[5]), .Z(n6644));
Q_AN02 U1608 ( .A0(n6720), .A1(ofifoAddr0N[4]), .Z(n6643));
Q_AN02 U1609 ( .A0(n6720), .A1(ofifoAddr0N[3]), .Z(n6642));
Q_AN02 U1610 ( .A0(n6720), .A1(ofifoAddr0N[2]), .Z(n6641));
Q_AN02 U1611 ( .A0(n6720), .A1(ofifoAddr0N[1]), .Z(n6640));
Q_AN02 U1612 ( .A0(n6720), .A1(ofifoAddr0N[0]), .Z(n6639));
Q_AN02 U1613 ( .A0(n6720), .A1(ofifoAddr1N[14]), .Z(n6638));
Q_AN02 U1614 ( .A0(n6720), .A1(ofifoAddr1N[13]), .Z(n6637));
Q_AN02 U1615 ( .A0(n6720), .A1(ofifoAddr1N[12]), .Z(n6636));
Q_AN02 U1616 ( .A0(n6720), .A1(ofifoAddr1N[11]), .Z(n6635));
Q_AN02 U1617 ( .A0(n6720), .A1(ofifoAddr1N[10]), .Z(n6634));
Q_AN02 U1618 ( .A0(n6720), .A1(ofifoAddr1N[9]), .Z(n6633));
Q_AN02 U1619 ( .A0(n6720), .A1(ofifoAddr1N[8]), .Z(n6632));
Q_AN02 U1620 ( .A0(n6720), .A1(ofifoAddr1N[7]), .Z(n6631));
Q_AN02 U1621 ( .A0(n6720), .A1(ofifoAddr1N[6]), .Z(n6630));
Q_AN02 U1622 ( .A0(n6720), .A1(ofifoAddr1N[5]), .Z(n6629));
Q_AN02 U1623 ( .A0(n6720), .A1(ofifoAddr1N[4]), .Z(n6628));
Q_AN02 U1624 ( .A0(n6720), .A1(ofifoAddr1N[3]), .Z(n6627));
Q_AN02 U1625 ( .A0(n6720), .A1(ofifoAddr1N[2]), .Z(n6626));
Q_AN02 U1626 ( .A0(n6720), .A1(ofifoAddr1N[1]), .Z(n6625));
Q_AN02 U1627 ( .A0(n6720), .A1(ofifoAddr2N[14]), .Z(n6624));
Q_AN02 U1628 ( .A0(n6720), .A1(ofifoAddr2N[13]), .Z(n6623));
Q_AN02 U1629 ( .A0(n6720), .A1(ofifoAddr2N[12]), .Z(n6622));
Q_AN02 U1630 ( .A0(n6720), .A1(ofifoAddr2N[11]), .Z(n6621));
Q_AN02 U1631 ( .A0(n6720), .A1(ofifoAddr2N[10]), .Z(n6620));
Q_AN02 U1632 ( .A0(n6720), .A1(ofifoAddr2N[9]), .Z(n6619));
Q_AN02 U1633 ( .A0(n6720), .A1(ofifoAddr2N[8]), .Z(n6618));
Q_AN02 U1634 ( .A0(n6720), .A1(ofifoAddr2N[7]), .Z(n6617));
Q_AN02 U1635 ( .A0(n6720), .A1(ofifoAddr2N[6]), .Z(n6616));
Q_AN02 U1636 ( .A0(n6720), .A1(ofifoAddr2N[5]), .Z(n6615));
Q_AN02 U1637 ( .A0(n6720), .A1(ofifoAddr2N[4]), .Z(n6614));
Q_AN02 U1638 ( .A0(n6720), .A1(ofifoAddr2N[3]), .Z(n6613));
Q_AN02 U1639 ( .A0(n6720), .A1(ofifoAddr2N[2]), .Z(n6612));
Q_AN02 U1640 ( .A0(n6720), .A1(ofifoDataN[767]), .Z(n6611));
Q_AN02 U1641 ( .A0(n6720), .A1(ofifoDataN[766]), .Z(n6610));
Q_AN02 U1642 ( .A0(n6720), .A1(ofifoDataN[765]), .Z(n6609));
Q_AN02 U1643 ( .A0(n6720), .A1(ofifoDataN[764]), .Z(n6608));
Q_AN02 U1644 ( .A0(n6720), .A1(ofifoDataN[763]), .Z(n6607));
Q_AN02 U1645 ( .A0(n6720), .A1(ofifoDataN[762]), .Z(n6606));
Q_AN02 U1646 ( .A0(n6720), .A1(ofifoDataN[761]), .Z(n6605));
Q_AN02 U1647 ( .A0(n6720), .A1(ofifoDataN[760]), .Z(n6604));
Q_AN02 U1648 ( .A0(n6720), .A1(ofifoDataN[759]), .Z(n6603));
Q_AN02 U1649 ( .A0(n6720), .A1(ofifoDataN[758]), .Z(n6602));
Q_AN02 U1650 ( .A0(n6720), .A1(ofifoDataN[757]), .Z(n6601));
Q_AN02 U1651 ( .A0(n6720), .A1(ofifoDataN[756]), .Z(n6600));
Q_AN02 U1652 ( .A0(n6720), .A1(ofifoDataN[755]), .Z(n6599));
Q_AN02 U1653 ( .A0(n6720), .A1(ofifoDataN[754]), .Z(n6598));
Q_AN02 U1654 ( .A0(n6720), .A1(ofifoDataN[753]), .Z(n6597));
Q_AN02 U1655 ( .A0(n6720), .A1(ofifoDataN[752]), .Z(n6596));
Q_AN02 U1656 ( .A0(n6720), .A1(ofifoDataN[751]), .Z(n6595));
Q_AN02 U1657 ( .A0(n6720), .A1(ofifoDataN[750]), .Z(n6594));
Q_AN02 U1658 ( .A0(n6720), .A1(ofifoDataN[749]), .Z(n6593));
Q_AN02 U1659 ( .A0(n6720), .A1(ofifoDataN[748]), .Z(n6592));
Q_AN02 U1660 ( .A0(n6720), .A1(ofifoDataN[747]), .Z(n6591));
Q_AN02 U1661 ( .A0(n6720), .A1(ofifoDataN[746]), .Z(n6590));
Q_AN02 U1662 ( .A0(n6720), .A1(ofifoDataN[745]), .Z(n6589));
Q_AN02 U1663 ( .A0(n6720), .A1(ofifoDataN[744]), .Z(n6588));
Q_AN02 U1664 ( .A0(n6720), .A1(ofifoDataN[743]), .Z(n6587));
Q_AN02 U1665 ( .A0(n6720), .A1(ofifoDataN[742]), .Z(n6586));
Q_AN02 U1666 ( .A0(n6720), .A1(ofifoDataN[741]), .Z(n6585));
Q_AN02 U1667 ( .A0(n6720), .A1(ofifoDataN[740]), .Z(n6584));
Q_AN02 U1668 ( .A0(n6720), .A1(ofifoDataN[739]), .Z(n6583));
Q_AN02 U1669 ( .A0(n6720), .A1(ofifoDataN[738]), .Z(n6582));
Q_AN02 U1670 ( .A0(n6720), .A1(ofifoDataN[737]), .Z(n6581));
Q_AN02 U1671 ( .A0(n6720), .A1(ofifoDataN[736]), .Z(n6580));
Q_AN02 U1672 ( .A0(n6720), .A1(ofifoDataN[735]), .Z(n6579));
Q_AN02 U1673 ( .A0(n6720), .A1(ofifoDataN[734]), .Z(n6578));
Q_AN02 U1674 ( .A0(n6720), .A1(ofifoDataN[733]), .Z(n6577));
Q_AN02 U1675 ( .A0(n6720), .A1(ofifoDataN[732]), .Z(n6576));
Q_AN02 U1676 ( .A0(n6720), .A1(ofifoDataN[731]), .Z(n6575));
Q_AN02 U1677 ( .A0(n6720), .A1(ofifoDataN[730]), .Z(n6574));
Q_AN02 U1678 ( .A0(n6720), .A1(ofifoDataN[729]), .Z(n6573));
Q_AN02 U1679 ( .A0(n6720), .A1(ofifoDataN[728]), .Z(n6572));
Q_AN02 U1680 ( .A0(n6720), .A1(ofifoDataN[727]), .Z(n6571));
Q_AN02 U1681 ( .A0(n6720), .A1(ofifoDataN[726]), .Z(n6570));
Q_AN02 U1682 ( .A0(n6720), .A1(ofifoDataN[725]), .Z(n6569));
Q_AN02 U1683 ( .A0(n6720), .A1(ofifoDataN[724]), .Z(n6568));
Q_AN02 U1684 ( .A0(n6720), .A1(ofifoDataN[723]), .Z(n6567));
Q_AN02 U1685 ( .A0(n6720), .A1(ofifoDataN[722]), .Z(n6566));
Q_AN02 U1686 ( .A0(n6720), .A1(ofifoDataN[721]), .Z(n6565));
Q_AN02 U1687 ( .A0(n6720), .A1(ofifoDataN[720]), .Z(n6564));
Q_AN02 U1688 ( .A0(n6720), .A1(ofifoDataN[719]), .Z(n6563));
Q_AN02 U1689 ( .A0(n6720), .A1(ofifoDataN[718]), .Z(n6562));
Q_AN02 U1690 ( .A0(n6720), .A1(ofifoDataN[717]), .Z(n6561));
Q_AN02 U1691 ( .A0(n6720), .A1(ofifoDataN[716]), .Z(n6560));
Q_AN02 U1692 ( .A0(n6720), .A1(ofifoDataN[715]), .Z(n6559));
Q_AN02 U1693 ( .A0(n6720), .A1(ofifoDataN[714]), .Z(n6558));
Q_AN02 U1694 ( .A0(n6720), .A1(ofifoDataN[713]), .Z(n6557));
Q_AN02 U1695 ( .A0(n6720), .A1(ofifoDataN[712]), .Z(n6556));
Q_AN02 U1696 ( .A0(n6720), .A1(ofifoDataN[711]), .Z(n6555));
Q_AN02 U1697 ( .A0(n6720), .A1(ofifoDataN[710]), .Z(n6554));
Q_AN02 U1698 ( .A0(n6720), .A1(ofifoDataN[709]), .Z(n6553));
Q_AN02 U1699 ( .A0(n6720), .A1(ofifoDataN[708]), .Z(n6552));
Q_AN02 U1700 ( .A0(n6720), .A1(ofifoDataN[707]), .Z(n6551));
Q_AN02 U1701 ( .A0(n6720), .A1(ofifoDataN[706]), .Z(n6550));
Q_AN02 U1702 ( .A0(n6720), .A1(ofifoDataN[705]), .Z(n6549));
Q_AN02 U1703 ( .A0(n6720), .A1(ofifoDataN[704]), .Z(n6548));
Q_AN02 U1704 ( .A0(n6720), .A1(ofifoDataN[703]), .Z(n6547));
Q_AN02 U1705 ( .A0(n6720), .A1(ofifoDataN[702]), .Z(n6546));
Q_AN02 U1706 ( .A0(n6720), .A1(ofifoDataN[701]), .Z(n6545));
Q_AN02 U1707 ( .A0(n6720), .A1(ofifoDataN[700]), .Z(n6544));
Q_AN02 U1708 ( .A0(n6720), .A1(ofifoDataN[699]), .Z(n6543));
Q_AN02 U1709 ( .A0(n6720), .A1(ofifoDataN[698]), .Z(n6542));
Q_AN02 U1710 ( .A0(n6720), .A1(ofifoDataN[697]), .Z(n6541));
Q_AN02 U1711 ( .A0(n6720), .A1(ofifoDataN[696]), .Z(n6540));
Q_AN02 U1712 ( .A0(n6720), .A1(ofifoDataN[695]), .Z(n6539));
Q_AN02 U1713 ( .A0(n6720), .A1(ofifoDataN[694]), .Z(n6538));
Q_AN02 U1714 ( .A0(n6720), .A1(ofifoDataN[693]), .Z(n6537));
Q_AN02 U1715 ( .A0(n6720), .A1(ofifoDataN[692]), .Z(n6536));
Q_AN02 U1716 ( .A0(n6720), .A1(ofifoDataN[691]), .Z(n6535));
Q_AN02 U1717 ( .A0(n6720), .A1(ofifoDataN[690]), .Z(n6534));
Q_AN02 U1718 ( .A0(n6720), .A1(ofifoDataN[689]), .Z(n6533));
Q_AN02 U1719 ( .A0(n6720), .A1(ofifoDataN[688]), .Z(n6532));
Q_AN02 U1720 ( .A0(n6720), .A1(ofifoDataN[687]), .Z(n6531));
Q_AN02 U1721 ( .A0(n6720), .A1(ofifoDataN[686]), .Z(n6530));
Q_AN02 U1722 ( .A0(n6720), .A1(ofifoDataN[685]), .Z(n6529));
Q_AN02 U1723 ( .A0(n6720), .A1(ofifoDataN[684]), .Z(n6528));
Q_AN02 U1724 ( .A0(n6720), .A1(ofifoDataN[683]), .Z(n6527));
Q_AN02 U1725 ( .A0(n6720), .A1(ofifoDataN[682]), .Z(n6526));
Q_AN02 U1726 ( .A0(n6720), .A1(ofifoDataN[681]), .Z(n6525));
Q_AN02 U1727 ( .A0(n6720), .A1(ofifoDataN[680]), .Z(n6524));
Q_AN02 U1728 ( .A0(n6720), .A1(ofifoDataN[679]), .Z(n6523));
Q_AN02 U1729 ( .A0(n6720), .A1(ofifoDataN[678]), .Z(n6522));
Q_AN02 U1730 ( .A0(n6720), .A1(ofifoDataN[677]), .Z(n6521));
Q_AN02 U1731 ( .A0(n6720), .A1(ofifoDataN[676]), .Z(n6520));
Q_AN02 U1732 ( .A0(n6720), .A1(ofifoDataN[675]), .Z(n6519));
Q_AN02 U1733 ( .A0(n6720), .A1(ofifoDataN[674]), .Z(n6518));
Q_AN02 U1734 ( .A0(n6720), .A1(ofifoDataN[673]), .Z(n6517));
Q_AN02 U1735 ( .A0(n6720), .A1(ofifoDataN[672]), .Z(n6516));
Q_AN02 U1736 ( .A0(n6720), .A1(ofifoDataN[671]), .Z(n6515));
Q_AN02 U1737 ( .A0(n6720), .A1(ofifoDataN[670]), .Z(n6514));
Q_AN02 U1738 ( .A0(n6720), .A1(ofifoDataN[669]), .Z(n6513));
Q_AN02 U1739 ( .A0(n6720), .A1(ofifoDataN[668]), .Z(n6512));
Q_AN02 U1740 ( .A0(n6720), .A1(ofifoDataN[667]), .Z(n6511));
Q_AN02 U1741 ( .A0(n6720), .A1(ofifoDataN[666]), .Z(n6510));
Q_AN02 U1742 ( .A0(n6720), .A1(ofifoDataN[665]), .Z(n6509));
Q_AN02 U1743 ( .A0(n6720), .A1(ofifoDataN[664]), .Z(n6508));
Q_AN02 U1744 ( .A0(n6720), .A1(ofifoDataN[663]), .Z(n6507));
Q_AN02 U1745 ( .A0(n6720), .A1(ofifoDataN[662]), .Z(n6506));
Q_AN02 U1746 ( .A0(n6720), .A1(ofifoDataN[661]), .Z(n6505));
Q_AN02 U1747 ( .A0(n6720), .A1(ofifoDataN[660]), .Z(n6504));
Q_AN02 U1748 ( .A0(n6720), .A1(ofifoDataN[659]), .Z(n6503));
Q_AN02 U1749 ( .A0(n6720), .A1(ofifoDataN[658]), .Z(n6502));
Q_AN02 U1750 ( .A0(n6720), .A1(ofifoDataN[657]), .Z(n6501));
Q_AN02 U1751 ( .A0(n6720), .A1(ofifoDataN[656]), .Z(n6500));
Q_AN02 U1752 ( .A0(n6720), .A1(ofifoDataN[655]), .Z(n6499));
Q_AN02 U1753 ( .A0(n6720), .A1(ofifoDataN[654]), .Z(n6498));
Q_AN02 U1754 ( .A0(n6720), .A1(ofifoDataN[653]), .Z(n6497));
Q_AN02 U1755 ( .A0(n6720), .A1(ofifoDataN[652]), .Z(n6496));
Q_AN02 U1756 ( .A0(n6720), .A1(ofifoDataN[651]), .Z(n6495));
Q_AN02 U1757 ( .A0(n6720), .A1(ofifoDataN[650]), .Z(n6494));
Q_AN02 U1758 ( .A0(n6720), .A1(ofifoDataN[649]), .Z(n6493));
Q_AN02 U1759 ( .A0(n6720), .A1(ofifoDataN[648]), .Z(n6492));
Q_AN02 U1760 ( .A0(n6720), .A1(ofifoDataN[647]), .Z(n6491));
Q_AN02 U1761 ( .A0(n6720), .A1(ofifoDataN[646]), .Z(n6490));
Q_AN02 U1762 ( .A0(n6720), .A1(ofifoDataN[645]), .Z(n6489));
Q_AN02 U1763 ( .A0(n6720), .A1(ofifoDataN[644]), .Z(n6488));
Q_AN02 U1764 ( .A0(n6720), .A1(ofifoDataN[643]), .Z(n6487));
Q_AN02 U1765 ( .A0(n6720), .A1(ofifoDataN[642]), .Z(n6486));
Q_AN02 U1766 ( .A0(n6720), .A1(ofifoDataN[641]), .Z(n6485));
Q_AN02 U1767 ( .A0(n6720), .A1(ofifoDataN[640]), .Z(n6484));
Q_AN02 U1768 ( .A0(n6720), .A1(ofifoDataN[639]), .Z(n6483));
Q_AN02 U1769 ( .A0(n6720), .A1(ofifoDataN[638]), .Z(n6482));
Q_AN02 U1770 ( .A0(n6720), .A1(ofifoDataN[637]), .Z(n6481));
Q_AN02 U1771 ( .A0(n6720), .A1(ofifoDataN[636]), .Z(n6480));
Q_AN02 U1772 ( .A0(n6720), .A1(ofifoDataN[635]), .Z(n6479));
Q_AN02 U1773 ( .A0(n6720), .A1(ofifoDataN[634]), .Z(n6478));
Q_AN02 U1774 ( .A0(n6720), .A1(ofifoDataN[633]), .Z(n6477));
Q_AN02 U1775 ( .A0(n6720), .A1(ofifoDataN[632]), .Z(n6476));
Q_AN02 U1776 ( .A0(n6720), .A1(ofifoDataN[631]), .Z(n6475));
Q_AN02 U1777 ( .A0(n6720), .A1(ofifoDataN[630]), .Z(n6474));
Q_AN02 U1778 ( .A0(n6720), .A1(ofifoDataN[629]), .Z(n6473));
Q_AN02 U1779 ( .A0(n6720), .A1(ofifoDataN[628]), .Z(n6472));
Q_AN02 U1780 ( .A0(n6720), .A1(ofifoDataN[627]), .Z(n6471));
Q_AN02 U1781 ( .A0(n6720), .A1(ofifoDataN[626]), .Z(n6470));
Q_AN02 U1782 ( .A0(n6720), .A1(ofifoDataN[625]), .Z(n6469));
Q_AN02 U1783 ( .A0(n6720), .A1(ofifoDataN[624]), .Z(n6468));
Q_AN02 U1784 ( .A0(n6720), .A1(ofifoDataN[623]), .Z(n6467));
Q_AN02 U1785 ( .A0(n6720), .A1(ofifoDataN[622]), .Z(n6466));
Q_AN02 U1786 ( .A0(n6720), .A1(ofifoDataN[621]), .Z(n6465));
Q_AN02 U1787 ( .A0(n6720), .A1(ofifoDataN[620]), .Z(n6464));
Q_AN02 U1788 ( .A0(n6720), .A1(ofifoDataN[619]), .Z(n6463));
Q_AN02 U1789 ( .A0(n6720), .A1(ofifoDataN[618]), .Z(n6462));
Q_AN02 U1790 ( .A0(n6720), .A1(ofifoDataN[617]), .Z(n6461));
Q_AN02 U1791 ( .A0(n6720), .A1(ofifoDataN[616]), .Z(n6460));
Q_AN02 U1792 ( .A0(n6720), .A1(ofifoDataN[615]), .Z(n6459));
Q_AN02 U1793 ( .A0(n6720), .A1(ofifoDataN[614]), .Z(n6458));
Q_AN02 U1794 ( .A0(n6720), .A1(ofifoDataN[613]), .Z(n6457));
Q_AN02 U1795 ( .A0(n6720), .A1(ofifoDataN[612]), .Z(n6456));
Q_AN02 U1796 ( .A0(n6720), .A1(ofifoDataN[611]), .Z(n6455));
Q_AN02 U1797 ( .A0(n6720), .A1(ofifoDataN[610]), .Z(n6454));
Q_AN02 U1798 ( .A0(n6720), .A1(ofifoDataN[609]), .Z(n6453));
Q_AN02 U1799 ( .A0(n6720), .A1(ofifoDataN[608]), .Z(n6452));
Q_AN02 U1800 ( .A0(n6720), .A1(ofifoDataN[607]), .Z(n6451));
Q_AN02 U1801 ( .A0(n6720), .A1(ofifoDataN[606]), .Z(n6450));
Q_AN02 U1802 ( .A0(n6720), .A1(ofifoDataN[605]), .Z(n6449));
Q_AN02 U1803 ( .A0(n6720), .A1(ofifoDataN[604]), .Z(n6448));
Q_AN02 U1804 ( .A0(n6720), .A1(ofifoDataN[603]), .Z(n6447));
Q_AN02 U1805 ( .A0(n6720), .A1(ofifoDataN[602]), .Z(n6446));
Q_AN02 U1806 ( .A0(n6720), .A1(ofifoDataN[601]), .Z(n6445));
Q_AN02 U1807 ( .A0(n6720), .A1(ofifoDataN[600]), .Z(n6444));
Q_AN02 U1808 ( .A0(n6720), .A1(ofifoDataN[599]), .Z(n6443));
Q_AN02 U1809 ( .A0(n6720), .A1(ofifoDataN[598]), .Z(n6442));
Q_AN02 U1810 ( .A0(n6720), .A1(ofifoDataN[597]), .Z(n6441));
Q_AN02 U1811 ( .A0(n6720), .A1(ofifoDataN[596]), .Z(n6440));
Q_AN02 U1812 ( .A0(n6720), .A1(ofifoDataN[595]), .Z(n6439));
Q_AN02 U1813 ( .A0(n6720), .A1(ofifoDataN[594]), .Z(n6438));
Q_AN02 U1814 ( .A0(n6720), .A1(ofifoDataN[593]), .Z(n6437));
Q_AN02 U1815 ( .A0(n6720), .A1(ofifoDataN[592]), .Z(n6436));
Q_AN02 U1816 ( .A0(n6720), .A1(ofifoDataN[591]), .Z(n6435));
Q_AN02 U1817 ( .A0(n6720), .A1(ofifoDataN[590]), .Z(n6434));
Q_AN02 U1818 ( .A0(n6720), .A1(ofifoDataN[589]), .Z(n6433));
Q_AN02 U1819 ( .A0(n6720), .A1(ofifoDataN[588]), .Z(n6432));
Q_AN02 U1820 ( .A0(n6720), .A1(ofifoDataN[587]), .Z(n6431));
Q_AN02 U1821 ( .A0(n6720), .A1(ofifoDataN[586]), .Z(n6430));
Q_AN02 U1822 ( .A0(n6720), .A1(ofifoDataN[585]), .Z(n6429));
Q_AN02 U1823 ( .A0(n6720), .A1(ofifoDataN[584]), .Z(n6428));
Q_AN02 U1824 ( .A0(n6720), .A1(ofifoDataN[583]), .Z(n6427));
Q_AN02 U1825 ( .A0(n6720), .A1(ofifoDataN[582]), .Z(n6426));
Q_AN02 U1826 ( .A0(n6720), .A1(ofifoDataN[581]), .Z(n6425));
Q_AN02 U1827 ( .A0(n6720), .A1(ofifoDataN[580]), .Z(n6424));
Q_AN02 U1828 ( .A0(n6720), .A1(ofifoDataN[579]), .Z(n6423));
Q_AN02 U1829 ( .A0(n6720), .A1(ofifoDataN[578]), .Z(n6422));
Q_AN02 U1830 ( .A0(n6720), .A1(ofifoDataN[577]), .Z(n6421));
Q_AN02 U1831 ( .A0(n6720), .A1(ofifoDataN[576]), .Z(n6420));
Q_AN02 U1832 ( .A0(n6720), .A1(ofifoDataN[575]), .Z(n6419));
Q_AN02 U1833 ( .A0(n6720), .A1(ofifoDataN[574]), .Z(n6418));
Q_AN02 U1834 ( .A0(n6720), .A1(ofifoDataN[573]), .Z(n6417));
Q_AN02 U1835 ( .A0(n6720), .A1(ofifoDataN[572]), .Z(n6416));
Q_AN02 U1836 ( .A0(n6720), .A1(ofifoDataN[571]), .Z(n6415));
Q_AN02 U1837 ( .A0(n6720), .A1(ofifoDataN[570]), .Z(n6414));
Q_AN02 U1838 ( .A0(n6720), .A1(ofifoDataN[569]), .Z(n6413));
Q_AN02 U1839 ( .A0(n6720), .A1(ofifoDataN[568]), .Z(n6412));
Q_AN02 U1840 ( .A0(n6720), .A1(ofifoDataN[567]), .Z(n6411));
Q_AN02 U1841 ( .A0(n6720), .A1(ofifoDataN[566]), .Z(n6410));
Q_AN02 U1842 ( .A0(n6720), .A1(ofifoDataN[565]), .Z(n6409));
Q_AN02 U1843 ( .A0(n6720), .A1(ofifoDataN[564]), .Z(n6408));
Q_AN02 U1844 ( .A0(n6720), .A1(ofifoDataN[563]), .Z(n6407));
Q_AN02 U1845 ( .A0(n6720), .A1(ofifoDataN[562]), .Z(n6406));
Q_AN02 U1846 ( .A0(n6720), .A1(ofifoDataN[561]), .Z(n6405));
Q_AN02 U1847 ( .A0(n6720), .A1(ofifoDataN[560]), .Z(n6404));
Q_AN02 U1848 ( .A0(n6720), .A1(ofifoDataN[559]), .Z(n6403));
Q_AN02 U1849 ( .A0(n6720), .A1(ofifoDataN[558]), .Z(n6402));
Q_AN02 U1850 ( .A0(n6720), .A1(ofifoDataN[557]), .Z(n6401));
Q_AN02 U1851 ( .A0(n6720), .A1(ofifoDataN[556]), .Z(n6400));
Q_AN02 U1852 ( .A0(n6720), .A1(ofifoDataN[555]), .Z(n6399));
Q_AN02 U1853 ( .A0(n6720), .A1(ofifoDataN[554]), .Z(n6398));
Q_AN02 U1854 ( .A0(n6720), .A1(ofifoDataN[553]), .Z(n6397));
Q_AN02 U1855 ( .A0(n6720), .A1(ofifoDataN[552]), .Z(n6396));
Q_AN02 U1856 ( .A0(n6720), .A1(ofifoDataN[551]), .Z(n6395));
Q_AN02 U1857 ( .A0(n6720), .A1(ofifoDataN[550]), .Z(n6394));
Q_AN02 U1858 ( .A0(n6720), .A1(ofifoDataN[549]), .Z(n6393));
Q_AN02 U1859 ( .A0(n6720), .A1(ofifoDataN[548]), .Z(n6392));
Q_AN02 U1860 ( .A0(n6720), .A1(ofifoDataN[547]), .Z(n6391));
Q_AN02 U1861 ( .A0(n6720), .A1(ofifoDataN[546]), .Z(n6390));
Q_AN02 U1862 ( .A0(n6720), .A1(ofifoDataN[545]), .Z(n6389));
Q_AN02 U1863 ( .A0(n6720), .A1(ofifoDataN[544]), .Z(n6388));
Q_AN02 U1864 ( .A0(n6720), .A1(ofifoDataN[543]), .Z(n6387));
Q_AN02 U1865 ( .A0(n6720), .A1(ofifoDataN[542]), .Z(n6386));
Q_AN02 U1866 ( .A0(n6720), .A1(ofifoDataN[541]), .Z(n6385));
Q_AN02 U1867 ( .A0(n6720), .A1(ofifoDataN[540]), .Z(n6384));
Q_AN02 U1868 ( .A0(n6720), .A1(ofifoDataN[539]), .Z(n6383));
Q_AN02 U1869 ( .A0(n6720), .A1(ofifoDataN[538]), .Z(n6382));
Q_AN02 U1870 ( .A0(n6720), .A1(ofifoDataN[537]), .Z(n6381));
Q_AN02 U1871 ( .A0(n6720), .A1(ofifoDataN[536]), .Z(n6380));
Q_AN02 U1872 ( .A0(n6720), .A1(ofifoDataN[535]), .Z(n6379));
Q_AN02 U1873 ( .A0(n6720), .A1(ofifoDataN[534]), .Z(n6378));
Q_AN02 U1874 ( .A0(n6720), .A1(ofifoDataN[533]), .Z(n6377));
Q_AN02 U1875 ( .A0(n6720), .A1(ofifoDataN[532]), .Z(n6376));
Q_AN02 U1876 ( .A0(n6720), .A1(ofifoDataN[531]), .Z(n6375));
Q_AN02 U1877 ( .A0(n6720), .A1(ofifoDataN[530]), .Z(n6374));
Q_AN02 U1878 ( .A0(n6720), .A1(ofifoDataN[529]), .Z(n6373));
Q_AN02 U1879 ( .A0(n6720), .A1(ofifoDataN[528]), .Z(n6372));
Q_AN02 U1880 ( .A0(n6720), .A1(ofifoDataN[527]), .Z(n6371));
Q_AN02 U1881 ( .A0(n6720), .A1(ofifoDataN[526]), .Z(n6370));
Q_AN02 U1882 ( .A0(n6720), .A1(ofifoDataN[525]), .Z(n6369));
Q_AN02 U1883 ( .A0(n6720), .A1(ofifoDataN[524]), .Z(n6368));
Q_AN02 U1884 ( .A0(n6720), .A1(ofifoDataN[523]), .Z(n6367));
Q_AN02 U1885 ( .A0(n6720), .A1(ofifoDataN[522]), .Z(n6366));
Q_AN02 U1886 ( .A0(n6720), .A1(ofifoDataN[521]), .Z(n6365));
Q_AN02 U1887 ( .A0(n6720), .A1(ofifoDataN[520]), .Z(n6364));
Q_AN02 U1888 ( .A0(n6720), .A1(ofifoDataN[519]), .Z(n6363));
Q_AN02 U1889 ( .A0(n6720), .A1(ofifoDataN[518]), .Z(n6362));
Q_AN02 U1890 ( .A0(n6720), .A1(ofifoDataN[517]), .Z(n6361));
Q_AN02 U1891 ( .A0(n6720), .A1(ofifoDataN[516]), .Z(n6360));
Q_AN02 U1892 ( .A0(n6720), .A1(ofifoDataN[515]), .Z(n6359));
Q_AN02 U1893 ( .A0(n6720), .A1(ofifoDataN[514]), .Z(n6358));
Q_AN02 U1894 ( .A0(n6720), .A1(ofifoDataN[513]), .Z(n6357));
Q_AN02 U1895 ( .A0(n6720), .A1(ofifoDataN[512]), .Z(n6356));
Q_AN02 U1896 ( .A0(n6720), .A1(ofifoDataN[511]), .Z(n6355));
Q_AN02 U1897 ( .A0(n6720), .A1(ofifoDataN[510]), .Z(n6354));
Q_AN02 U1898 ( .A0(n6720), .A1(ofifoDataN[509]), .Z(n6353));
Q_AN02 U1899 ( .A0(n6720), .A1(ofifoDataN[508]), .Z(n6352));
Q_AN02 U1900 ( .A0(n6720), .A1(ofifoDataN[507]), .Z(n6351));
Q_AN02 U1901 ( .A0(n6720), .A1(ofifoDataN[506]), .Z(n6350));
Q_AN02 U1902 ( .A0(n6720), .A1(ofifoDataN[505]), .Z(n6349));
Q_AN02 U1903 ( .A0(n6720), .A1(ofifoDataN[504]), .Z(n6348));
Q_AN02 U1904 ( .A0(n6720), .A1(ofifoDataN[503]), .Z(n6347));
Q_AN02 U1905 ( .A0(n6720), .A1(ofifoDataN[502]), .Z(n6346));
Q_AN02 U1906 ( .A0(n6720), .A1(ofifoDataN[501]), .Z(n6345));
Q_AN02 U1907 ( .A0(n6720), .A1(ofifoDataN[500]), .Z(n6344));
Q_AN02 U1908 ( .A0(n6720), .A1(ofifoDataN[499]), .Z(n6343));
Q_AN02 U1909 ( .A0(n6720), .A1(ofifoDataN[498]), .Z(n6342));
Q_AN02 U1910 ( .A0(n6720), .A1(ofifoDataN[497]), .Z(n6341));
Q_AN02 U1911 ( .A0(n6720), .A1(ofifoDataN[496]), .Z(n6340));
Q_AN02 U1912 ( .A0(n6720), .A1(ofifoDataN[495]), .Z(n6339));
Q_AN02 U1913 ( .A0(n6720), .A1(ofifoDataN[494]), .Z(n6338));
Q_AN02 U1914 ( .A0(n6720), .A1(ofifoDataN[493]), .Z(n6337));
Q_AN02 U1915 ( .A0(n6720), .A1(ofifoDataN[492]), .Z(n6336));
Q_AN02 U1916 ( .A0(n6720), .A1(ofifoDataN[491]), .Z(n6335));
Q_AN02 U1917 ( .A0(n6720), .A1(ofifoDataN[490]), .Z(n6334));
Q_AN02 U1918 ( .A0(n6720), .A1(ofifoDataN[489]), .Z(n6333));
Q_AN02 U1919 ( .A0(n6720), .A1(ofifoDataN[488]), .Z(n6332));
Q_AN02 U1920 ( .A0(n6720), .A1(ofifoDataN[487]), .Z(n6331));
Q_AN02 U1921 ( .A0(n6720), .A1(ofifoDataN[486]), .Z(n6330));
Q_AN02 U1922 ( .A0(n6720), .A1(ofifoDataN[485]), .Z(n6329));
Q_AN02 U1923 ( .A0(n6720), .A1(ofifoDataN[484]), .Z(n6328));
Q_AN02 U1924 ( .A0(n6720), .A1(ofifoDataN[483]), .Z(n6327));
Q_AN02 U1925 ( .A0(n6720), .A1(ofifoDataN[482]), .Z(n6326));
Q_AN02 U1926 ( .A0(n6720), .A1(ofifoDataN[481]), .Z(n6325));
Q_AN02 U1927 ( .A0(n6720), .A1(ofifoDataN[480]), .Z(n6324));
Q_AN02 U1928 ( .A0(n6720), .A1(ofifoDataN[479]), .Z(n6323));
Q_AN02 U1929 ( .A0(n6720), .A1(ofifoDataN[478]), .Z(n6322));
Q_AN02 U1930 ( .A0(n6720), .A1(ofifoDataN[477]), .Z(n6321));
Q_AN02 U1931 ( .A0(n6720), .A1(ofifoDataN[476]), .Z(n6320));
Q_AN02 U1932 ( .A0(n6720), .A1(ofifoDataN[475]), .Z(n6319));
Q_AN02 U1933 ( .A0(n6720), .A1(ofifoDataN[474]), .Z(n6318));
Q_AN02 U1934 ( .A0(n6720), .A1(ofifoDataN[473]), .Z(n6317));
Q_AN02 U1935 ( .A0(n6720), .A1(ofifoDataN[472]), .Z(n6316));
Q_AN02 U1936 ( .A0(n6720), .A1(ofifoDataN[471]), .Z(n6315));
Q_AN02 U1937 ( .A0(n6720), .A1(ofifoDataN[470]), .Z(n6314));
Q_AN02 U1938 ( .A0(n6720), .A1(ofifoDataN[469]), .Z(n6313));
Q_AN02 U1939 ( .A0(n6720), .A1(ofifoDataN[468]), .Z(n6312));
Q_AN02 U1940 ( .A0(n6720), .A1(ofifoDataN[467]), .Z(n6311));
Q_AN02 U1941 ( .A0(n6720), .A1(ofifoDataN[466]), .Z(n6310));
Q_AN02 U1942 ( .A0(n6720), .A1(ofifoDataN[465]), .Z(n6309));
Q_AN02 U1943 ( .A0(n6720), .A1(ofifoDataN[464]), .Z(n6308));
Q_AN02 U1944 ( .A0(n6720), .A1(ofifoDataN[463]), .Z(n6307));
Q_AN02 U1945 ( .A0(n6720), .A1(ofifoDataN[462]), .Z(n6306));
Q_AN02 U1946 ( .A0(n6720), .A1(ofifoDataN[461]), .Z(n6305));
Q_AN02 U1947 ( .A0(n6720), .A1(ofifoDataN[460]), .Z(n6304));
Q_AN02 U1948 ( .A0(n6720), .A1(ofifoDataN[459]), .Z(n6303));
Q_AN02 U1949 ( .A0(n6720), .A1(ofifoDataN[458]), .Z(n6302));
Q_AN02 U1950 ( .A0(n6720), .A1(ofifoDataN[457]), .Z(n6301));
Q_AN02 U1951 ( .A0(n6720), .A1(ofifoDataN[456]), .Z(n6300));
Q_AN02 U1952 ( .A0(n6720), .A1(ofifoDataN[455]), .Z(n6299));
Q_AN02 U1953 ( .A0(n6720), .A1(ofifoDataN[454]), .Z(n6298));
Q_AN02 U1954 ( .A0(n6720), .A1(ofifoDataN[453]), .Z(n6297));
Q_AN02 U1955 ( .A0(n6720), .A1(ofifoDataN[452]), .Z(n6296));
Q_AN02 U1956 ( .A0(n6720), .A1(ofifoDataN[451]), .Z(n6295));
Q_AN02 U1957 ( .A0(n6720), .A1(ofifoDataN[450]), .Z(n6294));
Q_AN02 U1958 ( .A0(n6720), .A1(ofifoDataN[449]), .Z(n6293));
Q_AN02 U1959 ( .A0(n6720), .A1(ofifoDataN[448]), .Z(n6292));
Q_AN02 U1960 ( .A0(n6720), .A1(ofifoDataN[447]), .Z(n6291));
Q_AN02 U1961 ( .A0(n6720), .A1(ofifoDataN[446]), .Z(n6290));
Q_AN02 U1962 ( .A0(n6720), .A1(ofifoDataN[445]), .Z(n6289));
Q_AN02 U1963 ( .A0(n6720), .A1(ofifoDataN[444]), .Z(n6288));
Q_AN02 U1964 ( .A0(n6720), .A1(ofifoDataN[443]), .Z(n6287));
Q_AN02 U1965 ( .A0(n6720), .A1(ofifoDataN[442]), .Z(n6286));
Q_AN02 U1966 ( .A0(n6720), .A1(ofifoDataN[441]), .Z(n6285));
Q_AN02 U1967 ( .A0(n6720), .A1(ofifoDataN[440]), .Z(n6284));
Q_AN02 U1968 ( .A0(n6720), .A1(ofifoDataN[439]), .Z(n6283));
Q_AN02 U1969 ( .A0(n6720), .A1(ofifoDataN[438]), .Z(n6282));
Q_AN02 U1970 ( .A0(n6720), .A1(ofifoDataN[437]), .Z(n6281));
Q_AN02 U1971 ( .A0(n6720), .A1(ofifoDataN[436]), .Z(n6280));
Q_AN02 U1972 ( .A0(n6720), .A1(ofifoDataN[435]), .Z(n6279));
Q_AN02 U1973 ( .A0(n6720), .A1(ofifoDataN[434]), .Z(n6278));
Q_AN02 U1974 ( .A0(n6720), .A1(ofifoDataN[433]), .Z(n6277));
Q_AN02 U1975 ( .A0(n6720), .A1(ofifoDataN[432]), .Z(n6276));
Q_AN02 U1976 ( .A0(n6720), .A1(ofifoDataN[431]), .Z(n6275));
Q_AN02 U1977 ( .A0(n6720), .A1(ofifoDataN[430]), .Z(n6274));
Q_AN02 U1978 ( .A0(n6720), .A1(ofifoDataN[429]), .Z(n6273));
Q_AN02 U1979 ( .A0(n6720), .A1(ofifoDataN[428]), .Z(n6272));
Q_AN02 U1980 ( .A0(n6720), .A1(ofifoDataN[427]), .Z(n6271));
Q_AN02 U1981 ( .A0(n6720), .A1(ofifoDataN[426]), .Z(n6270));
Q_AN02 U1982 ( .A0(n6720), .A1(ofifoDataN[425]), .Z(n6269));
Q_AN02 U1983 ( .A0(n6720), .A1(ofifoDataN[424]), .Z(n6268));
Q_AN02 U1984 ( .A0(n6720), .A1(ofifoDataN[423]), .Z(n6267));
Q_AN02 U1985 ( .A0(n6720), .A1(ofifoDataN[422]), .Z(n6266));
Q_AN02 U1986 ( .A0(n6720), .A1(ofifoDataN[421]), .Z(n6265));
Q_AN02 U1987 ( .A0(n6720), .A1(ofifoDataN[420]), .Z(n6264));
Q_AN02 U1988 ( .A0(n6720), .A1(ofifoDataN[419]), .Z(n6263));
Q_AN02 U1989 ( .A0(n6720), .A1(ofifoDataN[418]), .Z(n6262));
Q_AN02 U1990 ( .A0(n6720), .A1(ofifoDataN[417]), .Z(n6261));
Q_AN02 U1991 ( .A0(n6720), .A1(ofifoDataN[416]), .Z(n6260));
Q_AN02 U1992 ( .A0(n6720), .A1(ofifoDataN[415]), .Z(n6259));
Q_AN02 U1993 ( .A0(n6720), .A1(ofifoDataN[414]), .Z(n6258));
Q_AN02 U1994 ( .A0(n6720), .A1(ofifoDataN[413]), .Z(n6257));
Q_AN02 U1995 ( .A0(n6720), .A1(ofifoDataN[412]), .Z(n6256));
Q_AN02 U1996 ( .A0(n6720), .A1(ofifoDataN[411]), .Z(n6255));
Q_AN02 U1997 ( .A0(n6720), .A1(ofifoDataN[410]), .Z(n6254));
Q_AN02 U1998 ( .A0(n6720), .A1(ofifoDataN[409]), .Z(n6253));
Q_AN02 U1999 ( .A0(n6720), .A1(ofifoDataN[408]), .Z(n6252));
Q_AN02 U2000 ( .A0(n6720), .A1(ofifoDataN[407]), .Z(n6251));
Q_AN02 U2001 ( .A0(n6720), .A1(ofifoDataN[406]), .Z(n6250));
Q_AN02 U2002 ( .A0(n6720), .A1(ofifoDataN[405]), .Z(n6249));
Q_AN02 U2003 ( .A0(n6720), .A1(ofifoDataN[404]), .Z(n6248));
Q_AN02 U2004 ( .A0(n6720), .A1(ofifoDataN[403]), .Z(n6247));
Q_AN02 U2005 ( .A0(n6720), .A1(ofifoDataN[402]), .Z(n6246));
Q_AN02 U2006 ( .A0(n6720), .A1(ofifoDataN[401]), .Z(n6245));
Q_AN02 U2007 ( .A0(n6720), .A1(ofifoDataN[400]), .Z(n6244));
Q_AN02 U2008 ( .A0(n6720), .A1(ofifoDataN[399]), .Z(n6243));
Q_AN02 U2009 ( .A0(n6720), .A1(ofifoDataN[398]), .Z(n6242));
Q_AN02 U2010 ( .A0(n6720), .A1(ofifoDataN[397]), .Z(n6241));
Q_AN02 U2011 ( .A0(n6720), .A1(ofifoDataN[396]), .Z(n6240));
Q_AN02 U2012 ( .A0(n6720), .A1(ofifoDataN[395]), .Z(n6239));
Q_AN02 U2013 ( .A0(n6720), .A1(ofifoDataN[394]), .Z(n6238));
Q_AN02 U2014 ( .A0(n6720), .A1(ofifoDataN[393]), .Z(n6237));
Q_AN02 U2015 ( .A0(n6720), .A1(ofifoDataN[392]), .Z(n6236));
Q_AN02 U2016 ( .A0(n6720), .A1(ofifoDataN[391]), .Z(n6235));
Q_AN02 U2017 ( .A0(n6720), .A1(ofifoDataN[390]), .Z(n6234));
Q_AN02 U2018 ( .A0(n6720), .A1(ofifoDataN[389]), .Z(n6233));
Q_AN02 U2019 ( .A0(n6720), .A1(ofifoDataN[388]), .Z(n6232));
Q_AN02 U2020 ( .A0(n6720), .A1(ofifoDataN[387]), .Z(n6231));
Q_AN02 U2021 ( .A0(n6720), .A1(ofifoDataN[386]), .Z(n6230));
Q_AN02 U2022 ( .A0(n6720), .A1(ofifoDataN[385]), .Z(n6229));
Q_AN02 U2023 ( .A0(n6720), .A1(ofifoDataN[384]), .Z(n6228));
Q_AN02 U2024 ( .A0(n6720), .A1(ofifoDataN[383]), .Z(n6227));
Q_AN02 U2025 ( .A0(n6720), .A1(ofifoDataN[382]), .Z(n6226));
Q_AN02 U2026 ( .A0(n6720), .A1(ofifoDataN[381]), .Z(n6225));
Q_AN02 U2027 ( .A0(n6720), .A1(ofifoDataN[380]), .Z(n6224));
Q_AN02 U2028 ( .A0(n6720), .A1(ofifoDataN[379]), .Z(n6223));
Q_AN02 U2029 ( .A0(n6720), .A1(ofifoDataN[378]), .Z(n6222));
Q_AN02 U2030 ( .A0(n6720), .A1(ofifoDataN[377]), .Z(n6221));
Q_AN02 U2031 ( .A0(n6720), .A1(ofifoDataN[376]), .Z(n6220));
Q_AN02 U2032 ( .A0(n6720), .A1(ofifoDataN[375]), .Z(n6219));
Q_AN02 U2033 ( .A0(n6720), .A1(ofifoDataN[374]), .Z(n6218));
Q_AN02 U2034 ( .A0(n6720), .A1(ofifoDataN[373]), .Z(n6217));
Q_AN02 U2035 ( .A0(n6720), .A1(ofifoDataN[372]), .Z(n6216));
Q_AN02 U2036 ( .A0(n6720), .A1(ofifoDataN[371]), .Z(n6215));
Q_AN02 U2037 ( .A0(n6720), .A1(ofifoDataN[370]), .Z(n6214));
Q_AN02 U2038 ( .A0(n6720), .A1(ofifoDataN[369]), .Z(n6213));
Q_AN02 U2039 ( .A0(n6720), .A1(ofifoDataN[368]), .Z(n6212));
Q_AN02 U2040 ( .A0(n6720), .A1(ofifoDataN[367]), .Z(n6211));
Q_AN02 U2041 ( .A0(n6720), .A1(ofifoDataN[366]), .Z(n6210));
Q_AN02 U2042 ( .A0(n6720), .A1(ofifoDataN[365]), .Z(n6209));
Q_AN02 U2043 ( .A0(n6720), .A1(ofifoDataN[364]), .Z(n6208));
Q_AN02 U2044 ( .A0(n6720), .A1(ofifoDataN[363]), .Z(n6207));
Q_AN02 U2045 ( .A0(n6720), .A1(ofifoDataN[362]), .Z(n6206));
Q_AN02 U2046 ( .A0(n6720), .A1(ofifoDataN[361]), .Z(n6205));
Q_AN02 U2047 ( .A0(n6720), .A1(ofifoDataN[360]), .Z(n6204));
Q_AN02 U2048 ( .A0(n6720), .A1(ofifoDataN[359]), .Z(n6203));
Q_AN02 U2049 ( .A0(n6720), .A1(ofifoDataN[358]), .Z(n6202));
Q_AN02 U2050 ( .A0(n6720), .A1(ofifoDataN[357]), .Z(n6201));
Q_AN02 U2051 ( .A0(n6720), .A1(ofifoDataN[356]), .Z(n6200));
Q_AN02 U2052 ( .A0(n6720), .A1(ofifoDataN[355]), .Z(n6199));
Q_AN02 U2053 ( .A0(n6720), .A1(ofifoDataN[354]), .Z(n6198));
Q_AN02 U2054 ( .A0(n6720), .A1(ofifoDataN[353]), .Z(n6197));
Q_AN02 U2055 ( .A0(n6720), .A1(ofifoDataN[352]), .Z(n6196));
Q_AN02 U2056 ( .A0(n6720), .A1(ofifoDataN[351]), .Z(n6195));
Q_AN02 U2057 ( .A0(n6720), .A1(ofifoDataN[350]), .Z(n6194));
Q_AN02 U2058 ( .A0(n6720), .A1(ofifoDataN[349]), .Z(n6193));
Q_AN02 U2059 ( .A0(n6720), .A1(ofifoDataN[348]), .Z(n6192));
Q_AN02 U2060 ( .A0(n6720), .A1(ofifoDataN[347]), .Z(n6191));
Q_AN02 U2061 ( .A0(n6720), .A1(ofifoDataN[346]), .Z(n6190));
Q_AN02 U2062 ( .A0(n6720), .A1(ofifoDataN[345]), .Z(n6189));
Q_AN02 U2063 ( .A0(n6720), .A1(ofifoDataN[344]), .Z(n6188));
Q_AN02 U2064 ( .A0(n6720), .A1(ofifoDataN[343]), .Z(n6187));
Q_AN02 U2065 ( .A0(n6720), .A1(ofifoDataN[342]), .Z(n6186));
Q_AN02 U2066 ( .A0(n6720), .A1(ofifoDataN[341]), .Z(n6185));
Q_AN02 U2067 ( .A0(n6720), .A1(ofifoDataN[340]), .Z(n6184));
Q_AN02 U2068 ( .A0(n6720), .A1(ofifoDataN[339]), .Z(n6183));
Q_AN02 U2069 ( .A0(n6720), .A1(ofifoDataN[338]), .Z(n6182));
Q_AN02 U2070 ( .A0(n6720), .A1(ofifoDataN[337]), .Z(n6181));
Q_AN02 U2071 ( .A0(n6720), .A1(ofifoDataN[336]), .Z(n6180));
Q_AN02 U2072 ( .A0(n6720), .A1(ofifoDataN[335]), .Z(n6179));
Q_AN02 U2073 ( .A0(n6720), .A1(ofifoDataN[334]), .Z(n6178));
Q_AN02 U2074 ( .A0(n6720), .A1(ofifoDataN[333]), .Z(n6177));
Q_AN02 U2075 ( .A0(n6720), .A1(ofifoDataN[332]), .Z(n6176));
Q_AN02 U2076 ( .A0(n6720), .A1(ofifoDataN[331]), .Z(n6175));
Q_AN02 U2077 ( .A0(n6720), .A1(ofifoDataN[330]), .Z(n6174));
Q_AN02 U2078 ( .A0(n6720), .A1(ofifoDataN[329]), .Z(n6173));
Q_AN02 U2079 ( .A0(n6720), .A1(ofifoDataN[328]), .Z(n6172));
Q_AN02 U2080 ( .A0(n6720), .A1(ofifoDataN[327]), .Z(n6171));
Q_AN02 U2081 ( .A0(n6720), .A1(ofifoDataN[326]), .Z(n6170));
Q_AN02 U2082 ( .A0(n6720), .A1(ofifoDataN[325]), .Z(n6169));
Q_AN02 U2083 ( .A0(n6720), .A1(ofifoDataN[324]), .Z(n6168));
Q_AN02 U2084 ( .A0(n6720), .A1(ofifoDataN[323]), .Z(n6167));
Q_AN02 U2085 ( .A0(n6720), .A1(ofifoDataN[322]), .Z(n6166));
Q_AN02 U2086 ( .A0(n6720), .A1(ofifoDataN[321]), .Z(n6165));
Q_AN02 U2087 ( .A0(n6720), .A1(ofifoDataN[320]), .Z(n6164));
Q_AN02 U2088 ( .A0(n6720), .A1(ofifoDataN[319]), .Z(n6163));
Q_AN02 U2089 ( .A0(n6720), .A1(ofifoDataN[318]), .Z(n6162));
Q_AN02 U2090 ( .A0(n6720), .A1(ofifoDataN[317]), .Z(n6161));
Q_AN02 U2091 ( .A0(n6720), .A1(ofifoDataN[316]), .Z(n6160));
Q_AN02 U2092 ( .A0(n6720), .A1(ofifoDataN[315]), .Z(n6159));
Q_AN02 U2093 ( .A0(n6720), .A1(ofifoDataN[314]), .Z(n6158));
Q_AN02 U2094 ( .A0(n6720), .A1(ofifoDataN[313]), .Z(n6157));
Q_AN02 U2095 ( .A0(n6720), .A1(ofifoDataN[312]), .Z(n6156));
Q_AN02 U2096 ( .A0(n6720), .A1(ofifoDataN[311]), .Z(n6155));
Q_AN02 U2097 ( .A0(n6720), .A1(ofifoDataN[310]), .Z(n6154));
Q_AN02 U2098 ( .A0(n6720), .A1(ofifoDataN[309]), .Z(n6153));
Q_AN02 U2099 ( .A0(n6720), .A1(ofifoDataN[308]), .Z(n6152));
Q_AN02 U2100 ( .A0(n6720), .A1(ofifoDataN[307]), .Z(n6151));
Q_AN02 U2101 ( .A0(n6720), .A1(ofifoDataN[306]), .Z(n6150));
Q_AN02 U2102 ( .A0(n6720), .A1(ofifoDataN[305]), .Z(n6149));
Q_AN02 U2103 ( .A0(n6720), .A1(ofifoDataN[304]), .Z(n6148));
Q_AN02 U2104 ( .A0(n6720), .A1(ofifoDataN[303]), .Z(n6147));
Q_AN02 U2105 ( .A0(n6720), .A1(ofifoDataN[302]), .Z(n6146));
Q_AN02 U2106 ( .A0(n6720), .A1(ofifoDataN[301]), .Z(n6145));
Q_AN02 U2107 ( .A0(n6720), .A1(ofifoDataN[300]), .Z(n6144));
Q_AN02 U2108 ( .A0(n6720), .A1(ofifoDataN[299]), .Z(n6143));
Q_AN02 U2109 ( .A0(n6720), .A1(ofifoDataN[298]), .Z(n6142));
Q_AN02 U2110 ( .A0(n6720), .A1(ofifoDataN[297]), .Z(n6141));
Q_AN02 U2111 ( .A0(n6720), .A1(ofifoDataN[296]), .Z(n6140));
Q_AN02 U2112 ( .A0(n6720), .A1(ofifoDataN[295]), .Z(n6139));
Q_AN02 U2113 ( .A0(n6720), .A1(ofifoDataN[294]), .Z(n6138));
Q_AN02 U2114 ( .A0(n6720), .A1(ofifoDataN[293]), .Z(n6137));
Q_AN02 U2115 ( .A0(n6720), .A1(ofifoDataN[292]), .Z(n6136));
Q_AN02 U2116 ( .A0(n6720), .A1(ofifoDataN[291]), .Z(n6135));
Q_AN02 U2117 ( .A0(n6720), .A1(ofifoDataN[290]), .Z(n6134));
Q_AN02 U2118 ( .A0(n6720), .A1(ofifoDataN[289]), .Z(n6133));
Q_AN02 U2119 ( .A0(n6720), .A1(ofifoDataN[288]), .Z(n6132));
Q_AN02 U2120 ( .A0(n6720), .A1(ofifoDataN[287]), .Z(n6131));
Q_AN02 U2121 ( .A0(n6720), .A1(ofifoDataN[286]), .Z(n6130));
Q_AN02 U2122 ( .A0(n6720), .A1(ofifoDataN[285]), .Z(n6129));
Q_AN02 U2123 ( .A0(n6720), .A1(ofifoDataN[284]), .Z(n6128));
Q_AN02 U2124 ( .A0(n6720), .A1(ofifoDataN[283]), .Z(n6127));
Q_AN02 U2125 ( .A0(n6720), .A1(ofifoDataN[282]), .Z(n6126));
Q_AN02 U2126 ( .A0(n6720), .A1(ofifoDataN[281]), .Z(n6125));
Q_AN02 U2127 ( .A0(n6720), .A1(ofifoDataN[280]), .Z(n6124));
Q_AN02 U2128 ( .A0(n6720), .A1(ofifoDataN[279]), .Z(n6123));
Q_AN02 U2129 ( .A0(n6720), .A1(ofifoDataN[278]), .Z(n6122));
Q_AN02 U2130 ( .A0(n6720), .A1(ofifoDataN[277]), .Z(n6121));
Q_AN02 U2131 ( .A0(n6720), .A1(ofifoDataN[276]), .Z(n6120));
Q_AN02 U2132 ( .A0(n6720), .A1(ofifoDataN[275]), .Z(n6119));
Q_AN02 U2133 ( .A0(n6720), .A1(ofifoDataN[274]), .Z(n6118));
Q_AN02 U2134 ( .A0(n6720), .A1(ofifoDataN[273]), .Z(n6117));
Q_AN02 U2135 ( .A0(n6720), .A1(ofifoDataN[272]), .Z(n6116));
Q_AN02 U2136 ( .A0(n6720), .A1(ofifoDataN[271]), .Z(n6115));
Q_AN02 U2137 ( .A0(n6720), .A1(ofifoDataN[270]), .Z(n6114));
Q_AN02 U2138 ( .A0(n6720), .A1(ofifoDataN[269]), .Z(n6113));
Q_AN02 U2139 ( .A0(n6720), .A1(ofifoDataN[268]), .Z(n6112));
Q_AN02 U2140 ( .A0(n6720), .A1(ofifoDataN[267]), .Z(n6111));
Q_AN02 U2141 ( .A0(n6720), .A1(ofifoDataN[266]), .Z(n6110));
Q_AN02 U2142 ( .A0(n6720), .A1(ofifoDataN[265]), .Z(n6109));
Q_AN02 U2143 ( .A0(n6720), .A1(ofifoDataN[264]), .Z(n6108));
Q_AN02 U2144 ( .A0(n6720), .A1(ofifoDataN[263]), .Z(n6107));
Q_AN02 U2145 ( .A0(n6720), .A1(ofifoDataN[262]), .Z(n6106));
Q_AN02 U2146 ( .A0(n6720), .A1(ofifoDataN[261]), .Z(n6105));
Q_AN02 U2147 ( .A0(n6720), .A1(ofifoDataN[260]), .Z(n6104));
Q_AN02 U2148 ( .A0(n6720), .A1(ofifoDataN[259]), .Z(n6103));
Q_AN02 U2149 ( .A0(n6720), .A1(ofifoDataN[258]), .Z(n6102));
Q_AN02 U2150 ( .A0(n6720), .A1(ofifoDataN[257]), .Z(n6101));
Q_AN02 U2151 ( .A0(n6720), .A1(ofifoDataN[256]), .Z(n6100));
Q_AN02 U2152 ( .A0(n6720), .A1(ofifoDataN[255]), .Z(n6099));
Q_AN02 U2153 ( .A0(n6720), .A1(ofifoDataN[254]), .Z(n6098));
Q_AN02 U2154 ( .A0(n6720), .A1(ofifoDataN[253]), .Z(n6097));
Q_AN02 U2155 ( .A0(n6720), .A1(ofifoDataN[252]), .Z(n6096));
Q_AN02 U2156 ( .A0(n6720), .A1(ofifoDataN[251]), .Z(n6095));
Q_AN02 U2157 ( .A0(n6720), .A1(ofifoDataN[250]), .Z(n6094));
Q_AN02 U2158 ( .A0(n6720), .A1(ofifoDataN[249]), .Z(n6093));
Q_AN02 U2159 ( .A0(n6720), .A1(ofifoDataN[248]), .Z(n6092));
Q_AN02 U2160 ( .A0(n6720), .A1(ofifoDataN[247]), .Z(n6091));
Q_AN02 U2161 ( .A0(n6720), .A1(ofifoDataN[246]), .Z(n6090));
Q_AN02 U2162 ( .A0(n6720), .A1(ofifoDataN[245]), .Z(n6089));
Q_AN02 U2163 ( .A0(n6720), .A1(ofifoDataN[244]), .Z(n6088));
Q_AN02 U2164 ( .A0(n6720), .A1(ofifoDataN[243]), .Z(n6087));
Q_AN02 U2165 ( .A0(n6720), .A1(ofifoDataN[242]), .Z(n6086));
Q_AN02 U2166 ( .A0(n6720), .A1(ofifoDataN[241]), .Z(n6085));
Q_AN02 U2167 ( .A0(n6720), .A1(ofifoDataN[240]), .Z(n6084));
Q_AN02 U2168 ( .A0(n6720), .A1(ofifoDataN[239]), .Z(n6083));
Q_AN02 U2169 ( .A0(n6720), .A1(ofifoDataN[238]), .Z(n6082));
Q_AN02 U2170 ( .A0(n6720), .A1(ofifoDataN[237]), .Z(n6081));
Q_AN02 U2171 ( .A0(n6720), .A1(ofifoDataN[236]), .Z(n6080));
Q_AN02 U2172 ( .A0(n6720), .A1(ofifoDataN[235]), .Z(n6079));
Q_AN02 U2173 ( .A0(n6720), .A1(ofifoDataN[234]), .Z(n6078));
Q_AN02 U2174 ( .A0(n6720), .A1(ofifoDataN[233]), .Z(n6077));
Q_AN02 U2175 ( .A0(n6720), .A1(ofifoDataN[232]), .Z(n6076));
Q_AN02 U2176 ( .A0(n6720), .A1(ofifoDataN[231]), .Z(n6075));
Q_AN02 U2177 ( .A0(n6720), .A1(ofifoDataN[230]), .Z(n6074));
Q_AN02 U2178 ( .A0(n6720), .A1(ofifoDataN[229]), .Z(n6073));
Q_AN02 U2179 ( .A0(n6720), .A1(ofifoDataN[228]), .Z(n6072));
Q_AN02 U2180 ( .A0(n6720), .A1(ofifoDataN[227]), .Z(n6071));
Q_AN02 U2181 ( .A0(n6720), .A1(ofifoDataN[226]), .Z(n6070));
Q_AN02 U2182 ( .A0(n6720), .A1(ofifoDataN[225]), .Z(n6069));
Q_AN02 U2183 ( .A0(n6720), .A1(ofifoDataN[224]), .Z(n6068));
Q_AN02 U2184 ( .A0(n6720), .A1(ofifoDataN[223]), .Z(n6067));
Q_AN02 U2185 ( .A0(n6720), .A1(ofifoDataN[222]), .Z(n6066));
Q_AN02 U2186 ( .A0(n6720), .A1(ofifoDataN[221]), .Z(n6065));
Q_AN02 U2187 ( .A0(n6720), .A1(ofifoDataN[220]), .Z(n6064));
Q_AN02 U2188 ( .A0(n6720), .A1(ofifoDataN[219]), .Z(n6063));
Q_AN02 U2189 ( .A0(n6720), .A1(ofifoDataN[218]), .Z(n6062));
Q_AN02 U2190 ( .A0(n6720), .A1(ofifoDataN[217]), .Z(n6061));
Q_AN02 U2191 ( .A0(n6720), .A1(ofifoDataN[216]), .Z(n6060));
Q_AN02 U2192 ( .A0(n6720), .A1(ofifoDataN[215]), .Z(n6059));
Q_AN02 U2193 ( .A0(n6720), .A1(ofifoDataN[214]), .Z(n6058));
Q_AN02 U2194 ( .A0(n6720), .A1(ofifoDataN[213]), .Z(n6057));
Q_AN02 U2195 ( .A0(n6720), .A1(ofifoDataN[212]), .Z(n6056));
Q_AN02 U2196 ( .A0(n6720), .A1(ofifoDataN[211]), .Z(n6055));
Q_AN02 U2197 ( .A0(n6720), .A1(ofifoDataN[210]), .Z(n6054));
Q_AN02 U2198 ( .A0(n6720), .A1(ofifoDataN[209]), .Z(n6053));
Q_AN02 U2199 ( .A0(n6720), .A1(ofifoDataN[208]), .Z(n6052));
Q_AN02 U2200 ( .A0(n6720), .A1(ofifoDataN[207]), .Z(n6051));
Q_AN02 U2201 ( .A0(n6720), .A1(ofifoDataN[206]), .Z(n6050));
Q_AN02 U2202 ( .A0(n6720), .A1(ofifoDataN[205]), .Z(n6049));
Q_AN02 U2203 ( .A0(n6720), .A1(ofifoDataN[204]), .Z(n6048));
Q_AN02 U2204 ( .A0(n6720), .A1(ofifoDataN[203]), .Z(n6047));
Q_AN02 U2205 ( .A0(n6720), .A1(ofifoDataN[202]), .Z(n6046));
Q_AN02 U2206 ( .A0(n6720), .A1(ofifoDataN[201]), .Z(n6045));
Q_AN02 U2207 ( .A0(n6720), .A1(ofifoDataN[200]), .Z(n6044));
Q_AN02 U2208 ( .A0(n6720), .A1(ofifoDataN[199]), .Z(n6043));
Q_AN02 U2209 ( .A0(n6720), .A1(ofifoDataN[198]), .Z(n6042));
Q_AN02 U2210 ( .A0(n6720), .A1(ofifoDataN[197]), .Z(n6041));
Q_AN02 U2211 ( .A0(n6720), .A1(ofifoDataN[196]), .Z(n6040));
Q_AN02 U2212 ( .A0(n6720), .A1(ofifoDataN[195]), .Z(n6039));
Q_AN02 U2213 ( .A0(n6720), .A1(ofifoDataN[194]), .Z(n6038));
Q_AN02 U2214 ( .A0(n6720), .A1(ofifoDataN[193]), .Z(n6037));
Q_AN02 U2215 ( .A0(n6720), .A1(ofifoDataN[192]), .Z(n6036));
Q_AN02 U2216 ( .A0(n6720), .A1(ofifoDataN[191]), .Z(n6035));
Q_AN02 U2217 ( .A0(n6720), .A1(ofifoDataN[190]), .Z(n6034));
Q_AN02 U2218 ( .A0(n6720), .A1(ofifoDataN[189]), .Z(n6033));
Q_AN02 U2219 ( .A0(n6720), .A1(ofifoDataN[188]), .Z(n6032));
Q_AN02 U2220 ( .A0(n6720), .A1(ofifoDataN[187]), .Z(n6031));
Q_AN02 U2221 ( .A0(n6720), .A1(ofifoDataN[186]), .Z(n6030));
Q_AN02 U2222 ( .A0(n6720), .A1(ofifoDataN[185]), .Z(n6029));
Q_AN02 U2223 ( .A0(n6720), .A1(ofifoDataN[184]), .Z(n6028));
Q_AN02 U2224 ( .A0(n6720), .A1(ofifoDataN[183]), .Z(n6027));
Q_AN02 U2225 ( .A0(n6720), .A1(ofifoDataN[182]), .Z(n6026));
Q_AN02 U2226 ( .A0(n6720), .A1(ofifoDataN[181]), .Z(n6025));
Q_AN02 U2227 ( .A0(n6720), .A1(ofifoDataN[180]), .Z(n6024));
Q_AN02 U2228 ( .A0(n6720), .A1(ofifoDataN[179]), .Z(n6023));
Q_AN02 U2229 ( .A0(n6720), .A1(ofifoDataN[178]), .Z(n6022));
Q_AN02 U2230 ( .A0(n6720), .A1(ofifoDataN[177]), .Z(n6021));
Q_AN02 U2231 ( .A0(n6720), .A1(ofifoDataN[176]), .Z(n6020));
Q_AN02 U2232 ( .A0(n6720), .A1(ofifoDataN[175]), .Z(n6019));
Q_AN02 U2233 ( .A0(n6720), .A1(ofifoDataN[174]), .Z(n6018));
Q_AN02 U2234 ( .A0(n6720), .A1(ofifoDataN[173]), .Z(n6017));
Q_AN02 U2235 ( .A0(n6720), .A1(ofifoDataN[172]), .Z(n6016));
Q_AN02 U2236 ( .A0(n6720), .A1(ofifoDataN[171]), .Z(n6015));
Q_AN02 U2237 ( .A0(n6720), .A1(ofifoDataN[170]), .Z(n6014));
Q_AN02 U2238 ( .A0(n6720), .A1(ofifoDataN[169]), .Z(n6013));
Q_AN02 U2239 ( .A0(n6720), .A1(ofifoDataN[168]), .Z(n6012));
Q_AN02 U2240 ( .A0(n6720), .A1(ofifoDataN[167]), .Z(n6011));
Q_AN02 U2241 ( .A0(n6720), .A1(ofifoDataN[166]), .Z(n6010));
Q_AN02 U2242 ( .A0(n6720), .A1(ofifoDataN[165]), .Z(n6009));
Q_AN02 U2243 ( .A0(n6720), .A1(ofifoDataN[164]), .Z(n6008));
Q_AN02 U2244 ( .A0(n6720), .A1(ofifoDataN[163]), .Z(n6007));
Q_AN02 U2245 ( .A0(n6720), .A1(ofifoDataN[162]), .Z(n6006));
Q_AN02 U2246 ( .A0(n6720), .A1(ofifoDataN[161]), .Z(n6005));
Q_AN02 U2247 ( .A0(n6720), .A1(ofifoDataN[160]), .Z(n6004));
Q_AN02 U2248 ( .A0(n6720), .A1(ofifoDataN[159]), .Z(n6003));
Q_AN02 U2249 ( .A0(n6720), .A1(ofifoDataN[158]), .Z(n6002));
Q_AN02 U2250 ( .A0(n6720), .A1(ofifoDataN[157]), .Z(n6001));
Q_AN02 U2251 ( .A0(n6720), .A1(ofifoDataN[156]), .Z(n6000));
Q_AN02 U2252 ( .A0(n6720), .A1(ofifoDataN[155]), .Z(n5999));
Q_AN02 U2253 ( .A0(n6720), .A1(ofifoDataN[154]), .Z(n5998));
Q_AN02 U2254 ( .A0(n6720), .A1(ofifoDataN[153]), .Z(n5997));
Q_AN02 U2255 ( .A0(n6720), .A1(ofifoDataN[152]), .Z(n5996));
Q_AN02 U2256 ( .A0(n6720), .A1(ofifoDataN[151]), .Z(n5995));
Q_AN02 U2257 ( .A0(n6720), .A1(ofifoDataN[150]), .Z(n5994));
Q_AN02 U2258 ( .A0(n6720), .A1(ofifoDataN[149]), .Z(n5993));
Q_AN02 U2259 ( .A0(n6720), .A1(ofifoDataN[148]), .Z(n5992));
Q_AN02 U2260 ( .A0(n6720), .A1(ofifoDataN[147]), .Z(n5991));
Q_AN02 U2261 ( .A0(n6720), .A1(ofifoDataN[146]), .Z(n5990));
Q_AN02 U2262 ( .A0(n6720), .A1(ofifoDataN[145]), .Z(n5989));
Q_AN02 U2263 ( .A0(n6720), .A1(ofifoDataN[144]), .Z(n5988));
Q_AN02 U2264 ( .A0(n6720), .A1(ofifoDataN[143]), .Z(n5987));
Q_AN02 U2265 ( .A0(n6720), .A1(ofifoDataN[142]), .Z(n5986));
Q_AN02 U2266 ( .A0(n6720), .A1(ofifoDataN[141]), .Z(n5985));
Q_AN02 U2267 ( .A0(n6720), .A1(ofifoDataN[140]), .Z(n5984));
Q_AN02 U2268 ( .A0(n6720), .A1(ofifoDataN[139]), .Z(n5983));
Q_AN02 U2269 ( .A0(n6720), .A1(ofifoDataN[138]), .Z(n5982));
Q_AN02 U2270 ( .A0(n6720), .A1(ofifoDataN[137]), .Z(n5981));
Q_AN02 U2271 ( .A0(n6720), .A1(ofifoDataN[136]), .Z(n5980));
Q_AN02 U2272 ( .A0(n6720), .A1(ofifoDataN[135]), .Z(n5979));
Q_AN02 U2273 ( .A0(n6720), .A1(ofifoDataN[134]), .Z(n5978));
Q_AN02 U2274 ( .A0(n6720), .A1(ofifoDataN[133]), .Z(n5977));
Q_AN02 U2275 ( .A0(n6720), .A1(ofifoDataN[132]), .Z(n5976));
Q_AN02 U2276 ( .A0(n6720), .A1(ofifoDataN[131]), .Z(n5975));
Q_AN02 U2277 ( .A0(n6720), .A1(ofifoDataN[130]), .Z(n5974));
Q_AN02 U2278 ( .A0(n6720), .A1(ofifoDataN[129]), .Z(n5973));
Q_AN02 U2279 ( .A0(n6720), .A1(ofifoDataN[128]), .Z(n5972));
Q_AN02 U2280 ( .A0(n6720), .A1(ofifoDataN[127]), .Z(n5971));
Q_AN02 U2281 ( .A0(n6720), .A1(ofifoDataN[126]), .Z(n5970));
Q_AN02 U2282 ( .A0(n6720), .A1(ofifoDataN[125]), .Z(n5969));
Q_AN02 U2283 ( .A0(n6720), .A1(ofifoDataN[124]), .Z(n5968));
Q_AN02 U2284 ( .A0(n6720), .A1(ofifoDataN[123]), .Z(n5967));
Q_AN02 U2285 ( .A0(n6720), .A1(ofifoDataN[122]), .Z(n5966));
Q_AN02 U2286 ( .A0(n6720), .A1(ofifoDataN[121]), .Z(n5965));
Q_AN02 U2287 ( .A0(n6720), .A1(ofifoDataN[120]), .Z(n5964));
Q_AN02 U2288 ( .A0(n6720), .A1(ofifoDataN[119]), .Z(n5963));
Q_AN02 U2289 ( .A0(n6720), .A1(ofifoDataN[118]), .Z(n5962));
Q_AN02 U2290 ( .A0(n6720), .A1(ofifoDataN[117]), .Z(n5961));
Q_AN02 U2291 ( .A0(n6720), .A1(ofifoDataN[116]), .Z(n5960));
Q_AN02 U2292 ( .A0(n6720), .A1(ofifoDataN[115]), .Z(n5959));
Q_AN02 U2293 ( .A0(n6720), .A1(ofifoDataN[114]), .Z(n5958));
Q_AN02 U2294 ( .A0(n6720), .A1(ofifoDataN[113]), .Z(n5957));
Q_AN02 U2295 ( .A0(n6720), .A1(ofifoDataN[112]), .Z(n5956));
Q_AN02 U2296 ( .A0(n6720), .A1(ofifoDataN[111]), .Z(n5955));
Q_AN02 U2297 ( .A0(n6720), .A1(ofifoDataN[110]), .Z(n5954));
Q_AN02 U2298 ( .A0(n6720), .A1(ofifoDataN[109]), .Z(n5953));
Q_AN02 U2299 ( .A0(n6720), .A1(ofifoDataN[108]), .Z(n5952));
Q_AN02 U2300 ( .A0(n6720), .A1(ofifoDataN[107]), .Z(n5951));
Q_AN02 U2301 ( .A0(n6720), .A1(ofifoDataN[106]), .Z(n5950));
Q_AN02 U2302 ( .A0(n6720), .A1(ofifoDataN[105]), .Z(n5949));
Q_AN02 U2303 ( .A0(n6720), .A1(ofifoDataN[104]), .Z(n5948));
Q_AN02 U2304 ( .A0(n6720), .A1(ofifoDataN[103]), .Z(n5947));
Q_AN02 U2305 ( .A0(n6720), .A1(ofifoDataN[102]), .Z(n5946));
Q_AN02 U2306 ( .A0(n6720), .A1(ofifoDataN[101]), .Z(n5945));
Q_AN02 U2307 ( .A0(n6720), .A1(ofifoDataN[100]), .Z(n5944));
Q_AN02 U2308 ( .A0(n6720), .A1(ofifoDataN[99]), .Z(n5943));
Q_AN02 U2309 ( .A0(n6720), .A1(ofifoDataN[98]), .Z(n5942));
Q_AN02 U2310 ( .A0(n6720), .A1(ofifoDataN[97]), .Z(n5941));
Q_AN02 U2311 ( .A0(n6720), .A1(ofifoDataN[96]), .Z(n5940));
Q_AN02 U2312 ( .A0(n6720), .A1(ofifoDataN[95]), .Z(n5939));
Q_AN02 U2313 ( .A0(n6720), .A1(ofifoDataN[94]), .Z(n5938));
Q_AN02 U2314 ( .A0(n6720), .A1(ofifoDataN[93]), .Z(n5937));
Q_AN02 U2315 ( .A0(n6720), .A1(ofifoDataN[92]), .Z(n5936));
Q_AN02 U2316 ( .A0(n6720), .A1(ofifoDataN[91]), .Z(n5935));
Q_AN02 U2317 ( .A0(n6720), .A1(ofifoDataN[90]), .Z(n5934));
Q_AN02 U2318 ( .A0(n6720), .A1(ofifoDataN[89]), .Z(n5933));
Q_AN02 U2319 ( .A0(n6720), .A1(ofifoDataN[88]), .Z(n5932));
Q_AN02 U2320 ( .A0(n6720), .A1(ofifoDataN[87]), .Z(n5931));
Q_AN02 U2321 ( .A0(n6720), .A1(ofifoDataN[86]), .Z(n5930));
Q_AN02 U2322 ( .A0(n6720), .A1(ofifoDataN[85]), .Z(n5929));
Q_AN02 U2323 ( .A0(n6720), .A1(ofifoDataN[84]), .Z(n5928));
Q_AN02 U2324 ( .A0(n6720), .A1(ofifoDataN[83]), .Z(n5927));
Q_AN02 U2325 ( .A0(n6720), .A1(ofifoDataN[82]), .Z(n5926));
Q_AN02 U2326 ( .A0(n6720), .A1(ofifoDataN[81]), .Z(n5925));
Q_AN02 U2327 ( .A0(n6720), .A1(ofifoDataN[80]), .Z(n5924));
Q_AN02 U2328 ( .A0(n6720), .A1(ofifoDataN[79]), .Z(n5923));
Q_AN02 U2329 ( .A0(n6720), .A1(ofifoDataN[78]), .Z(n5922));
Q_AN02 U2330 ( .A0(n6720), .A1(ofifoDataN[77]), .Z(n5921));
Q_AN02 U2331 ( .A0(n6720), .A1(ofifoDataN[76]), .Z(n5920));
Q_AN02 U2332 ( .A0(n6720), .A1(ofifoDataN[75]), .Z(n5919));
Q_AN02 U2333 ( .A0(n6720), .A1(ofifoDataN[74]), .Z(n5918));
Q_AN02 U2334 ( .A0(n6720), .A1(ofifoDataN[73]), .Z(n5917));
Q_AN02 U2335 ( .A0(n6720), .A1(ofifoDataN[72]), .Z(n5916));
Q_AN02 U2336 ( .A0(n6720), .A1(ofifoDataN[71]), .Z(n5915));
Q_AN02 U2337 ( .A0(n6720), .A1(ofifoDataN[70]), .Z(n5914));
Q_AN02 U2338 ( .A0(n6720), .A1(ofifoDataN[69]), .Z(n5913));
Q_AN02 U2339 ( .A0(n6720), .A1(ofifoDataN[68]), .Z(n5912));
Q_AN02 U2340 ( .A0(n6720), .A1(ofifoDataN[67]), .Z(n5911));
Q_AN02 U2341 ( .A0(n6720), .A1(ofifoDataN[66]), .Z(n5910));
Q_AN02 U2342 ( .A0(n6720), .A1(ofifoDataN[65]), .Z(n5909));
Q_AN02 U2343 ( .A0(n6720), .A1(ofifoDataN[64]), .Z(n5908));
Q_AN02 U2344 ( .A0(n6720), .A1(ofifoDataN[63]), .Z(n5907));
Q_AN02 U2345 ( .A0(n6720), .A1(ofifoDataN[62]), .Z(n5906));
Q_AN02 U2346 ( .A0(n6720), .A1(ofifoDataN[61]), .Z(n5905));
Q_AN02 U2347 ( .A0(n6720), .A1(ofifoDataN[60]), .Z(n5904));
Q_AN02 U2348 ( .A0(n6720), .A1(ofifoDataN[59]), .Z(n5903));
Q_AN02 U2349 ( .A0(n6720), .A1(ofifoDataN[58]), .Z(n5902));
Q_AN02 U2350 ( .A0(n6720), .A1(ofifoDataN[57]), .Z(n5901));
Q_AN02 U2351 ( .A0(n6720), .A1(ofifoDataN[56]), .Z(n5900));
Q_AN02 U2352 ( .A0(n6720), .A1(ofifoDataN[55]), .Z(n5899));
Q_AN02 U2353 ( .A0(n6720), .A1(ofifoDataN[54]), .Z(n5898));
Q_AN02 U2354 ( .A0(n6720), .A1(ofifoDataN[53]), .Z(n5897));
Q_AN02 U2355 ( .A0(n6720), .A1(ofifoDataN[52]), .Z(n5896));
Q_AN02 U2356 ( .A0(n6720), .A1(ofifoDataN[51]), .Z(n5895));
Q_AN02 U2357 ( .A0(n6720), .A1(ofifoDataN[50]), .Z(n5894));
Q_AN02 U2358 ( .A0(n6720), .A1(ofifoDataN[49]), .Z(n5893));
Q_AN02 U2359 ( .A0(n6720), .A1(ofifoDataN[48]), .Z(n5892));
Q_AN02 U2360 ( .A0(n6720), .A1(ofifoDataN[47]), .Z(n5891));
Q_AN02 U2361 ( .A0(n6720), .A1(ofifoDataN[46]), .Z(n5890));
Q_AN02 U2362 ( .A0(n6720), .A1(ofifoDataN[45]), .Z(n5889));
Q_AN02 U2363 ( .A0(n6720), .A1(ofifoDataN[44]), .Z(n5888));
Q_AN02 U2364 ( .A0(n6720), .A1(ofifoDataN[43]), .Z(n5887));
Q_AN02 U2365 ( .A0(n6720), .A1(ofifoDataN[42]), .Z(n5886));
Q_AN02 U2366 ( .A0(n6720), .A1(ofifoDataN[41]), .Z(n5885));
Q_AN02 U2367 ( .A0(n6720), .A1(ofifoDataN[40]), .Z(n5884));
Q_AN02 U2368 ( .A0(n6720), .A1(ofifoDataN[39]), .Z(n5883));
Q_AN02 U2369 ( .A0(n6720), .A1(ofifoDataN[38]), .Z(n5882));
Q_AN02 U2370 ( .A0(n6720), .A1(ofifoDataN[37]), .Z(n5881));
Q_AN02 U2371 ( .A0(n6720), .A1(ofifoDataN[36]), .Z(n5880));
Q_AN02 U2372 ( .A0(n6720), .A1(ofifoDataN[35]), .Z(n5879));
Q_AN02 U2373 ( .A0(n6720), .A1(ofifoDataN[34]), .Z(n5878));
Q_AN02 U2374 ( .A0(n6720), .A1(ofifoDataN[33]), .Z(n5877));
Q_AN02 U2375 ( .A0(n6720), .A1(ofifoDataN[32]), .Z(n5876));
Q_AN02 U2376 ( .A0(n6720), .A1(ofifoDataN[31]), .Z(n5875));
Q_AN02 U2377 ( .A0(n6720), .A1(ofifoDataN[30]), .Z(n5874));
Q_AN02 U2378 ( .A0(n6720), .A1(ofifoDataN[29]), .Z(n5873));
Q_AN02 U2379 ( .A0(n6720), .A1(ofifoDataN[28]), .Z(n5872));
Q_AN02 U2380 ( .A0(n6720), .A1(ofifoDataN[27]), .Z(n5871));
Q_AN02 U2381 ( .A0(n6720), .A1(ofifoDataN[26]), .Z(n5870));
Q_AN02 U2382 ( .A0(n6720), .A1(ofifoDataN[25]), .Z(n5869));
Q_AN02 U2383 ( .A0(n6720), .A1(ofifoDataN[24]), .Z(n5868));
Q_AN02 U2384 ( .A0(n6720), .A1(ofifoDataN[23]), .Z(n5867));
Q_AN02 U2385 ( .A0(n6720), .A1(ofifoDataN[22]), .Z(n5866));
Q_AN02 U2386 ( .A0(n6720), .A1(ofifoDataN[21]), .Z(n5865));
Q_AN02 U2387 ( .A0(n6720), .A1(ofifoDataN[20]), .Z(n5864));
Q_AN02 U2388 ( .A0(n6720), .A1(ofifoDataN[19]), .Z(n5863));
Q_AN02 U2389 ( .A0(n6720), .A1(ofifoDataN[18]), .Z(n5862));
Q_AN02 U2390 ( .A0(n6720), .A1(ofifoDataN[17]), .Z(n5861));
Q_AN02 U2391 ( .A0(n6720), .A1(ofifoDataN[16]), .Z(n5860));
Q_AN02 U2392 ( .A0(n6720), .A1(ofifoDataN[15]), .Z(n5859));
Q_AN02 U2393 ( .A0(n6720), .A1(ofifoDataN[14]), .Z(n5858));
Q_AN02 U2394 ( .A0(n6720), .A1(ofifoDataN[13]), .Z(n5857));
Q_AN02 U2395 ( .A0(n6720), .A1(ofifoDataN[12]), .Z(n5856));
Q_AN02 U2396 ( .A0(n6720), .A1(ofifoDataN[11]), .Z(n5855));
Q_AN02 U2397 ( .A0(n6720), .A1(ofifoDataN[10]), .Z(n5854));
Q_AN02 U2398 ( .A0(n6720), .A1(ofifoDataN[9]), .Z(n5853));
Q_AN02 U2399 ( .A0(n6720), .A1(ofifoDataN[8]), .Z(n5852));
Q_AN02 U2400 ( .A0(n6720), .A1(ofifoDataN[7]), .Z(n5851));
Q_AN02 U2401 ( .A0(n6720), .A1(ofifoDataN[6]), .Z(n5850));
Q_AN02 U2402 ( .A0(n6720), .A1(ofifoDataN[5]), .Z(n5849));
Q_AN02 U2403 ( .A0(n6720), .A1(ofifoDataN[4]), .Z(n5848));
Q_AN02 U2404 ( .A0(n6720), .A1(ofifoDataN[3]), .Z(n5847));
Q_AN02 U2405 ( .A0(n6720), .A1(ofifoDataN[2]), .Z(n5846));
Q_AN02 U2406 ( .A0(n6720), .A1(ofifoDataN[1]), .Z(n5845));
Q_AN02 U2407 ( .A0(n6720), .A1(ofifoDataN[0]), .Z(n5844));
Q_AN02 U2408 ( .A0(n6720), .A1(oFillN[4]), .Z(n5843));
Q_AN02 U2409 ( .A0(n6720), .A1(oFillN[3]), .Z(n5842));
Q_AN02 U2410 ( .A0(n6720), .A1(oFillN[2]), .Z(n5841));
Q_AN02 U2411 ( .A0(n6720), .A1(oFillN[1]), .Z(n5840));
Q_AN02 U2412 ( .A0(n6720), .A1(oFillN[0]), .Z(n5839));
Q_AN02 U2413 ( .A0(n6720), .A1(ofifoWptrN[14]), .Z(n5838));
Q_AN02 U2414 ( .A0(n6720), .A1(ofifoWptrN[13]), .Z(n5837));
Q_AN02 U2415 ( .A0(n6720), .A1(ofifoWptrN[12]), .Z(n5836));
Q_AN02 U2416 ( .A0(n6720), .A1(ofifoWptrN[11]), .Z(n5835));
Q_AN02 U2417 ( .A0(n6720), .A1(ofifoWptrN[10]), .Z(n5834));
Q_AN02 U2418 ( .A0(n6720), .A1(ofifoWptrN[9]), .Z(n5833));
Q_AN02 U2419 ( .A0(n6720), .A1(ofifoWptrN[8]), .Z(n5832));
Q_AN02 U2420 ( .A0(n6720), .A1(ofifoWptrN[7]), .Z(n5831));
Q_AN02 U2421 ( .A0(n6720), .A1(ofifoWptrN[6]), .Z(n5830));
Q_AN02 U2422 ( .A0(n6720), .A1(ofifoWptrN[5]), .Z(n5829));
Q_AN02 U2423 ( .A0(n6720), .A1(ofifoWptrN[4]), .Z(n5828));
Q_AN02 U2424 ( .A0(n6720), .A1(ofifoWptrN[3]), .Z(n5827));
Q_AN02 U2425 ( .A0(n6720), .A1(ofifoWptrN[2]), .Z(n5826));
Q_AN02 U2426 ( .A0(n6720), .A1(ofifoWptrN[1]), .Z(n5825));
Q_AN02 U2427 ( .A0(n6720), .A1(ofifoWptrN[0]), .Z(n5824));
Q_INV U2428 ( .A(n5822), .Z(n5811));
Q_OA21 U2429 ( .A0(n5811), .A1(n5823), .B0(n6720), .Z(n5810));
Q_INV U2430 ( .A(n5821), .Z(n5806));
Q_NR02 U2431 ( .A0(xc_top.GFReset), .A1(n5821), .Z(n5809));
Q_AN02 U2432 ( .A0(n5809), .A1(n3683), .Z(n5808));
Q_AN02 U2433 ( .A0(n6720), .A1(n5822), .Z(n5819));
Q_AN03 U2434 ( .A0(n5822), .A1(n5816), .A2(n6720), .Z(n5817));
Q_OR02 U2435 ( .A0(n5817), .A1(xc_top.GFReset), .Z(n5807));
Q_AN03 U2436 ( .A0(n5822), .A1(n3699), .A2(n6720), .Z(n5818));
Q_INV U2437 ( .A(n5823), .Z(n5815));
Q_NR02 U2438 ( .A0(n5821), .A1(n3683), .Z(n5813));
Q_AN02 U2439 ( .A0(n5806), .A1(n3683), .Z(n5812));
Q_MX02 U2440 ( .S(n5819), .A0(argLen[0]), .A1(n4424), .Z(n5805));
Q_FDP0UA U2441 ( .D(n5805), .QTFCLK( ), .Q(argLen[0]));
Q_MX02 U2442 ( .S(n5819), .A0(argLen[1]), .A1(n4425), .Z(n5804));
Q_FDP0UA U2443 ( .D(n5804), .QTFCLK( ), .Q(argLen[1]));
Q_MX02 U2444 ( .S(n5819), .A0(argLen[2]), .A1(n4426), .Z(n5803));
Q_FDP0UA U2445 ( .D(n5803), .QTFCLK( ), .Q(argLen[2]));
Q_MX02 U2446 ( .S(n5819), .A0(argLen[3]), .A1(n4427), .Z(n5802));
Q_FDP0UA U2447 ( .D(n5802), .QTFCLK( ), .Q(argLen[3]));
Q_MX02 U2448 ( .S(n5819), .A0(argLen[4]), .A1(n4428), .Z(n5801));
Q_FDP0UA U2449 ( .D(n5801), .QTFCLK( ), .Q(argLen[4]));
Q_MX02 U2450 ( .S(n5819), .A0(argLen[5]), .A1(n4429), .Z(n5800));
Q_FDP0UA U2451 ( .D(n5800), .QTFCLK( ), .Q(argLen[5]));
Q_MX02 U2452 ( .S(n5819), .A0(argLen[6]), .A1(n4430), .Z(n5799));
Q_FDP0UA U2453 ( .D(n5799), .QTFCLK( ), .Q(argLen[6]));
Q_MX02 U2454 ( .S(n5819), .A0(argLen[7]), .A1(n4431), .Z(n5798));
Q_FDP0UA U2455 ( .D(n5798), .QTFCLK( ), .Q(argLen[7]));
Q_MX02 U2456 ( .S(n5819), .A0(argLen[8]), .A1(n4432), .Z(n5797));
Q_FDP0UA U2457 ( .D(n5797), .QTFCLK( ), .Q(argLen[8]));
Q_MX02 U2458 ( .S(n5819), .A0(argLen[9]), .A1(n4433), .Z(n5796));
Q_FDP0UA U2459 ( .D(n5796), .QTFCLK( ), .Q(argLen[9]));
Q_MX02 U2460 ( .S(n5819), .A0(argLen[10]), .A1(n4434), .Z(n5795));
Q_FDP0UA U2461 ( .D(n5795), .QTFCLK( ), .Q(argLen[10]));
Q_MX02 U2462 ( .S(n5819), .A0(argLen[11]), .A1(n4435), .Z(n5794));
Q_FDP0UA U2463 ( .D(n5794), .QTFCLK( ), .Q(argLen[11]));
Q_FDP0UA U2464 ( .D(n5692), .QTFCLK( ), .Q(wLen[0]));
Q_FDP0UA U2465 ( .D(n5694), .QTFCLK( ), .Q(wLen[1]));
Q_FDP0UA U2466 ( .D(n5696), .QTFCLK( ), .Q(wLen[2]));
Q_FDP0UA U2467 ( .D(n5698), .QTFCLK( ), .Q(wLen[3]));
Q_FDP0UA U2468 ( .D(n5700), .QTFCLK( ), .Q(wLen[4]));
Q_FDP0UA U2469 ( .D(n5702), .QTFCLK( ), .Q(wLen[5]));
Q_FDP0UA U2470 ( .D(n5704), .QTFCLK( ), .Q(wLen[6]));
Q_FDP0UA U2471 ( .D(n5706), .QTFCLK( ), .Q(wLen[7]));
Q_FDP0UA U2472 ( .D(n5708), .QTFCLK( ), .Q(wLen[8]));
Q_FDP0UA U2473 ( .D(n5710), .QTFCLK( ), .Q(wLen[9]));
Q_FDP0UA U2474 ( .D(n5712), .QTFCLK( ), .Q(wLen[10]));
Q_FDP0UA U2475 ( .D(n5714), .QTFCLK( ), .Q(wLen[11]));
Q_FDP0UA U2476 ( .D(n5716), .QTFCLK( ), .Q(wLen[12]));
Q_FDP0UA U2477 ( .D(n5718), .QTFCLK( ), .Q(wLen[13]));
Q_FDP0UA U2478 ( .D(n5720), .QTFCLK( ), .Q(wLen[14]));
Q_FDP0UA U2479 ( .D(n5722), .QTFCLK( ), .Q(wLen[15]));
Q_FDP0UA U2480 ( .D(n5724), .QTFCLK( ), .Q(wLen[16]));
Q_FDP0UA U2481 ( .D(n5726), .QTFCLK( ), .Q(wLen[17]));
Q_FDP0UA U2482 ( .D(n5728), .QTFCLK( ), .Q(wLen[18]));
Q_FDP0UA U2483 ( .D(n4559), .QTFCLK( ), .Q(writeLen[0]));
Q_FDP0UA U2484 ( .D(n4561), .QTFCLK( ), .Q(writeLen[1]));
Q_FDP0UA U2485 ( .D(n4563), .QTFCLK( ), .Q(writeLen[2]));
Q_FDP0UA U2486 ( .D(n4565), .QTFCLK( ), .Q(writeLen[3]));
Q_FDP0UA U2487 ( .D(n4567), .QTFCLK( ), .Q(writeLen[4]));
Q_FDP0UA U2488 ( .D(n4569), .QTFCLK( ), .Q(writeLen[5]));
Q_MX02 U2489 ( .S(n5810), .A0(n4570), .A1(wrtCnt[0]), .Z(n5793));
Q_FDP0UA U2490 ( .D(n5793), .QTFCLK( ), .Q(wrtCnt[0]));
Q_MX02 U2491 ( .S(n5810), .A0(n4571), .A1(wrtCnt[1]), .Z(n5792));
Q_FDP0UA U2492 ( .D(n5792), .QTFCLK( ), .Q(wrtCnt[1]));
Q_MX02 U2493 ( .S(n5810), .A0(n4572), .A1(wrtCnt[2]), .Z(n5791));
Q_FDP0UA U2494 ( .D(n5791), .QTFCLK( ), .Q(wrtCnt[2]));
Q_MX02 U2495 ( .S(n5810), .A0(n4573), .A1(wrtCnt[3]), .Z(n5790));
Q_FDP0UA U2496 ( .D(n5790), .QTFCLK( ), .Q(wrtCnt[3]));
Q_MX02 U2497 ( .S(n5810), .A0(n4574), .A1(wrtCnt[4]), .Z(n5789));
Q_FDP0UA U2498 ( .D(n5789), .QTFCLK( ), .Q(wrtCnt[4]));
Q_MX02 U2499 ( .S(n5810), .A0(n4575), .A1(wrtCnt[5]), .Z(n5788));
Q_FDP0UA U2500 ( .D(n5788), .QTFCLK( ), .Q(wrtCnt[5]));
Q_MX02 U2501 ( .S(n5810), .A0(n4576), .A1(wrtCnt[6]), .Z(n5787));
Q_FDP0UA U2502 ( .D(n5787), .QTFCLK( ), .Q(wrtCnt[6]));
Q_MX02 U2503 ( .S(n5810), .A0(n4577), .A1(wrtCnt[7]), .Z(n5786));
Q_FDP0UA U2504 ( .D(n5786), .QTFCLK( ), .Q(wrtCnt[7]));
Q_MX02 U2505 ( .S(n5810), .A0(n4578), .A1(wrtCnt[8]), .Z(n5785));
Q_FDP0UA U2506 ( .D(n5785), .QTFCLK( ), .Q(wrtCnt[8]));
Q_MX02 U2507 ( .S(n5810), .A0(n4579), .A1(wrtCnt[9]), .Z(n5784));
Q_FDP0UA U2508 ( .D(n5784), .QTFCLK( ), .Q(wrtCnt[9]));
Q_MX02 U2509 ( .S(n5810), .A0(n4580), .A1(wrtCnt[10]), .Z(n5783));
Q_FDP0UA U2510 ( .D(n5783), .QTFCLK( ), .Q(wrtCnt[10]));
Q_MX02 U2511 ( .S(n5810), .A0(n4581), .A1(wrtCnt[11]), .Z(n5782));
Q_FDP0UA U2512 ( .D(n5782), .QTFCLK( ), .Q(wrtCnt[11]));
Q_MX02 U2513 ( .S(n5810), .A0(n4582), .A1(wrtCnt[12]), .Z(n5781));
Q_FDP0UA U2514 ( .D(n5781), .QTFCLK( ), .Q(wrtCnt[12]));
Q_MX02 U2515 ( .S(n5810), .A0(n4583), .A1(wrtCnt[13]), .Z(n5780));
Q_FDP0UA U2516 ( .D(n5780), .QTFCLK( ), .Q(wrtCnt[13]));
Q_MX02 U2517 ( .S(n5810), .A0(n4584), .A1(wrtCnt[14]), .Z(n5779));
Q_FDP0UA U2518 ( .D(n5779), .QTFCLK( ), .Q(wrtCnt[14]));
Q_MX02 U2519 ( .S(n5810), .A0(n4585), .A1(wrtCnt[15]), .Z(n5778));
Q_FDP0UA U2520 ( .D(n5778), .QTFCLK( ), .Q(wrtCnt[15]));
Q_MX02 U2521 ( .S(n5810), .A0(n4586), .A1(wrtCnt[16]), .Z(n5777));
Q_FDP0UA U2522 ( .D(n5777), .QTFCLK( ), .Q(wrtCnt[16]));
Q_MX02 U2523 ( .S(n5810), .A0(n4587), .A1(wrtCnt[17]), .Z(n5776));
Q_FDP0UA U2524 ( .D(n5776), .QTFCLK( ), .Q(wrtCnt[17]));
Q_MX02 U2525 ( .S(n5810), .A0(n4588), .A1(wrtCnt[18]), .Z(n5775));
Q_FDP0UA U2526 ( .D(n5775), .QTFCLK( ), .Q(wrtCnt[18]));
Q_MX02 U2527 ( .S(n5810), .A0(n4589), .A1(wrtCnt[19]), .Z(n5774));
Q_FDP0UA U2528 ( .D(n5774), .QTFCLK( ), .Q(wrtCnt[19]));
Q_MX02 U2529 ( .S(n5810), .A0(n4590), .A1(wrtCnt[20]), .Z(n5773));
Q_FDP0UA U2530 ( .D(n5773), .QTFCLK( ), .Q(wrtCnt[20]));
Q_MX02 U2531 ( .S(n5810), .A0(n4591), .A1(wrtCnt[21]), .Z(n5772));
Q_FDP0UA U2532 ( .D(n5772), .QTFCLK( ), .Q(wrtCnt[21]));
Q_MX02 U2533 ( .S(n5810), .A0(n4592), .A1(wrtCnt[22]), .Z(n5771));
Q_FDP0UA U2534 ( .D(n5771), .QTFCLK( ), .Q(wrtCnt[22]));
Q_MX02 U2535 ( .S(n5810), .A0(n4593), .A1(wrtCnt[23]), .Z(n5770));
Q_FDP0UA U2536 ( .D(n5770), .QTFCLK( ), .Q(wrtCnt[23]));
Q_MX02 U2537 ( .S(n5810), .A0(n4594), .A1(wrtCnt[24]), .Z(n5769));
Q_FDP0UA U2538 ( .D(n5769), .QTFCLK( ), .Q(wrtCnt[24]));
Q_MX02 U2539 ( .S(n5810), .A0(n4595), .A1(wrtCnt[25]), .Z(n5768));
Q_FDP0UA U2540 ( .D(n5768), .QTFCLK( ), .Q(wrtCnt[25]));
Q_MX02 U2541 ( .S(n5810), .A0(n4596), .A1(wrtCnt[26]), .Z(n5767));
Q_FDP0UA U2542 ( .D(n5767), .QTFCLK( ), .Q(wrtCnt[26]));
Q_MX02 U2543 ( .S(n5810), .A0(n4597), .A1(wrtCnt[27]), .Z(n5766));
Q_FDP0UA U2544 ( .D(n5766), .QTFCLK( ), .Q(wrtCnt[27]));
Q_MX02 U2545 ( .S(n5810), .A0(n4598), .A1(wrtCnt[28]), .Z(n5765));
Q_FDP0UA U2546 ( .D(n5765), .QTFCLK( ), .Q(wrtCnt[28]));
Q_MX02 U2547 ( .S(n5810), .A0(n4599), .A1(wrtCnt[29]), .Z(n5764));
Q_FDP0UA U2548 ( .D(n5764), .QTFCLK( ), .Q(wrtCnt[29]));
Q_MX02 U2549 ( .S(n5810), .A0(n4600), .A1(wrtCnt[30]), .Z(n5763));
Q_FDP0UA U2550 ( .D(n5763), .QTFCLK( ), .Q(wrtCnt[30]));
Q_MX02 U2551 ( .S(n5810), .A0(n4601), .A1(wrtCnt[31]), .Z(n5762));
Q_FDP0UA U2552 ( .D(n5762), .QTFCLK( ), .Q(wrtCnt[31]));
Q_MX02 U2553 ( .S(n5810), .A0(n4602), .A1(wrtCnt[32]), .Z(n5761));
Q_FDP0UA U2554 ( .D(n5761), .QTFCLK( ), .Q(wrtCnt[32]));
Q_MX02 U2555 ( .S(n5810), .A0(n4603), .A1(wrtCnt[33]), .Z(n5760));
Q_FDP0UA U2556 ( .D(n5760), .QTFCLK( ), .Q(wrtCnt[33]));
Q_MX02 U2557 ( .S(n5810), .A0(n4604), .A1(wrtCnt[34]), .Z(n5759));
Q_FDP0UA U2558 ( .D(n5759), .QTFCLK( ), .Q(wrtCnt[34]));
Q_MX02 U2559 ( .S(n5810), .A0(n4605), .A1(wrtCnt[35]), .Z(n5758));
Q_FDP0UA U2560 ( .D(n5758), .QTFCLK( ), .Q(wrtCnt[35]));
Q_MX02 U2561 ( .S(n5810), .A0(n4606), .A1(wrtCnt[36]), .Z(n5757));
Q_FDP0UA U2562 ( .D(n5757), .QTFCLK( ), .Q(wrtCnt[36]));
Q_MX02 U2563 ( .S(n5810), .A0(n4607), .A1(wrtCnt[37]), .Z(n5756));
Q_FDP0UA U2564 ( .D(n5756), .QTFCLK( ), .Q(wrtCnt[37]));
Q_MX02 U2565 ( .S(n5810), .A0(n4608), .A1(wrtCnt[38]), .Z(n5755));
Q_FDP0UA U2566 ( .D(n5755), .QTFCLK( ), .Q(wrtCnt[38]));
Q_MX02 U2567 ( .S(n5810), .A0(n4609), .A1(wrtCnt[39]), .Z(n5754));
Q_FDP0UA U2568 ( .D(n5754), .QTFCLK( ), .Q(wrtCnt[39]));
Q_MX02 U2569 ( .S(n5810), .A0(n4610), .A1(wrtCnt[40]), .Z(n5753));
Q_FDP0UA U2570 ( .D(n5753), .QTFCLK( ), .Q(wrtCnt[40]));
Q_MX02 U2571 ( .S(n5810), .A0(n4611), .A1(wrtCnt[41]), .Z(n5752));
Q_FDP0UA U2572 ( .D(n5752), .QTFCLK( ), .Q(wrtCnt[41]));
Q_MX02 U2573 ( .S(n5810), .A0(n4612), .A1(wrtCnt[42]), .Z(n5751));
Q_FDP0UA U2574 ( .D(n5751), .QTFCLK( ), .Q(wrtCnt[42]));
Q_MX02 U2575 ( .S(n5810), .A0(n4613), .A1(wrtCnt[43]), .Z(n5750));
Q_FDP0UA U2576 ( .D(n5750), .QTFCLK( ), .Q(wrtCnt[43]));
Q_MX02 U2577 ( .S(n5810), .A0(n4614), .A1(wrtCnt[44]), .Z(n5749));
Q_FDP0UA U2578 ( .D(n5749), .QTFCLK( ), .Q(wrtCnt[44]));
Q_MX02 U2579 ( .S(n5810), .A0(n4615), .A1(wrtCnt[45]), .Z(n5748));
Q_FDP0UA U2580 ( .D(n5748), .QTFCLK( ), .Q(wrtCnt[45]));
Q_MX02 U2581 ( .S(n5810), .A0(n4616), .A1(wrtCnt[46]), .Z(n5747));
Q_FDP0UA U2582 ( .D(n5747), .QTFCLK( ), .Q(wrtCnt[46]));
Q_MX02 U2583 ( .S(n5810), .A0(n4617), .A1(wrtCnt[47]), .Z(n5746));
Q_FDP0UA U2584 ( .D(n5746), .QTFCLK( ), .Q(wrtCnt[47]));
Q_MX02 U2585 ( .S(n5810), .A0(n4618), .A1(wrtCnt[48]), .Z(n5745));
Q_FDP0UA U2586 ( .D(n5745), .QTFCLK( ), .Q(wrtCnt[48]));
Q_MX02 U2587 ( .S(n5810), .A0(n4619), .A1(wrtCnt[49]), .Z(n5744));
Q_FDP0UA U2588 ( .D(n5744), .QTFCLK( ), .Q(wrtCnt[49]));
Q_MX02 U2589 ( .S(n5810), .A0(n4620), .A1(wrtCnt[50]), .Z(n5743));
Q_FDP0UA U2590 ( .D(n5743), .QTFCLK( ), .Q(wrtCnt[50]));
Q_MX02 U2591 ( .S(n5810), .A0(n4621), .A1(wrtCnt[51]), .Z(n5742));
Q_FDP0UA U2592 ( .D(n5742), .QTFCLK( ), .Q(wrtCnt[51]));
Q_MX02 U2593 ( .S(n5810), .A0(n4622), .A1(wrtCnt[52]), .Z(n5741));
Q_FDP0UA U2594 ( .D(n5741), .QTFCLK( ), .Q(wrtCnt[52]));
Q_MX02 U2595 ( .S(n5810), .A0(n4623), .A1(wrtCnt[53]), .Z(n5740));
Q_FDP0UA U2596 ( .D(n5740), .QTFCLK( ), .Q(wrtCnt[53]));
Q_MX02 U2597 ( .S(n5810), .A0(n4624), .A1(wrtCnt[54]), .Z(n5739));
Q_FDP0UA U2598 ( .D(n5739), .QTFCLK( ), .Q(wrtCnt[54]));
Q_MX02 U2599 ( .S(n5810), .A0(n4625), .A1(wrtCnt[55]), .Z(n5738));
Q_FDP0UA U2600 ( .D(n5738), .QTFCLK( ), .Q(wrtCnt[55]));
Q_MX02 U2601 ( .S(n5810), .A0(n4626), .A1(wrtCnt[56]), .Z(n5737));
Q_FDP0UA U2602 ( .D(n5737), .QTFCLK( ), .Q(wrtCnt[56]));
Q_MX02 U2603 ( .S(n5810), .A0(n4627), .A1(wrtCnt[57]), .Z(n5736));
Q_FDP0UA U2604 ( .D(n5736), .QTFCLK( ), .Q(wrtCnt[57]));
Q_MX02 U2605 ( .S(n5810), .A0(n4628), .A1(wrtCnt[58]), .Z(n5735));
Q_FDP0UA U2606 ( .D(n5735), .QTFCLK( ), .Q(wrtCnt[58]));
Q_MX02 U2607 ( .S(n5810), .A0(n4629), .A1(wrtCnt[59]), .Z(n5734));
Q_FDP0UA U2608 ( .D(n5734), .QTFCLK( ), .Q(wrtCnt[59]));
Q_MX02 U2609 ( .S(n5810), .A0(n4630), .A1(wrtCnt[60]), .Z(n5733));
Q_FDP0UA U2610 ( .D(n5733), .QTFCLK( ), .Q(wrtCnt[60]));
Q_MX02 U2611 ( .S(n5810), .A0(n4631), .A1(wrtCnt[61]), .Z(n5732));
Q_FDP0UA U2612 ( .D(n5732), .QTFCLK( ), .Q(wrtCnt[61]));
Q_MX02 U2613 ( .S(n5810), .A0(n4632), .A1(wrtCnt[62]), .Z(n5731));
Q_FDP0UA U2614 ( .D(n5731), .QTFCLK( ), .Q(wrtCnt[62]));
Q_MX02 U2615 ( .S(n5810), .A0(n4633), .A1(wrtCnt[63]), .Z(n5730));
Q_FDP0UA U2616 ( .D(n5730), .QTFCLK( ), .Q(wrtCnt[63]));
Q_FDP0UA U2617 ( .D(n4635), .QTFCLK( ), .Q(xdata[0]));
Q_FDP0UA U2618 ( .D(n4637), .QTFCLK( ), .Q(xdata[1]));
Q_FDP0UA U2619 ( .D(n4639), .QTFCLK( ), .Q(xdata[2]));
Q_FDP0UA U2620 ( .D(n4641), .QTFCLK( ), .Q(xdata[3]));
Q_FDP0UA U2621 ( .D(n4643), .QTFCLK( ), .Q(xdata[4]));
Q_FDP0UA U2622 ( .D(n4645), .QTFCLK( ), .Q(xdata[5]));
Q_FDP0UA U2623 ( .D(n4647), .QTFCLK( ), .Q(xdata[6]));
Q_FDP0UA U2624 ( .D(n4649), .QTFCLK( ), .Q(xdata[7]));
Q_FDP0UA U2625 ( .D(n4651), .QTFCLK( ), .Q(xdata[8]));
Q_FDP0UA U2626 ( .D(n4653), .QTFCLK( ), .Q(xdata[9]));
Q_FDP0UA U2627 ( .D(n4655), .QTFCLK( ), .Q(xdata[10]));
Q_FDP0UA U2628 ( .D(n4657), .QTFCLK( ), .Q(xdata[11]));
Q_FDP0UA U2629 ( .D(n4659), .QTFCLK( ), .Q(xdata[12]));
Q_FDP0UA U2630 ( .D(n4661), .QTFCLK( ), .Q(xdata[13]));
Q_FDP0UA U2631 ( .D(n4663), .QTFCLK( ), .Q(xdata[14]));
Q_FDP0UA U2632 ( .D(n4665), .QTFCLK( ), .Q(xdata[15]));
Q_FDP0UA U2633 ( .D(n4667), .QTFCLK( ), .Q(xdata[16]));
Q_FDP0UA U2634 ( .D(n4669), .QTFCLK( ), .Q(xdata[17]));
Q_FDP0UA U2635 ( .D(n4671), .QTFCLK( ), .Q(xdata[18]));
Q_FDP0UA U2636 ( .D(n4673), .QTFCLK( ), .Q(xdata[19]));
Q_FDP0UA U2637 ( .D(n4675), .QTFCLK( ), .Q(xdata[20]));
Q_FDP0UA U2638 ( .D(n4677), .QTFCLK( ), .Q(xdata[21]));
Q_FDP0UA U2639 ( .D(n4679), .QTFCLK( ), .Q(xdata[22]));
Q_FDP0UA U2640 ( .D(n4681), .QTFCLK( ), .Q(xdata[23]));
Q_FDP0UA U2641 ( .D(n4683), .QTFCLK( ), .Q(xdata[24]));
Q_FDP0UA U2642 ( .D(n4685), .QTFCLK( ), .Q(xdata[25]));
Q_FDP0UA U2643 ( .D(n4687), .QTFCLK( ), .Q(xdata[26]));
Q_FDP0UA U2644 ( .D(n4689), .QTFCLK( ), .Q(xdata[27]));
Q_FDP0UA U2645 ( .D(n4691), .QTFCLK( ), .Q(xdata[28]));
Q_FDP0UA U2646 ( .D(n4693), .QTFCLK( ), .Q(xdata[29]));
Q_FDP0UA U2647 ( .D(n4695), .QTFCLK( ), .Q(xdata[30]));
Q_FDP0UA U2648 ( .D(n4697), .QTFCLK( ), .Q(xdata[31]));
Q_FDP0UA U2649 ( .D(n4699), .QTFCLK( ), .Q(xdata[32]));
Q_FDP0UA U2650 ( .D(n4701), .QTFCLK( ), .Q(xdata[33]));
Q_FDP0UA U2651 ( .D(n4703), .QTFCLK( ), .Q(xdata[34]));
Q_FDP0UA U2652 ( .D(n4705), .QTFCLK( ), .Q(xdata[35]));
Q_FDP0UA U2653 ( .D(n4707), .QTFCLK( ), .Q(xdata[36]));
Q_FDP0UA U2654 ( .D(n4709), .QTFCLK( ), .Q(xdata[37]));
Q_FDP0UA U2655 ( .D(n4711), .QTFCLK( ), .Q(xdata[38]));
Q_FDP0UA U2656 ( .D(n4713), .QTFCLK( ), .Q(xdata[39]));
Q_FDP0UA U2657 ( .D(n4715), .QTFCLK( ), .Q(xdata[40]));
Q_FDP0UA U2658 ( .D(n4717), .QTFCLK( ), .Q(xdata[41]));
Q_FDP0UA U2659 ( .D(n4719), .QTFCLK( ), .Q(xdata[42]));
Q_FDP0UA U2660 ( .D(n4721), .QTFCLK( ), .Q(xdata[43]));
Q_FDP0UA U2661 ( .D(n4723), .QTFCLK( ), .Q(xdata[44]));
Q_FDP0UA U2662 ( .D(n4725), .QTFCLK( ), .Q(xdata[45]));
Q_FDP0UA U2663 ( .D(n4727), .QTFCLK( ), .Q(xdata[46]));
Q_FDP0UA U2664 ( .D(n4729), .QTFCLK( ), .Q(xdata[47]));
Q_FDP0UA U2665 ( .D(n4731), .QTFCLK( ), .Q(xdata[48]));
Q_FDP0UA U2666 ( .D(n4733), .QTFCLK( ), .Q(xdata[49]));
Q_FDP0UA U2667 ( .D(n4735), .QTFCLK( ), .Q(xdata[50]));
Q_FDP0UA U2668 ( .D(n4737), .QTFCLK( ), .Q(xdata[51]));
Q_FDP0UA U2669 ( .D(n4739), .QTFCLK( ), .Q(xdata[52]));
Q_FDP0UA U2670 ( .D(n4741), .QTFCLK( ), .Q(xdata[53]));
Q_FDP0UA U2671 ( .D(n4743), .QTFCLK( ), .Q(xdata[54]));
Q_FDP0UA U2672 ( .D(n4745), .QTFCLK( ), .Q(xdata[55]));
Q_FDP0UA U2673 ( .D(n4747), .QTFCLK( ), .Q(xdata[56]));
Q_FDP0UA U2674 ( .D(n4749), .QTFCLK( ), .Q(xdata[57]));
Q_FDP0UA U2675 ( .D(n4751), .QTFCLK( ), .Q(xdata[58]));
Q_FDP0UA U2676 ( .D(n4753), .QTFCLK( ), .Q(xdata[59]));
Q_FDP0UA U2677 ( .D(n4755), .QTFCLK( ), .Q(xdata[60]));
Q_FDP0UA U2678 ( .D(n4757), .QTFCLK( ), .Q(xdata[61]));
Q_FDP0UA U2679 ( .D(n4759), .QTFCLK( ), .Q(xdata[62]));
Q_FDP0UA U2680 ( .D(n4761), .QTFCLK( ), .Q(xdata[63]));
Q_FDP0UA U2681 ( .D(n4763), .QTFCLK( ), .Q(xdata[64]));
Q_FDP0UA U2682 ( .D(n4765), .QTFCLK( ), .Q(xdata[65]));
Q_FDP0UA U2683 ( .D(n4767), .QTFCLK( ), .Q(xdata[66]));
Q_FDP0UA U2684 ( .D(n4769), .QTFCLK( ), .Q(xdata[67]));
Q_FDP0UA U2685 ( .D(n4771), .QTFCLK( ), .Q(xdata[68]));
Q_FDP0UA U2686 ( .D(n4773), .QTFCLK( ), .Q(xdata[69]));
Q_FDP0UA U2687 ( .D(n4775), .QTFCLK( ), .Q(xdata[70]));
Q_FDP0UA U2688 ( .D(n4777), .QTFCLK( ), .Q(xdata[71]));
Q_FDP0UA U2689 ( .D(n4779), .QTFCLK( ), .Q(xdata[72]));
Q_FDP0UA U2690 ( .D(n4781), .QTFCLK( ), .Q(xdata[73]));
Q_FDP0UA U2691 ( .D(n4783), .QTFCLK( ), .Q(xdata[74]));
Q_FDP0UA U2692 ( .D(n4785), .QTFCLK( ), .Q(xdata[75]));
Q_FDP0UA U2693 ( .D(n4787), .QTFCLK( ), .Q(xdata[76]));
Q_FDP0UA U2694 ( .D(n4789), .QTFCLK( ), .Q(xdata[77]));
Q_FDP0UA U2695 ( .D(n4791), .QTFCLK( ), .Q(xdata[78]));
Q_FDP0UA U2696 ( .D(n4793), .QTFCLK( ), .Q(xdata[79]));
Q_FDP0UA U2697 ( .D(n4795), .QTFCLK( ), .Q(xdata[80]));
Q_FDP0UA U2698 ( .D(n4797), .QTFCLK( ), .Q(xdata[81]));
Q_FDP0UA U2699 ( .D(n4799), .QTFCLK( ), .Q(xdata[82]));
Q_FDP0UA U2700 ( .D(n4801), .QTFCLK( ), .Q(xdata[83]));
Q_FDP0UA U2701 ( .D(n4803), .QTFCLK( ), .Q(xdata[84]));
Q_FDP0UA U2702 ( .D(n4805), .QTFCLK( ), .Q(xdata[85]));
Q_FDP0UA U2703 ( .D(n4807), .QTFCLK( ), .Q(xdata[86]));
Q_FDP0UA U2704 ( .D(n4809), .QTFCLK( ), .Q(xdata[87]));
Q_FDP0UA U2705 ( .D(n4811), .QTFCLK( ), .Q(xdata[88]));
Q_FDP0UA U2706 ( .D(n4813), .QTFCLK( ), .Q(xdata[89]));
Q_FDP0UA U2707 ( .D(n4815), .QTFCLK( ), .Q(xdata[90]));
Q_FDP0UA U2708 ( .D(n4817), .QTFCLK( ), .Q(xdata[91]));
Q_FDP0UA U2709 ( .D(n4819), .QTFCLK( ), .Q(xdata[92]));
Q_FDP0UA U2710 ( .D(n4821), .QTFCLK( ), .Q(xdata[93]));
Q_FDP0UA U2711 ( .D(n4823), .QTFCLK( ), .Q(xdata[94]));
Q_FDP0UA U2712 ( .D(n4825), .QTFCLK( ), .Q(xdata[95]));
Q_FDP0UA U2713 ( .D(n4827), .QTFCLK( ), .Q(xdata[96]));
Q_FDP0UA U2714 ( .D(n4829), .QTFCLK( ), .Q(xdata[97]));
Q_FDP0UA U2715 ( .D(n4831), .QTFCLK( ), .Q(xdata[98]));
Q_FDP0UA U2716 ( .D(n4833), .QTFCLK( ), .Q(xdata[99]));
Q_FDP0UA U2717 ( .D(n4835), .QTFCLK( ), .Q(xdata[100]));
Q_FDP0UA U2718 ( .D(n4837), .QTFCLK( ), .Q(xdata[101]));
Q_FDP0UA U2719 ( .D(n4839), .QTFCLK( ), .Q(xdata[102]));
Q_FDP0UA U2720 ( .D(n4841), .QTFCLK( ), .Q(xdata[103]));
Q_FDP0UA U2721 ( .D(n4843), .QTFCLK( ), .Q(xdata[104]));
Q_FDP0UA U2722 ( .D(n4845), .QTFCLK( ), .Q(xdata[105]));
Q_FDP0UA U2723 ( .D(n4847), .QTFCLK( ), .Q(xdata[106]));
Q_FDP0UA U2724 ( .D(n4849), .QTFCLK( ), .Q(xdata[107]));
Q_FDP0UA U2725 ( .D(n4851), .QTFCLK( ), .Q(xdata[108]));
Q_FDP0UA U2726 ( .D(n4853), .QTFCLK( ), .Q(xdata[109]));
Q_FDP0UA U2727 ( .D(n4855), .QTFCLK( ), .Q(xdata[110]));
Q_FDP0UA U2728 ( .D(n4857), .QTFCLK( ), .Q(xdata[111]));
Q_FDP0UA U2729 ( .D(n4859), .QTFCLK( ), .Q(xdata[112]));
Q_FDP0UA U2730 ( .D(n4861), .QTFCLK( ), .Q(xdata[113]));
Q_FDP0UA U2731 ( .D(n4863), .QTFCLK( ), .Q(xdata[114]));
Q_FDP0UA U2732 ( .D(n4865), .QTFCLK( ), .Q(xdata[115]));
Q_FDP0UA U2733 ( .D(n4867), .QTFCLK( ), .Q(xdata[116]));
Q_FDP0UA U2734 ( .D(n4869), .QTFCLK( ), .Q(xdata[117]));
Q_FDP0UA U2735 ( .D(n4871), .QTFCLK( ), .Q(xdata[118]));
Q_FDP0UA U2736 ( .D(n4873), .QTFCLK( ), .Q(xdata[119]));
Q_FDP0UA U2737 ( .D(n4875), .QTFCLK( ), .Q(xdata[120]));
Q_FDP0UA U2738 ( .D(n4877), .QTFCLK( ), .Q(xdata[121]));
Q_FDP0UA U2739 ( .D(n4879), .QTFCLK( ), .Q(xdata[122]));
Q_FDP0UA U2740 ( .D(n4881), .QTFCLK( ), .Q(xdata[123]));
Q_FDP0UA U2741 ( .D(n4883), .QTFCLK( ), .Q(xdata[124]));
Q_FDP0UA U2742 ( .D(n4885), .QTFCLK( ), .Q(xdata[125]));
Q_FDP0UA U2743 ( .D(n4887), .QTFCLK( ), .Q(xdata[126]));
Q_FDP0UA U2744 ( .D(n4889), .QTFCLK( ), .Q(xdata[127]));
Q_FDP0UA U2745 ( .D(n4891), .QTFCLK( ), .Q(xdata[128]));
Q_FDP0UA U2746 ( .D(n4893), .QTFCLK( ), .Q(xdata[129]));
Q_FDP0UA U2747 ( .D(n4895), .QTFCLK( ), .Q(xdata[130]));
Q_FDP0UA U2748 ( .D(n4897), .QTFCLK( ), .Q(xdata[131]));
Q_FDP0UA U2749 ( .D(n4899), .QTFCLK( ), .Q(xdata[132]));
Q_FDP0UA U2750 ( .D(n4901), .QTFCLK( ), .Q(xdata[133]));
Q_FDP0UA U2751 ( .D(n4903), .QTFCLK( ), .Q(xdata[134]));
Q_FDP0UA U2752 ( .D(n4905), .QTFCLK( ), .Q(xdata[135]));
Q_FDP0UA U2753 ( .D(n4907), .QTFCLK( ), .Q(xdata[136]));
Q_FDP0UA U2754 ( .D(n4909), .QTFCLK( ), .Q(xdata[137]));
Q_FDP0UA U2755 ( .D(n4911), .QTFCLK( ), .Q(xdata[138]));
Q_FDP0UA U2756 ( .D(n4913), .QTFCLK( ), .Q(xdata[139]));
Q_FDP0UA U2757 ( .D(n4915), .QTFCLK( ), .Q(xdata[140]));
Q_FDP0UA U2758 ( .D(n4917), .QTFCLK( ), .Q(xdata[141]));
Q_FDP0UA U2759 ( .D(n4919), .QTFCLK( ), .Q(xdata[142]));
Q_FDP0UA U2760 ( .D(n4921), .QTFCLK( ), .Q(xdata[143]));
Q_FDP0UA U2761 ( .D(n4923), .QTFCLK( ), .Q(xdata[144]));
Q_FDP0UA U2762 ( .D(n4925), .QTFCLK( ), .Q(xdata[145]));
Q_FDP0UA U2763 ( .D(n4927), .QTFCLK( ), .Q(xdata[146]));
Q_FDP0UA U2764 ( .D(n4929), .QTFCLK( ), .Q(xdata[147]));
Q_FDP0UA U2765 ( .D(n4931), .QTFCLK( ), .Q(xdata[148]));
Q_FDP0UA U2766 ( .D(n4933), .QTFCLK( ), .Q(xdata[149]));
Q_FDP0UA U2767 ( .D(n4935), .QTFCLK( ), .Q(xdata[150]));
Q_FDP0UA U2768 ( .D(n4937), .QTFCLK( ), .Q(xdata[151]));
Q_FDP0UA U2769 ( .D(n4939), .QTFCLK( ), .Q(xdata[152]));
Q_FDP0UA U2770 ( .D(n4941), .QTFCLK( ), .Q(xdata[153]));
Q_FDP0UA U2771 ( .D(n4943), .QTFCLK( ), .Q(xdata[154]));
Q_FDP0UA U2772 ( .D(n4945), .QTFCLK( ), .Q(xdata[155]));
Q_FDP0UA U2773 ( .D(n4947), .QTFCLK( ), .Q(xdata[156]));
Q_FDP0UA U2774 ( .D(n4949), .QTFCLK( ), .Q(xdata[157]));
Q_FDP0UA U2775 ( .D(n4951), .QTFCLK( ), .Q(xdata[158]));
Q_FDP0UA U2776 ( .D(n4953), .QTFCLK( ), .Q(xdata[159]));
Q_FDP0UA U2777 ( .D(n4955), .QTFCLK( ), .Q(xdata[160]));
Q_FDP0UA U2778 ( .D(n4957), .QTFCLK( ), .Q(xdata[161]));
Q_FDP0UA U2779 ( .D(n4959), .QTFCLK( ), .Q(xdata[162]));
Q_FDP0UA U2780 ( .D(n4961), .QTFCLK( ), .Q(xdata[163]));
Q_FDP0UA U2781 ( .D(n4963), .QTFCLK( ), .Q(xdata[164]));
Q_FDP0UA U2782 ( .D(n4965), .QTFCLK( ), .Q(xdata[165]));
Q_FDP0UA U2783 ( .D(n4967), .QTFCLK( ), .Q(xdata[166]));
Q_FDP0UA U2784 ( .D(n4969), .QTFCLK( ), .Q(xdata[167]));
Q_FDP0UA U2785 ( .D(n4971), .QTFCLK( ), .Q(xdata[168]));
Q_FDP0UA U2786 ( .D(n4973), .QTFCLK( ), .Q(xdata[169]));
Q_FDP0UA U2787 ( .D(n4975), .QTFCLK( ), .Q(xdata[170]));
Q_FDP0UA U2788 ( .D(n4977), .QTFCLK( ), .Q(xdata[171]));
Q_FDP0UA U2789 ( .D(n4979), .QTFCLK( ), .Q(xdata[172]));
Q_FDP0UA U2790 ( .D(n4981), .QTFCLK( ), .Q(xdata[173]));
Q_FDP0UA U2791 ( .D(n4983), .QTFCLK( ), .Q(xdata[174]));
Q_FDP0UA U2792 ( .D(n4985), .QTFCLK( ), .Q(xdata[175]));
Q_FDP0UA U2793 ( .D(n4987), .QTFCLK( ), .Q(xdata[176]));
Q_FDP0UA U2794 ( .D(n4989), .QTFCLK( ), .Q(xdata[177]));
Q_FDP0UA U2795 ( .D(n4991), .QTFCLK( ), .Q(xdata[178]));
Q_FDP0UA U2796 ( .D(n4993), .QTFCLK( ), .Q(xdata[179]));
Q_FDP0UA U2797 ( .D(n4995), .QTFCLK( ), .Q(xdata[180]));
Q_FDP0UA U2798 ( .D(n4997), .QTFCLK( ), .Q(xdata[181]));
Q_FDP0UA U2799 ( .D(n4999), .QTFCLK( ), .Q(xdata[182]));
Q_FDP0UA U2800 ( .D(n5001), .QTFCLK( ), .Q(xdata[183]));
Q_FDP0UA U2801 ( .D(n5003), .QTFCLK( ), .Q(xdata[184]));
Q_FDP0UA U2802 ( .D(n5005), .QTFCLK( ), .Q(xdata[185]));
Q_FDP0UA U2803 ( .D(n5007), .QTFCLK( ), .Q(xdata[186]));
Q_FDP0UA U2804 ( .D(n5009), .QTFCLK( ), .Q(xdata[187]));
Q_FDP0UA U2805 ( .D(n5011), .QTFCLK( ), .Q(xdata[188]));
Q_FDP0UA U2806 ( .D(n5013), .QTFCLK( ), .Q(xdata[189]));
Q_FDP0UA U2807 ( .D(n5015), .QTFCLK( ), .Q(xdata[190]));
Q_FDP0UA U2808 ( .D(n5017), .QTFCLK( ), .Q(xdata[191]));
Q_FDP0UA U2809 ( .D(n5019), .QTFCLK( ), .Q(xdata[192]));
Q_FDP0UA U2810 ( .D(n5021), .QTFCLK( ), .Q(xdata[193]));
Q_FDP0UA U2811 ( .D(n5023), .QTFCLK( ), .Q(xdata[194]));
Q_FDP0UA U2812 ( .D(n5025), .QTFCLK( ), .Q(xdata[195]));
Q_FDP0UA U2813 ( .D(n5027), .QTFCLK( ), .Q(xdata[196]));
Q_FDP0UA U2814 ( .D(n5029), .QTFCLK( ), .Q(xdata[197]));
Q_FDP0UA U2815 ( .D(n5031), .QTFCLK( ), .Q(xdata[198]));
Q_FDP0UA U2816 ( .D(n5033), .QTFCLK( ), .Q(xdata[199]));
Q_FDP0UA U2817 ( .D(n5035), .QTFCLK( ), .Q(xdata[200]));
Q_FDP0UA U2818 ( .D(n5037), .QTFCLK( ), .Q(xdata[201]));
Q_FDP0UA U2819 ( .D(n5039), .QTFCLK( ), .Q(xdata[202]));
Q_FDP0UA U2820 ( .D(n5041), .QTFCLK( ), .Q(xdata[203]));
Q_FDP0UA U2821 ( .D(n5043), .QTFCLK( ), .Q(xdata[204]));
Q_FDP0UA U2822 ( .D(n5045), .QTFCLK( ), .Q(xdata[205]));
Q_FDP0UA U2823 ( .D(n5047), .QTFCLK( ), .Q(xdata[206]));
Q_FDP0UA U2824 ( .D(n5049), .QTFCLK( ), .Q(xdata[207]));
Q_FDP0UA U2825 ( .D(n5051), .QTFCLK( ), .Q(xdata[208]));
Q_FDP0UA U2826 ( .D(n5053), .QTFCLK( ), .Q(xdata[209]));
Q_FDP0UA U2827 ( .D(n5055), .QTFCLK( ), .Q(xdata[210]));
Q_FDP0UA U2828 ( .D(n5057), .QTFCLK( ), .Q(xdata[211]));
Q_FDP0UA U2829 ( .D(n5059), .QTFCLK( ), .Q(xdata[212]));
Q_FDP0UA U2830 ( .D(n5061), .QTFCLK( ), .Q(xdata[213]));
Q_FDP0UA U2831 ( .D(n5063), .QTFCLK( ), .Q(xdata[214]));
Q_FDP0UA U2832 ( .D(n5065), .QTFCLK( ), .Q(xdata[215]));
Q_FDP0UA U2833 ( .D(n5067), .QTFCLK( ), .Q(xdata[216]));
Q_FDP0UA U2834 ( .D(n5069), .QTFCLK( ), .Q(xdata[217]));
Q_FDP0UA U2835 ( .D(n5071), .QTFCLK( ), .Q(xdata[218]));
Q_FDP0UA U2836 ( .D(n5073), .QTFCLK( ), .Q(xdata[219]));
Q_FDP0UA U2837 ( .D(n5075), .QTFCLK( ), .Q(xdata[220]));
Q_FDP0UA U2838 ( .D(n5077), .QTFCLK( ), .Q(xdata[221]));
Q_FDP0UA U2839 ( .D(n5079), .QTFCLK( ), .Q(xdata[222]));
Q_FDP0UA U2840 ( .D(n5081), .QTFCLK( ), .Q(xdata[223]));
Q_FDP0UA U2841 ( .D(n5083), .QTFCLK( ), .Q(xdata[224]));
Q_FDP0UA U2842 ( .D(n5085), .QTFCLK( ), .Q(xdata[225]));
Q_FDP0UA U2843 ( .D(n5087), .QTFCLK( ), .Q(xdata[226]));
Q_FDP0UA U2844 ( .D(n5089), .QTFCLK( ), .Q(xdata[227]));
Q_FDP0UA U2845 ( .D(n5091), .QTFCLK( ), .Q(xdata[228]));
Q_FDP0UA U2846 ( .D(n5093), .QTFCLK( ), .Q(xdata[229]));
Q_FDP0UA U2847 ( .D(n5095), .QTFCLK( ), .Q(xdata[230]));
Q_FDP0UA U2848 ( .D(n5097), .QTFCLK( ), .Q(xdata[231]));
Q_FDP0UA U2849 ( .D(n5099), .QTFCLK( ), .Q(xdata[232]));
Q_FDP0UA U2850 ( .D(n5101), .QTFCLK( ), .Q(xdata[233]));
Q_FDP0UA U2851 ( .D(n5103), .QTFCLK( ), .Q(xdata[234]));
Q_FDP0UA U2852 ( .D(n5105), .QTFCLK( ), .Q(xdata[235]));
Q_FDP0UA U2853 ( .D(n5107), .QTFCLK( ), .Q(xdata[236]));
Q_FDP0UA U2854 ( .D(n5109), .QTFCLK( ), .Q(xdata[237]));
Q_FDP0UA U2855 ( .D(n5111), .QTFCLK( ), .Q(xdata[238]));
Q_FDP0UA U2856 ( .D(n5113), .QTFCLK( ), .Q(xdata[239]));
Q_FDP0UA U2857 ( .D(n5115), .QTFCLK( ), .Q(xdata[240]));
Q_FDP0UA U2858 ( .D(n5117), .QTFCLK( ), .Q(xdata[241]));
Q_FDP0UA U2859 ( .D(n5119), .QTFCLK( ), .Q(xdata[242]));
Q_FDP0UA U2860 ( .D(n5121), .QTFCLK( ), .Q(xdata[243]));
Q_FDP0UA U2861 ( .D(n5123), .QTFCLK( ), .Q(xdata[244]));
Q_FDP0UA U2862 ( .D(n5125), .QTFCLK( ), .Q(xdata[245]));
Q_FDP0UA U2863 ( .D(n5127), .QTFCLK( ), .Q(xdata[246]));
Q_FDP0UA U2864 ( .D(n5129), .QTFCLK( ), .Q(xdata[247]));
Q_FDP0UA U2865 ( .D(n5131), .QTFCLK( ), .Q(xdata[248]));
Q_FDP0UA U2866 ( .D(n5133), .QTFCLK( ), .Q(xdata[249]));
Q_FDP0UA U2867 ( .D(n5135), .QTFCLK( ), .Q(xdata[250]));
Q_FDP0UA U2868 ( .D(n5137), .QTFCLK( ), .Q(xdata[251]));
Q_FDP0UA U2869 ( .D(n5139), .QTFCLK( ), .Q(xdata[252]));
Q_FDP0UA U2870 ( .D(n5141), .QTFCLK( ), .Q(xdata[253]));
Q_FDP0UA U2871 ( .D(n5143), .QTFCLK( ), .Q(xdata[254]));
Q_FDP0UA U2872 ( .D(n5145), .QTFCLK( ), .Q(xdata[255]));
Q_FDP0UA U2873 ( .D(n5147), .QTFCLK( ), .Q(xdata[256]));
Q_FDP0UA U2874 ( .D(n5149), .QTFCLK( ), .Q(xdata[257]));
Q_FDP0UA U2875 ( .D(n5151), .QTFCLK( ), .Q(xdata[258]));
Q_FDP0UA U2876 ( .D(n5153), .QTFCLK( ), .Q(xdata[259]));
Q_FDP0UA U2877 ( .D(n5155), .QTFCLK( ), .Q(xdata[260]));
Q_FDP0UA U2878 ( .D(n5157), .QTFCLK( ), .Q(xdata[261]));
Q_FDP0UA U2879 ( .D(n5159), .QTFCLK( ), .Q(xdata[262]));
Q_FDP0UA U2880 ( .D(n5161), .QTFCLK( ), .Q(xdata[263]));
Q_FDP0UA U2881 ( .D(n5163), .QTFCLK( ), .Q(xdata[264]));
Q_FDP0UA U2882 ( .D(n5165), .QTFCLK( ), .Q(xdata[265]));
Q_FDP0UA U2883 ( .D(n5167), .QTFCLK( ), .Q(xdata[266]));
Q_FDP0UA U2884 ( .D(n5169), .QTFCLK( ), .Q(xdata[267]));
Q_FDP0UA U2885 ( .D(n5171), .QTFCLK( ), .Q(xdata[268]));
Q_FDP0UA U2886 ( .D(n5173), .QTFCLK( ), .Q(xdata[269]));
Q_FDP0UA U2887 ( .D(n5175), .QTFCLK( ), .Q(xdata[270]));
Q_FDP0UA U2888 ( .D(n5177), .QTFCLK( ), .Q(xdata[271]));
Q_FDP0UA U2889 ( .D(n5179), .QTFCLK( ), .Q(xdata[272]));
Q_FDP0UA U2890 ( .D(n5181), .QTFCLK( ), .Q(xdata[273]));
Q_FDP0UA U2891 ( .D(n5183), .QTFCLK( ), .Q(xdata[274]));
Q_FDP0UA U2892 ( .D(n5185), .QTFCLK( ), .Q(xdata[275]));
Q_FDP0UA U2893 ( .D(n5187), .QTFCLK( ), .Q(xdata[276]));
Q_FDP0UA U2894 ( .D(n5189), .QTFCLK( ), .Q(xdata[277]));
Q_FDP0UA U2895 ( .D(n5191), .QTFCLK( ), .Q(xdata[278]));
Q_FDP0UA U2896 ( .D(n5193), .QTFCLK( ), .Q(xdata[279]));
Q_FDP0UA U2897 ( .D(n5195), .QTFCLK( ), .Q(xdata[280]));
Q_FDP0UA U2898 ( .D(n5197), .QTFCLK( ), .Q(xdata[281]));
Q_FDP0UA U2899 ( .D(n5199), .QTFCLK( ), .Q(xdata[282]));
Q_FDP0UA U2900 ( .D(n5201), .QTFCLK( ), .Q(xdata[283]));
Q_FDP0UA U2901 ( .D(n5203), .QTFCLK( ), .Q(xdata[284]));
Q_FDP0UA U2902 ( .D(n5205), .QTFCLK( ), .Q(xdata[285]));
Q_FDP0UA U2903 ( .D(n5207), .QTFCLK( ), .Q(xdata[286]));
Q_FDP0UA U2904 ( .D(n5209), .QTFCLK( ), .Q(xdata[287]));
Q_FDP0UA U2905 ( .D(n5211), .QTFCLK( ), .Q(xdata[288]));
Q_FDP0UA U2906 ( .D(n5213), .QTFCLK( ), .Q(xdata[289]));
Q_FDP0UA U2907 ( .D(n5215), .QTFCLK( ), .Q(xdata[290]));
Q_FDP0UA U2908 ( .D(n5217), .QTFCLK( ), .Q(xdata[291]));
Q_FDP0UA U2909 ( .D(n5219), .QTFCLK( ), .Q(xdata[292]));
Q_FDP0UA U2910 ( .D(n5221), .QTFCLK( ), .Q(xdata[293]));
Q_FDP0UA U2911 ( .D(n5223), .QTFCLK( ), .Q(xdata[294]));
Q_FDP0UA U2912 ( .D(n5225), .QTFCLK( ), .Q(xdata[295]));
Q_FDP0UA U2913 ( .D(n5227), .QTFCLK( ), .Q(xdata[296]));
Q_FDP0UA U2914 ( .D(n5229), .QTFCLK( ), .Q(xdata[297]));
Q_FDP0UA U2915 ( .D(n5231), .QTFCLK( ), .Q(xdata[298]));
Q_FDP0UA U2916 ( .D(n5233), .QTFCLK( ), .Q(xdata[299]));
Q_FDP0UA U2917 ( .D(n5235), .QTFCLK( ), .Q(xdata[300]));
Q_FDP0UA U2918 ( .D(n5237), .QTFCLK( ), .Q(xdata[301]));
Q_FDP0UA U2919 ( .D(n5239), .QTFCLK( ), .Q(xdata[302]));
Q_FDP0UA U2920 ( .D(n5241), .QTFCLK( ), .Q(xdata[303]));
Q_FDP0UA U2921 ( .D(n5243), .QTFCLK( ), .Q(xdata[304]));
Q_FDP0UA U2922 ( .D(n5245), .QTFCLK( ), .Q(xdata[305]));
Q_FDP0UA U2923 ( .D(n5247), .QTFCLK( ), .Q(xdata[306]));
Q_FDP0UA U2924 ( .D(n5249), .QTFCLK( ), .Q(xdata[307]));
Q_FDP0UA U2925 ( .D(n5251), .QTFCLK( ), .Q(xdata[308]));
Q_FDP0UA U2926 ( .D(n5253), .QTFCLK( ), .Q(xdata[309]));
Q_FDP0UA U2927 ( .D(n5255), .QTFCLK( ), .Q(xdata[310]));
Q_FDP0UA U2928 ( .D(n5257), .QTFCLK( ), .Q(xdata[311]));
Q_FDP0UA U2929 ( .D(n5259), .QTFCLK( ), .Q(xdata[312]));
Q_FDP0UA U2930 ( .D(n5261), .QTFCLK( ), .Q(xdata[313]));
Q_FDP0UA U2931 ( .D(n5263), .QTFCLK( ), .Q(xdata[314]));
Q_FDP0UA U2932 ( .D(n5265), .QTFCLK( ), .Q(xdata[315]));
Q_FDP0UA U2933 ( .D(n5267), .QTFCLK( ), .Q(xdata[316]));
Q_FDP0UA U2934 ( .D(n5269), .QTFCLK( ), .Q(xdata[317]));
Q_FDP0UA U2935 ( .D(n5271), .QTFCLK( ), .Q(xdata[318]));
Q_FDP0UA U2936 ( .D(n5273), .QTFCLK( ), .Q(xdata[319]));
Q_FDP0UA U2937 ( .D(n5275), .QTFCLK( ), .Q(xdata[320]));
Q_FDP0UA U2938 ( .D(n5277), .QTFCLK( ), .Q(xdata[321]));
Q_FDP0UA U2939 ( .D(n5279), .QTFCLK( ), .Q(xdata[322]));
Q_FDP0UA U2940 ( .D(n5281), .QTFCLK( ), .Q(xdata[323]));
Q_FDP0UA U2941 ( .D(n5283), .QTFCLK( ), .Q(xdata[324]));
Q_FDP0UA U2942 ( .D(n5285), .QTFCLK( ), .Q(xdata[325]));
Q_FDP0UA U2943 ( .D(n5287), .QTFCLK( ), .Q(xdata[326]));
Q_FDP0UA U2944 ( .D(n5289), .QTFCLK( ), .Q(xdata[327]));
Q_FDP0UA U2945 ( .D(n5291), .QTFCLK( ), .Q(xdata[328]));
Q_FDP0UA U2946 ( .D(n5293), .QTFCLK( ), .Q(xdata[329]));
Q_FDP0UA U2947 ( .D(n5295), .QTFCLK( ), .Q(xdata[330]));
Q_FDP0UA U2948 ( .D(n5297), .QTFCLK( ), .Q(xdata[331]));
Q_FDP0UA U2949 ( .D(n5299), .QTFCLK( ), .Q(xdata[332]));
Q_FDP0UA U2950 ( .D(n5301), .QTFCLK( ), .Q(xdata[333]));
Q_FDP0UA U2951 ( .D(n5303), .QTFCLK( ), .Q(xdata[334]));
Q_FDP0UA U2952 ( .D(n5305), .QTFCLK( ), .Q(xdata[335]));
Q_FDP0UA U2953 ( .D(n5307), .QTFCLK( ), .Q(xdata[336]));
Q_FDP0UA U2954 ( .D(n5309), .QTFCLK( ), .Q(xdata[337]));
Q_FDP0UA U2955 ( .D(n5311), .QTFCLK( ), .Q(xdata[338]));
Q_FDP0UA U2956 ( .D(n5313), .QTFCLK( ), .Q(xdata[339]));
Q_FDP0UA U2957 ( .D(n5315), .QTFCLK( ), .Q(xdata[340]));
Q_FDP0UA U2958 ( .D(n5317), .QTFCLK( ), .Q(xdata[341]));
Q_FDP0UA U2959 ( .D(n5319), .QTFCLK( ), .Q(xdata[342]));
Q_FDP0UA U2960 ( .D(n5321), .QTFCLK( ), .Q(xdata[343]));
Q_FDP0UA U2961 ( .D(n5323), .QTFCLK( ), .Q(xdata[344]));
Q_FDP0UA U2962 ( .D(n5325), .QTFCLK( ), .Q(xdata[345]));
Q_FDP0UA U2963 ( .D(n5327), .QTFCLK( ), .Q(xdata[346]));
Q_FDP0UA U2964 ( .D(n5329), .QTFCLK( ), .Q(xdata[347]));
Q_FDP0UA U2965 ( .D(n5331), .QTFCLK( ), .Q(xdata[348]));
Q_FDP0UA U2966 ( .D(n5333), .QTFCLK( ), .Q(xdata[349]));
Q_FDP0UA U2967 ( .D(n5335), .QTFCLK( ), .Q(xdata[350]));
Q_FDP0UA U2968 ( .D(n5337), .QTFCLK( ), .Q(xdata[351]));
Q_FDP0UA U2969 ( .D(n5339), .QTFCLK( ), .Q(xdata[352]));
Q_FDP0UA U2970 ( .D(n5341), .QTFCLK( ), .Q(xdata[353]));
Q_FDP0UA U2971 ( .D(n5343), .QTFCLK( ), .Q(xdata[354]));
Q_FDP0UA U2972 ( .D(n5345), .QTFCLK( ), .Q(xdata[355]));
Q_FDP0UA U2973 ( .D(n5347), .QTFCLK( ), .Q(xdata[356]));
Q_FDP0UA U2974 ( .D(n5349), .QTFCLK( ), .Q(xdata[357]));
Q_FDP0UA U2975 ( .D(n5351), .QTFCLK( ), .Q(xdata[358]));
Q_FDP0UA U2976 ( .D(n5353), .QTFCLK( ), .Q(xdata[359]));
Q_FDP0UA U2977 ( .D(n5355), .QTFCLK( ), .Q(xdata[360]));
Q_FDP0UA U2978 ( .D(n5357), .QTFCLK( ), .Q(xdata[361]));
Q_FDP0UA U2979 ( .D(n5359), .QTFCLK( ), .Q(xdata[362]));
Q_FDP0UA U2980 ( .D(n5361), .QTFCLK( ), .Q(xdata[363]));
Q_FDP0UA U2981 ( .D(n5363), .QTFCLK( ), .Q(xdata[364]));
Q_FDP0UA U2982 ( .D(n5365), .QTFCLK( ), .Q(xdata[365]));
Q_FDP0UA U2983 ( .D(n5367), .QTFCLK( ), .Q(xdata[366]));
Q_FDP0UA U2984 ( .D(n5369), .QTFCLK( ), .Q(xdata[367]));
Q_FDP0UA U2985 ( .D(n5371), .QTFCLK( ), .Q(xdata[368]));
Q_FDP0UA U2986 ( .D(n5373), .QTFCLK( ), .Q(xdata[369]));
Q_FDP0UA U2987 ( .D(n5375), .QTFCLK( ), .Q(xdata[370]));
Q_FDP0UA U2988 ( .D(n5377), .QTFCLK( ), .Q(xdata[371]));
Q_FDP0UA U2989 ( .D(n5379), .QTFCLK( ), .Q(xdata[372]));
Q_FDP0UA U2990 ( .D(n5381), .QTFCLK( ), .Q(xdata[373]));
Q_FDP0UA U2991 ( .D(n5383), .QTFCLK( ), .Q(xdata[374]));
Q_FDP0UA U2992 ( .D(n5385), .QTFCLK( ), .Q(xdata[375]));
Q_FDP0UA U2993 ( .D(n5387), .QTFCLK( ), .Q(xdata[376]));
Q_FDP0UA U2994 ( .D(n5389), .QTFCLK( ), .Q(xdata[377]));
Q_FDP0UA U2995 ( .D(n5391), .QTFCLK( ), .Q(xdata[378]));
Q_FDP0UA U2996 ( .D(n5393), .QTFCLK( ), .Q(xdata[379]));
Q_FDP0UA U2997 ( .D(n5395), .QTFCLK( ), .Q(xdata[380]));
Q_FDP0UA U2998 ( .D(n5397), .QTFCLK( ), .Q(xdata[381]));
Q_FDP0UA U2999 ( .D(n5399), .QTFCLK( ), .Q(xdata[382]));
Q_FDP0UA U3000 ( .D(n5401), .QTFCLK( ), .Q(xdata[383]));
Q_FDP0UA U3001 ( .D(n5403), .QTFCLK( ), .Q(xdata[384]));
Q_FDP0UA U3002 ( .D(n5405), .QTFCLK( ), .Q(xdata[385]));
Q_FDP0UA U3003 ( .D(n5407), .QTFCLK( ), .Q(xdata[386]));
Q_FDP0UA U3004 ( .D(n5409), .QTFCLK( ), .Q(xdata[387]));
Q_FDP0UA U3005 ( .D(n5411), .QTFCLK( ), .Q(xdata[388]));
Q_FDP0UA U3006 ( .D(n5413), .QTFCLK( ), .Q(xdata[389]));
Q_FDP0UA U3007 ( .D(n5415), .QTFCLK( ), .Q(xdata[390]));
Q_FDP0UA U3008 ( .D(n5417), .QTFCLK( ), .Q(xdata[391]));
Q_FDP0UA U3009 ( .D(n5419), .QTFCLK( ), .Q(xdata[392]));
Q_FDP0UA U3010 ( .D(n5421), .QTFCLK( ), .Q(xdata[393]));
Q_FDP0UA U3011 ( .D(n5423), .QTFCLK( ), .Q(xdata[394]));
Q_FDP0UA U3012 ( .D(n5425), .QTFCLK( ), .Q(xdata[395]));
Q_FDP0UA U3013 ( .D(n5427), .QTFCLK( ), .Q(xdata[396]));
Q_FDP0UA U3014 ( .D(n5429), .QTFCLK( ), .Q(xdata[397]));
Q_FDP0UA U3015 ( .D(n5431), .QTFCLK( ), .Q(xdata[398]));
Q_FDP0UA U3016 ( .D(n5433), .QTFCLK( ), .Q(xdata[399]));
Q_FDP0UA U3017 ( .D(n5435), .QTFCLK( ), .Q(xdata[400]));
Q_FDP0UA U3018 ( .D(n5437), .QTFCLK( ), .Q(xdata[401]));
Q_FDP0UA U3019 ( .D(n5439), .QTFCLK( ), .Q(xdata[402]));
Q_FDP0UA U3020 ( .D(n5441), .QTFCLK( ), .Q(xdata[403]));
Q_FDP0UA U3021 ( .D(n5443), .QTFCLK( ), .Q(xdata[404]));
Q_FDP0UA U3022 ( .D(n5445), .QTFCLK( ), .Q(xdata[405]));
Q_FDP0UA U3023 ( .D(n5447), .QTFCLK( ), .Q(xdata[406]));
Q_FDP0UA U3024 ( .D(n5449), .QTFCLK( ), .Q(xdata[407]));
Q_FDP0UA U3025 ( .D(n5451), .QTFCLK( ), .Q(xdata[408]));
Q_FDP0UA U3026 ( .D(n5453), .QTFCLK( ), .Q(xdata[409]));
Q_FDP0UA U3027 ( .D(n5455), .QTFCLK( ), .Q(xdata[410]));
Q_FDP0UA U3028 ( .D(n5457), .QTFCLK( ), .Q(xdata[411]));
Q_FDP0UA U3029 ( .D(n5459), .QTFCLK( ), .Q(xdata[412]));
Q_FDP0UA U3030 ( .D(n5461), .QTFCLK( ), .Q(xdata[413]));
Q_FDP0UA U3031 ( .D(n5463), .QTFCLK( ), .Q(xdata[414]));
Q_FDP0UA U3032 ( .D(n5465), .QTFCLK( ), .Q(xdata[415]));
Q_FDP0UA U3033 ( .D(n5467), .QTFCLK( ), .Q(xdata[416]));
Q_FDP0UA U3034 ( .D(n5469), .QTFCLK( ), .Q(xdata[417]));
Q_FDP0UA U3035 ( .D(n5471), .QTFCLK( ), .Q(xdata[418]));
Q_FDP0UA U3036 ( .D(n5473), .QTFCLK( ), .Q(xdata[419]));
Q_FDP0UA U3037 ( .D(n5475), .QTFCLK( ), .Q(xdata[420]));
Q_FDP0UA U3038 ( .D(n5477), .QTFCLK( ), .Q(xdata[421]));
Q_FDP0UA U3039 ( .D(n5479), .QTFCLK( ), .Q(xdata[422]));
Q_FDP0UA U3040 ( .D(n5481), .QTFCLK( ), .Q(xdata[423]));
Q_FDP0UA U3041 ( .D(n5483), .QTFCLK( ), .Q(xdata[424]));
Q_FDP0UA U3042 ( .D(n5485), .QTFCLK( ), .Q(xdata[425]));
Q_FDP0UA U3043 ( .D(n5487), .QTFCLK( ), .Q(xdata[426]));
Q_FDP0UA U3044 ( .D(n5489), .QTFCLK( ), .Q(xdata[427]));
Q_FDP0UA U3045 ( .D(n5491), .QTFCLK( ), .Q(xdata[428]));
Q_FDP0UA U3046 ( .D(n5493), .QTFCLK( ), .Q(xdata[429]));
Q_FDP0UA U3047 ( .D(n5495), .QTFCLK( ), .Q(xdata[430]));
Q_FDP0UA U3048 ( .D(n5497), .QTFCLK( ), .Q(xdata[431]));
Q_FDP0UA U3049 ( .D(n5499), .QTFCLK( ), .Q(xdata[432]));
Q_FDP0UA U3050 ( .D(n5501), .QTFCLK( ), .Q(xdata[433]));
Q_FDP0UA U3051 ( .D(n5503), .QTFCLK( ), .Q(xdata[434]));
Q_FDP0UA U3052 ( .D(n5505), .QTFCLK( ), .Q(xdata[435]));
Q_FDP0UA U3053 ( .D(n5507), .QTFCLK( ), .Q(xdata[436]));
Q_FDP0UA U3054 ( .D(n5509), .QTFCLK( ), .Q(xdata[437]));
Q_FDP0UA U3055 ( .D(n5511), .QTFCLK( ), .Q(xdata[438]));
Q_FDP0UA U3056 ( .D(n5513), .QTFCLK( ), .Q(xdata[439]));
Q_FDP0UA U3057 ( .D(n5515), .QTFCLK( ), .Q(xdata[440]));
Q_FDP0UA U3058 ( .D(n5517), .QTFCLK( ), .Q(xdata[441]));
Q_FDP0UA U3059 ( .D(n5519), .QTFCLK( ), .Q(xdata[442]));
Q_FDP0UA U3060 ( .D(n5521), .QTFCLK( ), .Q(xdata[443]));
Q_FDP0UA U3061 ( .D(n5523), .QTFCLK( ), .Q(xdata[444]));
Q_FDP0UA U3062 ( .D(n5525), .QTFCLK( ), .Q(xdata[445]));
Q_FDP0UA U3063 ( .D(n5527), .QTFCLK( ), .Q(xdata[446]));
Q_FDP0UA U3064 ( .D(n5529), .QTFCLK( ), .Q(xdata[447]));
Q_FDP0UA U3065 ( .D(n5531), .QTFCLK( ), .Q(xdata[448]));
Q_FDP0UA U3066 ( .D(n5533), .QTFCLK( ), .Q(xdata[449]));
Q_FDP0UA U3067 ( .D(n5535), .QTFCLK( ), .Q(xdata[450]));
Q_FDP0UA U3068 ( .D(n5537), .QTFCLK( ), .Q(xdata[451]));
Q_FDP0UA U3069 ( .D(n5539), .QTFCLK( ), .Q(xdata[452]));
Q_FDP0UA U3070 ( .D(n5541), .QTFCLK( ), .Q(xdata[453]));
Q_FDP0UA U3071 ( .D(n5543), .QTFCLK( ), .Q(xdata[454]));
Q_FDP0UA U3072 ( .D(n5545), .QTFCLK( ), .Q(xdata[455]));
Q_FDP0UA U3073 ( .D(n5547), .QTFCLK( ), .Q(xdata[456]));
Q_FDP0UA U3074 ( .D(n5549), .QTFCLK( ), .Q(xdata[457]));
Q_FDP0UA U3075 ( .D(n5551), .QTFCLK( ), .Q(xdata[458]));
Q_FDP0UA U3076 ( .D(n5553), .QTFCLK( ), .Q(xdata[459]));
Q_FDP0UA U3077 ( .D(n5555), .QTFCLK( ), .Q(xdata[460]));
Q_FDP0UA U3078 ( .D(n5557), .QTFCLK( ), .Q(xdata[461]));
Q_FDP0UA U3079 ( .D(n5559), .QTFCLK( ), .Q(xdata[462]));
Q_FDP0UA U3080 ( .D(n5561), .QTFCLK( ), .Q(xdata[463]));
Q_FDP0UA U3081 ( .D(n5563), .QTFCLK( ), .Q(xdata[464]));
Q_FDP0UA U3082 ( .D(n5565), .QTFCLK( ), .Q(xdata[465]));
Q_FDP0UA U3083 ( .D(n5567), .QTFCLK( ), .Q(xdata[466]));
Q_FDP0UA U3084 ( .D(n5569), .QTFCLK( ), .Q(xdata[467]));
Q_FDP0UA U3085 ( .D(n5571), .QTFCLK( ), .Q(xdata[468]));
Q_FDP0UA U3086 ( .D(n5573), .QTFCLK( ), .Q(xdata[469]));
Q_FDP0UA U3087 ( .D(n5575), .QTFCLK( ), .Q(xdata[470]));
Q_FDP0UA U3088 ( .D(n5577), .QTFCLK( ), .Q(xdata[471]));
Q_FDP0UA U3089 ( .D(n5579), .QTFCLK( ), .Q(xdata[472]));
Q_FDP0UA U3090 ( .D(n5581), .QTFCLK( ), .Q(xdata[473]));
Q_FDP0UA U3091 ( .D(n5583), .QTFCLK( ), .Q(xdata[474]));
Q_FDP0UA U3092 ( .D(n5585), .QTFCLK( ), .Q(xdata[475]));
Q_FDP0UA U3093 ( .D(n5587), .QTFCLK( ), .Q(xdata[476]));
Q_FDP0UA U3094 ( .D(n5589), .QTFCLK( ), .Q(xdata[477]));
Q_FDP0UA U3095 ( .D(n5591), .QTFCLK( ), .Q(xdata[478]));
Q_FDP0UA U3096 ( .D(n5593), .QTFCLK( ), .Q(xdata[479]));
Q_FDP0UA U3097 ( .D(n5595), .QTFCLK( ), .Q(xdata[480]));
Q_FDP0UA U3098 ( .D(n5597), .QTFCLK( ), .Q(xdata[481]));
Q_FDP0UA U3099 ( .D(n5599), .QTFCLK( ), .Q(xdata[482]));
Q_FDP0UA U3100 ( .D(n5601), .QTFCLK( ), .Q(xdata[483]));
Q_FDP0UA U3101 ( .D(n5603), .QTFCLK( ), .Q(xdata[484]));
Q_FDP0UA U3102 ( .D(n5605), .QTFCLK( ), .Q(xdata[485]));
Q_FDP0UA U3103 ( .D(n5607), .QTFCLK( ), .Q(xdata[486]));
Q_FDP0UA U3104 ( .D(n5609), .QTFCLK( ), .Q(xdata[487]));
Q_FDP0UA U3105 ( .D(n5611), .QTFCLK( ), .Q(xdata[488]));
Q_FDP0UA U3106 ( .D(n5613), .QTFCLK( ), .Q(xdata[489]));
Q_FDP0UA U3107 ( .D(n5615), .QTFCLK( ), .Q(xdata[490]));
Q_FDP0UA U3108 ( .D(n5617), .QTFCLK( ), .Q(xdata[491]));
Q_FDP0UA U3109 ( .D(n5619), .QTFCLK( ), .Q(xdata[492]));
Q_FDP0UA U3110 ( .D(n5621), .QTFCLK( ), .Q(xdata[493]));
Q_FDP0UA U3111 ( .D(n5623), .QTFCLK( ), .Q(xdata[494]));
Q_FDP0UA U3112 ( .D(n5625), .QTFCLK( ), .Q(xdata[495]));
Q_FDP0UA U3113 ( .D(n5627), .QTFCLK( ), .Q(xdata[496]));
Q_FDP0UA U3114 ( .D(n5629), .QTFCLK( ), .Q(xdata[497]));
Q_FDP0UA U3115 ( .D(n5631), .QTFCLK( ), .Q(xdata[498]));
Q_FDP0UA U3116 ( .D(n5633), .QTFCLK( ), .Q(xdata[499]));
Q_FDP0UA U3117 ( .D(n5635), .QTFCLK( ), .Q(xdata[500]));
Q_FDP0UA U3118 ( .D(n5637), .QTFCLK( ), .Q(xdata[501]));
Q_FDP0UA U3119 ( .D(n5639), .QTFCLK( ), .Q(xdata[502]));
Q_FDP0UA U3120 ( .D(n5641), .QTFCLK( ), .Q(xdata[503]));
Q_FDP0UA U3121 ( .D(n5643), .QTFCLK( ), .Q(xdata[504]));
Q_FDP0UA U3122 ( .D(n5645), .QTFCLK( ), .Q(xdata[505]));
Q_FDP0UA U3123 ( .D(n5647), .QTFCLK( ), .Q(xdata[506]));
Q_FDP0UA U3124 ( .D(n5649), .QTFCLK( ), .Q(xdata[507]));
Q_FDP0UA U3125 ( .D(n5651), .QTFCLK( ), .Q(xdata[508]));
Q_FDP0UA U3126 ( .D(n5653), .QTFCLK( ), .Q(xdata[509]));
Q_FDP0UA U3127 ( .D(n5655), .QTFCLK( ), .Q(xdata[510]));
Q_FDP0UA U3128 ( .D(n5657), .QTFCLK( ), .Q(xdata[511]));
Q_FDP0UA U3129 ( .D(n5658), .QTFCLK( ), .Q(xdata[512]));
Q_FDP0UA U3130 ( .D(n5659), .QTFCLK( ), .Q(xdata[513]));
Q_FDP0UA U3131 ( .D(n5660), .QTFCLK( ), .Q(xdata[514]));
Q_FDP0UA U3132 ( .D(n5661), .QTFCLK( ), .Q(xdata[515]));
Q_FDP0UA U3133 ( .D(n5662), .QTFCLK( ), .Q(xdata[516]));
Q_FDP0UA U3134 ( .D(n5663), .QTFCLK( ), .Q(xdata[517]));
Q_FDP0UA U3135 ( .D(n5664), .QTFCLK( ), .Q(xdata[518]));
Q_FDP0UA U3136 ( .D(n5665), .QTFCLK( ), .Q(xdata[519]));
Q_FDP0UA U3137 ( .D(n5666), .QTFCLK( ), .Q(xdata[520]));
Q_FDP0UA U3138 ( .D(n5667), .QTFCLK( ), .Q(xdata[521]));
Q_FDP0UA U3139 ( .D(n5668), .QTFCLK( ), .Q(xdata[522]));
Q_FDP0UA U3140 ( .D(n5669), .QTFCLK( ), .Q(xdata[523]));
Q_FDP0UA U3141 ( .D(n5670), .QTFCLK( ), .Q(xdata[524]));
Q_FDP0UA U3142 ( .D(n5671), .QTFCLK( ), .Q(xdata[525]));
Q_FDP0UA U3143 ( .D(n5672), .QTFCLK( ), .Q(xdata[526]));
Q_FDP0UA U3144 ( .D(n5673), .QTFCLK( ), .Q(xdata[527]));
Q_FDP0UA U3145 ( .D(n5674), .QTFCLK( ), .Q(xdata[528]));
Q_FDP0UA U3146 ( .D(n5675), .QTFCLK( ), .Q(xdata[529]));
Q_FDP0UA U3147 ( .D(n5676), .QTFCLK( ), .Q(xdata[530]));
Q_FDP0UA U3148 ( .D(n5677), .QTFCLK( ), .Q(xdata[531]));
Q_FDP0UA U3149 ( .D(n5678), .QTFCLK( ), .Q(xdata[532]));
Q_FDP0UA U3150 ( .D(n5679), .QTFCLK( ), .Q(xdata[533]));
Q_FDP0UA U3151 ( .D(n5680), .QTFCLK( ), .Q(xdata[534]));
Q_FDP0UA U3152 ( .D(n5681), .QTFCLK( ), .Q(xdata[535]));
Q_FDP0UA U3153 ( .D(n5682), .QTFCLK( ), .Q(xdata[536]));
Q_FDP0UA U3154 ( .D(n5683), .QTFCLK( ), .Q(xdata[537]));
Q_FDP0UA U3155 ( .D(n5684), .QTFCLK( ), .Q(xdata[538]));
Q_FDP0UA U3156 ( .D(n5685), .QTFCLK( ), .Q(xdata[539]));
Q_FDP0UA U3157 ( .D(n5686), .QTFCLK( ), .Q(xdata[540]));
Q_FDP0UA U3158 ( .D(n5687), .QTFCLK( ), .Q(xdata[541]));
Q_FDP0UA U3159 ( .D(n5688), .QTFCLK( ), .Q(xdata[542]));
Q_FDP0UA U3160 ( .D(n5689), .QTFCLK( ), .Q(xdata[543]));
Q_MX02 U3161 ( .S(n5808), .A0(n5690), .A1(rSync), .Z(n5729));
Q_FDP0UA U3162 ( .D(n5729), .QTFCLK( ), .Q(rSync));
Q_MX02 U3163 ( .S(n5807), .A0(n3862), .A1(n5727), .Z(n5728));
Q_AN02 U3164 ( .A0(n5817), .A1(n3894), .Z(n5727));
Q_MX02 U3165 ( .S(n5807), .A0(n3860), .A1(n5725), .Z(n5726));
Q_AN02 U3166 ( .A0(n5817), .A1(n3892), .Z(n5725));
Q_MX02 U3167 ( .S(n5807), .A0(n3858), .A1(n5723), .Z(n5724));
Q_AN02 U3168 ( .A0(n5817), .A1(n3890), .Z(n5723));
Q_MX02 U3169 ( .S(n5807), .A0(n3856), .A1(n5721), .Z(n5722));
Q_AN02 U3170 ( .A0(n5817), .A1(n3888), .Z(n5721));
Q_MX02 U3171 ( .S(n5807), .A0(n3854), .A1(n5719), .Z(n5720));
Q_AN02 U3172 ( .A0(n5817), .A1(n3886), .Z(n5719));
Q_MX02 U3173 ( .S(n5807), .A0(n3852), .A1(n5717), .Z(n5718));
Q_AN02 U3174 ( .A0(n5817), .A1(n3884), .Z(n5717));
Q_MX02 U3175 ( .S(n5807), .A0(n3850), .A1(n5715), .Z(n5716));
Q_AN02 U3176 ( .A0(n5817), .A1(n3882), .Z(n5715));
Q_MX02 U3177 ( .S(n5807), .A0(n3848), .A1(n5713), .Z(n5714));
Q_AN02 U3178 ( .A0(n5817), .A1(n3880), .Z(n5713));
Q_MX02 U3179 ( .S(n5807), .A0(n3846), .A1(n5711), .Z(n5712));
Q_AN02 U3180 ( .A0(n5817), .A1(n3879), .Z(n5711));
Q_MX02 U3181 ( .S(n5807), .A0(n3844), .A1(n5709), .Z(n5710));
Q_AN02 U3182 ( .A0(n5817), .A1(n3877), .Z(n5709));
Q_MX02 U3183 ( .S(n5807), .A0(n3842), .A1(n5707), .Z(n5708));
Q_AN02 U3184 ( .A0(n5817), .A1(n3876), .Z(n5707));
Q_MX02 U3185 ( .S(n5807), .A0(n3840), .A1(n5705), .Z(n5706));
Q_AN02 U3186 ( .A0(n5817), .A1(n3874), .Z(n5705));
Q_MX02 U3187 ( .S(n5807), .A0(n3838), .A1(n5703), .Z(n5704));
Q_AN02 U3188 ( .A0(n5817), .A1(n3873), .Z(n5703));
Q_MX02 U3189 ( .S(n5807), .A0(n3836), .A1(n5701), .Z(n5702));
Q_AN02 U3190 ( .A0(n5817), .A1(n3871), .Z(n5701));
Q_MX02 U3191 ( .S(n5807), .A0(n3834), .A1(n5699), .Z(n5700));
Q_AN02 U3192 ( .A0(n5817), .A1(n3870), .Z(n5699));
Q_MX02 U3193 ( .S(n5807), .A0(n3832), .A1(n5697), .Z(n5698));
Q_AN02 U3194 ( .A0(n5817), .A1(n3868), .Z(n5697));
Q_MX02 U3195 ( .S(n5807), .A0(n3830), .A1(n5695), .Z(n5696));
Q_AN02 U3196 ( .A0(n5817), .A1(n3867), .Z(n5695));
Q_MX02 U3197 ( .S(n5807), .A0(n3828), .A1(n5693), .Z(n5694));
Q_AN02 U3198 ( .A0(n5817), .A1(n3865), .Z(n5693));
Q_MX02 U3199 ( .S(n5807), .A0(n3826), .A1(n5691), .Z(n5692));
Q_AN02 U3200 ( .A0(n5817), .A1(n3863), .Z(n5691));
Q_AN02 U3201 ( .A0(n6720), .A1(wSync), .Z(n5690));
Q_MX02 U3202 ( .S(n5817), .A0(n5656), .A1(n4407), .Z(n5657));
Q_AN02 U3203 ( .A0(n5818), .A1(GFidata[511]), .Z(n5656));
Q_MX02 U3204 ( .S(n5817), .A0(n5654), .A1(n4406), .Z(n5655));
Q_AN02 U3205 ( .A0(n5818), .A1(GFidata[510]), .Z(n5654));
Q_MX02 U3206 ( .S(n5817), .A0(n5652), .A1(n4405), .Z(n5653));
Q_AN02 U3207 ( .A0(n5818), .A1(GFidata[509]), .Z(n5652));
Q_MX02 U3208 ( .S(n5817), .A0(n5650), .A1(n4404), .Z(n5651));
Q_AN02 U3209 ( .A0(n5818), .A1(GFidata[508]), .Z(n5650));
Q_MX02 U3210 ( .S(n5817), .A0(n5648), .A1(n4403), .Z(n5649));
Q_AN02 U3211 ( .A0(n5818), .A1(GFidata[507]), .Z(n5648));
Q_MX02 U3212 ( .S(n5817), .A0(n5646), .A1(n4402), .Z(n5647));
Q_AN02 U3213 ( .A0(n5818), .A1(GFidata[506]), .Z(n5646));
Q_MX02 U3214 ( .S(n5817), .A0(n5644), .A1(n4401), .Z(n5645));
Q_AN02 U3215 ( .A0(n5818), .A1(GFidata[505]), .Z(n5644));
Q_MX02 U3216 ( .S(n5817), .A0(n5642), .A1(n4400), .Z(n5643));
Q_AN02 U3217 ( .A0(n5818), .A1(GFidata[504]), .Z(n5642));
Q_MX02 U3218 ( .S(n5817), .A0(n5640), .A1(n4399), .Z(n5641));
Q_AN02 U3219 ( .A0(n5818), .A1(GFidata[503]), .Z(n5640));
Q_MX02 U3220 ( .S(n5817), .A0(n5638), .A1(n4398), .Z(n5639));
Q_AN02 U3221 ( .A0(n5818), .A1(GFidata[502]), .Z(n5638));
Q_MX02 U3222 ( .S(n5817), .A0(n5636), .A1(n4397), .Z(n5637));
Q_AN02 U3223 ( .A0(n5818), .A1(GFidata[501]), .Z(n5636));
Q_MX02 U3224 ( .S(n5817), .A0(n5634), .A1(n4396), .Z(n5635));
Q_AN02 U3225 ( .A0(n5818), .A1(GFidata[500]), .Z(n5634));
Q_MX02 U3226 ( .S(n5817), .A0(n5632), .A1(n4395), .Z(n5633));
Q_AN02 U3227 ( .A0(n5818), .A1(GFidata[499]), .Z(n5632));
Q_MX02 U3228 ( .S(n5817), .A0(n5630), .A1(n4394), .Z(n5631));
Q_AN02 U3229 ( .A0(n5818), .A1(GFidata[498]), .Z(n5630));
Q_MX02 U3230 ( .S(n5817), .A0(n5628), .A1(n4393), .Z(n5629));
Q_AN02 U3231 ( .A0(n5818), .A1(GFidata[497]), .Z(n5628));
Q_MX02 U3232 ( .S(n5817), .A0(n5626), .A1(n4392), .Z(n5627));
Q_AN02 U3233 ( .A0(n5818), .A1(GFidata[496]), .Z(n5626));
Q_MX02 U3234 ( .S(n5817), .A0(n5624), .A1(n4391), .Z(n5625));
Q_AN02 U3235 ( .A0(n5818), .A1(GFidata[495]), .Z(n5624));
Q_MX02 U3236 ( .S(n5817), .A0(n5622), .A1(n4390), .Z(n5623));
Q_AN02 U3237 ( .A0(n5818), .A1(GFidata[494]), .Z(n5622));
Q_MX02 U3238 ( .S(n5817), .A0(n5620), .A1(n4389), .Z(n5621));
Q_AN02 U3239 ( .A0(n5818), .A1(GFidata[493]), .Z(n5620));
Q_MX02 U3240 ( .S(n5817), .A0(n5618), .A1(n4388), .Z(n5619));
Q_AN02 U3241 ( .A0(n5818), .A1(GFidata[492]), .Z(n5618));
Q_MX02 U3242 ( .S(n5817), .A0(n5616), .A1(n4387), .Z(n5617));
Q_AN02 U3243 ( .A0(n5818), .A1(GFidata[491]), .Z(n5616));
Q_MX02 U3244 ( .S(n5817), .A0(n5614), .A1(n4386), .Z(n5615));
Q_AN02 U3245 ( .A0(n5818), .A1(GFidata[490]), .Z(n5614));
Q_MX02 U3246 ( .S(n5817), .A0(n5612), .A1(n4385), .Z(n5613));
Q_AN02 U3247 ( .A0(n5818), .A1(GFidata[489]), .Z(n5612));
Q_MX02 U3248 ( .S(n5817), .A0(n5610), .A1(n4384), .Z(n5611));
Q_AN02 U3249 ( .A0(n5818), .A1(GFidata[488]), .Z(n5610));
Q_MX02 U3250 ( .S(n5817), .A0(n5608), .A1(n4383), .Z(n5609));
Q_AN02 U3251 ( .A0(n5818), .A1(GFidata[487]), .Z(n5608));
Q_MX02 U3252 ( .S(n5817), .A0(n5606), .A1(n4382), .Z(n5607));
Q_AN02 U3253 ( .A0(n5818), .A1(GFidata[486]), .Z(n5606));
Q_MX02 U3254 ( .S(n5817), .A0(n5604), .A1(n4381), .Z(n5605));
Q_AN02 U3255 ( .A0(n5818), .A1(GFidata[485]), .Z(n5604));
Q_MX02 U3256 ( .S(n5817), .A0(n5602), .A1(n4380), .Z(n5603));
Q_AN02 U3257 ( .A0(n5818), .A1(GFidata[484]), .Z(n5602));
Q_MX02 U3258 ( .S(n5817), .A0(n5600), .A1(n4379), .Z(n5601));
Q_AN02 U3259 ( .A0(n5818), .A1(GFidata[483]), .Z(n5600));
Q_MX02 U3260 ( .S(n5817), .A0(n5598), .A1(n4378), .Z(n5599));
Q_AN02 U3261 ( .A0(n5818), .A1(GFidata[482]), .Z(n5598));
Q_MX02 U3262 ( .S(n5817), .A0(n5596), .A1(n4377), .Z(n5597));
Q_AN02 U3263 ( .A0(n5818), .A1(GFidata[481]), .Z(n5596));
Q_MX02 U3264 ( .S(n5817), .A0(n5594), .A1(n4376), .Z(n5595));
Q_AN02 U3265 ( .A0(n5818), .A1(GFidata[480]), .Z(n5594));
Q_MX02 U3266 ( .S(n5817), .A0(n5592), .A1(n4375), .Z(n5593));
Q_AN02 U3267 ( .A0(n5818), .A1(GFidata[479]), .Z(n5592));
Q_MX02 U3268 ( .S(n5817), .A0(n5590), .A1(n4374), .Z(n5591));
Q_AN02 U3269 ( .A0(n5818), .A1(GFidata[478]), .Z(n5590));
Q_MX02 U3270 ( .S(n5817), .A0(n5588), .A1(n4373), .Z(n5589));
Q_AN02 U3271 ( .A0(n5818), .A1(GFidata[477]), .Z(n5588));
Q_MX02 U3272 ( .S(n5817), .A0(n5586), .A1(n4372), .Z(n5587));
Q_AN02 U3273 ( .A0(n5818), .A1(GFidata[476]), .Z(n5586));
Q_MX02 U3274 ( .S(n5817), .A0(n5584), .A1(n4371), .Z(n5585));
Q_AN02 U3275 ( .A0(n5818), .A1(GFidata[475]), .Z(n5584));
Q_MX02 U3276 ( .S(n5817), .A0(n5582), .A1(n4370), .Z(n5583));
Q_AN02 U3277 ( .A0(n5818), .A1(GFidata[474]), .Z(n5582));
Q_MX02 U3278 ( .S(n5817), .A0(n5580), .A1(n4369), .Z(n5581));
Q_AN02 U3279 ( .A0(n5818), .A1(GFidata[473]), .Z(n5580));
Q_MX02 U3280 ( .S(n5817), .A0(n5578), .A1(n4368), .Z(n5579));
Q_AN02 U3281 ( .A0(n5818), .A1(GFidata[472]), .Z(n5578));
Q_MX02 U3282 ( .S(n5817), .A0(n5576), .A1(n4367), .Z(n5577));
Q_AN02 U3283 ( .A0(n5818), .A1(GFidata[471]), .Z(n5576));
Q_MX02 U3284 ( .S(n5817), .A0(n5574), .A1(n4366), .Z(n5575));
Q_AN02 U3285 ( .A0(n5818), .A1(GFidata[470]), .Z(n5574));
Q_MX02 U3286 ( .S(n5817), .A0(n5572), .A1(n4365), .Z(n5573));
Q_AN02 U3287 ( .A0(n5818), .A1(GFidata[469]), .Z(n5572));
Q_MX02 U3288 ( .S(n5817), .A0(n5570), .A1(n4364), .Z(n5571));
Q_AN02 U3289 ( .A0(n5818), .A1(GFidata[468]), .Z(n5570));
Q_MX02 U3290 ( .S(n5817), .A0(n5568), .A1(n4363), .Z(n5569));
Q_AN02 U3291 ( .A0(n5818), .A1(GFidata[467]), .Z(n5568));
Q_MX02 U3292 ( .S(n5817), .A0(n5566), .A1(n4362), .Z(n5567));
Q_AN02 U3293 ( .A0(n5818), .A1(GFidata[466]), .Z(n5566));
Q_MX02 U3294 ( .S(n5817), .A0(n5564), .A1(n4361), .Z(n5565));
Q_AN02 U3295 ( .A0(n5818), .A1(GFidata[465]), .Z(n5564));
Q_MX02 U3296 ( .S(n5817), .A0(n5562), .A1(n4360), .Z(n5563));
Q_AN02 U3297 ( .A0(n5818), .A1(GFidata[464]), .Z(n5562));
Q_MX02 U3298 ( .S(n5817), .A0(n5560), .A1(n4359), .Z(n5561));
Q_AN02 U3299 ( .A0(n5818), .A1(GFidata[463]), .Z(n5560));
Q_MX02 U3300 ( .S(n5817), .A0(n5558), .A1(n4358), .Z(n5559));
Q_AN02 U3301 ( .A0(n5818), .A1(GFidata[462]), .Z(n5558));
Q_MX02 U3302 ( .S(n5817), .A0(n5556), .A1(n4357), .Z(n5557));
Q_AN02 U3303 ( .A0(n5818), .A1(GFidata[461]), .Z(n5556));
Q_MX02 U3304 ( .S(n5817), .A0(n5554), .A1(n4356), .Z(n5555));
Q_AN02 U3305 ( .A0(n5818), .A1(GFidata[460]), .Z(n5554));
Q_MX02 U3306 ( .S(n5817), .A0(n5552), .A1(n4355), .Z(n5553));
Q_AN02 U3307 ( .A0(n5818), .A1(GFidata[459]), .Z(n5552));
Q_MX02 U3308 ( .S(n5817), .A0(n5550), .A1(n4354), .Z(n5551));
Q_AN02 U3309 ( .A0(n5818), .A1(GFidata[458]), .Z(n5550));
Q_MX02 U3310 ( .S(n5817), .A0(n5548), .A1(n4353), .Z(n5549));
Q_AN02 U3311 ( .A0(n5818), .A1(GFidata[457]), .Z(n5548));
Q_MX02 U3312 ( .S(n5817), .A0(n5546), .A1(n4352), .Z(n5547));
Q_AN02 U3313 ( .A0(n5818), .A1(GFidata[456]), .Z(n5546));
Q_MX02 U3314 ( .S(n5817), .A0(n5544), .A1(n4351), .Z(n5545));
Q_AN02 U3315 ( .A0(n5818), .A1(GFidata[455]), .Z(n5544));
Q_MX02 U3316 ( .S(n5817), .A0(n5542), .A1(n4350), .Z(n5543));
Q_AN02 U3317 ( .A0(n5818), .A1(GFidata[454]), .Z(n5542));
Q_MX02 U3318 ( .S(n5817), .A0(n5540), .A1(n4349), .Z(n5541));
Q_AN02 U3319 ( .A0(n5818), .A1(GFidata[453]), .Z(n5540));
Q_MX02 U3320 ( .S(n5817), .A0(n5538), .A1(n4348), .Z(n5539));
Q_AN02 U3321 ( .A0(n5818), .A1(GFidata[452]), .Z(n5538));
Q_MX02 U3322 ( .S(n5817), .A0(n5536), .A1(n4347), .Z(n5537));
Q_AN02 U3323 ( .A0(n5818), .A1(GFidata[451]), .Z(n5536));
Q_MX02 U3324 ( .S(n5817), .A0(n5534), .A1(n4346), .Z(n5535));
Q_AN02 U3325 ( .A0(n5818), .A1(GFidata[450]), .Z(n5534));
Q_MX02 U3326 ( .S(n5817), .A0(n5532), .A1(n4345), .Z(n5533));
Q_AN02 U3327 ( .A0(n5818), .A1(GFidata[449]), .Z(n5532));
Q_MX02 U3328 ( .S(n5817), .A0(n5530), .A1(n4344), .Z(n5531));
Q_AN02 U3329 ( .A0(n5818), .A1(GFidata[448]), .Z(n5530));
Q_MX02 U3330 ( .S(n5817), .A0(n5528), .A1(n4343), .Z(n5529));
Q_AN02 U3331 ( .A0(n5818), .A1(GFidata[447]), .Z(n5528));
Q_MX02 U3332 ( .S(n5817), .A0(n5526), .A1(n4342), .Z(n5527));
Q_AN02 U3333 ( .A0(n5818), .A1(GFidata[446]), .Z(n5526));
Q_MX02 U3334 ( .S(n5817), .A0(n5524), .A1(n4341), .Z(n5525));
Q_AN02 U3335 ( .A0(n5818), .A1(GFidata[445]), .Z(n5524));
Q_MX02 U3336 ( .S(n5817), .A0(n5522), .A1(n4340), .Z(n5523));
Q_AN02 U3337 ( .A0(n5818), .A1(GFidata[444]), .Z(n5522));
Q_MX02 U3338 ( .S(n5817), .A0(n5520), .A1(n4339), .Z(n5521));
Q_AN02 U3339 ( .A0(n5818), .A1(GFidata[443]), .Z(n5520));
Q_MX02 U3340 ( .S(n5817), .A0(n5518), .A1(n4338), .Z(n5519));
Q_AN02 U3341 ( .A0(n5818), .A1(GFidata[442]), .Z(n5518));
Q_MX02 U3342 ( .S(n5817), .A0(n5516), .A1(n4337), .Z(n5517));
Q_AN02 U3343 ( .A0(n5818), .A1(GFidata[441]), .Z(n5516));
Q_MX02 U3344 ( .S(n5817), .A0(n5514), .A1(n4336), .Z(n5515));
Q_AN02 U3345 ( .A0(n5818), .A1(GFidata[440]), .Z(n5514));
Q_MX02 U3346 ( .S(n5817), .A0(n5512), .A1(n4335), .Z(n5513));
Q_AN02 U3347 ( .A0(n5818), .A1(GFidata[439]), .Z(n5512));
Q_MX02 U3348 ( .S(n5817), .A0(n5510), .A1(n4334), .Z(n5511));
Q_AN02 U3349 ( .A0(n5818), .A1(GFidata[438]), .Z(n5510));
Q_MX02 U3350 ( .S(n5817), .A0(n5508), .A1(n4333), .Z(n5509));
Q_AN02 U3351 ( .A0(n5818), .A1(GFidata[437]), .Z(n5508));
Q_MX02 U3352 ( .S(n5817), .A0(n5506), .A1(n4332), .Z(n5507));
Q_AN02 U3353 ( .A0(n5818), .A1(GFidata[436]), .Z(n5506));
Q_MX02 U3354 ( .S(n5817), .A0(n5504), .A1(n4331), .Z(n5505));
Q_AN02 U3355 ( .A0(n5818), .A1(GFidata[435]), .Z(n5504));
Q_MX02 U3356 ( .S(n5817), .A0(n5502), .A1(n4330), .Z(n5503));
Q_AN02 U3357 ( .A0(n5818), .A1(GFidata[434]), .Z(n5502));
Q_MX02 U3358 ( .S(n5817), .A0(n5500), .A1(n4329), .Z(n5501));
Q_AN02 U3359 ( .A0(n5818), .A1(GFidata[433]), .Z(n5500));
Q_MX02 U3360 ( .S(n5817), .A0(n5498), .A1(n4328), .Z(n5499));
Q_AN02 U3361 ( .A0(n5818), .A1(GFidata[432]), .Z(n5498));
Q_MX02 U3362 ( .S(n5817), .A0(n5496), .A1(n4327), .Z(n5497));
Q_AN02 U3363 ( .A0(n5818), .A1(GFidata[431]), .Z(n5496));
Q_MX02 U3364 ( .S(n5817), .A0(n5494), .A1(n4326), .Z(n5495));
Q_AN02 U3365 ( .A0(n5818), .A1(GFidata[430]), .Z(n5494));
Q_MX02 U3366 ( .S(n5817), .A0(n5492), .A1(n4325), .Z(n5493));
Q_AN02 U3367 ( .A0(n5818), .A1(GFidata[429]), .Z(n5492));
Q_MX02 U3368 ( .S(n5817), .A0(n5490), .A1(n4324), .Z(n5491));
Q_AN02 U3369 ( .A0(n5818), .A1(GFidata[428]), .Z(n5490));
Q_MX02 U3370 ( .S(n5817), .A0(n5488), .A1(n4323), .Z(n5489));
Q_AN02 U3371 ( .A0(n5818), .A1(GFidata[427]), .Z(n5488));
Q_MX02 U3372 ( .S(n5817), .A0(n5486), .A1(n4322), .Z(n5487));
Q_AN02 U3373 ( .A0(n5818), .A1(GFidata[426]), .Z(n5486));
Q_MX02 U3374 ( .S(n5817), .A0(n5484), .A1(n4321), .Z(n5485));
Q_AN02 U3375 ( .A0(n5818), .A1(GFidata[425]), .Z(n5484));
Q_MX02 U3376 ( .S(n5817), .A0(n5482), .A1(n4320), .Z(n5483));
Q_AN02 U3377 ( .A0(n5818), .A1(GFidata[424]), .Z(n5482));
Q_MX02 U3378 ( .S(n5817), .A0(n5480), .A1(n4319), .Z(n5481));
Q_AN02 U3379 ( .A0(n5818), .A1(GFidata[423]), .Z(n5480));
Q_MX02 U3380 ( .S(n5817), .A0(n5478), .A1(n4318), .Z(n5479));
Q_AN02 U3381 ( .A0(n5818), .A1(GFidata[422]), .Z(n5478));
Q_MX02 U3382 ( .S(n5817), .A0(n5476), .A1(n4317), .Z(n5477));
Q_AN02 U3383 ( .A0(n5818), .A1(GFidata[421]), .Z(n5476));
Q_MX02 U3384 ( .S(n5817), .A0(n5474), .A1(n4316), .Z(n5475));
Q_AN02 U3385 ( .A0(n5818), .A1(GFidata[420]), .Z(n5474));
Q_MX02 U3386 ( .S(n5817), .A0(n5472), .A1(n4315), .Z(n5473));
Q_AN02 U3387 ( .A0(n5818), .A1(GFidata[419]), .Z(n5472));
Q_MX02 U3388 ( .S(n5817), .A0(n5470), .A1(n4314), .Z(n5471));
Q_AN02 U3389 ( .A0(n5818), .A1(GFidata[418]), .Z(n5470));
Q_MX02 U3390 ( .S(n5817), .A0(n5468), .A1(n4313), .Z(n5469));
Q_AN02 U3391 ( .A0(n5818), .A1(GFidata[417]), .Z(n5468));
Q_MX02 U3392 ( .S(n5817), .A0(n5466), .A1(n4312), .Z(n5467));
Q_AN02 U3393 ( .A0(n5818), .A1(GFidata[416]), .Z(n5466));
Q_MX02 U3394 ( .S(n5817), .A0(n5464), .A1(n4311), .Z(n5465));
Q_AN02 U3395 ( .A0(n5818), .A1(GFidata[415]), .Z(n5464));
Q_MX02 U3396 ( .S(n5817), .A0(n5462), .A1(n4310), .Z(n5463));
Q_AN02 U3397 ( .A0(n5818), .A1(GFidata[414]), .Z(n5462));
Q_MX02 U3398 ( .S(n5817), .A0(n5460), .A1(n4309), .Z(n5461));
Q_AN02 U3399 ( .A0(n5818), .A1(GFidata[413]), .Z(n5460));
Q_MX02 U3400 ( .S(n5817), .A0(n5458), .A1(n4308), .Z(n5459));
Q_AN02 U3401 ( .A0(n5818), .A1(GFidata[412]), .Z(n5458));
Q_MX02 U3402 ( .S(n5817), .A0(n5456), .A1(n4307), .Z(n5457));
Q_AN02 U3403 ( .A0(n5818), .A1(GFidata[411]), .Z(n5456));
Q_MX02 U3404 ( .S(n5817), .A0(n5454), .A1(n4306), .Z(n5455));
Q_AN02 U3405 ( .A0(n5818), .A1(GFidata[410]), .Z(n5454));
Q_MX02 U3406 ( .S(n5817), .A0(n5452), .A1(n4305), .Z(n5453));
Q_AN02 U3407 ( .A0(n5818), .A1(GFidata[409]), .Z(n5452));
Q_MX02 U3408 ( .S(n5817), .A0(n5450), .A1(n4304), .Z(n5451));
Q_AN02 U3409 ( .A0(n5818), .A1(GFidata[408]), .Z(n5450));
Q_MX02 U3410 ( .S(n5817), .A0(n5448), .A1(n4303), .Z(n5449));
Q_AN02 U3411 ( .A0(n5818), .A1(GFidata[407]), .Z(n5448));
Q_MX02 U3412 ( .S(n5817), .A0(n5446), .A1(n4302), .Z(n5447));
Q_AN02 U3413 ( .A0(n5818), .A1(GFidata[406]), .Z(n5446));
Q_MX02 U3414 ( .S(n5817), .A0(n5444), .A1(n4301), .Z(n5445));
Q_AN02 U3415 ( .A0(n5818), .A1(GFidata[405]), .Z(n5444));
Q_MX02 U3416 ( .S(n5817), .A0(n5442), .A1(n4300), .Z(n5443));
Q_AN02 U3417 ( .A0(n5818), .A1(GFidata[404]), .Z(n5442));
Q_MX02 U3418 ( .S(n5817), .A0(n5440), .A1(n4299), .Z(n5441));
Q_AN02 U3419 ( .A0(n5818), .A1(GFidata[403]), .Z(n5440));
Q_MX02 U3420 ( .S(n5817), .A0(n5438), .A1(n4298), .Z(n5439));
Q_AN02 U3421 ( .A0(n5818), .A1(GFidata[402]), .Z(n5438));
Q_MX02 U3422 ( .S(n5817), .A0(n5436), .A1(n4297), .Z(n5437));
Q_AN02 U3423 ( .A0(n5818), .A1(GFidata[401]), .Z(n5436));
Q_MX02 U3424 ( .S(n5817), .A0(n5434), .A1(n4296), .Z(n5435));
Q_AN02 U3425 ( .A0(n5818), .A1(GFidata[400]), .Z(n5434));
Q_MX02 U3426 ( .S(n5817), .A0(n5432), .A1(n4295), .Z(n5433));
Q_AN02 U3427 ( .A0(n5818), .A1(GFidata[399]), .Z(n5432));
Q_MX02 U3428 ( .S(n5817), .A0(n5430), .A1(n4294), .Z(n5431));
Q_AN02 U3429 ( .A0(n5818), .A1(GFidata[398]), .Z(n5430));
Q_MX02 U3430 ( .S(n5817), .A0(n5428), .A1(n4293), .Z(n5429));
Q_AN02 U3431 ( .A0(n5818), .A1(GFidata[397]), .Z(n5428));
Q_MX02 U3432 ( .S(n5817), .A0(n5426), .A1(n4292), .Z(n5427));
Q_AN02 U3433 ( .A0(n5818), .A1(GFidata[396]), .Z(n5426));
Q_MX02 U3434 ( .S(n5817), .A0(n5424), .A1(n4291), .Z(n5425));
Q_AN02 U3435 ( .A0(n5818), .A1(GFidata[395]), .Z(n5424));
Q_MX02 U3436 ( .S(n5817), .A0(n5422), .A1(n4290), .Z(n5423));
Q_AN02 U3437 ( .A0(n5818), .A1(GFidata[394]), .Z(n5422));
Q_MX02 U3438 ( .S(n5817), .A0(n5420), .A1(n4289), .Z(n5421));
Q_AN02 U3439 ( .A0(n5818), .A1(GFidata[393]), .Z(n5420));
Q_MX02 U3440 ( .S(n5817), .A0(n5418), .A1(n4288), .Z(n5419));
Q_AN02 U3441 ( .A0(n5818), .A1(GFidata[392]), .Z(n5418));
Q_MX02 U3442 ( .S(n5817), .A0(n5416), .A1(n4287), .Z(n5417));
Q_AN02 U3443 ( .A0(n5818), .A1(GFidata[391]), .Z(n5416));
Q_MX02 U3444 ( .S(n5817), .A0(n5414), .A1(n4286), .Z(n5415));
Q_AN02 U3445 ( .A0(n5818), .A1(GFidata[390]), .Z(n5414));
Q_MX02 U3446 ( .S(n5817), .A0(n5412), .A1(n4285), .Z(n5413));
Q_AN02 U3447 ( .A0(n5818), .A1(GFidata[389]), .Z(n5412));
Q_MX02 U3448 ( .S(n5817), .A0(n5410), .A1(n4284), .Z(n5411));
Q_AN02 U3449 ( .A0(n5818), .A1(GFidata[388]), .Z(n5410));
Q_MX02 U3450 ( .S(n5817), .A0(n5408), .A1(n4283), .Z(n5409));
Q_AN02 U3451 ( .A0(n5818), .A1(GFidata[387]), .Z(n5408));
Q_MX02 U3452 ( .S(n5817), .A0(n5406), .A1(n4282), .Z(n5407));
Q_AN02 U3453 ( .A0(n5818), .A1(GFidata[386]), .Z(n5406));
Q_MX02 U3454 ( .S(n5817), .A0(n5404), .A1(n4281), .Z(n5405));
Q_AN02 U3455 ( .A0(n5818), .A1(GFidata[385]), .Z(n5404));
Q_MX02 U3456 ( .S(n5817), .A0(n5402), .A1(n4280), .Z(n5403));
Q_AN02 U3457 ( .A0(n5818), .A1(GFidata[384]), .Z(n5402));
Q_MX02 U3458 ( .S(n5817), .A0(n5400), .A1(n4279), .Z(n5401));
Q_AN02 U3459 ( .A0(n5818), .A1(GFidata[383]), .Z(n5400));
Q_MX02 U3460 ( .S(n5817), .A0(n5398), .A1(n4278), .Z(n5399));
Q_AN02 U3461 ( .A0(n5818), .A1(GFidata[382]), .Z(n5398));
Q_MX02 U3462 ( .S(n5817), .A0(n5396), .A1(n4277), .Z(n5397));
Q_AN02 U3463 ( .A0(n5818), .A1(GFidata[381]), .Z(n5396));
Q_MX02 U3464 ( .S(n5817), .A0(n5394), .A1(n4276), .Z(n5395));
Q_AN02 U3465 ( .A0(n5818), .A1(GFidata[380]), .Z(n5394));
Q_MX02 U3466 ( .S(n5817), .A0(n5392), .A1(n4275), .Z(n5393));
Q_AN02 U3467 ( .A0(n5818), .A1(GFidata[379]), .Z(n5392));
Q_MX02 U3468 ( .S(n5817), .A0(n5390), .A1(n4274), .Z(n5391));
Q_AN02 U3469 ( .A0(n5818), .A1(GFidata[378]), .Z(n5390));
Q_MX02 U3470 ( .S(n5817), .A0(n5388), .A1(n4273), .Z(n5389));
Q_AN02 U3471 ( .A0(n5818), .A1(GFidata[377]), .Z(n5388));
Q_MX02 U3472 ( .S(n5817), .A0(n5386), .A1(n4272), .Z(n5387));
Q_AN02 U3473 ( .A0(n5818), .A1(GFidata[376]), .Z(n5386));
Q_MX02 U3474 ( .S(n5817), .A0(n5384), .A1(n4271), .Z(n5385));
Q_AN02 U3475 ( .A0(n5818), .A1(GFidata[375]), .Z(n5384));
Q_MX02 U3476 ( .S(n5817), .A0(n5382), .A1(n4270), .Z(n5383));
Q_AN02 U3477 ( .A0(n5818), .A1(GFidata[374]), .Z(n5382));
Q_MX02 U3478 ( .S(n5817), .A0(n5380), .A1(n4269), .Z(n5381));
Q_AN02 U3479 ( .A0(n5818), .A1(GFidata[373]), .Z(n5380));
Q_MX02 U3480 ( .S(n5817), .A0(n5378), .A1(n4268), .Z(n5379));
Q_AN02 U3481 ( .A0(n5818), .A1(GFidata[372]), .Z(n5378));
Q_MX02 U3482 ( .S(n5817), .A0(n5376), .A1(n4267), .Z(n5377));
Q_AN02 U3483 ( .A0(n5818), .A1(GFidata[371]), .Z(n5376));
Q_MX02 U3484 ( .S(n5817), .A0(n5374), .A1(n4266), .Z(n5375));
Q_AN02 U3485 ( .A0(n5818), .A1(GFidata[370]), .Z(n5374));
Q_MX02 U3486 ( .S(n5817), .A0(n5372), .A1(n4265), .Z(n5373));
Q_AN02 U3487 ( .A0(n5818), .A1(GFidata[369]), .Z(n5372));
Q_MX02 U3488 ( .S(n5817), .A0(n5370), .A1(n4264), .Z(n5371));
Q_AN02 U3489 ( .A0(n5818), .A1(GFidata[368]), .Z(n5370));
Q_MX02 U3490 ( .S(n5817), .A0(n5368), .A1(n4263), .Z(n5369));
Q_AN02 U3491 ( .A0(n5818), .A1(GFidata[367]), .Z(n5368));
Q_MX02 U3492 ( .S(n5817), .A0(n5366), .A1(n4262), .Z(n5367));
Q_AN02 U3493 ( .A0(n5818), .A1(GFidata[366]), .Z(n5366));
Q_MX02 U3494 ( .S(n5817), .A0(n5364), .A1(n4261), .Z(n5365));
Q_AN02 U3495 ( .A0(n5818), .A1(GFidata[365]), .Z(n5364));
Q_MX02 U3496 ( .S(n5817), .A0(n5362), .A1(n4260), .Z(n5363));
Q_AN02 U3497 ( .A0(n5818), .A1(GFidata[364]), .Z(n5362));
Q_MX02 U3498 ( .S(n5817), .A0(n5360), .A1(n4259), .Z(n5361));
Q_AN02 U3499 ( .A0(n5818), .A1(GFidata[363]), .Z(n5360));
Q_MX02 U3500 ( .S(n5817), .A0(n5358), .A1(n4258), .Z(n5359));
Q_AN02 U3501 ( .A0(n5818), .A1(GFidata[362]), .Z(n5358));
Q_MX02 U3502 ( .S(n5817), .A0(n5356), .A1(n4257), .Z(n5357));
Q_AN02 U3503 ( .A0(n5818), .A1(GFidata[361]), .Z(n5356));
Q_MX02 U3504 ( .S(n5817), .A0(n5354), .A1(n4256), .Z(n5355));
Q_AN02 U3505 ( .A0(n5818), .A1(GFidata[360]), .Z(n5354));
Q_MX02 U3506 ( .S(n5817), .A0(n5352), .A1(n4255), .Z(n5353));
Q_AN02 U3507 ( .A0(n5818), .A1(GFidata[359]), .Z(n5352));
Q_MX02 U3508 ( .S(n5817), .A0(n5350), .A1(n4254), .Z(n5351));
Q_AN02 U3509 ( .A0(n5818), .A1(GFidata[358]), .Z(n5350));
Q_MX02 U3510 ( .S(n5817), .A0(n5348), .A1(n4253), .Z(n5349));
Q_AN02 U3511 ( .A0(n5818), .A1(GFidata[357]), .Z(n5348));
Q_MX02 U3512 ( .S(n5817), .A0(n5346), .A1(n4252), .Z(n5347));
Q_AN02 U3513 ( .A0(n5818), .A1(GFidata[356]), .Z(n5346));
Q_MX02 U3514 ( .S(n5817), .A0(n5344), .A1(n4251), .Z(n5345));
Q_AN02 U3515 ( .A0(n5818), .A1(GFidata[355]), .Z(n5344));
Q_MX02 U3516 ( .S(n5817), .A0(n5342), .A1(n4250), .Z(n5343));
Q_AN02 U3517 ( .A0(n5818), .A1(GFidata[354]), .Z(n5342));
Q_MX02 U3518 ( .S(n5817), .A0(n5340), .A1(n4249), .Z(n5341));
Q_AN02 U3519 ( .A0(n5818), .A1(GFidata[353]), .Z(n5340));
Q_MX02 U3520 ( .S(n5817), .A0(n5338), .A1(n4248), .Z(n5339));
Q_AN02 U3521 ( .A0(n5818), .A1(GFidata[352]), .Z(n5338));
Q_MX02 U3522 ( .S(n5817), .A0(n5336), .A1(n4247), .Z(n5337));
Q_AN02 U3523 ( .A0(n5818), .A1(GFidata[351]), .Z(n5336));
Q_MX02 U3524 ( .S(n5817), .A0(n5334), .A1(n4246), .Z(n5335));
Q_AN02 U3525 ( .A0(n5818), .A1(GFidata[350]), .Z(n5334));
Q_MX02 U3526 ( .S(n5817), .A0(n5332), .A1(n4245), .Z(n5333));
Q_AN02 U3527 ( .A0(n5818), .A1(GFidata[349]), .Z(n5332));
Q_MX02 U3528 ( .S(n5817), .A0(n5330), .A1(n4244), .Z(n5331));
Q_AN02 U3529 ( .A0(n5818), .A1(GFidata[348]), .Z(n5330));
Q_MX02 U3530 ( .S(n5817), .A0(n5328), .A1(n4243), .Z(n5329));
Q_AN02 U3531 ( .A0(n5818), .A1(GFidata[347]), .Z(n5328));
Q_MX02 U3532 ( .S(n5817), .A0(n5326), .A1(n4242), .Z(n5327));
Q_AN02 U3533 ( .A0(n5818), .A1(GFidata[346]), .Z(n5326));
Q_MX02 U3534 ( .S(n5817), .A0(n5324), .A1(n4241), .Z(n5325));
Q_AN02 U3535 ( .A0(n5818), .A1(GFidata[345]), .Z(n5324));
Q_MX02 U3536 ( .S(n5817), .A0(n5322), .A1(n4240), .Z(n5323));
Q_AN02 U3537 ( .A0(n5818), .A1(GFidata[344]), .Z(n5322));
Q_MX02 U3538 ( .S(n5817), .A0(n5320), .A1(n4239), .Z(n5321));
Q_AN02 U3539 ( .A0(n5818), .A1(GFidata[343]), .Z(n5320));
Q_MX02 U3540 ( .S(n5817), .A0(n5318), .A1(n4238), .Z(n5319));
Q_AN02 U3541 ( .A0(n5818), .A1(GFidata[342]), .Z(n5318));
Q_MX02 U3542 ( .S(n5817), .A0(n5316), .A1(n4237), .Z(n5317));
Q_AN02 U3543 ( .A0(n5818), .A1(GFidata[341]), .Z(n5316));
Q_MX02 U3544 ( .S(n5817), .A0(n5314), .A1(n4236), .Z(n5315));
Q_AN02 U3545 ( .A0(n5818), .A1(GFidata[340]), .Z(n5314));
Q_MX02 U3546 ( .S(n5817), .A0(n5312), .A1(n4235), .Z(n5313));
Q_AN02 U3547 ( .A0(n5818), .A1(GFidata[339]), .Z(n5312));
Q_MX02 U3548 ( .S(n5817), .A0(n5310), .A1(n4234), .Z(n5311));
Q_AN02 U3549 ( .A0(n5818), .A1(GFidata[338]), .Z(n5310));
Q_MX02 U3550 ( .S(n5817), .A0(n5308), .A1(n4233), .Z(n5309));
Q_AN02 U3551 ( .A0(n5818), .A1(GFidata[337]), .Z(n5308));
Q_MX02 U3552 ( .S(n5817), .A0(n5306), .A1(n4232), .Z(n5307));
Q_AN02 U3553 ( .A0(n5818), .A1(GFidata[336]), .Z(n5306));
Q_MX02 U3554 ( .S(n5817), .A0(n5304), .A1(n4231), .Z(n5305));
Q_AN02 U3555 ( .A0(n5818), .A1(GFidata[335]), .Z(n5304));
Q_MX02 U3556 ( .S(n5817), .A0(n5302), .A1(n4230), .Z(n5303));
Q_AN02 U3557 ( .A0(n5818), .A1(GFidata[334]), .Z(n5302));
Q_MX02 U3558 ( .S(n5817), .A0(n5300), .A1(n4229), .Z(n5301));
Q_AN02 U3559 ( .A0(n5818), .A1(GFidata[333]), .Z(n5300));
Q_MX02 U3560 ( .S(n5817), .A0(n5298), .A1(n4228), .Z(n5299));
Q_AN02 U3561 ( .A0(n5818), .A1(GFidata[332]), .Z(n5298));
Q_MX02 U3562 ( .S(n5817), .A0(n5296), .A1(n4227), .Z(n5297));
Q_AN02 U3563 ( .A0(n5818), .A1(GFidata[331]), .Z(n5296));
Q_MX02 U3564 ( .S(n5817), .A0(n5294), .A1(n4226), .Z(n5295));
Q_AN02 U3565 ( .A0(n5818), .A1(GFidata[330]), .Z(n5294));
Q_MX02 U3566 ( .S(n5817), .A0(n5292), .A1(n4225), .Z(n5293));
Q_AN02 U3567 ( .A0(n5818), .A1(GFidata[329]), .Z(n5292));
Q_MX02 U3568 ( .S(n5817), .A0(n5290), .A1(n4224), .Z(n5291));
Q_AN02 U3569 ( .A0(n5818), .A1(GFidata[328]), .Z(n5290));
Q_MX02 U3570 ( .S(n5817), .A0(n5288), .A1(n4223), .Z(n5289));
Q_AN02 U3571 ( .A0(n5818), .A1(GFidata[327]), .Z(n5288));
Q_MX02 U3572 ( .S(n5817), .A0(n5286), .A1(n4222), .Z(n5287));
Q_AN02 U3573 ( .A0(n5818), .A1(GFidata[326]), .Z(n5286));
Q_MX02 U3574 ( .S(n5817), .A0(n5284), .A1(n4221), .Z(n5285));
Q_AN02 U3575 ( .A0(n5818), .A1(GFidata[325]), .Z(n5284));
Q_MX02 U3576 ( .S(n5817), .A0(n5282), .A1(n4220), .Z(n5283));
Q_AN02 U3577 ( .A0(n5818), .A1(GFidata[324]), .Z(n5282));
Q_MX02 U3578 ( .S(n5817), .A0(n5280), .A1(n4219), .Z(n5281));
Q_AN02 U3579 ( .A0(n5818), .A1(GFidata[323]), .Z(n5280));
Q_MX02 U3580 ( .S(n5817), .A0(n5278), .A1(n4218), .Z(n5279));
Q_AN02 U3581 ( .A0(n5818), .A1(GFidata[322]), .Z(n5278));
Q_MX02 U3582 ( .S(n5817), .A0(n5276), .A1(n4217), .Z(n5277));
Q_AN02 U3583 ( .A0(n5818), .A1(GFidata[321]), .Z(n5276));
Q_MX02 U3584 ( .S(n5817), .A0(n5274), .A1(n4216), .Z(n5275));
Q_AN02 U3585 ( .A0(n5818), .A1(GFidata[320]), .Z(n5274));
Q_MX02 U3586 ( .S(n5817), .A0(n5272), .A1(n4215), .Z(n5273));
Q_AN02 U3587 ( .A0(n5818), .A1(GFidata[319]), .Z(n5272));
Q_MX02 U3588 ( .S(n5817), .A0(n5270), .A1(n4214), .Z(n5271));
Q_AN02 U3589 ( .A0(n5818), .A1(GFidata[318]), .Z(n5270));
Q_MX02 U3590 ( .S(n5817), .A0(n5268), .A1(n4213), .Z(n5269));
Q_AN02 U3591 ( .A0(n5818), .A1(GFidata[317]), .Z(n5268));
Q_MX02 U3592 ( .S(n5817), .A0(n5266), .A1(n4212), .Z(n5267));
Q_AN02 U3593 ( .A0(n5818), .A1(GFidata[316]), .Z(n5266));
Q_MX02 U3594 ( .S(n5817), .A0(n5264), .A1(n4211), .Z(n5265));
Q_AN02 U3595 ( .A0(n5818), .A1(GFidata[315]), .Z(n5264));
Q_MX02 U3596 ( .S(n5817), .A0(n5262), .A1(n4210), .Z(n5263));
Q_AN02 U3597 ( .A0(n5818), .A1(GFidata[314]), .Z(n5262));
Q_MX02 U3598 ( .S(n5817), .A0(n5260), .A1(n4209), .Z(n5261));
Q_AN02 U3599 ( .A0(n5818), .A1(GFidata[313]), .Z(n5260));
Q_MX02 U3600 ( .S(n5817), .A0(n5258), .A1(n4208), .Z(n5259));
Q_AN02 U3601 ( .A0(n5818), .A1(GFidata[312]), .Z(n5258));
Q_MX02 U3602 ( .S(n5817), .A0(n5256), .A1(n4207), .Z(n5257));
Q_AN02 U3603 ( .A0(n5818), .A1(GFidata[311]), .Z(n5256));
Q_MX02 U3604 ( .S(n5817), .A0(n5254), .A1(n4206), .Z(n5255));
Q_AN02 U3605 ( .A0(n5818), .A1(GFidata[310]), .Z(n5254));
Q_MX02 U3606 ( .S(n5817), .A0(n5252), .A1(n4205), .Z(n5253));
Q_AN02 U3607 ( .A0(n5818), .A1(GFidata[309]), .Z(n5252));
Q_MX02 U3608 ( .S(n5817), .A0(n5250), .A1(n4204), .Z(n5251));
Q_AN02 U3609 ( .A0(n5818), .A1(GFidata[308]), .Z(n5250));
Q_MX02 U3610 ( .S(n5817), .A0(n5248), .A1(n4203), .Z(n5249));
Q_AN02 U3611 ( .A0(n5818), .A1(GFidata[307]), .Z(n5248));
Q_MX02 U3612 ( .S(n5817), .A0(n5246), .A1(n4202), .Z(n5247));
Q_AN02 U3613 ( .A0(n5818), .A1(GFidata[306]), .Z(n5246));
Q_MX02 U3614 ( .S(n5817), .A0(n5244), .A1(n4201), .Z(n5245));
Q_AN02 U3615 ( .A0(n5818), .A1(GFidata[305]), .Z(n5244));
Q_MX02 U3616 ( .S(n5817), .A0(n5242), .A1(n4200), .Z(n5243));
Q_AN02 U3617 ( .A0(n5818), .A1(GFidata[304]), .Z(n5242));
Q_MX02 U3618 ( .S(n5817), .A0(n5240), .A1(n4199), .Z(n5241));
Q_AN02 U3619 ( .A0(n5818), .A1(GFidata[303]), .Z(n5240));
Q_MX02 U3620 ( .S(n5817), .A0(n5238), .A1(n4198), .Z(n5239));
Q_AN02 U3621 ( .A0(n5818), .A1(GFidata[302]), .Z(n5238));
Q_MX02 U3622 ( .S(n5817), .A0(n5236), .A1(n4197), .Z(n5237));
Q_AN02 U3623 ( .A0(n5818), .A1(GFidata[301]), .Z(n5236));
Q_MX02 U3624 ( .S(n5817), .A0(n5234), .A1(n4196), .Z(n5235));
Q_AN02 U3625 ( .A0(n5818), .A1(GFidata[300]), .Z(n5234));
Q_MX02 U3626 ( .S(n5817), .A0(n5232), .A1(n4195), .Z(n5233));
Q_AN02 U3627 ( .A0(n5818), .A1(GFidata[299]), .Z(n5232));
Q_MX02 U3628 ( .S(n5817), .A0(n5230), .A1(n4194), .Z(n5231));
Q_AN02 U3629 ( .A0(n5818), .A1(GFidata[298]), .Z(n5230));
Q_MX02 U3630 ( .S(n5817), .A0(n5228), .A1(n4193), .Z(n5229));
Q_AN02 U3631 ( .A0(n5818), .A1(GFidata[297]), .Z(n5228));
Q_MX02 U3632 ( .S(n5817), .A0(n5226), .A1(n4192), .Z(n5227));
Q_AN02 U3633 ( .A0(n5818), .A1(GFidata[296]), .Z(n5226));
Q_MX02 U3634 ( .S(n5817), .A0(n5224), .A1(n4191), .Z(n5225));
Q_AN02 U3635 ( .A0(n5818), .A1(GFidata[295]), .Z(n5224));
Q_MX02 U3636 ( .S(n5817), .A0(n5222), .A1(n4190), .Z(n5223));
Q_AN02 U3637 ( .A0(n5818), .A1(GFidata[294]), .Z(n5222));
Q_MX02 U3638 ( .S(n5817), .A0(n5220), .A1(n4189), .Z(n5221));
Q_AN02 U3639 ( .A0(n5818), .A1(GFidata[293]), .Z(n5220));
Q_MX02 U3640 ( .S(n5817), .A0(n5218), .A1(n4188), .Z(n5219));
Q_AN02 U3641 ( .A0(n5818), .A1(GFidata[292]), .Z(n5218));
Q_MX02 U3642 ( .S(n5817), .A0(n5216), .A1(n4187), .Z(n5217));
Q_AN02 U3643 ( .A0(n5818), .A1(GFidata[291]), .Z(n5216));
Q_MX02 U3644 ( .S(n5817), .A0(n5214), .A1(n4186), .Z(n5215));
Q_AN02 U3645 ( .A0(n5818), .A1(GFidata[290]), .Z(n5214));
Q_MX02 U3646 ( .S(n5817), .A0(n5212), .A1(n4185), .Z(n5213));
Q_AN02 U3647 ( .A0(n5818), .A1(GFidata[289]), .Z(n5212));
Q_MX02 U3648 ( .S(n5817), .A0(n5210), .A1(n4184), .Z(n5211));
Q_AN02 U3649 ( .A0(n5818), .A1(GFidata[288]), .Z(n5210));
Q_MX02 U3650 ( .S(n5817), .A0(n5208), .A1(n4183), .Z(n5209));
Q_AN02 U3651 ( .A0(n5818), .A1(GFidata[287]), .Z(n5208));
Q_MX02 U3652 ( .S(n5817), .A0(n5206), .A1(n4182), .Z(n5207));
Q_AN02 U3653 ( .A0(n5818), .A1(GFidata[286]), .Z(n5206));
Q_MX02 U3654 ( .S(n5817), .A0(n5204), .A1(n4181), .Z(n5205));
Q_AN02 U3655 ( .A0(n5818), .A1(GFidata[285]), .Z(n5204));
Q_MX02 U3656 ( .S(n5817), .A0(n5202), .A1(n4180), .Z(n5203));
Q_AN02 U3657 ( .A0(n5818), .A1(GFidata[284]), .Z(n5202));
Q_MX02 U3658 ( .S(n5817), .A0(n5200), .A1(n4179), .Z(n5201));
Q_AN02 U3659 ( .A0(n5818), .A1(GFidata[283]), .Z(n5200));
Q_MX02 U3660 ( .S(n5817), .A0(n5198), .A1(n4178), .Z(n5199));
Q_AN02 U3661 ( .A0(n5818), .A1(GFidata[282]), .Z(n5198));
Q_MX02 U3662 ( .S(n5817), .A0(n5196), .A1(n4177), .Z(n5197));
Q_AN02 U3663 ( .A0(n5818), .A1(GFidata[281]), .Z(n5196));
Q_MX02 U3664 ( .S(n5817), .A0(n5194), .A1(n4176), .Z(n5195));
Q_AN02 U3665 ( .A0(n5818), .A1(GFidata[280]), .Z(n5194));
Q_MX02 U3666 ( .S(n5817), .A0(n5192), .A1(n4175), .Z(n5193));
Q_AN02 U3667 ( .A0(n5818), .A1(GFidata[279]), .Z(n5192));
Q_MX02 U3668 ( .S(n5817), .A0(n5190), .A1(n4174), .Z(n5191));
Q_AN02 U3669 ( .A0(n5818), .A1(GFidata[278]), .Z(n5190));
Q_MX02 U3670 ( .S(n5817), .A0(n5188), .A1(n4173), .Z(n5189));
Q_AN02 U3671 ( .A0(n5818), .A1(GFidata[277]), .Z(n5188));
Q_MX02 U3672 ( .S(n5817), .A0(n5186), .A1(n4172), .Z(n5187));
Q_AN02 U3673 ( .A0(n5818), .A1(GFidata[276]), .Z(n5186));
Q_MX02 U3674 ( .S(n5817), .A0(n5184), .A1(n4171), .Z(n5185));
Q_AN02 U3675 ( .A0(n5818), .A1(GFidata[275]), .Z(n5184));
Q_MX02 U3676 ( .S(n5817), .A0(n5182), .A1(n4170), .Z(n5183));
Q_AN02 U3677 ( .A0(n5818), .A1(GFidata[274]), .Z(n5182));
Q_MX02 U3678 ( .S(n5817), .A0(n5180), .A1(n4169), .Z(n5181));
Q_AN02 U3679 ( .A0(n5818), .A1(GFidata[273]), .Z(n5180));
Q_MX02 U3680 ( .S(n5817), .A0(n5178), .A1(n4168), .Z(n5179));
Q_AN02 U3681 ( .A0(n5818), .A1(GFidata[272]), .Z(n5178));
Q_MX02 U3682 ( .S(n5817), .A0(n5176), .A1(n4167), .Z(n5177));
Q_AN02 U3683 ( .A0(n5818), .A1(GFidata[271]), .Z(n5176));
Q_MX02 U3684 ( .S(n5817), .A0(n5174), .A1(n4166), .Z(n5175));
Q_AN02 U3685 ( .A0(n5818), .A1(GFidata[270]), .Z(n5174));
Q_MX02 U3686 ( .S(n5817), .A0(n5172), .A1(n4165), .Z(n5173));
Q_AN02 U3687 ( .A0(n5818), .A1(GFidata[269]), .Z(n5172));
Q_MX02 U3688 ( .S(n5817), .A0(n5170), .A1(n4164), .Z(n5171));
Q_AN02 U3689 ( .A0(n5818), .A1(GFidata[268]), .Z(n5170));
Q_MX02 U3690 ( .S(n5817), .A0(n5168), .A1(n4163), .Z(n5169));
Q_AN02 U3691 ( .A0(n5818), .A1(GFidata[267]), .Z(n5168));
Q_MX02 U3692 ( .S(n5817), .A0(n5166), .A1(n4162), .Z(n5167));
Q_AN02 U3693 ( .A0(n5818), .A1(GFidata[266]), .Z(n5166));
Q_MX02 U3694 ( .S(n5817), .A0(n5164), .A1(n4161), .Z(n5165));
Q_AN02 U3695 ( .A0(n5818), .A1(GFidata[265]), .Z(n5164));
Q_MX02 U3696 ( .S(n5817), .A0(n5162), .A1(n4160), .Z(n5163));
Q_AN02 U3697 ( .A0(n5818), .A1(GFidata[264]), .Z(n5162));
Q_MX02 U3698 ( .S(n5817), .A0(n5160), .A1(n4159), .Z(n5161));
Q_AN02 U3699 ( .A0(n5818), .A1(GFidata[263]), .Z(n5160));
Q_MX02 U3700 ( .S(n5817), .A0(n5158), .A1(n4158), .Z(n5159));
Q_AN02 U3701 ( .A0(n5818), .A1(GFidata[262]), .Z(n5158));
Q_MX02 U3702 ( .S(n5817), .A0(n5156), .A1(n4157), .Z(n5157));
Q_AN02 U3703 ( .A0(n5818), .A1(GFidata[261]), .Z(n5156));
Q_MX02 U3704 ( .S(n5817), .A0(n5154), .A1(n4156), .Z(n5155));
Q_AN02 U3705 ( .A0(n5818), .A1(GFidata[260]), .Z(n5154));
Q_MX02 U3706 ( .S(n5817), .A0(n5152), .A1(n4155), .Z(n5153));
Q_AN02 U3707 ( .A0(n5818), .A1(GFidata[259]), .Z(n5152));
Q_MX02 U3708 ( .S(n5817), .A0(n5150), .A1(n4154), .Z(n5151));
Q_AN02 U3709 ( .A0(n5818), .A1(GFidata[258]), .Z(n5150));
Q_MX02 U3710 ( .S(n5817), .A0(n5148), .A1(n4153), .Z(n5149));
Q_AN02 U3711 ( .A0(n5818), .A1(GFidata[257]), .Z(n5148));
Q_MX02 U3712 ( .S(n5817), .A0(n5146), .A1(n4152), .Z(n5147));
Q_AN02 U3713 ( .A0(n5818), .A1(GFidata[256]), .Z(n5146));
Q_MX02 U3714 ( .S(n5817), .A0(n5144), .A1(n4151), .Z(n5145));
Q_AN02 U3715 ( .A0(n5818), .A1(GFidata[255]), .Z(n5144));
Q_MX02 U3716 ( .S(n5817), .A0(n5142), .A1(n4150), .Z(n5143));
Q_AN02 U3717 ( .A0(n5818), .A1(GFidata[254]), .Z(n5142));
Q_MX02 U3718 ( .S(n5817), .A0(n5140), .A1(n4149), .Z(n5141));
Q_AN02 U3719 ( .A0(n5818), .A1(GFidata[253]), .Z(n5140));
Q_MX02 U3720 ( .S(n5817), .A0(n5138), .A1(n4148), .Z(n5139));
Q_AN02 U3721 ( .A0(n5818), .A1(GFidata[252]), .Z(n5138));
Q_MX02 U3722 ( .S(n5817), .A0(n5136), .A1(n4147), .Z(n5137));
Q_AN02 U3723 ( .A0(n5818), .A1(GFidata[251]), .Z(n5136));
Q_MX02 U3724 ( .S(n5817), .A0(n5134), .A1(n4146), .Z(n5135));
Q_AN02 U3725 ( .A0(n5818), .A1(GFidata[250]), .Z(n5134));
Q_MX02 U3726 ( .S(n5817), .A0(n5132), .A1(n4145), .Z(n5133));
Q_AN02 U3727 ( .A0(n5818), .A1(GFidata[249]), .Z(n5132));
Q_MX02 U3728 ( .S(n5817), .A0(n5130), .A1(n4144), .Z(n5131));
Q_AN02 U3729 ( .A0(n5818), .A1(GFidata[248]), .Z(n5130));
Q_MX02 U3730 ( .S(n5817), .A0(n5128), .A1(n4143), .Z(n5129));
Q_AN02 U3731 ( .A0(n5818), .A1(GFidata[247]), .Z(n5128));
Q_MX02 U3732 ( .S(n5817), .A0(n5126), .A1(n4142), .Z(n5127));
Q_AN02 U3733 ( .A0(n5818), .A1(GFidata[246]), .Z(n5126));
Q_MX02 U3734 ( .S(n5817), .A0(n5124), .A1(n4141), .Z(n5125));
Q_AN02 U3735 ( .A0(n5818), .A1(GFidata[245]), .Z(n5124));
Q_MX02 U3736 ( .S(n5817), .A0(n5122), .A1(n4140), .Z(n5123));
Q_AN02 U3737 ( .A0(n5818), .A1(GFidata[244]), .Z(n5122));
Q_MX02 U3738 ( .S(n5817), .A0(n5120), .A1(n4139), .Z(n5121));
Q_AN02 U3739 ( .A0(n5818), .A1(GFidata[243]), .Z(n5120));
Q_MX02 U3740 ( .S(n5817), .A0(n5118), .A1(n4138), .Z(n5119));
Q_AN02 U3741 ( .A0(n5818), .A1(GFidata[242]), .Z(n5118));
Q_MX02 U3742 ( .S(n5817), .A0(n5116), .A1(n4137), .Z(n5117));
Q_AN02 U3743 ( .A0(n5818), .A1(GFidata[241]), .Z(n5116));
Q_MX02 U3744 ( .S(n5817), .A0(n5114), .A1(n4136), .Z(n5115));
Q_AN02 U3745 ( .A0(n5818), .A1(GFidata[240]), .Z(n5114));
Q_MX02 U3746 ( .S(n5817), .A0(n5112), .A1(n4135), .Z(n5113));
Q_AN02 U3747 ( .A0(n5818), .A1(GFidata[239]), .Z(n5112));
Q_MX02 U3748 ( .S(n5817), .A0(n5110), .A1(n4134), .Z(n5111));
Q_AN02 U3749 ( .A0(n5818), .A1(GFidata[238]), .Z(n5110));
Q_MX02 U3750 ( .S(n5817), .A0(n5108), .A1(n4133), .Z(n5109));
Q_AN02 U3751 ( .A0(n5818), .A1(GFidata[237]), .Z(n5108));
Q_MX02 U3752 ( .S(n5817), .A0(n5106), .A1(n4132), .Z(n5107));
Q_AN02 U3753 ( .A0(n5818), .A1(GFidata[236]), .Z(n5106));
Q_MX02 U3754 ( .S(n5817), .A0(n5104), .A1(n4131), .Z(n5105));
Q_AN02 U3755 ( .A0(n5818), .A1(GFidata[235]), .Z(n5104));
Q_MX02 U3756 ( .S(n5817), .A0(n5102), .A1(n4130), .Z(n5103));
Q_AN02 U3757 ( .A0(n5818), .A1(GFidata[234]), .Z(n5102));
Q_MX02 U3758 ( .S(n5817), .A0(n5100), .A1(n4129), .Z(n5101));
Q_AN02 U3759 ( .A0(n5818), .A1(GFidata[233]), .Z(n5100));
Q_MX02 U3760 ( .S(n5817), .A0(n5098), .A1(n4128), .Z(n5099));
Q_AN02 U3761 ( .A0(n5818), .A1(GFidata[232]), .Z(n5098));
Q_MX02 U3762 ( .S(n5817), .A0(n5096), .A1(n4127), .Z(n5097));
Q_AN02 U3763 ( .A0(n5818), .A1(GFidata[231]), .Z(n5096));
Q_MX02 U3764 ( .S(n5817), .A0(n5094), .A1(n4126), .Z(n5095));
Q_AN02 U3765 ( .A0(n5818), .A1(GFidata[230]), .Z(n5094));
Q_MX02 U3766 ( .S(n5817), .A0(n5092), .A1(n4125), .Z(n5093));
Q_AN02 U3767 ( .A0(n5818), .A1(GFidata[229]), .Z(n5092));
Q_MX02 U3768 ( .S(n5817), .A0(n5090), .A1(n4124), .Z(n5091));
Q_AN02 U3769 ( .A0(n5818), .A1(GFidata[228]), .Z(n5090));
Q_MX02 U3770 ( .S(n5817), .A0(n5088), .A1(n4123), .Z(n5089));
Q_AN02 U3771 ( .A0(n5818), .A1(GFidata[227]), .Z(n5088));
Q_MX02 U3772 ( .S(n5817), .A0(n5086), .A1(n4122), .Z(n5087));
Q_AN02 U3773 ( .A0(n5818), .A1(GFidata[226]), .Z(n5086));
Q_MX02 U3774 ( .S(n5817), .A0(n5084), .A1(n4121), .Z(n5085));
Q_AN02 U3775 ( .A0(n5818), .A1(GFidata[225]), .Z(n5084));
Q_MX02 U3776 ( .S(n5817), .A0(n5082), .A1(n4120), .Z(n5083));
Q_AN02 U3777 ( .A0(n5818), .A1(GFidata[224]), .Z(n5082));
Q_MX02 U3778 ( .S(n5817), .A0(n5080), .A1(n4119), .Z(n5081));
Q_AN02 U3779 ( .A0(n5818), .A1(GFidata[223]), .Z(n5080));
Q_MX02 U3780 ( .S(n5817), .A0(n5078), .A1(n4118), .Z(n5079));
Q_AN02 U3781 ( .A0(n5818), .A1(GFidata[222]), .Z(n5078));
Q_MX02 U3782 ( .S(n5817), .A0(n5076), .A1(n4117), .Z(n5077));
Q_AN02 U3783 ( .A0(n5818), .A1(GFidata[221]), .Z(n5076));
Q_MX02 U3784 ( .S(n5817), .A0(n5074), .A1(n4116), .Z(n5075));
Q_AN02 U3785 ( .A0(n5818), .A1(GFidata[220]), .Z(n5074));
Q_MX02 U3786 ( .S(n5817), .A0(n5072), .A1(n4115), .Z(n5073));
Q_AN02 U3787 ( .A0(n5818), .A1(GFidata[219]), .Z(n5072));
Q_MX02 U3788 ( .S(n5817), .A0(n5070), .A1(n4114), .Z(n5071));
Q_AN02 U3789 ( .A0(n5818), .A1(GFidata[218]), .Z(n5070));
Q_MX02 U3790 ( .S(n5817), .A0(n5068), .A1(n4113), .Z(n5069));
Q_AN02 U3791 ( .A0(n5818), .A1(GFidata[217]), .Z(n5068));
Q_MX02 U3792 ( .S(n5817), .A0(n5066), .A1(n4112), .Z(n5067));
Q_AN02 U3793 ( .A0(n5818), .A1(GFidata[216]), .Z(n5066));
Q_MX02 U3794 ( .S(n5817), .A0(n5064), .A1(n4111), .Z(n5065));
Q_AN02 U3795 ( .A0(n5818), .A1(GFidata[215]), .Z(n5064));
Q_MX02 U3796 ( .S(n5817), .A0(n5062), .A1(n4110), .Z(n5063));
Q_AN02 U3797 ( .A0(n5818), .A1(GFidata[214]), .Z(n5062));
Q_MX02 U3798 ( .S(n5817), .A0(n5060), .A1(n4109), .Z(n5061));
Q_AN02 U3799 ( .A0(n5818), .A1(GFidata[213]), .Z(n5060));
Q_MX02 U3800 ( .S(n5817), .A0(n5058), .A1(n4108), .Z(n5059));
Q_AN02 U3801 ( .A0(n5818), .A1(GFidata[212]), .Z(n5058));
Q_MX02 U3802 ( .S(n5817), .A0(n5056), .A1(n4107), .Z(n5057));
Q_AN02 U3803 ( .A0(n5818), .A1(GFidata[211]), .Z(n5056));
Q_MX02 U3804 ( .S(n5817), .A0(n5054), .A1(n4106), .Z(n5055));
Q_AN02 U3805 ( .A0(n5818), .A1(GFidata[210]), .Z(n5054));
Q_MX02 U3806 ( .S(n5817), .A0(n5052), .A1(n4105), .Z(n5053));
Q_AN02 U3807 ( .A0(n5818), .A1(GFidata[209]), .Z(n5052));
Q_MX02 U3808 ( .S(n5817), .A0(n5050), .A1(n4104), .Z(n5051));
Q_AN02 U3809 ( .A0(n5818), .A1(GFidata[208]), .Z(n5050));
Q_MX02 U3810 ( .S(n5817), .A0(n5048), .A1(n4103), .Z(n5049));
Q_AN02 U3811 ( .A0(n5818), .A1(GFidata[207]), .Z(n5048));
Q_MX02 U3812 ( .S(n5817), .A0(n5046), .A1(n4102), .Z(n5047));
Q_AN02 U3813 ( .A0(n5818), .A1(GFidata[206]), .Z(n5046));
Q_MX02 U3814 ( .S(n5817), .A0(n5044), .A1(n4101), .Z(n5045));
Q_AN02 U3815 ( .A0(n5818), .A1(GFidata[205]), .Z(n5044));
Q_MX02 U3816 ( .S(n5817), .A0(n5042), .A1(n4100), .Z(n5043));
Q_AN02 U3817 ( .A0(n5818), .A1(GFidata[204]), .Z(n5042));
Q_MX02 U3818 ( .S(n5817), .A0(n5040), .A1(n4099), .Z(n5041));
Q_AN02 U3819 ( .A0(n5818), .A1(GFidata[203]), .Z(n5040));
Q_MX02 U3820 ( .S(n5817), .A0(n5038), .A1(n4098), .Z(n5039));
Q_AN02 U3821 ( .A0(n5818), .A1(GFidata[202]), .Z(n5038));
Q_MX02 U3822 ( .S(n5817), .A0(n5036), .A1(n4097), .Z(n5037));
Q_AN02 U3823 ( .A0(n5818), .A1(GFidata[201]), .Z(n5036));
Q_MX02 U3824 ( .S(n5817), .A0(n5034), .A1(n4096), .Z(n5035));
Q_AN02 U3825 ( .A0(n5818), .A1(GFidata[200]), .Z(n5034));
Q_MX02 U3826 ( .S(n5817), .A0(n5032), .A1(n4095), .Z(n5033));
Q_AN02 U3827 ( .A0(n5818), .A1(GFidata[199]), .Z(n5032));
Q_MX02 U3828 ( .S(n5817), .A0(n5030), .A1(n4094), .Z(n5031));
Q_AN02 U3829 ( .A0(n5818), .A1(GFidata[198]), .Z(n5030));
Q_MX02 U3830 ( .S(n5817), .A0(n5028), .A1(n4093), .Z(n5029));
Q_AN02 U3831 ( .A0(n5818), .A1(GFidata[197]), .Z(n5028));
Q_MX02 U3832 ( .S(n5817), .A0(n5026), .A1(n4092), .Z(n5027));
Q_AN02 U3833 ( .A0(n5818), .A1(GFidata[196]), .Z(n5026));
Q_MX02 U3834 ( .S(n5817), .A0(n5024), .A1(n4091), .Z(n5025));
Q_AN02 U3835 ( .A0(n5818), .A1(GFidata[195]), .Z(n5024));
Q_MX02 U3836 ( .S(n5817), .A0(n5022), .A1(n4090), .Z(n5023));
Q_AN02 U3837 ( .A0(n5818), .A1(GFidata[194]), .Z(n5022));
Q_MX02 U3838 ( .S(n5817), .A0(n5020), .A1(n4089), .Z(n5021));
Q_AN02 U3839 ( .A0(n5818), .A1(GFidata[193]), .Z(n5020));
Q_MX02 U3840 ( .S(n5817), .A0(n5018), .A1(n4088), .Z(n5019));
Q_AN02 U3841 ( .A0(n5818), .A1(GFidata[192]), .Z(n5018));
Q_MX02 U3842 ( .S(n5817), .A0(n5016), .A1(n4087), .Z(n5017));
Q_AN02 U3843 ( .A0(n5818), .A1(GFidata[191]), .Z(n5016));
Q_MX02 U3844 ( .S(n5817), .A0(n5014), .A1(n4086), .Z(n5015));
Q_AN02 U3845 ( .A0(n5818), .A1(GFidata[190]), .Z(n5014));
Q_MX02 U3846 ( .S(n5817), .A0(n5012), .A1(n4085), .Z(n5013));
Q_AN02 U3847 ( .A0(n5818), .A1(GFidata[189]), .Z(n5012));
Q_MX02 U3848 ( .S(n5817), .A0(n5010), .A1(n4084), .Z(n5011));
Q_AN02 U3849 ( .A0(n5818), .A1(GFidata[188]), .Z(n5010));
Q_MX02 U3850 ( .S(n5817), .A0(n5008), .A1(n4083), .Z(n5009));
Q_AN02 U3851 ( .A0(n5818), .A1(GFidata[187]), .Z(n5008));
Q_MX02 U3852 ( .S(n5817), .A0(n5006), .A1(n4082), .Z(n5007));
Q_AN02 U3853 ( .A0(n5818), .A1(GFidata[186]), .Z(n5006));
Q_MX02 U3854 ( .S(n5817), .A0(n5004), .A1(n4081), .Z(n5005));
Q_AN02 U3855 ( .A0(n5818), .A1(GFidata[185]), .Z(n5004));
Q_MX02 U3856 ( .S(n5817), .A0(n5002), .A1(n4080), .Z(n5003));
Q_AN02 U3857 ( .A0(n5818), .A1(GFidata[184]), .Z(n5002));
Q_MX02 U3858 ( .S(n5817), .A0(n5000), .A1(n4079), .Z(n5001));
Q_AN02 U3859 ( .A0(n5818), .A1(GFidata[183]), .Z(n5000));
Q_MX02 U3860 ( .S(n5817), .A0(n4998), .A1(n4078), .Z(n4999));
Q_AN02 U3861 ( .A0(n5818), .A1(GFidata[182]), .Z(n4998));
Q_MX02 U3862 ( .S(n5817), .A0(n4996), .A1(n4077), .Z(n4997));
Q_AN02 U3863 ( .A0(n5818), .A1(GFidata[181]), .Z(n4996));
Q_MX02 U3864 ( .S(n5817), .A0(n4994), .A1(n4076), .Z(n4995));
Q_AN02 U3865 ( .A0(n5818), .A1(GFidata[180]), .Z(n4994));
Q_MX02 U3866 ( .S(n5817), .A0(n4992), .A1(n4075), .Z(n4993));
Q_AN02 U3867 ( .A0(n5818), .A1(GFidata[179]), .Z(n4992));
Q_MX02 U3868 ( .S(n5817), .A0(n4990), .A1(n4074), .Z(n4991));
Q_AN02 U3869 ( .A0(n5818), .A1(GFidata[178]), .Z(n4990));
Q_MX02 U3870 ( .S(n5817), .A0(n4988), .A1(n4073), .Z(n4989));
Q_AN02 U3871 ( .A0(n5818), .A1(GFidata[177]), .Z(n4988));
Q_MX02 U3872 ( .S(n5817), .A0(n4986), .A1(n4072), .Z(n4987));
Q_AN02 U3873 ( .A0(n5818), .A1(GFidata[176]), .Z(n4986));
Q_MX02 U3874 ( .S(n5817), .A0(n4984), .A1(n4071), .Z(n4985));
Q_AN02 U3875 ( .A0(n5818), .A1(GFidata[175]), .Z(n4984));
Q_MX02 U3876 ( .S(n5817), .A0(n4982), .A1(n4070), .Z(n4983));
Q_AN02 U3877 ( .A0(n5818), .A1(GFidata[174]), .Z(n4982));
Q_MX02 U3878 ( .S(n5817), .A0(n4980), .A1(n4069), .Z(n4981));
Q_AN02 U3879 ( .A0(n5818), .A1(GFidata[173]), .Z(n4980));
Q_MX02 U3880 ( .S(n5817), .A0(n4978), .A1(n4068), .Z(n4979));
Q_AN02 U3881 ( .A0(n5818), .A1(GFidata[172]), .Z(n4978));
Q_MX02 U3882 ( .S(n5817), .A0(n4976), .A1(n4067), .Z(n4977));
Q_AN02 U3883 ( .A0(n5818), .A1(GFidata[171]), .Z(n4976));
Q_MX02 U3884 ( .S(n5817), .A0(n4974), .A1(n4066), .Z(n4975));
Q_AN02 U3885 ( .A0(n5818), .A1(GFidata[170]), .Z(n4974));
Q_MX02 U3886 ( .S(n5817), .A0(n4972), .A1(n4065), .Z(n4973));
Q_AN02 U3887 ( .A0(n5818), .A1(GFidata[169]), .Z(n4972));
Q_MX02 U3888 ( .S(n5817), .A0(n4970), .A1(n4064), .Z(n4971));
Q_AN02 U3889 ( .A0(n5818), .A1(GFidata[168]), .Z(n4970));
Q_MX02 U3890 ( .S(n5817), .A0(n4968), .A1(n4063), .Z(n4969));
Q_AN02 U3891 ( .A0(n5818), .A1(GFidata[167]), .Z(n4968));
Q_MX02 U3892 ( .S(n5817), .A0(n4966), .A1(n4062), .Z(n4967));
Q_AN02 U3893 ( .A0(n5818), .A1(GFidata[166]), .Z(n4966));
Q_MX02 U3894 ( .S(n5817), .A0(n4964), .A1(n4061), .Z(n4965));
Q_AN02 U3895 ( .A0(n5818), .A1(GFidata[165]), .Z(n4964));
Q_MX02 U3896 ( .S(n5817), .A0(n4962), .A1(n4060), .Z(n4963));
Q_AN02 U3897 ( .A0(n5818), .A1(GFidata[164]), .Z(n4962));
Q_MX02 U3898 ( .S(n5817), .A0(n4960), .A1(n4059), .Z(n4961));
Q_AN02 U3899 ( .A0(n5818), .A1(GFidata[163]), .Z(n4960));
Q_MX02 U3900 ( .S(n5817), .A0(n4958), .A1(n4058), .Z(n4959));
Q_AN02 U3901 ( .A0(n5818), .A1(GFidata[162]), .Z(n4958));
Q_MX02 U3902 ( .S(n5817), .A0(n4956), .A1(n4057), .Z(n4957));
Q_AN02 U3903 ( .A0(n5818), .A1(GFidata[161]), .Z(n4956));
Q_MX02 U3904 ( .S(n5817), .A0(n4954), .A1(n4056), .Z(n4955));
Q_AN02 U3905 ( .A0(n5818), .A1(GFidata[160]), .Z(n4954));
Q_MX02 U3906 ( .S(n5817), .A0(n4952), .A1(n4055), .Z(n4953));
Q_AN02 U3907 ( .A0(n5818), .A1(GFidata[159]), .Z(n4952));
Q_MX02 U3908 ( .S(n5817), .A0(n4950), .A1(n4054), .Z(n4951));
Q_AN02 U3909 ( .A0(n5818), .A1(GFidata[158]), .Z(n4950));
Q_MX02 U3910 ( .S(n5817), .A0(n4948), .A1(n4053), .Z(n4949));
Q_AN02 U3911 ( .A0(n5818), .A1(GFidata[157]), .Z(n4948));
Q_MX02 U3912 ( .S(n5817), .A0(n4946), .A1(n4052), .Z(n4947));
Q_AN02 U3913 ( .A0(n5818), .A1(GFidata[156]), .Z(n4946));
Q_MX02 U3914 ( .S(n5817), .A0(n4944), .A1(n4051), .Z(n4945));
Q_AN02 U3915 ( .A0(n5818), .A1(GFidata[155]), .Z(n4944));
Q_MX02 U3916 ( .S(n5817), .A0(n4942), .A1(n4050), .Z(n4943));
Q_AN02 U3917 ( .A0(n5818), .A1(GFidata[154]), .Z(n4942));
Q_MX02 U3918 ( .S(n5817), .A0(n4940), .A1(n4049), .Z(n4941));
Q_AN02 U3919 ( .A0(n5818), .A1(GFidata[153]), .Z(n4940));
Q_MX02 U3920 ( .S(n5817), .A0(n4938), .A1(n4048), .Z(n4939));
Q_AN02 U3921 ( .A0(n5818), .A1(GFidata[152]), .Z(n4938));
Q_MX02 U3922 ( .S(n5817), .A0(n4936), .A1(n4047), .Z(n4937));
Q_AN02 U3923 ( .A0(n5818), .A1(GFidata[151]), .Z(n4936));
Q_MX02 U3924 ( .S(n5817), .A0(n4934), .A1(n4046), .Z(n4935));
Q_AN02 U3925 ( .A0(n5818), .A1(GFidata[150]), .Z(n4934));
Q_MX02 U3926 ( .S(n5817), .A0(n4932), .A1(n4045), .Z(n4933));
Q_AN02 U3927 ( .A0(n5818), .A1(GFidata[149]), .Z(n4932));
Q_MX02 U3928 ( .S(n5817), .A0(n4930), .A1(n4044), .Z(n4931));
Q_AN02 U3929 ( .A0(n5818), .A1(GFidata[148]), .Z(n4930));
Q_MX02 U3930 ( .S(n5817), .A0(n4928), .A1(n4043), .Z(n4929));
Q_AN02 U3931 ( .A0(n5818), .A1(GFidata[147]), .Z(n4928));
Q_MX02 U3932 ( .S(n5817), .A0(n4926), .A1(n4042), .Z(n4927));
Q_AN02 U3933 ( .A0(n5818), .A1(GFidata[146]), .Z(n4926));
Q_MX02 U3934 ( .S(n5817), .A0(n4924), .A1(n4041), .Z(n4925));
Q_AN02 U3935 ( .A0(n5818), .A1(GFidata[145]), .Z(n4924));
Q_MX02 U3936 ( .S(n5817), .A0(n4922), .A1(n4040), .Z(n4923));
Q_AN02 U3937 ( .A0(n5818), .A1(GFidata[144]), .Z(n4922));
Q_MX02 U3938 ( .S(n5817), .A0(n4920), .A1(n4039), .Z(n4921));
Q_AN02 U3939 ( .A0(n5818), .A1(GFidata[143]), .Z(n4920));
Q_MX02 U3940 ( .S(n5817), .A0(n4918), .A1(n4038), .Z(n4919));
Q_AN02 U3941 ( .A0(n5818), .A1(GFidata[142]), .Z(n4918));
Q_MX02 U3942 ( .S(n5817), .A0(n4916), .A1(n4037), .Z(n4917));
Q_AN02 U3943 ( .A0(n5818), .A1(GFidata[141]), .Z(n4916));
Q_MX02 U3944 ( .S(n5817), .A0(n4914), .A1(n4036), .Z(n4915));
Q_AN02 U3945 ( .A0(n5818), .A1(GFidata[140]), .Z(n4914));
Q_MX02 U3946 ( .S(n5817), .A0(n4912), .A1(n4035), .Z(n4913));
Q_AN02 U3947 ( .A0(n5818), .A1(GFidata[139]), .Z(n4912));
Q_MX02 U3948 ( .S(n5817), .A0(n4910), .A1(n4034), .Z(n4911));
Q_AN02 U3949 ( .A0(n5818), .A1(GFidata[138]), .Z(n4910));
Q_MX02 U3950 ( .S(n5817), .A0(n4908), .A1(n4033), .Z(n4909));
Q_AN02 U3951 ( .A0(n5818), .A1(GFidata[137]), .Z(n4908));
Q_MX02 U3952 ( .S(n5817), .A0(n4906), .A1(n4032), .Z(n4907));
Q_AN02 U3953 ( .A0(n5818), .A1(GFidata[136]), .Z(n4906));
Q_MX02 U3954 ( .S(n5817), .A0(n4904), .A1(n4031), .Z(n4905));
Q_AN02 U3955 ( .A0(n5818), .A1(GFidata[135]), .Z(n4904));
Q_MX02 U3956 ( .S(n5817), .A0(n4902), .A1(n4030), .Z(n4903));
Q_AN02 U3957 ( .A0(n5818), .A1(GFidata[134]), .Z(n4902));
Q_MX02 U3958 ( .S(n5817), .A0(n4900), .A1(n4029), .Z(n4901));
Q_AN02 U3959 ( .A0(n5818), .A1(GFidata[133]), .Z(n4900));
Q_MX02 U3960 ( .S(n5817), .A0(n4898), .A1(n4028), .Z(n4899));
Q_AN02 U3961 ( .A0(n5818), .A1(GFidata[132]), .Z(n4898));
Q_MX02 U3962 ( .S(n5817), .A0(n4896), .A1(n4027), .Z(n4897));
Q_AN02 U3963 ( .A0(n5818), .A1(GFidata[131]), .Z(n4896));
Q_MX02 U3964 ( .S(n5817), .A0(n4894), .A1(n4026), .Z(n4895));
Q_AN02 U3965 ( .A0(n5818), .A1(GFidata[130]), .Z(n4894));
Q_MX02 U3966 ( .S(n5817), .A0(n4892), .A1(n4025), .Z(n4893));
Q_AN02 U3967 ( .A0(n5818), .A1(GFidata[129]), .Z(n4892));
Q_MX02 U3968 ( .S(n5817), .A0(n4890), .A1(n4024), .Z(n4891));
Q_AN02 U3969 ( .A0(n5818), .A1(GFidata[128]), .Z(n4890));
Q_MX02 U3970 ( .S(n5817), .A0(n4888), .A1(n4023), .Z(n4889));
Q_AN02 U3971 ( .A0(n5818), .A1(GFidata[127]), .Z(n4888));
Q_MX02 U3972 ( .S(n5817), .A0(n4886), .A1(n4022), .Z(n4887));
Q_AN02 U3973 ( .A0(n5818), .A1(GFidata[126]), .Z(n4886));
Q_MX02 U3974 ( .S(n5817), .A0(n4884), .A1(n4021), .Z(n4885));
Q_AN02 U3975 ( .A0(n5818), .A1(GFidata[125]), .Z(n4884));
Q_MX02 U3976 ( .S(n5817), .A0(n4882), .A1(n4020), .Z(n4883));
Q_AN02 U3977 ( .A0(n5818), .A1(GFidata[124]), .Z(n4882));
Q_MX02 U3978 ( .S(n5817), .A0(n4880), .A1(n4019), .Z(n4881));
Q_AN02 U3979 ( .A0(n5818), .A1(GFidata[123]), .Z(n4880));
Q_MX02 U3980 ( .S(n5817), .A0(n4878), .A1(n4018), .Z(n4879));
Q_AN02 U3981 ( .A0(n5818), .A1(GFidata[122]), .Z(n4878));
Q_MX02 U3982 ( .S(n5817), .A0(n4876), .A1(n4017), .Z(n4877));
Q_AN02 U3983 ( .A0(n5818), .A1(GFidata[121]), .Z(n4876));
Q_MX02 U3984 ( .S(n5817), .A0(n4874), .A1(n4016), .Z(n4875));
Q_AN02 U3985 ( .A0(n5818), .A1(GFidata[120]), .Z(n4874));
Q_MX02 U3986 ( .S(n5817), .A0(n4872), .A1(n4015), .Z(n4873));
Q_AN02 U3987 ( .A0(n5818), .A1(GFidata[119]), .Z(n4872));
Q_MX02 U3988 ( .S(n5817), .A0(n4870), .A1(n4014), .Z(n4871));
Q_AN02 U3989 ( .A0(n5818), .A1(GFidata[118]), .Z(n4870));
Q_MX02 U3990 ( .S(n5817), .A0(n4868), .A1(n4013), .Z(n4869));
Q_AN02 U3991 ( .A0(n5818), .A1(GFidata[117]), .Z(n4868));
Q_MX02 U3992 ( .S(n5817), .A0(n4866), .A1(n4012), .Z(n4867));
Q_AN02 U3993 ( .A0(n5818), .A1(GFidata[116]), .Z(n4866));
Q_MX02 U3994 ( .S(n5817), .A0(n4864), .A1(n4011), .Z(n4865));
Q_AN02 U3995 ( .A0(n5818), .A1(GFidata[115]), .Z(n4864));
Q_MX02 U3996 ( .S(n5817), .A0(n4862), .A1(n4010), .Z(n4863));
Q_AN02 U3997 ( .A0(n5818), .A1(GFidata[114]), .Z(n4862));
Q_MX02 U3998 ( .S(n5817), .A0(n4860), .A1(n4009), .Z(n4861));
Q_AN02 U3999 ( .A0(n5818), .A1(GFidata[113]), .Z(n4860));
Q_MX02 U4000 ( .S(n5817), .A0(n4858), .A1(n4008), .Z(n4859));
Q_AN02 U4001 ( .A0(n5818), .A1(GFidata[112]), .Z(n4858));
Q_MX02 U4002 ( .S(n5817), .A0(n4856), .A1(n4007), .Z(n4857));
Q_AN02 U4003 ( .A0(n5818), .A1(GFidata[111]), .Z(n4856));
Q_MX02 U4004 ( .S(n5817), .A0(n4854), .A1(n4006), .Z(n4855));
Q_AN02 U4005 ( .A0(n5818), .A1(GFidata[110]), .Z(n4854));
Q_MX02 U4006 ( .S(n5817), .A0(n4852), .A1(n4005), .Z(n4853));
Q_AN02 U4007 ( .A0(n5818), .A1(GFidata[109]), .Z(n4852));
Q_MX02 U4008 ( .S(n5817), .A0(n4850), .A1(n4004), .Z(n4851));
Q_AN02 U4009 ( .A0(n5818), .A1(GFidata[108]), .Z(n4850));
Q_MX02 U4010 ( .S(n5817), .A0(n4848), .A1(n4003), .Z(n4849));
Q_AN02 U4011 ( .A0(n5818), .A1(GFidata[107]), .Z(n4848));
Q_MX02 U4012 ( .S(n5817), .A0(n4846), .A1(n4002), .Z(n4847));
Q_AN02 U4013 ( .A0(n5818), .A1(GFidata[106]), .Z(n4846));
Q_MX02 U4014 ( .S(n5817), .A0(n4844), .A1(n4001), .Z(n4845));
Q_AN02 U4015 ( .A0(n5818), .A1(GFidata[105]), .Z(n4844));
Q_MX02 U4016 ( .S(n5817), .A0(n4842), .A1(n4000), .Z(n4843));
Q_AN02 U4017 ( .A0(n5818), .A1(GFidata[104]), .Z(n4842));
Q_MX02 U4018 ( .S(n5817), .A0(n4840), .A1(n3999), .Z(n4841));
Q_AN02 U4019 ( .A0(n5818), .A1(GFidata[103]), .Z(n4840));
Q_MX02 U4020 ( .S(n5817), .A0(n4838), .A1(n3998), .Z(n4839));
Q_AN02 U4021 ( .A0(n5818), .A1(GFidata[102]), .Z(n4838));
Q_MX02 U4022 ( .S(n5817), .A0(n4836), .A1(n3997), .Z(n4837));
Q_AN02 U4023 ( .A0(n5818), .A1(GFidata[101]), .Z(n4836));
Q_MX02 U4024 ( .S(n5817), .A0(n4834), .A1(n3996), .Z(n4835));
Q_AN02 U4025 ( .A0(n5818), .A1(GFidata[100]), .Z(n4834));
Q_MX02 U4026 ( .S(n5817), .A0(n4832), .A1(n3995), .Z(n4833));
Q_AN02 U4027 ( .A0(n5818), .A1(GFidata[99]), .Z(n4832));
Q_MX02 U4028 ( .S(n5817), .A0(n4830), .A1(n3994), .Z(n4831));
Q_AN02 U4029 ( .A0(n5818), .A1(GFidata[98]), .Z(n4830));
Q_MX02 U4030 ( .S(n5817), .A0(n4828), .A1(n3993), .Z(n4829));
Q_AN02 U4031 ( .A0(n5818), .A1(GFidata[97]), .Z(n4828));
Q_MX02 U4032 ( .S(n5817), .A0(n4826), .A1(n3992), .Z(n4827));
Q_AN02 U4033 ( .A0(n5818), .A1(GFidata[96]), .Z(n4826));
Q_MX02 U4034 ( .S(n5817), .A0(n4824), .A1(n3991), .Z(n4825));
Q_AN02 U4035 ( .A0(n5818), .A1(GFidata[95]), .Z(n4824));
Q_MX02 U4036 ( .S(n5817), .A0(n4822), .A1(n3990), .Z(n4823));
Q_AN02 U4037 ( .A0(n5818), .A1(GFidata[94]), .Z(n4822));
Q_MX02 U4038 ( .S(n5817), .A0(n4820), .A1(n3989), .Z(n4821));
Q_AN02 U4039 ( .A0(n5818), .A1(GFidata[93]), .Z(n4820));
Q_MX02 U4040 ( .S(n5817), .A0(n4818), .A1(n3988), .Z(n4819));
Q_AN02 U4041 ( .A0(n5818), .A1(GFidata[92]), .Z(n4818));
Q_MX02 U4042 ( .S(n5817), .A0(n4816), .A1(n3987), .Z(n4817));
Q_AN02 U4043 ( .A0(n5818), .A1(GFidata[91]), .Z(n4816));
Q_MX02 U4044 ( .S(n5817), .A0(n4814), .A1(n3986), .Z(n4815));
Q_AN02 U4045 ( .A0(n5818), .A1(GFidata[90]), .Z(n4814));
Q_MX02 U4046 ( .S(n5817), .A0(n4812), .A1(n3985), .Z(n4813));
Q_AN02 U4047 ( .A0(n5818), .A1(GFidata[89]), .Z(n4812));
Q_MX02 U4048 ( .S(n5817), .A0(n4810), .A1(n3984), .Z(n4811));
Q_AN02 U4049 ( .A0(n5818), .A1(GFidata[88]), .Z(n4810));
Q_MX02 U4050 ( .S(n5817), .A0(n4808), .A1(n3983), .Z(n4809));
Q_AN02 U4051 ( .A0(n5818), .A1(GFidata[87]), .Z(n4808));
Q_MX02 U4052 ( .S(n5817), .A0(n4806), .A1(n3982), .Z(n4807));
Q_AN02 U4053 ( .A0(n5818), .A1(GFidata[86]), .Z(n4806));
Q_MX02 U4054 ( .S(n5817), .A0(n4804), .A1(n3981), .Z(n4805));
Q_AN02 U4055 ( .A0(n5818), .A1(GFidata[85]), .Z(n4804));
Q_MX02 U4056 ( .S(n5817), .A0(n4802), .A1(n3980), .Z(n4803));
Q_AN02 U4057 ( .A0(n5818), .A1(GFidata[84]), .Z(n4802));
Q_MX02 U4058 ( .S(n5817), .A0(n4800), .A1(n3979), .Z(n4801));
Q_AN02 U4059 ( .A0(n5818), .A1(GFidata[83]), .Z(n4800));
Q_MX02 U4060 ( .S(n5817), .A0(n4798), .A1(n3978), .Z(n4799));
Q_AN02 U4061 ( .A0(n5818), .A1(GFidata[82]), .Z(n4798));
Q_MX02 U4062 ( .S(n5817), .A0(n4796), .A1(n3977), .Z(n4797));
Q_AN02 U4063 ( .A0(n5818), .A1(GFidata[81]), .Z(n4796));
Q_MX02 U4064 ( .S(n5817), .A0(n4794), .A1(n3976), .Z(n4795));
Q_AN02 U4065 ( .A0(n5818), .A1(GFidata[80]), .Z(n4794));
Q_MX02 U4066 ( .S(n5817), .A0(n4792), .A1(n3975), .Z(n4793));
Q_AN02 U4067 ( .A0(n5818), .A1(GFidata[79]), .Z(n4792));
Q_MX02 U4068 ( .S(n5817), .A0(n4790), .A1(n3974), .Z(n4791));
Q_AN02 U4069 ( .A0(n5818), .A1(GFidata[78]), .Z(n4790));
Q_MX02 U4070 ( .S(n5817), .A0(n4788), .A1(n3973), .Z(n4789));
Q_AN02 U4071 ( .A0(n5818), .A1(GFidata[77]), .Z(n4788));
Q_MX02 U4072 ( .S(n5817), .A0(n4786), .A1(n3972), .Z(n4787));
Q_AN02 U4073 ( .A0(n5818), .A1(GFidata[76]), .Z(n4786));
Q_MX02 U4074 ( .S(n5817), .A0(n4784), .A1(n3971), .Z(n4785));
Q_AN02 U4075 ( .A0(n5818), .A1(GFidata[75]), .Z(n4784));
Q_MX02 U4076 ( .S(n5817), .A0(n4782), .A1(n3970), .Z(n4783));
Q_AN02 U4077 ( .A0(n5818), .A1(GFidata[74]), .Z(n4782));
Q_MX02 U4078 ( .S(n5817), .A0(n4780), .A1(n3969), .Z(n4781));
Q_AN02 U4079 ( .A0(n5818), .A1(GFidata[73]), .Z(n4780));
Q_MX02 U4080 ( .S(n5817), .A0(n4778), .A1(n3968), .Z(n4779));
Q_AN02 U4081 ( .A0(n5818), .A1(GFidata[72]), .Z(n4778));
Q_MX02 U4082 ( .S(n5817), .A0(n4776), .A1(n3967), .Z(n4777));
Q_AN02 U4083 ( .A0(n5818), .A1(GFidata[71]), .Z(n4776));
Q_MX02 U4084 ( .S(n5817), .A0(n4774), .A1(n3966), .Z(n4775));
Q_AN02 U4085 ( .A0(n5818), .A1(GFidata[70]), .Z(n4774));
Q_MX02 U4086 ( .S(n5817), .A0(n4772), .A1(n3965), .Z(n4773));
Q_AN02 U4087 ( .A0(n5818), .A1(GFidata[69]), .Z(n4772));
Q_MX02 U4088 ( .S(n5817), .A0(n4770), .A1(n3964), .Z(n4771));
Q_AN02 U4089 ( .A0(n5818), .A1(GFidata[68]), .Z(n4770));
Q_MX02 U4090 ( .S(n5817), .A0(n4768), .A1(n3963), .Z(n4769));
Q_AN02 U4091 ( .A0(n5818), .A1(GFidata[67]), .Z(n4768));
Q_MX02 U4092 ( .S(n5817), .A0(n4766), .A1(n3962), .Z(n4767));
Q_AN02 U4093 ( .A0(n5818), .A1(GFidata[66]), .Z(n4766));
Q_MX02 U4094 ( .S(n5817), .A0(n4764), .A1(n3961), .Z(n4765));
Q_AN02 U4095 ( .A0(n5818), .A1(GFidata[65]), .Z(n4764));
Q_MX02 U4096 ( .S(n5817), .A0(n4762), .A1(n3960), .Z(n4763));
Q_AN02 U4097 ( .A0(n5818), .A1(GFidata[64]), .Z(n4762));
Q_MX02 U4098 ( .S(n5817), .A0(n4760), .A1(n3958), .Z(n4761));
Q_AN02 U4099 ( .A0(n5818), .A1(GFidata[63]), .Z(n4760));
Q_MX02 U4100 ( .S(n5817), .A0(n4758), .A1(n3957), .Z(n4759));
Q_AN02 U4101 ( .A0(n5818), .A1(GFidata[62]), .Z(n4758));
Q_MX02 U4102 ( .S(n5817), .A0(n4756), .A1(n3956), .Z(n4757));
Q_AN02 U4103 ( .A0(n5818), .A1(GFidata[61]), .Z(n4756));
Q_MX02 U4104 ( .S(n5817), .A0(n4754), .A1(n3955), .Z(n4755));
Q_AN02 U4105 ( .A0(n5818), .A1(GFidata[60]), .Z(n4754));
Q_MX02 U4106 ( .S(n5817), .A0(n4752), .A1(n3954), .Z(n4753));
Q_AN02 U4107 ( .A0(n5818), .A1(GFidata[59]), .Z(n4752));
Q_MX02 U4108 ( .S(n5817), .A0(n4750), .A1(n3953), .Z(n4751));
Q_AN02 U4109 ( .A0(n5818), .A1(GFidata[58]), .Z(n4750));
Q_MX02 U4110 ( .S(n5817), .A0(n4748), .A1(n3952), .Z(n4749));
Q_AN02 U4111 ( .A0(n5818), .A1(GFidata[57]), .Z(n4748));
Q_MX02 U4112 ( .S(n5817), .A0(n4746), .A1(n3951), .Z(n4747));
Q_AN02 U4113 ( .A0(n5818), .A1(GFidata[56]), .Z(n4746));
Q_MX02 U4114 ( .S(n5817), .A0(n4744), .A1(n3950), .Z(n4745));
Q_AN02 U4115 ( .A0(n5818), .A1(GFidata[55]), .Z(n4744));
Q_MX02 U4116 ( .S(n5817), .A0(n4742), .A1(n3949), .Z(n4743));
Q_AN02 U4117 ( .A0(n5818), .A1(GFidata[54]), .Z(n4742));
Q_MX02 U4118 ( .S(n5817), .A0(n4740), .A1(n3948), .Z(n4741));
Q_AN02 U4119 ( .A0(n5818), .A1(GFidata[53]), .Z(n4740));
Q_MX02 U4120 ( .S(n5817), .A0(n4738), .A1(n3947), .Z(n4739));
Q_AN02 U4121 ( .A0(n5818), .A1(GFidata[52]), .Z(n4738));
Q_MX02 U4122 ( .S(n5817), .A0(n4736), .A1(n3946), .Z(n4737));
Q_AN02 U4123 ( .A0(n5818), .A1(GFidata[51]), .Z(n4736));
Q_MX02 U4124 ( .S(n5817), .A0(n4734), .A1(n3945), .Z(n4735));
Q_AN02 U4125 ( .A0(n5818), .A1(GFidata[50]), .Z(n4734));
Q_MX02 U4126 ( .S(n5817), .A0(n4732), .A1(n3944), .Z(n4733));
Q_AN02 U4127 ( .A0(n5818), .A1(GFidata[49]), .Z(n4732));
Q_MX02 U4128 ( .S(n5817), .A0(n4730), .A1(n3943), .Z(n4731));
Q_AN02 U4129 ( .A0(n5818), .A1(GFidata[48]), .Z(n4730));
Q_MX02 U4130 ( .S(n5817), .A0(n4728), .A1(n3942), .Z(n4729));
Q_AN02 U4131 ( .A0(n5818), .A1(GFidata[47]), .Z(n4728));
Q_MX02 U4132 ( .S(n5817), .A0(n4726), .A1(n3941), .Z(n4727));
Q_AN02 U4133 ( .A0(n5818), .A1(GFidata[46]), .Z(n4726));
Q_MX02 U4134 ( .S(n5817), .A0(n4724), .A1(n3940), .Z(n4725));
Q_AN02 U4135 ( .A0(n5818), .A1(GFidata[45]), .Z(n4724));
Q_MX02 U4136 ( .S(n5817), .A0(n4722), .A1(n3939), .Z(n4723));
Q_AN02 U4137 ( .A0(n5818), .A1(GFidata[44]), .Z(n4722));
Q_MX02 U4138 ( .S(n5817), .A0(n4720), .A1(n3938), .Z(n4721));
Q_AN02 U4139 ( .A0(n5818), .A1(GFidata[43]), .Z(n4720));
Q_MX02 U4140 ( .S(n5817), .A0(n4718), .A1(n3937), .Z(n4719));
Q_AN02 U4141 ( .A0(n5818), .A1(GFidata[42]), .Z(n4718));
Q_MX02 U4142 ( .S(n5817), .A0(n4716), .A1(n3936), .Z(n4717));
Q_AN02 U4143 ( .A0(n5818), .A1(GFidata[41]), .Z(n4716));
Q_MX02 U4144 ( .S(n5817), .A0(n4714), .A1(n3935), .Z(n4715));
Q_AN02 U4145 ( .A0(n5818), .A1(GFidata[40]), .Z(n4714));
Q_MX02 U4146 ( .S(n5817), .A0(n4712), .A1(n3934), .Z(n4713));
Q_AN02 U4147 ( .A0(n5818), .A1(GFidata[39]), .Z(n4712));
Q_MX02 U4148 ( .S(n5817), .A0(n4710), .A1(n3933), .Z(n4711));
Q_AN02 U4149 ( .A0(n5818), .A1(GFidata[38]), .Z(n4710));
Q_MX02 U4150 ( .S(n5817), .A0(n4708), .A1(n3932), .Z(n4709));
Q_AN02 U4151 ( .A0(n5818), .A1(GFidata[37]), .Z(n4708));
Q_MX02 U4152 ( .S(n5817), .A0(n4706), .A1(n3931), .Z(n4707));
Q_AN02 U4153 ( .A0(n5818), .A1(GFidata[36]), .Z(n4706));
Q_MX02 U4154 ( .S(n5817), .A0(n4704), .A1(n3930), .Z(n4705));
Q_AN02 U4155 ( .A0(n5818), .A1(GFidata[35]), .Z(n4704));
Q_MX02 U4156 ( .S(n5817), .A0(n4702), .A1(n3929), .Z(n4703));
Q_AN02 U4157 ( .A0(n5818), .A1(GFidata[34]), .Z(n4702));
Q_MX02 U4158 ( .S(n5817), .A0(n4700), .A1(n3928), .Z(n4701));
Q_AN02 U4159 ( .A0(n5818), .A1(GFidata[33]), .Z(n4700));
Q_MX02 U4160 ( .S(n5817), .A0(n4698), .A1(n3927), .Z(n4699));
Q_AN02 U4161 ( .A0(n5818), .A1(GFidata[32]), .Z(n4698));
Q_MX02 U4162 ( .S(n5817), .A0(n4696), .A1(n3926), .Z(n4697));
Q_AN02 U4163 ( .A0(n5818), .A1(GFidata[31]), .Z(n4696));
Q_MX02 U4164 ( .S(n5817), .A0(n4694), .A1(n3925), .Z(n4695));
Q_AN02 U4165 ( .A0(n5818), .A1(GFidata[30]), .Z(n4694));
Q_MX02 U4166 ( .S(n5817), .A0(n4692), .A1(n3924), .Z(n4693));
Q_AN02 U4167 ( .A0(n5818), .A1(GFidata[29]), .Z(n4692));
Q_MX02 U4168 ( .S(n5817), .A0(n4690), .A1(n3923), .Z(n4691));
Q_AN02 U4169 ( .A0(n5818), .A1(GFidata[28]), .Z(n4690));
Q_MX02 U4170 ( .S(n5817), .A0(n4688), .A1(n3922), .Z(n4689));
Q_AN02 U4171 ( .A0(n5818), .A1(GFidata[27]), .Z(n4688));
Q_MX02 U4172 ( .S(n5817), .A0(n4686), .A1(n3921), .Z(n4687));
Q_AN02 U4173 ( .A0(n5818), .A1(GFidata[26]), .Z(n4686));
Q_MX02 U4174 ( .S(n5817), .A0(n4684), .A1(n3920), .Z(n4685));
Q_AN02 U4175 ( .A0(n5818), .A1(GFidata[25]), .Z(n4684));
Q_MX02 U4176 ( .S(n5817), .A0(n4682), .A1(n3919), .Z(n4683));
Q_AN02 U4177 ( .A0(n5818), .A1(GFidata[24]), .Z(n4682));
Q_MX02 U4178 ( .S(n5817), .A0(n4680), .A1(n3918), .Z(n4681));
Q_AN02 U4179 ( .A0(n5818), .A1(GFidata[23]), .Z(n4680));
Q_MX02 U4180 ( .S(n5817), .A0(n4678), .A1(n3917), .Z(n4679));
Q_AN02 U4181 ( .A0(n5818), .A1(GFidata[22]), .Z(n4678));
Q_MX02 U4182 ( .S(n5817), .A0(n4676), .A1(n3916), .Z(n4677));
Q_AN02 U4183 ( .A0(n5818), .A1(GFidata[21]), .Z(n4676));
Q_MX02 U4184 ( .S(n5817), .A0(n4674), .A1(n3915), .Z(n4675));
Q_AN02 U4185 ( .A0(n5818), .A1(GFidata[20]), .Z(n4674));
Q_MX02 U4186 ( .S(n5817), .A0(n4672), .A1(n3914), .Z(n4673));
Q_AN02 U4187 ( .A0(n5818), .A1(GFidata[19]), .Z(n4672));
Q_MX02 U4188 ( .S(n5817), .A0(n4670), .A1(n3913), .Z(n4671));
Q_AN02 U4189 ( .A0(n5818), .A1(GFidata[18]), .Z(n4670));
Q_MX02 U4190 ( .S(n5817), .A0(n4668), .A1(n3912), .Z(n4669));
Q_AN02 U4191 ( .A0(n5818), .A1(GFidata[17]), .Z(n4668));
Q_MX02 U4192 ( .S(n5817), .A0(n4666), .A1(n3911), .Z(n4667));
Q_AN02 U4193 ( .A0(n5818), .A1(GFidata[16]), .Z(n4666));
Q_MX02 U4194 ( .S(n5817), .A0(n4664), .A1(n3910), .Z(n4665));
Q_AN02 U4195 ( .A0(n5818), .A1(GFidata[15]), .Z(n4664));
Q_MX02 U4196 ( .S(n5817), .A0(n4662), .A1(n3909), .Z(n4663));
Q_AN02 U4197 ( .A0(n5818), .A1(GFidata[14]), .Z(n4662));
Q_MX02 U4198 ( .S(n5817), .A0(n4660), .A1(n3908), .Z(n4661));
Q_AN02 U4199 ( .A0(n5818), .A1(GFidata[13]), .Z(n4660));
Q_MX02 U4200 ( .S(n5817), .A0(n4658), .A1(n3907), .Z(n4659));
Q_AN02 U4201 ( .A0(n5818), .A1(GFidata[12]), .Z(n4658));
Q_MX02 U4202 ( .S(n5817), .A0(n4656), .A1(n3906), .Z(n4657));
Q_AN02 U4203 ( .A0(n5818), .A1(GFidata[11]), .Z(n4656));
Q_MX02 U4204 ( .S(n5817), .A0(n4654), .A1(n3905), .Z(n4655));
Q_AN02 U4205 ( .A0(n5818), .A1(GFidata[10]), .Z(n4654));
Q_MX02 U4206 ( .S(n5817), .A0(n4652), .A1(n3904), .Z(n4653));
Q_AN02 U4207 ( .A0(n5818), .A1(GFidata[9]), .Z(n4652));
Q_MX02 U4208 ( .S(n5817), .A0(n4650), .A1(n3903), .Z(n4651));
Q_AN02 U4209 ( .A0(n5818), .A1(GFidata[8]), .Z(n4650));
Q_MX02 U4210 ( .S(n5817), .A0(n4648), .A1(n3902), .Z(n4649));
Q_AN02 U4211 ( .A0(n5818), .A1(GFidata[7]), .Z(n4648));
Q_MX02 U4212 ( .S(n5817), .A0(n4646), .A1(n3901), .Z(n4647));
Q_AN02 U4213 ( .A0(n5818), .A1(GFidata[6]), .Z(n4646));
Q_MX02 U4214 ( .S(n5817), .A0(n4644), .A1(n3900), .Z(n4645));
Q_AN02 U4215 ( .A0(n5818), .A1(GFidata[5]), .Z(n4644));
Q_MX02 U4216 ( .S(n5817), .A0(n4642), .A1(n3899), .Z(n4643));
Q_AN02 U4217 ( .A0(n5818), .A1(GFidata[4]), .Z(n4642));
Q_MX02 U4218 ( .S(n5817), .A0(n4640), .A1(n3898), .Z(n4641));
Q_AN02 U4219 ( .A0(n5818), .A1(GFidata[3]), .Z(n4640));
Q_MX02 U4220 ( .S(n5817), .A0(n4638), .A1(n3897), .Z(n4639));
Q_AN02 U4221 ( .A0(n5818), .A1(GFidata[2]), .Z(n4638));
Q_MX02 U4222 ( .S(n5817), .A0(n4636), .A1(n3896), .Z(n4637));
Q_AN02 U4223 ( .A0(n5818), .A1(GFidata[1]), .Z(n4636));
Q_MX02 U4224 ( .S(n5817), .A0(n4634), .A1(n3895), .Z(n4635));
Q_AN02 U4225 ( .A0(n5818), .A1(GFidata[0]), .Z(n4634));
Q_AN02 U4226 ( .A0(n6720), .A1(n4557), .Z(n4633));
Q_AN02 U4227 ( .A0(n6720), .A1(n4555), .Z(n4632));
Q_AN02 U4228 ( .A0(n6720), .A1(n4553), .Z(n4631));
Q_AN02 U4229 ( .A0(n6720), .A1(n4551), .Z(n4630));
Q_AN02 U4230 ( .A0(n6720), .A1(n4549), .Z(n4629));
Q_AN02 U4231 ( .A0(n6720), .A1(n4547), .Z(n4628));
Q_AN02 U4232 ( .A0(n6720), .A1(n4545), .Z(n4627));
Q_AN02 U4233 ( .A0(n6720), .A1(n4543), .Z(n4626));
Q_AN02 U4234 ( .A0(n6720), .A1(n4541), .Z(n4625));
Q_AN02 U4235 ( .A0(n6720), .A1(n4539), .Z(n4624));
Q_AN02 U4236 ( .A0(n6720), .A1(n4537), .Z(n4623));
Q_AN02 U4237 ( .A0(n6720), .A1(n4535), .Z(n4622));
Q_AN02 U4238 ( .A0(n6720), .A1(n4533), .Z(n4621));
Q_AN02 U4239 ( .A0(n6720), .A1(n4531), .Z(n4620));
Q_AN02 U4240 ( .A0(n6720), .A1(n4529), .Z(n4619));
Q_AN02 U4241 ( .A0(n6720), .A1(n4527), .Z(n4618));
Q_AN02 U4242 ( .A0(n6720), .A1(n4525), .Z(n4617));
Q_AN02 U4243 ( .A0(n6720), .A1(n4523), .Z(n4616));
Q_AN02 U4244 ( .A0(n6720), .A1(n4521), .Z(n4615));
Q_AN02 U4245 ( .A0(n6720), .A1(n4519), .Z(n4614));
Q_AN02 U4246 ( .A0(n6720), .A1(n4517), .Z(n4613));
Q_AN02 U4247 ( .A0(n6720), .A1(n4515), .Z(n4612));
Q_AN02 U4248 ( .A0(n6720), .A1(n4513), .Z(n4611));
Q_AN02 U4249 ( .A0(n6720), .A1(n4511), .Z(n4610));
Q_AN02 U4250 ( .A0(n6720), .A1(n4509), .Z(n4609));
Q_AN02 U4251 ( .A0(n6720), .A1(n4507), .Z(n4608));
Q_AN02 U4252 ( .A0(n6720), .A1(n4505), .Z(n4607));
Q_AN02 U4253 ( .A0(n6720), .A1(n4503), .Z(n4606));
Q_AN02 U4254 ( .A0(n6720), .A1(n4501), .Z(n4605));
Q_AN02 U4255 ( .A0(n6720), .A1(n4499), .Z(n4604));
Q_AN02 U4256 ( .A0(n6720), .A1(n4497), .Z(n4603));
Q_AN02 U4257 ( .A0(n6720), .A1(n4495), .Z(n4602));
Q_AN02 U4258 ( .A0(n6720), .A1(n4493), .Z(n4601));
Q_AN02 U4259 ( .A0(n6720), .A1(n4491), .Z(n4600));
Q_AN02 U4260 ( .A0(n6720), .A1(n4489), .Z(n4599));
Q_AN02 U4261 ( .A0(n6720), .A1(n4487), .Z(n4598));
Q_AN02 U4262 ( .A0(n6720), .A1(n4485), .Z(n4597));
Q_AN02 U4263 ( .A0(n6720), .A1(n4483), .Z(n4596));
Q_AN02 U4264 ( .A0(n6720), .A1(n4481), .Z(n4595));
Q_AN02 U4265 ( .A0(n6720), .A1(n4479), .Z(n4594));
Q_AN02 U4266 ( .A0(n6720), .A1(n4477), .Z(n4593));
Q_AN02 U4267 ( .A0(n6720), .A1(n4475), .Z(n4592));
Q_AN02 U4268 ( .A0(n6720), .A1(n4473), .Z(n4591));
Q_AN02 U4269 ( .A0(n6720), .A1(n4471), .Z(n4590));
Q_AN02 U4270 ( .A0(n6720), .A1(n4469), .Z(n4589));
Q_AN02 U4271 ( .A0(n6720), .A1(n4467), .Z(n4588));
Q_AN02 U4272 ( .A0(n6720), .A1(n4465), .Z(n4587));
Q_AN02 U4273 ( .A0(n6720), .A1(n4463), .Z(n4586));
Q_AN02 U4274 ( .A0(n6720), .A1(n4461), .Z(n4585));
Q_AN02 U4275 ( .A0(n6720), .A1(n4459), .Z(n4584));
Q_AN02 U4276 ( .A0(n6720), .A1(n4457), .Z(n4583));
Q_AN02 U4277 ( .A0(n6720), .A1(n4455), .Z(n4582));
Q_AN02 U4278 ( .A0(n6720), .A1(n4453), .Z(n4581));
Q_AN02 U4279 ( .A0(n6720), .A1(n4452), .Z(n4580));
Q_AN02 U4280 ( .A0(n6720), .A1(n4450), .Z(n4579));
Q_AN02 U4281 ( .A0(n6720), .A1(n4449), .Z(n4578));
Q_AN02 U4282 ( .A0(n6720), .A1(n4447), .Z(n4577));
Q_AN02 U4283 ( .A0(n6720), .A1(n4446), .Z(n4576));
Q_AN02 U4284 ( .A0(n6720), .A1(n4444), .Z(n4575));
Q_AN02 U4285 ( .A0(n6720), .A1(n4443), .Z(n4574));
Q_AN02 U4286 ( .A0(n6720), .A1(n4441), .Z(n4573));
Q_AN02 U4287 ( .A0(n6720), .A1(n4440), .Z(n4572));
Q_AN02 U4288 ( .A0(n6720), .A1(n4438), .Z(n4571));
Q_AN02 U4289 ( .A0(n6720), .A1(n4436), .Z(n4570));
Q_MX02 U4290 ( .S(n5818), .A0(n4568), .A1(n4423), .Z(n4569));
Q_AN02 U4291 ( .A0(n5817), .A1(n4417), .Z(n4568));
Q_MX02 U4292 ( .S(n5818), .A0(n4566), .A1(n4422), .Z(n4567));
Q_AN02 U4293 ( .A0(n5817), .A1(n4415), .Z(n4566));
Q_MX02 U4294 ( .S(n5818), .A0(n4564), .A1(n4421), .Z(n4565));
Q_AN02 U4295 ( .A0(n5817), .A1(n4413), .Z(n4564));
Q_MX02 U4296 ( .S(n5818), .A0(n4562), .A1(n4420), .Z(n4563));
Q_AN02 U4297 ( .A0(n5817), .A1(n4411), .Z(n4562));
Q_MX02 U4298 ( .S(n5818), .A0(n4560), .A1(n4419), .Z(n4561));
Q_AN02 U4299 ( .A0(n5817), .A1(n4409), .Z(n4560));
Q_MX02 U4300 ( .S(n5818), .A0(n4558), .A1(n4418), .Z(n4559));
Q_AN02 U4301 ( .A0(n5817), .A1(n4408), .Z(n4558));
Q_XOR2 U4302 ( .A0(wrtCnt[63]), .A1(n4556), .Z(n4557));
Q_AD01HF U4303 ( .A0(wrtCnt[62]), .B0(n4554), .S(n4555), .CO(n4556));
Q_AD01HF U4304 ( .A0(wrtCnt[61]), .B0(n4552), .S(n4553), .CO(n4554));
Q_AD01HF U4305 ( .A0(wrtCnt[60]), .B0(n4550), .S(n4551), .CO(n4552));
Q_AD01HF U4306 ( .A0(wrtCnt[59]), .B0(n4548), .S(n4549), .CO(n4550));
Q_AD01HF U4307 ( .A0(wrtCnt[58]), .B0(n4546), .S(n4547), .CO(n4548));
Q_AD01HF U4308 ( .A0(wrtCnt[57]), .B0(n4544), .S(n4545), .CO(n4546));
Q_AD01HF U4309 ( .A0(wrtCnt[56]), .B0(n4542), .S(n4543), .CO(n4544));
Q_AD01HF U4310 ( .A0(wrtCnt[55]), .B0(n4540), .S(n4541), .CO(n4542));
Q_AD01HF U4311 ( .A0(wrtCnt[54]), .B0(n4538), .S(n4539), .CO(n4540));
Q_AD01HF U4312 ( .A0(wrtCnt[53]), .B0(n4536), .S(n4537), .CO(n4538));
Q_AD01HF U4313 ( .A0(wrtCnt[52]), .B0(n4534), .S(n4535), .CO(n4536));
Q_AD01HF U4314 ( .A0(wrtCnt[51]), .B0(n4532), .S(n4533), .CO(n4534));
Q_AD01HF U4315 ( .A0(wrtCnt[50]), .B0(n4530), .S(n4531), .CO(n4532));
Q_AD01HF U4316 ( .A0(wrtCnt[49]), .B0(n4528), .S(n4529), .CO(n4530));
Q_AD01HF U4317 ( .A0(wrtCnt[48]), .B0(n4526), .S(n4527), .CO(n4528));
Q_AD01HF U4318 ( .A0(wrtCnt[47]), .B0(n4524), .S(n4525), .CO(n4526));
Q_AD01HF U4319 ( .A0(wrtCnt[46]), .B0(n4522), .S(n4523), .CO(n4524));
Q_AD01HF U4320 ( .A0(wrtCnt[45]), .B0(n4520), .S(n4521), .CO(n4522));
Q_AD01HF U4321 ( .A0(wrtCnt[44]), .B0(n4518), .S(n4519), .CO(n4520));
Q_AD01HF U4322 ( .A0(wrtCnt[43]), .B0(n4516), .S(n4517), .CO(n4518));
Q_AD01HF U4323 ( .A0(wrtCnt[42]), .B0(n4514), .S(n4515), .CO(n4516));
Q_AD01HF U4324 ( .A0(wrtCnt[41]), .B0(n4512), .S(n4513), .CO(n4514));
Q_AD01HF U4325 ( .A0(wrtCnt[40]), .B0(n4510), .S(n4511), .CO(n4512));
Q_AD01HF U4326 ( .A0(wrtCnt[39]), .B0(n4508), .S(n4509), .CO(n4510));
Q_AD01HF U4327 ( .A0(wrtCnt[38]), .B0(n4506), .S(n4507), .CO(n4508));
Q_AD01HF U4328 ( .A0(wrtCnt[37]), .B0(n4504), .S(n4505), .CO(n4506));
Q_AD01HF U4329 ( .A0(wrtCnt[36]), .B0(n4502), .S(n4503), .CO(n4504));
Q_AD01HF U4330 ( .A0(wrtCnt[35]), .B0(n4500), .S(n4501), .CO(n4502));
Q_AD01HF U4331 ( .A0(wrtCnt[34]), .B0(n4498), .S(n4499), .CO(n4500));
Q_AD01HF U4332 ( .A0(wrtCnt[33]), .B0(n4496), .S(n4497), .CO(n4498));
Q_AD01HF U4333 ( .A0(wrtCnt[32]), .B0(n4494), .S(n4495), .CO(n4496));
Q_AD01HF U4334 ( .A0(wrtCnt[31]), .B0(n4492), .S(n4493), .CO(n4494));
Q_AD01HF U4335 ( .A0(wrtCnt[30]), .B0(n4490), .S(n4491), .CO(n4492));
Q_AD01HF U4336 ( .A0(wrtCnt[29]), .B0(n4488), .S(n4489), .CO(n4490));
Q_AD01HF U4337 ( .A0(wrtCnt[28]), .B0(n4486), .S(n4487), .CO(n4488));
Q_AD01HF U4338 ( .A0(wrtCnt[27]), .B0(n4484), .S(n4485), .CO(n4486));
Q_AD01HF U4339 ( .A0(wrtCnt[26]), .B0(n4482), .S(n4483), .CO(n4484));
Q_AD01HF U4340 ( .A0(wrtCnt[25]), .B0(n4480), .S(n4481), .CO(n4482));
Q_AD01HF U4341 ( .A0(wrtCnt[24]), .B0(n4478), .S(n4479), .CO(n4480));
Q_AD01HF U4342 ( .A0(wrtCnt[23]), .B0(n4476), .S(n4477), .CO(n4478));
Q_AD01HF U4343 ( .A0(wrtCnt[22]), .B0(n4474), .S(n4475), .CO(n4476));
Q_AD01HF U4344 ( .A0(wrtCnt[21]), .B0(n4472), .S(n4473), .CO(n4474));
Q_AD01HF U4345 ( .A0(wrtCnt[20]), .B0(n4470), .S(n4471), .CO(n4472));
Q_AD01HF U4346 ( .A0(wrtCnt[19]), .B0(n4468), .S(n4469), .CO(n4470));
Q_AD01HF U4347 ( .A0(wrtCnt[18]), .B0(n4466), .S(n4467), .CO(n4468));
Q_AD01HF U4348 ( .A0(wrtCnt[17]), .B0(n4464), .S(n4465), .CO(n4466));
Q_AD01HF U4349 ( .A0(wrtCnt[16]), .B0(n4462), .S(n4463), .CO(n4464));
Q_AD01HF U4350 ( .A0(wrtCnt[15]), .B0(n4460), .S(n4461), .CO(n4462));
Q_AD01HF U4351 ( .A0(wrtCnt[14]), .B0(n4458), .S(n4459), .CO(n4460));
Q_AD01HF U4352 ( .A0(wrtCnt[13]), .B0(n4456), .S(n4457), .CO(n4458));
Q_AD01HF U4353 ( .A0(wrtCnt[12]), .B0(n4454), .S(n4455), .CO(n4456));
Q_AD02 U4354 ( .CI(n4451), .A0(wrtCnt[10]), .A1(wrtCnt[11]), .B0(n4434), .B1(n4435), .S0(n4452), .S1(n4453), .CO(n4454));
Q_AD02 U4355 ( .CI(n4448), .A0(wrtCnt[8]), .A1(wrtCnt[9]), .B0(n4432), .B1(n4433), .S0(n4449), .S1(n4450), .CO(n4451));
Q_AD02 U4356 ( .CI(n4445), .A0(wrtCnt[6]), .A1(wrtCnt[7]), .B0(n4430), .B1(n4431), .S0(n4446), .S1(n4447), .CO(n4448));
Q_AD02 U4357 ( .CI(n4442), .A0(wrtCnt[4]), .A1(wrtCnt[5]), .B0(n4428), .B1(n4429), .S0(n4443), .S1(n4444), .CO(n4445));
Q_AD02 U4358 ( .CI(n4439), .A0(wrtCnt[2]), .A1(wrtCnt[3]), .B0(n4426), .B1(n4427), .S0(n4440), .S1(n4441), .CO(n4442));
Q_AD01 U4359 ( .CI(n4437), .A0(wrtCnt[1]), .B0(n4425), .S(n4438), .CO(n4439));
Q_OR02 U4360 ( .A0(wrtCnt[0]), .A1(n4424), .Z(n4437));
Q_XNR2 U4361 ( .A0(wrtCnt[0]), .A1(n4424), .Z(n4436));
Q_MX02 U4362 ( .S(n3699), .A0(GFlen[11]), .A1(argLen[11]), .Z(n4435));
Q_MX02 U4363 ( .S(n3699), .A0(GFlen[10]), .A1(argLen[10]), .Z(n4434));
Q_MX02 U4364 ( .S(n3699), .A0(GFlen[9]), .A1(argLen[9]), .Z(n4433));
Q_MX02 U4365 ( .S(n3699), .A0(GFlen[8]), .A1(argLen[8]), .Z(n4432));
Q_MX02 U4366 ( .S(n3699), .A0(GFlen[7]), .A1(argLen[7]), .Z(n4431));
Q_MX02 U4367 ( .S(n3699), .A0(GFlen[6]), .A1(argLen[6]), .Z(n4430));
Q_MX02 U4368 ( .S(n3699), .A0(GFlen[5]), .A1(argLen[5]), .Z(n4429));
Q_MX02 U4369 ( .S(n3699), .A0(GFlen[4]), .A1(argLen[4]), .Z(n4428));
Q_MX02 U4370 ( .S(n3699), .A0(GFlen[3]), .A1(argLen[3]), .Z(n4427));
Q_MX02 U4371 ( .S(n3699), .A0(GFlen[2]), .A1(argLen[2]), .Z(n4426));
Q_MX02 U4372 ( .S(n3699), .A0(GFlen[1]), .A1(argLen[1]), .Z(n4425));
Q_MX02 U4373 ( .S(n3699), .A0(GFlen[0]), .A1(argLen[0]), .Z(n4424));
Q_AN02 U4374 ( .A0(n5815), .A1(GFlen[5]), .Z(n4423));
Q_OR02 U4375 ( .A0(n5823), .A1(GFlen[4]), .Z(n4422));
Q_AN02 U4376 ( .A0(n5815), .A1(GFlen[3]), .Z(n4421));
Q_AN02 U4377 ( .A0(n5815), .A1(GFlen[2]), .Z(n4420));
Q_AN02 U4378 ( .A0(n5815), .A1(GFlen[1]), .Z(n4419));
Q_AN02 U4379 ( .A0(n5815), .A1(GFlen[0]), .Z(n4418));
Q_AD01HF U4380 ( .A0(n4414), .B0(n4422), .S(n4415), .CO(n4416));
Q_AD01HF U4381 ( .A0(n4412), .B0(n4421), .S(n4413), .CO(n4414));
Q_AD01HF U4382 ( .A0(n4410), .B0(n4420), .S(n4411), .CO(n4412));
Q_AD01HF U4383 ( .A0(n4419), .B0(n4418), .S(n4409), .CO(n4410));
Q_INV U4384 ( .A(n4418), .Z(n4408));
Q_AN03 U4385 ( .A0(n3959), .A1(GFidata[511]), .A2(n5817), .Z(n5689));
Q_AN03 U4386 ( .A0(n3959), .A1(GFidata[510]), .A2(n5817), .Z(n5688));
Q_AN03 U4387 ( .A0(n3959), .A1(GFidata[509]), .A2(n5817), .Z(n5687));
Q_AN03 U4388 ( .A0(n3959), .A1(GFidata[508]), .A2(n5817), .Z(n5686));
Q_AN03 U4389 ( .A0(n3959), .A1(GFidata[507]), .A2(n5817), .Z(n5685));
Q_AN03 U4390 ( .A0(n3959), .A1(GFidata[506]), .A2(n5817), .Z(n5684));
Q_AN03 U4391 ( .A0(n3959), .A1(GFidata[505]), .A2(n5817), .Z(n5683));
Q_AN03 U4392 ( .A0(n3959), .A1(GFidata[504]), .A2(n5817), .Z(n5682));
Q_AN03 U4393 ( .A0(n3959), .A1(GFidata[503]), .A2(n5817), .Z(n5681));
Q_AN03 U4394 ( .A0(n3959), .A1(GFidata[502]), .A2(n5817), .Z(n5680));
Q_AN03 U4395 ( .A0(n3959), .A1(GFidata[501]), .A2(n5817), .Z(n5679));
Q_AN03 U4396 ( .A0(n3959), .A1(GFidata[500]), .A2(n5817), .Z(n5678));
Q_AN03 U4397 ( .A0(n3959), .A1(GFidata[499]), .A2(n5817), .Z(n5677));
Q_AN03 U4398 ( .A0(n3959), .A1(GFidata[498]), .A2(n5817), .Z(n5676));
Q_AN03 U4399 ( .A0(n3959), .A1(GFidata[497]), .A2(n5817), .Z(n5675));
Q_AN03 U4400 ( .A0(n3959), .A1(GFidata[496]), .A2(n5817), .Z(n5674));
Q_AN03 U4401 ( .A0(n3959), .A1(GFidata[495]), .A2(n5817), .Z(n5673));
Q_AN03 U4402 ( .A0(n3959), .A1(GFidata[494]), .A2(n5817), .Z(n5672));
Q_AN03 U4403 ( .A0(n3959), .A1(GFidata[493]), .A2(n5817), .Z(n5671));
Q_AN03 U4404 ( .A0(n3959), .A1(GFidata[492]), .A2(n5817), .Z(n5670));
Q_AN03 U4405 ( .A0(n3959), .A1(GFidata[491]), .A2(n5817), .Z(n5669));
Q_AN03 U4406 ( .A0(n3959), .A1(GFidata[490]), .A2(n5817), .Z(n5668));
Q_AN03 U4407 ( .A0(n3959), .A1(GFidata[489]), .A2(n5817), .Z(n5667));
Q_AN03 U4408 ( .A0(n3959), .A1(GFidata[488]), .A2(n5817), .Z(n5666));
Q_AN03 U4409 ( .A0(n3959), .A1(GFidata[487]), .A2(n5817), .Z(n5665));
Q_AN03 U4410 ( .A0(n3959), .A1(GFidata[486]), .A2(n5817), .Z(n5664));
Q_AN03 U4411 ( .A0(n3959), .A1(GFidata[485]), .A2(n5817), .Z(n5663));
Q_AN03 U4412 ( .A0(n3959), .A1(GFidata[484]), .A2(n5817), .Z(n5662));
Q_AN03 U4413 ( .A0(n3959), .A1(GFidata[483]), .A2(n5817), .Z(n5661));
Q_AN03 U4414 ( .A0(n3959), .A1(GFidata[482]), .A2(n5817), .Z(n5660));
Q_AN03 U4415 ( .A0(n3959), .A1(GFidata[481]), .A2(n5817), .Z(n5659));
Q_AN03 U4416 ( .A0(n3959), .A1(GFidata[480]), .A2(n5817), .Z(n5658));
Q_AN02 U4417 ( .A0(n3959), .A1(GFidata[479]), .Z(n4407));
Q_AN02 U4418 ( .A0(n3959), .A1(GFidata[478]), .Z(n4406));
Q_AN02 U4419 ( .A0(n3959), .A1(GFidata[477]), .Z(n4405));
Q_AN02 U4420 ( .A0(n3959), .A1(GFidata[476]), .Z(n4404));
Q_AN02 U4421 ( .A0(n3959), .A1(GFidata[475]), .Z(n4403));
Q_AN02 U4422 ( .A0(n3959), .A1(GFidata[474]), .Z(n4402));
Q_AN02 U4423 ( .A0(n3959), .A1(GFidata[473]), .Z(n4401));
Q_AN02 U4424 ( .A0(n3959), .A1(GFidata[472]), .Z(n4400));
Q_AN02 U4425 ( .A0(n3959), .A1(GFidata[471]), .Z(n4399));
Q_AN02 U4426 ( .A0(n3959), .A1(GFidata[470]), .Z(n4398));
Q_AN02 U4427 ( .A0(n3959), .A1(GFidata[469]), .Z(n4397));
Q_AN02 U4428 ( .A0(n3959), .A1(GFidata[468]), .Z(n4396));
Q_AN02 U4429 ( .A0(n3959), .A1(GFidata[467]), .Z(n4395));
Q_AN02 U4430 ( .A0(n3959), .A1(GFidata[466]), .Z(n4394));
Q_AN02 U4431 ( .A0(n3959), .A1(GFidata[465]), .Z(n4393));
Q_AN02 U4432 ( .A0(n3959), .A1(GFidata[464]), .Z(n4392));
Q_AN02 U4433 ( .A0(n3959), .A1(GFidata[463]), .Z(n4391));
Q_AN02 U4434 ( .A0(n3959), .A1(GFidata[462]), .Z(n4390));
Q_AN02 U4435 ( .A0(n3959), .A1(GFidata[461]), .Z(n4389));
Q_AN02 U4436 ( .A0(n3959), .A1(GFidata[460]), .Z(n4388));
Q_AN02 U4437 ( .A0(n3959), .A1(GFidata[459]), .Z(n4387));
Q_AN02 U4438 ( .A0(n3959), .A1(GFidata[458]), .Z(n4386));
Q_AN02 U4439 ( .A0(n3959), .A1(GFidata[457]), .Z(n4385));
Q_AN02 U4440 ( .A0(n3959), .A1(GFidata[456]), .Z(n4384));
Q_AN02 U4441 ( .A0(n3959), .A1(GFidata[455]), .Z(n4383));
Q_AN02 U4442 ( .A0(n3959), .A1(GFidata[454]), .Z(n4382));
Q_AN02 U4443 ( .A0(n3959), .A1(GFidata[453]), .Z(n4381));
Q_AN02 U4444 ( .A0(n3959), .A1(GFidata[452]), .Z(n4380));
Q_AN02 U4445 ( .A0(n3959), .A1(GFidata[451]), .Z(n4379));
Q_AN02 U4446 ( .A0(n3959), .A1(GFidata[450]), .Z(n4378));
Q_AN02 U4447 ( .A0(n3959), .A1(GFidata[449]), .Z(n4377));
Q_AN02 U4448 ( .A0(n3959), .A1(GFidata[448]), .Z(n4376));
Q_AN02 U4449 ( .A0(n3959), .A1(GFidata[447]), .Z(n4375));
Q_AN02 U4450 ( .A0(n3959), .A1(GFidata[446]), .Z(n4374));
Q_AN02 U4451 ( .A0(n3959), .A1(GFidata[445]), .Z(n4373));
Q_AN02 U4452 ( .A0(n3959), .A1(GFidata[444]), .Z(n4372));
Q_AN02 U4453 ( .A0(n3959), .A1(GFidata[443]), .Z(n4371));
Q_AN02 U4454 ( .A0(n3959), .A1(GFidata[442]), .Z(n4370));
Q_AN02 U4455 ( .A0(n3959), .A1(GFidata[441]), .Z(n4369));
Q_AN02 U4456 ( .A0(n3959), .A1(GFidata[440]), .Z(n4368));
Q_AN02 U4457 ( .A0(n3959), .A1(GFidata[439]), .Z(n4367));
Q_AN02 U4458 ( .A0(n3959), .A1(GFidata[438]), .Z(n4366));
Q_AN02 U4459 ( .A0(n3959), .A1(GFidata[437]), .Z(n4365));
Q_AN02 U4460 ( .A0(n3959), .A1(GFidata[436]), .Z(n4364));
Q_AN02 U4461 ( .A0(n3959), .A1(GFidata[435]), .Z(n4363));
Q_AN02 U4462 ( .A0(n3959), .A1(GFidata[434]), .Z(n4362));
Q_AN02 U4463 ( .A0(n3959), .A1(GFidata[433]), .Z(n4361));
Q_AN02 U4464 ( .A0(n3959), .A1(GFidata[432]), .Z(n4360));
Q_AN02 U4465 ( .A0(n3959), .A1(GFidata[431]), .Z(n4359));
Q_AN02 U4466 ( .A0(n3959), .A1(GFidata[430]), .Z(n4358));
Q_AN02 U4467 ( .A0(n3959), .A1(GFidata[429]), .Z(n4357));
Q_AN02 U4468 ( .A0(n3959), .A1(GFidata[428]), .Z(n4356));
Q_AN02 U4469 ( .A0(n3959), .A1(GFidata[427]), .Z(n4355));
Q_AN02 U4470 ( .A0(n3959), .A1(GFidata[426]), .Z(n4354));
Q_AN02 U4471 ( .A0(n3959), .A1(GFidata[425]), .Z(n4353));
Q_AN02 U4472 ( .A0(n3959), .A1(GFidata[424]), .Z(n4352));
Q_AN02 U4473 ( .A0(n3959), .A1(GFidata[423]), .Z(n4351));
Q_AN02 U4474 ( .A0(n3959), .A1(GFidata[422]), .Z(n4350));
Q_AN02 U4475 ( .A0(n3959), .A1(GFidata[421]), .Z(n4349));
Q_AN02 U4476 ( .A0(n3959), .A1(GFidata[420]), .Z(n4348));
Q_AN02 U4477 ( .A0(n3959), .A1(GFidata[419]), .Z(n4347));
Q_AN02 U4478 ( .A0(n3959), .A1(GFidata[418]), .Z(n4346));
Q_AN02 U4479 ( .A0(n3959), .A1(GFidata[417]), .Z(n4345));
Q_AN02 U4480 ( .A0(n3959), .A1(GFidata[416]), .Z(n4344));
Q_AN02 U4481 ( .A0(n3959), .A1(GFidata[415]), .Z(n4343));
Q_AN02 U4482 ( .A0(n3959), .A1(GFidata[414]), .Z(n4342));
Q_AN02 U4483 ( .A0(n3959), .A1(GFidata[413]), .Z(n4341));
Q_AN02 U4484 ( .A0(n3959), .A1(GFidata[412]), .Z(n4340));
Q_AN02 U4485 ( .A0(n3959), .A1(GFidata[411]), .Z(n4339));
Q_AN02 U4486 ( .A0(n3959), .A1(GFidata[410]), .Z(n4338));
Q_AN02 U4487 ( .A0(n3959), .A1(GFidata[409]), .Z(n4337));
Q_AN02 U4488 ( .A0(n3959), .A1(GFidata[408]), .Z(n4336));
Q_AN02 U4489 ( .A0(n3959), .A1(GFidata[407]), .Z(n4335));
Q_AN02 U4490 ( .A0(n3959), .A1(GFidata[406]), .Z(n4334));
Q_AN02 U4491 ( .A0(n3959), .A1(GFidata[405]), .Z(n4333));
Q_AN02 U4492 ( .A0(n3959), .A1(GFidata[404]), .Z(n4332));
Q_AN02 U4493 ( .A0(n3959), .A1(GFidata[403]), .Z(n4331));
Q_AN02 U4494 ( .A0(n3959), .A1(GFidata[402]), .Z(n4330));
Q_AN02 U4495 ( .A0(n3959), .A1(GFidata[401]), .Z(n4329));
Q_AN02 U4496 ( .A0(n3959), .A1(GFidata[400]), .Z(n4328));
Q_AN02 U4497 ( .A0(n3959), .A1(GFidata[399]), .Z(n4327));
Q_AN02 U4498 ( .A0(n3959), .A1(GFidata[398]), .Z(n4326));
Q_AN02 U4499 ( .A0(n3959), .A1(GFidata[397]), .Z(n4325));
Q_AN02 U4500 ( .A0(n3959), .A1(GFidata[396]), .Z(n4324));
Q_AN02 U4501 ( .A0(n3959), .A1(GFidata[395]), .Z(n4323));
Q_AN02 U4502 ( .A0(n3959), .A1(GFidata[394]), .Z(n4322));
Q_AN02 U4503 ( .A0(n3959), .A1(GFidata[393]), .Z(n4321));
Q_AN02 U4504 ( .A0(n3959), .A1(GFidata[392]), .Z(n4320));
Q_AN02 U4505 ( .A0(n3959), .A1(GFidata[391]), .Z(n4319));
Q_AN02 U4506 ( .A0(n3959), .A1(GFidata[390]), .Z(n4318));
Q_AN02 U4507 ( .A0(n3959), .A1(GFidata[389]), .Z(n4317));
Q_AN02 U4508 ( .A0(n3959), .A1(GFidata[388]), .Z(n4316));
Q_AN02 U4509 ( .A0(n3959), .A1(GFidata[387]), .Z(n4315));
Q_AN02 U4510 ( .A0(n3959), .A1(GFidata[386]), .Z(n4314));
Q_AN02 U4511 ( .A0(n3959), .A1(GFidata[385]), .Z(n4313));
Q_AN02 U4512 ( .A0(n3959), .A1(GFidata[384]), .Z(n4312));
Q_AN02 U4513 ( .A0(n3959), .A1(GFidata[383]), .Z(n4311));
Q_AN02 U4514 ( .A0(n3959), .A1(GFidata[382]), .Z(n4310));
Q_AN02 U4515 ( .A0(n3959), .A1(GFidata[381]), .Z(n4309));
Q_AN02 U4516 ( .A0(n3959), .A1(GFidata[380]), .Z(n4308));
Q_AN02 U4517 ( .A0(n3959), .A1(GFidata[379]), .Z(n4307));
Q_AN02 U4518 ( .A0(n3959), .A1(GFidata[378]), .Z(n4306));
Q_AN02 U4519 ( .A0(n3959), .A1(GFidata[377]), .Z(n4305));
Q_AN02 U4520 ( .A0(n3959), .A1(GFidata[376]), .Z(n4304));
Q_AN02 U4521 ( .A0(n3959), .A1(GFidata[375]), .Z(n4303));
Q_AN02 U4522 ( .A0(n3959), .A1(GFidata[374]), .Z(n4302));
Q_AN02 U4523 ( .A0(n3959), .A1(GFidata[373]), .Z(n4301));
Q_AN02 U4524 ( .A0(n3959), .A1(GFidata[372]), .Z(n4300));
Q_AN02 U4525 ( .A0(n3959), .A1(GFidata[371]), .Z(n4299));
Q_AN02 U4526 ( .A0(n3959), .A1(GFidata[370]), .Z(n4298));
Q_AN02 U4527 ( .A0(n3959), .A1(GFidata[369]), .Z(n4297));
Q_AN02 U4528 ( .A0(n3959), .A1(GFidata[368]), .Z(n4296));
Q_AN02 U4529 ( .A0(n3959), .A1(GFidata[367]), .Z(n4295));
Q_AN02 U4530 ( .A0(n3959), .A1(GFidata[366]), .Z(n4294));
Q_AN02 U4531 ( .A0(n3959), .A1(GFidata[365]), .Z(n4293));
Q_AN02 U4532 ( .A0(n3959), .A1(GFidata[364]), .Z(n4292));
Q_AN02 U4533 ( .A0(n3959), .A1(GFidata[363]), .Z(n4291));
Q_AN02 U4534 ( .A0(n3959), .A1(GFidata[362]), .Z(n4290));
Q_AN02 U4535 ( .A0(n3959), .A1(GFidata[361]), .Z(n4289));
Q_AN02 U4536 ( .A0(n3959), .A1(GFidata[360]), .Z(n4288));
Q_AN02 U4537 ( .A0(n3959), .A1(GFidata[359]), .Z(n4287));
Q_AN02 U4538 ( .A0(n3959), .A1(GFidata[358]), .Z(n4286));
Q_AN02 U4539 ( .A0(n3959), .A1(GFidata[357]), .Z(n4285));
Q_AN02 U4540 ( .A0(n3959), .A1(GFidata[356]), .Z(n4284));
Q_AN02 U4541 ( .A0(n3959), .A1(GFidata[355]), .Z(n4283));
Q_AN02 U4542 ( .A0(n3959), .A1(GFidata[354]), .Z(n4282));
Q_AN02 U4543 ( .A0(n3959), .A1(GFidata[353]), .Z(n4281));
Q_AN02 U4544 ( .A0(n3959), .A1(GFidata[352]), .Z(n4280));
Q_AN02 U4545 ( .A0(n3959), .A1(GFidata[351]), .Z(n4279));
Q_AN02 U4546 ( .A0(n3959), .A1(GFidata[350]), .Z(n4278));
Q_AN02 U4547 ( .A0(n3959), .A1(GFidata[349]), .Z(n4277));
Q_AN02 U4548 ( .A0(n3959), .A1(GFidata[348]), .Z(n4276));
Q_AN02 U4549 ( .A0(n3959), .A1(GFidata[347]), .Z(n4275));
Q_AN02 U4550 ( .A0(n3959), .A1(GFidata[346]), .Z(n4274));
Q_AN02 U4551 ( .A0(n3959), .A1(GFidata[345]), .Z(n4273));
Q_AN02 U4552 ( .A0(n3959), .A1(GFidata[344]), .Z(n4272));
Q_AN02 U4553 ( .A0(n3959), .A1(GFidata[343]), .Z(n4271));
Q_AN02 U4554 ( .A0(n3959), .A1(GFidata[342]), .Z(n4270));
Q_AN02 U4555 ( .A0(n3959), .A1(GFidata[341]), .Z(n4269));
Q_AN02 U4556 ( .A0(n3959), .A1(GFidata[340]), .Z(n4268));
Q_AN02 U4557 ( .A0(n3959), .A1(GFidata[339]), .Z(n4267));
Q_AN02 U4558 ( .A0(n3959), .A1(GFidata[338]), .Z(n4266));
Q_AN02 U4559 ( .A0(n3959), .A1(GFidata[337]), .Z(n4265));
Q_AN02 U4560 ( .A0(n3959), .A1(GFidata[336]), .Z(n4264));
Q_AN02 U4561 ( .A0(n3959), .A1(GFidata[335]), .Z(n4263));
Q_AN02 U4562 ( .A0(n3959), .A1(GFidata[334]), .Z(n4262));
Q_AN02 U4563 ( .A0(n3959), .A1(GFidata[333]), .Z(n4261));
Q_AN02 U4564 ( .A0(n3959), .A1(GFidata[332]), .Z(n4260));
Q_AN02 U4565 ( .A0(n3959), .A1(GFidata[331]), .Z(n4259));
Q_AN02 U4566 ( .A0(n3959), .A1(GFidata[330]), .Z(n4258));
Q_AN02 U4567 ( .A0(n3959), .A1(GFidata[329]), .Z(n4257));
Q_AN02 U4568 ( .A0(n3959), .A1(GFidata[328]), .Z(n4256));
Q_AN02 U4569 ( .A0(n3959), .A1(GFidata[327]), .Z(n4255));
Q_AN02 U4570 ( .A0(n3959), .A1(GFidata[326]), .Z(n4254));
Q_AN02 U4571 ( .A0(n3959), .A1(GFidata[325]), .Z(n4253));
Q_AN02 U4572 ( .A0(n3959), .A1(GFidata[324]), .Z(n4252));
Q_AN02 U4573 ( .A0(n3959), .A1(GFidata[323]), .Z(n4251));
Q_AN02 U4574 ( .A0(n3959), .A1(GFidata[322]), .Z(n4250));
Q_AN02 U4575 ( .A0(n3959), .A1(GFidata[321]), .Z(n4249));
Q_AN02 U4576 ( .A0(n3959), .A1(GFidata[320]), .Z(n4248));
Q_AN02 U4577 ( .A0(n3959), .A1(GFidata[319]), .Z(n4247));
Q_AN02 U4578 ( .A0(n3959), .A1(GFidata[318]), .Z(n4246));
Q_AN02 U4579 ( .A0(n3959), .A1(GFidata[317]), .Z(n4245));
Q_AN02 U4580 ( .A0(n3959), .A1(GFidata[316]), .Z(n4244));
Q_AN02 U4581 ( .A0(n3959), .A1(GFidata[315]), .Z(n4243));
Q_AN02 U4582 ( .A0(n3959), .A1(GFidata[314]), .Z(n4242));
Q_AN02 U4583 ( .A0(n3959), .A1(GFidata[313]), .Z(n4241));
Q_AN02 U4584 ( .A0(n3959), .A1(GFidata[312]), .Z(n4240));
Q_AN02 U4585 ( .A0(n3959), .A1(GFidata[311]), .Z(n4239));
Q_AN02 U4586 ( .A0(n3959), .A1(GFidata[310]), .Z(n4238));
Q_AN02 U4587 ( .A0(n3959), .A1(GFidata[309]), .Z(n4237));
Q_AN02 U4588 ( .A0(n3959), .A1(GFidata[308]), .Z(n4236));
Q_AN02 U4589 ( .A0(n3959), .A1(GFidata[307]), .Z(n4235));
Q_AN02 U4590 ( .A0(n3959), .A1(GFidata[306]), .Z(n4234));
Q_AN02 U4591 ( .A0(n3959), .A1(GFidata[305]), .Z(n4233));
Q_AN02 U4592 ( .A0(n3959), .A1(GFidata[304]), .Z(n4232));
Q_AN02 U4593 ( .A0(n3959), .A1(GFidata[303]), .Z(n4231));
Q_AN02 U4594 ( .A0(n3959), .A1(GFidata[302]), .Z(n4230));
Q_AN02 U4595 ( .A0(n3959), .A1(GFidata[301]), .Z(n4229));
Q_AN02 U4596 ( .A0(n3959), .A1(GFidata[300]), .Z(n4228));
Q_AN02 U4597 ( .A0(n3959), .A1(GFidata[299]), .Z(n4227));
Q_AN02 U4598 ( .A0(n3959), .A1(GFidata[298]), .Z(n4226));
Q_AN02 U4599 ( .A0(n3959), .A1(GFidata[297]), .Z(n4225));
Q_AN02 U4600 ( .A0(n3959), .A1(GFidata[296]), .Z(n4224));
Q_AN02 U4601 ( .A0(n3959), .A1(GFidata[295]), .Z(n4223));
Q_AN02 U4602 ( .A0(n3959), .A1(GFidata[294]), .Z(n4222));
Q_AN02 U4603 ( .A0(n3959), .A1(GFidata[293]), .Z(n4221));
Q_AN02 U4604 ( .A0(n3959), .A1(GFidata[292]), .Z(n4220));
Q_AN02 U4605 ( .A0(n3959), .A1(GFidata[291]), .Z(n4219));
Q_AN02 U4606 ( .A0(n3959), .A1(GFidata[290]), .Z(n4218));
Q_AN02 U4607 ( .A0(n3959), .A1(GFidata[289]), .Z(n4217));
Q_AN02 U4608 ( .A0(n3959), .A1(GFidata[288]), .Z(n4216));
Q_AN02 U4609 ( .A0(n3959), .A1(GFidata[287]), .Z(n4215));
Q_AN02 U4610 ( .A0(n3959), .A1(GFidata[286]), .Z(n4214));
Q_AN02 U4611 ( .A0(n3959), .A1(GFidata[285]), .Z(n4213));
Q_AN02 U4612 ( .A0(n3959), .A1(GFidata[284]), .Z(n4212));
Q_AN02 U4613 ( .A0(n3959), .A1(GFidata[283]), .Z(n4211));
Q_AN02 U4614 ( .A0(n3959), .A1(GFidata[282]), .Z(n4210));
Q_AN02 U4615 ( .A0(n3959), .A1(GFidata[281]), .Z(n4209));
Q_AN02 U4616 ( .A0(n3959), .A1(GFidata[280]), .Z(n4208));
Q_AN02 U4617 ( .A0(n3959), .A1(GFidata[279]), .Z(n4207));
Q_AN02 U4618 ( .A0(n3959), .A1(GFidata[278]), .Z(n4206));
Q_AN02 U4619 ( .A0(n3959), .A1(GFidata[277]), .Z(n4205));
Q_AN02 U4620 ( .A0(n3959), .A1(GFidata[276]), .Z(n4204));
Q_AN02 U4621 ( .A0(n3959), .A1(GFidata[275]), .Z(n4203));
Q_AN02 U4622 ( .A0(n3959), .A1(GFidata[274]), .Z(n4202));
Q_AN02 U4623 ( .A0(n3959), .A1(GFidata[273]), .Z(n4201));
Q_AN02 U4624 ( .A0(n3959), .A1(GFidata[272]), .Z(n4200));
Q_AN02 U4625 ( .A0(n3959), .A1(GFidata[271]), .Z(n4199));
Q_AN02 U4626 ( .A0(n3959), .A1(GFidata[270]), .Z(n4198));
Q_AN02 U4627 ( .A0(n3959), .A1(GFidata[269]), .Z(n4197));
Q_AN02 U4628 ( .A0(n3959), .A1(GFidata[268]), .Z(n4196));
Q_AN02 U4629 ( .A0(n3959), .A1(GFidata[267]), .Z(n4195));
Q_AN02 U4630 ( .A0(n3959), .A1(GFidata[266]), .Z(n4194));
Q_AN02 U4631 ( .A0(n3959), .A1(GFidata[265]), .Z(n4193));
Q_AN02 U4632 ( .A0(n3959), .A1(GFidata[264]), .Z(n4192));
Q_AN02 U4633 ( .A0(n3959), .A1(GFidata[263]), .Z(n4191));
Q_AN02 U4634 ( .A0(n3959), .A1(GFidata[262]), .Z(n4190));
Q_AN02 U4635 ( .A0(n3959), .A1(GFidata[261]), .Z(n4189));
Q_AN02 U4636 ( .A0(n3959), .A1(GFidata[260]), .Z(n4188));
Q_AN02 U4637 ( .A0(n3959), .A1(GFidata[259]), .Z(n4187));
Q_AN02 U4638 ( .A0(n3959), .A1(GFidata[258]), .Z(n4186));
Q_AN02 U4639 ( .A0(n3959), .A1(GFidata[257]), .Z(n4185));
Q_AN02 U4640 ( .A0(n3959), .A1(GFidata[256]), .Z(n4184));
Q_AN02 U4641 ( .A0(n3959), .A1(GFidata[255]), .Z(n4183));
Q_AN02 U4642 ( .A0(n3959), .A1(GFidata[254]), .Z(n4182));
Q_AN02 U4643 ( .A0(n3959), .A1(GFidata[253]), .Z(n4181));
Q_AN02 U4644 ( .A0(n3959), .A1(GFidata[252]), .Z(n4180));
Q_AN02 U4645 ( .A0(n3959), .A1(GFidata[251]), .Z(n4179));
Q_AN02 U4646 ( .A0(n3959), .A1(GFidata[250]), .Z(n4178));
Q_AN02 U4647 ( .A0(n3959), .A1(GFidata[249]), .Z(n4177));
Q_AN02 U4648 ( .A0(n3959), .A1(GFidata[248]), .Z(n4176));
Q_AN02 U4649 ( .A0(n3959), .A1(GFidata[247]), .Z(n4175));
Q_AN02 U4650 ( .A0(n3959), .A1(GFidata[246]), .Z(n4174));
Q_AN02 U4651 ( .A0(n3959), .A1(GFidata[245]), .Z(n4173));
Q_AN02 U4652 ( .A0(n3959), .A1(GFidata[244]), .Z(n4172));
Q_AN02 U4653 ( .A0(n3959), .A1(GFidata[243]), .Z(n4171));
Q_AN02 U4654 ( .A0(n3959), .A1(GFidata[242]), .Z(n4170));
Q_AN02 U4655 ( .A0(n3959), .A1(GFidata[241]), .Z(n4169));
Q_AN02 U4656 ( .A0(n3959), .A1(GFidata[240]), .Z(n4168));
Q_AN02 U4657 ( .A0(n3959), .A1(GFidata[239]), .Z(n4167));
Q_AN02 U4658 ( .A0(n3959), .A1(GFidata[238]), .Z(n4166));
Q_AN02 U4659 ( .A0(n3959), .A1(GFidata[237]), .Z(n4165));
Q_AN02 U4660 ( .A0(n3959), .A1(GFidata[236]), .Z(n4164));
Q_AN02 U4661 ( .A0(n3959), .A1(GFidata[235]), .Z(n4163));
Q_AN02 U4662 ( .A0(n3959), .A1(GFidata[234]), .Z(n4162));
Q_AN02 U4663 ( .A0(n3959), .A1(GFidata[233]), .Z(n4161));
Q_AN02 U4664 ( .A0(n3959), .A1(GFidata[232]), .Z(n4160));
Q_AN02 U4665 ( .A0(n3959), .A1(GFidata[231]), .Z(n4159));
Q_AN02 U4666 ( .A0(n3959), .A1(GFidata[230]), .Z(n4158));
Q_AN02 U4667 ( .A0(n3959), .A1(GFidata[229]), .Z(n4157));
Q_AN02 U4668 ( .A0(n3959), .A1(GFidata[228]), .Z(n4156));
Q_AN02 U4669 ( .A0(n3959), .A1(GFidata[227]), .Z(n4155));
Q_AN02 U4670 ( .A0(n3959), .A1(GFidata[226]), .Z(n4154));
Q_AN02 U4671 ( .A0(n3959), .A1(GFidata[225]), .Z(n4153));
Q_AN02 U4672 ( .A0(n3959), .A1(GFidata[224]), .Z(n4152));
Q_AN02 U4673 ( .A0(n3959), .A1(GFidata[223]), .Z(n4151));
Q_AN02 U4674 ( .A0(n3959), .A1(GFidata[222]), .Z(n4150));
Q_AN02 U4675 ( .A0(n3959), .A1(GFidata[221]), .Z(n4149));
Q_AN02 U4676 ( .A0(n3959), .A1(GFidata[220]), .Z(n4148));
Q_AN02 U4677 ( .A0(n3959), .A1(GFidata[219]), .Z(n4147));
Q_AN02 U4678 ( .A0(n3959), .A1(GFidata[218]), .Z(n4146));
Q_AN02 U4679 ( .A0(n3959), .A1(GFidata[217]), .Z(n4145));
Q_AN02 U4680 ( .A0(n3959), .A1(GFidata[216]), .Z(n4144));
Q_AN02 U4681 ( .A0(n3959), .A1(GFidata[215]), .Z(n4143));
Q_AN02 U4682 ( .A0(n3959), .A1(GFidata[214]), .Z(n4142));
Q_AN02 U4683 ( .A0(n3959), .A1(GFidata[213]), .Z(n4141));
Q_AN02 U4684 ( .A0(n3959), .A1(GFidata[212]), .Z(n4140));
Q_AN02 U4685 ( .A0(n3959), .A1(GFidata[211]), .Z(n4139));
Q_AN02 U4686 ( .A0(n3959), .A1(GFidata[210]), .Z(n4138));
Q_AN02 U4687 ( .A0(n3959), .A1(GFidata[209]), .Z(n4137));
Q_AN02 U4688 ( .A0(n3959), .A1(GFidata[208]), .Z(n4136));
Q_AN02 U4689 ( .A0(n3959), .A1(GFidata[207]), .Z(n4135));
Q_AN02 U4690 ( .A0(n3959), .A1(GFidata[206]), .Z(n4134));
Q_AN02 U4691 ( .A0(n3959), .A1(GFidata[205]), .Z(n4133));
Q_AN02 U4692 ( .A0(n3959), .A1(GFidata[204]), .Z(n4132));
Q_AN02 U4693 ( .A0(n3959), .A1(GFidata[203]), .Z(n4131));
Q_AN02 U4694 ( .A0(n3959), .A1(GFidata[202]), .Z(n4130));
Q_AN02 U4695 ( .A0(n3959), .A1(GFidata[201]), .Z(n4129));
Q_AN02 U4696 ( .A0(n3959), .A1(GFidata[200]), .Z(n4128));
Q_AN02 U4697 ( .A0(n3959), .A1(GFidata[199]), .Z(n4127));
Q_AN02 U4698 ( .A0(n3959), .A1(GFidata[198]), .Z(n4126));
Q_AN02 U4699 ( .A0(n3959), .A1(GFidata[197]), .Z(n4125));
Q_AN02 U4700 ( .A0(n3959), .A1(GFidata[196]), .Z(n4124));
Q_AN02 U4701 ( .A0(n3959), .A1(GFidata[195]), .Z(n4123));
Q_AN02 U4702 ( .A0(n3959), .A1(GFidata[194]), .Z(n4122));
Q_AN02 U4703 ( .A0(n3959), .A1(GFidata[193]), .Z(n4121));
Q_AN02 U4704 ( .A0(n3959), .A1(GFidata[192]), .Z(n4120));
Q_AN02 U4705 ( .A0(n3959), .A1(GFidata[191]), .Z(n4119));
Q_AN02 U4706 ( .A0(n3959), .A1(GFidata[190]), .Z(n4118));
Q_AN02 U4707 ( .A0(n3959), .A1(GFidata[189]), .Z(n4117));
Q_AN02 U4708 ( .A0(n3959), .A1(GFidata[188]), .Z(n4116));
Q_AN02 U4709 ( .A0(n3959), .A1(GFidata[187]), .Z(n4115));
Q_AN02 U4710 ( .A0(n3959), .A1(GFidata[186]), .Z(n4114));
Q_AN02 U4711 ( .A0(n3959), .A1(GFidata[185]), .Z(n4113));
Q_AN02 U4712 ( .A0(n3959), .A1(GFidata[184]), .Z(n4112));
Q_AN02 U4713 ( .A0(n3959), .A1(GFidata[183]), .Z(n4111));
Q_AN02 U4714 ( .A0(n3959), .A1(GFidata[182]), .Z(n4110));
Q_AN02 U4715 ( .A0(n3959), .A1(GFidata[181]), .Z(n4109));
Q_AN02 U4716 ( .A0(n3959), .A1(GFidata[180]), .Z(n4108));
Q_AN02 U4717 ( .A0(n3959), .A1(GFidata[179]), .Z(n4107));
Q_AN02 U4718 ( .A0(n3959), .A1(GFidata[178]), .Z(n4106));
Q_AN02 U4719 ( .A0(n3959), .A1(GFidata[177]), .Z(n4105));
Q_AN02 U4720 ( .A0(n3959), .A1(GFidata[176]), .Z(n4104));
Q_AN02 U4721 ( .A0(n3959), .A1(GFidata[175]), .Z(n4103));
Q_AN02 U4722 ( .A0(n3959), .A1(GFidata[174]), .Z(n4102));
Q_AN02 U4723 ( .A0(n3959), .A1(GFidata[173]), .Z(n4101));
Q_AN02 U4724 ( .A0(n3959), .A1(GFidata[172]), .Z(n4100));
Q_AN02 U4725 ( .A0(n3959), .A1(GFidata[171]), .Z(n4099));
Q_AN02 U4726 ( .A0(n3959), .A1(GFidata[170]), .Z(n4098));
Q_AN02 U4727 ( .A0(n3959), .A1(GFidata[169]), .Z(n4097));
Q_AN02 U4728 ( .A0(n3959), .A1(GFidata[168]), .Z(n4096));
Q_AN02 U4729 ( .A0(n3959), .A1(GFidata[167]), .Z(n4095));
Q_AN02 U4730 ( .A0(n3959), .A1(GFidata[166]), .Z(n4094));
Q_AN02 U4731 ( .A0(n3959), .A1(GFidata[165]), .Z(n4093));
Q_AN02 U4732 ( .A0(n3959), .A1(GFidata[164]), .Z(n4092));
Q_AN02 U4733 ( .A0(n3959), .A1(GFidata[163]), .Z(n4091));
Q_AN02 U4734 ( .A0(n3959), .A1(GFidata[162]), .Z(n4090));
Q_AN02 U4735 ( .A0(n3959), .A1(GFidata[161]), .Z(n4089));
Q_AN02 U4736 ( .A0(n3959), .A1(GFidata[160]), .Z(n4088));
Q_AN02 U4737 ( .A0(n3959), .A1(GFidata[159]), .Z(n4087));
Q_AN02 U4738 ( .A0(n3959), .A1(GFidata[158]), .Z(n4086));
Q_AN02 U4739 ( .A0(n3959), .A1(GFidata[157]), .Z(n4085));
Q_AN02 U4740 ( .A0(n3959), .A1(GFidata[156]), .Z(n4084));
Q_AN02 U4741 ( .A0(n3959), .A1(GFidata[155]), .Z(n4083));
Q_AN02 U4742 ( .A0(n3959), .A1(GFidata[154]), .Z(n4082));
Q_AN02 U4743 ( .A0(n3959), .A1(GFidata[153]), .Z(n4081));
Q_AN02 U4744 ( .A0(n3959), .A1(GFidata[152]), .Z(n4080));
Q_AN02 U4745 ( .A0(n3959), .A1(GFidata[151]), .Z(n4079));
Q_AN02 U4746 ( .A0(n3959), .A1(GFidata[150]), .Z(n4078));
Q_AN02 U4747 ( .A0(n3959), .A1(GFidata[149]), .Z(n4077));
Q_AN02 U4748 ( .A0(n3959), .A1(GFidata[148]), .Z(n4076));
Q_AN02 U4749 ( .A0(n3959), .A1(GFidata[147]), .Z(n4075));
Q_AN02 U4750 ( .A0(n3959), .A1(GFidata[146]), .Z(n4074));
Q_AN02 U4751 ( .A0(n3959), .A1(GFidata[145]), .Z(n4073));
Q_AN02 U4752 ( .A0(n3959), .A1(GFidata[144]), .Z(n4072));
Q_AN02 U4753 ( .A0(n3959), .A1(GFidata[143]), .Z(n4071));
Q_AN02 U4754 ( .A0(n3959), .A1(GFidata[142]), .Z(n4070));
Q_AN02 U4755 ( .A0(n3959), .A1(GFidata[141]), .Z(n4069));
Q_AN02 U4756 ( .A0(n3959), .A1(GFidata[140]), .Z(n4068));
Q_AN02 U4757 ( .A0(n3959), .A1(GFidata[139]), .Z(n4067));
Q_AN02 U4758 ( .A0(n3959), .A1(GFidata[138]), .Z(n4066));
Q_AN02 U4759 ( .A0(n3959), .A1(GFidata[137]), .Z(n4065));
Q_AN02 U4760 ( .A0(n3959), .A1(GFidata[136]), .Z(n4064));
Q_AN02 U4761 ( .A0(n3959), .A1(GFidata[135]), .Z(n4063));
Q_AN02 U4762 ( .A0(n3959), .A1(GFidata[134]), .Z(n4062));
Q_AN02 U4763 ( .A0(n3959), .A1(GFidata[133]), .Z(n4061));
Q_AN02 U4764 ( .A0(n3959), .A1(GFidata[132]), .Z(n4060));
Q_AN02 U4765 ( .A0(n3959), .A1(GFidata[131]), .Z(n4059));
Q_AN02 U4766 ( .A0(n3959), .A1(GFidata[130]), .Z(n4058));
Q_AN02 U4767 ( .A0(n3959), .A1(GFidata[129]), .Z(n4057));
Q_AN02 U4768 ( .A0(n3959), .A1(GFidata[128]), .Z(n4056));
Q_AN02 U4769 ( .A0(n3959), .A1(GFidata[127]), .Z(n4055));
Q_AN02 U4770 ( .A0(n3959), .A1(GFidata[126]), .Z(n4054));
Q_AN02 U4771 ( .A0(n3959), .A1(GFidata[125]), .Z(n4053));
Q_AN02 U4772 ( .A0(n3959), .A1(GFidata[124]), .Z(n4052));
Q_AN02 U4773 ( .A0(n3959), .A1(GFidata[123]), .Z(n4051));
Q_AN02 U4774 ( .A0(n3959), .A1(GFidata[122]), .Z(n4050));
Q_AN02 U4775 ( .A0(n3959), .A1(GFidata[121]), .Z(n4049));
Q_AN02 U4776 ( .A0(n3959), .A1(GFidata[120]), .Z(n4048));
Q_AN02 U4777 ( .A0(n3959), .A1(GFidata[119]), .Z(n4047));
Q_AN02 U4778 ( .A0(n3959), .A1(GFidata[118]), .Z(n4046));
Q_AN02 U4779 ( .A0(n3959), .A1(GFidata[117]), .Z(n4045));
Q_AN02 U4780 ( .A0(n3959), .A1(GFidata[116]), .Z(n4044));
Q_AN02 U4781 ( .A0(n3959), .A1(GFidata[115]), .Z(n4043));
Q_AN02 U4782 ( .A0(n3959), .A1(GFidata[114]), .Z(n4042));
Q_AN02 U4783 ( .A0(n3959), .A1(GFidata[113]), .Z(n4041));
Q_AN02 U4784 ( .A0(n3959), .A1(GFidata[112]), .Z(n4040));
Q_AN02 U4785 ( .A0(n3959), .A1(GFidata[111]), .Z(n4039));
Q_AN02 U4786 ( .A0(n3959), .A1(GFidata[110]), .Z(n4038));
Q_AN02 U4787 ( .A0(n3959), .A1(GFidata[109]), .Z(n4037));
Q_AN02 U4788 ( .A0(n3959), .A1(GFidata[108]), .Z(n4036));
Q_AN02 U4789 ( .A0(n3959), .A1(GFidata[107]), .Z(n4035));
Q_AN02 U4790 ( .A0(n3959), .A1(GFidata[106]), .Z(n4034));
Q_AN02 U4791 ( .A0(n3959), .A1(GFidata[105]), .Z(n4033));
Q_AN02 U4792 ( .A0(n3959), .A1(GFidata[104]), .Z(n4032));
Q_AN02 U4793 ( .A0(n3959), .A1(GFidata[103]), .Z(n4031));
Q_AN02 U4794 ( .A0(n3959), .A1(GFidata[102]), .Z(n4030));
Q_AN02 U4795 ( .A0(n3959), .A1(GFidata[101]), .Z(n4029));
Q_AN02 U4796 ( .A0(n3959), .A1(GFidata[100]), .Z(n4028));
Q_AN02 U4797 ( .A0(n3959), .A1(GFidata[99]), .Z(n4027));
Q_AN02 U4798 ( .A0(n3959), .A1(GFidata[98]), .Z(n4026));
Q_AN02 U4799 ( .A0(n3959), .A1(GFidata[97]), .Z(n4025));
Q_AN02 U4800 ( .A0(n3959), .A1(GFidata[96]), .Z(n4024));
Q_AN02 U4801 ( .A0(n3959), .A1(GFidata[95]), .Z(n4023));
Q_AN02 U4802 ( .A0(n3959), .A1(GFidata[94]), .Z(n4022));
Q_AN02 U4803 ( .A0(n3959), .A1(GFidata[93]), .Z(n4021));
Q_AN02 U4804 ( .A0(n3959), .A1(GFidata[92]), .Z(n4020));
Q_AN02 U4805 ( .A0(n3959), .A1(GFidata[91]), .Z(n4019));
Q_AN02 U4806 ( .A0(n3959), .A1(GFidata[90]), .Z(n4018));
Q_AN02 U4807 ( .A0(n3959), .A1(GFidata[89]), .Z(n4017));
Q_AN02 U4808 ( .A0(n3959), .A1(GFidata[88]), .Z(n4016));
Q_AN02 U4809 ( .A0(n3959), .A1(GFidata[87]), .Z(n4015));
Q_AN02 U4810 ( .A0(n3959), .A1(GFidata[86]), .Z(n4014));
Q_AN02 U4811 ( .A0(n3959), .A1(GFidata[85]), .Z(n4013));
Q_AN02 U4812 ( .A0(n3959), .A1(GFidata[84]), .Z(n4012));
Q_AN02 U4813 ( .A0(n3959), .A1(GFidata[83]), .Z(n4011));
Q_AN02 U4814 ( .A0(n3959), .A1(GFidata[82]), .Z(n4010));
Q_AN02 U4815 ( .A0(n3959), .A1(GFidata[81]), .Z(n4009));
Q_AN02 U4816 ( .A0(n3959), .A1(GFidata[80]), .Z(n4008));
Q_AN02 U4817 ( .A0(n3959), .A1(GFidata[79]), .Z(n4007));
Q_AN02 U4818 ( .A0(n3959), .A1(GFidata[78]), .Z(n4006));
Q_AN02 U4819 ( .A0(n3959), .A1(GFidata[77]), .Z(n4005));
Q_AN02 U4820 ( .A0(n3959), .A1(GFidata[76]), .Z(n4004));
Q_AN02 U4821 ( .A0(n3959), .A1(GFidata[75]), .Z(n4003));
Q_AN02 U4822 ( .A0(n3959), .A1(GFidata[74]), .Z(n4002));
Q_AN02 U4823 ( .A0(n3959), .A1(GFidata[73]), .Z(n4001));
Q_AN02 U4824 ( .A0(n3959), .A1(GFidata[72]), .Z(n4000));
Q_AN02 U4825 ( .A0(n3959), .A1(GFidata[71]), .Z(n3999));
Q_AN02 U4826 ( .A0(n3959), .A1(GFidata[70]), .Z(n3998));
Q_AN02 U4827 ( .A0(n3959), .A1(GFidata[69]), .Z(n3997));
Q_AN02 U4828 ( .A0(n3959), .A1(GFidata[68]), .Z(n3996));
Q_AN02 U4829 ( .A0(n3959), .A1(GFidata[67]), .Z(n3995));
Q_AN02 U4830 ( .A0(n3959), .A1(GFidata[66]), .Z(n3994));
Q_AN02 U4831 ( .A0(n3959), .A1(GFidata[65]), .Z(n3993));
Q_AN02 U4832 ( .A0(n3959), .A1(GFidata[64]), .Z(n3992));
Q_AN02 U4833 ( .A0(n3959), .A1(GFidata[63]), .Z(n3991));
Q_AN02 U4834 ( .A0(n3959), .A1(GFidata[62]), .Z(n3990));
Q_AN02 U4835 ( .A0(n3959), .A1(GFidata[61]), .Z(n3989));
Q_AN02 U4836 ( .A0(n3959), .A1(GFidata[60]), .Z(n3988));
Q_AN02 U4837 ( .A0(n3959), .A1(GFidata[59]), .Z(n3987));
Q_AN02 U4838 ( .A0(n3959), .A1(GFidata[58]), .Z(n3986));
Q_AN02 U4839 ( .A0(n3959), .A1(GFidata[57]), .Z(n3985));
Q_AN02 U4840 ( .A0(n3959), .A1(GFidata[56]), .Z(n3984));
Q_AN02 U4841 ( .A0(n3959), .A1(GFidata[55]), .Z(n3983));
Q_AN02 U4842 ( .A0(n3959), .A1(GFidata[54]), .Z(n3982));
Q_AN02 U4843 ( .A0(n3959), .A1(GFidata[53]), .Z(n3981));
Q_AN02 U4844 ( .A0(n3959), .A1(GFidata[52]), .Z(n3980));
Q_AN02 U4845 ( .A0(n3959), .A1(GFidata[51]), .Z(n3979));
Q_AN02 U4846 ( .A0(n3959), .A1(GFidata[50]), .Z(n3978));
Q_AN02 U4847 ( .A0(n3959), .A1(GFidata[49]), .Z(n3977));
Q_AN02 U4848 ( .A0(n3959), .A1(GFidata[48]), .Z(n3976));
Q_AN02 U4849 ( .A0(n3959), .A1(GFidata[47]), .Z(n3975));
Q_AN02 U4850 ( .A0(n3959), .A1(GFidata[46]), .Z(n3974));
Q_AN02 U4851 ( .A0(n3959), .A1(GFidata[45]), .Z(n3973));
Q_AN02 U4852 ( .A0(n3959), .A1(GFidata[44]), .Z(n3972));
Q_AN02 U4853 ( .A0(n3959), .A1(GFidata[43]), .Z(n3971));
Q_AN02 U4854 ( .A0(n3959), .A1(GFidata[42]), .Z(n3970));
Q_AN02 U4855 ( .A0(n3959), .A1(GFidata[41]), .Z(n3969));
Q_AN02 U4856 ( .A0(n3959), .A1(GFidata[40]), .Z(n3968));
Q_AN02 U4857 ( .A0(n3959), .A1(GFidata[39]), .Z(n3967));
Q_AN02 U4858 ( .A0(n3959), .A1(GFidata[38]), .Z(n3966));
Q_AN02 U4859 ( .A0(n3959), .A1(GFidata[37]), .Z(n3965));
Q_AN02 U4860 ( .A0(n3959), .A1(GFidata[36]), .Z(n3964));
Q_AN02 U4861 ( .A0(n3959), .A1(GFidata[35]), .Z(n3963));
Q_AN02 U4862 ( .A0(n3959), .A1(GFidata[34]), .Z(n3962));
Q_AN02 U4863 ( .A0(n3959), .A1(GFidata[33]), .Z(n3961));
Q_AN02 U4864 ( .A0(n3959), .A1(GFidata[32]), .Z(n3960));
Q_INV U4865 ( .A(n5814), .Z(n3959));
Q_MX02 U4866 ( .S(n5814), .A0(GFidata[31]), .A1(timeStampPkt[63]), .Z(n3958));
Q_MX02 U4867 ( .S(n5814), .A0(GFidata[30]), .A1(timeStampPkt[62]), .Z(n3957));
Q_MX02 U4868 ( .S(n5814), .A0(GFidata[29]), .A1(timeStampPkt[61]), .Z(n3956));
Q_MX02 U4869 ( .S(n5814), .A0(GFidata[28]), .A1(timeStampPkt[60]), .Z(n3955));
Q_MX02 U4870 ( .S(n5814), .A0(GFidata[27]), .A1(timeStampPkt[59]), .Z(n3954));
Q_MX02 U4871 ( .S(n5814), .A0(GFidata[26]), .A1(timeStampPkt[58]), .Z(n3953));
Q_MX02 U4872 ( .S(n5814), .A0(GFidata[25]), .A1(timeStampPkt[57]), .Z(n3952));
Q_MX02 U4873 ( .S(n5814), .A0(GFidata[24]), .A1(timeStampPkt[56]), .Z(n3951));
Q_MX02 U4874 ( .S(n5814), .A0(GFidata[23]), .A1(timeStampPkt[55]), .Z(n3950));
Q_MX02 U4875 ( .S(n5814), .A0(GFidata[22]), .A1(timeStampPkt[54]), .Z(n3949));
Q_MX02 U4876 ( .S(n5814), .A0(GFidata[21]), .A1(timeStampPkt[53]), .Z(n3948));
Q_MX02 U4877 ( .S(n5814), .A0(GFidata[20]), .A1(timeStampPkt[52]), .Z(n3947));
Q_MX02 U4878 ( .S(n5814), .A0(GFidata[19]), .A1(timeStampPkt[51]), .Z(n3946));
Q_MX02 U4879 ( .S(n5814), .A0(GFidata[18]), .A1(timeStampPkt[50]), .Z(n3945));
Q_MX02 U4880 ( .S(n5814), .A0(GFidata[17]), .A1(timeStampPkt[49]), .Z(n3944));
Q_MX02 U4881 ( .S(n5814), .A0(GFidata[16]), .A1(timeStampPkt[48]), .Z(n3943));
Q_MX02 U4882 ( .S(n5814), .A0(GFidata[15]), .A1(timeStampPkt[47]), .Z(n3942));
Q_MX02 U4883 ( .S(n5814), .A0(GFidata[14]), .A1(timeStampPkt[46]), .Z(n3941));
Q_MX02 U4884 ( .S(n5814), .A0(GFidata[13]), .A1(timeStampPkt[45]), .Z(n3940));
Q_MX02 U4885 ( .S(n5814), .A0(GFidata[12]), .A1(timeStampPkt[44]), .Z(n3939));
Q_MX02 U4886 ( .S(n5814), .A0(GFidata[11]), .A1(timeStampPkt[43]), .Z(n3938));
Q_MX02 U4887 ( .S(n5814), .A0(GFidata[10]), .A1(timeStampPkt[42]), .Z(n3937));
Q_MX02 U4888 ( .S(n5814), .A0(GFidata[9]), .A1(timeStampPkt[41]), .Z(n3936));
Q_MX02 U4889 ( .S(n5814), .A0(GFidata[8]), .A1(timeStampPkt[40]), .Z(n3935));
Q_MX02 U4890 ( .S(n5814), .A0(GFidata[7]), .A1(timeStampPkt[39]), .Z(n3934));
Q_MX02 U4891 ( .S(n5814), .A0(GFidata[6]), .A1(timeStampPkt[38]), .Z(n3933));
Q_MX02 U4892 ( .S(n5814), .A0(GFidata[5]), .A1(timeStampPkt[37]), .Z(n3932));
Q_MX02 U4893 ( .S(n5814), .A0(GFidata[4]), .A1(timeStampPkt[36]), .Z(n3931));
Q_MX02 U4894 ( .S(n5814), .A0(GFidata[3]), .A1(timeStampPkt[35]), .Z(n3930));
Q_MX02 U4895 ( .S(n5814), .A0(GFidata[2]), .A1(timeStampPkt[34]), .Z(n3929));
Q_MX02 U4896 ( .S(n5814), .A0(GFidata[1]), .A1(timeStampPkt[33]), .Z(n3928));
Q_MX02 U4897 ( .S(n5814), .A0(GFidata[0]), .A1(timeStampPkt[32]), .Z(n3927));
Q_MX02 U4898 ( .S(n5814), .A0(GFlen[10]), .A1(timeStampPkt[30]), .Z(n3925));
Q_MX02 U4899 ( .S(n5814), .A0(GFlen[9]), .A1(timeStampPkt[29]), .Z(n3924));
Q_MX02 U4900 ( .S(n5814), .A0(GFlen[8]), .A1(timeStampPkt[28]), .Z(n3923));
Q_MX02 U4901 ( .S(n5814), .A0(GFlen[7]), .A1(timeStampPkt[27]), .Z(n3922));
Q_MX02 U4902 ( .S(n5814), .A0(GFlen[6]), .A1(timeStampPkt[26]), .Z(n3921));
Q_MX02 U4903 ( .S(n5814), .A0(GFlen[5]), .A1(timeStampPkt[25]), .Z(n3920));
Q_MX02 U4904 ( .S(n5814), .A0(GFlen[4]), .A1(timeStampPkt[24]), .Z(n3919));
Q_MX02 U4905 ( .S(n5814), .A0(GFlen[3]), .A1(timeStampPkt[23]), .Z(n3918));
Q_MX02 U4906 ( .S(n5814), .A0(GFlen[2]), .A1(timeStampPkt[22]), .Z(n3917));
Q_MX02 U4907 ( .S(n5814), .A0(GFlen[1]), .A1(timeStampPkt[21]), .Z(n3916));
Q_MX02 U4908 ( .S(n5814), .A0(GFlen[0]), .A1(timeStampPkt[20]), .Z(n3915));
Q_MX02 U4909 ( .S(n5814), .A0(GFcbid[19]), .A1(timeStampPkt[19]), .Z(n3914));
Q_MX02 U4910 ( .S(n5814), .A0(GFcbid[18]), .A1(timeStampPkt[18]), .Z(n3913));
Q_MX02 U4911 ( .S(n5814), .A0(GFcbid[17]), .A1(timeStampPkt[17]), .Z(n3912));
Q_MX02 U4912 ( .S(n5814), .A0(GFcbid[16]), .A1(timeStampPkt[16]), .Z(n3911));
Q_MX02 U4913 ( .S(n5814), .A0(GFcbid[15]), .A1(timeStampPkt[15]), .Z(n3910));
Q_MX02 U4914 ( .S(n5814), .A0(GFcbid[14]), .A1(timeStampPkt[14]), .Z(n3909));
Q_MX02 U4915 ( .S(n5814), .A0(GFcbid[13]), .A1(timeStampPkt[13]), .Z(n3908));
Q_MX02 U4916 ( .S(n5814), .A0(GFcbid[12]), .A1(timeStampPkt[12]), .Z(n3907));
Q_MX02 U4917 ( .S(n5814), .A0(GFcbid[11]), .A1(timeStampPkt[11]), .Z(n3906));
Q_MX02 U4918 ( .S(n5814), .A0(GFcbid[10]), .A1(timeStampPkt[10]), .Z(n3905));
Q_MX02 U4919 ( .S(n5814), .A0(GFcbid[9]), .A1(timeStampPkt[9]), .Z(n3904));
Q_MX02 U4920 ( .S(n5814), .A0(GFcbid[8]), .A1(timeStampPkt[8]), .Z(n3903));
Q_MX02 U4921 ( .S(n5814), .A0(GFcbid[7]), .A1(timeStampPkt[7]), .Z(n3902));
Q_MX02 U4922 ( .S(n5814), .A0(GFcbid[6]), .A1(timeStampPkt[6]), .Z(n3901));
Q_MX02 U4923 ( .S(n5814), .A0(GFcbid[5]), .A1(timeStampPkt[5]), .Z(n3900));
Q_MX02 U4924 ( .S(n5814), .A0(GFcbid[4]), .A1(timeStampPkt[4]), .Z(n3899));
Q_MX02 U4925 ( .S(n5814), .A0(GFcbid[3]), .A1(timeStampPkt[3]), .Z(n3898));
Q_MX02 U4926 ( .S(n5814), .A0(GFcbid[2]), .A1(timeStampPkt[2]), .Z(n3897));
Q_MX02 U4927 ( .S(n5814), .A0(GFcbid[1]), .A1(timeStampPkt[1]), .Z(n3896));
Q_MX02 U4928 ( .S(n5814), .A0(GFcbid[0]), .A1(timeStampPkt[0]), .Z(n3895));
Q_AD01HF U4929 ( .A0(n3891), .B0(n3860), .S(n3892), .CO(n3893));
Q_AD01HF U4930 ( .A0(n3889), .B0(n3858), .S(n3890), .CO(n3891));
Q_AD01HF U4931 ( .A0(n3887), .B0(n3856), .S(n3888), .CO(n3889));
Q_AD01HF U4932 ( .A0(n3885), .B0(n3854), .S(n3886), .CO(n3887));
Q_AD01HF U4933 ( .A0(n3883), .B0(n3852), .S(n3884), .CO(n3885));
Q_AD01HF U4934 ( .A0(n3850), .B0(n3881), .S(n3882), .CO(n3883));
Q_AD02 U4935 ( .CI(n3878), .A0(GFlen[10]), .A1(GFlen[11]), .B0(n3846), .B1(n3848), .S0(n3879), .S1(n3880), .CO(n3881));
Q_AD02 U4936 ( .CI(n3875), .A0(GFlen[8]), .A1(GFlen[9]), .B0(n3842), .B1(n3844), .S0(n3876), .S1(n3877), .CO(n3878));
Q_AD02 U4937 ( .CI(n3872), .A0(GFlen[6]), .A1(GFlen[7]), .B0(n3838), .B1(n3840), .S0(n3873), .S1(n3874), .CO(n3875));
Q_AD02 U4938 ( .CI(n3869), .A0(GFlen[4]), .A1(GFlen[5]), .B0(n3834), .B1(n3836), .S0(n3870), .S1(n3871), .CO(n3872));
Q_AD02 U4939 ( .CI(n3866), .A0(GFlen[2]), .A1(GFlen[3]), .B0(n3830), .B1(n3832), .S0(n3867), .S1(n3868), .CO(n3869));
Q_AD01 U4940 ( .CI(n3828), .A0(GFlen[1]), .B0(n3864), .S(n3865), .CO(n3866));
Q_OR02 U4941 ( .A0(GFlen[0]), .A1(n3826), .Z(n3864));
Q_XNR2 U4942 ( .A0(GFlen[0]), .A1(n3826), .Z(n3863));
Q_MX02 U4943 ( .S(n5813), .A0(n3861), .A1(n3824), .Z(n3862));
Q_AN02 U4944 ( .A0(n5812), .A1(wLen[18]), .Z(n3861));
Q_MX02 U4945 ( .S(n5813), .A0(n3859), .A1(n3822), .Z(n3860));
Q_AN02 U4946 ( .A0(n5812), .A1(wLen[17]), .Z(n3859));
Q_MX02 U4947 ( .S(n5813), .A0(n3857), .A1(n3821), .Z(n3858));
Q_AN02 U4948 ( .A0(n5812), .A1(wLen[16]), .Z(n3857));
Q_MX02 U4949 ( .S(n5813), .A0(n3855), .A1(n3819), .Z(n3856));
Q_AN02 U4950 ( .A0(n5812), .A1(wLen[15]), .Z(n3855));
Q_MX02 U4951 ( .S(n5813), .A0(n3853), .A1(n3818), .Z(n3854));
Q_AN02 U4952 ( .A0(n5812), .A1(wLen[14]), .Z(n3853));
Q_MX02 U4953 ( .S(n5813), .A0(n3851), .A1(n3816), .Z(n3852));
Q_AN02 U4954 ( .A0(n5812), .A1(wLen[13]), .Z(n3851));
Q_MX02 U4955 ( .S(n5813), .A0(n3849), .A1(n3815), .Z(n3850));
Q_AN02 U4956 ( .A0(n5812), .A1(wLen[12]), .Z(n3849));
Q_MX02 U4957 ( .S(n5813), .A0(n3847), .A1(n3813), .Z(n3848));
Q_AN02 U4958 ( .A0(n5812), .A1(wLen[11]), .Z(n3847));
Q_MX02 U4959 ( .S(n5813), .A0(n3845), .A1(n3812), .Z(n3846));
Q_AN02 U4960 ( .A0(n5812), .A1(wLen[10]), .Z(n3845));
Q_MX02 U4961 ( .S(n5813), .A0(n3843), .A1(n3810), .Z(n3844));
Q_AN02 U4962 ( .A0(n5812), .A1(wLen[9]), .Z(n3843));
Q_MX02 U4963 ( .S(n5813), .A0(n3841), .A1(n3809), .Z(n3842));
Q_AN02 U4964 ( .A0(n5812), .A1(wLen[8]), .Z(n3841));
Q_MX02 U4965 ( .S(n5813), .A0(n3839), .A1(n3807), .Z(n3840));
Q_AN02 U4966 ( .A0(n5812), .A1(wLen[7]), .Z(n3839));
Q_MX02 U4967 ( .S(n5813), .A0(n3837), .A1(n3806), .Z(n3838));
Q_AN02 U4968 ( .A0(n5812), .A1(wLen[6]), .Z(n3837));
Q_MX02 U4969 ( .S(n5813), .A0(n3835), .A1(n3804), .Z(n3836));
Q_AN02 U4970 ( .A0(n5812), .A1(wLen[5]), .Z(n3835));
Q_MX02 U4971 ( .S(n5813), .A0(n3833), .A1(n3803), .Z(n3834));
Q_AN02 U4972 ( .A0(n5812), .A1(wLen[4]), .Z(n3833));
Q_MX02 U4973 ( .S(n5813), .A0(n3831), .A1(n3801), .Z(n3832));
Q_AN02 U4974 ( .A0(n5812), .A1(wLen[3]), .Z(n3831));
Q_MX02 U4975 ( .S(n5813), .A0(n3829), .A1(n3800), .Z(n3830));
Q_AN02 U4976 ( .A0(n5812), .A1(wLen[2]), .Z(n3829));
Q_MX02 U4977 ( .S(n5813), .A0(n3827), .A1(n3798), .Z(n3828));
Q_AN02 U4978 ( .A0(n5812), .A1(wLen[1]), .Z(n3827));
Q_MX02 U4979 ( .S(n5813), .A0(n3825), .A1(n3796), .Z(n3826));
Q_AN02 U4980 ( .A0(n5812), .A1(wLen[0]), .Z(n3825));
Q_XOR2 U4981 ( .A0(n3706), .A1(n3823), .Z(n3824));
Q_AD02 U4982 ( .CI(n3820), .A0(wLen[16]), .A1(wLen[17]), .B0(n3794), .B1(n3795), .S0(n3821), .S1(n3822), .CO(n3823));
Q_AD02 U4983 ( .CI(n3817), .A0(wLen[14]), .A1(wLen[15]), .B0(n3792), .B1(n3793), .S0(n3818), .S1(n3819), .CO(n3820));
Q_AD02 U4984 ( .CI(n3814), .A0(wLen[12]), .A1(wLen[13]), .B0(n3790), .B1(n3791), .S0(n3815), .S1(n3816), .CO(n3817));
Q_AD02 U4985 ( .CI(n3811), .A0(wLen[10]), .A1(wLen[11]), .B0(n3788), .B1(n3789), .S0(n3812), .S1(n3813), .CO(n3814));
Q_AD02 U4986 ( .CI(n3808), .A0(wLen[8]), .A1(wLen[9]), .B0(n3786), .B1(n3787), .S0(n3809), .S1(n3810), .CO(n3811));
Q_AD02 U4987 ( .CI(n3805), .A0(wLen[6]), .A1(wLen[7]), .B0(n3784), .B1(n3785), .S0(n3806), .S1(n3807), .CO(n3808));
Q_AD02 U4988 ( .CI(n3802), .A0(wLen[4]), .A1(wLen[5]), .B0(n3782), .B1(n3783), .S0(n3803), .S1(n3804), .CO(n3805));
Q_AD02 U4989 ( .CI(n3799), .A0(wLen[2]), .A1(wLen[3]), .B0(n3780), .B1(n3781), .S0(n3800), .S1(n3801), .CO(n3802));
Q_AD01 U4990 ( .CI(n3797), .A0(wLen[1]), .B0(n3779), .S(n3798), .CO(n3799));
Q_OR02 U4991 ( .A0(wLen[0]), .A1(n3778), .Z(n3797));
Q_XNR2 U4992 ( .A0(wLen[0]), .A1(n3778), .Z(n3796));
Q_ND02 U4993 ( .A0(n5820), .A1(rLen[17]), .Z(n3795));
Q_ND02 U4994 ( .A0(n5820), .A1(rLen[16]), .Z(n3794));
Q_ND02 U4995 ( .A0(n5820), .A1(rLen[15]), .Z(n3793));
Q_ND02 U4996 ( .A0(n5820), .A1(rLen[14]), .Z(n3792));
Q_ND02 U4997 ( .A0(n5820), .A1(rLen[13]), .Z(n3791));
Q_ND02 U4998 ( .A0(n5820), .A1(rLen[12]), .Z(n3790));
Q_ND02 U4999 ( .A0(n5820), .A1(rLen[11]), .Z(n3789));
Q_ND02 U5000 ( .A0(n5820), .A1(rLen[10]), .Z(n3788));
Q_ND02 U5001 ( .A0(n5820), .A1(rLen[9]), .Z(n3787));
Q_ND02 U5002 ( .A0(n5820), .A1(rLen[8]), .Z(n3786));
Q_ND02 U5003 ( .A0(n5820), .A1(rLen[7]), .Z(n3785));
Q_ND02 U5004 ( .A0(n5820), .A1(rLen[6]), .Z(n3784));
Q_ND02 U5005 ( .A0(n5820), .A1(rLen[5]), .Z(n3783));
Q_ND02 U5006 ( .A0(n5820), .A1(rLen[4]), .Z(n3782));
Q_ND02 U5007 ( .A0(n5820), .A1(rLen[3]), .Z(n3781));
Q_ND02 U5008 ( .A0(n5820), .A1(rLen[2]), .Z(n3780));
Q_ND02 U5009 ( .A0(n5820), .A1(rLen[1]), .Z(n3779));
Q_ND02 U5010 ( .A0(n5820), .A1(rLen[0]), .Z(n3778));
Q_INV U5011 ( .A(n3777), .Z(n5820));
Q_AO21 U5012 ( .A0(n3776), .A1(n3769), .B0(n3775), .Z(n3777));
Q_OR03 U5013 ( .A0(n3716), .A1(n3774), .A2(n3773), .Z(n3775));
Q_AO21 U5014 ( .A0(n3770), .A1(n3745), .B0(n3772), .Z(n3773));
Q_OR03 U5015 ( .A0(n3761), .A1(n3768), .A2(n3767), .Z(n3769));
Q_AN03 U5016 ( .A0(n3762), .A1(n3764), .A2(n3766), .Z(n3767));
Q_AN02 U5017 ( .A0(rLen[0]), .A1(n3765), .Z(n3766));
Q_INV U5018 ( .A(wLen[0]), .Z(n3765));
Q_OR02 U5019 ( .A0(rLen[1]), .A1(n3763), .Z(n3764));
Q_AN03 U5020 ( .A0(rLen[1]), .A1(n3763), .A2(n3762), .Z(n3768));
Q_INV U5021 ( .A(wLen[1]), .Z(n3763));
Q_OR02 U5022 ( .A0(rLen[2]), .A1(n3760), .Z(n3762));
Q_AN02 U5023 ( .A0(rLen[2]), .A1(n3760), .Z(n3761));
Q_INV U5024 ( .A(wLen[2]), .Z(n3760));
Q_AN03 U5025 ( .A0(n3756), .A1(n3754), .A2(n3771), .Z(n3776));
Q_OA21 U5026 ( .A0(n3759), .A1(n3758), .B0(n3771), .Z(n3772));
Q_AO21 U5027 ( .A0(n3748), .A1(n3750), .B0(n3747), .Z(n3759));
Q_AO21 U5028 ( .A0(n3755), .A1(n3752), .B0(n3757), .Z(n3758));
Q_OR02 U5029 ( .A0(rLen[3]), .A1(n3753), .Z(n3754));
Q_AN03 U5030 ( .A0(rLen[3]), .A1(n3753), .A2(n3756), .Z(n3757));
Q_INV U5031 ( .A(wLen[3]), .Z(n3753));
Q_OA21 U5032 ( .A0(rLen[4]), .A1(n3751), .B0(n3755), .Z(n3756));
Q_AN02 U5033 ( .A0(rLen[4]), .A1(n3751), .Z(n3752));
Q_INV U5034 ( .A(wLen[4]), .Z(n3751));
Q_OA21 U5035 ( .A0(rLen[5]), .A1(n3749), .B0(n3748), .Z(n3755));
Q_AN02 U5036 ( .A0(rLen[5]), .A1(n3749), .Z(n3750));
Q_INV U5037 ( .A(wLen[5]), .Z(n3749));
Q_OR02 U5038 ( .A0(rLen[6]), .A1(n3746), .Z(n3748));
Q_AN02 U5039 ( .A0(rLen[6]), .A1(n3746), .Z(n3747));
Q_INV U5040 ( .A(wLen[6]), .Z(n3746));
Q_AN03 U5041 ( .A0(n3741), .A1(n3739), .A2(n3770), .Z(n3771));
Q_OR03 U5042 ( .A0(n3733), .A1(n3744), .A2(n3743), .Z(n3745));
Q_AO21 U5043 ( .A0(n3740), .A1(n3737), .B0(n3742), .Z(n3743));
Q_OR02 U5044 ( .A0(rLen[7]), .A1(n3738), .Z(n3739));
Q_AN03 U5045 ( .A0(rLen[7]), .A1(n3738), .A2(n3741), .Z(n3742));
Q_INV U5046 ( .A(wLen[7]), .Z(n3738));
Q_OA21 U5047 ( .A0(rLen[8]), .A1(n3736), .B0(n3740), .Z(n3741));
Q_AN02 U5048 ( .A0(rLen[8]), .A1(n3736), .Z(n3737));
Q_INV U5049 ( .A(wLen[8]), .Z(n3736));
Q_OA21 U5050 ( .A0(rLen[9]), .A1(n3735), .B0(n3734), .Z(n3740));
Q_AN03 U5051 ( .A0(rLen[9]), .A1(n3735), .A2(n3734), .Z(n3744));
Q_INV U5052 ( .A(wLen[9]), .Z(n3735));
Q_OR02 U5053 ( .A0(rLen[10]), .A1(n3732), .Z(n3734));
Q_AN02 U5054 ( .A0(rLen[10]), .A1(n3732), .Z(n3733));
Q_INV U5055 ( .A(wLen[10]), .Z(n3732));
Q_AN03 U5056 ( .A0(n3728), .A1(n3726), .A2(n3717), .Z(n3770));
Q_OA21 U5057 ( .A0(n3731), .A1(n3730), .B0(n3717), .Z(n3774));
Q_AO21 U5058 ( .A0(n3720), .A1(n3722), .B0(n3719), .Z(n3731));
Q_AO21 U5059 ( .A0(n3727), .A1(n3724), .B0(n3729), .Z(n3730));
Q_OR02 U5060 ( .A0(rLen[11]), .A1(n3725), .Z(n3726));
Q_AN03 U5061 ( .A0(rLen[11]), .A1(n3725), .A2(n3728), .Z(n3729));
Q_INV U5062 ( .A(wLen[11]), .Z(n3725));
Q_OA21 U5063 ( .A0(rLen[12]), .A1(n3723), .B0(n3727), .Z(n3728));
Q_AN02 U5064 ( .A0(rLen[12]), .A1(n3723), .Z(n3724));
Q_INV U5065 ( .A(wLen[12]), .Z(n3723));
Q_OA21 U5066 ( .A0(rLen[13]), .A1(n3721), .B0(n3720), .Z(n3727));
Q_AN02 U5067 ( .A0(rLen[13]), .A1(n3721), .Z(n3722));
Q_INV U5068 ( .A(wLen[13]), .Z(n3721));
Q_OR02 U5069 ( .A0(rLen[14]), .A1(n3718), .Z(n3720));
Q_AN02 U5070 ( .A0(rLen[14]), .A1(n3718), .Z(n3719));
Q_INV U5071 ( .A(wLen[14]), .Z(n3718));
Q_AO21 U5072 ( .A0(n3706), .A1(n3708), .B0(n3715), .Z(n3716));
Q_AO21 U5073 ( .A0(n3712), .A1(n3710), .B0(n3714), .Z(n3715));
Q_OA21 U5074 ( .A0(rLen[15]), .A1(n3711), .B0(n3713), .Z(n3717));
Q_AN03 U5075 ( .A0(rLen[15]), .A1(n3711), .A2(n3713), .Z(n3714));
Q_INV U5076 ( .A(wLen[15]), .Z(n3711));
Q_OA21 U5077 ( .A0(rLen[16]), .A1(n3709), .B0(n3712), .Z(n3713));
Q_AN02 U5078 ( .A0(rLen[16]), .A1(n3709), .Z(n3710));
Q_INV U5079 ( .A(wLen[16]), .Z(n3709));
Q_OA21 U5080 ( .A0(rLen[17]), .A1(n3707), .B0(n3706), .Z(n3712));
Q_AN02 U5081 ( .A0(rLen[17]), .A1(n3707), .Z(n3708));
Q_INV U5082 ( .A(wLen[17]), .Z(n3707));
Q_INV U5083 ( .A(wLen[18]), .Z(n3706));
Q_OR03 U5084 ( .A0(n3701), .A1(n3702), .A2(n3705), .Z(n5823));
Q_OA21 U5085 ( .A0(n3704), .A1(n3703), .B0(GFlen[4]), .Z(n3705));
Q_OR02 U5086 ( .A0(GFlen[3]), .A1(GFlen[2]), .Z(n3704));
Q_OR02 U5087 ( .A0(GFlen[1]), .A1(GFlen[0]), .Z(n3703));
Q_OR03 U5088 ( .A0(GFlen[7]), .A1(GFlen[6]), .A2(GFlen[5]), .Z(n3702));
Q_OR03 U5089 ( .A0(GFlen[11]), .A1(GFlen[10]), .A2(n3700), .Z(n3701));
Q_OR02 U5090 ( .A0(GFlen[9]), .A1(GFlen[8]), .Z(n3700));
Q_INV U5091 ( .A(n3699), .Z(n5816));
Q_AN02 U5092 ( .A0(n3697), .A1(n3698), .Z(n3699));
Q_AN03 U5093 ( .A0(n3694), .A1(n3695), .A2(n3696), .Z(n3698));
Q_AN03 U5094 ( .A0(n3691), .A1(n3692), .A2(n3693), .Z(n3697));
Q_AN03 U5095 ( .A0(GFcbid[1]), .A1(GFcbid[0]), .A2(n3690), .Z(n3696));
Q_AN03 U5096 ( .A0(GFcbid[4]), .A1(GFcbid[3]), .A2(GFcbid[2]), .Z(n3695));
Q_AN03 U5097 ( .A0(GFcbid[7]), .A1(GFcbid[6]), .A2(GFcbid[5]), .Z(n3694));
Q_AN03 U5098 ( .A0(GFcbid[10]), .A1(GFcbid[9]), .A2(GFcbid[8]), .Z(n3693));
Q_AN03 U5099 ( .A0(GFcbid[13]), .A1(GFcbid[12]), .A2(GFcbid[11]), .Z(n3692));
Q_AN03 U5100 ( .A0(GFcbid[16]), .A1(GFcbid[15]), .A2(GFcbid[14]), .Z(n3691));
Q_AN03 U5101 ( .A0(GFcbid[19]), .A1(GFcbid[18]), .A2(GFcbid[17]), .Z(n3690));
Q_AN03 U5102 ( .A0(n3684), .A1(n3685), .A2(n3689), .Z(n5822));
Q_ND02 U5103 ( .A0(n3697), .A1(n3688), .Z(n3689));
Q_AN03 U5104 ( .A0(n3694), .A1(n3695), .A2(n3687), .Z(n3688));
Q_AN03 U5105 ( .A0(n3686), .A1(GFcbid[0]), .A2(n3690), .Z(n3687));
Q_INV U5106 ( .A(GFcbid[1]), .Z(n3686));
Q_INV U5107 ( .A(xc_top.GFLock2), .Z(n3685));
Q_OR02 U5108 ( .A0(reqD), .A1(GFtsAdd), .Z(n3684));
Q_XNR2 U5109 ( .A0(rSync), .A1(wSync), .Z(n3683));
Q_AN02 U5110 ( .A0(n3697), .A1(n3682), .Z(n5814));
Q_AN03 U5111 ( .A0(n3694), .A1(n3695), .A2(n3681), .Z(n3682));
Q_AN03 U5112 ( .A0(GFcbid[1]), .A1(n3680), .A2(n3690), .Z(n3681));
Q_INV U5113 ( .A(GFcbid[0]), .Z(n3680));
Q_AN03 U5114 ( .A0(xc_top.anyStop), .A1(LBempty), .A2(n6717), .Z(n5821));
Q_AN02 U5115 ( .A0(n6720), .A1(hasMultiLevelGFIFO), .Z(n3679));
Q_NR02 U5116 ( .A0(xc_top.GFReset), .A1(hasMultiLevelGFIFO), .Z(n3678));
Q_FDP0UA U5117 ( .D(n3675), .QTFCLK( ), .Q(GFfullD));
Q_FDP0UA U5118 ( .D(n3677), .QTFCLK( ), .Q(reqD));
Q_MX02 U5119 ( .S(n3679), .A0(n3676), .A1(n3673), .Z(n3677));
Q_AN02 U5120 ( .A0(n6720), .A1(GFfull), .Z(n3675));
Q_AN03 U5121 ( .A0(GFreq), .A1(n3674), .A2(n3678), .Z(n3676));
Q_INV U5122 ( .A(GFfull), .Z(n3674));
Q_AN02 U5123 ( .A0(GFreq), .A1(n3672), .Z(n3673));
Q_INV U5124 ( .A(GFfullD), .Z(n3672));
Q_FDP0UA U5125 ( .D(n3671), .QTFCLK( ), .Q(ackClk));
Q_INV U5126 ( .A(n3670), .Z(n3671));
Q_AN02 U5127 ( .A0(n3668), .A1(n3669), .Z(n3670));
Q_AN03 U5128 ( .A0(n3660), .A1(n3659), .A2(n3667), .Z(n3669));
Q_AN03 U5129 ( .A0(n3663), .A1(n3662), .A2(n3661), .Z(n3668));
Q_AN03 U5130 ( .A0(n3666), .A1(n3665), .A2(n3664), .Z(n3667));
Q_XNR2 U5131 ( .A0(ackIdNew[7]), .A1(ackId[7]), .Z(n3666));
Q_XNR2 U5132 ( .A0(ackIdNew[6]), .A1(ackId[6]), .Z(n3665));
Q_XNR2 U5133 ( .A0(ackIdNew[5]), .A1(ackId[5]), .Z(n3664));
Q_XNR2 U5134 ( .A0(ackIdNew[4]), .A1(ackId[4]), .Z(n3663));
Q_XNR2 U5135 ( .A0(ackIdNew[3]), .A1(ackId[3]), .Z(n3662));
Q_XNR2 U5136 ( .A0(ackIdNew[2]), .A1(ackId[2]), .Z(n3661));
Q_XNR2 U5137 ( .A0(ackIdNew[1]), .A1(ackId[1]), .Z(n3660));
Q_XNR2 U5138 ( .A0(ackIdNew[0]), .A1(ackId[0]), .Z(n3659));
Q_MX02 U5139 ( .S(n3670), .A0(ackIdNew[0]), .A1(ackId[0]), .Z(n3658));
Q_FDP0UA U5140 ( .D(n3658), .QTFCLK( ), .Q(ackId[0]));
Q_MX02 U5141 ( .S(n3670), .A0(ackIdNew[1]), .A1(ackId[1]), .Z(n3657));
Q_FDP0UA U5142 ( .D(n3657), .QTFCLK( ), .Q(ackId[1]));
Q_MX02 U5143 ( .S(n3670), .A0(ackIdNew[2]), .A1(ackId[2]), .Z(n3656));
Q_FDP0UA U5144 ( .D(n3656), .QTFCLK( ), .Q(ackId[2]));
Q_MX02 U5145 ( .S(n3670), .A0(ackIdNew[3]), .A1(ackId[3]), .Z(n3655));
Q_FDP0UA U5146 ( .D(n3655), .QTFCLK( ), .Q(ackId[3]));
Q_MX02 U5147 ( .S(n3670), .A0(ackIdNew[4]), .A1(ackId[4]), .Z(n3654));
Q_FDP0UA U5148 ( .D(n3654), .QTFCLK( ), .Q(ackId[4]));
Q_MX02 U5149 ( .S(n3670), .A0(ackIdNew[5]), .A1(ackId[5]), .Z(n3653));
Q_FDP0UA U5150 ( .D(n3653), .QTFCLK( ), .Q(ackId[5]));
Q_MX02 U5151 ( .S(n3670), .A0(ackIdNew[6]), .A1(ackId[6]), .Z(n3652));
Q_FDP0UA U5152 ( .D(n3652), .QTFCLK( ), .Q(ackId[6]));
Q_MX02 U5153 ( .S(n3670), .A0(ackIdNew[7]), .A1(ackId[7]), .Z(n3651));
Q_FDP0UA U5154 ( .D(n3651), .QTFCLK( ), .Q(ackId[7]));
Q_FDP0UA U5155 ( .D(wrtCnt[63]), .QTFCLK( ), .Q(wrtCntD[63]));
Q_FDP0UA U5156 ( .D(wrtCnt[62]), .QTFCLK( ), .Q(wrtCntD[62]));
Q_FDP0UA U5157 ( .D(wrtCnt[61]), .QTFCLK( ), .Q(wrtCntD[61]));
Q_FDP0UA U5158 ( .D(wrtCnt[60]), .QTFCLK( ), .Q(wrtCntD[60]));
Q_FDP0UA U5159 ( .D(wrtCnt[59]), .QTFCLK( ), .Q(wrtCntD[59]));
Q_FDP0UA U5160 ( .D(wrtCnt[58]), .QTFCLK( ), .Q(wrtCntD[58]));
Q_FDP0UA U5161 ( .D(wrtCnt[57]), .QTFCLK( ), .Q(wrtCntD[57]));
Q_FDP0UA U5162 ( .D(wrtCnt[56]), .QTFCLK( ), .Q(wrtCntD[56]));
Q_FDP0UA U5163 ( .D(wrtCnt[55]), .QTFCLK( ), .Q(wrtCntD[55]));
Q_FDP0UA U5164 ( .D(wrtCnt[54]), .QTFCLK( ), .Q(wrtCntD[54]));
Q_FDP0UA U5165 ( .D(wrtCnt[53]), .QTFCLK( ), .Q(wrtCntD[53]));
Q_FDP0UA U5166 ( .D(wrtCnt[52]), .QTFCLK( ), .Q(wrtCntD[52]));
Q_FDP0UA U5167 ( .D(wrtCnt[51]), .QTFCLK( ), .Q(wrtCntD[51]));
Q_FDP0UA U5168 ( .D(wrtCnt[50]), .QTFCLK( ), .Q(wrtCntD[50]));
Q_FDP0UA U5169 ( .D(wrtCnt[49]), .QTFCLK( ), .Q(wrtCntD[49]));
Q_FDP0UA U5170 ( .D(wrtCnt[48]), .QTFCLK( ), .Q(wrtCntD[48]));
Q_FDP0UA U5171 ( .D(wrtCnt[47]), .QTFCLK( ), .Q(wrtCntD[47]));
Q_FDP0UA U5172 ( .D(wrtCnt[46]), .QTFCLK( ), .Q(wrtCntD[46]));
Q_FDP0UA U5173 ( .D(wrtCnt[45]), .QTFCLK( ), .Q(wrtCntD[45]));
Q_FDP0UA U5174 ( .D(wrtCnt[44]), .QTFCLK( ), .Q(wrtCntD[44]));
Q_FDP0UA U5175 ( .D(wrtCnt[43]), .QTFCLK( ), .Q(wrtCntD[43]));
Q_FDP0UA U5176 ( .D(wrtCnt[42]), .QTFCLK( ), .Q(wrtCntD[42]));
Q_FDP0UA U5177 ( .D(wrtCnt[41]), .QTFCLK( ), .Q(wrtCntD[41]));
Q_FDP0UA U5178 ( .D(wrtCnt[40]), .QTFCLK( ), .Q(wrtCntD[40]));
Q_FDP0UA U5179 ( .D(wrtCnt[39]), .QTFCLK( ), .Q(wrtCntD[39]));
Q_FDP0UA U5180 ( .D(wrtCnt[38]), .QTFCLK( ), .Q(wrtCntD[38]));
Q_FDP0UA U5181 ( .D(wrtCnt[37]), .QTFCLK( ), .Q(wrtCntD[37]));
Q_FDP0UA U5182 ( .D(wrtCnt[36]), .QTFCLK( ), .Q(wrtCntD[36]));
Q_FDP0UA U5183 ( .D(wrtCnt[35]), .QTFCLK( ), .Q(wrtCntD[35]));
Q_FDP0UA U5184 ( .D(wrtCnt[34]), .QTFCLK( ), .Q(wrtCntD[34]));
Q_FDP0UA U5185 ( .D(wrtCnt[33]), .QTFCLK( ), .Q(wrtCntD[33]));
Q_FDP0UA U5186 ( .D(wrtCnt[32]), .QTFCLK( ), .Q(wrtCntD[32]));
Q_FDP0UA U5187 ( .D(wrtCnt[31]), .QTFCLK( ), .Q(wrtCntD[31]));
Q_FDP0UA U5188 ( .D(wrtCnt[30]), .QTFCLK( ), .Q(wrtCntD[30]));
Q_FDP0UA U5189 ( .D(wrtCnt[29]), .QTFCLK( ), .Q(wrtCntD[29]));
Q_FDP0UA U5190 ( .D(wrtCnt[28]), .QTFCLK( ), .Q(wrtCntD[28]));
Q_FDP0UA U5191 ( .D(wrtCnt[27]), .QTFCLK( ), .Q(wrtCntD[27]));
Q_FDP0UA U5192 ( .D(wrtCnt[26]), .QTFCLK( ), .Q(wrtCntD[26]));
Q_FDP0UA U5193 ( .D(wrtCnt[25]), .QTFCLK( ), .Q(wrtCntD[25]));
Q_FDP0UA U5194 ( .D(wrtCnt[24]), .QTFCLK( ), .Q(wrtCntD[24]));
Q_FDP0UA U5195 ( .D(wrtCnt[23]), .QTFCLK( ), .Q(wrtCntD[23]));
Q_FDP0UA U5196 ( .D(wrtCnt[22]), .QTFCLK( ), .Q(wrtCntD[22]));
Q_FDP0UA U5197 ( .D(wrtCnt[21]), .QTFCLK( ), .Q(wrtCntD[21]));
Q_FDP0UA U5198 ( .D(wrtCnt[20]), .QTFCLK( ), .Q(wrtCntD[20]));
Q_FDP0UA U5199 ( .D(wrtCnt[19]), .QTFCLK( ), .Q(wrtCntD[19]));
Q_FDP0UA U5200 ( .D(wrtCnt[18]), .QTFCLK( ), .Q(wrtCntD[18]));
Q_FDP0UA U5201 ( .D(wrtCnt[17]), .QTFCLK( ), .Q(wrtCntD[17]));
Q_FDP0UA U5202 ( .D(wrtCnt[16]), .QTFCLK( ), .Q(wrtCntD[16]));
Q_FDP0UA U5203 ( .D(wrtCnt[15]), .QTFCLK( ), .Q(wrtCntD[15]));
Q_FDP0UA U5204 ( .D(wrtCnt[14]), .QTFCLK( ), .Q(wrtCntD[14]));
Q_FDP0UA U5205 ( .D(wrtCnt[13]), .QTFCLK( ), .Q(wrtCntD[13]));
Q_FDP0UA U5206 ( .D(wrtCnt[12]), .QTFCLK( ), .Q(wrtCntD[12]));
Q_FDP0UA U5207 ( .D(wrtCnt[11]), .QTFCLK( ), .Q(wrtCntD[11]));
Q_FDP0UA U5208 ( .D(wrtCnt[10]), .QTFCLK( ), .Q(wrtCntD[10]));
Q_FDP0UA U5209 ( .D(wrtCnt[9]), .QTFCLK( ), .Q(wrtCntD[9]));
Q_FDP0UA U5210 ( .D(wrtCnt[8]), .QTFCLK( ), .Q(wrtCntD[8]));
Q_FDP0UA U5211 ( .D(wrtCnt[7]), .QTFCLK( ), .Q(wrtCntD[7]));
Q_FDP0UA U5212 ( .D(wrtCnt[6]), .QTFCLK( ), .Q(wrtCntD[6]));
Q_FDP0UA U5213 ( .D(wrtCnt[5]), .QTFCLK( ), .Q(wrtCntD[5]));
Q_FDP0UA U5214 ( .D(wrtCnt[4]), .QTFCLK( ), .Q(wrtCntD[4]));
Q_FDP0UA U5215 ( .D(wrtCnt[3]), .QTFCLK( ), .Q(wrtCntD[3]));
Q_FDP0UA U5216 ( .D(wrtCnt[2]), .QTFCLK( ), .Q(wrtCntD[2]));
Q_FDP0UA U5217 ( .D(wrtCnt[1]), .QTFCLK( ), .Q(wrtCntD[1]));
Q_FDP0UA U5218 ( .D(wrtCnt[0]), .QTFCLK( ), .Q(wrtCntD[0]));
Q_AN02 U5219 ( .A0(n1610), .A1(LBwrI[3]), .Z(LBwr[3]));
Q_OR02 U5220 ( .A0(LBfull), .A1(LBwrI[2]), .Z(LBwr[2]));
Q_INV U5221 ( .A(n1610), .Z(LBfull));
Q_AN02 U5222 ( .A0(n1610), .A1(LBwrI[1]), .Z(LBwr[1]));
Q_AN02 U5223 ( .A0(n1610), .A1(LBwrI[0]), .Z(LBwr[0]));
Q_AN02 U5224 ( .A0(LBreq), .A1(LBempty), .Z(n3649));
Q_OA21 U5225 ( .A0(gfTsEn), .A1(n3649), .B0(gfTsReqO), .Z(GFtsAdd));
Q_INV U5226 ( .A(LBwr[3]), .Z(n3648));
Q_INV U5227 ( .A(ofifoAddr0N[0]), .Z(ofifoAddr1N[0]));
Q_AD01HF U5228 ( .A0(ofifoAddr0N[1]), .B0(ofifoAddr0N[0]), .S(ofifoAddr1N[1]), .CO(n3647));
Q_AD01HF U5229 ( .A0(ofifoAddr0N[2]), .B0(n3647), .S(ofifoAddr1N[2]), .CO(n3646));
Q_AD01HF U5230 ( .A0(ofifoAddr0N[3]), .B0(n3646), .S(ofifoAddr1N[3]), .CO(n3645));
Q_AD01HF U5231 ( .A0(ofifoAddr0N[4]), .B0(n3645), .S(ofifoAddr1N[4]), .CO(n3644));
Q_AD01HF U5232 ( .A0(ofifoAddr0N[5]), .B0(n3644), .S(ofifoAddr1N[5]), .CO(n3643));
Q_AD01HF U5233 ( .A0(ofifoAddr0N[6]), .B0(n3643), .S(ofifoAddr1N[6]), .CO(n3642));
Q_AD01HF U5234 ( .A0(ofifoAddr0N[7]), .B0(n3642), .S(ofifoAddr1N[7]), .CO(n3641));
Q_AD01HF U5235 ( .A0(ofifoAddr0N[8]), .B0(n3641), .S(ofifoAddr1N[8]), .CO(n3640));
Q_AD01HF U5236 ( .A0(ofifoAddr0N[9]), .B0(n3640), .S(ofifoAddr1N[9]), .CO(n3639));
Q_AD01HF U5237 ( .A0(ofifoAddr0N[10]), .B0(n3639), .S(ofifoAddr1N[10]), .CO(n3638));
Q_AD01HF U5238 ( .A0(ofifoAddr0N[11]), .B0(n3638), .S(ofifoAddr1N[11]), .CO(n3637));
Q_AD01HF U5239 ( .A0(ofifoAddr0N[12]), .B0(n3637), .S(ofifoAddr1N[12]), .CO(n3636));
Q_AD01HF U5240 ( .A0(ofifoAddr0N[13]), .B0(n3636), .S(ofifoAddr1N[13]), .CO(n3635));
Q_XOR2 U5241 ( .A0(ofifoAddr0N[14]), .A1(n3635), .Z(ofifoAddr1N[14]));
Q_INV U5242 ( .A(ofifoAddr0N[1]), .Z(ofifoAddr2N[1]));
Q_AD01HF U5243 ( .A0(ofifoAddr0N[2]), .B0(ofifoAddr0N[1]), .S(ofifoAddr2N[2]), .CO(n3634));
Q_AD01HF U5244 ( .A0(ofifoAddr0N[3]), .B0(n3634), .S(ofifoAddr2N[3]), .CO(n3633));
Q_AD01HF U5245 ( .A0(ofifoAddr0N[4]), .B0(n3633), .S(ofifoAddr2N[4]), .CO(n3632));
Q_AD01HF U5246 ( .A0(ofifoAddr0N[5]), .B0(n3632), .S(ofifoAddr2N[5]), .CO(n3631));
Q_AD01HF U5247 ( .A0(ofifoAddr0N[6]), .B0(n3631), .S(ofifoAddr2N[6]), .CO(n3630));
Q_AD01HF U5248 ( .A0(ofifoAddr0N[7]), .B0(n3630), .S(ofifoAddr2N[7]), .CO(n3629));
Q_AD01HF U5249 ( .A0(ofifoAddr0N[8]), .B0(n3629), .S(ofifoAddr2N[8]), .CO(n3628));
Q_AD01HF U5250 ( .A0(ofifoAddr0N[9]), .B0(n3628), .S(ofifoAddr2N[9]), .CO(n3627));
Q_AD01HF U5251 ( .A0(ofifoAddr0N[10]), .B0(n3627), .S(ofifoAddr2N[10]), .CO(n3626));
Q_AD01HF U5252 ( .A0(ofifoAddr0N[11]), .B0(n3626), .S(ofifoAddr2N[11]), .CO(n3625));
Q_AD01HF U5253 ( .A0(ofifoAddr0N[12]), .B0(n3625), .S(ofifoAddr2N[12]), .CO(n3624));
Q_AD01HF U5254 ( .A0(ofifoAddr0N[13]), .B0(n3624), .S(ofifoAddr2N[13]), .CO(n3623));
Q_XOR2 U5255 ( .A0(ofifoAddr0N[14]), .A1(n3623), .Z(ofifoAddr2N[14]));
Q_AN02 U5256 ( .A0(shiftCount[5]), .A1(xdata[543]), .Z(n3622));
Q_AN02 U5257 ( .A0(shiftCount[5]), .A1(xdata[542]), .Z(n3621));
Q_AN02 U5258 ( .A0(shiftCount[5]), .A1(xdata[541]), .Z(n3620));
Q_AN02 U5259 ( .A0(shiftCount[5]), .A1(xdata[540]), .Z(n3619));
Q_AN02 U5260 ( .A0(shiftCount[5]), .A1(xdata[539]), .Z(n3618));
Q_AN02 U5261 ( .A0(shiftCount[5]), .A1(xdata[538]), .Z(n3617));
Q_AN02 U5262 ( .A0(shiftCount[5]), .A1(xdata[537]), .Z(n3616));
Q_AN02 U5263 ( .A0(shiftCount[5]), .A1(xdata[536]), .Z(n3615));
Q_AN02 U5264 ( .A0(shiftCount[5]), .A1(xdata[535]), .Z(n3614));
Q_AN02 U5265 ( .A0(shiftCount[5]), .A1(xdata[534]), .Z(n3613));
Q_AN02 U5266 ( .A0(shiftCount[5]), .A1(xdata[533]), .Z(n3612));
Q_AN02 U5267 ( .A0(shiftCount[5]), .A1(xdata[532]), .Z(n3611));
Q_AN02 U5268 ( .A0(shiftCount[5]), .A1(xdata[531]), .Z(n3610));
Q_AN02 U5269 ( .A0(shiftCount[5]), .A1(xdata[530]), .Z(n3609));
Q_AN02 U5270 ( .A0(shiftCount[5]), .A1(xdata[529]), .Z(n3608));
Q_AN02 U5271 ( .A0(shiftCount[5]), .A1(xdata[528]), .Z(n3607));
Q_AN02 U5272 ( .A0(shiftCount[5]), .A1(xdata[527]), .Z(n3606));
Q_AN02 U5273 ( .A0(shiftCount[5]), .A1(xdata[526]), .Z(n3605));
Q_AN02 U5274 ( .A0(shiftCount[5]), .A1(xdata[525]), .Z(n3604));
Q_AN02 U5275 ( .A0(shiftCount[5]), .A1(xdata[524]), .Z(n3603));
Q_AN02 U5276 ( .A0(shiftCount[5]), .A1(xdata[523]), .Z(n3602));
Q_AN02 U5277 ( .A0(shiftCount[5]), .A1(xdata[522]), .Z(n3601));
Q_AN02 U5278 ( .A0(shiftCount[5]), .A1(xdata[521]), .Z(n3600));
Q_AN02 U5279 ( .A0(shiftCount[5]), .A1(xdata[520]), .Z(n3599));
Q_AN02 U5280 ( .A0(shiftCount[5]), .A1(xdata[519]), .Z(n3598));
Q_AN02 U5281 ( .A0(shiftCount[5]), .A1(xdata[518]), .Z(n3597));
Q_AN02 U5282 ( .A0(shiftCount[5]), .A1(xdata[517]), .Z(n3596));
Q_AN02 U5283 ( .A0(shiftCount[5]), .A1(xdata[516]), .Z(n3595));
Q_AN02 U5284 ( .A0(shiftCount[5]), .A1(xdata[515]), .Z(n3594));
Q_AN02 U5285 ( .A0(shiftCount[5]), .A1(xdata[514]), .Z(n3593));
Q_AN02 U5286 ( .A0(shiftCount[5]), .A1(xdata[513]), .Z(n3592));
Q_AN02 U5287 ( .A0(shiftCount[5]), .A1(xdata[512]), .Z(n3591));
Q_MX02 U5288 ( .S(shiftCount[5]), .A0(xdata[543]), .A1(xdata[511]), .Z(n3590));
Q_MX02 U5289 ( .S(shiftCount[5]), .A0(xdata[542]), .A1(xdata[510]), .Z(n3589));
Q_MX02 U5290 ( .S(shiftCount[5]), .A0(xdata[541]), .A1(xdata[509]), .Z(n3588));
Q_MX02 U5291 ( .S(shiftCount[5]), .A0(xdata[540]), .A1(xdata[508]), .Z(n3587));
Q_MX02 U5292 ( .S(shiftCount[5]), .A0(xdata[539]), .A1(xdata[507]), .Z(n3586));
Q_MX02 U5293 ( .S(shiftCount[5]), .A0(xdata[538]), .A1(xdata[506]), .Z(n3585));
Q_MX02 U5294 ( .S(shiftCount[5]), .A0(xdata[537]), .A1(xdata[505]), .Z(n3584));
Q_MX02 U5295 ( .S(shiftCount[5]), .A0(xdata[536]), .A1(xdata[504]), .Z(n3583));
Q_MX02 U5296 ( .S(shiftCount[5]), .A0(xdata[535]), .A1(xdata[503]), .Z(n3582));
Q_MX02 U5297 ( .S(shiftCount[5]), .A0(xdata[534]), .A1(xdata[502]), .Z(n3581));
Q_MX02 U5298 ( .S(shiftCount[5]), .A0(xdata[533]), .A1(xdata[501]), .Z(n3580));
Q_MX02 U5299 ( .S(shiftCount[5]), .A0(xdata[532]), .A1(xdata[500]), .Z(n3579));
Q_MX02 U5300 ( .S(shiftCount[5]), .A0(xdata[531]), .A1(xdata[499]), .Z(n3578));
Q_MX02 U5301 ( .S(shiftCount[5]), .A0(xdata[530]), .A1(xdata[498]), .Z(n3577));
Q_MX02 U5302 ( .S(shiftCount[5]), .A0(xdata[529]), .A1(xdata[497]), .Z(n3576));
Q_MX02 U5303 ( .S(shiftCount[5]), .A0(xdata[528]), .A1(xdata[496]), .Z(n3575));
Q_MX02 U5304 ( .S(shiftCount[5]), .A0(xdata[527]), .A1(xdata[495]), .Z(n3574));
Q_MX02 U5305 ( .S(shiftCount[5]), .A0(xdata[526]), .A1(xdata[494]), .Z(n3573));
Q_MX02 U5306 ( .S(shiftCount[5]), .A0(xdata[525]), .A1(xdata[493]), .Z(n3572));
Q_MX02 U5307 ( .S(shiftCount[5]), .A0(xdata[524]), .A1(xdata[492]), .Z(n3571));
Q_MX02 U5308 ( .S(shiftCount[5]), .A0(xdata[523]), .A1(xdata[491]), .Z(n3570));
Q_MX02 U5309 ( .S(shiftCount[5]), .A0(xdata[522]), .A1(xdata[490]), .Z(n3569));
Q_MX02 U5310 ( .S(shiftCount[5]), .A0(xdata[521]), .A1(xdata[489]), .Z(n3568));
Q_MX02 U5311 ( .S(shiftCount[5]), .A0(xdata[520]), .A1(xdata[488]), .Z(n3567));
Q_MX02 U5312 ( .S(shiftCount[5]), .A0(xdata[519]), .A1(xdata[487]), .Z(n3566));
Q_MX02 U5313 ( .S(shiftCount[5]), .A0(xdata[518]), .A1(xdata[486]), .Z(n3565));
Q_MX02 U5314 ( .S(shiftCount[5]), .A0(xdata[517]), .A1(xdata[485]), .Z(n3564));
Q_MX02 U5315 ( .S(shiftCount[5]), .A0(xdata[516]), .A1(xdata[484]), .Z(n3563));
Q_MX02 U5316 ( .S(shiftCount[5]), .A0(xdata[515]), .A1(xdata[483]), .Z(n3562));
Q_MX02 U5317 ( .S(shiftCount[5]), .A0(xdata[514]), .A1(xdata[482]), .Z(n3561));
Q_MX02 U5318 ( .S(shiftCount[5]), .A0(xdata[513]), .A1(xdata[481]), .Z(n3560));
Q_MX02 U5319 ( .S(shiftCount[5]), .A0(xdata[512]), .A1(xdata[480]), .Z(n3559));
Q_MX02 U5320 ( .S(shiftCount[5]), .A0(xdata[511]), .A1(xdata[479]), .Z(n3558));
Q_MX02 U5321 ( .S(shiftCount[5]), .A0(xdata[510]), .A1(xdata[478]), .Z(n3557));
Q_MX02 U5322 ( .S(shiftCount[5]), .A0(xdata[509]), .A1(xdata[477]), .Z(n3556));
Q_MX02 U5323 ( .S(shiftCount[5]), .A0(xdata[508]), .A1(xdata[476]), .Z(n3555));
Q_MX02 U5324 ( .S(shiftCount[5]), .A0(xdata[507]), .A1(xdata[475]), .Z(n3554));
Q_MX02 U5325 ( .S(shiftCount[5]), .A0(xdata[506]), .A1(xdata[474]), .Z(n3553));
Q_MX02 U5326 ( .S(shiftCount[5]), .A0(xdata[505]), .A1(xdata[473]), .Z(n3552));
Q_MX02 U5327 ( .S(shiftCount[5]), .A0(xdata[504]), .A1(xdata[472]), .Z(n3551));
Q_MX02 U5328 ( .S(shiftCount[5]), .A0(xdata[503]), .A1(xdata[471]), .Z(n3550));
Q_MX02 U5329 ( .S(shiftCount[5]), .A0(xdata[502]), .A1(xdata[470]), .Z(n3549));
Q_MX02 U5330 ( .S(shiftCount[5]), .A0(xdata[501]), .A1(xdata[469]), .Z(n3548));
Q_MX02 U5331 ( .S(shiftCount[5]), .A0(xdata[500]), .A1(xdata[468]), .Z(n3547));
Q_MX02 U5332 ( .S(shiftCount[5]), .A0(xdata[499]), .A1(xdata[467]), .Z(n3546));
Q_MX02 U5333 ( .S(shiftCount[5]), .A0(xdata[498]), .A1(xdata[466]), .Z(n3545));
Q_MX02 U5334 ( .S(shiftCount[5]), .A0(xdata[497]), .A1(xdata[465]), .Z(n3544));
Q_MX02 U5335 ( .S(shiftCount[5]), .A0(xdata[496]), .A1(xdata[464]), .Z(n3543));
Q_MX02 U5336 ( .S(shiftCount[5]), .A0(xdata[495]), .A1(xdata[463]), .Z(n3542));
Q_MX02 U5337 ( .S(shiftCount[5]), .A0(xdata[494]), .A1(xdata[462]), .Z(n3541));
Q_MX02 U5338 ( .S(shiftCount[5]), .A0(xdata[493]), .A1(xdata[461]), .Z(n3540));
Q_MX02 U5339 ( .S(shiftCount[5]), .A0(xdata[492]), .A1(xdata[460]), .Z(n3539));
Q_MX02 U5340 ( .S(shiftCount[5]), .A0(xdata[491]), .A1(xdata[459]), .Z(n3538));
Q_MX02 U5341 ( .S(shiftCount[5]), .A0(xdata[490]), .A1(xdata[458]), .Z(n3537));
Q_MX02 U5342 ( .S(shiftCount[5]), .A0(xdata[489]), .A1(xdata[457]), .Z(n3536));
Q_MX02 U5343 ( .S(shiftCount[5]), .A0(xdata[488]), .A1(xdata[456]), .Z(n3535));
Q_MX02 U5344 ( .S(shiftCount[5]), .A0(xdata[487]), .A1(xdata[455]), .Z(n3534));
Q_MX02 U5345 ( .S(shiftCount[5]), .A0(xdata[486]), .A1(xdata[454]), .Z(n3533));
Q_MX02 U5346 ( .S(shiftCount[5]), .A0(xdata[485]), .A1(xdata[453]), .Z(n3532));
Q_MX02 U5347 ( .S(shiftCount[5]), .A0(xdata[484]), .A1(xdata[452]), .Z(n3531));
Q_MX02 U5348 ( .S(shiftCount[5]), .A0(xdata[483]), .A1(xdata[451]), .Z(n3530));
Q_MX02 U5349 ( .S(shiftCount[5]), .A0(xdata[482]), .A1(xdata[450]), .Z(n3529));
Q_MX02 U5350 ( .S(shiftCount[5]), .A0(xdata[481]), .A1(xdata[449]), .Z(n3528));
Q_MX02 U5351 ( .S(shiftCount[5]), .A0(xdata[480]), .A1(xdata[448]), .Z(n3527));
Q_MX02 U5352 ( .S(shiftCount[5]), .A0(xdata[479]), .A1(xdata[447]), .Z(n3526));
Q_MX02 U5353 ( .S(shiftCount[5]), .A0(xdata[478]), .A1(xdata[446]), .Z(n3525));
Q_MX02 U5354 ( .S(shiftCount[5]), .A0(xdata[477]), .A1(xdata[445]), .Z(n3524));
Q_MX02 U5355 ( .S(shiftCount[5]), .A0(xdata[476]), .A1(xdata[444]), .Z(n3523));
Q_MX02 U5356 ( .S(shiftCount[5]), .A0(xdata[475]), .A1(xdata[443]), .Z(n3522));
Q_MX02 U5357 ( .S(shiftCount[5]), .A0(xdata[474]), .A1(xdata[442]), .Z(n3521));
Q_MX02 U5358 ( .S(shiftCount[5]), .A0(xdata[473]), .A1(xdata[441]), .Z(n3520));
Q_MX02 U5359 ( .S(shiftCount[5]), .A0(xdata[472]), .A1(xdata[440]), .Z(n3519));
Q_MX02 U5360 ( .S(shiftCount[5]), .A0(xdata[471]), .A1(xdata[439]), .Z(n3518));
Q_MX02 U5361 ( .S(shiftCount[5]), .A0(xdata[470]), .A1(xdata[438]), .Z(n3517));
Q_MX02 U5362 ( .S(shiftCount[5]), .A0(xdata[469]), .A1(xdata[437]), .Z(n3516));
Q_MX02 U5363 ( .S(shiftCount[5]), .A0(xdata[468]), .A1(xdata[436]), .Z(n3515));
Q_MX02 U5364 ( .S(shiftCount[5]), .A0(xdata[467]), .A1(xdata[435]), .Z(n3514));
Q_MX02 U5365 ( .S(shiftCount[5]), .A0(xdata[466]), .A1(xdata[434]), .Z(n3513));
Q_MX02 U5366 ( .S(shiftCount[5]), .A0(xdata[465]), .A1(xdata[433]), .Z(n3512));
Q_MX02 U5367 ( .S(shiftCount[5]), .A0(xdata[464]), .A1(xdata[432]), .Z(n3511));
Q_MX02 U5368 ( .S(shiftCount[5]), .A0(xdata[463]), .A1(xdata[431]), .Z(n3510));
Q_MX02 U5369 ( .S(shiftCount[5]), .A0(xdata[462]), .A1(xdata[430]), .Z(n3509));
Q_MX02 U5370 ( .S(shiftCount[5]), .A0(xdata[461]), .A1(xdata[429]), .Z(n3508));
Q_MX02 U5371 ( .S(shiftCount[5]), .A0(xdata[460]), .A1(xdata[428]), .Z(n3507));
Q_MX02 U5372 ( .S(shiftCount[5]), .A0(xdata[459]), .A1(xdata[427]), .Z(n3506));
Q_MX02 U5373 ( .S(shiftCount[5]), .A0(xdata[458]), .A1(xdata[426]), .Z(n3505));
Q_MX02 U5374 ( .S(shiftCount[5]), .A0(xdata[457]), .A1(xdata[425]), .Z(n3504));
Q_MX02 U5375 ( .S(shiftCount[5]), .A0(xdata[456]), .A1(xdata[424]), .Z(n3503));
Q_MX02 U5376 ( .S(shiftCount[5]), .A0(xdata[455]), .A1(xdata[423]), .Z(n3502));
Q_MX02 U5377 ( .S(shiftCount[5]), .A0(xdata[454]), .A1(xdata[422]), .Z(n3501));
Q_MX02 U5378 ( .S(shiftCount[5]), .A0(xdata[453]), .A1(xdata[421]), .Z(n3500));
Q_MX02 U5379 ( .S(shiftCount[5]), .A0(xdata[452]), .A1(xdata[420]), .Z(n3499));
Q_MX02 U5380 ( .S(shiftCount[5]), .A0(xdata[451]), .A1(xdata[419]), .Z(n3498));
Q_MX02 U5381 ( .S(shiftCount[5]), .A0(xdata[450]), .A1(xdata[418]), .Z(n3497));
Q_MX02 U5382 ( .S(shiftCount[5]), .A0(xdata[449]), .A1(xdata[417]), .Z(n3496));
Q_MX02 U5383 ( .S(shiftCount[5]), .A0(xdata[448]), .A1(xdata[416]), .Z(n3495));
Q_MX02 U5384 ( .S(shiftCount[5]), .A0(xdata[447]), .A1(xdata[415]), .Z(n3494));
Q_MX02 U5385 ( .S(shiftCount[5]), .A0(xdata[446]), .A1(xdata[414]), .Z(n3493));
Q_MX02 U5386 ( .S(shiftCount[5]), .A0(xdata[445]), .A1(xdata[413]), .Z(n3492));
Q_MX02 U5387 ( .S(shiftCount[5]), .A0(xdata[444]), .A1(xdata[412]), .Z(n3491));
Q_MX02 U5388 ( .S(shiftCount[5]), .A0(xdata[443]), .A1(xdata[411]), .Z(n3490));
Q_MX02 U5389 ( .S(shiftCount[5]), .A0(xdata[442]), .A1(xdata[410]), .Z(n3489));
Q_MX02 U5390 ( .S(shiftCount[5]), .A0(xdata[441]), .A1(xdata[409]), .Z(n3488));
Q_MX02 U5391 ( .S(shiftCount[5]), .A0(xdata[440]), .A1(xdata[408]), .Z(n3487));
Q_MX02 U5392 ( .S(shiftCount[5]), .A0(xdata[439]), .A1(xdata[407]), .Z(n3486));
Q_MX02 U5393 ( .S(shiftCount[5]), .A0(xdata[438]), .A1(xdata[406]), .Z(n3485));
Q_MX02 U5394 ( .S(shiftCount[5]), .A0(xdata[437]), .A1(xdata[405]), .Z(n3484));
Q_MX02 U5395 ( .S(shiftCount[5]), .A0(xdata[436]), .A1(xdata[404]), .Z(n3483));
Q_MX02 U5396 ( .S(shiftCount[5]), .A0(xdata[435]), .A1(xdata[403]), .Z(n3482));
Q_MX02 U5397 ( .S(shiftCount[5]), .A0(xdata[434]), .A1(xdata[402]), .Z(n3481));
Q_MX02 U5398 ( .S(shiftCount[5]), .A0(xdata[433]), .A1(xdata[401]), .Z(n3480));
Q_MX02 U5399 ( .S(shiftCount[5]), .A0(xdata[432]), .A1(xdata[400]), .Z(n3479));
Q_MX02 U5400 ( .S(shiftCount[5]), .A0(xdata[431]), .A1(xdata[399]), .Z(n3478));
Q_MX02 U5401 ( .S(shiftCount[5]), .A0(xdata[430]), .A1(xdata[398]), .Z(n3477));
Q_MX02 U5402 ( .S(shiftCount[5]), .A0(xdata[429]), .A1(xdata[397]), .Z(n3476));
Q_MX02 U5403 ( .S(shiftCount[5]), .A0(xdata[428]), .A1(xdata[396]), .Z(n3475));
Q_MX02 U5404 ( .S(shiftCount[5]), .A0(xdata[427]), .A1(xdata[395]), .Z(n3474));
Q_MX02 U5405 ( .S(shiftCount[5]), .A0(xdata[426]), .A1(xdata[394]), .Z(n3473));
Q_MX02 U5406 ( .S(shiftCount[5]), .A0(xdata[425]), .A1(xdata[393]), .Z(n3472));
Q_MX02 U5407 ( .S(shiftCount[5]), .A0(xdata[424]), .A1(xdata[392]), .Z(n3471));
Q_MX02 U5408 ( .S(shiftCount[5]), .A0(xdata[423]), .A1(xdata[391]), .Z(n3470));
Q_MX02 U5409 ( .S(shiftCount[5]), .A0(xdata[422]), .A1(xdata[390]), .Z(n3469));
Q_MX02 U5410 ( .S(shiftCount[5]), .A0(xdata[421]), .A1(xdata[389]), .Z(n3468));
Q_MX02 U5411 ( .S(shiftCount[5]), .A0(xdata[420]), .A1(xdata[388]), .Z(n3467));
Q_MX02 U5412 ( .S(shiftCount[5]), .A0(xdata[419]), .A1(xdata[387]), .Z(n3466));
Q_MX02 U5413 ( .S(shiftCount[5]), .A0(xdata[418]), .A1(xdata[386]), .Z(n3465));
Q_MX02 U5414 ( .S(shiftCount[5]), .A0(xdata[417]), .A1(xdata[385]), .Z(n3464));
Q_MX02 U5415 ( .S(shiftCount[5]), .A0(xdata[416]), .A1(xdata[384]), .Z(n3463));
Q_MX02 U5416 ( .S(shiftCount[5]), .A0(xdata[415]), .A1(xdata[383]), .Z(n3462));
Q_MX02 U5417 ( .S(shiftCount[5]), .A0(xdata[414]), .A1(xdata[382]), .Z(n3461));
Q_MX02 U5418 ( .S(shiftCount[5]), .A0(xdata[413]), .A1(xdata[381]), .Z(n3460));
Q_MX02 U5419 ( .S(shiftCount[5]), .A0(xdata[412]), .A1(xdata[380]), .Z(n3459));
Q_MX02 U5420 ( .S(shiftCount[5]), .A0(xdata[411]), .A1(xdata[379]), .Z(n3458));
Q_MX02 U5421 ( .S(shiftCount[5]), .A0(xdata[410]), .A1(xdata[378]), .Z(n3457));
Q_MX02 U5422 ( .S(shiftCount[5]), .A0(xdata[409]), .A1(xdata[377]), .Z(n3456));
Q_MX02 U5423 ( .S(shiftCount[5]), .A0(xdata[408]), .A1(xdata[376]), .Z(n3455));
Q_MX02 U5424 ( .S(shiftCount[5]), .A0(xdata[407]), .A1(xdata[375]), .Z(n3454));
Q_MX02 U5425 ( .S(shiftCount[5]), .A0(xdata[406]), .A1(xdata[374]), .Z(n3453));
Q_MX02 U5426 ( .S(shiftCount[5]), .A0(xdata[405]), .A1(xdata[373]), .Z(n3452));
Q_MX02 U5427 ( .S(shiftCount[5]), .A0(xdata[404]), .A1(xdata[372]), .Z(n3451));
Q_MX02 U5428 ( .S(shiftCount[5]), .A0(xdata[403]), .A1(xdata[371]), .Z(n3450));
Q_MX02 U5429 ( .S(shiftCount[5]), .A0(xdata[402]), .A1(xdata[370]), .Z(n3449));
Q_MX02 U5430 ( .S(shiftCount[5]), .A0(xdata[401]), .A1(xdata[369]), .Z(n3448));
Q_MX02 U5431 ( .S(shiftCount[5]), .A0(xdata[400]), .A1(xdata[368]), .Z(n3447));
Q_MX02 U5432 ( .S(shiftCount[5]), .A0(xdata[399]), .A1(xdata[367]), .Z(n3446));
Q_MX02 U5433 ( .S(shiftCount[5]), .A0(xdata[398]), .A1(xdata[366]), .Z(n3445));
Q_MX02 U5434 ( .S(shiftCount[5]), .A0(xdata[397]), .A1(xdata[365]), .Z(n3444));
Q_MX02 U5435 ( .S(shiftCount[5]), .A0(xdata[396]), .A1(xdata[364]), .Z(n3443));
Q_MX02 U5436 ( .S(shiftCount[5]), .A0(xdata[395]), .A1(xdata[363]), .Z(n3442));
Q_MX02 U5437 ( .S(shiftCount[5]), .A0(xdata[394]), .A1(xdata[362]), .Z(n3441));
Q_MX02 U5438 ( .S(shiftCount[5]), .A0(xdata[393]), .A1(xdata[361]), .Z(n3440));
Q_MX02 U5439 ( .S(shiftCount[5]), .A0(xdata[392]), .A1(xdata[360]), .Z(n3439));
Q_MX02 U5440 ( .S(shiftCount[5]), .A0(xdata[391]), .A1(xdata[359]), .Z(n3438));
Q_MX02 U5441 ( .S(shiftCount[5]), .A0(xdata[390]), .A1(xdata[358]), .Z(n3437));
Q_MX02 U5442 ( .S(shiftCount[5]), .A0(xdata[389]), .A1(xdata[357]), .Z(n3436));
Q_MX02 U5443 ( .S(shiftCount[5]), .A0(xdata[388]), .A1(xdata[356]), .Z(n3435));
Q_MX02 U5444 ( .S(shiftCount[5]), .A0(xdata[387]), .A1(xdata[355]), .Z(n3434));
Q_MX02 U5445 ( .S(shiftCount[5]), .A0(xdata[386]), .A1(xdata[354]), .Z(n3433));
Q_MX02 U5446 ( .S(shiftCount[5]), .A0(xdata[385]), .A1(xdata[353]), .Z(n3432));
Q_MX02 U5447 ( .S(shiftCount[5]), .A0(xdata[384]), .A1(xdata[352]), .Z(n3431));
Q_MX02 U5448 ( .S(shiftCount[5]), .A0(xdata[383]), .A1(xdata[351]), .Z(n3430));
Q_MX02 U5449 ( .S(shiftCount[5]), .A0(xdata[382]), .A1(xdata[350]), .Z(n3429));
Q_MX02 U5450 ( .S(shiftCount[5]), .A0(xdata[381]), .A1(xdata[349]), .Z(n3428));
Q_MX02 U5451 ( .S(shiftCount[5]), .A0(xdata[380]), .A1(xdata[348]), .Z(n3427));
Q_MX02 U5452 ( .S(shiftCount[5]), .A0(xdata[379]), .A1(xdata[347]), .Z(n3426));
Q_MX02 U5453 ( .S(shiftCount[5]), .A0(xdata[378]), .A1(xdata[346]), .Z(n3425));
Q_MX02 U5454 ( .S(shiftCount[5]), .A0(xdata[377]), .A1(xdata[345]), .Z(n3424));
Q_MX02 U5455 ( .S(shiftCount[5]), .A0(xdata[376]), .A1(xdata[344]), .Z(n3423));
Q_MX02 U5456 ( .S(shiftCount[5]), .A0(xdata[375]), .A1(xdata[343]), .Z(n3422));
Q_MX02 U5457 ( .S(shiftCount[5]), .A0(xdata[374]), .A1(xdata[342]), .Z(n3421));
Q_MX02 U5458 ( .S(shiftCount[5]), .A0(xdata[373]), .A1(xdata[341]), .Z(n3420));
Q_MX02 U5459 ( .S(shiftCount[5]), .A0(xdata[372]), .A1(xdata[340]), .Z(n3419));
Q_MX02 U5460 ( .S(shiftCount[5]), .A0(xdata[371]), .A1(xdata[339]), .Z(n3418));
Q_MX02 U5461 ( .S(shiftCount[5]), .A0(xdata[370]), .A1(xdata[338]), .Z(n3417));
Q_MX02 U5462 ( .S(shiftCount[5]), .A0(xdata[369]), .A1(xdata[337]), .Z(n3416));
Q_MX02 U5463 ( .S(shiftCount[5]), .A0(xdata[368]), .A1(xdata[336]), .Z(n3415));
Q_MX02 U5464 ( .S(shiftCount[5]), .A0(xdata[367]), .A1(xdata[335]), .Z(n3414));
Q_MX02 U5465 ( .S(shiftCount[5]), .A0(xdata[366]), .A1(xdata[334]), .Z(n3413));
Q_MX02 U5466 ( .S(shiftCount[5]), .A0(xdata[365]), .A1(xdata[333]), .Z(n3412));
Q_MX02 U5467 ( .S(shiftCount[5]), .A0(xdata[364]), .A1(xdata[332]), .Z(n3411));
Q_MX02 U5468 ( .S(shiftCount[5]), .A0(xdata[363]), .A1(xdata[331]), .Z(n3410));
Q_MX02 U5469 ( .S(shiftCount[5]), .A0(xdata[362]), .A1(xdata[330]), .Z(n3409));
Q_MX02 U5470 ( .S(shiftCount[5]), .A0(xdata[361]), .A1(xdata[329]), .Z(n3408));
Q_MX02 U5471 ( .S(shiftCount[5]), .A0(xdata[360]), .A1(xdata[328]), .Z(n3407));
Q_MX02 U5472 ( .S(shiftCount[5]), .A0(xdata[359]), .A1(xdata[327]), .Z(n3406));
Q_MX02 U5473 ( .S(shiftCount[5]), .A0(xdata[358]), .A1(xdata[326]), .Z(n3405));
Q_MX02 U5474 ( .S(shiftCount[5]), .A0(xdata[357]), .A1(xdata[325]), .Z(n3404));
Q_MX02 U5475 ( .S(shiftCount[5]), .A0(xdata[356]), .A1(xdata[324]), .Z(n3403));
Q_MX02 U5476 ( .S(shiftCount[5]), .A0(xdata[355]), .A1(xdata[323]), .Z(n3402));
Q_MX02 U5477 ( .S(shiftCount[5]), .A0(xdata[354]), .A1(xdata[322]), .Z(n3401));
Q_MX02 U5478 ( .S(shiftCount[5]), .A0(xdata[353]), .A1(xdata[321]), .Z(n3400));
Q_MX02 U5479 ( .S(shiftCount[5]), .A0(xdata[352]), .A1(xdata[320]), .Z(n3399));
Q_MX02 U5480 ( .S(shiftCount[5]), .A0(xdata[351]), .A1(xdata[319]), .Z(n3398));
Q_MX02 U5481 ( .S(shiftCount[5]), .A0(xdata[350]), .A1(xdata[318]), .Z(n3397));
Q_MX02 U5482 ( .S(shiftCount[5]), .A0(xdata[349]), .A1(xdata[317]), .Z(n3396));
Q_MX02 U5483 ( .S(shiftCount[5]), .A0(xdata[348]), .A1(xdata[316]), .Z(n3395));
Q_MX02 U5484 ( .S(shiftCount[5]), .A0(xdata[347]), .A1(xdata[315]), .Z(n3394));
Q_MX02 U5485 ( .S(shiftCount[5]), .A0(xdata[346]), .A1(xdata[314]), .Z(n3393));
Q_MX02 U5486 ( .S(shiftCount[5]), .A0(xdata[345]), .A1(xdata[313]), .Z(n3392));
Q_MX02 U5487 ( .S(shiftCount[5]), .A0(xdata[344]), .A1(xdata[312]), .Z(n3391));
Q_MX02 U5488 ( .S(shiftCount[5]), .A0(xdata[343]), .A1(xdata[311]), .Z(n3390));
Q_MX02 U5489 ( .S(shiftCount[5]), .A0(xdata[342]), .A1(xdata[310]), .Z(n3389));
Q_MX02 U5490 ( .S(shiftCount[5]), .A0(xdata[341]), .A1(xdata[309]), .Z(n3388));
Q_MX02 U5491 ( .S(shiftCount[5]), .A0(xdata[340]), .A1(xdata[308]), .Z(n3387));
Q_MX02 U5492 ( .S(shiftCount[5]), .A0(xdata[339]), .A1(xdata[307]), .Z(n3386));
Q_MX02 U5493 ( .S(shiftCount[5]), .A0(xdata[338]), .A1(xdata[306]), .Z(n3385));
Q_MX02 U5494 ( .S(shiftCount[5]), .A0(xdata[337]), .A1(xdata[305]), .Z(n3384));
Q_MX02 U5495 ( .S(shiftCount[5]), .A0(xdata[336]), .A1(xdata[304]), .Z(n3383));
Q_MX02 U5496 ( .S(shiftCount[5]), .A0(xdata[335]), .A1(xdata[303]), .Z(n3382));
Q_MX02 U5497 ( .S(shiftCount[5]), .A0(xdata[334]), .A1(xdata[302]), .Z(n3381));
Q_MX02 U5498 ( .S(shiftCount[5]), .A0(xdata[333]), .A1(xdata[301]), .Z(n3380));
Q_MX02 U5499 ( .S(shiftCount[5]), .A0(xdata[332]), .A1(xdata[300]), .Z(n3379));
Q_MX02 U5500 ( .S(shiftCount[5]), .A0(xdata[331]), .A1(xdata[299]), .Z(n3378));
Q_MX02 U5501 ( .S(shiftCount[5]), .A0(xdata[330]), .A1(xdata[298]), .Z(n3377));
Q_MX02 U5502 ( .S(shiftCount[5]), .A0(xdata[329]), .A1(xdata[297]), .Z(n3376));
Q_MX02 U5503 ( .S(shiftCount[5]), .A0(xdata[328]), .A1(xdata[296]), .Z(n3375));
Q_MX02 U5504 ( .S(shiftCount[5]), .A0(xdata[327]), .A1(xdata[295]), .Z(n3374));
Q_MX02 U5505 ( .S(shiftCount[5]), .A0(xdata[326]), .A1(xdata[294]), .Z(n3373));
Q_MX02 U5506 ( .S(shiftCount[5]), .A0(xdata[325]), .A1(xdata[293]), .Z(n3372));
Q_MX02 U5507 ( .S(shiftCount[5]), .A0(xdata[324]), .A1(xdata[292]), .Z(n3371));
Q_MX02 U5508 ( .S(shiftCount[5]), .A0(xdata[323]), .A1(xdata[291]), .Z(n3370));
Q_MX02 U5509 ( .S(shiftCount[5]), .A0(xdata[322]), .A1(xdata[290]), .Z(n3369));
Q_MX02 U5510 ( .S(shiftCount[5]), .A0(xdata[321]), .A1(xdata[289]), .Z(n3368));
Q_MX02 U5511 ( .S(shiftCount[5]), .A0(xdata[320]), .A1(xdata[288]), .Z(n3367));
Q_MX02 U5512 ( .S(shiftCount[5]), .A0(xdata[319]), .A1(xdata[287]), .Z(n3366));
Q_MX02 U5513 ( .S(shiftCount[5]), .A0(xdata[318]), .A1(xdata[286]), .Z(n3365));
Q_MX02 U5514 ( .S(shiftCount[5]), .A0(xdata[317]), .A1(xdata[285]), .Z(n3364));
Q_MX02 U5515 ( .S(shiftCount[5]), .A0(xdata[316]), .A1(xdata[284]), .Z(n3363));
Q_MX02 U5516 ( .S(shiftCount[5]), .A0(xdata[315]), .A1(xdata[283]), .Z(n3362));
Q_MX02 U5517 ( .S(shiftCount[5]), .A0(xdata[314]), .A1(xdata[282]), .Z(n3361));
Q_MX02 U5518 ( .S(shiftCount[5]), .A0(xdata[313]), .A1(xdata[281]), .Z(n3360));
Q_MX02 U5519 ( .S(shiftCount[5]), .A0(xdata[312]), .A1(xdata[280]), .Z(n3359));
Q_MX02 U5520 ( .S(shiftCount[5]), .A0(xdata[311]), .A1(xdata[279]), .Z(n3358));
Q_MX02 U5521 ( .S(shiftCount[5]), .A0(xdata[310]), .A1(xdata[278]), .Z(n3357));
Q_MX02 U5522 ( .S(shiftCount[5]), .A0(xdata[309]), .A1(xdata[277]), .Z(n3356));
Q_MX02 U5523 ( .S(shiftCount[5]), .A0(xdata[308]), .A1(xdata[276]), .Z(n3355));
Q_MX02 U5524 ( .S(shiftCount[5]), .A0(xdata[307]), .A1(xdata[275]), .Z(n3354));
Q_MX02 U5525 ( .S(shiftCount[5]), .A0(xdata[306]), .A1(xdata[274]), .Z(n3353));
Q_MX02 U5526 ( .S(shiftCount[5]), .A0(xdata[305]), .A1(xdata[273]), .Z(n3352));
Q_MX02 U5527 ( .S(shiftCount[5]), .A0(xdata[304]), .A1(xdata[272]), .Z(n3351));
Q_MX02 U5528 ( .S(shiftCount[5]), .A0(xdata[303]), .A1(xdata[271]), .Z(n3350));
Q_MX02 U5529 ( .S(shiftCount[5]), .A0(xdata[302]), .A1(xdata[270]), .Z(n3349));
Q_MX02 U5530 ( .S(shiftCount[5]), .A0(xdata[301]), .A1(xdata[269]), .Z(n3348));
Q_MX02 U5531 ( .S(shiftCount[5]), .A0(xdata[300]), .A1(xdata[268]), .Z(n3347));
Q_MX02 U5532 ( .S(shiftCount[5]), .A0(xdata[299]), .A1(xdata[267]), .Z(n3346));
Q_MX02 U5533 ( .S(shiftCount[5]), .A0(xdata[298]), .A1(xdata[266]), .Z(n3345));
Q_MX02 U5534 ( .S(shiftCount[5]), .A0(xdata[297]), .A1(xdata[265]), .Z(n3344));
Q_MX02 U5535 ( .S(shiftCount[5]), .A0(xdata[296]), .A1(xdata[264]), .Z(n3343));
Q_MX02 U5536 ( .S(shiftCount[5]), .A0(xdata[295]), .A1(xdata[263]), .Z(n3342));
Q_MX02 U5537 ( .S(shiftCount[5]), .A0(xdata[294]), .A1(xdata[262]), .Z(n3341));
Q_MX02 U5538 ( .S(shiftCount[5]), .A0(xdata[293]), .A1(xdata[261]), .Z(n3340));
Q_MX02 U5539 ( .S(shiftCount[5]), .A0(xdata[292]), .A1(xdata[260]), .Z(n3339));
Q_MX02 U5540 ( .S(shiftCount[5]), .A0(xdata[291]), .A1(xdata[259]), .Z(n3338));
Q_MX02 U5541 ( .S(shiftCount[5]), .A0(xdata[290]), .A1(xdata[258]), .Z(n3337));
Q_MX02 U5542 ( .S(shiftCount[5]), .A0(xdata[289]), .A1(xdata[257]), .Z(n3336));
Q_MX02 U5543 ( .S(shiftCount[5]), .A0(xdata[288]), .A1(xdata[256]), .Z(n3335));
Q_MX02 U5544 ( .S(shiftCount[5]), .A0(xdata[287]), .A1(xdata[255]), .Z(n3334));
Q_MX02 U5545 ( .S(shiftCount[5]), .A0(xdata[286]), .A1(xdata[254]), .Z(n3333));
Q_MX02 U5546 ( .S(shiftCount[5]), .A0(xdata[285]), .A1(xdata[253]), .Z(n3332));
Q_MX02 U5547 ( .S(shiftCount[5]), .A0(xdata[284]), .A1(xdata[252]), .Z(n3331));
Q_MX02 U5548 ( .S(shiftCount[5]), .A0(xdata[283]), .A1(xdata[251]), .Z(n3330));
Q_MX02 U5549 ( .S(shiftCount[5]), .A0(xdata[282]), .A1(xdata[250]), .Z(n3329));
Q_MX02 U5550 ( .S(shiftCount[5]), .A0(xdata[281]), .A1(xdata[249]), .Z(n3328));
Q_MX02 U5551 ( .S(shiftCount[5]), .A0(xdata[280]), .A1(xdata[248]), .Z(n3327));
Q_MX02 U5552 ( .S(shiftCount[5]), .A0(xdata[279]), .A1(xdata[247]), .Z(n3326));
Q_MX02 U5553 ( .S(shiftCount[5]), .A0(xdata[278]), .A1(xdata[246]), .Z(n3325));
Q_MX02 U5554 ( .S(shiftCount[5]), .A0(xdata[277]), .A1(xdata[245]), .Z(n3324));
Q_MX02 U5555 ( .S(shiftCount[5]), .A0(xdata[276]), .A1(xdata[244]), .Z(n3323));
Q_MX02 U5556 ( .S(shiftCount[5]), .A0(xdata[275]), .A1(xdata[243]), .Z(n3322));
Q_MX02 U5557 ( .S(shiftCount[5]), .A0(xdata[274]), .A1(xdata[242]), .Z(n3321));
Q_MX02 U5558 ( .S(shiftCount[5]), .A0(xdata[273]), .A1(xdata[241]), .Z(n3320));
Q_MX02 U5559 ( .S(shiftCount[5]), .A0(xdata[272]), .A1(xdata[240]), .Z(n3319));
Q_MX02 U5560 ( .S(shiftCount[5]), .A0(xdata[271]), .A1(xdata[239]), .Z(n3318));
Q_MX02 U5561 ( .S(shiftCount[5]), .A0(xdata[270]), .A1(xdata[238]), .Z(n3317));
Q_MX02 U5562 ( .S(shiftCount[5]), .A0(xdata[269]), .A1(xdata[237]), .Z(n3316));
Q_MX02 U5563 ( .S(shiftCount[5]), .A0(xdata[268]), .A1(xdata[236]), .Z(n3315));
Q_MX02 U5564 ( .S(shiftCount[5]), .A0(xdata[267]), .A1(xdata[235]), .Z(n3314));
Q_MX02 U5565 ( .S(shiftCount[5]), .A0(xdata[266]), .A1(xdata[234]), .Z(n3313));
Q_MX02 U5566 ( .S(shiftCount[5]), .A0(xdata[265]), .A1(xdata[233]), .Z(n3312));
Q_MX02 U5567 ( .S(shiftCount[5]), .A0(xdata[264]), .A1(xdata[232]), .Z(n3311));
Q_MX02 U5568 ( .S(shiftCount[5]), .A0(xdata[263]), .A1(xdata[231]), .Z(n3310));
Q_MX02 U5569 ( .S(shiftCount[5]), .A0(xdata[262]), .A1(xdata[230]), .Z(n3309));
Q_MX02 U5570 ( .S(shiftCount[5]), .A0(xdata[261]), .A1(xdata[229]), .Z(n3308));
Q_MX02 U5571 ( .S(shiftCount[5]), .A0(xdata[260]), .A1(xdata[228]), .Z(n3307));
Q_MX02 U5572 ( .S(shiftCount[5]), .A0(xdata[259]), .A1(xdata[227]), .Z(n3306));
Q_MX02 U5573 ( .S(shiftCount[5]), .A0(xdata[258]), .A1(xdata[226]), .Z(n3305));
Q_MX02 U5574 ( .S(shiftCount[5]), .A0(xdata[257]), .A1(xdata[225]), .Z(n3304));
Q_MX02 U5575 ( .S(shiftCount[5]), .A0(xdata[256]), .A1(xdata[224]), .Z(n3303));
Q_MX02 U5576 ( .S(shiftCount[5]), .A0(xdata[255]), .A1(xdata[223]), .Z(n3302));
Q_MX02 U5577 ( .S(shiftCount[5]), .A0(xdata[254]), .A1(xdata[222]), .Z(n3301));
Q_MX02 U5578 ( .S(shiftCount[5]), .A0(xdata[253]), .A1(xdata[221]), .Z(n3300));
Q_MX02 U5579 ( .S(shiftCount[5]), .A0(xdata[252]), .A1(xdata[220]), .Z(n3299));
Q_MX02 U5580 ( .S(shiftCount[5]), .A0(xdata[251]), .A1(xdata[219]), .Z(n3298));
Q_MX02 U5581 ( .S(shiftCount[5]), .A0(xdata[250]), .A1(xdata[218]), .Z(n3297));
Q_MX02 U5582 ( .S(shiftCount[5]), .A0(xdata[249]), .A1(xdata[217]), .Z(n3296));
Q_MX02 U5583 ( .S(shiftCount[5]), .A0(xdata[248]), .A1(xdata[216]), .Z(n3295));
Q_MX02 U5584 ( .S(shiftCount[5]), .A0(xdata[247]), .A1(xdata[215]), .Z(n3294));
Q_MX02 U5585 ( .S(shiftCount[5]), .A0(xdata[246]), .A1(xdata[214]), .Z(n3293));
Q_MX02 U5586 ( .S(shiftCount[5]), .A0(xdata[245]), .A1(xdata[213]), .Z(n3292));
Q_MX02 U5587 ( .S(shiftCount[5]), .A0(xdata[244]), .A1(xdata[212]), .Z(n3291));
Q_MX02 U5588 ( .S(shiftCount[5]), .A0(xdata[243]), .A1(xdata[211]), .Z(n3290));
Q_MX02 U5589 ( .S(shiftCount[5]), .A0(xdata[242]), .A1(xdata[210]), .Z(n3289));
Q_MX02 U5590 ( .S(shiftCount[5]), .A0(xdata[241]), .A1(xdata[209]), .Z(n3288));
Q_MX02 U5591 ( .S(shiftCount[5]), .A0(xdata[240]), .A1(xdata[208]), .Z(n3287));
Q_MX02 U5592 ( .S(shiftCount[5]), .A0(xdata[239]), .A1(xdata[207]), .Z(n3286));
Q_MX02 U5593 ( .S(shiftCount[5]), .A0(xdata[238]), .A1(xdata[206]), .Z(n3285));
Q_MX02 U5594 ( .S(shiftCount[5]), .A0(xdata[237]), .A1(xdata[205]), .Z(n3284));
Q_MX02 U5595 ( .S(shiftCount[5]), .A0(xdata[236]), .A1(xdata[204]), .Z(n3283));
Q_MX02 U5596 ( .S(shiftCount[5]), .A0(xdata[235]), .A1(xdata[203]), .Z(n3282));
Q_MX02 U5597 ( .S(shiftCount[5]), .A0(xdata[234]), .A1(xdata[202]), .Z(n3281));
Q_MX02 U5598 ( .S(shiftCount[5]), .A0(xdata[233]), .A1(xdata[201]), .Z(n3280));
Q_MX02 U5599 ( .S(shiftCount[5]), .A0(xdata[232]), .A1(xdata[200]), .Z(n3279));
Q_MX02 U5600 ( .S(shiftCount[5]), .A0(xdata[231]), .A1(xdata[199]), .Z(n3278));
Q_MX02 U5601 ( .S(shiftCount[5]), .A0(xdata[230]), .A1(xdata[198]), .Z(n3277));
Q_MX02 U5602 ( .S(shiftCount[5]), .A0(xdata[229]), .A1(xdata[197]), .Z(n3276));
Q_MX02 U5603 ( .S(shiftCount[5]), .A0(xdata[228]), .A1(xdata[196]), .Z(n3275));
Q_MX02 U5604 ( .S(shiftCount[5]), .A0(xdata[227]), .A1(xdata[195]), .Z(n3274));
Q_MX02 U5605 ( .S(shiftCount[5]), .A0(xdata[226]), .A1(xdata[194]), .Z(n3273));
Q_MX02 U5606 ( .S(shiftCount[5]), .A0(xdata[225]), .A1(xdata[193]), .Z(n3272));
Q_MX02 U5607 ( .S(shiftCount[5]), .A0(xdata[224]), .A1(xdata[192]), .Z(n3271));
Q_MX02 U5608 ( .S(shiftCount[5]), .A0(xdata[223]), .A1(xdata[191]), .Z(n3270));
Q_MX02 U5609 ( .S(shiftCount[5]), .A0(xdata[222]), .A1(xdata[190]), .Z(n3269));
Q_MX02 U5610 ( .S(shiftCount[5]), .A0(xdata[221]), .A1(xdata[189]), .Z(n3268));
Q_MX02 U5611 ( .S(shiftCount[5]), .A0(xdata[220]), .A1(xdata[188]), .Z(n3267));
Q_MX02 U5612 ( .S(shiftCount[5]), .A0(xdata[219]), .A1(xdata[187]), .Z(n3266));
Q_MX02 U5613 ( .S(shiftCount[5]), .A0(xdata[218]), .A1(xdata[186]), .Z(n3265));
Q_MX02 U5614 ( .S(shiftCount[5]), .A0(xdata[217]), .A1(xdata[185]), .Z(n3264));
Q_MX02 U5615 ( .S(shiftCount[5]), .A0(xdata[216]), .A1(xdata[184]), .Z(n3263));
Q_MX02 U5616 ( .S(shiftCount[5]), .A0(xdata[215]), .A1(xdata[183]), .Z(n3262));
Q_MX02 U5617 ( .S(shiftCount[5]), .A0(xdata[214]), .A1(xdata[182]), .Z(n3261));
Q_MX02 U5618 ( .S(shiftCount[5]), .A0(xdata[213]), .A1(xdata[181]), .Z(n3260));
Q_MX02 U5619 ( .S(shiftCount[5]), .A0(xdata[212]), .A1(xdata[180]), .Z(n3259));
Q_MX02 U5620 ( .S(shiftCount[5]), .A0(xdata[211]), .A1(xdata[179]), .Z(n3258));
Q_MX02 U5621 ( .S(shiftCount[5]), .A0(xdata[210]), .A1(xdata[178]), .Z(n3257));
Q_MX02 U5622 ( .S(shiftCount[5]), .A0(xdata[209]), .A1(xdata[177]), .Z(n3256));
Q_MX02 U5623 ( .S(shiftCount[5]), .A0(xdata[208]), .A1(xdata[176]), .Z(n3255));
Q_MX02 U5624 ( .S(shiftCount[5]), .A0(xdata[207]), .A1(xdata[175]), .Z(n3254));
Q_MX02 U5625 ( .S(shiftCount[5]), .A0(xdata[206]), .A1(xdata[174]), .Z(n3253));
Q_MX02 U5626 ( .S(shiftCount[5]), .A0(xdata[205]), .A1(xdata[173]), .Z(n3252));
Q_MX02 U5627 ( .S(shiftCount[5]), .A0(xdata[204]), .A1(xdata[172]), .Z(n3251));
Q_MX02 U5628 ( .S(shiftCount[5]), .A0(xdata[203]), .A1(xdata[171]), .Z(n3250));
Q_MX02 U5629 ( .S(shiftCount[5]), .A0(xdata[202]), .A1(xdata[170]), .Z(n3249));
Q_MX02 U5630 ( .S(shiftCount[5]), .A0(xdata[201]), .A1(xdata[169]), .Z(n3248));
Q_MX02 U5631 ( .S(shiftCount[5]), .A0(xdata[200]), .A1(xdata[168]), .Z(n3247));
Q_MX02 U5632 ( .S(shiftCount[5]), .A0(xdata[199]), .A1(xdata[167]), .Z(n3246));
Q_MX02 U5633 ( .S(shiftCount[5]), .A0(xdata[198]), .A1(xdata[166]), .Z(n3245));
Q_MX02 U5634 ( .S(shiftCount[5]), .A0(xdata[197]), .A1(xdata[165]), .Z(n3244));
Q_MX02 U5635 ( .S(shiftCount[5]), .A0(xdata[196]), .A1(xdata[164]), .Z(n3243));
Q_MX02 U5636 ( .S(shiftCount[5]), .A0(xdata[195]), .A1(xdata[163]), .Z(n3242));
Q_MX02 U5637 ( .S(shiftCount[5]), .A0(xdata[194]), .A1(xdata[162]), .Z(n3241));
Q_MX02 U5638 ( .S(shiftCount[5]), .A0(xdata[193]), .A1(xdata[161]), .Z(n3240));
Q_MX02 U5639 ( .S(shiftCount[5]), .A0(xdata[192]), .A1(xdata[160]), .Z(n3239));
Q_MX02 U5640 ( .S(shiftCount[5]), .A0(xdata[191]), .A1(xdata[159]), .Z(n3238));
Q_MX02 U5641 ( .S(shiftCount[5]), .A0(xdata[190]), .A1(xdata[158]), .Z(n3237));
Q_MX02 U5642 ( .S(shiftCount[5]), .A0(xdata[189]), .A1(xdata[157]), .Z(n3236));
Q_MX02 U5643 ( .S(shiftCount[5]), .A0(xdata[188]), .A1(xdata[156]), .Z(n3235));
Q_MX02 U5644 ( .S(shiftCount[5]), .A0(xdata[187]), .A1(xdata[155]), .Z(n3234));
Q_MX02 U5645 ( .S(shiftCount[5]), .A0(xdata[186]), .A1(xdata[154]), .Z(n3233));
Q_MX02 U5646 ( .S(shiftCount[5]), .A0(xdata[185]), .A1(xdata[153]), .Z(n3232));
Q_MX02 U5647 ( .S(shiftCount[5]), .A0(xdata[184]), .A1(xdata[152]), .Z(n3231));
Q_MX02 U5648 ( .S(shiftCount[5]), .A0(xdata[183]), .A1(xdata[151]), .Z(n3230));
Q_MX02 U5649 ( .S(shiftCount[5]), .A0(xdata[182]), .A1(xdata[150]), .Z(n3229));
Q_MX02 U5650 ( .S(shiftCount[5]), .A0(xdata[181]), .A1(xdata[149]), .Z(n3228));
Q_MX02 U5651 ( .S(shiftCount[5]), .A0(xdata[180]), .A1(xdata[148]), .Z(n3227));
Q_MX02 U5652 ( .S(shiftCount[5]), .A0(xdata[179]), .A1(xdata[147]), .Z(n3226));
Q_MX02 U5653 ( .S(shiftCount[5]), .A0(xdata[178]), .A1(xdata[146]), .Z(n3225));
Q_MX02 U5654 ( .S(shiftCount[5]), .A0(xdata[177]), .A1(xdata[145]), .Z(n3224));
Q_MX02 U5655 ( .S(shiftCount[5]), .A0(xdata[176]), .A1(xdata[144]), .Z(n3223));
Q_MX02 U5656 ( .S(shiftCount[5]), .A0(xdata[175]), .A1(xdata[143]), .Z(n3222));
Q_MX02 U5657 ( .S(shiftCount[5]), .A0(xdata[174]), .A1(xdata[142]), .Z(n3221));
Q_MX02 U5658 ( .S(shiftCount[5]), .A0(xdata[173]), .A1(xdata[141]), .Z(n3220));
Q_MX02 U5659 ( .S(shiftCount[5]), .A0(xdata[172]), .A1(xdata[140]), .Z(n3219));
Q_MX02 U5660 ( .S(shiftCount[5]), .A0(xdata[171]), .A1(xdata[139]), .Z(n3218));
Q_MX02 U5661 ( .S(shiftCount[5]), .A0(xdata[170]), .A1(xdata[138]), .Z(n3217));
Q_MX02 U5662 ( .S(shiftCount[5]), .A0(xdata[169]), .A1(xdata[137]), .Z(n3216));
Q_MX02 U5663 ( .S(shiftCount[5]), .A0(xdata[168]), .A1(xdata[136]), .Z(n3215));
Q_MX02 U5664 ( .S(shiftCount[5]), .A0(xdata[167]), .A1(xdata[135]), .Z(n3214));
Q_MX02 U5665 ( .S(shiftCount[5]), .A0(xdata[166]), .A1(xdata[134]), .Z(n3213));
Q_MX02 U5666 ( .S(shiftCount[5]), .A0(xdata[165]), .A1(xdata[133]), .Z(n3212));
Q_MX02 U5667 ( .S(shiftCount[5]), .A0(xdata[164]), .A1(xdata[132]), .Z(n3211));
Q_MX02 U5668 ( .S(shiftCount[5]), .A0(xdata[163]), .A1(xdata[131]), .Z(n3210));
Q_MX02 U5669 ( .S(shiftCount[5]), .A0(xdata[162]), .A1(xdata[130]), .Z(n3209));
Q_MX02 U5670 ( .S(shiftCount[5]), .A0(xdata[161]), .A1(xdata[129]), .Z(n3208));
Q_MX02 U5671 ( .S(shiftCount[5]), .A0(xdata[160]), .A1(xdata[128]), .Z(n3207));
Q_MX02 U5672 ( .S(shiftCount[5]), .A0(xdata[159]), .A1(xdata[127]), .Z(n3206));
Q_MX02 U5673 ( .S(shiftCount[5]), .A0(xdata[158]), .A1(xdata[126]), .Z(n3205));
Q_MX02 U5674 ( .S(shiftCount[5]), .A0(xdata[157]), .A1(xdata[125]), .Z(n3204));
Q_MX02 U5675 ( .S(shiftCount[5]), .A0(xdata[156]), .A1(xdata[124]), .Z(n3203));
Q_MX02 U5676 ( .S(shiftCount[5]), .A0(xdata[155]), .A1(xdata[123]), .Z(n3202));
Q_MX02 U5677 ( .S(shiftCount[5]), .A0(xdata[154]), .A1(xdata[122]), .Z(n3201));
Q_MX02 U5678 ( .S(shiftCount[5]), .A0(xdata[153]), .A1(xdata[121]), .Z(n3200));
Q_MX02 U5679 ( .S(shiftCount[5]), .A0(xdata[152]), .A1(xdata[120]), .Z(n3199));
Q_MX02 U5680 ( .S(shiftCount[5]), .A0(xdata[151]), .A1(xdata[119]), .Z(n3198));
Q_MX02 U5681 ( .S(shiftCount[5]), .A0(xdata[150]), .A1(xdata[118]), .Z(n3197));
Q_MX02 U5682 ( .S(shiftCount[5]), .A0(xdata[149]), .A1(xdata[117]), .Z(n3196));
Q_MX02 U5683 ( .S(shiftCount[5]), .A0(xdata[148]), .A1(xdata[116]), .Z(n3195));
Q_MX02 U5684 ( .S(shiftCount[5]), .A0(xdata[147]), .A1(xdata[115]), .Z(n3194));
Q_MX02 U5685 ( .S(shiftCount[5]), .A0(xdata[146]), .A1(xdata[114]), .Z(n3193));
Q_MX02 U5686 ( .S(shiftCount[5]), .A0(xdata[145]), .A1(xdata[113]), .Z(n3192));
Q_MX02 U5687 ( .S(shiftCount[5]), .A0(xdata[144]), .A1(xdata[112]), .Z(n3191));
Q_MX02 U5688 ( .S(shiftCount[5]), .A0(xdata[143]), .A1(xdata[111]), .Z(n3190));
Q_MX02 U5689 ( .S(shiftCount[5]), .A0(xdata[142]), .A1(xdata[110]), .Z(n3189));
Q_MX02 U5690 ( .S(shiftCount[5]), .A0(xdata[141]), .A1(xdata[109]), .Z(n3188));
Q_MX02 U5691 ( .S(shiftCount[5]), .A0(xdata[140]), .A1(xdata[108]), .Z(n3187));
Q_MX02 U5692 ( .S(shiftCount[5]), .A0(xdata[139]), .A1(xdata[107]), .Z(n3186));
Q_MX02 U5693 ( .S(shiftCount[5]), .A0(xdata[138]), .A1(xdata[106]), .Z(n3185));
Q_MX02 U5694 ( .S(shiftCount[5]), .A0(xdata[137]), .A1(xdata[105]), .Z(n3184));
Q_MX02 U5695 ( .S(shiftCount[5]), .A0(xdata[136]), .A1(xdata[104]), .Z(n3183));
Q_MX02 U5696 ( .S(shiftCount[5]), .A0(xdata[135]), .A1(xdata[103]), .Z(n3182));
Q_MX02 U5697 ( .S(shiftCount[5]), .A0(xdata[134]), .A1(xdata[102]), .Z(n3181));
Q_MX02 U5698 ( .S(shiftCount[5]), .A0(xdata[133]), .A1(xdata[101]), .Z(n3180));
Q_MX02 U5699 ( .S(shiftCount[5]), .A0(xdata[132]), .A1(xdata[100]), .Z(n3179));
Q_MX02 U5700 ( .S(shiftCount[5]), .A0(xdata[131]), .A1(xdata[99]), .Z(n3178));
Q_MX02 U5701 ( .S(shiftCount[5]), .A0(xdata[130]), .A1(xdata[98]), .Z(n3177));
Q_MX02 U5702 ( .S(shiftCount[5]), .A0(xdata[129]), .A1(xdata[97]), .Z(n3176));
Q_MX02 U5703 ( .S(shiftCount[5]), .A0(xdata[128]), .A1(xdata[96]), .Z(n3175));
Q_MX02 U5704 ( .S(shiftCount[5]), .A0(xdata[127]), .A1(xdata[95]), .Z(n3174));
Q_MX02 U5705 ( .S(shiftCount[5]), .A0(xdata[126]), .A1(xdata[94]), .Z(n3173));
Q_MX02 U5706 ( .S(shiftCount[5]), .A0(xdata[125]), .A1(xdata[93]), .Z(n3172));
Q_MX02 U5707 ( .S(shiftCount[5]), .A0(xdata[124]), .A1(xdata[92]), .Z(n3171));
Q_MX02 U5708 ( .S(shiftCount[5]), .A0(xdata[123]), .A1(xdata[91]), .Z(n3170));
Q_MX02 U5709 ( .S(shiftCount[5]), .A0(xdata[122]), .A1(xdata[90]), .Z(n3169));
Q_MX02 U5710 ( .S(shiftCount[5]), .A0(xdata[121]), .A1(xdata[89]), .Z(n3168));
Q_MX02 U5711 ( .S(shiftCount[5]), .A0(xdata[120]), .A1(xdata[88]), .Z(n3167));
Q_MX02 U5712 ( .S(shiftCount[5]), .A0(xdata[119]), .A1(xdata[87]), .Z(n3166));
Q_MX02 U5713 ( .S(shiftCount[5]), .A0(xdata[118]), .A1(xdata[86]), .Z(n3165));
Q_MX02 U5714 ( .S(shiftCount[5]), .A0(xdata[117]), .A1(xdata[85]), .Z(n3164));
Q_MX02 U5715 ( .S(shiftCount[5]), .A0(xdata[116]), .A1(xdata[84]), .Z(n3163));
Q_MX02 U5716 ( .S(shiftCount[5]), .A0(xdata[115]), .A1(xdata[83]), .Z(n3162));
Q_MX02 U5717 ( .S(shiftCount[5]), .A0(xdata[114]), .A1(xdata[82]), .Z(n3161));
Q_MX02 U5718 ( .S(shiftCount[5]), .A0(xdata[113]), .A1(xdata[81]), .Z(n3160));
Q_MX02 U5719 ( .S(shiftCount[5]), .A0(xdata[112]), .A1(xdata[80]), .Z(n3159));
Q_MX02 U5720 ( .S(shiftCount[5]), .A0(xdata[111]), .A1(xdata[79]), .Z(n3158));
Q_MX02 U5721 ( .S(shiftCount[5]), .A0(xdata[110]), .A1(xdata[78]), .Z(n3157));
Q_MX02 U5722 ( .S(shiftCount[5]), .A0(xdata[109]), .A1(xdata[77]), .Z(n3156));
Q_MX02 U5723 ( .S(shiftCount[5]), .A0(xdata[108]), .A1(xdata[76]), .Z(n3155));
Q_MX02 U5724 ( .S(shiftCount[5]), .A0(xdata[107]), .A1(xdata[75]), .Z(n3154));
Q_MX02 U5725 ( .S(shiftCount[5]), .A0(xdata[106]), .A1(xdata[74]), .Z(n3153));
Q_MX02 U5726 ( .S(shiftCount[5]), .A0(xdata[105]), .A1(xdata[73]), .Z(n3152));
Q_MX02 U5727 ( .S(shiftCount[5]), .A0(xdata[104]), .A1(xdata[72]), .Z(n3151));
Q_MX02 U5728 ( .S(shiftCount[5]), .A0(xdata[103]), .A1(xdata[71]), .Z(n3150));
Q_MX02 U5729 ( .S(shiftCount[5]), .A0(xdata[102]), .A1(xdata[70]), .Z(n3149));
Q_MX02 U5730 ( .S(shiftCount[5]), .A0(xdata[101]), .A1(xdata[69]), .Z(n3148));
Q_MX02 U5731 ( .S(shiftCount[5]), .A0(xdata[100]), .A1(xdata[68]), .Z(n3147));
Q_MX02 U5732 ( .S(shiftCount[5]), .A0(xdata[99]), .A1(xdata[67]), .Z(n3146));
Q_MX02 U5733 ( .S(shiftCount[5]), .A0(xdata[98]), .A1(xdata[66]), .Z(n3145));
Q_MX02 U5734 ( .S(shiftCount[5]), .A0(xdata[97]), .A1(xdata[65]), .Z(n3144));
Q_MX02 U5735 ( .S(shiftCount[5]), .A0(xdata[96]), .A1(xdata[64]), .Z(n3143));
Q_MX02 U5736 ( .S(shiftCount[5]), .A0(xdata[95]), .A1(xdata[63]), .Z(n3142));
Q_MX02 U5737 ( .S(shiftCount[5]), .A0(xdata[94]), .A1(xdata[62]), .Z(n3141));
Q_MX02 U5738 ( .S(shiftCount[5]), .A0(xdata[93]), .A1(xdata[61]), .Z(n3140));
Q_MX02 U5739 ( .S(shiftCount[5]), .A0(xdata[92]), .A1(xdata[60]), .Z(n3139));
Q_MX02 U5740 ( .S(shiftCount[5]), .A0(xdata[91]), .A1(xdata[59]), .Z(n3138));
Q_MX02 U5741 ( .S(shiftCount[5]), .A0(xdata[90]), .A1(xdata[58]), .Z(n3137));
Q_MX02 U5742 ( .S(shiftCount[5]), .A0(xdata[89]), .A1(xdata[57]), .Z(n3136));
Q_MX02 U5743 ( .S(shiftCount[5]), .A0(xdata[88]), .A1(xdata[56]), .Z(n3135));
Q_MX02 U5744 ( .S(shiftCount[5]), .A0(xdata[87]), .A1(xdata[55]), .Z(n3134));
Q_MX02 U5745 ( .S(shiftCount[5]), .A0(xdata[86]), .A1(xdata[54]), .Z(n3133));
Q_MX02 U5746 ( .S(shiftCount[5]), .A0(xdata[85]), .A1(xdata[53]), .Z(n3132));
Q_MX02 U5747 ( .S(shiftCount[5]), .A0(xdata[84]), .A1(xdata[52]), .Z(n3131));
Q_MX02 U5748 ( .S(shiftCount[5]), .A0(xdata[83]), .A1(xdata[51]), .Z(n3130));
Q_MX02 U5749 ( .S(shiftCount[5]), .A0(xdata[82]), .A1(xdata[50]), .Z(n3129));
Q_MX02 U5750 ( .S(shiftCount[5]), .A0(xdata[81]), .A1(xdata[49]), .Z(n3128));
Q_MX02 U5751 ( .S(shiftCount[5]), .A0(xdata[80]), .A1(xdata[48]), .Z(n3127));
Q_MX02 U5752 ( .S(shiftCount[5]), .A0(xdata[79]), .A1(xdata[47]), .Z(n3126));
Q_MX02 U5753 ( .S(shiftCount[5]), .A0(xdata[78]), .A1(xdata[46]), .Z(n3125));
Q_MX02 U5754 ( .S(shiftCount[5]), .A0(xdata[77]), .A1(xdata[45]), .Z(n3124));
Q_MX02 U5755 ( .S(shiftCount[5]), .A0(xdata[76]), .A1(xdata[44]), .Z(n3123));
Q_MX02 U5756 ( .S(shiftCount[5]), .A0(xdata[75]), .A1(xdata[43]), .Z(n3122));
Q_MX02 U5757 ( .S(shiftCount[5]), .A0(xdata[74]), .A1(xdata[42]), .Z(n3121));
Q_MX02 U5758 ( .S(shiftCount[5]), .A0(xdata[73]), .A1(xdata[41]), .Z(n3120));
Q_MX02 U5759 ( .S(shiftCount[5]), .A0(xdata[72]), .A1(xdata[40]), .Z(n3119));
Q_MX02 U5760 ( .S(shiftCount[5]), .A0(xdata[71]), .A1(xdata[39]), .Z(n3118));
Q_MX02 U5761 ( .S(shiftCount[5]), .A0(xdata[70]), .A1(xdata[38]), .Z(n3117));
Q_MX02 U5762 ( .S(shiftCount[5]), .A0(xdata[69]), .A1(xdata[37]), .Z(n3116));
Q_MX02 U5763 ( .S(shiftCount[5]), .A0(xdata[68]), .A1(xdata[36]), .Z(n3115));
Q_MX02 U5764 ( .S(shiftCount[5]), .A0(xdata[67]), .A1(xdata[35]), .Z(n3114));
Q_MX02 U5765 ( .S(shiftCount[5]), .A0(xdata[66]), .A1(xdata[34]), .Z(n3113));
Q_MX02 U5766 ( .S(shiftCount[5]), .A0(xdata[65]), .A1(xdata[33]), .Z(n3112));
Q_MX02 U5767 ( .S(shiftCount[5]), .A0(xdata[64]), .A1(xdata[32]), .Z(n3111));
Q_MX02 U5768 ( .S(shiftCount[5]), .A0(xdata[63]), .A1(xdata[31]), .Z(n3110));
Q_MX02 U5769 ( .S(shiftCount[5]), .A0(xdata[62]), .A1(xdata[30]), .Z(n3109));
Q_MX02 U5770 ( .S(shiftCount[5]), .A0(xdata[61]), .A1(xdata[29]), .Z(n3108));
Q_MX02 U5771 ( .S(shiftCount[5]), .A0(xdata[60]), .A1(xdata[28]), .Z(n3107));
Q_MX02 U5772 ( .S(shiftCount[5]), .A0(xdata[59]), .A1(xdata[27]), .Z(n3106));
Q_MX02 U5773 ( .S(shiftCount[5]), .A0(xdata[58]), .A1(xdata[26]), .Z(n3105));
Q_MX02 U5774 ( .S(shiftCount[5]), .A0(xdata[57]), .A1(xdata[25]), .Z(n3104));
Q_MX02 U5775 ( .S(shiftCount[5]), .A0(xdata[56]), .A1(xdata[24]), .Z(n3103));
Q_MX02 U5776 ( .S(shiftCount[5]), .A0(xdata[55]), .A1(xdata[23]), .Z(n3102));
Q_MX02 U5777 ( .S(shiftCount[5]), .A0(xdata[54]), .A1(xdata[22]), .Z(n3101));
Q_MX02 U5778 ( .S(shiftCount[5]), .A0(xdata[53]), .A1(xdata[21]), .Z(n3100));
Q_MX02 U5779 ( .S(shiftCount[5]), .A0(xdata[52]), .A1(xdata[20]), .Z(n3099));
Q_MX02 U5780 ( .S(shiftCount[5]), .A0(xdata[51]), .A1(xdata[19]), .Z(n3098));
Q_MX02 U5781 ( .S(shiftCount[5]), .A0(xdata[50]), .A1(xdata[18]), .Z(n3097));
Q_MX02 U5782 ( .S(shiftCount[5]), .A0(xdata[49]), .A1(xdata[17]), .Z(n3096));
Q_MX02 U5783 ( .S(shiftCount[5]), .A0(xdata[48]), .A1(xdata[16]), .Z(n3095));
Q_MX02 U5784 ( .S(shiftCount[5]), .A0(xdata[47]), .A1(xdata[15]), .Z(n3094));
Q_MX02 U5785 ( .S(shiftCount[5]), .A0(xdata[46]), .A1(xdata[14]), .Z(n3093));
Q_MX02 U5786 ( .S(shiftCount[5]), .A0(xdata[45]), .A1(xdata[13]), .Z(n3092));
Q_MX02 U5787 ( .S(shiftCount[5]), .A0(xdata[44]), .A1(xdata[12]), .Z(n3091));
Q_MX02 U5788 ( .S(shiftCount[5]), .A0(xdata[43]), .A1(xdata[11]), .Z(n3090));
Q_MX02 U5789 ( .S(shiftCount[5]), .A0(xdata[42]), .A1(xdata[10]), .Z(n3089));
Q_MX02 U5790 ( .S(shiftCount[5]), .A0(xdata[41]), .A1(xdata[9]), .Z(n3088));
Q_MX02 U5791 ( .S(shiftCount[5]), .A0(xdata[40]), .A1(xdata[8]), .Z(n3087));
Q_MX02 U5792 ( .S(shiftCount[5]), .A0(xdata[39]), .A1(xdata[7]), .Z(n3086));
Q_MX02 U5793 ( .S(shiftCount[5]), .A0(xdata[38]), .A1(xdata[6]), .Z(n3085));
Q_MX02 U5794 ( .S(shiftCount[5]), .A0(xdata[37]), .A1(xdata[5]), .Z(n3084));
Q_MX02 U5795 ( .S(shiftCount[5]), .A0(xdata[36]), .A1(xdata[4]), .Z(n3083));
Q_MX02 U5796 ( .S(shiftCount[5]), .A0(xdata[35]), .A1(xdata[3]), .Z(n3082));
Q_MX02 U5797 ( .S(shiftCount[5]), .A0(xdata[34]), .A1(xdata[2]), .Z(n3081));
Q_MX02 U5798 ( .S(shiftCount[5]), .A0(xdata[33]), .A1(xdata[1]), .Z(n3080));
Q_MX02 U5799 ( .S(shiftCount[5]), .A0(xdata[32]), .A1(xdata[0]), .Z(n3079));
Q_INV U5800 ( .A(shiftCount[5]), .Z(n3078));
Q_AN02 U5801 ( .A0(n3078), .A1(xdata[31]), .Z(n3077));
Q_AN02 U5802 ( .A0(n3078), .A1(xdata[30]), .Z(n3076));
Q_AN02 U5803 ( .A0(n3078), .A1(xdata[29]), .Z(n3075));
Q_AN02 U5804 ( .A0(n3078), .A1(xdata[28]), .Z(n3074));
Q_AN02 U5805 ( .A0(n3078), .A1(xdata[27]), .Z(n3073));
Q_AN02 U5806 ( .A0(n3078), .A1(xdata[26]), .Z(n3072));
Q_AN02 U5807 ( .A0(n3078), .A1(xdata[25]), .Z(n3071));
Q_AN02 U5808 ( .A0(n3078), .A1(xdata[24]), .Z(n3070));
Q_AN02 U5809 ( .A0(n3078), .A1(xdata[23]), .Z(n3069));
Q_AN02 U5810 ( .A0(n3078), .A1(xdata[22]), .Z(n3068));
Q_AN02 U5811 ( .A0(n3078), .A1(xdata[21]), .Z(n3067));
Q_AN02 U5812 ( .A0(n3078), .A1(xdata[20]), .Z(n3066));
Q_AN02 U5813 ( .A0(n3078), .A1(xdata[19]), .Z(n3065));
Q_AN02 U5814 ( .A0(n3078), .A1(xdata[18]), .Z(n3064));
Q_AN02 U5815 ( .A0(n3078), .A1(xdata[17]), .Z(n3063));
Q_AN02 U5816 ( .A0(n3078), .A1(xdata[16]), .Z(n3062));
Q_AN02 U5817 ( .A0(n3078), .A1(xdata[15]), .Z(n3061));
Q_AN02 U5818 ( .A0(n3078), .A1(xdata[14]), .Z(n3060));
Q_AN02 U5819 ( .A0(n3078), .A1(xdata[13]), .Z(n3059));
Q_AN02 U5820 ( .A0(n3078), .A1(xdata[12]), .Z(n3058));
Q_AN02 U5821 ( .A0(n3078), .A1(xdata[11]), .Z(n3057));
Q_AN02 U5822 ( .A0(n3078), .A1(xdata[10]), .Z(n3056));
Q_AN02 U5823 ( .A0(n3078), .A1(xdata[9]), .Z(n3055));
Q_AN02 U5824 ( .A0(n3078), .A1(xdata[8]), .Z(n3054));
Q_AN02 U5825 ( .A0(n3078), .A1(xdata[7]), .Z(n3053));
Q_AN02 U5826 ( .A0(n3078), .A1(xdata[6]), .Z(n3052));
Q_AN02 U5827 ( .A0(n3078), .A1(xdata[5]), .Z(n3051));
Q_AN02 U5828 ( .A0(n3078), .A1(xdata[4]), .Z(n3050));
Q_AN02 U5829 ( .A0(n3078), .A1(xdata[3]), .Z(n3049));
Q_AN02 U5830 ( .A0(n3078), .A1(xdata[2]), .Z(n3048));
Q_AN02 U5831 ( .A0(n3078), .A1(xdata[1]), .Z(n3047));
Q_AN02 U5832 ( .A0(n3078), .A1(xdata[0]), .Z(n3046));
Q_AN02 U5833 ( .A0(shiftCount[6]), .A1(n3622), .Z(n3045));
Q_AN02 U5834 ( .A0(shiftCount[6]), .A1(n3621), .Z(n3044));
Q_AN02 U5835 ( .A0(shiftCount[6]), .A1(n3620), .Z(n3043));
Q_AN02 U5836 ( .A0(shiftCount[6]), .A1(n3619), .Z(n3042));
Q_AN02 U5837 ( .A0(shiftCount[6]), .A1(n3618), .Z(n3041));
Q_AN02 U5838 ( .A0(shiftCount[6]), .A1(n3617), .Z(n3040));
Q_AN02 U5839 ( .A0(shiftCount[6]), .A1(n3616), .Z(n3039));
Q_AN02 U5840 ( .A0(shiftCount[6]), .A1(n3615), .Z(n3038));
Q_AN02 U5841 ( .A0(shiftCount[6]), .A1(n3614), .Z(n3037));
Q_AN02 U5842 ( .A0(shiftCount[6]), .A1(n3613), .Z(n3036));
Q_AN02 U5843 ( .A0(shiftCount[6]), .A1(n3612), .Z(n3035));
Q_AN02 U5844 ( .A0(shiftCount[6]), .A1(n3611), .Z(n3034));
Q_AN02 U5845 ( .A0(shiftCount[6]), .A1(n3610), .Z(n3033));
Q_AN02 U5846 ( .A0(shiftCount[6]), .A1(n3609), .Z(n3032));
Q_AN02 U5847 ( .A0(shiftCount[6]), .A1(n3608), .Z(n3031));
Q_AN02 U5848 ( .A0(shiftCount[6]), .A1(n3607), .Z(n3030));
Q_AN02 U5849 ( .A0(shiftCount[6]), .A1(n3606), .Z(n3029));
Q_AN02 U5850 ( .A0(shiftCount[6]), .A1(n3605), .Z(n3028));
Q_AN02 U5851 ( .A0(shiftCount[6]), .A1(n3604), .Z(n3027));
Q_AN02 U5852 ( .A0(shiftCount[6]), .A1(n3603), .Z(n3026));
Q_AN02 U5853 ( .A0(shiftCount[6]), .A1(n3602), .Z(n3025));
Q_AN02 U5854 ( .A0(shiftCount[6]), .A1(n3601), .Z(n3024));
Q_AN02 U5855 ( .A0(shiftCount[6]), .A1(n3600), .Z(n3023));
Q_AN02 U5856 ( .A0(shiftCount[6]), .A1(n3599), .Z(n3022));
Q_AN02 U5857 ( .A0(shiftCount[6]), .A1(n3598), .Z(n3021));
Q_AN02 U5858 ( .A0(shiftCount[6]), .A1(n3597), .Z(n3020));
Q_AN02 U5859 ( .A0(shiftCount[6]), .A1(n3596), .Z(n3019));
Q_AN02 U5860 ( .A0(shiftCount[6]), .A1(n3595), .Z(n3018));
Q_AN02 U5861 ( .A0(shiftCount[6]), .A1(n3594), .Z(n3017));
Q_AN02 U5862 ( .A0(shiftCount[6]), .A1(n3593), .Z(n3016));
Q_AN02 U5863 ( .A0(shiftCount[6]), .A1(n3592), .Z(n3015));
Q_AN02 U5864 ( .A0(shiftCount[6]), .A1(n3591), .Z(n3014));
Q_AN02 U5865 ( .A0(shiftCount[6]), .A1(n3590), .Z(n3013));
Q_AN02 U5866 ( .A0(shiftCount[6]), .A1(n3589), .Z(n3012));
Q_AN02 U5867 ( .A0(shiftCount[6]), .A1(n3588), .Z(n3011));
Q_AN02 U5868 ( .A0(shiftCount[6]), .A1(n3587), .Z(n3010));
Q_AN02 U5869 ( .A0(shiftCount[6]), .A1(n3586), .Z(n3009));
Q_AN02 U5870 ( .A0(shiftCount[6]), .A1(n3585), .Z(n3008));
Q_AN02 U5871 ( .A0(shiftCount[6]), .A1(n3584), .Z(n3007));
Q_AN02 U5872 ( .A0(shiftCount[6]), .A1(n3583), .Z(n3006));
Q_AN02 U5873 ( .A0(shiftCount[6]), .A1(n3582), .Z(n3005));
Q_AN02 U5874 ( .A0(shiftCount[6]), .A1(n3581), .Z(n3004));
Q_AN02 U5875 ( .A0(shiftCount[6]), .A1(n3580), .Z(n3003));
Q_AN02 U5876 ( .A0(shiftCount[6]), .A1(n3579), .Z(n3002));
Q_AN02 U5877 ( .A0(shiftCount[6]), .A1(n3578), .Z(n3001));
Q_AN02 U5878 ( .A0(shiftCount[6]), .A1(n3577), .Z(n3000));
Q_AN02 U5879 ( .A0(shiftCount[6]), .A1(n3576), .Z(n2999));
Q_AN02 U5880 ( .A0(shiftCount[6]), .A1(n3575), .Z(n2998));
Q_AN02 U5881 ( .A0(shiftCount[6]), .A1(n3574), .Z(n2997));
Q_AN02 U5882 ( .A0(shiftCount[6]), .A1(n3573), .Z(n2996));
Q_AN02 U5883 ( .A0(shiftCount[6]), .A1(n3572), .Z(n2995));
Q_AN02 U5884 ( .A0(shiftCount[6]), .A1(n3571), .Z(n2994));
Q_AN02 U5885 ( .A0(shiftCount[6]), .A1(n3570), .Z(n2993));
Q_AN02 U5886 ( .A0(shiftCount[6]), .A1(n3569), .Z(n2992));
Q_AN02 U5887 ( .A0(shiftCount[6]), .A1(n3568), .Z(n2991));
Q_AN02 U5888 ( .A0(shiftCount[6]), .A1(n3567), .Z(n2990));
Q_AN02 U5889 ( .A0(shiftCount[6]), .A1(n3566), .Z(n2989));
Q_AN02 U5890 ( .A0(shiftCount[6]), .A1(n3565), .Z(n2988));
Q_AN02 U5891 ( .A0(shiftCount[6]), .A1(n3564), .Z(n2987));
Q_AN02 U5892 ( .A0(shiftCount[6]), .A1(n3563), .Z(n2986));
Q_AN02 U5893 ( .A0(shiftCount[6]), .A1(n3562), .Z(n2985));
Q_AN02 U5894 ( .A0(shiftCount[6]), .A1(n3561), .Z(n2984));
Q_AN02 U5895 ( .A0(shiftCount[6]), .A1(n3560), .Z(n2983));
Q_AN02 U5896 ( .A0(shiftCount[6]), .A1(n3559), .Z(n2982));
Q_MX02 U5897 ( .S(shiftCount[6]), .A0(n3622), .A1(n3558), .Z(n2981));
Q_MX02 U5898 ( .S(shiftCount[6]), .A0(n3621), .A1(n3557), .Z(n2980));
Q_MX02 U5899 ( .S(shiftCount[6]), .A0(n3620), .A1(n3556), .Z(n2979));
Q_MX02 U5900 ( .S(shiftCount[6]), .A0(n3619), .A1(n3555), .Z(n2978));
Q_MX02 U5901 ( .S(shiftCount[6]), .A0(n3618), .A1(n3554), .Z(n2977));
Q_MX02 U5902 ( .S(shiftCount[6]), .A0(n3617), .A1(n3553), .Z(n2976));
Q_MX02 U5903 ( .S(shiftCount[6]), .A0(n3616), .A1(n3552), .Z(n2975));
Q_MX02 U5904 ( .S(shiftCount[6]), .A0(n3615), .A1(n3551), .Z(n2974));
Q_MX02 U5905 ( .S(shiftCount[6]), .A0(n3614), .A1(n3550), .Z(n2973));
Q_MX02 U5906 ( .S(shiftCount[6]), .A0(n3613), .A1(n3549), .Z(n2972));
Q_MX02 U5907 ( .S(shiftCount[6]), .A0(n3612), .A1(n3548), .Z(n2971));
Q_MX02 U5908 ( .S(shiftCount[6]), .A0(n3611), .A1(n3547), .Z(n2970));
Q_MX02 U5909 ( .S(shiftCount[6]), .A0(n3610), .A1(n3546), .Z(n2969));
Q_MX02 U5910 ( .S(shiftCount[6]), .A0(n3609), .A1(n3545), .Z(n2968));
Q_MX02 U5911 ( .S(shiftCount[6]), .A0(n3608), .A1(n3544), .Z(n2967));
Q_MX02 U5912 ( .S(shiftCount[6]), .A0(n3607), .A1(n3543), .Z(n2966));
Q_MX02 U5913 ( .S(shiftCount[6]), .A0(n3606), .A1(n3542), .Z(n2965));
Q_MX02 U5914 ( .S(shiftCount[6]), .A0(n3605), .A1(n3541), .Z(n2964));
Q_MX02 U5915 ( .S(shiftCount[6]), .A0(n3604), .A1(n3540), .Z(n2963));
Q_MX02 U5916 ( .S(shiftCount[6]), .A0(n3603), .A1(n3539), .Z(n2962));
Q_MX02 U5917 ( .S(shiftCount[6]), .A0(n3602), .A1(n3538), .Z(n2961));
Q_MX02 U5918 ( .S(shiftCount[6]), .A0(n3601), .A1(n3537), .Z(n2960));
Q_MX02 U5919 ( .S(shiftCount[6]), .A0(n3600), .A1(n3536), .Z(n2959));
Q_MX02 U5920 ( .S(shiftCount[6]), .A0(n3599), .A1(n3535), .Z(n2958));
Q_MX02 U5921 ( .S(shiftCount[6]), .A0(n3598), .A1(n3534), .Z(n2957));
Q_MX02 U5922 ( .S(shiftCount[6]), .A0(n3597), .A1(n3533), .Z(n2956));
Q_MX02 U5923 ( .S(shiftCount[6]), .A0(n3596), .A1(n3532), .Z(n2955));
Q_MX02 U5924 ( .S(shiftCount[6]), .A0(n3595), .A1(n3531), .Z(n2954));
Q_MX02 U5925 ( .S(shiftCount[6]), .A0(n3594), .A1(n3530), .Z(n2953));
Q_MX02 U5926 ( .S(shiftCount[6]), .A0(n3593), .A1(n3529), .Z(n2952));
Q_MX02 U5927 ( .S(shiftCount[6]), .A0(n3592), .A1(n3528), .Z(n2951));
Q_MX02 U5928 ( .S(shiftCount[6]), .A0(n3591), .A1(n3527), .Z(n2950));
Q_MX02 U5929 ( .S(shiftCount[6]), .A0(n3590), .A1(n3526), .Z(n2949));
Q_MX02 U5930 ( .S(shiftCount[6]), .A0(n3589), .A1(n3525), .Z(n2948));
Q_MX02 U5931 ( .S(shiftCount[6]), .A0(n3588), .A1(n3524), .Z(n2947));
Q_MX02 U5932 ( .S(shiftCount[6]), .A0(n3587), .A1(n3523), .Z(n2946));
Q_MX02 U5933 ( .S(shiftCount[6]), .A0(n3586), .A1(n3522), .Z(n2945));
Q_MX02 U5934 ( .S(shiftCount[6]), .A0(n3585), .A1(n3521), .Z(n2944));
Q_MX02 U5935 ( .S(shiftCount[6]), .A0(n3584), .A1(n3520), .Z(n2943));
Q_MX02 U5936 ( .S(shiftCount[6]), .A0(n3583), .A1(n3519), .Z(n2942));
Q_MX02 U5937 ( .S(shiftCount[6]), .A0(n3582), .A1(n3518), .Z(n2941));
Q_MX02 U5938 ( .S(shiftCount[6]), .A0(n3581), .A1(n3517), .Z(n2940));
Q_MX02 U5939 ( .S(shiftCount[6]), .A0(n3580), .A1(n3516), .Z(n2939));
Q_MX02 U5940 ( .S(shiftCount[6]), .A0(n3579), .A1(n3515), .Z(n2938));
Q_MX02 U5941 ( .S(shiftCount[6]), .A0(n3578), .A1(n3514), .Z(n2937));
Q_MX02 U5942 ( .S(shiftCount[6]), .A0(n3577), .A1(n3513), .Z(n2936));
Q_MX02 U5943 ( .S(shiftCount[6]), .A0(n3576), .A1(n3512), .Z(n2935));
Q_MX02 U5944 ( .S(shiftCount[6]), .A0(n3575), .A1(n3511), .Z(n2934));
Q_MX02 U5945 ( .S(shiftCount[6]), .A0(n3574), .A1(n3510), .Z(n2933));
Q_MX02 U5946 ( .S(shiftCount[6]), .A0(n3573), .A1(n3509), .Z(n2932));
Q_MX02 U5947 ( .S(shiftCount[6]), .A0(n3572), .A1(n3508), .Z(n2931));
Q_MX02 U5948 ( .S(shiftCount[6]), .A0(n3571), .A1(n3507), .Z(n2930));
Q_MX02 U5949 ( .S(shiftCount[6]), .A0(n3570), .A1(n3506), .Z(n2929));
Q_MX02 U5950 ( .S(shiftCount[6]), .A0(n3569), .A1(n3505), .Z(n2928));
Q_MX02 U5951 ( .S(shiftCount[6]), .A0(n3568), .A1(n3504), .Z(n2927));
Q_MX02 U5952 ( .S(shiftCount[6]), .A0(n3567), .A1(n3503), .Z(n2926));
Q_MX02 U5953 ( .S(shiftCount[6]), .A0(n3566), .A1(n3502), .Z(n2925));
Q_MX02 U5954 ( .S(shiftCount[6]), .A0(n3565), .A1(n3501), .Z(n2924));
Q_MX02 U5955 ( .S(shiftCount[6]), .A0(n3564), .A1(n3500), .Z(n2923));
Q_MX02 U5956 ( .S(shiftCount[6]), .A0(n3563), .A1(n3499), .Z(n2922));
Q_MX02 U5957 ( .S(shiftCount[6]), .A0(n3562), .A1(n3498), .Z(n2921));
Q_MX02 U5958 ( .S(shiftCount[6]), .A0(n3561), .A1(n3497), .Z(n2920));
Q_MX02 U5959 ( .S(shiftCount[6]), .A0(n3560), .A1(n3496), .Z(n2919));
Q_MX02 U5960 ( .S(shiftCount[6]), .A0(n3559), .A1(n3495), .Z(n2918));
Q_MX02 U5961 ( .S(shiftCount[6]), .A0(n3558), .A1(n3494), .Z(n2917));
Q_MX02 U5962 ( .S(shiftCount[6]), .A0(n3557), .A1(n3493), .Z(n2916));
Q_MX02 U5963 ( .S(shiftCount[6]), .A0(n3556), .A1(n3492), .Z(n2915));
Q_MX02 U5964 ( .S(shiftCount[6]), .A0(n3555), .A1(n3491), .Z(n2914));
Q_MX02 U5965 ( .S(shiftCount[6]), .A0(n3554), .A1(n3490), .Z(n2913));
Q_MX02 U5966 ( .S(shiftCount[6]), .A0(n3553), .A1(n3489), .Z(n2912));
Q_MX02 U5967 ( .S(shiftCount[6]), .A0(n3552), .A1(n3488), .Z(n2911));
Q_MX02 U5968 ( .S(shiftCount[6]), .A0(n3551), .A1(n3487), .Z(n2910));
Q_MX02 U5969 ( .S(shiftCount[6]), .A0(n3550), .A1(n3486), .Z(n2909));
Q_MX02 U5970 ( .S(shiftCount[6]), .A0(n3549), .A1(n3485), .Z(n2908));
Q_MX02 U5971 ( .S(shiftCount[6]), .A0(n3548), .A1(n3484), .Z(n2907));
Q_MX02 U5972 ( .S(shiftCount[6]), .A0(n3547), .A1(n3483), .Z(n2906));
Q_MX02 U5973 ( .S(shiftCount[6]), .A0(n3546), .A1(n3482), .Z(n2905));
Q_MX02 U5974 ( .S(shiftCount[6]), .A0(n3545), .A1(n3481), .Z(n2904));
Q_MX02 U5975 ( .S(shiftCount[6]), .A0(n3544), .A1(n3480), .Z(n2903));
Q_MX02 U5976 ( .S(shiftCount[6]), .A0(n3543), .A1(n3479), .Z(n2902));
Q_MX02 U5977 ( .S(shiftCount[6]), .A0(n3542), .A1(n3478), .Z(n2901));
Q_MX02 U5978 ( .S(shiftCount[6]), .A0(n3541), .A1(n3477), .Z(n2900));
Q_MX02 U5979 ( .S(shiftCount[6]), .A0(n3540), .A1(n3476), .Z(n2899));
Q_MX02 U5980 ( .S(shiftCount[6]), .A0(n3539), .A1(n3475), .Z(n2898));
Q_MX02 U5981 ( .S(shiftCount[6]), .A0(n3538), .A1(n3474), .Z(n2897));
Q_MX02 U5982 ( .S(shiftCount[6]), .A0(n3537), .A1(n3473), .Z(n2896));
Q_MX02 U5983 ( .S(shiftCount[6]), .A0(n3536), .A1(n3472), .Z(n2895));
Q_MX02 U5984 ( .S(shiftCount[6]), .A0(n3535), .A1(n3471), .Z(n2894));
Q_MX02 U5985 ( .S(shiftCount[6]), .A0(n3534), .A1(n3470), .Z(n2893));
Q_MX02 U5986 ( .S(shiftCount[6]), .A0(n3533), .A1(n3469), .Z(n2892));
Q_MX02 U5987 ( .S(shiftCount[6]), .A0(n3532), .A1(n3468), .Z(n2891));
Q_MX02 U5988 ( .S(shiftCount[6]), .A0(n3531), .A1(n3467), .Z(n2890));
Q_MX02 U5989 ( .S(shiftCount[6]), .A0(n3530), .A1(n3466), .Z(n2889));
Q_MX02 U5990 ( .S(shiftCount[6]), .A0(n3529), .A1(n3465), .Z(n2888));
Q_MX02 U5991 ( .S(shiftCount[6]), .A0(n3528), .A1(n3464), .Z(n2887));
Q_MX02 U5992 ( .S(shiftCount[6]), .A0(n3527), .A1(n3463), .Z(n2886));
Q_MX02 U5993 ( .S(shiftCount[6]), .A0(n3526), .A1(n3462), .Z(n2885));
Q_MX02 U5994 ( .S(shiftCount[6]), .A0(n3525), .A1(n3461), .Z(n2884));
Q_MX02 U5995 ( .S(shiftCount[6]), .A0(n3524), .A1(n3460), .Z(n2883));
Q_MX02 U5996 ( .S(shiftCount[6]), .A0(n3523), .A1(n3459), .Z(n2882));
Q_MX02 U5997 ( .S(shiftCount[6]), .A0(n3522), .A1(n3458), .Z(n2881));
Q_MX02 U5998 ( .S(shiftCount[6]), .A0(n3521), .A1(n3457), .Z(n2880));
Q_MX02 U5999 ( .S(shiftCount[6]), .A0(n3520), .A1(n3456), .Z(n2879));
Q_MX02 U6000 ( .S(shiftCount[6]), .A0(n3519), .A1(n3455), .Z(n2878));
Q_MX02 U6001 ( .S(shiftCount[6]), .A0(n3518), .A1(n3454), .Z(n2877));
Q_MX02 U6002 ( .S(shiftCount[6]), .A0(n3517), .A1(n3453), .Z(n2876));
Q_MX02 U6003 ( .S(shiftCount[6]), .A0(n3516), .A1(n3452), .Z(n2875));
Q_MX02 U6004 ( .S(shiftCount[6]), .A0(n3515), .A1(n3451), .Z(n2874));
Q_MX02 U6005 ( .S(shiftCount[6]), .A0(n3514), .A1(n3450), .Z(n2873));
Q_MX02 U6006 ( .S(shiftCount[6]), .A0(n3513), .A1(n3449), .Z(n2872));
Q_MX02 U6007 ( .S(shiftCount[6]), .A0(n3512), .A1(n3448), .Z(n2871));
Q_MX02 U6008 ( .S(shiftCount[6]), .A0(n3511), .A1(n3447), .Z(n2870));
Q_MX02 U6009 ( .S(shiftCount[6]), .A0(n3510), .A1(n3446), .Z(n2869));
Q_MX02 U6010 ( .S(shiftCount[6]), .A0(n3509), .A1(n3445), .Z(n2868));
Q_MX02 U6011 ( .S(shiftCount[6]), .A0(n3508), .A1(n3444), .Z(n2867));
Q_MX02 U6012 ( .S(shiftCount[6]), .A0(n3507), .A1(n3443), .Z(n2866));
Q_MX02 U6013 ( .S(shiftCount[6]), .A0(n3506), .A1(n3442), .Z(n2865));
Q_MX02 U6014 ( .S(shiftCount[6]), .A0(n3505), .A1(n3441), .Z(n2864));
Q_MX02 U6015 ( .S(shiftCount[6]), .A0(n3504), .A1(n3440), .Z(n2863));
Q_MX02 U6016 ( .S(shiftCount[6]), .A0(n3503), .A1(n3439), .Z(n2862));
Q_MX02 U6017 ( .S(shiftCount[6]), .A0(n3502), .A1(n3438), .Z(n2861));
Q_MX02 U6018 ( .S(shiftCount[6]), .A0(n3501), .A1(n3437), .Z(n2860));
Q_MX02 U6019 ( .S(shiftCount[6]), .A0(n3500), .A1(n3436), .Z(n2859));
Q_MX02 U6020 ( .S(shiftCount[6]), .A0(n3499), .A1(n3435), .Z(n2858));
Q_MX02 U6021 ( .S(shiftCount[6]), .A0(n3498), .A1(n3434), .Z(n2857));
Q_MX02 U6022 ( .S(shiftCount[6]), .A0(n3497), .A1(n3433), .Z(n2856));
Q_MX02 U6023 ( .S(shiftCount[6]), .A0(n3496), .A1(n3432), .Z(n2855));
Q_MX02 U6024 ( .S(shiftCount[6]), .A0(n3495), .A1(n3431), .Z(n2854));
Q_MX02 U6025 ( .S(shiftCount[6]), .A0(n3494), .A1(n3430), .Z(n2853));
Q_MX02 U6026 ( .S(shiftCount[6]), .A0(n3493), .A1(n3429), .Z(n2852));
Q_MX02 U6027 ( .S(shiftCount[6]), .A0(n3492), .A1(n3428), .Z(n2851));
Q_MX02 U6028 ( .S(shiftCount[6]), .A0(n3491), .A1(n3427), .Z(n2850));
Q_MX02 U6029 ( .S(shiftCount[6]), .A0(n3490), .A1(n3426), .Z(n2849));
Q_MX02 U6030 ( .S(shiftCount[6]), .A0(n3489), .A1(n3425), .Z(n2848));
Q_MX02 U6031 ( .S(shiftCount[6]), .A0(n3488), .A1(n3424), .Z(n2847));
Q_MX02 U6032 ( .S(shiftCount[6]), .A0(n3487), .A1(n3423), .Z(n2846));
Q_MX02 U6033 ( .S(shiftCount[6]), .A0(n3486), .A1(n3422), .Z(n2845));
Q_MX02 U6034 ( .S(shiftCount[6]), .A0(n3485), .A1(n3421), .Z(n2844));
Q_MX02 U6035 ( .S(shiftCount[6]), .A0(n3484), .A1(n3420), .Z(n2843));
Q_MX02 U6036 ( .S(shiftCount[6]), .A0(n3483), .A1(n3419), .Z(n2842));
Q_MX02 U6037 ( .S(shiftCount[6]), .A0(n3482), .A1(n3418), .Z(n2841));
Q_MX02 U6038 ( .S(shiftCount[6]), .A0(n3481), .A1(n3417), .Z(n2840));
Q_MX02 U6039 ( .S(shiftCount[6]), .A0(n3480), .A1(n3416), .Z(n2839));
Q_MX02 U6040 ( .S(shiftCount[6]), .A0(n3479), .A1(n3415), .Z(n2838));
Q_MX02 U6041 ( .S(shiftCount[6]), .A0(n3478), .A1(n3414), .Z(n2837));
Q_MX02 U6042 ( .S(shiftCount[6]), .A0(n3477), .A1(n3413), .Z(n2836));
Q_MX02 U6043 ( .S(shiftCount[6]), .A0(n3476), .A1(n3412), .Z(n2835));
Q_MX02 U6044 ( .S(shiftCount[6]), .A0(n3475), .A1(n3411), .Z(n2834));
Q_MX02 U6045 ( .S(shiftCount[6]), .A0(n3474), .A1(n3410), .Z(n2833));
Q_MX02 U6046 ( .S(shiftCount[6]), .A0(n3473), .A1(n3409), .Z(n2832));
Q_MX02 U6047 ( .S(shiftCount[6]), .A0(n3472), .A1(n3408), .Z(n2831));
Q_MX02 U6048 ( .S(shiftCount[6]), .A0(n3471), .A1(n3407), .Z(n2830));
Q_MX02 U6049 ( .S(shiftCount[6]), .A0(n3470), .A1(n3406), .Z(n2829));
Q_MX02 U6050 ( .S(shiftCount[6]), .A0(n3469), .A1(n3405), .Z(n2828));
Q_MX02 U6051 ( .S(shiftCount[6]), .A0(n3468), .A1(n3404), .Z(n2827));
Q_MX02 U6052 ( .S(shiftCount[6]), .A0(n3467), .A1(n3403), .Z(n2826));
Q_MX02 U6053 ( .S(shiftCount[6]), .A0(n3466), .A1(n3402), .Z(n2825));
Q_MX02 U6054 ( .S(shiftCount[6]), .A0(n3465), .A1(n3401), .Z(n2824));
Q_MX02 U6055 ( .S(shiftCount[6]), .A0(n3464), .A1(n3400), .Z(n2823));
Q_MX02 U6056 ( .S(shiftCount[6]), .A0(n3463), .A1(n3399), .Z(n2822));
Q_MX02 U6057 ( .S(shiftCount[6]), .A0(n3462), .A1(n3398), .Z(n2821));
Q_MX02 U6058 ( .S(shiftCount[6]), .A0(n3461), .A1(n3397), .Z(n2820));
Q_MX02 U6059 ( .S(shiftCount[6]), .A0(n3460), .A1(n3396), .Z(n2819));
Q_MX02 U6060 ( .S(shiftCount[6]), .A0(n3459), .A1(n3395), .Z(n2818));
Q_MX02 U6061 ( .S(shiftCount[6]), .A0(n3458), .A1(n3394), .Z(n2817));
Q_MX02 U6062 ( .S(shiftCount[6]), .A0(n3457), .A1(n3393), .Z(n2816));
Q_MX02 U6063 ( .S(shiftCount[6]), .A0(n3456), .A1(n3392), .Z(n2815));
Q_MX02 U6064 ( .S(shiftCount[6]), .A0(n3455), .A1(n3391), .Z(n2814));
Q_MX02 U6065 ( .S(shiftCount[6]), .A0(n3454), .A1(n3390), .Z(n2813));
Q_MX02 U6066 ( .S(shiftCount[6]), .A0(n3453), .A1(n3389), .Z(n2812));
Q_MX02 U6067 ( .S(shiftCount[6]), .A0(n3452), .A1(n3388), .Z(n2811));
Q_MX02 U6068 ( .S(shiftCount[6]), .A0(n3451), .A1(n3387), .Z(n2810));
Q_MX02 U6069 ( .S(shiftCount[6]), .A0(n3450), .A1(n3386), .Z(n2809));
Q_MX02 U6070 ( .S(shiftCount[6]), .A0(n3449), .A1(n3385), .Z(n2808));
Q_MX02 U6071 ( .S(shiftCount[6]), .A0(n3448), .A1(n3384), .Z(n2807));
Q_MX02 U6072 ( .S(shiftCount[6]), .A0(n3447), .A1(n3383), .Z(n2806));
Q_MX02 U6073 ( .S(shiftCount[6]), .A0(n3446), .A1(n3382), .Z(n2805));
Q_MX02 U6074 ( .S(shiftCount[6]), .A0(n3445), .A1(n3381), .Z(n2804));
Q_MX02 U6075 ( .S(shiftCount[6]), .A0(n3444), .A1(n3380), .Z(n2803));
Q_MX02 U6076 ( .S(shiftCount[6]), .A0(n3443), .A1(n3379), .Z(n2802));
Q_MX02 U6077 ( .S(shiftCount[6]), .A0(n3442), .A1(n3378), .Z(n2801));
Q_MX02 U6078 ( .S(shiftCount[6]), .A0(n3441), .A1(n3377), .Z(n2800));
Q_MX02 U6079 ( .S(shiftCount[6]), .A0(n3440), .A1(n3376), .Z(n2799));
Q_MX02 U6080 ( .S(shiftCount[6]), .A0(n3439), .A1(n3375), .Z(n2798));
Q_MX02 U6081 ( .S(shiftCount[6]), .A0(n3438), .A1(n3374), .Z(n2797));
Q_MX02 U6082 ( .S(shiftCount[6]), .A0(n3437), .A1(n3373), .Z(n2796));
Q_MX02 U6083 ( .S(shiftCount[6]), .A0(n3436), .A1(n3372), .Z(n2795));
Q_MX02 U6084 ( .S(shiftCount[6]), .A0(n3435), .A1(n3371), .Z(n2794));
Q_MX02 U6085 ( .S(shiftCount[6]), .A0(n3434), .A1(n3370), .Z(n2793));
Q_MX02 U6086 ( .S(shiftCount[6]), .A0(n3433), .A1(n3369), .Z(n2792));
Q_MX02 U6087 ( .S(shiftCount[6]), .A0(n3432), .A1(n3368), .Z(n2791));
Q_MX02 U6088 ( .S(shiftCount[6]), .A0(n3431), .A1(n3367), .Z(n2790));
Q_MX02 U6089 ( .S(shiftCount[6]), .A0(n3430), .A1(n3366), .Z(n2789));
Q_MX02 U6090 ( .S(shiftCount[6]), .A0(n3429), .A1(n3365), .Z(n2788));
Q_MX02 U6091 ( .S(shiftCount[6]), .A0(n3428), .A1(n3364), .Z(n2787));
Q_MX02 U6092 ( .S(shiftCount[6]), .A0(n3427), .A1(n3363), .Z(n2786));
Q_MX02 U6093 ( .S(shiftCount[6]), .A0(n3426), .A1(n3362), .Z(n2785));
Q_MX02 U6094 ( .S(shiftCount[6]), .A0(n3425), .A1(n3361), .Z(n2784));
Q_MX02 U6095 ( .S(shiftCount[6]), .A0(n3424), .A1(n3360), .Z(n2783));
Q_MX02 U6096 ( .S(shiftCount[6]), .A0(n3423), .A1(n3359), .Z(n2782));
Q_MX02 U6097 ( .S(shiftCount[6]), .A0(n3422), .A1(n3358), .Z(n2781));
Q_MX02 U6098 ( .S(shiftCount[6]), .A0(n3421), .A1(n3357), .Z(n2780));
Q_MX02 U6099 ( .S(shiftCount[6]), .A0(n3420), .A1(n3356), .Z(n2779));
Q_MX02 U6100 ( .S(shiftCount[6]), .A0(n3419), .A1(n3355), .Z(n2778));
Q_MX02 U6101 ( .S(shiftCount[6]), .A0(n3418), .A1(n3354), .Z(n2777));
Q_MX02 U6102 ( .S(shiftCount[6]), .A0(n3417), .A1(n3353), .Z(n2776));
Q_MX02 U6103 ( .S(shiftCount[6]), .A0(n3416), .A1(n3352), .Z(n2775));
Q_MX02 U6104 ( .S(shiftCount[6]), .A0(n3415), .A1(n3351), .Z(n2774));
Q_MX02 U6105 ( .S(shiftCount[6]), .A0(n3414), .A1(n3350), .Z(n2773));
Q_MX02 U6106 ( .S(shiftCount[6]), .A0(n3413), .A1(n3349), .Z(n2772));
Q_MX02 U6107 ( .S(shiftCount[6]), .A0(n3412), .A1(n3348), .Z(n2771));
Q_MX02 U6108 ( .S(shiftCount[6]), .A0(n3411), .A1(n3347), .Z(n2770));
Q_MX02 U6109 ( .S(shiftCount[6]), .A0(n3410), .A1(n3346), .Z(n2769));
Q_MX02 U6110 ( .S(shiftCount[6]), .A0(n3409), .A1(n3345), .Z(n2768));
Q_MX02 U6111 ( .S(shiftCount[6]), .A0(n3408), .A1(n3344), .Z(n2767));
Q_MX02 U6112 ( .S(shiftCount[6]), .A0(n3407), .A1(n3343), .Z(n2766));
Q_MX02 U6113 ( .S(shiftCount[6]), .A0(n3406), .A1(n3342), .Z(n2765));
Q_MX02 U6114 ( .S(shiftCount[6]), .A0(n3405), .A1(n3341), .Z(n2764));
Q_MX02 U6115 ( .S(shiftCount[6]), .A0(n3404), .A1(n3340), .Z(n2763));
Q_MX02 U6116 ( .S(shiftCount[6]), .A0(n3403), .A1(n3339), .Z(n2762));
Q_MX02 U6117 ( .S(shiftCount[6]), .A0(n3402), .A1(n3338), .Z(n2761));
Q_MX02 U6118 ( .S(shiftCount[6]), .A0(n3401), .A1(n3337), .Z(n2760));
Q_MX02 U6119 ( .S(shiftCount[6]), .A0(n3400), .A1(n3336), .Z(n2759));
Q_MX02 U6120 ( .S(shiftCount[6]), .A0(n3399), .A1(n3335), .Z(n2758));
Q_MX02 U6121 ( .S(shiftCount[6]), .A0(n3398), .A1(n3334), .Z(n2757));
Q_MX02 U6122 ( .S(shiftCount[6]), .A0(n3397), .A1(n3333), .Z(n2756));
Q_MX02 U6123 ( .S(shiftCount[6]), .A0(n3396), .A1(n3332), .Z(n2755));
Q_MX02 U6124 ( .S(shiftCount[6]), .A0(n3395), .A1(n3331), .Z(n2754));
Q_MX02 U6125 ( .S(shiftCount[6]), .A0(n3394), .A1(n3330), .Z(n2753));
Q_MX02 U6126 ( .S(shiftCount[6]), .A0(n3393), .A1(n3329), .Z(n2752));
Q_MX02 U6127 ( .S(shiftCount[6]), .A0(n3392), .A1(n3328), .Z(n2751));
Q_MX02 U6128 ( .S(shiftCount[6]), .A0(n3391), .A1(n3327), .Z(n2750));
Q_MX02 U6129 ( .S(shiftCount[6]), .A0(n3390), .A1(n3326), .Z(n2749));
Q_MX02 U6130 ( .S(shiftCount[6]), .A0(n3389), .A1(n3325), .Z(n2748));
Q_MX02 U6131 ( .S(shiftCount[6]), .A0(n3388), .A1(n3324), .Z(n2747));
Q_MX02 U6132 ( .S(shiftCount[6]), .A0(n3387), .A1(n3323), .Z(n2746));
Q_MX02 U6133 ( .S(shiftCount[6]), .A0(n3386), .A1(n3322), .Z(n2745));
Q_MX02 U6134 ( .S(shiftCount[6]), .A0(n3385), .A1(n3321), .Z(n2744));
Q_MX02 U6135 ( .S(shiftCount[6]), .A0(n3384), .A1(n3320), .Z(n2743));
Q_MX02 U6136 ( .S(shiftCount[6]), .A0(n3383), .A1(n3319), .Z(n2742));
Q_MX02 U6137 ( .S(shiftCount[6]), .A0(n3382), .A1(n3318), .Z(n2741));
Q_MX02 U6138 ( .S(shiftCount[6]), .A0(n3381), .A1(n3317), .Z(n2740));
Q_MX02 U6139 ( .S(shiftCount[6]), .A0(n3380), .A1(n3316), .Z(n2739));
Q_MX02 U6140 ( .S(shiftCount[6]), .A0(n3379), .A1(n3315), .Z(n2738));
Q_MX02 U6141 ( .S(shiftCount[6]), .A0(n3378), .A1(n3314), .Z(n2737));
Q_MX02 U6142 ( .S(shiftCount[6]), .A0(n3377), .A1(n3313), .Z(n2736));
Q_MX02 U6143 ( .S(shiftCount[6]), .A0(n3376), .A1(n3312), .Z(n2735));
Q_MX02 U6144 ( .S(shiftCount[6]), .A0(n3375), .A1(n3311), .Z(n2734));
Q_MX02 U6145 ( .S(shiftCount[6]), .A0(n3374), .A1(n3310), .Z(n2733));
Q_MX02 U6146 ( .S(shiftCount[6]), .A0(n3373), .A1(n3309), .Z(n2732));
Q_MX02 U6147 ( .S(shiftCount[6]), .A0(n3372), .A1(n3308), .Z(n2731));
Q_MX02 U6148 ( .S(shiftCount[6]), .A0(n3371), .A1(n3307), .Z(n2730));
Q_MX02 U6149 ( .S(shiftCount[6]), .A0(n3370), .A1(n3306), .Z(n2729));
Q_MX02 U6150 ( .S(shiftCount[6]), .A0(n3369), .A1(n3305), .Z(n2728));
Q_MX02 U6151 ( .S(shiftCount[6]), .A0(n3368), .A1(n3304), .Z(n2727));
Q_MX02 U6152 ( .S(shiftCount[6]), .A0(n3367), .A1(n3303), .Z(n2726));
Q_MX02 U6153 ( .S(shiftCount[6]), .A0(n3366), .A1(n3302), .Z(n2725));
Q_MX02 U6154 ( .S(shiftCount[6]), .A0(n3365), .A1(n3301), .Z(n2724));
Q_MX02 U6155 ( .S(shiftCount[6]), .A0(n3364), .A1(n3300), .Z(n2723));
Q_MX02 U6156 ( .S(shiftCount[6]), .A0(n3363), .A1(n3299), .Z(n2722));
Q_MX02 U6157 ( .S(shiftCount[6]), .A0(n3362), .A1(n3298), .Z(n2721));
Q_MX02 U6158 ( .S(shiftCount[6]), .A0(n3361), .A1(n3297), .Z(n2720));
Q_MX02 U6159 ( .S(shiftCount[6]), .A0(n3360), .A1(n3296), .Z(n2719));
Q_MX02 U6160 ( .S(shiftCount[6]), .A0(n3359), .A1(n3295), .Z(n2718));
Q_MX02 U6161 ( .S(shiftCount[6]), .A0(n3358), .A1(n3294), .Z(n2717));
Q_MX02 U6162 ( .S(shiftCount[6]), .A0(n3357), .A1(n3293), .Z(n2716));
Q_MX02 U6163 ( .S(shiftCount[6]), .A0(n3356), .A1(n3292), .Z(n2715));
Q_MX02 U6164 ( .S(shiftCount[6]), .A0(n3355), .A1(n3291), .Z(n2714));
Q_MX02 U6165 ( .S(shiftCount[6]), .A0(n3354), .A1(n3290), .Z(n2713));
Q_MX02 U6166 ( .S(shiftCount[6]), .A0(n3353), .A1(n3289), .Z(n2712));
Q_MX02 U6167 ( .S(shiftCount[6]), .A0(n3352), .A1(n3288), .Z(n2711));
Q_MX02 U6168 ( .S(shiftCount[6]), .A0(n3351), .A1(n3287), .Z(n2710));
Q_MX02 U6169 ( .S(shiftCount[6]), .A0(n3350), .A1(n3286), .Z(n2709));
Q_MX02 U6170 ( .S(shiftCount[6]), .A0(n3349), .A1(n3285), .Z(n2708));
Q_MX02 U6171 ( .S(shiftCount[6]), .A0(n3348), .A1(n3284), .Z(n2707));
Q_MX02 U6172 ( .S(shiftCount[6]), .A0(n3347), .A1(n3283), .Z(n2706));
Q_MX02 U6173 ( .S(shiftCount[6]), .A0(n3346), .A1(n3282), .Z(n2705));
Q_MX02 U6174 ( .S(shiftCount[6]), .A0(n3345), .A1(n3281), .Z(n2704));
Q_MX02 U6175 ( .S(shiftCount[6]), .A0(n3344), .A1(n3280), .Z(n2703));
Q_MX02 U6176 ( .S(shiftCount[6]), .A0(n3343), .A1(n3279), .Z(n2702));
Q_MX02 U6177 ( .S(shiftCount[6]), .A0(n3342), .A1(n3278), .Z(n2701));
Q_MX02 U6178 ( .S(shiftCount[6]), .A0(n3341), .A1(n3277), .Z(n2700));
Q_MX02 U6179 ( .S(shiftCount[6]), .A0(n3340), .A1(n3276), .Z(n2699));
Q_MX02 U6180 ( .S(shiftCount[6]), .A0(n3339), .A1(n3275), .Z(n2698));
Q_MX02 U6181 ( .S(shiftCount[6]), .A0(n3338), .A1(n3274), .Z(n2697));
Q_MX02 U6182 ( .S(shiftCount[6]), .A0(n3337), .A1(n3273), .Z(n2696));
Q_MX02 U6183 ( .S(shiftCount[6]), .A0(n3336), .A1(n3272), .Z(n2695));
Q_MX02 U6184 ( .S(shiftCount[6]), .A0(n3335), .A1(n3271), .Z(n2694));
Q_MX02 U6185 ( .S(shiftCount[6]), .A0(n3334), .A1(n3270), .Z(n2693));
Q_MX02 U6186 ( .S(shiftCount[6]), .A0(n3333), .A1(n3269), .Z(n2692));
Q_MX02 U6187 ( .S(shiftCount[6]), .A0(n3332), .A1(n3268), .Z(n2691));
Q_MX02 U6188 ( .S(shiftCount[6]), .A0(n3331), .A1(n3267), .Z(n2690));
Q_MX02 U6189 ( .S(shiftCount[6]), .A0(n3330), .A1(n3266), .Z(n2689));
Q_MX02 U6190 ( .S(shiftCount[6]), .A0(n3329), .A1(n3265), .Z(n2688));
Q_MX02 U6191 ( .S(shiftCount[6]), .A0(n3328), .A1(n3264), .Z(n2687));
Q_MX02 U6192 ( .S(shiftCount[6]), .A0(n3327), .A1(n3263), .Z(n2686));
Q_MX02 U6193 ( .S(shiftCount[6]), .A0(n3326), .A1(n3262), .Z(n2685));
Q_MX02 U6194 ( .S(shiftCount[6]), .A0(n3325), .A1(n3261), .Z(n2684));
Q_MX02 U6195 ( .S(shiftCount[6]), .A0(n3324), .A1(n3260), .Z(n2683));
Q_MX02 U6196 ( .S(shiftCount[6]), .A0(n3323), .A1(n3259), .Z(n2682));
Q_MX02 U6197 ( .S(shiftCount[6]), .A0(n3322), .A1(n3258), .Z(n2681));
Q_MX02 U6198 ( .S(shiftCount[6]), .A0(n3321), .A1(n3257), .Z(n2680));
Q_MX02 U6199 ( .S(shiftCount[6]), .A0(n3320), .A1(n3256), .Z(n2679));
Q_MX02 U6200 ( .S(shiftCount[6]), .A0(n3319), .A1(n3255), .Z(n2678));
Q_MX02 U6201 ( .S(shiftCount[6]), .A0(n3318), .A1(n3254), .Z(n2677));
Q_MX02 U6202 ( .S(shiftCount[6]), .A0(n3317), .A1(n3253), .Z(n2676));
Q_MX02 U6203 ( .S(shiftCount[6]), .A0(n3316), .A1(n3252), .Z(n2675));
Q_MX02 U6204 ( .S(shiftCount[6]), .A0(n3315), .A1(n3251), .Z(n2674));
Q_MX02 U6205 ( .S(shiftCount[6]), .A0(n3314), .A1(n3250), .Z(n2673));
Q_MX02 U6206 ( .S(shiftCount[6]), .A0(n3313), .A1(n3249), .Z(n2672));
Q_MX02 U6207 ( .S(shiftCount[6]), .A0(n3312), .A1(n3248), .Z(n2671));
Q_MX02 U6208 ( .S(shiftCount[6]), .A0(n3311), .A1(n3247), .Z(n2670));
Q_MX02 U6209 ( .S(shiftCount[6]), .A0(n3310), .A1(n3246), .Z(n2669));
Q_MX02 U6210 ( .S(shiftCount[6]), .A0(n3309), .A1(n3245), .Z(n2668));
Q_MX02 U6211 ( .S(shiftCount[6]), .A0(n3308), .A1(n3244), .Z(n2667));
Q_MX02 U6212 ( .S(shiftCount[6]), .A0(n3307), .A1(n3243), .Z(n2666));
Q_MX02 U6213 ( .S(shiftCount[6]), .A0(n3306), .A1(n3242), .Z(n2665));
Q_MX02 U6214 ( .S(shiftCount[6]), .A0(n3305), .A1(n3241), .Z(n2664));
Q_MX02 U6215 ( .S(shiftCount[6]), .A0(n3304), .A1(n3240), .Z(n2663));
Q_MX02 U6216 ( .S(shiftCount[6]), .A0(n3303), .A1(n3239), .Z(n2662));
Q_MX02 U6217 ( .S(shiftCount[6]), .A0(n3302), .A1(n3238), .Z(n2661));
Q_MX02 U6218 ( .S(shiftCount[6]), .A0(n3301), .A1(n3237), .Z(n2660));
Q_MX02 U6219 ( .S(shiftCount[6]), .A0(n3300), .A1(n3236), .Z(n2659));
Q_MX02 U6220 ( .S(shiftCount[6]), .A0(n3299), .A1(n3235), .Z(n2658));
Q_MX02 U6221 ( .S(shiftCount[6]), .A0(n3298), .A1(n3234), .Z(n2657));
Q_MX02 U6222 ( .S(shiftCount[6]), .A0(n3297), .A1(n3233), .Z(n2656));
Q_MX02 U6223 ( .S(shiftCount[6]), .A0(n3296), .A1(n3232), .Z(n2655));
Q_MX02 U6224 ( .S(shiftCount[6]), .A0(n3295), .A1(n3231), .Z(n2654));
Q_MX02 U6225 ( .S(shiftCount[6]), .A0(n3294), .A1(n3230), .Z(n2653));
Q_MX02 U6226 ( .S(shiftCount[6]), .A0(n3293), .A1(n3229), .Z(n2652));
Q_MX02 U6227 ( .S(shiftCount[6]), .A0(n3292), .A1(n3228), .Z(n2651));
Q_MX02 U6228 ( .S(shiftCount[6]), .A0(n3291), .A1(n3227), .Z(n2650));
Q_MX02 U6229 ( .S(shiftCount[6]), .A0(n3290), .A1(n3226), .Z(n2649));
Q_MX02 U6230 ( .S(shiftCount[6]), .A0(n3289), .A1(n3225), .Z(n2648));
Q_MX02 U6231 ( .S(shiftCount[6]), .A0(n3288), .A1(n3224), .Z(n2647));
Q_MX02 U6232 ( .S(shiftCount[6]), .A0(n3287), .A1(n3223), .Z(n2646));
Q_MX02 U6233 ( .S(shiftCount[6]), .A0(n3286), .A1(n3222), .Z(n2645));
Q_MX02 U6234 ( .S(shiftCount[6]), .A0(n3285), .A1(n3221), .Z(n2644));
Q_MX02 U6235 ( .S(shiftCount[6]), .A0(n3284), .A1(n3220), .Z(n2643));
Q_MX02 U6236 ( .S(shiftCount[6]), .A0(n3283), .A1(n3219), .Z(n2642));
Q_MX02 U6237 ( .S(shiftCount[6]), .A0(n3282), .A1(n3218), .Z(n2641));
Q_MX02 U6238 ( .S(shiftCount[6]), .A0(n3281), .A1(n3217), .Z(n2640));
Q_MX02 U6239 ( .S(shiftCount[6]), .A0(n3280), .A1(n3216), .Z(n2639));
Q_MX02 U6240 ( .S(shiftCount[6]), .A0(n3279), .A1(n3215), .Z(n2638));
Q_MX02 U6241 ( .S(shiftCount[6]), .A0(n3278), .A1(n3214), .Z(n2637));
Q_MX02 U6242 ( .S(shiftCount[6]), .A0(n3277), .A1(n3213), .Z(n2636));
Q_MX02 U6243 ( .S(shiftCount[6]), .A0(n3276), .A1(n3212), .Z(n2635));
Q_MX02 U6244 ( .S(shiftCount[6]), .A0(n3275), .A1(n3211), .Z(n2634));
Q_MX02 U6245 ( .S(shiftCount[6]), .A0(n3274), .A1(n3210), .Z(n2633));
Q_MX02 U6246 ( .S(shiftCount[6]), .A0(n3273), .A1(n3209), .Z(n2632));
Q_MX02 U6247 ( .S(shiftCount[6]), .A0(n3272), .A1(n3208), .Z(n2631));
Q_MX02 U6248 ( .S(shiftCount[6]), .A0(n3271), .A1(n3207), .Z(n2630));
Q_MX02 U6249 ( .S(shiftCount[6]), .A0(n3270), .A1(n3206), .Z(n2629));
Q_MX02 U6250 ( .S(shiftCount[6]), .A0(n3269), .A1(n3205), .Z(n2628));
Q_MX02 U6251 ( .S(shiftCount[6]), .A0(n3268), .A1(n3204), .Z(n2627));
Q_MX02 U6252 ( .S(shiftCount[6]), .A0(n3267), .A1(n3203), .Z(n2626));
Q_MX02 U6253 ( .S(shiftCount[6]), .A0(n3266), .A1(n3202), .Z(n2625));
Q_MX02 U6254 ( .S(shiftCount[6]), .A0(n3265), .A1(n3201), .Z(n2624));
Q_MX02 U6255 ( .S(shiftCount[6]), .A0(n3264), .A1(n3200), .Z(n2623));
Q_MX02 U6256 ( .S(shiftCount[6]), .A0(n3263), .A1(n3199), .Z(n2622));
Q_MX02 U6257 ( .S(shiftCount[6]), .A0(n3262), .A1(n3198), .Z(n2621));
Q_MX02 U6258 ( .S(shiftCount[6]), .A0(n3261), .A1(n3197), .Z(n2620));
Q_MX02 U6259 ( .S(shiftCount[6]), .A0(n3260), .A1(n3196), .Z(n2619));
Q_MX02 U6260 ( .S(shiftCount[6]), .A0(n3259), .A1(n3195), .Z(n2618));
Q_MX02 U6261 ( .S(shiftCount[6]), .A0(n3258), .A1(n3194), .Z(n2617));
Q_MX02 U6262 ( .S(shiftCount[6]), .A0(n3257), .A1(n3193), .Z(n2616));
Q_MX02 U6263 ( .S(shiftCount[6]), .A0(n3256), .A1(n3192), .Z(n2615));
Q_MX02 U6264 ( .S(shiftCount[6]), .A0(n3255), .A1(n3191), .Z(n2614));
Q_MX02 U6265 ( .S(shiftCount[6]), .A0(n3254), .A1(n3190), .Z(n2613));
Q_MX02 U6266 ( .S(shiftCount[6]), .A0(n3253), .A1(n3189), .Z(n2612));
Q_MX02 U6267 ( .S(shiftCount[6]), .A0(n3252), .A1(n3188), .Z(n2611));
Q_MX02 U6268 ( .S(shiftCount[6]), .A0(n3251), .A1(n3187), .Z(n2610));
Q_MX02 U6269 ( .S(shiftCount[6]), .A0(n3250), .A1(n3186), .Z(n2609));
Q_MX02 U6270 ( .S(shiftCount[6]), .A0(n3249), .A1(n3185), .Z(n2608));
Q_MX02 U6271 ( .S(shiftCount[6]), .A0(n3248), .A1(n3184), .Z(n2607));
Q_MX02 U6272 ( .S(shiftCount[6]), .A0(n3247), .A1(n3183), .Z(n2606));
Q_MX02 U6273 ( .S(shiftCount[6]), .A0(n3246), .A1(n3182), .Z(n2605));
Q_MX02 U6274 ( .S(shiftCount[6]), .A0(n3245), .A1(n3181), .Z(n2604));
Q_MX02 U6275 ( .S(shiftCount[6]), .A0(n3244), .A1(n3180), .Z(n2603));
Q_MX02 U6276 ( .S(shiftCount[6]), .A0(n3243), .A1(n3179), .Z(n2602));
Q_MX02 U6277 ( .S(shiftCount[6]), .A0(n3242), .A1(n3178), .Z(n2601));
Q_MX02 U6278 ( .S(shiftCount[6]), .A0(n3241), .A1(n3177), .Z(n2600));
Q_MX02 U6279 ( .S(shiftCount[6]), .A0(n3240), .A1(n3176), .Z(n2599));
Q_MX02 U6280 ( .S(shiftCount[6]), .A0(n3239), .A1(n3175), .Z(n2598));
Q_MX02 U6281 ( .S(shiftCount[6]), .A0(n3238), .A1(n3174), .Z(n2597));
Q_MX02 U6282 ( .S(shiftCount[6]), .A0(n3237), .A1(n3173), .Z(n2596));
Q_MX02 U6283 ( .S(shiftCount[6]), .A0(n3236), .A1(n3172), .Z(n2595));
Q_MX02 U6284 ( .S(shiftCount[6]), .A0(n3235), .A1(n3171), .Z(n2594));
Q_MX02 U6285 ( .S(shiftCount[6]), .A0(n3234), .A1(n3170), .Z(n2593));
Q_MX02 U6286 ( .S(shiftCount[6]), .A0(n3233), .A1(n3169), .Z(n2592));
Q_MX02 U6287 ( .S(shiftCount[6]), .A0(n3232), .A1(n3168), .Z(n2591));
Q_MX02 U6288 ( .S(shiftCount[6]), .A0(n3231), .A1(n3167), .Z(n2590));
Q_MX02 U6289 ( .S(shiftCount[6]), .A0(n3230), .A1(n3166), .Z(n2589));
Q_MX02 U6290 ( .S(shiftCount[6]), .A0(n3229), .A1(n3165), .Z(n2588));
Q_MX02 U6291 ( .S(shiftCount[6]), .A0(n3228), .A1(n3164), .Z(n2587));
Q_MX02 U6292 ( .S(shiftCount[6]), .A0(n3227), .A1(n3163), .Z(n2586));
Q_MX02 U6293 ( .S(shiftCount[6]), .A0(n3226), .A1(n3162), .Z(n2585));
Q_MX02 U6294 ( .S(shiftCount[6]), .A0(n3225), .A1(n3161), .Z(n2584));
Q_MX02 U6295 ( .S(shiftCount[6]), .A0(n3224), .A1(n3160), .Z(n2583));
Q_MX02 U6296 ( .S(shiftCount[6]), .A0(n3223), .A1(n3159), .Z(n2582));
Q_MX02 U6297 ( .S(shiftCount[6]), .A0(n3222), .A1(n3158), .Z(n2581));
Q_MX02 U6298 ( .S(shiftCount[6]), .A0(n3221), .A1(n3157), .Z(n2580));
Q_MX02 U6299 ( .S(shiftCount[6]), .A0(n3220), .A1(n3156), .Z(n2579));
Q_MX02 U6300 ( .S(shiftCount[6]), .A0(n3219), .A1(n3155), .Z(n2578));
Q_MX02 U6301 ( .S(shiftCount[6]), .A0(n3218), .A1(n3154), .Z(n2577));
Q_MX02 U6302 ( .S(shiftCount[6]), .A0(n3217), .A1(n3153), .Z(n2576));
Q_MX02 U6303 ( .S(shiftCount[6]), .A0(n3216), .A1(n3152), .Z(n2575));
Q_MX02 U6304 ( .S(shiftCount[6]), .A0(n3215), .A1(n3151), .Z(n2574));
Q_MX02 U6305 ( .S(shiftCount[6]), .A0(n3214), .A1(n3150), .Z(n2573));
Q_MX02 U6306 ( .S(shiftCount[6]), .A0(n3213), .A1(n3149), .Z(n2572));
Q_MX02 U6307 ( .S(shiftCount[6]), .A0(n3212), .A1(n3148), .Z(n2571));
Q_MX02 U6308 ( .S(shiftCount[6]), .A0(n3211), .A1(n3147), .Z(n2570));
Q_MX02 U6309 ( .S(shiftCount[6]), .A0(n3210), .A1(n3146), .Z(n2569));
Q_MX02 U6310 ( .S(shiftCount[6]), .A0(n3209), .A1(n3145), .Z(n2568));
Q_MX02 U6311 ( .S(shiftCount[6]), .A0(n3208), .A1(n3144), .Z(n2567));
Q_MX02 U6312 ( .S(shiftCount[6]), .A0(n3207), .A1(n3143), .Z(n2566));
Q_MX02 U6313 ( .S(shiftCount[6]), .A0(n3206), .A1(n3142), .Z(n2565));
Q_MX02 U6314 ( .S(shiftCount[6]), .A0(n3205), .A1(n3141), .Z(n2564));
Q_MX02 U6315 ( .S(shiftCount[6]), .A0(n3204), .A1(n3140), .Z(n2563));
Q_MX02 U6316 ( .S(shiftCount[6]), .A0(n3203), .A1(n3139), .Z(n2562));
Q_MX02 U6317 ( .S(shiftCount[6]), .A0(n3202), .A1(n3138), .Z(n2561));
Q_MX02 U6318 ( .S(shiftCount[6]), .A0(n3201), .A1(n3137), .Z(n2560));
Q_MX02 U6319 ( .S(shiftCount[6]), .A0(n3200), .A1(n3136), .Z(n2559));
Q_MX02 U6320 ( .S(shiftCount[6]), .A0(n3199), .A1(n3135), .Z(n2558));
Q_MX02 U6321 ( .S(shiftCount[6]), .A0(n3198), .A1(n3134), .Z(n2557));
Q_MX02 U6322 ( .S(shiftCount[6]), .A0(n3197), .A1(n3133), .Z(n2556));
Q_MX02 U6323 ( .S(shiftCount[6]), .A0(n3196), .A1(n3132), .Z(n2555));
Q_MX02 U6324 ( .S(shiftCount[6]), .A0(n3195), .A1(n3131), .Z(n2554));
Q_MX02 U6325 ( .S(shiftCount[6]), .A0(n3194), .A1(n3130), .Z(n2553));
Q_MX02 U6326 ( .S(shiftCount[6]), .A0(n3193), .A1(n3129), .Z(n2552));
Q_MX02 U6327 ( .S(shiftCount[6]), .A0(n3192), .A1(n3128), .Z(n2551));
Q_MX02 U6328 ( .S(shiftCount[6]), .A0(n3191), .A1(n3127), .Z(n2550));
Q_MX02 U6329 ( .S(shiftCount[6]), .A0(n3190), .A1(n3126), .Z(n2549));
Q_MX02 U6330 ( .S(shiftCount[6]), .A0(n3189), .A1(n3125), .Z(n2548));
Q_MX02 U6331 ( .S(shiftCount[6]), .A0(n3188), .A1(n3124), .Z(n2547));
Q_MX02 U6332 ( .S(shiftCount[6]), .A0(n3187), .A1(n3123), .Z(n2546));
Q_MX02 U6333 ( .S(shiftCount[6]), .A0(n3186), .A1(n3122), .Z(n2545));
Q_MX02 U6334 ( .S(shiftCount[6]), .A0(n3185), .A1(n3121), .Z(n2544));
Q_MX02 U6335 ( .S(shiftCount[6]), .A0(n3184), .A1(n3120), .Z(n2543));
Q_MX02 U6336 ( .S(shiftCount[6]), .A0(n3183), .A1(n3119), .Z(n2542));
Q_MX02 U6337 ( .S(shiftCount[6]), .A0(n3182), .A1(n3118), .Z(n2541));
Q_MX02 U6338 ( .S(shiftCount[6]), .A0(n3181), .A1(n3117), .Z(n2540));
Q_MX02 U6339 ( .S(shiftCount[6]), .A0(n3180), .A1(n3116), .Z(n2539));
Q_MX02 U6340 ( .S(shiftCount[6]), .A0(n3179), .A1(n3115), .Z(n2538));
Q_MX02 U6341 ( .S(shiftCount[6]), .A0(n3178), .A1(n3114), .Z(n2537));
Q_MX02 U6342 ( .S(shiftCount[6]), .A0(n3177), .A1(n3113), .Z(n2536));
Q_MX02 U6343 ( .S(shiftCount[6]), .A0(n3176), .A1(n3112), .Z(n2535));
Q_MX02 U6344 ( .S(shiftCount[6]), .A0(n3175), .A1(n3111), .Z(n2534));
Q_MX02 U6345 ( .S(shiftCount[6]), .A0(n3174), .A1(n3110), .Z(n2533));
Q_MX02 U6346 ( .S(shiftCount[6]), .A0(n3173), .A1(n3109), .Z(n2532));
Q_MX02 U6347 ( .S(shiftCount[6]), .A0(n3172), .A1(n3108), .Z(n2531));
Q_MX02 U6348 ( .S(shiftCount[6]), .A0(n3171), .A1(n3107), .Z(n2530));
Q_MX02 U6349 ( .S(shiftCount[6]), .A0(n3170), .A1(n3106), .Z(n2529));
Q_MX02 U6350 ( .S(shiftCount[6]), .A0(n3169), .A1(n3105), .Z(n2528));
Q_MX02 U6351 ( .S(shiftCount[6]), .A0(n3168), .A1(n3104), .Z(n2527));
Q_MX02 U6352 ( .S(shiftCount[6]), .A0(n3167), .A1(n3103), .Z(n2526));
Q_MX02 U6353 ( .S(shiftCount[6]), .A0(n3166), .A1(n3102), .Z(n2525));
Q_MX02 U6354 ( .S(shiftCount[6]), .A0(n3165), .A1(n3101), .Z(n2524));
Q_MX02 U6355 ( .S(shiftCount[6]), .A0(n3164), .A1(n3100), .Z(n2523));
Q_MX02 U6356 ( .S(shiftCount[6]), .A0(n3163), .A1(n3099), .Z(n2522));
Q_MX02 U6357 ( .S(shiftCount[6]), .A0(n3162), .A1(n3098), .Z(n2521));
Q_MX02 U6358 ( .S(shiftCount[6]), .A0(n3161), .A1(n3097), .Z(n2520));
Q_MX02 U6359 ( .S(shiftCount[6]), .A0(n3160), .A1(n3096), .Z(n2519));
Q_MX02 U6360 ( .S(shiftCount[6]), .A0(n3159), .A1(n3095), .Z(n2518));
Q_MX02 U6361 ( .S(shiftCount[6]), .A0(n3158), .A1(n3094), .Z(n2517));
Q_MX02 U6362 ( .S(shiftCount[6]), .A0(n3157), .A1(n3093), .Z(n2516));
Q_MX02 U6363 ( .S(shiftCount[6]), .A0(n3156), .A1(n3092), .Z(n2515));
Q_MX02 U6364 ( .S(shiftCount[6]), .A0(n3155), .A1(n3091), .Z(n2514));
Q_MX02 U6365 ( .S(shiftCount[6]), .A0(n3154), .A1(n3090), .Z(n2513));
Q_MX02 U6366 ( .S(shiftCount[6]), .A0(n3153), .A1(n3089), .Z(n2512));
Q_MX02 U6367 ( .S(shiftCount[6]), .A0(n3152), .A1(n3088), .Z(n2511));
Q_MX02 U6368 ( .S(shiftCount[6]), .A0(n3151), .A1(n3087), .Z(n2510));
Q_MX02 U6369 ( .S(shiftCount[6]), .A0(n3150), .A1(n3086), .Z(n2509));
Q_MX02 U6370 ( .S(shiftCount[6]), .A0(n3149), .A1(n3085), .Z(n2508));
Q_MX02 U6371 ( .S(shiftCount[6]), .A0(n3148), .A1(n3084), .Z(n2507));
Q_MX02 U6372 ( .S(shiftCount[6]), .A0(n3147), .A1(n3083), .Z(n2506));
Q_MX02 U6373 ( .S(shiftCount[6]), .A0(n3146), .A1(n3082), .Z(n2505));
Q_MX02 U6374 ( .S(shiftCount[6]), .A0(n3145), .A1(n3081), .Z(n2504));
Q_MX02 U6375 ( .S(shiftCount[6]), .A0(n3144), .A1(n3080), .Z(n2503));
Q_MX02 U6376 ( .S(shiftCount[6]), .A0(n3143), .A1(n3079), .Z(n2502));
Q_MX02 U6377 ( .S(shiftCount[6]), .A0(n3142), .A1(n3077), .Z(n2501));
Q_MX02 U6378 ( .S(shiftCount[6]), .A0(n3141), .A1(n3076), .Z(n2500));
Q_MX02 U6379 ( .S(shiftCount[6]), .A0(n3140), .A1(n3075), .Z(n2499));
Q_MX02 U6380 ( .S(shiftCount[6]), .A0(n3139), .A1(n3074), .Z(n2498));
Q_MX02 U6381 ( .S(shiftCount[6]), .A0(n3138), .A1(n3073), .Z(n2497));
Q_MX02 U6382 ( .S(shiftCount[6]), .A0(n3137), .A1(n3072), .Z(n2496));
Q_MX02 U6383 ( .S(shiftCount[6]), .A0(n3136), .A1(n3071), .Z(n2495));
Q_MX02 U6384 ( .S(shiftCount[6]), .A0(n3135), .A1(n3070), .Z(n2494));
Q_MX02 U6385 ( .S(shiftCount[6]), .A0(n3134), .A1(n3069), .Z(n2493));
Q_MX02 U6386 ( .S(shiftCount[6]), .A0(n3133), .A1(n3068), .Z(n2492));
Q_MX02 U6387 ( .S(shiftCount[6]), .A0(n3132), .A1(n3067), .Z(n2491));
Q_MX02 U6388 ( .S(shiftCount[6]), .A0(n3131), .A1(n3066), .Z(n2490));
Q_MX02 U6389 ( .S(shiftCount[6]), .A0(n3130), .A1(n3065), .Z(n2489));
Q_MX02 U6390 ( .S(shiftCount[6]), .A0(n3129), .A1(n3064), .Z(n2488));
Q_MX02 U6391 ( .S(shiftCount[6]), .A0(n3128), .A1(n3063), .Z(n2487));
Q_MX02 U6392 ( .S(shiftCount[6]), .A0(n3127), .A1(n3062), .Z(n2486));
Q_MX02 U6393 ( .S(shiftCount[6]), .A0(n3126), .A1(n3061), .Z(n2485));
Q_MX02 U6394 ( .S(shiftCount[6]), .A0(n3125), .A1(n3060), .Z(n2484));
Q_MX02 U6395 ( .S(shiftCount[6]), .A0(n3124), .A1(n3059), .Z(n2483));
Q_MX02 U6396 ( .S(shiftCount[6]), .A0(n3123), .A1(n3058), .Z(n2482));
Q_MX02 U6397 ( .S(shiftCount[6]), .A0(n3122), .A1(n3057), .Z(n2481));
Q_MX02 U6398 ( .S(shiftCount[6]), .A0(n3121), .A1(n3056), .Z(n2480));
Q_MX02 U6399 ( .S(shiftCount[6]), .A0(n3120), .A1(n3055), .Z(n2479));
Q_MX02 U6400 ( .S(shiftCount[6]), .A0(n3119), .A1(n3054), .Z(n2478));
Q_MX02 U6401 ( .S(shiftCount[6]), .A0(n3118), .A1(n3053), .Z(n2477));
Q_MX02 U6402 ( .S(shiftCount[6]), .A0(n3117), .A1(n3052), .Z(n2476));
Q_MX02 U6403 ( .S(shiftCount[6]), .A0(n3116), .A1(n3051), .Z(n2475));
Q_MX02 U6404 ( .S(shiftCount[6]), .A0(n3115), .A1(n3050), .Z(n2474));
Q_MX02 U6405 ( .S(shiftCount[6]), .A0(n3114), .A1(n3049), .Z(n2473));
Q_MX02 U6406 ( .S(shiftCount[6]), .A0(n3113), .A1(n3048), .Z(n2472));
Q_MX02 U6407 ( .S(shiftCount[6]), .A0(n3112), .A1(n3047), .Z(n2471));
Q_MX02 U6408 ( .S(shiftCount[6]), .A0(n3111), .A1(n3046), .Z(n2470));
Q_INV U6409 ( .A(shiftCount[6]), .Z(n2469));
Q_AN02 U6410 ( .A0(n2469), .A1(n3110), .Z(n2468));
Q_AN02 U6411 ( .A0(n2469), .A1(n3109), .Z(n2467));
Q_AN02 U6412 ( .A0(n2469), .A1(n3108), .Z(n2466));
Q_AN02 U6413 ( .A0(n2469), .A1(n3107), .Z(n2465));
Q_AN02 U6414 ( .A0(n2469), .A1(n3106), .Z(n2464));
Q_AN02 U6415 ( .A0(n2469), .A1(n3105), .Z(n2463));
Q_AN02 U6416 ( .A0(n2469), .A1(n3104), .Z(n2462));
Q_AN02 U6417 ( .A0(n2469), .A1(n3103), .Z(n2461));
Q_AN02 U6418 ( .A0(n2469), .A1(n3102), .Z(n2460));
Q_AN02 U6419 ( .A0(n2469), .A1(n3101), .Z(n2459));
Q_AN02 U6420 ( .A0(n2469), .A1(n3100), .Z(n2458));
Q_AN02 U6421 ( .A0(n2469), .A1(n3099), .Z(n2457));
Q_AN02 U6422 ( .A0(n2469), .A1(n3098), .Z(n2456));
Q_AN02 U6423 ( .A0(n2469), .A1(n3097), .Z(n2455));
Q_AN02 U6424 ( .A0(n2469), .A1(n3096), .Z(n2454));
Q_AN02 U6425 ( .A0(n2469), .A1(n3095), .Z(n2453));
Q_AN02 U6426 ( .A0(n2469), .A1(n3094), .Z(n2452));
Q_AN02 U6427 ( .A0(n2469), .A1(n3093), .Z(n2451));
Q_AN02 U6428 ( .A0(n2469), .A1(n3092), .Z(n2450));
Q_AN02 U6429 ( .A0(n2469), .A1(n3091), .Z(n2449));
Q_AN02 U6430 ( .A0(n2469), .A1(n3090), .Z(n2448));
Q_AN02 U6431 ( .A0(n2469), .A1(n3089), .Z(n2447));
Q_AN02 U6432 ( .A0(n2469), .A1(n3088), .Z(n2446));
Q_AN02 U6433 ( .A0(n2469), .A1(n3087), .Z(n2445));
Q_AN02 U6434 ( .A0(n2469), .A1(n3086), .Z(n2444));
Q_AN02 U6435 ( .A0(n2469), .A1(n3085), .Z(n2443));
Q_AN02 U6436 ( .A0(n2469), .A1(n3084), .Z(n2442));
Q_AN02 U6437 ( .A0(n2469), .A1(n3083), .Z(n2441));
Q_AN02 U6438 ( .A0(n2469), .A1(n3082), .Z(n2440));
Q_AN02 U6439 ( .A0(n2469), .A1(n3081), .Z(n2439));
Q_AN02 U6440 ( .A0(n2469), .A1(n3080), .Z(n2438));
Q_AN02 U6441 ( .A0(n2469), .A1(n3079), .Z(n2437));
Q_AN02 U6442 ( .A0(n2469), .A1(n3077), .Z(n2436));
Q_AN02 U6443 ( .A0(n2469), .A1(n3076), .Z(n2435));
Q_AN02 U6444 ( .A0(n2469), .A1(n3075), .Z(n2434));
Q_AN02 U6445 ( .A0(n2469), .A1(n3074), .Z(n2433));
Q_AN02 U6446 ( .A0(n2469), .A1(n3073), .Z(n2432));
Q_AN02 U6447 ( .A0(n2469), .A1(n3072), .Z(n2431));
Q_AN02 U6448 ( .A0(n2469), .A1(n3071), .Z(n2430));
Q_AN02 U6449 ( .A0(n2469), .A1(n3070), .Z(n2429));
Q_AN02 U6450 ( .A0(n2469), .A1(n3069), .Z(n2428));
Q_AN02 U6451 ( .A0(n2469), .A1(n3068), .Z(n2427));
Q_AN02 U6452 ( .A0(n2469), .A1(n3067), .Z(n2426));
Q_AN02 U6453 ( .A0(n2469), .A1(n3066), .Z(n2425));
Q_AN02 U6454 ( .A0(n2469), .A1(n3065), .Z(n2424));
Q_AN02 U6455 ( .A0(n2469), .A1(n3064), .Z(n2423));
Q_AN02 U6456 ( .A0(n2469), .A1(n3063), .Z(n2422));
Q_AN02 U6457 ( .A0(n2469), .A1(n3062), .Z(n2421));
Q_AN02 U6458 ( .A0(n2469), .A1(n3061), .Z(n2420));
Q_AN02 U6459 ( .A0(n2469), .A1(n3060), .Z(n2419));
Q_AN02 U6460 ( .A0(n2469), .A1(n3059), .Z(n2418));
Q_AN02 U6461 ( .A0(n2469), .A1(n3058), .Z(n2417));
Q_AN02 U6462 ( .A0(n2469), .A1(n3057), .Z(n2416));
Q_AN02 U6463 ( .A0(n2469), .A1(n3056), .Z(n2415));
Q_AN02 U6464 ( .A0(n2469), .A1(n3055), .Z(n2414));
Q_AN02 U6465 ( .A0(n2469), .A1(n3054), .Z(n2413));
Q_AN02 U6466 ( .A0(n2469), .A1(n3053), .Z(n2412));
Q_AN02 U6467 ( .A0(n2469), .A1(n3052), .Z(n2411));
Q_AN02 U6468 ( .A0(n2469), .A1(n3051), .Z(n2410));
Q_AN02 U6469 ( .A0(n2469), .A1(n3050), .Z(n2409));
Q_AN02 U6470 ( .A0(n2469), .A1(n3049), .Z(n2408));
Q_AN02 U6471 ( .A0(n2469), .A1(n3048), .Z(n2407));
Q_AN02 U6472 ( .A0(n2469), .A1(n3047), .Z(n2406));
Q_AN02 U6473 ( .A0(n2469), .A1(n3046), .Z(n2405));
Q_AN02 U6474 ( .A0(shiftCount[7]), .A1(n3045), .Z(shiftedXdata[767]));
Q_AN02 U6475 ( .A0(shiftCount[7]), .A1(n3044), .Z(shiftedXdata[766]));
Q_AN02 U6476 ( .A0(shiftCount[7]), .A1(n3043), .Z(shiftedXdata[765]));
Q_AN02 U6477 ( .A0(shiftCount[7]), .A1(n3042), .Z(shiftedXdata[764]));
Q_AN02 U6478 ( .A0(shiftCount[7]), .A1(n3041), .Z(shiftedXdata[763]));
Q_AN02 U6479 ( .A0(shiftCount[7]), .A1(n3040), .Z(shiftedXdata[762]));
Q_AN02 U6480 ( .A0(shiftCount[7]), .A1(n3039), .Z(shiftedXdata[761]));
Q_AN02 U6481 ( .A0(shiftCount[7]), .A1(n3038), .Z(shiftedXdata[760]));
Q_AN02 U6482 ( .A0(shiftCount[7]), .A1(n3037), .Z(shiftedXdata[759]));
Q_AN02 U6483 ( .A0(shiftCount[7]), .A1(n3036), .Z(shiftedXdata[758]));
Q_AN02 U6484 ( .A0(shiftCount[7]), .A1(n3035), .Z(shiftedXdata[757]));
Q_AN02 U6485 ( .A0(shiftCount[7]), .A1(n3034), .Z(shiftedXdata[756]));
Q_AN02 U6486 ( .A0(shiftCount[7]), .A1(n3033), .Z(shiftedXdata[755]));
Q_AN02 U6487 ( .A0(shiftCount[7]), .A1(n3032), .Z(shiftedXdata[754]));
Q_AN02 U6488 ( .A0(shiftCount[7]), .A1(n3031), .Z(shiftedXdata[753]));
Q_AN02 U6489 ( .A0(shiftCount[7]), .A1(n3030), .Z(shiftedXdata[752]));
Q_AN02 U6490 ( .A0(shiftCount[7]), .A1(n3029), .Z(shiftedXdata[751]));
Q_AN02 U6491 ( .A0(shiftCount[7]), .A1(n3028), .Z(shiftedXdata[750]));
Q_AN02 U6492 ( .A0(shiftCount[7]), .A1(n3027), .Z(shiftedXdata[749]));
Q_AN02 U6493 ( .A0(shiftCount[7]), .A1(n3026), .Z(shiftedXdata[748]));
Q_AN02 U6494 ( .A0(shiftCount[7]), .A1(n3025), .Z(shiftedXdata[747]));
Q_AN02 U6495 ( .A0(shiftCount[7]), .A1(n3024), .Z(shiftedXdata[746]));
Q_AN02 U6496 ( .A0(shiftCount[7]), .A1(n3023), .Z(shiftedXdata[745]));
Q_AN02 U6497 ( .A0(shiftCount[7]), .A1(n3022), .Z(shiftedXdata[744]));
Q_AN02 U6498 ( .A0(shiftCount[7]), .A1(n3021), .Z(shiftedXdata[743]));
Q_AN02 U6499 ( .A0(shiftCount[7]), .A1(n3020), .Z(shiftedXdata[742]));
Q_AN02 U6500 ( .A0(shiftCount[7]), .A1(n3019), .Z(shiftedXdata[741]));
Q_AN02 U6501 ( .A0(shiftCount[7]), .A1(n3018), .Z(shiftedXdata[740]));
Q_AN02 U6502 ( .A0(shiftCount[7]), .A1(n3017), .Z(shiftedXdata[739]));
Q_AN02 U6503 ( .A0(shiftCount[7]), .A1(n3016), .Z(shiftedXdata[738]));
Q_AN02 U6504 ( .A0(shiftCount[7]), .A1(n3015), .Z(shiftedXdata[737]));
Q_AN02 U6505 ( .A0(shiftCount[7]), .A1(n3014), .Z(shiftedXdata[736]));
Q_AN02 U6506 ( .A0(shiftCount[7]), .A1(n3013), .Z(shiftedXdata[735]));
Q_AN02 U6507 ( .A0(shiftCount[7]), .A1(n3012), .Z(shiftedXdata[734]));
Q_AN02 U6508 ( .A0(shiftCount[7]), .A1(n3011), .Z(shiftedXdata[733]));
Q_AN02 U6509 ( .A0(shiftCount[7]), .A1(n3010), .Z(shiftedXdata[732]));
Q_AN02 U6510 ( .A0(shiftCount[7]), .A1(n3009), .Z(shiftedXdata[731]));
Q_AN02 U6511 ( .A0(shiftCount[7]), .A1(n3008), .Z(shiftedXdata[730]));
Q_AN02 U6512 ( .A0(shiftCount[7]), .A1(n3007), .Z(shiftedXdata[729]));
Q_AN02 U6513 ( .A0(shiftCount[7]), .A1(n3006), .Z(shiftedXdata[728]));
Q_AN02 U6514 ( .A0(shiftCount[7]), .A1(n3005), .Z(shiftedXdata[727]));
Q_AN02 U6515 ( .A0(shiftCount[7]), .A1(n3004), .Z(shiftedXdata[726]));
Q_AN02 U6516 ( .A0(shiftCount[7]), .A1(n3003), .Z(shiftedXdata[725]));
Q_AN02 U6517 ( .A0(shiftCount[7]), .A1(n3002), .Z(shiftedXdata[724]));
Q_AN02 U6518 ( .A0(shiftCount[7]), .A1(n3001), .Z(shiftedXdata[723]));
Q_AN02 U6519 ( .A0(shiftCount[7]), .A1(n3000), .Z(shiftedXdata[722]));
Q_AN02 U6520 ( .A0(shiftCount[7]), .A1(n2999), .Z(shiftedXdata[721]));
Q_AN02 U6521 ( .A0(shiftCount[7]), .A1(n2998), .Z(shiftedXdata[720]));
Q_AN02 U6522 ( .A0(shiftCount[7]), .A1(n2997), .Z(shiftedXdata[719]));
Q_AN02 U6523 ( .A0(shiftCount[7]), .A1(n2996), .Z(shiftedXdata[718]));
Q_AN02 U6524 ( .A0(shiftCount[7]), .A1(n2995), .Z(shiftedXdata[717]));
Q_AN02 U6525 ( .A0(shiftCount[7]), .A1(n2994), .Z(shiftedXdata[716]));
Q_AN02 U6526 ( .A0(shiftCount[7]), .A1(n2993), .Z(shiftedXdata[715]));
Q_AN02 U6527 ( .A0(shiftCount[7]), .A1(n2992), .Z(shiftedXdata[714]));
Q_AN02 U6528 ( .A0(shiftCount[7]), .A1(n2991), .Z(shiftedXdata[713]));
Q_AN02 U6529 ( .A0(shiftCount[7]), .A1(n2990), .Z(shiftedXdata[712]));
Q_AN02 U6530 ( .A0(shiftCount[7]), .A1(n2989), .Z(shiftedXdata[711]));
Q_AN02 U6531 ( .A0(shiftCount[7]), .A1(n2988), .Z(shiftedXdata[710]));
Q_AN02 U6532 ( .A0(shiftCount[7]), .A1(n2987), .Z(shiftedXdata[709]));
Q_AN02 U6533 ( .A0(shiftCount[7]), .A1(n2986), .Z(shiftedXdata[708]));
Q_AN02 U6534 ( .A0(shiftCount[7]), .A1(n2985), .Z(shiftedXdata[707]));
Q_AN02 U6535 ( .A0(shiftCount[7]), .A1(n2984), .Z(shiftedXdata[706]));
Q_AN02 U6536 ( .A0(shiftCount[7]), .A1(n2983), .Z(shiftedXdata[705]));
Q_AN02 U6537 ( .A0(shiftCount[7]), .A1(n2982), .Z(shiftedXdata[704]));
Q_AN02 U6538 ( .A0(shiftCount[7]), .A1(n2981), .Z(shiftedXdata[703]));
Q_AN02 U6539 ( .A0(shiftCount[7]), .A1(n2980), .Z(shiftedXdata[702]));
Q_AN02 U6540 ( .A0(shiftCount[7]), .A1(n2979), .Z(shiftedXdata[701]));
Q_AN02 U6541 ( .A0(shiftCount[7]), .A1(n2978), .Z(shiftedXdata[700]));
Q_AN02 U6542 ( .A0(shiftCount[7]), .A1(n2977), .Z(shiftedXdata[699]));
Q_AN02 U6543 ( .A0(shiftCount[7]), .A1(n2976), .Z(shiftedXdata[698]));
Q_AN02 U6544 ( .A0(shiftCount[7]), .A1(n2975), .Z(shiftedXdata[697]));
Q_AN02 U6545 ( .A0(shiftCount[7]), .A1(n2974), .Z(shiftedXdata[696]));
Q_AN02 U6546 ( .A0(shiftCount[7]), .A1(n2973), .Z(shiftedXdata[695]));
Q_AN02 U6547 ( .A0(shiftCount[7]), .A1(n2972), .Z(shiftedXdata[694]));
Q_AN02 U6548 ( .A0(shiftCount[7]), .A1(n2971), .Z(shiftedXdata[693]));
Q_AN02 U6549 ( .A0(shiftCount[7]), .A1(n2970), .Z(shiftedXdata[692]));
Q_AN02 U6550 ( .A0(shiftCount[7]), .A1(n2969), .Z(shiftedXdata[691]));
Q_AN02 U6551 ( .A0(shiftCount[7]), .A1(n2968), .Z(shiftedXdata[690]));
Q_AN02 U6552 ( .A0(shiftCount[7]), .A1(n2967), .Z(shiftedXdata[689]));
Q_AN02 U6553 ( .A0(shiftCount[7]), .A1(n2966), .Z(shiftedXdata[688]));
Q_AN02 U6554 ( .A0(shiftCount[7]), .A1(n2965), .Z(shiftedXdata[687]));
Q_AN02 U6555 ( .A0(shiftCount[7]), .A1(n2964), .Z(shiftedXdata[686]));
Q_AN02 U6556 ( .A0(shiftCount[7]), .A1(n2963), .Z(shiftedXdata[685]));
Q_AN02 U6557 ( .A0(shiftCount[7]), .A1(n2962), .Z(shiftedXdata[684]));
Q_AN02 U6558 ( .A0(shiftCount[7]), .A1(n2961), .Z(shiftedXdata[683]));
Q_AN02 U6559 ( .A0(shiftCount[7]), .A1(n2960), .Z(shiftedXdata[682]));
Q_AN02 U6560 ( .A0(shiftCount[7]), .A1(n2959), .Z(shiftedXdata[681]));
Q_AN02 U6561 ( .A0(shiftCount[7]), .A1(n2958), .Z(shiftedXdata[680]));
Q_AN02 U6562 ( .A0(shiftCount[7]), .A1(n2957), .Z(shiftedXdata[679]));
Q_AN02 U6563 ( .A0(shiftCount[7]), .A1(n2956), .Z(shiftedXdata[678]));
Q_AN02 U6564 ( .A0(shiftCount[7]), .A1(n2955), .Z(shiftedXdata[677]));
Q_AN02 U6565 ( .A0(shiftCount[7]), .A1(n2954), .Z(shiftedXdata[676]));
Q_AN02 U6566 ( .A0(shiftCount[7]), .A1(n2953), .Z(shiftedXdata[675]));
Q_AN02 U6567 ( .A0(shiftCount[7]), .A1(n2952), .Z(shiftedXdata[674]));
Q_AN02 U6568 ( .A0(shiftCount[7]), .A1(n2951), .Z(shiftedXdata[673]));
Q_AN02 U6569 ( .A0(shiftCount[7]), .A1(n2950), .Z(shiftedXdata[672]));
Q_AN02 U6570 ( .A0(shiftCount[7]), .A1(n2949), .Z(shiftedXdata[671]));
Q_AN02 U6571 ( .A0(shiftCount[7]), .A1(n2948), .Z(shiftedXdata[670]));
Q_AN02 U6572 ( .A0(shiftCount[7]), .A1(n2947), .Z(shiftedXdata[669]));
Q_AN02 U6573 ( .A0(shiftCount[7]), .A1(n2946), .Z(shiftedXdata[668]));
Q_AN02 U6574 ( .A0(shiftCount[7]), .A1(n2945), .Z(shiftedXdata[667]));
Q_AN02 U6575 ( .A0(shiftCount[7]), .A1(n2944), .Z(shiftedXdata[666]));
Q_AN02 U6576 ( .A0(shiftCount[7]), .A1(n2943), .Z(shiftedXdata[665]));
Q_AN02 U6577 ( .A0(shiftCount[7]), .A1(n2942), .Z(shiftedXdata[664]));
Q_AN02 U6578 ( .A0(shiftCount[7]), .A1(n2941), .Z(shiftedXdata[663]));
Q_AN02 U6579 ( .A0(shiftCount[7]), .A1(n2940), .Z(shiftedXdata[662]));
Q_AN02 U6580 ( .A0(shiftCount[7]), .A1(n2939), .Z(shiftedXdata[661]));
Q_AN02 U6581 ( .A0(shiftCount[7]), .A1(n2938), .Z(shiftedXdata[660]));
Q_AN02 U6582 ( .A0(shiftCount[7]), .A1(n2937), .Z(shiftedXdata[659]));
Q_AN02 U6583 ( .A0(shiftCount[7]), .A1(n2936), .Z(shiftedXdata[658]));
Q_AN02 U6584 ( .A0(shiftCount[7]), .A1(n2935), .Z(shiftedXdata[657]));
Q_AN02 U6585 ( .A0(shiftCount[7]), .A1(n2934), .Z(shiftedXdata[656]));
Q_AN02 U6586 ( .A0(shiftCount[7]), .A1(n2933), .Z(shiftedXdata[655]));
Q_AN02 U6587 ( .A0(shiftCount[7]), .A1(n2932), .Z(shiftedXdata[654]));
Q_AN02 U6588 ( .A0(shiftCount[7]), .A1(n2931), .Z(shiftedXdata[653]));
Q_AN02 U6589 ( .A0(shiftCount[7]), .A1(n2930), .Z(shiftedXdata[652]));
Q_AN02 U6590 ( .A0(shiftCount[7]), .A1(n2929), .Z(shiftedXdata[651]));
Q_AN02 U6591 ( .A0(shiftCount[7]), .A1(n2928), .Z(shiftedXdata[650]));
Q_AN02 U6592 ( .A0(shiftCount[7]), .A1(n2927), .Z(shiftedXdata[649]));
Q_AN02 U6593 ( .A0(shiftCount[7]), .A1(n2926), .Z(shiftedXdata[648]));
Q_AN02 U6594 ( .A0(shiftCount[7]), .A1(n2925), .Z(shiftedXdata[647]));
Q_AN02 U6595 ( .A0(shiftCount[7]), .A1(n2924), .Z(shiftedXdata[646]));
Q_AN02 U6596 ( .A0(shiftCount[7]), .A1(n2923), .Z(shiftedXdata[645]));
Q_AN02 U6597 ( .A0(shiftCount[7]), .A1(n2922), .Z(shiftedXdata[644]));
Q_AN02 U6598 ( .A0(shiftCount[7]), .A1(n2921), .Z(shiftedXdata[643]));
Q_AN02 U6599 ( .A0(shiftCount[7]), .A1(n2920), .Z(shiftedXdata[642]));
Q_AN02 U6600 ( .A0(shiftCount[7]), .A1(n2919), .Z(shiftedXdata[641]));
Q_AN02 U6601 ( .A0(shiftCount[7]), .A1(n2918), .Z(shiftedXdata[640]));
Q_MX02 U6602 ( .S(shiftCount[7]), .A0(n3045), .A1(n2917), .Z(shiftedXdata[639]));
Q_MX02 U6603 ( .S(shiftCount[7]), .A0(n3044), .A1(n2916), .Z(shiftedXdata[638]));
Q_MX02 U6604 ( .S(shiftCount[7]), .A0(n3043), .A1(n2915), .Z(shiftedXdata[637]));
Q_MX02 U6605 ( .S(shiftCount[7]), .A0(n3042), .A1(n2914), .Z(shiftedXdata[636]));
Q_MX02 U6606 ( .S(shiftCount[7]), .A0(n3041), .A1(n2913), .Z(shiftedXdata[635]));
Q_MX02 U6607 ( .S(shiftCount[7]), .A0(n3040), .A1(n2912), .Z(shiftedXdata[634]));
Q_MX02 U6608 ( .S(shiftCount[7]), .A0(n3039), .A1(n2911), .Z(shiftedXdata[633]));
Q_MX02 U6609 ( .S(shiftCount[7]), .A0(n3038), .A1(n2910), .Z(shiftedXdata[632]));
Q_MX02 U6610 ( .S(shiftCount[7]), .A0(n3037), .A1(n2909), .Z(shiftedXdata[631]));
Q_MX02 U6611 ( .S(shiftCount[7]), .A0(n3036), .A1(n2908), .Z(shiftedXdata[630]));
Q_MX02 U6612 ( .S(shiftCount[7]), .A0(n3035), .A1(n2907), .Z(shiftedXdata[629]));
Q_MX02 U6613 ( .S(shiftCount[7]), .A0(n3034), .A1(n2906), .Z(shiftedXdata[628]));
Q_MX02 U6614 ( .S(shiftCount[7]), .A0(n3033), .A1(n2905), .Z(shiftedXdata[627]));
Q_MX02 U6615 ( .S(shiftCount[7]), .A0(n3032), .A1(n2904), .Z(shiftedXdata[626]));
Q_MX02 U6616 ( .S(shiftCount[7]), .A0(n3031), .A1(n2903), .Z(shiftedXdata[625]));
Q_MX02 U6617 ( .S(shiftCount[7]), .A0(n3030), .A1(n2902), .Z(shiftedXdata[624]));
Q_MX02 U6618 ( .S(shiftCount[7]), .A0(n3029), .A1(n2901), .Z(shiftedXdata[623]));
Q_MX02 U6619 ( .S(shiftCount[7]), .A0(n3028), .A1(n2900), .Z(shiftedXdata[622]));
Q_MX02 U6620 ( .S(shiftCount[7]), .A0(n3027), .A1(n2899), .Z(shiftedXdata[621]));
Q_MX02 U6621 ( .S(shiftCount[7]), .A0(n3026), .A1(n2898), .Z(shiftedXdata[620]));
Q_MX02 U6622 ( .S(shiftCount[7]), .A0(n3025), .A1(n2897), .Z(shiftedXdata[619]));
Q_MX02 U6623 ( .S(shiftCount[7]), .A0(n3024), .A1(n2896), .Z(shiftedXdata[618]));
Q_MX02 U6624 ( .S(shiftCount[7]), .A0(n3023), .A1(n2895), .Z(shiftedXdata[617]));
Q_MX02 U6625 ( .S(shiftCount[7]), .A0(n3022), .A1(n2894), .Z(shiftedXdata[616]));
Q_MX02 U6626 ( .S(shiftCount[7]), .A0(n3021), .A1(n2893), .Z(shiftedXdata[615]));
Q_MX02 U6627 ( .S(shiftCount[7]), .A0(n3020), .A1(n2892), .Z(shiftedXdata[614]));
Q_MX02 U6628 ( .S(shiftCount[7]), .A0(n3019), .A1(n2891), .Z(shiftedXdata[613]));
Q_MX02 U6629 ( .S(shiftCount[7]), .A0(n3018), .A1(n2890), .Z(shiftedXdata[612]));
Q_MX02 U6630 ( .S(shiftCount[7]), .A0(n3017), .A1(n2889), .Z(shiftedXdata[611]));
Q_MX02 U6631 ( .S(shiftCount[7]), .A0(n3016), .A1(n2888), .Z(shiftedXdata[610]));
Q_MX02 U6632 ( .S(shiftCount[7]), .A0(n3015), .A1(n2887), .Z(shiftedXdata[609]));
Q_MX02 U6633 ( .S(shiftCount[7]), .A0(n3014), .A1(n2886), .Z(shiftedXdata[608]));
Q_MX02 U6634 ( .S(shiftCount[7]), .A0(n3013), .A1(n2885), .Z(shiftedXdata[607]));
Q_MX02 U6635 ( .S(shiftCount[7]), .A0(n3012), .A1(n2884), .Z(shiftedXdata[606]));
Q_MX02 U6636 ( .S(shiftCount[7]), .A0(n3011), .A1(n2883), .Z(shiftedXdata[605]));
Q_MX02 U6637 ( .S(shiftCount[7]), .A0(n3010), .A1(n2882), .Z(shiftedXdata[604]));
Q_MX02 U6638 ( .S(shiftCount[7]), .A0(n3009), .A1(n2881), .Z(shiftedXdata[603]));
Q_MX02 U6639 ( .S(shiftCount[7]), .A0(n3008), .A1(n2880), .Z(shiftedXdata[602]));
Q_MX02 U6640 ( .S(shiftCount[7]), .A0(n3007), .A1(n2879), .Z(shiftedXdata[601]));
Q_MX02 U6641 ( .S(shiftCount[7]), .A0(n3006), .A1(n2878), .Z(shiftedXdata[600]));
Q_MX02 U6642 ( .S(shiftCount[7]), .A0(n3005), .A1(n2877), .Z(shiftedXdata[599]));
Q_MX02 U6643 ( .S(shiftCount[7]), .A0(n3004), .A1(n2876), .Z(shiftedXdata[598]));
Q_MX02 U6644 ( .S(shiftCount[7]), .A0(n3003), .A1(n2875), .Z(shiftedXdata[597]));
Q_MX02 U6645 ( .S(shiftCount[7]), .A0(n3002), .A1(n2874), .Z(shiftedXdata[596]));
Q_MX02 U6646 ( .S(shiftCount[7]), .A0(n3001), .A1(n2873), .Z(shiftedXdata[595]));
Q_MX02 U6647 ( .S(shiftCount[7]), .A0(n3000), .A1(n2872), .Z(shiftedXdata[594]));
Q_MX02 U6648 ( .S(shiftCount[7]), .A0(n2999), .A1(n2871), .Z(shiftedXdata[593]));
Q_MX02 U6649 ( .S(shiftCount[7]), .A0(n2998), .A1(n2870), .Z(shiftedXdata[592]));
Q_MX02 U6650 ( .S(shiftCount[7]), .A0(n2997), .A1(n2869), .Z(shiftedXdata[591]));
Q_MX02 U6651 ( .S(shiftCount[7]), .A0(n2996), .A1(n2868), .Z(shiftedXdata[590]));
Q_MX02 U6652 ( .S(shiftCount[7]), .A0(n2995), .A1(n2867), .Z(shiftedXdata[589]));
Q_MX02 U6653 ( .S(shiftCount[7]), .A0(n2994), .A1(n2866), .Z(shiftedXdata[588]));
Q_MX02 U6654 ( .S(shiftCount[7]), .A0(n2993), .A1(n2865), .Z(shiftedXdata[587]));
Q_MX02 U6655 ( .S(shiftCount[7]), .A0(n2992), .A1(n2864), .Z(shiftedXdata[586]));
Q_MX02 U6656 ( .S(shiftCount[7]), .A0(n2991), .A1(n2863), .Z(shiftedXdata[585]));
Q_MX02 U6657 ( .S(shiftCount[7]), .A0(n2990), .A1(n2862), .Z(shiftedXdata[584]));
Q_MX02 U6658 ( .S(shiftCount[7]), .A0(n2989), .A1(n2861), .Z(shiftedXdata[583]));
Q_MX02 U6659 ( .S(shiftCount[7]), .A0(n2988), .A1(n2860), .Z(shiftedXdata[582]));
Q_MX02 U6660 ( .S(shiftCount[7]), .A0(n2987), .A1(n2859), .Z(shiftedXdata[581]));
Q_MX02 U6661 ( .S(shiftCount[7]), .A0(n2986), .A1(n2858), .Z(shiftedXdata[580]));
Q_MX02 U6662 ( .S(shiftCount[7]), .A0(n2985), .A1(n2857), .Z(shiftedXdata[579]));
Q_MX02 U6663 ( .S(shiftCount[7]), .A0(n2984), .A1(n2856), .Z(shiftedXdata[578]));
Q_MX02 U6664 ( .S(shiftCount[7]), .A0(n2983), .A1(n2855), .Z(shiftedXdata[577]));
Q_MX02 U6665 ( .S(shiftCount[7]), .A0(n2982), .A1(n2854), .Z(shiftedXdata[576]));
Q_MX02 U6666 ( .S(shiftCount[7]), .A0(n2981), .A1(n2853), .Z(shiftedXdata[575]));
Q_MX02 U6667 ( .S(shiftCount[7]), .A0(n2980), .A1(n2852), .Z(shiftedXdata[574]));
Q_MX02 U6668 ( .S(shiftCount[7]), .A0(n2979), .A1(n2851), .Z(shiftedXdata[573]));
Q_MX02 U6669 ( .S(shiftCount[7]), .A0(n2978), .A1(n2850), .Z(shiftedXdata[572]));
Q_MX02 U6670 ( .S(shiftCount[7]), .A0(n2977), .A1(n2849), .Z(shiftedXdata[571]));
Q_MX02 U6671 ( .S(shiftCount[7]), .A0(n2976), .A1(n2848), .Z(shiftedXdata[570]));
Q_MX02 U6672 ( .S(shiftCount[7]), .A0(n2975), .A1(n2847), .Z(shiftedXdata[569]));
Q_MX02 U6673 ( .S(shiftCount[7]), .A0(n2974), .A1(n2846), .Z(shiftedXdata[568]));
Q_MX02 U6674 ( .S(shiftCount[7]), .A0(n2973), .A1(n2845), .Z(shiftedXdata[567]));
Q_MX02 U6675 ( .S(shiftCount[7]), .A0(n2972), .A1(n2844), .Z(shiftedXdata[566]));
Q_MX02 U6676 ( .S(shiftCount[7]), .A0(n2971), .A1(n2843), .Z(shiftedXdata[565]));
Q_MX02 U6677 ( .S(shiftCount[7]), .A0(n2970), .A1(n2842), .Z(shiftedXdata[564]));
Q_MX02 U6678 ( .S(shiftCount[7]), .A0(n2969), .A1(n2841), .Z(shiftedXdata[563]));
Q_MX02 U6679 ( .S(shiftCount[7]), .A0(n2968), .A1(n2840), .Z(shiftedXdata[562]));
Q_MX02 U6680 ( .S(shiftCount[7]), .A0(n2967), .A1(n2839), .Z(shiftedXdata[561]));
Q_MX02 U6681 ( .S(shiftCount[7]), .A0(n2966), .A1(n2838), .Z(shiftedXdata[560]));
Q_MX02 U6682 ( .S(shiftCount[7]), .A0(n2965), .A1(n2837), .Z(shiftedXdata[559]));
Q_MX02 U6683 ( .S(shiftCount[7]), .A0(n2964), .A1(n2836), .Z(shiftedXdata[558]));
Q_MX02 U6684 ( .S(shiftCount[7]), .A0(n2963), .A1(n2835), .Z(shiftedXdata[557]));
Q_MX02 U6685 ( .S(shiftCount[7]), .A0(n2962), .A1(n2834), .Z(shiftedXdata[556]));
Q_MX02 U6686 ( .S(shiftCount[7]), .A0(n2961), .A1(n2833), .Z(shiftedXdata[555]));
Q_MX02 U6687 ( .S(shiftCount[7]), .A0(n2960), .A1(n2832), .Z(shiftedXdata[554]));
Q_MX02 U6688 ( .S(shiftCount[7]), .A0(n2959), .A1(n2831), .Z(shiftedXdata[553]));
Q_MX02 U6689 ( .S(shiftCount[7]), .A0(n2958), .A1(n2830), .Z(shiftedXdata[552]));
Q_MX02 U6690 ( .S(shiftCount[7]), .A0(n2957), .A1(n2829), .Z(shiftedXdata[551]));
Q_MX02 U6691 ( .S(shiftCount[7]), .A0(n2956), .A1(n2828), .Z(shiftedXdata[550]));
Q_MX02 U6692 ( .S(shiftCount[7]), .A0(n2955), .A1(n2827), .Z(shiftedXdata[549]));
Q_MX02 U6693 ( .S(shiftCount[7]), .A0(n2954), .A1(n2826), .Z(shiftedXdata[548]));
Q_MX02 U6694 ( .S(shiftCount[7]), .A0(n2953), .A1(n2825), .Z(shiftedXdata[547]));
Q_MX02 U6695 ( .S(shiftCount[7]), .A0(n2952), .A1(n2824), .Z(shiftedXdata[546]));
Q_MX02 U6696 ( .S(shiftCount[7]), .A0(n2951), .A1(n2823), .Z(shiftedXdata[545]));
Q_MX02 U6697 ( .S(shiftCount[7]), .A0(n2950), .A1(n2822), .Z(shiftedXdata[544]));
Q_MX02 U6698 ( .S(shiftCount[7]), .A0(n2949), .A1(n2821), .Z(shiftedXdata[543]));
Q_MX02 U6699 ( .S(shiftCount[7]), .A0(n2948), .A1(n2820), .Z(shiftedXdata[542]));
Q_MX02 U6700 ( .S(shiftCount[7]), .A0(n2947), .A1(n2819), .Z(shiftedXdata[541]));
Q_MX02 U6701 ( .S(shiftCount[7]), .A0(n2946), .A1(n2818), .Z(shiftedXdata[540]));
Q_MX02 U6702 ( .S(shiftCount[7]), .A0(n2945), .A1(n2817), .Z(shiftedXdata[539]));
Q_MX02 U6703 ( .S(shiftCount[7]), .A0(n2944), .A1(n2816), .Z(shiftedXdata[538]));
Q_MX02 U6704 ( .S(shiftCount[7]), .A0(n2943), .A1(n2815), .Z(shiftedXdata[537]));
Q_MX02 U6705 ( .S(shiftCount[7]), .A0(n2942), .A1(n2814), .Z(shiftedXdata[536]));
Q_MX02 U6706 ( .S(shiftCount[7]), .A0(n2941), .A1(n2813), .Z(shiftedXdata[535]));
Q_MX02 U6707 ( .S(shiftCount[7]), .A0(n2940), .A1(n2812), .Z(shiftedXdata[534]));
Q_MX02 U6708 ( .S(shiftCount[7]), .A0(n2939), .A1(n2811), .Z(shiftedXdata[533]));
Q_MX02 U6709 ( .S(shiftCount[7]), .A0(n2938), .A1(n2810), .Z(shiftedXdata[532]));
Q_MX02 U6710 ( .S(shiftCount[7]), .A0(n2937), .A1(n2809), .Z(shiftedXdata[531]));
Q_MX02 U6711 ( .S(shiftCount[7]), .A0(n2936), .A1(n2808), .Z(shiftedXdata[530]));
Q_MX02 U6712 ( .S(shiftCount[7]), .A0(n2935), .A1(n2807), .Z(shiftedXdata[529]));
Q_MX02 U6713 ( .S(shiftCount[7]), .A0(n2934), .A1(n2806), .Z(shiftedXdata[528]));
Q_MX02 U6714 ( .S(shiftCount[7]), .A0(n2933), .A1(n2805), .Z(shiftedXdata[527]));
Q_MX02 U6715 ( .S(shiftCount[7]), .A0(n2932), .A1(n2804), .Z(shiftedXdata[526]));
Q_MX02 U6716 ( .S(shiftCount[7]), .A0(n2931), .A1(n2803), .Z(shiftedXdata[525]));
Q_MX02 U6717 ( .S(shiftCount[7]), .A0(n2930), .A1(n2802), .Z(shiftedXdata[524]));
Q_MX02 U6718 ( .S(shiftCount[7]), .A0(n2929), .A1(n2801), .Z(shiftedXdata[523]));
Q_MX02 U6719 ( .S(shiftCount[7]), .A0(n2928), .A1(n2800), .Z(shiftedXdata[522]));
Q_MX02 U6720 ( .S(shiftCount[7]), .A0(n2927), .A1(n2799), .Z(shiftedXdata[521]));
Q_MX02 U6721 ( .S(shiftCount[7]), .A0(n2926), .A1(n2798), .Z(shiftedXdata[520]));
Q_MX02 U6722 ( .S(shiftCount[7]), .A0(n2925), .A1(n2797), .Z(shiftedXdata[519]));
Q_MX02 U6723 ( .S(shiftCount[7]), .A0(n2924), .A1(n2796), .Z(shiftedXdata[518]));
Q_MX02 U6724 ( .S(shiftCount[7]), .A0(n2923), .A1(n2795), .Z(shiftedXdata[517]));
Q_MX02 U6725 ( .S(shiftCount[7]), .A0(n2922), .A1(n2794), .Z(shiftedXdata[516]));
Q_MX02 U6726 ( .S(shiftCount[7]), .A0(n2921), .A1(n2793), .Z(shiftedXdata[515]));
Q_MX02 U6727 ( .S(shiftCount[7]), .A0(n2920), .A1(n2792), .Z(shiftedXdata[514]));
Q_MX02 U6728 ( .S(shiftCount[7]), .A0(n2919), .A1(n2791), .Z(shiftedXdata[513]));
Q_MX02 U6729 ( .S(shiftCount[7]), .A0(n2918), .A1(n2790), .Z(shiftedXdata[512]));
Q_MX02 U6730 ( .S(shiftCount[7]), .A0(n2917), .A1(n2789), .Z(shiftedXdata[511]));
Q_MX02 U6731 ( .S(shiftCount[7]), .A0(n2916), .A1(n2788), .Z(shiftedXdata[510]));
Q_MX02 U6732 ( .S(shiftCount[7]), .A0(n2915), .A1(n2787), .Z(shiftedXdata[509]));
Q_MX02 U6733 ( .S(shiftCount[7]), .A0(n2914), .A1(n2786), .Z(shiftedXdata[508]));
Q_MX02 U6734 ( .S(shiftCount[7]), .A0(n2913), .A1(n2785), .Z(shiftedXdata[507]));
Q_MX02 U6735 ( .S(shiftCount[7]), .A0(n2912), .A1(n2784), .Z(shiftedXdata[506]));
Q_MX02 U6736 ( .S(shiftCount[7]), .A0(n2911), .A1(n2783), .Z(shiftedXdata[505]));
Q_MX02 U6737 ( .S(shiftCount[7]), .A0(n2910), .A1(n2782), .Z(shiftedXdata[504]));
Q_MX02 U6738 ( .S(shiftCount[7]), .A0(n2909), .A1(n2781), .Z(shiftedXdata[503]));
Q_MX02 U6739 ( .S(shiftCount[7]), .A0(n2908), .A1(n2780), .Z(shiftedXdata[502]));
Q_MX02 U6740 ( .S(shiftCount[7]), .A0(n2907), .A1(n2779), .Z(shiftedXdata[501]));
Q_MX02 U6741 ( .S(shiftCount[7]), .A0(n2906), .A1(n2778), .Z(shiftedXdata[500]));
Q_MX02 U6742 ( .S(shiftCount[7]), .A0(n2905), .A1(n2777), .Z(shiftedXdata[499]));
Q_MX02 U6743 ( .S(shiftCount[7]), .A0(n2904), .A1(n2776), .Z(shiftedXdata[498]));
Q_MX02 U6744 ( .S(shiftCount[7]), .A0(n2903), .A1(n2775), .Z(shiftedXdata[497]));
Q_MX02 U6745 ( .S(shiftCount[7]), .A0(n2902), .A1(n2774), .Z(shiftedXdata[496]));
Q_MX02 U6746 ( .S(shiftCount[7]), .A0(n2901), .A1(n2773), .Z(shiftedXdata[495]));
Q_MX02 U6747 ( .S(shiftCount[7]), .A0(n2900), .A1(n2772), .Z(shiftedXdata[494]));
Q_MX02 U6748 ( .S(shiftCount[7]), .A0(n2899), .A1(n2771), .Z(shiftedXdata[493]));
Q_MX02 U6749 ( .S(shiftCount[7]), .A0(n2898), .A1(n2770), .Z(shiftedXdata[492]));
Q_MX02 U6750 ( .S(shiftCount[7]), .A0(n2897), .A1(n2769), .Z(shiftedXdata[491]));
Q_MX02 U6751 ( .S(shiftCount[7]), .A0(n2896), .A1(n2768), .Z(shiftedXdata[490]));
Q_MX02 U6752 ( .S(shiftCount[7]), .A0(n2895), .A1(n2767), .Z(shiftedXdata[489]));
Q_MX02 U6753 ( .S(shiftCount[7]), .A0(n2894), .A1(n2766), .Z(shiftedXdata[488]));
Q_MX02 U6754 ( .S(shiftCount[7]), .A0(n2893), .A1(n2765), .Z(shiftedXdata[487]));
Q_MX02 U6755 ( .S(shiftCount[7]), .A0(n2892), .A1(n2764), .Z(shiftedXdata[486]));
Q_MX02 U6756 ( .S(shiftCount[7]), .A0(n2891), .A1(n2763), .Z(shiftedXdata[485]));
Q_MX02 U6757 ( .S(shiftCount[7]), .A0(n2890), .A1(n2762), .Z(shiftedXdata[484]));
Q_MX02 U6758 ( .S(shiftCount[7]), .A0(n2889), .A1(n2761), .Z(shiftedXdata[483]));
Q_MX02 U6759 ( .S(shiftCount[7]), .A0(n2888), .A1(n2760), .Z(shiftedXdata[482]));
Q_MX02 U6760 ( .S(shiftCount[7]), .A0(n2887), .A1(n2759), .Z(shiftedXdata[481]));
Q_MX02 U6761 ( .S(shiftCount[7]), .A0(n2886), .A1(n2758), .Z(shiftedXdata[480]));
Q_MX02 U6762 ( .S(shiftCount[7]), .A0(n2885), .A1(n2757), .Z(shiftedXdata[479]));
Q_MX02 U6763 ( .S(shiftCount[7]), .A0(n2884), .A1(n2756), .Z(shiftedXdata[478]));
Q_MX02 U6764 ( .S(shiftCount[7]), .A0(n2883), .A1(n2755), .Z(shiftedXdata[477]));
Q_MX02 U6765 ( .S(shiftCount[7]), .A0(n2882), .A1(n2754), .Z(shiftedXdata[476]));
Q_MX02 U6766 ( .S(shiftCount[7]), .A0(n2881), .A1(n2753), .Z(shiftedXdata[475]));
Q_MX02 U6767 ( .S(shiftCount[7]), .A0(n2880), .A1(n2752), .Z(shiftedXdata[474]));
Q_MX02 U6768 ( .S(shiftCount[7]), .A0(n2879), .A1(n2751), .Z(shiftedXdata[473]));
Q_MX02 U6769 ( .S(shiftCount[7]), .A0(n2878), .A1(n2750), .Z(shiftedXdata[472]));
Q_MX02 U6770 ( .S(shiftCount[7]), .A0(n2877), .A1(n2749), .Z(shiftedXdata[471]));
Q_MX02 U6771 ( .S(shiftCount[7]), .A0(n2876), .A1(n2748), .Z(shiftedXdata[470]));
Q_MX02 U6772 ( .S(shiftCount[7]), .A0(n2875), .A1(n2747), .Z(shiftedXdata[469]));
Q_MX02 U6773 ( .S(shiftCount[7]), .A0(n2874), .A1(n2746), .Z(shiftedXdata[468]));
Q_MX02 U6774 ( .S(shiftCount[7]), .A0(n2873), .A1(n2745), .Z(shiftedXdata[467]));
Q_MX02 U6775 ( .S(shiftCount[7]), .A0(n2872), .A1(n2744), .Z(shiftedXdata[466]));
Q_MX02 U6776 ( .S(shiftCount[7]), .A0(n2871), .A1(n2743), .Z(shiftedXdata[465]));
Q_MX02 U6777 ( .S(shiftCount[7]), .A0(n2870), .A1(n2742), .Z(shiftedXdata[464]));
Q_MX02 U6778 ( .S(shiftCount[7]), .A0(n2869), .A1(n2741), .Z(shiftedXdata[463]));
Q_MX02 U6779 ( .S(shiftCount[7]), .A0(n2868), .A1(n2740), .Z(shiftedXdata[462]));
Q_MX02 U6780 ( .S(shiftCount[7]), .A0(n2867), .A1(n2739), .Z(shiftedXdata[461]));
Q_MX02 U6781 ( .S(shiftCount[7]), .A0(n2866), .A1(n2738), .Z(shiftedXdata[460]));
Q_MX02 U6782 ( .S(shiftCount[7]), .A0(n2865), .A1(n2737), .Z(shiftedXdata[459]));
Q_MX02 U6783 ( .S(shiftCount[7]), .A0(n2864), .A1(n2736), .Z(shiftedXdata[458]));
Q_MX02 U6784 ( .S(shiftCount[7]), .A0(n2863), .A1(n2735), .Z(shiftedXdata[457]));
Q_MX02 U6785 ( .S(shiftCount[7]), .A0(n2862), .A1(n2734), .Z(shiftedXdata[456]));
Q_MX02 U6786 ( .S(shiftCount[7]), .A0(n2861), .A1(n2733), .Z(shiftedXdata[455]));
Q_MX02 U6787 ( .S(shiftCount[7]), .A0(n2860), .A1(n2732), .Z(shiftedXdata[454]));
Q_MX02 U6788 ( .S(shiftCount[7]), .A0(n2859), .A1(n2731), .Z(shiftedXdata[453]));
Q_MX02 U6789 ( .S(shiftCount[7]), .A0(n2858), .A1(n2730), .Z(shiftedXdata[452]));
Q_MX02 U6790 ( .S(shiftCount[7]), .A0(n2857), .A1(n2729), .Z(shiftedXdata[451]));
Q_MX02 U6791 ( .S(shiftCount[7]), .A0(n2856), .A1(n2728), .Z(shiftedXdata[450]));
Q_MX02 U6792 ( .S(shiftCount[7]), .A0(n2855), .A1(n2727), .Z(shiftedXdata[449]));
Q_MX02 U6793 ( .S(shiftCount[7]), .A0(n2854), .A1(n2726), .Z(shiftedXdata[448]));
Q_MX02 U6794 ( .S(shiftCount[7]), .A0(n2853), .A1(n2725), .Z(shiftedXdata[447]));
Q_MX02 U6795 ( .S(shiftCount[7]), .A0(n2852), .A1(n2724), .Z(shiftedXdata[446]));
Q_MX02 U6796 ( .S(shiftCount[7]), .A0(n2851), .A1(n2723), .Z(shiftedXdata[445]));
Q_MX02 U6797 ( .S(shiftCount[7]), .A0(n2850), .A1(n2722), .Z(shiftedXdata[444]));
Q_MX02 U6798 ( .S(shiftCount[7]), .A0(n2849), .A1(n2721), .Z(shiftedXdata[443]));
Q_MX02 U6799 ( .S(shiftCount[7]), .A0(n2848), .A1(n2720), .Z(shiftedXdata[442]));
Q_MX02 U6800 ( .S(shiftCount[7]), .A0(n2847), .A1(n2719), .Z(shiftedXdata[441]));
Q_MX02 U6801 ( .S(shiftCount[7]), .A0(n2846), .A1(n2718), .Z(shiftedXdata[440]));
Q_MX02 U6802 ( .S(shiftCount[7]), .A0(n2845), .A1(n2717), .Z(shiftedXdata[439]));
Q_MX02 U6803 ( .S(shiftCount[7]), .A0(n2844), .A1(n2716), .Z(shiftedXdata[438]));
Q_MX02 U6804 ( .S(shiftCount[7]), .A0(n2843), .A1(n2715), .Z(shiftedXdata[437]));
Q_MX02 U6805 ( .S(shiftCount[7]), .A0(n2842), .A1(n2714), .Z(shiftedXdata[436]));
Q_MX02 U6806 ( .S(shiftCount[7]), .A0(n2841), .A1(n2713), .Z(shiftedXdata[435]));
Q_MX02 U6807 ( .S(shiftCount[7]), .A0(n2840), .A1(n2712), .Z(shiftedXdata[434]));
Q_MX02 U6808 ( .S(shiftCount[7]), .A0(n2839), .A1(n2711), .Z(shiftedXdata[433]));
Q_MX02 U6809 ( .S(shiftCount[7]), .A0(n2838), .A1(n2710), .Z(shiftedXdata[432]));
Q_MX02 U6810 ( .S(shiftCount[7]), .A0(n2837), .A1(n2709), .Z(shiftedXdata[431]));
Q_MX02 U6811 ( .S(shiftCount[7]), .A0(n2836), .A1(n2708), .Z(shiftedXdata[430]));
Q_MX02 U6812 ( .S(shiftCount[7]), .A0(n2835), .A1(n2707), .Z(shiftedXdata[429]));
Q_MX02 U6813 ( .S(shiftCount[7]), .A0(n2834), .A1(n2706), .Z(shiftedXdata[428]));
Q_MX02 U6814 ( .S(shiftCount[7]), .A0(n2833), .A1(n2705), .Z(shiftedXdata[427]));
Q_MX02 U6815 ( .S(shiftCount[7]), .A0(n2832), .A1(n2704), .Z(shiftedXdata[426]));
Q_MX02 U6816 ( .S(shiftCount[7]), .A0(n2831), .A1(n2703), .Z(shiftedXdata[425]));
Q_MX02 U6817 ( .S(shiftCount[7]), .A0(n2830), .A1(n2702), .Z(shiftedXdata[424]));
Q_MX02 U6818 ( .S(shiftCount[7]), .A0(n2829), .A1(n2701), .Z(shiftedXdata[423]));
Q_MX02 U6819 ( .S(shiftCount[7]), .A0(n2828), .A1(n2700), .Z(shiftedXdata[422]));
Q_MX02 U6820 ( .S(shiftCount[7]), .A0(n2827), .A1(n2699), .Z(shiftedXdata[421]));
Q_MX02 U6821 ( .S(shiftCount[7]), .A0(n2826), .A1(n2698), .Z(shiftedXdata[420]));
Q_MX02 U6822 ( .S(shiftCount[7]), .A0(n2825), .A1(n2697), .Z(shiftedXdata[419]));
Q_MX02 U6823 ( .S(shiftCount[7]), .A0(n2824), .A1(n2696), .Z(shiftedXdata[418]));
Q_MX02 U6824 ( .S(shiftCount[7]), .A0(n2823), .A1(n2695), .Z(shiftedXdata[417]));
Q_MX02 U6825 ( .S(shiftCount[7]), .A0(n2822), .A1(n2694), .Z(shiftedXdata[416]));
Q_MX02 U6826 ( .S(shiftCount[7]), .A0(n2821), .A1(n2693), .Z(shiftedXdata[415]));
Q_MX02 U6827 ( .S(shiftCount[7]), .A0(n2820), .A1(n2692), .Z(shiftedXdata[414]));
Q_MX02 U6828 ( .S(shiftCount[7]), .A0(n2819), .A1(n2691), .Z(shiftedXdata[413]));
Q_MX02 U6829 ( .S(shiftCount[7]), .A0(n2818), .A1(n2690), .Z(shiftedXdata[412]));
Q_MX02 U6830 ( .S(shiftCount[7]), .A0(n2817), .A1(n2689), .Z(shiftedXdata[411]));
Q_MX02 U6831 ( .S(shiftCount[7]), .A0(n2816), .A1(n2688), .Z(shiftedXdata[410]));
Q_MX02 U6832 ( .S(shiftCount[7]), .A0(n2815), .A1(n2687), .Z(shiftedXdata[409]));
Q_MX02 U6833 ( .S(shiftCount[7]), .A0(n2814), .A1(n2686), .Z(shiftedXdata[408]));
Q_MX02 U6834 ( .S(shiftCount[7]), .A0(n2813), .A1(n2685), .Z(shiftedXdata[407]));
Q_MX02 U6835 ( .S(shiftCount[7]), .A0(n2812), .A1(n2684), .Z(shiftedXdata[406]));
Q_MX02 U6836 ( .S(shiftCount[7]), .A0(n2811), .A1(n2683), .Z(shiftedXdata[405]));
Q_MX02 U6837 ( .S(shiftCount[7]), .A0(n2810), .A1(n2682), .Z(shiftedXdata[404]));
Q_MX02 U6838 ( .S(shiftCount[7]), .A0(n2809), .A1(n2681), .Z(shiftedXdata[403]));
Q_MX02 U6839 ( .S(shiftCount[7]), .A0(n2808), .A1(n2680), .Z(shiftedXdata[402]));
Q_MX02 U6840 ( .S(shiftCount[7]), .A0(n2807), .A1(n2679), .Z(shiftedXdata[401]));
Q_MX02 U6841 ( .S(shiftCount[7]), .A0(n2806), .A1(n2678), .Z(shiftedXdata[400]));
Q_MX02 U6842 ( .S(shiftCount[7]), .A0(n2805), .A1(n2677), .Z(shiftedXdata[399]));
Q_MX02 U6843 ( .S(shiftCount[7]), .A0(n2804), .A1(n2676), .Z(shiftedXdata[398]));
Q_MX02 U6844 ( .S(shiftCount[7]), .A0(n2803), .A1(n2675), .Z(shiftedXdata[397]));
Q_MX02 U6845 ( .S(shiftCount[7]), .A0(n2802), .A1(n2674), .Z(shiftedXdata[396]));
Q_MX02 U6846 ( .S(shiftCount[7]), .A0(n2801), .A1(n2673), .Z(shiftedXdata[395]));
Q_MX02 U6847 ( .S(shiftCount[7]), .A0(n2800), .A1(n2672), .Z(shiftedXdata[394]));
Q_MX02 U6848 ( .S(shiftCount[7]), .A0(n2799), .A1(n2671), .Z(shiftedXdata[393]));
Q_MX02 U6849 ( .S(shiftCount[7]), .A0(n2798), .A1(n2670), .Z(shiftedXdata[392]));
Q_MX02 U6850 ( .S(shiftCount[7]), .A0(n2797), .A1(n2669), .Z(shiftedXdata[391]));
Q_MX02 U6851 ( .S(shiftCount[7]), .A0(n2796), .A1(n2668), .Z(shiftedXdata[390]));
Q_MX02 U6852 ( .S(shiftCount[7]), .A0(n2795), .A1(n2667), .Z(shiftedXdata[389]));
Q_MX02 U6853 ( .S(shiftCount[7]), .A0(n2794), .A1(n2666), .Z(shiftedXdata[388]));
Q_MX02 U6854 ( .S(shiftCount[7]), .A0(n2793), .A1(n2665), .Z(shiftedXdata[387]));
Q_MX02 U6855 ( .S(shiftCount[7]), .A0(n2792), .A1(n2664), .Z(shiftedXdata[386]));
Q_MX02 U6856 ( .S(shiftCount[7]), .A0(n2791), .A1(n2663), .Z(shiftedXdata[385]));
Q_MX02 U6857 ( .S(shiftCount[7]), .A0(n2790), .A1(n2662), .Z(shiftedXdata[384]));
Q_MX02 U6858 ( .S(shiftCount[7]), .A0(n2789), .A1(n2661), .Z(shiftedXdata[383]));
Q_MX02 U6859 ( .S(shiftCount[7]), .A0(n2788), .A1(n2660), .Z(shiftedXdata[382]));
Q_MX02 U6860 ( .S(shiftCount[7]), .A0(n2787), .A1(n2659), .Z(shiftedXdata[381]));
Q_MX02 U6861 ( .S(shiftCount[7]), .A0(n2786), .A1(n2658), .Z(shiftedXdata[380]));
Q_MX02 U6862 ( .S(shiftCount[7]), .A0(n2785), .A1(n2657), .Z(shiftedXdata[379]));
Q_MX02 U6863 ( .S(shiftCount[7]), .A0(n2784), .A1(n2656), .Z(shiftedXdata[378]));
Q_MX02 U6864 ( .S(shiftCount[7]), .A0(n2783), .A1(n2655), .Z(shiftedXdata[377]));
Q_MX02 U6865 ( .S(shiftCount[7]), .A0(n2782), .A1(n2654), .Z(shiftedXdata[376]));
Q_MX02 U6866 ( .S(shiftCount[7]), .A0(n2781), .A1(n2653), .Z(shiftedXdata[375]));
Q_MX02 U6867 ( .S(shiftCount[7]), .A0(n2780), .A1(n2652), .Z(shiftedXdata[374]));
Q_MX02 U6868 ( .S(shiftCount[7]), .A0(n2779), .A1(n2651), .Z(shiftedXdata[373]));
Q_MX02 U6869 ( .S(shiftCount[7]), .A0(n2778), .A1(n2650), .Z(shiftedXdata[372]));
Q_MX02 U6870 ( .S(shiftCount[7]), .A0(n2777), .A1(n2649), .Z(shiftedXdata[371]));
Q_MX02 U6871 ( .S(shiftCount[7]), .A0(n2776), .A1(n2648), .Z(shiftedXdata[370]));
Q_MX02 U6872 ( .S(shiftCount[7]), .A0(n2775), .A1(n2647), .Z(shiftedXdata[369]));
Q_MX02 U6873 ( .S(shiftCount[7]), .A0(n2774), .A1(n2646), .Z(shiftedXdata[368]));
Q_MX02 U6874 ( .S(shiftCount[7]), .A0(n2773), .A1(n2645), .Z(shiftedXdata[367]));
Q_MX02 U6875 ( .S(shiftCount[7]), .A0(n2772), .A1(n2644), .Z(shiftedXdata[366]));
Q_MX02 U6876 ( .S(shiftCount[7]), .A0(n2771), .A1(n2643), .Z(shiftedXdata[365]));
Q_MX02 U6877 ( .S(shiftCount[7]), .A0(n2770), .A1(n2642), .Z(shiftedXdata[364]));
Q_MX02 U6878 ( .S(shiftCount[7]), .A0(n2769), .A1(n2641), .Z(shiftedXdata[363]));
Q_MX02 U6879 ( .S(shiftCount[7]), .A0(n2768), .A1(n2640), .Z(shiftedXdata[362]));
Q_MX02 U6880 ( .S(shiftCount[7]), .A0(n2767), .A1(n2639), .Z(shiftedXdata[361]));
Q_MX02 U6881 ( .S(shiftCount[7]), .A0(n2766), .A1(n2638), .Z(shiftedXdata[360]));
Q_MX02 U6882 ( .S(shiftCount[7]), .A0(n2765), .A1(n2637), .Z(shiftedXdata[359]));
Q_MX02 U6883 ( .S(shiftCount[7]), .A0(n2764), .A1(n2636), .Z(shiftedXdata[358]));
Q_MX02 U6884 ( .S(shiftCount[7]), .A0(n2763), .A1(n2635), .Z(shiftedXdata[357]));
Q_MX02 U6885 ( .S(shiftCount[7]), .A0(n2762), .A1(n2634), .Z(shiftedXdata[356]));
Q_MX02 U6886 ( .S(shiftCount[7]), .A0(n2761), .A1(n2633), .Z(shiftedXdata[355]));
Q_MX02 U6887 ( .S(shiftCount[7]), .A0(n2760), .A1(n2632), .Z(shiftedXdata[354]));
Q_MX02 U6888 ( .S(shiftCount[7]), .A0(n2759), .A1(n2631), .Z(shiftedXdata[353]));
Q_MX02 U6889 ( .S(shiftCount[7]), .A0(n2758), .A1(n2630), .Z(shiftedXdata[352]));
Q_MX02 U6890 ( .S(shiftCount[7]), .A0(n2757), .A1(n2629), .Z(shiftedXdata[351]));
Q_MX02 U6891 ( .S(shiftCount[7]), .A0(n2756), .A1(n2628), .Z(shiftedXdata[350]));
Q_MX02 U6892 ( .S(shiftCount[7]), .A0(n2755), .A1(n2627), .Z(shiftedXdata[349]));
Q_MX02 U6893 ( .S(shiftCount[7]), .A0(n2754), .A1(n2626), .Z(shiftedXdata[348]));
Q_MX02 U6894 ( .S(shiftCount[7]), .A0(n2753), .A1(n2625), .Z(shiftedXdata[347]));
Q_MX02 U6895 ( .S(shiftCount[7]), .A0(n2752), .A1(n2624), .Z(shiftedXdata[346]));
Q_MX02 U6896 ( .S(shiftCount[7]), .A0(n2751), .A1(n2623), .Z(shiftedXdata[345]));
Q_MX02 U6897 ( .S(shiftCount[7]), .A0(n2750), .A1(n2622), .Z(shiftedXdata[344]));
Q_MX02 U6898 ( .S(shiftCount[7]), .A0(n2749), .A1(n2621), .Z(shiftedXdata[343]));
Q_MX02 U6899 ( .S(shiftCount[7]), .A0(n2748), .A1(n2620), .Z(shiftedXdata[342]));
Q_MX02 U6900 ( .S(shiftCount[7]), .A0(n2747), .A1(n2619), .Z(shiftedXdata[341]));
Q_MX02 U6901 ( .S(shiftCount[7]), .A0(n2746), .A1(n2618), .Z(shiftedXdata[340]));
Q_MX02 U6902 ( .S(shiftCount[7]), .A0(n2745), .A1(n2617), .Z(shiftedXdata[339]));
Q_MX02 U6903 ( .S(shiftCount[7]), .A0(n2744), .A1(n2616), .Z(shiftedXdata[338]));
Q_MX02 U6904 ( .S(shiftCount[7]), .A0(n2743), .A1(n2615), .Z(shiftedXdata[337]));
Q_MX02 U6905 ( .S(shiftCount[7]), .A0(n2742), .A1(n2614), .Z(shiftedXdata[336]));
Q_MX02 U6906 ( .S(shiftCount[7]), .A0(n2741), .A1(n2613), .Z(shiftedXdata[335]));
Q_MX02 U6907 ( .S(shiftCount[7]), .A0(n2740), .A1(n2612), .Z(shiftedXdata[334]));
Q_MX02 U6908 ( .S(shiftCount[7]), .A0(n2739), .A1(n2611), .Z(shiftedXdata[333]));
Q_MX02 U6909 ( .S(shiftCount[7]), .A0(n2738), .A1(n2610), .Z(shiftedXdata[332]));
Q_MX02 U6910 ( .S(shiftCount[7]), .A0(n2737), .A1(n2609), .Z(shiftedXdata[331]));
Q_MX02 U6911 ( .S(shiftCount[7]), .A0(n2736), .A1(n2608), .Z(shiftedXdata[330]));
Q_MX02 U6912 ( .S(shiftCount[7]), .A0(n2735), .A1(n2607), .Z(shiftedXdata[329]));
Q_MX02 U6913 ( .S(shiftCount[7]), .A0(n2734), .A1(n2606), .Z(shiftedXdata[328]));
Q_MX02 U6914 ( .S(shiftCount[7]), .A0(n2733), .A1(n2605), .Z(shiftedXdata[327]));
Q_MX02 U6915 ( .S(shiftCount[7]), .A0(n2732), .A1(n2604), .Z(shiftedXdata[326]));
Q_MX02 U6916 ( .S(shiftCount[7]), .A0(n2731), .A1(n2603), .Z(shiftedXdata[325]));
Q_MX02 U6917 ( .S(shiftCount[7]), .A0(n2730), .A1(n2602), .Z(shiftedXdata[324]));
Q_MX02 U6918 ( .S(shiftCount[7]), .A0(n2729), .A1(n2601), .Z(shiftedXdata[323]));
Q_MX02 U6919 ( .S(shiftCount[7]), .A0(n2728), .A1(n2600), .Z(shiftedXdata[322]));
Q_MX02 U6920 ( .S(shiftCount[7]), .A0(n2727), .A1(n2599), .Z(shiftedXdata[321]));
Q_MX02 U6921 ( .S(shiftCount[7]), .A0(n2726), .A1(n2598), .Z(shiftedXdata[320]));
Q_MX02 U6922 ( .S(shiftCount[7]), .A0(n2725), .A1(n2597), .Z(shiftedXdata[319]));
Q_MX02 U6923 ( .S(shiftCount[7]), .A0(n2724), .A1(n2596), .Z(shiftedXdata[318]));
Q_MX02 U6924 ( .S(shiftCount[7]), .A0(n2723), .A1(n2595), .Z(shiftedXdata[317]));
Q_MX02 U6925 ( .S(shiftCount[7]), .A0(n2722), .A1(n2594), .Z(shiftedXdata[316]));
Q_MX02 U6926 ( .S(shiftCount[7]), .A0(n2721), .A1(n2593), .Z(shiftedXdata[315]));
Q_MX02 U6927 ( .S(shiftCount[7]), .A0(n2720), .A1(n2592), .Z(shiftedXdata[314]));
Q_MX02 U6928 ( .S(shiftCount[7]), .A0(n2719), .A1(n2591), .Z(shiftedXdata[313]));
Q_MX02 U6929 ( .S(shiftCount[7]), .A0(n2718), .A1(n2590), .Z(shiftedXdata[312]));
Q_MX02 U6930 ( .S(shiftCount[7]), .A0(n2717), .A1(n2589), .Z(shiftedXdata[311]));
Q_MX02 U6931 ( .S(shiftCount[7]), .A0(n2716), .A1(n2588), .Z(shiftedXdata[310]));
Q_MX02 U6932 ( .S(shiftCount[7]), .A0(n2715), .A1(n2587), .Z(shiftedXdata[309]));
Q_MX02 U6933 ( .S(shiftCount[7]), .A0(n2714), .A1(n2586), .Z(shiftedXdata[308]));
Q_MX02 U6934 ( .S(shiftCount[7]), .A0(n2713), .A1(n2585), .Z(shiftedXdata[307]));
Q_MX02 U6935 ( .S(shiftCount[7]), .A0(n2712), .A1(n2584), .Z(shiftedXdata[306]));
Q_MX02 U6936 ( .S(shiftCount[7]), .A0(n2711), .A1(n2583), .Z(shiftedXdata[305]));
Q_MX02 U6937 ( .S(shiftCount[7]), .A0(n2710), .A1(n2582), .Z(shiftedXdata[304]));
Q_MX02 U6938 ( .S(shiftCount[7]), .A0(n2709), .A1(n2581), .Z(shiftedXdata[303]));
Q_MX02 U6939 ( .S(shiftCount[7]), .A0(n2708), .A1(n2580), .Z(shiftedXdata[302]));
Q_MX02 U6940 ( .S(shiftCount[7]), .A0(n2707), .A1(n2579), .Z(shiftedXdata[301]));
Q_MX02 U6941 ( .S(shiftCount[7]), .A0(n2706), .A1(n2578), .Z(shiftedXdata[300]));
Q_MX02 U6942 ( .S(shiftCount[7]), .A0(n2705), .A1(n2577), .Z(shiftedXdata[299]));
Q_MX02 U6943 ( .S(shiftCount[7]), .A0(n2704), .A1(n2576), .Z(shiftedXdata[298]));
Q_MX02 U6944 ( .S(shiftCount[7]), .A0(n2703), .A1(n2575), .Z(shiftedXdata[297]));
Q_MX02 U6945 ( .S(shiftCount[7]), .A0(n2702), .A1(n2574), .Z(shiftedXdata[296]));
Q_MX02 U6946 ( .S(shiftCount[7]), .A0(n2701), .A1(n2573), .Z(shiftedXdata[295]));
Q_MX02 U6947 ( .S(shiftCount[7]), .A0(n2700), .A1(n2572), .Z(shiftedXdata[294]));
Q_MX02 U6948 ( .S(shiftCount[7]), .A0(n2699), .A1(n2571), .Z(shiftedXdata[293]));
Q_MX02 U6949 ( .S(shiftCount[7]), .A0(n2698), .A1(n2570), .Z(shiftedXdata[292]));
Q_MX02 U6950 ( .S(shiftCount[7]), .A0(n2697), .A1(n2569), .Z(shiftedXdata[291]));
Q_MX02 U6951 ( .S(shiftCount[7]), .A0(n2696), .A1(n2568), .Z(shiftedXdata[290]));
Q_MX02 U6952 ( .S(shiftCount[7]), .A0(n2695), .A1(n2567), .Z(shiftedXdata[289]));
Q_MX02 U6953 ( .S(shiftCount[7]), .A0(n2694), .A1(n2566), .Z(shiftedXdata[288]));
Q_MX02 U6954 ( .S(shiftCount[7]), .A0(n2693), .A1(n2565), .Z(shiftedXdata[287]));
Q_MX02 U6955 ( .S(shiftCount[7]), .A0(n2692), .A1(n2564), .Z(shiftedXdata[286]));
Q_MX02 U6956 ( .S(shiftCount[7]), .A0(n2691), .A1(n2563), .Z(shiftedXdata[285]));
Q_MX02 U6957 ( .S(shiftCount[7]), .A0(n2690), .A1(n2562), .Z(shiftedXdata[284]));
Q_MX02 U6958 ( .S(shiftCount[7]), .A0(n2689), .A1(n2561), .Z(shiftedXdata[283]));
Q_MX02 U6959 ( .S(shiftCount[7]), .A0(n2688), .A1(n2560), .Z(shiftedXdata[282]));
Q_MX02 U6960 ( .S(shiftCount[7]), .A0(n2687), .A1(n2559), .Z(shiftedXdata[281]));
Q_MX02 U6961 ( .S(shiftCount[7]), .A0(n2686), .A1(n2558), .Z(shiftedXdata[280]));
Q_MX02 U6962 ( .S(shiftCount[7]), .A0(n2685), .A1(n2557), .Z(shiftedXdata[279]));
Q_MX02 U6963 ( .S(shiftCount[7]), .A0(n2684), .A1(n2556), .Z(shiftedXdata[278]));
Q_MX02 U6964 ( .S(shiftCount[7]), .A0(n2683), .A1(n2555), .Z(shiftedXdata[277]));
Q_MX02 U6965 ( .S(shiftCount[7]), .A0(n2682), .A1(n2554), .Z(shiftedXdata[276]));
Q_MX02 U6966 ( .S(shiftCount[7]), .A0(n2681), .A1(n2553), .Z(shiftedXdata[275]));
Q_MX02 U6967 ( .S(shiftCount[7]), .A0(n2680), .A1(n2552), .Z(shiftedXdata[274]));
Q_MX02 U6968 ( .S(shiftCount[7]), .A0(n2679), .A1(n2551), .Z(shiftedXdata[273]));
Q_MX02 U6969 ( .S(shiftCount[7]), .A0(n2678), .A1(n2550), .Z(shiftedXdata[272]));
Q_MX02 U6970 ( .S(shiftCount[7]), .A0(n2677), .A1(n2549), .Z(shiftedXdata[271]));
Q_MX02 U6971 ( .S(shiftCount[7]), .A0(n2676), .A1(n2548), .Z(shiftedXdata[270]));
Q_MX02 U6972 ( .S(shiftCount[7]), .A0(n2675), .A1(n2547), .Z(shiftedXdata[269]));
Q_MX02 U6973 ( .S(shiftCount[7]), .A0(n2674), .A1(n2546), .Z(shiftedXdata[268]));
Q_MX02 U6974 ( .S(shiftCount[7]), .A0(n2673), .A1(n2545), .Z(shiftedXdata[267]));
Q_MX02 U6975 ( .S(shiftCount[7]), .A0(n2672), .A1(n2544), .Z(shiftedXdata[266]));
Q_MX02 U6976 ( .S(shiftCount[7]), .A0(n2671), .A1(n2543), .Z(shiftedXdata[265]));
Q_MX02 U6977 ( .S(shiftCount[7]), .A0(n2670), .A1(n2542), .Z(shiftedXdata[264]));
Q_MX02 U6978 ( .S(shiftCount[7]), .A0(n2669), .A1(n2541), .Z(shiftedXdata[263]));
Q_MX02 U6979 ( .S(shiftCount[7]), .A0(n2668), .A1(n2540), .Z(shiftedXdata[262]));
Q_MX02 U6980 ( .S(shiftCount[7]), .A0(n2667), .A1(n2539), .Z(shiftedXdata[261]));
Q_MX02 U6981 ( .S(shiftCount[7]), .A0(n2666), .A1(n2538), .Z(shiftedXdata[260]));
Q_MX02 U6982 ( .S(shiftCount[7]), .A0(n2665), .A1(n2537), .Z(shiftedXdata[259]));
Q_MX02 U6983 ( .S(shiftCount[7]), .A0(n2664), .A1(n2536), .Z(shiftedXdata[258]));
Q_MX02 U6984 ( .S(shiftCount[7]), .A0(n2663), .A1(n2535), .Z(shiftedXdata[257]));
Q_MX02 U6985 ( .S(shiftCount[7]), .A0(n2662), .A1(n2534), .Z(shiftedXdata[256]));
Q_MX02 U6986 ( .S(shiftCount[7]), .A0(n2661), .A1(n2533), .Z(shiftedXdata[255]));
Q_MX02 U6987 ( .S(shiftCount[7]), .A0(n2660), .A1(n2532), .Z(shiftedXdata[254]));
Q_MX02 U6988 ( .S(shiftCount[7]), .A0(n2659), .A1(n2531), .Z(shiftedXdata[253]));
Q_MX02 U6989 ( .S(shiftCount[7]), .A0(n2658), .A1(n2530), .Z(shiftedXdata[252]));
Q_MX02 U6990 ( .S(shiftCount[7]), .A0(n2657), .A1(n2529), .Z(shiftedXdata[251]));
Q_MX02 U6991 ( .S(shiftCount[7]), .A0(n2656), .A1(n2528), .Z(shiftedXdata[250]));
Q_MX02 U6992 ( .S(shiftCount[7]), .A0(n2655), .A1(n2527), .Z(shiftedXdata[249]));
Q_MX02 U6993 ( .S(shiftCount[7]), .A0(n2654), .A1(n2526), .Z(shiftedXdata[248]));
Q_MX02 U6994 ( .S(shiftCount[7]), .A0(n2653), .A1(n2525), .Z(shiftedXdata[247]));
Q_MX02 U6995 ( .S(shiftCount[7]), .A0(n2652), .A1(n2524), .Z(shiftedXdata[246]));
Q_MX02 U6996 ( .S(shiftCount[7]), .A0(n2651), .A1(n2523), .Z(shiftedXdata[245]));
Q_MX02 U6997 ( .S(shiftCount[7]), .A0(n2650), .A1(n2522), .Z(shiftedXdata[244]));
Q_MX02 U6998 ( .S(shiftCount[7]), .A0(n2649), .A1(n2521), .Z(shiftedXdata[243]));
Q_MX02 U6999 ( .S(shiftCount[7]), .A0(n2648), .A1(n2520), .Z(shiftedXdata[242]));
Q_MX02 U7000 ( .S(shiftCount[7]), .A0(n2647), .A1(n2519), .Z(shiftedXdata[241]));
Q_MX02 U7001 ( .S(shiftCount[7]), .A0(n2646), .A1(n2518), .Z(shiftedXdata[240]));
Q_MX02 U7002 ( .S(shiftCount[7]), .A0(n2645), .A1(n2517), .Z(shiftedXdata[239]));
Q_MX02 U7003 ( .S(shiftCount[7]), .A0(n2644), .A1(n2516), .Z(shiftedXdata[238]));
Q_MX02 U7004 ( .S(shiftCount[7]), .A0(n2643), .A1(n2515), .Z(shiftedXdata[237]));
Q_MX02 U7005 ( .S(shiftCount[7]), .A0(n2642), .A1(n2514), .Z(shiftedXdata[236]));
Q_MX02 U7006 ( .S(shiftCount[7]), .A0(n2641), .A1(n2513), .Z(shiftedXdata[235]));
Q_MX02 U7007 ( .S(shiftCount[7]), .A0(n2640), .A1(n2512), .Z(shiftedXdata[234]));
Q_MX02 U7008 ( .S(shiftCount[7]), .A0(n2639), .A1(n2511), .Z(shiftedXdata[233]));
Q_MX02 U7009 ( .S(shiftCount[7]), .A0(n2638), .A1(n2510), .Z(shiftedXdata[232]));
Q_MX02 U7010 ( .S(shiftCount[7]), .A0(n2637), .A1(n2509), .Z(shiftedXdata[231]));
Q_MX02 U7011 ( .S(shiftCount[7]), .A0(n2636), .A1(n2508), .Z(shiftedXdata[230]));
Q_MX02 U7012 ( .S(shiftCount[7]), .A0(n2635), .A1(n2507), .Z(shiftedXdata[229]));
Q_MX02 U7013 ( .S(shiftCount[7]), .A0(n2634), .A1(n2506), .Z(shiftedXdata[228]));
Q_MX02 U7014 ( .S(shiftCount[7]), .A0(n2633), .A1(n2505), .Z(shiftedXdata[227]));
Q_MX02 U7015 ( .S(shiftCount[7]), .A0(n2632), .A1(n2504), .Z(shiftedXdata[226]));
Q_MX02 U7016 ( .S(shiftCount[7]), .A0(n2631), .A1(n2503), .Z(shiftedXdata[225]));
Q_MX02 U7017 ( .S(shiftCount[7]), .A0(n2630), .A1(n2502), .Z(shiftedXdata[224]));
Q_MX02 U7018 ( .S(shiftCount[7]), .A0(n2629), .A1(n2501), .Z(shiftedXdata[223]));
Q_MX02 U7019 ( .S(shiftCount[7]), .A0(n2628), .A1(n2500), .Z(shiftedXdata[222]));
Q_MX02 U7020 ( .S(shiftCount[7]), .A0(n2627), .A1(n2499), .Z(shiftedXdata[221]));
Q_MX02 U7021 ( .S(shiftCount[7]), .A0(n2626), .A1(n2498), .Z(shiftedXdata[220]));
Q_MX02 U7022 ( .S(shiftCount[7]), .A0(n2625), .A1(n2497), .Z(shiftedXdata[219]));
Q_MX02 U7023 ( .S(shiftCount[7]), .A0(n2624), .A1(n2496), .Z(shiftedXdata[218]));
Q_MX02 U7024 ( .S(shiftCount[7]), .A0(n2623), .A1(n2495), .Z(shiftedXdata[217]));
Q_MX02 U7025 ( .S(shiftCount[7]), .A0(n2622), .A1(n2494), .Z(shiftedXdata[216]));
Q_MX02 U7026 ( .S(shiftCount[7]), .A0(n2621), .A1(n2493), .Z(shiftedXdata[215]));
Q_MX02 U7027 ( .S(shiftCount[7]), .A0(n2620), .A1(n2492), .Z(shiftedXdata[214]));
Q_MX02 U7028 ( .S(shiftCount[7]), .A0(n2619), .A1(n2491), .Z(shiftedXdata[213]));
Q_MX02 U7029 ( .S(shiftCount[7]), .A0(n2618), .A1(n2490), .Z(shiftedXdata[212]));
Q_MX02 U7030 ( .S(shiftCount[7]), .A0(n2617), .A1(n2489), .Z(shiftedXdata[211]));
Q_MX02 U7031 ( .S(shiftCount[7]), .A0(n2616), .A1(n2488), .Z(shiftedXdata[210]));
Q_MX02 U7032 ( .S(shiftCount[7]), .A0(n2615), .A1(n2487), .Z(shiftedXdata[209]));
Q_MX02 U7033 ( .S(shiftCount[7]), .A0(n2614), .A1(n2486), .Z(shiftedXdata[208]));
Q_MX02 U7034 ( .S(shiftCount[7]), .A0(n2613), .A1(n2485), .Z(shiftedXdata[207]));
Q_MX02 U7035 ( .S(shiftCount[7]), .A0(n2612), .A1(n2484), .Z(shiftedXdata[206]));
Q_MX02 U7036 ( .S(shiftCount[7]), .A0(n2611), .A1(n2483), .Z(shiftedXdata[205]));
Q_MX02 U7037 ( .S(shiftCount[7]), .A0(n2610), .A1(n2482), .Z(shiftedXdata[204]));
Q_MX02 U7038 ( .S(shiftCount[7]), .A0(n2609), .A1(n2481), .Z(shiftedXdata[203]));
Q_MX02 U7039 ( .S(shiftCount[7]), .A0(n2608), .A1(n2480), .Z(shiftedXdata[202]));
Q_MX02 U7040 ( .S(shiftCount[7]), .A0(n2607), .A1(n2479), .Z(shiftedXdata[201]));
Q_MX02 U7041 ( .S(shiftCount[7]), .A0(n2606), .A1(n2478), .Z(shiftedXdata[200]));
Q_MX02 U7042 ( .S(shiftCount[7]), .A0(n2605), .A1(n2477), .Z(shiftedXdata[199]));
Q_MX02 U7043 ( .S(shiftCount[7]), .A0(n2604), .A1(n2476), .Z(shiftedXdata[198]));
Q_MX02 U7044 ( .S(shiftCount[7]), .A0(n2603), .A1(n2475), .Z(shiftedXdata[197]));
Q_MX02 U7045 ( .S(shiftCount[7]), .A0(n2602), .A1(n2474), .Z(shiftedXdata[196]));
Q_MX02 U7046 ( .S(shiftCount[7]), .A0(n2601), .A1(n2473), .Z(shiftedXdata[195]));
Q_MX02 U7047 ( .S(shiftCount[7]), .A0(n2600), .A1(n2472), .Z(shiftedXdata[194]));
Q_MX02 U7048 ( .S(shiftCount[7]), .A0(n2599), .A1(n2471), .Z(shiftedXdata[193]));
Q_MX02 U7049 ( .S(shiftCount[7]), .A0(n2598), .A1(n2470), .Z(shiftedXdata[192]));
Q_MX02 U7050 ( .S(shiftCount[7]), .A0(n2597), .A1(n2468), .Z(shiftedXdata[191]));
Q_MX02 U7051 ( .S(shiftCount[7]), .A0(n2596), .A1(n2467), .Z(shiftedXdata[190]));
Q_MX02 U7052 ( .S(shiftCount[7]), .A0(n2595), .A1(n2466), .Z(shiftedXdata[189]));
Q_MX02 U7053 ( .S(shiftCount[7]), .A0(n2594), .A1(n2465), .Z(shiftedXdata[188]));
Q_MX02 U7054 ( .S(shiftCount[7]), .A0(n2593), .A1(n2464), .Z(shiftedXdata[187]));
Q_MX02 U7055 ( .S(shiftCount[7]), .A0(n2592), .A1(n2463), .Z(shiftedXdata[186]));
Q_MX02 U7056 ( .S(shiftCount[7]), .A0(n2591), .A1(n2462), .Z(shiftedXdata[185]));
Q_MX02 U7057 ( .S(shiftCount[7]), .A0(n2590), .A1(n2461), .Z(shiftedXdata[184]));
Q_MX02 U7058 ( .S(shiftCount[7]), .A0(n2589), .A1(n2460), .Z(shiftedXdata[183]));
Q_MX02 U7059 ( .S(shiftCount[7]), .A0(n2588), .A1(n2459), .Z(shiftedXdata[182]));
Q_MX02 U7060 ( .S(shiftCount[7]), .A0(n2587), .A1(n2458), .Z(shiftedXdata[181]));
Q_MX02 U7061 ( .S(shiftCount[7]), .A0(n2586), .A1(n2457), .Z(shiftedXdata[180]));
Q_MX02 U7062 ( .S(shiftCount[7]), .A0(n2585), .A1(n2456), .Z(shiftedXdata[179]));
Q_MX02 U7063 ( .S(shiftCount[7]), .A0(n2584), .A1(n2455), .Z(shiftedXdata[178]));
Q_MX02 U7064 ( .S(shiftCount[7]), .A0(n2583), .A1(n2454), .Z(shiftedXdata[177]));
Q_MX02 U7065 ( .S(shiftCount[7]), .A0(n2582), .A1(n2453), .Z(shiftedXdata[176]));
Q_MX02 U7066 ( .S(shiftCount[7]), .A0(n2581), .A1(n2452), .Z(shiftedXdata[175]));
Q_MX02 U7067 ( .S(shiftCount[7]), .A0(n2580), .A1(n2451), .Z(shiftedXdata[174]));
Q_MX02 U7068 ( .S(shiftCount[7]), .A0(n2579), .A1(n2450), .Z(shiftedXdata[173]));
Q_MX02 U7069 ( .S(shiftCount[7]), .A0(n2578), .A1(n2449), .Z(shiftedXdata[172]));
Q_MX02 U7070 ( .S(shiftCount[7]), .A0(n2577), .A1(n2448), .Z(shiftedXdata[171]));
Q_MX02 U7071 ( .S(shiftCount[7]), .A0(n2576), .A1(n2447), .Z(shiftedXdata[170]));
Q_MX02 U7072 ( .S(shiftCount[7]), .A0(n2575), .A1(n2446), .Z(shiftedXdata[169]));
Q_MX02 U7073 ( .S(shiftCount[7]), .A0(n2574), .A1(n2445), .Z(shiftedXdata[168]));
Q_MX02 U7074 ( .S(shiftCount[7]), .A0(n2573), .A1(n2444), .Z(shiftedXdata[167]));
Q_MX02 U7075 ( .S(shiftCount[7]), .A0(n2572), .A1(n2443), .Z(shiftedXdata[166]));
Q_MX02 U7076 ( .S(shiftCount[7]), .A0(n2571), .A1(n2442), .Z(shiftedXdata[165]));
Q_MX02 U7077 ( .S(shiftCount[7]), .A0(n2570), .A1(n2441), .Z(shiftedXdata[164]));
Q_MX02 U7078 ( .S(shiftCount[7]), .A0(n2569), .A1(n2440), .Z(shiftedXdata[163]));
Q_MX02 U7079 ( .S(shiftCount[7]), .A0(n2568), .A1(n2439), .Z(shiftedXdata[162]));
Q_MX02 U7080 ( .S(shiftCount[7]), .A0(n2567), .A1(n2438), .Z(shiftedXdata[161]));
Q_MX02 U7081 ( .S(shiftCount[7]), .A0(n2566), .A1(n2437), .Z(shiftedXdata[160]));
Q_MX02 U7082 ( .S(shiftCount[7]), .A0(n2565), .A1(n2436), .Z(shiftedXdata[159]));
Q_MX02 U7083 ( .S(shiftCount[7]), .A0(n2564), .A1(n2435), .Z(shiftedXdata[158]));
Q_MX02 U7084 ( .S(shiftCount[7]), .A0(n2563), .A1(n2434), .Z(shiftedXdata[157]));
Q_MX02 U7085 ( .S(shiftCount[7]), .A0(n2562), .A1(n2433), .Z(shiftedXdata[156]));
Q_MX02 U7086 ( .S(shiftCount[7]), .A0(n2561), .A1(n2432), .Z(shiftedXdata[155]));
Q_MX02 U7087 ( .S(shiftCount[7]), .A0(n2560), .A1(n2431), .Z(shiftedXdata[154]));
Q_MX02 U7088 ( .S(shiftCount[7]), .A0(n2559), .A1(n2430), .Z(shiftedXdata[153]));
Q_MX02 U7089 ( .S(shiftCount[7]), .A0(n2558), .A1(n2429), .Z(shiftedXdata[152]));
Q_MX02 U7090 ( .S(shiftCount[7]), .A0(n2557), .A1(n2428), .Z(shiftedXdata[151]));
Q_MX02 U7091 ( .S(shiftCount[7]), .A0(n2556), .A1(n2427), .Z(shiftedXdata[150]));
Q_MX02 U7092 ( .S(shiftCount[7]), .A0(n2555), .A1(n2426), .Z(shiftedXdata[149]));
Q_MX02 U7093 ( .S(shiftCount[7]), .A0(n2554), .A1(n2425), .Z(shiftedXdata[148]));
Q_MX02 U7094 ( .S(shiftCount[7]), .A0(n2553), .A1(n2424), .Z(shiftedXdata[147]));
Q_MX02 U7095 ( .S(shiftCount[7]), .A0(n2552), .A1(n2423), .Z(shiftedXdata[146]));
Q_MX02 U7096 ( .S(shiftCount[7]), .A0(n2551), .A1(n2422), .Z(shiftedXdata[145]));
Q_MX02 U7097 ( .S(shiftCount[7]), .A0(n2550), .A1(n2421), .Z(shiftedXdata[144]));
Q_MX02 U7098 ( .S(shiftCount[7]), .A0(n2549), .A1(n2420), .Z(shiftedXdata[143]));
Q_MX02 U7099 ( .S(shiftCount[7]), .A0(n2548), .A1(n2419), .Z(shiftedXdata[142]));
Q_MX02 U7100 ( .S(shiftCount[7]), .A0(n2547), .A1(n2418), .Z(shiftedXdata[141]));
Q_MX02 U7101 ( .S(shiftCount[7]), .A0(n2546), .A1(n2417), .Z(shiftedXdata[140]));
Q_MX02 U7102 ( .S(shiftCount[7]), .A0(n2545), .A1(n2416), .Z(shiftedXdata[139]));
Q_MX02 U7103 ( .S(shiftCount[7]), .A0(n2544), .A1(n2415), .Z(shiftedXdata[138]));
Q_MX02 U7104 ( .S(shiftCount[7]), .A0(n2543), .A1(n2414), .Z(shiftedXdata[137]));
Q_MX02 U7105 ( .S(shiftCount[7]), .A0(n2542), .A1(n2413), .Z(shiftedXdata[136]));
Q_MX02 U7106 ( .S(shiftCount[7]), .A0(n2541), .A1(n2412), .Z(shiftedXdata[135]));
Q_MX02 U7107 ( .S(shiftCount[7]), .A0(n2540), .A1(n2411), .Z(shiftedXdata[134]));
Q_MX02 U7108 ( .S(shiftCount[7]), .A0(n2539), .A1(n2410), .Z(shiftedXdata[133]));
Q_MX02 U7109 ( .S(shiftCount[7]), .A0(n2538), .A1(n2409), .Z(shiftedXdata[132]));
Q_MX02 U7110 ( .S(shiftCount[7]), .A0(n2537), .A1(n2408), .Z(shiftedXdata[131]));
Q_MX02 U7111 ( .S(shiftCount[7]), .A0(n2536), .A1(n2407), .Z(shiftedXdata[130]));
Q_MX02 U7112 ( .S(shiftCount[7]), .A0(n2535), .A1(n2406), .Z(shiftedXdata[129]));
Q_MX02 U7113 ( .S(shiftCount[7]), .A0(n2534), .A1(n2405), .Z(shiftedXdata[128]));
Q_INV U7114 ( .A(shiftCount[7]), .Z(n2404));
Q_AN02 U7115 ( .A0(n2404), .A1(n2533), .Z(shiftedXdata[127]));
Q_AN02 U7116 ( .A0(n2404), .A1(n2532), .Z(shiftedXdata[126]));
Q_AN02 U7117 ( .A0(n2404), .A1(n2531), .Z(shiftedXdata[125]));
Q_AN02 U7118 ( .A0(n2404), .A1(n2530), .Z(shiftedXdata[124]));
Q_AN02 U7119 ( .A0(n2404), .A1(n2529), .Z(shiftedXdata[123]));
Q_AN02 U7120 ( .A0(n2404), .A1(n2528), .Z(shiftedXdata[122]));
Q_AN02 U7121 ( .A0(n2404), .A1(n2527), .Z(shiftedXdata[121]));
Q_AN02 U7122 ( .A0(n2404), .A1(n2526), .Z(shiftedXdata[120]));
Q_AN02 U7123 ( .A0(n2404), .A1(n2525), .Z(shiftedXdata[119]));
Q_AN02 U7124 ( .A0(n2404), .A1(n2524), .Z(shiftedXdata[118]));
Q_AN02 U7125 ( .A0(n2404), .A1(n2523), .Z(shiftedXdata[117]));
Q_AN02 U7126 ( .A0(n2404), .A1(n2522), .Z(shiftedXdata[116]));
Q_AN02 U7127 ( .A0(n2404), .A1(n2521), .Z(shiftedXdata[115]));
Q_AN02 U7128 ( .A0(n2404), .A1(n2520), .Z(shiftedXdata[114]));
Q_AN02 U7129 ( .A0(n2404), .A1(n2519), .Z(shiftedXdata[113]));
Q_AN02 U7130 ( .A0(n2404), .A1(n2518), .Z(shiftedXdata[112]));
Q_AN02 U7131 ( .A0(n2404), .A1(n2517), .Z(shiftedXdata[111]));
Q_AN02 U7132 ( .A0(n2404), .A1(n2516), .Z(shiftedXdata[110]));
Q_AN02 U7133 ( .A0(n2404), .A1(n2515), .Z(shiftedXdata[109]));
Q_AN02 U7134 ( .A0(n2404), .A1(n2514), .Z(shiftedXdata[108]));
Q_AN02 U7135 ( .A0(n2404), .A1(n2513), .Z(shiftedXdata[107]));
Q_AN02 U7136 ( .A0(n2404), .A1(n2512), .Z(shiftedXdata[106]));
Q_AN02 U7137 ( .A0(n2404), .A1(n2511), .Z(shiftedXdata[105]));
Q_AN02 U7138 ( .A0(n2404), .A1(n2510), .Z(shiftedXdata[104]));
Q_AN02 U7139 ( .A0(n2404), .A1(n2509), .Z(shiftedXdata[103]));
Q_AN02 U7140 ( .A0(n2404), .A1(n2508), .Z(shiftedXdata[102]));
Q_AN02 U7141 ( .A0(n2404), .A1(n2507), .Z(shiftedXdata[101]));
Q_AN02 U7142 ( .A0(n2404), .A1(n2506), .Z(shiftedXdata[100]));
Q_AN02 U7143 ( .A0(n2404), .A1(n2505), .Z(shiftedXdata[99]));
Q_AN02 U7144 ( .A0(n2404), .A1(n2504), .Z(shiftedXdata[98]));
Q_AN02 U7145 ( .A0(n2404), .A1(n2503), .Z(shiftedXdata[97]));
Q_AN02 U7146 ( .A0(n2404), .A1(n2502), .Z(shiftedXdata[96]));
Q_AN02 U7147 ( .A0(n2404), .A1(n2501), .Z(shiftedXdata[95]));
Q_AN02 U7148 ( .A0(n2404), .A1(n2500), .Z(shiftedXdata[94]));
Q_AN02 U7149 ( .A0(n2404), .A1(n2499), .Z(shiftedXdata[93]));
Q_AN02 U7150 ( .A0(n2404), .A1(n2498), .Z(shiftedXdata[92]));
Q_AN02 U7151 ( .A0(n2404), .A1(n2497), .Z(shiftedXdata[91]));
Q_AN02 U7152 ( .A0(n2404), .A1(n2496), .Z(shiftedXdata[90]));
Q_AN02 U7153 ( .A0(n2404), .A1(n2495), .Z(shiftedXdata[89]));
Q_AN02 U7154 ( .A0(n2404), .A1(n2494), .Z(shiftedXdata[88]));
Q_AN02 U7155 ( .A0(n2404), .A1(n2493), .Z(shiftedXdata[87]));
Q_AN02 U7156 ( .A0(n2404), .A1(n2492), .Z(shiftedXdata[86]));
Q_AN02 U7157 ( .A0(n2404), .A1(n2491), .Z(shiftedXdata[85]));
Q_AN02 U7158 ( .A0(n2404), .A1(n2490), .Z(shiftedXdata[84]));
Q_AN02 U7159 ( .A0(n2404), .A1(n2489), .Z(shiftedXdata[83]));
Q_AN02 U7160 ( .A0(n2404), .A1(n2488), .Z(shiftedXdata[82]));
Q_AN02 U7161 ( .A0(n2404), .A1(n2487), .Z(shiftedXdata[81]));
Q_AN02 U7162 ( .A0(n2404), .A1(n2486), .Z(shiftedXdata[80]));
Q_AN02 U7163 ( .A0(n2404), .A1(n2485), .Z(shiftedXdata[79]));
Q_AN02 U7164 ( .A0(n2404), .A1(n2484), .Z(shiftedXdata[78]));
Q_AN02 U7165 ( .A0(n2404), .A1(n2483), .Z(shiftedXdata[77]));
Q_AN02 U7166 ( .A0(n2404), .A1(n2482), .Z(shiftedXdata[76]));
Q_AN02 U7167 ( .A0(n2404), .A1(n2481), .Z(shiftedXdata[75]));
Q_AN02 U7168 ( .A0(n2404), .A1(n2480), .Z(shiftedXdata[74]));
Q_AN02 U7169 ( .A0(n2404), .A1(n2479), .Z(shiftedXdata[73]));
Q_AN02 U7170 ( .A0(n2404), .A1(n2478), .Z(shiftedXdata[72]));
Q_AN02 U7171 ( .A0(n2404), .A1(n2477), .Z(shiftedXdata[71]));
Q_AN02 U7172 ( .A0(n2404), .A1(n2476), .Z(shiftedXdata[70]));
Q_AN02 U7173 ( .A0(n2404), .A1(n2475), .Z(shiftedXdata[69]));
Q_AN02 U7174 ( .A0(n2404), .A1(n2474), .Z(shiftedXdata[68]));
Q_AN02 U7175 ( .A0(n2404), .A1(n2473), .Z(shiftedXdata[67]));
Q_AN02 U7176 ( .A0(n2404), .A1(n2472), .Z(shiftedXdata[66]));
Q_AN02 U7177 ( .A0(n2404), .A1(n2471), .Z(shiftedXdata[65]));
Q_AN02 U7178 ( .A0(n2404), .A1(n2470), .Z(shiftedXdata[64]));
Q_AN02 U7179 ( .A0(n2404), .A1(n2468), .Z(shiftedXdata[63]));
Q_AN02 U7180 ( .A0(n2404), .A1(n2467), .Z(shiftedXdata[62]));
Q_AN02 U7181 ( .A0(n2404), .A1(n2466), .Z(shiftedXdata[61]));
Q_AN02 U7182 ( .A0(n2404), .A1(n2465), .Z(shiftedXdata[60]));
Q_AN02 U7183 ( .A0(n2404), .A1(n2464), .Z(shiftedXdata[59]));
Q_AN02 U7184 ( .A0(n2404), .A1(n2463), .Z(shiftedXdata[58]));
Q_AN02 U7185 ( .A0(n2404), .A1(n2462), .Z(shiftedXdata[57]));
Q_AN02 U7186 ( .A0(n2404), .A1(n2461), .Z(shiftedXdata[56]));
Q_AN02 U7187 ( .A0(n2404), .A1(n2460), .Z(shiftedXdata[55]));
Q_AN02 U7188 ( .A0(n2404), .A1(n2459), .Z(shiftedXdata[54]));
Q_AN02 U7189 ( .A0(n2404), .A1(n2458), .Z(shiftedXdata[53]));
Q_AN02 U7190 ( .A0(n2404), .A1(n2457), .Z(shiftedXdata[52]));
Q_AN02 U7191 ( .A0(n2404), .A1(n2456), .Z(shiftedXdata[51]));
Q_AN02 U7192 ( .A0(n2404), .A1(n2455), .Z(shiftedXdata[50]));
Q_AN02 U7193 ( .A0(n2404), .A1(n2454), .Z(shiftedXdata[49]));
Q_AN02 U7194 ( .A0(n2404), .A1(n2453), .Z(shiftedXdata[48]));
Q_AN02 U7195 ( .A0(n2404), .A1(n2452), .Z(shiftedXdata[47]));
Q_AN02 U7196 ( .A0(n2404), .A1(n2451), .Z(shiftedXdata[46]));
Q_AN02 U7197 ( .A0(n2404), .A1(n2450), .Z(shiftedXdata[45]));
Q_AN02 U7198 ( .A0(n2404), .A1(n2449), .Z(shiftedXdata[44]));
Q_AN02 U7199 ( .A0(n2404), .A1(n2448), .Z(shiftedXdata[43]));
Q_AN02 U7200 ( .A0(n2404), .A1(n2447), .Z(shiftedXdata[42]));
Q_AN02 U7201 ( .A0(n2404), .A1(n2446), .Z(shiftedXdata[41]));
Q_AN02 U7202 ( .A0(n2404), .A1(n2445), .Z(shiftedXdata[40]));
Q_AN02 U7203 ( .A0(n2404), .A1(n2444), .Z(shiftedXdata[39]));
Q_AN02 U7204 ( .A0(n2404), .A1(n2443), .Z(shiftedXdata[38]));
Q_AN02 U7205 ( .A0(n2404), .A1(n2442), .Z(shiftedXdata[37]));
Q_AN02 U7206 ( .A0(n2404), .A1(n2441), .Z(shiftedXdata[36]));
Q_AN02 U7207 ( .A0(n2404), .A1(n2440), .Z(shiftedXdata[35]));
Q_AN02 U7208 ( .A0(n2404), .A1(n2439), .Z(shiftedXdata[34]));
Q_AN02 U7209 ( .A0(n2404), .A1(n2438), .Z(shiftedXdata[33]));
Q_AN02 U7210 ( .A0(n2404), .A1(n2437), .Z(shiftedXdata[32]));
Q_AN02 U7211 ( .A0(n2404), .A1(n2436), .Z(shiftedXdata[31]));
Q_AN02 U7212 ( .A0(n2404), .A1(n2435), .Z(shiftedXdata[30]));
Q_AN02 U7213 ( .A0(n2404), .A1(n2434), .Z(shiftedXdata[29]));
Q_AN02 U7214 ( .A0(n2404), .A1(n2433), .Z(shiftedXdata[28]));
Q_AN02 U7215 ( .A0(n2404), .A1(n2432), .Z(shiftedXdata[27]));
Q_AN02 U7216 ( .A0(n2404), .A1(n2431), .Z(shiftedXdata[26]));
Q_AN02 U7217 ( .A0(n2404), .A1(n2430), .Z(shiftedXdata[25]));
Q_AN02 U7218 ( .A0(n2404), .A1(n2429), .Z(shiftedXdata[24]));
Q_AN02 U7219 ( .A0(n2404), .A1(n2428), .Z(shiftedXdata[23]));
Q_AN02 U7220 ( .A0(n2404), .A1(n2427), .Z(shiftedXdata[22]));
Q_AN02 U7221 ( .A0(n2404), .A1(n2426), .Z(shiftedXdata[21]));
Q_AN02 U7222 ( .A0(n2404), .A1(n2425), .Z(shiftedXdata[20]));
Q_AN02 U7223 ( .A0(n2404), .A1(n2424), .Z(shiftedXdata[19]));
Q_AN02 U7224 ( .A0(n2404), .A1(n2423), .Z(shiftedXdata[18]));
Q_AN02 U7225 ( .A0(n2404), .A1(n2422), .Z(shiftedXdata[17]));
Q_AN02 U7226 ( .A0(n2404), .A1(n2421), .Z(shiftedXdata[16]));
Q_AN02 U7227 ( .A0(n2404), .A1(n2420), .Z(shiftedXdata[15]));
Q_AN02 U7228 ( .A0(n2404), .A1(n2419), .Z(shiftedXdata[14]));
Q_AN02 U7229 ( .A0(n2404), .A1(n2418), .Z(shiftedXdata[13]));
Q_AN02 U7230 ( .A0(n2404), .A1(n2417), .Z(shiftedXdata[12]));
Q_AN02 U7231 ( .A0(n2404), .A1(n2416), .Z(shiftedXdata[11]));
Q_AN02 U7232 ( .A0(n2404), .A1(n2415), .Z(shiftedXdata[10]));
Q_AN02 U7233 ( .A0(n2404), .A1(n2414), .Z(shiftedXdata[9]));
Q_AN02 U7234 ( .A0(n2404), .A1(n2413), .Z(shiftedXdata[8]));
Q_AN02 U7235 ( .A0(n2404), .A1(n2412), .Z(shiftedXdata[7]));
Q_AN02 U7236 ( .A0(n2404), .A1(n2411), .Z(shiftedXdata[6]));
Q_AN02 U7237 ( .A0(n2404), .A1(n2410), .Z(shiftedXdata[5]));
Q_AN02 U7238 ( .A0(n2404), .A1(n2409), .Z(shiftedXdata[4]));
Q_AN02 U7239 ( .A0(n2404), .A1(n2408), .Z(shiftedXdata[3]));
Q_AN02 U7240 ( .A0(n2404), .A1(n2407), .Z(shiftedXdata[2]));
Q_AN02 U7241 ( .A0(n2404), .A1(n2406), .Z(shiftedXdata[1]));
Q_AN02 U7242 ( .A0(n2404), .A1(n2405), .Z(shiftedXdata[0]));
Q_AO21 U7243 ( .A0(oFill[3]), .A1(oFill[4]), .B0(xc_top.GFReset), .Z(n2141));
Q_INV U7244 ( .A(oFill[3]), .Z(n2403));
Q_AN02 U7245 ( .A0(n2403), .A1(oFill[4]), .Z(n2402));
Q_OR02 U7246 ( .A0(n2401), .A1(shiftedXdata[0]), .Z(n2142));
Q_OR02 U7247 ( .A0(n2400), .A1(shiftedXdata[1]), .Z(n2139));
Q_OR02 U7248 ( .A0(n2399), .A1(shiftedXdata[2]), .Z(n2137));
Q_OR02 U7249 ( .A0(n2398), .A1(shiftedXdata[3]), .Z(n2135));
Q_OR02 U7250 ( .A0(n2397), .A1(shiftedXdata[4]), .Z(n2133));
Q_OR02 U7251 ( .A0(n2396), .A1(shiftedXdata[5]), .Z(n2131));
Q_OR02 U7252 ( .A0(n2395), .A1(shiftedXdata[6]), .Z(n2129));
Q_OR02 U7253 ( .A0(n2394), .A1(shiftedXdata[7]), .Z(n2127));
Q_OR02 U7254 ( .A0(n2393), .A1(shiftedXdata[8]), .Z(n2125));
Q_OR02 U7255 ( .A0(n2392), .A1(shiftedXdata[9]), .Z(n2123));
Q_OR02 U7256 ( .A0(n2391), .A1(shiftedXdata[10]), .Z(n2121));
Q_OR02 U7257 ( .A0(n2390), .A1(shiftedXdata[11]), .Z(n2119));
Q_OR02 U7258 ( .A0(n2389), .A1(shiftedXdata[12]), .Z(n2117));
Q_OR02 U7259 ( .A0(n2388), .A1(shiftedXdata[13]), .Z(n2115));
Q_OR02 U7260 ( .A0(n2387), .A1(shiftedXdata[14]), .Z(n2113));
Q_OR02 U7261 ( .A0(n2386), .A1(shiftedXdata[15]), .Z(n2111));
Q_OR02 U7262 ( .A0(n2385), .A1(shiftedXdata[16]), .Z(n2109));
Q_OR02 U7263 ( .A0(n2384), .A1(shiftedXdata[17]), .Z(n2107));
Q_OR02 U7264 ( .A0(n2383), .A1(shiftedXdata[18]), .Z(n2105));
Q_OR02 U7265 ( .A0(n2382), .A1(shiftedXdata[19]), .Z(n2103));
Q_OR02 U7266 ( .A0(n2381), .A1(shiftedXdata[20]), .Z(n2101));
Q_OR02 U7267 ( .A0(n2380), .A1(shiftedXdata[21]), .Z(n2099));
Q_OR02 U7268 ( .A0(n2379), .A1(shiftedXdata[22]), .Z(n2097));
Q_OR02 U7269 ( .A0(n2378), .A1(shiftedXdata[23]), .Z(n2095));
Q_OR02 U7270 ( .A0(n2377), .A1(shiftedXdata[24]), .Z(n2093));
Q_OR02 U7271 ( .A0(n2376), .A1(shiftedXdata[25]), .Z(n2091));
Q_OR02 U7272 ( .A0(n2375), .A1(shiftedXdata[26]), .Z(n2089));
Q_OR02 U7273 ( .A0(n2374), .A1(shiftedXdata[27]), .Z(n2087));
Q_OR02 U7274 ( .A0(n2373), .A1(shiftedXdata[28]), .Z(n2085));
Q_OR02 U7275 ( .A0(n2372), .A1(shiftedXdata[29]), .Z(n2083));
Q_OR02 U7276 ( .A0(n2371), .A1(shiftedXdata[30]), .Z(n2081));
Q_OR02 U7277 ( .A0(n2370), .A1(shiftedXdata[31]), .Z(n2079));
Q_OR02 U7278 ( .A0(n2369), .A1(shiftedXdata[32]), .Z(n2077));
Q_OR02 U7279 ( .A0(n2368), .A1(shiftedXdata[33]), .Z(n2075));
Q_OR02 U7280 ( .A0(n2367), .A1(shiftedXdata[34]), .Z(n2073));
Q_OR02 U7281 ( .A0(n2366), .A1(shiftedXdata[35]), .Z(n2071));
Q_OR02 U7282 ( .A0(n2365), .A1(shiftedXdata[36]), .Z(n2069));
Q_OR02 U7283 ( .A0(n2364), .A1(shiftedXdata[37]), .Z(n2067));
Q_OR02 U7284 ( .A0(n2363), .A1(shiftedXdata[38]), .Z(n2065));
Q_OR02 U7285 ( .A0(n2362), .A1(shiftedXdata[39]), .Z(n2063));
Q_OR02 U7286 ( .A0(n2361), .A1(shiftedXdata[40]), .Z(n2061));
Q_OR02 U7287 ( .A0(n2360), .A1(shiftedXdata[41]), .Z(n2059));
Q_OR02 U7288 ( .A0(n2359), .A1(shiftedXdata[42]), .Z(n2057));
Q_OR02 U7289 ( .A0(n2358), .A1(shiftedXdata[43]), .Z(n2055));
Q_OR02 U7290 ( .A0(n2357), .A1(shiftedXdata[44]), .Z(n2053));
Q_OR02 U7291 ( .A0(n2356), .A1(shiftedXdata[45]), .Z(n2051));
Q_OR02 U7292 ( .A0(n2355), .A1(shiftedXdata[46]), .Z(n2049));
Q_OR02 U7293 ( .A0(n2354), .A1(shiftedXdata[47]), .Z(n2047));
Q_OR02 U7294 ( .A0(n2353), .A1(shiftedXdata[48]), .Z(n2045));
Q_OR02 U7295 ( .A0(n2352), .A1(shiftedXdata[49]), .Z(n2043));
Q_OR02 U7296 ( .A0(n2351), .A1(shiftedXdata[50]), .Z(n2041));
Q_OR02 U7297 ( .A0(n2350), .A1(shiftedXdata[51]), .Z(n2039));
Q_OR02 U7298 ( .A0(n2349), .A1(shiftedXdata[52]), .Z(n2037));
Q_OR02 U7299 ( .A0(n2348), .A1(shiftedXdata[53]), .Z(n2035));
Q_OR02 U7300 ( .A0(n2347), .A1(shiftedXdata[54]), .Z(n2033));
Q_OR02 U7301 ( .A0(n2346), .A1(shiftedXdata[55]), .Z(n2031));
Q_OR02 U7302 ( .A0(n2345), .A1(shiftedXdata[56]), .Z(n2029));
Q_OR02 U7303 ( .A0(n2344), .A1(shiftedXdata[57]), .Z(n2027));
Q_OR02 U7304 ( .A0(n2343), .A1(shiftedXdata[58]), .Z(n2025));
Q_OR02 U7305 ( .A0(n2342), .A1(shiftedXdata[59]), .Z(n2023));
Q_OR02 U7306 ( .A0(n2341), .A1(shiftedXdata[60]), .Z(n2021));
Q_OR02 U7307 ( .A0(n2340), .A1(shiftedXdata[61]), .Z(n2019));
Q_OR02 U7308 ( .A0(n2339), .A1(shiftedXdata[62]), .Z(n2017));
Q_OR02 U7309 ( .A0(n2338), .A1(shiftedXdata[63]), .Z(n2015));
Q_OR02 U7310 ( .A0(n2337), .A1(shiftedXdata[64]), .Z(n2013));
Q_OR02 U7311 ( .A0(n2336), .A1(shiftedXdata[65]), .Z(n2011));
Q_OR02 U7312 ( .A0(n2335), .A1(shiftedXdata[66]), .Z(n2009));
Q_OR02 U7313 ( .A0(n2334), .A1(shiftedXdata[67]), .Z(n2007));
Q_OR02 U7314 ( .A0(n2333), .A1(shiftedXdata[68]), .Z(n2005));
Q_OR02 U7315 ( .A0(n2332), .A1(shiftedXdata[69]), .Z(n2003));
Q_OR02 U7316 ( .A0(n2331), .A1(shiftedXdata[70]), .Z(n2001));
Q_OR02 U7317 ( .A0(n2330), .A1(shiftedXdata[71]), .Z(n1999));
Q_OR02 U7318 ( .A0(n2329), .A1(shiftedXdata[72]), .Z(n1997));
Q_OR02 U7319 ( .A0(n2328), .A1(shiftedXdata[73]), .Z(n1995));
Q_OR02 U7320 ( .A0(n2327), .A1(shiftedXdata[74]), .Z(n1993));
Q_OR02 U7321 ( .A0(n2326), .A1(shiftedXdata[75]), .Z(n1991));
Q_OR02 U7322 ( .A0(n2325), .A1(shiftedXdata[76]), .Z(n1989));
Q_OR02 U7323 ( .A0(n2324), .A1(shiftedXdata[77]), .Z(n1987));
Q_OR02 U7324 ( .A0(n2323), .A1(shiftedXdata[78]), .Z(n1985));
Q_OR02 U7325 ( .A0(n2322), .A1(shiftedXdata[79]), .Z(n1983));
Q_OR02 U7326 ( .A0(n2321), .A1(shiftedXdata[80]), .Z(n1981));
Q_OR02 U7327 ( .A0(n2320), .A1(shiftedXdata[81]), .Z(n1979));
Q_OR02 U7328 ( .A0(n2319), .A1(shiftedXdata[82]), .Z(n1977));
Q_OR02 U7329 ( .A0(n2318), .A1(shiftedXdata[83]), .Z(n1975));
Q_OR02 U7330 ( .A0(n2317), .A1(shiftedXdata[84]), .Z(n1973));
Q_OR02 U7331 ( .A0(n2316), .A1(shiftedXdata[85]), .Z(n1971));
Q_OR02 U7332 ( .A0(n2315), .A1(shiftedXdata[86]), .Z(n1969));
Q_OR02 U7333 ( .A0(n2314), .A1(shiftedXdata[87]), .Z(n1967));
Q_OR02 U7334 ( .A0(n2313), .A1(shiftedXdata[88]), .Z(n1965));
Q_OR02 U7335 ( .A0(n2312), .A1(shiftedXdata[89]), .Z(n1963));
Q_OR02 U7336 ( .A0(n2311), .A1(shiftedXdata[90]), .Z(n1961));
Q_OR02 U7337 ( .A0(n2310), .A1(shiftedXdata[91]), .Z(n1959));
Q_OR02 U7338 ( .A0(n2309), .A1(shiftedXdata[92]), .Z(n1957));
Q_OR02 U7339 ( .A0(n2308), .A1(shiftedXdata[93]), .Z(n1955));
Q_OR02 U7340 ( .A0(n2307), .A1(shiftedXdata[94]), .Z(n1953));
Q_OR02 U7341 ( .A0(n2306), .A1(shiftedXdata[95]), .Z(n1951));
Q_OR02 U7342 ( .A0(n2305), .A1(shiftedXdata[96]), .Z(n1949));
Q_OR02 U7343 ( .A0(n2304), .A1(shiftedXdata[97]), .Z(n1947));
Q_OR02 U7344 ( .A0(n2303), .A1(shiftedXdata[98]), .Z(n1945));
Q_OR02 U7345 ( .A0(n2302), .A1(shiftedXdata[99]), .Z(n1943));
Q_OR02 U7346 ( .A0(n2301), .A1(shiftedXdata[100]), .Z(n1941));
Q_OR02 U7347 ( .A0(n2300), .A1(shiftedXdata[101]), .Z(n1939));
Q_OR02 U7348 ( .A0(n2299), .A1(shiftedXdata[102]), .Z(n1937));
Q_OR02 U7349 ( .A0(n2298), .A1(shiftedXdata[103]), .Z(n1935));
Q_OR02 U7350 ( .A0(n2297), .A1(shiftedXdata[104]), .Z(n1933));
Q_OR02 U7351 ( .A0(n2296), .A1(shiftedXdata[105]), .Z(n1931));
Q_OR02 U7352 ( .A0(n2295), .A1(shiftedXdata[106]), .Z(n1929));
Q_OR02 U7353 ( .A0(n2294), .A1(shiftedXdata[107]), .Z(n1927));
Q_OR02 U7354 ( .A0(n2293), .A1(shiftedXdata[108]), .Z(n1925));
Q_OR02 U7355 ( .A0(n2292), .A1(shiftedXdata[109]), .Z(n1923));
Q_OR02 U7356 ( .A0(n2291), .A1(shiftedXdata[110]), .Z(n1921));
Q_OR02 U7357 ( .A0(n2290), .A1(shiftedXdata[111]), .Z(n1919));
Q_OR02 U7358 ( .A0(n2289), .A1(shiftedXdata[112]), .Z(n1917));
Q_OR02 U7359 ( .A0(n2288), .A1(shiftedXdata[113]), .Z(n1915));
Q_OR02 U7360 ( .A0(n2287), .A1(shiftedXdata[114]), .Z(n1913));
Q_OR02 U7361 ( .A0(n2286), .A1(shiftedXdata[115]), .Z(n1911));
Q_OR02 U7362 ( .A0(n2285), .A1(shiftedXdata[116]), .Z(n1909));
Q_OR02 U7363 ( .A0(n2284), .A1(shiftedXdata[117]), .Z(n1907));
Q_OR02 U7364 ( .A0(n2283), .A1(shiftedXdata[118]), .Z(n1905));
Q_OR02 U7365 ( .A0(n2282), .A1(shiftedXdata[119]), .Z(n1903));
Q_OR02 U7366 ( .A0(n2281), .A1(shiftedXdata[120]), .Z(n1901));
Q_OR02 U7367 ( .A0(n2280), .A1(shiftedXdata[121]), .Z(n1899));
Q_OR02 U7368 ( .A0(n2279), .A1(shiftedXdata[122]), .Z(n1897));
Q_OR02 U7369 ( .A0(n2278), .A1(shiftedXdata[123]), .Z(n1895));
Q_OR02 U7370 ( .A0(n2277), .A1(shiftedXdata[124]), .Z(n1893));
Q_OR02 U7371 ( .A0(n2276), .A1(shiftedXdata[125]), .Z(n1891));
Q_OR02 U7372 ( .A0(n2275), .A1(shiftedXdata[126]), .Z(n1889));
Q_OR02 U7373 ( .A0(n2274), .A1(shiftedXdata[127]), .Z(n1887));
Q_OR02 U7374 ( .A0(n2273), .A1(shiftedXdata[128]), .Z(n1885));
Q_OR02 U7375 ( .A0(n2272), .A1(shiftedXdata[129]), .Z(n1883));
Q_OR02 U7376 ( .A0(n2271), .A1(shiftedXdata[130]), .Z(n1881));
Q_OR02 U7377 ( .A0(n2270), .A1(shiftedXdata[131]), .Z(n1879));
Q_OR02 U7378 ( .A0(n2269), .A1(shiftedXdata[132]), .Z(n1877));
Q_OR02 U7379 ( .A0(n2268), .A1(shiftedXdata[133]), .Z(n1875));
Q_OR02 U7380 ( .A0(n2267), .A1(shiftedXdata[134]), .Z(n1873));
Q_OR02 U7381 ( .A0(n2266), .A1(shiftedXdata[135]), .Z(n1871));
Q_OR02 U7382 ( .A0(n2265), .A1(shiftedXdata[136]), .Z(n1869));
Q_OR02 U7383 ( .A0(n2264), .A1(shiftedXdata[137]), .Z(n1867));
Q_OR02 U7384 ( .A0(n2263), .A1(shiftedXdata[138]), .Z(n1865));
Q_OR02 U7385 ( .A0(n2262), .A1(shiftedXdata[139]), .Z(n1863));
Q_OR02 U7386 ( .A0(n2261), .A1(shiftedXdata[140]), .Z(n1861));
Q_OR02 U7387 ( .A0(n2260), .A1(shiftedXdata[141]), .Z(n1859));
Q_OR02 U7388 ( .A0(n2259), .A1(shiftedXdata[142]), .Z(n1857));
Q_OR02 U7389 ( .A0(n2258), .A1(shiftedXdata[143]), .Z(n1855));
Q_OR02 U7390 ( .A0(n2257), .A1(shiftedXdata[144]), .Z(n1853));
Q_OR02 U7391 ( .A0(n2256), .A1(shiftedXdata[145]), .Z(n1851));
Q_OR02 U7392 ( .A0(n2255), .A1(shiftedXdata[146]), .Z(n1849));
Q_OR02 U7393 ( .A0(n2254), .A1(shiftedXdata[147]), .Z(n1847));
Q_OR02 U7394 ( .A0(n2253), .A1(shiftedXdata[148]), .Z(n1845));
Q_OR02 U7395 ( .A0(n2252), .A1(shiftedXdata[149]), .Z(n1843));
Q_OR02 U7396 ( .A0(n2251), .A1(shiftedXdata[150]), .Z(n1841));
Q_OR02 U7397 ( .A0(n2250), .A1(shiftedXdata[151]), .Z(n1839));
Q_OR02 U7398 ( .A0(n2249), .A1(shiftedXdata[152]), .Z(n1837));
Q_OR02 U7399 ( .A0(n2248), .A1(shiftedXdata[153]), .Z(n1835));
Q_OR02 U7400 ( .A0(n2247), .A1(shiftedXdata[154]), .Z(n1833));
Q_OR02 U7401 ( .A0(n2246), .A1(shiftedXdata[155]), .Z(n1831));
Q_OR02 U7402 ( .A0(n2245), .A1(shiftedXdata[156]), .Z(n1829));
Q_OR02 U7403 ( .A0(n2244), .A1(shiftedXdata[157]), .Z(n1827));
Q_OR02 U7404 ( .A0(n2243), .A1(shiftedXdata[158]), .Z(n1825));
Q_OR02 U7405 ( .A0(n2242), .A1(shiftedXdata[159]), .Z(n1823));
Q_OR02 U7406 ( .A0(n2241), .A1(shiftedXdata[160]), .Z(n1821));
Q_OR02 U7407 ( .A0(n2240), .A1(shiftedXdata[161]), .Z(n1819));
Q_OR02 U7408 ( .A0(n2239), .A1(shiftedXdata[162]), .Z(n1817));
Q_OR02 U7409 ( .A0(n2238), .A1(shiftedXdata[163]), .Z(n1815));
Q_OR02 U7410 ( .A0(n2237), .A1(shiftedXdata[164]), .Z(n1813));
Q_OR02 U7411 ( .A0(n2236), .A1(shiftedXdata[165]), .Z(n1811));
Q_OR02 U7412 ( .A0(n2235), .A1(shiftedXdata[166]), .Z(n1809));
Q_OR02 U7413 ( .A0(n2234), .A1(shiftedXdata[167]), .Z(n1807));
Q_OR02 U7414 ( .A0(n2233), .A1(shiftedXdata[168]), .Z(n1805));
Q_OR02 U7415 ( .A0(n2232), .A1(shiftedXdata[169]), .Z(n1803));
Q_OR02 U7416 ( .A0(n2231), .A1(shiftedXdata[170]), .Z(n1801));
Q_OR02 U7417 ( .A0(n2230), .A1(shiftedXdata[171]), .Z(n1799));
Q_OR02 U7418 ( .A0(n2229), .A1(shiftedXdata[172]), .Z(n1797));
Q_OR02 U7419 ( .A0(n2228), .A1(shiftedXdata[173]), .Z(n1795));
Q_OR02 U7420 ( .A0(n2227), .A1(shiftedXdata[174]), .Z(n1793));
Q_OR02 U7421 ( .A0(n2226), .A1(shiftedXdata[175]), .Z(n1791));
Q_OR02 U7422 ( .A0(n2225), .A1(shiftedXdata[176]), .Z(n1789));
Q_OR02 U7423 ( .A0(n2224), .A1(shiftedXdata[177]), .Z(n1787));
Q_OR02 U7424 ( .A0(n2223), .A1(shiftedXdata[178]), .Z(n1785));
Q_OR02 U7425 ( .A0(n2222), .A1(shiftedXdata[179]), .Z(n1783));
Q_OR02 U7426 ( .A0(n2221), .A1(shiftedXdata[180]), .Z(n1781));
Q_OR02 U7427 ( .A0(n2220), .A1(shiftedXdata[181]), .Z(n1779));
Q_OR02 U7428 ( .A0(n2219), .A1(shiftedXdata[182]), .Z(n1777));
Q_OR02 U7429 ( .A0(n2218), .A1(shiftedXdata[183]), .Z(n1775));
Q_OR02 U7430 ( .A0(n2217), .A1(shiftedXdata[184]), .Z(n1773));
Q_OR02 U7431 ( .A0(n2216), .A1(shiftedXdata[185]), .Z(n1771));
Q_OR02 U7432 ( .A0(n2215), .A1(shiftedXdata[186]), .Z(n1769));
Q_OR02 U7433 ( .A0(n2214), .A1(shiftedXdata[187]), .Z(n1767));
Q_OR02 U7434 ( .A0(n2213), .A1(shiftedXdata[188]), .Z(n1765));
Q_OR02 U7435 ( .A0(n2212), .A1(shiftedXdata[189]), .Z(n1763));
Q_OR02 U7436 ( .A0(n2211), .A1(shiftedXdata[190]), .Z(n1761));
Q_OR02 U7437 ( .A0(n2210), .A1(shiftedXdata[191]), .Z(n1759));
Q_OR02 U7438 ( .A0(n2209), .A1(shiftedXdata[192]), .Z(n1757));
Q_OR02 U7439 ( .A0(n2208), .A1(shiftedXdata[193]), .Z(n1755));
Q_OR02 U7440 ( .A0(n2207), .A1(shiftedXdata[194]), .Z(n1753));
Q_OR02 U7441 ( .A0(n2206), .A1(shiftedXdata[195]), .Z(n1751));
Q_OR02 U7442 ( .A0(n2205), .A1(shiftedXdata[196]), .Z(n1749));
Q_OR02 U7443 ( .A0(n2204), .A1(shiftedXdata[197]), .Z(n1747));
Q_OR02 U7444 ( .A0(n2203), .A1(shiftedXdata[198]), .Z(n1745));
Q_OR02 U7445 ( .A0(n2202), .A1(shiftedXdata[199]), .Z(n1743));
Q_OR02 U7446 ( .A0(n2201), .A1(shiftedXdata[200]), .Z(n1741));
Q_OR02 U7447 ( .A0(n2200), .A1(shiftedXdata[201]), .Z(n1739));
Q_OR02 U7448 ( .A0(n2199), .A1(shiftedXdata[202]), .Z(n1737));
Q_OR02 U7449 ( .A0(n2198), .A1(shiftedXdata[203]), .Z(n1735));
Q_OR02 U7450 ( .A0(n2197), .A1(shiftedXdata[204]), .Z(n1733));
Q_OR02 U7451 ( .A0(n2196), .A1(shiftedXdata[205]), .Z(n1731));
Q_OR02 U7452 ( .A0(n2195), .A1(shiftedXdata[206]), .Z(n1729));
Q_OR02 U7453 ( .A0(n2194), .A1(shiftedXdata[207]), .Z(n1727));
Q_OR02 U7454 ( .A0(n2193), .A1(shiftedXdata[208]), .Z(n1725));
Q_OR02 U7455 ( .A0(n2192), .A1(shiftedXdata[209]), .Z(n1723));
Q_OR02 U7456 ( .A0(n2191), .A1(shiftedXdata[210]), .Z(n1721));
Q_OR02 U7457 ( .A0(n2190), .A1(shiftedXdata[211]), .Z(n1719));
Q_OR02 U7458 ( .A0(n2189), .A1(shiftedXdata[212]), .Z(n1717));
Q_OR02 U7459 ( .A0(n2188), .A1(shiftedXdata[213]), .Z(n1715));
Q_OR02 U7460 ( .A0(n2187), .A1(shiftedXdata[214]), .Z(n1713));
Q_OR02 U7461 ( .A0(n2186), .A1(shiftedXdata[215]), .Z(n1711));
Q_OR02 U7462 ( .A0(n2185), .A1(shiftedXdata[216]), .Z(n1709));
Q_OR02 U7463 ( .A0(n2184), .A1(shiftedXdata[217]), .Z(n1707));
Q_OR02 U7464 ( .A0(n2183), .A1(shiftedXdata[218]), .Z(n1705));
Q_OR02 U7465 ( .A0(n2182), .A1(shiftedXdata[219]), .Z(n1703));
Q_OR02 U7466 ( .A0(n2181), .A1(shiftedXdata[220]), .Z(n1701));
Q_OR02 U7467 ( .A0(n2180), .A1(shiftedXdata[221]), .Z(n1699));
Q_OR02 U7468 ( .A0(n2179), .A1(shiftedXdata[222]), .Z(n1697));
Q_OR02 U7469 ( .A0(n2178), .A1(shiftedXdata[223]), .Z(n1695));
Q_OR02 U7470 ( .A0(n2177), .A1(shiftedXdata[224]), .Z(n1693));
Q_OR02 U7471 ( .A0(n2176), .A1(shiftedXdata[225]), .Z(n1691));
Q_OR02 U7472 ( .A0(n2175), .A1(shiftedXdata[226]), .Z(n1689));
Q_OR02 U7473 ( .A0(n2174), .A1(shiftedXdata[227]), .Z(n1687));
Q_OR02 U7474 ( .A0(n2173), .A1(shiftedXdata[228]), .Z(n1685));
Q_OR02 U7475 ( .A0(n2172), .A1(shiftedXdata[229]), .Z(n1683));
Q_OR02 U7476 ( .A0(n2171), .A1(shiftedXdata[230]), .Z(n1681));
Q_OR02 U7477 ( .A0(n2170), .A1(shiftedXdata[231]), .Z(n1679));
Q_OR02 U7478 ( .A0(n2169), .A1(shiftedXdata[232]), .Z(n1677));
Q_OR02 U7479 ( .A0(n2168), .A1(shiftedXdata[233]), .Z(n1675));
Q_OR02 U7480 ( .A0(n2167), .A1(shiftedXdata[234]), .Z(n1673));
Q_OR02 U7481 ( .A0(n2166), .A1(shiftedXdata[235]), .Z(n1671));
Q_OR02 U7482 ( .A0(n2165), .A1(shiftedXdata[236]), .Z(n1669));
Q_OR02 U7483 ( .A0(n2164), .A1(shiftedXdata[237]), .Z(n1667));
Q_OR02 U7484 ( .A0(n2163), .A1(shiftedXdata[238]), .Z(n1665));
Q_OR02 U7485 ( .A0(n2162), .A1(shiftedXdata[239]), .Z(n1663));
Q_OR02 U7486 ( .A0(n2161), .A1(shiftedXdata[240]), .Z(n1661));
Q_OR02 U7487 ( .A0(n2160), .A1(shiftedXdata[241]), .Z(n1659));
Q_OR02 U7488 ( .A0(n2159), .A1(shiftedXdata[242]), .Z(n1657));
Q_OR02 U7489 ( .A0(n2158), .A1(shiftedXdata[243]), .Z(n1655));
Q_OR02 U7490 ( .A0(n2157), .A1(shiftedXdata[244]), .Z(n1653));
Q_OR02 U7491 ( .A0(n2156), .A1(shiftedXdata[245]), .Z(n1651));
Q_OR02 U7492 ( .A0(n2155), .A1(shiftedXdata[246]), .Z(n1649));
Q_OR02 U7493 ( .A0(n2154), .A1(shiftedXdata[247]), .Z(n1647));
Q_OR02 U7494 ( .A0(n2153), .A1(shiftedXdata[248]), .Z(n1645));
Q_OR02 U7495 ( .A0(n2152), .A1(shiftedXdata[249]), .Z(n1643));
Q_OR02 U7496 ( .A0(n2151), .A1(shiftedXdata[250]), .Z(n1641));
Q_OR02 U7497 ( .A0(n2150), .A1(shiftedXdata[251]), .Z(n1639));
Q_OR02 U7498 ( .A0(n2149), .A1(shiftedXdata[252]), .Z(n1637));
Q_OR02 U7499 ( .A0(n2148), .A1(shiftedXdata[253]), .Z(n1635));
Q_OR02 U7500 ( .A0(n2147), .A1(shiftedXdata[254]), .Z(n1633));
Q_OR02 U7501 ( .A0(n2146), .A1(shiftedXdata[255]), .Z(n1631));
Q_INV U7502 ( .A(oFill[4]), .Z(n2145));
Q_AN02 U7503 ( .A0(oFill[3]), .A1(n2145), .Z(n2144));
Q_AN02 U7504 ( .A0(n6720), .A1(shiftedXdata[0]), .Z(n2143));
Q_MX03 U7505 ( .S0(n2144), .S1(n2402), .A0(ofifoData[0]), .A1(ofifoData[256]), .A2(ofifoData[512]), .Z(n2401));
Q_MX02 U7506 ( .S(n2141), .A0(n2142), .A1(n2143), .Z(ofifoDataN[0]));
Q_AN02 U7507 ( .A0(n6720), .A1(shiftedXdata[1]), .Z(n2140));
Q_MX03 U7508 ( .S0(n2144), .S1(n2402), .A0(ofifoData[1]), .A1(ofifoData[257]), .A2(ofifoData[513]), .Z(n2400));
Q_MX02 U7509 ( .S(n2141), .A0(n2139), .A1(n2140), .Z(ofifoDataN[1]));
Q_AN02 U7510 ( .A0(n6720), .A1(shiftedXdata[2]), .Z(n2138));
Q_MX03 U7511 ( .S0(n2144), .S1(n2402), .A0(ofifoData[2]), .A1(ofifoData[258]), .A2(ofifoData[514]), .Z(n2399));
Q_MX02 U7512 ( .S(n2141), .A0(n2137), .A1(n2138), .Z(ofifoDataN[2]));
Q_AN02 U7513 ( .A0(n6720), .A1(shiftedXdata[3]), .Z(n2136));
Q_MX03 U7514 ( .S0(n2144), .S1(n2402), .A0(ofifoData[3]), .A1(ofifoData[259]), .A2(ofifoData[515]), .Z(n2398));
Q_MX02 U7515 ( .S(n2141), .A0(n2135), .A1(n2136), .Z(ofifoDataN[3]));
Q_AN02 U7516 ( .A0(n6720), .A1(shiftedXdata[4]), .Z(n2134));
Q_MX03 U7517 ( .S0(n2144), .S1(n2402), .A0(ofifoData[4]), .A1(ofifoData[260]), .A2(ofifoData[516]), .Z(n2397));
Q_MX02 U7518 ( .S(n2141), .A0(n2133), .A1(n2134), .Z(ofifoDataN[4]));
Q_AN02 U7519 ( .A0(n6720), .A1(shiftedXdata[5]), .Z(n2132));
Q_MX03 U7520 ( .S0(n2144), .S1(n2402), .A0(ofifoData[5]), .A1(ofifoData[261]), .A2(ofifoData[517]), .Z(n2396));
Q_MX02 U7521 ( .S(n2141), .A0(n2131), .A1(n2132), .Z(ofifoDataN[5]));
Q_AN02 U7522 ( .A0(n6720), .A1(shiftedXdata[6]), .Z(n2130));
Q_MX03 U7523 ( .S0(n2144), .S1(n2402), .A0(ofifoData[6]), .A1(ofifoData[262]), .A2(ofifoData[518]), .Z(n2395));
Q_MX02 U7524 ( .S(n2141), .A0(n2129), .A1(n2130), .Z(ofifoDataN[6]));
Q_AN02 U7525 ( .A0(n6720), .A1(shiftedXdata[7]), .Z(n2128));
Q_MX03 U7526 ( .S0(n2144), .S1(n2402), .A0(ofifoData[7]), .A1(ofifoData[263]), .A2(ofifoData[519]), .Z(n2394));
Q_MX02 U7527 ( .S(n2141), .A0(n2127), .A1(n2128), .Z(ofifoDataN[7]));
Q_AN02 U7528 ( .A0(n6720), .A1(shiftedXdata[8]), .Z(n2126));
Q_MX03 U7529 ( .S0(n2144), .S1(n2402), .A0(ofifoData[8]), .A1(ofifoData[264]), .A2(ofifoData[520]), .Z(n2393));
Q_MX02 U7530 ( .S(n2141), .A0(n2125), .A1(n2126), .Z(ofifoDataN[8]));
Q_AN02 U7531 ( .A0(n6720), .A1(shiftedXdata[9]), .Z(n2124));
Q_MX03 U7532 ( .S0(n2144), .S1(n2402), .A0(ofifoData[9]), .A1(ofifoData[265]), .A2(ofifoData[521]), .Z(n2392));
Q_MX02 U7533 ( .S(n2141), .A0(n2123), .A1(n2124), .Z(ofifoDataN[9]));
Q_AN02 U7534 ( .A0(n6720), .A1(shiftedXdata[10]), .Z(n2122));
Q_MX03 U7535 ( .S0(n2144), .S1(n2402), .A0(ofifoData[10]), .A1(ofifoData[266]), .A2(ofifoData[522]), .Z(n2391));
Q_MX02 U7536 ( .S(n2141), .A0(n2121), .A1(n2122), .Z(ofifoDataN[10]));
Q_AN02 U7537 ( .A0(n6720), .A1(shiftedXdata[11]), .Z(n2120));
Q_MX03 U7538 ( .S0(n2144), .S1(n2402), .A0(ofifoData[11]), .A1(ofifoData[267]), .A2(ofifoData[523]), .Z(n2390));
Q_MX02 U7539 ( .S(n2141), .A0(n2119), .A1(n2120), .Z(ofifoDataN[11]));
Q_AN02 U7540 ( .A0(n6720), .A1(shiftedXdata[12]), .Z(n2118));
Q_MX03 U7541 ( .S0(n2144), .S1(n2402), .A0(ofifoData[12]), .A1(ofifoData[268]), .A2(ofifoData[524]), .Z(n2389));
Q_MX02 U7542 ( .S(n2141), .A0(n2117), .A1(n2118), .Z(ofifoDataN[12]));
Q_AN02 U7543 ( .A0(n6720), .A1(shiftedXdata[13]), .Z(n2116));
Q_MX03 U7544 ( .S0(n2144), .S1(n2402), .A0(ofifoData[13]), .A1(ofifoData[269]), .A2(ofifoData[525]), .Z(n2388));
Q_MX02 U7545 ( .S(n2141), .A0(n2115), .A1(n2116), .Z(ofifoDataN[13]));
Q_AN02 U7546 ( .A0(n6720), .A1(shiftedXdata[14]), .Z(n2114));
Q_MX03 U7547 ( .S0(n2144), .S1(n2402), .A0(ofifoData[14]), .A1(ofifoData[270]), .A2(ofifoData[526]), .Z(n2387));
Q_MX02 U7548 ( .S(n2141), .A0(n2113), .A1(n2114), .Z(ofifoDataN[14]));
Q_AN02 U7549 ( .A0(n6720), .A1(shiftedXdata[15]), .Z(n2112));
Q_MX03 U7550 ( .S0(n2144), .S1(n2402), .A0(ofifoData[15]), .A1(ofifoData[271]), .A2(ofifoData[527]), .Z(n2386));
Q_MX02 U7551 ( .S(n2141), .A0(n2111), .A1(n2112), .Z(ofifoDataN[15]));
Q_AN02 U7552 ( .A0(n6720), .A1(shiftedXdata[16]), .Z(n2110));
Q_MX03 U7553 ( .S0(n2144), .S1(n2402), .A0(ofifoData[16]), .A1(ofifoData[272]), .A2(ofifoData[528]), .Z(n2385));
Q_MX02 U7554 ( .S(n2141), .A0(n2109), .A1(n2110), .Z(ofifoDataN[16]));
Q_AN02 U7555 ( .A0(n6720), .A1(shiftedXdata[17]), .Z(n2108));
Q_MX03 U7556 ( .S0(n2144), .S1(n2402), .A0(ofifoData[17]), .A1(ofifoData[273]), .A2(ofifoData[529]), .Z(n2384));
Q_MX02 U7557 ( .S(n2141), .A0(n2107), .A1(n2108), .Z(ofifoDataN[17]));
Q_AN02 U7558 ( .A0(n6720), .A1(shiftedXdata[18]), .Z(n2106));
Q_MX03 U7559 ( .S0(n2144), .S1(n2402), .A0(ofifoData[18]), .A1(ofifoData[274]), .A2(ofifoData[530]), .Z(n2383));
Q_MX02 U7560 ( .S(n2141), .A0(n2105), .A1(n2106), .Z(ofifoDataN[18]));
Q_AN02 U7561 ( .A0(n6720), .A1(shiftedXdata[19]), .Z(n2104));
Q_MX03 U7562 ( .S0(n2144), .S1(n2402), .A0(ofifoData[19]), .A1(ofifoData[275]), .A2(ofifoData[531]), .Z(n2382));
Q_MX02 U7563 ( .S(n2141), .A0(n2103), .A1(n2104), .Z(ofifoDataN[19]));
Q_AN02 U7564 ( .A0(n6720), .A1(shiftedXdata[20]), .Z(n2102));
Q_MX03 U7565 ( .S0(n2144), .S1(n2402), .A0(ofifoData[20]), .A1(ofifoData[276]), .A2(ofifoData[532]), .Z(n2381));
Q_MX02 U7566 ( .S(n2141), .A0(n2101), .A1(n2102), .Z(ofifoDataN[20]));
Q_AN02 U7567 ( .A0(n6720), .A1(shiftedXdata[21]), .Z(n2100));
Q_MX03 U7568 ( .S0(n2144), .S1(n2402), .A0(ofifoData[21]), .A1(ofifoData[277]), .A2(ofifoData[533]), .Z(n2380));
Q_MX02 U7569 ( .S(n2141), .A0(n2099), .A1(n2100), .Z(ofifoDataN[21]));
Q_AN02 U7570 ( .A0(n6720), .A1(shiftedXdata[22]), .Z(n2098));
Q_MX03 U7571 ( .S0(n2144), .S1(n2402), .A0(ofifoData[22]), .A1(ofifoData[278]), .A2(ofifoData[534]), .Z(n2379));
Q_MX02 U7572 ( .S(n2141), .A0(n2097), .A1(n2098), .Z(ofifoDataN[22]));
Q_AN02 U7573 ( .A0(n6720), .A1(shiftedXdata[23]), .Z(n2096));
Q_MX03 U7574 ( .S0(n2144), .S1(n2402), .A0(ofifoData[23]), .A1(ofifoData[279]), .A2(ofifoData[535]), .Z(n2378));
Q_MX02 U7575 ( .S(n2141), .A0(n2095), .A1(n2096), .Z(ofifoDataN[23]));
Q_AN02 U7576 ( .A0(n6720), .A1(shiftedXdata[24]), .Z(n2094));
Q_MX03 U7577 ( .S0(n2144), .S1(n2402), .A0(ofifoData[24]), .A1(ofifoData[280]), .A2(ofifoData[536]), .Z(n2377));
Q_MX02 U7578 ( .S(n2141), .A0(n2093), .A1(n2094), .Z(ofifoDataN[24]));
Q_AN02 U7579 ( .A0(n6720), .A1(shiftedXdata[25]), .Z(n2092));
Q_MX03 U7580 ( .S0(n2144), .S1(n2402), .A0(ofifoData[25]), .A1(ofifoData[281]), .A2(ofifoData[537]), .Z(n2376));
Q_MX02 U7581 ( .S(n2141), .A0(n2091), .A1(n2092), .Z(ofifoDataN[25]));
Q_AN02 U7582 ( .A0(n6720), .A1(shiftedXdata[26]), .Z(n2090));
Q_MX03 U7583 ( .S0(n2144), .S1(n2402), .A0(ofifoData[26]), .A1(ofifoData[282]), .A2(ofifoData[538]), .Z(n2375));
Q_MX02 U7584 ( .S(n2141), .A0(n2089), .A1(n2090), .Z(ofifoDataN[26]));
Q_AN02 U7585 ( .A0(n6720), .A1(shiftedXdata[27]), .Z(n2088));
Q_MX03 U7586 ( .S0(n2144), .S1(n2402), .A0(ofifoData[27]), .A1(ofifoData[283]), .A2(ofifoData[539]), .Z(n2374));
Q_MX02 U7587 ( .S(n2141), .A0(n2087), .A1(n2088), .Z(ofifoDataN[27]));
Q_AN02 U7588 ( .A0(n6720), .A1(shiftedXdata[28]), .Z(n2086));
Q_MX03 U7589 ( .S0(n2144), .S1(n2402), .A0(ofifoData[28]), .A1(ofifoData[284]), .A2(ofifoData[540]), .Z(n2373));
Q_MX02 U7590 ( .S(n2141), .A0(n2085), .A1(n2086), .Z(ofifoDataN[28]));
Q_AN02 U7591 ( .A0(n6720), .A1(shiftedXdata[29]), .Z(n2084));
Q_MX03 U7592 ( .S0(n2144), .S1(n2402), .A0(ofifoData[29]), .A1(ofifoData[285]), .A2(ofifoData[541]), .Z(n2372));
Q_MX02 U7593 ( .S(n2141), .A0(n2083), .A1(n2084), .Z(ofifoDataN[29]));
Q_AN02 U7594 ( .A0(n6720), .A1(shiftedXdata[30]), .Z(n2082));
Q_MX03 U7595 ( .S0(n2144), .S1(n2402), .A0(ofifoData[30]), .A1(ofifoData[286]), .A2(ofifoData[542]), .Z(n2371));
Q_MX02 U7596 ( .S(n2141), .A0(n2081), .A1(n2082), .Z(ofifoDataN[30]));
Q_AN02 U7597 ( .A0(n6720), .A1(shiftedXdata[31]), .Z(n2080));
Q_MX03 U7598 ( .S0(n2144), .S1(n2402), .A0(ofifoData[31]), .A1(ofifoData[287]), .A2(ofifoData[543]), .Z(n2370));
Q_MX02 U7599 ( .S(n2141), .A0(n2079), .A1(n2080), .Z(ofifoDataN[31]));
Q_AN02 U7600 ( .A0(n6720), .A1(shiftedXdata[32]), .Z(n2078));
Q_MX03 U7601 ( .S0(n2144), .S1(n2402), .A0(ofifoData[32]), .A1(ofifoData[288]), .A2(ofifoData[544]), .Z(n2369));
Q_MX02 U7602 ( .S(n2141), .A0(n2077), .A1(n2078), .Z(ofifoDataN[32]));
Q_AN02 U7603 ( .A0(n6720), .A1(shiftedXdata[33]), .Z(n2076));
Q_MX03 U7604 ( .S0(n2144), .S1(n2402), .A0(ofifoData[33]), .A1(ofifoData[289]), .A2(ofifoData[545]), .Z(n2368));
Q_MX02 U7605 ( .S(n2141), .A0(n2075), .A1(n2076), .Z(ofifoDataN[33]));
Q_AN02 U7606 ( .A0(n6720), .A1(shiftedXdata[34]), .Z(n2074));
Q_MX03 U7607 ( .S0(n2144), .S1(n2402), .A0(ofifoData[34]), .A1(ofifoData[290]), .A2(ofifoData[546]), .Z(n2367));
Q_MX02 U7608 ( .S(n2141), .A0(n2073), .A1(n2074), .Z(ofifoDataN[34]));
Q_AN02 U7609 ( .A0(n6720), .A1(shiftedXdata[35]), .Z(n2072));
Q_MX03 U7610 ( .S0(n2144), .S1(n2402), .A0(ofifoData[35]), .A1(ofifoData[291]), .A2(ofifoData[547]), .Z(n2366));
Q_MX02 U7611 ( .S(n2141), .A0(n2071), .A1(n2072), .Z(ofifoDataN[35]));
Q_AN02 U7612 ( .A0(n6720), .A1(shiftedXdata[36]), .Z(n2070));
Q_MX03 U7613 ( .S0(n2144), .S1(n2402), .A0(ofifoData[36]), .A1(ofifoData[292]), .A2(ofifoData[548]), .Z(n2365));
Q_MX02 U7614 ( .S(n2141), .A0(n2069), .A1(n2070), .Z(ofifoDataN[36]));
Q_AN02 U7615 ( .A0(n6720), .A1(shiftedXdata[37]), .Z(n2068));
Q_MX03 U7616 ( .S0(n2144), .S1(n2402), .A0(ofifoData[37]), .A1(ofifoData[293]), .A2(ofifoData[549]), .Z(n2364));
Q_MX02 U7617 ( .S(n2141), .A0(n2067), .A1(n2068), .Z(ofifoDataN[37]));
Q_AN02 U7618 ( .A0(n6720), .A1(shiftedXdata[38]), .Z(n2066));
Q_MX03 U7619 ( .S0(n2144), .S1(n2402), .A0(ofifoData[38]), .A1(ofifoData[294]), .A2(ofifoData[550]), .Z(n2363));
Q_MX02 U7620 ( .S(n2141), .A0(n2065), .A1(n2066), .Z(ofifoDataN[38]));
Q_AN02 U7621 ( .A0(n6720), .A1(shiftedXdata[39]), .Z(n2064));
Q_MX03 U7622 ( .S0(n2144), .S1(n2402), .A0(ofifoData[39]), .A1(ofifoData[295]), .A2(ofifoData[551]), .Z(n2362));
Q_MX02 U7623 ( .S(n2141), .A0(n2063), .A1(n2064), .Z(ofifoDataN[39]));
Q_AN02 U7624 ( .A0(n6720), .A1(shiftedXdata[40]), .Z(n2062));
Q_MX03 U7625 ( .S0(n2144), .S1(n2402), .A0(ofifoData[40]), .A1(ofifoData[296]), .A2(ofifoData[552]), .Z(n2361));
Q_MX02 U7626 ( .S(n2141), .A0(n2061), .A1(n2062), .Z(ofifoDataN[40]));
Q_AN02 U7627 ( .A0(n6720), .A1(shiftedXdata[41]), .Z(n2060));
Q_MX03 U7628 ( .S0(n2144), .S1(n2402), .A0(ofifoData[41]), .A1(ofifoData[297]), .A2(ofifoData[553]), .Z(n2360));
Q_MX02 U7629 ( .S(n2141), .A0(n2059), .A1(n2060), .Z(ofifoDataN[41]));
Q_AN02 U7630 ( .A0(n6720), .A1(shiftedXdata[42]), .Z(n2058));
Q_MX03 U7631 ( .S0(n2144), .S1(n2402), .A0(ofifoData[42]), .A1(ofifoData[298]), .A2(ofifoData[554]), .Z(n2359));
Q_MX02 U7632 ( .S(n2141), .A0(n2057), .A1(n2058), .Z(ofifoDataN[42]));
Q_AN02 U7633 ( .A0(n6720), .A1(shiftedXdata[43]), .Z(n2056));
Q_MX03 U7634 ( .S0(n2144), .S1(n2402), .A0(ofifoData[43]), .A1(ofifoData[299]), .A2(ofifoData[555]), .Z(n2358));
Q_MX02 U7635 ( .S(n2141), .A0(n2055), .A1(n2056), .Z(ofifoDataN[43]));
Q_AN02 U7636 ( .A0(n6720), .A1(shiftedXdata[44]), .Z(n2054));
Q_MX03 U7637 ( .S0(n2144), .S1(n2402), .A0(ofifoData[44]), .A1(ofifoData[300]), .A2(ofifoData[556]), .Z(n2357));
Q_MX02 U7638 ( .S(n2141), .A0(n2053), .A1(n2054), .Z(ofifoDataN[44]));
Q_AN02 U7639 ( .A0(n6720), .A1(shiftedXdata[45]), .Z(n2052));
Q_MX03 U7640 ( .S0(n2144), .S1(n2402), .A0(ofifoData[45]), .A1(ofifoData[301]), .A2(ofifoData[557]), .Z(n2356));
Q_MX02 U7641 ( .S(n2141), .A0(n2051), .A1(n2052), .Z(ofifoDataN[45]));
Q_AN02 U7642 ( .A0(n6720), .A1(shiftedXdata[46]), .Z(n2050));
Q_MX03 U7643 ( .S0(n2144), .S1(n2402), .A0(ofifoData[46]), .A1(ofifoData[302]), .A2(ofifoData[558]), .Z(n2355));
Q_MX02 U7644 ( .S(n2141), .A0(n2049), .A1(n2050), .Z(ofifoDataN[46]));
Q_AN02 U7645 ( .A0(n6720), .A1(shiftedXdata[47]), .Z(n2048));
Q_MX03 U7646 ( .S0(n2144), .S1(n2402), .A0(ofifoData[47]), .A1(ofifoData[303]), .A2(ofifoData[559]), .Z(n2354));
Q_MX02 U7647 ( .S(n2141), .A0(n2047), .A1(n2048), .Z(ofifoDataN[47]));
Q_AN02 U7648 ( .A0(n6720), .A1(shiftedXdata[48]), .Z(n2046));
Q_MX03 U7649 ( .S0(n2144), .S1(n2402), .A0(ofifoData[48]), .A1(ofifoData[304]), .A2(ofifoData[560]), .Z(n2353));
Q_MX02 U7650 ( .S(n2141), .A0(n2045), .A1(n2046), .Z(ofifoDataN[48]));
Q_AN02 U7651 ( .A0(n6720), .A1(shiftedXdata[49]), .Z(n2044));
Q_MX03 U7652 ( .S0(n2144), .S1(n2402), .A0(ofifoData[49]), .A1(ofifoData[305]), .A2(ofifoData[561]), .Z(n2352));
Q_MX02 U7653 ( .S(n2141), .A0(n2043), .A1(n2044), .Z(ofifoDataN[49]));
Q_AN02 U7654 ( .A0(n6720), .A1(shiftedXdata[50]), .Z(n2042));
Q_MX03 U7655 ( .S0(n2144), .S1(n2402), .A0(ofifoData[50]), .A1(ofifoData[306]), .A2(ofifoData[562]), .Z(n2351));
Q_MX02 U7656 ( .S(n2141), .A0(n2041), .A1(n2042), .Z(ofifoDataN[50]));
Q_AN02 U7657 ( .A0(n6720), .A1(shiftedXdata[51]), .Z(n2040));
Q_MX03 U7658 ( .S0(n2144), .S1(n2402), .A0(ofifoData[51]), .A1(ofifoData[307]), .A2(ofifoData[563]), .Z(n2350));
Q_MX02 U7659 ( .S(n2141), .A0(n2039), .A1(n2040), .Z(ofifoDataN[51]));
Q_AN02 U7660 ( .A0(n6720), .A1(shiftedXdata[52]), .Z(n2038));
Q_MX03 U7661 ( .S0(n2144), .S1(n2402), .A0(ofifoData[52]), .A1(ofifoData[308]), .A2(ofifoData[564]), .Z(n2349));
Q_MX02 U7662 ( .S(n2141), .A0(n2037), .A1(n2038), .Z(ofifoDataN[52]));
Q_AN02 U7663 ( .A0(n6720), .A1(shiftedXdata[53]), .Z(n2036));
Q_MX03 U7664 ( .S0(n2144), .S1(n2402), .A0(ofifoData[53]), .A1(ofifoData[309]), .A2(ofifoData[565]), .Z(n2348));
Q_MX02 U7665 ( .S(n2141), .A0(n2035), .A1(n2036), .Z(ofifoDataN[53]));
Q_AN02 U7666 ( .A0(n6720), .A1(shiftedXdata[54]), .Z(n2034));
Q_MX03 U7667 ( .S0(n2144), .S1(n2402), .A0(ofifoData[54]), .A1(ofifoData[310]), .A2(ofifoData[566]), .Z(n2347));
Q_MX02 U7668 ( .S(n2141), .A0(n2033), .A1(n2034), .Z(ofifoDataN[54]));
Q_AN02 U7669 ( .A0(n6720), .A1(shiftedXdata[55]), .Z(n2032));
Q_MX03 U7670 ( .S0(n2144), .S1(n2402), .A0(ofifoData[55]), .A1(ofifoData[311]), .A2(ofifoData[567]), .Z(n2346));
Q_MX02 U7671 ( .S(n2141), .A0(n2031), .A1(n2032), .Z(ofifoDataN[55]));
Q_AN02 U7672 ( .A0(n6720), .A1(shiftedXdata[56]), .Z(n2030));
Q_MX03 U7673 ( .S0(n2144), .S1(n2402), .A0(ofifoData[56]), .A1(ofifoData[312]), .A2(ofifoData[568]), .Z(n2345));
Q_MX02 U7674 ( .S(n2141), .A0(n2029), .A1(n2030), .Z(ofifoDataN[56]));
Q_AN02 U7675 ( .A0(n6720), .A1(shiftedXdata[57]), .Z(n2028));
Q_MX03 U7676 ( .S0(n2144), .S1(n2402), .A0(ofifoData[57]), .A1(ofifoData[313]), .A2(ofifoData[569]), .Z(n2344));
Q_MX02 U7677 ( .S(n2141), .A0(n2027), .A1(n2028), .Z(ofifoDataN[57]));
Q_AN02 U7678 ( .A0(n6720), .A1(shiftedXdata[58]), .Z(n2026));
Q_MX03 U7679 ( .S0(n2144), .S1(n2402), .A0(ofifoData[58]), .A1(ofifoData[314]), .A2(ofifoData[570]), .Z(n2343));
Q_MX02 U7680 ( .S(n2141), .A0(n2025), .A1(n2026), .Z(ofifoDataN[58]));
Q_AN02 U7681 ( .A0(n6720), .A1(shiftedXdata[59]), .Z(n2024));
Q_MX03 U7682 ( .S0(n2144), .S1(n2402), .A0(ofifoData[59]), .A1(ofifoData[315]), .A2(ofifoData[571]), .Z(n2342));
Q_MX02 U7683 ( .S(n2141), .A0(n2023), .A1(n2024), .Z(ofifoDataN[59]));
Q_AN02 U7684 ( .A0(n6720), .A1(shiftedXdata[60]), .Z(n2022));
Q_MX03 U7685 ( .S0(n2144), .S1(n2402), .A0(ofifoData[60]), .A1(ofifoData[316]), .A2(ofifoData[572]), .Z(n2341));
Q_MX02 U7686 ( .S(n2141), .A0(n2021), .A1(n2022), .Z(ofifoDataN[60]));
Q_AN02 U7687 ( .A0(n6720), .A1(shiftedXdata[61]), .Z(n2020));
Q_MX03 U7688 ( .S0(n2144), .S1(n2402), .A0(ofifoData[61]), .A1(ofifoData[317]), .A2(ofifoData[573]), .Z(n2340));
Q_MX02 U7689 ( .S(n2141), .A0(n2019), .A1(n2020), .Z(ofifoDataN[61]));
Q_AN02 U7690 ( .A0(n6720), .A1(shiftedXdata[62]), .Z(n2018));
Q_MX03 U7691 ( .S0(n2144), .S1(n2402), .A0(ofifoData[62]), .A1(ofifoData[318]), .A2(ofifoData[574]), .Z(n2339));
Q_MX02 U7692 ( .S(n2141), .A0(n2017), .A1(n2018), .Z(ofifoDataN[62]));
Q_AN02 U7693 ( .A0(n6720), .A1(shiftedXdata[63]), .Z(n2016));
Q_MX03 U7694 ( .S0(n2144), .S1(n2402), .A0(ofifoData[63]), .A1(ofifoData[319]), .A2(ofifoData[575]), .Z(n2338));
Q_MX02 U7695 ( .S(n2141), .A0(n2015), .A1(n2016), .Z(ofifoDataN[63]));
Q_AN02 U7696 ( .A0(n6720), .A1(shiftedXdata[64]), .Z(n2014));
Q_MX03 U7697 ( .S0(n2144), .S1(n2402), .A0(ofifoData[64]), .A1(ofifoData[320]), .A2(ofifoData[576]), .Z(n2337));
Q_MX02 U7698 ( .S(n2141), .A0(n2013), .A1(n2014), .Z(ofifoDataN[64]));
Q_AN02 U7699 ( .A0(n6720), .A1(shiftedXdata[65]), .Z(n2012));
Q_MX03 U7700 ( .S0(n2144), .S1(n2402), .A0(ofifoData[65]), .A1(ofifoData[321]), .A2(ofifoData[577]), .Z(n2336));
Q_MX02 U7701 ( .S(n2141), .A0(n2011), .A1(n2012), .Z(ofifoDataN[65]));
Q_AN02 U7702 ( .A0(n6720), .A1(shiftedXdata[66]), .Z(n2010));
Q_MX03 U7703 ( .S0(n2144), .S1(n2402), .A0(ofifoData[66]), .A1(ofifoData[322]), .A2(ofifoData[578]), .Z(n2335));
Q_MX02 U7704 ( .S(n2141), .A0(n2009), .A1(n2010), .Z(ofifoDataN[66]));
Q_AN02 U7705 ( .A0(n6720), .A1(shiftedXdata[67]), .Z(n2008));
Q_MX03 U7706 ( .S0(n2144), .S1(n2402), .A0(ofifoData[67]), .A1(ofifoData[323]), .A2(ofifoData[579]), .Z(n2334));
Q_MX02 U7707 ( .S(n2141), .A0(n2007), .A1(n2008), .Z(ofifoDataN[67]));
Q_AN02 U7708 ( .A0(n6720), .A1(shiftedXdata[68]), .Z(n2006));
Q_MX03 U7709 ( .S0(n2144), .S1(n2402), .A0(ofifoData[68]), .A1(ofifoData[324]), .A2(ofifoData[580]), .Z(n2333));
Q_MX02 U7710 ( .S(n2141), .A0(n2005), .A1(n2006), .Z(ofifoDataN[68]));
Q_AN02 U7711 ( .A0(n6720), .A1(shiftedXdata[69]), .Z(n2004));
Q_MX03 U7712 ( .S0(n2144), .S1(n2402), .A0(ofifoData[69]), .A1(ofifoData[325]), .A2(ofifoData[581]), .Z(n2332));
Q_MX02 U7713 ( .S(n2141), .A0(n2003), .A1(n2004), .Z(ofifoDataN[69]));
Q_AN02 U7714 ( .A0(n6720), .A1(shiftedXdata[70]), .Z(n2002));
Q_MX03 U7715 ( .S0(n2144), .S1(n2402), .A0(ofifoData[70]), .A1(ofifoData[326]), .A2(ofifoData[582]), .Z(n2331));
Q_MX02 U7716 ( .S(n2141), .A0(n2001), .A1(n2002), .Z(ofifoDataN[70]));
Q_AN02 U7717 ( .A0(n6720), .A1(shiftedXdata[71]), .Z(n2000));
Q_MX03 U7718 ( .S0(n2144), .S1(n2402), .A0(ofifoData[71]), .A1(ofifoData[327]), .A2(ofifoData[583]), .Z(n2330));
Q_MX02 U7719 ( .S(n2141), .A0(n1999), .A1(n2000), .Z(ofifoDataN[71]));
Q_AN02 U7720 ( .A0(n6720), .A1(shiftedXdata[72]), .Z(n1998));
Q_MX03 U7721 ( .S0(n2144), .S1(n2402), .A0(ofifoData[72]), .A1(ofifoData[328]), .A2(ofifoData[584]), .Z(n2329));
Q_MX02 U7722 ( .S(n2141), .A0(n1997), .A1(n1998), .Z(ofifoDataN[72]));
Q_AN02 U7723 ( .A0(n6720), .A1(shiftedXdata[73]), .Z(n1996));
Q_MX03 U7724 ( .S0(n2144), .S1(n2402), .A0(ofifoData[73]), .A1(ofifoData[329]), .A2(ofifoData[585]), .Z(n2328));
Q_MX02 U7725 ( .S(n2141), .A0(n1995), .A1(n1996), .Z(ofifoDataN[73]));
Q_AN02 U7726 ( .A0(n6720), .A1(shiftedXdata[74]), .Z(n1994));
Q_MX03 U7727 ( .S0(n2144), .S1(n2402), .A0(ofifoData[74]), .A1(ofifoData[330]), .A2(ofifoData[586]), .Z(n2327));
Q_MX02 U7728 ( .S(n2141), .A0(n1993), .A1(n1994), .Z(ofifoDataN[74]));
Q_AN02 U7729 ( .A0(n6720), .A1(shiftedXdata[75]), .Z(n1992));
Q_MX03 U7730 ( .S0(n2144), .S1(n2402), .A0(ofifoData[75]), .A1(ofifoData[331]), .A2(ofifoData[587]), .Z(n2326));
Q_MX02 U7731 ( .S(n2141), .A0(n1991), .A1(n1992), .Z(ofifoDataN[75]));
Q_AN02 U7732 ( .A0(n6720), .A1(shiftedXdata[76]), .Z(n1990));
Q_MX03 U7733 ( .S0(n2144), .S1(n2402), .A0(ofifoData[76]), .A1(ofifoData[332]), .A2(ofifoData[588]), .Z(n2325));
Q_MX02 U7734 ( .S(n2141), .A0(n1989), .A1(n1990), .Z(ofifoDataN[76]));
Q_AN02 U7735 ( .A0(n6720), .A1(shiftedXdata[77]), .Z(n1988));
Q_MX03 U7736 ( .S0(n2144), .S1(n2402), .A0(ofifoData[77]), .A1(ofifoData[333]), .A2(ofifoData[589]), .Z(n2324));
Q_MX02 U7737 ( .S(n2141), .A0(n1987), .A1(n1988), .Z(ofifoDataN[77]));
Q_AN02 U7738 ( .A0(n6720), .A1(shiftedXdata[78]), .Z(n1986));
Q_MX03 U7739 ( .S0(n2144), .S1(n2402), .A0(ofifoData[78]), .A1(ofifoData[334]), .A2(ofifoData[590]), .Z(n2323));
Q_MX02 U7740 ( .S(n2141), .A0(n1985), .A1(n1986), .Z(ofifoDataN[78]));
Q_AN02 U7741 ( .A0(n6720), .A1(shiftedXdata[79]), .Z(n1984));
Q_MX03 U7742 ( .S0(n2144), .S1(n2402), .A0(ofifoData[79]), .A1(ofifoData[335]), .A2(ofifoData[591]), .Z(n2322));
Q_MX02 U7743 ( .S(n2141), .A0(n1983), .A1(n1984), .Z(ofifoDataN[79]));
Q_AN02 U7744 ( .A0(n6720), .A1(shiftedXdata[80]), .Z(n1982));
Q_MX03 U7745 ( .S0(n2144), .S1(n2402), .A0(ofifoData[80]), .A1(ofifoData[336]), .A2(ofifoData[592]), .Z(n2321));
Q_MX02 U7746 ( .S(n2141), .A0(n1981), .A1(n1982), .Z(ofifoDataN[80]));
Q_AN02 U7747 ( .A0(n6720), .A1(shiftedXdata[81]), .Z(n1980));
Q_MX03 U7748 ( .S0(n2144), .S1(n2402), .A0(ofifoData[81]), .A1(ofifoData[337]), .A2(ofifoData[593]), .Z(n2320));
Q_MX02 U7749 ( .S(n2141), .A0(n1979), .A1(n1980), .Z(ofifoDataN[81]));
Q_AN02 U7750 ( .A0(n6720), .A1(shiftedXdata[82]), .Z(n1978));
Q_MX03 U7751 ( .S0(n2144), .S1(n2402), .A0(ofifoData[82]), .A1(ofifoData[338]), .A2(ofifoData[594]), .Z(n2319));
Q_MX02 U7752 ( .S(n2141), .A0(n1977), .A1(n1978), .Z(ofifoDataN[82]));
Q_AN02 U7753 ( .A0(n6720), .A1(shiftedXdata[83]), .Z(n1976));
Q_MX03 U7754 ( .S0(n2144), .S1(n2402), .A0(ofifoData[83]), .A1(ofifoData[339]), .A2(ofifoData[595]), .Z(n2318));
Q_MX02 U7755 ( .S(n2141), .A0(n1975), .A1(n1976), .Z(ofifoDataN[83]));
Q_AN02 U7756 ( .A0(n6720), .A1(shiftedXdata[84]), .Z(n1974));
Q_MX03 U7757 ( .S0(n2144), .S1(n2402), .A0(ofifoData[84]), .A1(ofifoData[340]), .A2(ofifoData[596]), .Z(n2317));
Q_MX02 U7758 ( .S(n2141), .A0(n1973), .A1(n1974), .Z(ofifoDataN[84]));
Q_AN02 U7759 ( .A0(n6720), .A1(shiftedXdata[85]), .Z(n1972));
Q_MX03 U7760 ( .S0(n2144), .S1(n2402), .A0(ofifoData[85]), .A1(ofifoData[341]), .A2(ofifoData[597]), .Z(n2316));
Q_MX02 U7761 ( .S(n2141), .A0(n1971), .A1(n1972), .Z(ofifoDataN[85]));
Q_AN02 U7762 ( .A0(n6720), .A1(shiftedXdata[86]), .Z(n1970));
Q_MX03 U7763 ( .S0(n2144), .S1(n2402), .A0(ofifoData[86]), .A1(ofifoData[342]), .A2(ofifoData[598]), .Z(n2315));
Q_MX02 U7764 ( .S(n2141), .A0(n1969), .A1(n1970), .Z(ofifoDataN[86]));
Q_AN02 U7765 ( .A0(n6720), .A1(shiftedXdata[87]), .Z(n1968));
Q_MX03 U7766 ( .S0(n2144), .S1(n2402), .A0(ofifoData[87]), .A1(ofifoData[343]), .A2(ofifoData[599]), .Z(n2314));
Q_MX02 U7767 ( .S(n2141), .A0(n1967), .A1(n1968), .Z(ofifoDataN[87]));
Q_AN02 U7768 ( .A0(n6720), .A1(shiftedXdata[88]), .Z(n1966));
Q_MX03 U7769 ( .S0(n2144), .S1(n2402), .A0(ofifoData[88]), .A1(ofifoData[344]), .A2(ofifoData[600]), .Z(n2313));
Q_MX02 U7770 ( .S(n2141), .A0(n1965), .A1(n1966), .Z(ofifoDataN[88]));
Q_AN02 U7771 ( .A0(n6720), .A1(shiftedXdata[89]), .Z(n1964));
Q_MX03 U7772 ( .S0(n2144), .S1(n2402), .A0(ofifoData[89]), .A1(ofifoData[345]), .A2(ofifoData[601]), .Z(n2312));
Q_MX02 U7773 ( .S(n2141), .A0(n1963), .A1(n1964), .Z(ofifoDataN[89]));
Q_AN02 U7774 ( .A0(n6720), .A1(shiftedXdata[90]), .Z(n1962));
Q_MX03 U7775 ( .S0(n2144), .S1(n2402), .A0(ofifoData[90]), .A1(ofifoData[346]), .A2(ofifoData[602]), .Z(n2311));
Q_MX02 U7776 ( .S(n2141), .A0(n1961), .A1(n1962), .Z(ofifoDataN[90]));
Q_AN02 U7777 ( .A0(n6720), .A1(shiftedXdata[91]), .Z(n1960));
Q_MX03 U7778 ( .S0(n2144), .S1(n2402), .A0(ofifoData[91]), .A1(ofifoData[347]), .A2(ofifoData[603]), .Z(n2310));
Q_MX02 U7779 ( .S(n2141), .A0(n1959), .A1(n1960), .Z(ofifoDataN[91]));
Q_AN02 U7780 ( .A0(n6720), .A1(shiftedXdata[92]), .Z(n1958));
Q_MX03 U7781 ( .S0(n2144), .S1(n2402), .A0(ofifoData[92]), .A1(ofifoData[348]), .A2(ofifoData[604]), .Z(n2309));
Q_MX02 U7782 ( .S(n2141), .A0(n1957), .A1(n1958), .Z(ofifoDataN[92]));
Q_AN02 U7783 ( .A0(n6720), .A1(shiftedXdata[93]), .Z(n1956));
Q_MX03 U7784 ( .S0(n2144), .S1(n2402), .A0(ofifoData[93]), .A1(ofifoData[349]), .A2(ofifoData[605]), .Z(n2308));
Q_MX02 U7785 ( .S(n2141), .A0(n1955), .A1(n1956), .Z(ofifoDataN[93]));
Q_AN02 U7786 ( .A0(n6720), .A1(shiftedXdata[94]), .Z(n1954));
Q_MX03 U7787 ( .S0(n2144), .S1(n2402), .A0(ofifoData[94]), .A1(ofifoData[350]), .A2(ofifoData[606]), .Z(n2307));
Q_MX02 U7788 ( .S(n2141), .A0(n1953), .A1(n1954), .Z(ofifoDataN[94]));
Q_AN02 U7789 ( .A0(n6720), .A1(shiftedXdata[95]), .Z(n1952));
Q_MX03 U7790 ( .S0(n2144), .S1(n2402), .A0(ofifoData[95]), .A1(ofifoData[351]), .A2(ofifoData[607]), .Z(n2306));
Q_MX02 U7791 ( .S(n2141), .A0(n1951), .A1(n1952), .Z(ofifoDataN[95]));
Q_AN02 U7792 ( .A0(n6720), .A1(shiftedXdata[96]), .Z(n1950));
Q_MX03 U7793 ( .S0(n2144), .S1(n2402), .A0(ofifoData[96]), .A1(ofifoData[352]), .A2(ofifoData[608]), .Z(n2305));
Q_MX02 U7794 ( .S(n2141), .A0(n1949), .A1(n1950), .Z(ofifoDataN[96]));
Q_AN02 U7795 ( .A0(n6720), .A1(shiftedXdata[97]), .Z(n1948));
Q_MX03 U7796 ( .S0(n2144), .S1(n2402), .A0(ofifoData[97]), .A1(ofifoData[353]), .A2(ofifoData[609]), .Z(n2304));
Q_MX02 U7797 ( .S(n2141), .A0(n1947), .A1(n1948), .Z(ofifoDataN[97]));
Q_AN02 U7798 ( .A0(n6720), .A1(shiftedXdata[98]), .Z(n1946));
Q_MX03 U7799 ( .S0(n2144), .S1(n2402), .A0(ofifoData[98]), .A1(ofifoData[354]), .A2(ofifoData[610]), .Z(n2303));
Q_MX02 U7800 ( .S(n2141), .A0(n1945), .A1(n1946), .Z(ofifoDataN[98]));
Q_AN02 U7801 ( .A0(n6720), .A1(shiftedXdata[99]), .Z(n1944));
Q_MX03 U7802 ( .S0(n2144), .S1(n2402), .A0(ofifoData[99]), .A1(ofifoData[355]), .A2(ofifoData[611]), .Z(n2302));
Q_MX02 U7803 ( .S(n2141), .A0(n1943), .A1(n1944), .Z(ofifoDataN[99]));
Q_AN02 U7804 ( .A0(n6720), .A1(shiftedXdata[100]), .Z(n1942));
Q_MX03 U7805 ( .S0(n2144), .S1(n2402), .A0(ofifoData[100]), .A1(ofifoData[356]), .A2(ofifoData[612]), .Z(n2301));
Q_MX02 U7806 ( .S(n2141), .A0(n1941), .A1(n1942), .Z(ofifoDataN[100]));
Q_AN02 U7807 ( .A0(n6720), .A1(shiftedXdata[101]), .Z(n1940));
Q_MX03 U7808 ( .S0(n2144), .S1(n2402), .A0(ofifoData[101]), .A1(ofifoData[357]), .A2(ofifoData[613]), .Z(n2300));
Q_MX02 U7809 ( .S(n2141), .A0(n1939), .A1(n1940), .Z(ofifoDataN[101]));
Q_AN02 U7810 ( .A0(n6720), .A1(shiftedXdata[102]), .Z(n1938));
Q_MX03 U7811 ( .S0(n2144), .S1(n2402), .A0(ofifoData[102]), .A1(ofifoData[358]), .A2(ofifoData[614]), .Z(n2299));
Q_MX02 U7812 ( .S(n2141), .A0(n1937), .A1(n1938), .Z(ofifoDataN[102]));
Q_AN02 U7813 ( .A0(n6720), .A1(shiftedXdata[103]), .Z(n1936));
Q_MX03 U7814 ( .S0(n2144), .S1(n2402), .A0(ofifoData[103]), .A1(ofifoData[359]), .A2(ofifoData[615]), .Z(n2298));
Q_MX02 U7815 ( .S(n2141), .A0(n1935), .A1(n1936), .Z(ofifoDataN[103]));
Q_AN02 U7816 ( .A0(n6720), .A1(shiftedXdata[104]), .Z(n1934));
Q_MX03 U7817 ( .S0(n2144), .S1(n2402), .A0(ofifoData[104]), .A1(ofifoData[360]), .A2(ofifoData[616]), .Z(n2297));
Q_MX02 U7818 ( .S(n2141), .A0(n1933), .A1(n1934), .Z(ofifoDataN[104]));
Q_AN02 U7819 ( .A0(n6720), .A1(shiftedXdata[105]), .Z(n1932));
Q_MX03 U7820 ( .S0(n2144), .S1(n2402), .A0(ofifoData[105]), .A1(ofifoData[361]), .A2(ofifoData[617]), .Z(n2296));
Q_MX02 U7821 ( .S(n2141), .A0(n1931), .A1(n1932), .Z(ofifoDataN[105]));
Q_AN02 U7822 ( .A0(n6720), .A1(shiftedXdata[106]), .Z(n1930));
Q_MX03 U7823 ( .S0(n2144), .S1(n2402), .A0(ofifoData[106]), .A1(ofifoData[362]), .A2(ofifoData[618]), .Z(n2295));
Q_MX02 U7824 ( .S(n2141), .A0(n1929), .A1(n1930), .Z(ofifoDataN[106]));
Q_AN02 U7825 ( .A0(n6720), .A1(shiftedXdata[107]), .Z(n1928));
Q_MX03 U7826 ( .S0(n2144), .S1(n2402), .A0(ofifoData[107]), .A1(ofifoData[363]), .A2(ofifoData[619]), .Z(n2294));
Q_MX02 U7827 ( .S(n2141), .A0(n1927), .A1(n1928), .Z(ofifoDataN[107]));
Q_AN02 U7828 ( .A0(n6720), .A1(shiftedXdata[108]), .Z(n1926));
Q_MX03 U7829 ( .S0(n2144), .S1(n2402), .A0(ofifoData[108]), .A1(ofifoData[364]), .A2(ofifoData[620]), .Z(n2293));
Q_MX02 U7830 ( .S(n2141), .A0(n1925), .A1(n1926), .Z(ofifoDataN[108]));
Q_AN02 U7831 ( .A0(n6720), .A1(shiftedXdata[109]), .Z(n1924));
Q_MX03 U7832 ( .S0(n2144), .S1(n2402), .A0(ofifoData[109]), .A1(ofifoData[365]), .A2(ofifoData[621]), .Z(n2292));
Q_MX02 U7833 ( .S(n2141), .A0(n1923), .A1(n1924), .Z(ofifoDataN[109]));
Q_AN02 U7834 ( .A0(n6720), .A1(shiftedXdata[110]), .Z(n1922));
Q_MX03 U7835 ( .S0(n2144), .S1(n2402), .A0(ofifoData[110]), .A1(ofifoData[366]), .A2(ofifoData[622]), .Z(n2291));
Q_MX02 U7836 ( .S(n2141), .A0(n1921), .A1(n1922), .Z(ofifoDataN[110]));
Q_AN02 U7837 ( .A0(n6720), .A1(shiftedXdata[111]), .Z(n1920));
Q_MX03 U7838 ( .S0(n2144), .S1(n2402), .A0(ofifoData[111]), .A1(ofifoData[367]), .A2(ofifoData[623]), .Z(n2290));
Q_MX02 U7839 ( .S(n2141), .A0(n1919), .A1(n1920), .Z(ofifoDataN[111]));
Q_AN02 U7840 ( .A0(n6720), .A1(shiftedXdata[112]), .Z(n1918));
Q_MX03 U7841 ( .S0(n2144), .S1(n2402), .A0(ofifoData[112]), .A1(ofifoData[368]), .A2(ofifoData[624]), .Z(n2289));
Q_MX02 U7842 ( .S(n2141), .A0(n1917), .A1(n1918), .Z(ofifoDataN[112]));
Q_AN02 U7843 ( .A0(n6720), .A1(shiftedXdata[113]), .Z(n1916));
Q_MX03 U7844 ( .S0(n2144), .S1(n2402), .A0(ofifoData[113]), .A1(ofifoData[369]), .A2(ofifoData[625]), .Z(n2288));
Q_MX02 U7845 ( .S(n2141), .A0(n1915), .A1(n1916), .Z(ofifoDataN[113]));
Q_AN02 U7846 ( .A0(n6720), .A1(shiftedXdata[114]), .Z(n1914));
Q_MX03 U7847 ( .S0(n2144), .S1(n2402), .A0(ofifoData[114]), .A1(ofifoData[370]), .A2(ofifoData[626]), .Z(n2287));
Q_MX02 U7848 ( .S(n2141), .A0(n1913), .A1(n1914), .Z(ofifoDataN[114]));
Q_AN02 U7849 ( .A0(n6720), .A1(shiftedXdata[115]), .Z(n1912));
Q_MX03 U7850 ( .S0(n2144), .S1(n2402), .A0(ofifoData[115]), .A1(ofifoData[371]), .A2(ofifoData[627]), .Z(n2286));
Q_MX02 U7851 ( .S(n2141), .A0(n1911), .A1(n1912), .Z(ofifoDataN[115]));
Q_AN02 U7852 ( .A0(n6720), .A1(shiftedXdata[116]), .Z(n1910));
Q_MX03 U7853 ( .S0(n2144), .S1(n2402), .A0(ofifoData[116]), .A1(ofifoData[372]), .A2(ofifoData[628]), .Z(n2285));
Q_MX02 U7854 ( .S(n2141), .A0(n1909), .A1(n1910), .Z(ofifoDataN[116]));
Q_AN02 U7855 ( .A0(n6720), .A1(shiftedXdata[117]), .Z(n1908));
Q_MX03 U7856 ( .S0(n2144), .S1(n2402), .A0(ofifoData[117]), .A1(ofifoData[373]), .A2(ofifoData[629]), .Z(n2284));
Q_MX02 U7857 ( .S(n2141), .A0(n1907), .A1(n1908), .Z(ofifoDataN[117]));
Q_AN02 U7858 ( .A0(n6720), .A1(shiftedXdata[118]), .Z(n1906));
Q_MX03 U7859 ( .S0(n2144), .S1(n2402), .A0(ofifoData[118]), .A1(ofifoData[374]), .A2(ofifoData[630]), .Z(n2283));
Q_MX02 U7860 ( .S(n2141), .A0(n1905), .A1(n1906), .Z(ofifoDataN[118]));
Q_AN02 U7861 ( .A0(n6720), .A1(shiftedXdata[119]), .Z(n1904));
Q_MX03 U7862 ( .S0(n2144), .S1(n2402), .A0(ofifoData[119]), .A1(ofifoData[375]), .A2(ofifoData[631]), .Z(n2282));
Q_MX02 U7863 ( .S(n2141), .A0(n1903), .A1(n1904), .Z(ofifoDataN[119]));
Q_AN02 U7864 ( .A0(n6720), .A1(shiftedXdata[120]), .Z(n1902));
Q_MX03 U7865 ( .S0(n2144), .S1(n2402), .A0(ofifoData[120]), .A1(ofifoData[376]), .A2(ofifoData[632]), .Z(n2281));
Q_MX02 U7866 ( .S(n2141), .A0(n1901), .A1(n1902), .Z(ofifoDataN[120]));
Q_AN02 U7867 ( .A0(n6720), .A1(shiftedXdata[121]), .Z(n1900));
Q_MX03 U7868 ( .S0(n2144), .S1(n2402), .A0(ofifoData[121]), .A1(ofifoData[377]), .A2(ofifoData[633]), .Z(n2280));
Q_MX02 U7869 ( .S(n2141), .A0(n1899), .A1(n1900), .Z(ofifoDataN[121]));
Q_AN02 U7870 ( .A0(n6720), .A1(shiftedXdata[122]), .Z(n1898));
Q_MX03 U7871 ( .S0(n2144), .S1(n2402), .A0(ofifoData[122]), .A1(ofifoData[378]), .A2(ofifoData[634]), .Z(n2279));
Q_MX02 U7872 ( .S(n2141), .A0(n1897), .A1(n1898), .Z(ofifoDataN[122]));
Q_AN02 U7873 ( .A0(n6720), .A1(shiftedXdata[123]), .Z(n1896));
Q_MX03 U7874 ( .S0(n2144), .S1(n2402), .A0(ofifoData[123]), .A1(ofifoData[379]), .A2(ofifoData[635]), .Z(n2278));
Q_MX02 U7875 ( .S(n2141), .A0(n1895), .A1(n1896), .Z(ofifoDataN[123]));
Q_AN02 U7876 ( .A0(n6720), .A1(shiftedXdata[124]), .Z(n1894));
Q_MX03 U7877 ( .S0(n2144), .S1(n2402), .A0(ofifoData[124]), .A1(ofifoData[380]), .A2(ofifoData[636]), .Z(n2277));
Q_MX02 U7878 ( .S(n2141), .A0(n1893), .A1(n1894), .Z(ofifoDataN[124]));
Q_AN02 U7879 ( .A0(n6720), .A1(shiftedXdata[125]), .Z(n1892));
Q_MX03 U7880 ( .S0(n2144), .S1(n2402), .A0(ofifoData[125]), .A1(ofifoData[381]), .A2(ofifoData[637]), .Z(n2276));
Q_MX02 U7881 ( .S(n2141), .A0(n1891), .A1(n1892), .Z(ofifoDataN[125]));
Q_AN02 U7882 ( .A0(n6720), .A1(shiftedXdata[126]), .Z(n1890));
Q_MX03 U7883 ( .S0(n2144), .S1(n2402), .A0(ofifoData[126]), .A1(ofifoData[382]), .A2(ofifoData[638]), .Z(n2275));
Q_MX02 U7884 ( .S(n2141), .A0(n1889), .A1(n1890), .Z(ofifoDataN[126]));
Q_AN02 U7885 ( .A0(n6720), .A1(shiftedXdata[127]), .Z(n1888));
Q_MX03 U7886 ( .S0(n2144), .S1(n2402), .A0(ofifoData[127]), .A1(ofifoData[383]), .A2(ofifoData[639]), .Z(n2274));
Q_MX02 U7887 ( .S(n2141), .A0(n1887), .A1(n1888), .Z(ofifoDataN[127]));
Q_AN02 U7888 ( .A0(n6720), .A1(shiftedXdata[128]), .Z(n1886));
Q_MX03 U7889 ( .S0(n2144), .S1(n2402), .A0(ofifoData[128]), .A1(ofifoData[384]), .A2(ofifoData[640]), .Z(n2273));
Q_MX02 U7890 ( .S(n2141), .A0(n1885), .A1(n1886), .Z(ofifoDataN[128]));
Q_AN02 U7891 ( .A0(n6720), .A1(shiftedXdata[129]), .Z(n1884));
Q_MX03 U7892 ( .S0(n2144), .S1(n2402), .A0(ofifoData[129]), .A1(ofifoData[385]), .A2(ofifoData[641]), .Z(n2272));
Q_MX02 U7893 ( .S(n2141), .A0(n1883), .A1(n1884), .Z(ofifoDataN[129]));
Q_AN02 U7894 ( .A0(n6720), .A1(shiftedXdata[130]), .Z(n1882));
Q_MX03 U7895 ( .S0(n2144), .S1(n2402), .A0(ofifoData[130]), .A1(ofifoData[386]), .A2(ofifoData[642]), .Z(n2271));
Q_MX02 U7896 ( .S(n2141), .A0(n1881), .A1(n1882), .Z(ofifoDataN[130]));
Q_AN02 U7897 ( .A0(n6720), .A1(shiftedXdata[131]), .Z(n1880));
Q_MX03 U7898 ( .S0(n2144), .S1(n2402), .A0(ofifoData[131]), .A1(ofifoData[387]), .A2(ofifoData[643]), .Z(n2270));
Q_MX02 U7899 ( .S(n2141), .A0(n1879), .A1(n1880), .Z(ofifoDataN[131]));
Q_AN02 U7900 ( .A0(n6720), .A1(shiftedXdata[132]), .Z(n1878));
Q_MX03 U7901 ( .S0(n2144), .S1(n2402), .A0(ofifoData[132]), .A1(ofifoData[388]), .A2(ofifoData[644]), .Z(n2269));
Q_MX02 U7902 ( .S(n2141), .A0(n1877), .A1(n1878), .Z(ofifoDataN[132]));
Q_AN02 U7903 ( .A0(n6720), .A1(shiftedXdata[133]), .Z(n1876));
Q_MX03 U7904 ( .S0(n2144), .S1(n2402), .A0(ofifoData[133]), .A1(ofifoData[389]), .A2(ofifoData[645]), .Z(n2268));
Q_MX02 U7905 ( .S(n2141), .A0(n1875), .A1(n1876), .Z(ofifoDataN[133]));
Q_AN02 U7906 ( .A0(n6720), .A1(shiftedXdata[134]), .Z(n1874));
Q_MX03 U7907 ( .S0(n2144), .S1(n2402), .A0(ofifoData[134]), .A1(ofifoData[390]), .A2(ofifoData[646]), .Z(n2267));
Q_MX02 U7908 ( .S(n2141), .A0(n1873), .A1(n1874), .Z(ofifoDataN[134]));
Q_AN02 U7909 ( .A0(n6720), .A1(shiftedXdata[135]), .Z(n1872));
Q_MX03 U7910 ( .S0(n2144), .S1(n2402), .A0(ofifoData[135]), .A1(ofifoData[391]), .A2(ofifoData[647]), .Z(n2266));
Q_MX02 U7911 ( .S(n2141), .A0(n1871), .A1(n1872), .Z(ofifoDataN[135]));
Q_AN02 U7912 ( .A0(n6720), .A1(shiftedXdata[136]), .Z(n1870));
Q_MX03 U7913 ( .S0(n2144), .S1(n2402), .A0(ofifoData[136]), .A1(ofifoData[392]), .A2(ofifoData[648]), .Z(n2265));
Q_MX02 U7914 ( .S(n2141), .A0(n1869), .A1(n1870), .Z(ofifoDataN[136]));
Q_AN02 U7915 ( .A0(n6720), .A1(shiftedXdata[137]), .Z(n1868));
Q_MX03 U7916 ( .S0(n2144), .S1(n2402), .A0(ofifoData[137]), .A1(ofifoData[393]), .A2(ofifoData[649]), .Z(n2264));
Q_MX02 U7917 ( .S(n2141), .A0(n1867), .A1(n1868), .Z(ofifoDataN[137]));
Q_AN02 U7918 ( .A0(n6720), .A1(shiftedXdata[138]), .Z(n1866));
Q_MX03 U7919 ( .S0(n2144), .S1(n2402), .A0(ofifoData[138]), .A1(ofifoData[394]), .A2(ofifoData[650]), .Z(n2263));
Q_MX02 U7920 ( .S(n2141), .A0(n1865), .A1(n1866), .Z(ofifoDataN[138]));
Q_AN02 U7921 ( .A0(n6720), .A1(shiftedXdata[139]), .Z(n1864));
Q_MX03 U7922 ( .S0(n2144), .S1(n2402), .A0(ofifoData[139]), .A1(ofifoData[395]), .A2(ofifoData[651]), .Z(n2262));
Q_MX02 U7923 ( .S(n2141), .A0(n1863), .A1(n1864), .Z(ofifoDataN[139]));
Q_AN02 U7924 ( .A0(n6720), .A1(shiftedXdata[140]), .Z(n1862));
Q_MX03 U7925 ( .S0(n2144), .S1(n2402), .A0(ofifoData[140]), .A1(ofifoData[396]), .A2(ofifoData[652]), .Z(n2261));
Q_MX02 U7926 ( .S(n2141), .A0(n1861), .A1(n1862), .Z(ofifoDataN[140]));
Q_AN02 U7927 ( .A0(n6720), .A1(shiftedXdata[141]), .Z(n1860));
Q_MX03 U7928 ( .S0(n2144), .S1(n2402), .A0(ofifoData[141]), .A1(ofifoData[397]), .A2(ofifoData[653]), .Z(n2260));
Q_MX02 U7929 ( .S(n2141), .A0(n1859), .A1(n1860), .Z(ofifoDataN[141]));
Q_AN02 U7930 ( .A0(n6720), .A1(shiftedXdata[142]), .Z(n1858));
Q_MX03 U7931 ( .S0(n2144), .S1(n2402), .A0(ofifoData[142]), .A1(ofifoData[398]), .A2(ofifoData[654]), .Z(n2259));
Q_MX02 U7932 ( .S(n2141), .A0(n1857), .A1(n1858), .Z(ofifoDataN[142]));
Q_AN02 U7933 ( .A0(n6720), .A1(shiftedXdata[143]), .Z(n1856));
Q_MX03 U7934 ( .S0(n2144), .S1(n2402), .A0(ofifoData[143]), .A1(ofifoData[399]), .A2(ofifoData[655]), .Z(n2258));
Q_MX02 U7935 ( .S(n2141), .A0(n1855), .A1(n1856), .Z(ofifoDataN[143]));
Q_AN02 U7936 ( .A0(n6720), .A1(shiftedXdata[144]), .Z(n1854));
Q_MX03 U7937 ( .S0(n2144), .S1(n2402), .A0(ofifoData[144]), .A1(ofifoData[400]), .A2(ofifoData[656]), .Z(n2257));
Q_MX02 U7938 ( .S(n2141), .A0(n1853), .A1(n1854), .Z(ofifoDataN[144]));
Q_AN02 U7939 ( .A0(n6720), .A1(shiftedXdata[145]), .Z(n1852));
Q_MX03 U7940 ( .S0(n2144), .S1(n2402), .A0(ofifoData[145]), .A1(ofifoData[401]), .A2(ofifoData[657]), .Z(n2256));
Q_MX02 U7941 ( .S(n2141), .A0(n1851), .A1(n1852), .Z(ofifoDataN[145]));
Q_AN02 U7942 ( .A0(n6720), .A1(shiftedXdata[146]), .Z(n1850));
Q_MX03 U7943 ( .S0(n2144), .S1(n2402), .A0(ofifoData[146]), .A1(ofifoData[402]), .A2(ofifoData[658]), .Z(n2255));
Q_MX02 U7944 ( .S(n2141), .A0(n1849), .A1(n1850), .Z(ofifoDataN[146]));
Q_AN02 U7945 ( .A0(n6720), .A1(shiftedXdata[147]), .Z(n1848));
Q_MX03 U7946 ( .S0(n2144), .S1(n2402), .A0(ofifoData[147]), .A1(ofifoData[403]), .A2(ofifoData[659]), .Z(n2254));
Q_MX02 U7947 ( .S(n2141), .A0(n1847), .A1(n1848), .Z(ofifoDataN[147]));
Q_AN02 U7948 ( .A0(n6720), .A1(shiftedXdata[148]), .Z(n1846));
Q_MX03 U7949 ( .S0(n2144), .S1(n2402), .A0(ofifoData[148]), .A1(ofifoData[404]), .A2(ofifoData[660]), .Z(n2253));
Q_MX02 U7950 ( .S(n2141), .A0(n1845), .A1(n1846), .Z(ofifoDataN[148]));
Q_AN02 U7951 ( .A0(n6720), .A1(shiftedXdata[149]), .Z(n1844));
Q_MX03 U7952 ( .S0(n2144), .S1(n2402), .A0(ofifoData[149]), .A1(ofifoData[405]), .A2(ofifoData[661]), .Z(n2252));
Q_MX02 U7953 ( .S(n2141), .A0(n1843), .A1(n1844), .Z(ofifoDataN[149]));
Q_AN02 U7954 ( .A0(n6720), .A1(shiftedXdata[150]), .Z(n1842));
Q_MX03 U7955 ( .S0(n2144), .S1(n2402), .A0(ofifoData[150]), .A1(ofifoData[406]), .A2(ofifoData[662]), .Z(n2251));
Q_MX02 U7956 ( .S(n2141), .A0(n1841), .A1(n1842), .Z(ofifoDataN[150]));
Q_AN02 U7957 ( .A0(n6720), .A1(shiftedXdata[151]), .Z(n1840));
Q_MX03 U7958 ( .S0(n2144), .S1(n2402), .A0(ofifoData[151]), .A1(ofifoData[407]), .A2(ofifoData[663]), .Z(n2250));
Q_MX02 U7959 ( .S(n2141), .A0(n1839), .A1(n1840), .Z(ofifoDataN[151]));
Q_AN02 U7960 ( .A0(n6720), .A1(shiftedXdata[152]), .Z(n1838));
Q_MX03 U7961 ( .S0(n2144), .S1(n2402), .A0(ofifoData[152]), .A1(ofifoData[408]), .A2(ofifoData[664]), .Z(n2249));
Q_MX02 U7962 ( .S(n2141), .A0(n1837), .A1(n1838), .Z(ofifoDataN[152]));
Q_AN02 U7963 ( .A0(n6720), .A1(shiftedXdata[153]), .Z(n1836));
Q_MX03 U7964 ( .S0(n2144), .S1(n2402), .A0(ofifoData[153]), .A1(ofifoData[409]), .A2(ofifoData[665]), .Z(n2248));
Q_MX02 U7965 ( .S(n2141), .A0(n1835), .A1(n1836), .Z(ofifoDataN[153]));
Q_AN02 U7966 ( .A0(n6720), .A1(shiftedXdata[154]), .Z(n1834));
Q_MX03 U7967 ( .S0(n2144), .S1(n2402), .A0(ofifoData[154]), .A1(ofifoData[410]), .A2(ofifoData[666]), .Z(n2247));
Q_MX02 U7968 ( .S(n2141), .A0(n1833), .A1(n1834), .Z(ofifoDataN[154]));
Q_AN02 U7969 ( .A0(n6720), .A1(shiftedXdata[155]), .Z(n1832));
Q_MX03 U7970 ( .S0(n2144), .S1(n2402), .A0(ofifoData[155]), .A1(ofifoData[411]), .A2(ofifoData[667]), .Z(n2246));
Q_MX02 U7971 ( .S(n2141), .A0(n1831), .A1(n1832), .Z(ofifoDataN[155]));
Q_AN02 U7972 ( .A0(n6720), .A1(shiftedXdata[156]), .Z(n1830));
Q_MX03 U7973 ( .S0(n2144), .S1(n2402), .A0(ofifoData[156]), .A1(ofifoData[412]), .A2(ofifoData[668]), .Z(n2245));
Q_MX02 U7974 ( .S(n2141), .A0(n1829), .A1(n1830), .Z(ofifoDataN[156]));
Q_AN02 U7975 ( .A0(n6720), .A1(shiftedXdata[157]), .Z(n1828));
Q_MX03 U7976 ( .S0(n2144), .S1(n2402), .A0(ofifoData[157]), .A1(ofifoData[413]), .A2(ofifoData[669]), .Z(n2244));
Q_MX02 U7977 ( .S(n2141), .A0(n1827), .A1(n1828), .Z(ofifoDataN[157]));
Q_AN02 U7978 ( .A0(n6720), .A1(shiftedXdata[158]), .Z(n1826));
Q_MX03 U7979 ( .S0(n2144), .S1(n2402), .A0(ofifoData[158]), .A1(ofifoData[414]), .A2(ofifoData[670]), .Z(n2243));
Q_MX02 U7980 ( .S(n2141), .A0(n1825), .A1(n1826), .Z(ofifoDataN[158]));
Q_AN02 U7981 ( .A0(n6720), .A1(shiftedXdata[159]), .Z(n1824));
Q_MX03 U7982 ( .S0(n2144), .S1(n2402), .A0(ofifoData[159]), .A1(ofifoData[415]), .A2(ofifoData[671]), .Z(n2242));
Q_MX02 U7983 ( .S(n2141), .A0(n1823), .A1(n1824), .Z(ofifoDataN[159]));
Q_AN02 U7984 ( .A0(n6720), .A1(shiftedXdata[160]), .Z(n1822));
Q_MX03 U7985 ( .S0(n2144), .S1(n2402), .A0(ofifoData[160]), .A1(ofifoData[416]), .A2(ofifoData[672]), .Z(n2241));
Q_MX02 U7986 ( .S(n2141), .A0(n1821), .A1(n1822), .Z(ofifoDataN[160]));
Q_AN02 U7987 ( .A0(n6720), .A1(shiftedXdata[161]), .Z(n1820));
Q_MX03 U7988 ( .S0(n2144), .S1(n2402), .A0(ofifoData[161]), .A1(ofifoData[417]), .A2(ofifoData[673]), .Z(n2240));
Q_MX02 U7989 ( .S(n2141), .A0(n1819), .A1(n1820), .Z(ofifoDataN[161]));
Q_AN02 U7990 ( .A0(n6720), .A1(shiftedXdata[162]), .Z(n1818));
Q_MX03 U7991 ( .S0(n2144), .S1(n2402), .A0(ofifoData[162]), .A1(ofifoData[418]), .A2(ofifoData[674]), .Z(n2239));
Q_MX02 U7992 ( .S(n2141), .A0(n1817), .A1(n1818), .Z(ofifoDataN[162]));
Q_AN02 U7993 ( .A0(n6720), .A1(shiftedXdata[163]), .Z(n1816));
Q_MX03 U7994 ( .S0(n2144), .S1(n2402), .A0(ofifoData[163]), .A1(ofifoData[419]), .A2(ofifoData[675]), .Z(n2238));
Q_MX02 U7995 ( .S(n2141), .A0(n1815), .A1(n1816), .Z(ofifoDataN[163]));
Q_AN02 U7996 ( .A0(n6720), .A1(shiftedXdata[164]), .Z(n1814));
Q_MX03 U7997 ( .S0(n2144), .S1(n2402), .A0(ofifoData[164]), .A1(ofifoData[420]), .A2(ofifoData[676]), .Z(n2237));
Q_MX02 U7998 ( .S(n2141), .A0(n1813), .A1(n1814), .Z(ofifoDataN[164]));
Q_AN02 U7999 ( .A0(n6720), .A1(shiftedXdata[165]), .Z(n1812));
Q_MX03 U8000 ( .S0(n2144), .S1(n2402), .A0(ofifoData[165]), .A1(ofifoData[421]), .A2(ofifoData[677]), .Z(n2236));
Q_MX02 U8001 ( .S(n2141), .A0(n1811), .A1(n1812), .Z(ofifoDataN[165]));
Q_AN02 U8002 ( .A0(n6720), .A1(shiftedXdata[166]), .Z(n1810));
Q_MX03 U8003 ( .S0(n2144), .S1(n2402), .A0(ofifoData[166]), .A1(ofifoData[422]), .A2(ofifoData[678]), .Z(n2235));
Q_MX02 U8004 ( .S(n2141), .A0(n1809), .A1(n1810), .Z(ofifoDataN[166]));
Q_AN02 U8005 ( .A0(n6720), .A1(shiftedXdata[167]), .Z(n1808));
Q_MX03 U8006 ( .S0(n2144), .S1(n2402), .A0(ofifoData[167]), .A1(ofifoData[423]), .A2(ofifoData[679]), .Z(n2234));
Q_MX02 U8007 ( .S(n2141), .A0(n1807), .A1(n1808), .Z(ofifoDataN[167]));
Q_AN02 U8008 ( .A0(n6720), .A1(shiftedXdata[168]), .Z(n1806));
Q_MX03 U8009 ( .S0(n2144), .S1(n2402), .A0(ofifoData[168]), .A1(ofifoData[424]), .A2(ofifoData[680]), .Z(n2233));
Q_MX02 U8010 ( .S(n2141), .A0(n1805), .A1(n1806), .Z(ofifoDataN[168]));
Q_AN02 U8011 ( .A0(n6720), .A1(shiftedXdata[169]), .Z(n1804));
Q_MX03 U8012 ( .S0(n2144), .S1(n2402), .A0(ofifoData[169]), .A1(ofifoData[425]), .A2(ofifoData[681]), .Z(n2232));
Q_MX02 U8013 ( .S(n2141), .A0(n1803), .A1(n1804), .Z(ofifoDataN[169]));
Q_AN02 U8014 ( .A0(n6720), .A1(shiftedXdata[170]), .Z(n1802));
Q_MX03 U8015 ( .S0(n2144), .S1(n2402), .A0(ofifoData[170]), .A1(ofifoData[426]), .A2(ofifoData[682]), .Z(n2231));
Q_MX02 U8016 ( .S(n2141), .A0(n1801), .A1(n1802), .Z(ofifoDataN[170]));
Q_AN02 U8017 ( .A0(n6720), .A1(shiftedXdata[171]), .Z(n1800));
Q_MX03 U8018 ( .S0(n2144), .S1(n2402), .A0(ofifoData[171]), .A1(ofifoData[427]), .A2(ofifoData[683]), .Z(n2230));
Q_MX02 U8019 ( .S(n2141), .A0(n1799), .A1(n1800), .Z(ofifoDataN[171]));
Q_AN02 U8020 ( .A0(n6720), .A1(shiftedXdata[172]), .Z(n1798));
Q_MX03 U8021 ( .S0(n2144), .S1(n2402), .A0(ofifoData[172]), .A1(ofifoData[428]), .A2(ofifoData[684]), .Z(n2229));
Q_MX02 U8022 ( .S(n2141), .A0(n1797), .A1(n1798), .Z(ofifoDataN[172]));
Q_AN02 U8023 ( .A0(n6720), .A1(shiftedXdata[173]), .Z(n1796));
Q_MX03 U8024 ( .S0(n2144), .S1(n2402), .A0(ofifoData[173]), .A1(ofifoData[429]), .A2(ofifoData[685]), .Z(n2228));
Q_MX02 U8025 ( .S(n2141), .A0(n1795), .A1(n1796), .Z(ofifoDataN[173]));
Q_AN02 U8026 ( .A0(n6720), .A1(shiftedXdata[174]), .Z(n1794));
Q_MX03 U8027 ( .S0(n2144), .S1(n2402), .A0(ofifoData[174]), .A1(ofifoData[430]), .A2(ofifoData[686]), .Z(n2227));
Q_MX02 U8028 ( .S(n2141), .A0(n1793), .A1(n1794), .Z(ofifoDataN[174]));
Q_AN02 U8029 ( .A0(n6720), .A1(shiftedXdata[175]), .Z(n1792));
Q_MX03 U8030 ( .S0(n2144), .S1(n2402), .A0(ofifoData[175]), .A1(ofifoData[431]), .A2(ofifoData[687]), .Z(n2226));
Q_MX02 U8031 ( .S(n2141), .A0(n1791), .A1(n1792), .Z(ofifoDataN[175]));
Q_AN02 U8032 ( .A0(n6720), .A1(shiftedXdata[176]), .Z(n1790));
Q_MX03 U8033 ( .S0(n2144), .S1(n2402), .A0(ofifoData[176]), .A1(ofifoData[432]), .A2(ofifoData[688]), .Z(n2225));
Q_MX02 U8034 ( .S(n2141), .A0(n1789), .A1(n1790), .Z(ofifoDataN[176]));
Q_AN02 U8035 ( .A0(n6720), .A1(shiftedXdata[177]), .Z(n1788));
Q_MX03 U8036 ( .S0(n2144), .S1(n2402), .A0(ofifoData[177]), .A1(ofifoData[433]), .A2(ofifoData[689]), .Z(n2224));
Q_MX02 U8037 ( .S(n2141), .A0(n1787), .A1(n1788), .Z(ofifoDataN[177]));
Q_AN02 U8038 ( .A0(n6720), .A1(shiftedXdata[178]), .Z(n1786));
Q_MX03 U8039 ( .S0(n2144), .S1(n2402), .A0(ofifoData[178]), .A1(ofifoData[434]), .A2(ofifoData[690]), .Z(n2223));
Q_MX02 U8040 ( .S(n2141), .A0(n1785), .A1(n1786), .Z(ofifoDataN[178]));
Q_AN02 U8041 ( .A0(n6720), .A1(shiftedXdata[179]), .Z(n1784));
Q_MX03 U8042 ( .S0(n2144), .S1(n2402), .A0(ofifoData[179]), .A1(ofifoData[435]), .A2(ofifoData[691]), .Z(n2222));
Q_MX02 U8043 ( .S(n2141), .A0(n1783), .A1(n1784), .Z(ofifoDataN[179]));
Q_AN02 U8044 ( .A0(n6720), .A1(shiftedXdata[180]), .Z(n1782));
Q_MX03 U8045 ( .S0(n2144), .S1(n2402), .A0(ofifoData[180]), .A1(ofifoData[436]), .A2(ofifoData[692]), .Z(n2221));
Q_MX02 U8046 ( .S(n2141), .A0(n1781), .A1(n1782), .Z(ofifoDataN[180]));
Q_AN02 U8047 ( .A0(n6720), .A1(shiftedXdata[181]), .Z(n1780));
Q_MX03 U8048 ( .S0(n2144), .S1(n2402), .A0(ofifoData[181]), .A1(ofifoData[437]), .A2(ofifoData[693]), .Z(n2220));
Q_MX02 U8049 ( .S(n2141), .A0(n1779), .A1(n1780), .Z(ofifoDataN[181]));
Q_AN02 U8050 ( .A0(n6720), .A1(shiftedXdata[182]), .Z(n1778));
Q_MX03 U8051 ( .S0(n2144), .S1(n2402), .A0(ofifoData[182]), .A1(ofifoData[438]), .A2(ofifoData[694]), .Z(n2219));
Q_MX02 U8052 ( .S(n2141), .A0(n1777), .A1(n1778), .Z(ofifoDataN[182]));
Q_AN02 U8053 ( .A0(n6720), .A1(shiftedXdata[183]), .Z(n1776));
Q_MX03 U8054 ( .S0(n2144), .S1(n2402), .A0(ofifoData[183]), .A1(ofifoData[439]), .A2(ofifoData[695]), .Z(n2218));
Q_MX02 U8055 ( .S(n2141), .A0(n1775), .A1(n1776), .Z(ofifoDataN[183]));
Q_AN02 U8056 ( .A0(n6720), .A1(shiftedXdata[184]), .Z(n1774));
Q_MX03 U8057 ( .S0(n2144), .S1(n2402), .A0(ofifoData[184]), .A1(ofifoData[440]), .A2(ofifoData[696]), .Z(n2217));
Q_MX02 U8058 ( .S(n2141), .A0(n1773), .A1(n1774), .Z(ofifoDataN[184]));
Q_AN02 U8059 ( .A0(n6720), .A1(shiftedXdata[185]), .Z(n1772));
Q_MX03 U8060 ( .S0(n2144), .S1(n2402), .A0(ofifoData[185]), .A1(ofifoData[441]), .A2(ofifoData[697]), .Z(n2216));
Q_MX02 U8061 ( .S(n2141), .A0(n1771), .A1(n1772), .Z(ofifoDataN[185]));
Q_AN02 U8062 ( .A0(n6720), .A1(shiftedXdata[186]), .Z(n1770));
Q_MX03 U8063 ( .S0(n2144), .S1(n2402), .A0(ofifoData[186]), .A1(ofifoData[442]), .A2(ofifoData[698]), .Z(n2215));
Q_MX02 U8064 ( .S(n2141), .A0(n1769), .A1(n1770), .Z(ofifoDataN[186]));
Q_AN02 U8065 ( .A0(n6720), .A1(shiftedXdata[187]), .Z(n1768));
Q_MX03 U8066 ( .S0(n2144), .S1(n2402), .A0(ofifoData[187]), .A1(ofifoData[443]), .A2(ofifoData[699]), .Z(n2214));
Q_MX02 U8067 ( .S(n2141), .A0(n1767), .A1(n1768), .Z(ofifoDataN[187]));
Q_AN02 U8068 ( .A0(n6720), .A1(shiftedXdata[188]), .Z(n1766));
Q_MX03 U8069 ( .S0(n2144), .S1(n2402), .A0(ofifoData[188]), .A1(ofifoData[444]), .A2(ofifoData[700]), .Z(n2213));
Q_MX02 U8070 ( .S(n2141), .A0(n1765), .A1(n1766), .Z(ofifoDataN[188]));
Q_AN02 U8071 ( .A0(n6720), .A1(shiftedXdata[189]), .Z(n1764));
Q_MX03 U8072 ( .S0(n2144), .S1(n2402), .A0(ofifoData[189]), .A1(ofifoData[445]), .A2(ofifoData[701]), .Z(n2212));
Q_MX02 U8073 ( .S(n2141), .A0(n1763), .A1(n1764), .Z(ofifoDataN[189]));
Q_AN02 U8074 ( .A0(n6720), .A1(shiftedXdata[190]), .Z(n1762));
Q_MX03 U8075 ( .S0(n2144), .S1(n2402), .A0(ofifoData[190]), .A1(ofifoData[446]), .A2(ofifoData[702]), .Z(n2211));
Q_MX02 U8076 ( .S(n2141), .A0(n1761), .A1(n1762), .Z(ofifoDataN[190]));
Q_AN02 U8077 ( .A0(n6720), .A1(shiftedXdata[191]), .Z(n1760));
Q_MX03 U8078 ( .S0(n2144), .S1(n2402), .A0(ofifoData[191]), .A1(ofifoData[447]), .A2(ofifoData[703]), .Z(n2210));
Q_MX02 U8079 ( .S(n2141), .A0(n1759), .A1(n1760), .Z(ofifoDataN[191]));
Q_AN02 U8080 ( .A0(n6720), .A1(shiftedXdata[192]), .Z(n1758));
Q_MX03 U8081 ( .S0(n2144), .S1(n2402), .A0(ofifoData[192]), .A1(ofifoData[448]), .A2(ofifoData[704]), .Z(n2209));
Q_MX02 U8082 ( .S(n2141), .A0(n1757), .A1(n1758), .Z(ofifoDataN[192]));
Q_AN02 U8083 ( .A0(n6720), .A1(shiftedXdata[193]), .Z(n1756));
Q_MX03 U8084 ( .S0(n2144), .S1(n2402), .A0(ofifoData[193]), .A1(ofifoData[449]), .A2(ofifoData[705]), .Z(n2208));
Q_MX02 U8085 ( .S(n2141), .A0(n1755), .A1(n1756), .Z(ofifoDataN[193]));
Q_AN02 U8086 ( .A0(n6720), .A1(shiftedXdata[194]), .Z(n1754));
Q_MX03 U8087 ( .S0(n2144), .S1(n2402), .A0(ofifoData[194]), .A1(ofifoData[450]), .A2(ofifoData[706]), .Z(n2207));
Q_MX02 U8088 ( .S(n2141), .A0(n1753), .A1(n1754), .Z(ofifoDataN[194]));
Q_AN02 U8089 ( .A0(n6720), .A1(shiftedXdata[195]), .Z(n1752));
Q_MX03 U8090 ( .S0(n2144), .S1(n2402), .A0(ofifoData[195]), .A1(ofifoData[451]), .A2(ofifoData[707]), .Z(n2206));
Q_MX02 U8091 ( .S(n2141), .A0(n1751), .A1(n1752), .Z(ofifoDataN[195]));
Q_AN02 U8092 ( .A0(n6720), .A1(shiftedXdata[196]), .Z(n1750));
Q_MX03 U8093 ( .S0(n2144), .S1(n2402), .A0(ofifoData[196]), .A1(ofifoData[452]), .A2(ofifoData[708]), .Z(n2205));
Q_MX02 U8094 ( .S(n2141), .A0(n1749), .A1(n1750), .Z(ofifoDataN[196]));
Q_AN02 U8095 ( .A0(n6720), .A1(shiftedXdata[197]), .Z(n1748));
Q_MX03 U8096 ( .S0(n2144), .S1(n2402), .A0(ofifoData[197]), .A1(ofifoData[453]), .A2(ofifoData[709]), .Z(n2204));
Q_MX02 U8097 ( .S(n2141), .A0(n1747), .A1(n1748), .Z(ofifoDataN[197]));
Q_AN02 U8098 ( .A0(n6720), .A1(shiftedXdata[198]), .Z(n1746));
Q_MX03 U8099 ( .S0(n2144), .S1(n2402), .A0(ofifoData[198]), .A1(ofifoData[454]), .A2(ofifoData[710]), .Z(n2203));
Q_MX02 U8100 ( .S(n2141), .A0(n1745), .A1(n1746), .Z(ofifoDataN[198]));
Q_AN02 U8101 ( .A0(n6720), .A1(shiftedXdata[199]), .Z(n1744));
Q_MX03 U8102 ( .S0(n2144), .S1(n2402), .A0(ofifoData[199]), .A1(ofifoData[455]), .A2(ofifoData[711]), .Z(n2202));
Q_MX02 U8103 ( .S(n2141), .A0(n1743), .A1(n1744), .Z(ofifoDataN[199]));
Q_AN02 U8104 ( .A0(n6720), .A1(shiftedXdata[200]), .Z(n1742));
Q_MX03 U8105 ( .S0(n2144), .S1(n2402), .A0(ofifoData[200]), .A1(ofifoData[456]), .A2(ofifoData[712]), .Z(n2201));
Q_MX02 U8106 ( .S(n2141), .A0(n1741), .A1(n1742), .Z(ofifoDataN[200]));
Q_AN02 U8107 ( .A0(n6720), .A1(shiftedXdata[201]), .Z(n1740));
Q_MX03 U8108 ( .S0(n2144), .S1(n2402), .A0(ofifoData[201]), .A1(ofifoData[457]), .A2(ofifoData[713]), .Z(n2200));
Q_MX02 U8109 ( .S(n2141), .A0(n1739), .A1(n1740), .Z(ofifoDataN[201]));
Q_AN02 U8110 ( .A0(n6720), .A1(shiftedXdata[202]), .Z(n1738));
Q_MX03 U8111 ( .S0(n2144), .S1(n2402), .A0(ofifoData[202]), .A1(ofifoData[458]), .A2(ofifoData[714]), .Z(n2199));
Q_MX02 U8112 ( .S(n2141), .A0(n1737), .A1(n1738), .Z(ofifoDataN[202]));
Q_AN02 U8113 ( .A0(n6720), .A1(shiftedXdata[203]), .Z(n1736));
Q_MX03 U8114 ( .S0(n2144), .S1(n2402), .A0(ofifoData[203]), .A1(ofifoData[459]), .A2(ofifoData[715]), .Z(n2198));
Q_MX02 U8115 ( .S(n2141), .A0(n1735), .A1(n1736), .Z(ofifoDataN[203]));
Q_AN02 U8116 ( .A0(n6720), .A1(shiftedXdata[204]), .Z(n1734));
Q_MX03 U8117 ( .S0(n2144), .S1(n2402), .A0(ofifoData[204]), .A1(ofifoData[460]), .A2(ofifoData[716]), .Z(n2197));
Q_MX02 U8118 ( .S(n2141), .A0(n1733), .A1(n1734), .Z(ofifoDataN[204]));
Q_AN02 U8119 ( .A0(n6720), .A1(shiftedXdata[205]), .Z(n1732));
Q_MX03 U8120 ( .S0(n2144), .S1(n2402), .A0(ofifoData[205]), .A1(ofifoData[461]), .A2(ofifoData[717]), .Z(n2196));
Q_MX02 U8121 ( .S(n2141), .A0(n1731), .A1(n1732), .Z(ofifoDataN[205]));
Q_AN02 U8122 ( .A0(n6720), .A1(shiftedXdata[206]), .Z(n1730));
Q_MX03 U8123 ( .S0(n2144), .S1(n2402), .A0(ofifoData[206]), .A1(ofifoData[462]), .A2(ofifoData[718]), .Z(n2195));
Q_MX02 U8124 ( .S(n2141), .A0(n1729), .A1(n1730), .Z(ofifoDataN[206]));
Q_AN02 U8125 ( .A0(n6720), .A1(shiftedXdata[207]), .Z(n1728));
Q_MX03 U8126 ( .S0(n2144), .S1(n2402), .A0(ofifoData[207]), .A1(ofifoData[463]), .A2(ofifoData[719]), .Z(n2194));
Q_MX02 U8127 ( .S(n2141), .A0(n1727), .A1(n1728), .Z(ofifoDataN[207]));
Q_AN02 U8128 ( .A0(n6720), .A1(shiftedXdata[208]), .Z(n1726));
Q_MX03 U8129 ( .S0(n2144), .S1(n2402), .A0(ofifoData[208]), .A1(ofifoData[464]), .A2(ofifoData[720]), .Z(n2193));
Q_MX02 U8130 ( .S(n2141), .A0(n1725), .A1(n1726), .Z(ofifoDataN[208]));
Q_AN02 U8131 ( .A0(n6720), .A1(shiftedXdata[209]), .Z(n1724));
Q_MX03 U8132 ( .S0(n2144), .S1(n2402), .A0(ofifoData[209]), .A1(ofifoData[465]), .A2(ofifoData[721]), .Z(n2192));
Q_MX02 U8133 ( .S(n2141), .A0(n1723), .A1(n1724), .Z(ofifoDataN[209]));
Q_AN02 U8134 ( .A0(n6720), .A1(shiftedXdata[210]), .Z(n1722));
Q_MX03 U8135 ( .S0(n2144), .S1(n2402), .A0(ofifoData[210]), .A1(ofifoData[466]), .A2(ofifoData[722]), .Z(n2191));
Q_MX02 U8136 ( .S(n2141), .A0(n1721), .A1(n1722), .Z(ofifoDataN[210]));
Q_AN02 U8137 ( .A0(n6720), .A1(shiftedXdata[211]), .Z(n1720));
Q_MX03 U8138 ( .S0(n2144), .S1(n2402), .A0(ofifoData[211]), .A1(ofifoData[467]), .A2(ofifoData[723]), .Z(n2190));
Q_MX02 U8139 ( .S(n2141), .A0(n1719), .A1(n1720), .Z(ofifoDataN[211]));
Q_AN02 U8140 ( .A0(n6720), .A1(shiftedXdata[212]), .Z(n1718));
Q_MX03 U8141 ( .S0(n2144), .S1(n2402), .A0(ofifoData[212]), .A1(ofifoData[468]), .A2(ofifoData[724]), .Z(n2189));
Q_MX02 U8142 ( .S(n2141), .A0(n1717), .A1(n1718), .Z(ofifoDataN[212]));
Q_AN02 U8143 ( .A0(n6720), .A1(shiftedXdata[213]), .Z(n1716));
Q_MX03 U8144 ( .S0(n2144), .S1(n2402), .A0(ofifoData[213]), .A1(ofifoData[469]), .A2(ofifoData[725]), .Z(n2188));
Q_MX02 U8145 ( .S(n2141), .A0(n1715), .A1(n1716), .Z(ofifoDataN[213]));
Q_AN02 U8146 ( .A0(n6720), .A1(shiftedXdata[214]), .Z(n1714));
Q_MX03 U8147 ( .S0(n2144), .S1(n2402), .A0(ofifoData[214]), .A1(ofifoData[470]), .A2(ofifoData[726]), .Z(n2187));
Q_MX02 U8148 ( .S(n2141), .A0(n1713), .A1(n1714), .Z(ofifoDataN[214]));
Q_AN02 U8149 ( .A0(n6720), .A1(shiftedXdata[215]), .Z(n1712));
Q_MX03 U8150 ( .S0(n2144), .S1(n2402), .A0(ofifoData[215]), .A1(ofifoData[471]), .A2(ofifoData[727]), .Z(n2186));
Q_MX02 U8151 ( .S(n2141), .A0(n1711), .A1(n1712), .Z(ofifoDataN[215]));
Q_AN02 U8152 ( .A0(n6720), .A1(shiftedXdata[216]), .Z(n1710));
Q_MX03 U8153 ( .S0(n2144), .S1(n2402), .A0(ofifoData[216]), .A1(ofifoData[472]), .A2(ofifoData[728]), .Z(n2185));
Q_MX02 U8154 ( .S(n2141), .A0(n1709), .A1(n1710), .Z(ofifoDataN[216]));
Q_AN02 U8155 ( .A0(n6720), .A1(shiftedXdata[217]), .Z(n1708));
Q_MX03 U8156 ( .S0(n2144), .S1(n2402), .A0(ofifoData[217]), .A1(ofifoData[473]), .A2(ofifoData[729]), .Z(n2184));
Q_MX02 U8157 ( .S(n2141), .A0(n1707), .A1(n1708), .Z(ofifoDataN[217]));
Q_AN02 U8158 ( .A0(n6720), .A1(shiftedXdata[218]), .Z(n1706));
Q_MX03 U8159 ( .S0(n2144), .S1(n2402), .A0(ofifoData[218]), .A1(ofifoData[474]), .A2(ofifoData[730]), .Z(n2183));
Q_MX02 U8160 ( .S(n2141), .A0(n1705), .A1(n1706), .Z(ofifoDataN[218]));
Q_AN02 U8161 ( .A0(n6720), .A1(shiftedXdata[219]), .Z(n1704));
Q_MX03 U8162 ( .S0(n2144), .S1(n2402), .A0(ofifoData[219]), .A1(ofifoData[475]), .A2(ofifoData[731]), .Z(n2182));
Q_MX02 U8163 ( .S(n2141), .A0(n1703), .A1(n1704), .Z(ofifoDataN[219]));
Q_AN02 U8164 ( .A0(n6720), .A1(shiftedXdata[220]), .Z(n1702));
Q_MX03 U8165 ( .S0(n2144), .S1(n2402), .A0(ofifoData[220]), .A1(ofifoData[476]), .A2(ofifoData[732]), .Z(n2181));
Q_MX02 U8166 ( .S(n2141), .A0(n1701), .A1(n1702), .Z(ofifoDataN[220]));
Q_AN02 U8167 ( .A0(n6720), .A1(shiftedXdata[221]), .Z(n1700));
Q_MX03 U8168 ( .S0(n2144), .S1(n2402), .A0(ofifoData[221]), .A1(ofifoData[477]), .A2(ofifoData[733]), .Z(n2180));
Q_MX02 U8169 ( .S(n2141), .A0(n1699), .A1(n1700), .Z(ofifoDataN[221]));
Q_AN02 U8170 ( .A0(n6720), .A1(shiftedXdata[222]), .Z(n1698));
Q_MX03 U8171 ( .S0(n2144), .S1(n2402), .A0(ofifoData[222]), .A1(ofifoData[478]), .A2(ofifoData[734]), .Z(n2179));
Q_MX02 U8172 ( .S(n2141), .A0(n1697), .A1(n1698), .Z(ofifoDataN[222]));
Q_AN02 U8173 ( .A0(n6720), .A1(shiftedXdata[223]), .Z(n1696));
Q_MX03 U8174 ( .S0(n2144), .S1(n2402), .A0(ofifoData[223]), .A1(ofifoData[479]), .A2(ofifoData[735]), .Z(n2178));
Q_MX02 U8175 ( .S(n2141), .A0(n1695), .A1(n1696), .Z(ofifoDataN[223]));
Q_AN02 U8176 ( .A0(n6720), .A1(shiftedXdata[224]), .Z(n1694));
Q_MX03 U8177 ( .S0(n2144), .S1(n2402), .A0(ofifoData[224]), .A1(ofifoData[480]), .A2(ofifoData[736]), .Z(n2177));
Q_MX02 U8178 ( .S(n2141), .A0(n1693), .A1(n1694), .Z(ofifoDataN[224]));
Q_AN02 U8179 ( .A0(n6720), .A1(shiftedXdata[225]), .Z(n1692));
Q_MX03 U8180 ( .S0(n2144), .S1(n2402), .A0(ofifoData[225]), .A1(ofifoData[481]), .A2(ofifoData[737]), .Z(n2176));
Q_MX02 U8181 ( .S(n2141), .A0(n1691), .A1(n1692), .Z(ofifoDataN[225]));
Q_AN02 U8182 ( .A0(n6720), .A1(shiftedXdata[226]), .Z(n1690));
Q_MX03 U8183 ( .S0(n2144), .S1(n2402), .A0(ofifoData[226]), .A1(ofifoData[482]), .A2(ofifoData[738]), .Z(n2175));
Q_MX02 U8184 ( .S(n2141), .A0(n1689), .A1(n1690), .Z(ofifoDataN[226]));
Q_AN02 U8185 ( .A0(n6720), .A1(shiftedXdata[227]), .Z(n1688));
Q_MX03 U8186 ( .S0(n2144), .S1(n2402), .A0(ofifoData[227]), .A1(ofifoData[483]), .A2(ofifoData[739]), .Z(n2174));
Q_MX02 U8187 ( .S(n2141), .A0(n1687), .A1(n1688), .Z(ofifoDataN[227]));
Q_AN02 U8188 ( .A0(n6720), .A1(shiftedXdata[228]), .Z(n1686));
Q_MX03 U8189 ( .S0(n2144), .S1(n2402), .A0(ofifoData[228]), .A1(ofifoData[484]), .A2(ofifoData[740]), .Z(n2173));
Q_MX02 U8190 ( .S(n2141), .A0(n1685), .A1(n1686), .Z(ofifoDataN[228]));
Q_AN02 U8191 ( .A0(n6720), .A1(shiftedXdata[229]), .Z(n1684));
Q_MX03 U8192 ( .S0(n2144), .S1(n2402), .A0(ofifoData[229]), .A1(ofifoData[485]), .A2(ofifoData[741]), .Z(n2172));
Q_MX02 U8193 ( .S(n2141), .A0(n1683), .A1(n1684), .Z(ofifoDataN[229]));
Q_AN02 U8194 ( .A0(n6720), .A1(shiftedXdata[230]), .Z(n1682));
Q_MX03 U8195 ( .S0(n2144), .S1(n2402), .A0(ofifoData[230]), .A1(ofifoData[486]), .A2(ofifoData[742]), .Z(n2171));
Q_MX02 U8196 ( .S(n2141), .A0(n1681), .A1(n1682), .Z(ofifoDataN[230]));
Q_AN02 U8197 ( .A0(n6720), .A1(shiftedXdata[231]), .Z(n1680));
Q_MX03 U8198 ( .S0(n2144), .S1(n2402), .A0(ofifoData[231]), .A1(ofifoData[487]), .A2(ofifoData[743]), .Z(n2170));
Q_MX02 U8199 ( .S(n2141), .A0(n1679), .A1(n1680), .Z(ofifoDataN[231]));
Q_AN02 U8200 ( .A0(n6720), .A1(shiftedXdata[232]), .Z(n1678));
Q_MX03 U8201 ( .S0(n2144), .S1(n2402), .A0(ofifoData[232]), .A1(ofifoData[488]), .A2(ofifoData[744]), .Z(n2169));
Q_MX02 U8202 ( .S(n2141), .A0(n1677), .A1(n1678), .Z(ofifoDataN[232]));
Q_AN02 U8203 ( .A0(n6720), .A1(shiftedXdata[233]), .Z(n1676));
Q_MX03 U8204 ( .S0(n2144), .S1(n2402), .A0(ofifoData[233]), .A1(ofifoData[489]), .A2(ofifoData[745]), .Z(n2168));
Q_MX02 U8205 ( .S(n2141), .A0(n1675), .A1(n1676), .Z(ofifoDataN[233]));
Q_AN02 U8206 ( .A0(n6720), .A1(shiftedXdata[234]), .Z(n1674));
Q_MX03 U8207 ( .S0(n2144), .S1(n2402), .A0(ofifoData[234]), .A1(ofifoData[490]), .A2(ofifoData[746]), .Z(n2167));
Q_MX02 U8208 ( .S(n2141), .A0(n1673), .A1(n1674), .Z(ofifoDataN[234]));
Q_AN02 U8209 ( .A0(n6720), .A1(shiftedXdata[235]), .Z(n1672));
Q_MX03 U8210 ( .S0(n2144), .S1(n2402), .A0(ofifoData[235]), .A1(ofifoData[491]), .A2(ofifoData[747]), .Z(n2166));
Q_MX02 U8211 ( .S(n2141), .A0(n1671), .A1(n1672), .Z(ofifoDataN[235]));
Q_AN02 U8212 ( .A0(n6720), .A1(shiftedXdata[236]), .Z(n1670));
Q_MX03 U8213 ( .S0(n2144), .S1(n2402), .A0(ofifoData[236]), .A1(ofifoData[492]), .A2(ofifoData[748]), .Z(n2165));
Q_MX02 U8214 ( .S(n2141), .A0(n1669), .A1(n1670), .Z(ofifoDataN[236]));
Q_AN02 U8215 ( .A0(n6720), .A1(shiftedXdata[237]), .Z(n1668));
Q_MX03 U8216 ( .S0(n2144), .S1(n2402), .A0(ofifoData[237]), .A1(ofifoData[493]), .A2(ofifoData[749]), .Z(n2164));
Q_MX02 U8217 ( .S(n2141), .A0(n1667), .A1(n1668), .Z(ofifoDataN[237]));
Q_AN02 U8218 ( .A0(n6720), .A1(shiftedXdata[238]), .Z(n1666));
Q_MX03 U8219 ( .S0(n2144), .S1(n2402), .A0(ofifoData[238]), .A1(ofifoData[494]), .A2(ofifoData[750]), .Z(n2163));
Q_MX02 U8220 ( .S(n2141), .A0(n1665), .A1(n1666), .Z(ofifoDataN[238]));
Q_AN02 U8221 ( .A0(n6720), .A1(shiftedXdata[239]), .Z(n1664));
Q_MX03 U8222 ( .S0(n2144), .S1(n2402), .A0(ofifoData[239]), .A1(ofifoData[495]), .A2(ofifoData[751]), .Z(n2162));
Q_MX02 U8223 ( .S(n2141), .A0(n1663), .A1(n1664), .Z(ofifoDataN[239]));
Q_AN02 U8224 ( .A0(n6720), .A1(shiftedXdata[240]), .Z(n1662));
Q_MX03 U8225 ( .S0(n2144), .S1(n2402), .A0(ofifoData[240]), .A1(ofifoData[496]), .A2(ofifoData[752]), .Z(n2161));
Q_MX02 U8226 ( .S(n2141), .A0(n1661), .A1(n1662), .Z(ofifoDataN[240]));
Q_AN02 U8227 ( .A0(n6720), .A1(shiftedXdata[241]), .Z(n1660));
Q_MX03 U8228 ( .S0(n2144), .S1(n2402), .A0(ofifoData[241]), .A1(ofifoData[497]), .A2(ofifoData[753]), .Z(n2160));
Q_MX02 U8229 ( .S(n2141), .A0(n1659), .A1(n1660), .Z(ofifoDataN[241]));
Q_AN02 U8230 ( .A0(n6720), .A1(shiftedXdata[242]), .Z(n1658));
Q_MX03 U8231 ( .S0(n2144), .S1(n2402), .A0(ofifoData[242]), .A1(ofifoData[498]), .A2(ofifoData[754]), .Z(n2159));
Q_MX02 U8232 ( .S(n2141), .A0(n1657), .A1(n1658), .Z(ofifoDataN[242]));
Q_AN02 U8233 ( .A0(n6720), .A1(shiftedXdata[243]), .Z(n1656));
Q_MX03 U8234 ( .S0(n2144), .S1(n2402), .A0(ofifoData[243]), .A1(ofifoData[499]), .A2(ofifoData[755]), .Z(n2158));
Q_MX02 U8235 ( .S(n2141), .A0(n1655), .A1(n1656), .Z(ofifoDataN[243]));
Q_AN02 U8236 ( .A0(n6720), .A1(shiftedXdata[244]), .Z(n1654));
Q_MX03 U8237 ( .S0(n2144), .S1(n2402), .A0(ofifoData[244]), .A1(ofifoData[500]), .A2(ofifoData[756]), .Z(n2157));
Q_MX02 U8238 ( .S(n2141), .A0(n1653), .A1(n1654), .Z(ofifoDataN[244]));
Q_AN02 U8239 ( .A0(n6720), .A1(shiftedXdata[245]), .Z(n1652));
Q_MX03 U8240 ( .S0(n2144), .S1(n2402), .A0(ofifoData[245]), .A1(ofifoData[501]), .A2(ofifoData[757]), .Z(n2156));
Q_MX02 U8241 ( .S(n2141), .A0(n1651), .A1(n1652), .Z(ofifoDataN[245]));
Q_AN02 U8242 ( .A0(n6720), .A1(shiftedXdata[246]), .Z(n1650));
Q_MX03 U8243 ( .S0(n2144), .S1(n2402), .A0(ofifoData[246]), .A1(ofifoData[502]), .A2(ofifoData[758]), .Z(n2155));
Q_MX02 U8244 ( .S(n2141), .A0(n1649), .A1(n1650), .Z(ofifoDataN[246]));
Q_AN02 U8245 ( .A0(n6720), .A1(shiftedXdata[247]), .Z(n1648));
Q_MX03 U8246 ( .S0(n2144), .S1(n2402), .A0(ofifoData[247]), .A1(ofifoData[503]), .A2(ofifoData[759]), .Z(n2154));
Q_MX02 U8247 ( .S(n2141), .A0(n1647), .A1(n1648), .Z(ofifoDataN[247]));
Q_AN02 U8248 ( .A0(n6720), .A1(shiftedXdata[248]), .Z(n1646));
Q_MX03 U8249 ( .S0(n2144), .S1(n2402), .A0(ofifoData[248]), .A1(ofifoData[504]), .A2(ofifoData[760]), .Z(n2153));
Q_MX02 U8250 ( .S(n2141), .A0(n1645), .A1(n1646), .Z(ofifoDataN[248]));
Q_AN02 U8251 ( .A0(n6720), .A1(shiftedXdata[249]), .Z(n1644));
Q_MX03 U8252 ( .S0(n2144), .S1(n2402), .A0(ofifoData[249]), .A1(ofifoData[505]), .A2(ofifoData[761]), .Z(n2152));
Q_MX02 U8253 ( .S(n2141), .A0(n1643), .A1(n1644), .Z(ofifoDataN[249]));
Q_AN02 U8254 ( .A0(n6720), .A1(shiftedXdata[250]), .Z(n1642));
Q_MX03 U8255 ( .S0(n2144), .S1(n2402), .A0(ofifoData[250]), .A1(ofifoData[506]), .A2(ofifoData[762]), .Z(n2151));
Q_MX02 U8256 ( .S(n2141), .A0(n1641), .A1(n1642), .Z(ofifoDataN[250]));
Q_AN02 U8257 ( .A0(n6720), .A1(shiftedXdata[251]), .Z(n1640));
Q_MX03 U8258 ( .S0(n2144), .S1(n2402), .A0(ofifoData[251]), .A1(ofifoData[507]), .A2(ofifoData[763]), .Z(n2150));
Q_MX02 U8259 ( .S(n2141), .A0(n1639), .A1(n1640), .Z(ofifoDataN[251]));
Q_AN02 U8260 ( .A0(n6720), .A1(shiftedXdata[252]), .Z(n1638));
Q_MX03 U8261 ( .S0(n2144), .S1(n2402), .A0(ofifoData[252]), .A1(ofifoData[508]), .A2(ofifoData[764]), .Z(n2149));
Q_MX02 U8262 ( .S(n2141), .A0(n1637), .A1(n1638), .Z(ofifoDataN[252]));
Q_AN02 U8263 ( .A0(n6720), .A1(shiftedXdata[253]), .Z(n1636));
Q_MX03 U8264 ( .S0(n2144), .S1(n2402), .A0(ofifoData[253]), .A1(ofifoData[509]), .A2(ofifoData[765]), .Z(n2148));
Q_MX02 U8265 ( .S(n2141), .A0(n1635), .A1(n1636), .Z(ofifoDataN[253]));
Q_AN02 U8266 ( .A0(n6720), .A1(shiftedXdata[254]), .Z(n1634));
Q_MX03 U8267 ( .S0(n2144), .S1(n2402), .A0(ofifoData[254]), .A1(ofifoData[510]), .A2(ofifoData[766]), .Z(n2147));
Q_MX02 U8268 ( .S(n2141), .A0(n1633), .A1(n1634), .Z(ofifoDataN[254]));
Q_AN02 U8269 ( .A0(n6720), .A1(shiftedXdata[255]), .Z(n1632));
Q_MX03 U8270 ( .S0(n2144), .S1(n2402), .A0(ofifoData[255]), .A1(ofifoData[511]), .A2(ofifoData[767]), .Z(n2146));
Q_MX02 U8271 ( .S(n2141), .A0(n1631), .A1(n1632), .Z(ofifoDataN[255]));
Q_AN02 U8272 ( .A0(n6720), .A1(shiftedXdata[256]), .Z(ofifoDataN[256]));
Q_AN02 U8273 ( .A0(n6720), .A1(shiftedXdata[257]), .Z(ofifoDataN[257]));
Q_AN02 U8274 ( .A0(n6720), .A1(shiftedXdata[258]), .Z(ofifoDataN[258]));
Q_AN02 U8275 ( .A0(n6720), .A1(shiftedXdata[259]), .Z(ofifoDataN[259]));
Q_AN02 U8276 ( .A0(n6720), .A1(shiftedXdata[260]), .Z(ofifoDataN[260]));
Q_AN02 U8277 ( .A0(n6720), .A1(shiftedXdata[261]), .Z(ofifoDataN[261]));
Q_AN02 U8278 ( .A0(n6720), .A1(shiftedXdata[262]), .Z(ofifoDataN[262]));
Q_AN02 U8279 ( .A0(n6720), .A1(shiftedXdata[263]), .Z(ofifoDataN[263]));
Q_AN02 U8280 ( .A0(n6720), .A1(shiftedXdata[264]), .Z(ofifoDataN[264]));
Q_AN02 U8281 ( .A0(n6720), .A1(shiftedXdata[265]), .Z(ofifoDataN[265]));
Q_AN02 U8282 ( .A0(n6720), .A1(shiftedXdata[266]), .Z(ofifoDataN[266]));
Q_AN02 U8283 ( .A0(n6720), .A1(shiftedXdata[267]), .Z(ofifoDataN[267]));
Q_AN02 U8284 ( .A0(n6720), .A1(shiftedXdata[268]), .Z(ofifoDataN[268]));
Q_AN02 U8285 ( .A0(n6720), .A1(shiftedXdata[269]), .Z(ofifoDataN[269]));
Q_AN02 U8286 ( .A0(n6720), .A1(shiftedXdata[270]), .Z(ofifoDataN[270]));
Q_AN02 U8287 ( .A0(n6720), .A1(shiftedXdata[271]), .Z(ofifoDataN[271]));
Q_AN02 U8288 ( .A0(n6720), .A1(shiftedXdata[272]), .Z(ofifoDataN[272]));
Q_AN02 U8289 ( .A0(n6720), .A1(shiftedXdata[273]), .Z(ofifoDataN[273]));
Q_AN02 U8290 ( .A0(n6720), .A1(shiftedXdata[274]), .Z(ofifoDataN[274]));
Q_AN02 U8291 ( .A0(n6720), .A1(shiftedXdata[275]), .Z(ofifoDataN[275]));
Q_AN02 U8292 ( .A0(n6720), .A1(shiftedXdata[276]), .Z(ofifoDataN[276]));
Q_AN02 U8293 ( .A0(n6720), .A1(shiftedXdata[277]), .Z(ofifoDataN[277]));
Q_AN02 U8294 ( .A0(n6720), .A1(shiftedXdata[278]), .Z(ofifoDataN[278]));
Q_AN02 U8295 ( .A0(n6720), .A1(shiftedXdata[279]), .Z(ofifoDataN[279]));
Q_AN02 U8296 ( .A0(n6720), .A1(shiftedXdata[280]), .Z(ofifoDataN[280]));
Q_AN02 U8297 ( .A0(n6720), .A1(shiftedXdata[281]), .Z(ofifoDataN[281]));
Q_AN02 U8298 ( .A0(n6720), .A1(shiftedXdata[282]), .Z(ofifoDataN[282]));
Q_AN02 U8299 ( .A0(n6720), .A1(shiftedXdata[283]), .Z(ofifoDataN[283]));
Q_AN02 U8300 ( .A0(n6720), .A1(shiftedXdata[284]), .Z(ofifoDataN[284]));
Q_AN02 U8301 ( .A0(n6720), .A1(shiftedXdata[285]), .Z(ofifoDataN[285]));
Q_AN02 U8302 ( .A0(n6720), .A1(shiftedXdata[286]), .Z(ofifoDataN[286]));
Q_AN02 U8303 ( .A0(n6720), .A1(shiftedXdata[287]), .Z(ofifoDataN[287]));
Q_AN02 U8304 ( .A0(n6720), .A1(shiftedXdata[288]), .Z(ofifoDataN[288]));
Q_AN02 U8305 ( .A0(n6720), .A1(shiftedXdata[289]), .Z(ofifoDataN[289]));
Q_AN02 U8306 ( .A0(n6720), .A1(shiftedXdata[290]), .Z(ofifoDataN[290]));
Q_AN02 U8307 ( .A0(n6720), .A1(shiftedXdata[291]), .Z(ofifoDataN[291]));
Q_AN02 U8308 ( .A0(n6720), .A1(shiftedXdata[292]), .Z(ofifoDataN[292]));
Q_AN02 U8309 ( .A0(n6720), .A1(shiftedXdata[293]), .Z(ofifoDataN[293]));
Q_AN02 U8310 ( .A0(n6720), .A1(shiftedXdata[294]), .Z(ofifoDataN[294]));
Q_AN02 U8311 ( .A0(n6720), .A1(shiftedXdata[295]), .Z(ofifoDataN[295]));
Q_AN02 U8312 ( .A0(n6720), .A1(shiftedXdata[296]), .Z(ofifoDataN[296]));
Q_AN02 U8313 ( .A0(n6720), .A1(shiftedXdata[297]), .Z(ofifoDataN[297]));
Q_AN02 U8314 ( .A0(n6720), .A1(shiftedXdata[298]), .Z(ofifoDataN[298]));
Q_AN02 U8315 ( .A0(n6720), .A1(shiftedXdata[299]), .Z(ofifoDataN[299]));
Q_AN02 U8316 ( .A0(n6720), .A1(shiftedXdata[300]), .Z(ofifoDataN[300]));
Q_AN02 U8317 ( .A0(n6720), .A1(shiftedXdata[301]), .Z(ofifoDataN[301]));
Q_AN02 U8318 ( .A0(n6720), .A1(shiftedXdata[302]), .Z(ofifoDataN[302]));
Q_AN02 U8319 ( .A0(n6720), .A1(shiftedXdata[303]), .Z(ofifoDataN[303]));
Q_AN02 U8320 ( .A0(n6720), .A1(shiftedXdata[304]), .Z(ofifoDataN[304]));
Q_AN02 U8321 ( .A0(n6720), .A1(shiftedXdata[305]), .Z(ofifoDataN[305]));
Q_AN02 U8322 ( .A0(n6720), .A1(shiftedXdata[306]), .Z(ofifoDataN[306]));
Q_AN02 U8323 ( .A0(n6720), .A1(shiftedXdata[307]), .Z(ofifoDataN[307]));
Q_AN02 U8324 ( .A0(n6720), .A1(shiftedXdata[308]), .Z(ofifoDataN[308]));
Q_AN02 U8325 ( .A0(n6720), .A1(shiftedXdata[309]), .Z(ofifoDataN[309]));
Q_AN02 U8326 ( .A0(n6720), .A1(shiftedXdata[310]), .Z(ofifoDataN[310]));
Q_AN02 U8327 ( .A0(n6720), .A1(shiftedXdata[311]), .Z(ofifoDataN[311]));
Q_AN02 U8328 ( .A0(n6720), .A1(shiftedXdata[312]), .Z(ofifoDataN[312]));
Q_AN02 U8329 ( .A0(n6720), .A1(shiftedXdata[313]), .Z(ofifoDataN[313]));
Q_AN02 U8330 ( .A0(n6720), .A1(shiftedXdata[314]), .Z(ofifoDataN[314]));
Q_AN02 U8331 ( .A0(n6720), .A1(shiftedXdata[315]), .Z(ofifoDataN[315]));
Q_AN02 U8332 ( .A0(n6720), .A1(shiftedXdata[316]), .Z(ofifoDataN[316]));
Q_AN02 U8333 ( .A0(n6720), .A1(shiftedXdata[317]), .Z(ofifoDataN[317]));
Q_AN02 U8334 ( .A0(n6720), .A1(shiftedXdata[318]), .Z(ofifoDataN[318]));
Q_AN02 U8335 ( .A0(n6720), .A1(shiftedXdata[319]), .Z(ofifoDataN[319]));
Q_AN02 U8336 ( .A0(n6720), .A1(shiftedXdata[320]), .Z(ofifoDataN[320]));
Q_AN02 U8337 ( .A0(n6720), .A1(shiftedXdata[321]), .Z(ofifoDataN[321]));
Q_AN02 U8338 ( .A0(n6720), .A1(shiftedXdata[322]), .Z(ofifoDataN[322]));
Q_AN02 U8339 ( .A0(n6720), .A1(shiftedXdata[323]), .Z(ofifoDataN[323]));
Q_AN02 U8340 ( .A0(n6720), .A1(shiftedXdata[324]), .Z(ofifoDataN[324]));
Q_AN02 U8341 ( .A0(n6720), .A1(shiftedXdata[325]), .Z(ofifoDataN[325]));
Q_AN02 U8342 ( .A0(n6720), .A1(shiftedXdata[326]), .Z(ofifoDataN[326]));
Q_AN02 U8343 ( .A0(n6720), .A1(shiftedXdata[327]), .Z(ofifoDataN[327]));
Q_AN02 U8344 ( .A0(n6720), .A1(shiftedXdata[328]), .Z(ofifoDataN[328]));
Q_AN02 U8345 ( .A0(n6720), .A1(shiftedXdata[329]), .Z(ofifoDataN[329]));
Q_AN02 U8346 ( .A0(n6720), .A1(shiftedXdata[330]), .Z(ofifoDataN[330]));
Q_AN02 U8347 ( .A0(n6720), .A1(shiftedXdata[331]), .Z(ofifoDataN[331]));
Q_AN02 U8348 ( .A0(n6720), .A1(shiftedXdata[332]), .Z(ofifoDataN[332]));
Q_AN02 U8349 ( .A0(n6720), .A1(shiftedXdata[333]), .Z(ofifoDataN[333]));
Q_AN02 U8350 ( .A0(n6720), .A1(shiftedXdata[334]), .Z(ofifoDataN[334]));
Q_AN02 U8351 ( .A0(n6720), .A1(shiftedXdata[335]), .Z(ofifoDataN[335]));
Q_AN02 U8352 ( .A0(n6720), .A1(shiftedXdata[336]), .Z(ofifoDataN[336]));
Q_AN02 U8353 ( .A0(n6720), .A1(shiftedXdata[337]), .Z(ofifoDataN[337]));
Q_AN02 U8354 ( .A0(n6720), .A1(shiftedXdata[338]), .Z(ofifoDataN[338]));
Q_AN02 U8355 ( .A0(n6720), .A1(shiftedXdata[339]), .Z(ofifoDataN[339]));
Q_AN02 U8356 ( .A0(n6720), .A1(shiftedXdata[340]), .Z(ofifoDataN[340]));
Q_AN02 U8357 ( .A0(n6720), .A1(shiftedXdata[341]), .Z(ofifoDataN[341]));
Q_AN02 U8358 ( .A0(n6720), .A1(shiftedXdata[342]), .Z(ofifoDataN[342]));
Q_AN02 U8359 ( .A0(n6720), .A1(shiftedXdata[343]), .Z(ofifoDataN[343]));
Q_AN02 U8360 ( .A0(n6720), .A1(shiftedXdata[344]), .Z(ofifoDataN[344]));
Q_AN02 U8361 ( .A0(n6720), .A1(shiftedXdata[345]), .Z(ofifoDataN[345]));
Q_AN02 U8362 ( .A0(n6720), .A1(shiftedXdata[346]), .Z(ofifoDataN[346]));
Q_AN02 U8363 ( .A0(n6720), .A1(shiftedXdata[347]), .Z(ofifoDataN[347]));
Q_AN02 U8364 ( .A0(n6720), .A1(shiftedXdata[348]), .Z(ofifoDataN[348]));
Q_AN02 U8365 ( .A0(n6720), .A1(shiftedXdata[349]), .Z(ofifoDataN[349]));
Q_AN02 U8366 ( .A0(n6720), .A1(shiftedXdata[350]), .Z(ofifoDataN[350]));
Q_AN02 U8367 ( .A0(n6720), .A1(shiftedXdata[351]), .Z(ofifoDataN[351]));
Q_AN02 U8368 ( .A0(n6720), .A1(shiftedXdata[352]), .Z(ofifoDataN[352]));
Q_AN02 U8369 ( .A0(n6720), .A1(shiftedXdata[353]), .Z(ofifoDataN[353]));
Q_AN02 U8370 ( .A0(n6720), .A1(shiftedXdata[354]), .Z(ofifoDataN[354]));
Q_AN02 U8371 ( .A0(n6720), .A1(shiftedXdata[355]), .Z(ofifoDataN[355]));
Q_AN02 U8372 ( .A0(n6720), .A1(shiftedXdata[356]), .Z(ofifoDataN[356]));
Q_AN02 U8373 ( .A0(n6720), .A1(shiftedXdata[357]), .Z(ofifoDataN[357]));
Q_AN02 U8374 ( .A0(n6720), .A1(shiftedXdata[358]), .Z(ofifoDataN[358]));
Q_AN02 U8375 ( .A0(n6720), .A1(shiftedXdata[359]), .Z(ofifoDataN[359]));
Q_AN02 U8376 ( .A0(n6720), .A1(shiftedXdata[360]), .Z(ofifoDataN[360]));
Q_AN02 U8377 ( .A0(n6720), .A1(shiftedXdata[361]), .Z(ofifoDataN[361]));
Q_AN02 U8378 ( .A0(n6720), .A1(shiftedXdata[362]), .Z(ofifoDataN[362]));
Q_AN02 U8379 ( .A0(n6720), .A1(shiftedXdata[363]), .Z(ofifoDataN[363]));
Q_AN02 U8380 ( .A0(n6720), .A1(shiftedXdata[364]), .Z(ofifoDataN[364]));
Q_AN02 U8381 ( .A0(n6720), .A1(shiftedXdata[365]), .Z(ofifoDataN[365]));
Q_AN02 U8382 ( .A0(n6720), .A1(shiftedXdata[366]), .Z(ofifoDataN[366]));
Q_AN02 U8383 ( .A0(n6720), .A1(shiftedXdata[367]), .Z(ofifoDataN[367]));
Q_AN02 U8384 ( .A0(n6720), .A1(shiftedXdata[368]), .Z(ofifoDataN[368]));
Q_AN02 U8385 ( .A0(n6720), .A1(shiftedXdata[369]), .Z(ofifoDataN[369]));
Q_AN02 U8386 ( .A0(n6720), .A1(shiftedXdata[370]), .Z(ofifoDataN[370]));
Q_AN02 U8387 ( .A0(n6720), .A1(shiftedXdata[371]), .Z(ofifoDataN[371]));
Q_AN02 U8388 ( .A0(n6720), .A1(shiftedXdata[372]), .Z(ofifoDataN[372]));
Q_AN02 U8389 ( .A0(n6720), .A1(shiftedXdata[373]), .Z(ofifoDataN[373]));
Q_AN02 U8390 ( .A0(n6720), .A1(shiftedXdata[374]), .Z(ofifoDataN[374]));
Q_AN02 U8391 ( .A0(n6720), .A1(shiftedXdata[375]), .Z(ofifoDataN[375]));
Q_AN02 U8392 ( .A0(n6720), .A1(shiftedXdata[376]), .Z(ofifoDataN[376]));
Q_AN02 U8393 ( .A0(n6720), .A1(shiftedXdata[377]), .Z(ofifoDataN[377]));
Q_AN02 U8394 ( .A0(n6720), .A1(shiftedXdata[378]), .Z(ofifoDataN[378]));
Q_AN02 U8395 ( .A0(n6720), .A1(shiftedXdata[379]), .Z(ofifoDataN[379]));
Q_AN02 U8396 ( .A0(n6720), .A1(shiftedXdata[380]), .Z(ofifoDataN[380]));
Q_AN02 U8397 ( .A0(n6720), .A1(shiftedXdata[381]), .Z(ofifoDataN[381]));
Q_AN02 U8398 ( .A0(n6720), .A1(shiftedXdata[382]), .Z(ofifoDataN[382]));
Q_AN02 U8399 ( .A0(n6720), .A1(shiftedXdata[383]), .Z(ofifoDataN[383]));
Q_AN02 U8400 ( .A0(n6720), .A1(shiftedXdata[384]), .Z(ofifoDataN[384]));
Q_AN02 U8401 ( .A0(n6720), .A1(shiftedXdata[385]), .Z(ofifoDataN[385]));
Q_AN02 U8402 ( .A0(n6720), .A1(shiftedXdata[386]), .Z(ofifoDataN[386]));
Q_AN02 U8403 ( .A0(n6720), .A1(shiftedXdata[387]), .Z(ofifoDataN[387]));
Q_AN02 U8404 ( .A0(n6720), .A1(shiftedXdata[388]), .Z(ofifoDataN[388]));
Q_AN02 U8405 ( .A0(n6720), .A1(shiftedXdata[389]), .Z(ofifoDataN[389]));
Q_AN02 U8406 ( .A0(n6720), .A1(shiftedXdata[390]), .Z(ofifoDataN[390]));
Q_AN02 U8407 ( .A0(n6720), .A1(shiftedXdata[391]), .Z(ofifoDataN[391]));
Q_AN02 U8408 ( .A0(n6720), .A1(shiftedXdata[392]), .Z(ofifoDataN[392]));
Q_AN02 U8409 ( .A0(n6720), .A1(shiftedXdata[393]), .Z(ofifoDataN[393]));
Q_AN02 U8410 ( .A0(n6720), .A1(shiftedXdata[394]), .Z(ofifoDataN[394]));
Q_AN02 U8411 ( .A0(n6720), .A1(shiftedXdata[395]), .Z(ofifoDataN[395]));
Q_AN02 U8412 ( .A0(n6720), .A1(shiftedXdata[396]), .Z(ofifoDataN[396]));
Q_AN02 U8413 ( .A0(n6720), .A1(shiftedXdata[397]), .Z(ofifoDataN[397]));
Q_AN02 U8414 ( .A0(n6720), .A1(shiftedXdata[398]), .Z(ofifoDataN[398]));
Q_AN02 U8415 ( .A0(n6720), .A1(shiftedXdata[399]), .Z(ofifoDataN[399]));
Q_AN02 U8416 ( .A0(n6720), .A1(shiftedXdata[400]), .Z(ofifoDataN[400]));
Q_AN02 U8417 ( .A0(n6720), .A1(shiftedXdata[401]), .Z(ofifoDataN[401]));
Q_AN02 U8418 ( .A0(n6720), .A1(shiftedXdata[402]), .Z(ofifoDataN[402]));
Q_AN02 U8419 ( .A0(n6720), .A1(shiftedXdata[403]), .Z(ofifoDataN[403]));
Q_AN02 U8420 ( .A0(n6720), .A1(shiftedXdata[404]), .Z(ofifoDataN[404]));
Q_AN02 U8421 ( .A0(n6720), .A1(shiftedXdata[405]), .Z(ofifoDataN[405]));
Q_AN02 U8422 ( .A0(n6720), .A1(shiftedXdata[406]), .Z(ofifoDataN[406]));
Q_AN02 U8423 ( .A0(n6720), .A1(shiftedXdata[407]), .Z(ofifoDataN[407]));
Q_AN02 U8424 ( .A0(n6720), .A1(shiftedXdata[408]), .Z(ofifoDataN[408]));
Q_AN02 U8425 ( .A0(n6720), .A1(shiftedXdata[409]), .Z(ofifoDataN[409]));
Q_AN02 U8426 ( .A0(n6720), .A1(shiftedXdata[410]), .Z(ofifoDataN[410]));
Q_AN02 U8427 ( .A0(n6720), .A1(shiftedXdata[411]), .Z(ofifoDataN[411]));
Q_AN02 U8428 ( .A0(n6720), .A1(shiftedXdata[412]), .Z(ofifoDataN[412]));
Q_AN02 U8429 ( .A0(n6720), .A1(shiftedXdata[413]), .Z(ofifoDataN[413]));
Q_AN02 U8430 ( .A0(n6720), .A1(shiftedXdata[414]), .Z(ofifoDataN[414]));
Q_AN02 U8431 ( .A0(n6720), .A1(shiftedXdata[415]), .Z(ofifoDataN[415]));
Q_AN02 U8432 ( .A0(n6720), .A1(shiftedXdata[416]), .Z(ofifoDataN[416]));
Q_AN02 U8433 ( .A0(n6720), .A1(shiftedXdata[417]), .Z(ofifoDataN[417]));
Q_AN02 U8434 ( .A0(n6720), .A1(shiftedXdata[418]), .Z(ofifoDataN[418]));
Q_AN02 U8435 ( .A0(n6720), .A1(shiftedXdata[419]), .Z(ofifoDataN[419]));
Q_AN02 U8436 ( .A0(n6720), .A1(shiftedXdata[420]), .Z(ofifoDataN[420]));
Q_AN02 U8437 ( .A0(n6720), .A1(shiftedXdata[421]), .Z(ofifoDataN[421]));
Q_AN02 U8438 ( .A0(n6720), .A1(shiftedXdata[422]), .Z(ofifoDataN[422]));
Q_AN02 U8439 ( .A0(n6720), .A1(shiftedXdata[423]), .Z(ofifoDataN[423]));
Q_AN02 U8440 ( .A0(n6720), .A1(shiftedXdata[424]), .Z(ofifoDataN[424]));
Q_AN02 U8441 ( .A0(n6720), .A1(shiftedXdata[425]), .Z(ofifoDataN[425]));
Q_AN02 U8442 ( .A0(n6720), .A1(shiftedXdata[426]), .Z(ofifoDataN[426]));
Q_AN02 U8443 ( .A0(n6720), .A1(shiftedXdata[427]), .Z(ofifoDataN[427]));
Q_AN02 U8444 ( .A0(n6720), .A1(shiftedXdata[428]), .Z(ofifoDataN[428]));
Q_AN02 U8445 ( .A0(n6720), .A1(shiftedXdata[429]), .Z(ofifoDataN[429]));
Q_AN02 U8446 ( .A0(n6720), .A1(shiftedXdata[430]), .Z(ofifoDataN[430]));
Q_AN02 U8447 ( .A0(n6720), .A1(shiftedXdata[431]), .Z(ofifoDataN[431]));
Q_AN02 U8448 ( .A0(n6720), .A1(shiftedXdata[432]), .Z(ofifoDataN[432]));
Q_AN02 U8449 ( .A0(n6720), .A1(shiftedXdata[433]), .Z(ofifoDataN[433]));
Q_AN02 U8450 ( .A0(n6720), .A1(shiftedXdata[434]), .Z(ofifoDataN[434]));
Q_AN02 U8451 ( .A0(n6720), .A1(shiftedXdata[435]), .Z(ofifoDataN[435]));
Q_AN02 U8452 ( .A0(n6720), .A1(shiftedXdata[436]), .Z(ofifoDataN[436]));
Q_AN02 U8453 ( .A0(n6720), .A1(shiftedXdata[437]), .Z(ofifoDataN[437]));
Q_AN02 U8454 ( .A0(n6720), .A1(shiftedXdata[438]), .Z(ofifoDataN[438]));
Q_AN02 U8455 ( .A0(n6720), .A1(shiftedXdata[439]), .Z(ofifoDataN[439]));
Q_AN02 U8456 ( .A0(n6720), .A1(shiftedXdata[440]), .Z(ofifoDataN[440]));
Q_AN02 U8457 ( .A0(n6720), .A1(shiftedXdata[441]), .Z(ofifoDataN[441]));
Q_AN02 U8458 ( .A0(n6720), .A1(shiftedXdata[442]), .Z(ofifoDataN[442]));
Q_AN02 U8459 ( .A0(n6720), .A1(shiftedXdata[443]), .Z(ofifoDataN[443]));
Q_AN02 U8460 ( .A0(n6720), .A1(shiftedXdata[444]), .Z(ofifoDataN[444]));
Q_AN02 U8461 ( .A0(n6720), .A1(shiftedXdata[445]), .Z(ofifoDataN[445]));
Q_AN02 U8462 ( .A0(n6720), .A1(shiftedXdata[446]), .Z(ofifoDataN[446]));
Q_AN02 U8463 ( .A0(n6720), .A1(shiftedXdata[447]), .Z(ofifoDataN[447]));
Q_AN02 U8464 ( .A0(n6720), .A1(shiftedXdata[448]), .Z(ofifoDataN[448]));
Q_AN02 U8465 ( .A0(n6720), .A1(shiftedXdata[449]), .Z(ofifoDataN[449]));
Q_AN02 U8466 ( .A0(n6720), .A1(shiftedXdata[450]), .Z(ofifoDataN[450]));
Q_AN02 U8467 ( .A0(n6720), .A1(shiftedXdata[451]), .Z(ofifoDataN[451]));
Q_AN02 U8468 ( .A0(n6720), .A1(shiftedXdata[452]), .Z(ofifoDataN[452]));
Q_AN02 U8469 ( .A0(n6720), .A1(shiftedXdata[453]), .Z(ofifoDataN[453]));
Q_AN02 U8470 ( .A0(n6720), .A1(shiftedXdata[454]), .Z(ofifoDataN[454]));
Q_AN02 U8471 ( .A0(n6720), .A1(shiftedXdata[455]), .Z(ofifoDataN[455]));
Q_AN02 U8472 ( .A0(n6720), .A1(shiftedXdata[456]), .Z(ofifoDataN[456]));
Q_AN02 U8473 ( .A0(n6720), .A1(shiftedXdata[457]), .Z(ofifoDataN[457]));
Q_AN02 U8474 ( .A0(n6720), .A1(shiftedXdata[458]), .Z(ofifoDataN[458]));
Q_AN02 U8475 ( .A0(n6720), .A1(shiftedXdata[459]), .Z(ofifoDataN[459]));
Q_AN02 U8476 ( .A0(n6720), .A1(shiftedXdata[460]), .Z(ofifoDataN[460]));
Q_AN02 U8477 ( .A0(n6720), .A1(shiftedXdata[461]), .Z(ofifoDataN[461]));
Q_AN02 U8478 ( .A0(n6720), .A1(shiftedXdata[462]), .Z(ofifoDataN[462]));
Q_AN02 U8479 ( .A0(n6720), .A1(shiftedXdata[463]), .Z(ofifoDataN[463]));
Q_AN02 U8480 ( .A0(n6720), .A1(shiftedXdata[464]), .Z(ofifoDataN[464]));
Q_AN02 U8481 ( .A0(n6720), .A1(shiftedXdata[465]), .Z(ofifoDataN[465]));
Q_AN02 U8482 ( .A0(n6720), .A1(shiftedXdata[466]), .Z(ofifoDataN[466]));
Q_AN02 U8483 ( .A0(n6720), .A1(shiftedXdata[467]), .Z(ofifoDataN[467]));
Q_AN02 U8484 ( .A0(n6720), .A1(shiftedXdata[468]), .Z(ofifoDataN[468]));
Q_AN02 U8485 ( .A0(n6720), .A1(shiftedXdata[469]), .Z(ofifoDataN[469]));
Q_AN02 U8486 ( .A0(n6720), .A1(shiftedXdata[470]), .Z(ofifoDataN[470]));
Q_AN02 U8487 ( .A0(n6720), .A1(shiftedXdata[471]), .Z(ofifoDataN[471]));
Q_AN02 U8488 ( .A0(n6720), .A1(shiftedXdata[472]), .Z(ofifoDataN[472]));
Q_AN02 U8489 ( .A0(n6720), .A1(shiftedXdata[473]), .Z(ofifoDataN[473]));
Q_AN02 U8490 ( .A0(n6720), .A1(shiftedXdata[474]), .Z(ofifoDataN[474]));
Q_AN02 U8491 ( .A0(n6720), .A1(shiftedXdata[475]), .Z(ofifoDataN[475]));
Q_AN02 U8492 ( .A0(n6720), .A1(shiftedXdata[476]), .Z(ofifoDataN[476]));
Q_AN02 U8493 ( .A0(n6720), .A1(shiftedXdata[477]), .Z(ofifoDataN[477]));
Q_AN02 U8494 ( .A0(n6720), .A1(shiftedXdata[478]), .Z(ofifoDataN[478]));
Q_AN02 U8495 ( .A0(n6720), .A1(shiftedXdata[479]), .Z(ofifoDataN[479]));
Q_AN02 U8496 ( .A0(n6720), .A1(shiftedXdata[480]), .Z(ofifoDataN[480]));
Q_AN02 U8497 ( .A0(n6720), .A1(shiftedXdata[481]), .Z(ofifoDataN[481]));
Q_AN02 U8498 ( .A0(n6720), .A1(shiftedXdata[482]), .Z(ofifoDataN[482]));
Q_AN02 U8499 ( .A0(n6720), .A1(shiftedXdata[483]), .Z(ofifoDataN[483]));
Q_AN02 U8500 ( .A0(n6720), .A1(shiftedXdata[484]), .Z(ofifoDataN[484]));
Q_AN02 U8501 ( .A0(n6720), .A1(shiftedXdata[485]), .Z(ofifoDataN[485]));
Q_AN02 U8502 ( .A0(n6720), .A1(shiftedXdata[486]), .Z(ofifoDataN[486]));
Q_AN02 U8503 ( .A0(n6720), .A1(shiftedXdata[487]), .Z(ofifoDataN[487]));
Q_AN02 U8504 ( .A0(n6720), .A1(shiftedXdata[488]), .Z(ofifoDataN[488]));
Q_AN02 U8505 ( .A0(n6720), .A1(shiftedXdata[489]), .Z(ofifoDataN[489]));
Q_AN02 U8506 ( .A0(n6720), .A1(shiftedXdata[490]), .Z(ofifoDataN[490]));
Q_AN02 U8507 ( .A0(n6720), .A1(shiftedXdata[491]), .Z(ofifoDataN[491]));
Q_AN02 U8508 ( .A0(n6720), .A1(shiftedXdata[492]), .Z(ofifoDataN[492]));
Q_AN02 U8509 ( .A0(n6720), .A1(shiftedXdata[493]), .Z(ofifoDataN[493]));
Q_AN02 U8510 ( .A0(n6720), .A1(shiftedXdata[494]), .Z(ofifoDataN[494]));
Q_AN02 U8511 ( .A0(n6720), .A1(shiftedXdata[495]), .Z(ofifoDataN[495]));
Q_AN02 U8512 ( .A0(n6720), .A1(shiftedXdata[496]), .Z(ofifoDataN[496]));
Q_AN02 U8513 ( .A0(n6720), .A1(shiftedXdata[497]), .Z(ofifoDataN[497]));
Q_AN02 U8514 ( .A0(n6720), .A1(shiftedXdata[498]), .Z(ofifoDataN[498]));
Q_AN02 U8515 ( .A0(n6720), .A1(shiftedXdata[499]), .Z(ofifoDataN[499]));
Q_AN02 U8516 ( .A0(n6720), .A1(shiftedXdata[500]), .Z(ofifoDataN[500]));
Q_AN02 U8517 ( .A0(n6720), .A1(shiftedXdata[501]), .Z(ofifoDataN[501]));
Q_AN02 U8518 ( .A0(n6720), .A1(shiftedXdata[502]), .Z(ofifoDataN[502]));
Q_AN02 U8519 ( .A0(n6720), .A1(shiftedXdata[503]), .Z(ofifoDataN[503]));
Q_AN02 U8520 ( .A0(n6720), .A1(shiftedXdata[504]), .Z(ofifoDataN[504]));
Q_AN02 U8521 ( .A0(n6720), .A1(shiftedXdata[505]), .Z(ofifoDataN[505]));
Q_AN02 U8522 ( .A0(n6720), .A1(shiftedXdata[506]), .Z(ofifoDataN[506]));
Q_AN02 U8523 ( .A0(n6720), .A1(shiftedXdata[507]), .Z(ofifoDataN[507]));
Q_AN02 U8524 ( .A0(n6720), .A1(shiftedXdata[508]), .Z(ofifoDataN[508]));
Q_AN02 U8525 ( .A0(n6720), .A1(shiftedXdata[509]), .Z(ofifoDataN[509]));
Q_AN02 U8526 ( .A0(n6720), .A1(shiftedXdata[510]), .Z(ofifoDataN[510]));
Q_AN02 U8527 ( .A0(n6720), .A1(shiftedXdata[511]), .Z(ofifoDataN[511]));
Q_AN02 U8528 ( .A0(n6720), .A1(shiftedXdata[512]), .Z(ofifoDataN[512]));
Q_AN02 U8529 ( .A0(n6720), .A1(shiftedXdata[513]), .Z(ofifoDataN[513]));
Q_AN02 U8530 ( .A0(n6720), .A1(shiftedXdata[514]), .Z(ofifoDataN[514]));
Q_AN02 U8531 ( .A0(n6720), .A1(shiftedXdata[515]), .Z(ofifoDataN[515]));
Q_AN02 U8532 ( .A0(n6720), .A1(shiftedXdata[516]), .Z(ofifoDataN[516]));
Q_AN02 U8533 ( .A0(n6720), .A1(shiftedXdata[517]), .Z(ofifoDataN[517]));
Q_AN02 U8534 ( .A0(n6720), .A1(shiftedXdata[518]), .Z(ofifoDataN[518]));
Q_AN02 U8535 ( .A0(n6720), .A1(shiftedXdata[519]), .Z(ofifoDataN[519]));
Q_AN02 U8536 ( .A0(n6720), .A1(shiftedXdata[520]), .Z(ofifoDataN[520]));
Q_AN02 U8537 ( .A0(n6720), .A1(shiftedXdata[521]), .Z(ofifoDataN[521]));
Q_AN02 U8538 ( .A0(n6720), .A1(shiftedXdata[522]), .Z(ofifoDataN[522]));
Q_AN02 U8539 ( .A0(n6720), .A1(shiftedXdata[523]), .Z(ofifoDataN[523]));
Q_AN02 U8540 ( .A0(n6720), .A1(shiftedXdata[524]), .Z(ofifoDataN[524]));
Q_AN02 U8541 ( .A0(n6720), .A1(shiftedXdata[525]), .Z(ofifoDataN[525]));
Q_AN02 U8542 ( .A0(n6720), .A1(shiftedXdata[526]), .Z(ofifoDataN[526]));
Q_AN02 U8543 ( .A0(n6720), .A1(shiftedXdata[527]), .Z(ofifoDataN[527]));
Q_AN02 U8544 ( .A0(n6720), .A1(shiftedXdata[528]), .Z(ofifoDataN[528]));
Q_AN02 U8545 ( .A0(n6720), .A1(shiftedXdata[529]), .Z(ofifoDataN[529]));
Q_AN02 U8546 ( .A0(n6720), .A1(shiftedXdata[530]), .Z(ofifoDataN[530]));
Q_AN02 U8547 ( .A0(n6720), .A1(shiftedXdata[531]), .Z(ofifoDataN[531]));
Q_AN02 U8548 ( .A0(n6720), .A1(shiftedXdata[532]), .Z(ofifoDataN[532]));
Q_AN02 U8549 ( .A0(n6720), .A1(shiftedXdata[533]), .Z(ofifoDataN[533]));
Q_AN02 U8550 ( .A0(n6720), .A1(shiftedXdata[534]), .Z(ofifoDataN[534]));
Q_AN02 U8551 ( .A0(n6720), .A1(shiftedXdata[535]), .Z(ofifoDataN[535]));
Q_AN02 U8552 ( .A0(n6720), .A1(shiftedXdata[536]), .Z(ofifoDataN[536]));
Q_AN02 U8553 ( .A0(n6720), .A1(shiftedXdata[537]), .Z(ofifoDataN[537]));
Q_AN02 U8554 ( .A0(n6720), .A1(shiftedXdata[538]), .Z(ofifoDataN[538]));
Q_AN02 U8555 ( .A0(n6720), .A1(shiftedXdata[539]), .Z(ofifoDataN[539]));
Q_AN02 U8556 ( .A0(n6720), .A1(shiftedXdata[540]), .Z(ofifoDataN[540]));
Q_AN02 U8557 ( .A0(n6720), .A1(shiftedXdata[541]), .Z(ofifoDataN[541]));
Q_AN02 U8558 ( .A0(n6720), .A1(shiftedXdata[542]), .Z(ofifoDataN[542]));
Q_AN02 U8559 ( .A0(n6720), .A1(shiftedXdata[543]), .Z(ofifoDataN[543]));
Q_AN02 U8560 ( .A0(n6720), .A1(shiftedXdata[544]), .Z(ofifoDataN[544]));
Q_AN02 U8561 ( .A0(n6720), .A1(shiftedXdata[545]), .Z(ofifoDataN[545]));
Q_AN02 U8562 ( .A0(n6720), .A1(shiftedXdata[546]), .Z(ofifoDataN[546]));
Q_AN02 U8563 ( .A0(n6720), .A1(shiftedXdata[547]), .Z(ofifoDataN[547]));
Q_AN02 U8564 ( .A0(n6720), .A1(shiftedXdata[548]), .Z(ofifoDataN[548]));
Q_AN02 U8565 ( .A0(n6720), .A1(shiftedXdata[549]), .Z(ofifoDataN[549]));
Q_AN02 U8566 ( .A0(n6720), .A1(shiftedXdata[550]), .Z(ofifoDataN[550]));
Q_AN02 U8567 ( .A0(n6720), .A1(shiftedXdata[551]), .Z(ofifoDataN[551]));
Q_AN02 U8568 ( .A0(n6720), .A1(shiftedXdata[552]), .Z(ofifoDataN[552]));
Q_AN02 U8569 ( .A0(n6720), .A1(shiftedXdata[553]), .Z(ofifoDataN[553]));
Q_AN02 U8570 ( .A0(n6720), .A1(shiftedXdata[554]), .Z(ofifoDataN[554]));
Q_AN02 U8571 ( .A0(n6720), .A1(shiftedXdata[555]), .Z(ofifoDataN[555]));
Q_AN02 U8572 ( .A0(n6720), .A1(shiftedXdata[556]), .Z(ofifoDataN[556]));
Q_AN02 U8573 ( .A0(n6720), .A1(shiftedXdata[557]), .Z(ofifoDataN[557]));
Q_AN02 U8574 ( .A0(n6720), .A1(shiftedXdata[558]), .Z(ofifoDataN[558]));
Q_AN02 U8575 ( .A0(n6720), .A1(shiftedXdata[559]), .Z(ofifoDataN[559]));
Q_AN02 U8576 ( .A0(n6720), .A1(shiftedXdata[560]), .Z(ofifoDataN[560]));
Q_AN02 U8577 ( .A0(n6720), .A1(shiftedXdata[561]), .Z(ofifoDataN[561]));
Q_AN02 U8578 ( .A0(n6720), .A1(shiftedXdata[562]), .Z(ofifoDataN[562]));
Q_AN02 U8579 ( .A0(n6720), .A1(shiftedXdata[563]), .Z(ofifoDataN[563]));
Q_AN02 U8580 ( .A0(n6720), .A1(shiftedXdata[564]), .Z(ofifoDataN[564]));
Q_AN02 U8581 ( .A0(n6720), .A1(shiftedXdata[565]), .Z(ofifoDataN[565]));
Q_AN02 U8582 ( .A0(n6720), .A1(shiftedXdata[566]), .Z(ofifoDataN[566]));
Q_AN02 U8583 ( .A0(n6720), .A1(shiftedXdata[567]), .Z(ofifoDataN[567]));
Q_AN02 U8584 ( .A0(n6720), .A1(shiftedXdata[568]), .Z(ofifoDataN[568]));
Q_AN02 U8585 ( .A0(n6720), .A1(shiftedXdata[569]), .Z(ofifoDataN[569]));
Q_AN02 U8586 ( .A0(n6720), .A1(shiftedXdata[570]), .Z(ofifoDataN[570]));
Q_AN02 U8587 ( .A0(n6720), .A1(shiftedXdata[571]), .Z(ofifoDataN[571]));
Q_AN02 U8588 ( .A0(n6720), .A1(shiftedXdata[572]), .Z(ofifoDataN[572]));
Q_AN02 U8589 ( .A0(n6720), .A1(shiftedXdata[573]), .Z(ofifoDataN[573]));
Q_AN02 U8590 ( .A0(n6720), .A1(shiftedXdata[574]), .Z(ofifoDataN[574]));
Q_AN02 U8591 ( .A0(n6720), .A1(shiftedXdata[575]), .Z(ofifoDataN[575]));
Q_AN02 U8592 ( .A0(n6720), .A1(shiftedXdata[576]), .Z(ofifoDataN[576]));
Q_AN02 U8593 ( .A0(n6720), .A1(shiftedXdata[577]), .Z(ofifoDataN[577]));
Q_AN02 U8594 ( .A0(n6720), .A1(shiftedXdata[578]), .Z(ofifoDataN[578]));
Q_AN02 U8595 ( .A0(n6720), .A1(shiftedXdata[579]), .Z(ofifoDataN[579]));
Q_AN02 U8596 ( .A0(n6720), .A1(shiftedXdata[580]), .Z(ofifoDataN[580]));
Q_AN02 U8597 ( .A0(n6720), .A1(shiftedXdata[581]), .Z(ofifoDataN[581]));
Q_AN02 U8598 ( .A0(n6720), .A1(shiftedXdata[582]), .Z(ofifoDataN[582]));
Q_AN02 U8599 ( .A0(n6720), .A1(shiftedXdata[583]), .Z(ofifoDataN[583]));
Q_AN02 U8600 ( .A0(n6720), .A1(shiftedXdata[584]), .Z(ofifoDataN[584]));
Q_AN02 U8601 ( .A0(n6720), .A1(shiftedXdata[585]), .Z(ofifoDataN[585]));
Q_AN02 U8602 ( .A0(n6720), .A1(shiftedXdata[586]), .Z(ofifoDataN[586]));
Q_AN02 U8603 ( .A0(n6720), .A1(shiftedXdata[587]), .Z(ofifoDataN[587]));
Q_AN02 U8604 ( .A0(n6720), .A1(shiftedXdata[588]), .Z(ofifoDataN[588]));
Q_AN02 U8605 ( .A0(n6720), .A1(shiftedXdata[589]), .Z(ofifoDataN[589]));
Q_AN02 U8606 ( .A0(n6720), .A1(shiftedXdata[590]), .Z(ofifoDataN[590]));
Q_AN02 U8607 ( .A0(n6720), .A1(shiftedXdata[591]), .Z(ofifoDataN[591]));
Q_AN02 U8608 ( .A0(n6720), .A1(shiftedXdata[592]), .Z(ofifoDataN[592]));
Q_AN02 U8609 ( .A0(n6720), .A1(shiftedXdata[593]), .Z(ofifoDataN[593]));
Q_AN02 U8610 ( .A0(n6720), .A1(shiftedXdata[594]), .Z(ofifoDataN[594]));
Q_AN02 U8611 ( .A0(n6720), .A1(shiftedXdata[595]), .Z(ofifoDataN[595]));
Q_AN02 U8612 ( .A0(n6720), .A1(shiftedXdata[596]), .Z(ofifoDataN[596]));
Q_AN02 U8613 ( .A0(n6720), .A1(shiftedXdata[597]), .Z(ofifoDataN[597]));
Q_AN02 U8614 ( .A0(n6720), .A1(shiftedXdata[598]), .Z(ofifoDataN[598]));
Q_AN02 U8615 ( .A0(n6720), .A1(shiftedXdata[599]), .Z(ofifoDataN[599]));
Q_AN02 U8616 ( .A0(n6720), .A1(shiftedXdata[600]), .Z(ofifoDataN[600]));
Q_AN02 U8617 ( .A0(n6720), .A1(shiftedXdata[601]), .Z(ofifoDataN[601]));
Q_AN02 U8618 ( .A0(n6720), .A1(shiftedXdata[602]), .Z(ofifoDataN[602]));
Q_AN02 U8619 ( .A0(n6720), .A1(shiftedXdata[603]), .Z(ofifoDataN[603]));
Q_AN02 U8620 ( .A0(n6720), .A1(shiftedXdata[604]), .Z(ofifoDataN[604]));
Q_AN02 U8621 ( .A0(n6720), .A1(shiftedXdata[605]), .Z(ofifoDataN[605]));
Q_AN02 U8622 ( .A0(n6720), .A1(shiftedXdata[606]), .Z(ofifoDataN[606]));
Q_AN02 U8623 ( .A0(n6720), .A1(shiftedXdata[607]), .Z(ofifoDataN[607]));
Q_AN02 U8624 ( .A0(n6720), .A1(shiftedXdata[608]), .Z(ofifoDataN[608]));
Q_AN02 U8625 ( .A0(n6720), .A1(shiftedXdata[609]), .Z(ofifoDataN[609]));
Q_AN02 U8626 ( .A0(n6720), .A1(shiftedXdata[610]), .Z(ofifoDataN[610]));
Q_AN02 U8627 ( .A0(n6720), .A1(shiftedXdata[611]), .Z(ofifoDataN[611]));
Q_AN02 U8628 ( .A0(n6720), .A1(shiftedXdata[612]), .Z(ofifoDataN[612]));
Q_AN02 U8629 ( .A0(n6720), .A1(shiftedXdata[613]), .Z(ofifoDataN[613]));
Q_AN02 U8630 ( .A0(n6720), .A1(shiftedXdata[614]), .Z(ofifoDataN[614]));
Q_AN02 U8631 ( .A0(n6720), .A1(shiftedXdata[615]), .Z(ofifoDataN[615]));
Q_AN02 U8632 ( .A0(n6720), .A1(shiftedXdata[616]), .Z(ofifoDataN[616]));
Q_AN02 U8633 ( .A0(n6720), .A1(shiftedXdata[617]), .Z(ofifoDataN[617]));
Q_AN02 U8634 ( .A0(n6720), .A1(shiftedXdata[618]), .Z(ofifoDataN[618]));
Q_AN02 U8635 ( .A0(n6720), .A1(shiftedXdata[619]), .Z(ofifoDataN[619]));
Q_AN02 U8636 ( .A0(n6720), .A1(shiftedXdata[620]), .Z(ofifoDataN[620]));
Q_AN02 U8637 ( .A0(n6720), .A1(shiftedXdata[621]), .Z(ofifoDataN[621]));
Q_AN02 U8638 ( .A0(n6720), .A1(shiftedXdata[622]), .Z(ofifoDataN[622]));
Q_AN02 U8639 ( .A0(n6720), .A1(shiftedXdata[623]), .Z(ofifoDataN[623]));
Q_AN02 U8640 ( .A0(n6720), .A1(shiftedXdata[624]), .Z(ofifoDataN[624]));
Q_AN02 U8641 ( .A0(n6720), .A1(shiftedXdata[625]), .Z(ofifoDataN[625]));
Q_AN02 U8642 ( .A0(n6720), .A1(shiftedXdata[626]), .Z(ofifoDataN[626]));
Q_AN02 U8643 ( .A0(n6720), .A1(shiftedXdata[627]), .Z(ofifoDataN[627]));
Q_AN02 U8644 ( .A0(n6720), .A1(shiftedXdata[628]), .Z(ofifoDataN[628]));
Q_AN02 U8645 ( .A0(n6720), .A1(shiftedXdata[629]), .Z(ofifoDataN[629]));
Q_AN02 U8646 ( .A0(n6720), .A1(shiftedXdata[630]), .Z(ofifoDataN[630]));
Q_AN02 U8647 ( .A0(n6720), .A1(shiftedXdata[631]), .Z(ofifoDataN[631]));
Q_AN02 U8648 ( .A0(n6720), .A1(shiftedXdata[632]), .Z(ofifoDataN[632]));
Q_AN02 U8649 ( .A0(n6720), .A1(shiftedXdata[633]), .Z(ofifoDataN[633]));
Q_AN02 U8650 ( .A0(n6720), .A1(shiftedXdata[634]), .Z(ofifoDataN[634]));
Q_AN02 U8651 ( .A0(n6720), .A1(shiftedXdata[635]), .Z(ofifoDataN[635]));
Q_AN02 U8652 ( .A0(n6720), .A1(shiftedXdata[636]), .Z(ofifoDataN[636]));
Q_AN02 U8653 ( .A0(n6720), .A1(shiftedXdata[637]), .Z(ofifoDataN[637]));
Q_AN02 U8654 ( .A0(n6720), .A1(shiftedXdata[638]), .Z(ofifoDataN[638]));
Q_AN02 U8655 ( .A0(n6720), .A1(shiftedXdata[639]), .Z(ofifoDataN[639]));
Q_AN02 U8656 ( .A0(n6720), .A1(shiftedXdata[640]), .Z(ofifoDataN[640]));
Q_AN02 U8657 ( .A0(n6720), .A1(shiftedXdata[641]), .Z(ofifoDataN[641]));
Q_AN02 U8658 ( .A0(n6720), .A1(shiftedXdata[642]), .Z(ofifoDataN[642]));
Q_AN02 U8659 ( .A0(n6720), .A1(shiftedXdata[643]), .Z(ofifoDataN[643]));
Q_AN02 U8660 ( .A0(n6720), .A1(shiftedXdata[644]), .Z(ofifoDataN[644]));
Q_AN02 U8661 ( .A0(n6720), .A1(shiftedXdata[645]), .Z(ofifoDataN[645]));
Q_AN02 U8662 ( .A0(n6720), .A1(shiftedXdata[646]), .Z(ofifoDataN[646]));
Q_AN02 U8663 ( .A0(n6720), .A1(shiftedXdata[647]), .Z(ofifoDataN[647]));
Q_AN02 U8664 ( .A0(n6720), .A1(shiftedXdata[648]), .Z(ofifoDataN[648]));
Q_AN02 U8665 ( .A0(n6720), .A1(shiftedXdata[649]), .Z(ofifoDataN[649]));
Q_AN02 U8666 ( .A0(n6720), .A1(shiftedXdata[650]), .Z(ofifoDataN[650]));
Q_AN02 U8667 ( .A0(n6720), .A1(shiftedXdata[651]), .Z(ofifoDataN[651]));
Q_AN02 U8668 ( .A0(n6720), .A1(shiftedXdata[652]), .Z(ofifoDataN[652]));
Q_AN02 U8669 ( .A0(n6720), .A1(shiftedXdata[653]), .Z(ofifoDataN[653]));
Q_AN02 U8670 ( .A0(n6720), .A1(shiftedXdata[654]), .Z(ofifoDataN[654]));
Q_AN02 U8671 ( .A0(n6720), .A1(shiftedXdata[655]), .Z(ofifoDataN[655]));
Q_AN02 U8672 ( .A0(n6720), .A1(shiftedXdata[656]), .Z(ofifoDataN[656]));
Q_AN02 U8673 ( .A0(n6720), .A1(shiftedXdata[657]), .Z(ofifoDataN[657]));
Q_AN02 U8674 ( .A0(n6720), .A1(shiftedXdata[658]), .Z(ofifoDataN[658]));
Q_AN02 U8675 ( .A0(n6720), .A1(shiftedXdata[659]), .Z(ofifoDataN[659]));
Q_AN02 U8676 ( .A0(n6720), .A1(shiftedXdata[660]), .Z(ofifoDataN[660]));
Q_AN02 U8677 ( .A0(n6720), .A1(shiftedXdata[661]), .Z(ofifoDataN[661]));
Q_AN02 U8678 ( .A0(n6720), .A1(shiftedXdata[662]), .Z(ofifoDataN[662]));
Q_AN02 U8679 ( .A0(n6720), .A1(shiftedXdata[663]), .Z(ofifoDataN[663]));
Q_AN02 U8680 ( .A0(n6720), .A1(shiftedXdata[664]), .Z(ofifoDataN[664]));
Q_AN02 U8681 ( .A0(n6720), .A1(shiftedXdata[665]), .Z(ofifoDataN[665]));
Q_AN02 U8682 ( .A0(n6720), .A1(shiftedXdata[666]), .Z(ofifoDataN[666]));
Q_AN02 U8683 ( .A0(n6720), .A1(shiftedXdata[667]), .Z(ofifoDataN[667]));
Q_AN02 U8684 ( .A0(n6720), .A1(shiftedXdata[668]), .Z(ofifoDataN[668]));
Q_AN02 U8685 ( .A0(n6720), .A1(shiftedXdata[669]), .Z(ofifoDataN[669]));
Q_AN02 U8686 ( .A0(n6720), .A1(shiftedXdata[670]), .Z(ofifoDataN[670]));
Q_AN02 U8687 ( .A0(n6720), .A1(shiftedXdata[671]), .Z(ofifoDataN[671]));
Q_AN02 U8688 ( .A0(n6720), .A1(shiftedXdata[672]), .Z(ofifoDataN[672]));
Q_AN02 U8689 ( .A0(n6720), .A1(shiftedXdata[673]), .Z(ofifoDataN[673]));
Q_AN02 U8690 ( .A0(n6720), .A1(shiftedXdata[674]), .Z(ofifoDataN[674]));
Q_AN02 U8691 ( .A0(n6720), .A1(shiftedXdata[675]), .Z(ofifoDataN[675]));
Q_AN02 U8692 ( .A0(n6720), .A1(shiftedXdata[676]), .Z(ofifoDataN[676]));
Q_AN02 U8693 ( .A0(n6720), .A1(shiftedXdata[677]), .Z(ofifoDataN[677]));
Q_AN02 U8694 ( .A0(n6720), .A1(shiftedXdata[678]), .Z(ofifoDataN[678]));
Q_AN02 U8695 ( .A0(n6720), .A1(shiftedXdata[679]), .Z(ofifoDataN[679]));
Q_AN02 U8696 ( .A0(n6720), .A1(shiftedXdata[680]), .Z(ofifoDataN[680]));
Q_AN02 U8697 ( .A0(n6720), .A1(shiftedXdata[681]), .Z(ofifoDataN[681]));
Q_AN02 U8698 ( .A0(n6720), .A1(shiftedXdata[682]), .Z(ofifoDataN[682]));
Q_AN02 U8699 ( .A0(n6720), .A1(shiftedXdata[683]), .Z(ofifoDataN[683]));
Q_AN02 U8700 ( .A0(n6720), .A1(shiftedXdata[684]), .Z(ofifoDataN[684]));
Q_AN02 U8701 ( .A0(n6720), .A1(shiftedXdata[685]), .Z(ofifoDataN[685]));
Q_AN02 U8702 ( .A0(n6720), .A1(shiftedXdata[686]), .Z(ofifoDataN[686]));
Q_AN02 U8703 ( .A0(n6720), .A1(shiftedXdata[687]), .Z(ofifoDataN[687]));
Q_AN02 U8704 ( .A0(n6720), .A1(shiftedXdata[688]), .Z(ofifoDataN[688]));
Q_AN02 U8705 ( .A0(n6720), .A1(shiftedXdata[689]), .Z(ofifoDataN[689]));
Q_AN02 U8706 ( .A0(n6720), .A1(shiftedXdata[690]), .Z(ofifoDataN[690]));
Q_AN02 U8707 ( .A0(n6720), .A1(shiftedXdata[691]), .Z(ofifoDataN[691]));
Q_AN02 U8708 ( .A0(n6720), .A1(shiftedXdata[692]), .Z(ofifoDataN[692]));
Q_AN02 U8709 ( .A0(n6720), .A1(shiftedXdata[693]), .Z(ofifoDataN[693]));
Q_AN02 U8710 ( .A0(n6720), .A1(shiftedXdata[694]), .Z(ofifoDataN[694]));
Q_AN02 U8711 ( .A0(n6720), .A1(shiftedXdata[695]), .Z(ofifoDataN[695]));
Q_AN02 U8712 ( .A0(n6720), .A1(shiftedXdata[696]), .Z(ofifoDataN[696]));
Q_AN02 U8713 ( .A0(n6720), .A1(shiftedXdata[697]), .Z(ofifoDataN[697]));
Q_AN02 U8714 ( .A0(n6720), .A1(shiftedXdata[698]), .Z(ofifoDataN[698]));
Q_AN02 U8715 ( .A0(n6720), .A1(shiftedXdata[699]), .Z(ofifoDataN[699]));
Q_AN02 U8716 ( .A0(n6720), .A1(shiftedXdata[700]), .Z(ofifoDataN[700]));
Q_AN02 U8717 ( .A0(n6720), .A1(shiftedXdata[701]), .Z(ofifoDataN[701]));
Q_AN02 U8718 ( .A0(n6720), .A1(shiftedXdata[702]), .Z(ofifoDataN[702]));
Q_AN02 U8719 ( .A0(n6720), .A1(shiftedXdata[703]), .Z(ofifoDataN[703]));
Q_AN02 U8720 ( .A0(n6720), .A1(shiftedXdata[704]), .Z(ofifoDataN[704]));
Q_AN02 U8721 ( .A0(n6720), .A1(shiftedXdata[705]), .Z(ofifoDataN[705]));
Q_AN02 U8722 ( .A0(n6720), .A1(shiftedXdata[706]), .Z(ofifoDataN[706]));
Q_AN02 U8723 ( .A0(n6720), .A1(shiftedXdata[707]), .Z(ofifoDataN[707]));
Q_AN02 U8724 ( .A0(n6720), .A1(shiftedXdata[708]), .Z(ofifoDataN[708]));
Q_AN02 U8725 ( .A0(n6720), .A1(shiftedXdata[709]), .Z(ofifoDataN[709]));
Q_AN02 U8726 ( .A0(n6720), .A1(shiftedXdata[710]), .Z(ofifoDataN[710]));
Q_AN02 U8727 ( .A0(n6720), .A1(shiftedXdata[711]), .Z(ofifoDataN[711]));
Q_AN02 U8728 ( .A0(n6720), .A1(shiftedXdata[712]), .Z(ofifoDataN[712]));
Q_AN02 U8729 ( .A0(n6720), .A1(shiftedXdata[713]), .Z(ofifoDataN[713]));
Q_AN02 U8730 ( .A0(n6720), .A1(shiftedXdata[714]), .Z(ofifoDataN[714]));
Q_AN02 U8731 ( .A0(n6720), .A1(shiftedXdata[715]), .Z(ofifoDataN[715]));
Q_AN02 U8732 ( .A0(n6720), .A1(shiftedXdata[716]), .Z(ofifoDataN[716]));
Q_AN02 U8733 ( .A0(n6720), .A1(shiftedXdata[717]), .Z(ofifoDataN[717]));
Q_AN02 U8734 ( .A0(n6720), .A1(shiftedXdata[718]), .Z(ofifoDataN[718]));
Q_AN02 U8735 ( .A0(n6720), .A1(shiftedXdata[719]), .Z(ofifoDataN[719]));
Q_AN02 U8736 ( .A0(n6720), .A1(shiftedXdata[720]), .Z(ofifoDataN[720]));
Q_AN02 U8737 ( .A0(n6720), .A1(shiftedXdata[721]), .Z(ofifoDataN[721]));
Q_AN02 U8738 ( .A0(n6720), .A1(shiftedXdata[722]), .Z(ofifoDataN[722]));
Q_AN02 U8739 ( .A0(n6720), .A1(shiftedXdata[723]), .Z(ofifoDataN[723]));
Q_AN02 U8740 ( .A0(n6720), .A1(shiftedXdata[724]), .Z(ofifoDataN[724]));
Q_AN02 U8741 ( .A0(n6720), .A1(shiftedXdata[725]), .Z(ofifoDataN[725]));
Q_AN02 U8742 ( .A0(n6720), .A1(shiftedXdata[726]), .Z(ofifoDataN[726]));
Q_AN02 U8743 ( .A0(n6720), .A1(shiftedXdata[727]), .Z(ofifoDataN[727]));
Q_AN02 U8744 ( .A0(n6720), .A1(shiftedXdata[728]), .Z(ofifoDataN[728]));
Q_AN02 U8745 ( .A0(n6720), .A1(shiftedXdata[729]), .Z(ofifoDataN[729]));
Q_AN02 U8746 ( .A0(n6720), .A1(shiftedXdata[730]), .Z(ofifoDataN[730]));
Q_AN02 U8747 ( .A0(n6720), .A1(shiftedXdata[731]), .Z(ofifoDataN[731]));
Q_AN02 U8748 ( .A0(n6720), .A1(shiftedXdata[732]), .Z(ofifoDataN[732]));
Q_AN02 U8749 ( .A0(n6720), .A1(shiftedXdata[733]), .Z(ofifoDataN[733]));
Q_AN02 U8750 ( .A0(n6720), .A1(shiftedXdata[734]), .Z(ofifoDataN[734]));
Q_AN02 U8751 ( .A0(n6720), .A1(shiftedXdata[735]), .Z(ofifoDataN[735]));
Q_AN02 U8752 ( .A0(n6720), .A1(shiftedXdata[736]), .Z(ofifoDataN[736]));
Q_AN02 U8753 ( .A0(n6720), .A1(shiftedXdata[737]), .Z(ofifoDataN[737]));
Q_AN02 U8754 ( .A0(n6720), .A1(shiftedXdata[738]), .Z(ofifoDataN[738]));
Q_AN02 U8755 ( .A0(n6720), .A1(shiftedXdata[739]), .Z(ofifoDataN[739]));
Q_AN02 U8756 ( .A0(n6720), .A1(shiftedXdata[740]), .Z(ofifoDataN[740]));
Q_AN02 U8757 ( .A0(n6720), .A1(shiftedXdata[741]), .Z(ofifoDataN[741]));
Q_AN02 U8758 ( .A0(n6720), .A1(shiftedXdata[742]), .Z(ofifoDataN[742]));
Q_AN02 U8759 ( .A0(n6720), .A1(shiftedXdata[743]), .Z(ofifoDataN[743]));
Q_AN02 U8760 ( .A0(n6720), .A1(shiftedXdata[744]), .Z(ofifoDataN[744]));
Q_AN02 U8761 ( .A0(n6720), .A1(shiftedXdata[745]), .Z(ofifoDataN[745]));
Q_AN02 U8762 ( .A0(n6720), .A1(shiftedXdata[746]), .Z(ofifoDataN[746]));
Q_AN02 U8763 ( .A0(n6720), .A1(shiftedXdata[747]), .Z(ofifoDataN[747]));
Q_AN02 U8764 ( .A0(n6720), .A1(shiftedXdata[748]), .Z(ofifoDataN[748]));
Q_AN02 U8765 ( .A0(n6720), .A1(shiftedXdata[749]), .Z(ofifoDataN[749]));
Q_AN02 U8766 ( .A0(n6720), .A1(shiftedXdata[750]), .Z(ofifoDataN[750]));
Q_AN02 U8767 ( .A0(n6720), .A1(shiftedXdata[751]), .Z(ofifoDataN[751]));
Q_AN02 U8768 ( .A0(n6720), .A1(shiftedXdata[752]), .Z(ofifoDataN[752]));
Q_AN02 U8769 ( .A0(n6720), .A1(shiftedXdata[753]), .Z(ofifoDataN[753]));
Q_AN02 U8770 ( .A0(n6720), .A1(shiftedXdata[754]), .Z(ofifoDataN[754]));
Q_AN02 U8771 ( .A0(n6720), .A1(shiftedXdata[755]), .Z(ofifoDataN[755]));
Q_AN02 U8772 ( .A0(n6720), .A1(shiftedXdata[756]), .Z(ofifoDataN[756]));
Q_AN02 U8773 ( .A0(n6720), .A1(shiftedXdata[757]), .Z(ofifoDataN[757]));
Q_AN02 U8774 ( .A0(n6720), .A1(shiftedXdata[758]), .Z(ofifoDataN[758]));
Q_AN02 U8775 ( .A0(n6720), .A1(shiftedXdata[759]), .Z(ofifoDataN[759]));
Q_AN02 U8776 ( .A0(n6720), .A1(shiftedXdata[760]), .Z(ofifoDataN[760]));
Q_AN02 U8777 ( .A0(n6720), .A1(shiftedXdata[761]), .Z(ofifoDataN[761]));
Q_AN02 U8778 ( .A0(n6720), .A1(shiftedXdata[762]), .Z(ofifoDataN[762]));
Q_AN02 U8779 ( .A0(n6720), .A1(shiftedXdata[763]), .Z(ofifoDataN[763]));
Q_AN02 U8780 ( .A0(n6720), .A1(shiftedXdata[764]), .Z(ofifoDataN[764]));
Q_AN02 U8781 ( .A0(n6720), .A1(shiftedXdata[765]), .Z(ofifoDataN[765]));
Q_AN02 U8782 ( .A0(n6720), .A1(shiftedXdata[766]), .Z(ofifoDataN[766]));
Q_AN02 U8783 ( .A0(n6720), .A1(shiftedXdata[767]), .Z(ofifoDataN[767]));
Q_AD01HF U8784 ( .A0(shiftCount[5]), .B0(writeLen[0]), .S(oFillN[0]), .CO(n1630));
Q_AD02 U8785 ( .CI(n1630), .A0(shiftCount[6]), .A1(shiftCount[7]), .B0(writeLen[1]), .B1(writeLen[2]), .S0(oFillN[1]), .S1(oFillN[2]), .CO(n1629));
Q_AD01HF U8786 ( .A0(writeLen[3]), .B0(n1629), .S(oFillN[3]), .CO(n1628));
Q_AD01HF U8787 ( .A0(ofifoAddr0N[0]), .B0(oFillN[3]), .S(ofifoWptrN[0]), .CO(n1627));
Q_AD01 U8788 ( .CI(oFillN[4]), .A0(ofifoAddr0N[1]), .B0(n1627), .S(ofifoWptrN[1]), .CO(n1626));
Q_AD01HF U8789 ( .A0(ofifoAddr0N[2]), .B0(n1626), .S(ofifoWptrN[2]), .CO(n1625));
Q_AD01HF U8790 ( .A0(ofifoAddr0N[3]), .B0(n1625), .S(ofifoWptrN[3]), .CO(n1624));
Q_AD01HF U8791 ( .A0(ofifoAddr0N[4]), .B0(n1624), .S(ofifoWptrN[4]), .CO(n1623));
Q_AD01HF U8792 ( .A0(ofifoAddr0N[5]), .B0(n1623), .S(ofifoWptrN[5]), .CO(n1622));
Q_AD01HF U8793 ( .A0(ofifoAddr0N[6]), .B0(n1622), .S(ofifoWptrN[6]), .CO(n1621));
Q_AD01HF U8794 ( .A0(ofifoAddr0N[7]), .B0(n1621), .S(ofifoWptrN[7]), .CO(n1620));
Q_AD01HF U8795 ( .A0(ofifoAddr0N[8]), .B0(n1620), .S(ofifoWptrN[8]), .CO(n1619));
Q_AD01HF U8796 ( .A0(ofifoAddr0N[9]), .B0(n1619), .S(ofifoWptrN[9]), .CO(n1618));
Q_AD01HF U8797 ( .A0(ofifoAddr0N[10]), .B0(n1618), .S(ofifoWptrN[10]), .CO(n1617));
Q_AD01HF U8798 ( .A0(ofifoAddr0N[11]), .B0(n1617), .S(ofifoWptrN[11]), .CO(n1616));
Q_AD01HF U8799 ( .A0(ofifoAddr0N[12]), .B0(n1616), .S(ofifoWptrN[12]), .CO(n1615));
Q_AD01HF U8800 ( .A0(ofifoAddr0N[13]), .B0(n1615), .S(ofifoWptrN[13]), .CO(n1614));
Q_XOR2 U8801 ( .A0(ofifoAddr0N[14]), .A1(n1614), .Z(ofifoWptrN[14]));
Q_FDP0 \rLen_REG[17] ( .CK(ackClk), .D(ackLen[17]), .Q(rLen[17]), .QN( ));
Q_FDP0 \rLen_REG[16] ( .CK(ackClk), .D(ackLen[16]), .Q(rLen[16]), .QN( ));
Q_FDP0 \rLen_REG[15] ( .CK(ackClk), .D(ackLen[15]), .Q(rLen[15]), .QN( ));
Q_FDP0 \rLen_REG[14] ( .CK(ackClk), .D(ackLen[14]), .Q(rLen[14]), .QN( ));
Q_FDP0 \rLen_REG[13] ( .CK(ackClk), .D(ackLen[13]), .Q(rLen[13]), .QN( ));
Q_FDP0 \rLen_REG[12] ( .CK(ackClk), .D(ackLen[12]), .Q(rLen[12]), .QN( ));
Q_FDP0 \rLen_REG[11] ( .CK(ackClk), .D(ackLen[11]), .Q(rLen[11]), .QN( ));
Q_FDP0 \rLen_REG[10] ( .CK(ackClk), .D(ackLen[10]), .Q(rLen[10]), .QN( ));
Q_FDP0 \rLen_REG[9] ( .CK(ackClk), .D(ackLen[9]), .Q(rLen[9]), .QN( ));
Q_FDP0 \rLen_REG[8] ( .CK(ackClk), .D(ackLen[8]), .Q(rLen[8]), .QN( ));
Q_FDP0 \rLen_REG[7] ( .CK(ackClk), .D(ackLen[7]), .Q(rLen[7]), .QN( ));
Q_FDP0 \rLen_REG[6] ( .CK(ackClk), .D(ackLen[6]), .Q(rLen[6]), .QN( ));
Q_FDP0 \rLen_REG[5] ( .CK(ackClk), .D(ackLen[5]), .Q(rLen[5]), .QN( ));
Q_FDP0 \rLen_REG[4] ( .CK(ackClk), .D(ackLen[4]), .Q(rLen[4]), .QN( ));
Q_FDP0 \rLen_REG[3] ( .CK(ackClk), .D(ackLen[3]), .Q(rLen[3]), .QN( ));
Q_FDP0 \rLen_REG[2] ( .CK(ackClk), .D(ackLen[2]), .Q(rLen[2]), .QN( ));
Q_FDP0 \rLen_REG[1] ( .CK(ackClk), .D(ackLen[1]), .Q(rLen[1]), .QN( ));
Q_FDP0 \rLen_REG[0] ( .CK(ackClk), .D(ackLen[0]), .Q(rLen[0]), .QN( ));
Q_FDP0 wSync_REG  ( .CK(ackClk), .D(n1613), .Q(wSync), .QN(n1613));
Q_INV U8821 ( .A(svGFbusy1), .Z(LBempty));
Q_OR02 U8822 ( .A0(svGFbusy1), .A1(svGFbusy2), .Z(n1612));
Q_BUFZP U8823 ( .OE(n1612), .A(n1572), .Z(xc_top.svGFbusy));
Q_BUFZP U8824 ( .OE(GFfull), .A(n1572), .Z(xc_top.GFGBfull));
Q_BUFZP U8825 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[11]));
Q_BUFZP U8826 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[10]));
Q_BUFZP U8827 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[9]));
Q_BUFZP U8828 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[8]));
Q_BUFZP U8829 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[7]));
Q_BUFZP U8830 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[6]));
Q_BUFZP U8831 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[5]));
Q_BUFZP U8832 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[4]));
Q_BUFZP U8833 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[3]));
Q_BUFZP U8834 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[2]));
Q_BUFZP U8835 ( .OE(GFtsAdd), .A(n1611), .Z(GFlen[1]));
Q_BUFZP U8836 ( .OE(GFtsAdd), .A(n1572), .Z(GFlen[0]));
Q_BUFZP U8837 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[19]));
Q_BUFZP U8838 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[18]));
Q_BUFZP U8839 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[17]));
Q_BUFZP U8840 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[16]));
Q_BUFZP U8841 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[15]));
Q_BUFZP U8842 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[14]));
Q_BUFZP U8843 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[13]));
Q_BUFZP U8844 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[12]));
Q_BUFZP U8845 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[11]));
Q_BUFZP U8846 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[10]));
Q_BUFZP U8847 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[9]));
Q_BUFZP U8848 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[8]));
Q_BUFZP U8849 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[7]));
Q_BUFZP U8850 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[6]));
Q_BUFZP U8851 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[5]));
Q_BUFZP U8852 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[4]));
Q_BUFZP U8853 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[3]));
Q_BUFZP U8854 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[2]));
Q_BUFZP U8855 ( .OE(GFtsAdd), .A(n1572), .Z(GFcbid[1]));
Q_BUFZP U8856 ( .OE(GFtsAdd), .A(n1611), .Z(GFcbid[0]));
Q_BUFZP U8857 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[31]));
Q_BUFZP U8858 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[30]));
Q_BUFZP U8859 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[29]));
Q_BUFZP U8860 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[28]));
Q_BUFZP U8861 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[27]));
Q_BUFZP U8862 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[26]));
Q_BUFZP U8863 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[25]));
Q_BUFZP U8864 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[24]));
Q_BUFZP U8865 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[23]));
Q_BUFZP U8866 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[22]));
Q_BUFZP U8867 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[21]));
Q_BUFZP U8868 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[20]));
Q_BUFZP U8869 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[19]));
Q_BUFZP U8870 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[18]));
Q_BUFZP U8871 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[17]));
Q_BUFZP U8872 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[16]));
Q_BUFZP U8873 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[15]));
Q_BUFZP U8874 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[14]));
Q_BUFZP U8875 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[13]));
Q_BUFZP U8876 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[12]));
Q_BUFZP U8877 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[11]));
Q_BUFZP U8878 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[10]));
Q_BUFZP U8879 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[9]));
Q_BUFZP U8880 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[8]));
Q_BUFZP U8881 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[7]));
Q_BUFZP U8882 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[6]));
Q_BUFZP U8883 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[5]));
Q_BUFZP U8884 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[4]));
Q_BUFZP U8885 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[3]));
Q_BUFZP U8886 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[2]));
Q_BUFZP U8887 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[1]));
Q_BUFZP U8888 ( .OE(GFtsAdd), .A(n1611), .Z(GFidata[0]));
Q_BUFZN U8889 ( .OE(n3670), .A(n1572), .Z(xc_top.GFAck));
Q_RDN U8890 ( .Z(GFcbid[19]));
Q_RDN U8891 ( .Z(GFcbid[18]));
Q_RDN U8892 ( .Z(GFcbid[17]));
Q_RDN U8893 ( .Z(GFcbid[16]));
Q_RDN U8894 ( .Z(GFcbid[15]));
Q_RDN U8895 ( .Z(GFcbid[14]));
Q_RDN U8896 ( .Z(GFcbid[13]));
Q_RDN U8897 ( .Z(GFcbid[12]));
Q_RDN U8898 ( .Z(GFcbid[11]));
Q_RDN U8899 ( .Z(GFcbid[10]));
Q_RDN U8900 ( .Z(GFcbid[9]));
Q_RDN U8901 ( .Z(GFcbid[8]));
Q_RDN U8902 ( .Z(GFcbid[7]));
Q_RDN U8903 ( .Z(GFcbid[6]));
Q_RDN U8904 ( .Z(GFcbid[5]));
Q_RDN U8905 ( .Z(GFcbid[4]));
Q_RDN U8906 ( .Z(GFcbid[3]));
Q_RDN U8907 ( .Z(GFcbid[2]));
Q_RDN U8908 ( .Z(GFcbid[1]));
Q_RDN U8909 ( .Z(GFcbid[0]));
Q_RDN U8910 ( .Z(GFlen[11]));
Q_RDN U8911 ( .Z(GFlen[10]));
Q_RDN U8912 ( .Z(GFlen[9]));
Q_RDN U8913 ( .Z(GFlen[8]));
Q_RDN U8914 ( .Z(GFlen[7]));
Q_RDN U8915 ( .Z(GFlen[6]));
Q_RDN U8916 ( .Z(GFlen[5]));
Q_RDN U8917 ( .Z(GFlen[4]));
Q_RDN U8918 ( .Z(GFlen[3]));
Q_RDN U8919 ( .Z(GFlen[2]));
Q_RDN U8920 ( .Z(GFlen[1]));
Q_RDN U8921 ( .Z(GFlen[0]));
Q_RDN U8922 ( .Z(GFidata[511]));
Q_RDN U8923 ( .Z(GFidata[510]));
Q_RDN U8924 ( .Z(GFidata[509]));
Q_RDN U8925 ( .Z(GFidata[508]));
Q_RDN U8926 ( .Z(GFidata[507]));
Q_RDN U8927 ( .Z(GFidata[506]));
Q_RDN U8928 ( .Z(GFidata[505]));
Q_RDN U8929 ( .Z(GFidata[504]));
Q_RDN U8930 ( .Z(GFidata[503]));
Q_RDN U8931 ( .Z(GFidata[502]));
Q_RDN U8932 ( .Z(GFidata[501]));
Q_RDN U8933 ( .Z(GFidata[500]));
Q_RDN U8934 ( .Z(GFidata[499]));
Q_RDN U8935 ( .Z(GFidata[498]));
Q_RDN U8936 ( .Z(GFidata[497]));
Q_RDN U8937 ( .Z(GFidata[496]));
Q_RDN U8938 ( .Z(GFidata[495]));
Q_RDN U8939 ( .Z(GFidata[494]));
Q_RDN U8940 ( .Z(GFidata[493]));
Q_RDN U8941 ( .Z(GFidata[492]));
Q_RDN U8942 ( .Z(GFidata[491]));
Q_RDN U8943 ( .Z(GFidata[490]));
Q_RDN U8944 ( .Z(GFidata[489]));
Q_RDN U8945 ( .Z(GFidata[488]));
Q_RDN U8946 ( .Z(GFidata[487]));
Q_RDN U8947 ( .Z(GFidata[486]));
Q_RDN U8948 ( .Z(GFidata[485]));
Q_RDN U8949 ( .Z(GFidata[484]));
Q_RDN U8950 ( .Z(GFidata[483]));
Q_RDN U8951 ( .Z(GFidata[482]));
Q_RDN U8952 ( .Z(GFidata[481]));
Q_RDN U8953 ( .Z(GFidata[480]));
Q_RDN U8954 ( .Z(GFidata[479]));
Q_RDN U8955 ( .Z(GFidata[478]));
Q_RDN U8956 ( .Z(GFidata[477]));
Q_RDN U8957 ( .Z(GFidata[476]));
Q_RDN U8958 ( .Z(GFidata[475]));
Q_RDN U8959 ( .Z(GFidata[474]));
Q_RDN U8960 ( .Z(GFidata[473]));
Q_RDN U8961 ( .Z(GFidata[472]));
Q_RDN U8962 ( .Z(GFidata[471]));
Q_RDN U8963 ( .Z(GFidata[470]));
Q_RDN U8964 ( .Z(GFidata[469]));
Q_RDN U8965 ( .Z(GFidata[468]));
Q_RDN U8966 ( .Z(GFidata[467]));
Q_RDN U8967 ( .Z(GFidata[466]));
Q_RDN U8968 ( .Z(GFidata[465]));
Q_RDN U8969 ( .Z(GFidata[464]));
Q_RDN U8970 ( .Z(GFidata[463]));
Q_RDN U8971 ( .Z(GFidata[462]));
Q_RDN U8972 ( .Z(GFidata[461]));
Q_RDN U8973 ( .Z(GFidata[460]));
Q_RDN U8974 ( .Z(GFidata[459]));
Q_RDN U8975 ( .Z(GFidata[458]));
Q_RDN U8976 ( .Z(GFidata[457]));
Q_RDN U8977 ( .Z(GFidata[456]));
Q_RDN U8978 ( .Z(GFidata[455]));
Q_RDN U8979 ( .Z(GFidata[454]));
Q_RDN U8980 ( .Z(GFidata[453]));
Q_RDN U8981 ( .Z(GFidata[452]));
Q_RDN U8982 ( .Z(GFidata[451]));
Q_RDN U8983 ( .Z(GFidata[450]));
Q_RDN U8984 ( .Z(GFidata[449]));
Q_RDN U8985 ( .Z(GFidata[448]));
Q_RDN U8986 ( .Z(GFidata[447]));
Q_RDN U8987 ( .Z(GFidata[446]));
Q_RDN U8988 ( .Z(GFidata[445]));
Q_RDN U8989 ( .Z(GFidata[444]));
Q_RDN U8990 ( .Z(GFidata[443]));
Q_RDN U8991 ( .Z(GFidata[442]));
Q_RDN U8992 ( .Z(GFidata[441]));
Q_RDN U8993 ( .Z(GFidata[440]));
Q_RDN U8994 ( .Z(GFidata[439]));
Q_RDN U8995 ( .Z(GFidata[438]));
Q_RDN U8996 ( .Z(GFidata[437]));
Q_RDN U8997 ( .Z(GFidata[436]));
Q_RDN U8998 ( .Z(GFidata[435]));
Q_RDN U8999 ( .Z(GFidata[434]));
Q_RDN U9000 ( .Z(GFidata[433]));
Q_RDN U9001 ( .Z(GFidata[432]));
Q_RDN U9002 ( .Z(GFidata[431]));
Q_RDN U9003 ( .Z(GFidata[430]));
Q_RDN U9004 ( .Z(GFidata[429]));
Q_RDN U9005 ( .Z(GFidata[428]));
Q_RDN U9006 ( .Z(GFidata[427]));
Q_RDN U9007 ( .Z(GFidata[426]));
Q_RDN U9008 ( .Z(GFidata[425]));
Q_RDN U9009 ( .Z(GFidata[424]));
Q_RDN U9010 ( .Z(GFidata[423]));
Q_RDN U9011 ( .Z(GFidata[422]));
Q_RDN U9012 ( .Z(GFidata[421]));
Q_RDN U9013 ( .Z(GFidata[420]));
Q_RDN U9014 ( .Z(GFidata[419]));
Q_RDN U9015 ( .Z(GFidata[418]));
Q_RDN U9016 ( .Z(GFidata[417]));
Q_RDN U9017 ( .Z(GFidata[416]));
Q_RDN U9018 ( .Z(GFidata[415]));
Q_RDN U9019 ( .Z(GFidata[414]));
Q_RDN U9020 ( .Z(GFidata[413]));
Q_RDN U9021 ( .Z(GFidata[412]));
Q_RDN U9022 ( .Z(GFidata[411]));
Q_RDN U9023 ( .Z(GFidata[410]));
Q_RDN U9024 ( .Z(GFidata[409]));
Q_RDN U9025 ( .Z(GFidata[408]));
Q_RDN U9026 ( .Z(GFidata[407]));
Q_RDN U9027 ( .Z(GFidata[406]));
Q_RDN U9028 ( .Z(GFidata[405]));
Q_RDN U9029 ( .Z(GFidata[404]));
Q_RDN U9030 ( .Z(GFidata[403]));
Q_RDN U9031 ( .Z(GFidata[402]));
Q_RDN U9032 ( .Z(GFidata[401]));
Q_RDN U9033 ( .Z(GFidata[400]));
Q_RDN U9034 ( .Z(GFidata[399]));
Q_RDN U9035 ( .Z(GFidata[398]));
Q_RDN U9036 ( .Z(GFidata[397]));
Q_RDN U9037 ( .Z(GFidata[396]));
Q_RDN U9038 ( .Z(GFidata[395]));
Q_RDN U9039 ( .Z(GFidata[394]));
Q_RDN U9040 ( .Z(GFidata[393]));
Q_RDN U9041 ( .Z(GFidata[392]));
Q_RDN U9042 ( .Z(GFidata[391]));
Q_RDN U9043 ( .Z(GFidata[390]));
Q_RDN U9044 ( .Z(GFidata[389]));
Q_RDN U9045 ( .Z(GFidata[388]));
Q_RDN U9046 ( .Z(GFidata[387]));
Q_RDN U9047 ( .Z(GFidata[386]));
Q_RDN U9048 ( .Z(GFidata[385]));
Q_RDN U9049 ( .Z(GFidata[384]));
Q_RDN U9050 ( .Z(GFidata[383]));
Q_RDN U9051 ( .Z(GFidata[382]));
Q_RDN U9052 ( .Z(GFidata[381]));
Q_RDN U9053 ( .Z(GFidata[380]));
Q_RDN U9054 ( .Z(GFidata[379]));
Q_RDN U9055 ( .Z(GFidata[378]));
Q_RDN U9056 ( .Z(GFidata[377]));
Q_RDN U9057 ( .Z(GFidata[376]));
Q_RDN U9058 ( .Z(GFidata[375]));
Q_RDN U9059 ( .Z(GFidata[374]));
Q_RDN U9060 ( .Z(GFidata[373]));
Q_RDN U9061 ( .Z(GFidata[372]));
Q_RDN U9062 ( .Z(GFidata[371]));
Q_RDN U9063 ( .Z(GFidata[370]));
Q_RDN U9064 ( .Z(GFidata[369]));
Q_RDN U9065 ( .Z(GFidata[368]));
Q_RDN U9066 ( .Z(GFidata[367]));
Q_RDN U9067 ( .Z(GFidata[366]));
Q_RDN U9068 ( .Z(GFidata[365]));
Q_RDN U9069 ( .Z(GFidata[364]));
Q_RDN U9070 ( .Z(GFidata[363]));
Q_RDN U9071 ( .Z(GFidata[362]));
Q_RDN U9072 ( .Z(GFidata[361]));
Q_RDN U9073 ( .Z(GFidata[360]));
Q_RDN U9074 ( .Z(GFidata[359]));
Q_RDN U9075 ( .Z(GFidata[358]));
Q_RDN U9076 ( .Z(GFidata[357]));
Q_RDN U9077 ( .Z(GFidata[356]));
Q_RDN U9078 ( .Z(GFidata[355]));
Q_RDN U9079 ( .Z(GFidata[354]));
Q_RDN U9080 ( .Z(GFidata[353]));
Q_RDN U9081 ( .Z(GFidata[352]));
Q_RDN U9082 ( .Z(GFidata[351]));
Q_RDN U9083 ( .Z(GFidata[350]));
Q_RDN U9084 ( .Z(GFidata[349]));
Q_RDN U9085 ( .Z(GFidata[348]));
Q_RDN U9086 ( .Z(GFidata[347]));
Q_RDN U9087 ( .Z(GFidata[346]));
Q_RDN U9088 ( .Z(GFidata[345]));
Q_RDN U9089 ( .Z(GFidata[344]));
Q_RDN U9090 ( .Z(GFidata[343]));
Q_RDN U9091 ( .Z(GFidata[342]));
Q_RDN U9092 ( .Z(GFidata[341]));
Q_RDN U9093 ( .Z(GFidata[340]));
Q_RDN U9094 ( .Z(GFidata[339]));
Q_RDN U9095 ( .Z(GFidata[338]));
Q_RDN U9096 ( .Z(GFidata[337]));
Q_RDN U9097 ( .Z(GFidata[336]));
Q_RDN U9098 ( .Z(GFidata[335]));
Q_RDN U9099 ( .Z(GFidata[334]));
Q_RDN U9100 ( .Z(GFidata[333]));
Q_RDN U9101 ( .Z(GFidata[332]));
Q_RDN U9102 ( .Z(GFidata[331]));
Q_RDN U9103 ( .Z(GFidata[330]));
Q_RDN U9104 ( .Z(GFidata[329]));
Q_RDN U9105 ( .Z(GFidata[328]));
Q_RDN U9106 ( .Z(GFidata[327]));
Q_RDN U9107 ( .Z(GFidata[326]));
Q_RDN U9108 ( .Z(GFidata[325]));
Q_RDN U9109 ( .Z(GFidata[324]));
Q_RDN U9110 ( .Z(GFidata[323]));
Q_RDN U9111 ( .Z(GFidata[322]));
Q_RDN U9112 ( .Z(GFidata[321]));
Q_RDN U9113 ( .Z(GFidata[320]));
Q_RDN U9114 ( .Z(GFidata[319]));
Q_RDN U9115 ( .Z(GFidata[318]));
Q_RDN U9116 ( .Z(GFidata[317]));
Q_RDN U9117 ( .Z(GFidata[316]));
Q_RDN U9118 ( .Z(GFidata[315]));
Q_RDN U9119 ( .Z(GFidata[314]));
Q_RDN U9120 ( .Z(GFidata[313]));
Q_RDN U9121 ( .Z(GFidata[312]));
Q_RDN U9122 ( .Z(GFidata[311]));
Q_RDN U9123 ( .Z(GFidata[310]));
Q_RDN U9124 ( .Z(GFidata[309]));
Q_RDN U9125 ( .Z(GFidata[308]));
Q_RDN U9126 ( .Z(GFidata[307]));
Q_RDN U9127 ( .Z(GFidata[306]));
Q_RDN U9128 ( .Z(GFidata[305]));
Q_RDN U9129 ( .Z(GFidata[304]));
Q_RDN U9130 ( .Z(GFidata[303]));
Q_RDN U9131 ( .Z(GFidata[302]));
Q_RDN U9132 ( .Z(GFidata[301]));
Q_RDN U9133 ( .Z(GFidata[300]));
Q_RDN U9134 ( .Z(GFidata[299]));
Q_RDN U9135 ( .Z(GFidata[298]));
Q_RDN U9136 ( .Z(GFidata[297]));
Q_RDN U9137 ( .Z(GFidata[296]));
Q_RDN U9138 ( .Z(GFidata[295]));
Q_RDN U9139 ( .Z(GFidata[294]));
Q_RDN U9140 ( .Z(GFidata[293]));
Q_RDN U9141 ( .Z(GFidata[292]));
Q_RDN U9142 ( .Z(GFidata[291]));
Q_RDN U9143 ( .Z(GFidata[290]));
Q_RDN U9144 ( .Z(GFidata[289]));
Q_RDN U9145 ( .Z(GFidata[288]));
Q_RDN U9146 ( .Z(GFidata[287]));
Q_RDN U9147 ( .Z(GFidata[286]));
Q_RDN U9148 ( .Z(GFidata[285]));
Q_RDN U9149 ( .Z(GFidata[284]));
Q_RDN U9150 ( .Z(GFidata[283]));
Q_RDN U9151 ( .Z(GFidata[282]));
Q_RDN U9152 ( .Z(GFidata[281]));
Q_RDN U9153 ( .Z(GFidata[280]));
Q_RDN U9154 ( .Z(GFidata[279]));
Q_RDN U9155 ( .Z(GFidata[278]));
Q_RDN U9156 ( .Z(GFidata[277]));
Q_RDN U9157 ( .Z(GFidata[276]));
Q_RDN U9158 ( .Z(GFidata[275]));
Q_RDN U9159 ( .Z(GFidata[274]));
Q_RDN U9160 ( .Z(GFidata[273]));
Q_RDN U9161 ( .Z(GFidata[272]));
Q_RDN U9162 ( .Z(GFidata[271]));
Q_RDN U9163 ( .Z(GFidata[270]));
Q_RDN U9164 ( .Z(GFidata[269]));
Q_RDN U9165 ( .Z(GFidata[268]));
Q_RDN U9166 ( .Z(GFidata[267]));
Q_RDN U9167 ( .Z(GFidata[266]));
Q_RDN U9168 ( .Z(GFidata[265]));
Q_RDN U9169 ( .Z(GFidata[264]));
Q_RDN U9170 ( .Z(GFidata[263]));
Q_RDN U9171 ( .Z(GFidata[262]));
Q_RDN U9172 ( .Z(GFidata[261]));
Q_RDN U9173 ( .Z(GFidata[260]));
Q_RDN U9174 ( .Z(GFidata[259]));
Q_RDN U9175 ( .Z(GFidata[258]));
Q_RDN U9176 ( .Z(GFidata[257]));
Q_RDN U9177 ( .Z(GFidata[256]));
Q_RDN U9178 ( .Z(GFidata[255]));
Q_RDN U9179 ( .Z(GFidata[254]));
Q_RDN U9180 ( .Z(GFidata[253]));
Q_RDN U9181 ( .Z(GFidata[252]));
Q_RDN U9182 ( .Z(GFidata[251]));
Q_RDN U9183 ( .Z(GFidata[250]));
Q_RDN U9184 ( .Z(GFidata[249]));
Q_RDN U9185 ( .Z(GFidata[248]));
Q_RDN U9186 ( .Z(GFidata[247]));
Q_RDN U9187 ( .Z(GFidata[246]));
Q_RDN U9188 ( .Z(GFidata[245]));
Q_RDN U9189 ( .Z(GFidata[244]));
Q_RDN U9190 ( .Z(GFidata[243]));
Q_RDN U9191 ( .Z(GFidata[242]));
Q_RDN U9192 ( .Z(GFidata[241]));
Q_RDN U9193 ( .Z(GFidata[240]));
Q_RDN U9194 ( .Z(GFidata[239]));
Q_RDN U9195 ( .Z(GFidata[238]));
Q_RDN U9196 ( .Z(GFidata[237]));
Q_RDN U9197 ( .Z(GFidata[236]));
Q_RDN U9198 ( .Z(GFidata[235]));
Q_RDN U9199 ( .Z(GFidata[234]));
Q_RDN U9200 ( .Z(GFidata[233]));
Q_RDN U9201 ( .Z(GFidata[232]));
Q_RDN U9202 ( .Z(GFidata[231]));
Q_RDN U9203 ( .Z(GFidata[230]));
Q_RDN U9204 ( .Z(GFidata[229]));
Q_RDN U9205 ( .Z(GFidata[228]));
Q_RDN U9206 ( .Z(GFidata[227]));
Q_RDN U9207 ( .Z(GFidata[226]));
Q_RDN U9208 ( .Z(GFidata[225]));
Q_RDN U9209 ( .Z(GFidata[224]));
Q_RDN U9210 ( .Z(GFidata[223]));
Q_RDN U9211 ( .Z(GFidata[222]));
Q_RDN U9212 ( .Z(GFidata[221]));
Q_RDN U9213 ( .Z(GFidata[220]));
Q_RDN U9214 ( .Z(GFidata[219]));
Q_RDN U9215 ( .Z(GFidata[218]));
Q_RDN U9216 ( .Z(GFidata[217]));
Q_RDN U9217 ( .Z(GFidata[216]));
Q_RDN U9218 ( .Z(GFidata[215]));
Q_RDN U9219 ( .Z(GFidata[214]));
Q_RDN U9220 ( .Z(GFidata[213]));
Q_RDN U9221 ( .Z(GFidata[212]));
Q_RDN U9222 ( .Z(GFidata[211]));
Q_RDN U9223 ( .Z(GFidata[210]));
Q_RDN U9224 ( .Z(GFidata[209]));
Q_RDN U9225 ( .Z(GFidata[208]));
Q_RDN U9226 ( .Z(GFidata[207]));
Q_RDN U9227 ( .Z(GFidata[206]));
Q_RDN U9228 ( .Z(GFidata[205]));
Q_RDN U9229 ( .Z(GFidata[204]));
Q_RDN U9230 ( .Z(GFidata[203]));
Q_RDN U9231 ( .Z(GFidata[202]));
Q_RDN U9232 ( .Z(GFidata[201]));
Q_RDN U9233 ( .Z(GFidata[200]));
Q_RDN U9234 ( .Z(GFidata[199]));
Q_RDN U9235 ( .Z(GFidata[198]));
Q_RDN U9236 ( .Z(GFidata[197]));
Q_RDN U9237 ( .Z(GFidata[196]));
Q_RDN U9238 ( .Z(GFidata[195]));
Q_RDN U9239 ( .Z(GFidata[194]));
Q_RDN U9240 ( .Z(GFidata[193]));
Q_RDN U9241 ( .Z(GFidata[192]));
Q_RDN U9242 ( .Z(GFidata[191]));
Q_RDN U9243 ( .Z(GFidata[190]));
Q_RDN U9244 ( .Z(GFidata[189]));
Q_RDN U9245 ( .Z(GFidata[188]));
Q_RDN U9246 ( .Z(GFidata[187]));
Q_RDN U9247 ( .Z(GFidata[186]));
Q_RDN U9248 ( .Z(GFidata[185]));
Q_RDN U9249 ( .Z(GFidata[184]));
Q_RDN U9250 ( .Z(GFidata[183]));
Q_RDN U9251 ( .Z(GFidata[182]));
Q_RDN U9252 ( .Z(GFidata[181]));
Q_RDN U9253 ( .Z(GFidata[180]));
Q_RDN U9254 ( .Z(GFidata[179]));
Q_RDN U9255 ( .Z(GFidata[178]));
Q_RDN U9256 ( .Z(GFidata[177]));
Q_RDN U9257 ( .Z(GFidata[176]));
Q_RDN U9258 ( .Z(GFidata[175]));
Q_RDN U9259 ( .Z(GFidata[174]));
Q_RDN U9260 ( .Z(GFidata[173]));
Q_RDN U9261 ( .Z(GFidata[172]));
Q_RDN U9262 ( .Z(GFidata[171]));
Q_RDN U9263 ( .Z(GFidata[170]));
Q_RDN U9264 ( .Z(GFidata[169]));
Q_RDN U9265 ( .Z(GFidata[168]));
Q_RDN U9266 ( .Z(GFidata[167]));
Q_RDN U9267 ( .Z(GFidata[166]));
Q_RDN U9268 ( .Z(GFidata[165]));
Q_RDN U9269 ( .Z(GFidata[164]));
Q_RDN U9270 ( .Z(GFidata[163]));
Q_RDN U9271 ( .Z(GFidata[162]));
Q_RDN U9272 ( .Z(GFidata[161]));
Q_RDN U9273 ( .Z(GFidata[160]));
Q_RDN U9274 ( .Z(GFidata[159]));
Q_RDN U9275 ( .Z(GFidata[158]));
Q_RDN U9276 ( .Z(GFidata[157]));
Q_RDN U9277 ( .Z(GFidata[156]));
Q_RDN U9278 ( .Z(GFidata[155]));
Q_RDN U9279 ( .Z(GFidata[154]));
Q_RDN U9280 ( .Z(GFidata[153]));
Q_RDN U9281 ( .Z(GFidata[152]));
Q_RDN U9282 ( .Z(GFidata[151]));
Q_RDN U9283 ( .Z(GFidata[150]));
Q_RDN U9284 ( .Z(GFidata[149]));
Q_RDN U9285 ( .Z(GFidata[148]));
Q_RDN U9286 ( .Z(GFidata[147]));
Q_RDN U9287 ( .Z(GFidata[146]));
Q_RDN U9288 ( .Z(GFidata[145]));
Q_RDN U9289 ( .Z(GFidata[144]));
Q_RDN U9290 ( .Z(GFidata[143]));
Q_RDN U9291 ( .Z(GFidata[142]));
Q_RDN U9292 ( .Z(GFidata[141]));
Q_RDN U9293 ( .Z(GFidata[140]));
Q_RDN U9294 ( .Z(GFidata[139]));
Q_RDN U9295 ( .Z(GFidata[138]));
Q_RDN U9296 ( .Z(GFidata[137]));
Q_RDN U9297 ( .Z(GFidata[136]));
Q_RDN U9298 ( .Z(GFidata[135]));
Q_RDN U9299 ( .Z(GFidata[134]));
Q_RDN U9300 ( .Z(GFidata[133]));
Q_RDN U9301 ( .Z(GFidata[132]));
Q_RDN U9302 ( .Z(GFidata[131]));
Q_RDN U9303 ( .Z(GFidata[130]));
Q_RDN U9304 ( .Z(GFidata[129]));
Q_RDN U9305 ( .Z(GFidata[128]));
Q_RDN U9306 ( .Z(GFidata[127]));
Q_RDN U9307 ( .Z(GFidata[126]));
Q_RDN U9308 ( .Z(GFidata[125]));
Q_RDN U9309 ( .Z(GFidata[124]));
Q_RDN U9310 ( .Z(GFidata[123]));
Q_RDN U9311 ( .Z(GFidata[122]));
Q_RDN U9312 ( .Z(GFidata[121]));
Q_RDN U9313 ( .Z(GFidata[120]));
Q_RDN U9314 ( .Z(GFidata[119]));
Q_RDN U9315 ( .Z(GFidata[118]));
Q_RDN U9316 ( .Z(GFidata[117]));
Q_RDN U9317 ( .Z(GFidata[116]));
Q_RDN U9318 ( .Z(GFidata[115]));
Q_RDN U9319 ( .Z(GFidata[114]));
Q_RDN U9320 ( .Z(GFidata[113]));
Q_RDN U9321 ( .Z(GFidata[112]));
Q_RDN U9322 ( .Z(GFidata[111]));
Q_RDN U9323 ( .Z(GFidata[110]));
Q_RDN U9324 ( .Z(GFidata[109]));
Q_RDN U9325 ( .Z(GFidata[108]));
Q_RDN U9326 ( .Z(GFidata[107]));
Q_RDN U9327 ( .Z(GFidata[106]));
Q_RDN U9328 ( .Z(GFidata[105]));
Q_RDN U9329 ( .Z(GFidata[104]));
Q_RDN U9330 ( .Z(GFidata[103]));
Q_RDN U9331 ( .Z(GFidata[102]));
Q_RDN U9332 ( .Z(GFidata[101]));
Q_RDN U9333 ( .Z(GFidata[100]));
Q_RDN U9334 ( .Z(GFidata[99]));
Q_RDN U9335 ( .Z(GFidata[98]));
Q_RDN U9336 ( .Z(GFidata[97]));
Q_RDN U9337 ( .Z(GFidata[96]));
Q_RDN U9338 ( .Z(GFidata[95]));
Q_RDN U9339 ( .Z(GFidata[94]));
Q_RDN U9340 ( .Z(GFidata[93]));
Q_RDN U9341 ( .Z(GFidata[92]));
Q_RDN U9342 ( .Z(GFidata[91]));
Q_RDN U9343 ( .Z(GFidata[90]));
Q_RDN U9344 ( .Z(GFidata[89]));
Q_RDN U9345 ( .Z(GFidata[88]));
Q_RDN U9346 ( .Z(GFidata[87]));
Q_RDN U9347 ( .Z(GFidata[86]));
Q_RDN U9348 ( .Z(GFidata[85]));
Q_RDN U9349 ( .Z(GFidata[84]));
Q_RDN U9350 ( .Z(GFidata[83]));
Q_RDN U9351 ( .Z(GFidata[82]));
Q_RDN U9352 ( .Z(GFidata[81]));
Q_RDN U9353 ( .Z(GFidata[80]));
Q_RDN U9354 ( .Z(GFidata[79]));
Q_RDN U9355 ( .Z(GFidata[78]));
Q_RDN U9356 ( .Z(GFidata[77]));
Q_RDN U9357 ( .Z(GFidata[76]));
Q_RDN U9358 ( .Z(GFidata[75]));
Q_RDN U9359 ( .Z(GFidata[74]));
Q_RDN U9360 ( .Z(GFidata[73]));
Q_RDN U9361 ( .Z(GFidata[72]));
Q_RDN U9362 ( .Z(GFidata[71]));
Q_RDN U9363 ( .Z(GFidata[70]));
Q_RDN U9364 ( .Z(GFidata[69]));
Q_RDN U9365 ( .Z(GFidata[68]));
Q_RDN U9366 ( .Z(GFidata[67]));
Q_RDN U9367 ( .Z(GFidata[66]));
Q_RDN U9368 ( .Z(GFidata[65]));
Q_RDN U9369 ( .Z(GFidata[64]));
Q_RDN U9370 ( .Z(GFidata[63]));
Q_RDN U9371 ( .Z(GFidata[62]));
Q_RDN U9372 ( .Z(GFidata[61]));
Q_RDN U9373 ( .Z(GFidata[60]));
Q_RDN U9374 ( .Z(GFidata[59]));
Q_RDN U9375 ( .Z(GFidata[58]));
Q_RDN U9376 ( .Z(GFidata[57]));
Q_RDN U9377 ( .Z(GFidata[56]));
Q_RDN U9378 ( .Z(GFidata[55]));
Q_RDN U9379 ( .Z(GFidata[54]));
Q_RDN U9380 ( .Z(GFidata[53]));
Q_RDN U9381 ( .Z(GFidata[52]));
Q_RDN U9382 ( .Z(GFidata[51]));
Q_RDN U9383 ( .Z(GFidata[50]));
Q_RDN U9384 ( .Z(GFidata[49]));
Q_RDN U9385 ( .Z(GFidata[48]));
Q_RDN U9386 ( .Z(GFidata[47]));
Q_RDN U9387 ( .Z(GFidata[46]));
Q_RDN U9388 ( .Z(GFidata[45]));
Q_RDN U9389 ( .Z(GFidata[44]));
Q_RDN U9390 ( .Z(GFidata[43]));
Q_RDN U9391 ( .Z(GFidata[42]));
Q_RDN U9392 ( .Z(GFidata[41]));
Q_RDN U9393 ( .Z(GFidata[40]));
Q_RDN U9394 ( .Z(GFidata[39]));
Q_RDN U9395 ( .Z(GFidata[38]));
Q_RDN U9396 ( .Z(GFidata[37]));
Q_RDN U9397 ( .Z(GFidata[36]));
Q_RDN U9398 ( .Z(GFidata[35]));
Q_RDN U9399 ( .Z(GFidata[34]));
Q_RDN U9400 ( .Z(GFidata[33]));
Q_RDN U9401 ( .Z(GFidata[32]));
Q_RDN U9402 ( .Z(GFidata[31]));
Q_RDN U9403 ( .Z(GFidata[30]));
Q_RDN U9404 ( .Z(GFidata[29]));
Q_RDN U9405 ( .Z(GFidata[28]));
Q_RDN U9406 ( .Z(GFidata[27]));
Q_RDN U9407 ( .Z(GFidata[26]));
Q_RDN U9408 ( .Z(GFidata[25]));
Q_RDN U9409 ( .Z(GFidata[24]));
Q_RDN U9410 ( .Z(GFidata[23]));
Q_RDN U9411 ( .Z(GFidata[22]));
Q_RDN U9412 ( .Z(GFidata[21]));
Q_RDN U9413 ( .Z(GFidata[20]));
Q_RDN U9414 ( .Z(GFidata[19]));
Q_RDN U9415 ( .Z(GFidata[18]));
Q_RDN U9416 ( .Z(GFidata[17]));
Q_RDN U9417 ( .Z(GFidata[16]));
Q_RDN U9418 ( .Z(GFidata[15]));
Q_RDN U9419 ( .Z(GFidata[14]));
Q_RDN U9420 ( .Z(GFidata[13]));
Q_RDN U9421 ( .Z(GFidata[12]));
Q_RDN U9422 ( .Z(GFidata[11]));
Q_RDN U9423 ( .Z(GFidata[10]));
Q_RDN U9424 ( .Z(GFidata[9]));
Q_RDN U9425 ( .Z(GFidata[8]));
Q_RDN U9426 ( .Z(GFidata[7]));
Q_RDN U9427 ( .Z(GFidata[6]));
Q_RDN U9428 ( .Z(GFidata[5]));
Q_RDN U9429 ( .Z(GFidata[4]));
Q_RDN U9430 ( .Z(GFidata[3]));
Q_RDN U9431 ( .Z(GFidata[2]));
Q_RDN U9432 ( .Z(GFidata[1]));
Q_RDN U9433 ( .Z(GFidata[0]));
Q_RDN U9434 ( .Z(LBreq));
Q_RDN U9435 ( .Z(GFtsReq));
Q_AN03 U9436 ( .A0(wLen[17]), .A1(wLen[16]), .A2(wLen[15]), .Z(n1573));
Q_AN03 U9437 ( .A0(wLen[14]), .A1(wLen[13]), .A2(wLen[12]), .Z(n1574));
Q_AN03 U9438 ( .A0(n1574), .A1(wLen[11]), .A2(n1573), .Z(n1582));
Q_OR02 U9439 ( .A0(wLen[8]), .A1(wLen[7]), .Z(n1575));
Q_OR03 U9440 ( .A0(wLen[10]), .A1(wLen[9]), .A2(n1575), .Z(n1576));
Q_OR02 U9441 ( .A0(wLen[4]), .A1(wLen[3]), .Z(n1577));
Q_OR03 U9442 ( .A0(wLen[6]), .A1(wLen[5]), .A2(n1577), .Z(n1578));
Q_OR03 U9443 ( .A0(wLen[2]), .A1(wLen[1]), .A2(wLen[0]), .Z(n1579));
Q_AN02 U9444 ( .A0(n1573), .A1(n1574), .Z(n1580));
Q_OA21 U9445 ( .A0(n1576), .A1(n1578), .B0(n1580), .Z(n1581));
Q_OR03 U9446 ( .A0(wLen[18]), .A1(n1582), .A2(n1581), .Z(n1583));
Q_AO21 U9447 ( .A0(n1580), .A1(n1579), .B0(n1583), .Z(GFfull));
axis_tbcall_BP_1 tbcx ( flushTbc, n1584, flushTbc_x$tbc, n1585);
Q_XOR3 U9449 ( .A0(timeStampPkt[63]), .A1(timeStampPkt[62]), .A2(timeStampPkt[61]), .Z(n1586));
Q_XOR3 U9450 ( .A0(timeStampPkt[60]), .A1(timeStampPkt[59]), .A2(timeStampPkt[58]), .Z(n1587));
Q_XOR3 U9451 ( .A0(timeStampPkt[57]), .A1(timeStampPkt[56]), .A2(n1586), .Z(n1588));
Q_XOR2 U9452 ( .A0(n1587), .A1(n1588), .Z(timeStampPkt[30]));
Q_XOR3 U9453 ( .A0(timeStampPkt[55]), .A1(timeStampPkt[54]), .A2(timeStampPkt[53]), .Z(n1589));
Q_XOR3 U9454 ( .A0(timeStampPkt[52]), .A1(timeStampPkt[51]), .A2(timeStampPkt[50]), .Z(n1590));
Q_XOR3 U9455 ( .A0(timeStampPkt[49]), .A1(timeStampPkt[48]), .A2(n1589), .Z(n1591));
Q_XOR2 U9456 ( .A0(n1590), .A1(n1591), .Z(timeStampPkt[29]));
Q_XOR3 U9457 ( .A0(timeStampPkt[47]), .A1(timeStampPkt[46]), .A2(timeStampPkt[45]), .Z(n1592));
Q_XOR3 U9458 ( .A0(timeStampPkt[44]), .A1(timeStampPkt[43]), .A2(timeStampPkt[42]), .Z(n1593));
Q_XOR3 U9459 ( .A0(timeStampPkt[41]), .A1(timeStampPkt[40]), .A2(n1592), .Z(n1594));
Q_XOR2 U9460 ( .A0(n1593), .A1(n1594), .Z(timeStampPkt[28]));
Q_XOR3 U9461 ( .A0(timeStampPkt[39]), .A1(timeStampPkt[38]), .A2(timeStampPkt[37]), .Z(n1595));
Q_XOR3 U9462 ( .A0(timeStampPkt[36]), .A1(timeStampPkt[35]), .A2(timeStampPkt[34]), .Z(n1596));
Q_XOR3 U9463 ( .A0(timeStampPkt[33]), .A1(timeStampPkt[32]), .A2(n1595), .Z(n1597));
Q_XOR2 U9464 ( .A0(n1596), .A1(n1597), .Z(timeStampPkt[27]));
Q_XOR3 U9465 ( .A0(timeStampPkt[23]), .A1(timeStampPkt[22]), .A2(timeStampPkt[21]), .Z(n1598));
Q_XOR3 U9466 ( .A0(timeStampPkt[20]), .A1(timeStampPkt[19]), .A2(timeStampPkt[18]), .Z(n1599));
Q_XOR3 U9467 ( .A0(timeStampPkt[17]), .A1(timeStampPkt[16]), .A2(n1598), .Z(n1600));
Q_XOR2 U9468 ( .A0(n1599), .A1(n1600), .Z(timeStampPkt[26]));
Q_XOR3 U9469 ( .A0(timeStampPkt[15]), .A1(timeStampPkt[14]), .A2(timeStampPkt[13]), .Z(n1601));
Q_XOR3 U9470 ( .A0(timeStampPkt[12]), .A1(timeStampPkt[11]), .A2(timeStampPkt[10]), .Z(n1602));
Q_XOR3 U9471 ( .A0(timeStampPkt[9]), .A1(timeStampPkt[8]), .A2(n1601), .Z(n1603));
Q_XOR2 U9472 ( .A0(n1602), .A1(n1603), .Z(timeStampPkt[25]));
Q_XOR3 U9473 ( .A0(timeStampPkt[7]), .A1(timeStampPkt[6]), .A2(timeStampPkt[5]), .Z(n1604));
Q_XOR3 U9474 ( .A0(timeStampPkt[4]), .A1(timeStampPkt[3]), .A2(timeStampPkt[2]), .Z(n1605));
Q_XOR3 U9475 ( .A0(timeStampPkt[1]), .A1(timeStampPkt[0]), .A2(n1604), .Z(n1606));
Q_XOR2 U9476 ( .A0(n1605), .A1(n1606), .Z(timeStampPkt[24]));
Q_OR03 U9477 ( .A0(LBfill[3]), .A1(LBfill[2]), .A2(LBfill[1]), .Z(n1607));
Q_OR02 U9478 ( .A0(LBfill[0]), .A1(n1607), .Z(svGFbusy1));
Q_INV U9479 ( .A(LBfill[2]), .Z(n1608));
Q_OR03 U9480 ( .A0(LBfill[3]), .A1(n1608), .A2(LBfill[1]), .Z(n1609));
Q_OR02 U9481 ( .A0(LBfill[0]), .A1(n1609), .Z(n1610));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_INV U9483 ( .A(n6639), .Z(n1570));
Q_INV U9484 ( .A(n6640), .Z(n1569));
`ifdef CBV

reg [255:0] ixc_gfm_ofifo [0:32767];
always @(ofifoAddr0N[14] or ofifoAddr0N[13] or ofifoAddr0N[12] or ofifoAddr0N[11] or ofifoAddr0N[10]
 or ofifoAddr0N[9] or ofifoAddr0N[8] or ofifoAddr0N[7] or ofifoAddr0N[6] or ofifoAddr0N[5] or ofifoAddr0N[4] or ofifoAddr0N[3] or ofifoAddr0N[2]
 or ofifoAddr0N[1] or ofifoAddr0N[0] or ofifoDataN[255] or ofifoDataN[254] or ofifoDataN[253] or ofifoDataN[252] or ofifoDataN[251] or ofifoDataN[250]
 or ofifoDataN[249] or ofifoDataN[248] or ofifoDataN[247] or ofifoDataN[246] or ofifoDataN[245] or ofifoDataN[244] or ofifoDataN[243] or ofifoDataN[242]
 or ofifoDataN[241] or ofifoDataN[240] or ofifoDataN[239] or ofifoDataN[238] or ofifoDataN[237] or ofifoDataN[236] or ofifoDataN[235] or ofifoDataN[234]
 or ofifoDataN[233] or ofifoDataN[232] or ofifoDataN[231] or ofifoDataN[230] or ofifoDataN[229] or ofifoDataN[228] or ofifoDataN[227] or ofifoDataN[226]
 or ofifoDataN[225] or ofifoDataN[224] or ofifoDataN[223] or ofifoDataN[222] or ofifoDataN[221] or ofifoDataN[220] or ofifoDataN[219] or ofifoDataN[218]
 or ofifoDataN[217] or ofifoDataN[216] or ofifoDataN[215] or ofifoDataN[214] or ofifoDataN[213] or ofifoDataN[212] or ofifoDataN[211] or ofifoDataN[210]
 or ofifoDataN[209] or ofifoDataN[208] or ofifoDataN[207] or ofifoDataN[206] or ofifoDataN[205] or ofifoDataN[204] or ofifoDataN[203] or ofifoDataN[202]
 or ofifoDataN[201] or ofifoDataN[200] or ofifoDataN[199] or ofifoDataN[198] or ofifoDataN[197] or ofifoDataN[196] or ofifoDataN[195] or ofifoDataN[194]
 or ofifoDataN[193] or ofifoDataN[192] or ofifoDataN[191] or ofifoDataN[190] or ofifoDataN[189] or ofifoDataN[188] or ofifoDataN[187] or ofifoDataN[186]
 or ofifoDataN[185] or ofifoDataN[184] or ofifoDataN[183] or ofifoDataN[182] or ofifoDataN[181] or ofifoDataN[180] or ofifoDataN[179] or ofifoDataN[178]
 or ofifoDataN[177] or ofifoDataN[176] or ofifoDataN[175] or ofifoDataN[174] or ofifoDataN[173] or ofifoDataN[172] or ofifoDataN[171] or ofifoDataN[170]
 or ofifoDataN[169] or ofifoDataN[168] or ofifoDataN[167] or ofifoDataN[166] or ofifoDataN[165] or ofifoDataN[164] or ofifoDataN[163] or ofifoDataN[162]
 or ofifoDataN[161] or ofifoDataN[160] or ofifoDataN[159] or ofifoDataN[158] or ofifoDataN[157] or ofifoDataN[156] or ofifoDataN[155] or ofifoDataN[154]
 or ofifoDataN[153] or ofifoDataN[152] or ofifoDataN[151] or ofifoDataN[150] or ofifoDataN[149] or ofifoDataN[148] or ofifoDataN[147] or ofifoDataN[146]
 or ofifoDataN[145] or ofifoDataN[144] or ofifoDataN[143] or ofifoDataN[142] or ofifoDataN[141] or ofifoDataN[140] or ofifoDataN[139] or ofifoDataN[138]
 or ofifoDataN[137] or ofifoDataN[136] or ofifoDataN[135] or ofifoDataN[134] or ofifoDataN[133] or ofifoDataN[132] or ofifoDataN[131] or ofifoDataN[130]
 or ofifoDataN[129] or ofifoDataN[128] or ofifoDataN[127] or ofifoDataN[126] or ofifoDataN[125] or ofifoDataN[124] or ofifoDataN[123] or ofifoDataN[122]
 or ofifoDataN[121] or ofifoDataN[120] or ofifoDataN[119] or ofifoDataN[118] or ofifoDataN[117] or ofifoDataN[116] or ofifoDataN[115] or ofifoDataN[114]
 or ofifoDataN[113] or ofifoDataN[112] or ofifoDataN[111] or ofifoDataN[110] or ofifoDataN[109] or ofifoDataN[108] or ofifoDataN[107] or ofifoDataN[106]
 or ofifoDataN[105] or ofifoDataN[104] or ofifoDataN[103] or ofifoDataN[102] or ofifoDataN[101] or ofifoDataN[100] or ofifoDataN[99] or ofifoDataN[98]
 or ofifoDataN[97] or ofifoDataN[96] or ofifoDataN[95] or ofifoDataN[94] or ofifoDataN[93] or ofifoDataN[92] or ofifoDataN[91] or ofifoDataN[90]
 or ofifoDataN[89] or ofifoDataN[88] or ofifoDataN[87] or ofifoDataN[86] or ofifoDataN[85] or ofifoDataN[84] or ofifoDataN[83] or ofifoDataN[82]
 or ofifoDataN[81] or ofifoDataN[80] or ofifoDataN[79] or ofifoDataN[78] or ofifoDataN[77] or ofifoDataN[76] or ofifoDataN[75] or ofifoDataN[74]
 or ofifoDataN[73] or ofifoDataN[72] or ofifoDataN[71] or ofifoDataN[70] or ofifoDataN[69] or ofifoDataN[68] or ofifoDataN[67] or ofifoDataN[66]
 or ofifoDataN[65] or ofifoDataN[64] or ofifoDataN[63] or ofifoDataN[62] or ofifoDataN[61] or ofifoDataN[60] or ofifoDataN[59] or ofifoDataN[58]
 or ofifoDataN[57] or ofifoDataN[56] or ofifoDataN[55] or ofifoDataN[54] or ofifoDataN[53] or ofifoDataN[52] or ofifoDataN[51] or ofifoDataN[50]
 or ofifoDataN[49] or ofifoDataN[48] or ofifoDataN[47] or ofifoDataN[46] or ofifoDataN[45] or ofifoDataN[44] or ofifoDataN[43] or ofifoDataN[42]
 or ofifoDataN[41] or ofifoDataN[40] or ofifoDataN[39] or ofifoDataN[38] or ofifoDataN[37] or ofifoDataN[36] or ofifoDataN[35] or ofifoDataN[34]
 or ofifoDataN[33] or ofifoDataN[32] or ofifoDataN[31] or ofifoDataN[30] or ofifoDataN[29] or ofifoDataN[28] or ofifoDataN[27] or ofifoDataN[26]
 or ofifoDataN[25] or ofifoDataN[24] or ofifoDataN[23] or ofifoDataN[22] or ofifoDataN[21] or ofifoDataN[20] or ofifoDataN[19] or ofifoDataN[18]
 or ofifoDataN[17] or ofifoDataN[16] or ofifoDataN[15] or ofifoDataN[14] or ofifoDataN[13] or ofifoDataN[12] or ofifoDataN[11] or ofifoDataN[10]
 or ofifoDataN[9] or ofifoDataN[8] or ofifoDataN[7] or ofifoDataN[6] or ofifoDataN[5] or ofifoDataN[4] or ofifoDataN[3] or ofifoDataN[2]
 or ofifoDataN[1] or ofifoDataN[0] or n1572 or ofifoAddr1N[14] or ofifoAddr1N[13] or ofifoAddr1N[12] or ofifoAddr1N[11] or ofifoAddr1N[10]
 or ofifoAddr1N[9] or ofifoAddr1N[8] or ofifoAddr1N[7] or ofifoAddr1N[6] or ofifoAddr1N[5] or ofifoAddr1N[4] or ofifoAddr1N[3] or ofifoAddr1N[2]
 or ofifoAddr1N[1] or ofifoAddr1N[0] or ofifoDataN[511] or ofifoDataN[510] or ofifoDataN[509] or ofifoDataN[508] or ofifoDataN[507] or ofifoDataN[506]
 or ofifoDataN[505] or ofifoDataN[504] or ofifoDataN[503] or ofifoDataN[502] or ofifoDataN[501] or ofifoDataN[500] or ofifoDataN[499] or ofifoDataN[498]
 or ofifoDataN[497] or ofifoDataN[496] or ofifoDataN[495] or ofifoDataN[494] or ofifoDataN[493] or ofifoDataN[492] or ofifoDataN[491] or ofifoDataN[490]
 or ofifoDataN[489] or ofifoDataN[488] or ofifoDataN[487] or ofifoDataN[486] or ofifoDataN[485] or ofifoDataN[484] or ofifoDataN[483] or ofifoDataN[482]
 or ofifoDataN[481] or ofifoDataN[480] or ofifoDataN[479] or ofifoDataN[478] or ofifoDataN[477] or ofifoDataN[476] or ofifoDataN[475] or ofifoDataN[474]
 or ofifoDataN[473] or ofifoDataN[472] or ofifoDataN[471] or ofifoDataN[470] or ofifoDataN[469] or ofifoDataN[468] or ofifoDataN[467] or ofifoDataN[466]
 or ofifoDataN[465] or ofifoDataN[464] or ofifoDataN[463] or ofifoDataN[462] or ofifoDataN[461] or ofifoDataN[460] or ofifoDataN[459] or ofifoDataN[458]
 or ofifoDataN[457] or ofifoDataN[456] or ofifoDataN[455] or ofifoDataN[454] or ofifoDataN[453] or ofifoDataN[452] or ofifoDataN[451] or ofifoDataN[450]
 or ofifoDataN[449] or ofifoDataN[448] or ofifoDataN[447] or ofifoDataN[446] or ofifoDataN[445] or ofifoDataN[444] or ofifoDataN[443] or ofifoDataN[442]
 or ofifoDataN[441] or ofifoDataN[440] or ofifoDataN[439] or ofifoDataN[438] or ofifoDataN[437] or ofifoDataN[436] or ofifoDataN[435] or ofifoDataN[434]
 or ofifoDataN[433] or ofifoDataN[432] or ofifoDataN[431] or ofifoDataN[430] or ofifoDataN[429] or ofifoDataN[428] or ofifoDataN[427] or ofifoDataN[426]
 or ofifoDataN[425] or ofifoDataN[424] or ofifoDataN[423] or ofifoDataN[422] or ofifoDataN[421] or ofifoDataN[420] or ofifoDataN[419] or ofifoDataN[418]
 or ofifoDataN[417] or ofifoDataN[416] or ofifoDataN[415] or ofifoDataN[414] or ofifoDataN[413] or ofifoDataN[412] or ofifoDataN[411] or ofifoDataN[410]
 or ofifoDataN[409] or ofifoDataN[408] or ofifoDataN[407] or ofifoDataN[406] or ofifoDataN[405] or ofifoDataN[404] or ofifoDataN[403] or ofifoDataN[402]
 or ofifoDataN[401] or ofifoDataN[400] or ofifoDataN[399] or ofifoDataN[398] or ofifoDataN[397] or ofifoDataN[396] or ofifoDataN[395] or ofifoDataN[394]
 or ofifoDataN[393] or ofifoDataN[392] or ofifoDataN[391] or ofifoDataN[390] or ofifoDataN[389] or ofifoDataN[388] or ofifoDataN[387] or ofifoDataN[386]
 or ofifoDataN[385] or ofifoDataN[384] or ofifoDataN[383] or ofifoDataN[382] or ofifoDataN[381] or ofifoDataN[380] or ofifoDataN[379] or ofifoDataN[378]
 or ofifoDataN[377] or ofifoDataN[376] or ofifoDataN[375] or ofifoDataN[374] or ofifoDataN[373] or ofifoDataN[372] or ofifoDataN[371] or ofifoDataN[370]
 or ofifoDataN[369] or ofifoDataN[368] or ofifoDataN[367] or ofifoDataN[366] or ofifoDataN[365] or ofifoDataN[364] or ofifoDataN[363] or ofifoDataN[362]
 or ofifoDataN[361] or ofifoDataN[360] or ofifoDataN[359] or ofifoDataN[358] or ofifoDataN[357] or ofifoDataN[356] or ofifoDataN[355] or ofifoDataN[354]
 or ofifoDataN[353] or ofifoDataN[352] or ofifoDataN[351] or ofifoDataN[350] or ofifoDataN[349] or ofifoDataN[348] or ofifoDataN[347] or ofifoDataN[346]
 or ofifoDataN[345] or ofifoDataN[344] or ofifoDataN[343] or ofifoDataN[342] or ofifoDataN[341] or ofifoDataN[340] or ofifoDataN[339] or ofifoDataN[338]
 or ofifoDataN[337] or ofifoDataN[336] or ofifoDataN[335] or ofifoDataN[334] or ofifoDataN[333] or ofifoDataN[332] or ofifoDataN[331] or ofifoDataN[330]
 or ofifoDataN[329] or ofifoDataN[328] or ofifoDataN[327] or ofifoDataN[326] or ofifoDataN[325] or ofifoDataN[324] or ofifoDataN[323] or ofifoDataN[322]
 or ofifoDataN[321] or ofifoDataN[320] or ofifoDataN[319] or ofifoDataN[318] or ofifoDataN[317] or ofifoDataN[316] or ofifoDataN[315] or ofifoDataN[314]
 or ofifoDataN[313] or ofifoDataN[312] or ofifoDataN[311] or ofifoDataN[310] or ofifoDataN[309] or ofifoDataN[308] or ofifoDataN[307] or ofifoDataN[306]
 or ofifoDataN[305] or ofifoDataN[304] or ofifoDataN[303] or ofifoDataN[302] or ofifoDataN[301] or ofifoDataN[300] or ofifoDataN[299] or ofifoDataN[298]
 or ofifoDataN[297] or ofifoDataN[296] or ofifoDataN[295] or ofifoDataN[294] or ofifoDataN[293] or ofifoDataN[292] or ofifoDataN[291] or ofifoDataN[290]
 or ofifoDataN[289] or ofifoDataN[288] or ofifoDataN[287] or ofifoDataN[286] or ofifoDataN[285] or ofifoDataN[284] or ofifoDataN[283] or ofifoDataN[282]
 or ofifoDataN[281] or ofifoDataN[280] or ofifoDataN[279] or ofifoDataN[278] or ofifoDataN[277] or ofifoDataN[276] or ofifoDataN[275] or ofifoDataN[274]
 or ofifoDataN[273] or ofifoDataN[272] or ofifoDataN[271] or ofifoDataN[270] or ofifoDataN[269] or ofifoDataN[268] or ofifoDataN[267] or ofifoDataN[266]
 or ofifoDataN[265] or ofifoDataN[264] or ofifoDataN[263] or ofifoDataN[262] or ofifoDataN[261] or ofifoDataN[260] or ofifoDataN[259] or ofifoDataN[258]
 or ofifoDataN[257] or ofifoDataN[256] or ofifoAddr2N[14] or ofifoAddr2N[13] or ofifoAddr2N[12] or ofifoAddr2N[11] or ofifoAddr2N[10] or ofifoAddr2N[9]
 or ofifoAddr2N[8] or ofifoAddr2N[7] or ofifoAddr2N[6] or ofifoAddr2N[5] or ofifoAddr2N[4] or ofifoAddr2N[3] or ofifoAddr2N[2] or ofifoAddr2N[1]
 or ofifoDataN[767] or ofifoDataN[766] or ofifoDataN[765] or ofifoDataN[764] or ofifoDataN[763] or ofifoDataN[762] or ofifoDataN[761] or ofifoDataN[760]
 or ofifoDataN[759] or ofifoDataN[758] or ofifoDataN[757] or ofifoDataN[756] or ofifoDataN[755] or ofifoDataN[754] or ofifoDataN[753] or ofifoDataN[752]
 or ofifoDataN[751] or ofifoDataN[750] or ofifoDataN[749] or ofifoDataN[748] or ofifoDataN[747] or ofifoDataN[746] or ofifoDataN[745] or ofifoDataN[744]
 or ofifoDataN[743] or ofifoDataN[742] or ofifoDataN[741] or ofifoDataN[740] or ofifoDataN[739] or ofifoDataN[738] or ofifoDataN[737] or ofifoDataN[736]
 or ofifoDataN[735] or ofifoDataN[734] or ofifoDataN[733] or ofifoDataN[732] or ofifoDataN[731] or ofifoDataN[730] or ofifoDataN[729] or ofifoDataN[728]
 or ofifoDataN[727] or ofifoDataN[726] or ofifoDataN[725] or ofifoDataN[724] or ofifoDataN[723] or ofifoDataN[722] or ofifoDataN[721] or ofifoDataN[720]
 or ofifoDataN[719] or ofifoDataN[718] or ofifoDataN[717] or ofifoDataN[716] or ofifoDataN[715] or ofifoDataN[714] or ofifoDataN[713] or ofifoDataN[712]
 or ofifoDataN[711] or ofifoDataN[710] or ofifoDataN[709] or ofifoDataN[708] or ofifoDataN[707] or ofifoDataN[706] or ofifoDataN[705] or ofifoDataN[704]
 or ofifoDataN[703] or ofifoDataN[702] or ofifoDataN[701] or ofifoDataN[700] or ofifoDataN[699] or ofifoDataN[698] or ofifoDataN[697] or ofifoDataN[696]
 or ofifoDataN[695] or ofifoDataN[694] or ofifoDataN[693] or ofifoDataN[692] or ofifoDataN[691] or ofifoDataN[690] or ofifoDataN[689] or ofifoDataN[688]
 or ofifoDataN[687] or ofifoDataN[686] or ofifoDataN[685] or ofifoDataN[684] or ofifoDataN[683] or ofifoDataN[682] or ofifoDataN[681] or ofifoDataN[680]
 or ofifoDataN[679] or ofifoDataN[678] or ofifoDataN[677] or ofifoDataN[676] or ofifoDataN[675] or ofifoDataN[674] or ofifoDataN[673] or ofifoDataN[672]
 or ofifoDataN[671] or ofifoDataN[670] or ofifoDataN[669] or ofifoDataN[668] or ofifoDataN[667] or ofifoDataN[666] or ofifoDataN[665] or ofifoDataN[664]
 or ofifoDataN[663] or ofifoDataN[662] or ofifoDataN[661] or ofifoDataN[660] or ofifoDataN[659] or ofifoDataN[658] or ofifoDataN[657] or ofifoDataN[656]
 or ofifoDataN[655] or ofifoDataN[654] or ofifoDataN[653] or ofifoDataN[652] or ofifoDataN[651] or ofifoDataN[650] or ofifoDataN[649] or ofifoDataN[648]
 or ofifoDataN[647] or ofifoDataN[646] or ofifoDataN[645] or ofifoDataN[644] or ofifoDataN[643] or ofifoDataN[642] or ofifoDataN[641] or ofifoDataN[640]
 or ofifoDataN[639] or ofifoDataN[638] or ofifoDataN[637] or ofifoDataN[636] or ofifoDataN[635] or ofifoDataN[634] or ofifoDataN[633] or ofifoDataN[632]
 or ofifoDataN[631] or ofifoDataN[630] or ofifoDataN[629] or ofifoDataN[628] or ofifoDataN[627] or ofifoDataN[626] or ofifoDataN[625] or ofifoDataN[624]
 or ofifoDataN[623] or ofifoDataN[622] or ofifoDataN[621] or ofifoDataN[620] or ofifoDataN[619] or ofifoDataN[618] or ofifoDataN[617] or ofifoDataN[616]
 or ofifoDataN[615] or ofifoDataN[614] or ofifoDataN[613] or ofifoDataN[612] or ofifoDataN[611] or ofifoDataN[610] or ofifoDataN[609] or ofifoDataN[608]
 or ofifoDataN[607] or ofifoDataN[606] or ofifoDataN[605] or ofifoDataN[604] or ofifoDataN[603] or ofifoDataN[602] or ofifoDataN[601] or ofifoDataN[600]
 or ofifoDataN[599] or ofifoDataN[598] or ofifoDataN[597] or ofifoDataN[596] or ofifoDataN[595] or ofifoDataN[594] or ofifoDataN[593] or ofifoDataN[592]
 or ofifoDataN[591] or ofifoDataN[590] or ofifoDataN[589] or ofifoDataN[588] or ofifoDataN[587] or ofifoDataN[586] or ofifoDataN[585] or ofifoDataN[584]
 or ofifoDataN[583] or ofifoDataN[582] or ofifoDataN[581] or ofifoDataN[580] or ofifoDataN[579] or ofifoDataN[578] or ofifoDataN[577] or ofifoDataN[576]
 or ofifoDataN[575] or ofifoDataN[574] or ofifoDataN[573] or ofifoDataN[572] or ofifoDataN[571] or ofifoDataN[570] or ofifoDataN[569] or ofifoDataN[568]
 or ofifoDataN[567] or ofifoDataN[566] or ofifoDataN[565] or ofifoDataN[564] or ofifoDataN[563] or ofifoDataN[562] or ofifoDataN[561] or ofifoDataN[560]
 or ofifoDataN[559] or ofifoDataN[558] or ofifoDataN[557] or ofifoDataN[556] or ofifoDataN[555] or ofifoDataN[554] or ofifoDataN[553] or ofifoDataN[552]
 or ofifoDataN[551] or ofifoDataN[550] or ofifoDataN[549] or ofifoDataN[548] or ofifoDataN[547] or ofifoDataN[546] or ofifoDataN[545] or ofifoDataN[544]
 or ofifoDataN[543] or ofifoDataN[542] or ofifoDataN[541] or ofifoDataN[540] or ofifoDataN[539] or ofifoDataN[538] or ofifoDataN[537] or ofifoDataN[536]
 or ofifoDataN[535] or ofifoDataN[534] or ofifoDataN[533] or ofifoDataN[532] or ofifoDataN[531] or ofifoDataN[530] or ofifoDataN[529] or ofifoDataN[528]
 or ofifoDataN[527] or ofifoDataN[526] or ofifoDataN[525] or ofifoDataN[524] or ofifoDataN[523] or ofifoDataN[522] or ofifoDataN[521] or ofifoDataN[520]
 or ofifoDataN[519] or ofifoDataN[518] or ofifoDataN[517] or ofifoDataN[516] or ofifoDataN[515] or ofifoDataN[514] or ofifoDataN[513] or ofifoDataN[512])
#0 begin
if (n1572)
ixc_gfm_ofifo[{ofifoAddr0N[14], ofifoAddr0N[13], ofifoAddr0N[12], ofifoAddr0N[11], ofifoAddr0N[10],
 ofifoAddr0N[9], ofifoAddr0N[8], ofifoAddr0N[7], ofifoAddr0N[6], ofifoAddr0N[5], ofifoAddr0N[4], ofifoAddr0N[3], ofifoAddr0N[2],
 ofifoAddr0N[1], ofifoAddr0N[0]}] =
{ofifoDataN[255], ofifoDataN[254], ofifoDataN[253], ofifoDataN[252], ofifoDataN[251],
 ofifoDataN[250], ofifoDataN[249], ofifoDataN[248], ofifoDataN[247], ofifoDataN[246], ofifoDataN[245], ofifoDataN[244], ofifoDataN[243],
 ofifoDataN[242], ofifoDataN[241], ofifoDataN[240], ofifoDataN[239], ofifoDataN[238], ofifoDataN[237], ofifoDataN[236], ofifoDataN[235],
 ofifoDataN[234], ofifoDataN[233], ofifoDataN[232], ofifoDataN[231], ofifoDataN[230], ofifoDataN[229], ofifoDataN[228], ofifoDataN[227],
 ofifoDataN[226], ofifoDataN[225], ofifoDataN[224], ofifoDataN[223], ofifoDataN[222], ofifoDataN[221], ofifoDataN[220], ofifoDataN[219],
 ofifoDataN[218], ofifoDataN[217], ofifoDataN[216], ofifoDataN[215], ofifoDataN[214], ofifoDataN[213], ofifoDataN[212], ofifoDataN[211],
 ofifoDataN[210], ofifoDataN[209], ofifoDataN[208], ofifoDataN[207], ofifoDataN[206], ofifoDataN[205], ofifoDataN[204], ofifoDataN[203],
 ofifoDataN[202], ofifoDataN[201], ofifoDataN[200], ofifoDataN[199], ofifoDataN[198], ofifoDataN[197], ofifoDataN[196], ofifoDataN[195],
 ofifoDataN[194], ofifoDataN[193], ofifoDataN[192], ofifoDataN[191], ofifoDataN[190], ofifoDataN[189], ofifoDataN[188], ofifoDataN[187],
 ofifoDataN[186], ofifoDataN[185], ofifoDataN[184], ofifoDataN[183], ofifoDataN[182], ofifoDataN[181], ofifoDataN[180], ofifoDataN[179],
 ofifoDataN[178], ofifoDataN[177], ofifoDataN[176], ofifoDataN[175], ofifoDataN[174], ofifoDataN[173], ofifoDataN[172], ofifoDataN[171],
 ofifoDataN[170], ofifoDataN[169], ofifoDataN[168], ofifoDataN[167], ofifoDataN[166], ofifoDataN[165], ofifoDataN[164], ofifoDataN[163],
 ofifoDataN[162], ofifoDataN[161], ofifoDataN[160], ofifoDataN[159], ofifoDataN[158], ofifoDataN[157], ofifoDataN[156], ofifoDataN[155],
 ofifoDataN[154], ofifoDataN[153], ofifoDataN[152], ofifoDataN[151], ofifoDataN[150], ofifoDataN[149], ofifoDataN[148], ofifoDataN[147],
 ofifoDataN[146], ofifoDataN[145], ofifoDataN[144], ofifoDataN[143], ofifoDataN[142], ofifoDataN[141], ofifoDataN[140], ofifoDataN[139],
 ofifoDataN[138], ofifoDataN[137], ofifoDataN[136], ofifoDataN[135], ofifoDataN[134], ofifoDataN[133], ofifoDataN[132], ofifoDataN[131],
 ofifoDataN[130], ofifoDataN[129], ofifoDataN[128], ofifoDataN[127], ofifoDataN[126], ofifoDataN[125], ofifoDataN[124], ofifoDataN[123],
 ofifoDataN[122], ofifoDataN[121], ofifoDataN[120], ofifoDataN[119], ofifoDataN[118], ofifoDataN[117], ofifoDataN[116], ofifoDataN[115],
 ofifoDataN[114], ofifoDataN[113], ofifoDataN[112], ofifoDataN[111], ofifoDataN[110], ofifoDataN[109], ofifoDataN[108], ofifoDataN[107],
 ofifoDataN[106], ofifoDataN[105], ofifoDataN[104], ofifoDataN[103], ofifoDataN[102], ofifoDataN[101], ofifoDataN[100], ofifoDataN[99],
 ofifoDataN[98], ofifoDataN[97], ofifoDataN[96], ofifoDataN[95], ofifoDataN[94], ofifoDataN[93], ofifoDataN[92], ofifoDataN[91],
 ofifoDataN[90], ofifoDataN[89], ofifoDataN[88], ofifoDataN[87], ofifoDataN[86], ofifoDataN[85], ofifoDataN[84], ofifoDataN[83],
 ofifoDataN[82], ofifoDataN[81], ofifoDataN[80], ofifoDataN[79], ofifoDataN[78], ofifoDataN[77], ofifoDataN[76], ofifoDataN[75],
 ofifoDataN[74], ofifoDataN[73], ofifoDataN[72], ofifoDataN[71], ofifoDataN[70], ofifoDataN[69], ofifoDataN[68], ofifoDataN[67],
 ofifoDataN[66], ofifoDataN[65], ofifoDataN[64], ofifoDataN[63], ofifoDataN[62], ofifoDataN[61], ofifoDataN[60], ofifoDataN[59],
 ofifoDataN[58], ofifoDataN[57], ofifoDataN[56], ofifoDataN[55], ofifoDataN[54], ofifoDataN[53], ofifoDataN[52], ofifoDataN[51],
 ofifoDataN[50], ofifoDataN[49], ofifoDataN[48], ofifoDataN[47], ofifoDataN[46], ofifoDataN[45], ofifoDataN[44], ofifoDataN[43],
 ofifoDataN[42], ofifoDataN[41], ofifoDataN[40], ofifoDataN[39], ofifoDataN[38], ofifoDataN[37], ofifoDataN[36], ofifoDataN[35],
 ofifoDataN[34], ofifoDataN[33], ofifoDataN[32], ofifoDataN[31], ofifoDataN[30], ofifoDataN[29], ofifoDataN[28], ofifoDataN[27],
 ofifoDataN[26], ofifoDataN[25], ofifoDataN[24], ofifoDataN[23], ofifoDataN[22], ofifoDataN[21], ofifoDataN[20], ofifoDataN[19],
 ofifoDataN[18], ofifoDataN[17], ofifoDataN[16], ofifoDataN[15], ofifoDataN[14], ofifoDataN[13], ofifoDataN[12], ofifoDataN[11],
 ofifoDataN[10], ofifoDataN[9], ofifoDataN[8], ofifoDataN[7], ofifoDataN[6], ofifoDataN[5], ofifoDataN[4], ofifoDataN[3],
 ofifoDataN[2], ofifoDataN[1], ofifoDataN[0]};
if (n1572)
ixc_gfm_ofifo[{ofifoAddr1N[14], ofifoAddr1N[13], ofifoAddr1N[12], ofifoAddr1N[11], ofifoAddr1N[10],
 ofifoAddr1N[9], ofifoAddr1N[8], ofifoAddr1N[7], ofifoAddr1N[6], ofifoAddr1N[5], ofifoAddr1N[4], ofifoAddr1N[3], ofifoAddr1N[2],
 ofifoAddr1N[1], ofifoAddr1N[0]}] =
{ofifoDataN[511], ofifoDataN[510], ofifoDataN[509], ofifoDataN[508], ofifoDataN[507],
 ofifoDataN[506], ofifoDataN[505], ofifoDataN[504], ofifoDataN[503], ofifoDataN[502], ofifoDataN[501], ofifoDataN[500], ofifoDataN[499],
 ofifoDataN[498], ofifoDataN[497], ofifoDataN[496], ofifoDataN[495], ofifoDataN[494], ofifoDataN[493], ofifoDataN[492], ofifoDataN[491],
 ofifoDataN[490], ofifoDataN[489], ofifoDataN[488], ofifoDataN[487], ofifoDataN[486], ofifoDataN[485], ofifoDataN[484], ofifoDataN[483],
 ofifoDataN[482], ofifoDataN[481], ofifoDataN[480], ofifoDataN[479], ofifoDataN[478], ofifoDataN[477], ofifoDataN[476], ofifoDataN[475],
 ofifoDataN[474], ofifoDataN[473], ofifoDataN[472], ofifoDataN[471], ofifoDataN[470], ofifoDataN[469], ofifoDataN[468], ofifoDataN[467],
 ofifoDataN[466], ofifoDataN[465], ofifoDataN[464], ofifoDataN[463], ofifoDataN[462], ofifoDataN[461], ofifoDataN[460], ofifoDataN[459],
 ofifoDataN[458], ofifoDataN[457], ofifoDataN[456], ofifoDataN[455], ofifoDataN[454], ofifoDataN[453], ofifoDataN[452], ofifoDataN[451],
 ofifoDataN[450], ofifoDataN[449], ofifoDataN[448], ofifoDataN[447], ofifoDataN[446], ofifoDataN[445], ofifoDataN[444], ofifoDataN[443],
 ofifoDataN[442], ofifoDataN[441], ofifoDataN[440], ofifoDataN[439], ofifoDataN[438], ofifoDataN[437], ofifoDataN[436], ofifoDataN[435],
 ofifoDataN[434], ofifoDataN[433], ofifoDataN[432], ofifoDataN[431], ofifoDataN[430], ofifoDataN[429], ofifoDataN[428], ofifoDataN[427],
 ofifoDataN[426], ofifoDataN[425], ofifoDataN[424], ofifoDataN[423], ofifoDataN[422], ofifoDataN[421], ofifoDataN[420], ofifoDataN[419],
 ofifoDataN[418], ofifoDataN[417], ofifoDataN[416], ofifoDataN[415], ofifoDataN[414], ofifoDataN[413], ofifoDataN[412], ofifoDataN[411],
 ofifoDataN[410], ofifoDataN[409], ofifoDataN[408], ofifoDataN[407], ofifoDataN[406], ofifoDataN[405], ofifoDataN[404], ofifoDataN[403],
 ofifoDataN[402], ofifoDataN[401], ofifoDataN[400], ofifoDataN[399], ofifoDataN[398], ofifoDataN[397], ofifoDataN[396], ofifoDataN[395],
 ofifoDataN[394], ofifoDataN[393], ofifoDataN[392], ofifoDataN[391], ofifoDataN[390], ofifoDataN[389], ofifoDataN[388], ofifoDataN[387],
 ofifoDataN[386], ofifoDataN[385], ofifoDataN[384], ofifoDataN[383], ofifoDataN[382], ofifoDataN[381], ofifoDataN[380], ofifoDataN[379],
 ofifoDataN[378], ofifoDataN[377], ofifoDataN[376], ofifoDataN[375], ofifoDataN[374], ofifoDataN[373], ofifoDataN[372], ofifoDataN[371],
 ofifoDataN[370], ofifoDataN[369], ofifoDataN[368], ofifoDataN[367], ofifoDataN[366], ofifoDataN[365], ofifoDataN[364], ofifoDataN[363],
 ofifoDataN[362], ofifoDataN[361], ofifoDataN[360], ofifoDataN[359], ofifoDataN[358], ofifoDataN[357], ofifoDataN[356], ofifoDataN[355],
 ofifoDataN[354], ofifoDataN[353], ofifoDataN[352], ofifoDataN[351], ofifoDataN[350], ofifoDataN[349], ofifoDataN[348], ofifoDataN[347],
 ofifoDataN[346], ofifoDataN[345], ofifoDataN[344], ofifoDataN[343], ofifoDataN[342], ofifoDataN[341], ofifoDataN[340], ofifoDataN[339],
 ofifoDataN[338], ofifoDataN[337], ofifoDataN[336], ofifoDataN[335], ofifoDataN[334], ofifoDataN[333], ofifoDataN[332], ofifoDataN[331],
 ofifoDataN[330], ofifoDataN[329], ofifoDataN[328], ofifoDataN[327], ofifoDataN[326], ofifoDataN[325], ofifoDataN[324], ofifoDataN[323],
 ofifoDataN[322], ofifoDataN[321], ofifoDataN[320], ofifoDataN[319], ofifoDataN[318], ofifoDataN[317], ofifoDataN[316], ofifoDataN[315],
 ofifoDataN[314], ofifoDataN[313], ofifoDataN[312], ofifoDataN[311], ofifoDataN[310], ofifoDataN[309], ofifoDataN[308], ofifoDataN[307],
 ofifoDataN[306], ofifoDataN[305], ofifoDataN[304], ofifoDataN[303], ofifoDataN[302], ofifoDataN[301], ofifoDataN[300], ofifoDataN[299],
 ofifoDataN[298], ofifoDataN[297], ofifoDataN[296], ofifoDataN[295], ofifoDataN[294], ofifoDataN[293], ofifoDataN[292], ofifoDataN[291],
 ofifoDataN[290], ofifoDataN[289], ofifoDataN[288], ofifoDataN[287], ofifoDataN[286], ofifoDataN[285], ofifoDataN[284], ofifoDataN[283],
 ofifoDataN[282], ofifoDataN[281], ofifoDataN[280], ofifoDataN[279], ofifoDataN[278], ofifoDataN[277], ofifoDataN[276], ofifoDataN[275],
 ofifoDataN[274], ofifoDataN[273], ofifoDataN[272], ofifoDataN[271], ofifoDataN[270], ofifoDataN[269], ofifoDataN[268], ofifoDataN[267],
 ofifoDataN[266], ofifoDataN[265], ofifoDataN[264], ofifoDataN[263], ofifoDataN[262], ofifoDataN[261], ofifoDataN[260], ofifoDataN[259],
 ofifoDataN[258], ofifoDataN[257], ofifoDataN[256]};
if (n1572)
ixc_gfm_ofifo[{ofifoAddr2N[14], ofifoAddr2N[13], ofifoAddr2N[12], ofifoAddr2N[11], ofifoAddr2N[10],
 ofifoAddr2N[9], ofifoAddr2N[8], ofifoAddr2N[7], ofifoAddr2N[6], ofifoAddr2N[5], ofifoAddr2N[4], ofifoAddr2N[3], ofifoAddr2N[2],
 ofifoAddr2N[1], ofifoAddr0N[0]}] =
{ofifoDataN[767], ofifoDataN[766], ofifoDataN[765], ofifoDataN[764], ofifoDataN[763],
 ofifoDataN[762], ofifoDataN[761], ofifoDataN[760], ofifoDataN[759], ofifoDataN[758], ofifoDataN[757], ofifoDataN[756], ofifoDataN[755],
 ofifoDataN[754], ofifoDataN[753], ofifoDataN[752], ofifoDataN[751], ofifoDataN[750], ofifoDataN[749], ofifoDataN[748], ofifoDataN[747],
 ofifoDataN[746], ofifoDataN[745], ofifoDataN[744], ofifoDataN[743], ofifoDataN[742], ofifoDataN[741], ofifoDataN[740], ofifoDataN[739],
 ofifoDataN[738], ofifoDataN[737], ofifoDataN[736], ofifoDataN[735], ofifoDataN[734], ofifoDataN[733], ofifoDataN[732], ofifoDataN[731],
 ofifoDataN[730], ofifoDataN[729], ofifoDataN[728], ofifoDataN[727], ofifoDataN[726], ofifoDataN[725], ofifoDataN[724], ofifoDataN[723],
 ofifoDataN[722], ofifoDataN[721], ofifoDataN[720], ofifoDataN[719], ofifoDataN[718], ofifoDataN[717], ofifoDataN[716], ofifoDataN[715],
 ofifoDataN[714], ofifoDataN[713], ofifoDataN[712], ofifoDataN[711], ofifoDataN[710], ofifoDataN[709], ofifoDataN[708], ofifoDataN[707],
 ofifoDataN[706], ofifoDataN[705], ofifoDataN[704], ofifoDataN[703], ofifoDataN[702], ofifoDataN[701], ofifoDataN[700], ofifoDataN[699],
 ofifoDataN[698], ofifoDataN[697], ofifoDataN[696], ofifoDataN[695], ofifoDataN[694], ofifoDataN[693], ofifoDataN[692], ofifoDataN[691],
 ofifoDataN[690], ofifoDataN[689], ofifoDataN[688], ofifoDataN[687], ofifoDataN[686], ofifoDataN[685], ofifoDataN[684], ofifoDataN[683],
 ofifoDataN[682], ofifoDataN[681], ofifoDataN[680], ofifoDataN[679], ofifoDataN[678], ofifoDataN[677], ofifoDataN[676], ofifoDataN[675],
 ofifoDataN[674], ofifoDataN[673], ofifoDataN[672], ofifoDataN[671], ofifoDataN[670], ofifoDataN[669], ofifoDataN[668], ofifoDataN[667],
 ofifoDataN[666], ofifoDataN[665], ofifoDataN[664], ofifoDataN[663], ofifoDataN[662], ofifoDataN[661], ofifoDataN[660], ofifoDataN[659],
 ofifoDataN[658], ofifoDataN[657], ofifoDataN[656], ofifoDataN[655], ofifoDataN[654], ofifoDataN[653], ofifoDataN[652], ofifoDataN[651],
 ofifoDataN[650], ofifoDataN[649], ofifoDataN[648], ofifoDataN[647], ofifoDataN[646], ofifoDataN[645], ofifoDataN[644], ofifoDataN[643],
 ofifoDataN[642], ofifoDataN[641], ofifoDataN[640], ofifoDataN[639], ofifoDataN[638], ofifoDataN[637], ofifoDataN[636], ofifoDataN[635],
 ofifoDataN[634], ofifoDataN[633], ofifoDataN[632], ofifoDataN[631], ofifoDataN[630], ofifoDataN[629], ofifoDataN[628], ofifoDataN[627],
 ofifoDataN[626], ofifoDataN[625], ofifoDataN[624], ofifoDataN[623], ofifoDataN[622], ofifoDataN[621], ofifoDataN[620], ofifoDataN[619],
 ofifoDataN[618], ofifoDataN[617], ofifoDataN[616], ofifoDataN[615], ofifoDataN[614], ofifoDataN[613], ofifoDataN[612], ofifoDataN[611],
 ofifoDataN[610], ofifoDataN[609], ofifoDataN[608], ofifoDataN[607], ofifoDataN[606], ofifoDataN[605], ofifoDataN[604], ofifoDataN[603],
 ofifoDataN[602], ofifoDataN[601], ofifoDataN[600], ofifoDataN[599], ofifoDataN[598], ofifoDataN[597], ofifoDataN[596], ofifoDataN[595],
 ofifoDataN[594], ofifoDataN[593], ofifoDataN[592], ofifoDataN[591], ofifoDataN[590], ofifoDataN[589], ofifoDataN[588], ofifoDataN[587],
 ofifoDataN[586], ofifoDataN[585], ofifoDataN[584], ofifoDataN[583], ofifoDataN[582], ofifoDataN[581], ofifoDataN[580], ofifoDataN[579],
 ofifoDataN[578], ofifoDataN[577], ofifoDataN[576], ofifoDataN[575], ofifoDataN[574], ofifoDataN[573], ofifoDataN[572], ofifoDataN[571],
 ofifoDataN[570], ofifoDataN[569], ofifoDataN[568], ofifoDataN[567], ofifoDataN[566], ofifoDataN[565], ofifoDataN[564], ofifoDataN[563],
 ofifoDataN[562], ofifoDataN[561], ofifoDataN[560], ofifoDataN[559], ofifoDataN[558], ofifoDataN[557], ofifoDataN[556], ofifoDataN[555],
 ofifoDataN[554], ofifoDataN[553], ofifoDataN[552], ofifoDataN[551], ofifoDataN[550], ofifoDataN[549], ofifoDataN[548], ofifoDataN[547],
 ofifoDataN[546], ofifoDataN[545], ofifoDataN[544], ofifoDataN[543], ofifoDataN[542], ofifoDataN[541], ofifoDataN[540], ofifoDataN[539],
 ofifoDataN[538], ofifoDataN[537], ofifoDataN[536], ofifoDataN[535], ofifoDataN[534], ofifoDataN[533], ofifoDataN[532], ofifoDataN[531],
 ofifoDataN[530], ofifoDataN[529], ofifoDataN[528], ofifoDataN[527], ofifoDataN[526], ofifoDataN[525], ofifoDataN[524], ofifoDataN[523],
 ofifoDataN[522], ofifoDataN[521], ofifoDataN[520], ofifoDataN[519], ofifoDataN[518], ofifoDataN[517], ofifoDataN[516], ofifoDataN[515],
 ofifoDataN[514], ofifoDataN[513], ofifoDataN[512]};
end
`else

MPW32KX256 ixc_gfm_ofifo ( .A14(ofifoAddr0N[14]), .A13(ofifoAddr0N[13]), .A12(ofifoAddr0N[12]), .A11(ofifoAddr0N[11]), .A10(ofifoAddr0N[10]), .A9(ofifoAddr0N[9]),
 .A8(ofifoAddr0N[8]), .A7(ofifoAddr0N[7]), .A6(ofifoAddr0N[6]), .A5(ofifoAddr0N[5]), .A4(ofifoAddr0N[4]), .A3(ofifoAddr0N[3]), .A2(ofifoAddr0N[2]), .A1(ofifoAddr0N[1]),
 .A0(ofifoAddr0N[0]), .DI255(ofifoDataN[255]), .DI254(ofifoDataN[254]), .DI253(ofifoDataN[253]), .DI252(ofifoDataN[252]), .DI251(ofifoDataN[251]), .DI250(ofifoDataN[250]), .DI249(ofifoDataN[249]),
 .DI248(ofifoDataN[248]), .DI247(ofifoDataN[247]), .DI246(ofifoDataN[246]), .DI245(ofifoDataN[245]), .DI244(ofifoDataN[244]), .DI243(ofifoDataN[243]), .DI242(ofifoDataN[242]), .DI241(ofifoDataN[241]),
 .DI240(ofifoDataN[240]), .DI239(ofifoDataN[239]), .DI238(ofifoDataN[238]), .DI237(ofifoDataN[237]), .DI236(ofifoDataN[236]), .DI235(ofifoDataN[235]), .DI234(ofifoDataN[234]), .DI233(ofifoDataN[233]),
 .DI232(ofifoDataN[232]), .DI231(ofifoDataN[231]), .DI230(ofifoDataN[230]), .DI229(ofifoDataN[229]), .DI228(ofifoDataN[228]), .DI227(ofifoDataN[227]), .DI226(ofifoDataN[226]), .DI225(ofifoDataN[225]),
 .DI224(ofifoDataN[224]), .DI223(ofifoDataN[223]), .DI222(ofifoDataN[222]), .DI221(ofifoDataN[221]), .DI220(ofifoDataN[220]), .DI219(ofifoDataN[219]), .DI218(ofifoDataN[218]), .DI217(ofifoDataN[217]),
 .DI216(ofifoDataN[216]), .DI215(ofifoDataN[215]), .DI214(ofifoDataN[214]), .DI213(ofifoDataN[213]), .DI212(ofifoDataN[212]), .DI211(ofifoDataN[211]), .DI210(ofifoDataN[210]), .DI209(ofifoDataN[209]),
 .DI208(ofifoDataN[208]), .DI207(ofifoDataN[207]), .DI206(ofifoDataN[206]), .DI205(ofifoDataN[205]), .DI204(ofifoDataN[204]), .DI203(ofifoDataN[203]), .DI202(ofifoDataN[202]), .DI201(ofifoDataN[201]),
 .DI200(ofifoDataN[200]), .DI199(ofifoDataN[199]), .DI198(ofifoDataN[198]), .DI197(ofifoDataN[197]), .DI196(ofifoDataN[196]), .DI195(ofifoDataN[195]), .DI194(ofifoDataN[194]), .DI193(ofifoDataN[193]),
 .DI192(ofifoDataN[192]), .DI191(ofifoDataN[191]), .DI190(ofifoDataN[190]), .DI189(ofifoDataN[189]), .DI188(ofifoDataN[188]), .DI187(ofifoDataN[187]), .DI186(ofifoDataN[186]), .DI185(ofifoDataN[185]),
 .DI184(ofifoDataN[184]), .DI183(ofifoDataN[183]), .DI182(ofifoDataN[182]), .DI181(ofifoDataN[181]), .DI180(ofifoDataN[180]), .DI179(ofifoDataN[179]), .DI178(ofifoDataN[178]), .DI177(ofifoDataN[177]),
 .DI176(ofifoDataN[176]), .DI175(ofifoDataN[175]), .DI174(ofifoDataN[174]), .DI173(ofifoDataN[173]), .DI172(ofifoDataN[172]), .DI171(ofifoDataN[171]), .DI170(ofifoDataN[170]), .DI169(ofifoDataN[169]),
 .DI168(ofifoDataN[168]), .DI167(ofifoDataN[167]), .DI166(ofifoDataN[166]), .DI165(ofifoDataN[165]), .DI164(ofifoDataN[164]), .DI163(ofifoDataN[163]), .DI162(ofifoDataN[162]), .DI161(ofifoDataN[161]),
 .DI160(ofifoDataN[160]), .DI159(ofifoDataN[159]), .DI158(ofifoDataN[158]), .DI157(ofifoDataN[157]), .DI156(ofifoDataN[156]), .DI155(ofifoDataN[155]), .DI154(ofifoDataN[154]), .DI153(ofifoDataN[153]),
 .DI152(ofifoDataN[152]), .DI151(ofifoDataN[151]), .DI150(ofifoDataN[150]), .DI149(ofifoDataN[149]), .DI148(ofifoDataN[148]), .DI147(ofifoDataN[147]), .DI146(ofifoDataN[146]), .DI145(ofifoDataN[145]),
 .DI144(ofifoDataN[144]), .DI143(ofifoDataN[143]), .DI142(ofifoDataN[142]), .DI141(ofifoDataN[141]), .DI140(ofifoDataN[140]), .DI139(ofifoDataN[139]), .DI138(ofifoDataN[138]), .DI137(ofifoDataN[137]),
 .DI136(ofifoDataN[136]), .DI135(ofifoDataN[135]), .DI134(ofifoDataN[134]), .DI133(ofifoDataN[133]), .DI132(ofifoDataN[132]), .DI131(ofifoDataN[131]), .DI130(ofifoDataN[130]), .DI129(ofifoDataN[129]),
 .DI128(ofifoDataN[128]), .DI127(ofifoDataN[127]), .DI126(ofifoDataN[126]), .DI125(ofifoDataN[125]), .DI124(ofifoDataN[124]), .DI123(ofifoDataN[123]), .DI122(ofifoDataN[122]), .DI121(ofifoDataN[121]),
 .DI120(ofifoDataN[120]), .DI119(ofifoDataN[119]), .DI118(ofifoDataN[118]), .DI117(ofifoDataN[117]), .DI116(ofifoDataN[116]), .DI115(ofifoDataN[115]), .DI114(ofifoDataN[114]), .DI113(ofifoDataN[113]),
 .DI112(ofifoDataN[112]), .DI111(ofifoDataN[111]), .DI110(ofifoDataN[110]), .DI109(ofifoDataN[109]), .DI108(ofifoDataN[108]), .DI107(ofifoDataN[107]), .DI106(ofifoDataN[106]), .DI105(ofifoDataN[105]),
 .DI104(ofifoDataN[104]), .DI103(ofifoDataN[103]), .DI102(ofifoDataN[102]), .DI101(ofifoDataN[101]), .DI100(ofifoDataN[100]), .DI99(ofifoDataN[99]), .DI98(ofifoDataN[98]), .DI97(ofifoDataN[97]),
 .DI96(ofifoDataN[96]), .DI95(ofifoDataN[95]), .DI94(ofifoDataN[94]), .DI93(ofifoDataN[93]), .DI92(ofifoDataN[92]), .DI91(ofifoDataN[91]), .DI90(ofifoDataN[90]), .DI89(ofifoDataN[89]),
 .DI88(ofifoDataN[88]), .DI87(ofifoDataN[87]), .DI86(ofifoDataN[86]), .DI85(ofifoDataN[85]), .DI84(ofifoDataN[84]), .DI83(ofifoDataN[83]), .DI82(ofifoDataN[82]), .DI81(ofifoDataN[81]),
 .DI80(ofifoDataN[80]), .DI79(ofifoDataN[79]), .DI78(ofifoDataN[78]), .DI77(ofifoDataN[77]), .DI76(ofifoDataN[76]), .DI75(ofifoDataN[75]), .DI74(ofifoDataN[74]), .DI73(ofifoDataN[73]),
 .DI72(ofifoDataN[72]), .DI71(ofifoDataN[71]), .DI70(ofifoDataN[70]), .DI69(ofifoDataN[69]), .DI68(ofifoDataN[68]), .DI67(ofifoDataN[67]), .DI66(ofifoDataN[66]), .DI65(ofifoDataN[65]),
 .DI64(ofifoDataN[64]), .DI63(ofifoDataN[63]), .DI62(ofifoDataN[62]), .DI61(ofifoDataN[61]), .DI60(ofifoDataN[60]), .DI59(ofifoDataN[59]), .DI58(ofifoDataN[58]), .DI57(ofifoDataN[57]),
 .DI56(ofifoDataN[56]), .DI55(ofifoDataN[55]), .DI54(ofifoDataN[54]), .DI53(ofifoDataN[53]), .DI52(ofifoDataN[52]), .DI51(ofifoDataN[51]), .DI50(ofifoDataN[50]), .DI49(ofifoDataN[49]),
 .DI48(ofifoDataN[48]), .DI47(ofifoDataN[47]), .DI46(ofifoDataN[46]), .DI45(ofifoDataN[45]), .DI44(ofifoDataN[44]), .DI43(ofifoDataN[43]), .DI42(ofifoDataN[42]), .DI41(ofifoDataN[41]),
 .DI40(ofifoDataN[40]), .DI39(ofifoDataN[39]), .DI38(ofifoDataN[38]), .DI37(ofifoDataN[37]), .DI36(ofifoDataN[36]), .DI35(ofifoDataN[35]), .DI34(ofifoDataN[34]), .DI33(ofifoDataN[33]),
 .DI32(ofifoDataN[32]), .DI31(ofifoDataN[31]), .DI30(ofifoDataN[30]), .DI29(ofifoDataN[29]), .DI28(ofifoDataN[28]), .DI27(ofifoDataN[27]), .DI26(ofifoDataN[26]), .DI25(ofifoDataN[25]),
 .DI24(ofifoDataN[24]), .DI23(ofifoDataN[23]), .DI22(ofifoDataN[22]), .DI21(ofifoDataN[21]), .DI20(ofifoDataN[20]), .DI19(ofifoDataN[19]), .DI18(ofifoDataN[18]), .DI17(ofifoDataN[17]),
 .DI16(ofifoDataN[16]), .DI15(ofifoDataN[15]), .DI14(ofifoDataN[14]), .DI13(ofifoDataN[13]), .DI12(ofifoDataN[12]), .DI11(ofifoDataN[11]), .DI10(ofifoDataN[10]), .DI9(ofifoDataN[9]),
 .DI8(ofifoDataN[8]), .DI7(ofifoDataN[7]), .DI6(ofifoDataN[6]), .DI5(ofifoDataN[5]), .DI4(ofifoDataN[4]), .DI3(ofifoDataN[3]), .DI2(ofifoDataN[2]), .DI1(ofifoDataN[1]),
 .DI0(ofifoDataN[0]), .WE(n1572), .SYNC_IN(n1611), .SYNC_OUT(n6742));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ofifo" HDL_MEMORY_DECL "1 255 0 0 32767"
MPW32KX256 U9486 ( .A14(ofifoAddr1N[14]), .A13(ofifoAddr1N[13]), .A12(ofifoAddr1N[12]), .A11(ofifoAddr1N[11]), .A10(ofifoAddr1N[10]), .A9(ofifoAddr1N[9]),
 .A8(ofifoAddr1N[8]), .A7(ofifoAddr1N[7]), .A6(ofifoAddr1N[6]), .A5(ofifoAddr1N[5]), .A4(ofifoAddr1N[4]), .A3(ofifoAddr1N[3]), .A2(ofifoAddr1N[2]), .A1(ofifoAddr1N[1]),
 .A0(ofifoAddr1N[0]), .DI255(ofifoDataN[511]), .DI254(ofifoDataN[510]), .DI253(ofifoDataN[509]), .DI252(ofifoDataN[508]), .DI251(ofifoDataN[507]), .DI250(ofifoDataN[506]), .DI249(ofifoDataN[505]),
 .DI248(ofifoDataN[504]), .DI247(ofifoDataN[503]), .DI246(ofifoDataN[502]), .DI245(ofifoDataN[501]), .DI244(ofifoDataN[500]), .DI243(ofifoDataN[499]), .DI242(ofifoDataN[498]), .DI241(ofifoDataN[497]),
 .DI240(ofifoDataN[496]), .DI239(ofifoDataN[495]), .DI238(ofifoDataN[494]), .DI237(ofifoDataN[493]), .DI236(ofifoDataN[492]), .DI235(ofifoDataN[491]), .DI234(ofifoDataN[490]), .DI233(ofifoDataN[489]),
 .DI232(ofifoDataN[488]), .DI231(ofifoDataN[487]), .DI230(ofifoDataN[486]), .DI229(ofifoDataN[485]), .DI228(ofifoDataN[484]), .DI227(ofifoDataN[483]), .DI226(ofifoDataN[482]), .DI225(ofifoDataN[481]),
 .DI224(ofifoDataN[480]), .DI223(ofifoDataN[479]), .DI222(ofifoDataN[478]), .DI221(ofifoDataN[477]), .DI220(ofifoDataN[476]), .DI219(ofifoDataN[475]), .DI218(ofifoDataN[474]), .DI217(ofifoDataN[473]),
 .DI216(ofifoDataN[472]), .DI215(ofifoDataN[471]), .DI214(ofifoDataN[470]), .DI213(ofifoDataN[469]), .DI212(ofifoDataN[468]), .DI211(ofifoDataN[467]), .DI210(ofifoDataN[466]), .DI209(ofifoDataN[465]),
 .DI208(ofifoDataN[464]), .DI207(ofifoDataN[463]), .DI206(ofifoDataN[462]), .DI205(ofifoDataN[461]), .DI204(ofifoDataN[460]), .DI203(ofifoDataN[459]), .DI202(ofifoDataN[458]), .DI201(ofifoDataN[457]),
 .DI200(ofifoDataN[456]), .DI199(ofifoDataN[455]), .DI198(ofifoDataN[454]), .DI197(ofifoDataN[453]), .DI196(ofifoDataN[452]), .DI195(ofifoDataN[451]), .DI194(ofifoDataN[450]), .DI193(ofifoDataN[449]),
 .DI192(ofifoDataN[448]), .DI191(ofifoDataN[447]), .DI190(ofifoDataN[446]), .DI189(ofifoDataN[445]), .DI188(ofifoDataN[444]), .DI187(ofifoDataN[443]), .DI186(ofifoDataN[442]), .DI185(ofifoDataN[441]),
 .DI184(ofifoDataN[440]), .DI183(ofifoDataN[439]), .DI182(ofifoDataN[438]), .DI181(ofifoDataN[437]), .DI180(ofifoDataN[436]), .DI179(ofifoDataN[435]), .DI178(ofifoDataN[434]), .DI177(ofifoDataN[433]),
 .DI176(ofifoDataN[432]), .DI175(ofifoDataN[431]), .DI174(ofifoDataN[430]), .DI173(ofifoDataN[429]), .DI172(ofifoDataN[428]), .DI171(ofifoDataN[427]), .DI170(ofifoDataN[426]), .DI169(ofifoDataN[425]),
 .DI168(ofifoDataN[424]), .DI167(ofifoDataN[423]), .DI166(ofifoDataN[422]), .DI165(ofifoDataN[421]), .DI164(ofifoDataN[420]), .DI163(ofifoDataN[419]), .DI162(ofifoDataN[418]), .DI161(ofifoDataN[417]),
 .DI160(ofifoDataN[416]), .DI159(ofifoDataN[415]), .DI158(ofifoDataN[414]), .DI157(ofifoDataN[413]), .DI156(ofifoDataN[412]), .DI155(ofifoDataN[411]), .DI154(ofifoDataN[410]), .DI153(ofifoDataN[409]),
 .DI152(ofifoDataN[408]), .DI151(ofifoDataN[407]), .DI150(ofifoDataN[406]), .DI149(ofifoDataN[405]), .DI148(ofifoDataN[404]), .DI147(ofifoDataN[403]), .DI146(ofifoDataN[402]), .DI145(ofifoDataN[401]),
 .DI144(ofifoDataN[400]), .DI143(ofifoDataN[399]), .DI142(ofifoDataN[398]), .DI141(ofifoDataN[397]), .DI140(ofifoDataN[396]), .DI139(ofifoDataN[395]), .DI138(ofifoDataN[394]), .DI137(ofifoDataN[393]),
 .DI136(ofifoDataN[392]), .DI135(ofifoDataN[391]), .DI134(ofifoDataN[390]), .DI133(ofifoDataN[389]), .DI132(ofifoDataN[388]), .DI131(ofifoDataN[387]), .DI130(ofifoDataN[386]), .DI129(ofifoDataN[385]),
 .DI128(ofifoDataN[384]), .DI127(ofifoDataN[383]), .DI126(ofifoDataN[382]), .DI125(ofifoDataN[381]), .DI124(ofifoDataN[380]), .DI123(ofifoDataN[379]), .DI122(ofifoDataN[378]), .DI121(ofifoDataN[377]),
 .DI120(ofifoDataN[376]), .DI119(ofifoDataN[375]), .DI118(ofifoDataN[374]), .DI117(ofifoDataN[373]), .DI116(ofifoDataN[372]), .DI115(ofifoDataN[371]), .DI114(ofifoDataN[370]), .DI113(ofifoDataN[369]),
 .DI112(ofifoDataN[368]), .DI111(ofifoDataN[367]), .DI110(ofifoDataN[366]), .DI109(ofifoDataN[365]), .DI108(ofifoDataN[364]), .DI107(ofifoDataN[363]), .DI106(ofifoDataN[362]), .DI105(ofifoDataN[361]),
 .DI104(ofifoDataN[360]), .DI103(ofifoDataN[359]), .DI102(ofifoDataN[358]), .DI101(ofifoDataN[357]), .DI100(ofifoDataN[356]), .DI99(ofifoDataN[355]), .DI98(ofifoDataN[354]), .DI97(ofifoDataN[353]),
 .DI96(ofifoDataN[352]), .DI95(ofifoDataN[351]), .DI94(ofifoDataN[350]), .DI93(ofifoDataN[349]), .DI92(ofifoDataN[348]), .DI91(ofifoDataN[347]), .DI90(ofifoDataN[346]), .DI89(ofifoDataN[345]),
 .DI88(ofifoDataN[344]), .DI87(ofifoDataN[343]), .DI86(ofifoDataN[342]), .DI85(ofifoDataN[341]), .DI84(ofifoDataN[340]), .DI83(ofifoDataN[339]), .DI82(ofifoDataN[338]), .DI81(ofifoDataN[337]),
 .DI80(ofifoDataN[336]), .DI79(ofifoDataN[335]), .DI78(ofifoDataN[334]), .DI77(ofifoDataN[333]), .DI76(ofifoDataN[332]), .DI75(ofifoDataN[331]), .DI74(ofifoDataN[330]), .DI73(ofifoDataN[329]),
 .DI72(ofifoDataN[328]), .DI71(ofifoDataN[327]), .DI70(ofifoDataN[326]), .DI69(ofifoDataN[325]), .DI68(ofifoDataN[324]), .DI67(ofifoDataN[323]), .DI66(ofifoDataN[322]), .DI65(ofifoDataN[321]),
 .DI64(ofifoDataN[320]), .DI63(ofifoDataN[319]), .DI62(ofifoDataN[318]), .DI61(ofifoDataN[317]), .DI60(ofifoDataN[316]), .DI59(ofifoDataN[315]), .DI58(ofifoDataN[314]), .DI57(ofifoDataN[313]),
 .DI56(ofifoDataN[312]), .DI55(ofifoDataN[311]), .DI54(ofifoDataN[310]), .DI53(ofifoDataN[309]), .DI52(ofifoDataN[308]), .DI51(ofifoDataN[307]), .DI50(ofifoDataN[306]), .DI49(ofifoDataN[305]),
 .DI48(ofifoDataN[304]), .DI47(ofifoDataN[303]), .DI46(ofifoDataN[302]), .DI45(ofifoDataN[301]), .DI44(ofifoDataN[300]), .DI43(ofifoDataN[299]), .DI42(ofifoDataN[298]), .DI41(ofifoDataN[297]),
 .DI40(ofifoDataN[296]), .DI39(ofifoDataN[295]), .DI38(ofifoDataN[294]), .DI37(ofifoDataN[293]), .DI36(ofifoDataN[292]), .DI35(ofifoDataN[291]), .DI34(ofifoDataN[290]), .DI33(ofifoDataN[289]),
 .DI32(ofifoDataN[288]), .DI31(ofifoDataN[287]), .DI30(ofifoDataN[286]), .DI29(ofifoDataN[285]), .DI28(ofifoDataN[284]), .DI27(ofifoDataN[283]), .DI26(ofifoDataN[282]), .DI25(ofifoDataN[281]),
 .DI24(ofifoDataN[280]), .DI23(ofifoDataN[279]), .DI22(ofifoDataN[278]), .DI21(ofifoDataN[277]), .DI20(ofifoDataN[276]), .DI19(ofifoDataN[275]), .DI18(ofifoDataN[274]), .DI17(ofifoDataN[273]),
 .DI16(ofifoDataN[272]), .DI15(ofifoDataN[271]), .DI14(ofifoDataN[270]), .DI13(ofifoDataN[269]), .DI12(ofifoDataN[268]), .DI11(ofifoDataN[267]), .DI10(ofifoDataN[266]), .DI9(ofifoDataN[265]),
 .DI8(ofifoDataN[264]), .DI7(ofifoDataN[263]), .DI6(ofifoDataN[262]), .DI5(ofifoDataN[261]), .DI4(ofifoDataN[260]), .DI3(ofifoDataN[259]), .DI2(ofifoDataN[258]), .DI1(ofifoDataN[257]),
 .DI0(ofifoDataN[256]), .WE(n1572), .SYNC_IN(n6742), .SYNC_OUT(n6743));
MPW32KX256 U9487 ( .A14(ofifoAddr2N[14]), .A13(ofifoAddr2N[13]), .A12(ofifoAddr2N[12]), .A11(ofifoAddr2N[11]), .A10(ofifoAddr2N[10]), .A9(ofifoAddr2N[9]),
 .A8(ofifoAddr2N[8]), .A7(ofifoAddr2N[7]), .A6(ofifoAddr2N[6]), .A5(ofifoAddr2N[5]), .A4(ofifoAddr2N[4]), .A3(ofifoAddr2N[3]), .A2(ofifoAddr2N[2]), .A1(ofifoAddr2N[1]),
 .A0(ofifoAddr0N[0]), .DI255(ofifoDataN[767]), .DI254(ofifoDataN[766]), .DI253(ofifoDataN[765]), .DI252(ofifoDataN[764]), .DI251(ofifoDataN[763]), .DI250(ofifoDataN[762]), .DI249(ofifoDataN[761]),
 .DI248(ofifoDataN[760]), .DI247(ofifoDataN[759]), .DI246(ofifoDataN[758]), .DI245(ofifoDataN[757]), .DI244(ofifoDataN[756]), .DI243(ofifoDataN[755]), .DI242(ofifoDataN[754]), .DI241(ofifoDataN[753]),
 .DI240(ofifoDataN[752]), .DI239(ofifoDataN[751]), .DI238(ofifoDataN[750]), .DI237(ofifoDataN[749]), .DI236(ofifoDataN[748]), .DI235(ofifoDataN[747]), .DI234(ofifoDataN[746]), .DI233(ofifoDataN[745]),
 .DI232(ofifoDataN[744]), .DI231(ofifoDataN[743]), .DI230(ofifoDataN[742]), .DI229(ofifoDataN[741]), .DI228(ofifoDataN[740]), .DI227(ofifoDataN[739]), .DI226(ofifoDataN[738]), .DI225(ofifoDataN[737]),
 .DI224(ofifoDataN[736]), .DI223(ofifoDataN[735]), .DI222(ofifoDataN[734]), .DI221(ofifoDataN[733]), .DI220(ofifoDataN[732]), .DI219(ofifoDataN[731]), .DI218(ofifoDataN[730]), .DI217(ofifoDataN[729]),
 .DI216(ofifoDataN[728]), .DI215(ofifoDataN[727]), .DI214(ofifoDataN[726]), .DI213(ofifoDataN[725]), .DI212(ofifoDataN[724]), .DI211(ofifoDataN[723]), .DI210(ofifoDataN[722]), .DI209(ofifoDataN[721]),
 .DI208(ofifoDataN[720]), .DI207(ofifoDataN[719]), .DI206(ofifoDataN[718]), .DI205(ofifoDataN[717]), .DI204(ofifoDataN[716]), .DI203(ofifoDataN[715]), .DI202(ofifoDataN[714]), .DI201(ofifoDataN[713]),
 .DI200(ofifoDataN[712]), .DI199(ofifoDataN[711]), .DI198(ofifoDataN[710]), .DI197(ofifoDataN[709]), .DI196(ofifoDataN[708]), .DI195(ofifoDataN[707]), .DI194(ofifoDataN[706]), .DI193(ofifoDataN[705]),
 .DI192(ofifoDataN[704]), .DI191(ofifoDataN[703]), .DI190(ofifoDataN[702]), .DI189(ofifoDataN[701]), .DI188(ofifoDataN[700]), .DI187(ofifoDataN[699]), .DI186(ofifoDataN[698]), .DI185(ofifoDataN[697]),
 .DI184(ofifoDataN[696]), .DI183(ofifoDataN[695]), .DI182(ofifoDataN[694]), .DI181(ofifoDataN[693]), .DI180(ofifoDataN[692]), .DI179(ofifoDataN[691]), .DI178(ofifoDataN[690]), .DI177(ofifoDataN[689]),
 .DI176(ofifoDataN[688]), .DI175(ofifoDataN[687]), .DI174(ofifoDataN[686]), .DI173(ofifoDataN[685]), .DI172(ofifoDataN[684]), .DI171(ofifoDataN[683]), .DI170(ofifoDataN[682]), .DI169(ofifoDataN[681]),
 .DI168(ofifoDataN[680]), .DI167(ofifoDataN[679]), .DI166(ofifoDataN[678]), .DI165(ofifoDataN[677]), .DI164(ofifoDataN[676]), .DI163(ofifoDataN[675]), .DI162(ofifoDataN[674]), .DI161(ofifoDataN[673]),
 .DI160(ofifoDataN[672]), .DI159(ofifoDataN[671]), .DI158(ofifoDataN[670]), .DI157(ofifoDataN[669]), .DI156(ofifoDataN[668]), .DI155(ofifoDataN[667]), .DI154(ofifoDataN[666]), .DI153(ofifoDataN[665]),
 .DI152(ofifoDataN[664]), .DI151(ofifoDataN[663]), .DI150(ofifoDataN[662]), .DI149(ofifoDataN[661]), .DI148(ofifoDataN[660]), .DI147(ofifoDataN[659]), .DI146(ofifoDataN[658]), .DI145(ofifoDataN[657]),
 .DI144(ofifoDataN[656]), .DI143(ofifoDataN[655]), .DI142(ofifoDataN[654]), .DI141(ofifoDataN[653]), .DI140(ofifoDataN[652]), .DI139(ofifoDataN[651]), .DI138(ofifoDataN[650]), .DI137(ofifoDataN[649]),
 .DI136(ofifoDataN[648]), .DI135(ofifoDataN[647]), .DI134(ofifoDataN[646]), .DI133(ofifoDataN[645]), .DI132(ofifoDataN[644]), .DI131(ofifoDataN[643]), .DI130(ofifoDataN[642]), .DI129(ofifoDataN[641]),
 .DI128(ofifoDataN[640]), .DI127(ofifoDataN[639]), .DI126(ofifoDataN[638]), .DI125(ofifoDataN[637]), .DI124(ofifoDataN[636]), .DI123(ofifoDataN[635]), .DI122(ofifoDataN[634]), .DI121(ofifoDataN[633]),
 .DI120(ofifoDataN[632]), .DI119(ofifoDataN[631]), .DI118(ofifoDataN[630]), .DI117(ofifoDataN[629]), .DI116(ofifoDataN[628]), .DI115(ofifoDataN[627]), .DI114(ofifoDataN[626]), .DI113(ofifoDataN[625]),
 .DI112(ofifoDataN[624]), .DI111(ofifoDataN[623]), .DI110(ofifoDataN[622]), .DI109(ofifoDataN[621]), .DI108(ofifoDataN[620]), .DI107(ofifoDataN[619]), .DI106(ofifoDataN[618]), .DI105(ofifoDataN[617]),
 .DI104(ofifoDataN[616]), .DI103(ofifoDataN[615]), .DI102(ofifoDataN[614]), .DI101(ofifoDataN[613]), .DI100(ofifoDataN[612]), .DI99(ofifoDataN[611]), .DI98(ofifoDataN[610]), .DI97(ofifoDataN[609]),
 .DI96(ofifoDataN[608]), .DI95(ofifoDataN[607]), .DI94(ofifoDataN[606]), .DI93(ofifoDataN[605]), .DI92(ofifoDataN[604]), .DI91(ofifoDataN[603]), .DI90(ofifoDataN[602]), .DI89(ofifoDataN[601]),
 .DI88(ofifoDataN[600]), .DI87(ofifoDataN[599]), .DI86(ofifoDataN[598]), .DI85(ofifoDataN[597]), .DI84(ofifoDataN[596]), .DI83(ofifoDataN[595]), .DI82(ofifoDataN[594]), .DI81(ofifoDataN[593]),
 .DI80(ofifoDataN[592]), .DI79(ofifoDataN[591]), .DI78(ofifoDataN[590]), .DI77(ofifoDataN[589]), .DI76(ofifoDataN[588]), .DI75(ofifoDataN[587]), .DI74(ofifoDataN[586]), .DI73(ofifoDataN[585]),
 .DI72(ofifoDataN[584]), .DI71(ofifoDataN[583]), .DI70(ofifoDataN[582]), .DI69(ofifoDataN[581]), .DI68(ofifoDataN[580]), .DI67(ofifoDataN[579]), .DI66(ofifoDataN[578]), .DI65(ofifoDataN[577]),
 .DI64(ofifoDataN[576]), .DI63(ofifoDataN[575]), .DI62(ofifoDataN[574]), .DI61(ofifoDataN[573]), .DI60(ofifoDataN[572]), .DI59(ofifoDataN[571]), .DI58(ofifoDataN[570]), .DI57(ofifoDataN[569]),
 .DI56(ofifoDataN[568]), .DI55(ofifoDataN[567]), .DI54(ofifoDataN[566]), .DI53(ofifoDataN[565]), .DI52(ofifoDataN[564]), .DI51(ofifoDataN[563]), .DI50(ofifoDataN[562]), .DI49(ofifoDataN[561]),
 .DI48(ofifoDataN[560]), .DI47(ofifoDataN[559]), .DI46(ofifoDataN[558]), .DI45(ofifoDataN[557]), .DI44(ofifoDataN[556]), .DI43(ofifoDataN[555]), .DI42(ofifoDataN[554]), .DI41(ofifoDataN[553]),
 .DI40(ofifoDataN[552]), .DI39(ofifoDataN[551]), .DI38(ofifoDataN[550]), .DI37(ofifoDataN[549]), .DI36(ofifoDataN[548]), .DI35(ofifoDataN[547]), .DI34(ofifoDataN[546]), .DI33(ofifoDataN[545]),
 .DI32(ofifoDataN[544]), .DI31(ofifoDataN[543]), .DI30(ofifoDataN[542]), .DI29(ofifoDataN[541]), .DI28(ofifoDataN[540]), .DI27(ofifoDataN[539]), .DI26(ofifoDataN[538]), .DI25(ofifoDataN[537]),
 .DI24(ofifoDataN[536]), .DI23(ofifoDataN[535]), .DI22(ofifoDataN[534]), .DI21(ofifoDataN[533]), .DI20(ofifoDataN[532]), .DI19(ofifoDataN[531]), .DI18(ofifoDataN[530]), .DI17(ofifoDataN[529]),
 .DI16(ofifoDataN[528]), .DI15(ofifoDataN[527]), .DI14(ofifoDataN[526]), .DI13(ofifoDataN[525]), .DI12(ofifoDataN[524]), .DI11(ofifoDataN[523]), .DI10(ofifoDataN[522]), .DI9(ofifoDataN[521]),
 .DI8(ofifoDataN[520]), .DI7(ofifoDataN[519]), .DI6(ofifoDataN[518]), .DI5(ofifoDataN[517]), .DI4(ofifoDataN[516]), .DI3(ofifoDataN[515]), .DI2(ofifoDataN[514]), .DI1(ofifoDataN[513]),
 .DI0(ofifoDataN[512]), .WE(n1572), .SYNC_IN(n6743), .SYNC_OUT( ));
`endif
`ifdef CBV

reg [63:0] ixc_gfm_ctl [0:3];
always @(n1611 or wrtCntD[62] or wrtCntD[61] or wrtCntD[60] or wrtCntD[59]
 or wrtCntD[58] or wrtCntD[57] or wrtCntD[56] or wrtCntD[55] or wrtCntD[54] or wrtCntD[53] or wrtCntD[52] or wrtCntD[51]
 or wrtCntD[50] or wrtCntD[49] or wrtCntD[48] or wrtCntD[47] or wrtCntD[46] or wrtCntD[45] or wrtCntD[44] or wrtCntD[43]
 or wrtCntD[42] or wrtCntD[41] or wrtCntD[40] or wrtCntD[39] or wrtCntD[38] or wrtCntD[37] or wrtCntD[36] or wrtCntD[35]
 or wrtCntD[34] or wrtCntD[33] or wrtCntD[32] or wrtCntD[31] or wrtCntD[30] or wrtCntD[29] or wrtCntD[28] or wrtCntD[27]
 or wrtCntD[26] or wrtCntD[25] or wrtCntD[24] or wrtCntD[23] or wrtCntD[22] or wrtCntD[21] or wrtCntD[20] or wrtCntD[19]
 or wrtCntD[18] or wrtCntD[17] or wrtCntD[16] or wrtCntD[15] or wrtCntD[14] or wrtCntD[13] or wrtCntD[12] or wrtCntD[11]
 or wrtCntD[10] or wrtCntD[9] or wrtCntD[8] or wrtCntD[7] or wrtCntD[6] or wrtCntD[5] or wrtCntD[4] or wrtCntD[3]
 or wrtCntD[2] or wrtCntD[1] or wrtCntD[0] or xc_top.svGFbusy or n1572 or rdCnt[63] or rdCnt[62] or rdCnt[61]
 or rdCnt[60] or rdCnt[59] or rdCnt[58] or rdCnt[57] or rdCnt[56] or rdCnt[55] or rdCnt[54] or rdCnt[53]
 or rdCnt[52] or rdCnt[51] or rdCnt[50] or rdCnt[49] or rdCnt[48] or rdCnt[47] or rdCnt[46] or rdCnt[45]
 or rdCnt[44] or rdCnt[43] or rdCnt[42] or rdCnt[41] or rdCnt[40] or rdCnt[39] or rdCnt[38] or rdCnt[37]
 or rdCnt[36] or rdCnt[35] or rdCnt[34] or rdCnt[33] or rdCnt[32] or rdCnt[31] or rdCnt[30] or rdCnt[29]
 or rdCnt[28] or rdCnt[27] or rdCnt[26] or rdCnt[25] or rdCnt[24] or rdCnt[23] or rdCnt[22] or rdCnt[21]
 or rdCnt[20] or rdCnt[19] or rdCnt[18] or rdCnt[17] or rdCnt[16] or rdCnt[15] or rdCnt[14] or rdCnt[13]
 or rdCnt[12] or rdCnt[11] or rdCnt[10] or rdCnt[9] or rdCnt[8] or rdCnt[7] or rdCnt[6] or rdCnt[5]
 or rdCnt[4] or rdCnt[3] or rdCnt[2] or rdCnt[1] or rdCnt[0] or xc_top.ixcSimTime[62] or xc_top.ixcSimTime[61] or xc_top.ixcSimTime[60]
 or xc_top.ixcSimTime[59] or xc_top.ixcSimTime[58] or xc_top.ixcSimTime[57] or xc_top.ixcSimTime[56] or xc_top.ixcSimTime[55] or xc_top.ixcSimTime[54] or xc_top.ixcSimTime[53] or xc_top.ixcSimTime[52]
 or xc_top.ixcSimTime[51] or xc_top.ixcSimTime[50] or xc_top.ixcSimTime[49] or xc_top.ixcSimTime[48] or xc_top.ixcSimTime[47] or xc_top.ixcSimTime[46] or xc_top.ixcSimTime[45] or xc_top.ixcSimTime[44]
 or xc_top.ixcSimTime[43] or xc_top.ixcSimTime[42] or xc_top.ixcSimTime[41] or xc_top.ixcSimTime[40] or xc_top.ixcSimTime[39] or xc_top.ixcSimTime[38] or xc_top.ixcSimTime[37] or xc_top.ixcSimTime[36]
 or xc_top.ixcSimTime[35] or xc_top.ixcSimTime[34] or xc_top.ixcSimTime[33] or xc_top.ixcSimTime[32] or xc_top.ixcSimTime[31] or xc_top.ixcSimTime[30] or xc_top.ixcSimTime[29] or xc_top.ixcSimTime[28]
 or xc_top.ixcSimTime[27] or xc_top.ixcSimTime[26] or xc_top.ixcSimTime[25] or xc_top.ixcSimTime[24] or xc_top.ixcSimTime[23] or xc_top.ixcSimTime[22] or xc_top.ixcSimTime[21] or xc_top.ixcSimTime[20]
 or xc_top.ixcSimTime[19] or xc_top.ixcSimTime[18] or xc_top.ixcSimTime[17] or xc_top.ixcSimTime[16] or xc_top.ixcSimTime[15] or xc_top.ixcSimTime[14] or xc_top.ixcSimTime[13] or xc_top.ixcSimTime[12]
 or xc_top.ixcSimTime[11] or xc_top.ixcSimTime[10] or xc_top.ixcSimTime[9] or xc_top.ixcSimTime[8] or xc_top.ixcSimTime[7] or xc_top.ixcSimTime[6] or xc_top.ixcSimTime[5] or xc_top.ixcSimTime[4]
 or xc_top.ixcSimTime[3] or xc_top.ixcSimTime[2] or xc_top.ixcSimTime[1] or xc_top.ixcSimTime[0] or xc_top.tbcPO or ackId[7] or ackId[6] or ackId[5]
 or ackId[4] or ackId[3] or ackId[2] or ackId[1] or ackId[0])
#0 begin
if (n1572)
ixc_gfm_ctl[{n1611, n1611}] =
{wrtCntD[62], wrtCntD[61], wrtCntD[60], wrtCntD[59], wrtCntD[58],
 wrtCntD[57], wrtCntD[56], wrtCntD[55], wrtCntD[54], wrtCntD[53], wrtCntD[52], wrtCntD[51], wrtCntD[50],
 wrtCntD[49], wrtCntD[48], wrtCntD[47], wrtCntD[46], wrtCntD[45], wrtCntD[44], wrtCntD[43], wrtCntD[42],
 wrtCntD[41], wrtCntD[40], wrtCntD[39], wrtCntD[38], wrtCntD[37], wrtCntD[36], wrtCntD[35], wrtCntD[34],
 wrtCntD[33], wrtCntD[32], wrtCntD[31], wrtCntD[30], wrtCntD[29], wrtCntD[28], wrtCntD[27], wrtCntD[26],
 wrtCntD[25], wrtCntD[24], wrtCntD[23], wrtCntD[22], wrtCntD[21], wrtCntD[20], wrtCntD[19], wrtCntD[18],
 wrtCntD[17], wrtCntD[16], wrtCntD[15], wrtCntD[14], wrtCntD[13], wrtCntD[12], wrtCntD[11], wrtCntD[10],
 wrtCntD[9], wrtCntD[8], wrtCntD[7], wrtCntD[6], wrtCntD[5], wrtCntD[4], wrtCntD[3], wrtCntD[2],
 wrtCntD[1], wrtCntD[0], xc_top.svGFbusy};
if (n1572)
ixc_gfm_ctl[{n1611, n1572}] =
{rdCnt[63], rdCnt[62], rdCnt[61], rdCnt[60], rdCnt[59],
 rdCnt[58], rdCnt[57], rdCnt[56], rdCnt[55], rdCnt[54], rdCnt[53], rdCnt[52], rdCnt[51],
 rdCnt[50], rdCnt[49], rdCnt[48], rdCnt[47], rdCnt[46], rdCnt[45], rdCnt[44], rdCnt[43],
 rdCnt[42], rdCnt[41], rdCnt[40], rdCnt[39], rdCnt[38], rdCnt[37], rdCnt[36], rdCnt[35],
 rdCnt[34], rdCnt[33], rdCnt[32], rdCnt[31], rdCnt[30], rdCnt[29], rdCnt[28], rdCnt[27],
 rdCnt[26], rdCnt[25], rdCnt[24], rdCnt[23], rdCnt[22], rdCnt[21], rdCnt[20], rdCnt[19],
 rdCnt[18], rdCnt[17], rdCnt[16], rdCnt[15], rdCnt[14], rdCnt[13], rdCnt[12], rdCnt[11],
 rdCnt[10], rdCnt[9], rdCnt[8], rdCnt[7], rdCnt[6], rdCnt[5], rdCnt[4], rdCnt[3],
 rdCnt[2], rdCnt[1], rdCnt[0]};
if (n1572)
ixc_gfm_ctl[{n1572, n1611}] =
{xc_top.ixcSimTime[62], xc_top.ixcSimTime[61], xc_top.ixcSimTime[60], xc_top.ixcSimTime[59], xc_top.ixcSimTime[58],
 xc_top.ixcSimTime[57], xc_top.ixcSimTime[56], xc_top.ixcSimTime[55], xc_top.ixcSimTime[54], xc_top.ixcSimTime[53], xc_top.ixcSimTime[52], xc_top.ixcSimTime[51], xc_top.ixcSimTime[50],
 xc_top.ixcSimTime[49], xc_top.ixcSimTime[48], xc_top.ixcSimTime[47], xc_top.ixcSimTime[46], xc_top.ixcSimTime[45], xc_top.ixcSimTime[44], xc_top.ixcSimTime[43], xc_top.ixcSimTime[42],
 xc_top.ixcSimTime[41], xc_top.ixcSimTime[40], xc_top.ixcSimTime[39], xc_top.ixcSimTime[38], xc_top.ixcSimTime[37], xc_top.ixcSimTime[36], xc_top.ixcSimTime[35], xc_top.ixcSimTime[34],
 xc_top.ixcSimTime[33], xc_top.ixcSimTime[32], xc_top.ixcSimTime[31], xc_top.ixcSimTime[30], xc_top.ixcSimTime[29], xc_top.ixcSimTime[28], xc_top.ixcSimTime[27], xc_top.ixcSimTime[26],
 xc_top.ixcSimTime[25], xc_top.ixcSimTime[24], xc_top.ixcSimTime[23], xc_top.ixcSimTime[22], xc_top.ixcSimTime[21], xc_top.ixcSimTime[20], xc_top.ixcSimTime[19], xc_top.ixcSimTime[18],
 xc_top.ixcSimTime[17], xc_top.ixcSimTime[16], xc_top.ixcSimTime[15], xc_top.ixcSimTime[14], xc_top.ixcSimTime[13], xc_top.ixcSimTime[12], xc_top.ixcSimTime[11], xc_top.ixcSimTime[10],
 xc_top.ixcSimTime[9], xc_top.ixcSimTime[8], xc_top.ixcSimTime[7], xc_top.ixcSimTime[6], xc_top.ixcSimTime[5], xc_top.ixcSimTime[4], xc_top.ixcSimTime[3], xc_top.ixcSimTime[2],
 xc_top.ixcSimTime[1], xc_top.ixcSimTime[0], xc_top.tbcPO};
if (n1572)
ixc_gfm_ctl[{n1572, n1572}] =
{n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, n1611, n1611, n1611, n1611, n1611,
 n1611, n1611, n1611, ackId[7], ackId[6], ackId[5], ackId[4], ackId[3],
 ackId[2], ackId[1], ackId[0]};
end
`else

MPW4X64 ixc_gfm_ctl ( .A1(n1611), .A0(n1611), .DI63(wrtCntD[62]), .DI62(wrtCntD[61]), .DI61(wrtCntD[60]), .DI60(wrtCntD[59]),
 .DI59(wrtCntD[58]), .DI58(wrtCntD[57]), .DI57(wrtCntD[56]), .DI56(wrtCntD[55]), .DI55(wrtCntD[54]), .DI54(wrtCntD[53]), .DI53(wrtCntD[52]), .DI52(wrtCntD[51]),
 .DI51(wrtCntD[50]), .DI50(wrtCntD[49]), .DI49(wrtCntD[48]), .DI48(wrtCntD[47]), .DI47(wrtCntD[46]), .DI46(wrtCntD[45]), .DI45(wrtCntD[44]), .DI44(wrtCntD[43]),
 .DI43(wrtCntD[42]), .DI42(wrtCntD[41]), .DI41(wrtCntD[40]), .DI40(wrtCntD[39]), .DI39(wrtCntD[38]), .DI38(wrtCntD[37]), .DI37(wrtCntD[36]), .DI36(wrtCntD[35]),
 .DI35(wrtCntD[34]), .DI34(wrtCntD[33]), .DI33(wrtCntD[32]), .DI32(wrtCntD[31]), .DI31(wrtCntD[30]), .DI30(wrtCntD[29]), .DI29(wrtCntD[28]), .DI28(wrtCntD[27]),
 .DI27(wrtCntD[26]), .DI26(wrtCntD[25]), .DI25(wrtCntD[24]), .DI24(wrtCntD[23]), .DI23(wrtCntD[22]), .DI22(wrtCntD[21]), .DI21(wrtCntD[20]), .DI20(wrtCntD[19]),
 .DI19(wrtCntD[18]), .DI18(wrtCntD[17]), .DI17(wrtCntD[16]), .DI16(wrtCntD[15]), .DI15(wrtCntD[14]), .DI14(wrtCntD[13]), .DI13(wrtCntD[12]), .DI12(wrtCntD[11]),
 .DI11(wrtCntD[10]), .DI10(wrtCntD[9]), .DI9(wrtCntD[8]), .DI8(wrtCntD[7]), .DI7(wrtCntD[6]), .DI6(wrtCntD[5]), .DI5(wrtCntD[4]), .DI4(wrtCntD[3]),
 .DI3(wrtCntD[2]), .DI2(wrtCntD[1]), .DI1(wrtCntD[0]), .DI0(xc_top.svGFbusy), .WE(n1572), .SYNC_IN(n1611), .SYNC_OUT(n6744));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ctl" HDL_MEMORY_DECL "1 63 0 0 3"
MPW4X64 U9489 ( .A1(n1611), .A0(n1572), .DI63(rdCnt[63]), .DI62(rdCnt[62]), .DI61(rdCnt[61]), .DI60(rdCnt[60]),
 .DI59(rdCnt[59]), .DI58(rdCnt[58]), .DI57(rdCnt[57]), .DI56(rdCnt[56]), .DI55(rdCnt[55]), .DI54(rdCnt[54]), .DI53(rdCnt[53]), .DI52(rdCnt[52]),
 .DI51(rdCnt[51]), .DI50(rdCnt[50]), .DI49(rdCnt[49]), .DI48(rdCnt[48]), .DI47(rdCnt[47]), .DI46(rdCnt[46]), .DI45(rdCnt[45]), .DI44(rdCnt[44]),
 .DI43(rdCnt[43]), .DI42(rdCnt[42]), .DI41(rdCnt[41]), .DI40(rdCnt[40]), .DI39(rdCnt[39]), .DI38(rdCnt[38]), .DI37(rdCnt[37]), .DI36(rdCnt[36]),
 .DI35(rdCnt[35]), .DI34(rdCnt[34]), .DI33(rdCnt[33]), .DI32(rdCnt[32]), .DI31(rdCnt[31]), .DI30(rdCnt[30]), .DI29(rdCnt[29]), .DI28(rdCnt[28]),
 .DI27(rdCnt[27]), .DI26(rdCnt[26]), .DI25(rdCnt[25]), .DI24(rdCnt[24]), .DI23(rdCnt[23]), .DI22(rdCnt[22]), .DI21(rdCnt[21]), .DI20(rdCnt[20]),
 .DI19(rdCnt[19]), .DI18(rdCnt[18]), .DI17(rdCnt[17]), .DI16(rdCnt[16]), .DI15(rdCnt[15]), .DI14(rdCnt[14]), .DI13(rdCnt[13]), .DI12(rdCnt[12]),
 .DI11(rdCnt[11]), .DI10(rdCnt[10]), .DI9(rdCnt[9]), .DI8(rdCnt[8]), .DI7(rdCnt[7]), .DI6(rdCnt[6]), .DI5(rdCnt[5]), .DI4(rdCnt[4]),
 .DI3(rdCnt[3]), .DI2(rdCnt[2]), .DI1(rdCnt[1]), .DI0(rdCnt[0]), .WE(n1572), .SYNC_IN(n6744), .SYNC_OUT(n6745));
MPW4X64 U9490 ( .A1(n1572), .A0(n1611), .DI63(xc_top.ixcSimTime[62]), .DI62(xc_top.ixcSimTime[61]), .DI61(xc_top.ixcSimTime[60]), .DI60(xc_top.ixcSimTime[59]),
 .DI59(xc_top.ixcSimTime[58]), .DI58(xc_top.ixcSimTime[57]), .DI57(xc_top.ixcSimTime[56]), .DI56(xc_top.ixcSimTime[55]), .DI55(xc_top.ixcSimTime[54]), .DI54(xc_top.ixcSimTime[53]), .DI53(xc_top.ixcSimTime[52]), .DI52(xc_top.ixcSimTime[51]),
 .DI51(xc_top.ixcSimTime[50]), .DI50(xc_top.ixcSimTime[49]), .DI49(xc_top.ixcSimTime[48]), .DI48(xc_top.ixcSimTime[47]), .DI47(xc_top.ixcSimTime[46]), .DI46(xc_top.ixcSimTime[45]), .DI45(xc_top.ixcSimTime[44]), .DI44(xc_top.ixcSimTime[43]),
 .DI43(xc_top.ixcSimTime[42]), .DI42(xc_top.ixcSimTime[41]), .DI41(xc_top.ixcSimTime[40]), .DI40(xc_top.ixcSimTime[39]), .DI39(xc_top.ixcSimTime[38]), .DI38(xc_top.ixcSimTime[37]), .DI37(xc_top.ixcSimTime[36]), .DI36(xc_top.ixcSimTime[35]),
 .DI35(xc_top.ixcSimTime[34]), .DI34(xc_top.ixcSimTime[33]), .DI33(xc_top.ixcSimTime[32]), .DI32(xc_top.ixcSimTime[31]), .DI31(xc_top.ixcSimTime[30]), .DI30(xc_top.ixcSimTime[29]), .DI29(xc_top.ixcSimTime[28]), .DI28(xc_top.ixcSimTime[27]),
 .DI27(xc_top.ixcSimTime[26]), .DI26(xc_top.ixcSimTime[25]), .DI25(xc_top.ixcSimTime[24]), .DI24(xc_top.ixcSimTime[23]), .DI23(xc_top.ixcSimTime[22]), .DI22(xc_top.ixcSimTime[21]), .DI21(xc_top.ixcSimTime[20]), .DI20(xc_top.ixcSimTime[19]),
 .DI19(xc_top.ixcSimTime[18]), .DI18(xc_top.ixcSimTime[17]), .DI17(xc_top.ixcSimTime[16]), .DI16(xc_top.ixcSimTime[15]), .DI15(xc_top.ixcSimTime[14]), .DI14(xc_top.ixcSimTime[13]), .DI13(xc_top.ixcSimTime[12]), .DI12(xc_top.ixcSimTime[11]),
 .DI11(xc_top.ixcSimTime[10]), .DI10(xc_top.ixcSimTime[9]), .DI9(xc_top.ixcSimTime[8]), .DI8(xc_top.ixcSimTime[7]), .DI7(xc_top.ixcSimTime[6]), .DI6(xc_top.ixcSimTime[5]), .DI5(xc_top.ixcSimTime[4]), .DI4(xc_top.ixcSimTime[3]),
 .DI3(xc_top.ixcSimTime[2]), .DI2(xc_top.ixcSimTime[1]), .DI1(xc_top.ixcSimTime[0]), .DI0(xc_top.tbcPO), .WE(n1572), .SYNC_IN(n6745), .SYNC_OUT(n6746));
MPW4X64 U9491 ( .A1(n1572), .A0(n1572), .DI63(n1611), .DI62(n1611), .DI61(n1611), .DI60(n1611),
 .DI59(n1611), .DI58(n1611), .DI57(n1611), .DI56(n1611), .DI55(n1611), .DI54(n1611), .DI53(n1611), .DI52(n1611),
 .DI51(n1611), .DI50(n1611), .DI49(n1611), .DI48(n1611), .DI47(n1611), .DI46(n1611), .DI45(n1611), .DI44(n1611),
 .DI43(n1611), .DI42(n1611), .DI41(n1611), .DI40(n1611), .DI39(n1611), .DI38(n1611), .DI37(n1611), .DI36(n1611),
 .DI35(n1611), .DI34(n1611), .DI33(n1611), .DI32(n1611), .DI31(n1611), .DI30(n1611), .DI29(n1611), .DI28(n1611),
 .DI27(n1611), .DI26(n1611), .DI25(n1611), .DI24(n1611), .DI23(n1611), .DI22(n1611), .DI21(n1611), .DI20(n1611),
 .DI19(n1611), .DI18(n1611), .DI17(n1611), .DI16(n1611), .DI15(n1611), .DI14(n1611), .DI13(n1611), .DI12(n1611),
 .DI11(n1611), .DI10(n1611), .DI9(n1611), .DI8(n1611), .DI7(ackId[7]), .DI6(ackId[6]), .DI5(ackId[5]), .DI4(ackId[4]),
 .DI3(ackId[3]), .DI2(ackId[2]), .DI1(ackId[1]), .DI0(ackId[0]), .WE(n1572), .SYNC_IN(n6746), .SYNC_OUT( ));
`endif
`ifdef CBV

reg [63:0] ixc_gfm_ack [0:0];
initial begin: U9492
  integer j;
  for (j=0; j<=0; j=j+1) ixc_gfm_ack[j] =
`ifdef CBV_MEM_INIT1
  {64{1'b1}};
`else
  64'b0;
`endif
end
reg [63:0] n6747;
buf(ackLen[17], n6747[25]);
buf(ackLen[16], n6747[24]);
buf(ackLen[15], n6747[23]);
buf(ackLen[14], n6747[22]);
buf(ackLen[13], n6747[21]);
buf(ackLen[12], n6747[20]);
buf(ackLen[11], n6747[19]);
buf(ackLen[10], n6747[18]);
buf(ackLen[9], n6747[17]);
buf(ackLen[8], n6747[16]);
buf(ackLen[7], n6747[15]);
buf(ackLen[6], n6747[14]);
buf(ackLen[5], n6747[13]);
buf(ackLen[4], n6747[12]);
buf(ackLen[3], n6747[11]);
buf(ackLen[2], n6747[10]);
buf(ackLen[1], n6747[9]);
buf(ackLen[0], n6747[8]);
buf(ackIdNew[7], n6747[7]);
buf(ackIdNew[6], n6747[6]);
buf(ackIdNew[5], n6747[5]);
buf(ackIdNew[4], n6747[4]);
buf(ackIdNew[3], n6747[3]);
buf(ackIdNew[2], n6747[2]);
buf(ackIdNew[1], n6747[1]);
buf(ackIdNew[0], n6747[0]);
always @(n1611)
#0 begin
n6747 = ixc_gfm_ack[{n1611}];
end
`else

MPR2X64 ixc_gfm_ack ( .A0(n1611), .SYNC_IN(n1611), .DO63( ), .DO62( ), .DO61( ), .DO60( ),
 .DO59( ), .DO58( ), .DO57( ), .DO56( ), .DO55( ), .DO54( ), .DO53( ), .DO52( ),
 .DO51( ), .DO50( ), .DO49( ), .DO48( ), .DO47( ), .DO46( ), .DO45( ), .DO44( ),
 .DO43( ), .DO42( ), .DO41( ), .DO40( ), .DO39( ), .DO38( ), .DO37( ), .DO36( ),
 .DO35( ), .DO34( ), .DO33( ), .DO32( ), .DO31( ), .DO30( ), .DO29( ), .DO28( ),
 .DO27( ), .DO26( ), .DO25(ackLen[17]), .DO24(ackLen[16]), .DO23(ackLen[15]), .DO22(ackLen[14]), .DO21(ackLen[13]), .DO20(ackLen[12]),
 .DO19(ackLen[11]), .DO18(ackLen[10]), .DO17(ackLen[9]), .DO16(ackLen[8]), .DO15(ackLen[7]), .DO14(ackLen[6]), .DO13(ackLen[5]), .DO12(ackLen[4]),
 .DO11(ackLen[3]), .DO10(ackLen[2]), .DO9(ackLen[1]), .DO8(ackLen[0]), .DO7(ackIdNew[7]), .DO6(ackIdNew[6]), .DO5(ackIdNew[5]), .DO4(ackIdNew[4]),
 .DO3(ackIdNew[3]), .DO2(ackIdNew[2]), .DO1(ackIdNew[1]), .DO0(ackIdNew[0]), .SYNC_OUT( ));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ack" HDL_MEMORY_DECL "1 63 0 0 0"
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "TsBuf 1 64 0 0 7"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "ixc_gfm_ofifo 1 255 0 0 32767"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "ixc_gfm_ctl 1 63 0 0 3"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "ixc_gfm_ack 1 63 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "3"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW2X64_MPR2X64
`else
module MPW2X64( A0, DI63, DI62, DI61, DI60, DI59, DI58,
 DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42,
 DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34,
 DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26,
 DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18,
 DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2,
 DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A0, DI63, DI62, DI61, DI60, DI59, DI58, DI57,
 DI56, DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48, DI47,
 DI46, DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37,
 DI36, DI35, DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18, DI17,
 DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8, DI7,
 DI6, DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR2X64_
`else
module MPR2X64( A0, SYNC_IN, DO63, DO62, DO61, DO60, DO59,
 DO58, DO57, DO56, DO55, DO54, DO53, DO52, DO51,
 DO50, DO49, DO48, DO47, DO46, DO45, DO44, DO43,
 DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35,
 DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27,
 DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19,
 DO18, DO17, DO16, DO15, DO14, DO13, DO12, DO11,
 DO10, DO9, DO8, DO7, DO6, DO5, DO4, DO3,
 DO2, DO1, DO0, SYNC_OUT);
input  A0, SYNC_IN;
output  DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56,
 DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26,
 DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16,
 DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR2X64_
`endif
`define MPW2X64_MPR2X64
`endif
`ifdef MPW4X64_MPR4X64
`else
module MPW4X64( A1, A0, DI63, DI62, DI61, DI60, DI59,
 DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51,
 DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19,
 DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11,
 DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A1, A0, DI63, DI62, DI61, DI60, DI59, DI58,
 DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48,
 DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38,
 DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30, DI29, DI28,
 DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18,
 DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8,
 DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR4X64_
`else
module MPR4X64( A1, A0, SYNC_IN, DO63, DO62, DO61, DO60,
 DO59, DO58, DO57, DO56, DO55, DO54, DO53, DO52,
 DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12,
 DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT);
input  A1, A0, SYNC_IN;
output  DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56,
 DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26,
 DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16,
 DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR4X64_
`endif
`define MPW4X64_MPR4X64
`endif
`ifdef MPW32KX256_MPR32KX256
`else
module MPW32KX256( A14, A13, A12, A11, A10, A9, A8,
 A7, A6, A5, A4, A3, A2, A1, A0,
 DI255, DI254, DI253, DI252, DI251, DI250, DI249, DI248,
 DI247, DI246, DI245, DI244, DI243, DI242, DI241, DI240,
 DI239, DI238, DI237, DI236, DI235, DI234, DI233, DI232,
 DI231, DI230, DI229, DI228, DI227, DI226, DI225, DI224,
 DI223, DI222, DI221, DI220, DI219, DI218, DI217, DI216,
 DI215, DI214, DI213, DI212, DI211, DI210, DI209, DI208,
 DI207, DI206, DI205, DI204, DI203, DI202, DI201, DI200,
 DI199, DI198, DI197, DI196, DI195, DI194, DI193, DI192,
 DI191, DI190, DI189, DI188, DI187, DI186, DI185, DI184,
 DI183, DI182, DI181, DI180, DI179, DI178, DI177, DI176,
 DI175, DI174, DI173, DI172, DI171, DI170, DI169, DI168,
 DI167, DI166, DI165, DI164, DI163, DI162, DI161, DI160,
 DI159, DI158, DI157, DI156, DI155, DI154, DI153, DI152,
 DI151, DI150, DI149, DI148, DI147, DI146, DI145, DI144,
 DI143, DI142, DI141, DI140, DI139, DI138, DI137, DI136,
 DI135, DI134, DI133, DI132, DI131, DI130, DI129, DI128,
 DI127, DI126, DI125, DI124, DI123, DI122, DI121, DI120,
 DI119, DI118, DI117, DI116, DI115, DI114, DI113, DI112,
 DI111, DI110, DI109, DI108, DI107, DI106, DI105, DI104,
 DI103, DI102, DI101, DI100, DI99, DI98, DI97, DI96,
 DI95, DI94, DI93, DI92, DI91, DI90, DI89, DI88,
 DI87, DI86, DI85, DI84, DI83, DI82, DI81, DI80,
 DI79, DI78, DI77, DI76, DI75, DI74, DI73, DI72,
 DI71, DI70, DI69, DI68, DI67, DI66, DI65, DI64,
 DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56,
 DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48,
 DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32,
 DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24,
 DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16,
 DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8,
 DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN, SYNC_OUT);
input  A14, A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, DI255, DI254, DI253,
 DI252, DI251, DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235, DI234, DI233,
 DI232, DI231, DI230, DI229, DI228, DI227, DI226, DI225, DI224, DI223,
 DI222, DI221, DI220, DI219, DI218, DI217, DI216, DI215, DI214, DI213,
 DI212, DI211, DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195, DI194, DI193,
 DI192, DI191, DI190, DI189, DI188, DI187, DI186, DI185, DI184, DI183,
 DI182, DI181, DI180, DI179, DI178, DI177, DI176, DI175, DI174, DI173,
 DI172, DI171, DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155, DI154, DI153,
 DI152, DI151, DI150, DI149, DI148, DI147, DI146, DI145, DI144, DI143,
 DI142, DI141, DI140, DI139, DI138, DI137, DI136, DI135, DI134, DI133,
 DI132, DI131, DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115, DI114, DI113,
 DI112, DI111, DI110, DI109, DI108, DI107, DI106, DI105, DI104, DI103,
 DI102, DI101, DI100, DI99, DI98, DI97, DI96, DI95, DI94, DI93,
 DI92, DI91, DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75, DI74, DI73,
 DI72, DI71, DI70, DI69, DI68, DI67, DI66, DI65, DI64, DI63,
 DI62, DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54, DI53,
 DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34, DI33,
 DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24, DI23,
 DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR32KX256_
`else
module MPR32KX256( A14, A13, A12, A11, A10, A9, A8,
 A7, A6, A5, A4, A3, A2, A1, A0,
 SYNC_IN, DO255, DO254, DO253, DO252, DO251, DO250, DO249,
 DO248, DO247, DO246, DO245, DO244, DO243, DO242, DO241,
 DO240, DO239, DO238, DO237, DO236, DO235, DO234, DO233,
 DO232, DO231, DO230, DO229, DO228, DO227, DO226, DO225,
 DO224, DO223, DO222, DO221, DO220, DO219, DO218, DO217,
 DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209,
 DO208, DO207, DO206, DO205, DO204, DO203, DO202, DO201,
 DO200, DO199, DO198, DO197, DO196, DO195, DO194, DO193,
 DO192, DO191, DO190, DO189, DO188, DO187, DO186, DO185,
 DO184, DO183, DO182, DO181, DO180, DO179, DO178, DO177,
 DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169,
 DO168, DO167, DO166, DO165, DO164, DO163, DO162, DO161,
 DO160, DO159, DO158, DO157, DO156, DO155, DO154, DO153,
 DO152, DO151, DO150, DO149, DO148, DO147, DO146, DO145,
 DO144, DO143, DO142, DO141, DO140, DO139, DO138, DO137,
 DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129,
 DO128, DO127, DO126, DO125, DO124, DO123, DO122, DO121,
 DO120, DO119, DO118, DO117, DO116, DO115, DO114, DO113,
 DO112, DO111, DO110, DO109, DO108, DO107, DO106, DO105,
 DO104, DO103, DO102, DO101, DO100, DO99, DO98, DO97,
 DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89,
 DO88, DO87, DO86, DO85, DO84, DO83, DO82, DO81,
 DO80, DO79, DO78, DO77, DO76, DO75, DO74, DO73,
 DO72, DO71, DO70, DO69, DO68, DO67, DO66, DO65,
 DO64, DO63, DO62, DO61, DO60, DO59, DO58, DO57,
 DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49,
 DO48, DO47, DO46, DO45, DO44, DO43, DO42, DO41,
 DO40, DO39, DO38, DO37, DO36, DO35, DO34, DO33,
 DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25,
 DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17,
 DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9,
 DO8, DO7, DO6, DO5, DO4, DO3, DO2, DO1,
 DO0, SYNC_OUT);
input  A14, A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, SYNC_IN;
output  DO255, DO254, DO253, DO252, DO251, DO250, DO249, DO248,
 DO247, DO246, DO245, DO244, DO243, DO242, DO241, DO240, DO239, DO238,
 DO237, DO236, DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220, DO219, DO218,
 DO217, DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209, DO208,
 DO207, DO206, DO205, DO204, DO203, DO202, DO201, DO200, DO199, DO198,
 DO197, DO196, DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180, DO179, DO178,
 DO177, DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169, DO168,
 DO167, DO166, DO165, DO164, DO163, DO162, DO161, DO160, DO159, DO158,
 DO157, DO156, DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140, DO139, DO138,
 DO137, DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129, DO128,
 DO127, DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119, DO118,
 DO117, DO116, DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99, DO98,
 DO97, DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89, DO88,
 DO87, DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79, DO78,
 DO77, DO76, DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59, DO58,
 DO57, DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48,
 DO47, DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18,
 DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8,
 DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR32KX256_
`endif
`define MPW32KX256_MPR32KX256
`endif
`endif
