
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_ckv_reader ( ckvreader_kimreader_ack, ckvreader_kopassigner_valid, 
	.ckvreader_kopassigner_data( {\ckvreader_kopassigner_data.sot [0], 
	\ckvreader_kopassigner_data.eoi [0], 
	\ckvreader_kopassigner_data.eot [0], 
	\ckvreader_kopassigner_data.id [3], 
	\ckvreader_kopassigner_data.id [2], 
	\ckvreader_kopassigner_data.id [1], 
	\ckvreader_kopassigner_data.id [0], 
	\ckvreader_kopassigner_data.tdata [63], 
	\ckvreader_kopassigner_data.tdata [62], 
	\ckvreader_kopassigner_data.tdata [61], 
	\ckvreader_kopassigner_data.tdata [60], 
	\ckvreader_kopassigner_data.tdata [59], 
	\ckvreader_kopassigner_data.tdata [58], 
	\ckvreader_kopassigner_data.tdata [57], 
	\ckvreader_kopassigner_data.tdata [56], 
	\ckvreader_kopassigner_data.tdata [55], 
	\ckvreader_kopassigner_data.tdata [54], 
	\ckvreader_kopassigner_data.tdata [53], 
	\ckvreader_kopassigner_data.tdata [52], 
	\ckvreader_kopassigner_data.tdata [51], 
	\ckvreader_kopassigner_data.tdata [50], 
	\ckvreader_kopassigner_data.tdata [49], 
	\ckvreader_kopassigner_data.tdata [48], 
	\ckvreader_kopassigner_data.tdata [47], 
	\ckvreader_kopassigner_data.tdata [46], 
	\ckvreader_kopassigner_data.tdata [45], 
	\ckvreader_kopassigner_data.tdata [44], 
	\ckvreader_kopassigner_data.tdata [43], 
	\ckvreader_kopassigner_data.tdata [42], 
	\ckvreader_kopassigner_data.tdata [41], 
	\ckvreader_kopassigner_data.tdata [40], 
	\ckvreader_kopassigner_data.tdata [39], 
	\ckvreader_kopassigner_data.tdata [38], 
	\ckvreader_kopassigner_data.tdata [37], 
	\ckvreader_kopassigner_data.tdata [36], 
	\ckvreader_kopassigner_data.tdata [35], 
	\ckvreader_kopassigner_data.tdata [34], 
	\ckvreader_kopassigner_data.tdata [33], 
	\ckvreader_kopassigner_data.tdata [32], 
	\ckvreader_kopassigner_data.tdata [31], 
	\ckvreader_kopassigner_data.tdata [30], 
	\ckvreader_kopassigner_data.tdata [29], 
	\ckvreader_kopassigner_data.tdata [28], 
	\ckvreader_kopassigner_data.tdata [27], 
	\ckvreader_kopassigner_data.tdata [26], 
	\ckvreader_kopassigner_data.tdata [25], 
	\ckvreader_kopassigner_data.tdata [24], 
	\ckvreader_kopassigner_data.tdata [23], 
	\ckvreader_kopassigner_data.tdata [22], 
	\ckvreader_kopassigner_data.tdata [21], 
	\ckvreader_kopassigner_data.tdata [20], 
	\ckvreader_kopassigner_data.tdata [19], 
	\ckvreader_kopassigner_data.tdata [18], 
	\ckvreader_kopassigner_data.tdata [17], 
	\ckvreader_kopassigner_data.tdata [16], 
	\ckvreader_kopassigner_data.tdata [15], 
	\ckvreader_kopassigner_data.tdata [14], 
	\ckvreader_kopassigner_data.tdata [13], 
	\ckvreader_kopassigner_data.tdata [12], 
	\ckvreader_kopassigner_data.tdata [11], 
	\ckvreader_kopassigner_data.tdata [10], 
	\ckvreader_kopassigner_data.tdata [9], 
	\ckvreader_kopassigner_data.tdata [8], 
	\ckvreader_kopassigner_data.tdata [7], 
	\ckvreader_kopassigner_data.tdata [6], 
	\ckvreader_kopassigner_data.tdata [5], 
	\ckvreader_kopassigner_data.tdata [4], 
	\ckvreader_kopassigner_data.tdata [3], 
	\ckvreader_kopassigner_data.tdata [2], 
	\ckvreader_kopassigner_data.tdata [1], 
	\ckvreader_kopassigner_data.tdata [0]} ), ckv_rd, ckv_addr, clk, 
	rst_n, kimreader_ckvreader_valid, .kimreader_ckvreader_data( {
	\kimreader_ckvreader_data.sot [0], \kimreader_ckvreader_data.eoi [0], 
	\kimreader_ckvreader_data.eot [0], \kimreader_ckvreader_data.id [3], 
	\kimreader_ckvreader_data.id [2], \kimreader_ckvreader_data.id [1], 
	\kimreader_ckvreader_data.id [0], 
	\kimreader_ckvreader_data.tdata [63], 
	\kimreader_ckvreader_data.tdata [62], 
	\kimreader_ckvreader_data.tdata [61], 
	\kimreader_ckvreader_data.tdata [60], 
	\kimreader_ckvreader_data.tdata [59], 
	\kimreader_ckvreader_data.tdata [58], 
	\kimreader_ckvreader_data.tdata [57], 
	\kimreader_ckvreader_data.tdata [56], 
	\kimreader_ckvreader_data.tdata [55], 
	\kimreader_ckvreader_data.tdata [54], 
	\kimreader_ckvreader_data.tdata [53], 
	\kimreader_ckvreader_data.tdata [52], 
	\kimreader_ckvreader_data.tdata [51], 
	\kimreader_ckvreader_data.tdata [50], 
	\kimreader_ckvreader_data.tdata [49], 
	\kimreader_ckvreader_data.tdata [48], 
	\kimreader_ckvreader_data.tdata [47], 
	\kimreader_ckvreader_data.tdata [46], 
	\kimreader_ckvreader_data.tdata [45], 
	\kimreader_ckvreader_data.tdata [44], 
	\kimreader_ckvreader_data.tdata [43], 
	\kimreader_ckvreader_data.tdata [42], 
	\kimreader_ckvreader_data.tdata [41], 
	\kimreader_ckvreader_data.tdata [40], 
	\kimreader_ckvreader_data.tdata [39], 
	\kimreader_ckvreader_data.tdata [38], 
	\kimreader_ckvreader_data.tdata [37], 
	\kimreader_ckvreader_data.tdata [36], 
	\kimreader_ckvreader_data.tdata [35], 
	\kimreader_ckvreader_data.tdata [34], 
	\kimreader_ckvreader_data.tdata [33], 
	\kimreader_ckvreader_data.tdata [32], 
	\kimreader_ckvreader_data.tdata [31], 
	\kimreader_ckvreader_data.tdata [30], 
	\kimreader_ckvreader_data.tdata [29], 
	\kimreader_ckvreader_data.tdata [28], 
	\kimreader_ckvreader_data.tdata [27], 
	\kimreader_ckvreader_data.tdata [26], 
	\kimreader_ckvreader_data.tdata [25], 
	\kimreader_ckvreader_data.tdata [24], 
	\kimreader_ckvreader_data.tdata [23], 
	\kimreader_ckvreader_data.tdata [22], 
	\kimreader_ckvreader_data.tdata [21], 
	\kimreader_ckvreader_data.tdata [20], 
	\kimreader_ckvreader_data.tdata [19], 
	\kimreader_ckvreader_data.tdata [18], 
	\kimreader_ckvreader_data.tdata [17], 
	\kimreader_ckvreader_data.tdata [16], 
	\kimreader_ckvreader_data.tdata [15], 
	\kimreader_ckvreader_data.tdata [14], 
	\kimreader_ckvreader_data.tdata [13], 
	\kimreader_ckvreader_data.tdata [12], 
	\kimreader_ckvreader_data.tdata [11], 
	\kimreader_ckvreader_data.tdata [10], 
	\kimreader_ckvreader_data.tdata [9], 
	\kimreader_ckvreader_data.tdata [8], 
	\kimreader_ckvreader_data.tdata [7], 
	\kimreader_ckvreader_data.tdata [6], 
	\kimreader_ckvreader_data.tdata [5], 
	\kimreader_ckvreader_data.tdata [4], 
	\kimreader_ckvreader_data.tdata [3], 
	\kimreader_ckvreader_data.tdata [2], 
	\kimreader_ckvreader_data.tdata [1], 
	\kimreader_ckvreader_data.tdata [0]} ), kopassigner_ckvreader_ack, 
	ckv_dout, ckv_mbe);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output ckvreader_kimreader_ack;
output ckvreader_kopassigner_valid;
output [0:0] \ckvreader_kopassigner_data.sot ;
output [0:0] \ckvreader_kopassigner_data.eoi ;
output [0:0] \ckvreader_kopassigner_data.eot ;
output [3:0] \ckvreader_kopassigner_data.id ;
output [63:0] \ckvreader_kopassigner_data.tdata ;
wire [70:0] ckvreader_kopassigner_data;
output ckv_rd;
output [14:0] ckv_addr;
input clk;
input rst_n;
input kimreader_ckvreader_valid;
input [0:0] \kimreader_ckvreader_data.sot ;
input [0:0] \kimreader_ckvreader_data.eoi ;
input [0:0] \kimreader_ckvreader_data.eot ;
input [3:0] \kimreader_ckvreader_data.id ;
input [63:0] \kimreader_ckvreader_data.tdata ;
wire [70:0] kimreader_ckvreader_data;
input kopassigner_ckvreader_ack;
input [63:0] ckv_dout;
input ckv_mbe;
wire fifo_out_mbe;
wire [63:0] fifo_out;
wire fifo_out_valid;
wire fifo_in_stall;
wire _zy_simnet_ckvreader_kimreader_ack_0_w$;
wire _zy_simnet_ckvreader_kopassigner_valid_1_w$;
wire [0:70] _zy_simnet_ckvreader_kopassigner_data_2_w$;
wire _zy_simnet_ckv_rd_3_w$;
wire [0:14] _zy_simnet_ckv_addr_4_w$;
wire _zy_simnet_dio_5;
wire _zy_simnet_dio_6;
wire _zy_simnet_ckv_rd_q_7_w$;
wire _zy_simnet_fifo_out_ack_8_w$;
wire _zy_simnet_cio_9;
wire _zy_sva_brcm_dek_key_1_reset_or;
wire _zy_sva_brcm_dak_key_2_reset_or;
wire _zy_sva_brcm_dek_key_3_reset_or;
wire _zy_sva_brcm_dak_key_4_reset_or;
wire _zy_sva_brcm_dek_key_5_reset_or;
wire _zy_sva_brcm_dak_key_6_reset_or;
wire _zy_sva_brcm_dek_key_7_reset_or;
wire _zy_sva_brcm_dak_key_8_reset_or;
wire _zy_sva_b0_t;
wire _zy_sva_b1_t;
wire _zy_sva_b2_t;
wire _zy_sva_b3_t;
wire _zy_sva_b4_t;
wire _zy_sva_b5_t;
wire _zy_sva_b6_t;
wire _zy_sva_b7_t;
wire [0:0] cur_state;
wire [0:0] nxt_state;
wire ckv_rd_q;
wire half_dek;
wire [63:0] tlv_word0;
wire [55:0] tlv_word42;
wire [63:0] tlv_word8;
wire [63:0] nxt_tlv_word8;
wire [63:0] tlv_word9;
wire [63:0] nxt_tlv_word9;
wire [31:0] aux_key_ctrl;
wire fifo_out_ack;
wire report_kme_error;
wire [3:0] ckv_read_num;
wire ktype_is_aux_key_only;
wire nxt_ktype_is_aux_key_only;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_1_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_1_cpass;
`_2_ wire _zy_sva_b0;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_2_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_2_cpass;
`_2_ wire _zy_sva_b1;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_3_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_3_cpass;
`_2_ wire _zy_sva_b2;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_4_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_4_cpass;
`_2_ wire _zy_sva_b3;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_5_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_5_cpass;
`_2_ wire _zy_sva_b4;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_6_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_6_cpass;
`_2_ wire _zy_sva_b5;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_7_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dek_key_7_cpass;
`_2_ wire _zy_sva_b6;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_8_ccheck;
`_2_ wire [0:0] _zy_sva_brcm_dak_key_8_cpass;
`_2_ wire _zy_sva_b7;
supply1 n1;
supply0 n2;
wire [1:0] \tlv_word0.tlv_bip2 ;
wire [12:0] \tlv_word0.resv0 ;
wire [0:0] \tlv_word0.kdf_dek_iter ;
wire [0:0] \tlv_word0.keyless_algos ;
wire [0:0] \tlv_word0.needs_dek ;
wire [0:0] \tlv_word0.needs_dak ;
wire [5:0] \tlv_word0.key_type ;
wire [10:0] \tlv_word0.tlv_frame_num ;
wire [3:0] \tlv_word0.tlv_eng_id ;
wire [7:0] \tlv_word0.tlv_seq_num ;
wire [7:0] \tlv_word0.tlv_len ;
wire [7:0] \tlv_word0.tlv_type ;
wire [0:0] \tlv_word42.corrupt_crc32 ;
wire [46:0] \tlv_word42.unused ;
wire [7:0] \tlv_word42.error_code ;
wire [0:0] \tlv_word8.dek_kim_entry.valid ;
wire [2:0] \tlv_word8.dek_kim_entry.label_index ;
wire [1:0] \tlv_word8.dek_kim_entry.ckv_length ;
wire [14:0] \tlv_word8.dek_kim_entry.ckv_pointer ;
wire [3:0] \tlv_word8.dek_kim_entry.pf_num ;
wire [11:0] \tlv_word8.dek_kim_entry.vf_num ;
wire [0:0] \tlv_word8.dek_kim_entry.vf_valid ;
wire [5:0] \tlv_word8.unused ;
wire [0:0] \tlv_word8.missing_iv ;
wire [0:0] \tlv_word8.missing_guid ;
wire [0:0] \tlv_word8.validate_dek ;
wire [0:0] \tlv_word8.vf_valid ;
wire [3:0] \tlv_word8.pf_num ;
wire [11:0] \tlv_word8.vf_num ;
wire [0:0] \nxt_tlv_word8.dek_kim_entry.valid ;
wire [2:0] \nxt_tlv_word8.dek_kim_entry.label_index ;
wire [1:0] \nxt_tlv_word8.dek_kim_entry.ckv_length ;
wire [14:0] \nxt_tlv_word8.dek_kim_entry.ckv_pointer ;
wire [3:0] \nxt_tlv_word8.dek_kim_entry.pf_num ;
wire [11:0] \nxt_tlv_word8.dek_kim_entry.vf_num ;
wire [0:0] \nxt_tlv_word8.dek_kim_entry.vf_valid ;
wire [5:0] \nxt_tlv_word8.unused ;
wire [0:0] \nxt_tlv_word8.missing_iv ;
wire [0:0] \nxt_tlv_word8.missing_guid ;
wire [0:0] \nxt_tlv_word8.validate_dek ;
wire [0:0] \nxt_tlv_word8.vf_valid ;
wire [3:0] \nxt_tlv_word8.pf_num ;
wire [11:0] \nxt_tlv_word8.vf_num ;
wire [0:0] \tlv_word9.dak_kim_entry.valid ;
wire [2:0] \tlv_word9.dak_kim_entry.label_index ;
wire [1:0] \tlv_word9.dak_kim_entry.ckv_length ;
wire [14:0] \tlv_word9.dak_kim_entry.ckv_pointer ;
wire [3:0] \tlv_word9.dak_kim_entry.pf_num ;
wire [11:0] \tlv_word9.dak_kim_entry.vf_num ;
wire [0:0] \tlv_word9.dak_kim_entry.vf_valid ;
wire [7:0] \tlv_word9.unused ;
wire [0:0] \tlv_word9.validate_dak ;
wire [0:0] \tlv_word9.vf_valid ;
wire [3:0] \tlv_word9.pf_num ;
wire [11:0] \tlv_word9.vf_num ;
wire [0:0] \nxt_tlv_word9.dak_kim_entry.valid ;
wire [2:0] \nxt_tlv_word9.dak_kim_entry.label_index ;
wire [1:0] \nxt_tlv_word9.dak_kim_entry.ckv_length ;
wire [14:0] \nxt_tlv_word9.dak_kim_entry.ckv_pointer ;
wire [3:0] \nxt_tlv_word9.dak_kim_entry.pf_num ;
wire [11:0] \nxt_tlv_word9.dak_kim_entry.vf_num ;
wire [0:0] \nxt_tlv_word9.dak_kim_entry.vf_valid ;
wire [7:0] \nxt_tlv_word9.unused ;
wire [0:0] \nxt_tlv_word9.validate_dak ;
wire [0:0] \nxt_tlv_word9.vf_valid ;
wire [3:0] \nxt_tlv_word9.pf_num ;
wire [11:0] \nxt_tlv_word9.vf_num ;
wire [0:0] \aux_key_ctrl.dak_key_op ;
wire [13:0] \aux_key_ctrl.dak_key_ref ;
wire [1:0] \aux_key_ctrl.kdf_mode ;
wire [0:0] \aux_key_ctrl.dek_key_op ;
wire [13:0] \aux_key_ctrl.dek_key_ref ;
tran (ckvreader_kopassigner_data[70], \ckvreader_kopassigner_data.sot [0]);
tran (ckvreader_kopassigner_data[69], \ckvreader_kopassigner_data.eoi [0]);
tran (ckvreader_kopassigner_data[68], \ckvreader_kopassigner_data.eot [0]);
tran (ckvreader_kopassigner_data[67], \ckvreader_kopassigner_data.id [3]);
tran (ckvreader_kopassigner_data[66], \ckvreader_kopassigner_data.id [2]);
tran (ckvreader_kopassigner_data[65], \ckvreader_kopassigner_data.id [1]);
tran (ckvreader_kopassigner_data[64], \ckvreader_kopassigner_data.id [0]);
tran (ckvreader_kopassigner_data[63], \ckvreader_kopassigner_data.tdata [63]);
tran (ckvreader_kopassigner_data[62], \ckvreader_kopassigner_data.tdata [62]);
tran (ckvreader_kopassigner_data[61], \ckvreader_kopassigner_data.tdata [61]);
tran (ckvreader_kopassigner_data[60], \ckvreader_kopassigner_data.tdata [60]);
tran (ckvreader_kopassigner_data[59], \ckvreader_kopassigner_data.tdata [59]);
tran (ckvreader_kopassigner_data[58], \ckvreader_kopassigner_data.tdata [58]);
tran (ckvreader_kopassigner_data[57], \ckvreader_kopassigner_data.tdata [57]);
tran (ckvreader_kopassigner_data[56], \ckvreader_kopassigner_data.tdata [56]);
tran (ckvreader_kopassigner_data[55], \ckvreader_kopassigner_data.tdata [55]);
tran (ckvreader_kopassigner_data[54], \ckvreader_kopassigner_data.tdata [54]);
tran (ckvreader_kopassigner_data[53], \ckvreader_kopassigner_data.tdata [53]);
tran (ckvreader_kopassigner_data[52], \ckvreader_kopassigner_data.tdata [52]);
tran (ckvreader_kopassigner_data[51], \ckvreader_kopassigner_data.tdata [51]);
tran (ckvreader_kopassigner_data[50], \ckvreader_kopassigner_data.tdata [50]);
tran (ckvreader_kopassigner_data[49], \ckvreader_kopassigner_data.tdata [49]);
tran (ckvreader_kopassigner_data[48], \ckvreader_kopassigner_data.tdata [48]);
tran (ckvreader_kopassigner_data[47], \ckvreader_kopassigner_data.tdata [47]);
tran (ckvreader_kopassigner_data[46], \ckvreader_kopassigner_data.tdata [46]);
tran (ckvreader_kopassigner_data[45], \ckvreader_kopassigner_data.tdata [45]);
tran (ckvreader_kopassigner_data[44], \ckvreader_kopassigner_data.tdata [44]);
tran (ckvreader_kopassigner_data[43], \ckvreader_kopassigner_data.tdata [43]);
tran (ckvreader_kopassigner_data[42], \ckvreader_kopassigner_data.tdata [42]);
tran (ckvreader_kopassigner_data[41], \ckvreader_kopassigner_data.tdata [41]);
tran (ckvreader_kopassigner_data[40], \ckvreader_kopassigner_data.tdata [40]);
tran (ckvreader_kopassigner_data[39], \ckvreader_kopassigner_data.tdata [39]);
tran (ckvreader_kopassigner_data[38], \ckvreader_kopassigner_data.tdata [38]);
tran (ckvreader_kopassigner_data[37], \ckvreader_kopassigner_data.tdata [37]);
tran (ckvreader_kopassigner_data[36], \ckvreader_kopassigner_data.tdata [36]);
tran (ckvreader_kopassigner_data[35], \ckvreader_kopassigner_data.tdata [35]);
tran (ckvreader_kopassigner_data[34], \ckvreader_kopassigner_data.tdata [34]);
tran (ckvreader_kopassigner_data[33], \ckvreader_kopassigner_data.tdata [33]);
tran (ckvreader_kopassigner_data[32], \ckvreader_kopassigner_data.tdata [32]);
tran (ckvreader_kopassigner_data[31], \ckvreader_kopassigner_data.tdata [31]);
tran (ckvreader_kopassigner_data[30], \ckvreader_kopassigner_data.tdata [30]);
tran (ckvreader_kopassigner_data[29], \ckvreader_kopassigner_data.tdata [29]);
tran (ckvreader_kopassigner_data[28], \ckvreader_kopassigner_data.tdata [28]);
tran (ckvreader_kopassigner_data[27], \ckvreader_kopassigner_data.tdata [27]);
tran (ckvreader_kopassigner_data[26], \ckvreader_kopassigner_data.tdata [26]);
tran (ckvreader_kopassigner_data[25], \ckvreader_kopassigner_data.tdata [25]);
tran (ckvreader_kopassigner_data[24], \ckvreader_kopassigner_data.tdata [24]);
tran (ckvreader_kopassigner_data[23], \ckvreader_kopassigner_data.tdata [23]);
tran (ckvreader_kopassigner_data[22], \ckvreader_kopassigner_data.tdata [22]);
tran (ckvreader_kopassigner_data[21], \ckvreader_kopassigner_data.tdata [21]);
tran (ckvreader_kopassigner_data[20], \ckvreader_kopassigner_data.tdata [20]);
tran (ckvreader_kopassigner_data[19], \ckvreader_kopassigner_data.tdata [19]);
tran (ckvreader_kopassigner_data[18], \ckvreader_kopassigner_data.tdata [18]);
tran (ckvreader_kopassigner_data[17], \ckvreader_kopassigner_data.tdata [17]);
tran (ckvreader_kopassigner_data[16], \ckvreader_kopassigner_data.tdata [16]);
tran (ckvreader_kopassigner_data[15], \ckvreader_kopassigner_data.tdata [15]);
tran (ckvreader_kopassigner_data[14], \ckvreader_kopassigner_data.tdata [14]);
tran (ckvreader_kopassigner_data[13], \ckvreader_kopassigner_data.tdata [13]);
tran (ckvreader_kopassigner_data[12], \ckvreader_kopassigner_data.tdata [12]);
tran (ckvreader_kopassigner_data[11], \ckvreader_kopassigner_data.tdata [11]);
tran (ckvreader_kopassigner_data[10], \ckvreader_kopassigner_data.tdata [10]);
tran (ckvreader_kopassigner_data[9], \ckvreader_kopassigner_data.tdata [9]);
tran (ckvreader_kopassigner_data[8], \ckvreader_kopassigner_data.tdata [8]);
tran (ckvreader_kopassigner_data[7], \ckvreader_kopassigner_data.tdata [7]);
tran (ckvreader_kopassigner_data[6], \ckvreader_kopassigner_data.tdata [6]);
tran (ckvreader_kopassigner_data[5], \ckvreader_kopassigner_data.tdata [5]);
tran (ckvreader_kopassigner_data[4], \ckvreader_kopassigner_data.tdata [4]);
tran (ckvreader_kopassigner_data[3], \ckvreader_kopassigner_data.tdata [3]);
tran (ckvreader_kopassigner_data[2], \ckvreader_kopassigner_data.tdata [2]);
tran (ckvreader_kopassigner_data[1], \ckvreader_kopassigner_data.tdata [1]);
tran (ckvreader_kopassigner_data[0], \ckvreader_kopassigner_data.tdata [0]);
tran (kimreader_ckvreader_data[70], \kimreader_ckvreader_data.sot [0]);
tran (kimreader_ckvreader_data[69], \kimreader_ckvreader_data.eoi [0]);
tran (kimreader_ckvreader_data[68], \kimreader_ckvreader_data.eot [0]);
tran (kimreader_ckvreader_data[67], \kimreader_ckvreader_data.id [3]);
tran (kimreader_ckvreader_data[66], \kimreader_ckvreader_data.id [2]);
tran (kimreader_ckvreader_data[65], \kimreader_ckvreader_data.id [1]);
tran (kimreader_ckvreader_data[64], \kimreader_ckvreader_data.id [0]);
tran (kimreader_ckvreader_data[63], \kimreader_ckvreader_data.tdata [63]);
tran (kimreader_ckvreader_data[62], \kimreader_ckvreader_data.tdata [62]);
tran (kimreader_ckvreader_data[61], \kimreader_ckvreader_data.tdata [61]);
tran (kimreader_ckvreader_data[60], \kimreader_ckvreader_data.tdata [60]);
tran (kimreader_ckvreader_data[59], \kimreader_ckvreader_data.tdata [59]);
tran (kimreader_ckvreader_data[58], \kimreader_ckvreader_data.tdata [58]);
tran (kimreader_ckvreader_data[57], \kimreader_ckvreader_data.tdata [57]);
tran (kimreader_ckvreader_data[56], \kimreader_ckvreader_data.tdata [56]);
tran (kimreader_ckvreader_data[55], \kimreader_ckvreader_data.tdata [55]);
tran (kimreader_ckvreader_data[54], \kimreader_ckvreader_data.tdata [54]);
tran (kimreader_ckvreader_data[53], \kimreader_ckvreader_data.tdata [53]);
tran (kimreader_ckvreader_data[52], \kimreader_ckvreader_data.tdata [52]);
tran (kimreader_ckvreader_data[51], \kimreader_ckvreader_data.tdata [51]);
tran (kimreader_ckvreader_data[50], \kimreader_ckvreader_data.tdata [50]);
tran (kimreader_ckvreader_data[49], \kimreader_ckvreader_data.tdata [49]);
tran (kimreader_ckvreader_data[48], \kimreader_ckvreader_data.tdata [48]);
tran (kimreader_ckvreader_data[47], \kimreader_ckvreader_data.tdata [47]);
tran (kimreader_ckvreader_data[46], \kimreader_ckvreader_data.tdata [46]);
tran (kimreader_ckvreader_data[45], \kimreader_ckvreader_data.tdata [45]);
tran (kimreader_ckvreader_data[44], \kimreader_ckvreader_data.tdata [44]);
tran (kimreader_ckvreader_data[43], \kimreader_ckvreader_data.tdata [43]);
tran (kimreader_ckvreader_data[42], \kimreader_ckvreader_data.tdata [42]);
tran (kimreader_ckvreader_data[41], \kimreader_ckvreader_data.tdata [41]);
tran (kimreader_ckvreader_data[40], \kimreader_ckvreader_data.tdata [40]);
tran (kimreader_ckvreader_data[39], \kimreader_ckvreader_data.tdata [39]);
tran (kimreader_ckvreader_data[38], \kimreader_ckvreader_data.tdata [38]);
tran (kimreader_ckvreader_data[37], \kimreader_ckvreader_data.tdata [37]);
tran (kimreader_ckvreader_data[36], \kimreader_ckvreader_data.tdata [36]);
tran (kimreader_ckvreader_data[35], \kimreader_ckvreader_data.tdata [35]);
tran (kimreader_ckvreader_data[34], \kimreader_ckvreader_data.tdata [34]);
tran (kimreader_ckvreader_data[33], \kimreader_ckvreader_data.tdata [33]);
tran (kimreader_ckvreader_data[32], \kimreader_ckvreader_data.tdata [32]);
tran (kimreader_ckvreader_data[31], \kimreader_ckvreader_data.tdata [31]);
tran (kimreader_ckvreader_data[30], \kimreader_ckvreader_data.tdata [30]);
tran (kimreader_ckvreader_data[29], \kimreader_ckvreader_data.tdata [29]);
tran (kimreader_ckvreader_data[28], \kimreader_ckvreader_data.tdata [28]);
tran (kimreader_ckvreader_data[27], \kimreader_ckvreader_data.tdata [27]);
tran (kimreader_ckvreader_data[26], \kimreader_ckvreader_data.tdata [26]);
tran (kimreader_ckvreader_data[25], \kimreader_ckvreader_data.tdata [25]);
tran (kimreader_ckvreader_data[24], \kimreader_ckvreader_data.tdata [24]);
tran (kimreader_ckvreader_data[23], \kimreader_ckvreader_data.tdata [23]);
tran (kimreader_ckvreader_data[22], \kimreader_ckvreader_data.tdata [22]);
tran (kimreader_ckvreader_data[21], \kimreader_ckvreader_data.tdata [21]);
tran (kimreader_ckvreader_data[20], \kimreader_ckvreader_data.tdata [20]);
tran (kimreader_ckvreader_data[19], \kimreader_ckvreader_data.tdata [19]);
tran (kimreader_ckvreader_data[18], \kimreader_ckvreader_data.tdata [18]);
tran (kimreader_ckvreader_data[17], \kimreader_ckvreader_data.tdata [17]);
tran (kimreader_ckvreader_data[16], \kimreader_ckvreader_data.tdata [16]);
tran (kimreader_ckvreader_data[15], \kimreader_ckvreader_data.tdata [15]);
tran (kimreader_ckvreader_data[14], \kimreader_ckvreader_data.tdata [14]);
tran (kimreader_ckvreader_data[13], \kimreader_ckvreader_data.tdata [13]);
tran (kimreader_ckvreader_data[12], \kimreader_ckvreader_data.tdata [12]);
tran (kimreader_ckvreader_data[11], \kimreader_ckvreader_data.tdata [11]);
tran (kimreader_ckvreader_data[10], \kimreader_ckvreader_data.tdata [10]);
tran (kimreader_ckvreader_data[9], \kimreader_ckvreader_data.tdata [9]);
tran (kimreader_ckvreader_data[8], \kimreader_ckvreader_data.tdata [8]);
tran (kimreader_ckvreader_data[7], \kimreader_ckvreader_data.tdata [7]);
tran (kimreader_ckvreader_data[6], \kimreader_ckvreader_data.tdata [6]);
tran (kimreader_ckvreader_data[5], \kimreader_ckvreader_data.tdata [5]);
tran (kimreader_ckvreader_data[4], \kimreader_ckvreader_data.tdata [4]);
tran (kimreader_ckvreader_data[3], \kimreader_ckvreader_data.tdata [3]);
tran (kimreader_ckvreader_data[2], \kimreader_ckvreader_data.tdata [2]);
tran (kimreader_ckvreader_data[1], \kimreader_ckvreader_data.tdata [1]);
tran (kimreader_ckvreader_data[0], \kimreader_ckvreader_data.tdata [0]);
tran (tlv_word0[63], \tlv_word0.tlv_bip2 [1]);
tran (tlv_word0[62], \tlv_word0.tlv_bip2 [0]);
tran (tlv_word0[61], \tlv_word0.resv0 [12]);
tran (tlv_word0[60], \tlv_word0.resv0 [11]);
tran (tlv_word0[59], \tlv_word0.resv0 [10]);
tran (tlv_word0[58], \tlv_word0.resv0 [9]);
tran (tlv_word0[57], \tlv_word0.resv0 [8]);
tran (tlv_word0[56], \tlv_word0.resv0 [7]);
tran (tlv_word0[55], \tlv_word0.resv0 [6]);
tran (tlv_word42[55], \tlv_word42.corrupt_crc32 [0]);
tran (tlv_word0[54], \tlv_word0.resv0 [5]);
tran (tlv_word42[54], \tlv_word42.unused [46]);
tran (tlv_word0[53], \tlv_word0.resv0 [4]);
tran (tlv_word42[53], \tlv_word42.unused [45]);
tran (tlv_word0[52], \tlv_word0.resv0 [3]);
tran (tlv_word42[52], \tlv_word42.unused [44]);
tran (tlv_word0[51], \tlv_word0.resv0 [2]);
tran (tlv_word42[51], \tlv_word42.unused [43]);
tran (tlv_word0[50], \tlv_word0.resv0 [1]);
tran (tlv_word42[50], \tlv_word42.unused [42]);
tran (tlv_word0[49], \tlv_word0.resv0 [0]);
tran (tlv_word42[49], \tlv_word42.unused [41]);
tran (tlv_word0[48], \tlv_word0.kdf_dek_iter [0]);
tran (tlv_word42[48], \tlv_word42.unused [40]);
tran (tlv_word0[47], \tlv_word0.keyless_algos [0]);
tran (tlv_word42[47], \tlv_word42.unused [39]);
tran (tlv_word0[46], \tlv_word0.needs_dek [0]);
tran (tlv_word42[46], \tlv_word42.unused [38]);
tran (tlv_word0[45], \tlv_word0.needs_dak [0]);
tran (tlv_word42[45], \tlv_word42.unused [37]);
tran (tlv_word0[44], \tlv_word0.key_type [5]);
tran (tlv_word42[44], \tlv_word42.unused [36]);
tran (tlv_word0[43], \tlv_word0.key_type [4]);
tran (tlv_word42[43], \tlv_word42.unused [35]);
tran (tlv_word0[42], \tlv_word0.key_type [3]);
tran (tlv_word42[42], \tlv_word42.unused [34]);
tran (tlv_word0[41], \tlv_word0.key_type [2]);
tran (tlv_word42[41], \tlv_word42.unused [33]);
tran (tlv_word0[40], \tlv_word0.key_type [1]);
tran (tlv_word42[40], \tlv_word42.unused [32]);
tran (tlv_word0[39], \tlv_word0.key_type [0]);
tran (tlv_word42[39], \tlv_word42.unused [31]);
tran (tlv_word0[38], \tlv_word0.tlv_frame_num [10]);
tran (tlv_word42[38], \tlv_word42.unused [30]);
tran (tlv_word0[37], \tlv_word0.tlv_frame_num [9]);
tran (tlv_word42[37], \tlv_word42.unused [29]);
tran (tlv_word0[36], \tlv_word0.tlv_frame_num [8]);
tran (tlv_word42[36], \tlv_word42.unused [28]);
tran (tlv_word0[35], \tlv_word0.tlv_frame_num [7]);
tran (tlv_word42[35], \tlv_word42.unused [27]);
tran (tlv_word0[34], \tlv_word0.tlv_frame_num [6]);
tran (tlv_word42[34], \tlv_word42.unused [26]);
tran (tlv_word0[33], \tlv_word0.tlv_frame_num [5]);
tran (tlv_word42[33], \tlv_word42.unused [25]);
tran (tlv_word0[32], \tlv_word0.tlv_frame_num [4]);
tran (tlv_word42[32], \tlv_word42.unused [24]);
tran (tlv_word0[31], \tlv_word0.tlv_frame_num [3]);
tran (tlv_word42[31], \tlv_word42.unused [23]);
tran (aux_key_ctrl[31], \aux_key_ctrl.dak_key_op [0]);
tran (tlv_word0[30], \tlv_word0.tlv_frame_num [2]);
tran (tlv_word42[30], \tlv_word42.unused [22]);
tran (aux_key_ctrl[30], \aux_key_ctrl.dak_key_ref [13]);
tran (tlv_word0[29], \tlv_word0.tlv_frame_num [1]);
tran (tlv_word42[29], \tlv_word42.unused [21]);
tran (aux_key_ctrl[29], \aux_key_ctrl.dak_key_ref [12]);
tran (tlv_word0[28], \tlv_word0.tlv_frame_num [0]);
tran (tlv_word42[28], \tlv_word42.unused [20]);
tran (aux_key_ctrl[28], \aux_key_ctrl.dak_key_ref [11]);
tran (tlv_word0[27], \tlv_word0.tlv_eng_id [3]);
tran (tlv_word42[27], \tlv_word42.unused [19]);
tran (aux_key_ctrl[27], \aux_key_ctrl.dak_key_ref [10]);
tran (tlv_word0[26], \tlv_word0.tlv_eng_id [2]);
tran (tlv_word42[26], \tlv_word42.unused [18]);
tran (aux_key_ctrl[26], \aux_key_ctrl.dak_key_ref [9]);
tran (tlv_word0[25], \tlv_word0.tlv_eng_id [1]);
tran (tlv_word42[25], \tlv_word42.unused [17]);
tran (aux_key_ctrl[25], \aux_key_ctrl.dak_key_ref [8]);
tran (tlv_word0[24], \tlv_word0.tlv_eng_id [0]);
tran (tlv_word42[24], \tlv_word42.unused [16]);
tran (aux_key_ctrl[24], \aux_key_ctrl.dak_key_ref [7]);
tran (tlv_word0[23], \tlv_word0.tlv_seq_num [7]);
tran (tlv_word42[23], \tlv_word42.unused [15]);
tran (aux_key_ctrl[23], \aux_key_ctrl.dak_key_ref [6]);
tran (tlv_word0[22], \tlv_word0.tlv_seq_num [6]);
tran (tlv_word42[22], \tlv_word42.unused [14]);
tran (aux_key_ctrl[22], \aux_key_ctrl.dak_key_ref [5]);
tran (tlv_word0[21], \tlv_word0.tlv_seq_num [5]);
tran (tlv_word42[21], \tlv_word42.unused [13]);
tran (aux_key_ctrl[21], \aux_key_ctrl.dak_key_ref [4]);
tran (tlv_word0[20], \tlv_word0.tlv_seq_num [4]);
tran (tlv_word42[20], \tlv_word42.unused [12]);
tran (aux_key_ctrl[20], \aux_key_ctrl.dak_key_ref [3]);
tran (tlv_word0[19], \tlv_word0.tlv_seq_num [3]);
tran (tlv_word42[19], \tlv_word42.unused [11]);
tran (aux_key_ctrl[19], \aux_key_ctrl.dak_key_ref [2]);
tran (tlv_word0[18], \tlv_word0.tlv_seq_num [2]);
tran (tlv_word42[18], \tlv_word42.unused [10]);
tran (aux_key_ctrl[18], \aux_key_ctrl.dak_key_ref [1]);
tran (tlv_word0[17], \tlv_word0.tlv_seq_num [1]);
tran (tlv_word42[17], \tlv_word42.unused [9]);
tran (aux_key_ctrl[17], \aux_key_ctrl.dak_key_ref [0]);
tran (tlv_word0[16], \tlv_word0.tlv_seq_num [0]);
tran (tlv_word42[16], \tlv_word42.unused [8]);
tran (aux_key_ctrl[16], \aux_key_ctrl.kdf_mode [1]);
tran (tlv_word0[15], \tlv_word0.tlv_len [7]);
tran (tlv_word42[15], \tlv_word42.unused [7]);
tran (aux_key_ctrl[15], \aux_key_ctrl.kdf_mode [0]);
tran (tlv_word0[14], \tlv_word0.tlv_len [6]);
tran (tlv_word42[14], \tlv_word42.unused [6]);
tran (aux_key_ctrl[14], \aux_key_ctrl.dek_key_op [0]);
tran (tlv_word0[13], \tlv_word0.tlv_len [5]);
tran (tlv_word42[13], \tlv_word42.unused [5]);
tran (aux_key_ctrl[13], \aux_key_ctrl.dek_key_ref [13]);
tran (tlv_word0[12], \tlv_word0.tlv_len [4]);
tran (tlv_word42[12], \tlv_word42.unused [4]);
tran (aux_key_ctrl[12], \aux_key_ctrl.dek_key_ref [12]);
tran (tlv_word0[11], \tlv_word0.tlv_len [3]);
tran (tlv_word42[11], \tlv_word42.unused [3]);
tran (aux_key_ctrl[11], \aux_key_ctrl.dek_key_ref [11]);
tran (tlv_word0[10], \tlv_word0.tlv_len [2]);
tran (tlv_word42[10], \tlv_word42.unused [2]);
tran (aux_key_ctrl[10], \aux_key_ctrl.dek_key_ref [10]);
tran (tlv_word0[9], \tlv_word0.tlv_len [1]);
tran (tlv_word42[9], \tlv_word42.unused [1]);
tran (aux_key_ctrl[9], \aux_key_ctrl.dek_key_ref [9]);
tran (tlv_word0[8], \tlv_word0.tlv_len [0]);
tran (tlv_word42[8], \tlv_word42.unused [0]);
tran (aux_key_ctrl[8], \aux_key_ctrl.dek_key_ref [8]);
tran (tlv_word0[7], \tlv_word0.tlv_type [7]);
tran (aux_key_ctrl[7], \aux_key_ctrl.dek_key_ref [7]);
tran (tlv_word0[6], \tlv_word0.tlv_type [6]);
tran (aux_key_ctrl[6], \aux_key_ctrl.dek_key_ref [6]);
tran (tlv_word0[5], \tlv_word0.tlv_type [5]);
tran (aux_key_ctrl[5], \aux_key_ctrl.dek_key_ref [5]);
tran (tlv_word0[4], \tlv_word0.tlv_type [4]);
tran (aux_key_ctrl[4], \aux_key_ctrl.dek_key_ref [4]);
tran (tlv_word0[3], \tlv_word0.tlv_type [3]);
tran (aux_key_ctrl[3], \aux_key_ctrl.dek_key_ref [3]);
tran (tlv_word0[2], \tlv_word0.tlv_type [2]);
tran (aux_key_ctrl[2], \aux_key_ctrl.dek_key_ref [2]);
tran (tlv_word0[1], \tlv_word0.tlv_type [1]);
tran (aux_key_ctrl[1], \aux_key_ctrl.dek_key_ref [1]);
tran (tlv_word0[0], \tlv_word0.tlv_type [0]);
tran (aux_key_ctrl[0], \aux_key_ctrl.dek_key_ref [0]);
tran (tlv_word9[17], \tlv_word9.validate_dak [0]);
tran (tlv_word8[17], \tlv_word8.validate_dek [0]);
tran (nxt_tlv_word9[0], \nxt_tlv_word9.vf_num [0]);
tran (nxt_tlv_word9[1], \nxt_tlv_word9.vf_num [1]);
tran (nxt_tlv_word9[2], \nxt_tlv_word9.vf_num [2]);
tran (nxt_tlv_word9[3], \nxt_tlv_word9.vf_num [3]);
tran (nxt_tlv_word9[4], \nxt_tlv_word9.vf_num [4]);
tran (nxt_tlv_word9[5], \nxt_tlv_word9.vf_num [5]);
tran (nxt_tlv_word9[6], \nxt_tlv_word9.vf_num [6]);
tran (nxt_tlv_word9[7], \nxt_tlv_word9.vf_num [7]);
tran (nxt_tlv_word9[8], \nxt_tlv_word9.vf_num [8]);
tran (nxt_tlv_word9[9], \nxt_tlv_word9.vf_num [9]);
tran (nxt_tlv_word9[10], \nxt_tlv_word9.vf_num [10]);
tran (nxt_tlv_word9[11], \nxt_tlv_word9.vf_num [11]);
tran (nxt_tlv_word9[12], \nxt_tlv_word9.pf_num [0]);
tran (nxt_tlv_word9[13], \nxt_tlv_word9.pf_num [1]);
tran (nxt_tlv_word9[14], \nxt_tlv_word9.pf_num [2]);
tran (nxt_tlv_word9[15], \nxt_tlv_word9.pf_num [3]);
tran (nxt_tlv_word9[16], \nxt_tlv_word9.vf_valid [0]);
tran (nxt_tlv_word9[17], \nxt_tlv_word9.validate_dak [0]);
tran (nxt_tlv_word9[18], \nxt_tlv_word9.unused [0]);
tran (nxt_tlv_word9[19], \nxt_tlv_word9.unused [1]);
tran (nxt_tlv_word9[20], \nxt_tlv_word9.unused [2]);
tran (nxt_tlv_word9[21], \nxt_tlv_word9.unused [3]);
tran (nxt_tlv_word9[22], \nxt_tlv_word9.unused [4]);
tran (nxt_tlv_word9[23], \nxt_tlv_word9.unused [5]);
tran (nxt_tlv_word9[24], \nxt_tlv_word9.unused [6]);
tran (nxt_tlv_word9[25], \nxt_tlv_word9.unused [7]);
tran (nxt_tlv_word9[26], \nxt_tlv_word9.dak_kim_entry.vf_valid [0]);
tran (nxt_tlv_word9[27], \nxt_tlv_word9.dak_kim_entry.vf_num [0]);
tran (nxt_tlv_word9[28], \nxt_tlv_word9.dak_kim_entry.vf_num [1]);
tran (nxt_tlv_word9[29], \nxt_tlv_word9.dak_kim_entry.vf_num [2]);
tran (nxt_tlv_word9[30], \nxt_tlv_word9.dak_kim_entry.vf_num [3]);
tran (nxt_tlv_word9[31], \nxt_tlv_word9.dak_kim_entry.vf_num [4]);
tran (nxt_tlv_word9[32], \nxt_tlv_word9.dak_kim_entry.vf_num [5]);
tran (nxt_tlv_word9[33], \nxt_tlv_word9.dak_kim_entry.vf_num [6]);
tran (nxt_tlv_word9[34], \nxt_tlv_word9.dak_kim_entry.vf_num [7]);
tran (nxt_tlv_word9[35], \nxt_tlv_word9.dak_kim_entry.vf_num [8]);
tran (nxt_tlv_word9[36], \nxt_tlv_word9.dak_kim_entry.vf_num [9]);
tran (nxt_tlv_word9[37], \nxt_tlv_word9.dak_kim_entry.vf_num [10]);
tran (nxt_tlv_word9[38], \nxt_tlv_word9.dak_kim_entry.vf_num [11]);
tran (nxt_tlv_word9[39], \nxt_tlv_word9.dak_kim_entry.pf_num [0]);
tran (nxt_tlv_word9[40], \nxt_tlv_word9.dak_kim_entry.pf_num [1]);
tran (nxt_tlv_word9[41], \nxt_tlv_word9.dak_kim_entry.pf_num [2]);
tran (nxt_tlv_word9[42], \nxt_tlv_word9.dak_kim_entry.pf_num [3]);
tran (nxt_tlv_word9[43], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [0]);
tran (nxt_tlv_word9[44], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [1]);
tran (nxt_tlv_word9[45], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [2]);
tran (nxt_tlv_word9[46], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [3]);
tran (nxt_tlv_word9[47], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [4]);
tran (nxt_tlv_word9[48], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [5]);
tran (nxt_tlv_word9[49], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [6]);
tran (nxt_tlv_word9[50], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [7]);
tran (nxt_tlv_word9[51], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [8]);
tran (nxt_tlv_word9[52], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [9]);
tran (nxt_tlv_word9[53], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [10]);
tran (nxt_tlv_word9[54], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [11]);
tran (nxt_tlv_word9[55], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [12]);
tran (nxt_tlv_word9[56], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [13]);
tran (nxt_tlv_word9[57], \nxt_tlv_word9.dak_kim_entry.ckv_pointer [14]);
tran (nxt_tlv_word9[58], \nxt_tlv_word9.dak_kim_entry.ckv_length [0]);
tran (nxt_tlv_word9[59], \nxt_tlv_word9.dak_kim_entry.ckv_length [1]);
tran (nxt_tlv_word9[60], \nxt_tlv_word9.dak_kim_entry.label_index [0]);
tran (nxt_tlv_word9[61], \nxt_tlv_word9.dak_kim_entry.label_index [1]);
tran (nxt_tlv_word9[62], \nxt_tlv_word9.dak_kim_entry.label_index [2]);
tran (nxt_tlv_word9[63], \nxt_tlv_word9.dak_kim_entry.valid [0]);
tran (nxt_tlv_word8[0], \nxt_tlv_word8.vf_num [0]);
tran (nxt_tlv_word8[1], \nxt_tlv_word8.vf_num [1]);
tran (nxt_tlv_word8[2], \nxt_tlv_word8.vf_num [2]);
tran (nxt_tlv_word8[3], \nxt_tlv_word8.vf_num [3]);
tran (nxt_tlv_word8[4], \nxt_tlv_word8.vf_num [4]);
tran (nxt_tlv_word8[5], \nxt_tlv_word8.vf_num [5]);
tran (nxt_tlv_word8[6], \nxt_tlv_word8.vf_num [6]);
tran (nxt_tlv_word8[7], \nxt_tlv_word8.vf_num [7]);
tran (nxt_tlv_word8[8], \nxt_tlv_word8.vf_num [8]);
tran (nxt_tlv_word8[9], \nxt_tlv_word8.vf_num [9]);
tran (nxt_tlv_word8[10], \nxt_tlv_word8.vf_num [10]);
tran (nxt_tlv_word8[11], \nxt_tlv_word8.vf_num [11]);
tran (nxt_tlv_word8[12], \nxt_tlv_word8.pf_num [0]);
tran (nxt_tlv_word8[13], \nxt_tlv_word8.pf_num [1]);
tran (nxt_tlv_word8[14], \nxt_tlv_word8.pf_num [2]);
tran (nxt_tlv_word8[15], \nxt_tlv_word8.pf_num [3]);
tran (nxt_tlv_word8[16], \nxt_tlv_word8.vf_valid [0]);
tran (nxt_tlv_word8[17], \nxt_tlv_word8.validate_dek [0]);
tran (nxt_tlv_word8[18], \nxt_tlv_word8.missing_guid [0]);
tran (nxt_tlv_word8[19], \nxt_tlv_word8.missing_iv [0]);
tran (nxt_tlv_word8[20], \nxt_tlv_word8.unused [0]);
tran (nxt_tlv_word8[21], \nxt_tlv_word8.unused [1]);
tran (nxt_tlv_word8[22], \nxt_tlv_word8.unused [2]);
tran (nxt_tlv_word8[23], \nxt_tlv_word8.unused [3]);
tran (nxt_tlv_word8[24], \nxt_tlv_word8.unused [4]);
tran (nxt_tlv_word8[25], \nxt_tlv_word8.unused [5]);
tran (nxt_tlv_word8[26], \nxt_tlv_word8.dek_kim_entry.vf_valid [0]);
tran (nxt_tlv_word8[27], \nxt_tlv_word8.dek_kim_entry.vf_num [0]);
tran (nxt_tlv_word8[28], \nxt_tlv_word8.dek_kim_entry.vf_num [1]);
tran (nxt_tlv_word8[29], \nxt_tlv_word8.dek_kim_entry.vf_num [2]);
tran (nxt_tlv_word8[30], \nxt_tlv_word8.dek_kim_entry.vf_num [3]);
tran (nxt_tlv_word8[31], \nxt_tlv_word8.dek_kim_entry.vf_num [4]);
tran (nxt_tlv_word8[32], \nxt_tlv_word8.dek_kim_entry.vf_num [5]);
tran (nxt_tlv_word8[33], \nxt_tlv_word8.dek_kim_entry.vf_num [6]);
tran (nxt_tlv_word8[34], \nxt_tlv_word8.dek_kim_entry.vf_num [7]);
tran (nxt_tlv_word8[35], \nxt_tlv_word8.dek_kim_entry.vf_num [8]);
tran (nxt_tlv_word8[36], \nxt_tlv_word8.dek_kim_entry.vf_num [9]);
tran (nxt_tlv_word8[37], \nxt_tlv_word8.dek_kim_entry.vf_num [10]);
tran (nxt_tlv_word8[38], \nxt_tlv_word8.dek_kim_entry.vf_num [11]);
tran (nxt_tlv_word8[39], \nxt_tlv_word8.dek_kim_entry.pf_num [0]);
tran (nxt_tlv_word8[40], \nxt_tlv_word8.dek_kim_entry.pf_num [1]);
tran (nxt_tlv_word8[41], \nxt_tlv_word8.dek_kim_entry.pf_num [2]);
tran (nxt_tlv_word8[42], \nxt_tlv_word8.dek_kim_entry.pf_num [3]);
tran (nxt_tlv_word8[43], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [0]);
tran (nxt_tlv_word8[44], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [1]);
tran (nxt_tlv_word8[45], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [2]);
tran (nxt_tlv_word8[46], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [3]);
tran (nxt_tlv_word8[47], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [4]);
tran (nxt_tlv_word8[48], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [5]);
tran (nxt_tlv_word8[49], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [6]);
tran (nxt_tlv_word8[50], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [7]);
tran (nxt_tlv_word8[51], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [8]);
tran (nxt_tlv_word8[52], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [9]);
tran (nxt_tlv_word8[53], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [10]);
tran (nxt_tlv_word8[54], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [11]);
tran (nxt_tlv_word8[55], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [12]);
tran (nxt_tlv_word8[56], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [13]);
tran (nxt_tlv_word8[57], \nxt_tlv_word8.dek_kim_entry.ckv_pointer [14]);
tran (nxt_tlv_word8[58], \nxt_tlv_word8.dek_kim_entry.ckv_length [0]);
tran (nxt_tlv_word8[59], \nxt_tlv_word8.dek_kim_entry.ckv_length [1]);
tran (nxt_tlv_word8[60], \nxt_tlv_word8.dek_kim_entry.label_index [0]);
tran (nxt_tlv_word8[61], \nxt_tlv_word8.dek_kim_entry.label_index [1]);
tran (nxt_tlv_word8[62], \nxt_tlv_word8.dek_kim_entry.label_index [2]);
tran (nxt_tlv_word8[63], \nxt_tlv_word8.dek_kim_entry.valid [0]);
tran (tlv_word42[0], \tlv_word42.error_code [0]);
tran (tlv_word42[1], \tlv_word42.error_code [1]);
tran (tlv_word42[2], \tlv_word42.error_code [2]);
tran (tlv_word42[3], \tlv_word42.error_code [3]);
tran (tlv_word42[4], \tlv_word42.error_code [4]);
tran (tlv_word42[5], \tlv_word42.error_code [5]);
tran (tlv_word42[6], \tlv_word42.error_code [6]);
tran (tlv_word42[7], \tlv_word42.error_code [7]);
tran (tlv_word9[0], \tlv_word9.vf_num [0]);
tran (tlv_word9[1], \tlv_word9.vf_num [1]);
tran (tlv_word9[2], \tlv_word9.vf_num [2]);
tran (tlv_word9[3], \tlv_word9.vf_num [3]);
tran (tlv_word9[4], \tlv_word9.vf_num [4]);
tran (tlv_word9[5], \tlv_word9.vf_num [5]);
tran (tlv_word9[6], \tlv_word9.vf_num [6]);
tran (tlv_word9[7], \tlv_word9.vf_num [7]);
tran (tlv_word9[8], \tlv_word9.vf_num [8]);
tran (tlv_word9[9], \tlv_word9.vf_num [9]);
tran (tlv_word9[10], \tlv_word9.vf_num [10]);
tran (tlv_word9[11], \tlv_word9.vf_num [11]);
tran (tlv_word9[12], \tlv_word9.pf_num [0]);
tran (tlv_word9[13], \tlv_word9.pf_num [1]);
tran (tlv_word9[14], \tlv_word9.pf_num [2]);
tran (tlv_word9[15], \tlv_word9.pf_num [3]);
tran (tlv_word9[16], \tlv_word9.vf_valid [0]);
tran (tlv_word9[18], \tlv_word9.unused [0]);
tran (tlv_word9[19], \tlv_word9.unused [1]);
tran (tlv_word9[20], \tlv_word9.unused [2]);
tran (tlv_word9[21], \tlv_word9.unused [3]);
tran (tlv_word9[22], \tlv_word9.unused [4]);
tran (tlv_word9[23], \tlv_word9.unused [5]);
tran (tlv_word9[24], \tlv_word9.unused [6]);
tran (tlv_word9[25], \tlv_word9.unused [7]);
tran (tlv_word9[26], \tlv_word9.dak_kim_entry.vf_valid [0]);
tran (tlv_word9[27], \tlv_word9.dak_kim_entry.vf_num [0]);
tran (tlv_word9[28], \tlv_word9.dak_kim_entry.vf_num [1]);
tran (tlv_word9[29], \tlv_word9.dak_kim_entry.vf_num [2]);
tran (tlv_word9[30], \tlv_word9.dak_kim_entry.vf_num [3]);
tran (tlv_word9[31], \tlv_word9.dak_kim_entry.vf_num [4]);
tran (tlv_word9[32], \tlv_word9.dak_kim_entry.vf_num [5]);
tran (tlv_word9[33], \tlv_word9.dak_kim_entry.vf_num [6]);
tran (tlv_word9[34], \tlv_word9.dak_kim_entry.vf_num [7]);
tran (tlv_word9[35], \tlv_word9.dak_kim_entry.vf_num [8]);
tran (tlv_word9[36], \tlv_word9.dak_kim_entry.vf_num [9]);
tran (tlv_word9[37], \tlv_word9.dak_kim_entry.vf_num [10]);
tran (tlv_word9[38], \tlv_word9.dak_kim_entry.vf_num [11]);
tran (tlv_word9[39], \tlv_word9.dak_kim_entry.pf_num [0]);
tran (tlv_word9[40], \tlv_word9.dak_kim_entry.pf_num [1]);
tran (tlv_word9[41], \tlv_word9.dak_kim_entry.pf_num [2]);
tran (tlv_word9[42], \tlv_word9.dak_kim_entry.pf_num [3]);
tran (tlv_word9[43], \tlv_word9.dak_kim_entry.ckv_pointer [0]);
tran (tlv_word9[44], \tlv_word9.dak_kim_entry.ckv_pointer [1]);
tran (tlv_word9[45], \tlv_word9.dak_kim_entry.ckv_pointer [2]);
tran (tlv_word9[46], \tlv_word9.dak_kim_entry.ckv_pointer [3]);
tran (tlv_word9[47], \tlv_word9.dak_kim_entry.ckv_pointer [4]);
tran (tlv_word9[48], \tlv_word9.dak_kim_entry.ckv_pointer [5]);
tran (tlv_word9[49], \tlv_word9.dak_kim_entry.ckv_pointer [6]);
tran (tlv_word9[50], \tlv_word9.dak_kim_entry.ckv_pointer [7]);
tran (tlv_word9[51], \tlv_word9.dak_kim_entry.ckv_pointer [8]);
tran (tlv_word9[52], \tlv_word9.dak_kim_entry.ckv_pointer [9]);
tran (tlv_word9[53], \tlv_word9.dak_kim_entry.ckv_pointer [10]);
tran (tlv_word9[54], \tlv_word9.dak_kim_entry.ckv_pointer [11]);
tran (tlv_word9[55], \tlv_word9.dak_kim_entry.ckv_pointer [12]);
tran (tlv_word9[56], \tlv_word9.dak_kim_entry.ckv_pointer [13]);
tran (tlv_word9[57], \tlv_word9.dak_kim_entry.ckv_pointer [14]);
tran (tlv_word9[58], \tlv_word9.dak_kim_entry.ckv_length [0]);
tran (tlv_word9[59], \tlv_word9.dak_kim_entry.ckv_length [1]);
tran (tlv_word9[60], \tlv_word9.dak_kim_entry.label_index [0]);
tran (tlv_word9[61], \tlv_word9.dak_kim_entry.label_index [1]);
tran (tlv_word9[62], \tlv_word9.dak_kim_entry.label_index [2]);
tran (tlv_word9[63], \tlv_word9.dak_kim_entry.valid [0]);
tran (tlv_word8[0], \tlv_word8.vf_num [0]);
tran (tlv_word8[1], \tlv_word8.vf_num [1]);
tran (tlv_word8[2], \tlv_word8.vf_num [2]);
tran (tlv_word8[3], \tlv_word8.vf_num [3]);
tran (tlv_word8[4], \tlv_word8.vf_num [4]);
tran (tlv_word8[5], \tlv_word8.vf_num [5]);
tran (tlv_word8[6], \tlv_word8.vf_num [6]);
tran (tlv_word8[7], \tlv_word8.vf_num [7]);
tran (tlv_word8[8], \tlv_word8.vf_num [8]);
tran (tlv_word8[9], \tlv_word8.vf_num [9]);
tran (tlv_word8[10], \tlv_word8.vf_num [10]);
tran (tlv_word8[11], \tlv_word8.vf_num [11]);
tran (tlv_word8[12], \tlv_word8.pf_num [0]);
tran (tlv_word8[13], \tlv_word8.pf_num [1]);
tran (tlv_word8[14], \tlv_word8.pf_num [2]);
tran (tlv_word8[15], \tlv_word8.pf_num [3]);
tran (tlv_word8[16], \tlv_word8.vf_valid [0]);
tran (tlv_word8[18], \tlv_word8.missing_guid [0]);
tran (tlv_word8[19], \tlv_word8.missing_iv [0]);
tran (tlv_word8[20], \tlv_word8.unused [0]);
tran (tlv_word8[21], \tlv_word8.unused [1]);
tran (tlv_word8[22], \tlv_word8.unused [2]);
tran (tlv_word8[23], \tlv_word8.unused [3]);
tran (tlv_word8[24], \tlv_word8.unused [4]);
tran (tlv_word8[25], \tlv_word8.unused [5]);
tran (tlv_word8[26], \tlv_word8.dek_kim_entry.vf_valid [0]);
tran (tlv_word8[27], \tlv_word8.dek_kim_entry.vf_num [0]);
tran (tlv_word8[28], \tlv_word8.dek_kim_entry.vf_num [1]);
tran (tlv_word8[29], \tlv_word8.dek_kim_entry.vf_num [2]);
tran (tlv_word8[30], \tlv_word8.dek_kim_entry.vf_num [3]);
tran (tlv_word8[31], \tlv_word8.dek_kim_entry.vf_num [4]);
tran (tlv_word8[32], \tlv_word8.dek_kim_entry.vf_num [5]);
tran (tlv_word8[33], \tlv_word8.dek_kim_entry.vf_num [6]);
tran (tlv_word8[34], \tlv_word8.dek_kim_entry.vf_num [7]);
tran (tlv_word8[35], \tlv_word8.dek_kim_entry.vf_num [8]);
tran (tlv_word8[36], \tlv_word8.dek_kim_entry.vf_num [9]);
tran (tlv_word8[37], \tlv_word8.dek_kim_entry.vf_num [10]);
tran (tlv_word8[38], \tlv_word8.dek_kim_entry.vf_num [11]);
tran (tlv_word8[39], \tlv_word8.dek_kim_entry.pf_num [0]);
tran (tlv_word8[40], \tlv_word8.dek_kim_entry.pf_num [1]);
tran (tlv_word8[41], \tlv_word8.dek_kim_entry.pf_num [2]);
tran (tlv_word8[42], \tlv_word8.dek_kim_entry.pf_num [3]);
tran (tlv_word8[43], \tlv_word8.dek_kim_entry.ckv_pointer [0]);
tran (tlv_word8[44], \tlv_word8.dek_kim_entry.ckv_pointer [1]);
tran (tlv_word8[45], \tlv_word8.dek_kim_entry.ckv_pointer [2]);
tran (tlv_word8[46], \tlv_word8.dek_kim_entry.ckv_pointer [3]);
tran (tlv_word8[47], \tlv_word8.dek_kim_entry.ckv_pointer [4]);
tran (tlv_word8[48], \tlv_word8.dek_kim_entry.ckv_pointer [5]);
tran (tlv_word8[49], \tlv_word8.dek_kim_entry.ckv_pointer [6]);
tran (tlv_word8[50], \tlv_word8.dek_kim_entry.ckv_pointer [7]);
tran (tlv_word8[51], \tlv_word8.dek_kim_entry.ckv_pointer [8]);
tran (tlv_word8[52], \tlv_word8.dek_kim_entry.ckv_pointer [9]);
tran (tlv_word8[53], \tlv_word8.dek_kim_entry.ckv_pointer [10]);
tran (tlv_word8[54], \tlv_word8.dek_kim_entry.ckv_pointer [11]);
tran (tlv_word8[55], \tlv_word8.dek_kim_entry.ckv_pointer [12]);
tran (tlv_word8[56], \tlv_word8.dek_kim_entry.ckv_pointer [13]);
tran (tlv_word8[57], \tlv_word8.dek_kim_entry.ckv_pointer [14]);
tran (tlv_word8[58], \tlv_word8.dek_kim_entry.ckv_length [0]);
tran (tlv_word8[59], \tlv_word8.dek_kim_entry.ckv_length [1]);
tran (tlv_word8[60], \tlv_word8.dek_kim_entry.label_index [0]);
tran (tlv_word8[61], \tlv_word8.dek_kim_entry.label_index [1]);
tran (tlv_word8[62], \tlv_word8.dek_kim_entry.label_index [2]);
tran (tlv_word8[63], \tlv_word8.dek_kim_entry.valid [0]);
Q_BUF U0 ( .A(n2), .Z(_zy_simnet_cio_9));
Q_ASSIGN U1 ( .B(kimreader_ckvreader_data[63]), .A(tlv_word0[63]));
Q_ASSIGN U2 ( .B(kimreader_ckvreader_data[62]), .A(tlv_word0[62]));
Q_ASSIGN U3 ( .B(kimreader_ckvreader_data[61]), .A(tlv_word0[61]));
Q_ASSIGN U4 ( .B(kimreader_ckvreader_data[60]), .A(tlv_word0[60]));
Q_ASSIGN U5 ( .B(kimreader_ckvreader_data[59]), .A(tlv_word0[59]));
Q_ASSIGN U6 ( .B(kimreader_ckvreader_data[58]), .A(tlv_word0[58]));
Q_ASSIGN U7 ( .B(kimreader_ckvreader_data[57]), .A(tlv_word0[57]));
Q_ASSIGN U8 ( .B(kimreader_ckvreader_data[56]), .A(tlv_word0[56]));
Q_ASSIGN U9 ( .B(kimreader_ckvreader_data[55]), .A(tlv_word0[55]));
Q_ASSIGN U10 ( .B(kimreader_ckvreader_data[55]), .A(tlv_word42[55]));
Q_ASSIGN U11 ( .B(kimreader_ckvreader_data[54]), .A(tlv_word0[54]));
Q_ASSIGN U12 ( .B(kimreader_ckvreader_data[54]), .A(tlv_word42[54]));
Q_ASSIGN U13 ( .B(kimreader_ckvreader_data[53]), .A(tlv_word0[53]));
Q_ASSIGN U14 ( .B(kimreader_ckvreader_data[53]), .A(tlv_word42[53]));
Q_ASSIGN U15 ( .B(kimreader_ckvreader_data[52]), .A(tlv_word0[52]));
Q_ASSIGN U16 ( .B(kimreader_ckvreader_data[52]), .A(tlv_word42[52]));
Q_ASSIGN U17 ( .B(kimreader_ckvreader_data[51]), .A(tlv_word0[51]));
Q_ASSIGN U18 ( .B(kimreader_ckvreader_data[51]), .A(tlv_word42[51]));
Q_ASSIGN U19 ( .B(kimreader_ckvreader_data[50]), .A(tlv_word0[50]));
Q_ASSIGN U20 ( .B(kimreader_ckvreader_data[50]), .A(tlv_word42[50]));
Q_ASSIGN U21 ( .B(kimreader_ckvreader_data[49]), .A(tlv_word0[49]));
Q_ASSIGN U22 ( .B(kimreader_ckvreader_data[49]), .A(tlv_word42[49]));
Q_ASSIGN U23 ( .B(kimreader_ckvreader_data[48]), .A(tlv_word0[48]));
Q_ASSIGN U24 ( .B(kimreader_ckvreader_data[48]), .A(tlv_word42[48]));
Q_ASSIGN U25 ( .B(kimreader_ckvreader_data[47]), .A(tlv_word0[47]));
Q_ASSIGN U26 ( .B(kimreader_ckvreader_data[47]), .A(tlv_word42[47]));
Q_ASSIGN U27 ( .B(kimreader_ckvreader_data[46]), .A(tlv_word0[46]));
Q_ASSIGN U28 ( .B(kimreader_ckvreader_data[46]), .A(tlv_word42[46]));
Q_ASSIGN U29 ( .B(kimreader_ckvreader_data[45]), .A(tlv_word0[45]));
Q_ASSIGN U30 ( .B(kimreader_ckvreader_data[45]), .A(tlv_word42[45]));
Q_ASSIGN U31 ( .B(kimreader_ckvreader_data[44]), .A(tlv_word0[44]));
Q_ASSIGN U32 ( .B(kimreader_ckvreader_data[44]), .A(tlv_word42[44]));
Q_ASSIGN U33 ( .B(kimreader_ckvreader_data[43]), .A(tlv_word0[43]));
Q_ASSIGN U34 ( .B(kimreader_ckvreader_data[43]), .A(tlv_word42[43]));
Q_ASSIGN U35 ( .B(kimreader_ckvreader_data[42]), .A(tlv_word0[42]));
Q_ASSIGN U36 ( .B(kimreader_ckvreader_data[42]), .A(tlv_word42[42]));
Q_ASSIGN U37 ( .B(kimreader_ckvreader_data[41]), .A(tlv_word0[41]));
Q_ASSIGN U38 ( .B(kimreader_ckvreader_data[41]), .A(tlv_word42[41]));
Q_ASSIGN U39 ( .B(kimreader_ckvreader_data[40]), .A(tlv_word0[40]));
Q_ASSIGN U40 ( .B(kimreader_ckvreader_data[40]), .A(tlv_word42[40]));
Q_ASSIGN U41 ( .B(kimreader_ckvreader_data[39]), .A(tlv_word0[39]));
Q_ASSIGN U42 ( .B(kimreader_ckvreader_data[39]), .A(tlv_word42[39]));
Q_ASSIGN U43 ( .B(kimreader_ckvreader_data[38]), .A(tlv_word0[38]));
Q_ASSIGN U44 ( .B(kimreader_ckvreader_data[38]), .A(tlv_word42[38]));
Q_ASSIGN U45 ( .B(kimreader_ckvreader_data[37]), .A(tlv_word0[37]));
Q_ASSIGN U46 ( .B(kimreader_ckvreader_data[37]), .A(tlv_word42[37]));
Q_ASSIGN U47 ( .B(kimreader_ckvreader_data[36]), .A(tlv_word0[36]));
Q_ASSIGN U48 ( .B(kimreader_ckvreader_data[36]), .A(tlv_word42[36]));
Q_ASSIGN U49 ( .B(kimreader_ckvreader_data[35]), .A(tlv_word0[35]));
Q_ASSIGN U50 ( .B(kimreader_ckvreader_data[35]), .A(tlv_word42[35]));
Q_ASSIGN U51 ( .B(kimreader_ckvreader_data[34]), .A(tlv_word0[34]));
Q_ASSIGN U52 ( .B(kimreader_ckvreader_data[34]), .A(tlv_word42[34]));
Q_ASSIGN U53 ( .B(kimreader_ckvreader_data[33]), .A(tlv_word0[33]));
Q_ASSIGN U54 ( .B(kimreader_ckvreader_data[33]), .A(tlv_word42[33]));
Q_ASSIGN U55 ( .B(kimreader_ckvreader_data[32]), .A(tlv_word0[32]));
Q_ASSIGN U56 ( .B(kimreader_ckvreader_data[32]), .A(tlv_word42[32]));
Q_ASSIGN U57 ( .B(kimreader_ckvreader_data[31]), .A(tlv_word0[31]));
Q_ASSIGN U58 ( .B(kimreader_ckvreader_data[31]), .A(tlv_word42[31]));
Q_ASSIGN U59 ( .B(kimreader_ckvreader_data[31]), .A(aux_key_ctrl[31]));
Q_ASSIGN U60 ( .B(kimreader_ckvreader_data[30]), .A(tlv_word0[30]));
Q_ASSIGN U61 ( .B(kimreader_ckvreader_data[30]), .A(tlv_word42[30]));
Q_ASSIGN U62 ( .B(kimreader_ckvreader_data[30]), .A(aux_key_ctrl[30]));
Q_ASSIGN U63 ( .B(kimreader_ckvreader_data[29]), .A(tlv_word0[29]));
Q_ASSIGN U64 ( .B(kimreader_ckvreader_data[29]), .A(tlv_word42[29]));
Q_ASSIGN U65 ( .B(kimreader_ckvreader_data[29]), .A(aux_key_ctrl[29]));
Q_ASSIGN U66 ( .B(kimreader_ckvreader_data[28]), .A(tlv_word0[28]));
Q_ASSIGN U67 ( .B(kimreader_ckvreader_data[28]), .A(tlv_word42[28]));
Q_ASSIGN U68 ( .B(kimreader_ckvreader_data[28]), .A(aux_key_ctrl[28]));
Q_ASSIGN U69 ( .B(kimreader_ckvreader_data[27]), .A(tlv_word0[27]));
Q_ASSIGN U70 ( .B(kimreader_ckvreader_data[27]), .A(tlv_word42[27]));
Q_ASSIGN U71 ( .B(kimreader_ckvreader_data[27]), .A(aux_key_ctrl[27]));
Q_ASSIGN U72 ( .B(kimreader_ckvreader_data[26]), .A(tlv_word0[26]));
Q_ASSIGN U73 ( .B(kimreader_ckvreader_data[26]), .A(tlv_word42[26]));
Q_ASSIGN U74 ( .B(kimreader_ckvreader_data[26]), .A(aux_key_ctrl[26]));
Q_ASSIGN U75 ( .B(kimreader_ckvreader_data[25]), .A(tlv_word0[25]));
Q_ASSIGN U76 ( .B(kimreader_ckvreader_data[25]), .A(tlv_word42[25]));
Q_ASSIGN U77 ( .B(kimreader_ckvreader_data[25]), .A(aux_key_ctrl[25]));
Q_ASSIGN U78 ( .B(kimreader_ckvreader_data[24]), .A(tlv_word0[24]));
Q_ASSIGN U79 ( .B(kimreader_ckvreader_data[24]), .A(tlv_word42[24]));
Q_ASSIGN U80 ( .B(kimreader_ckvreader_data[24]), .A(aux_key_ctrl[24]));
Q_ASSIGN U81 ( .B(kimreader_ckvreader_data[23]), .A(tlv_word0[23]));
Q_ASSIGN U82 ( .B(kimreader_ckvreader_data[23]), .A(tlv_word42[23]));
Q_ASSIGN U83 ( .B(kimreader_ckvreader_data[23]), .A(aux_key_ctrl[23]));
Q_ASSIGN U84 ( .B(kimreader_ckvreader_data[22]), .A(tlv_word0[22]));
Q_ASSIGN U85 ( .B(kimreader_ckvreader_data[22]), .A(tlv_word42[22]));
Q_ASSIGN U86 ( .B(kimreader_ckvreader_data[22]), .A(aux_key_ctrl[22]));
Q_ASSIGN U87 ( .B(kimreader_ckvreader_data[21]), .A(tlv_word0[21]));
Q_ASSIGN U88 ( .B(kimreader_ckvreader_data[21]), .A(tlv_word42[21]));
Q_ASSIGN U89 ( .B(kimreader_ckvreader_data[21]), .A(aux_key_ctrl[21]));
Q_ASSIGN U90 ( .B(kimreader_ckvreader_data[20]), .A(tlv_word0[20]));
Q_ASSIGN U91 ( .B(kimreader_ckvreader_data[20]), .A(tlv_word42[20]));
Q_ASSIGN U92 ( .B(kimreader_ckvreader_data[20]), .A(aux_key_ctrl[20]));
Q_ASSIGN U93 ( .B(kimreader_ckvreader_data[19]), .A(tlv_word0[19]));
Q_ASSIGN U94 ( .B(kimreader_ckvreader_data[19]), .A(tlv_word42[19]));
Q_ASSIGN U95 ( .B(kimreader_ckvreader_data[19]), .A(aux_key_ctrl[19]));
Q_ASSIGN U96 ( .B(kimreader_ckvreader_data[18]), .A(tlv_word0[18]));
Q_ASSIGN U97 ( .B(kimreader_ckvreader_data[18]), .A(tlv_word42[18]));
Q_ASSIGN U98 ( .B(kimreader_ckvreader_data[18]), .A(aux_key_ctrl[18]));
Q_ASSIGN U99 ( .B(kimreader_ckvreader_data[17]), .A(tlv_word0[17]));
Q_ASSIGN U100 ( .B(kimreader_ckvreader_data[17]), .A(tlv_word42[17]));
Q_ASSIGN U101 ( .B(kimreader_ckvreader_data[17]), .A(aux_key_ctrl[17]));
Q_ASSIGN U102 ( .B(kimreader_ckvreader_data[16]), .A(tlv_word0[16]));
Q_ASSIGN U103 ( .B(kimreader_ckvreader_data[16]), .A(tlv_word42[16]));
Q_ASSIGN U104 ( .B(kimreader_ckvreader_data[16]), .A(aux_key_ctrl[16]));
Q_ASSIGN U105 ( .B(kimreader_ckvreader_data[15]), .A(tlv_word0[15]));
Q_ASSIGN U106 ( .B(kimreader_ckvreader_data[15]), .A(tlv_word42[15]));
Q_ASSIGN U107 ( .B(kimreader_ckvreader_data[15]), .A(aux_key_ctrl[15]));
Q_ASSIGN U108 ( .B(kimreader_ckvreader_data[14]), .A(tlv_word0[14]));
Q_ASSIGN U109 ( .B(kimreader_ckvreader_data[14]), .A(tlv_word42[14]));
Q_ASSIGN U110 ( .B(kimreader_ckvreader_data[14]), .A(aux_key_ctrl[14]));
Q_ASSIGN U111 ( .B(kimreader_ckvreader_data[13]), .A(tlv_word0[13]));
Q_ASSIGN U112 ( .B(kimreader_ckvreader_data[13]), .A(tlv_word42[13]));
Q_ASSIGN U113 ( .B(kimreader_ckvreader_data[13]), .A(aux_key_ctrl[13]));
Q_ASSIGN U114 ( .B(kimreader_ckvreader_data[12]), .A(tlv_word0[12]));
Q_ASSIGN U115 ( .B(kimreader_ckvreader_data[12]), .A(tlv_word42[12]));
Q_ASSIGN U116 ( .B(kimreader_ckvreader_data[12]), .A(aux_key_ctrl[12]));
Q_ASSIGN U117 ( .B(kimreader_ckvreader_data[11]), .A(tlv_word0[11]));
Q_ASSIGN U118 ( .B(kimreader_ckvreader_data[11]), .A(tlv_word42[11]));
Q_ASSIGN U119 ( .B(kimreader_ckvreader_data[11]), .A(aux_key_ctrl[11]));
Q_ASSIGN U120 ( .B(kimreader_ckvreader_data[10]), .A(tlv_word0[10]));
Q_ASSIGN U121 ( .B(kimreader_ckvreader_data[10]), .A(tlv_word42[10]));
Q_ASSIGN U122 ( .B(kimreader_ckvreader_data[10]), .A(aux_key_ctrl[10]));
Q_ASSIGN U123 ( .B(kimreader_ckvreader_data[9]), .A(tlv_word0[9]));
Q_ASSIGN U124 ( .B(kimreader_ckvreader_data[9]), .A(tlv_word42[9]));
Q_ASSIGN U125 ( .B(kimreader_ckvreader_data[9]), .A(aux_key_ctrl[9]));
Q_ASSIGN U126 ( .B(kimreader_ckvreader_data[8]), .A(tlv_word0[8]));
Q_ASSIGN U127 ( .B(kimreader_ckvreader_data[8]), .A(tlv_word42[8]));
Q_ASSIGN U128 ( .B(kimreader_ckvreader_data[8]), .A(aux_key_ctrl[8]));
Q_ASSIGN U129 ( .B(kimreader_ckvreader_data[7]), .A(tlv_word0[7]));
Q_ASSIGN U130 ( .B(kimreader_ckvreader_data[7]), .A(aux_key_ctrl[7]));
Q_ASSIGN U131 ( .B(kimreader_ckvreader_data[6]), .A(tlv_word0[6]));
Q_ASSIGN U132 ( .B(kimreader_ckvreader_data[6]), .A(aux_key_ctrl[6]));
Q_ASSIGN U133 ( .B(kimreader_ckvreader_data[5]), .A(tlv_word0[5]));
Q_ASSIGN U134 ( .B(kimreader_ckvreader_data[5]), .A(aux_key_ctrl[5]));
Q_ASSIGN U135 ( .B(kimreader_ckvreader_data[4]), .A(tlv_word0[4]));
Q_ASSIGN U136 ( .B(kimreader_ckvreader_data[4]), .A(aux_key_ctrl[4]));
Q_ASSIGN U137 ( .B(kimreader_ckvreader_data[3]), .A(tlv_word0[3]));
Q_ASSIGN U138 ( .B(kimreader_ckvreader_data[3]), .A(aux_key_ctrl[3]));
Q_ASSIGN U139 ( .B(kimreader_ckvreader_data[2]), .A(tlv_word0[2]));
Q_ASSIGN U140 ( .B(kimreader_ckvreader_data[2]), .A(aux_key_ctrl[2]));
Q_ASSIGN U141 ( .B(kimreader_ckvreader_data[1]), .A(tlv_word0[1]));
Q_ASSIGN U142 ( .B(kimreader_ckvreader_data[1]), .A(aux_key_ctrl[1]));
Q_ASSIGN U143 ( .B(kimreader_ckvreader_data[0]), .A(tlv_word0[0]));
Q_ASSIGN U144 ( .B(kimreader_ckvreader_data[0]), .A(aux_key_ctrl[0]));
Q_BUF U145 ( .A(_zy_sva_brcm_dek_key_3_reset_or), .Z(_zy_sva_brcm_dak_key_2_reset_or));
Q_BUF U146 ( .A(_zy_sva_brcm_dak_key_4_reset_or), .Z(_zy_sva_brcm_dek_key_3_reset_or));
Q_BUF U147 ( .A(_zy_sva_brcm_dek_key_5_reset_or), .Z(_zy_sva_brcm_dak_key_4_reset_or));
Q_BUF U148 ( .A(_zy_sva_brcm_dak_key_6_reset_or), .Z(_zy_sva_brcm_dek_key_5_reset_or));
Q_BUF U149 ( .A(_zy_sva_brcm_dek_key_7_reset_or), .Z(_zy_sva_brcm_dak_key_6_reset_or));
Q_BUF U150 ( .A(_zy_sva_brcm_dak_key_8_reset_or), .Z(_zy_sva_brcm_dek_key_7_reset_or));
Q_BUF U151 ( .A(_zy_sva_brcm_dek_key_1_reset_or), .Z(_zy_sva_brcm_dak_key_8_reset_or));
Q_BUF U152 ( .A(kopassigner_ckvreader_ack), .Z(ckvreader_kimreader_ack));
Q_ASSIGN U153 ( .B(kimreader_ckvreader_data[70]), .A(ckvreader_kopassigner_data[70]));
Q_BUF U154 ( .A(kimreader_ckvreader_data[69]), .Z(ckvreader_kopassigner_data[69]));
Q_ASSIGN U155 ( .B(kimreader_ckvreader_data[68]), .A(ckvreader_kopassigner_data[68]));
Q_BUF U156 ( .A(kimreader_ckvreader_data[67]), .Z(ckvreader_kopassigner_data[67]));
Q_BUF U157 ( .A(kimreader_ckvreader_data[66]), .Z(ckvreader_kopassigner_data[66]));
Q_BUF U158 ( .A(kimreader_ckvreader_data[65]), .Z(ckvreader_kopassigner_data[65]));
Q_BUF U159 ( .A(kimreader_ckvreader_data[64]), .Z(ckvreader_kopassigner_data[64]));
Q_INV U160 ( .A(fifo_out_mbe), .Z(n4));
Q_MX02 U161 ( .S(fifo_out_ack), .A0(n3), .A1(n4), .Z(n5));
Q_ND02 U162 ( .A0(kopassigner_ckvreader_ack), .A1(n419), .Z(n3));
Q_AN02 U163 ( .A0(cur_state[0]), .A1(n385), .Z(n24));
Q_AN02 U164 ( .A0(kimreader_ckvreader_data[66]), .A1(kimreader_ckvreader_data[65]), .Z(n16));
Q_AN02 U165 ( .A0(kimreader_ckvreader_data[64]), .A1(n415), .Z(n15));
Q_AN03 U166 ( .A0(n16), .A1(n15), .A2(n24), .Z(n9));
Q_INV U167 ( .A(kimreader_ckvreader_data[64]), .Z(n17));
Q_AN02 U168 ( .A0(kimreader_ckvreader_data[65]), .A1(n17), .Z(n18));
Q_AO21 U169 ( .A0(n18), .A1(n418), .B0(n19), .Z(n20));
Q_INV U170 ( .A(kimreader_ckvreader_data[65]), .Z(n21));
Q_AN02 U171 ( .A0(kimreader_ckvreader_data[64]), .A1(n406), .Z(n22));
Q_AN02 U172 ( .A0(n21), .A1(n22), .Z(n19));
Q_AN03 U173 ( .A0(n24), .A1(kimreader_ckvreader_data[66]), .A2(n20), .Z(n10));
Q_AN02 U174 ( .A0(kimreader_ckvreader_data[66]), .A1(n21), .Z(n23));
Q_AN03 U175 ( .A0(n23), .A1(n22), .A2(n24), .Z(n26));
Q_AN03 U176 ( .A0(kimreader_ckvreader_valid), .A1(n419), .A2(n382), .Z(n25));
Q_NR03 U177 ( .A0(n9), .A1(n25), .A2(n26), .Z(n27));
Q_AN02 U178 ( .A0(n382), .A1(kimreader_ckvreader_valid), .Z(n34));
Q_AN02 U179 ( .A0(n34), .A1(n8), .Z(n11));
Q_NR02 U180 ( .A0(n8), .A1(n316), .Z(n28));
Q_OR02 U181 ( .A0(n28), .A1(n8), .Z(n29));
Q_ND02 U182 ( .A0(n34), .A1(n29), .Z(n30));
Q_AN02 U183 ( .A0(n34), .A1(n7), .Z(n12));
Q_NR02 U184 ( .A0(n7), .A1(n316), .Z(n31));
Q_OR02 U185 ( .A0(n31), .A1(n7), .Z(n32));
Q_ND02 U186 ( .A0(n34), .A1(n32), .Z(n33));
Q_AN02 U187 ( .A0(n34), .A1(n6), .Z(n13));
Q_MX03 U188 ( .S0(n10), .S1(n9), .A0(n35), .A1(n248), .A2(n184), .Z(ckvreader_kopassigner_data[63]));
Q_AN02 U189 ( .A0(n27), .A1(tlv_word0[63]), .Z(n35));
Q_MX03 U190 ( .S0(n10), .S1(n9), .A0(n36), .A1(n249), .A2(n185), .Z(ckvreader_kopassigner_data[62]));
Q_AN02 U191 ( .A0(n27), .A1(tlv_word0[62]), .Z(n36));
Q_MX03 U192 ( .S0(n10), .S1(n9), .A0(n37), .A1(n250), .A2(n186), .Z(ckvreader_kopassigner_data[61]));
Q_AN02 U193 ( .A0(n27), .A1(tlv_word0[61]), .Z(n37));
Q_MX03 U194 ( .S0(n10), .S1(n9), .A0(n38), .A1(n251), .A2(n187), .Z(ckvreader_kopassigner_data[60]));
Q_AN02 U195 ( .A0(n27), .A1(tlv_word0[60]), .Z(n38));
Q_MX03 U196 ( .S0(n10), .S1(n9), .A0(n39), .A1(n252), .A2(n188), .Z(ckvreader_kopassigner_data[59]));
Q_AN02 U197 ( .A0(n27), .A1(tlv_word0[59]), .Z(n39));
Q_MX03 U198 ( .S0(n10), .S1(n9), .A0(n40), .A1(n253), .A2(n189), .Z(ckvreader_kopassigner_data[58]));
Q_AN02 U199 ( .A0(n27), .A1(tlv_word0[58]), .Z(n40));
Q_MX03 U200 ( .S0(n10), .S1(n9), .A0(n41), .A1(n254), .A2(n190), .Z(ckvreader_kopassigner_data[57]));
Q_AN02 U201 ( .A0(n27), .A1(tlv_word0[57]), .Z(n41));
Q_MX03 U202 ( .S0(n10), .S1(n9), .A0(n42), .A1(n255), .A2(n191), .Z(ckvreader_kopassigner_data[56]));
Q_AN02 U203 ( .A0(n27), .A1(tlv_word0[56]), .Z(n42));
Q_MX03 U204 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[55]), .A1(n256), .A2(n192), .Z(ckvreader_kopassigner_data[55]));
Q_MX03 U205 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[54]), .A1(n257), .A2(n193), .Z(ckvreader_kopassigner_data[54]));
Q_MX03 U206 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[53]), .A1(n258), .A2(n194), .Z(ckvreader_kopassigner_data[53]));
Q_MX03 U207 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[52]), .A1(n259), .A2(n195), .Z(ckvreader_kopassigner_data[52]));
Q_MX03 U208 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[51]), .A1(n260), .A2(n196), .Z(ckvreader_kopassigner_data[51]));
Q_MX03 U209 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[50]), .A1(n261), .A2(n197), .Z(ckvreader_kopassigner_data[50]));
Q_MX03 U210 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[49]), .A1(n262), .A2(n198), .Z(ckvreader_kopassigner_data[49]));
Q_MX03 U211 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[48]), .A1(n263), .A2(n199), .Z(ckvreader_kopassigner_data[48]));
Q_MX03 U212 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[47]), .A1(n264), .A2(n200), .Z(ckvreader_kopassigner_data[47]));
Q_MX03 U213 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[46]), .A1(n265), .A2(n201), .Z(ckvreader_kopassigner_data[46]));
Q_MX03 U214 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[45]), .A1(n266), .A2(n202), .Z(ckvreader_kopassigner_data[45]));
Q_MX03 U215 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[44]), .A1(n267), .A2(n203), .Z(ckvreader_kopassigner_data[44]));
Q_MX03 U216 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[43]), .A1(n268), .A2(n204), .Z(ckvreader_kopassigner_data[43]));
Q_MX03 U217 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[42]), .A1(n269), .A2(n205), .Z(ckvreader_kopassigner_data[42]));
Q_MX03 U218 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[41]), .A1(n270), .A2(n206), .Z(ckvreader_kopassigner_data[41]));
Q_MX03 U219 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[40]), .A1(n271), .A2(n207), .Z(ckvreader_kopassigner_data[40]));
Q_MX03 U220 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[39]), .A1(n272), .A2(n208), .Z(ckvreader_kopassigner_data[39]));
Q_MX03 U221 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[38]), .A1(n273), .A2(n209), .Z(ckvreader_kopassigner_data[38]));
Q_MX03 U222 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[37]), .A1(n274), .A2(n210), .Z(ckvreader_kopassigner_data[37]));
Q_MX03 U223 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[36]), .A1(n275), .A2(n211), .Z(ckvreader_kopassigner_data[36]));
Q_MX03 U224 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[35]), .A1(n276), .A2(n212), .Z(ckvreader_kopassigner_data[35]));
Q_MX03 U225 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[34]), .A1(n277), .A2(n213), .Z(ckvreader_kopassigner_data[34]));
Q_MX03 U226 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[33]), .A1(n278), .A2(n214), .Z(ckvreader_kopassigner_data[33]));
Q_MX03 U227 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[32]), .A1(n279), .A2(n215), .Z(ckvreader_kopassigner_data[32]));
Q_MX03 U228 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[31]), .A1(n280), .A2(n216), .Z(ckvreader_kopassigner_data[31]));
Q_MX03 U229 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[30]), .A1(n281), .A2(n217), .Z(ckvreader_kopassigner_data[30]));
Q_MX03 U230 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[29]), .A1(n282), .A2(n218), .Z(ckvreader_kopassigner_data[29]));
Q_MX03 U231 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[28]), .A1(n283), .A2(n219), .Z(ckvreader_kopassigner_data[28]));
Q_MX03 U232 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[27]), .A1(n284), .A2(n220), .Z(ckvreader_kopassigner_data[27]));
Q_MX03 U233 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[26]), .A1(n285), .A2(n221), .Z(ckvreader_kopassigner_data[26]));
Q_MX03 U234 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[25]), .A1(n286), .A2(n222), .Z(ckvreader_kopassigner_data[25]));
Q_MX03 U235 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[24]), .A1(n287), .A2(n223), .Z(ckvreader_kopassigner_data[24]));
Q_MX03 U236 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[23]), .A1(n288), .A2(n224), .Z(ckvreader_kopassigner_data[23]));
Q_MX03 U237 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[22]), .A1(n289), .A2(n225), .Z(ckvreader_kopassigner_data[22]));
Q_MX03 U238 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[21]), .A1(n290), .A2(n226), .Z(ckvreader_kopassigner_data[21]));
Q_MX03 U239 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[20]), .A1(n291), .A2(n227), .Z(ckvreader_kopassigner_data[20]));
Q_MX03 U240 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[19]), .A1(n292), .A2(n228), .Z(ckvreader_kopassigner_data[19]));
Q_MX03 U241 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[18]), .A1(n293), .A2(n229), .Z(ckvreader_kopassigner_data[18]));
Q_MX03 U242 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[17]), .A1(n294), .A2(n230), .Z(ckvreader_kopassigner_data[17]));
Q_MX03 U243 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[16]), .A1(n295), .A2(n231), .Z(ckvreader_kopassigner_data[16]));
Q_MX03 U244 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[15]), .A1(n296), .A2(n232), .Z(ckvreader_kopassigner_data[15]));
Q_MX03 U245 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[14]), .A1(n297), .A2(n233), .Z(ckvreader_kopassigner_data[14]));
Q_MX03 U246 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[13]), .A1(n298), .A2(n234), .Z(ckvreader_kopassigner_data[13]));
Q_MX03 U247 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[12]), .A1(n299), .A2(n235), .Z(ckvreader_kopassigner_data[12]));
Q_MX03 U248 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[11]), .A1(n300), .A2(n236), .Z(ckvreader_kopassigner_data[11]));
Q_MX03 U249 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[10]), .A1(n301), .A2(n237), .Z(ckvreader_kopassigner_data[10]));
Q_MX03 U250 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[9]), .A1(n302), .A2(n238), .Z(ckvreader_kopassigner_data[9]));
Q_MX03 U251 ( .S0(n10), .S1(n9), .A0(kimreader_ckvreader_data[8]), .A1(n303), .A2(n239), .Z(ckvreader_kopassigner_data[8]));
Q_MX02 U252 ( .S(n9), .A0(n43), .A1(n240), .Z(ckvreader_kopassigner_data[7]));
Q_MX02 U253 ( .S(n9), .A0(n44), .A1(n241), .Z(ckvreader_kopassigner_data[6]));
Q_MX02 U254 ( .S(n9), .A0(n45), .A1(n242), .Z(ckvreader_kopassigner_data[5]));
Q_MX02 U255 ( .S(n9), .A0(n46), .A1(n243), .Z(ckvreader_kopassigner_data[4]));
Q_MX02 U256 ( .S(n9), .A0(n47), .A1(n244), .Z(ckvreader_kopassigner_data[3]));
Q_MX02 U257 ( .S(n9), .A0(n48), .A1(n245), .Z(ckvreader_kopassigner_data[2]));
Q_MX02 U258 ( .S(n9), .A0(n49), .A1(n246), .Z(ckvreader_kopassigner_data[1]));
Q_MX02 U259 ( .S(n9), .A0(n50), .A1(n247), .Z(ckvreader_kopassigner_data[0]));
Q_AN02 U260 ( .A0(cur_state[0]), .A1(n179), .Z(ckv_rd));
Q_MX02 U261 ( .S(n11), .A0(n51), .A1(tlv_word0[63]), .Z(nxt_tlv_word8[63]));
Q_AN02 U262 ( .A0(n30), .A1(tlv_word8[63]), .Z(n51));
Q_MX02 U263 ( .S(n11), .A0(n52), .A1(tlv_word0[62]), .Z(nxt_tlv_word8[62]));
Q_AN02 U264 ( .A0(n30), .A1(tlv_word8[62]), .Z(n52));
Q_MX02 U265 ( .S(n11), .A0(n53), .A1(tlv_word0[61]), .Z(nxt_tlv_word8[61]));
Q_AN02 U266 ( .A0(n30), .A1(tlv_word8[61]), .Z(n53));
Q_MX02 U267 ( .S(n11), .A0(n54), .A1(tlv_word0[60]), .Z(nxt_tlv_word8[60]));
Q_AN02 U268 ( .A0(n30), .A1(tlv_word8[60]), .Z(n54));
Q_MX02 U269 ( .S(n11), .A0(n55), .A1(tlv_word0[59]), .Z(nxt_tlv_word8[59]));
Q_AN02 U270 ( .A0(n30), .A1(tlv_word8[59]), .Z(n55));
Q_MX02 U271 ( .S(n11), .A0(n56), .A1(tlv_word0[58]), .Z(nxt_tlv_word8[58]));
Q_AN02 U272 ( .A0(n30), .A1(tlv_word8[58]), .Z(n56));
Q_MX02 U273 ( .S(n11), .A0(n57), .A1(tlv_word0[57]), .Z(nxt_tlv_word8[57]));
Q_AN02 U274 ( .A0(n30), .A1(tlv_word8[57]), .Z(n57));
Q_MX02 U275 ( .S(n11), .A0(n58), .A1(tlv_word0[56]), .Z(nxt_tlv_word8[56]));
Q_AN02 U276 ( .A0(n30), .A1(tlv_word8[56]), .Z(n58));
Q_MX02 U277 ( .S(n11), .A0(n59), .A1(kimreader_ckvreader_data[55]), .Z(nxt_tlv_word8[55]));
Q_AN02 U278 ( .A0(n30), .A1(tlv_word8[55]), .Z(n59));
Q_MX02 U279 ( .S(n11), .A0(n60), .A1(kimreader_ckvreader_data[54]), .Z(nxt_tlv_word8[54]));
Q_AN02 U280 ( .A0(n30), .A1(tlv_word8[54]), .Z(n60));
Q_MX02 U281 ( .S(n11), .A0(n61), .A1(kimreader_ckvreader_data[53]), .Z(nxt_tlv_word8[53]));
Q_AN02 U282 ( .A0(n30), .A1(tlv_word8[53]), .Z(n61));
Q_MX02 U283 ( .S(n11), .A0(n62), .A1(kimreader_ckvreader_data[52]), .Z(nxt_tlv_word8[52]));
Q_AN02 U284 ( .A0(n30), .A1(tlv_word8[52]), .Z(n62));
Q_MX02 U285 ( .S(n11), .A0(n63), .A1(kimreader_ckvreader_data[51]), .Z(nxt_tlv_word8[51]));
Q_AN02 U286 ( .A0(n30), .A1(tlv_word8[51]), .Z(n63));
Q_MX02 U287 ( .S(n11), .A0(n64), .A1(kimreader_ckvreader_data[50]), .Z(nxt_tlv_word8[50]));
Q_AN02 U288 ( .A0(n30), .A1(tlv_word8[50]), .Z(n64));
Q_MX02 U289 ( .S(n11), .A0(n65), .A1(kimreader_ckvreader_data[49]), .Z(nxt_tlv_word8[49]));
Q_AN02 U290 ( .A0(n30), .A1(tlv_word8[49]), .Z(n65));
Q_MX02 U291 ( .S(n11), .A0(n66), .A1(kimreader_ckvreader_data[48]), .Z(nxt_tlv_word8[48]));
Q_AN02 U292 ( .A0(n30), .A1(tlv_word8[48]), .Z(n66));
Q_MX02 U293 ( .S(n11), .A0(n67), .A1(kimreader_ckvreader_data[47]), .Z(nxt_tlv_word8[47]));
Q_AN02 U294 ( .A0(n30), .A1(tlv_word8[47]), .Z(n67));
Q_MX02 U295 ( .S(n11), .A0(n68), .A1(kimreader_ckvreader_data[46]), .Z(nxt_tlv_word8[46]));
Q_AN02 U296 ( .A0(n30), .A1(tlv_word8[46]), .Z(n68));
Q_MX02 U297 ( .S(n11), .A0(n69), .A1(kimreader_ckvreader_data[45]), .Z(nxt_tlv_word8[45]));
Q_AN02 U298 ( .A0(n30), .A1(tlv_word8[45]), .Z(n69));
Q_MX02 U299 ( .S(n11), .A0(n70), .A1(kimreader_ckvreader_data[44]), .Z(nxt_tlv_word8[44]));
Q_AN02 U300 ( .A0(n30), .A1(tlv_word8[44]), .Z(n70));
Q_MX02 U301 ( .S(n11), .A0(n71), .A1(kimreader_ckvreader_data[43]), .Z(nxt_tlv_word8[43]));
Q_AN02 U302 ( .A0(n30), .A1(tlv_word8[43]), .Z(n71));
Q_MX02 U303 ( .S(n11), .A0(n72), .A1(kimreader_ckvreader_data[42]), .Z(nxt_tlv_word8[42]));
Q_AN02 U304 ( .A0(n30), .A1(tlv_word8[42]), .Z(n72));
Q_MX02 U305 ( .S(n11), .A0(n73), .A1(kimreader_ckvreader_data[41]), .Z(nxt_tlv_word8[41]));
Q_AN02 U306 ( .A0(n30), .A1(tlv_word8[41]), .Z(n73));
Q_MX02 U307 ( .S(n11), .A0(n74), .A1(kimreader_ckvreader_data[40]), .Z(nxt_tlv_word8[40]));
Q_AN02 U308 ( .A0(n30), .A1(tlv_word8[40]), .Z(n74));
Q_MX02 U309 ( .S(n11), .A0(n75), .A1(kimreader_ckvreader_data[39]), .Z(nxt_tlv_word8[39]));
Q_AN02 U310 ( .A0(n30), .A1(tlv_word8[39]), .Z(n75));
Q_MX02 U311 ( .S(n11), .A0(n76), .A1(kimreader_ckvreader_data[38]), .Z(nxt_tlv_word8[38]));
Q_AN02 U312 ( .A0(n30), .A1(tlv_word8[38]), .Z(n76));
Q_MX02 U313 ( .S(n11), .A0(n77), .A1(kimreader_ckvreader_data[37]), .Z(nxt_tlv_word8[37]));
Q_AN02 U314 ( .A0(n30), .A1(tlv_word8[37]), .Z(n77));
Q_MX02 U315 ( .S(n11), .A0(n78), .A1(kimreader_ckvreader_data[36]), .Z(nxt_tlv_word8[36]));
Q_AN02 U316 ( .A0(n30), .A1(tlv_word8[36]), .Z(n78));
Q_MX02 U317 ( .S(n11), .A0(n79), .A1(kimreader_ckvreader_data[35]), .Z(nxt_tlv_word8[35]));
Q_AN02 U318 ( .A0(n30), .A1(tlv_word8[35]), .Z(n79));
Q_MX02 U319 ( .S(n11), .A0(n80), .A1(kimreader_ckvreader_data[34]), .Z(nxt_tlv_word8[34]));
Q_AN02 U320 ( .A0(n30), .A1(tlv_word8[34]), .Z(n80));
Q_MX02 U321 ( .S(n11), .A0(n81), .A1(kimreader_ckvreader_data[33]), .Z(nxt_tlv_word8[33]));
Q_AN02 U322 ( .A0(n30), .A1(tlv_word8[33]), .Z(n81));
Q_MX02 U323 ( .S(n11), .A0(n82), .A1(kimreader_ckvreader_data[32]), .Z(nxt_tlv_word8[32]));
Q_AN02 U324 ( .A0(n30), .A1(tlv_word8[32]), .Z(n82));
Q_MX02 U325 ( .S(n11), .A0(n83), .A1(kimreader_ckvreader_data[31]), .Z(nxt_tlv_word8[31]));
Q_AN02 U326 ( .A0(n30), .A1(tlv_word8[31]), .Z(n83));
Q_MX02 U327 ( .S(n11), .A0(n84), .A1(kimreader_ckvreader_data[30]), .Z(nxt_tlv_word8[30]));
Q_AN02 U328 ( .A0(n30), .A1(tlv_word8[30]), .Z(n84));
Q_MX02 U329 ( .S(n11), .A0(n85), .A1(kimreader_ckvreader_data[29]), .Z(nxt_tlv_word8[29]));
Q_AN02 U330 ( .A0(n30), .A1(tlv_word8[29]), .Z(n85));
Q_MX02 U331 ( .S(n11), .A0(n86), .A1(kimreader_ckvreader_data[28]), .Z(nxt_tlv_word8[28]));
Q_AN02 U332 ( .A0(n30), .A1(tlv_word8[28]), .Z(n86));
Q_MX02 U333 ( .S(n11), .A0(n87), .A1(kimreader_ckvreader_data[27]), .Z(nxt_tlv_word8[27]));
Q_AN02 U334 ( .A0(n30), .A1(tlv_word8[27]), .Z(n87));
Q_MX02 U335 ( .S(n11), .A0(n88), .A1(kimreader_ckvreader_data[26]), .Z(nxt_tlv_word8[26]));
Q_AN02 U336 ( .A0(n30), .A1(tlv_word8[26]), .Z(n88));
Q_MX02 U337 ( .S(n11), .A0(n89), .A1(kimreader_ckvreader_data[25]), .Z(nxt_tlv_word8[25]));
Q_AN02 U338 ( .A0(n30), .A1(tlv_word8[25]), .Z(n89));
Q_MX02 U339 ( .S(n11), .A0(n90), .A1(kimreader_ckvreader_data[24]), .Z(nxt_tlv_word8[24]));
Q_AN02 U340 ( .A0(n30), .A1(tlv_word8[24]), .Z(n90));
Q_MX02 U341 ( .S(n11), .A0(n91), .A1(kimreader_ckvreader_data[23]), .Z(nxt_tlv_word8[23]));
Q_AN02 U342 ( .A0(n30), .A1(tlv_word8[23]), .Z(n91));
Q_MX02 U343 ( .S(n11), .A0(n92), .A1(kimreader_ckvreader_data[22]), .Z(nxt_tlv_word8[22]));
Q_AN02 U344 ( .A0(n30), .A1(tlv_word8[22]), .Z(n92));
Q_MX02 U345 ( .S(n11), .A0(n93), .A1(kimreader_ckvreader_data[21]), .Z(nxt_tlv_word8[21]));
Q_AN02 U346 ( .A0(n30), .A1(tlv_word8[21]), .Z(n93));
Q_MX02 U347 ( .S(n11), .A0(n94), .A1(kimreader_ckvreader_data[20]), .Z(nxt_tlv_word8[20]));
Q_AN02 U348 ( .A0(n30), .A1(tlv_word8[20]), .Z(n94));
Q_MX02 U349 ( .S(n11), .A0(n95), .A1(kimreader_ckvreader_data[19]), .Z(nxt_tlv_word8[19]));
Q_AN02 U350 ( .A0(n30), .A1(tlv_word8[19]), .Z(n95));
Q_MX02 U351 ( .S(n11), .A0(n96), .A1(kimreader_ckvreader_data[18]), .Z(nxt_tlv_word8[18]));
Q_AN02 U352 ( .A0(n30), .A1(tlv_word8[18]), .Z(n96));
Q_MX02 U353 ( .S(n11), .A0(n97), .A1(kimreader_ckvreader_data[17]), .Z(nxt_tlv_word8[17]));
Q_AN02 U354 ( .A0(n30), .A1(tlv_word8[17]), .Z(n97));
Q_MX02 U355 ( .S(n11), .A0(n98), .A1(kimreader_ckvreader_data[16]), .Z(nxt_tlv_word8[16]));
Q_AN02 U356 ( .A0(n30), .A1(tlv_word8[16]), .Z(n98));
Q_MX02 U357 ( .S(n11), .A0(n99), .A1(kimreader_ckvreader_data[15]), .Z(nxt_tlv_word8[15]));
Q_AN02 U358 ( .A0(n30), .A1(tlv_word8[15]), .Z(n99));
Q_MX02 U359 ( .S(n11), .A0(n100), .A1(kimreader_ckvreader_data[14]), .Z(nxt_tlv_word8[14]));
Q_AN02 U360 ( .A0(n30), .A1(tlv_word8[14]), .Z(n100));
Q_MX02 U361 ( .S(n11), .A0(n101), .A1(kimreader_ckvreader_data[13]), .Z(nxt_tlv_word8[13]));
Q_AN02 U362 ( .A0(n30), .A1(tlv_word8[13]), .Z(n101));
Q_MX02 U363 ( .S(n11), .A0(n102), .A1(kimreader_ckvreader_data[12]), .Z(nxt_tlv_word8[12]));
Q_AN02 U364 ( .A0(n30), .A1(tlv_word8[12]), .Z(n102));
Q_MX02 U365 ( .S(n11), .A0(n103), .A1(kimreader_ckvreader_data[11]), .Z(nxt_tlv_word8[11]));
Q_AN02 U366 ( .A0(n30), .A1(tlv_word8[11]), .Z(n103));
Q_MX02 U367 ( .S(n11), .A0(n104), .A1(kimreader_ckvreader_data[10]), .Z(nxt_tlv_word8[10]));
Q_AN02 U368 ( .A0(n30), .A1(tlv_word8[10]), .Z(n104));
Q_MX02 U369 ( .S(n11), .A0(n105), .A1(kimreader_ckvreader_data[9]), .Z(nxt_tlv_word8[9]));
Q_AN02 U370 ( .A0(n30), .A1(tlv_word8[9]), .Z(n105));
Q_MX02 U371 ( .S(n11), .A0(n106), .A1(kimreader_ckvreader_data[8]), .Z(nxt_tlv_word8[8]));
Q_AN02 U372 ( .A0(n30), .A1(tlv_word8[8]), .Z(n106));
Q_MX02 U373 ( .S(n11), .A0(n107), .A1(kimreader_ckvreader_data[7]), .Z(nxt_tlv_word8[7]));
Q_AN02 U374 ( .A0(n30), .A1(tlv_word8[7]), .Z(n107));
Q_MX02 U375 ( .S(n11), .A0(n108), .A1(kimreader_ckvreader_data[6]), .Z(nxt_tlv_word8[6]));
Q_AN02 U376 ( .A0(n30), .A1(tlv_word8[6]), .Z(n108));
Q_MX02 U377 ( .S(n11), .A0(n109), .A1(kimreader_ckvreader_data[5]), .Z(nxt_tlv_word8[5]));
Q_AN02 U378 ( .A0(n30), .A1(tlv_word8[5]), .Z(n109));
Q_MX02 U379 ( .S(n11), .A0(n110), .A1(kimreader_ckvreader_data[4]), .Z(nxt_tlv_word8[4]));
Q_AN02 U380 ( .A0(n30), .A1(tlv_word8[4]), .Z(n110));
Q_MX02 U381 ( .S(n11), .A0(n111), .A1(kimreader_ckvreader_data[3]), .Z(nxt_tlv_word8[3]));
Q_AN02 U382 ( .A0(n30), .A1(tlv_word8[3]), .Z(n111));
Q_MX02 U383 ( .S(n11), .A0(n112), .A1(kimreader_ckvreader_data[2]), .Z(nxt_tlv_word8[2]));
Q_AN02 U384 ( .A0(n30), .A1(tlv_word8[2]), .Z(n112));
Q_MX02 U385 ( .S(n11), .A0(n113), .A1(kimreader_ckvreader_data[1]), .Z(nxt_tlv_word8[1]));
Q_AN02 U386 ( .A0(n30), .A1(tlv_word8[1]), .Z(n113));
Q_MX02 U387 ( .S(n11), .A0(n114), .A1(kimreader_ckvreader_data[0]), .Z(nxt_tlv_word8[0]));
Q_AN02 U388 ( .A0(n30), .A1(tlv_word8[0]), .Z(n114));
Q_MX02 U389 ( .S(n12), .A0(n115), .A1(tlv_word0[63]), .Z(nxt_tlv_word9[63]));
Q_AN02 U390 ( .A0(n33), .A1(tlv_word9[63]), .Z(n115));
Q_MX02 U391 ( .S(n12), .A0(n116), .A1(tlv_word0[62]), .Z(nxt_tlv_word9[62]));
Q_AN02 U392 ( .A0(n33), .A1(tlv_word9[62]), .Z(n116));
Q_MX02 U393 ( .S(n12), .A0(n117), .A1(tlv_word0[61]), .Z(nxt_tlv_word9[61]));
Q_AN02 U394 ( .A0(n33), .A1(tlv_word9[61]), .Z(n117));
Q_MX02 U395 ( .S(n12), .A0(n118), .A1(tlv_word0[60]), .Z(nxt_tlv_word9[60]));
Q_AN02 U396 ( .A0(n33), .A1(tlv_word9[60]), .Z(n118));
Q_MX02 U397 ( .S(n12), .A0(n119), .A1(tlv_word0[59]), .Z(nxt_tlv_word9[59]));
Q_AN02 U398 ( .A0(n33), .A1(tlv_word9[59]), .Z(n119));
Q_MX02 U399 ( .S(n12), .A0(n120), .A1(tlv_word0[58]), .Z(nxt_tlv_word9[58]));
Q_AN02 U400 ( .A0(n33), .A1(tlv_word9[58]), .Z(n120));
Q_MX02 U401 ( .S(n12), .A0(n121), .A1(tlv_word0[57]), .Z(nxt_tlv_word9[57]));
Q_AN02 U402 ( .A0(n33), .A1(tlv_word9[57]), .Z(n121));
Q_MX02 U403 ( .S(n12), .A0(n122), .A1(tlv_word0[56]), .Z(nxt_tlv_word9[56]));
Q_AN02 U404 ( .A0(n33), .A1(tlv_word9[56]), .Z(n122));
Q_MX02 U405 ( .S(n12), .A0(n123), .A1(kimreader_ckvreader_data[55]), .Z(nxt_tlv_word9[55]));
Q_AN02 U406 ( .A0(n33), .A1(tlv_word9[55]), .Z(n123));
Q_MX02 U407 ( .S(n12), .A0(n124), .A1(kimreader_ckvreader_data[54]), .Z(nxt_tlv_word9[54]));
Q_AN02 U408 ( .A0(n33), .A1(tlv_word9[54]), .Z(n124));
Q_MX02 U409 ( .S(n12), .A0(n125), .A1(kimreader_ckvreader_data[53]), .Z(nxt_tlv_word9[53]));
Q_AN02 U410 ( .A0(n33), .A1(tlv_word9[53]), .Z(n125));
Q_MX02 U411 ( .S(n12), .A0(n126), .A1(kimreader_ckvreader_data[52]), .Z(nxt_tlv_word9[52]));
Q_AN02 U412 ( .A0(n33), .A1(tlv_word9[52]), .Z(n126));
Q_MX02 U413 ( .S(n12), .A0(n127), .A1(kimreader_ckvreader_data[51]), .Z(nxt_tlv_word9[51]));
Q_AN02 U414 ( .A0(n33), .A1(tlv_word9[51]), .Z(n127));
Q_MX02 U415 ( .S(n12), .A0(n128), .A1(kimreader_ckvreader_data[50]), .Z(nxt_tlv_word9[50]));
Q_AN02 U416 ( .A0(n33), .A1(tlv_word9[50]), .Z(n128));
Q_MX02 U417 ( .S(n12), .A0(n129), .A1(kimreader_ckvreader_data[49]), .Z(nxt_tlv_word9[49]));
Q_AN02 U418 ( .A0(n33), .A1(tlv_word9[49]), .Z(n129));
Q_MX02 U419 ( .S(n12), .A0(n130), .A1(kimreader_ckvreader_data[48]), .Z(nxt_tlv_word9[48]));
Q_AN02 U420 ( .A0(n33), .A1(tlv_word9[48]), .Z(n130));
Q_MX02 U421 ( .S(n12), .A0(n131), .A1(kimreader_ckvreader_data[47]), .Z(nxt_tlv_word9[47]));
Q_AN02 U422 ( .A0(n33), .A1(tlv_word9[47]), .Z(n131));
Q_MX02 U423 ( .S(n12), .A0(n132), .A1(kimreader_ckvreader_data[46]), .Z(nxt_tlv_word9[46]));
Q_AN02 U424 ( .A0(n33), .A1(tlv_word9[46]), .Z(n132));
Q_MX02 U425 ( .S(n12), .A0(n133), .A1(kimreader_ckvreader_data[45]), .Z(nxt_tlv_word9[45]));
Q_AN02 U426 ( .A0(n33), .A1(tlv_word9[45]), .Z(n133));
Q_MX02 U427 ( .S(n12), .A0(n134), .A1(kimreader_ckvreader_data[44]), .Z(nxt_tlv_word9[44]));
Q_AN02 U428 ( .A0(n33), .A1(tlv_word9[44]), .Z(n134));
Q_MX02 U429 ( .S(n12), .A0(n135), .A1(kimreader_ckvreader_data[43]), .Z(nxt_tlv_word9[43]));
Q_AN02 U430 ( .A0(n33), .A1(tlv_word9[43]), .Z(n135));
Q_MX02 U431 ( .S(n12), .A0(n136), .A1(kimreader_ckvreader_data[42]), .Z(nxt_tlv_word9[42]));
Q_AN02 U432 ( .A0(n33), .A1(tlv_word9[42]), .Z(n136));
Q_MX02 U433 ( .S(n12), .A0(n137), .A1(kimreader_ckvreader_data[41]), .Z(nxt_tlv_word9[41]));
Q_AN02 U434 ( .A0(n33), .A1(tlv_word9[41]), .Z(n137));
Q_MX02 U435 ( .S(n12), .A0(n138), .A1(kimreader_ckvreader_data[40]), .Z(nxt_tlv_word9[40]));
Q_AN02 U436 ( .A0(n33), .A1(tlv_word9[40]), .Z(n138));
Q_MX02 U437 ( .S(n12), .A0(n139), .A1(kimreader_ckvreader_data[39]), .Z(nxt_tlv_word9[39]));
Q_AN02 U438 ( .A0(n33), .A1(tlv_word9[39]), .Z(n139));
Q_MX02 U439 ( .S(n12), .A0(n140), .A1(kimreader_ckvreader_data[38]), .Z(nxt_tlv_word9[38]));
Q_AN02 U440 ( .A0(n33), .A1(tlv_word9[38]), .Z(n140));
Q_MX02 U441 ( .S(n12), .A0(n141), .A1(kimreader_ckvreader_data[37]), .Z(nxt_tlv_word9[37]));
Q_AN02 U442 ( .A0(n33), .A1(tlv_word9[37]), .Z(n141));
Q_MX02 U443 ( .S(n12), .A0(n142), .A1(kimreader_ckvreader_data[36]), .Z(nxt_tlv_word9[36]));
Q_AN02 U444 ( .A0(n33), .A1(tlv_word9[36]), .Z(n142));
Q_MX02 U445 ( .S(n12), .A0(n143), .A1(kimreader_ckvreader_data[35]), .Z(nxt_tlv_word9[35]));
Q_AN02 U446 ( .A0(n33), .A1(tlv_word9[35]), .Z(n143));
Q_MX02 U447 ( .S(n12), .A0(n144), .A1(kimreader_ckvreader_data[34]), .Z(nxt_tlv_word9[34]));
Q_AN02 U448 ( .A0(n33), .A1(tlv_word9[34]), .Z(n144));
Q_MX02 U449 ( .S(n12), .A0(n145), .A1(kimreader_ckvreader_data[33]), .Z(nxt_tlv_word9[33]));
Q_AN02 U450 ( .A0(n33), .A1(tlv_word9[33]), .Z(n145));
Q_MX02 U451 ( .S(n12), .A0(n146), .A1(kimreader_ckvreader_data[32]), .Z(nxt_tlv_word9[32]));
Q_AN02 U452 ( .A0(n33), .A1(tlv_word9[32]), .Z(n146));
Q_MX02 U453 ( .S(n12), .A0(n147), .A1(kimreader_ckvreader_data[31]), .Z(nxt_tlv_word9[31]));
Q_AN02 U454 ( .A0(n33), .A1(tlv_word9[31]), .Z(n147));
Q_MX02 U455 ( .S(n12), .A0(n148), .A1(kimreader_ckvreader_data[30]), .Z(nxt_tlv_word9[30]));
Q_AN02 U456 ( .A0(n33), .A1(tlv_word9[30]), .Z(n148));
Q_MX02 U457 ( .S(n12), .A0(n149), .A1(kimreader_ckvreader_data[29]), .Z(nxt_tlv_word9[29]));
Q_AN02 U458 ( .A0(n33), .A1(tlv_word9[29]), .Z(n149));
Q_MX02 U459 ( .S(n12), .A0(n150), .A1(kimreader_ckvreader_data[28]), .Z(nxt_tlv_word9[28]));
Q_AN02 U460 ( .A0(n33), .A1(tlv_word9[28]), .Z(n150));
Q_MX02 U461 ( .S(n12), .A0(n151), .A1(kimreader_ckvreader_data[27]), .Z(nxt_tlv_word9[27]));
Q_AN02 U462 ( .A0(n33), .A1(tlv_word9[27]), .Z(n151));
Q_MX02 U463 ( .S(n12), .A0(n152), .A1(kimreader_ckvreader_data[26]), .Z(nxt_tlv_word9[26]));
Q_AN02 U464 ( .A0(n33), .A1(tlv_word9[26]), .Z(n152));
Q_MX02 U465 ( .S(n12), .A0(n153), .A1(kimreader_ckvreader_data[25]), .Z(nxt_tlv_word9[25]));
Q_AN02 U466 ( .A0(n33), .A1(tlv_word9[25]), .Z(n153));
Q_MX02 U467 ( .S(n12), .A0(n154), .A1(kimreader_ckvreader_data[24]), .Z(nxt_tlv_word9[24]));
Q_AN02 U468 ( .A0(n33), .A1(tlv_word9[24]), .Z(n154));
Q_MX02 U469 ( .S(n12), .A0(n155), .A1(kimreader_ckvreader_data[23]), .Z(nxt_tlv_word9[23]));
Q_AN02 U470 ( .A0(n33), .A1(tlv_word9[23]), .Z(n155));
Q_MX02 U471 ( .S(n12), .A0(n156), .A1(kimreader_ckvreader_data[22]), .Z(nxt_tlv_word9[22]));
Q_AN02 U472 ( .A0(n33), .A1(tlv_word9[22]), .Z(n156));
Q_MX02 U473 ( .S(n12), .A0(n157), .A1(kimreader_ckvreader_data[21]), .Z(nxt_tlv_word9[21]));
Q_AN02 U474 ( .A0(n33), .A1(tlv_word9[21]), .Z(n157));
Q_MX02 U475 ( .S(n12), .A0(n158), .A1(kimreader_ckvreader_data[20]), .Z(nxt_tlv_word9[20]));
Q_AN02 U476 ( .A0(n33), .A1(tlv_word9[20]), .Z(n158));
Q_MX02 U477 ( .S(n12), .A0(n159), .A1(kimreader_ckvreader_data[19]), .Z(nxt_tlv_word9[19]));
Q_AN02 U478 ( .A0(n33), .A1(tlv_word9[19]), .Z(n159));
Q_MX02 U479 ( .S(n12), .A0(n160), .A1(kimreader_ckvreader_data[18]), .Z(nxt_tlv_word9[18]));
Q_AN02 U480 ( .A0(n33), .A1(tlv_word9[18]), .Z(n160));
Q_MX02 U481 ( .S(n12), .A0(n161), .A1(kimreader_ckvreader_data[17]), .Z(nxt_tlv_word9[17]));
Q_AN02 U482 ( .A0(n33), .A1(tlv_word9[17]), .Z(n161));
Q_MX02 U483 ( .S(n12), .A0(n162), .A1(kimreader_ckvreader_data[16]), .Z(nxt_tlv_word9[16]));
Q_AN02 U484 ( .A0(n33), .A1(tlv_word9[16]), .Z(n162));
Q_MX02 U485 ( .S(n12), .A0(n163), .A1(kimreader_ckvreader_data[15]), .Z(nxt_tlv_word9[15]));
Q_AN02 U486 ( .A0(n33), .A1(tlv_word9[15]), .Z(n163));
Q_MX02 U487 ( .S(n12), .A0(n164), .A1(kimreader_ckvreader_data[14]), .Z(nxt_tlv_word9[14]));
Q_AN02 U488 ( .A0(n33), .A1(tlv_word9[14]), .Z(n164));
Q_MX02 U489 ( .S(n12), .A0(n165), .A1(kimreader_ckvreader_data[13]), .Z(nxt_tlv_word9[13]));
Q_AN02 U490 ( .A0(n33), .A1(tlv_word9[13]), .Z(n165));
Q_MX02 U491 ( .S(n12), .A0(n166), .A1(kimreader_ckvreader_data[12]), .Z(nxt_tlv_word9[12]));
Q_AN02 U492 ( .A0(n33), .A1(tlv_word9[12]), .Z(n166));
Q_MX02 U493 ( .S(n12), .A0(n167), .A1(kimreader_ckvreader_data[11]), .Z(nxt_tlv_word9[11]));
Q_AN02 U494 ( .A0(n33), .A1(tlv_word9[11]), .Z(n167));
Q_MX02 U495 ( .S(n12), .A0(n168), .A1(kimreader_ckvreader_data[10]), .Z(nxt_tlv_word9[10]));
Q_AN02 U496 ( .A0(n33), .A1(tlv_word9[10]), .Z(n168));
Q_MX02 U497 ( .S(n12), .A0(n169), .A1(kimreader_ckvreader_data[9]), .Z(nxt_tlv_word9[9]));
Q_AN02 U498 ( .A0(n33), .A1(tlv_word9[9]), .Z(n169));
Q_MX02 U499 ( .S(n12), .A0(n170), .A1(kimreader_ckvreader_data[8]), .Z(nxt_tlv_word9[8]));
Q_AN02 U500 ( .A0(n33), .A1(tlv_word9[8]), .Z(n170));
Q_MX02 U501 ( .S(n12), .A0(n171), .A1(kimreader_ckvreader_data[7]), .Z(nxt_tlv_word9[7]));
Q_AN02 U502 ( .A0(n33), .A1(tlv_word9[7]), .Z(n171));
Q_MX02 U503 ( .S(n12), .A0(n172), .A1(kimreader_ckvreader_data[6]), .Z(nxt_tlv_word9[6]));
Q_AN02 U504 ( .A0(n33), .A1(tlv_word9[6]), .Z(n172));
Q_MX02 U505 ( .S(n12), .A0(n173), .A1(kimreader_ckvreader_data[5]), .Z(nxt_tlv_word9[5]));
Q_AN02 U506 ( .A0(n33), .A1(tlv_word9[5]), .Z(n173));
Q_MX02 U507 ( .S(n12), .A0(n174), .A1(kimreader_ckvreader_data[4]), .Z(nxt_tlv_word9[4]));
Q_AN02 U508 ( .A0(n33), .A1(tlv_word9[4]), .Z(n174));
Q_MX02 U509 ( .S(n12), .A0(n175), .A1(kimreader_ckvreader_data[3]), .Z(nxt_tlv_word9[3]));
Q_AN02 U510 ( .A0(n33), .A1(tlv_word9[3]), .Z(n175));
Q_MX02 U511 ( .S(n12), .A0(n176), .A1(kimreader_ckvreader_data[2]), .Z(nxt_tlv_word9[2]));
Q_AN02 U512 ( .A0(n33), .A1(tlv_word9[2]), .Z(n176));
Q_MX02 U513 ( .S(n12), .A0(n177), .A1(kimreader_ckvreader_data[1]), .Z(nxt_tlv_word9[1]));
Q_AN02 U514 ( .A0(n33), .A1(tlv_word9[1]), .Z(n177));
Q_MX02 U515 ( .S(n12), .A0(n178), .A1(kimreader_ckvreader_data[0]), .Z(nxt_tlv_word9[0]));
Q_AN02 U516 ( .A0(n33), .A1(tlv_word9[0]), .Z(n178));
Q_MX02 U517 ( .S(n13), .A0(ktype_is_aux_key_only), .A1(n312), .Z(nxt_ktype_is_aux_key_only));
Q_AN02 U518 ( .A0(cur_state[0]), .A1(kopassigner_ckvreader_ack), .Z(fifo_out_ack));
Q_ND02 U519 ( .A0(n351), .A1(n181), .Z(n180));
Q_AN03 U520 ( .A0(ckv_read_num[3]), .A1(ckv_read_num[2]), .A2(n182), .Z(n181));
Q_OA21 U521 ( .A0(n183), .A1(kopassigner_ckvreader_ack), .B0(n180), .Z(n179));
Q_INV U522 ( .A(fifo_in_stall), .Z(n183));
Q_AN02 U523 ( .A0(tlv_word9[17]), .A1(fifo_out[63]), .Z(n184));
Q_AN02 U524 ( .A0(tlv_word9[17]), .A1(fifo_out[62]), .Z(n185));
Q_AN02 U525 ( .A0(tlv_word9[17]), .A1(fifo_out[61]), .Z(n186));
Q_AN02 U526 ( .A0(tlv_word9[17]), .A1(fifo_out[60]), .Z(n187));
Q_AN02 U527 ( .A0(tlv_word9[17]), .A1(fifo_out[59]), .Z(n188));
Q_AN02 U528 ( .A0(tlv_word9[17]), .A1(fifo_out[58]), .Z(n189));
Q_AN02 U529 ( .A0(tlv_word9[17]), .A1(fifo_out[57]), .Z(n190));
Q_AN02 U530 ( .A0(tlv_word9[17]), .A1(fifo_out[56]), .Z(n191));
Q_AN02 U531 ( .A0(tlv_word9[17]), .A1(fifo_out[55]), .Z(n192));
Q_AN02 U532 ( .A0(tlv_word9[17]), .A1(fifo_out[54]), .Z(n193));
Q_AN02 U533 ( .A0(tlv_word9[17]), .A1(fifo_out[53]), .Z(n194));
Q_AN02 U534 ( .A0(tlv_word9[17]), .A1(fifo_out[52]), .Z(n195));
Q_AN02 U535 ( .A0(tlv_word9[17]), .A1(fifo_out[51]), .Z(n196));
Q_AN02 U536 ( .A0(tlv_word9[17]), .A1(fifo_out[50]), .Z(n197));
Q_AN02 U537 ( .A0(tlv_word9[17]), .A1(fifo_out[49]), .Z(n198));
Q_AN02 U538 ( .A0(tlv_word9[17]), .A1(fifo_out[48]), .Z(n199));
Q_AN02 U539 ( .A0(tlv_word9[17]), .A1(fifo_out[47]), .Z(n200));
Q_AN02 U540 ( .A0(tlv_word9[17]), .A1(fifo_out[46]), .Z(n201));
Q_AN02 U541 ( .A0(tlv_word9[17]), .A1(fifo_out[45]), .Z(n202));
Q_AN02 U542 ( .A0(tlv_word9[17]), .A1(fifo_out[44]), .Z(n203));
Q_AN02 U543 ( .A0(tlv_word9[17]), .A1(fifo_out[43]), .Z(n204));
Q_AN02 U544 ( .A0(tlv_word9[17]), .A1(fifo_out[42]), .Z(n205));
Q_AN02 U545 ( .A0(tlv_word9[17]), .A1(fifo_out[41]), .Z(n206));
Q_AN02 U546 ( .A0(tlv_word9[17]), .A1(fifo_out[40]), .Z(n207));
Q_AN02 U547 ( .A0(tlv_word9[17]), .A1(fifo_out[39]), .Z(n208));
Q_AN02 U548 ( .A0(tlv_word9[17]), .A1(fifo_out[38]), .Z(n209));
Q_AN02 U549 ( .A0(tlv_word9[17]), .A1(fifo_out[37]), .Z(n210));
Q_AN02 U550 ( .A0(tlv_word9[17]), .A1(fifo_out[36]), .Z(n211));
Q_AN02 U551 ( .A0(tlv_word9[17]), .A1(fifo_out[35]), .Z(n212));
Q_AN02 U552 ( .A0(tlv_word9[17]), .A1(fifo_out[34]), .Z(n213));
Q_AN02 U553 ( .A0(tlv_word9[17]), .A1(fifo_out[33]), .Z(n214));
Q_AN02 U554 ( .A0(tlv_word9[17]), .A1(fifo_out[32]), .Z(n215));
Q_AN02 U555 ( .A0(tlv_word9[17]), .A1(fifo_out[31]), .Z(n216));
Q_AN02 U556 ( .A0(tlv_word9[17]), .A1(fifo_out[30]), .Z(n217));
Q_AN02 U557 ( .A0(tlv_word9[17]), .A1(fifo_out[29]), .Z(n218));
Q_AN02 U558 ( .A0(tlv_word9[17]), .A1(fifo_out[28]), .Z(n219));
Q_AN02 U559 ( .A0(tlv_word9[17]), .A1(fifo_out[27]), .Z(n220));
Q_AN02 U560 ( .A0(tlv_word9[17]), .A1(fifo_out[26]), .Z(n221));
Q_AN02 U561 ( .A0(tlv_word9[17]), .A1(fifo_out[25]), .Z(n222));
Q_AN02 U562 ( .A0(tlv_word9[17]), .A1(fifo_out[24]), .Z(n223));
Q_AN02 U563 ( .A0(tlv_word9[17]), .A1(fifo_out[23]), .Z(n224));
Q_AN02 U564 ( .A0(tlv_word9[17]), .A1(fifo_out[22]), .Z(n225));
Q_AN02 U565 ( .A0(tlv_word9[17]), .A1(fifo_out[21]), .Z(n226));
Q_AN02 U566 ( .A0(tlv_word9[17]), .A1(fifo_out[20]), .Z(n227));
Q_AN02 U567 ( .A0(tlv_word9[17]), .A1(fifo_out[19]), .Z(n228));
Q_AN02 U568 ( .A0(tlv_word9[17]), .A1(fifo_out[18]), .Z(n229));
Q_AN02 U569 ( .A0(tlv_word9[17]), .A1(fifo_out[17]), .Z(n230));
Q_AN02 U570 ( .A0(tlv_word9[17]), .A1(fifo_out[16]), .Z(n231));
Q_AN02 U571 ( .A0(tlv_word9[17]), .A1(fifo_out[15]), .Z(n232));
Q_AN02 U572 ( .A0(tlv_word9[17]), .A1(fifo_out[14]), .Z(n233));
Q_AN02 U573 ( .A0(tlv_word9[17]), .A1(fifo_out[13]), .Z(n234));
Q_AN02 U574 ( .A0(tlv_word9[17]), .A1(fifo_out[12]), .Z(n235));
Q_AN02 U575 ( .A0(tlv_word9[17]), .A1(fifo_out[11]), .Z(n236));
Q_AN02 U576 ( .A0(tlv_word9[17]), .A1(fifo_out[10]), .Z(n237));
Q_AN02 U577 ( .A0(tlv_word9[17]), .A1(fifo_out[9]), .Z(n238));
Q_AN02 U578 ( .A0(tlv_word9[17]), .A1(fifo_out[8]), .Z(n239));
Q_AN02 U579 ( .A0(tlv_word9[17]), .A1(fifo_out[7]), .Z(n240));
Q_AN02 U580 ( .A0(tlv_word9[17]), .A1(fifo_out[6]), .Z(n241));
Q_AN02 U581 ( .A0(tlv_word9[17]), .A1(fifo_out[5]), .Z(n242));
Q_AN02 U582 ( .A0(tlv_word9[17]), .A1(fifo_out[4]), .Z(n243));
Q_AN02 U583 ( .A0(tlv_word9[17]), .A1(fifo_out[3]), .Z(n244));
Q_AN02 U584 ( .A0(tlv_word9[17]), .A1(fifo_out[2]), .Z(n245));
Q_AN02 U585 ( .A0(tlv_word9[17]), .A1(fifo_out[1]), .Z(n246));
Q_AN02 U586 ( .A0(tlv_word9[17]), .A1(fifo_out[0]), .Z(n247));
Q_AN02 U587 ( .A0(tlv_word8[17]), .A1(fifo_out[63]), .Z(n248));
Q_AN02 U588 ( .A0(tlv_word8[17]), .A1(fifo_out[62]), .Z(n249));
Q_AN02 U589 ( .A0(tlv_word8[17]), .A1(fifo_out[61]), .Z(n250));
Q_AN02 U590 ( .A0(tlv_word8[17]), .A1(fifo_out[60]), .Z(n251));
Q_AN02 U591 ( .A0(tlv_word8[17]), .A1(fifo_out[59]), .Z(n252));
Q_AN02 U592 ( .A0(tlv_word8[17]), .A1(fifo_out[58]), .Z(n253));
Q_AN02 U593 ( .A0(tlv_word8[17]), .A1(fifo_out[57]), .Z(n254));
Q_AN02 U594 ( .A0(tlv_word8[17]), .A1(fifo_out[56]), .Z(n255));
Q_AN02 U595 ( .A0(tlv_word8[17]), .A1(fifo_out[55]), .Z(n256));
Q_AN02 U596 ( .A0(tlv_word8[17]), .A1(fifo_out[54]), .Z(n257));
Q_AN02 U597 ( .A0(tlv_word8[17]), .A1(fifo_out[53]), .Z(n258));
Q_AN02 U598 ( .A0(tlv_word8[17]), .A1(fifo_out[52]), .Z(n259));
Q_AN02 U599 ( .A0(tlv_word8[17]), .A1(fifo_out[51]), .Z(n260));
Q_AN02 U600 ( .A0(tlv_word8[17]), .A1(fifo_out[50]), .Z(n261));
Q_AN02 U601 ( .A0(tlv_word8[17]), .A1(fifo_out[49]), .Z(n262));
Q_AN02 U602 ( .A0(tlv_word8[17]), .A1(fifo_out[48]), .Z(n263));
Q_AN02 U603 ( .A0(tlv_word8[17]), .A1(fifo_out[47]), .Z(n264));
Q_AN02 U604 ( .A0(tlv_word8[17]), .A1(fifo_out[46]), .Z(n265));
Q_AN02 U605 ( .A0(tlv_word8[17]), .A1(fifo_out[45]), .Z(n266));
Q_AN02 U606 ( .A0(tlv_word8[17]), .A1(fifo_out[44]), .Z(n267));
Q_AN02 U607 ( .A0(tlv_word8[17]), .A1(fifo_out[43]), .Z(n268));
Q_AN02 U608 ( .A0(tlv_word8[17]), .A1(fifo_out[42]), .Z(n269));
Q_AN02 U609 ( .A0(tlv_word8[17]), .A1(fifo_out[41]), .Z(n270));
Q_AN02 U610 ( .A0(tlv_word8[17]), .A1(fifo_out[40]), .Z(n271));
Q_AN02 U611 ( .A0(tlv_word8[17]), .A1(fifo_out[39]), .Z(n272));
Q_AN02 U612 ( .A0(tlv_word8[17]), .A1(fifo_out[38]), .Z(n273));
Q_AN02 U613 ( .A0(tlv_word8[17]), .A1(fifo_out[37]), .Z(n274));
Q_AN02 U614 ( .A0(tlv_word8[17]), .A1(fifo_out[36]), .Z(n275));
Q_AN02 U615 ( .A0(tlv_word8[17]), .A1(fifo_out[35]), .Z(n276));
Q_AN02 U616 ( .A0(tlv_word8[17]), .A1(fifo_out[34]), .Z(n277));
Q_AN02 U617 ( .A0(tlv_word8[17]), .A1(fifo_out[33]), .Z(n278));
Q_AN02 U618 ( .A0(tlv_word8[17]), .A1(fifo_out[32]), .Z(n279));
Q_AN02 U619 ( .A0(tlv_word8[17]), .A1(fifo_out[31]), .Z(n280));
Q_AN02 U620 ( .A0(tlv_word8[17]), .A1(fifo_out[30]), .Z(n281));
Q_AN02 U621 ( .A0(tlv_word8[17]), .A1(fifo_out[29]), .Z(n282));
Q_AN02 U622 ( .A0(tlv_word8[17]), .A1(fifo_out[28]), .Z(n283));
Q_AN02 U623 ( .A0(tlv_word8[17]), .A1(fifo_out[27]), .Z(n284));
Q_AN02 U624 ( .A0(tlv_word8[17]), .A1(fifo_out[26]), .Z(n285));
Q_AN02 U625 ( .A0(tlv_word8[17]), .A1(fifo_out[25]), .Z(n286));
Q_AN02 U626 ( .A0(tlv_word8[17]), .A1(fifo_out[24]), .Z(n287));
Q_AN02 U627 ( .A0(tlv_word8[17]), .A1(fifo_out[23]), .Z(n288));
Q_AN02 U628 ( .A0(tlv_word8[17]), .A1(fifo_out[22]), .Z(n289));
Q_AN02 U629 ( .A0(tlv_word8[17]), .A1(fifo_out[21]), .Z(n290));
Q_AN02 U630 ( .A0(tlv_word8[17]), .A1(fifo_out[20]), .Z(n291));
Q_AN02 U631 ( .A0(tlv_word8[17]), .A1(fifo_out[19]), .Z(n292));
Q_AN02 U632 ( .A0(tlv_word8[17]), .A1(fifo_out[18]), .Z(n293));
Q_AN02 U633 ( .A0(tlv_word8[17]), .A1(fifo_out[17]), .Z(n294));
Q_AN02 U634 ( .A0(tlv_word8[17]), .A1(fifo_out[16]), .Z(n295));
Q_AN02 U635 ( .A0(tlv_word8[17]), .A1(fifo_out[15]), .Z(n296));
Q_AN02 U636 ( .A0(tlv_word8[17]), .A1(fifo_out[14]), .Z(n297));
Q_AN02 U637 ( .A0(tlv_word8[17]), .A1(fifo_out[13]), .Z(n298));
Q_AN02 U638 ( .A0(tlv_word8[17]), .A1(fifo_out[12]), .Z(n299));
Q_AN02 U639 ( .A0(tlv_word8[17]), .A1(fifo_out[11]), .Z(n300));
Q_AN02 U640 ( .A0(tlv_word8[17]), .A1(fifo_out[10]), .Z(n301));
Q_AN02 U641 ( .A0(tlv_word8[17]), .A1(fifo_out[9]), .Z(n302));
Q_AN02 U642 ( .A0(tlv_word8[17]), .A1(fifo_out[8]), .Z(n303));
Q_AN02 U643 ( .A0(tlv_word8[17]), .A1(fifo_out[7]), .Z(n304));
Q_AN02 U644 ( .A0(tlv_word8[17]), .A1(fifo_out[6]), .Z(n305));
Q_AN02 U645 ( .A0(tlv_word8[17]), .A1(fifo_out[5]), .Z(n306));
Q_AN02 U646 ( .A0(tlv_word8[17]), .A1(fifo_out[4]), .Z(n307));
Q_AN02 U647 ( .A0(tlv_word8[17]), .A1(fifo_out[3]), .Z(n308));
Q_AN02 U648 ( .A0(tlv_word8[17]), .A1(fifo_out[2]), .Z(n309));
Q_AN02 U649 ( .A0(tlv_word8[17]), .A1(fifo_out[1]), .Z(n310));
Q_AN02 U650 ( .A0(tlv_word8[17]), .A1(fifo_out[0]), .Z(n311));
Q_OR02 U651 ( .A0(report_kme_error), .A1(kimreader_ckvreader_data[7]), .Z(tlv_word42[7]));
Q_AN02 U652 ( .A0(n14), .A1(kimreader_ckvreader_data[6]), .Z(tlv_word42[6]));
Q_AN02 U653 ( .A0(n14), .A1(kimreader_ckvreader_data[5]), .Z(tlv_word42[5]));
Q_AN02 U654 ( .A0(n14), .A1(kimreader_ckvreader_data[4]), .Z(tlv_word42[4]));
Q_OR02 U655 ( .A0(report_kme_error), .A1(kimreader_ckvreader_data[3]), .Z(tlv_word42[3]));
Q_AN02 U656 ( .A0(n14), .A1(kimreader_ckvreader_data[2]), .Z(tlv_word42[2]));
Q_AN02 U657 ( .A0(n14), .A1(kimreader_ckvreader_data[1]), .Z(tlv_word42[1]));
Q_OR02 U658 ( .A0(report_kme_error), .A1(kimreader_ckvreader_data[0]), .Z(tlv_word42[0]));
Q_AN02 U659 ( .A0(tlv_word8[58]), .A1(n412), .Z(half_dek));
Q_NR02 U660 ( .A0(n314), .A1(n313), .Z(n312));
Q_OR03 U661 ( .A0(kimreader_ckvreader_data[41]), .A1(kimreader_ckvreader_data[40]), .A2(n315), .Z(n313));
Q_OR03 U662 ( .A0(kimreader_ckvreader_data[44]), .A1(kimreader_ckvreader_data[43]), .A2(kimreader_ckvreader_data[42]), .Z(n314));
Q_INV U663 ( .A(kimreader_ckvreader_data[39]), .Z(n315));
Q_AN02 U664 ( .A0(n386), .A1(kimreader_ckvreader_data[69]), .Z(n7));
Q_NR02 U665 ( .A0(n387), .A1(kimreader_ckvreader_data[69]), .Z(n8));
Q_INV U666 ( .A(n316), .Z(n6));
Q_OR02 U667 ( .A0(kimreader_ckvreader_data[64]), .A1(n317), .Z(n316));
Q_OR03 U668 ( .A0(kimreader_ckvreader_data[67]), .A1(kimreader_ckvreader_data[66]), .A2(kimreader_ckvreader_data[65]), .Z(n317));
Q_OR02 U669 ( .A0(n382), .A1(ckv_rd), .Z(n318));
Q_AN02 U670 ( .A0(ckv_read_num[1]), .A1(half_dek), .Z(n323));
Q_INV U671 ( .A(n323), .Z(n321));
Q_OR03 U672 ( .A0(ckv_read_num[3]), .A1(ckv_read_num[2]), .A2(n321), .Z(n322));
Q_OA21 U673 ( .A0(n351), .A1(n322), .B0(cur_state[0]), .Z(n319));
Q_MX02 U674 ( .S(ckv_read_num[2]), .A0(n323), .A1(ckv_read_num[1]), .Z(n324));
Q_INV U675 ( .A(n324), .Z(n326));
Q_OR02 U676 ( .A0(n351), .A1(ckv_read_num[3]), .Z(n325));
Q_OR03 U677 ( .A0(n382), .A1(n325), .A2(n326), .Z(n320));
Q_MX04 U678 ( .S0(n320), .S1(n319), .A0(tlv_word8[57]), .A1(nxt_tlv_word8[57]), .A2(tlv_word9[57]), .A3(n352), .Z(n327));
Q_MX04 U679 ( .S0(n320), .S1(n319), .A0(tlv_word8[56]), .A1(nxt_tlv_word8[56]), .A2(tlv_word9[56]), .A3(n354), .Z(n328));
Q_MX04 U680 ( .S0(n320), .S1(n319), .A0(tlv_word8[55]), .A1(nxt_tlv_word8[55]), .A2(tlv_word9[55]), .A3(n356), .Z(n329));
Q_MX04 U681 ( .S0(n320), .S1(n319), .A0(tlv_word8[54]), .A1(nxt_tlv_word8[54]), .A2(tlv_word9[54]), .A3(n358), .Z(n330));
Q_MX04 U682 ( .S0(n320), .S1(n319), .A0(tlv_word8[53]), .A1(nxt_tlv_word8[53]), .A2(tlv_word9[53]), .A3(n360), .Z(n331));
Q_MX04 U683 ( .S0(n320), .S1(n319), .A0(tlv_word8[52]), .A1(nxt_tlv_word8[52]), .A2(tlv_word9[52]), .A3(n362), .Z(n332));
Q_MX04 U684 ( .S0(n320), .S1(n319), .A0(tlv_word8[51]), .A1(nxt_tlv_word8[51]), .A2(tlv_word9[51]), .A3(n364), .Z(n333));
Q_MX04 U685 ( .S0(n320), .S1(n319), .A0(tlv_word8[50]), .A1(nxt_tlv_word8[50]), .A2(tlv_word9[50]), .A3(n366), .Z(n334));
Q_MX04 U686 ( .S0(n320), .S1(n319), .A0(tlv_word8[49]), .A1(nxt_tlv_word8[49]), .A2(tlv_word9[49]), .A3(n368), .Z(n335));
Q_MX04 U687 ( .S0(n320), .S1(n319), .A0(tlv_word8[48]), .A1(nxt_tlv_word8[48]), .A2(tlv_word9[48]), .A3(n370), .Z(n336));
Q_MX04 U688 ( .S0(n320), .S1(n319), .A0(tlv_word8[47]), .A1(nxt_tlv_word8[47]), .A2(tlv_word9[47]), .A3(n372), .Z(n337));
Q_MX04 U689 ( .S0(n320), .S1(n319), .A0(tlv_word8[46]), .A1(nxt_tlv_word8[46]), .A2(tlv_word9[46]), .A3(n374), .Z(n338));
Q_MX04 U690 ( .S0(n320), .S1(n319), .A0(tlv_word8[45]), .A1(nxt_tlv_word8[45]), .A2(tlv_word9[45]), .A3(n376), .Z(n339));
Q_MX04 U691 ( .S0(n320), .S1(n319), .A0(tlv_word8[44]), .A1(nxt_tlv_word8[44]), .A2(tlv_word9[44]), .A3(n378), .Z(n340));
Q_MX04 U692 ( .S0(n320), .S1(n319), .A0(tlv_word8[43]), .A1(nxt_tlv_word8[43]), .A2(tlv_word9[43]), .A3(n379), .Z(n341));
Q_AN02 U693 ( .A0(cur_state[0]), .A1(n346), .Z(n342));
Q_AN02 U694 ( .A0(cur_state[0]), .A1(n348), .Z(n343));
Q_AN02 U695 ( .A0(cur_state[0]), .A1(n350), .Z(n344));
Q_AN02 U696 ( .A0(cur_state[0]), .A1(n351), .Z(n345));
Q_XOR2 U697 ( .A0(ckv_read_num[3]), .A1(n347), .Z(n346));
Q_AD01HF U698 ( .A0(ckv_read_num[2]), .B0(n349), .S(n348), .CO(n347));
Q_AD01HF U699 ( .A0(ckv_read_num[1]), .B0(ckv_read_num[0]), .S(n350), .CO(n349));
Q_XOR2 U700 ( .A0(ckv_addr[14]), .A1(n353), .Z(n352));
Q_AD01HF U701 ( .A0(ckv_addr[13]), .B0(n355), .S(n354), .CO(n353));
Q_AD01HF U702 ( .A0(ckv_addr[12]), .B0(n357), .S(n356), .CO(n355));
Q_AD01HF U703 ( .A0(ckv_addr[11]), .B0(n359), .S(n358), .CO(n357));
Q_AD01HF U704 ( .A0(ckv_addr[10]), .B0(n361), .S(n360), .CO(n359));
Q_AD01HF U705 ( .A0(ckv_addr[9]), .B0(n363), .S(n362), .CO(n361));
Q_AD01HF U706 ( .A0(ckv_addr[8]), .B0(n365), .S(n364), .CO(n363));
Q_AD01HF U707 ( .A0(ckv_addr[7]), .B0(n367), .S(n366), .CO(n365));
Q_AD01HF U708 ( .A0(ckv_addr[6]), .B0(n369), .S(n368), .CO(n367));
Q_AD01HF U709 ( .A0(ckv_addr[5]), .B0(n371), .S(n370), .CO(n369));
Q_AD01HF U710 ( .A0(ckv_addr[4]), .B0(n373), .S(n372), .CO(n371));
Q_AD01HF U711 ( .A0(ckv_addr[3]), .B0(n375), .S(n374), .CO(n373));
Q_AD01HF U712 ( .A0(ckv_addr[2]), .B0(n377), .S(n376), .CO(n375));
Q_AD01HF U713 ( .A0(ckv_addr[1]), .B0(ckv_addr[0]), .S(n378), .CO(n377));
Q_MX02 U714 ( .S(cur_state[0]), .A0(n381), .A1(n380), .Z(nxt_state[0]));
Q_ND03 U715 ( .A0(kopassigner_ckvreader_ack), .A1(n383), .A2(kimreader_ckvreader_data[69]), .Z(n380));
Q_AN02 U716 ( .A0(kimreader_ckvreader_data[64]), .A1(n384), .Z(n383));
Q_AN03 U717 ( .A0(n385), .A1(kimreader_ckvreader_data[66]), .A2(kimreader_ckvreader_data[65]), .Z(n384));
Q_INV U718 ( .A(kimreader_ckvreader_data[67]), .Z(n385));
Q_AN03 U719 ( .A0(kopassigner_ckvreader_ack), .A1(n386), .A2(kimreader_ckvreader_data[69]), .Z(n381));
Q_INV U720 ( .A(n387), .Z(n386));
Q_OR02 U721 ( .A0(kimreader_ckvreader_data[64]), .A1(n388), .Z(n387));
Q_OR03 U722 ( .A0(kimreader_ckvreader_data[67]), .A1(n389), .A2(kimreader_ckvreader_data[65]), .Z(n388));
Q_INV U723 ( .A(kimreader_ckvreader_data[66]), .Z(n389));
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN(n382));
Q_FDP1 ckv_rd_q_REG  ( .CK(clk), .R(rst_n), .D(ckv_rd), .Q(ckv_rd_q), .QN( ));
Q_FDP1 \tlv_word8_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[63]), .Q(tlv_word8[63]), .QN( ));
Q_FDP1 \tlv_word8_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[62]), .Q(tlv_word8[62]), .QN( ));
Q_FDP1 \tlv_word8_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[61]), .Q(tlv_word8[61]), .QN( ));
Q_FDP1 \tlv_word8_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[60]), .Q(tlv_word8[60]), .QN( ));
Q_FDP1 \tlv_word8_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[59]), .Q(tlv_word8[59]), .QN(n412));
Q_FDP1 \tlv_word8_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[58]), .Q(tlv_word8[58]), .QN(n407));
Q_FDP1 \tlv_word8_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[57]), .Q(tlv_word8[57]), .QN( ));
Q_FDP1 \tlv_word8_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[56]), .Q(tlv_word8[56]), .QN( ));
Q_FDP1 \tlv_word8_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[55]), .Q(tlv_word8[55]), .QN( ));
Q_FDP1 \tlv_word8_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[54]), .Q(tlv_word8[54]), .QN( ));
Q_FDP1 \tlv_word8_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[53]), .Q(tlv_word8[53]), .QN( ));
Q_FDP1 \tlv_word8_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[52]), .Q(tlv_word8[52]), .QN( ));
Q_FDP1 \tlv_word8_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[51]), .Q(tlv_word8[51]), .QN( ));
Q_FDP1 \tlv_word8_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[50]), .Q(tlv_word8[50]), .QN( ));
Q_FDP1 \tlv_word8_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[49]), .Q(tlv_word8[49]), .QN( ));
Q_FDP1 \tlv_word8_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[48]), .Q(tlv_word8[48]), .QN( ));
Q_FDP1 \tlv_word8_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[47]), .Q(tlv_word8[47]), .QN( ));
Q_FDP1 \tlv_word8_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[46]), .Q(tlv_word8[46]), .QN( ));
Q_FDP1 \tlv_word8_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[45]), .Q(tlv_word8[45]), .QN( ));
Q_FDP1 \tlv_word8_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[44]), .Q(tlv_word8[44]), .QN( ));
Q_FDP1 \tlv_word8_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[43]), .Q(tlv_word8[43]), .QN( ));
Q_FDP1 \tlv_word8_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[42]), .Q(tlv_word8[42]), .QN( ));
Q_FDP1 \tlv_word8_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[41]), .Q(tlv_word8[41]), .QN( ));
Q_FDP1 \tlv_word8_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[40]), .Q(tlv_word8[40]), .QN( ));
Q_FDP1 \tlv_word8_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[39]), .Q(tlv_word8[39]), .QN( ));
Q_FDP1 \tlv_word8_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[38]), .Q(tlv_word8[38]), .QN( ));
Q_FDP1 \tlv_word8_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[37]), .Q(tlv_word8[37]), .QN( ));
Q_FDP1 \tlv_word8_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[36]), .Q(tlv_word8[36]), .QN( ));
Q_FDP1 \tlv_word8_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[35]), .Q(tlv_word8[35]), .QN( ));
Q_FDP1 \tlv_word8_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[34]), .Q(tlv_word8[34]), .QN( ));
Q_FDP1 \tlv_word8_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[33]), .Q(tlv_word8[33]), .QN( ));
Q_FDP1 \tlv_word8_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[32]), .Q(tlv_word8[32]), .QN( ));
Q_FDP1 \tlv_word8_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[31]), .Q(tlv_word8[31]), .QN( ));
Q_FDP1 \tlv_word8_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[30]), .Q(tlv_word8[30]), .QN( ));
Q_FDP1 \tlv_word8_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[29]), .Q(tlv_word8[29]), .QN( ));
Q_FDP1 \tlv_word8_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[28]), .Q(tlv_word8[28]), .QN( ));
Q_FDP1 \tlv_word8_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[27]), .Q(tlv_word8[27]), .QN( ));
Q_FDP1 \tlv_word8_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[26]), .Q(tlv_word8[26]), .QN( ));
Q_FDP1 \tlv_word8_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[25]), .Q(tlv_word8[25]), .QN( ));
Q_FDP1 \tlv_word8_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[24]), .Q(tlv_word8[24]), .QN( ));
Q_FDP1 \tlv_word8_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[23]), .Q(tlv_word8[23]), .QN( ));
Q_FDP1 \tlv_word8_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[22]), .Q(tlv_word8[22]), .QN( ));
Q_FDP1 \tlv_word8_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[21]), .Q(tlv_word8[21]), .QN( ));
Q_FDP1 \tlv_word8_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[20]), .Q(tlv_word8[20]), .QN( ));
Q_FDP1 \tlv_word8_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[19]), .Q(tlv_word8[19]), .QN( ));
Q_FDP1 \tlv_word8_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[18]), .Q(tlv_word8[18]), .QN( ));
Q_FDP1 \tlv_word8_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[17]), .Q(tlv_word8[17]), .QN( ));
Q_FDP1 \tlv_word8_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[16]), .Q(tlv_word8[16]), .QN( ));
Q_FDP1 \tlv_word8_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[15]), .Q(tlv_word8[15]), .QN( ));
Q_FDP1 \tlv_word8_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[14]), .Q(tlv_word8[14]), .QN( ));
Q_FDP1 \tlv_word8_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[13]), .Q(tlv_word8[13]), .QN( ));
Q_FDP1 \tlv_word8_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[12]), .Q(tlv_word8[12]), .QN( ));
Q_FDP1 \tlv_word8_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[11]), .Q(tlv_word8[11]), .QN( ));
Q_FDP1 \tlv_word8_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[10]), .Q(tlv_word8[10]), .QN( ));
Q_FDP1 \tlv_word8_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[9]), .Q(tlv_word8[9]), .QN( ));
Q_FDP1 \tlv_word8_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[8]), .Q(tlv_word8[8]), .QN( ));
Q_FDP1 \tlv_word8_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[7]), .Q(tlv_word8[7]), .QN( ));
Q_FDP1 \tlv_word8_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[6]), .Q(tlv_word8[6]), .QN( ));
Q_FDP1 \tlv_word8_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[5]), .Q(tlv_word8[5]), .QN( ));
Q_FDP1 \tlv_word8_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[4]), .Q(tlv_word8[4]), .QN( ));
Q_FDP1 \tlv_word8_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[3]), .Q(tlv_word8[3]), .QN( ));
Q_FDP1 \tlv_word8_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[2]), .Q(tlv_word8[2]), .QN( ));
Q_FDP1 \tlv_word8_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[1]), .Q(tlv_word8[1]), .QN( ));
Q_FDP1 \tlv_word8_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word8[0]), .Q(tlv_word8[0]), .QN( ));
Q_FDP1 \tlv_word9_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[63]), .Q(tlv_word9[63]), .QN( ));
Q_FDP1 \tlv_word9_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[62]), .Q(tlv_word9[62]), .QN( ));
Q_FDP1 \tlv_word9_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[61]), .Q(tlv_word9[61]), .QN( ));
Q_FDP1 \tlv_word9_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[60]), .Q(tlv_word9[60]), .QN( ));
Q_FDP1 \tlv_word9_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[59]), .Q(tlv_word9[59]), .QN(n410));
Q_FDP1 \tlv_word9_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[58]), .Q(tlv_word9[58]), .QN(n404));
Q_FDP1 \tlv_word9_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[57]), .Q(tlv_word9[57]), .QN( ));
Q_FDP1 \tlv_word9_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[56]), .Q(tlv_word9[56]), .QN( ));
Q_FDP1 \tlv_word9_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[55]), .Q(tlv_word9[55]), .QN( ));
Q_FDP1 \tlv_word9_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[54]), .Q(tlv_word9[54]), .QN( ));
Q_FDP1 \tlv_word9_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[53]), .Q(tlv_word9[53]), .QN( ));
Q_FDP1 \tlv_word9_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[52]), .Q(tlv_word9[52]), .QN( ));
Q_FDP1 \tlv_word9_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[51]), .Q(tlv_word9[51]), .QN( ));
Q_FDP1 \tlv_word9_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[50]), .Q(tlv_word9[50]), .QN( ));
Q_FDP1 \tlv_word9_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[49]), .Q(tlv_word9[49]), .QN( ));
Q_FDP1 \tlv_word9_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[48]), .Q(tlv_word9[48]), .QN( ));
Q_FDP1 \tlv_word9_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[47]), .Q(tlv_word9[47]), .QN( ));
Q_FDP1 \tlv_word9_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[46]), .Q(tlv_word9[46]), .QN( ));
Q_FDP1 \tlv_word9_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[45]), .Q(tlv_word9[45]), .QN( ));
Q_FDP1 \tlv_word9_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[44]), .Q(tlv_word9[44]), .QN( ));
Q_FDP1 \tlv_word9_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[43]), .Q(tlv_word9[43]), .QN( ));
Q_FDP1 \tlv_word9_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[42]), .Q(tlv_word9[42]), .QN( ));
Q_FDP1 \tlv_word9_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[41]), .Q(tlv_word9[41]), .QN( ));
Q_FDP1 \tlv_word9_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[40]), .Q(tlv_word9[40]), .QN( ));
Q_FDP1 \tlv_word9_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[39]), .Q(tlv_word9[39]), .QN( ));
Q_FDP1 \tlv_word9_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[38]), .Q(tlv_word9[38]), .QN( ));
Q_FDP1 \tlv_word9_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[37]), .Q(tlv_word9[37]), .QN( ));
Q_FDP1 \tlv_word9_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[36]), .Q(tlv_word9[36]), .QN( ));
Q_FDP1 \tlv_word9_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[35]), .Q(tlv_word9[35]), .QN( ));
Q_FDP1 \tlv_word9_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[34]), .Q(tlv_word9[34]), .QN( ));
Q_FDP1 \tlv_word9_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[33]), .Q(tlv_word9[33]), .QN( ));
Q_FDP1 \tlv_word9_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[32]), .Q(tlv_word9[32]), .QN( ));
Q_FDP1 \tlv_word9_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[31]), .Q(tlv_word9[31]), .QN( ));
Q_FDP1 \tlv_word9_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[30]), .Q(tlv_word9[30]), .QN( ));
Q_FDP1 \tlv_word9_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[29]), .Q(tlv_word9[29]), .QN( ));
Q_FDP1 \tlv_word9_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[28]), .Q(tlv_word9[28]), .QN( ));
Q_FDP1 \tlv_word9_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[27]), .Q(tlv_word9[27]), .QN( ));
Q_FDP1 \tlv_word9_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[26]), .Q(tlv_word9[26]), .QN( ));
Q_FDP1 \tlv_word9_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[25]), .Q(tlv_word9[25]), .QN( ));
Q_FDP1 \tlv_word9_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[24]), .Q(tlv_word9[24]), .QN( ));
Q_FDP1 \tlv_word9_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[23]), .Q(tlv_word9[23]), .QN( ));
Q_FDP1 \tlv_word9_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[22]), .Q(tlv_word9[22]), .QN( ));
Q_FDP1 \tlv_word9_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[21]), .Q(tlv_word9[21]), .QN( ));
Q_FDP1 \tlv_word9_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[20]), .Q(tlv_word9[20]), .QN( ));
Q_FDP1 \tlv_word9_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[19]), .Q(tlv_word9[19]), .QN( ));
Q_FDP1 \tlv_word9_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[18]), .Q(tlv_word9[18]), .QN( ));
Q_FDP1 \tlv_word9_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[17]), .Q(tlv_word9[17]), .QN( ));
Q_FDP1 \tlv_word9_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[16]), .Q(tlv_word9[16]), .QN( ));
Q_FDP1 \tlv_word9_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[15]), .Q(tlv_word9[15]), .QN( ));
Q_FDP1 \tlv_word9_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[14]), .Q(tlv_word9[14]), .QN( ));
Q_FDP1 \tlv_word9_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[13]), .Q(tlv_word9[13]), .QN( ));
Q_FDP1 \tlv_word9_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[12]), .Q(tlv_word9[12]), .QN( ));
Q_FDP1 \tlv_word9_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[11]), .Q(tlv_word9[11]), .QN( ));
Q_FDP1 \tlv_word9_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[10]), .Q(tlv_word9[10]), .QN( ));
Q_FDP1 \tlv_word9_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[9]), .Q(tlv_word9[9]), .QN( ));
Q_FDP1 \tlv_word9_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[8]), .Q(tlv_word9[8]), .QN( ));
Q_FDP1 \tlv_word9_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[7]), .Q(tlv_word9[7]), .QN( ));
Q_FDP1 \tlv_word9_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[6]), .Q(tlv_word9[6]), .QN( ));
Q_FDP1 \tlv_word9_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[5]), .Q(tlv_word9[5]), .QN( ));
Q_FDP1 \tlv_word9_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[4]), .Q(tlv_word9[4]), .QN( ));
Q_FDP1 \tlv_word9_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[3]), .Q(tlv_word9[3]), .QN( ));
Q_FDP1 \tlv_word9_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[2]), .Q(tlv_word9[2]), .QN( ));
Q_FDP1 \tlv_word9_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[1]), .Q(tlv_word9[1]), .QN( ));
Q_FDP1 \tlv_word9_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_tlv_word9[0]), .Q(tlv_word9[0]), .QN( ));
Q_FDP1 ktype_is_aux_key_only_REG  ( .CK(clk), .R(rst_n), .D(nxt_ktype_is_aux_key_only), .Q(ktype_is_aux_key_only), .QN( ));
Q_AN02 U855 ( .A0(rst_n), .A1(_zy_sva_b7), .Z(n390));
Q_AN02 U856 ( .A0(rst_n), .A1(_zy_sva_b6), .Z(n391));
Q_AN02 U857 ( .A0(rst_n), .A1(_zy_sva_b5), .Z(n392));
Q_AN02 U858 ( .A0(rst_n), .A1(_zy_sva_b4), .Z(n393));
Q_AN02 U859 ( .A0(rst_n), .A1(_zy_sva_b3), .Z(n394));
Q_AN02 U860 ( .A0(rst_n), .A1(_zy_sva_b2), .Z(n395));
Q_AN02 U861 ( .A0(rst_n), .A1(_zy_sva_b1), .Z(n396));
Q_AN02 U862 ( .A0(rst_n), .A1(_zy_sva_b0), .Z(n397));
ixc_assign _zz_strnp_0 ( _zy_simnet_ckvreader_kimreader_ack_0_w$, 
	kopassigner_ckvreader_ack);
ixc_assign _zz_strnp_1 ( _zy_simnet_ckvreader_kopassigner_valid_1_w$, 
	ckvreader_kopassigner_valid);
ixc_assign_71 _zz_strnp_2 ( _zy_simnet_ckvreader_kopassigner_data_2_w$[0:70], { 
	kimreader_ckvreader_data[70], kimreader_ckvreader_data[69], 
	kimreader_ckvreader_data[68], kimreader_ckvreader_data[67], 
	kimreader_ckvreader_data[66], kimreader_ckvreader_data[65], 
	kimreader_ckvreader_data[64], ckvreader_kopassigner_data[63], 
	ckvreader_kopassigner_data[62], ckvreader_kopassigner_data[61], 
	ckvreader_kopassigner_data[60], ckvreader_kopassigner_data[59], 
	ckvreader_kopassigner_data[58], ckvreader_kopassigner_data[57], 
	ckvreader_kopassigner_data[56], ckvreader_kopassigner_data[55], 
	ckvreader_kopassigner_data[54], ckvreader_kopassigner_data[53], 
	ckvreader_kopassigner_data[52], ckvreader_kopassigner_data[51], 
	ckvreader_kopassigner_data[50], ckvreader_kopassigner_data[49], 
	ckvreader_kopassigner_data[48], ckvreader_kopassigner_data[47], 
	ckvreader_kopassigner_data[46], ckvreader_kopassigner_data[45], 
	ckvreader_kopassigner_data[44], ckvreader_kopassigner_data[43], 
	ckvreader_kopassigner_data[42], ckvreader_kopassigner_data[41], 
	ckvreader_kopassigner_data[40], ckvreader_kopassigner_data[39], 
	ckvreader_kopassigner_data[38], ckvreader_kopassigner_data[37], 
	ckvreader_kopassigner_data[36], ckvreader_kopassigner_data[35], 
	ckvreader_kopassigner_data[34], ckvreader_kopassigner_data[33], 
	ckvreader_kopassigner_data[32], ckvreader_kopassigner_data[31], 
	ckvreader_kopassigner_data[30], ckvreader_kopassigner_data[29], 
	ckvreader_kopassigner_data[28], ckvreader_kopassigner_data[27], 
	ckvreader_kopassigner_data[26], ckvreader_kopassigner_data[25], 
	ckvreader_kopassigner_data[24], ckvreader_kopassigner_data[23], 
	ckvreader_kopassigner_data[22], ckvreader_kopassigner_data[21], 
	ckvreader_kopassigner_data[20], ckvreader_kopassigner_data[19], 
	ckvreader_kopassigner_data[18], ckvreader_kopassigner_data[17], 
	ckvreader_kopassigner_data[16], ckvreader_kopassigner_data[15], 
	ckvreader_kopassigner_data[14], ckvreader_kopassigner_data[13], 
	ckvreader_kopassigner_data[12], ckvreader_kopassigner_data[11], 
	ckvreader_kopassigner_data[10], ckvreader_kopassigner_data[9], 
	ckvreader_kopassigner_data[8], ckvreader_kopassigner_data[7], 
	ckvreader_kopassigner_data[6], ckvreader_kopassigner_data[5], 
	ckvreader_kopassigner_data[4], ckvreader_kopassigner_data[3], 
	ckvreader_kopassigner_data[2], ckvreader_kopassigner_data[1], 
	ckvreader_kopassigner_data[0]});
ixc_assign _zz_strnp_3 ( _zy_simnet_ckv_rd_3_w$, ckv_rd);
ixc_assign_15 _zz_strnp_4 ( _zy_simnet_ckv_addr_4_w$[0:14], ckv_addr[14:0]);
ixc_assign _zz_strnp_5 ( _zy_simnet_ckv_rd_q_7_w$, ckv_rd_q);
ixc_assign _zz_strnp_6 ( _zy_simnet_fifo_out_ack_8_w$, fifo_out_ack);
Q_INV U870 ( .A(rst_n), .Z(_zy_sva_brcm_dek_key_1_reset_or));
Q_AN03 U871 ( .A0(kimreader_ckvreader_data[67]), .A1(kimreader_ckvreader_data[66]), .A2(kimreader_ckvreader_data[65]), .Z(n420));
Q_AN02 U872 ( .A0(kimreader_ckvreader_data[64]), .A1(n420), .Z(n419));
Q_OR02 U873 ( .A0(tlv_word8[58]), .A1(tlv_word8[59]), .Z(n418));
Q_INV U874 ( .A(n418), .Z(n417));
Q_AN03 U875 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n417), .Z(n416));
Q_AN02 U876 ( .A0(n419), .A1(n416), .Z(_zy_sva_b0_t));
Q_OR02 U877 ( .A0(tlv_word9[58]), .A1(tlv_word9[59]), .Z(n415));
Q_INV U878 ( .A(n415), .Z(n414));
Q_AN03 U879 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n414), .Z(n413));
Q_AN02 U880 ( .A0(n419), .A1(n413), .Z(_zy_sva_b1_t));
Q_AN03 U881 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(half_dek), .Z(n411));
Q_AN02 U882 ( .A0(n419), .A1(n411), .Z(_zy_sva_b2_t));
Q_AN02 U883 ( .A0(tlv_word9[58]), .A1(n410), .Z(n409));
Q_AN03 U884 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n409), .Z(n408));
Q_AN02 U885 ( .A0(n419), .A1(n408), .Z(_zy_sva_b3_t));
Q_AN02 U886 ( .A0(n407), .A1(tlv_word8[59]), .Z(n406));
Q_AN03 U887 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n406), .Z(n405));
Q_AN02 U888 ( .A0(n419), .A1(n405), .Z(_zy_sva_b4_t));
Q_AN02 U889 ( .A0(n404), .A1(tlv_word9[59]), .Z(n403));
Q_AN03 U890 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n403), .Z(n402));
Q_AN02 U891 ( .A0(n419), .A1(n402), .Z(_zy_sva_b5_t));
Q_AN02 U892 ( .A0(tlv_word8[58]), .A1(tlv_word8[59]), .Z(n401));
Q_AN03 U893 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n401), .Z(n400));
Q_AN02 U894 ( .A0(n419), .A1(n400), .Z(_zy_sva_b6_t));
Q_AN02 U895 ( .A0(tlv_word9[58]), .A1(tlv_word9[59]), .Z(n399));
Q_AN03 U896 ( .A0(ktype_is_aux_key_only), .A1(ckvreader_kopassigner_valid), .A2(n399), .Z(n398));
Q_AN02 U897 ( .A0(n419), .A1(n398), .Z(_zy_sva_b7_t));
ixc_sample_logic_1_3 _zz_zy_sva_b0 ( _zy_sva_b0, _zy_sva_b0_t);
ixc_sample_logic_1_3 _zz_zy_sva_b1 ( _zy_sva_b1, _zy_sva_b1_t);
ixc_sample_logic_1_3 _zz_zy_sva_b2 ( _zy_sva_b2, _zy_sva_b2_t);
ixc_sample_logic_1_3 _zz_zy_sva_b3 ( _zy_sva_b3, _zy_sva_b3_t);
ixc_sample_logic_1_3 _zz_zy_sva_b4 ( _zy_sva_b4, _zy_sva_b4_t);
ixc_sample_logic_1_3 _zz_zy_sva_b5 ( _zy_sva_b5, _zy_sva_b5_t);
ixc_sample_logic_1_3 _zz_zy_sva_b6 ( _zy_sva_b6, _zy_sva_b6_t);
ixc_sample_logic_1_3 _zz_zy_sva_b7 ( _zy_sva_b7, _zy_sva_b7_t);
wire [2:0] n423 = 3'b000;
Q_ASSERT \ckv_len_0_.brcm_dek_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dek_key_1_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dek_key_1_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n423[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_0_.brcm_dek_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_0_.brcm_dek_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_0_.brcm_dek_key " ASSERT_LINE 296
wire [2:0] n424 = 3'b000;
Q_ASSERT \ckv_len_0_.brcm_dak_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dak_key_2_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dak_key_2_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n424[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_0_.brcm_dak_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_0_.brcm_dak_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_0_.brcm_dak_key " ASSERT_LINE 297
wire [2:0] n425 = 3'b000;
Q_ASSERT \ckv_len_1_.brcm_dek_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dek_key_3_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dek_key_3_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n425[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_1_.brcm_dek_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_1_.brcm_dek_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_1_.brcm_dek_key " ASSERT_LINE 296
wire [2:0] n426 = 3'b000;
Q_ASSERT \ckv_len_1_.brcm_dak_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dak_key_4_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dak_key_4_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n426[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_1_.brcm_dak_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_1_.brcm_dak_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_1_.brcm_dak_key " ASSERT_LINE 297
wire [2:0] n427 = 3'b000;
Q_ASSERT \ckv_len_2_.brcm_dek_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dek_key_5_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dek_key_5_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n427[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_2_.brcm_dek_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_2_.brcm_dek_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_2_.brcm_dek_key " ASSERT_LINE 296
wire [2:0] n428 = 3'b000;
Q_ASSERT \ckv_len_2_.brcm_dak_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dak_key_6_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dak_key_6_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n428[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_2_.brcm_dak_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_2_.brcm_dak_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_2_.brcm_dak_key " ASSERT_LINE 297
wire [2:0] n429 = 3'b000;
Q_ASSERT \ckv_len_3_.brcm_dek_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dek_key_7_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dek_key_7_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n429[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_3_.brcm_dek_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_3_.brcm_dek_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_3_.brcm_dek_key " ASSERT_LINE 296
wire [2:0] n430 = 3'b000;
Q_ASSERT \ckv_len_3_.brcm_dak_key  ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT(_zy_sva_brcm_dak_key_8_cpass[0]), .FAIL_COUNT( ), .CHECK_COUNT(_zy_sva_brcm_dak_key_8_ccheck[0]), .KILL_SIGNAL( ), .SEVERITY(n430[0]));
// pragma CVASTRPROP INSTANCE "\ckv_len_3_.brcm_dak_key " HDL_ASSERT "%"
// pragma CVASTRPROP INSTANCE "\ckv_len_3_.brcm_dak_key " ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/cr_kme/cr_kme_ckv_reader.v"
//pragma CVAINTPROP INSTANCE "\ckv_len_3_.brcm_dak_key " ASSERT_LINE 297
cr_kme_fifo_xcm57 ckv_data_fifo ( .fifo_in_stall( fifo_in_stall), .fifo_out( { 
	fifo_out_mbe, fifo_out[63], fifo_out[62], fifo_out[61], fifo_out[60], 
	fifo_out[59], fifo_out[58], fifo_out[57], fifo_out[56], fifo_out[55], 
	fifo_out[54], fifo_out[53], fifo_out[52], fifo_out[51], fifo_out[50], 
	fifo_out[49], fifo_out[48], fifo_out[47], fifo_out[46], fifo_out[45], 
	fifo_out[44], fifo_out[43], fifo_out[42], fifo_out[41], fifo_out[40], 
	fifo_out[39], fifo_out[38], fifo_out[37], fifo_out[36], fifo_out[35], 
	fifo_out[34], fifo_out[33], fifo_out[32], fifo_out[31], fifo_out[30], 
	fifo_out[29], fifo_out[28], fifo_out[27], fifo_out[26], fifo_out[25], 
	fifo_out[24], fifo_out[23], fifo_out[22], fifo_out[21], fifo_out[20], 
	fifo_out[19], fifo_out[18], fifo_out[17], fifo_out[16], fifo_out[15], 
	fifo_out[14], fifo_out[13], fifo_out[12], fifo_out[11], fifo_out[10], 
	fifo_out[9], fifo_out[8], fifo_out[7], fifo_out[6], fifo_out[5], 
	fifo_out[4], fifo_out[3], fifo_out[2], fifo_out[1], fifo_out[0]}), 
	.fifo_out_valid( fifo_out_valid), .fifo_overflow( _zy_simnet_dio_5), 
	.fifo_underflow( _zy_simnet_dio_6), .clk( clk), .rst_n( rst_n), 
	.fifo_in( { ckv_mbe, ckv_dout[63], ckv_dout[62], ckv_dout[61], 
	ckv_dout[60], ckv_dout[59], ckv_dout[58], ckv_dout[57], ckv_dout[56], 
	ckv_dout[55], ckv_dout[54], ckv_dout[53], ckv_dout[52], ckv_dout[51], 
	ckv_dout[50], ckv_dout[49], ckv_dout[48], ckv_dout[47], ckv_dout[46], 
	ckv_dout[45], ckv_dout[44], ckv_dout[43], ckv_dout[42], ckv_dout[41], 
	ckv_dout[40], ckv_dout[39], ckv_dout[38], ckv_dout[37], ckv_dout[36], 
	ckv_dout[35], ckv_dout[34], ckv_dout[33], ckv_dout[32], ckv_dout[31], 
	ckv_dout[30], ckv_dout[29], ckv_dout[28], ckv_dout[27], ckv_dout[26], 
	ckv_dout[25], ckv_dout[24], ckv_dout[23], ckv_dout[22], ckv_dout[21], 
	ckv_dout[20], ckv_dout[19], ckv_dout[18], ckv_dout[17], ckv_dout[16], 
	ckv_dout[15], ckv_dout[14], ckv_dout[13], ckv_dout[12], ckv_dout[11], 
	ckv_dout[10], ckv_dout[9], ckv_dout[8], ckv_dout[7], ckv_dout[6], 
	ckv_dout[5], ckv_dout[4], ckv_dout[3], ckv_dout[2], ckv_dout[1], 
	ckv_dout[0]}), .fifo_in_valid( _zy_simnet_ckv_rd_q_7_w$), 
	.fifo_out_ack( _zy_simnet_fifo_out_ack_8_w$), 
	.fifo_in_stall_override( _zy_simnet_cio_9));
Q_OA21 U915 ( .A0(fifo_out_valid), .A1(n382), .B0(kimreader_ckvreader_valid), .Z(ckvreader_kopassigner_valid));
Q_MX03 U916 ( .S0(n27), .S1(n10), .A0(tlv_word42[0]), .A1(kimreader_ckvreader_data[0]), .A2(n311), .Z(n50));
Q_MX03 U917 ( .S0(n27), .S1(n10), .A0(tlv_word42[1]), .A1(kimreader_ckvreader_data[1]), .A2(n310), .Z(n49));
Q_MX03 U918 ( .S0(n27), .S1(n10), .A0(tlv_word42[2]), .A1(kimreader_ckvreader_data[2]), .A2(n309), .Z(n48));
Q_MX03 U919 ( .S0(n27), .S1(n10), .A0(tlv_word42[3]), .A1(kimreader_ckvreader_data[3]), .A2(n308), .Z(n47));
Q_MX03 U920 ( .S0(n27), .S1(n10), .A0(tlv_word42[4]), .A1(kimreader_ckvreader_data[4]), .A2(n307), .Z(n46));
Q_MX03 U921 ( .S0(n27), .S1(n10), .A0(tlv_word42[5]), .A1(kimreader_ckvreader_data[5]), .A2(n306), .Z(n45));
Q_MX03 U922 ( .S0(n27), .S1(n10), .A0(tlv_word42[6]), .A1(kimreader_ckvreader_data[6]), .A2(n305), .Z(n44));
Q_MX03 U923 ( .S0(n27), .S1(n10), .A0(tlv_word42[7]), .A1(kimreader_ckvreader_data[7]), .A2(n304), .Z(n43));
Q_FDP4EP \_zy_sva_brcm_dek_key_1_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_1_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_1_cpass_REG[0] ( .CK(clk), .CE(n397), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_1_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_2_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_2_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_2_cpass_REG[0] ( .CK(clk), .CE(n396), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_2_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_3_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_3_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_3_cpass_REG[0] ( .CK(clk), .CE(n395), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_3_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_4_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_4_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_4_cpass_REG[0] ( .CK(clk), .CE(n394), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_4_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_5_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_5_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_5_cpass_REG[0] ( .CK(clk), .CE(n393), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_5_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_6_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_6_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_6_cpass_REG[0] ( .CK(clk), .CE(n392), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_6_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_7_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_7_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dek_key_7_cpass_REG[0] ( .CK(clk), .CE(n391), .R(n2), .D(n1), .Q(_zy_sva_brcm_dek_key_7_cpass[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_8_ccheck_REG[0] ( .CK(clk), .CE(rst_n), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_8_ccheck[0]));
Q_FDP4EP \_zy_sva_brcm_dak_key_8_cpass_REG[0] ( .CK(clk), .CE(n390), .R(n2), .D(n1), .Q(_zy_sva_brcm_dak_key_8_cpass[0]));
Q_FDP4EP \ckv_addr_REG[14] ( .CK(clk), .CE(n318), .R(n421), .D(n327), .Q(ckv_addr[14]));
Q_INV U941 ( .A(rst_n), .Z(n421));
Q_FDP4EP \ckv_addr_REG[13] ( .CK(clk), .CE(n318), .R(n421), .D(n328), .Q(ckv_addr[13]));
Q_FDP4EP \ckv_addr_REG[12] ( .CK(clk), .CE(n318), .R(n421), .D(n329), .Q(ckv_addr[12]));
Q_FDP4EP \ckv_addr_REG[11] ( .CK(clk), .CE(n318), .R(n421), .D(n330), .Q(ckv_addr[11]));
Q_FDP4EP \ckv_addr_REG[10] ( .CK(clk), .CE(n318), .R(n421), .D(n331), .Q(ckv_addr[10]));
Q_FDP4EP \ckv_addr_REG[9] ( .CK(clk), .CE(n318), .R(n421), .D(n332), .Q(ckv_addr[9]));
Q_FDP4EP \ckv_addr_REG[8] ( .CK(clk), .CE(n318), .R(n421), .D(n333), .Q(ckv_addr[8]));
Q_FDP4EP \ckv_addr_REG[7] ( .CK(clk), .CE(n318), .R(n421), .D(n334), .Q(ckv_addr[7]));
Q_FDP4EP \ckv_addr_REG[6] ( .CK(clk), .CE(n318), .R(n421), .D(n335), .Q(ckv_addr[6]));
Q_FDP4EP \ckv_addr_REG[5] ( .CK(clk), .CE(n318), .R(n421), .D(n336), .Q(ckv_addr[5]));
Q_FDP4EP \ckv_addr_REG[4] ( .CK(clk), .CE(n318), .R(n421), .D(n337), .Q(ckv_addr[4]));
Q_FDP4EP \ckv_addr_REG[3] ( .CK(clk), .CE(n318), .R(n421), .D(n338), .Q(ckv_addr[3]));
Q_FDP4EP \ckv_addr_REG[2] ( .CK(clk), .CE(n318), .R(n421), .D(n339), .Q(ckv_addr[2]));
Q_FDP4EP \ckv_addr_REG[1] ( .CK(clk), .CE(n318), .R(n421), .D(n340), .Q(ckv_addr[1]));
Q_FDP4EP \ckv_addr_REG[0] ( .CK(clk), .CE(n318), .R(n421), .D(n341), .Q(ckv_addr[0]));
Q_INV U956 ( .A(ckv_addr[0]), .Z(n379));
Q_FDP4EP \ckv_read_num_REG[3] ( .CK(clk), .CE(n318), .R(n421), .D(n342), .Q(ckv_read_num[3]));
Q_FDP4EP \ckv_read_num_REG[2] ( .CK(clk), .CE(n318), .R(n421), .D(n343), .Q(ckv_read_num[2]));
Q_FDP4EP \ckv_read_num_REG[1] ( .CK(clk), .CE(n318), .R(n421), .D(n344), .Q(ckv_read_num[1]));
Q_INV U960 ( .A(ckv_read_num[1]), .Z(n182));
Q_FDP4EP \ckv_read_num_REG[0] ( .CK(clk), .CE(n318), .R(n421), .D(n345), .Q(ckv_read_num[0]));
Q_INV U962 ( .A(ckv_read_num[0]), .Z(n351));
Q_INV U963 ( .A(n5), .Z(n422));
Q_FDP4EP report_kme_error_REG  ( .CK(clk), .CE(n422), .R(n421), .D(fifo_out_ack), .Q(report_kme_error));
Q_INV U965 ( .A(report_kme_error), .Z(n14));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\ckvreader_kopassigner_data.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\ckvreader_kopassigner_data.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\ckvreader_kopassigner_data.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\ckvreader_kopassigner_data.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\ckvreader_kopassigner_data.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\kimreader_ckvreader_data.sot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\kimreader_ckvreader_data.eoi  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\kimreader_ckvreader_data.eot  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\kimreader_ckvreader_data.id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\kimreader_ckvreader_data.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\tlv_word0.tlv_bip2  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\tlv_word0.resv0  (1,0) 1 12 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\tlv_word0.kdf_dek_iter  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\tlv_word0.keyless_algos  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\tlv_word0.needs_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\tlv_word0.needs_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\tlv_word0.key_type  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\tlv_word0.tlv_frame_num  (1,0) 1 10 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\tlv_word0.tlv_eng_id  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\tlv_word0.tlv_seq_num  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\tlv_word0.tlv_len  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\tlv_word0.tlv_type  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\tlv_word42.corrupt_crc32  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\tlv_word42.unused  (1,0) 1 46 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\tlv_word42.error_code  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\tlv_word8.dek_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\tlv_word8.dek_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\tlv_word8.dek_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\tlv_word8.dek_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\tlv_word8.dek_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\tlv_word8.dek_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\tlv_word8.dek_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\tlv_word8.unused  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\tlv_word8.missing_iv  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\tlv_word8.missing_guid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\tlv_word8.validate_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\tlv_word8.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\tlv_word8.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\tlv_word8.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\nxt_tlv_word8.dek_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\nxt_tlv_word8.dek_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\nxt_tlv_word8.dek_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\nxt_tlv_word8.dek_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\nxt_tlv_word8.dek_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\nxt_tlv_word8.dek_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\nxt_tlv_word8.dek_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\nxt_tlv_word8.unused  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\nxt_tlv_word8.missing_iv  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\nxt_tlv_word8.missing_guid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\nxt_tlv_word8.validate_dek  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\nxt_tlv_word8.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\nxt_tlv_word8.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\nxt_tlv_word8.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\tlv_word9.dak_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\tlv_word9.dak_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\tlv_word9.dak_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\tlv_word9.dak_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\tlv_word9.dak_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\tlv_word9.dak_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\tlv_word9.dak_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\tlv_word9.unused  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\tlv_word9.validate_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\tlv_word9.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\tlv_word9.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\tlv_word9.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\nxt_tlv_word9.dak_kim_entry.valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\nxt_tlv_word9.dak_kim_entry.label_index  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\nxt_tlv_word9.dak_kim_entry.ckv_length  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\nxt_tlv_word9.dak_kim_entry.ckv_pointer  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\nxt_tlv_word9.dak_kim_entry.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\nxt_tlv_word9.dak_kim_entry.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\nxt_tlv_word9.dak_kim_entry.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\nxt_tlv_word9.unused  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\nxt_tlv_word9.validate_dak  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\nxt_tlv_word9.vf_valid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\nxt_tlv_word9.pf_num  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\nxt_tlv_word9.vf_num  (1,0) 1 11 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m78 "\aux_key_ctrl.dak_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m79 "\aux_key_ctrl.dak_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m80 "\aux_key_ctrl.kdf_mode  (1,0) 1 1 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m81 "\aux_key_ctrl.dek_key_op  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m82 "\aux_key_ctrl.dek_key_ref  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "82"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "ckvreader_kopassigner_data 5 \ckvreader_kopassigner_data.sot  \ckvreader_kopassigner_data.eoi  \ckvreader_kopassigner_data.eot  \ckvreader_kopassigner_data.id  \ckvreader_kopassigner_data.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "kimreader_ckvreader_data 5 \kimreader_ckvreader_data.sot  \kimreader_ckvreader_data.eoi  \kimreader_ckvreader_data.eot  \kimreader_ckvreader_data.id  \kimreader_ckvreader_data.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "tlv_word0 12 \tlv_word0.tlv_bip2  \tlv_word0.resv0  \tlv_word0.kdf_dek_iter  \tlv_word0.keyless_algos  \tlv_word0.needs_dek  \tlv_word0.needs_dak  \tlv_word0.key_type  \tlv_word0.tlv_frame_num  \tlv_word0.tlv_eng_id  \tlv_word0.tlv_seq_num  \tlv_word0.tlv_len  \tlv_word0.tlv_type "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "tlv_word42 3 \tlv_word42.corrupt_crc32  \tlv_word42.unused  \tlv_word42.error_code "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "tlv_word8 8 \tlv_word8.dek_kim_entry  { \tlv_word8.dek_kim_entry.valid  \tlv_word8.dek_kim_entry.label_index  \tlv_word8.dek_kim_entry.ckv_length  \tlv_word8.dek_kim_entry.ckv_pointer  \tlv_word8.dek_kim_entry.pf_num  \tlv_word8.dek_kim_entry.vf_num  \tlv_word8.dek_kim_entry.vf_valid  } \tlv_word8.unused  \tlv_word8.missing_iv  \tlv_word8.missing_guid  \tlv_word8.validate_dek  \tlv_word8.vf_valid  \tlv_word8.pf_num  \tlv_word8.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "nxt_tlv_word8 8 \nxt_tlv_word8.dek_kim_entry  { \nxt_tlv_word8.dek_kim_entry.valid  \nxt_tlv_word8.dek_kim_entry.label_index  \nxt_tlv_word8.dek_kim_entry.ckv_length  \nxt_tlv_word8.dek_kim_entry.ckv_pointer  \nxt_tlv_word8.dek_kim_entry.pf_num  \nxt_tlv_word8.dek_kim_entry.vf_num  \nxt_tlv_word8.dek_kim_entry.vf_valid  } \nxt_tlv_word8.unused  \nxt_tlv_word8.missing_iv  \nxt_tlv_word8.missing_guid  \nxt_tlv_word8.validate_dek  \nxt_tlv_word8.vf_valid  \nxt_tlv_word8.pf_num  \nxt_tlv_word8.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "tlv_word9 6 \tlv_word9.dak_kim_entry  { \tlv_word9.dak_kim_entry.valid  \tlv_word9.dak_kim_entry.label_index  \tlv_word9.dak_kim_entry.ckv_length  \tlv_word9.dak_kim_entry.ckv_pointer  \tlv_word9.dak_kim_entry.pf_num  \tlv_word9.dak_kim_entry.vf_num  \tlv_word9.dak_kim_entry.vf_valid  } \tlv_word9.unused  \tlv_word9.validate_dak  \tlv_word9.vf_valid  \tlv_word9.pf_num  \tlv_word9.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "nxt_tlv_word9 6 \nxt_tlv_word9.dak_kim_entry  { \nxt_tlv_word9.dak_kim_entry.valid  \nxt_tlv_word9.dak_kim_entry.label_index  \nxt_tlv_word9.dak_kim_entry.ckv_length  \nxt_tlv_word9.dak_kim_entry.ckv_pointer  \nxt_tlv_word9.dak_kim_entry.pf_num  \nxt_tlv_word9.dak_kim_entry.vf_num  \nxt_tlv_word9.dak_kim_entry.vf_valid  } \nxt_tlv_word9.unused  \nxt_tlv_word9.validate_dak  \nxt_tlv_word9.vf_valid  \nxt_tlv_word9.pf_num  \nxt_tlv_word9.vf_num "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "aux_key_ctrl 5 \aux_key_ctrl.dak_key_op  \aux_key_ctrl.dak_key_ref  \aux_key_ctrl.kdf_mode  \aux_key_ctrl.dek_key_op  \aux_key_ctrl.dek_key_ref "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "9"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 ckv_len 0 3 "
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "ckv_len[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "ckv_len[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "ckv_len[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "ckv_len[0]"
endmodule
