
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_xcm27 ( empty, full, underflow, overflow, used_slots, free_slots, 
	rdata, clk, rst_n, wen, ren, clear, wdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output empty;
output full;
output underflow;
output overflow;
output [1:0] used_slots;
output [1:0] free_slots;
output [127:0] rdata;
input clk;
input rst_n;
input wen;
input ren;
input clear;
input [127:0] wdata;
wire _zy_simnet_underflow_0_w$;
wire _zy_simnet_overflow_1_w$;
wire \depth_n._zy_simnet_overflow_3_w$ ;
wire \depth_n._zy_simnet_underflow_2_w$ ;
wire [1:0] \depth_n.wptr ;
wire [1:0] \depth_n.rptr ;
supply0 n1;
ixc_assign \depth_n._zz_strnp_0 ( underflow, 
	\depth_n._zy_simnet_underflow_2_w$ );
ixc_assign \depth_n._zz_strnp_1 ( overflow, 
	\depth_n._zy_simnet_overflow_3_w$ );
nx_fifo_ctrl_xcm36 \depth_n.fifo_ctrl ( .empty( empty), .full( full), 
	.used_slots( used_slots[1:0]), .free_slots( free_slots[1:0]), 
	.rptr( \depth_n.rptr [1:0]), .wptr( \depth_n.wptr [1:0]), 
	.underflow( \depth_n._zy_simnet_underflow_2_w$ ), .overflow( 
	\depth_n._zy_simnet_overflow_3_w$ ), .clk( clk), .rst_n( rst_n), 
	.wen( wen), .ren( ren), .clear( clear));
Q_AN02 U3 ( .A0(wen), .A1(n2), .Z(n3));
Q_INV U4 ( .A(full), .Z(n2));
Q_AN02 U5 ( .A0(n4), .A1(n13), .Z(rdata[0]));
Q_AN02 U6 ( .A0(n4), .A1(n14), .Z(rdata[1]));
Q_AN02 U7 ( .A0(n4), .A1(n15), .Z(rdata[2]));
Q_AN02 U8 ( .A0(n4), .A1(n16), .Z(rdata[3]));
Q_AN02 U9 ( .A0(n4), .A1(n17), .Z(rdata[4]));
Q_AN02 U10 ( .A0(n4), .A1(n18), .Z(rdata[5]));
Q_AN02 U11 ( .A0(n4), .A1(n19), .Z(rdata[6]));
Q_AN02 U12 ( .A0(n4), .A1(n20), .Z(rdata[7]));
Q_AN02 U13 ( .A0(n4), .A1(n21), .Z(rdata[8]));
Q_AN02 U14 ( .A0(n4), .A1(n22), .Z(rdata[9]));
Q_AN02 U15 ( .A0(n4), .A1(n23), .Z(rdata[10]));
Q_AN02 U16 ( .A0(n4), .A1(n24), .Z(rdata[11]));
Q_AN02 U17 ( .A0(n4), .A1(n25), .Z(rdata[12]));
Q_AN02 U18 ( .A0(n4), .A1(n26), .Z(rdata[13]));
Q_AN02 U19 ( .A0(n4), .A1(n27), .Z(rdata[14]));
Q_AN02 U20 ( .A0(n4), .A1(n28), .Z(rdata[15]));
Q_AN02 U21 ( .A0(n4), .A1(n29), .Z(rdata[16]));
Q_AN02 U22 ( .A0(n4), .A1(n30), .Z(rdata[17]));
Q_AN02 U23 ( .A0(n4), .A1(n31), .Z(rdata[18]));
Q_AN02 U24 ( .A0(n4), .A1(n32), .Z(rdata[19]));
Q_AN02 U25 ( .A0(n4), .A1(n33), .Z(rdata[20]));
Q_AN02 U26 ( .A0(n4), .A1(n34), .Z(rdata[21]));
Q_AN02 U27 ( .A0(n4), .A1(n35), .Z(rdata[22]));
Q_AN02 U28 ( .A0(n4), .A1(n36), .Z(rdata[23]));
Q_AN02 U29 ( .A0(n4), .A1(n37), .Z(rdata[24]));
Q_AN02 U30 ( .A0(n4), .A1(n38), .Z(rdata[25]));
Q_AN02 U31 ( .A0(n4), .A1(n39), .Z(rdata[26]));
Q_AN02 U32 ( .A0(n4), .A1(n40), .Z(rdata[27]));
Q_AN02 U33 ( .A0(n4), .A1(n41), .Z(rdata[28]));
Q_AN02 U34 ( .A0(n4), .A1(n42), .Z(rdata[29]));
Q_AN02 U35 ( .A0(n4), .A1(n43), .Z(rdata[30]));
Q_AN02 U36 ( .A0(n4), .A1(n44), .Z(rdata[31]));
Q_AN02 U37 ( .A0(n4), .A1(n45), .Z(rdata[32]));
Q_AN02 U38 ( .A0(n4), .A1(n46), .Z(rdata[33]));
Q_AN02 U39 ( .A0(n4), .A1(n47), .Z(rdata[34]));
Q_AN02 U40 ( .A0(n4), .A1(n48), .Z(rdata[35]));
Q_AN02 U41 ( .A0(n4), .A1(n49), .Z(rdata[36]));
Q_AN02 U42 ( .A0(n4), .A1(n50), .Z(rdata[37]));
Q_AN02 U43 ( .A0(n4), .A1(n51), .Z(rdata[38]));
Q_AN02 U44 ( .A0(n4), .A1(n52), .Z(rdata[39]));
Q_AN02 U45 ( .A0(n4), .A1(n53), .Z(rdata[40]));
Q_AN02 U46 ( .A0(n4), .A1(n54), .Z(rdata[41]));
Q_AN02 U47 ( .A0(n4), .A1(n55), .Z(rdata[42]));
Q_AN02 U48 ( .A0(n4), .A1(n56), .Z(rdata[43]));
Q_AN02 U49 ( .A0(n4), .A1(n57), .Z(rdata[44]));
Q_AN02 U50 ( .A0(n4), .A1(n58), .Z(rdata[45]));
Q_AN02 U51 ( .A0(n4), .A1(n59), .Z(rdata[46]));
Q_AN02 U52 ( .A0(n4), .A1(n60), .Z(rdata[47]));
Q_AN02 U53 ( .A0(n4), .A1(n61), .Z(rdata[48]));
Q_AN02 U54 ( .A0(n4), .A1(n62), .Z(rdata[49]));
Q_AN02 U55 ( .A0(n4), .A1(n63), .Z(rdata[50]));
Q_AN02 U56 ( .A0(n4), .A1(n64), .Z(rdata[51]));
Q_AN02 U57 ( .A0(n4), .A1(n65), .Z(rdata[52]));
Q_AN02 U58 ( .A0(n4), .A1(n66), .Z(rdata[53]));
Q_AN02 U59 ( .A0(n4), .A1(n67), .Z(rdata[54]));
Q_AN02 U60 ( .A0(n4), .A1(n68), .Z(rdata[55]));
Q_AN02 U61 ( .A0(n4), .A1(n69), .Z(rdata[56]));
Q_AN02 U62 ( .A0(n4), .A1(n70), .Z(rdata[57]));
Q_AN02 U63 ( .A0(n4), .A1(n71), .Z(rdata[58]));
Q_AN02 U64 ( .A0(n4), .A1(n72), .Z(rdata[59]));
Q_AN02 U65 ( .A0(n4), .A1(n73), .Z(rdata[60]));
Q_AN02 U66 ( .A0(n4), .A1(n74), .Z(rdata[61]));
Q_AN02 U67 ( .A0(n4), .A1(n75), .Z(rdata[62]));
Q_AN02 U68 ( .A0(n4), .A1(n76), .Z(rdata[63]));
Q_AN02 U69 ( .A0(n4), .A1(n77), .Z(rdata[64]));
Q_AN02 U70 ( .A0(n4), .A1(n78), .Z(rdata[65]));
Q_AN02 U71 ( .A0(n4), .A1(n79), .Z(rdata[66]));
Q_AN02 U72 ( .A0(n4), .A1(n80), .Z(rdata[67]));
Q_AN02 U73 ( .A0(n4), .A1(n81), .Z(rdata[68]));
Q_AN02 U74 ( .A0(n4), .A1(n82), .Z(rdata[69]));
Q_AN02 U75 ( .A0(n4), .A1(n83), .Z(rdata[70]));
Q_AN02 U76 ( .A0(n4), .A1(n84), .Z(rdata[71]));
Q_AN02 U77 ( .A0(n4), .A1(n85), .Z(rdata[72]));
Q_AN02 U78 ( .A0(n4), .A1(n86), .Z(rdata[73]));
Q_AN02 U79 ( .A0(n4), .A1(n87), .Z(rdata[74]));
Q_AN02 U80 ( .A0(n4), .A1(n88), .Z(rdata[75]));
Q_AN02 U81 ( .A0(n4), .A1(n89), .Z(rdata[76]));
Q_AN02 U82 ( .A0(n4), .A1(n90), .Z(rdata[77]));
Q_AN02 U83 ( .A0(n4), .A1(n91), .Z(rdata[78]));
Q_AN02 U84 ( .A0(n4), .A1(n92), .Z(rdata[79]));
Q_AN02 U85 ( .A0(n4), .A1(n93), .Z(rdata[80]));
Q_AN02 U86 ( .A0(n4), .A1(n94), .Z(rdata[81]));
Q_AN02 U87 ( .A0(n4), .A1(n95), .Z(rdata[82]));
Q_AN02 U88 ( .A0(n4), .A1(n96), .Z(rdata[83]));
Q_AN02 U89 ( .A0(n4), .A1(n97), .Z(rdata[84]));
Q_AN02 U90 ( .A0(n4), .A1(n98), .Z(rdata[85]));
Q_AN02 U91 ( .A0(n4), .A1(n99), .Z(rdata[86]));
Q_AN02 U92 ( .A0(n4), .A1(n100), .Z(rdata[87]));
Q_AN02 U93 ( .A0(n4), .A1(n101), .Z(rdata[88]));
Q_AN02 U94 ( .A0(n4), .A1(n102), .Z(rdata[89]));
Q_AN02 U95 ( .A0(n4), .A1(n103), .Z(rdata[90]));
Q_AN02 U96 ( .A0(n4), .A1(n104), .Z(rdata[91]));
Q_AN02 U97 ( .A0(n4), .A1(n105), .Z(rdata[92]));
Q_AN02 U98 ( .A0(n4), .A1(n106), .Z(rdata[93]));
Q_AN02 U99 ( .A0(n4), .A1(n107), .Z(rdata[94]));
Q_AN02 U100 ( .A0(n4), .A1(n108), .Z(rdata[95]));
Q_AN02 U101 ( .A0(n4), .A1(n109), .Z(rdata[96]));
Q_AN02 U102 ( .A0(n4), .A1(n110), .Z(rdata[97]));
Q_AN02 U103 ( .A0(n4), .A1(n111), .Z(rdata[98]));
Q_AN02 U104 ( .A0(n4), .A1(n112), .Z(rdata[99]));
Q_AN02 U105 ( .A0(n4), .A1(n113), .Z(rdata[100]));
Q_AN02 U106 ( .A0(n4), .A1(n114), .Z(rdata[101]));
Q_AN02 U107 ( .A0(n4), .A1(n115), .Z(rdata[102]));
Q_AN02 U108 ( .A0(n4), .A1(n116), .Z(rdata[103]));
Q_AN02 U109 ( .A0(n4), .A1(n117), .Z(rdata[104]));
Q_AN02 U110 ( .A0(n4), .A1(n118), .Z(rdata[105]));
Q_AN02 U111 ( .A0(n4), .A1(n119), .Z(rdata[106]));
Q_AN02 U112 ( .A0(n4), .A1(n120), .Z(rdata[107]));
Q_AN02 U113 ( .A0(n4), .A1(n121), .Z(rdata[108]));
Q_AN02 U114 ( .A0(n4), .A1(n122), .Z(rdata[109]));
Q_AN02 U115 ( .A0(n4), .A1(n123), .Z(rdata[110]));
Q_AN02 U116 ( .A0(n4), .A1(n124), .Z(rdata[111]));
Q_AN02 U117 ( .A0(n4), .A1(n125), .Z(rdata[112]));
Q_AN02 U118 ( .A0(n4), .A1(n126), .Z(rdata[113]));
Q_AN02 U119 ( .A0(n4), .A1(n127), .Z(rdata[114]));
Q_AN02 U120 ( .A0(n4), .A1(n128), .Z(rdata[115]));
Q_AN02 U121 ( .A0(n4), .A1(n129), .Z(rdata[116]));
Q_AN02 U122 ( .A0(n4), .A1(n130), .Z(rdata[117]));
Q_AN02 U123 ( .A0(n4), .A1(n131), .Z(rdata[118]));
Q_AN02 U124 ( .A0(n4), .A1(n132), .Z(rdata[119]));
Q_AN02 U125 ( .A0(n4), .A1(n133), .Z(rdata[120]));
Q_AN02 U126 ( .A0(n4), .A1(n134), .Z(rdata[121]));
Q_AN02 U127 ( .A0(n4), .A1(n135), .Z(rdata[122]));
Q_AN02 U128 ( .A0(n4), .A1(n136), .Z(rdata[123]));
Q_AN02 U129 ( .A0(n4), .A1(n137), .Z(rdata[124]));
Q_AN02 U130 ( .A0(n4), .A1(n138), .Z(rdata[125]));
Q_AN02 U131 ( .A0(n4), .A1(n139), .Z(rdata[126]));
Q_AN02 U132 ( .A0(n4), .A1(n140), .Z(rdata[127]));
Q_INV U133 ( .A(empty), .Z(n4));
Q_AN02 U134 ( .A0(\depth_n.wptr [0]), .A1(n3), .Z(n5));
Q_AN02 U135 ( .A0(\depth_n.wptr [1]), .A1(n3), .Z(n6));
Q_INV U136 ( .A(n5), .Z(n7));
Q_INV U137 ( .A(n6), .Z(n8));
Q_NR02 U138 ( .A0(n6), .A1(n5), .Z(n9));
Q_AN02 U139 ( .A0(n8), .A1(n5), .Z(n10));
Q_AN02 U140 ( .A0(n6), .A1(n7), .Z(n11));
Q_AN02 U141 ( .A0(n9), .A1(n3), .Z(n12));
Q_MX03 U142 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][0] ), .A1(\depth_n.r_data[1][0] ), .A2(\depth_n.r_data[2][0] ), .Z(n13));
Q_MX03 U143 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][1] ), .A1(\depth_n.r_data[1][1] ), .A2(\depth_n.r_data[2][1] ), .Z(n14));
Q_MX03 U144 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][2] ), .A1(\depth_n.r_data[1][2] ), .A2(\depth_n.r_data[2][2] ), .Z(n15));
Q_MX03 U145 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][3] ), .A1(\depth_n.r_data[1][3] ), .A2(\depth_n.r_data[2][3] ), .Z(n16));
Q_MX03 U146 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][4] ), .A1(\depth_n.r_data[1][4] ), .A2(\depth_n.r_data[2][4] ), .Z(n17));
Q_MX03 U147 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][5] ), .A1(\depth_n.r_data[1][5] ), .A2(\depth_n.r_data[2][5] ), .Z(n18));
Q_MX03 U148 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][6] ), .A1(\depth_n.r_data[1][6] ), .A2(\depth_n.r_data[2][6] ), .Z(n19));
Q_MX03 U149 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][7] ), .A1(\depth_n.r_data[1][7] ), .A2(\depth_n.r_data[2][7] ), .Z(n20));
Q_MX03 U150 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][8] ), .A1(\depth_n.r_data[1][8] ), .A2(\depth_n.r_data[2][8] ), .Z(n21));
Q_MX03 U151 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][9] ), .A1(\depth_n.r_data[1][9] ), .A2(\depth_n.r_data[2][9] ), .Z(n22));
Q_MX03 U152 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][10] ), .A1(\depth_n.r_data[1][10] ), .A2(\depth_n.r_data[2][10] ), .Z(n23));
Q_MX03 U153 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][11] ), .A1(\depth_n.r_data[1][11] ), .A2(\depth_n.r_data[2][11] ), .Z(n24));
Q_MX03 U154 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][12] ), .A1(\depth_n.r_data[1][12] ), .A2(\depth_n.r_data[2][12] ), .Z(n25));
Q_MX03 U155 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][13] ), .A1(\depth_n.r_data[1][13] ), .A2(\depth_n.r_data[2][13] ), .Z(n26));
Q_MX03 U156 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][14] ), .A1(\depth_n.r_data[1][14] ), .A2(\depth_n.r_data[2][14] ), .Z(n27));
Q_MX03 U157 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][15] ), .A1(\depth_n.r_data[1][15] ), .A2(\depth_n.r_data[2][15] ), .Z(n28));
Q_MX03 U158 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][16] ), .A1(\depth_n.r_data[1][16] ), .A2(\depth_n.r_data[2][16] ), .Z(n29));
Q_MX03 U159 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][17] ), .A1(\depth_n.r_data[1][17] ), .A2(\depth_n.r_data[2][17] ), .Z(n30));
Q_MX03 U160 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][18] ), .A1(\depth_n.r_data[1][18] ), .A2(\depth_n.r_data[2][18] ), .Z(n31));
Q_MX03 U161 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][19] ), .A1(\depth_n.r_data[1][19] ), .A2(\depth_n.r_data[2][19] ), .Z(n32));
Q_MX03 U162 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][20] ), .A1(\depth_n.r_data[1][20] ), .A2(\depth_n.r_data[2][20] ), .Z(n33));
Q_MX03 U163 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][21] ), .A1(\depth_n.r_data[1][21] ), .A2(\depth_n.r_data[2][21] ), .Z(n34));
Q_MX03 U164 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][22] ), .A1(\depth_n.r_data[1][22] ), .A2(\depth_n.r_data[2][22] ), .Z(n35));
Q_MX03 U165 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][23] ), .A1(\depth_n.r_data[1][23] ), .A2(\depth_n.r_data[2][23] ), .Z(n36));
Q_MX03 U166 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][24] ), .A1(\depth_n.r_data[1][24] ), .A2(\depth_n.r_data[2][24] ), .Z(n37));
Q_MX03 U167 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][25] ), .A1(\depth_n.r_data[1][25] ), .A2(\depth_n.r_data[2][25] ), .Z(n38));
Q_MX03 U168 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][26] ), .A1(\depth_n.r_data[1][26] ), .A2(\depth_n.r_data[2][26] ), .Z(n39));
Q_MX03 U169 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][27] ), .A1(\depth_n.r_data[1][27] ), .A2(\depth_n.r_data[2][27] ), .Z(n40));
Q_MX03 U170 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][28] ), .A1(\depth_n.r_data[1][28] ), .A2(\depth_n.r_data[2][28] ), .Z(n41));
Q_MX03 U171 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][29] ), .A1(\depth_n.r_data[1][29] ), .A2(\depth_n.r_data[2][29] ), .Z(n42));
Q_MX03 U172 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][30] ), .A1(\depth_n.r_data[1][30] ), .A2(\depth_n.r_data[2][30] ), .Z(n43));
Q_MX03 U173 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][31] ), .A1(\depth_n.r_data[1][31] ), .A2(\depth_n.r_data[2][31] ), .Z(n44));
Q_MX03 U174 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][32] ), .A1(\depth_n.r_data[1][32] ), .A2(\depth_n.r_data[2][32] ), .Z(n45));
Q_MX03 U175 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][33] ), .A1(\depth_n.r_data[1][33] ), .A2(\depth_n.r_data[2][33] ), .Z(n46));
Q_MX03 U176 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][34] ), .A1(\depth_n.r_data[1][34] ), .A2(\depth_n.r_data[2][34] ), .Z(n47));
Q_MX03 U177 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][35] ), .A1(\depth_n.r_data[1][35] ), .A2(\depth_n.r_data[2][35] ), .Z(n48));
Q_MX03 U178 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][36] ), .A1(\depth_n.r_data[1][36] ), .A2(\depth_n.r_data[2][36] ), .Z(n49));
Q_MX03 U179 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][37] ), .A1(\depth_n.r_data[1][37] ), .A2(\depth_n.r_data[2][37] ), .Z(n50));
Q_MX03 U180 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][38] ), .A1(\depth_n.r_data[1][38] ), .A2(\depth_n.r_data[2][38] ), .Z(n51));
Q_MX03 U181 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][39] ), .A1(\depth_n.r_data[1][39] ), .A2(\depth_n.r_data[2][39] ), .Z(n52));
Q_MX03 U182 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][40] ), .A1(\depth_n.r_data[1][40] ), .A2(\depth_n.r_data[2][40] ), .Z(n53));
Q_MX03 U183 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][41] ), .A1(\depth_n.r_data[1][41] ), .A2(\depth_n.r_data[2][41] ), .Z(n54));
Q_MX03 U184 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][42] ), .A1(\depth_n.r_data[1][42] ), .A2(\depth_n.r_data[2][42] ), .Z(n55));
Q_MX03 U185 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][43] ), .A1(\depth_n.r_data[1][43] ), .A2(\depth_n.r_data[2][43] ), .Z(n56));
Q_MX03 U186 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][44] ), .A1(\depth_n.r_data[1][44] ), .A2(\depth_n.r_data[2][44] ), .Z(n57));
Q_MX03 U187 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][45] ), .A1(\depth_n.r_data[1][45] ), .A2(\depth_n.r_data[2][45] ), .Z(n58));
Q_MX03 U188 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][46] ), .A1(\depth_n.r_data[1][46] ), .A2(\depth_n.r_data[2][46] ), .Z(n59));
Q_MX03 U189 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][47] ), .A1(\depth_n.r_data[1][47] ), .A2(\depth_n.r_data[2][47] ), .Z(n60));
Q_MX03 U190 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][48] ), .A1(\depth_n.r_data[1][48] ), .A2(\depth_n.r_data[2][48] ), .Z(n61));
Q_MX03 U191 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][49] ), .A1(\depth_n.r_data[1][49] ), .A2(\depth_n.r_data[2][49] ), .Z(n62));
Q_MX03 U192 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][50] ), .A1(\depth_n.r_data[1][50] ), .A2(\depth_n.r_data[2][50] ), .Z(n63));
Q_MX03 U193 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][51] ), .A1(\depth_n.r_data[1][51] ), .A2(\depth_n.r_data[2][51] ), .Z(n64));
Q_MX03 U194 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][52] ), .A1(\depth_n.r_data[1][52] ), .A2(\depth_n.r_data[2][52] ), .Z(n65));
Q_MX03 U195 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][53] ), .A1(\depth_n.r_data[1][53] ), .A2(\depth_n.r_data[2][53] ), .Z(n66));
Q_MX03 U196 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][54] ), .A1(\depth_n.r_data[1][54] ), .A2(\depth_n.r_data[2][54] ), .Z(n67));
Q_MX03 U197 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][55] ), .A1(\depth_n.r_data[1][55] ), .A2(\depth_n.r_data[2][55] ), .Z(n68));
Q_MX03 U198 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][56] ), .A1(\depth_n.r_data[1][56] ), .A2(\depth_n.r_data[2][56] ), .Z(n69));
Q_MX03 U199 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][57] ), .A1(\depth_n.r_data[1][57] ), .A2(\depth_n.r_data[2][57] ), .Z(n70));
Q_MX03 U200 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][58] ), .A1(\depth_n.r_data[1][58] ), .A2(\depth_n.r_data[2][58] ), .Z(n71));
Q_MX03 U201 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][59] ), .A1(\depth_n.r_data[1][59] ), .A2(\depth_n.r_data[2][59] ), .Z(n72));
Q_MX03 U202 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][60] ), .A1(\depth_n.r_data[1][60] ), .A2(\depth_n.r_data[2][60] ), .Z(n73));
Q_MX03 U203 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][61] ), .A1(\depth_n.r_data[1][61] ), .A2(\depth_n.r_data[2][61] ), .Z(n74));
Q_MX03 U204 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][62] ), .A1(\depth_n.r_data[1][62] ), .A2(\depth_n.r_data[2][62] ), .Z(n75));
Q_MX03 U205 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][63] ), .A1(\depth_n.r_data[1][63] ), .A2(\depth_n.r_data[2][63] ), .Z(n76));
Q_MX03 U206 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][64] ), .A1(\depth_n.r_data[1][64] ), .A2(\depth_n.r_data[2][64] ), .Z(n77));
Q_MX03 U207 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][65] ), .A1(\depth_n.r_data[1][65] ), .A2(\depth_n.r_data[2][65] ), .Z(n78));
Q_MX03 U208 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][66] ), .A1(\depth_n.r_data[1][66] ), .A2(\depth_n.r_data[2][66] ), .Z(n79));
Q_MX03 U209 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][67] ), .A1(\depth_n.r_data[1][67] ), .A2(\depth_n.r_data[2][67] ), .Z(n80));
Q_MX03 U210 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][68] ), .A1(\depth_n.r_data[1][68] ), .A2(\depth_n.r_data[2][68] ), .Z(n81));
Q_MX03 U211 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][69] ), .A1(\depth_n.r_data[1][69] ), .A2(\depth_n.r_data[2][69] ), .Z(n82));
Q_MX03 U212 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][70] ), .A1(\depth_n.r_data[1][70] ), .A2(\depth_n.r_data[2][70] ), .Z(n83));
Q_MX03 U213 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][71] ), .A1(\depth_n.r_data[1][71] ), .A2(\depth_n.r_data[2][71] ), .Z(n84));
Q_MX03 U214 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][72] ), .A1(\depth_n.r_data[1][72] ), .A2(\depth_n.r_data[2][72] ), .Z(n85));
Q_MX03 U215 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][73] ), .A1(\depth_n.r_data[1][73] ), .A2(\depth_n.r_data[2][73] ), .Z(n86));
Q_MX03 U216 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][74] ), .A1(\depth_n.r_data[1][74] ), .A2(\depth_n.r_data[2][74] ), .Z(n87));
Q_MX03 U217 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][75] ), .A1(\depth_n.r_data[1][75] ), .A2(\depth_n.r_data[2][75] ), .Z(n88));
Q_MX03 U218 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][76] ), .A1(\depth_n.r_data[1][76] ), .A2(\depth_n.r_data[2][76] ), .Z(n89));
Q_MX03 U219 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][77] ), .A1(\depth_n.r_data[1][77] ), .A2(\depth_n.r_data[2][77] ), .Z(n90));
Q_MX03 U220 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][78] ), .A1(\depth_n.r_data[1][78] ), .A2(\depth_n.r_data[2][78] ), .Z(n91));
Q_MX03 U221 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][79] ), .A1(\depth_n.r_data[1][79] ), .A2(\depth_n.r_data[2][79] ), .Z(n92));
Q_MX03 U222 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][80] ), .A1(\depth_n.r_data[1][80] ), .A2(\depth_n.r_data[2][80] ), .Z(n93));
Q_MX03 U223 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][81] ), .A1(\depth_n.r_data[1][81] ), .A2(\depth_n.r_data[2][81] ), .Z(n94));
Q_MX03 U224 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][82] ), .A1(\depth_n.r_data[1][82] ), .A2(\depth_n.r_data[2][82] ), .Z(n95));
Q_MX03 U225 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][83] ), .A1(\depth_n.r_data[1][83] ), .A2(\depth_n.r_data[2][83] ), .Z(n96));
Q_MX03 U226 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][84] ), .A1(\depth_n.r_data[1][84] ), .A2(\depth_n.r_data[2][84] ), .Z(n97));
Q_MX03 U227 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][85] ), .A1(\depth_n.r_data[1][85] ), .A2(\depth_n.r_data[2][85] ), .Z(n98));
Q_MX03 U228 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][86] ), .A1(\depth_n.r_data[1][86] ), .A2(\depth_n.r_data[2][86] ), .Z(n99));
Q_MX03 U229 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][87] ), .A1(\depth_n.r_data[1][87] ), .A2(\depth_n.r_data[2][87] ), .Z(n100));
Q_MX03 U230 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][88] ), .A1(\depth_n.r_data[1][88] ), .A2(\depth_n.r_data[2][88] ), .Z(n101));
Q_MX03 U231 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][89] ), .A1(\depth_n.r_data[1][89] ), .A2(\depth_n.r_data[2][89] ), .Z(n102));
Q_MX03 U232 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][90] ), .A1(\depth_n.r_data[1][90] ), .A2(\depth_n.r_data[2][90] ), .Z(n103));
Q_MX03 U233 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][91] ), .A1(\depth_n.r_data[1][91] ), .A2(\depth_n.r_data[2][91] ), .Z(n104));
Q_MX03 U234 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][92] ), .A1(\depth_n.r_data[1][92] ), .A2(\depth_n.r_data[2][92] ), .Z(n105));
Q_MX03 U235 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][93] ), .A1(\depth_n.r_data[1][93] ), .A2(\depth_n.r_data[2][93] ), .Z(n106));
Q_MX03 U236 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][94] ), .A1(\depth_n.r_data[1][94] ), .A2(\depth_n.r_data[2][94] ), .Z(n107));
Q_MX03 U237 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][95] ), .A1(\depth_n.r_data[1][95] ), .A2(\depth_n.r_data[2][95] ), .Z(n108));
Q_MX03 U238 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][96] ), .A1(\depth_n.r_data[1][96] ), .A2(\depth_n.r_data[2][96] ), .Z(n109));
Q_MX03 U239 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][97] ), .A1(\depth_n.r_data[1][97] ), .A2(\depth_n.r_data[2][97] ), .Z(n110));
Q_MX03 U240 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][98] ), .A1(\depth_n.r_data[1][98] ), .A2(\depth_n.r_data[2][98] ), .Z(n111));
Q_MX03 U241 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][99] ), .A1(\depth_n.r_data[1][99] ), .A2(\depth_n.r_data[2][99] ), .Z(n112));
Q_MX03 U242 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][100] ), .A1(\depth_n.r_data[1][100] ), .A2(\depth_n.r_data[2][100] ), .Z(n113));
Q_MX03 U243 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][101] ), .A1(\depth_n.r_data[1][101] ), .A2(\depth_n.r_data[2][101] ), .Z(n114));
Q_MX03 U244 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][102] ), .A1(\depth_n.r_data[1][102] ), .A2(\depth_n.r_data[2][102] ), .Z(n115));
Q_MX03 U245 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][103] ), .A1(\depth_n.r_data[1][103] ), .A2(\depth_n.r_data[2][103] ), .Z(n116));
Q_MX03 U246 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][104] ), .A1(\depth_n.r_data[1][104] ), .A2(\depth_n.r_data[2][104] ), .Z(n117));
Q_MX03 U247 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][105] ), .A1(\depth_n.r_data[1][105] ), .A2(\depth_n.r_data[2][105] ), .Z(n118));
Q_MX03 U248 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][106] ), .A1(\depth_n.r_data[1][106] ), .A2(\depth_n.r_data[2][106] ), .Z(n119));
Q_MX03 U249 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][107] ), .A1(\depth_n.r_data[1][107] ), .A2(\depth_n.r_data[2][107] ), .Z(n120));
Q_MX03 U250 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][108] ), .A1(\depth_n.r_data[1][108] ), .A2(\depth_n.r_data[2][108] ), .Z(n121));
Q_MX03 U251 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][109] ), .A1(\depth_n.r_data[1][109] ), .A2(\depth_n.r_data[2][109] ), .Z(n122));
Q_MX03 U252 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][110] ), .A1(\depth_n.r_data[1][110] ), .A2(\depth_n.r_data[2][110] ), .Z(n123));
Q_MX03 U253 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][111] ), .A1(\depth_n.r_data[1][111] ), .A2(\depth_n.r_data[2][111] ), .Z(n124));
Q_MX03 U254 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][112] ), .A1(\depth_n.r_data[1][112] ), .A2(\depth_n.r_data[2][112] ), .Z(n125));
Q_MX03 U255 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][113] ), .A1(\depth_n.r_data[1][113] ), .A2(\depth_n.r_data[2][113] ), .Z(n126));
Q_MX03 U256 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][114] ), .A1(\depth_n.r_data[1][114] ), .A2(\depth_n.r_data[2][114] ), .Z(n127));
Q_MX03 U257 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][115] ), .A1(\depth_n.r_data[1][115] ), .A2(\depth_n.r_data[2][115] ), .Z(n128));
Q_MX03 U258 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][116] ), .A1(\depth_n.r_data[1][116] ), .A2(\depth_n.r_data[2][116] ), .Z(n129));
Q_MX03 U259 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][117] ), .A1(\depth_n.r_data[1][117] ), .A2(\depth_n.r_data[2][117] ), .Z(n130));
Q_MX03 U260 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][118] ), .A1(\depth_n.r_data[1][118] ), .A2(\depth_n.r_data[2][118] ), .Z(n131));
Q_MX03 U261 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][119] ), .A1(\depth_n.r_data[1][119] ), .A2(\depth_n.r_data[2][119] ), .Z(n132));
Q_MX03 U262 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][120] ), .A1(\depth_n.r_data[1][120] ), .A2(\depth_n.r_data[2][120] ), .Z(n133));
Q_MX03 U263 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][121] ), .A1(\depth_n.r_data[1][121] ), .A2(\depth_n.r_data[2][121] ), .Z(n134));
Q_MX03 U264 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][122] ), .A1(\depth_n.r_data[1][122] ), .A2(\depth_n.r_data[2][122] ), .Z(n135));
Q_MX03 U265 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][123] ), .A1(\depth_n.r_data[1][123] ), .A2(\depth_n.r_data[2][123] ), .Z(n136));
Q_MX03 U266 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][124] ), .A1(\depth_n.r_data[1][124] ), .A2(\depth_n.r_data[2][124] ), .Z(n137));
Q_MX03 U267 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][125] ), .A1(\depth_n.r_data[1][125] ), .A2(\depth_n.r_data[2][125] ), .Z(n138));
Q_MX03 U268 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][126] ), .A1(\depth_n.r_data[1][126] ), .A2(\depth_n.r_data[2][126] ), .Z(n139));
Q_MX03 U269 ( .S0(\depth_n.rptr [0]), .S1(\depth_n.rptr [1]), .A0(\depth_n.r_data[0][127] ), .A1(\depth_n.r_data[1][127] ), .A2(\depth_n.r_data[2][127] ), .Z(n140));
ixc_assign _zz_strnp_2 ( _zy_simnet_underflow_0_w$, underflow);
ixc_assign _zz_strnp_3 ( _zy_simnet_overflow_1_w$, overflow);
Q_FDP4EP \depth_n.r_data_REG[2][127] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[127]), .Q(\depth_n.r_data[2][127] ));
Q_FDP4EP \depth_n.r_data_REG[2][126] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[126]), .Q(\depth_n.r_data[2][126] ));
Q_FDP4EP \depth_n.r_data_REG[2][125] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[125]), .Q(\depth_n.r_data[2][125] ));
Q_FDP4EP \depth_n.r_data_REG[2][124] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[124]), .Q(\depth_n.r_data[2][124] ));
Q_FDP4EP \depth_n.r_data_REG[2][123] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[123]), .Q(\depth_n.r_data[2][123] ));
Q_FDP4EP \depth_n.r_data_REG[2][122] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[122]), .Q(\depth_n.r_data[2][122] ));
Q_FDP4EP \depth_n.r_data_REG[2][121] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[121]), .Q(\depth_n.r_data[2][121] ));
Q_FDP4EP \depth_n.r_data_REG[2][120] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[120]), .Q(\depth_n.r_data[2][120] ));
Q_FDP4EP \depth_n.r_data_REG[2][119] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[119]), .Q(\depth_n.r_data[2][119] ));
Q_FDP4EP \depth_n.r_data_REG[2][118] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[118]), .Q(\depth_n.r_data[2][118] ));
Q_FDP4EP \depth_n.r_data_REG[2][117] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[117]), .Q(\depth_n.r_data[2][117] ));
Q_FDP4EP \depth_n.r_data_REG[2][116] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[116]), .Q(\depth_n.r_data[2][116] ));
Q_FDP4EP \depth_n.r_data_REG[2][115] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[115]), .Q(\depth_n.r_data[2][115] ));
Q_FDP4EP \depth_n.r_data_REG[2][114] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[114]), .Q(\depth_n.r_data[2][114] ));
Q_FDP4EP \depth_n.r_data_REG[2][113] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[113]), .Q(\depth_n.r_data[2][113] ));
Q_FDP4EP \depth_n.r_data_REG[2][112] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[112]), .Q(\depth_n.r_data[2][112] ));
Q_FDP4EP \depth_n.r_data_REG[2][111] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[111]), .Q(\depth_n.r_data[2][111] ));
Q_FDP4EP \depth_n.r_data_REG[2][110] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[110]), .Q(\depth_n.r_data[2][110] ));
Q_FDP4EP \depth_n.r_data_REG[2][109] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[109]), .Q(\depth_n.r_data[2][109] ));
Q_FDP4EP \depth_n.r_data_REG[2][108] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[108]), .Q(\depth_n.r_data[2][108] ));
Q_FDP4EP \depth_n.r_data_REG[2][107] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[107]), .Q(\depth_n.r_data[2][107] ));
Q_FDP4EP \depth_n.r_data_REG[2][106] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[106]), .Q(\depth_n.r_data[2][106] ));
Q_FDP4EP \depth_n.r_data_REG[2][105] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[105]), .Q(\depth_n.r_data[2][105] ));
Q_FDP4EP \depth_n.r_data_REG[2][104] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[104]), .Q(\depth_n.r_data[2][104] ));
Q_FDP4EP \depth_n.r_data_REG[2][103] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[103]), .Q(\depth_n.r_data[2][103] ));
Q_FDP4EP \depth_n.r_data_REG[2][102] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[102]), .Q(\depth_n.r_data[2][102] ));
Q_FDP4EP \depth_n.r_data_REG[2][101] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[101]), .Q(\depth_n.r_data[2][101] ));
Q_FDP4EP \depth_n.r_data_REG[2][100] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[100]), .Q(\depth_n.r_data[2][100] ));
Q_FDP4EP \depth_n.r_data_REG[2][99] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[99]), .Q(\depth_n.r_data[2][99] ));
Q_FDP4EP \depth_n.r_data_REG[2][98] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[98]), .Q(\depth_n.r_data[2][98] ));
Q_FDP4EP \depth_n.r_data_REG[2][97] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[97]), .Q(\depth_n.r_data[2][97] ));
Q_FDP4EP \depth_n.r_data_REG[2][96] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[96]), .Q(\depth_n.r_data[2][96] ));
Q_FDP4EP \depth_n.r_data_REG[2][95] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[95]), .Q(\depth_n.r_data[2][95] ));
Q_FDP4EP \depth_n.r_data_REG[2][94] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[94]), .Q(\depth_n.r_data[2][94] ));
Q_FDP4EP \depth_n.r_data_REG[2][93] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[93]), .Q(\depth_n.r_data[2][93] ));
Q_FDP4EP \depth_n.r_data_REG[2][92] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[92]), .Q(\depth_n.r_data[2][92] ));
Q_FDP4EP \depth_n.r_data_REG[2][91] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[91]), .Q(\depth_n.r_data[2][91] ));
Q_FDP4EP \depth_n.r_data_REG[2][90] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[90]), .Q(\depth_n.r_data[2][90] ));
Q_FDP4EP \depth_n.r_data_REG[2][89] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[89]), .Q(\depth_n.r_data[2][89] ));
Q_FDP4EP \depth_n.r_data_REG[2][88] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[88]), .Q(\depth_n.r_data[2][88] ));
Q_FDP4EP \depth_n.r_data_REG[2][87] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[87]), .Q(\depth_n.r_data[2][87] ));
Q_FDP4EP \depth_n.r_data_REG[2][86] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[86]), .Q(\depth_n.r_data[2][86] ));
Q_FDP4EP \depth_n.r_data_REG[2][85] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[85]), .Q(\depth_n.r_data[2][85] ));
Q_FDP4EP \depth_n.r_data_REG[2][84] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[84]), .Q(\depth_n.r_data[2][84] ));
Q_FDP4EP \depth_n.r_data_REG[2][83] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[83]), .Q(\depth_n.r_data[2][83] ));
Q_FDP4EP \depth_n.r_data_REG[2][82] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[82]), .Q(\depth_n.r_data[2][82] ));
Q_FDP4EP \depth_n.r_data_REG[2][81] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[81]), .Q(\depth_n.r_data[2][81] ));
Q_FDP4EP \depth_n.r_data_REG[2][80] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[80]), .Q(\depth_n.r_data[2][80] ));
Q_FDP4EP \depth_n.r_data_REG[2][79] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[79]), .Q(\depth_n.r_data[2][79] ));
Q_FDP4EP \depth_n.r_data_REG[2][78] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[78]), .Q(\depth_n.r_data[2][78] ));
Q_FDP4EP \depth_n.r_data_REG[2][77] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[77]), .Q(\depth_n.r_data[2][77] ));
Q_FDP4EP \depth_n.r_data_REG[2][76] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[76]), .Q(\depth_n.r_data[2][76] ));
Q_FDP4EP \depth_n.r_data_REG[2][75] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[75]), .Q(\depth_n.r_data[2][75] ));
Q_FDP4EP \depth_n.r_data_REG[2][74] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[74]), .Q(\depth_n.r_data[2][74] ));
Q_FDP4EP \depth_n.r_data_REG[2][73] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[73]), .Q(\depth_n.r_data[2][73] ));
Q_FDP4EP \depth_n.r_data_REG[2][72] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[72]), .Q(\depth_n.r_data[2][72] ));
Q_FDP4EP \depth_n.r_data_REG[2][71] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[71]), .Q(\depth_n.r_data[2][71] ));
Q_FDP4EP \depth_n.r_data_REG[2][70] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[70]), .Q(\depth_n.r_data[2][70] ));
Q_FDP4EP \depth_n.r_data_REG[2][69] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[69]), .Q(\depth_n.r_data[2][69] ));
Q_FDP4EP \depth_n.r_data_REG[2][68] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[68]), .Q(\depth_n.r_data[2][68] ));
Q_FDP4EP \depth_n.r_data_REG[2][67] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[67]), .Q(\depth_n.r_data[2][67] ));
Q_FDP4EP \depth_n.r_data_REG[2][66] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[66]), .Q(\depth_n.r_data[2][66] ));
Q_FDP4EP \depth_n.r_data_REG[2][65] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[65]), .Q(\depth_n.r_data[2][65] ));
Q_FDP4EP \depth_n.r_data_REG[2][64] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[64]), .Q(\depth_n.r_data[2][64] ));
Q_FDP4EP \depth_n.r_data_REG[2][63] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[63]), .Q(\depth_n.r_data[2][63] ));
Q_FDP4EP \depth_n.r_data_REG[2][62] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[62]), .Q(\depth_n.r_data[2][62] ));
Q_FDP4EP \depth_n.r_data_REG[2][61] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[61]), .Q(\depth_n.r_data[2][61] ));
Q_FDP4EP \depth_n.r_data_REG[2][60] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[60]), .Q(\depth_n.r_data[2][60] ));
Q_FDP4EP \depth_n.r_data_REG[2][59] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[59]), .Q(\depth_n.r_data[2][59] ));
Q_FDP4EP \depth_n.r_data_REG[2][58] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[58]), .Q(\depth_n.r_data[2][58] ));
Q_FDP4EP \depth_n.r_data_REG[2][57] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[57]), .Q(\depth_n.r_data[2][57] ));
Q_FDP4EP \depth_n.r_data_REG[2][56] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[56]), .Q(\depth_n.r_data[2][56] ));
Q_FDP4EP \depth_n.r_data_REG[2][55] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[55]), .Q(\depth_n.r_data[2][55] ));
Q_FDP4EP \depth_n.r_data_REG[2][54] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[54]), .Q(\depth_n.r_data[2][54] ));
Q_FDP4EP \depth_n.r_data_REG[2][53] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[53]), .Q(\depth_n.r_data[2][53] ));
Q_FDP4EP \depth_n.r_data_REG[2][52] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[52]), .Q(\depth_n.r_data[2][52] ));
Q_FDP4EP \depth_n.r_data_REG[2][51] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[51]), .Q(\depth_n.r_data[2][51] ));
Q_FDP4EP \depth_n.r_data_REG[2][50] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[50]), .Q(\depth_n.r_data[2][50] ));
Q_FDP4EP \depth_n.r_data_REG[2][49] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[49]), .Q(\depth_n.r_data[2][49] ));
Q_FDP4EP \depth_n.r_data_REG[2][48] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[48]), .Q(\depth_n.r_data[2][48] ));
Q_FDP4EP \depth_n.r_data_REG[2][47] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[47]), .Q(\depth_n.r_data[2][47] ));
Q_FDP4EP \depth_n.r_data_REG[2][46] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[46]), .Q(\depth_n.r_data[2][46] ));
Q_FDP4EP \depth_n.r_data_REG[2][45] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[45]), .Q(\depth_n.r_data[2][45] ));
Q_FDP4EP \depth_n.r_data_REG[2][44] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[44]), .Q(\depth_n.r_data[2][44] ));
Q_FDP4EP \depth_n.r_data_REG[2][43] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[43]), .Q(\depth_n.r_data[2][43] ));
Q_FDP4EP \depth_n.r_data_REG[2][42] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[42]), .Q(\depth_n.r_data[2][42] ));
Q_FDP4EP \depth_n.r_data_REG[2][41] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[41]), .Q(\depth_n.r_data[2][41] ));
Q_FDP4EP \depth_n.r_data_REG[2][40] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[40]), .Q(\depth_n.r_data[2][40] ));
Q_FDP4EP \depth_n.r_data_REG[2][39] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[39]), .Q(\depth_n.r_data[2][39] ));
Q_FDP4EP \depth_n.r_data_REG[2][38] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[38]), .Q(\depth_n.r_data[2][38] ));
Q_FDP4EP \depth_n.r_data_REG[2][37] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[37]), .Q(\depth_n.r_data[2][37] ));
Q_FDP4EP \depth_n.r_data_REG[2][36] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[36]), .Q(\depth_n.r_data[2][36] ));
Q_FDP4EP \depth_n.r_data_REG[2][35] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[35]), .Q(\depth_n.r_data[2][35] ));
Q_FDP4EP \depth_n.r_data_REG[2][34] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[34]), .Q(\depth_n.r_data[2][34] ));
Q_FDP4EP \depth_n.r_data_REG[2][33] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[33]), .Q(\depth_n.r_data[2][33] ));
Q_FDP4EP \depth_n.r_data_REG[2][32] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[32]), .Q(\depth_n.r_data[2][32] ));
Q_FDP4EP \depth_n.r_data_REG[2][31] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[31]), .Q(\depth_n.r_data[2][31] ));
Q_FDP4EP \depth_n.r_data_REG[2][30] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[30]), .Q(\depth_n.r_data[2][30] ));
Q_FDP4EP \depth_n.r_data_REG[2][29] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[29]), .Q(\depth_n.r_data[2][29] ));
Q_FDP4EP \depth_n.r_data_REG[2][28] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[28]), .Q(\depth_n.r_data[2][28] ));
Q_FDP4EP \depth_n.r_data_REG[2][27] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[27]), .Q(\depth_n.r_data[2][27] ));
Q_FDP4EP \depth_n.r_data_REG[2][26] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[26]), .Q(\depth_n.r_data[2][26] ));
Q_FDP4EP \depth_n.r_data_REG[2][25] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[25]), .Q(\depth_n.r_data[2][25] ));
Q_FDP4EP \depth_n.r_data_REG[2][24] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[24]), .Q(\depth_n.r_data[2][24] ));
Q_FDP4EP \depth_n.r_data_REG[2][23] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[23]), .Q(\depth_n.r_data[2][23] ));
Q_FDP4EP \depth_n.r_data_REG[2][22] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[22]), .Q(\depth_n.r_data[2][22] ));
Q_FDP4EP \depth_n.r_data_REG[2][21] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[21]), .Q(\depth_n.r_data[2][21] ));
Q_FDP4EP \depth_n.r_data_REG[2][20] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[20]), .Q(\depth_n.r_data[2][20] ));
Q_FDP4EP \depth_n.r_data_REG[2][19] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[19]), .Q(\depth_n.r_data[2][19] ));
Q_FDP4EP \depth_n.r_data_REG[2][18] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[18]), .Q(\depth_n.r_data[2][18] ));
Q_FDP4EP \depth_n.r_data_REG[2][17] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[17]), .Q(\depth_n.r_data[2][17] ));
Q_FDP4EP \depth_n.r_data_REG[2][16] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[16]), .Q(\depth_n.r_data[2][16] ));
Q_FDP4EP \depth_n.r_data_REG[2][15] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[15]), .Q(\depth_n.r_data[2][15] ));
Q_FDP4EP \depth_n.r_data_REG[2][14] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[14]), .Q(\depth_n.r_data[2][14] ));
Q_FDP4EP \depth_n.r_data_REG[2][13] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[13]), .Q(\depth_n.r_data[2][13] ));
Q_FDP4EP \depth_n.r_data_REG[2][12] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[12]), .Q(\depth_n.r_data[2][12] ));
Q_FDP4EP \depth_n.r_data_REG[2][11] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[11]), .Q(\depth_n.r_data[2][11] ));
Q_FDP4EP \depth_n.r_data_REG[2][10] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[10]), .Q(\depth_n.r_data[2][10] ));
Q_FDP4EP \depth_n.r_data_REG[2][9] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[9]), .Q(\depth_n.r_data[2][9] ));
Q_FDP4EP \depth_n.r_data_REG[2][8] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[8]), .Q(\depth_n.r_data[2][8] ));
Q_FDP4EP \depth_n.r_data_REG[2][7] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[7]), .Q(\depth_n.r_data[2][7] ));
Q_FDP4EP \depth_n.r_data_REG[2][6] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[6]), .Q(\depth_n.r_data[2][6] ));
Q_FDP4EP \depth_n.r_data_REG[2][5] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[5]), .Q(\depth_n.r_data[2][5] ));
Q_FDP4EP \depth_n.r_data_REG[2][4] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[4]), .Q(\depth_n.r_data[2][4] ));
Q_FDP4EP \depth_n.r_data_REG[2][3] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[3]), .Q(\depth_n.r_data[2][3] ));
Q_FDP4EP \depth_n.r_data_REG[2][2] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[2]), .Q(\depth_n.r_data[2][2] ));
Q_FDP4EP \depth_n.r_data_REG[2][1] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[1]), .Q(\depth_n.r_data[2][1] ));
Q_FDP4EP \depth_n.r_data_REG[2][0] ( .CK(clk), .CE(n11), .R(n1), .D(wdata[0]), .Q(\depth_n.r_data[2][0] ));
Q_FDP4EP \depth_n.r_data_REG[1][127] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[127]), .Q(\depth_n.r_data[1][127] ));
Q_FDP4EP \depth_n.r_data_REG[1][126] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[126]), .Q(\depth_n.r_data[1][126] ));
Q_FDP4EP \depth_n.r_data_REG[1][125] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[125]), .Q(\depth_n.r_data[1][125] ));
Q_FDP4EP \depth_n.r_data_REG[1][124] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[124]), .Q(\depth_n.r_data[1][124] ));
Q_FDP4EP \depth_n.r_data_REG[1][123] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[123]), .Q(\depth_n.r_data[1][123] ));
Q_FDP4EP \depth_n.r_data_REG[1][122] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[122]), .Q(\depth_n.r_data[1][122] ));
Q_FDP4EP \depth_n.r_data_REG[1][121] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[121]), .Q(\depth_n.r_data[1][121] ));
Q_FDP4EP \depth_n.r_data_REG[1][120] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[120]), .Q(\depth_n.r_data[1][120] ));
Q_FDP4EP \depth_n.r_data_REG[1][119] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[119]), .Q(\depth_n.r_data[1][119] ));
Q_FDP4EP \depth_n.r_data_REG[1][118] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[118]), .Q(\depth_n.r_data[1][118] ));
Q_FDP4EP \depth_n.r_data_REG[1][117] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[117]), .Q(\depth_n.r_data[1][117] ));
Q_FDP4EP \depth_n.r_data_REG[1][116] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[116]), .Q(\depth_n.r_data[1][116] ));
Q_FDP4EP \depth_n.r_data_REG[1][115] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[115]), .Q(\depth_n.r_data[1][115] ));
Q_FDP4EP \depth_n.r_data_REG[1][114] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[114]), .Q(\depth_n.r_data[1][114] ));
Q_FDP4EP \depth_n.r_data_REG[1][113] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[113]), .Q(\depth_n.r_data[1][113] ));
Q_FDP4EP \depth_n.r_data_REG[1][112] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[112]), .Q(\depth_n.r_data[1][112] ));
Q_FDP4EP \depth_n.r_data_REG[1][111] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[111]), .Q(\depth_n.r_data[1][111] ));
Q_FDP4EP \depth_n.r_data_REG[1][110] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[110]), .Q(\depth_n.r_data[1][110] ));
Q_FDP4EP \depth_n.r_data_REG[1][109] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[109]), .Q(\depth_n.r_data[1][109] ));
Q_FDP4EP \depth_n.r_data_REG[1][108] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[108]), .Q(\depth_n.r_data[1][108] ));
Q_FDP4EP \depth_n.r_data_REG[1][107] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[107]), .Q(\depth_n.r_data[1][107] ));
Q_FDP4EP \depth_n.r_data_REG[1][106] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[106]), .Q(\depth_n.r_data[1][106] ));
Q_FDP4EP \depth_n.r_data_REG[1][105] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[105]), .Q(\depth_n.r_data[1][105] ));
Q_FDP4EP \depth_n.r_data_REG[1][104] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[104]), .Q(\depth_n.r_data[1][104] ));
Q_FDP4EP \depth_n.r_data_REG[1][103] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[103]), .Q(\depth_n.r_data[1][103] ));
Q_FDP4EP \depth_n.r_data_REG[1][102] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[102]), .Q(\depth_n.r_data[1][102] ));
Q_FDP4EP \depth_n.r_data_REG[1][101] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[101]), .Q(\depth_n.r_data[1][101] ));
Q_FDP4EP \depth_n.r_data_REG[1][100] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[100]), .Q(\depth_n.r_data[1][100] ));
Q_FDP4EP \depth_n.r_data_REG[1][99] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[99]), .Q(\depth_n.r_data[1][99] ));
Q_FDP4EP \depth_n.r_data_REG[1][98] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[98]), .Q(\depth_n.r_data[1][98] ));
Q_FDP4EP \depth_n.r_data_REG[1][97] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[97]), .Q(\depth_n.r_data[1][97] ));
Q_FDP4EP \depth_n.r_data_REG[1][96] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[96]), .Q(\depth_n.r_data[1][96] ));
Q_FDP4EP \depth_n.r_data_REG[1][95] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[95]), .Q(\depth_n.r_data[1][95] ));
Q_FDP4EP \depth_n.r_data_REG[1][94] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[94]), .Q(\depth_n.r_data[1][94] ));
Q_FDP4EP \depth_n.r_data_REG[1][93] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[93]), .Q(\depth_n.r_data[1][93] ));
Q_FDP4EP \depth_n.r_data_REG[1][92] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[92]), .Q(\depth_n.r_data[1][92] ));
Q_FDP4EP \depth_n.r_data_REG[1][91] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[91]), .Q(\depth_n.r_data[1][91] ));
Q_FDP4EP \depth_n.r_data_REG[1][90] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[90]), .Q(\depth_n.r_data[1][90] ));
Q_FDP4EP \depth_n.r_data_REG[1][89] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[89]), .Q(\depth_n.r_data[1][89] ));
Q_FDP4EP \depth_n.r_data_REG[1][88] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[88]), .Q(\depth_n.r_data[1][88] ));
Q_FDP4EP \depth_n.r_data_REG[1][87] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[87]), .Q(\depth_n.r_data[1][87] ));
Q_FDP4EP \depth_n.r_data_REG[1][86] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[86]), .Q(\depth_n.r_data[1][86] ));
Q_FDP4EP \depth_n.r_data_REG[1][85] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[85]), .Q(\depth_n.r_data[1][85] ));
Q_FDP4EP \depth_n.r_data_REG[1][84] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[84]), .Q(\depth_n.r_data[1][84] ));
Q_FDP4EP \depth_n.r_data_REG[1][83] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[83]), .Q(\depth_n.r_data[1][83] ));
Q_FDP4EP \depth_n.r_data_REG[1][82] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[82]), .Q(\depth_n.r_data[1][82] ));
Q_FDP4EP \depth_n.r_data_REG[1][81] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[81]), .Q(\depth_n.r_data[1][81] ));
Q_FDP4EP \depth_n.r_data_REG[1][80] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[80]), .Q(\depth_n.r_data[1][80] ));
Q_FDP4EP \depth_n.r_data_REG[1][79] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[79]), .Q(\depth_n.r_data[1][79] ));
Q_FDP4EP \depth_n.r_data_REG[1][78] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[78]), .Q(\depth_n.r_data[1][78] ));
Q_FDP4EP \depth_n.r_data_REG[1][77] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[77]), .Q(\depth_n.r_data[1][77] ));
Q_FDP4EP \depth_n.r_data_REG[1][76] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[76]), .Q(\depth_n.r_data[1][76] ));
Q_FDP4EP \depth_n.r_data_REG[1][75] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[75]), .Q(\depth_n.r_data[1][75] ));
Q_FDP4EP \depth_n.r_data_REG[1][74] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[74]), .Q(\depth_n.r_data[1][74] ));
Q_FDP4EP \depth_n.r_data_REG[1][73] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[73]), .Q(\depth_n.r_data[1][73] ));
Q_FDP4EP \depth_n.r_data_REG[1][72] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[72]), .Q(\depth_n.r_data[1][72] ));
Q_FDP4EP \depth_n.r_data_REG[1][71] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[71]), .Q(\depth_n.r_data[1][71] ));
Q_FDP4EP \depth_n.r_data_REG[1][70] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[70]), .Q(\depth_n.r_data[1][70] ));
Q_FDP4EP \depth_n.r_data_REG[1][69] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[69]), .Q(\depth_n.r_data[1][69] ));
Q_FDP4EP \depth_n.r_data_REG[1][68] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[68]), .Q(\depth_n.r_data[1][68] ));
Q_FDP4EP \depth_n.r_data_REG[1][67] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[67]), .Q(\depth_n.r_data[1][67] ));
Q_FDP4EP \depth_n.r_data_REG[1][66] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[66]), .Q(\depth_n.r_data[1][66] ));
Q_FDP4EP \depth_n.r_data_REG[1][65] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[65]), .Q(\depth_n.r_data[1][65] ));
Q_FDP4EP \depth_n.r_data_REG[1][64] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[64]), .Q(\depth_n.r_data[1][64] ));
Q_FDP4EP \depth_n.r_data_REG[1][63] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[63]), .Q(\depth_n.r_data[1][63] ));
Q_FDP4EP \depth_n.r_data_REG[1][62] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[62]), .Q(\depth_n.r_data[1][62] ));
Q_FDP4EP \depth_n.r_data_REG[1][61] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[61]), .Q(\depth_n.r_data[1][61] ));
Q_FDP4EP \depth_n.r_data_REG[1][60] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[60]), .Q(\depth_n.r_data[1][60] ));
Q_FDP4EP \depth_n.r_data_REG[1][59] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[59]), .Q(\depth_n.r_data[1][59] ));
Q_FDP4EP \depth_n.r_data_REG[1][58] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[58]), .Q(\depth_n.r_data[1][58] ));
Q_FDP4EP \depth_n.r_data_REG[1][57] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[57]), .Q(\depth_n.r_data[1][57] ));
Q_FDP4EP \depth_n.r_data_REG[1][56] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[56]), .Q(\depth_n.r_data[1][56] ));
Q_FDP4EP \depth_n.r_data_REG[1][55] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[55]), .Q(\depth_n.r_data[1][55] ));
Q_FDP4EP \depth_n.r_data_REG[1][54] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[54]), .Q(\depth_n.r_data[1][54] ));
Q_FDP4EP \depth_n.r_data_REG[1][53] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[53]), .Q(\depth_n.r_data[1][53] ));
Q_FDP4EP \depth_n.r_data_REG[1][52] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[52]), .Q(\depth_n.r_data[1][52] ));
Q_FDP4EP \depth_n.r_data_REG[1][51] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[51]), .Q(\depth_n.r_data[1][51] ));
Q_FDP4EP \depth_n.r_data_REG[1][50] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[50]), .Q(\depth_n.r_data[1][50] ));
Q_FDP4EP \depth_n.r_data_REG[1][49] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[49]), .Q(\depth_n.r_data[1][49] ));
Q_FDP4EP \depth_n.r_data_REG[1][48] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[48]), .Q(\depth_n.r_data[1][48] ));
Q_FDP4EP \depth_n.r_data_REG[1][47] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[47]), .Q(\depth_n.r_data[1][47] ));
Q_FDP4EP \depth_n.r_data_REG[1][46] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[46]), .Q(\depth_n.r_data[1][46] ));
Q_FDP4EP \depth_n.r_data_REG[1][45] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[45]), .Q(\depth_n.r_data[1][45] ));
Q_FDP4EP \depth_n.r_data_REG[1][44] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[44]), .Q(\depth_n.r_data[1][44] ));
Q_FDP4EP \depth_n.r_data_REG[1][43] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[43]), .Q(\depth_n.r_data[1][43] ));
Q_FDP4EP \depth_n.r_data_REG[1][42] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[42]), .Q(\depth_n.r_data[1][42] ));
Q_FDP4EP \depth_n.r_data_REG[1][41] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[41]), .Q(\depth_n.r_data[1][41] ));
Q_FDP4EP \depth_n.r_data_REG[1][40] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[40]), .Q(\depth_n.r_data[1][40] ));
Q_FDP4EP \depth_n.r_data_REG[1][39] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[39]), .Q(\depth_n.r_data[1][39] ));
Q_FDP4EP \depth_n.r_data_REG[1][38] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[38]), .Q(\depth_n.r_data[1][38] ));
Q_FDP4EP \depth_n.r_data_REG[1][37] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[37]), .Q(\depth_n.r_data[1][37] ));
Q_FDP4EP \depth_n.r_data_REG[1][36] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[36]), .Q(\depth_n.r_data[1][36] ));
Q_FDP4EP \depth_n.r_data_REG[1][35] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[35]), .Q(\depth_n.r_data[1][35] ));
Q_FDP4EP \depth_n.r_data_REG[1][34] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[34]), .Q(\depth_n.r_data[1][34] ));
Q_FDP4EP \depth_n.r_data_REG[1][33] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[33]), .Q(\depth_n.r_data[1][33] ));
Q_FDP4EP \depth_n.r_data_REG[1][32] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[32]), .Q(\depth_n.r_data[1][32] ));
Q_FDP4EP \depth_n.r_data_REG[1][31] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[31]), .Q(\depth_n.r_data[1][31] ));
Q_FDP4EP \depth_n.r_data_REG[1][30] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[30]), .Q(\depth_n.r_data[1][30] ));
Q_FDP4EP \depth_n.r_data_REG[1][29] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[29]), .Q(\depth_n.r_data[1][29] ));
Q_FDP4EP \depth_n.r_data_REG[1][28] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[28]), .Q(\depth_n.r_data[1][28] ));
Q_FDP4EP \depth_n.r_data_REG[1][27] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[27]), .Q(\depth_n.r_data[1][27] ));
Q_FDP4EP \depth_n.r_data_REG[1][26] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[26]), .Q(\depth_n.r_data[1][26] ));
Q_FDP4EP \depth_n.r_data_REG[1][25] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[25]), .Q(\depth_n.r_data[1][25] ));
Q_FDP4EP \depth_n.r_data_REG[1][24] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[24]), .Q(\depth_n.r_data[1][24] ));
Q_FDP4EP \depth_n.r_data_REG[1][23] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[23]), .Q(\depth_n.r_data[1][23] ));
Q_FDP4EP \depth_n.r_data_REG[1][22] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[22]), .Q(\depth_n.r_data[1][22] ));
Q_FDP4EP \depth_n.r_data_REG[1][21] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[21]), .Q(\depth_n.r_data[1][21] ));
Q_FDP4EP \depth_n.r_data_REG[1][20] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[20]), .Q(\depth_n.r_data[1][20] ));
Q_FDP4EP \depth_n.r_data_REG[1][19] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[19]), .Q(\depth_n.r_data[1][19] ));
Q_FDP4EP \depth_n.r_data_REG[1][18] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[18]), .Q(\depth_n.r_data[1][18] ));
Q_FDP4EP \depth_n.r_data_REG[1][17] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[17]), .Q(\depth_n.r_data[1][17] ));
Q_FDP4EP \depth_n.r_data_REG[1][16] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[16]), .Q(\depth_n.r_data[1][16] ));
Q_FDP4EP \depth_n.r_data_REG[1][15] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[15]), .Q(\depth_n.r_data[1][15] ));
Q_FDP4EP \depth_n.r_data_REG[1][14] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[14]), .Q(\depth_n.r_data[1][14] ));
Q_FDP4EP \depth_n.r_data_REG[1][13] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[13]), .Q(\depth_n.r_data[1][13] ));
Q_FDP4EP \depth_n.r_data_REG[1][12] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[12]), .Q(\depth_n.r_data[1][12] ));
Q_FDP4EP \depth_n.r_data_REG[1][11] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[11]), .Q(\depth_n.r_data[1][11] ));
Q_FDP4EP \depth_n.r_data_REG[1][10] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[10]), .Q(\depth_n.r_data[1][10] ));
Q_FDP4EP \depth_n.r_data_REG[1][9] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[9]), .Q(\depth_n.r_data[1][9] ));
Q_FDP4EP \depth_n.r_data_REG[1][8] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[8]), .Q(\depth_n.r_data[1][8] ));
Q_FDP4EP \depth_n.r_data_REG[1][7] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[7]), .Q(\depth_n.r_data[1][7] ));
Q_FDP4EP \depth_n.r_data_REG[1][6] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[6]), .Q(\depth_n.r_data[1][6] ));
Q_FDP4EP \depth_n.r_data_REG[1][5] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[5]), .Q(\depth_n.r_data[1][5] ));
Q_FDP4EP \depth_n.r_data_REG[1][4] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[4]), .Q(\depth_n.r_data[1][4] ));
Q_FDP4EP \depth_n.r_data_REG[1][3] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[3]), .Q(\depth_n.r_data[1][3] ));
Q_FDP4EP \depth_n.r_data_REG[1][2] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[2]), .Q(\depth_n.r_data[1][2] ));
Q_FDP4EP \depth_n.r_data_REG[1][1] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[1]), .Q(\depth_n.r_data[1][1] ));
Q_FDP4EP \depth_n.r_data_REG[1][0] ( .CK(clk), .CE(n10), .R(n1), .D(wdata[0]), .Q(\depth_n.r_data[1][0] ));
Q_FDP4EP \depth_n.r_data_REG[0][127] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[127]), .Q(\depth_n.r_data[0][127] ));
Q_FDP4EP \depth_n.r_data_REG[0][126] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[126]), .Q(\depth_n.r_data[0][126] ));
Q_FDP4EP \depth_n.r_data_REG[0][125] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[125]), .Q(\depth_n.r_data[0][125] ));
Q_FDP4EP \depth_n.r_data_REG[0][124] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[124]), .Q(\depth_n.r_data[0][124] ));
Q_FDP4EP \depth_n.r_data_REG[0][123] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[123]), .Q(\depth_n.r_data[0][123] ));
Q_FDP4EP \depth_n.r_data_REG[0][122] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[122]), .Q(\depth_n.r_data[0][122] ));
Q_FDP4EP \depth_n.r_data_REG[0][121] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[121]), .Q(\depth_n.r_data[0][121] ));
Q_FDP4EP \depth_n.r_data_REG[0][120] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[120]), .Q(\depth_n.r_data[0][120] ));
Q_FDP4EP \depth_n.r_data_REG[0][119] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[119]), .Q(\depth_n.r_data[0][119] ));
Q_FDP4EP \depth_n.r_data_REG[0][118] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[118]), .Q(\depth_n.r_data[0][118] ));
Q_FDP4EP \depth_n.r_data_REG[0][117] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[117]), .Q(\depth_n.r_data[0][117] ));
Q_FDP4EP \depth_n.r_data_REG[0][116] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[116]), .Q(\depth_n.r_data[0][116] ));
Q_FDP4EP \depth_n.r_data_REG[0][115] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[115]), .Q(\depth_n.r_data[0][115] ));
Q_FDP4EP \depth_n.r_data_REG[0][114] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[114]), .Q(\depth_n.r_data[0][114] ));
Q_FDP4EP \depth_n.r_data_REG[0][113] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[113]), .Q(\depth_n.r_data[0][113] ));
Q_FDP4EP \depth_n.r_data_REG[0][112] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[112]), .Q(\depth_n.r_data[0][112] ));
Q_FDP4EP \depth_n.r_data_REG[0][111] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[111]), .Q(\depth_n.r_data[0][111] ));
Q_FDP4EP \depth_n.r_data_REG[0][110] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[110]), .Q(\depth_n.r_data[0][110] ));
Q_FDP4EP \depth_n.r_data_REG[0][109] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[109]), .Q(\depth_n.r_data[0][109] ));
Q_FDP4EP \depth_n.r_data_REG[0][108] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[108]), .Q(\depth_n.r_data[0][108] ));
Q_FDP4EP \depth_n.r_data_REG[0][107] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[107]), .Q(\depth_n.r_data[0][107] ));
Q_FDP4EP \depth_n.r_data_REG[0][106] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[106]), .Q(\depth_n.r_data[0][106] ));
Q_FDP4EP \depth_n.r_data_REG[0][105] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[105]), .Q(\depth_n.r_data[0][105] ));
Q_FDP4EP \depth_n.r_data_REG[0][104] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[104]), .Q(\depth_n.r_data[0][104] ));
Q_FDP4EP \depth_n.r_data_REG[0][103] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[103]), .Q(\depth_n.r_data[0][103] ));
Q_FDP4EP \depth_n.r_data_REG[0][102] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[102]), .Q(\depth_n.r_data[0][102] ));
Q_FDP4EP \depth_n.r_data_REG[0][101] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[101]), .Q(\depth_n.r_data[0][101] ));
Q_FDP4EP \depth_n.r_data_REG[0][100] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[100]), .Q(\depth_n.r_data[0][100] ));
Q_FDP4EP \depth_n.r_data_REG[0][99] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[99]), .Q(\depth_n.r_data[0][99] ));
Q_FDP4EP \depth_n.r_data_REG[0][98] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[98]), .Q(\depth_n.r_data[0][98] ));
Q_FDP4EP \depth_n.r_data_REG[0][97] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[97]), .Q(\depth_n.r_data[0][97] ));
Q_FDP4EP \depth_n.r_data_REG[0][96] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[96]), .Q(\depth_n.r_data[0][96] ));
Q_FDP4EP \depth_n.r_data_REG[0][95] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[95]), .Q(\depth_n.r_data[0][95] ));
Q_FDP4EP \depth_n.r_data_REG[0][94] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[94]), .Q(\depth_n.r_data[0][94] ));
Q_FDP4EP \depth_n.r_data_REG[0][93] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[93]), .Q(\depth_n.r_data[0][93] ));
Q_FDP4EP \depth_n.r_data_REG[0][92] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[92]), .Q(\depth_n.r_data[0][92] ));
Q_FDP4EP \depth_n.r_data_REG[0][91] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[91]), .Q(\depth_n.r_data[0][91] ));
Q_FDP4EP \depth_n.r_data_REG[0][90] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[90]), .Q(\depth_n.r_data[0][90] ));
Q_FDP4EP \depth_n.r_data_REG[0][89] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[89]), .Q(\depth_n.r_data[0][89] ));
Q_FDP4EP \depth_n.r_data_REG[0][88] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[88]), .Q(\depth_n.r_data[0][88] ));
Q_FDP4EP \depth_n.r_data_REG[0][87] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[87]), .Q(\depth_n.r_data[0][87] ));
Q_FDP4EP \depth_n.r_data_REG[0][86] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[86]), .Q(\depth_n.r_data[0][86] ));
Q_FDP4EP \depth_n.r_data_REG[0][85] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[85]), .Q(\depth_n.r_data[0][85] ));
Q_FDP4EP \depth_n.r_data_REG[0][84] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[84]), .Q(\depth_n.r_data[0][84] ));
Q_FDP4EP \depth_n.r_data_REG[0][83] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[83]), .Q(\depth_n.r_data[0][83] ));
Q_FDP4EP \depth_n.r_data_REG[0][82] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[82]), .Q(\depth_n.r_data[0][82] ));
Q_FDP4EP \depth_n.r_data_REG[0][81] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[81]), .Q(\depth_n.r_data[0][81] ));
Q_FDP4EP \depth_n.r_data_REG[0][80] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[80]), .Q(\depth_n.r_data[0][80] ));
Q_FDP4EP \depth_n.r_data_REG[0][79] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[79]), .Q(\depth_n.r_data[0][79] ));
Q_FDP4EP \depth_n.r_data_REG[0][78] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[78]), .Q(\depth_n.r_data[0][78] ));
Q_FDP4EP \depth_n.r_data_REG[0][77] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[77]), .Q(\depth_n.r_data[0][77] ));
Q_FDP4EP \depth_n.r_data_REG[0][76] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[76]), .Q(\depth_n.r_data[0][76] ));
Q_FDP4EP \depth_n.r_data_REG[0][75] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[75]), .Q(\depth_n.r_data[0][75] ));
Q_FDP4EP \depth_n.r_data_REG[0][74] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[74]), .Q(\depth_n.r_data[0][74] ));
Q_FDP4EP \depth_n.r_data_REG[0][73] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[73]), .Q(\depth_n.r_data[0][73] ));
Q_FDP4EP \depth_n.r_data_REG[0][72] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[72]), .Q(\depth_n.r_data[0][72] ));
Q_FDP4EP \depth_n.r_data_REG[0][71] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[71]), .Q(\depth_n.r_data[0][71] ));
Q_FDP4EP \depth_n.r_data_REG[0][70] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[70]), .Q(\depth_n.r_data[0][70] ));
Q_FDP4EP \depth_n.r_data_REG[0][69] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[69]), .Q(\depth_n.r_data[0][69] ));
Q_FDP4EP \depth_n.r_data_REG[0][68] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[68]), .Q(\depth_n.r_data[0][68] ));
Q_FDP4EP \depth_n.r_data_REG[0][67] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[67]), .Q(\depth_n.r_data[0][67] ));
Q_FDP4EP \depth_n.r_data_REG[0][66] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[66]), .Q(\depth_n.r_data[0][66] ));
Q_FDP4EP \depth_n.r_data_REG[0][65] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[65]), .Q(\depth_n.r_data[0][65] ));
Q_FDP4EP \depth_n.r_data_REG[0][64] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[64]), .Q(\depth_n.r_data[0][64] ));
Q_FDP4EP \depth_n.r_data_REG[0][63] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[63]), .Q(\depth_n.r_data[0][63] ));
Q_FDP4EP \depth_n.r_data_REG[0][62] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[62]), .Q(\depth_n.r_data[0][62] ));
Q_FDP4EP \depth_n.r_data_REG[0][61] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[61]), .Q(\depth_n.r_data[0][61] ));
Q_FDP4EP \depth_n.r_data_REG[0][60] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[60]), .Q(\depth_n.r_data[0][60] ));
Q_FDP4EP \depth_n.r_data_REG[0][59] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[59]), .Q(\depth_n.r_data[0][59] ));
Q_FDP4EP \depth_n.r_data_REG[0][58] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[58]), .Q(\depth_n.r_data[0][58] ));
Q_FDP4EP \depth_n.r_data_REG[0][57] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[57]), .Q(\depth_n.r_data[0][57] ));
Q_FDP4EP \depth_n.r_data_REG[0][56] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[56]), .Q(\depth_n.r_data[0][56] ));
Q_FDP4EP \depth_n.r_data_REG[0][55] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[55]), .Q(\depth_n.r_data[0][55] ));
Q_FDP4EP \depth_n.r_data_REG[0][54] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[54]), .Q(\depth_n.r_data[0][54] ));
Q_FDP4EP \depth_n.r_data_REG[0][53] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[53]), .Q(\depth_n.r_data[0][53] ));
Q_FDP4EP \depth_n.r_data_REG[0][52] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[52]), .Q(\depth_n.r_data[0][52] ));
Q_FDP4EP \depth_n.r_data_REG[0][51] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[51]), .Q(\depth_n.r_data[0][51] ));
Q_FDP4EP \depth_n.r_data_REG[0][50] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[50]), .Q(\depth_n.r_data[0][50] ));
Q_FDP4EP \depth_n.r_data_REG[0][49] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[49]), .Q(\depth_n.r_data[0][49] ));
Q_FDP4EP \depth_n.r_data_REG[0][48] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[48]), .Q(\depth_n.r_data[0][48] ));
Q_FDP4EP \depth_n.r_data_REG[0][47] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[47]), .Q(\depth_n.r_data[0][47] ));
Q_FDP4EP \depth_n.r_data_REG[0][46] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[46]), .Q(\depth_n.r_data[0][46] ));
Q_FDP4EP \depth_n.r_data_REG[0][45] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[45]), .Q(\depth_n.r_data[0][45] ));
Q_FDP4EP \depth_n.r_data_REG[0][44] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[44]), .Q(\depth_n.r_data[0][44] ));
Q_FDP4EP \depth_n.r_data_REG[0][43] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[43]), .Q(\depth_n.r_data[0][43] ));
Q_FDP4EP \depth_n.r_data_REG[0][42] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[42]), .Q(\depth_n.r_data[0][42] ));
Q_FDP4EP \depth_n.r_data_REG[0][41] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[41]), .Q(\depth_n.r_data[0][41] ));
Q_FDP4EP \depth_n.r_data_REG[0][40] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[40]), .Q(\depth_n.r_data[0][40] ));
Q_FDP4EP \depth_n.r_data_REG[0][39] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[39]), .Q(\depth_n.r_data[0][39] ));
Q_FDP4EP \depth_n.r_data_REG[0][38] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[38]), .Q(\depth_n.r_data[0][38] ));
Q_FDP4EP \depth_n.r_data_REG[0][37] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[37]), .Q(\depth_n.r_data[0][37] ));
Q_FDP4EP \depth_n.r_data_REG[0][36] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[36]), .Q(\depth_n.r_data[0][36] ));
Q_FDP4EP \depth_n.r_data_REG[0][35] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[35]), .Q(\depth_n.r_data[0][35] ));
Q_FDP4EP \depth_n.r_data_REG[0][34] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[34]), .Q(\depth_n.r_data[0][34] ));
Q_FDP4EP \depth_n.r_data_REG[0][33] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[33]), .Q(\depth_n.r_data[0][33] ));
Q_FDP4EP \depth_n.r_data_REG[0][32] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[32]), .Q(\depth_n.r_data[0][32] ));
Q_FDP4EP \depth_n.r_data_REG[0][31] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[31]), .Q(\depth_n.r_data[0][31] ));
Q_FDP4EP \depth_n.r_data_REG[0][30] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[30]), .Q(\depth_n.r_data[0][30] ));
Q_FDP4EP \depth_n.r_data_REG[0][29] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[29]), .Q(\depth_n.r_data[0][29] ));
Q_FDP4EP \depth_n.r_data_REG[0][28] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[28]), .Q(\depth_n.r_data[0][28] ));
Q_FDP4EP \depth_n.r_data_REG[0][27] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[27]), .Q(\depth_n.r_data[0][27] ));
Q_FDP4EP \depth_n.r_data_REG[0][26] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[26]), .Q(\depth_n.r_data[0][26] ));
Q_FDP4EP \depth_n.r_data_REG[0][25] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[25]), .Q(\depth_n.r_data[0][25] ));
Q_FDP4EP \depth_n.r_data_REG[0][24] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[24]), .Q(\depth_n.r_data[0][24] ));
Q_FDP4EP \depth_n.r_data_REG[0][23] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[23]), .Q(\depth_n.r_data[0][23] ));
Q_FDP4EP \depth_n.r_data_REG[0][22] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[22]), .Q(\depth_n.r_data[0][22] ));
Q_FDP4EP \depth_n.r_data_REG[0][21] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[21]), .Q(\depth_n.r_data[0][21] ));
Q_FDP4EP \depth_n.r_data_REG[0][20] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[20]), .Q(\depth_n.r_data[0][20] ));
Q_FDP4EP \depth_n.r_data_REG[0][19] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[19]), .Q(\depth_n.r_data[0][19] ));
Q_FDP4EP \depth_n.r_data_REG[0][18] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[18]), .Q(\depth_n.r_data[0][18] ));
Q_FDP4EP \depth_n.r_data_REG[0][17] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[17]), .Q(\depth_n.r_data[0][17] ));
Q_FDP4EP \depth_n.r_data_REG[0][16] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[16]), .Q(\depth_n.r_data[0][16] ));
Q_FDP4EP \depth_n.r_data_REG[0][15] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[15]), .Q(\depth_n.r_data[0][15] ));
Q_FDP4EP \depth_n.r_data_REG[0][14] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[14]), .Q(\depth_n.r_data[0][14] ));
Q_FDP4EP \depth_n.r_data_REG[0][13] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[13]), .Q(\depth_n.r_data[0][13] ));
Q_FDP4EP \depth_n.r_data_REG[0][12] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[12]), .Q(\depth_n.r_data[0][12] ));
Q_FDP4EP \depth_n.r_data_REG[0][11] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[11]), .Q(\depth_n.r_data[0][11] ));
Q_FDP4EP \depth_n.r_data_REG[0][10] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[10]), .Q(\depth_n.r_data[0][10] ));
Q_FDP4EP \depth_n.r_data_REG[0][9] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[9]), .Q(\depth_n.r_data[0][9] ));
Q_FDP4EP \depth_n.r_data_REG[0][8] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[8]), .Q(\depth_n.r_data[0][8] ));
Q_FDP4EP \depth_n.r_data_REG[0][7] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[7]), .Q(\depth_n.r_data[0][7] ));
Q_FDP4EP \depth_n.r_data_REG[0][6] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[6]), .Q(\depth_n.r_data[0][6] ));
Q_FDP4EP \depth_n.r_data_REG[0][5] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[5]), .Q(\depth_n.r_data[0][5] ));
Q_FDP4EP \depth_n.r_data_REG[0][4] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[4]), .Q(\depth_n.r_data[0][4] ));
Q_FDP4EP \depth_n.r_data_REG[0][3] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[3]), .Q(\depth_n.r_data[0][3] ));
Q_FDP4EP \depth_n.r_data_REG[0][2] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[2]), .Q(\depth_n.r_data[0][2] ));
Q_FDP4EP \depth_n.r_data_REG[0][1] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[1]), .Q(\depth_n.r_data[0][1] ));
Q_FDP4EP \depth_n.r_data_REG[0][0] ( .CK(clk), .CE(n12), .R(n1), .D(wdata[0]), .Q(\depth_n.r_data[0][0] ));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "\depth_n.r_data  1 127 0 2 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 depth_n  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n.genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n"
endmodule
