
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_fifo_xcm21 ( empty, full, underflow, overflow, used_slots, free_slots, 
	rdata, clk, rst_n, wen, ren, clear, wdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output empty;
output full;
output underflow;
output overflow;
output [4:0] used_slots;
output [4:0] free_slots;
output [63:0] rdata;
input clk;
input rst_n;
input wen;
input ren;
input clear;
input [63:0] wdata;
wire _zy_simnet_underflow_0_w$;
wire _zy_simnet_overflow_1_w$;
wire \depth_n._zy_simnet_overflow_3_w$ ;
wire \depth_n._zy_simnet_underflow_2_w$ ;
wire [3:0] \depth_n.wptr ;
wire [3:0] \depth_n.rptr ;
supply0 n143;
ixc_assign _zz_strnp_3 ( _zy_simnet_overflow_1_w$, overflow);
ixc_assign _zz_strnp_2 ( _zy_simnet_underflow_0_w$, underflow);
Q_FDP0 U2 ( .CK(clk), .D(wdata[63]), .Q(n142), .QN( ));
Q_FDP0 U3 ( .CK(clk), .D(wdata[62]), .Q(n141), .QN( ));
Q_FDP0 U4 ( .CK(clk), .D(wdata[61]), .Q(n140), .QN( ));
Q_FDP0 U5 ( .CK(clk), .D(wdata[60]), .Q(n139), .QN( ));
Q_FDP0 U6 ( .CK(clk), .D(wdata[59]), .Q(n138), .QN( ));
Q_FDP0 U7 ( .CK(clk), .D(wdata[58]), .Q(n137), .QN( ));
Q_FDP0 U8 ( .CK(clk), .D(wdata[57]), .Q(n136), .QN( ));
Q_FDP0 U9 ( .CK(clk), .D(wdata[56]), .Q(n135), .QN( ));
Q_FDP0 U10 ( .CK(clk), .D(wdata[55]), .Q(n134), .QN( ));
Q_FDP0 U11 ( .CK(clk), .D(wdata[54]), .Q(n133), .QN( ));
Q_FDP0 U12 ( .CK(clk), .D(wdata[53]), .Q(n132), .QN( ));
Q_FDP0 U13 ( .CK(clk), .D(wdata[52]), .Q(n131), .QN( ));
Q_FDP0 U14 ( .CK(clk), .D(wdata[51]), .Q(n130), .QN( ));
Q_FDP0 U15 ( .CK(clk), .D(wdata[50]), .Q(n129), .QN( ));
Q_FDP0 U16 ( .CK(clk), .D(wdata[49]), .Q(n128), .QN( ));
Q_FDP0 U17 ( .CK(clk), .D(wdata[48]), .Q(n127), .QN( ));
Q_FDP0 U18 ( .CK(clk), .D(wdata[47]), .Q(n126), .QN( ));
Q_FDP0 U19 ( .CK(clk), .D(wdata[46]), .Q(n125), .QN( ));
Q_FDP0 U20 ( .CK(clk), .D(wdata[45]), .Q(n124), .QN( ));
Q_FDP0 U21 ( .CK(clk), .D(wdata[44]), .Q(n123), .QN( ));
Q_FDP0 U22 ( .CK(clk), .D(wdata[43]), .Q(n122), .QN( ));
Q_FDP0 U23 ( .CK(clk), .D(wdata[42]), .Q(n121), .QN( ));
Q_FDP0 U24 ( .CK(clk), .D(wdata[41]), .Q(n120), .QN( ));
Q_FDP0 U25 ( .CK(clk), .D(wdata[40]), .Q(n119), .QN( ));
Q_FDP0 U26 ( .CK(clk), .D(wdata[39]), .Q(n118), .QN( ));
Q_FDP0 U27 ( .CK(clk), .D(wdata[38]), .Q(n117), .QN( ));
Q_FDP0 U28 ( .CK(clk), .D(wdata[37]), .Q(n116), .QN( ));
Q_FDP0 U29 ( .CK(clk), .D(wdata[36]), .Q(n115), .QN( ));
Q_FDP0 U30 ( .CK(clk), .D(wdata[35]), .Q(n114), .QN( ));
Q_FDP0 U31 ( .CK(clk), .D(wdata[34]), .Q(n113), .QN( ));
Q_FDP0 U32 ( .CK(clk), .D(wdata[33]), .Q(n112), .QN( ));
Q_FDP0 U33 ( .CK(clk), .D(wdata[32]), .Q(n111), .QN( ));
Q_FDP0 U34 ( .CK(clk), .D(wdata[31]), .Q(n110), .QN( ));
Q_FDP0 U35 ( .CK(clk), .D(wdata[30]), .Q(n109), .QN( ));
Q_FDP0 U36 ( .CK(clk), .D(wdata[29]), .Q(n108), .QN( ));
Q_FDP0 U37 ( .CK(clk), .D(wdata[28]), .Q(n107), .QN( ));
Q_FDP0 U38 ( .CK(clk), .D(wdata[27]), .Q(n106), .QN( ));
Q_FDP0 U39 ( .CK(clk), .D(wdata[26]), .Q(n105), .QN( ));
Q_FDP0 U40 ( .CK(clk), .D(wdata[25]), .Q(n104), .QN( ));
Q_FDP0 U41 ( .CK(clk), .D(wdata[24]), .Q(n103), .QN( ));
Q_FDP0 U42 ( .CK(clk), .D(wdata[23]), .Q(n102), .QN( ));
Q_FDP0 U43 ( .CK(clk), .D(wdata[22]), .Q(n101), .QN( ));
Q_FDP0 U44 ( .CK(clk), .D(wdata[21]), .Q(n100), .QN( ));
Q_FDP0 U45 ( .CK(clk), .D(wdata[20]), .Q(n99), .QN( ));
Q_FDP0 U46 ( .CK(clk), .D(wdata[19]), .Q(n98), .QN( ));
Q_FDP0 U47 ( .CK(clk), .D(wdata[18]), .Q(n97), .QN( ));
Q_FDP0 U48 ( .CK(clk), .D(wdata[17]), .Q(n96), .QN( ));
Q_FDP0 U49 ( .CK(clk), .D(wdata[16]), .Q(n95), .QN( ));
Q_FDP0 U50 ( .CK(clk), .D(wdata[15]), .Q(n94), .QN( ));
Q_FDP0 U51 ( .CK(clk), .D(wdata[14]), .Q(n93), .QN( ));
Q_FDP0 U52 ( .CK(clk), .D(wdata[13]), .Q(n92), .QN( ));
Q_FDP0 U53 ( .CK(clk), .D(wdata[12]), .Q(n91), .QN( ));
Q_FDP0 U54 ( .CK(clk), .D(wdata[11]), .Q(n90), .QN( ));
Q_FDP0 U55 ( .CK(clk), .D(wdata[10]), .Q(n89), .QN( ));
Q_FDP0 U56 ( .CK(clk), .D(wdata[9]), .Q(n88), .QN( ));
Q_FDP0 U57 ( .CK(clk), .D(wdata[8]), .Q(n87), .QN( ));
Q_FDP0 U58 ( .CK(clk), .D(wdata[7]), .Q(n86), .QN( ));
Q_FDP0 U59 ( .CK(clk), .D(wdata[6]), .Q(n85), .QN( ));
Q_FDP0 U60 ( .CK(clk), .D(wdata[5]), .Q(n84), .QN( ));
Q_FDP0 U61 ( .CK(clk), .D(wdata[4]), .Q(n83), .QN( ));
Q_FDP0 U62 ( .CK(clk), .D(wdata[3]), .Q(n82), .QN( ));
Q_FDP0 U63 ( .CK(clk), .D(wdata[2]), .Q(n81), .QN( ));
Q_FDP0 U64 ( .CK(clk), .D(wdata[1]), .Q(n80), .QN( ));
Q_FDP0 U65 ( .CK(clk), .D(wdata[0]), .Q(n79), .QN( ));
Q_FDP0 U66 ( .CK(clk), .D(\depth_n.wptr [3]), .Q(n78), .QN( ));
Q_FDP0 U67 ( .CK(clk), .D(\depth_n.wptr [2]), .Q(n77), .QN( ));
Q_FDP0 U68 ( .CK(clk), .D(\depth_n.wptr [1]), .Q(n76), .QN( ));
Q_FDP0 U69 ( .CK(clk), .D(\depth_n.wptr [0]), .Q(n75), .QN( ));
Q_AN02 U70 ( .A0(n70), .A1(n73), .Z(n74));
Q_XOR2 U71 ( .A0(n69), .A1(n72), .Z(n73));
// pragma CVAINTPROP NET n69 _2_state_ 1
// pragma CVAINTPROP INSTANCE U71 NOBREAKS 1
Q_FDP0B U72 ( .D(n69), .QTFCLK( ), .Q(n72));
Q_FDP0 U73 ( .CK(clk), .D(n3), .Q(n70), .QN( ));
Q_FDP0 U74 ( .CK(clk), .D(n71), .Q(n69), .QN(n71));
Q_INV U75 ( .A(empty), .Z(n68));
Q_AN02 U76 ( .A0(n68), .A1(n4), .Z(rdata[63]));
Q_AN02 U77 ( .A0(n68), .A1(n5), .Z(rdata[62]));
Q_AN02 U78 ( .A0(n68), .A1(n6), .Z(rdata[61]));
Q_AN02 U79 ( .A0(n68), .A1(n7), .Z(rdata[60]));
Q_AN02 U80 ( .A0(n68), .A1(n8), .Z(rdata[59]));
Q_AN02 U81 ( .A0(n68), .A1(n9), .Z(rdata[58]));
Q_AN02 U82 ( .A0(n68), .A1(n10), .Z(rdata[57]));
Q_AN02 U83 ( .A0(n68), .A1(n11), .Z(rdata[56]));
Q_AN02 U84 ( .A0(n68), .A1(n12), .Z(rdata[55]));
Q_AN02 U85 ( .A0(n68), .A1(n13), .Z(rdata[54]));
Q_AN02 U86 ( .A0(n68), .A1(n14), .Z(rdata[53]));
Q_AN02 U87 ( .A0(n68), .A1(n15), .Z(rdata[52]));
Q_AN02 U88 ( .A0(n68), .A1(n16), .Z(rdata[51]));
Q_AN02 U89 ( .A0(n68), .A1(n17), .Z(rdata[50]));
Q_AN02 U90 ( .A0(n68), .A1(n18), .Z(rdata[49]));
Q_AN02 U91 ( .A0(n68), .A1(n19), .Z(rdata[48]));
Q_AN02 U92 ( .A0(n68), .A1(n20), .Z(rdata[47]));
Q_AN02 U93 ( .A0(n68), .A1(n21), .Z(rdata[46]));
Q_AN02 U94 ( .A0(n68), .A1(n22), .Z(rdata[45]));
Q_AN02 U95 ( .A0(n68), .A1(n23), .Z(rdata[44]));
Q_AN02 U96 ( .A0(n68), .A1(n24), .Z(rdata[43]));
Q_AN02 U97 ( .A0(n68), .A1(n25), .Z(rdata[42]));
Q_AN02 U98 ( .A0(n68), .A1(n26), .Z(rdata[41]));
Q_AN02 U99 ( .A0(n68), .A1(n27), .Z(rdata[40]));
Q_AN02 U100 ( .A0(n68), .A1(n28), .Z(rdata[39]));
Q_AN02 U101 ( .A0(n68), .A1(n29), .Z(rdata[38]));
Q_AN02 U102 ( .A0(n68), .A1(n30), .Z(rdata[37]));
Q_AN02 U103 ( .A0(n68), .A1(n31), .Z(rdata[36]));
Q_AN02 U104 ( .A0(n68), .A1(n32), .Z(rdata[35]));
Q_AN02 U105 ( .A0(n68), .A1(n33), .Z(rdata[34]));
Q_AN02 U106 ( .A0(n68), .A1(n34), .Z(rdata[33]));
Q_AN02 U107 ( .A0(n68), .A1(n35), .Z(rdata[32]));
Q_AN02 U108 ( .A0(n68), .A1(n36), .Z(rdata[31]));
Q_AN02 U109 ( .A0(n68), .A1(n37), .Z(rdata[30]));
Q_AN02 U110 ( .A0(n68), .A1(n38), .Z(rdata[29]));
Q_AN02 U111 ( .A0(n68), .A1(n39), .Z(rdata[28]));
Q_AN02 U112 ( .A0(n68), .A1(n40), .Z(rdata[27]));
Q_AN02 U113 ( .A0(n68), .A1(n41), .Z(rdata[26]));
Q_AN02 U114 ( .A0(n68), .A1(n42), .Z(rdata[25]));
Q_AN02 U115 ( .A0(n68), .A1(n43), .Z(rdata[24]));
Q_AN02 U116 ( .A0(n68), .A1(n44), .Z(rdata[23]));
Q_AN02 U117 ( .A0(n68), .A1(n45), .Z(rdata[22]));
Q_AN02 U118 ( .A0(n68), .A1(n46), .Z(rdata[21]));
Q_AN02 U119 ( .A0(n68), .A1(n47), .Z(rdata[20]));
Q_AN02 U120 ( .A0(n68), .A1(n48), .Z(rdata[19]));
Q_AN02 U121 ( .A0(n68), .A1(n49), .Z(rdata[18]));
Q_AN02 U122 ( .A0(n68), .A1(n50), .Z(rdata[17]));
Q_AN02 U123 ( .A0(n68), .A1(n51), .Z(rdata[16]));
Q_AN02 U124 ( .A0(n68), .A1(n52), .Z(rdata[15]));
Q_AN02 U125 ( .A0(n68), .A1(n53), .Z(rdata[14]));
Q_AN02 U126 ( .A0(n68), .A1(n54), .Z(rdata[13]));
Q_AN02 U127 ( .A0(n68), .A1(n55), .Z(rdata[12]));
Q_AN02 U128 ( .A0(n68), .A1(n56), .Z(rdata[11]));
Q_AN02 U129 ( .A0(n68), .A1(n57), .Z(rdata[10]));
Q_AN02 U130 ( .A0(n68), .A1(n58), .Z(rdata[9]));
Q_AN02 U131 ( .A0(n68), .A1(n59), .Z(rdata[8]));
Q_AN02 U132 ( .A0(n68), .A1(n60), .Z(rdata[7]));
Q_AN02 U133 ( .A0(n68), .A1(n61), .Z(rdata[6]));
Q_AN02 U134 ( .A0(n68), .A1(n62), .Z(rdata[5]));
Q_AN02 U135 ( .A0(n68), .A1(n63), .Z(rdata[4]));
Q_AN02 U136 ( .A0(n68), .A1(n64), .Z(rdata[3]));
Q_AN02 U137 ( .A0(n68), .A1(n65), .Z(rdata[2]));
Q_AN02 U138 ( .A0(n68), .A1(n66), .Z(rdata[1]));
Q_AN02 U139 ( .A0(n68), .A1(n67), .Z(rdata[0]));
Q_INV U140 ( .A(full), .Z(n2));
Q_AN02 U141 ( .A0(wen), .A1(n2), .Z(n3));
nx_fifo_ctrl_xcm37 \depth_n.fifo_ctrl ( .empty( empty), .full( full), 
	.used_slots( used_slots[4:0]), .free_slots( free_slots[4:0]), 
	.rptr( \depth_n.rptr [3:0]), .wptr( \depth_n.wptr [3:0]), 
	.underflow( \depth_n._zy_simnet_underflow_2_w$ ), .overflow( 
	\depth_n._zy_simnet_overflow_3_w$ ), .clk( clk), .rst_n( rst_n), 
	.wen( wen), .ren( ren), .clear( clear));
ixc_assign \depth_n._zz_strnp_1 ( overflow, 
	\depth_n._zy_simnet_overflow_3_w$ );
ixc_assign \depth_n._zz_strnp_0 ( underflow, 
	\depth_n._zy_simnet_underflow_2_w$ );
`ifdef CBV

reg [63:0] \depth_n.r_data  [15:0];
initial begin: U145
  integer i;
  for (i=15; i>=0; i=i-1) \depth_n.r_data [i] =
`ifdef CBV_MEM_INIT1
  {64{1'b1}};
`else
  64'b0;
`endif
end
reg [63:0] n144;
assign {n4, n5, n6, n7, n8, n9, n10,
n11, n12, n13, n14, n15, n16, n17, n18,
n19, n20, n21, n22, n23, n24, n25, n26,
n27, n28, n29, n30, n31, n32, n33, n34,
n35, n36, n37, n38, n39, n40, n41, n42,
n43, n44, n45, n46, n47, n48, n49, n50,
n51, n52, n53, n54, n55, n56, n57, n58,
n59, n60, n61, n62, n63, n64, n65, n66,
n67} = n144; 
always @(n78 or n77 or n76 or n75 or n142
 or n141 or n140 or n139 or n138 or n137 or n136 or n135 or n134
 or n133 or n132 or n131 or n130 or n129 or n128 or n127 or n126
 or n125 or n124 or n123 or n122 or n121 or n120 or n119 or n118
 or n117 or n116 or n115 or n114 or n113 or n112 or n111 or n110
 or n109 or n108 or n107 or n106 or n105 or n104 or n103 or n102
 or n101 or n100 or n99 or n98 or n97 or n96 or n95 or n94
 or n93 or n92 or n91 or n90 or n89 or n88 or n87 or n86
 or n85 or n84 or n83 or n82 or n81 or n80 or n79 or n74
 or \depth_n.rptr [3] or \depth_n.rptr [2] or \depth_n.rptr [1] or \depth_n.rptr [0])
#0 begin
if (n74)
\depth_n.r_data [{n78, n77, n76, n75}] =
{n142, n141, n140, n139, n138,
 n137, n136, n135, n134, n133, n132, n131, n130,
 n129, n128, n127, n126, n125, n124, n123, n122,
 n121, n120, n119, n118, n117, n116, n115, n114,
 n113, n112, n111, n110, n109, n108, n107, n106,
 n105, n104, n103, n102, n101, n100, n99, n98,
 n97, n96, n95, n94, n93, n92, n91, n90,
 n89, n88, n87, n86, n85, n84, n83, n82,
 n81, n80, n79};
n144 = \depth_n.r_data [{\depth_n.rptr [3], \depth_n.rptr [2], \depth_n.rptr [1], \depth_n.rptr [0]}];
end
`else

MPW16X64 \depth_n.r_data  ( .A3(n78), .A2(n77), .A1(n76), .A0(n75), .DI63(n142), .DI62(n141),
 .DI61(n140), .DI60(n139), .DI59(n138), .DI58(n137), .DI57(n136), .DI56(n135), .DI55(n134), .DI54(n133),
 .DI53(n132), .DI52(n131), .DI51(n130), .DI50(n129), .DI49(n128), .DI48(n127), .DI47(n126), .DI46(n125),
 .DI45(n124), .DI44(n123), .DI43(n122), .DI42(n121), .DI41(n120), .DI40(n119), .DI39(n118), .DI38(n117),
 .DI37(n116), .DI36(n115), .DI35(n114), .DI34(n113), .DI33(n112), .DI32(n111), .DI31(n110), .DI30(n109),
 .DI29(n108), .DI28(n107), .DI27(n106), .DI26(n105), .DI25(n104), .DI24(n103), .DI23(n102), .DI22(n101),
 .DI21(n100), .DI20(n99), .DI19(n98), .DI18(n97), .DI17(n96), .DI16(n95), .DI15(n94), .DI14(n93),
 .DI13(n92), .DI12(n91), .DI11(n90), .DI10(n89), .DI9(n88), .DI8(n87), .DI7(n86), .DI6(n85),
 .DI5(n84), .DI4(n83), .DI3(n82), .DI2(n81), .DI1(n80), .DI0(n79), .WE(n74), .SYNC_IN(n143),
 .SYNC_OUT(n144));
// pragma CVASTRPROP INSTANCE "\depth_n.r_data " HDL_MEMORY_DECL "1 63 0 15 0"
MPR16X64 U146 ( .A3(\depth_n.rptr [3]), .A2(\depth_n.rptr [2]), .A1(\depth_n.rptr [1]), .A0(\depth_n.rptr [0]), .SYNC_IN(n144), .DO63(n4),
 .DO62(n5), .DO61(n6), .DO60(n7), .DO59(n8), .DO58(n9), .DO57(n10), .DO56(n11), .DO55(n12),
 .DO54(n13), .DO53(n14), .DO52(n15), .DO51(n16), .DO50(n17), .DO49(n18), .DO48(n19), .DO47(n20),
 .DO46(n21), .DO45(n22), .DO44(n23), .DO43(n24), .DO42(n25), .DO41(n26), .DO40(n27), .DO39(n28),
 .DO38(n29), .DO37(n30), .DO36(n31), .DO35(n32), .DO34(n33), .DO33(n34), .DO32(n35), .DO31(n36),
 .DO30(n37), .DO29(n38), .DO28(n39), .DO27(n40), .DO26(n41), .DO25(n42), .DO24(n43), .DO23(n44),
 .DO22(n45), .DO21(n46), .DO20(n47), .DO19(n48), .DO18(n49), .DO17(n50), .DO16(n51), .DO15(n52),
 .DO14(n53), .DO13(n54), .DO12(n55), .DO11(n56), .DO10(n57), .DO9(n58), .DO8(n59), .DO7(n60),
 .DO6(n61), .DO5(n62), .DO4(n63), .DO3(n64), .DO2(n65), .DO1(n66), .DO0(n67), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\depth_n.r_data  1 63 0 15 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 depth_n  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n.genblk1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "depth_n"
endmodule
`ifdef CBV
`else
`ifdef MPW16X64_MPR16X64
`else
module MPW16X64( A3, A2, A1, A0, DI63, DI62, DI61,
 DI60, DI59, DI58, DI57, DI56, DI55, DI54, DI53,
 DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45,
 DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37,
 DI36, DI35, DI34, DI33, DI32, DI31, DI30, DI29,
 DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21,
 DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5,
 DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A3, A2, A1, A0, DI63, DI62, DI61, DI60,
 DI59, DI58, DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32, DI31, DI30,
 DI29, DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21, DI20,
 DI19, DI18, DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR16X64_
`else
module MPR16X64( A3, A2, A1, A0, SYNC_IN, DO63, DO62,
 DO61, DO60, DO59, DO58, DO57, DO56, DO55, DO54,
 DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30,
 DO29, DO28, DO27, DO26, DO25, DO24, DO23, DO22,
 DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT);
input  A3, A2, A1, A0, SYNC_IN;
output  DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56,
 DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26,
 DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16,
 DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR16X64_
`endif
`define MPW16X64_MPR16X64
`endif
`endif
