
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module IXC_SV_SFIFO_VXE_256 ( rdCnt, scgGFreq);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
`_2_ output [63:0] rdCnt;
input scgGFreq;
wire fclk;
wire [0:63] _zy_simnet_rdCnt_0_w$;
`_2_ wire [21:0] tId;
`_2_ wire [511:0] iData;
`_2_ wire [16:0] wptr;
`_2_ wire [16:0] wptrN;
`_2_ wire [16:0] xptr;
`_2_ wire [16:0] xptrN;
`_2_ wire [255:0] ififoXdata;
`_2_ wire [255:0] ififoXdataFinal;
`_2_ wire [16:0] rptr;
`_2_ wire [16:0] rptrN;
`_2_ wire [14:0] ififoRaddr0;
`_2_ wire [14:0] ififoRaddr1;
`_2_ wire [14:0] ififoRaddr2;
`_2_ wire [767:0] ififoRdata;
`_2_ wire [17:0] rdDelta;
`_2_ wire [3:0] markBits;
`_2_ wire [3:0] markBitsN;
`_2_ wire [3:0] newMarkBits;
`_2_ wire [3:0] newMarkBitsD;
`_2_ wire [3:0] dataBits;
`_2_ wire [23:0] offset;
`_2_ wire [23:0] offsetN;
`_2_ wire moveForward;
`_2_ wire moveForwardN;
`_2_ wire active;
`_2_ wire activeD;
`_2_ wire [63:0] xval;
`_2_ wire nps;
`_2_ wire eob;
`_2_ wire [31:0] i;
`_2_ wire [63:0] head;
`_2_ wire [63:0] xhead;
`_2_ wire [63:0] vhead;
`_2_ wire [15:0] pktl;
`_2_ wire [15:0] pktlN;
`_2_ wire [9:0] vlen;
`_2_ wire [9:0] vlenN;
`_2_ wire rstDone;
`_2_ wire rstDoneD;
`_2_ wire rstDoneD2;
`_2_ wire [11:0] odly;
`_2_ wire [11:0] odlyN;
`_2_ wire vmode;
`_2_ wire [575:0] tmpData;
wire oSt;
`_2_ wire [255:0] oMark;
`_2_ wire oDataEn;
`_2_ wire [3:0] oDataLen;
`_2_ wire [511:0] oData;
`_2_ wire [31:0] numRsts;
`_2_ wire [767:0] ofifoData;
`_2_ wire [3:0] oFill;
`_2_ wire [14:0] ofifoAddr0;
`_2_ wire [15:0] ofifoAddr1;
`_2_ wire [15:0] ofifoAddr2;
`_2_ wire [14:0] ofifoWptr;
`_2_ wire [7:0] shiftCount;
`_2_ wire [767:0] shiftedOData;
supply0 n5631;
supply1 n6882;
Q_BUF U0 ( .A(n6882), .Z(xc_top.hasSFIFO));
Q_BUF U1 ( .A(ififoXdata[255]), .Z(newMarkBits[3]));
Q_BUF U2 ( .A(ififoXdata[191]), .Z(newMarkBits[2]));
Q_BUF U3 ( .A(ififoXdata[127]), .Z(newMarkBits[1]));
Q_BUF U4 ( .A(ififoXdata[63]), .Z(newMarkBits[0]));
Q_BUF U5 ( .A(dataBits[3]), .Z(xval[35]));
Q_BUF U6 ( .A(dataBits[2]), .Z(xval[34]));
Q_BUF U7 ( .A(dataBits[1]), .Z(xval[33]));
Q_BUF U8 ( .A(dataBits[0]), .Z(xval[32]));
Q_BUF U9 ( .A(iData[511]), .Z(tmpData[575]));
Q_BUF U10 ( .A(iData[510]), .Z(tmpData[574]));
Q_BUF U11 ( .A(iData[509]), .Z(tmpData[573]));
Q_BUF U12 ( .A(iData[508]), .Z(tmpData[572]));
Q_BUF U13 ( .A(iData[507]), .Z(tmpData[571]));
Q_BUF U14 ( .A(iData[506]), .Z(tmpData[570]));
Q_BUF U15 ( .A(iData[505]), .Z(tmpData[569]));
Q_BUF U16 ( .A(iData[504]), .Z(tmpData[568]));
Q_BUF U17 ( .A(iData[503]), .Z(tmpData[567]));
Q_BUF U18 ( .A(iData[502]), .Z(tmpData[566]));
Q_BUF U19 ( .A(iData[501]), .Z(tmpData[565]));
Q_BUF U20 ( .A(iData[500]), .Z(tmpData[564]));
Q_BUF U21 ( .A(iData[499]), .Z(tmpData[563]));
Q_BUF U22 ( .A(iData[498]), .Z(tmpData[562]));
Q_BUF U23 ( .A(iData[497]), .Z(tmpData[561]));
Q_BUF U24 ( .A(iData[496]), .Z(tmpData[560]));
Q_BUF U25 ( .A(iData[495]), .Z(tmpData[559]));
Q_BUF U26 ( .A(iData[494]), .Z(tmpData[558]));
Q_BUF U27 ( .A(iData[493]), .Z(tmpData[557]));
Q_BUF U28 ( .A(iData[492]), .Z(tmpData[556]));
Q_BUF U29 ( .A(iData[491]), .Z(tmpData[555]));
Q_BUF U30 ( .A(iData[490]), .Z(tmpData[554]));
Q_BUF U31 ( .A(iData[489]), .Z(tmpData[553]));
Q_BUF U32 ( .A(iData[488]), .Z(tmpData[552]));
Q_BUF U33 ( .A(iData[487]), .Z(tmpData[551]));
Q_BUF U34 ( .A(iData[486]), .Z(tmpData[550]));
Q_BUF U35 ( .A(iData[485]), .Z(tmpData[549]));
Q_BUF U36 ( .A(iData[484]), .Z(tmpData[548]));
Q_BUF U37 ( .A(iData[483]), .Z(tmpData[547]));
Q_BUF U38 ( .A(iData[482]), .Z(tmpData[546]));
Q_BUF U39 ( .A(iData[481]), .Z(tmpData[545]));
Q_BUF U40 ( .A(iData[480]), .Z(tmpData[544]));
Q_BUF U41 ( .A(iData[479]), .Z(tmpData[543]));
Q_BUF U42 ( .A(iData[478]), .Z(tmpData[542]));
Q_BUF U43 ( .A(iData[477]), .Z(tmpData[541]));
Q_BUF U44 ( .A(iData[476]), .Z(tmpData[540]));
Q_BUF U45 ( .A(iData[475]), .Z(tmpData[539]));
Q_BUF U46 ( .A(iData[474]), .Z(tmpData[538]));
Q_BUF U47 ( .A(iData[473]), .Z(tmpData[537]));
Q_BUF U48 ( .A(iData[472]), .Z(tmpData[536]));
Q_BUF U49 ( .A(iData[471]), .Z(tmpData[535]));
Q_BUF U50 ( .A(iData[470]), .Z(tmpData[534]));
Q_BUF U51 ( .A(iData[469]), .Z(tmpData[533]));
Q_BUF U52 ( .A(iData[468]), .Z(tmpData[532]));
Q_BUF U53 ( .A(iData[467]), .Z(tmpData[531]));
Q_BUF U54 ( .A(iData[466]), .Z(tmpData[530]));
Q_BUF U55 ( .A(iData[465]), .Z(tmpData[529]));
Q_BUF U56 ( .A(iData[464]), .Z(tmpData[528]));
Q_BUF U57 ( .A(iData[463]), .Z(tmpData[527]));
Q_BUF U58 ( .A(iData[462]), .Z(tmpData[526]));
Q_BUF U59 ( .A(iData[461]), .Z(tmpData[525]));
Q_BUF U60 ( .A(iData[460]), .Z(tmpData[524]));
Q_BUF U61 ( .A(iData[459]), .Z(tmpData[523]));
Q_BUF U62 ( .A(iData[458]), .Z(tmpData[522]));
Q_BUF U63 ( .A(iData[457]), .Z(tmpData[521]));
Q_BUF U64 ( .A(iData[456]), .Z(tmpData[520]));
Q_BUF U65 ( .A(iData[455]), .Z(tmpData[519]));
Q_BUF U66 ( .A(iData[454]), .Z(tmpData[518]));
Q_BUF U67 ( .A(iData[453]), .Z(tmpData[517]));
Q_BUF U68 ( .A(iData[452]), .Z(tmpData[516]));
Q_BUF U69 ( .A(iData[451]), .Z(tmpData[515]));
Q_BUF U70 ( .A(iData[450]), .Z(tmpData[514]));
Q_BUF U71 ( .A(iData[449]), .Z(tmpData[513]));
Q_BUF U72 ( .A(iData[448]), .Z(tmpData[512]));
Q_BUF U73 ( .A(iData[447]), .Z(tmpData[511]));
Q_BUF U74 ( .A(iData[446]), .Z(tmpData[510]));
Q_BUF U75 ( .A(iData[445]), .Z(tmpData[509]));
Q_BUF U76 ( .A(iData[444]), .Z(tmpData[508]));
Q_BUF U77 ( .A(iData[443]), .Z(tmpData[507]));
Q_BUF U78 ( .A(iData[442]), .Z(tmpData[506]));
Q_BUF U79 ( .A(iData[441]), .Z(tmpData[505]));
Q_BUF U80 ( .A(iData[440]), .Z(tmpData[504]));
Q_BUF U81 ( .A(iData[439]), .Z(tmpData[503]));
Q_BUF U82 ( .A(iData[438]), .Z(tmpData[502]));
Q_BUF U83 ( .A(iData[437]), .Z(tmpData[501]));
Q_BUF U84 ( .A(iData[436]), .Z(tmpData[500]));
Q_BUF U85 ( .A(iData[435]), .Z(tmpData[499]));
Q_BUF U86 ( .A(iData[434]), .Z(tmpData[498]));
Q_BUF U87 ( .A(iData[433]), .Z(tmpData[497]));
Q_BUF U88 ( .A(iData[432]), .Z(tmpData[496]));
Q_BUF U89 ( .A(iData[431]), .Z(tmpData[495]));
Q_BUF U90 ( .A(iData[430]), .Z(tmpData[494]));
Q_BUF U91 ( .A(iData[429]), .Z(tmpData[493]));
Q_BUF U92 ( .A(iData[428]), .Z(tmpData[492]));
Q_BUF U93 ( .A(iData[427]), .Z(tmpData[491]));
Q_BUF U94 ( .A(iData[426]), .Z(tmpData[490]));
Q_BUF U95 ( .A(iData[425]), .Z(tmpData[489]));
Q_BUF U96 ( .A(iData[424]), .Z(tmpData[488]));
Q_BUF U97 ( .A(iData[423]), .Z(tmpData[487]));
Q_BUF U98 ( .A(iData[422]), .Z(tmpData[486]));
Q_BUF U99 ( .A(iData[421]), .Z(tmpData[485]));
Q_BUF U100 ( .A(iData[420]), .Z(tmpData[484]));
Q_BUF U101 ( .A(iData[419]), .Z(tmpData[483]));
Q_BUF U102 ( .A(iData[418]), .Z(tmpData[482]));
Q_BUF U103 ( .A(iData[417]), .Z(tmpData[481]));
Q_BUF U104 ( .A(iData[416]), .Z(tmpData[480]));
Q_BUF U105 ( .A(iData[415]), .Z(tmpData[479]));
Q_BUF U106 ( .A(iData[414]), .Z(tmpData[478]));
Q_BUF U107 ( .A(iData[413]), .Z(tmpData[477]));
Q_BUF U108 ( .A(iData[412]), .Z(tmpData[476]));
Q_BUF U109 ( .A(iData[411]), .Z(tmpData[475]));
Q_BUF U110 ( .A(iData[410]), .Z(tmpData[474]));
Q_BUF U111 ( .A(iData[409]), .Z(tmpData[473]));
Q_BUF U112 ( .A(iData[408]), .Z(tmpData[472]));
Q_BUF U113 ( .A(iData[407]), .Z(tmpData[471]));
Q_BUF U114 ( .A(iData[406]), .Z(tmpData[470]));
Q_BUF U115 ( .A(iData[405]), .Z(tmpData[469]));
Q_BUF U116 ( .A(iData[404]), .Z(tmpData[468]));
Q_BUF U117 ( .A(iData[403]), .Z(tmpData[467]));
Q_BUF U118 ( .A(iData[402]), .Z(tmpData[466]));
Q_BUF U119 ( .A(iData[401]), .Z(tmpData[465]));
Q_BUF U120 ( .A(iData[400]), .Z(tmpData[464]));
Q_BUF U121 ( .A(iData[399]), .Z(tmpData[463]));
Q_BUF U122 ( .A(iData[398]), .Z(tmpData[462]));
Q_BUF U123 ( .A(iData[397]), .Z(tmpData[461]));
Q_BUF U124 ( .A(iData[396]), .Z(tmpData[460]));
Q_BUF U125 ( .A(iData[395]), .Z(tmpData[459]));
Q_BUF U126 ( .A(iData[394]), .Z(tmpData[458]));
Q_BUF U127 ( .A(iData[393]), .Z(tmpData[457]));
Q_BUF U128 ( .A(iData[392]), .Z(tmpData[456]));
Q_BUF U129 ( .A(iData[391]), .Z(tmpData[455]));
Q_BUF U130 ( .A(iData[390]), .Z(tmpData[454]));
Q_BUF U131 ( .A(iData[389]), .Z(tmpData[453]));
Q_BUF U132 ( .A(iData[388]), .Z(tmpData[452]));
Q_BUF U133 ( .A(iData[387]), .Z(tmpData[451]));
Q_BUF U134 ( .A(iData[386]), .Z(tmpData[450]));
Q_BUF U135 ( .A(iData[385]), .Z(tmpData[449]));
Q_BUF U136 ( .A(iData[384]), .Z(tmpData[448]));
Q_BUF U137 ( .A(iData[383]), .Z(tmpData[447]));
Q_BUF U138 ( .A(iData[382]), .Z(tmpData[446]));
Q_BUF U139 ( .A(iData[381]), .Z(tmpData[445]));
Q_BUF U140 ( .A(iData[380]), .Z(tmpData[444]));
Q_BUF U141 ( .A(iData[379]), .Z(tmpData[443]));
Q_BUF U142 ( .A(iData[378]), .Z(tmpData[442]));
Q_BUF U143 ( .A(iData[377]), .Z(tmpData[441]));
Q_BUF U144 ( .A(iData[376]), .Z(tmpData[440]));
Q_BUF U145 ( .A(iData[375]), .Z(tmpData[439]));
Q_BUF U146 ( .A(iData[374]), .Z(tmpData[438]));
Q_BUF U147 ( .A(iData[373]), .Z(tmpData[437]));
Q_BUF U148 ( .A(iData[372]), .Z(tmpData[436]));
Q_BUF U149 ( .A(iData[371]), .Z(tmpData[435]));
Q_BUF U150 ( .A(iData[370]), .Z(tmpData[434]));
Q_BUF U151 ( .A(iData[369]), .Z(tmpData[433]));
Q_BUF U152 ( .A(iData[368]), .Z(tmpData[432]));
Q_BUF U153 ( .A(iData[367]), .Z(tmpData[431]));
Q_BUF U154 ( .A(iData[366]), .Z(tmpData[430]));
Q_BUF U155 ( .A(iData[365]), .Z(tmpData[429]));
Q_BUF U156 ( .A(iData[364]), .Z(tmpData[428]));
Q_BUF U157 ( .A(iData[363]), .Z(tmpData[427]));
Q_BUF U158 ( .A(iData[362]), .Z(tmpData[426]));
Q_BUF U159 ( .A(iData[361]), .Z(tmpData[425]));
Q_BUF U160 ( .A(iData[360]), .Z(tmpData[424]));
Q_BUF U161 ( .A(iData[359]), .Z(tmpData[423]));
Q_BUF U162 ( .A(iData[358]), .Z(tmpData[422]));
Q_BUF U163 ( .A(iData[357]), .Z(tmpData[421]));
Q_BUF U164 ( .A(iData[356]), .Z(tmpData[420]));
Q_BUF U165 ( .A(iData[355]), .Z(tmpData[419]));
Q_BUF U166 ( .A(iData[354]), .Z(tmpData[418]));
Q_BUF U167 ( .A(iData[353]), .Z(tmpData[417]));
Q_BUF U168 ( .A(iData[352]), .Z(tmpData[416]));
Q_BUF U169 ( .A(iData[351]), .Z(tmpData[415]));
Q_BUF U170 ( .A(iData[350]), .Z(tmpData[414]));
Q_BUF U171 ( .A(iData[349]), .Z(tmpData[413]));
Q_BUF U172 ( .A(iData[348]), .Z(tmpData[412]));
Q_BUF U173 ( .A(iData[347]), .Z(tmpData[411]));
Q_BUF U174 ( .A(iData[346]), .Z(tmpData[410]));
Q_BUF U175 ( .A(iData[345]), .Z(tmpData[409]));
Q_BUF U176 ( .A(iData[344]), .Z(tmpData[408]));
Q_BUF U177 ( .A(iData[343]), .Z(tmpData[407]));
Q_BUF U178 ( .A(iData[342]), .Z(tmpData[406]));
Q_BUF U179 ( .A(iData[341]), .Z(tmpData[405]));
Q_BUF U180 ( .A(iData[340]), .Z(tmpData[404]));
Q_BUF U181 ( .A(iData[339]), .Z(tmpData[403]));
Q_BUF U182 ( .A(iData[338]), .Z(tmpData[402]));
Q_BUF U183 ( .A(iData[337]), .Z(tmpData[401]));
Q_BUF U184 ( .A(iData[336]), .Z(tmpData[400]));
Q_BUF U185 ( .A(iData[335]), .Z(tmpData[399]));
Q_BUF U186 ( .A(iData[334]), .Z(tmpData[398]));
Q_BUF U187 ( .A(iData[333]), .Z(tmpData[397]));
Q_BUF U188 ( .A(iData[332]), .Z(tmpData[396]));
Q_BUF U189 ( .A(iData[331]), .Z(tmpData[395]));
Q_BUF U190 ( .A(iData[330]), .Z(tmpData[394]));
Q_BUF U191 ( .A(iData[329]), .Z(tmpData[393]));
Q_BUF U192 ( .A(iData[328]), .Z(tmpData[392]));
Q_BUF U193 ( .A(iData[327]), .Z(tmpData[391]));
Q_BUF U194 ( .A(iData[326]), .Z(tmpData[390]));
Q_BUF U195 ( .A(iData[325]), .Z(tmpData[389]));
Q_BUF U196 ( .A(iData[324]), .Z(tmpData[388]));
Q_BUF U197 ( .A(iData[323]), .Z(tmpData[387]));
Q_BUF U198 ( .A(iData[322]), .Z(tmpData[386]));
Q_BUF U199 ( .A(iData[321]), .Z(tmpData[385]));
Q_BUF U200 ( .A(iData[320]), .Z(tmpData[384]));
Q_BUF U201 ( .A(iData[319]), .Z(tmpData[383]));
Q_BUF U202 ( .A(iData[318]), .Z(tmpData[382]));
Q_BUF U203 ( .A(iData[317]), .Z(tmpData[381]));
Q_BUF U204 ( .A(iData[316]), .Z(tmpData[380]));
Q_BUF U205 ( .A(iData[315]), .Z(tmpData[379]));
Q_BUF U206 ( .A(iData[314]), .Z(tmpData[378]));
Q_BUF U207 ( .A(iData[313]), .Z(tmpData[377]));
Q_BUF U208 ( .A(iData[312]), .Z(tmpData[376]));
Q_BUF U209 ( .A(iData[311]), .Z(tmpData[375]));
Q_BUF U210 ( .A(iData[310]), .Z(tmpData[374]));
Q_BUF U211 ( .A(iData[309]), .Z(tmpData[373]));
Q_BUF U212 ( .A(iData[308]), .Z(tmpData[372]));
Q_BUF U213 ( .A(iData[307]), .Z(tmpData[371]));
Q_BUF U214 ( .A(iData[306]), .Z(tmpData[370]));
Q_BUF U215 ( .A(iData[305]), .Z(tmpData[369]));
Q_BUF U216 ( .A(iData[304]), .Z(tmpData[368]));
Q_BUF U217 ( .A(iData[303]), .Z(tmpData[367]));
Q_BUF U218 ( .A(iData[302]), .Z(tmpData[366]));
Q_BUF U219 ( .A(iData[301]), .Z(tmpData[365]));
Q_BUF U220 ( .A(iData[300]), .Z(tmpData[364]));
Q_BUF U221 ( .A(iData[299]), .Z(tmpData[363]));
Q_BUF U222 ( .A(iData[298]), .Z(tmpData[362]));
Q_BUF U223 ( .A(iData[297]), .Z(tmpData[361]));
Q_BUF U224 ( .A(iData[296]), .Z(tmpData[360]));
Q_BUF U225 ( .A(iData[295]), .Z(tmpData[359]));
Q_BUF U226 ( .A(iData[294]), .Z(tmpData[358]));
Q_BUF U227 ( .A(iData[293]), .Z(tmpData[357]));
Q_BUF U228 ( .A(iData[292]), .Z(tmpData[356]));
Q_BUF U229 ( .A(iData[291]), .Z(tmpData[355]));
Q_BUF U230 ( .A(iData[290]), .Z(tmpData[354]));
Q_BUF U231 ( .A(iData[289]), .Z(tmpData[353]));
Q_BUF U232 ( .A(iData[288]), .Z(tmpData[352]));
Q_BUF U233 ( .A(iData[287]), .Z(tmpData[351]));
Q_BUF U234 ( .A(iData[286]), .Z(tmpData[350]));
Q_BUF U235 ( .A(iData[285]), .Z(tmpData[349]));
Q_BUF U236 ( .A(iData[284]), .Z(tmpData[348]));
Q_BUF U237 ( .A(iData[283]), .Z(tmpData[347]));
Q_BUF U238 ( .A(iData[282]), .Z(tmpData[346]));
Q_BUF U239 ( .A(iData[281]), .Z(tmpData[345]));
Q_BUF U240 ( .A(iData[280]), .Z(tmpData[344]));
Q_BUF U241 ( .A(iData[279]), .Z(tmpData[343]));
Q_BUF U242 ( .A(iData[278]), .Z(tmpData[342]));
Q_BUF U243 ( .A(iData[277]), .Z(tmpData[341]));
Q_BUF U244 ( .A(iData[276]), .Z(tmpData[340]));
Q_BUF U245 ( .A(iData[275]), .Z(tmpData[339]));
Q_BUF U246 ( .A(iData[274]), .Z(tmpData[338]));
Q_BUF U247 ( .A(iData[273]), .Z(tmpData[337]));
Q_BUF U248 ( .A(iData[272]), .Z(tmpData[336]));
Q_BUF U249 ( .A(iData[271]), .Z(tmpData[335]));
Q_BUF U250 ( .A(iData[270]), .Z(tmpData[334]));
Q_BUF U251 ( .A(iData[269]), .Z(tmpData[333]));
Q_BUF U252 ( .A(iData[268]), .Z(tmpData[332]));
Q_BUF U253 ( .A(iData[267]), .Z(tmpData[331]));
Q_BUF U254 ( .A(iData[266]), .Z(tmpData[330]));
Q_BUF U255 ( .A(iData[265]), .Z(tmpData[329]));
Q_BUF U256 ( .A(iData[264]), .Z(tmpData[328]));
Q_BUF U257 ( .A(iData[263]), .Z(tmpData[327]));
Q_BUF U258 ( .A(iData[262]), .Z(tmpData[326]));
Q_BUF U259 ( .A(iData[261]), .Z(tmpData[325]));
Q_BUF U260 ( .A(iData[260]), .Z(tmpData[324]));
Q_BUF U261 ( .A(iData[259]), .Z(tmpData[323]));
Q_BUF U262 ( .A(iData[258]), .Z(tmpData[322]));
Q_BUF U263 ( .A(iData[257]), .Z(tmpData[321]));
Q_BUF U264 ( .A(iData[256]), .Z(tmpData[320]));
Q_BUF U265 ( .A(iData[255]), .Z(tmpData[319]));
Q_BUF U266 ( .A(iData[254]), .Z(tmpData[318]));
Q_BUF U267 ( .A(iData[253]), .Z(tmpData[317]));
Q_BUF U268 ( .A(iData[252]), .Z(tmpData[316]));
Q_BUF U269 ( .A(iData[251]), .Z(tmpData[315]));
Q_BUF U270 ( .A(iData[250]), .Z(tmpData[314]));
Q_BUF U271 ( .A(iData[249]), .Z(tmpData[313]));
Q_BUF U272 ( .A(iData[248]), .Z(tmpData[312]));
Q_BUF U273 ( .A(iData[247]), .Z(tmpData[311]));
Q_BUF U274 ( .A(iData[246]), .Z(tmpData[310]));
Q_BUF U275 ( .A(iData[245]), .Z(tmpData[309]));
Q_BUF U276 ( .A(iData[244]), .Z(tmpData[308]));
Q_BUF U277 ( .A(iData[243]), .Z(tmpData[307]));
Q_BUF U278 ( .A(iData[242]), .Z(tmpData[306]));
Q_BUF U279 ( .A(iData[241]), .Z(tmpData[305]));
Q_BUF U280 ( .A(iData[240]), .Z(tmpData[304]));
Q_BUF U281 ( .A(iData[239]), .Z(tmpData[303]));
Q_BUF U282 ( .A(iData[238]), .Z(tmpData[302]));
Q_BUF U283 ( .A(iData[237]), .Z(tmpData[301]));
Q_BUF U284 ( .A(iData[236]), .Z(tmpData[300]));
Q_BUF U285 ( .A(iData[235]), .Z(tmpData[299]));
Q_BUF U286 ( .A(iData[234]), .Z(tmpData[298]));
Q_BUF U287 ( .A(iData[233]), .Z(tmpData[297]));
Q_BUF U288 ( .A(iData[232]), .Z(tmpData[296]));
Q_BUF U289 ( .A(iData[231]), .Z(tmpData[295]));
Q_BUF U290 ( .A(iData[230]), .Z(tmpData[294]));
Q_BUF U291 ( .A(iData[229]), .Z(tmpData[293]));
Q_BUF U292 ( .A(iData[228]), .Z(tmpData[292]));
Q_BUF U293 ( .A(iData[227]), .Z(tmpData[291]));
Q_BUF U294 ( .A(iData[226]), .Z(tmpData[290]));
Q_BUF U295 ( .A(iData[225]), .Z(tmpData[289]));
Q_BUF U296 ( .A(iData[224]), .Z(tmpData[288]));
Q_BUF U297 ( .A(iData[223]), .Z(tmpData[287]));
Q_BUF U298 ( .A(iData[222]), .Z(tmpData[286]));
Q_BUF U299 ( .A(iData[221]), .Z(tmpData[285]));
Q_BUF U300 ( .A(iData[220]), .Z(tmpData[284]));
Q_BUF U301 ( .A(iData[219]), .Z(tmpData[283]));
Q_BUF U302 ( .A(iData[218]), .Z(tmpData[282]));
Q_BUF U303 ( .A(iData[217]), .Z(tmpData[281]));
Q_BUF U304 ( .A(iData[216]), .Z(tmpData[280]));
Q_BUF U305 ( .A(iData[215]), .Z(tmpData[279]));
Q_BUF U306 ( .A(iData[214]), .Z(tmpData[278]));
Q_BUF U307 ( .A(iData[213]), .Z(tmpData[277]));
Q_BUF U308 ( .A(iData[212]), .Z(tmpData[276]));
Q_BUF U309 ( .A(iData[211]), .Z(tmpData[275]));
Q_BUF U310 ( .A(iData[210]), .Z(tmpData[274]));
Q_BUF U311 ( .A(iData[209]), .Z(tmpData[273]));
Q_BUF U312 ( .A(iData[208]), .Z(tmpData[272]));
Q_BUF U313 ( .A(iData[207]), .Z(tmpData[271]));
Q_BUF U314 ( .A(iData[206]), .Z(tmpData[270]));
Q_BUF U315 ( .A(iData[205]), .Z(tmpData[269]));
Q_BUF U316 ( .A(iData[204]), .Z(tmpData[268]));
Q_BUF U317 ( .A(iData[203]), .Z(tmpData[267]));
Q_BUF U318 ( .A(iData[202]), .Z(tmpData[266]));
Q_BUF U319 ( .A(iData[201]), .Z(tmpData[265]));
Q_BUF U320 ( .A(iData[200]), .Z(tmpData[264]));
Q_BUF U321 ( .A(iData[199]), .Z(tmpData[263]));
Q_BUF U322 ( .A(iData[198]), .Z(tmpData[262]));
Q_BUF U323 ( .A(iData[197]), .Z(tmpData[261]));
Q_BUF U324 ( .A(iData[196]), .Z(tmpData[260]));
Q_BUF U325 ( .A(iData[195]), .Z(tmpData[259]));
Q_BUF U326 ( .A(iData[194]), .Z(tmpData[258]));
Q_BUF U327 ( .A(iData[193]), .Z(tmpData[257]));
Q_BUF U328 ( .A(iData[192]), .Z(tmpData[256]));
Q_BUF U329 ( .A(iData[191]), .Z(tmpData[255]));
Q_BUF U330 ( .A(iData[190]), .Z(tmpData[254]));
Q_BUF U331 ( .A(iData[189]), .Z(tmpData[253]));
Q_BUF U332 ( .A(iData[188]), .Z(tmpData[252]));
Q_BUF U333 ( .A(iData[187]), .Z(tmpData[251]));
Q_BUF U334 ( .A(iData[186]), .Z(tmpData[250]));
Q_BUF U335 ( .A(iData[185]), .Z(tmpData[249]));
Q_BUF U336 ( .A(iData[184]), .Z(tmpData[248]));
Q_BUF U337 ( .A(iData[183]), .Z(tmpData[247]));
Q_BUF U338 ( .A(iData[182]), .Z(tmpData[246]));
Q_BUF U339 ( .A(iData[181]), .Z(tmpData[245]));
Q_BUF U340 ( .A(iData[180]), .Z(tmpData[244]));
Q_BUF U341 ( .A(iData[179]), .Z(tmpData[243]));
Q_BUF U342 ( .A(iData[178]), .Z(tmpData[242]));
Q_BUF U343 ( .A(iData[177]), .Z(tmpData[241]));
Q_BUF U344 ( .A(iData[176]), .Z(tmpData[240]));
Q_BUF U345 ( .A(iData[175]), .Z(tmpData[239]));
Q_BUF U346 ( .A(iData[174]), .Z(tmpData[238]));
Q_BUF U347 ( .A(iData[173]), .Z(tmpData[237]));
Q_BUF U348 ( .A(iData[172]), .Z(tmpData[236]));
Q_BUF U349 ( .A(iData[171]), .Z(tmpData[235]));
Q_BUF U350 ( .A(iData[170]), .Z(tmpData[234]));
Q_BUF U351 ( .A(iData[169]), .Z(tmpData[233]));
Q_BUF U352 ( .A(iData[168]), .Z(tmpData[232]));
Q_BUF U353 ( .A(iData[167]), .Z(tmpData[231]));
Q_BUF U354 ( .A(iData[166]), .Z(tmpData[230]));
Q_BUF U355 ( .A(iData[165]), .Z(tmpData[229]));
Q_BUF U356 ( .A(iData[164]), .Z(tmpData[228]));
Q_BUF U357 ( .A(iData[163]), .Z(tmpData[227]));
Q_BUF U358 ( .A(iData[162]), .Z(tmpData[226]));
Q_BUF U359 ( .A(iData[161]), .Z(tmpData[225]));
Q_BUF U360 ( .A(iData[160]), .Z(tmpData[224]));
Q_BUF U361 ( .A(iData[159]), .Z(tmpData[223]));
Q_BUF U362 ( .A(iData[158]), .Z(tmpData[222]));
Q_BUF U363 ( .A(iData[157]), .Z(tmpData[221]));
Q_BUF U364 ( .A(iData[156]), .Z(tmpData[220]));
Q_BUF U365 ( .A(iData[155]), .Z(tmpData[219]));
Q_BUF U366 ( .A(iData[154]), .Z(tmpData[218]));
Q_BUF U367 ( .A(iData[153]), .Z(tmpData[217]));
Q_BUF U368 ( .A(iData[152]), .Z(tmpData[216]));
Q_BUF U369 ( .A(iData[151]), .Z(tmpData[215]));
Q_BUF U370 ( .A(iData[150]), .Z(tmpData[214]));
Q_BUF U371 ( .A(iData[149]), .Z(tmpData[213]));
Q_BUF U372 ( .A(iData[148]), .Z(tmpData[212]));
Q_BUF U373 ( .A(iData[147]), .Z(tmpData[211]));
Q_BUF U374 ( .A(iData[146]), .Z(tmpData[210]));
Q_BUF U375 ( .A(iData[145]), .Z(tmpData[209]));
Q_BUF U376 ( .A(iData[144]), .Z(tmpData[208]));
Q_BUF U377 ( .A(iData[143]), .Z(tmpData[207]));
Q_BUF U378 ( .A(iData[142]), .Z(tmpData[206]));
Q_BUF U379 ( .A(iData[141]), .Z(tmpData[205]));
Q_BUF U380 ( .A(iData[140]), .Z(tmpData[204]));
Q_BUF U381 ( .A(iData[139]), .Z(tmpData[203]));
Q_BUF U382 ( .A(iData[138]), .Z(tmpData[202]));
Q_BUF U383 ( .A(iData[137]), .Z(tmpData[201]));
Q_BUF U384 ( .A(iData[136]), .Z(tmpData[200]));
Q_BUF U385 ( .A(iData[135]), .Z(tmpData[199]));
Q_BUF U386 ( .A(iData[134]), .Z(tmpData[198]));
Q_BUF U387 ( .A(iData[133]), .Z(tmpData[197]));
Q_BUF U388 ( .A(iData[132]), .Z(tmpData[196]));
Q_BUF U389 ( .A(iData[131]), .Z(tmpData[195]));
Q_BUF U390 ( .A(iData[130]), .Z(tmpData[194]));
Q_BUF U391 ( .A(iData[129]), .Z(tmpData[193]));
Q_BUF U392 ( .A(iData[128]), .Z(tmpData[192]));
Q_BUF U393 ( .A(iData[127]), .Z(tmpData[191]));
Q_BUF U394 ( .A(iData[126]), .Z(tmpData[190]));
Q_BUF U395 ( .A(iData[125]), .Z(tmpData[189]));
Q_BUF U396 ( .A(iData[124]), .Z(tmpData[188]));
Q_BUF U397 ( .A(iData[123]), .Z(tmpData[187]));
Q_BUF U398 ( .A(iData[122]), .Z(tmpData[186]));
Q_BUF U399 ( .A(iData[121]), .Z(tmpData[185]));
Q_BUF U400 ( .A(iData[120]), .Z(tmpData[184]));
Q_BUF U401 ( .A(iData[119]), .Z(tmpData[183]));
Q_BUF U402 ( .A(iData[118]), .Z(tmpData[182]));
Q_BUF U403 ( .A(iData[117]), .Z(tmpData[181]));
Q_BUF U404 ( .A(iData[116]), .Z(tmpData[180]));
Q_BUF U405 ( .A(iData[115]), .Z(tmpData[179]));
Q_BUF U406 ( .A(iData[114]), .Z(tmpData[178]));
Q_BUF U407 ( .A(iData[113]), .Z(tmpData[177]));
Q_BUF U408 ( .A(iData[112]), .Z(tmpData[176]));
Q_BUF U409 ( .A(iData[111]), .Z(tmpData[175]));
Q_BUF U410 ( .A(iData[110]), .Z(tmpData[174]));
Q_BUF U411 ( .A(iData[109]), .Z(tmpData[173]));
Q_BUF U412 ( .A(iData[108]), .Z(tmpData[172]));
Q_BUF U413 ( .A(iData[107]), .Z(tmpData[171]));
Q_BUF U414 ( .A(iData[106]), .Z(tmpData[170]));
Q_BUF U415 ( .A(iData[105]), .Z(tmpData[169]));
Q_BUF U416 ( .A(iData[104]), .Z(tmpData[168]));
Q_BUF U417 ( .A(iData[103]), .Z(tmpData[167]));
Q_BUF U418 ( .A(iData[102]), .Z(tmpData[166]));
Q_BUF U419 ( .A(iData[101]), .Z(tmpData[165]));
Q_BUF U420 ( .A(iData[100]), .Z(tmpData[164]));
Q_BUF U421 ( .A(iData[99]), .Z(tmpData[163]));
Q_BUF U422 ( .A(iData[98]), .Z(tmpData[162]));
Q_BUF U423 ( .A(iData[97]), .Z(tmpData[161]));
Q_BUF U424 ( .A(iData[96]), .Z(tmpData[160]));
Q_BUF U425 ( .A(iData[95]), .Z(tmpData[159]));
Q_BUF U426 ( .A(iData[94]), .Z(tmpData[158]));
Q_BUF U427 ( .A(iData[93]), .Z(tmpData[157]));
Q_BUF U428 ( .A(iData[92]), .Z(tmpData[156]));
Q_BUF U429 ( .A(iData[91]), .Z(tmpData[155]));
Q_BUF U430 ( .A(iData[90]), .Z(tmpData[154]));
Q_BUF U431 ( .A(iData[89]), .Z(tmpData[153]));
Q_BUF U432 ( .A(iData[88]), .Z(tmpData[152]));
Q_BUF U433 ( .A(iData[87]), .Z(tmpData[151]));
Q_BUF U434 ( .A(iData[86]), .Z(tmpData[150]));
Q_BUF U435 ( .A(iData[85]), .Z(tmpData[149]));
Q_BUF U436 ( .A(iData[84]), .Z(tmpData[148]));
Q_BUF U437 ( .A(iData[83]), .Z(tmpData[147]));
Q_BUF U438 ( .A(iData[82]), .Z(tmpData[146]));
Q_BUF U439 ( .A(iData[81]), .Z(tmpData[145]));
Q_BUF U440 ( .A(iData[80]), .Z(tmpData[144]));
Q_BUF U441 ( .A(iData[79]), .Z(tmpData[143]));
Q_BUF U442 ( .A(iData[78]), .Z(tmpData[142]));
Q_BUF U443 ( .A(iData[77]), .Z(tmpData[141]));
Q_BUF U444 ( .A(iData[76]), .Z(tmpData[140]));
Q_BUF U445 ( .A(iData[75]), .Z(tmpData[139]));
Q_BUF U446 ( .A(iData[74]), .Z(tmpData[138]));
Q_BUF U447 ( .A(iData[73]), .Z(tmpData[137]));
Q_BUF U448 ( .A(iData[72]), .Z(tmpData[136]));
Q_BUF U449 ( .A(iData[71]), .Z(tmpData[135]));
Q_BUF U450 ( .A(iData[70]), .Z(tmpData[134]));
Q_BUF U451 ( .A(iData[69]), .Z(tmpData[133]));
Q_BUF U452 ( .A(iData[68]), .Z(tmpData[132]));
Q_BUF U453 ( .A(iData[67]), .Z(tmpData[131]));
Q_BUF U454 ( .A(iData[66]), .Z(tmpData[130]));
Q_BUF U455 ( .A(iData[65]), .Z(tmpData[129]));
Q_BUF U456 ( .A(iData[64]), .Z(tmpData[128]));
Q_BUF U457 ( .A(iData[63]), .Z(tmpData[127]));
Q_BUF U458 ( .A(iData[62]), .Z(tmpData[126]));
Q_BUF U459 ( .A(iData[61]), .Z(tmpData[125]));
Q_BUF U460 ( .A(iData[60]), .Z(tmpData[124]));
Q_BUF U461 ( .A(iData[59]), .Z(tmpData[123]));
Q_BUF U462 ( .A(iData[58]), .Z(tmpData[122]));
Q_BUF U463 ( .A(iData[57]), .Z(tmpData[121]));
Q_BUF U464 ( .A(iData[56]), .Z(tmpData[120]));
Q_BUF U465 ( .A(iData[55]), .Z(tmpData[119]));
Q_BUF U466 ( .A(iData[54]), .Z(tmpData[118]));
Q_BUF U467 ( .A(iData[53]), .Z(tmpData[117]));
Q_BUF U468 ( .A(iData[52]), .Z(tmpData[116]));
Q_BUF U469 ( .A(iData[51]), .Z(tmpData[115]));
Q_BUF U470 ( .A(iData[50]), .Z(tmpData[114]));
Q_BUF U471 ( .A(iData[49]), .Z(tmpData[113]));
Q_BUF U472 ( .A(iData[48]), .Z(tmpData[112]));
Q_BUF U473 ( .A(iData[47]), .Z(tmpData[111]));
Q_BUF U474 ( .A(iData[46]), .Z(tmpData[110]));
Q_BUF U475 ( .A(iData[45]), .Z(tmpData[109]));
Q_BUF U476 ( .A(iData[44]), .Z(tmpData[108]));
Q_BUF U477 ( .A(iData[43]), .Z(tmpData[107]));
Q_BUF U478 ( .A(iData[42]), .Z(tmpData[106]));
Q_BUF U479 ( .A(iData[41]), .Z(tmpData[105]));
Q_BUF U480 ( .A(iData[40]), .Z(tmpData[104]));
Q_BUF U481 ( .A(iData[39]), .Z(tmpData[103]));
Q_BUF U482 ( .A(iData[38]), .Z(tmpData[102]));
Q_BUF U483 ( .A(iData[37]), .Z(tmpData[101]));
Q_BUF U484 ( .A(iData[36]), .Z(tmpData[100]));
Q_BUF U485 ( .A(iData[35]), .Z(tmpData[99]));
Q_BUF U486 ( .A(iData[34]), .Z(tmpData[98]));
Q_BUF U487 ( .A(iData[33]), .Z(tmpData[97]));
Q_BUF U488 ( .A(iData[32]), .Z(tmpData[96]));
Q_BUF U489 ( .A(iData[31]), .Z(tmpData[95]));
Q_BUF U490 ( .A(iData[30]), .Z(tmpData[94]));
Q_BUF U491 ( .A(iData[29]), .Z(tmpData[93]));
Q_BUF U492 ( .A(iData[28]), .Z(tmpData[92]));
Q_BUF U493 ( .A(iData[27]), .Z(tmpData[91]));
Q_BUF U494 ( .A(iData[26]), .Z(tmpData[90]));
Q_BUF U495 ( .A(iData[25]), .Z(tmpData[89]));
Q_BUF U496 ( .A(iData[24]), .Z(tmpData[88]));
Q_BUF U497 ( .A(iData[23]), .Z(tmpData[87]));
Q_BUF U498 ( .A(iData[22]), .Z(tmpData[86]));
Q_BUF U499 ( .A(iData[21]), .Z(tmpData[85]));
Q_BUF U500 ( .A(iData[20]), .Z(tmpData[84]));
Q_BUF U501 ( .A(iData[19]), .Z(tmpData[83]));
Q_BUF U502 ( .A(iData[18]), .Z(tmpData[82]));
Q_BUF U503 ( .A(iData[17]), .Z(tmpData[81]));
Q_BUF U504 ( .A(iData[16]), .Z(tmpData[80]));
Q_BUF U505 ( .A(iData[15]), .Z(tmpData[79]));
Q_BUF U506 ( .A(iData[14]), .Z(tmpData[78]));
Q_BUF U507 ( .A(iData[13]), .Z(tmpData[77]));
Q_BUF U508 ( .A(iData[12]), .Z(tmpData[76]));
Q_BUF U509 ( .A(iData[11]), .Z(tmpData[75]));
Q_BUF U510 ( .A(iData[10]), .Z(tmpData[74]));
Q_BUF U511 ( .A(iData[9]), .Z(tmpData[73]));
Q_BUF U512 ( .A(iData[8]), .Z(tmpData[72]));
Q_BUF U513 ( .A(iData[7]), .Z(tmpData[71]));
Q_BUF U514 ( .A(iData[6]), .Z(tmpData[70]));
Q_BUF U515 ( .A(iData[5]), .Z(tmpData[69]));
Q_BUF U516 ( .A(iData[4]), .Z(tmpData[68]));
Q_BUF U517 ( .A(iData[3]), .Z(tmpData[67]));
Q_BUF U518 ( .A(iData[2]), .Z(tmpData[66]));
Q_BUF U519 ( .A(iData[1]), .Z(tmpData[65]));
Q_BUF U520 ( .A(iData[0]), .Z(tmpData[64]));
Q_BUF U521 ( .A(xhead[63]), .Z(tmpData[63]));
Q_BUF U522 ( .A(xhead[62]), .Z(tmpData[62]));
Q_BUF U523 ( .A(xhead[61]), .Z(tmpData[61]));
Q_BUF U524 ( .A(xhead[60]), .Z(tmpData[60]));
Q_BUF U525 ( .A(xhead[59]), .Z(tmpData[59]));
Q_BUF U526 ( .A(xhead[58]), .Z(tmpData[58]));
Q_BUF U527 ( .A(xhead[57]), .Z(tmpData[57]));
Q_BUF U528 ( .A(xhead[56]), .Z(tmpData[56]));
Q_BUF U529 ( .A(xhead[55]), .Z(tmpData[55]));
Q_BUF U530 ( .A(xhead[54]), .Z(tmpData[54]));
Q_BUF U531 ( .A(xhead[53]), .Z(tmpData[53]));
Q_BUF U532 ( .A(xhead[52]), .Z(tmpData[52]));
Q_BUF U533 ( .A(xhead[51]), .Z(tmpData[51]));
Q_BUF U534 ( .A(xhead[50]), .Z(tmpData[50]));
Q_BUF U535 ( .A(xhead[49]), .Z(tmpData[49]));
Q_BUF U536 ( .A(xhead[48]), .Z(tmpData[48]));
Q_BUF U537 ( .A(xhead[47]), .Z(tmpData[47]));
Q_BUF U538 ( .A(xhead[46]), .Z(tmpData[46]));
Q_BUF U539 ( .A(xhead[45]), .Z(tmpData[45]));
Q_BUF U540 ( .A(xhead[44]), .Z(tmpData[44]));
Q_BUF U541 ( .A(xhead[43]), .Z(tmpData[43]));
Q_BUF U542 ( .A(xhead[42]), .Z(tmpData[42]));
Q_BUF U543 ( .A(xhead[41]), .Z(tmpData[41]));
Q_BUF U544 ( .A(xhead[40]), .Z(tmpData[40]));
Q_BUF U545 ( .A(xhead[39]), .Z(tmpData[39]));
Q_BUF U546 ( .A(xhead[38]), .Z(tmpData[38]));
Q_BUF U547 ( .A(xhead[37]), .Z(tmpData[37]));
Q_BUF U548 ( .A(xhead[36]), .Z(tmpData[36]));
Q_BUF U549 ( .A(xhead[35]), .Z(tmpData[35]));
Q_BUF U550 ( .A(xhead[34]), .Z(tmpData[34]));
Q_BUF U551 ( .A(xhead[33]), .Z(tmpData[33]));
Q_BUF U552 ( .A(xhead[32]), .Z(tmpData[32]));
Q_BUF U553 ( .A(xhead[31]), .Z(tmpData[31]));
Q_BUF U554 ( .A(xhead[30]), .Z(tmpData[30]));
Q_BUF U555 ( .A(xhead[29]), .Z(tmpData[29]));
Q_BUF U556 ( .A(xhead[28]), .Z(tmpData[28]));
Q_BUF U557 ( .A(xhead[27]), .Z(tmpData[27]));
Q_BUF U558 ( .A(xhead[26]), .Z(tmpData[26]));
Q_BUF U559 ( .A(xhead[25]), .Z(tmpData[25]));
Q_BUF U560 ( .A(xhead[24]), .Z(tmpData[24]));
Q_BUF U561 ( .A(xhead[23]), .Z(tmpData[23]));
Q_BUF U562 ( .A(xhead[22]), .Z(tmpData[22]));
Q_BUF U563 ( .A(xhead[21]), .Z(tmpData[21]));
Q_BUF U564 ( .A(xhead[20]), .Z(tmpData[20]));
Q_BUF U565 ( .A(xhead[19]), .Z(tmpData[19]));
Q_BUF U566 ( .A(xhead[18]), .Z(tmpData[18]));
Q_BUF U567 ( .A(xhead[17]), .Z(tmpData[17]));
Q_BUF U568 ( .A(xhead[16]), .Z(tmpData[16]));
Q_BUF U569 ( .A(xhead[15]), .Z(tmpData[15]));
Q_BUF U570 ( .A(xhead[14]), .Z(tmpData[14]));
Q_BUF U571 ( .A(xhead[13]), .Z(tmpData[13]));
Q_BUF U572 ( .A(xhead[12]), .Z(tmpData[12]));
Q_BUF U573 ( .A(xhead[11]), .Z(tmpData[11]));
Q_BUF U574 ( .A(xhead[10]), .Z(tmpData[10]));
Q_BUF U575 ( .A(xhead[9]), .Z(tmpData[9]));
Q_BUF U576 ( .A(xhead[8]), .Z(tmpData[8]));
Q_BUF U577 ( .A(xhead[7]), .Z(tmpData[7]));
Q_BUF U578 ( .A(xhead[6]), .Z(tmpData[6]));
Q_BUF U579 ( .A(xhead[5]), .Z(tmpData[5]));
Q_BUF U580 ( .A(xhead[4]), .Z(tmpData[4]));
Q_BUF U581 ( .A(xhead[3]), .Z(tmpData[3]));
Q_BUF U582 ( .A(xhead[2]), .Z(tmpData[2]));
Q_BUF U583 ( .A(xhead[1]), .Z(tmpData[1]));
Q_BUF U584 ( .A(xhead[0]), .Z(tmpData[0]));
Q_INV U585 ( .A(n3271), .Z(n6887));
Q_INV U586 ( .A(n5216), .Z(n6886));
Q_INV U587 ( .A(n5217), .Z(n6885));
Q_NOT_TOUCH _zzqnthw ( .sig());
ixc_assign_64 _zz_strnp_0 ( _zy_simnet_rdCnt_0_w$[0:63], rdCnt[63:0]);
Q_XNR2 U590 ( .A0(newMarkBitsD[0]), .A1(newMarkBits[0]), .Z(n6881));
Q_XNR2 U591 ( .A0(newMarkBitsD[1]), .A1(newMarkBits[1]), .Z(n6880));
Q_XNR2 U592 ( .A0(newMarkBitsD[2]), .A1(newMarkBits[2]), .Z(n6879));
Q_XNR2 U593 ( .A0(newMarkBitsD[3]), .A1(newMarkBits[3]), .Z(n6878));
Q_AN03 U594 ( .A0(n6878), .A1(n6879), .A2(n6880), .Z(n6877));
Q_AN03 U595 ( .A0(n6881), .A1(n6877), .A2(n6868), .Z(n6876));
Q_BUFZP U596 ( .OE(n6874), .A(n6882), .Z(xc_top.svAsyncCall));
Q_ND03 U597 ( .A0(n5650), .A1(n6875), .A2(n6876), .Z(n6874));
Q_INV U598 ( .A(activeD), .Z(n6875));
Q_XOR2 U599 ( .A0(newMarkBits[0]), .A1(markBits[0]), .Z(n6873));
Q_XOR2 U600 ( .A0(newMarkBits[1]), .A1(markBits[1]), .Z(n6872));
Q_XOR2 U601 ( .A0(newMarkBits[2]), .A1(markBits[2]), .Z(n6871));
Q_XOR2 U602 ( .A0(newMarkBits[3]), .A1(markBits[3]), .Z(n6870));
Q_AN03 U603 ( .A0(n6870), .A1(n6871), .A2(n6872), .Z(n6869));
Q_AN03 U604 ( .A0(n6873), .A1(n6869), .A2(n6867), .Z(moveForwardN));
Q_INV U605 ( .A(moveForward), .Z(n6868));
Q_NR03 U606 ( .A0(xc_top.SFIFOLock2), .A1(xc_top.GFReset), .A2(moveForward), .Z(n6867));
Q_LDP0 \ififoXdataFinal_REG[254] ( .G(moveForwardN), .D(ififoXdata[254]), .Q(ififoXdataFinal[254]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[253] ( .G(moveForwardN), .D(ififoXdata[253]), .Q(ififoXdataFinal[253]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[252] ( .G(moveForwardN), .D(ififoXdata[252]), .Q(ififoXdataFinal[252]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[251] ( .G(moveForwardN), .D(ififoXdata[251]), .Q(ififoXdataFinal[251]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[250] ( .G(moveForwardN), .D(ififoXdata[250]), .Q(ififoXdataFinal[250]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[249] ( .G(moveForwardN), .D(ififoXdata[249]), .Q(ififoXdataFinal[249]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[248] ( .G(moveForwardN), .D(ififoXdata[248]), .Q(ififoXdataFinal[248]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[247] ( .G(moveForwardN), .D(ififoXdata[247]), .Q(ififoXdataFinal[247]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[246] ( .G(moveForwardN), .D(ififoXdata[246]), .Q(ififoXdataFinal[246]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[245] ( .G(moveForwardN), .D(ififoXdata[245]), .Q(ififoXdataFinal[245]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[244] ( .G(moveForwardN), .D(ififoXdata[244]), .Q(ififoXdataFinal[244]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[243] ( .G(moveForwardN), .D(ififoXdata[243]), .Q(ififoXdataFinal[243]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[242] ( .G(moveForwardN), .D(ififoXdata[242]), .Q(ififoXdataFinal[242]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[241] ( .G(moveForwardN), .D(ififoXdata[241]), .Q(ififoXdataFinal[241]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[240] ( .G(moveForwardN), .D(ififoXdata[240]), .Q(ififoXdataFinal[240]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[239] ( .G(moveForwardN), .D(ififoXdata[239]), .Q(ififoXdataFinal[239]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[238] ( .G(moveForwardN), .D(ififoXdata[238]), .Q(ififoXdataFinal[238]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[237] ( .G(moveForwardN), .D(ififoXdata[237]), .Q(ififoXdataFinal[237]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[236] ( .G(moveForwardN), .D(ififoXdata[236]), .Q(ififoXdataFinal[236]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[235] ( .G(moveForwardN), .D(ififoXdata[235]), .Q(ififoXdataFinal[235]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[234] ( .G(moveForwardN), .D(ififoXdata[234]), .Q(ififoXdataFinal[234]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[233] ( .G(moveForwardN), .D(ififoXdata[233]), .Q(ififoXdataFinal[233]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[232] ( .G(moveForwardN), .D(ififoXdata[232]), .Q(ififoXdataFinal[232]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[231] ( .G(moveForwardN), .D(ififoXdata[231]), .Q(ififoXdataFinal[231]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[230] ( .G(moveForwardN), .D(ififoXdata[230]), .Q(ififoXdataFinal[230]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[229] ( .G(moveForwardN), .D(ififoXdata[229]), .Q(ififoXdataFinal[229]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[228] ( .G(moveForwardN), .D(ififoXdata[228]), .Q(ififoXdataFinal[228]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[227] ( .G(moveForwardN), .D(ififoXdata[227]), .Q(ififoXdataFinal[227]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[226] ( .G(moveForwardN), .D(ififoXdata[226]), .Q(ififoXdataFinal[226]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[225] ( .G(moveForwardN), .D(ififoXdata[225]), .Q(ififoXdataFinal[225]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[224] ( .G(moveForwardN), .D(ififoXdata[224]), .Q(ififoXdataFinal[224]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[223] ( .G(moveForwardN), .D(ififoXdata[223]), .Q(ififoXdataFinal[223]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[222] ( .G(moveForwardN), .D(ififoXdata[222]), .Q(ififoXdataFinal[222]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[221] ( .G(moveForwardN), .D(ififoXdata[221]), .Q(ififoXdataFinal[221]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[220] ( .G(moveForwardN), .D(ififoXdata[220]), .Q(ififoXdataFinal[220]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[219] ( .G(moveForwardN), .D(ififoXdata[219]), .Q(ififoXdataFinal[219]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[218] ( .G(moveForwardN), .D(ififoXdata[218]), .Q(ififoXdataFinal[218]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[217] ( .G(moveForwardN), .D(ififoXdata[217]), .Q(ififoXdataFinal[217]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[216] ( .G(moveForwardN), .D(ififoXdata[216]), .Q(ififoXdataFinal[216]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[215] ( .G(moveForwardN), .D(ififoXdata[215]), .Q(ififoXdataFinal[215]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[214] ( .G(moveForwardN), .D(ififoXdata[214]), .Q(ififoXdataFinal[214]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[213] ( .G(moveForwardN), .D(ififoXdata[213]), .Q(ififoXdataFinal[213]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[212] ( .G(moveForwardN), .D(ififoXdata[212]), .Q(ififoXdataFinal[212]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[211] ( .G(moveForwardN), .D(ififoXdata[211]), .Q(ififoXdataFinal[211]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[210] ( .G(moveForwardN), .D(ififoXdata[210]), .Q(ififoXdataFinal[210]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[209] ( .G(moveForwardN), .D(ififoXdata[209]), .Q(ififoXdataFinal[209]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[208] ( .G(moveForwardN), .D(ififoXdata[208]), .Q(ififoXdataFinal[208]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[207] ( .G(moveForwardN), .D(ififoXdata[207]), .Q(ififoXdataFinal[207]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[206] ( .G(moveForwardN), .D(ififoXdata[206]), .Q(ififoXdataFinal[206]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[205] ( .G(moveForwardN), .D(ififoXdata[205]), .Q(ififoXdataFinal[205]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[204] ( .G(moveForwardN), .D(ififoXdata[204]), .Q(ififoXdataFinal[204]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[203] ( .G(moveForwardN), .D(ififoXdata[203]), .Q(ififoXdataFinal[203]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[202] ( .G(moveForwardN), .D(ififoXdata[202]), .Q(ififoXdataFinal[202]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[201] ( .G(moveForwardN), .D(ififoXdata[201]), .Q(ififoXdataFinal[201]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[200] ( .G(moveForwardN), .D(ififoXdata[200]), .Q(ififoXdataFinal[200]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[199] ( .G(moveForwardN), .D(ififoXdata[199]), .Q(ififoXdataFinal[199]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[198] ( .G(moveForwardN), .D(ififoXdata[198]), .Q(ififoXdataFinal[198]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[197] ( .G(moveForwardN), .D(ififoXdata[197]), .Q(ififoXdataFinal[197]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[196] ( .G(moveForwardN), .D(ififoXdata[196]), .Q(ififoXdataFinal[196]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[195] ( .G(moveForwardN), .D(ififoXdata[195]), .Q(ififoXdataFinal[195]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[194] ( .G(moveForwardN), .D(ififoXdata[194]), .Q(ififoXdataFinal[194]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[193] ( .G(moveForwardN), .D(ififoXdata[193]), .Q(ififoXdataFinal[193]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[192] ( .G(moveForwardN), .D(ififoXdata[192]), .Q(ififoXdataFinal[192]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[190] ( .G(moveForwardN), .D(ififoXdata[190]), .Q(ififoXdataFinal[190]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[189] ( .G(moveForwardN), .D(ififoXdata[189]), .Q(ififoXdataFinal[189]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[188] ( .G(moveForwardN), .D(ififoXdata[188]), .Q(ififoXdataFinal[188]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[187] ( .G(moveForwardN), .D(ififoXdata[187]), .Q(ififoXdataFinal[187]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[186] ( .G(moveForwardN), .D(ififoXdata[186]), .Q(ififoXdataFinal[186]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[185] ( .G(moveForwardN), .D(ififoXdata[185]), .Q(ififoXdataFinal[185]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[184] ( .G(moveForwardN), .D(ififoXdata[184]), .Q(ififoXdataFinal[184]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[183] ( .G(moveForwardN), .D(ififoXdata[183]), .Q(ififoXdataFinal[183]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[182] ( .G(moveForwardN), .D(ififoXdata[182]), .Q(ififoXdataFinal[182]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[181] ( .G(moveForwardN), .D(ififoXdata[181]), .Q(ififoXdataFinal[181]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[180] ( .G(moveForwardN), .D(ififoXdata[180]), .Q(ififoXdataFinal[180]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[179] ( .G(moveForwardN), .D(ififoXdata[179]), .Q(ififoXdataFinal[179]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[178] ( .G(moveForwardN), .D(ififoXdata[178]), .Q(ififoXdataFinal[178]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[177] ( .G(moveForwardN), .D(ififoXdata[177]), .Q(ififoXdataFinal[177]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[176] ( .G(moveForwardN), .D(ififoXdata[176]), .Q(ififoXdataFinal[176]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[175] ( .G(moveForwardN), .D(ififoXdata[175]), .Q(ififoXdataFinal[175]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[174] ( .G(moveForwardN), .D(ififoXdata[174]), .Q(ififoXdataFinal[174]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[173] ( .G(moveForwardN), .D(ififoXdata[173]), .Q(ififoXdataFinal[173]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[172] ( .G(moveForwardN), .D(ififoXdata[172]), .Q(ififoXdataFinal[172]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[171] ( .G(moveForwardN), .D(ififoXdata[171]), .Q(ififoXdataFinal[171]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[170] ( .G(moveForwardN), .D(ififoXdata[170]), .Q(ififoXdataFinal[170]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[169] ( .G(moveForwardN), .D(ififoXdata[169]), .Q(ififoXdataFinal[169]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[168] ( .G(moveForwardN), .D(ififoXdata[168]), .Q(ififoXdataFinal[168]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[167] ( .G(moveForwardN), .D(ififoXdata[167]), .Q(ififoXdataFinal[167]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[166] ( .G(moveForwardN), .D(ififoXdata[166]), .Q(ififoXdataFinal[166]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[165] ( .G(moveForwardN), .D(ififoXdata[165]), .Q(ififoXdataFinal[165]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[164] ( .G(moveForwardN), .D(ififoXdata[164]), .Q(ififoXdataFinal[164]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[163] ( .G(moveForwardN), .D(ififoXdata[163]), .Q(ififoXdataFinal[163]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[162] ( .G(moveForwardN), .D(ififoXdata[162]), .Q(ififoXdataFinal[162]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[161] ( .G(moveForwardN), .D(ififoXdata[161]), .Q(ififoXdataFinal[161]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[160] ( .G(moveForwardN), .D(ififoXdata[160]), .Q(ififoXdataFinal[160]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[159] ( .G(moveForwardN), .D(ififoXdata[159]), .Q(ififoXdataFinal[159]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[158] ( .G(moveForwardN), .D(ififoXdata[158]), .Q(ififoXdataFinal[158]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[157] ( .G(moveForwardN), .D(ififoXdata[157]), .Q(ififoXdataFinal[157]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[156] ( .G(moveForwardN), .D(ififoXdata[156]), .Q(ififoXdataFinal[156]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[155] ( .G(moveForwardN), .D(ififoXdata[155]), .Q(ififoXdataFinal[155]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[154] ( .G(moveForwardN), .D(ififoXdata[154]), .Q(ififoXdataFinal[154]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[153] ( .G(moveForwardN), .D(ififoXdata[153]), .Q(ififoXdataFinal[153]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[152] ( .G(moveForwardN), .D(ififoXdata[152]), .Q(ififoXdataFinal[152]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[151] ( .G(moveForwardN), .D(ififoXdata[151]), .Q(ififoXdataFinal[151]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[150] ( .G(moveForwardN), .D(ififoXdata[150]), .Q(ififoXdataFinal[150]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[149] ( .G(moveForwardN), .D(ififoXdata[149]), .Q(ififoXdataFinal[149]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[148] ( .G(moveForwardN), .D(ififoXdata[148]), .Q(ififoXdataFinal[148]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[147] ( .G(moveForwardN), .D(ififoXdata[147]), .Q(ififoXdataFinal[147]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[146] ( .G(moveForwardN), .D(ififoXdata[146]), .Q(ififoXdataFinal[146]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[145] ( .G(moveForwardN), .D(ififoXdata[145]), .Q(ififoXdataFinal[145]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[144] ( .G(moveForwardN), .D(ififoXdata[144]), .Q(ififoXdataFinal[144]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[143] ( .G(moveForwardN), .D(ififoXdata[143]), .Q(ififoXdataFinal[143]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[142] ( .G(moveForwardN), .D(ififoXdata[142]), .Q(ififoXdataFinal[142]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[141] ( .G(moveForwardN), .D(ififoXdata[141]), .Q(ififoXdataFinal[141]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[140] ( .G(moveForwardN), .D(ififoXdata[140]), .Q(ififoXdataFinal[140]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[139] ( .G(moveForwardN), .D(ififoXdata[139]), .Q(ififoXdataFinal[139]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[138] ( .G(moveForwardN), .D(ififoXdata[138]), .Q(ififoXdataFinal[138]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[137] ( .G(moveForwardN), .D(ififoXdata[137]), .Q(ififoXdataFinal[137]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[136] ( .G(moveForwardN), .D(ififoXdata[136]), .Q(ififoXdataFinal[136]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[135] ( .G(moveForwardN), .D(ififoXdata[135]), .Q(ififoXdataFinal[135]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[134] ( .G(moveForwardN), .D(ififoXdata[134]), .Q(ififoXdataFinal[134]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[133] ( .G(moveForwardN), .D(ififoXdata[133]), .Q(ififoXdataFinal[133]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[132] ( .G(moveForwardN), .D(ififoXdata[132]), .Q(ififoXdataFinal[132]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[131] ( .G(moveForwardN), .D(ififoXdata[131]), .Q(ififoXdataFinal[131]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[130] ( .G(moveForwardN), .D(ififoXdata[130]), .Q(ififoXdataFinal[130]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[129] ( .G(moveForwardN), .D(ififoXdata[129]), .Q(ififoXdataFinal[129]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[128] ( .G(moveForwardN), .D(ififoXdata[128]), .Q(ififoXdataFinal[128]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[126] ( .G(moveForwardN), .D(ififoXdata[126]), .Q(ififoXdataFinal[126]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[125] ( .G(moveForwardN), .D(ififoXdata[125]), .Q(ififoXdataFinal[125]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[124] ( .G(moveForwardN), .D(ififoXdata[124]), .Q(ififoXdataFinal[124]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[123] ( .G(moveForwardN), .D(ififoXdata[123]), .Q(ififoXdataFinal[123]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[122] ( .G(moveForwardN), .D(ififoXdata[122]), .Q(ififoXdataFinal[122]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[121] ( .G(moveForwardN), .D(ififoXdata[121]), .Q(ififoXdataFinal[121]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[120] ( .G(moveForwardN), .D(ififoXdata[120]), .Q(ififoXdataFinal[120]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[119] ( .G(moveForwardN), .D(ififoXdata[119]), .Q(ififoXdataFinal[119]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[118] ( .G(moveForwardN), .D(ififoXdata[118]), .Q(ififoXdataFinal[118]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[117] ( .G(moveForwardN), .D(ififoXdata[117]), .Q(ififoXdataFinal[117]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[116] ( .G(moveForwardN), .D(ififoXdata[116]), .Q(ififoXdataFinal[116]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[115] ( .G(moveForwardN), .D(ififoXdata[115]), .Q(ififoXdataFinal[115]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[114] ( .G(moveForwardN), .D(ififoXdata[114]), .Q(ififoXdataFinal[114]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[113] ( .G(moveForwardN), .D(ififoXdata[113]), .Q(ififoXdataFinal[113]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[112] ( .G(moveForwardN), .D(ififoXdata[112]), .Q(ififoXdataFinal[112]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[111] ( .G(moveForwardN), .D(ififoXdata[111]), .Q(ififoXdataFinal[111]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[110] ( .G(moveForwardN), .D(ififoXdata[110]), .Q(ififoXdataFinal[110]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[109] ( .G(moveForwardN), .D(ififoXdata[109]), .Q(ififoXdataFinal[109]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[108] ( .G(moveForwardN), .D(ififoXdata[108]), .Q(ififoXdataFinal[108]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[107] ( .G(moveForwardN), .D(ififoXdata[107]), .Q(ififoXdataFinal[107]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[106] ( .G(moveForwardN), .D(ififoXdata[106]), .Q(ififoXdataFinal[106]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[105] ( .G(moveForwardN), .D(ififoXdata[105]), .Q(ififoXdataFinal[105]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[104] ( .G(moveForwardN), .D(ififoXdata[104]), .Q(ififoXdataFinal[104]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[103] ( .G(moveForwardN), .D(ififoXdata[103]), .Q(ififoXdataFinal[103]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[102] ( .G(moveForwardN), .D(ififoXdata[102]), .Q(ififoXdataFinal[102]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[101] ( .G(moveForwardN), .D(ififoXdata[101]), .Q(ififoXdataFinal[101]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[100] ( .G(moveForwardN), .D(ififoXdata[100]), .Q(ififoXdataFinal[100]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[99] ( .G(moveForwardN), .D(ififoXdata[99]), .Q(ififoXdataFinal[99]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[98] ( .G(moveForwardN), .D(ififoXdata[98]), .Q(ififoXdataFinal[98]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[97] ( .G(moveForwardN), .D(ififoXdata[97]), .Q(ififoXdataFinal[97]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[96] ( .G(moveForwardN), .D(ififoXdata[96]), .Q(ififoXdataFinal[96]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[95] ( .G(moveForwardN), .D(ififoXdata[95]), .Q(ififoXdataFinal[95]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[94] ( .G(moveForwardN), .D(ififoXdata[94]), .Q(ififoXdataFinal[94]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[93] ( .G(moveForwardN), .D(ififoXdata[93]), .Q(ififoXdataFinal[93]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[92] ( .G(moveForwardN), .D(ififoXdata[92]), .Q(ififoXdataFinal[92]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[91] ( .G(moveForwardN), .D(ififoXdata[91]), .Q(ififoXdataFinal[91]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[90] ( .G(moveForwardN), .D(ififoXdata[90]), .Q(ififoXdataFinal[90]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[89] ( .G(moveForwardN), .D(ififoXdata[89]), .Q(ififoXdataFinal[89]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[88] ( .G(moveForwardN), .D(ififoXdata[88]), .Q(ififoXdataFinal[88]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[87] ( .G(moveForwardN), .D(ififoXdata[87]), .Q(ififoXdataFinal[87]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[86] ( .G(moveForwardN), .D(ififoXdata[86]), .Q(ififoXdataFinal[86]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[85] ( .G(moveForwardN), .D(ififoXdata[85]), .Q(ififoXdataFinal[85]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[84] ( .G(moveForwardN), .D(ififoXdata[84]), .Q(ififoXdataFinal[84]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[83] ( .G(moveForwardN), .D(ififoXdata[83]), .Q(ififoXdataFinal[83]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[82] ( .G(moveForwardN), .D(ififoXdata[82]), .Q(ififoXdataFinal[82]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[81] ( .G(moveForwardN), .D(ififoXdata[81]), .Q(ififoXdataFinal[81]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[80] ( .G(moveForwardN), .D(ififoXdata[80]), .Q(ififoXdataFinal[80]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[79] ( .G(moveForwardN), .D(ififoXdata[79]), .Q(ififoXdataFinal[79]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[78] ( .G(moveForwardN), .D(ififoXdata[78]), .Q(ififoXdataFinal[78]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[77] ( .G(moveForwardN), .D(ififoXdata[77]), .Q(ififoXdataFinal[77]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[76] ( .G(moveForwardN), .D(ififoXdata[76]), .Q(ififoXdataFinal[76]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[75] ( .G(moveForwardN), .D(ififoXdata[75]), .Q(ififoXdataFinal[75]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[74] ( .G(moveForwardN), .D(ififoXdata[74]), .Q(ififoXdataFinal[74]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[73] ( .G(moveForwardN), .D(ififoXdata[73]), .Q(ififoXdataFinal[73]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[72] ( .G(moveForwardN), .D(ififoXdata[72]), .Q(ififoXdataFinal[72]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[71] ( .G(moveForwardN), .D(ififoXdata[71]), .Q(ififoXdataFinal[71]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[70] ( .G(moveForwardN), .D(ififoXdata[70]), .Q(ififoXdataFinal[70]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[69] ( .G(moveForwardN), .D(ififoXdata[69]), .Q(ififoXdataFinal[69]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[68] ( .G(moveForwardN), .D(ififoXdata[68]), .Q(ififoXdataFinal[68]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[67] ( .G(moveForwardN), .D(ififoXdata[67]), .Q(ififoXdataFinal[67]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[66] ( .G(moveForwardN), .D(ififoXdata[66]), .Q(ififoXdataFinal[66]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[65] ( .G(moveForwardN), .D(ififoXdata[65]), .Q(ififoXdataFinal[65]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[64] ( .G(moveForwardN), .D(ififoXdata[64]), .Q(ififoXdataFinal[64]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[62] ( .G(moveForwardN), .D(ififoXdata[62]), .Q(ififoXdataFinal[62]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[61] ( .G(moveForwardN), .D(ififoXdata[61]), .Q(ififoXdataFinal[61]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[60] ( .G(moveForwardN), .D(ififoXdata[60]), .Q(ififoXdataFinal[60]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[59] ( .G(moveForwardN), .D(ififoXdata[59]), .Q(ififoXdataFinal[59]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[58] ( .G(moveForwardN), .D(ififoXdata[58]), .Q(ififoXdataFinal[58]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[57] ( .G(moveForwardN), .D(ififoXdata[57]), .Q(ififoXdataFinal[57]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[56] ( .G(moveForwardN), .D(ififoXdata[56]), .Q(ififoXdataFinal[56]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[55] ( .G(moveForwardN), .D(ififoXdata[55]), .Q(ififoXdataFinal[55]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[54] ( .G(moveForwardN), .D(ififoXdata[54]), .Q(ififoXdataFinal[54]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[53] ( .G(moveForwardN), .D(ififoXdata[53]), .Q(ififoXdataFinal[53]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[52] ( .G(moveForwardN), .D(ififoXdata[52]), .Q(ififoXdataFinal[52]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[51] ( .G(moveForwardN), .D(ififoXdata[51]), .Q(ififoXdataFinal[51]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[50] ( .G(moveForwardN), .D(ififoXdata[50]), .Q(ififoXdataFinal[50]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[49] ( .G(moveForwardN), .D(ififoXdata[49]), .Q(ififoXdataFinal[49]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[48] ( .G(moveForwardN), .D(ififoXdata[48]), .Q(ififoXdataFinal[48]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[47] ( .G(moveForwardN), .D(ififoXdata[47]), .Q(ififoXdataFinal[47]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[46] ( .G(moveForwardN), .D(ififoXdata[46]), .Q(ififoXdataFinal[46]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[45] ( .G(moveForwardN), .D(ififoXdata[45]), .Q(ififoXdataFinal[45]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[44] ( .G(moveForwardN), .D(ififoXdata[44]), .Q(ififoXdataFinal[44]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[43] ( .G(moveForwardN), .D(ififoXdata[43]), .Q(ififoXdataFinal[43]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[42] ( .G(moveForwardN), .D(ififoXdata[42]), .Q(ififoXdataFinal[42]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[41] ( .G(moveForwardN), .D(ififoXdata[41]), .Q(ififoXdataFinal[41]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[40] ( .G(moveForwardN), .D(ififoXdata[40]), .Q(ififoXdataFinal[40]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[39] ( .G(moveForwardN), .D(ififoXdata[39]), .Q(ififoXdataFinal[39]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[38] ( .G(moveForwardN), .D(ififoXdata[38]), .Q(ififoXdataFinal[38]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[37] ( .G(moveForwardN), .D(ififoXdata[37]), .Q(ififoXdataFinal[37]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[36] ( .G(moveForwardN), .D(ififoXdata[36]), .Q(ififoXdataFinal[36]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[35] ( .G(moveForwardN), .D(ififoXdata[35]), .Q(ififoXdataFinal[35]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[34] ( .G(moveForwardN), .D(ififoXdata[34]), .Q(ififoXdataFinal[34]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[33] ( .G(moveForwardN), .D(ififoXdata[33]), .Q(ififoXdataFinal[33]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[32] ( .G(moveForwardN), .D(ififoXdata[32]), .Q(ififoXdataFinal[32]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[31] ( .G(moveForwardN), .D(ififoXdata[31]), .Q(ififoXdataFinal[31]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[30] ( .G(moveForwardN), .D(ififoXdata[30]), .Q(ififoXdataFinal[30]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[29] ( .G(moveForwardN), .D(ififoXdata[29]), .Q(ififoXdataFinal[29]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[28] ( .G(moveForwardN), .D(ififoXdata[28]), .Q(ififoXdataFinal[28]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[27] ( .G(moveForwardN), .D(ififoXdata[27]), .Q(ififoXdataFinal[27]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[26] ( .G(moveForwardN), .D(ififoXdata[26]), .Q(ififoXdataFinal[26]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[25] ( .G(moveForwardN), .D(ififoXdata[25]), .Q(ififoXdataFinal[25]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[24] ( .G(moveForwardN), .D(ififoXdata[24]), .Q(ififoXdataFinal[24]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[23] ( .G(moveForwardN), .D(ififoXdata[23]), .Q(ififoXdataFinal[23]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[22] ( .G(moveForwardN), .D(ififoXdata[22]), .Q(ififoXdataFinal[22]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[21] ( .G(moveForwardN), .D(ififoXdata[21]), .Q(ififoXdataFinal[21]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[20] ( .G(moveForwardN), .D(ififoXdata[20]), .Q(ififoXdataFinal[20]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[19] ( .G(moveForwardN), .D(ififoXdata[19]), .Q(ififoXdataFinal[19]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[18] ( .G(moveForwardN), .D(ififoXdata[18]), .Q(ififoXdataFinal[18]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[17] ( .G(moveForwardN), .D(ififoXdata[17]), .Q(ififoXdataFinal[17]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[16] ( .G(moveForwardN), .D(ififoXdata[16]), .Q(ififoXdataFinal[16]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[15] ( .G(moveForwardN), .D(ififoXdata[15]), .Q(ififoXdataFinal[15]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[14] ( .G(moveForwardN), .D(ififoXdata[14]), .Q(ififoXdataFinal[14]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[13] ( .G(moveForwardN), .D(ififoXdata[13]), .Q(ififoXdataFinal[13]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[12] ( .G(moveForwardN), .D(ififoXdata[12]), .Q(ififoXdataFinal[12]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[11] ( .G(moveForwardN), .D(ififoXdata[11]), .Q(ififoXdataFinal[11]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[10] ( .G(moveForwardN), .D(ififoXdata[10]), .Q(ififoXdataFinal[10]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[9] ( .G(moveForwardN), .D(ififoXdata[9]), .Q(ififoXdataFinal[9]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[8] ( .G(moveForwardN), .D(ififoXdata[8]), .Q(ififoXdataFinal[8]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[7] ( .G(moveForwardN), .D(ififoXdata[7]), .Q(ififoXdataFinal[7]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[6] ( .G(moveForwardN), .D(ififoXdata[6]), .Q(ififoXdataFinal[6]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[5] ( .G(moveForwardN), .D(ififoXdata[5]), .Q(ififoXdataFinal[5]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[4] ( .G(moveForwardN), .D(ififoXdata[4]), .Q(ififoXdataFinal[4]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[3] ( .G(moveForwardN), .D(ififoXdata[3]), .Q(ififoXdataFinal[3]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[2] ( .G(moveForwardN), .D(ififoXdata[2]), .Q(ififoXdataFinal[2]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[1] ( .G(moveForwardN), .D(ififoXdata[1]), .Q(ififoXdataFinal[1]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[0] ( .G(moveForwardN), .D(ififoXdata[0]), .Q(ififoXdataFinal[0]), .QN( ));
Q_MX04 U859 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[0]), .A1(ififoXdata[64]), .A2(ififoXdata[128]), .A3(ififoXdata[192]), .Z(xval[0]));
Q_MX04 U860 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[1]), .A1(ififoXdata[65]), .A2(ififoXdata[129]), .A3(ififoXdata[193]), .Z(xval[1]));
Q_MX04 U861 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[2]), .A1(ififoXdata[66]), .A2(ififoXdata[130]), .A3(ififoXdata[194]), .Z(xval[2]));
Q_MX04 U862 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[3]), .A1(ififoXdata[67]), .A2(ififoXdata[131]), .A3(ififoXdata[195]), .Z(xval[3]));
Q_MX04 U863 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[4]), .A1(ififoXdata[68]), .A2(ififoXdata[132]), .A3(ififoXdata[196]), .Z(xval[4]));
Q_MX04 U864 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[5]), .A1(ififoXdata[69]), .A2(ififoXdata[133]), .A3(ififoXdata[197]), .Z(xval[5]));
Q_MX04 U865 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[6]), .A1(ififoXdata[70]), .A2(ififoXdata[134]), .A3(ififoXdata[198]), .Z(xval[6]));
Q_MX04 U866 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[7]), .A1(ififoXdata[71]), .A2(ififoXdata[135]), .A3(ififoXdata[199]), .Z(xval[7]));
Q_MX04 U867 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[8]), .A1(ififoXdata[72]), .A2(ififoXdata[136]), .A3(ififoXdata[200]), .Z(xval[8]));
Q_MX04 U868 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[9]), .A1(ififoXdata[73]), .A2(ififoXdata[137]), .A3(ififoXdata[201]), .Z(xval[9]));
Q_MX04 U869 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[10]), .A1(ififoXdata[74]), .A2(ififoXdata[138]), .A3(ififoXdata[202]), .Z(xval[10]));
Q_MX04 U870 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[11]), .A1(ififoXdata[75]), .A2(ififoXdata[139]), .A3(ififoXdata[203]), .Z(xval[11]));
Q_MX04 U871 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[12]), .A1(ififoXdata[76]), .A2(ififoXdata[140]), .A3(ififoXdata[204]), .Z(xval[12]));
Q_MX04 U872 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[13]), .A1(ififoXdata[77]), .A2(ififoXdata[141]), .A3(ififoXdata[205]), .Z(xval[13]));
Q_MX04 U873 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[14]), .A1(ififoXdata[78]), .A2(ififoXdata[142]), .A3(ififoXdata[206]), .Z(xval[14]));
Q_MX04 U874 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[15]), .A1(ififoXdata[79]), .A2(ififoXdata[143]), .A3(ififoXdata[207]), .Z(xval[15]));
Q_MX04 U875 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[16]), .A1(ififoXdata[80]), .A2(ififoXdata[144]), .A3(ififoXdata[208]), .Z(xval[16]));
Q_MX04 U876 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[17]), .A1(ififoXdata[81]), .A2(ififoXdata[145]), .A3(ififoXdata[209]), .Z(xval[17]));
Q_MX04 U877 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[18]), .A1(ififoXdata[82]), .A2(ififoXdata[146]), .A3(ififoXdata[210]), .Z(xval[18]));
Q_MX04 U878 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[19]), .A1(ififoXdata[83]), .A2(ififoXdata[147]), .A3(ififoXdata[211]), .Z(xval[19]));
Q_MX04 U879 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[20]), .A1(ififoXdata[84]), .A2(ififoXdata[148]), .A3(ififoXdata[212]), .Z(xval[20]));
Q_MX04 U880 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[21]), .A1(ififoXdata[85]), .A2(ififoXdata[149]), .A3(ififoXdata[213]), .Z(xval[21]));
Q_MX04 U881 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[22]), .A1(ififoXdata[86]), .A2(ififoXdata[150]), .A3(ififoXdata[214]), .Z(xval[22]));
Q_MX04 U882 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[23]), .A1(ififoXdata[87]), .A2(ififoXdata[151]), .A3(ififoXdata[215]), .Z(xval[23]));
Q_MX04 U883 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[24]), .A1(ififoXdata[88]), .A2(ififoXdata[152]), .A3(ififoXdata[216]), .Z(xval[24]));
Q_MX04 U884 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[25]), .A1(ififoXdata[89]), .A2(ififoXdata[153]), .A3(ififoXdata[217]), .Z(xval[25]));
Q_MX04 U885 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[26]), .A1(ififoXdata[90]), .A2(ififoXdata[154]), .A3(ififoXdata[218]), .Z(xval[26]));
Q_MX04 U886 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[27]), .A1(ififoXdata[91]), .A2(ififoXdata[155]), .A3(ififoXdata[219]), .Z(xval[27]));
Q_MX04 U887 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[28]), .A1(ififoXdata[92]), .A2(ififoXdata[156]), .A3(ififoXdata[220]), .Z(xval[28]));
Q_MX04 U888 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[29]), .A1(ififoXdata[93]), .A2(ififoXdata[157]), .A3(ififoXdata[221]), .Z(xval[29]));
Q_MX04 U889 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[30]), .A1(ififoXdata[94]), .A2(ififoXdata[158]), .A3(ififoXdata[222]), .Z(xval[30]));
Q_MX04 U890 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[31]), .A1(ififoXdata[95]), .A2(ififoXdata[159]), .A3(ififoXdata[223]), .Z(xval[31]));
Q_MX04 U891 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[32]), .A1(ififoXdata[96]), .A2(ififoXdata[160]), .A3(ififoXdata[224]), .Z(dataBits[0]));
Q_MX04 U892 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[33]), .A1(ififoXdata[97]), .A2(ififoXdata[161]), .A3(ififoXdata[225]), .Z(dataBits[1]));
Q_MX04 U893 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[34]), .A1(ififoXdata[98]), .A2(ififoXdata[162]), .A3(ififoXdata[226]), .Z(dataBits[2]));
Q_MX04 U894 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[35]), .A1(ififoXdata[99]), .A2(ififoXdata[163]), .A3(ififoXdata[227]), .Z(dataBits[3]));
Q_MX04 U895 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[36]), .A1(ififoXdata[100]), .A2(ififoXdata[164]), .A3(ififoXdata[228]), .Z(xval[36]));
Q_MX04 U896 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[37]), .A1(ififoXdata[101]), .A2(ififoXdata[165]), .A3(ififoXdata[229]), .Z(xval[37]));
Q_MX04 U897 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[38]), .A1(ififoXdata[102]), .A2(ififoXdata[166]), .A3(ififoXdata[230]), .Z(xval[38]));
Q_MX04 U898 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[39]), .A1(ififoXdata[103]), .A2(ififoXdata[167]), .A3(ififoXdata[231]), .Z(xval[39]));
Q_MX04 U899 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[40]), .A1(ififoXdata[104]), .A2(ififoXdata[168]), .A3(ififoXdata[232]), .Z(xval[40]));
Q_MX04 U900 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[41]), .A1(ififoXdata[105]), .A2(ififoXdata[169]), .A3(ififoXdata[233]), .Z(xval[41]));
Q_MX04 U901 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[42]), .A1(ififoXdata[106]), .A2(ififoXdata[170]), .A3(ififoXdata[234]), .Z(xval[42]));
Q_MX04 U902 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[43]), .A1(ififoXdata[107]), .A2(ififoXdata[171]), .A3(ififoXdata[235]), .Z(xval[43]));
Q_MX04 U903 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[44]), .A1(ififoXdata[108]), .A2(ififoXdata[172]), .A3(ififoXdata[236]), .Z(xval[44]));
Q_MX04 U904 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[45]), .A1(ififoXdata[109]), .A2(ififoXdata[173]), .A3(ififoXdata[237]), .Z(xval[45]));
Q_MX04 U905 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[46]), .A1(ififoXdata[110]), .A2(ififoXdata[174]), .A3(ififoXdata[238]), .Z(xval[46]));
Q_MX04 U906 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[47]), .A1(ififoXdata[111]), .A2(ififoXdata[175]), .A3(ififoXdata[239]), .Z(xval[47]));
Q_MX04 U907 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[48]), .A1(ififoXdata[112]), .A2(ififoXdata[176]), .A3(ififoXdata[240]), .Z(xval[48]));
Q_MX04 U908 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[49]), .A1(ififoXdata[113]), .A2(ififoXdata[177]), .A3(ififoXdata[241]), .Z(xval[49]));
Q_MX04 U909 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[50]), .A1(ififoXdata[114]), .A2(ififoXdata[178]), .A3(ififoXdata[242]), .Z(xval[50]));
Q_MX04 U910 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[51]), .A1(ififoXdata[115]), .A2(ififoXdata[179]), .A3(ififoXdata[243]), .Z(xval[51]));
Q_MX04 U911 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[52]), .A1(ififoXdata[116]), .A2(ififoXdata[180]), .A3(ififoXdata[244]), .Z(xval[52]));
Q_MX04 U912 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[53]), .A1(ififoXdata[117]), .A2(ififoXdata[181]), .A3(ififoXdata[245]), .Z(xval[53]));
Q_MX04 U913 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[54]), .A1(ififoXdata[118]), .A2(ififoXdata[182]), .A3(ififoXdata[246]), .Z(xval[54]));
Q_MX04 U914 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[55]), .A1(ififoXdata[119]), .A2(ififoXdata[183]), .A3(ififoXdata[247]), .Z(xval[55]));
Q_MX04 U915 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[56]), .A1(ififoXdata[120]), .A2(ififoXdata[184]), .A3(ififoXdata[248]), .Z(xval[56]));
Q_MX04 U916 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[57]), .A1(ififoXdata[121]), .A2(ififoXdata[185]), .A3(ififoXdata[249]), .Z(xval[57]));
Q_MX04 U917 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[58]), .A1(ififoXdata[122]), .A2(ififoXdata[186]), .A3(ififoXdata[250]), .Z(xval[58]));
Q_MX04 U918 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[59]), .A1(ififoXdata[123]), .A2(ififoXdata[187]), .A3(ififoXdata[251]), .Z(xval[59]));
Q_MX04 U919 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[60]), .A1(ififoXdata[124]), .A2(ififoXdata[188]), .A3(ififoXdata[252]), .Z(xval[60]));
Q_MX04 U920 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[61]), .A1(ififoXdata[125]), .A2(ififoXdata[189]), .A3(ififoXdata[253]), .Z(xval[61]));
Q_MX04 U921 ( .S0(xptr[0]), .S1(xptr[1]), .A0(ififoXdata[62]), .A1(ififoXdata[126]), .A2(ififoXdata[190]), .A3(ififoXdata[254]), .Z(xval[62]));
Q_MX04 U922 ( .S0(xptr[0]), .S1(xptr[1]), .A0(newMarkBits[0]), .A1(newMarkBits[1]), .A2(newMarkBits[2]), .A3(newMarkBits[3]), .Z(xval[63]));
Q_LDP0 \ififoXdataFinal_REG[255] ( .G(moveForwardN), .D(xval[35]), .Q(ififoXdataFinal[255]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[191] ( .G(moveForwardN), .D(xval[34]), .Q(ififoXdataFinal[191]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[127] ( .G(moveForwardN), .D(xval[33]), .Q(ififoXdataFinal[127]), .QN( ));
Q_LDP0 \ififoXdataFinal_REG[63] ( .G(moveForwardN), .D(xval[32]), .Q(ififoXdataFinal[63]), .QN( ));
Q_MX02 U927 ( .S(moveForward), .A0(markBits[0]), .A1(xval[0]), .Z(markBitsN[0]));
Q_MX02 U928 ( .S(moveForward), .A0(markBits[1]), .A1(xval[1]), .Z(markBitsN[1]));
Q_MX02 U929 ( .S(moveForward), .A0(markBits[2]), .A1(xval[2]), .Z(markBitsN[2]));
Q_MX02 U930 ( .S(moveForward), .A0(markBits[3]), .A1(xval[3]), .Z(markBitsN[3]));
Q_MX02 U931 ( .S(moveForward), .A0(xptr[0]), .A1(xval[40]), .Z(xptrN[0]));
Q_MX02 U932 ( .S(moveForward), .A0(xptr[1]), .A1(xval[41]), .Z(xptrN[1]));
Q_MX02 U933 ( .S(moveForward), .A0(xptr[2]), .A1(xval[42]), .Z(xptrN[2]));
Q_MX02 U934 ( .S(moveForward), .A0(xptr[3]), .A1(xval[43]), .Z(xptrN[3]));
Q_MX02 U935 ( .S(moveForward), .A0(xptr[4]), .A1(xval[44]), .Z(xptrN[4]));
Q_MX02 U936 ( .S(moveForward), .A0(xptr[5]), .A1(xval[45]), .Z(xptrN[5]));
Q_MX02 U937 ( .S(moveForward), .A0(xptr[6]), .A1(xval[46]), .Z(xptrN[6]));
Q_MX02 U938 ( .S(moveForward), .A0(xptr[7]), .A1(xval[47]), .Z(xptrN[7]));
Q_MX02 U939 ( .S(moveForward), .A0(xptr[8]), .A1(xval[48]), .Z(xptrN[8]));
Q_MX02 U940 ( .S(moveForward), .A0(xptr[9]), .A1(xval[49]), .Z(xptrN[9]));
Q_MX02 U941 ( .S(moveForward), .A0(xptr[10]), .A1(xval[50]), .Z(xptrN[10]));
Q_MX02 U942 ( .S(moveForward), .A0(xptr[11]), .A1(xval[51]), .Z(xptrN[11]));
Q_MX02 U943 ( .S(moveForward), .A0(xptr[12]), .A1(xval[52]), .Z(xptrN[12]));
Q_MX02 U944 ( .S(moveForward), .A0(xptr[13]), .A1(xval[53]), .Z(xptrN[13]));
Q_MX02 U945 ( .S(moveForward), .A0(xptr[14]), .A1(xval[54]), .Z(xptrN[14]));
Q_MX02 U946 ( .S(moveForward), .A0(xptr[15]), .A1(xval[55]), .Z(xptrN[15]));
Q_MX02 U947 ( .S(moveForward), .A0(xptr[16]), .A1(xval[56]), .Z(xptrN[16]));
Q_MX02 U948 ( .S(moveForward), .A0(wptr[0]), .A1(xptr[0]), .Z(wptrN[0]));
Q_MX02 U949 ( .S(moveForward), .A0(wptr[1]), .A1(xptr[1]), .Z(wptrN[1]));
Q_MX02 U950 ( .S(moveForward), .A0(wptr[2]), .A1(xptr[2]), .Z(wptrN[2]));
Q_MX02 U951 ( .S(moveForward), .A0(wptr[3]), .A1(xptr[3]), .Z(wptrN[3]));
Q_MX02 U952 ( .S(moveForward), .A0(wptr[4]), .A1(xptr[4]), .Z(wptrN[4]));
Q_MX02 U953 ( .S(moveForward), .A0(wptr[5]), .A1(xptr[5]), .Z(wptrN[5]));
Q_MX02 U954 ( .S(moveForward), .A0(wptr[6]), .A1(xptr[6]), .Z(wptrN[6]));
Q_MX02 U955 ( .S(moveForward), .A0(wptr[7]), .A1(xptr[7]), .Z(wptrN[7]));
Q_MX02 U956 ( .S(moveForward), .A0(wptr[8]), .A1(xptr[8]), .Z(wptrN[8]));
Q_MX02 U957 ( .S(moveForward), .A0(wptr[9]), .A1(xptr[9]), .Z(wptrN[9]));
Q_MX02 U958 ( .S(moveForward), .A0(wptr[10]), .A1(xptr[10]), .Z(wptrN[10]));
Q_MX02 U959 ( .S(moveForward), .A0(wptr[11]), .A1(xptr[11]), .Z(wptrN[11]));
Q_MX02 U960 ( .S(moveForward), .A0(wptr[12]), .A1(xptr[12]), .Z(wptrN[12]));
Q_MX02 U961 ( .S(moveForward), .A0(wptr[13]), .A1(xptr[13]), .Z(wptrN[13]));
Q_MX02 U962 ( .S(moveForward), .A0(wptr[14]), .A1(xptr[14]), .Z(wptrN[14]));
Q_MX02 U963 ( .S(moveForward), .A0(wptr[15]), .A1(xptr[15]), .Z(wptrN[15]));
Q_MX02 U964 ( .S(moveForward), .A0(wptr[16]), .A1(xptr[16]), .Z(wptrN[16]));
Q_MX02 U965 ( .S(rptr[1]), .A0(n6738), .A1(n6866), .Z(iData[511]));
Q_MX02 U966 ( .S(rptr[1]), .A0(n6737), .A1(n6865), .Z(iData[510]));
Q_MX02 U967 ( .S(rptr[1]), .A0(n6736), .A1(n6864), .Z(iData[509]));
Q_MX02 U968 ( .S(rptr[1]), .A0(n6735), .A1(n6863), .Z(iData[508]));
Q_MX02 U969 ( .S(rptr[1]), .A0(n6734), .A1(n6862), .Z(iData[507]));
Q_MX02 U970 ( .S(rptr[1]), .A0(n6733), .A1(n6861), .Z(iData[506]));
Q_MX02 U971 ( .S(rptr[1]), .A0(n6732), .A1(n6860), .Z(iData[505]));
Q_MX02 U972 ( .S(rptr[1]), .A0(n6731), .A1(n6859), .Z(iData[504]));
Q_MX02 U973 ( .S(rptr[1]), .A0(n6730), .A1(n6858), .Z(iData[503]));
Q_MX02 U974 ( .S(rptr[1]), .A0(n6729), .A1(n6857), .Z(iData[502]));
Q_MX02 U975 ( .S(rptr[1]), .A0(n6728), .A1(n6856), .Z(iData[501]));
Q_MX02 U976 ( .S(rptr[1]), .A0(n6727), .A1(n6855), .Z(iData[500]));
Q_MX02 U977 ( .S(rptr[1]), .A0(n6726), .A1(n6854), .Z(iData[499]));
Q_MX02 U978 ( .S(rptr[1]), .A0(n6725), .A1(n6853), .Z(iData[498]));
Q_MX02 U979 ( .S(rptr[1]), .A0(n6724), .A1(n6852), .Z(iData[497]));
Q_MX02 U980 ( .S(rptr[1]), .A0(n6723), .A1(n6851), .Z(iData[496]));
Q_MX02 U981 ( .S(rptr[1]), .A0(n6722), .A1(n6850), .Z(iData[495]));
Q_MX02 U982 ( .S(rptr[1]), .A0(n6721), .A1(n6849), .Z(iData[494]));
Q_MX02 U983 ( .S(rptr[1]), .A0(n6720), .A1(n6848), .Z(iData[493]));
Q_MX02 U984 ( .S(rptr[1]), .A0(n6719), .A1(n6847), .Z(iData[492]));
Q_MX02 U985 ( .S(rptr[1]), .A0(n6718), .A1(n6846), .Z(iData[491]));
Q_MX02 U986 ( .S(rptr[1]), .A0(n6717), .A1(n6845), .Z(iData[490]));
Q_MX02 U987 ( .S(rptr[1]), .A0(n6716), .A1(n6844), .Z(iData[489]));
Q_MX02 U988 ( .S(rptr[1]), .A0(n6715), .A1(n6843), .Z(iData[488]));
Q_MX02 U989 ( .S(rptr[1]), .A0(n6714), .A1(n6842), .Z(iData[487]));
Q_MX02 U990 ( .S(rptr[1]), .A0(n6713), .A1(n6841), .Z(iData[486]));
Q_MX02 U991 ( .S(rptr[1]), .A0(n6712), .A1(n6840), .Z(iData[485]));
Q_MX02 U992 ( .S(rptr[1]), .A0(n6711), .A1(n6839), .Z(iData[484]));
Q_MX02 U993 ( .S(rptr[1]), .A0(n6710), .A1(n6838), .Z(iData[483]));
Q_MX02 U994 ( .S(rptr[1]), .A0(n6709), .A1(n6837), .Z(iData[482]));
Q_MX02 U995 ( .S(rptr[1]), .A0(n6708), .A1(n6836), .Z(iData[481]));
Q_MX02 U996 ( .S(rptr[1]), .A0(n6707), .A1(n6835), .Z(iData[480]));
Q_MX02 U997 ( .S(rptr[1]), .A0(n6706), .A1(n6834), .Z(iData[479]));
Q_MX02 U998 ( .S(rptr[1]), .A0(n6705), .A1(n6833), .Z(iData[478]));
Q_MX02 U999 ( .S(rptr[1]), .A0(n6704), .A1(n6832), .Z(iData[477]));
Q_MX02 U1000 ( .S(rptr[1]), .A0(n6703), .A1(n6831), .Z(iData[476]));
Q_MX02 U1001 ( .S(rptr[1]), .A0(n6702), .A1(n6830), .Z(iData[475]));
Q_MX02 U1002 ( .S(rptr[1]), .A0(n6701), .A1(n6829), .Z(iData[474]));
Q_MX02 U1003 ( .S(rptr[1]), .A0(n6700), .A1(n6828), .Z(iData[473]));
Q_MX02 U1004 ( .S(rptr[1]), .A0(n6699), .A1(n6827), .Z(iData[472]));
Q_MX02 U1005 ( .S(rptr[1]), .A0(n6698), .A1(n6826), .Z(iData[471]));
Q_MX02 U1006 ( .S(rptr[1]), .A0(n6697), .A1(n6825), .Z(iData[470]));
Q_MX02 U1007 ( .S(rptr[1]), .A0(n6696), .A1(n6824), .Z(iData[469]));
Q_MX02 U1008 ( .S(rptr[1]), .A0(n6695), .A1(n6823), .Z(iData[468]));
Q_MX02 U1009 ( .S(rptr[1]), .A0(n6694), .A1(n6822), .Z(iData[467]));
Q_MX02 U1010 ( .S(rptr[1]), .A0(n6693), .A1(n6821), .Z(iData[466]));
Q_MX02 U1011 ( .S(rptr[1]), .A0(n6692), .A1(n6820), .Z(iData[465]));
Q_MX02 U1012 ( .S(rptr[1]), .A0(n6691), .A1(n6819), .Z(iData[464]));
Q_MX02 U1013 ( .S(rptr[1]), .A0(n6690), .A1(n6818), .Z(iData[463]));
Q_MX02 U1014 ( .S(rptr[1]), .A0(n6689), .A1(n6817), .Z(iData[462]));
Q_MX02 U1015 ( .S(rptr[1]), .A0(n6688), .A1(n6816), .Z(iData[461]));
Q_MX02 U1016 ( .S(rptr[1]), .A0(n6687), .A1(n6815), .Z(iData[460]));
Q_MX02 U1017 ( .S(rptr[1]), .A0(n6686), .A1(n6814), .Z(iData[459]));
Q_MX02 U1018 ( .S(rptr[1]), .A0(n6685), .A1(n6813), .Z(iData[458]));
Q_MX02 U1019 ( .S(rptr[1]), .A0(n6684), .A1(n6812), .Z(iData[457]));
Q_MX02 U1020 ( .S(rptr[1]), .A0(n6683), .A1(n6811), .Z(iData[456]));
Q_MX02 U1021 ( .S(rptr[1]), .A0(n6682), .A1(n6810), .Z(iData[455]));
Q_MX02 U1022 ( .S(rptr[1]), .A0(n6681), .A1(n6809), .Z(iData[454]));
Q_MX02 U1023 ( .S(rptr[1]), .A0(n6680), .A1(n6808), .Z(iData[453]));
Q_MX02 U1024 ( .S(rptr[1]), .A0(n6679), .A1(n6807), .Z(iData[452]));
Q_MX02 U1025 ( .S(rptr[1]), .A0(n6678), .A1(n6806), .Z(iData[451]));
Q_MX02 U1026 ( .S(rptr[1]), .A0(n6677), .A1(n6805), .Z(iData[450]));
Q_MX02 U1027 ( .S(rptr[1]), .A0(n6676), .A1(n6804), .Z(iData[449]));
Q_MX02 U1028 ( .S(rptr[1]), .A0(n6675), .A1(n6803), .Z(iData[448]));
Q_MX02 U1029 ( .S(rptr[1]), .A0(n6674), .A1(n6802), .Z(iData[447]));
Q_MX02 U1030 ( .S(rptr[1]), .A0(n6673), .A1(n6801), .Z(iData[446]));
Q_MX02 U1031 ( .S(rptr[1]), .A0(n6672), .A1(n6800), .Z(iData[445]));
Q_MX02 U1032 ( .S(rptr[1]), .A0(n6671), .A1(n6799), .Z(iData[444]));
Q_MX02 U1033 ( .S(rptr[1]), .A0(n6670), .A1(n6798), .Z(iData[443]));
Q_MX02 U1034 ( .S(rptr[1]), .A0(n6669), .A1(n6797), .Z(iData[442]));
Q_MX02 U1035 ( .S(rptr[1]), .A0(n6668), .A1(n6796), .Z(iData[441]));
Q_MX02 U1036 ( .S(rptr[1]), .A0(n6667), .A1(n6795), .Z(iData[440]));
Q_MX02 U1037 ( .S(rptr[1]), .A0(n6666), .A1(n6794), .Z(iData[439]));
Q_MX02 U1038 ( .S(rptr[1]), .A0(n6665), .A1(n6793), .Z(iData[438]));
Q_MX02 U1039 ( .S(rptr[1]), .A0(n6664), .A1(n6792), .Z(iData[437]));
Q_MX02 U1040 ( .S(rptr[1]), .A0(n6663), .A1(n6791), .Z(iData[436]));
Q_MX02 U1041 ( .S(rptr[1]), .A0(n6662), .A1(n6790), .Z(iData[435]));
Q_MX02 U1042 ( .S(rptr[1]), .A0(n6661), .A1(n6789), .Z(iData[434]));
Q_MX02 U1043 ( .S(rptr[1]), .A0(n6660), .A1(n6788), .Z(iData[433]));
Q_MX02 U1044 ( .S(rptr[1]), .A0(n6659), .A1(n6787), .Z(iData[432]));
Q_MX02 U1045 ( .S(rptr[1]), .A0(n6658), .A1(n6786), .Z(iData[431]));
Q_MX02 U1046 ( .S(rptr[1]), .A0(n6657), .A1(n6785), .Z(iData[430]));
Q_MX02 U1047 ( .S(rptr[1]), .A0(n6656), .A1(n6784), .Z(iData[429]));
Q_MX02 U1048 ( .S(rptr[1]), .A0(n6655), .A1(n6783), .Z(iData[428]));
Q_MX02 U1049 ( .S(rptr[1]), .A0(n6654), .A1(n6782), .Z(iData[427]));
Q_MX02 U1050 ( .S(rptr[1]), .A0(n6653), .A1(n6781), .Z(iData[426]));
Q_MX02 U1051 ( .S(rptr[1]), .A0(n6652), .A1(n6780), .Z(iData[425]));
Q_MX02 U1052 ( .S(rptr[1]), .A0(n6651), .A1(n6779), .Z(iData[424]));
Q_MX02 U1053 ( .S(rptr[1]), .A0(n6650), .A1(n6778), .Z(iData[423]));
Q_MX02 U1054 ( .S(rptr[1]), .A0(n6649), .A1(n6777), .Z(iData[422]));
Q_MX02 U1055 ( .S(rptr[1]), .A0(n6648), .A1(n6776), .Z(iData[421]));
Q_MX02 U1056 ( .S(rptr[1]), .A0(n6647), .A1(n6775), .Z(iData[420]));
Q_MX02 U1057 ( .S(rptr[1]), .A0(n6646), .A1(n6774), .Z(iData[419]));
Q_MX02 U1058 ( .S(rptr[1]), .A0(n6645), .A1(n6773), .Z(iData[418]));
Q_MX02 U1059 ( .S(rptr[1]), .A0(n6644), .A1(n6772), .Z(iData[417]));
Q_MX02 U1060 ( .S(rptr[1]), .A0(n6643), .A1(n6771), .Z(iData[416]));
Q_MX02 U1061 ( .S(rptr[1]), .A0(n6642), .A1(n6770), .Z(iData[415]));
Q_MX02 U1062 ( .S(rptr[1]), .A0(n6641), .A1(n6769), .Z(iData[414]));
Q_MX02 U1063 ( .S(rptr[1]), .A0(n6640), .A1(n6768), .Z(iData[413]));
Q_MX02 U1064 ( .S(rptr[1]), .A0(n6639), .A1(n6767), .Z(iData[412]));
Q_MX02 U1065 ( .S(rptr[1]), .A0(n6638), .A1(n6766), .Z(iData[411]));
Q_MX02 U1066 ( .S(rptr[1]), .A0(n6637), .A1(n6765), .Z(iData[410]));
Q_MX02 U1067 ( .S(rptr[1]), .A0(n6636), .A1(n6764), .Z(iData[409]));
Q_MX02 U1068 ( .S(rptr[1]), .A0(n6635), .A1(n6763), .Z(iData[408]));
Q_MX02 U1069 ( .S(rptr[1]), .A0(n6634), .A1(n6762), .Z(iData[407]));
Q_MX02 U1070 ( .S(rptr[1]), .A0(n6633), .A1(n6761), .Z(iData[406]));
Q_MX02 U1071 ( .S(rptr[1]), .A0(n6632), .A1(n6760), .Z(iData[405]));
Q_MX02 U1072 ( .S(rptr[1]), .A0(n6631), .A1(n6759), .Z(iData[404]));
Q_MX02 U1073 ( .S(rptr[1]), .A0(n6630), .A1(n6758), .Z(iData[403]));
Q_MX02 U1074 ( .S(rptr[1]), .A0(n6629), .A1(n6757), .Z(iData[402]));
Q_MX02 U1075 ( .S(rptr[1]), .A0(n6628), .A1(n6756), .Z(iData[401]));
Q_MX02 U1076 ( .S(rptr[1]), .A0(n6627), .A1(n6755), .Z(iData[400]));
Q_MX02 U1077 ( .S(rptr[1]), .A0(n6626), .A1(n6754), .Z(iData[399]));
Q_MX02 U1078 ( .S(rptr[1]), .A0(n6625), .A1(n6753), .Z(iData[398]));
Q_MX02 U1079 ( .S(rptr[1]), .A0(n6624), .A1(n6752), .Z(iData[397]));
Q_MX02 U1080 ( .S(rptr[1]), .A0(n6623), .A1(n6751), .Z(iData[396]));
Q_MX02 U1081 ( .S(rptr[1]), .A0(n6622), .A1(n6750), .Z(iData[395]));
Q_MX02 U1082 ( .S(rptr[1]), .A0(n6621), .A1(n6749), .Z(iData[394]));
Q_MX02 U1083 ( .S(rptr[1]), .A0(n6620), .A1(n6748), .Z(iData[393]));
Q_MX02 U1084 ( .S(rptr[1]), .A0(n6619), .A1(n6747), .Z(iData[392]));
Q_MX02 U1085 ( .S(rptr[1]), .A0(n6618), .A1(n6746), .Z(iData[391]));
Q_MX02 U1086 ( .S(rptr[1]), .A0(n6617), .A1(n6745), .Z(iData[390]));
Q_MX02 U1087 ( .S(rptr[1]), .A0(n6616), .A1(n6744), .Z(iData[389]));
Q_MX02 U1088 ( .S(rptr[1]), .A0(n6615), .A1(n6743), .Z(iData[388]));
Q_MX02 U1089 ( .S(rptr[1]), .A0(n6614), .A1(n6742), .Z(iData[387]));
Q_MX02 U1090 ( .S(rptr[1]), .A0(n6613), .A1(n6741), .Z(iData[386]));
Q_MX02 U1091 ( .S(rptr[1]), .A0(n6612), .A1(n6740), .Z(iData[385]));
Q_MX02 U1092 ( .S(rptr[1]), .A0(n6611), .A1(n6739), .Z(iData[384]));
Q_MX02 U1093 ( .S(rptr[1]), .A0(n6610), .A1(n6738), .Z(iData[383]));
Q_MX02 U1094 ( .S(rptr[1]), .A0(n6609), .A1(n6737), .Z(iData[382]));
Q_MX02 U1095 ( .S(rptr[1]), .A0(n6608), .A1(n6736), .Z(iData[381]));
Q_MX02 U1096 ( .S(rptr[1]), .A0(n6607), .A1(n6735), .Z(iData[380]));
Q_MX02 U1097 ( .S(rptr[1]), .A0(n6606), .A1(n6734), .Z(iData[379]));
Q_MX02 U1098 ( .S(rptr[1]), .A0(n6605), .A1(n6733), .Z(iData[378]));
Q_MX02 U1099 ( .S(rptr[1]), .A0(n6604), .A1(n6732), .Z(iData[377]));
Q_MX02 U1100 ( .S(rptr[1]), .A0(n6603), .A1(n6731), .Z(iData[376]));
Q_MX02 U1101 ( .S(rptr[1]), .A0(n6602), .A1(n6730), .Z(iData[375]));
Q_MX02 U1102 ( .S(rptr[1]), .A0(n6601), .A1(n6729), .Z(iData[374]));
Q_MX02 U1103 ( .S(rptr[1]), .A0(n6600), .A1(n6728), .Z(iData[373]));
Q_MX02 U1104 ( .S(rptr[1]), .A0(n6599), .A1(n6727), .Z(iData[372]));
Q_MX02 U1105 ( .S(rptr[1]), .A0(n6598), .A1(n6726), .Z(iData[371]));
Q_MX02 U1106 ( .S(rptr[1]), .A0(n6597), .A1(n6725), .Z(iData[370]));
Q_MX02 U1107 ( .S(rptr[1]), .A0(n6596), .A1(n6724), .Z(iData[369]));
Q_MX02 U1108 ( .S(rptr[1]), .A0(n6595), .A1(n6723), .Z(iData[368]));
Q_MX02 U1109 ( .S(rptr[1]), .A0(n6594), .A1(n6722), .Z(iData[367]));
Q_MX02 U1110 ( .S(rptr[1]), .A0(n6593), .A1(n6721), .Z(iData[366]));
Q_MX02 U1111 ( .S(rptr[1]), .A0(n6592), .A1(n6720), .Z(iData[365]));
Q_MX02 U1112 ( .S(rptr[1]), .A0(n6591), .A1(n6719), .Z(iData[364]));
Q_MX02 U1113 ( .S(rptr[1]), .A0(n6590), .A1(n6718), .Z(iData[363]));
Q_MX02 U1114 ( .S(rptr[1]), .A0(n6589), .A1(n6717), .Z(iData[362]));
Q_MX02 U1115 ( .S(rptr[1]), .A0(n6588), .A1(n6716), .Z(iData[361]));
Q_MX02 U1116 ( .S(rptr[1]), .A0(n6587), .A1(n6715), .Z(iData[360]));
Q_MX02 U1117 ( .S(rptr[1]), .A0(n6586), .A1(n6714), .Z(iData[359]));
Q_MX02 U1118 ( .S(rptr[1]), .A0(n6585), .A1(n6713), .Z(iData[358]));
Q_MX02 U1119 ( .S(rptr[1]), .A0(n6584), .A1(n6712), .Z(iData[357]));
Q_MX02 U1120 ( .S(rptr[1]), .A0(n6583), .A1(n6711), .Z(iData[356]));
Q_MX02 U1121 ( .S(rptr[1]), .A0(n6582), .A1(n6710), .Z(iData[355]));
Q_MX02 U1122 ( .S(rptr[1]), .A0(n6581), .A1(n6709), .Z(iData[354]));
Q_MX02 U1123 ( .S(rptr[1]), .A0(n6580), .A1(n6708), .Z(iData[353]));
Q_MX02 U1124 ( .S(rptr[1]), .A0(n6579), .A1(n6707), .Z(iData[352]));
Q_MX02 U1125 ( .S(rptr[1]), .A0(n6578), .A1(n6706), .Z(iData[351]));
Q_MX02 U1126 ( .S(rptr[1]), .A0(n6577), .A1(n6705), .Z(iData[350]));
Q_MX02 U1127 ( .S(rptr[1]), .A0(n6576), .A1(n6704), .Z(iData[349]));
Q_MX02 U1128 ( .S(rptr[1]), .A0(n6575), .A1(n6703), .Z(iData[348]));
Q_MX02 U1129 ( .S(rptr[1]), .A0(n6574), .A1(n6702), .Z(iData[347]));
Q_MX02 U1130 ( .S(rptr[1]), .A0(n6573), .A1(n6701), .Z(iData[346]));
Q_MX02 U1131 ( .S(rptr[1]), .A0(n6572), .A1(n6700), .Z(iData[345]));
Q_MX02 U1132 ( .S(rptr[1]), .A0(n6571), .A1(n6699), .Z(iData[344]));
Q_MX02 U1133 ( .S(rptr[1]), .A0(n6570), .A1(n6698), .Z(iData[343]));
Q_MX02 U1134 ( .S(rptr[1]), .A0(n6569), .A1(n6697), .Z(iData[342]));
Q_MX02 U1135 ( .S(rptr[1]), .A0(n6568), .A1(n6696), .Z(iData[341]));
Q_MX02 U1136 ( .S(rptr[1]), .A0(n6567), .A1(n6695), .Z(iData[340]));
Q_MX02 U1137 ( .S(rptr[1]), .A0(n6566), .A1(n6694), .Z(iData[339]));
Q_MX02 U1138 ( .S(rptr[1]), .A0(n6565), .A1(n6693), .Z(iData[338]));
Q_MX02 U1139 ( .S(rptr[1]), .A0(n6564), .A1(n6692), .Z(iData[337]));
Q_MX02 U1140 ( .S(rptr[1]), .A0(n6563), .A1(n6691), .Z(iData[336]));
Q_MX02 U1141 ( .S(rptr[1]), .A0(n6562), .A1(n6690), .Z(iData[335]));
Q_MX02 U1142 ( .S(rptr[1]), .A0(n6561), .A1(n6689), .Z(iData[334]));
Q_MX02 U1143 ( .S(rptr[1]), .A0(n6560), .A1(n6688), .Z(iData[333]));
Q_MX02 U1144 ( .S(rptr[1]), .A0(n6559), .A1(n6687), .Z(iData[332]));
Q_MX02 U1145 ( .S(rptr[1]), .A0(n6558), .A1(n6686), .Z(iData[331]));
Q_MX02 U1146 ( .S(rptr[1]), .A0(n6557), .A1(n6685), .Z(iData[330]));
Q_MX02 U1147 ( .S(rptr[1]), .A0(n6556), .A1(n6684), .Z(iData[329]));
Q_MX02 U1148 ( .S(rptr[1]), .A0(n6555), .A1(n6683), .Z(iData[328]));
Q_MX02 U1149 ( .S(rptr[1]), .A0(n6554), .A1(n6682), .Z(iData[327]));
Q_MX02 U1150 ( .S(rptr[1]), .A0(n6553), .A1(n6681), .Z(iData[326]));
Q_MX02 U1151 ( .S(rptr[1]), .A0(n6552), .A1(n6680), .Z(iData[325]));
Q_MX02 U1152 ( .S(rptr[1]), .A0(n6551), .A1(n6679), .Z(iData[324]));
Q_MX02 U1153 ( .S(rptr[1]), .A0(n6550), .A1(n6678), .Z(iData[323]));
Q_MX02 U1154 ( .S(rptr[1]), .A0(n6549), .A1(n6677), .Z(iData[322]));
Q_MX02 U1155 ( .S(rptr[1]), .A0(n6548), .A1(n6676), .Z(iData[321]));
Q_MX02 U1156 ( .S(rptr[1]), .A0(n6547), .A1(n6675), .Z(iData[320]));
Q_MX02 U1157 ( .S(rptr[1]), .A0(n6546), .A1(n6674), .Z(iData[319]));
Q_MX02 U1158 ( .S(rptr[1]), .A0(n6545), .A1(n6673), .Z(iData[318]));
Q_MX02 U1159 ( .S(rptr[1]), .A0(n6544), .A1(n6672), .Z(iData[317]));
Q_MX02 U1160 ( .S(rptr[1]), .A0(n6543), .A1(n6671), .Z(iData[316]));
Q_MX02 U1161 ( .S(rptr[1]), .A0(n6542), .A1(n6670), .Z(iData[315]));
Q_MX02 U1162 ( .S(rptr[1]), .A0(n6541), .A1(n6669), .Z(iData[314]));
Q_MX02 U1163 ( .S(rptr[1]), .A0(n6540), .A1(n6668), .Z(iData[313]));
Q_MX02 U1164 ( .S(rptr[1]), .A0(n6539), .A1(n6667), .Z(iData[312]));
Q_MX02 U1165 ( .S(rptr[1]), .A0(n6538), .A1(n6666), .Z(iData[311]));
Q_MX02 U1166 ( .S(rptr[1]), .A0(n6537), .A1(n6665), .Z(iData[310]));
Q_MX02 U1167 ( .S(rptr[1]), .A0(n6536), .A1(n6664), .Z(iData[309]));
Q_MX02 U1168 ( .S(rptr[1]), .A0(n6535), .A1(n6663), .Z(iData[308]));
Q_MX02 U1169 ( .S(rptr[1]), .A0(n6534), .A1(n6662), .Z(iData[307]));
Q_MX02 U1170 ( .S(rptr[1]), .A0(n6533), .A1(n6661), .Z(iData[306]));
Q_MX02 U1171 ( .S(rptr[1]), .A0(n6532), .A1(n6660), .Z(iData[305]));
Q_MX02 U1172 ( .S(rptr[1]), .A0(n6531), .A1(n6659), .Z(iData[304]));
Q_MX02 U1173 ( .S(rptr[1]), .A0(n6530), .A1(n6658), .Z(iData[303]));
Q_MX02 U1174 ( .S(rptr[1]), .A0(n6529), .A1(n6657), .Z(iData[302]));
Q_MX02 U1175 ( .S(rptr[1]), .A0(n6528), .A1(n6656), .Z(iData[301]));
Q_MX02 U1176 ( .S(rptr[1]), .A0(n6527), .A1(n6655), .Z(iData[300]));
Q_MX02 U1177 ( .S(rptr[1]), .A0(n6526), .A1(n6654), .Z(iData[299]));
Q_MX02 U1178 ( .S(rptr[1]), .A0(n6525), .A1(n6653), .Z(iData[298]));
Q_MX02 U1179 ( .S(rptr[1]), .A0(n6524), .A1(n6652), .Z(iData[297]));
Q_MX02 U1180 ( .S(rptr[1]), .A0(n6523), .A1(n6651), .Z(iData[296]));
Q_MX02 U1181 ( .S(rptr[1]), .A0(n6522), .A1(n6650), .Z(iData[295]));
Q_MX02 U1182 ( .S(rptr[1]), .A0(n6521), .A1(n6649), .Z(iData[294]));
Q_MX02 U1183 ( .S(rptr[1]), .A0(n6520), .A1(n6648), .Z(iData[293]));
Q_MX02 U1184 ( .S(rptr[1]), .A0(n6519), .A1(n6647), .Z(iData[292]));
Q_MX02 U1185 ( .S(rptr[1]), .A0(n6518), .A1(n6646), .Z(iData[291]));
Q_MX02 U1186 ( .S(rptr[1]), .A0(n6517), .A1(n6645), .Z(iData[290]));
Q_MX02 U1187 ( .S(rptr[1]), .A0(n6516), .A1(n6644), .Z(iData[289]));
Q_MX02 U1188 ( .S(rptr[1]), .A0(n6515), .A1(n6643), .Z(iData[288]));
Q_MX02 U1189 ( .S(rptr[1]), .A0(n6514), .A1(n6642), .Z(iData[287]));
Q_MX02 U1190 ( .S(rptr[1]), .A0(n6513), .A1(n6641), .Z(iData[286]));
Q_MX02 U1191 ( .S(rptr[1]), .A0(n6512), .A1(n6640), .Z(iData[285]));
Q_MX02 U1192 ( .S(rptr[1]), .A0(n6511), .A1(n6639), .Z(iData[284]));
Q_MX02 U1193 ( .S(rptr[1]), .A0(n6510), .A1(n6638), .Z(iData[283]));
Q_MX02 U1194 ( .S(rptr[1]), .A0(n6509), .A1(n6637), .Z(iData[282]));
Q_MX02 U1195 ( .S(rptr[1]), .A0(n6508), .A1(n6636), .Z(iData[281]));
Q_MX02 U1196 ( .S(rptr[1]), .A0(n6507), .A1(n6635), .Z(iData[280]));
Q_MX02 U1197 ( .S(rptr[1]), .A0(n6506), .A1(n6634), .Z(iData[279]));
Q_MX02 U1198 ( .S(rptr[1]), .A0(n6505), .A1(n6633), .Z(iData[278]));
Q_MX02 U1199 ( .S(rptr[1]), .A0(n6504), .A1(n6632), .Z(iData[277]));
Q_MX02 U1200 ( .S(rptr[1]), .A0(n6503), .A1(n6631), .Z(iData[276]));
Q_MX02 U1201 ( .S(rptr[1]), .A0(n6502), .A1(n6630), .Z(iData[275]));
Q_MX02 U1202 ( .S(rptr[1]), .A0(n6501), .A1(n6629), .Z(iData[274]));
Q_MX02 U1203 ( .S(rptr[1]), .A0(n6500), .A1(n6628), .Z(iData[273]));
Q_MX02 U1204 ( .S(rptr[1]), .A0(n6499), .A1(n6627), .Z(iData[272]));
Q_MX02 U1205 ( .S(rptr[1]), .A0(n6498), .A1(n6626), .Z(iData[271]));
Q_MX02 U1206 ( .S(rptr[1]), .A0(n6497), .A1(n6625), .Z(iData[270]));
Q_MX02 U1207 ( .S(rptr[1]), .A0(n6496), .A1(n6624), .Z(iData[269]));
Q_MX02 U1208 ( .S(rptr[1]), .A0(n6495), .A1(n6623), .Z(iData[268]));
Q_MX02 U1209 ( .S(rptr[1]), .A0(n6494), .A1(n6622), .Z(iData[267]));
Q_MX02 U1210 ( .S(rptr[1]), .A0(n6493), .A1(n6621), .Z(iData[266]));
Q_MX02 U1211 ( .S(rptr[1]), .A0(n6492), .A1(n6620), .Z(iData[265]));
Q_MX02 U1212 ( .S(rptr[1]), .A0(n6491), .A1(n6619), .Z(iData[264]));
Q_MX02 U1213 ( .S(rptr[1]), .A0(n6490), .A1(n6618), .Z(iData[263]));
Q_MX02 U1214 ( .S(rptr[1]), .A0(n6489), .A1(n6617), .Z(iData[262]));
Q_MX02 U1215 ( .S(rptr[1]), .A0(n6488), .A1(n6616), .Z(iData[261]));
Q_MX02 U1216 ( .S(rptr[1]), .A0(n6487), .A1(n6615), .Z(iData[260]));
Q_MX02 U1217 ( .S(rptr[1]), .A0(n6486), .A1(n6614), .Z(iData[259]));
Q_MX02 U1218 ( .S(rptr[1]), .A0(n6485), .A1(n6613), .Z(iData[258]));
Q_MX02 U1219 ( .S(rptr[1]), .A0(n6484), .A1(n6612), .Z(iData[257]));
Q_MX02 U1220 ( .S(rptr[1]), .A0(n6483), .A1(n6611), .Z(iData[256]));
Q_MX02 U1221 ( .S(rptr[1]), .A0(n6482), .A1(n6610), .Z(iData[255]));
Q_MX02 U1222 ( .S(rptr[1]), .A0(n6481), .A1(n6609), .Z(iData[254]));
Q_MX02 U1223 ( .S(rptr[1]), .A0(n6480), .A1(n6608), .Z(iData[253]));
Q_MX02 U1224 ( .S(rptr[1]), .A0(n6479), .A1(n6607), .Z(iData[252]));
Q_MX02 U1225 ( .S(rptr[1]), .A0(n6478), .A1(n6606), .Z(iData[251]));
Q_MX02 U1226 ( .S(rptr[1]), .A0(n6477), .A1(n6605), .Z(iData[250]));
Q_MX02 U1227 ( .S(rptr[1]), .A0(n6476), .A1(n6604), .Z(iData[249]));
Q_MX02 U1228 ( .S(rptr[1]), .A0(n6475), .A1(n6603), .Z(iData[248]));
Q_MX02 U1229 ( .S(rptr[1]), .A0(n6474), .A1(n6602), .Z(iData[247]));
Q_MX02 U1230 ( .S(rptr[1]), .A0(n6473), .A1(n6601), .Z(iData[246]));
Q_MX02 U1231 ( .S(rptr[1]), .A0(n6472), .A1(n6600), .Z(iData[245]));
Q_MX02 U1232 ( .S(rptr[1]), .A0(n6471), .A1(n6599), .Z(iData[244]));
Q_MX02 U1233 ( .S(rptr[1]), .A0(n6470), .A1(n6598), .Z(iData[243]));
Q_MX02 U1234 ( .S(rptr[1]), .A0(n6469), .A1(n6597), .Z(iData[242]));
Q_MX02 U1235 ( .S(rptr[1]), .A0(n6468), .A1(n6596), .Z(iData[241]));
Q_MX02 U1236 ( .S(rptr[1]), .A0(n6467), .A1(n6595), .Z(iData[240]));
Q_MX02 U1237 ( .S(rptr[1]), .A0(n6466), .A1(n6594), .Z(iData[239]));
Q_MX02 U1238 ( .S(rptr[1]), .A0(n6465), .A1(n6593), .Z(iData[238]));
Q_MX02 U1239 ( .S(rptr[1]), .A0(n6464), .A1(n6592), .Z(iData[237]));
Q_MX02 U1240 ( .S(rptr[1]), .A0(n6463), .A1(n6591), .Z(iData[236]));
Q_MX02 U1241 ( .S(rptr[1]), .A0(n6462), .A1(n6590), .Z(iData[235]));
Q_MX02 U1242 ( .S(rptr[1]), .A0(n6461), .A1(n6589), .Z(iData[234]));
Q_MX02 U1243 ( .S(rptr[1]), .A0(n6460), .A1(n6588), .Z(iData[233]));
Q_MX02 U1244 ( .S(rptr[1]), .A0(n6459), .A1(n6587), .Z(iData[232]));
Q_MX02 U1245 ( .S(rptr[1]), .A0(n6458), .A1(n6586), .Z(iData[231]));
Q_MX02 U1246 ( .S(rptr[1]), .A0(n6457), .A1(n6585), .Z(iData[230]));
Q_MX02 U1247 ( .S(rptr[1]), .A0(n6456), .A1(n6584), .Z(iData[229]));
Q_MX02 U1248 ( .S(rptr[1]), .A0(n6455), .A1(n6583), .Z(iData[228]));
Q_MX02 U1249 ( .S(rptr[1]), .A0(n6454), .A1(n6582), .Z(iData[227]));
Q_MX02 U1250 ( .S(rptr[1]), .A0(n6453), .A1(n6581), .Z(iData[226]));
Q_MX02 U1251 ( .S(rptr[1]), .A0(n6452), .A1(n6580), .Z(iData[225]));
Q_MX02 U1252 ( .S(rptr[1]), .A0(n6451), .A1(n6579), .Z(iData[224]));
Q_MX02 U1253 ( .S(rptr[1]), .A0(n6450), .A1(n6578), .Z(iData[223]));
Q_MX02 U1254 ( .S(rptr[1]), .A0(n6449), .A1(n6577), .Z(iData[222]));
Q_MX02 U1255 ( .S(rptr[1]), .A0(n6448), .A1(n6576), .Z(iData[221]));
Q_MX02 U1256 ( .S(rptr[1]), .A0(n6447), .A1(n6575), .Z(iData[220]));
Q_MX02 U1257 ( .S(rptr[1]), .A0(n6446), .A1(n6574), .Z(iData[219]));
Q_MX02 U1258 ( .S(rptr[1]), .A0(n6445), .A1(n6573), .Z(iData[218]));
Q_MX02 U1259 ( .S(rptr[1]), .A0(n6444), .A1(n6572), .Z(iData[217]));
Q_MX02 U1260 ( .S(rptr[1]), .A0(n6443), .A1(n6571), .Z(iData[216]));
Q_MX02 U1261 ( .S(rptr[1]), .A0(n6442), .A1(n6570), .Z(iData[215]));
Q_MX02 U1262 ( .S(rptr[1]), .A0(n6441), .A1(n6569), .Z(iData[214]));
Q_MX02 U1263 ( .S(rptr[1]), .A0(n6440), .A1(n6568), .Z(iData[213]));
Q_MX02 U1264 ( .S(rptr[1]), .A0(n6439), .A1(n6567), .Z(iData[212]));
Q_MX02 U1265 ( .S(rptr[1]), .A0(n6438), .A1(n6566), .Z(iData[211]));
Q_MX02 U1266 ( .S(rptr[1]), .A0(n6437), .A1(n6565), .Z(iData[210]));
Q_MX02 U1267 ( .S(rptr[1]), .A0(n6436), .A1(n6564), .Z(iData[209]));
Q_MX02 U1268 ( .S(rptr[1]), .A0(n6435), .A1(n6563), .Z(iData[208]));
Q_MX02 U1269 ( .S(rptr[1]), .A0(n6434), .A1(n6562), .Z(iData[207]));
Q_MX02 U1270 ( .S(rptr[1]), .A0(n6433), .A1(n6561), .Z(iData[206]));
Q_MX02 U1271 ( .S(rptr[1]), .A0(n6432), .A1(n6560), .Z(iData[205]));
Q_MX02 U1272 ( .S(rptr[1]), .A0(n6431), .A1(n6559), .Z(iData[204]));
Q_MX02 U1273 ( .S(rptr[1]), .A0(n6430), .A1(n6558), .Z(iData[203]));
Q_MX02 U1274 ( .S(rptr[1]), .A0(n6429), .A1(n6557), .Z(iData[202]));
Q_MX02 U1275 ( .S(rptr[1]), .A0(n6428), .A1(n6556), .Z(iData[201]));
Q_MX02 U1276 ( .S(rptr[1]), .A0(n6427), .A1(n6555), .Z(iData[200]));
Q_MX02 U1277 ( .S(rptr[1]), .A0(n6426), .A1(n6554), .Z(iData[199]));
Q_MX02 U1278 ( .S(rptr[1]), .A0(n6425), .A1(n6553), .Z(iData[198]));
Q_MX02 U1279 ( .S(rptr[1]), .A0(n6424), .A1(n6552), .Z(iData[197]));
Q_MX02 U1280 ( .S(rptr[1]), .A0(n6423), .A1(n6551), .Z(iData[196]));
Q_MX02 U1281 ( .S(rptr[1]), .A0(n6422), .A1(n6550), .Z(iData[195]));
Q_MX02 U1282 ( .S(rptr[1]), .A0(n6421), .A1(n6549), .Z(iData[194]));
Q_MX02 U1283 ( .S(rptr[1]), .A0(n6420), .A1(n6548), .Z(iData[193]));
Q_MX02 U1284 ( .S(rptr[1]), .A0(n6419), .A1(n6547), .Z(iData[192]));
Q_MX02 U1285 ( .S(rptr[1]), .A0(n6418), .A1(n6546), .Z(iData[191]));
Q_MX02 U1286 ( .S(rptr[1]), .A0(n6417), .A1(n6545), .Z(iData[190]));
Q_MX02 U1287 ( .S(rptr[1]), .A0(n6416), .A1(n6544), .Z(iData[189]));
Q_MX02 U1288 ( .S(rptr[1]), .A0(n6415), .A1(n6543), .Z(iData[188]));
Q_MX02 U1289 ( .S(rptr[1]), .A0(n6414), .A1(n6542), .Z(iData[187]));
Q_MX02 U1290 ( .S(rptr[1]), .A0(n6413), .A1(n6541), .Z(iData[186]));
Q_MX02 U1291 ( .S(rptr[1]), .A0(n6412), .A1(n6540), .Z(iData[185]));
Q_MX02 U1292 ( .S(rptr[1]), .A0(n6411), .A1(n6539), .Z(iData[184]));
Q_MX02 U1293 ( .S(rptr[1]), .A0(n6410), .A1(n6538), .Z(iData[183]));
Q_MX02 U1294 ( .S(rptr[1]), .A0(n6409), .A1(n6537), .Z(iData[182]));
Q_MX02 U1295 ( .S(rptr[1]), .A0(n6408), .A1(n6536), .Z(iData[181]));
Q_MX02 U1296 ( .S(rptr[1]), .A0(n6407), .A1(n6535), .Z(iData[180]));
Q_MX02 U1297 ( .S(rptr[1]), .A0(n6406), .A1(n6534), .Z(iData[179]));
Q_MX02 U1298 ( .S(rptr[1]), .A0(n6405), .A1(n6533), .Z(iData[178]));
Q_MX02 U1299 ( .S(rptr[1]), .A0(n6404), .A1(n6532), .Z(iData[177]));
Q_MX02 U1300 ( .S(rptr[1]), .A0(n6403), .A1(n6531), .Z(iData[176]));
Q_MX02 U1301 ( .S(rptr[1]), .A0(n6402), .A1(n6530), .Z(iData[175]));
Q_MX02 U1302 ( .S(rptr[1]), .A0(n6401), .A1(n6529), .Z(iData[174]));
Q_MX02 U1303 ( .S(rptr[1]), .A0(n6400), .A1(n6528), .Z(iData[173]));
Q_MX02 U1304 ( .S(rptr[1]), .A0(n6399), .A1(n6527), .Z(iData[172]));
Q_MX02 U1305 ( .S(rptr[1]), .A0(n6398), .A1(n6526), .Z(iData[171]));
Q_MX02 U1306 ( .S(rptr[1]), .A0(n6397), .A1(n6525), .Z(iData[170]));
Q_MX02 U1307 ( .S(rptr[1]), .A0(n6396), .A1(n6524), .Z(iData[169]));
Q_MX02 U1308 ( .S(rptr[1]), .A0(n6395), .A1(n6523), .Z(iData[168]));
Q_MX02 U1309 ( .S(rptr[1]), .A0(n6394), .A1(n6522), .Z(iData[167]));
Q_MX02 U1310 ( .S(rptr[1]), .A0(n6393), .A1(n6521), .Z(iData[166]));
Q_MX02 U1311 ( .S(rptr[1]), .A0(n6392), .A1(n6520), .Z(iData[165]));
Q_MX02 U1312 ( .S(rptr[1]), .A0(n6391), .A1(n6519), .Z(iData[164]));
Q_MX02 U1313 ( .S(rptr[1]), .A0(n6390), .A1(n6518), .Z(iData[163]));
Q_MX02 U1314 ( .S(rptr[1]), .A0(n6389), .A1(n6517), .Z(iData[162]));
Q_MX02 U1315 ( .S(rptr[1]), .A0(n6388), .A1(n6516), .Z(iData[161]));
Q_MX02 U1316 ( .S(rptr[1]), .A0(n6387), .A1(n6515), .Z(iData[160]));
Q_MX02 U1317 ( .S(rptr[1]), .A0(n6386), .A1(n6514), .Z(iData[159]));
Q_MX02 U1318 ( .S(rptr[1]), .A0(n6385), .A1(n6513), .Z(iData[158]));
Q_MX02 U1319 ( .S(rptr[1]), .A0(n6384), .A1(n6512), .Z(iData[157]));
Q_MX02 U1320 ( .S(rptr[1]), .A0(n6383), .A1(n6511), .Z(iData[156]));
Q_MX02 U1321 ( .S(rptr[1]), .A0(n6382), .A1(n6510), .Z(iData[155]));
Q_MX02 U1322 ( .S(rptr[1]), .A0(n6381), .A1(n6509), .Z(iData[154]));
Q_MX02 U1323 ( .S(rptr[1]), .A0(n6380), .A1(n6508), .Z(iData[153]));
Q_MX02 U1324 ( .S(rptr[1]), .A0(n6379), .A1(n6507), .Z(iData[152]));
Q_MX02 U1325 ( .S(rptr[1]), .A0(n6378), .A1(n6506), .Z(iData[151]));
Q_MX02 U1326 ( .S(rptr[1]), .A0(n6377), .A1(n6505), .Z(iData[150]));
Q_MX02 U1327 ( .S(rptr[1]), .A0(n6376), .A1(n6504), .Z(iData[149]));
Q_MX02 U1328 ( .S(rptr[1]), .A0(n6375), .A1(n6503), .Z(iData[148]));
Q_MX02 U1329 ( .S(rptr[1]), .A0(n6374), .A1(n6502), .Z(iData[147]));
Q_MX02 U1330 ( .S(rptr[1]), .A0(n6373), .A1(n6501), .Z(iData[146]));
Q_MX02 U1331 ( .S(rptr[1]), .A0(n6372), .A1(n6500), .Z(iData[145]));
Q_MX02 U1332 ( .S(rptr[1]), .A0(n6371), .A1(n6499), .Z(iData[144]));
Q_MX02 U1333 ( .S(rptr[1]), .A0(n6370), .A1(n6498), .Z(iData[143]));
Q_MX02 U1334 ( .S(rptr[1]), .A0(n6369), .A1(n6497), .Z(iData[142]));
Q_MX02 U1335 ( .S(rptr[1]), .A0(n6368), .A1(n6496), .Z(iData[141]));
Q_MX02 U1336 ( .S(rptr[1]), .A0(n6367), .A1(n6495), .Z(iData[140]));
Q_MX02 U1337 ( .S(rptr[1]), .A0(n6366), .A1(n6494), .Z(iData[139]));
Q_MX02 U1338 ( .S(rptr[1]), .A0(n6365), .A1(n6493), .Z(iData[138]));
Q_MX02 U1339 ( .S(rptr[1]), .A0(n6364), .A1(n6492), .Z(iData[137]));
Q_MX02 U1340 ( .S(rptr[1]), .A0(n6363), .A1(n6491), .Z(iData[136]));
Q_MX02 U1341 ( .S(rptr[1]), .A0(n6362), .A1(n6490), .Z(iData[135]));
Q_MX02 U1342 ( .S(rptr[1]), .A0(n6361), .A1(n6489), .Z(iData[134]));
Q_MX02 U1343 ( .S(rptr[1]), .A0(n6360), .A1(n6488), .Z(iData[133]));
Q_MX02 U1344 ( .S(rptr[1]), .A0(n6359), .A1(n6487), .Z(iData[132]));
Q_MX02 U1345 ( .S(rptr[1]), .A0(n6358), .A1(n6486), .Z(iData[131]));
Q_MX02 U1346 ( .S(rptr[1]), .A0(n6357), .A1(n6485), .Z(iData[130]));
Q_MX02 U1347 ( .S(rptr[1]), .A0(n6356), .A1(n6484), .Z(iData[129]));
Q_MX02 U1348 ( .S(rptr[1]), .A0(n6355), .A1(n6483), .Z(iData[128]));
Q_MX02 U1349 ( .S(rptr[1]), .A0(n6354), .A1(n6482), .Z(iData[127]));
Q_MX02 U1350 ( .S(rptr[1]), .A0(n6353), .A1(n6481), .Z(iData[126]));
Q_MX02 U1351 ( .S(rptr[1]), .A0(n6352), .A1(n6480), .Z(iData[125]));
Q_MX02 U1352 ( .S(rptr[1]), .A0(n6351), .A1(n6479), .Z(iData[124]));
Q_MX02 U1353 ( .S(rptr[1]), .A0(n6350), .A1(n6478), .Z(iData[123]));
Q_MX02 U1354 ( .S(rptr[1]), .A0(n6349), .A1(n6477), .Z(iData[122]));
Q_MX02 U1355 ( .S(rptr[1]), .A0(n6348), .A1(n6476), .Z(iData[121]));
Q_MX02 U1356 ( .S(rptr[1]), .A0(n6347), .A1(n6475), .Z(iData[120]));
Q_MX02 U1357 ( .S(rptr[1]), .A0(n6346), .A1(n6474), .Z(iData[119]));
Q_MX02 U1358 ( .S(rptr[1]), .A0(n6345), .A1(n6473), .Z(iData[118]));
Q_MX02 U1359 ( .S(rptr[1]), .A0(n6344), .A1(n6472), .Z(iData[117]));
Q_MX02 U1360 ( .S(rptr[1]), .A0(n6343), .A1(n6471), .Z(iData[116]));
Q_MX02 U1361 ( .S(rptr[1]), .A0(n6342), .A1(n6470), .Z(iData[115]));
Q_MX02 U1362 ( .S(rptr[1]), .A0(n6341), .A1(n6469), .Z(iData[114]));
Q_MX02 U1363 ( .S(rptr[1]), .A0(n6340), .A1(n6468), .Z(iData[113]));
Q_MX02 U1364 ( .S(rptr[1]), .A0(n6339), .A1(n6467), .Z(iData[112]));
Q_MX02 U1365 ( .S(rptr[1]), .A0(n6338), .A1(n6466), .Z(iData[111]));
Q_MX02 U1366 ( .S(rptr[1]), .A0(n6337), .A1(n6465), .Z(iData[110]));
Q_MX02 U1367 ( .S(rptr[1]), .A0(n6336), .A1(n6464), .Z(iData[109]));
Q_MX02 U1368 ( .S(rptr[1]), .A0(n6335), .A1(n6463), .Z(iData[108]));
Q_MX02 U1369 ( .S(rptr[1]), .A0(n6334), .A1(n6462), .Z(iData[107]));
Q_MX02 U1370 ( .S(rptr[1]), .A0(n6333), .A1(n6461), .Z(iData[106]));
Q_MX02 U1371 ( .S(rptr[1]), .A0(n6332), .A1(n6460), .Z(iData[105]));
Q_MX02 U1372 ( .S(rptr[1]), .A0(n6331), .A1(n6459), .Z(iData[104]));
Q_MX02 U1373 ( .S(rptr[1]), .A0(n6330), .A1(n6458), .Z(iData[103]));
Q_MX02 U1374 ( .S(rptr[1]), .A0(n6329), .A1(n6457), .Z(iData[102]));
Q_MX02 U1375 ( .S(rptr[1]), .A0(n6328), .A1(n6456), .Z(iData[101]));
Q_MX02 U1376 ( .S(rptr[1]), .A0(n6327), .A1(n6455), .Z(iData[100]));
Q_MX02 U1377 ( .S(rptr[1]), .A0(n6326), .A1(n6454), .Z(iData[99]));
Q_MX02 U1378 ( .S(rptr[1]), .A0(n6325), .A1(n6453), .Z(iData[98]));
Q_MX02 U1379 ( .S(rptr[1]), .A0(n6324), .A1(n6452), .Z(iData[97]));
Q_MX02 U1380 ( .S(rptr[1]), .A0(n6323), .A1(n6451), .Z(iData[96]));
Q_MX02 U1381 ( .S(rptr[1]), .A0(n6322), .A1(n6450), .Z(iData[95]));
Q_MX02 U1382 ( .S(rptr[1]), .A0(n6321), .A1(n6449), .Z(iData[94]));
Q_MX02 U1383 ( .S(rptr[1]), .A0(n6320), .A1(n6448), .Z(iData[93]));
Q_MX02 U1384 ( .S(rptr[1]), .A0(n6319), .A1(n6447), .Z(iData[92]));
Q_MX02 U1385 ( .S(rptr[1]), .A0(n6318), .A1(n6446), .Z(iData[91]));
Q_MX02 U1386 ( .S(rptr[1]), .A0(n6317), .A1(n6445), .Z(iData[90]));
Q_MX02 U1387 ( .S(rptr[1]), .A0(n6316), .A1(n6444), .Z(iData[89]));
Q_MX02 U1388 ( .S(rptr[1]), .A0(n6315), .A1(n6443), .Z(iData[88]));
Q_MX02 U1389 ( .S(rptr[1]), .A0(n6314), .A1(n6442), .Z(iData[87]));
Q_MX02 U1390 ( .S(rptr[1]), .A0(n6313), .A1(n6441), .Z(iData[86]));
Q_MX02 U1391 ( .S(rptr[1]), .A0(n6312), .A1(n6440), .Z(iData[85]));
Q_MX02 U1392 ( .S(rptr[1]), .A0(n6311), .A1(n6439), .Z(iData[84]));
Q_MX02 U1393 ( .S(rptr[1]), .A0(n6310), .A1(n6438), .Z(iData[83]));
Q_MX02 U1394 ( .S(rptr[1]), .A0(n6309), .A1(n6437), .Z(iData[82]));
Q_MX02 U1395 ( .S(rptr[1]), .A0(n6308), .A1(n6436), .Z(iData[81]));
Q_MX02 U1396 ( .S(rptr[1]), .A0(n6307), .A1(n6435), .Z(iData[80]));
Q_MX02 U1397 ( .S(rptr[1]), .A0(n6306), .A1(n6434), .Z(iData[79]));
Q_MX02 U1398 ( .S(rptr[1]), .A0(n6305), .A1(n6433), .Z(iData[78]));
Q_MX02 U1399 ( .S(rptr[1]), .A0(n6304), .A1(n6432), .Z(iData[77]));
Q_MX02 U1400 ( .S(rptr[1]), .A0(n6303), .A1(n6431), .Z(iData[76]));
Q_MX02 U1401 ( .S(rptr[1]), .A0(n6302), .A1(n6430), .Z(iData[75]));
Q_MX02 U1402 ( .S(rptr[1]), .A0(n6301), .A1(n6429), .Z(iData[74]));
Q_MX02 U1403 ( .S(rptr[1]), .A0(n6300), .A1(n6428), .Z(iData[73]));
Q_MX02 U1404 ( .S(rptr[1]), .A0(n6299), .A1(n6427), .Z(iData[72]));
Q_MX02 U1405 ( .S(rptr[1]), .A0(n6298), .A1(n6426), .Z(iData[71]));
Q_MX02 U1406 ( .S(rptr[1]), .A0(n6297), .A1(n6425), .Z(iData[70]));
Q_MX02 U1407 ( .S(rptr[1]), .A0(n6296), .A1(n6424), .Z(iData[69]));
Q_MX02 U1408 ( .S(rptr[1]), .A0(n6295), .A1(n6423), .Z(iData[68]));
Q_MX02 U1409 ( .S(rptr[1]), .A0(n6294), .A1(n6422), .Z(iData[67]));
Q_MX02 U1410 ( .S(rptr[1]), .A0(n6293), .A1(n6421), .Z(iData[66]));
Q_MX02 U1411 ( .S(rptr[1]), .A0(n6292), .A1(n6420), .Z(iData[65]));
Q_MX02 U1412 ( .S(rptr[1]), .A0(n6291), .A1(n6419), .Z(iData[64]));
Q_MX03 U1413 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[127]), .A1(ififoRdata[191]), .A2(n6418), .Z(iData[63]));
Q_MX03 U1414 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[126]), .A1(ififoRdata[190]), .A2(n6417), .Z(iData[62]));
Q_MX03 U1415 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[125]), .A1(ififoRdata[189]), .A2(n6416), .Z(iData[61]));
Q_MX03 U1416 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[124]), .A1(ififoRdata[188]), .A2(n6415), .Z(iData[60]));
Q_MX03 U1417 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[123]), .A1(ififoRdata[187]), .A2(n6414), .Z(iData[59]));
Q_MX03 U1418 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[122]), .A1(ififoRdata[186]), .A2(n6413), .Z(iData[58]));
Q_MX03 U1419 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[121]), .A1(ififoRdata[185]), .A2(n6412), .Z(iData[57]));
Q_MX03 U1420 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[120]), .A1(ififoRdata[184]), .A2(n6411), .Z(iData[56]));
Q_MX03 U1421 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[119]), .A1(ififoRdata[183]), .A2(n6410), .Z(iData[55]));
Q_MX03 U1422 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[118]), .A1(ififoRdata[182]), .A2(n6409), .Z(iData[54]));
Q_MX03 U1423 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[117]), .A1(ififoRdata[181]), .A2(n6408), .Z(iData[53]));
Q_MX03 U1424 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[116]), .A1(ififoRdata[180]), .A2(n6407), .Z(iData[52]));
Q_MX03 U1425 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[115]), .A1(ififoRdata[179]), .A2(n6406), .Z(iData[51]));
Q_MX03 U1426 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[114]), .A1(ififoRdata[178]), .A2(n6405), .Z(iData[50]));
Q_MX03 U1427 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[113]), .A1(ififoRdata[177]), .A2(n6404), .Z(iData[49]));
Q_MX03 U1428 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[112]), .A1(ififoRdata[176]), .A2(n6403), .Z(iData[48]));
Q_MX03 U1429 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[111]), .A1(ififoRdata[175]), .A2(n6402), .Z(iData[47]));
Q_MX03 U1430 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[110]), .A1(ififoRdata[174]), .A2(n6401), .Z(iData[46]));
Q_MX03 U1431 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[109]), .A1(ififoRdata[173]), .A2(n6400), .Z(iData[45]));
Q_MX03 U1432 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[108]), .A1(ififoRdata[172]), .A2(n6399), .Z(iData[44]));
Q_MX03 U1433 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[107]), .A1(ififoRdata[171]), .A2(n6398), .Z(iData[43]));
Q_MX03 U1434 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[106]), .A1(ififoRdata[170]), .A2(n6397), .Z(iData[42]));
Q_MX03 U1435 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[105]), .A1(ififoRdata[169]), .A2(n6396), .Z(iData[41]));
Q_MX03 U1436 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[104]), .A1(ififoRdata[168]), .A2(n6395), .Z(iData[40]));
Q_MX03 U1437 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[103]), .A1(ififoRdata[167]), .A2(n6394), .Z(iData[39]));
Q_MX03 U1438 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[102]), .A1(ififoRdata[166]), .A2(n6393), .Z(iData[38]));
Q_MX03 U1439 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[101]), .A1(ififoRdata[165]), .A2(n6392), .Z(iData[37]));
Q_MX03 U1440 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[100]), .A1(ififoRdata[164]), .A2(n6391), .Z(iData[36]));
Q_MX03 U1441 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[99]), .A1(ififoRdata[163]), .A2(n6390), .Z(iData[35]));
Q_MX03 U1442 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[98]), .A1(ififoRdata[162]), .A2(n6389), .Z(iData[34]));
Q_MX03 U1443 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[97]), .A1(ififoRdata[161]), .A2(n6388), .Z(iData[33]));
Q_MX03 U1444 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[96]), .A1(ififoRdata[160]), .A2(n6387), .Z(iData[32]));
Q_MX03 U1445 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[95]), .A1(ififoRdata[159]), .A2(n6386), .Z(iData[31]));
Q_MX03 U1446 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[94]), .A1(ififoRdata[158]), .A2(n6385), .Z(iData[30]));
Q_MX03 U1447 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[93]), .A1(ififoRdata[157]), .A2(n6384), .Z(iData[29]));
Q_MX03 U1448 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[92]), .A1(ififoRdata[156]), .A2(n6383), .Z(iData[28]));
Q_MX03 U1449 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[91]), .A1(ififoRdata[155]), .A2(n6382), .Z(iData[27]));
Q_MX03 U1450 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[90]), .A1(ififoRdata[154]), .A2(n6381), .Z(iData[26]));
Q_MX03 U1451 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[89]), .A1(ififoRdata[153]), .A2(n6380), .Z(iData[25]));
Q_MX03 U1452 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[88]), .A1(ififoRdata[152]), .A2(n6379), .Z(iData[24]));
Q_MX03 U1453 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[87]), .A1(ififoRdata[151]), .A2(n6378), .Z(iData[23]));
Q_MX03 U1454 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[86]), .A1(ififoRdata[150]), .A2(n6377), .Z(iData[22]));
Q_MX03 U1455 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[85]), .A1(ififoRdata[149]), .A2(n6376), .Z(iData[21]));
Q_MX03 U1456 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[84]), .A1(ififoRdata[148]), .A2(n6375), .Z(iData[20]));
Q_MX03 U1457 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[83]), .A1(ififoRdata[147]), .A2(n6374), .Z(iData[19]));
Q_MX03 U1458 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[82]), .A1(ififoRdata[146]), .A2(n6373), .Z(iData[18]));
Q_MX03 U1459 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[81]), .A1(ififoRdata[145]), .A2(n6372), .Z(iData[17]));
Q_MX03 U1460 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[80]), .A1(ififoRdata[144]), .A2(n6371), .Z(iData[16]));
Q_MX03 U1461 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[79]), .A1(ififoRdata[143]), .A2(n6370), .Z(iData[15]));
Q_MX03 U1462 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[78]), .A1(ififoRdata[142]), .A2(n6369), .Z(iData[14]));
Q_MX03 U1463 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[77]), .A1(ififoRdata[141]), .A2(n6368), .Z(iData[13]));
Q_MX03 U1464 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[76]), .A1(ififoRdata[140]), .A2(n6367), .Z(iData[12]));
Q_MX03 U1465 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[75]), .A1(ififoRdata[139]), .A2(n6366), .Z(iData[11]));
Q_MX03 U1466 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[74]), .A1(ififoRdata[138]), .A2(n6365), .Z(iData[10]));
Q_MX03 U1467 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[73]), .A1(ififoRdata[137]), .A2(n6364), .Z(iData[9]));
Q_MX03 U1468 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[72]), .A1(ififoRdata[136]), .A2(n6363), .Z(iData[8]));
Q_MX03 U1469 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[71]), .A1(ififoRdata[135]), .A2(n6362), .Z(iData[7]));
Q_MX03 U1470 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[70]), .A1(ififoRdata[134]), .A2(n6361), .Z(iData[6]));
Q_MX03 U1471 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[69]), .A1(ififoRdata[133]), .A2(n6360), .Z(iData[5]));
Q_MX03 U1472 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[68]), .A1(ififoRdata[132]), .A2(n6359), .Z(iData[4]));
Q_MX03 U1473 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[67]), .A1(ififoRdata[131]), .A2(n6358), .Z(iData[3]));
Q_MX03 U1474 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[66]), .A1(ififoRdata[130]), .A2(n6357), .Z(iData[2]));
Q_MX03 U1475 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[65]), .A1(ififoRdata[129]), .A2(n6356), .Z(iData[1]));
Q_MX03 U1476 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[64]), .A1(ififoRdata[128]), .A2(n6355), .Z(iData[0]));
Q_MX03 U1477 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[63]), .A1(ififoRdata[127]), .A2(n6354), .Z(xhead[63]));
Q_MX03 U1478 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[62]), .A1(ififoRdata[126]), .A2(n6353), .Z(xhead[62]));
Q_MX03 U1479 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[61]), .A1(ififoRdata[125]), .A2(n6352), .Z(xhead[61]));
Q_MX03 U1480 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[60]), .A1(ififoRdata[124]), .A2(n6351), .Z(xhead[60]));
Q_MX03 U1481 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[59]), .A1(ififoRdata[123]), .A2(n6350), .Z(xhead[59]));
Q_MX03 U1482 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[58]), .A1(ififoRdata[122]), .A2(n6349), .Z(xhead[58]));
Q_MX03 U1483 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[57]), .A1(ififoRdata[121]), .A2(n6348), .Z(xhead[57]));
Q_MX03 U1484 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[56]), .A1(ififoRdata[120]), .A2(n6347), .Z(xhead[56]));
Q_MX03 U1485 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[55]), .A1(ififoRdata[119]), .A2(n6346), .Z(xhead[55]));
Q_MX03 U1486 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[54]), .A1(ififoRdata[118]), .A2(n6345), .Z(xhead[54]));
Q_MX03 U1487 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[53]), .A1(ififoRdata[117]), .A2(n6344), .Z(xhead[53]));
Q_MX03 U1488 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[52]), .A1(ififoRdata[116]), .A2(n6343), .Z(xhead[52]));
Q_MX03 U1489 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[51]), .A1(ififoRdata[115]), .A2(n6342), .Z(xhead[51]));
Q_MX03 U1490 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[50]), .A1(ififoRdata[114]), .A2(n6341), .Z(xhead[50]));
Q_MX03 U1491 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[49]), .A1(ififoRdata[113]), .A2(n6340), .Z(xhead[49]));
Q_MX03 U1492 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[48]), .A1(ififoRdata[112]), .A2(n6339), .Z(xhead[48]));
Q_MX03 U1493 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[47]), .A1(ififoRdata[111]), .A2(n6338), .Z(xhead[47]));
Q_MX03 U1494 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[46]), .A1(ififoRdata[110]), .A2(n6337), .Z(xhead[46]));
Q_MX03 U1495 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[45]), .A1(ififoRdata[109]), .A2(n6336), .Z(xhead[45]));
Q_MX03 U1496 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[44]), .A1(ififoRdata[108]), .A2(n6335), .Z(xhead[44]));
Q_MX03 U1497 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[43]), .A1(ififoRdata[107]), .A2(n6334), .Z(xhead[43]));
Q_MX03 U1498 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[42]), .A1(ififoRdata[106]), .A2(n6333), .Z(xhead[42]));
Q_MX03 U1499 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[41]), .A1(ififoRdata[105]), .A2(n6332), .Z(xhead[41]));
Q_MX03 U1500 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[40]), .A1(ififoRdata[104]), .A2(n6331), .Z(xhead[40]));
Q_MX03 U1501 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[39]), .A1(ififoRdata[103]), .A2(n6330), .Z(xhead[39]));
Q_MX03 U1502 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[38]), .A1(ififoRdata[102]), .A2(n6329), .Z(xhead[38]));
Q_MX03 U1503 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[37]), .A1(ififoRdata[101]), .A2(n6328), .Z(xhead[37]));
Q_MX03 U1504 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[36]), .A1(ififoRdata[100]), .A2(n6327), .Z(xhead[36]));
Q_MX03 U1505 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[35]), .A1(ififoRdata[99]), .A2(n6326), .Z(xhead[35]));
Q_MX03 U1506 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[34]), .A1(ififoRdata[98]), .A2(n6325), .Z(xhead[34]));
Q_MX03 U1507 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[33]), .A1(ififoRdata[97]), .A2(n6324), .Z(xhead[33]));
Q_MX03 U1508 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[32]), .A1(ififoRdata[96]), .A2(n6323), .Z(xhead[32]));
Q_MX03 U1509 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[31]), .A1(ififoRdata[95]), .A2(n6322), .Z(xhead[31]));
Q_MX03 U1510 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[30]), .A1(ififoRdata[94]), .A2(n6321), .Z(xhead[30]));
Q_MX03 U1511 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[29]), .A1(ififoRdata[93]), .A2(n6320), .Z(xhead[29]));
Q_MX03 U1512 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[28]), .A1(ififoRdata[92]), .A2(n6319), .Z(xhead[28]));
Q_MX03 U1513 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[27]), .A1(ififoRdata[91]), .A2(n6318), .Z(xhead[27]));
Q_MX03 U1514 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[26]), .A1(ififoRdata[90]), .A2(n6317), .Z(xhead[26]));
Q_MX03 U1515 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[25]), .A1(ififoRdata[89]), .A2(n6316), .Z(xhead[25]));
Q_MX03 U1516 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[24]), .A1(ififoRdata[88]), .A2(n6315), .Z(xhead[24]));
Q_MX03 U1517 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[23]), .A1(ififoRdata[87]), .A2(n6314), .Z(xhead[23]));
Q_MX03 U1518 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[22]), .A1(ififoRdata[86]), .A2(n6313), .Z(xhead[22]));
Q_MX03 U1519 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[21]), .A1(ififoRdata[85]), .A2(n6312), .Z(xhead[21]));
Q_MX03 U1520 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[20]), .A1(ififoRdata[84]), .A2(n6311), .Z(xhead[20]));
Q_MX03 U1521 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[19]), .A1(ififoRdata[83]), .A2(n6310), .Z(xhead[19]));
Q_MX03 U1522 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[18]), .A1(ififoRdata[82]), .A2(n6309), .Z(xhead[18]));
Q_MX03 U1523 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[17]), .A1(ififoRdata[81]), .A2(n6308), .Z(xhead[17]));
Q_MX03 U1524 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[16]), .A1(ififoRdata[80]), .A2(n6307), .Z(xhead[16]));
Q_MX03 U1525 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[15]), .A1(ififoRdata[79]), .A2(n6306), .Z(xhead[15]));
Q_MX03 U1526 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[14]), .A1(ififoRdata[78]), .A2(n6305), .Z(xhead[14]));
Q_MX03 U1527 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[13]), .A1(ififoRdata[77]), .A2(n6304), .Z(xhead[13]));
Q_MX03 U1528 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[12]), .A1(ififoRdata[76]), .A2(n6303), .Z(xhead[12]));
Q_MX03 U1529 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[11]), .A1(ififoRdata[75]), .A2(n6302), .Z(xhead[11]));
Q_MX03 U1530 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[10]), .A1(ififoRdata[74]), .A2(n6301), .Z(xhead[10]));
Q_MX03 U1531 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[9]), .A1(ififoRdata[73]), .A2(n6300), .Z(xhead[9]));
Q_MX03 U1532 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[8]), .A1(ififoRdata[72]), .A2(n6299), .Z(xhead[8]));
Q_MX03 U1533 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[7]), .A1(ififoRdata[71]), .A2(n6298), .Z(xhead[7]));
Q_MX03 U1534 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[6]), .A1(ififoRdata[70]), .A2(n6297), .Z(xhead[6]));
Q_MX03 U1535 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[5]), .A1(ififoRdata[69]), .A2(n6296), .Z(xhead[5]));
Q_MX03 U1536 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[4]), .A1(ififoRdata[68]), .A2(n6295), .Z(xhead[4]));
Q_MX03 U1537 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[3]), .A1(ififoRdata[67]), .A2(n6294), .Z(xhead[3]));
Q_MX03 U1538 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[2]), .A1(ififoRdata[66]), .A2(n6293), .Z(xhead[2]));
Q_MX03 U1539 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[1]), .A1(ififoRdata[65]), .A2(n6292), .Z(xhead[1]));
Q_MX03 U1540 ( .S0(rptr[0]), .S1(rptr[1]), .A0(ififoRdata[0]), .A1(ififoRdata[64]), .A2(n6291), .Z(xhead[0]));
Q_MX02 U1541 ( .S(rptr[0]), .A0(ififoRdata[703]), .A1(ififoRdata[767]), .Z(n6866));
Q_MX02 U1542 ( .S(rptr[0]), .A0(ififoRdata[702]), .A1(ififoRdata[766]), .Z(n6865));
Q_MX02 U1543 ( .S(rptr[0]), .A0(ififoRdata[701]), .A1(ififoRdata[765]), .Z(n6864));
Q_MX02 U1544 ( .S(rptr[0]), .A0(ififoRdata[700]), .A1(ififoRdata[764]), .Z(n6863));
Q_MX02 U1545 ( .S(rptr[0]), .A0(ififoRdata[699]), .A1(ififoRdata[763]), .Z(n6862));
Q_MX02 U1546 ( .S(rptr[0]), .A0(ififoRdata[698]), .A1(ififoRdata[762]), .Z(n6861));
Q_MX02 U1547 ( .S(rptr[0]), .A0(ififoRdata[697]), .A1(ififoRdata[761]), .Z(n6860));
Q_MX02 U1548 ( .S(rptr[0]), .A0(ififoRdata[696]), .A1(ififoRdata[760]), .Z(n6859));
Q_MX02 U1549 ( .S(rptr[0]), .A0(ififoRdata[695]), .A1(ififoRdata[759]), .Z(n6858));
Q_MX02 U1550 ( .S(rptr[0]), .A0(ififoRdata[694]), .A1(ififoRdata[758]), .Z(n6857));
Q_MX02 U1551 ( .S(rptr[0]), .A0(ififoRdata[693]), .A1(ififoRdata[757]), .Z(n6856));
Q_MX02 U1552 ( .S(rptr[0]), .A0(ififoRdata[692]), .A1(ififoRdata[756]), .Z(n6855));
Q_MX02 U1553 ( .S(rptr[0]), .A0(ififoRdata[691]), .A1(ififoRdata[755]), .Z(n6854));
Q_MX02 U1554 ( .S(rptr[0]), .A0(ififoRdata[690]), .A1(ififoRdata[754]), .Z(n6853));
Q_MX02 U1555 ( .S(rptr[0]), .A0(ififoRdata[689]), .A1(ififoRdata[753]), .Z(n6852));
Q_MX02 U1556 ( .S(rptr[0]), .A0(ififoRdata[688]), .A1(ififoRdata[752]), .Z(n6851));
Q_MX02 U1557 ( .S(rptr[0]), .A0(ififoRdata[687]), .A1(ififoRdata[751]), .Z(n6850));
Q_MX02 U1558 ( .S(rptr[0]), .A0(ififoRdata[686]), .A1(ififoRdata[750]), .Z(n6849));
Q_MX02 U1559 ( .S(rptr[0]), .A0(ififoRdata[685]), .A1(ififoRdata[749]), .Z(n6848));
Q_MX02 U1560 ( .S(rptr[0]), .A0(ififoRdata[684]), .A1(ififoRdata[748]), .Z(n6847));
Q_MX02 U1561 ( .S(rptr[0]), .A0(ififoRdata[683]), .A1(ififoRdata[747]), .Z(n6846));
Q_MX02 U1562 ( .S(rptr[0]), .A0(ififoRdata[682]), .A1(ififoRdata[746]), .Z(n6845));
Q_MX02 U1563 ( .S(rptr[0]), .A0(ififoRdata[681]), .A1(ififoRdata[745]), .Z(n6844));
Q_MX02 U1564 ( .S(rptr[0]), .A0(ififoRdata[680]), .A1(ififoRdata[744]), .Z(n6843));
Q_MX02 U1565 ( .S(rptr[0]), .A0(ififoRdata[679]), .A1(ififoRdata[743]), .Z(n6842));
Q_MX02 U1566 ( .S(rptr[0]), .A0(ififoRdata[678]), .A1(ififoRdata[742]), .Z(n6841));
Q_MX02 U1567 ( .S(rptr[0]), .A0(ififoRdata[677]), .A1(ififoRdata[741]), .Z(n6840));
Q_MX02 U1568 ( .S(rptr[0]), .A0(ififoRdata[676]), .A1(ififoRdata[740]), .Z(n6839));
Q_MX02 U1569 ( .S(rptr[0]), .A0(ififoRdata[675]), .A1(ififoRdata[739]), .Z(n6838));
Q_MX02 U1570 ( .S(rptr[0]), .A0(ififoRdata[674]), .A1(ififoRdata[738]), .Z(n6837));
Q_MX02 U1571 ( .S(rptr[0]), .A0(ififoRdata[673]), .A1(ififoRdata[737]), .Z(n6836));
Q_MX02 U1572 ( .S(rptr[0]), .A0(ififoRdata[672]), .A1(ififoRdata[736]), .Z(n6835));
Q_MX02 U1573 ( .S(rptr[0]), .A0(ififoRdata[671]), .A1(ififoRdata[735]), .Z(n6834));
Q_MX02 U1574 ( .S(rptr[0]), .A0(ififoRdata[670]), .A1(ififoRdata[734]), .Z(n6833));
Q_MX02 U1575 ( .S(rptr[0]), .A0(ififoRdata[669]), .A1(ififoRdata[733]), .Z(n6832));
Q_MX02 U1576 ( .S(rptr[0]), .A0(ififoRdata[668]), .A1(ififoRdata[732]), .Z(n6831));
Q_MX02 U1577 ( .S(rptr[0]), .A0(ififoRdata[667]), .A1(ififoRdata[731]), .Z(n6830));
Q_MX02 U1578 ( .S(rptr[0]), .A0(ififoRdata[666]), .A1(ififoRdata[730]), .Z(n6829));
Q_MX02 U1579 ( .S(rptr[0]), .A0(ififoRdata[665]), .A1(ififoRdata[729]), .Z(n6828));
Q_MX02 U1580 ( .S(rptr[0]), .A0(ififoRdata[664]), .A1(ififoRdata[728]), .Z(n6827));
Q_MX02 U1581 ( .S(rptr[0]), .A0(ififoRdata[663]), .A1(ififoRdata[727]), .Z(n6826));
Q_MX02 U1582 ( .S(rptr[0]), .A0(ififoRdata[662]), .A1(ififoRdata[726]), .Z(n6825));
Q_MX02 U1583 ( .S(rptr[0]), .A0(ififoRdata[661]), .A1(ififoRdata[725]), .Z(n6824));
Q_MX02 U1584 ( .S(rptr[0]), .A0(ififoRdata[660]), .A1(ififoRdata[724]), .Z(n6823));
Q_MX02 U1585 ( .S(rptr[0]), .A0(ififoRdata[659]), .A1(ififoRdata[723]), .Z(n6822));
Q_MX02 U1586 ( .S(rptr[0]), .A0(ififoRdata[658]), .A1(ififoRdata[722]), .Z(n6821));
Q_MX02 U1587 ( .S(rptr[0]), .A0(ififoRdata[657]), .A1(ififoRdata[721]), .Z(n6820));
Q_MX02 U1588 ( .S(rptr[0]), .A0(ififoRdata[656]), .A1(ififoRdata[720]), .Z(n6819));
Q_MX02 U1589 ( .S(rptr[0]), .A0(ififoRdata[655]), .A1(ififoRdata[719]), .Z(n6818));
Q_MX02 U1590 ( .S(rptr[0]), .A0(ififoRdata[654]), .A1(ififoRdata[718]), .Z(n6817));
Q_MX02 U1591 ( .S(rptr[0]), .A0(ififoRdata[653]), .A1(ififoRdata[717]), .Z(n6816));
Q_MX02 U1592 ( .S(rptr[0]), .A0(ififoRdata[652]), .A1(ififoRdata[716]), .Z(n6815));
Q_MX02 U1593 ( .S(rptr[0]), .A0(ififoRdata[651]), .A1(ififoRdata[715]), .Z(n6814));
Q_MX02 U1594 ( .S(rptr[0]), .A0(ififoRdata[650]), .A1(ififoRdata[714]), .Z(n6813));
Q_MX02 U1595 ( .S(rptr[0]), .A0(ififoRdata[649]), .A1(ififoRdata[713]), .Z(n6812));
Q_MX02 U1596 ( .S(rptr[0]), .A0(ififoRdata[648]), .A1(ififoRdata[712]), .Z(n6811));
Q_MX02 U1597 ( .S(rptr[0]), .A0(ififoRdata[647]), .A1(ififoRdata[711]), .Z(n6810));
Q_MX02 U1598 ( .S(rptr[0]), .A0(ififoRdata[646]), .A1(ififoRdata[710]), .Z(n6809));
Q_MX02 U1599 ( .S(rptr[0]), .A0(ififoRdata[645]), .A1(ififoRdata[709]), .Z(n6808));
Q_MX02 U1600 ( .S(rptr[0]), .A0(ififoRdata[644]), .A1(ififoRdata[708]), .Z(n6807));
Q_MX02 U1601 ( .S(rptr[0]), .A0(ififoRdata[643]), .A1(ififoRdata[707]), .Z(n6806));
Q_MX02 U1602 ( .S(rptr[0]), .A0(ififoRdata[642]), .A1(ififoRdata[706]), .Z(n6805));
Q_MX02 U1603 ( .S(rptr[0]), .A0(ififoRdata[641]), .A1(ififoRdata[705]), .Z(n6804));
Q_MX02 U1604 ( .S(rptr[0]), .A0(ififoRdata[640]), .A1(ififoRdata[704]), .Z(n6803));
Q_MX02 U1605 ( .S(rptr[0]), .A0(ififoRdata[639]), .A1(ififoRdata[703]), .Z(n6802));
Q_MX02 U1606 ( .S(rptr[0]), .A0(ififoRdata[638]), .A1(ififoRdata[702]), .Z(n6801));
Q_MX02 U1607 ( .S(rptr[0]), .A0(ififoRdata[637]), .A1(ififoRdata[701]), .Z(n6800));
Q_MX02 U1608 ( .S(rptr[0]), .A0(ififoRdata[636]), .A1(ififoRdata[700]), .Z(n6799));
Q_MX02 U1609 ( .S(rptr[0]), .A0(ififoRdata[635]), .A1(ififoRdata[699]), .Z(n6798));
Q_MX02 U1610 ( .S(rptr[0]), .A0(ififoRdata[634]), .A1(ififoRdata[698]), .Z(n6797));
Q_MX02 U1611 ( .S(rptr[0]), .A0(ififoRdata[633]), .A1(ififoRdata[697]), .Z(n6796));
Q_MX02 U1612 ( .S(rptr[0]), .A0(ififoRdata[632]), .A1(ififoRdata[696]), .Z(n6795));
Q_MX02 U1613 ( .S(rptr[0]), .A0(ififoRdata[631]), .A1(ififoRdata[695]), .Z(n6794));
Q_MX02 U1614 ( .S(rptr[0]), .A0(ififoRdata[630]), .A1(ififoRdata[694]), .Z(n6793));
Q_MX02 U1615 ( .S(rptr[0]), .A0(ififoRdata[629]), .A1(ififoRdata[693]), .Z(n6792));
Q_MX02 U1616 ( .S(rptr[0]), .A0(ififoRdata[628]), .A1(ififoRdata[692]), .Z(n6791));
Q_MX02 U1617 ( .S(rptr[0]), .A0(ififoRdata[627]), .A1(ififoRdata[691]), .Z(n6790));
Q_MX02 U1618 ( .S(rptr[0]), .A0(ififoRdata[626]), .A1(ififoRdata[690]), .Z(n6789));
Q_MX02 U1619 ( .S(rptr[0]), .A0(ififoRdata[625]), .A1(ififoRdata[689]), .Z(n6788));
Q_MX02 U1620 ( .S(rptr[0]), .A0(ififoRdata[624]), .A1(ififoRdata[688]), .Z(n6787));
Q_MX02 U1621 ( .S(rptr[0]), .A0(ififoRdata[623]), .A1(ififoRdata[687]), .Z(n6786));
Q_MX02 U1622 ( .S(rptr[0]), .A0(ififoRdata[622]), .A1(ififoRdata[686]), .Z(n6785));
Q_MX02 U1623 ( .S(rptr[0]), .A0(ififoRdata[621]), .A1(ififoRdata[685]), .Z(n6784));
Q_MX02 U1624 ( .S(rptr[0]), .A0(ififoRdata[620]), .A1(ififoRdata[684]), .Z(n6783));
Q_MX02 U1625 ( .S(rptr[0]), .A0(ififoRdata[619]), .A1(ififoRdata[683]), .Z(n6782));
Q_MX02 U1626 ( .S(rptr[0]), .A0(ififoRdata[618]), .A1(ififoRdata[682]), .Z(n6781));
Q_MX02 U1627 ( .S(rptr[0]), .A0(ififoRdata[617]), .A1(ififoRdata[681]), .Z(n6780));
Q_MX02 U1628 ( .S(rptr[0]), .A0(ififoRdata[616]), .A1(ififoRdata[680]), .Z(n6779));
Q_MX02 U1629 ( .S(rptr[0]), .A0(ififoRdata[615]), .A1(ififoRdata[679]), .Z(n6778));
Q_MX02 U1630 ( .S(rptr[0]), .A0(ififoRdata[614]), .A1(ififoRdata[678]), .Z(n6777));
Q_MX02 U1631 ( .S(rptr[0]), .A0(ififoRdata[613]), .A1(ififoRdata[677]), .Z(n6776));
Q_MX02 U1632 ( .S(rptr[0]), .A0(ififoRdata[612]), .A1(ififoRdata[676]), .Z(n6775));
Q_MX02 U1633 ( .S(rptr[0]), .A0(ififoRdata[611]), .A1(ififoRdata[675]), .Z(n6774));
Q_MX02 U1634 ( .S(rptr[0]), .A0(ififoRdata[610]), .A1(ififoRdata[674]), .Z(n6773));
Q_MX02 U1635 ( .S(rptr[0]), .A0(ififoRdata[609]), .A1(ififoRdata[673]), .Z(n6772));
Q_MX02 U1636 ( .S(rptr[0]), .A0(ififoRdata[608]), .A1(ififoRdata[672]), .Z(n6771));
Q_MX02 U1637 ( .S(rptr[0]), .A0(ififoRdata[607]), .A1(ififoRdata[671]), .Z(n6770));
Q_MX02 U1638 ( .S(rptr[0]), .A0(ififoRdata[606]), .A1(ififoRdata[670]), .Z(n6769));
Q_MX02 U1639 ( .S(rptr[0]), .A0(ififoRdata[605]), .A1(ififoRdata[669]), .Z(n6768));
Q_MX02 U1640 ( .S(rptr[0]), .A0(ififoRdata[604]), .A1(ififoRdata[668]), .Z(n6767));
Q_MX02 U1641 ( .S(rptr[0]), .A0(ififoRdata[603]), .A1(ififoRdata[667]), .Z(n6766));
Q_MX02 U1642 ( .S(rptr[0]), .A0(ififoRdata[602]), .A1(ififoRdata[666]), .Z(n6765));
Q_MX02 U1643 ( .S(rptr[0]), .A0(ififoRdata[601]), .A1(ififoRdata[665]), .Z(n6764));
Q_MX02 U1644 ( .S(rptr[0]), .A0(ififoRdata[600]), .A1(ififoRdata[664]), .Z(n6763));
Q_MX02 U1645 ( .S(rptr[0]), .A0(ififoRdata[599]), .A1(ififoRdata[663]), .Z(n6762));
Q_MX02 U1646 ( .S(rptr[0]), .A0(ififoRdata[598]), .A1(ififoRdata[662]), .Z(n6761));
Q_MX02 U1647 ( .S(rptr[0]), .A0(ififoRdata[597]), .A1(ififoRdata[661]), .Z(n6760));
Q_MX02 U1648 ( .S(rptr[0]), .A0(ififoRdata[596]), .A1(ififoRdata[660]), .Z(n6759));
Q_MX02 U1649 ( .S(rptr[0]), .A0(ififoRdata[595]), .A1(ififoRdata[659]), .Z(n6758));
Q_MX02 U1650 ( .S(rptr[0]), .A0(ififoRdata[594]), .A1(ififoRdata[658]), .Z(n6757));
Q_MX02 U1651 ( .S(rptr[0]), .A0(ififoRdata[593]), .A1(ififoRdata[657]), .Z(n6756));
Q_MX02 U1652 ( .S(rptr[0]), .A0(ififoRdata[592]), .A1(ififoRdata[656]), .Z(n6755));
Q_MX02 U1653 ( .S(rptr[0]), .A0(ififoRdata[591]), .A1(ififoRdata[655]), .Z(n6754));
Q_MX02 U1654 ( .S(rptr[0]), .A0(ififoRdata[590]), .A1(ififoRdata[654]), .Z(n6753));
Q_MX02 U1655 ( .S(rptr[0]), .A0(ififoRdata[589]), .A1(ififoRdata[653]), .Z(n6752));
Q_MX02 U1656 ( .S(rptr[0]), .A0(ififoRdata[588]), .A1(ififoRdata[652]), .Z(n6751));
Q_MX02 U1657 ( .S(rptr[0]), .A0(ififoRdata[587]), .A1(ififoRdata[651]), .Z(n6750));
Q_MX02 U1658 ( .S(rptr[0]), .A0(ififoRdata[586]), .A1(ififoRdata[650]), .Z(n6749));
Q_MX02 U1659 ( .S(rptr[0]), .A0(ififoRdata[585]), .A1(ififoRdata[649]), .Z(n6748));
Q_MX02 U1660 ( .S(rptr[0]), .A0(ififoRdata[584]), .A1(ififoRdata[648]), .Z(n6747));
Q_MX02 U1661 ( .S(rptr[0]), .A0(ififoRdata[583]), .A1(ififoRdata[647]), .Z(n6746));
Q_MX02 U1662 ( .S(rptr[0]), .A0(ififoRdata[582]), .A1(ififoRdata[646]), .Z(n6745));
Q_MX02 U1663 ( .S(rptr[0]), .A0(ififoRdata[581]), .A1(ififoRdata[645]), .Z(n6744));
Q_MX02 U1664 ( .S(rptr[0]), .A0(ififoRdata[580]), .A1(ififoRdata[644]), .Z(n6743));
Q_MX02 U1665 ( .S(rptr[0]), .A0(ififoRdata[579]), .A1(ififoRdata[643]), .Z(n6742));
Q_MX02 U1666 ( .S(rptr[0]), .A0(ififoRdata[578]), .A1(ififoRdata[642]), .Z(n6741));
Q_MX02 U1667 ( .S(rptr[0]), .A0(ififoRdata[577]), .A1(ififoRdata[641]), .Z(n6740));
Q_MX02 U1668 ( .S(rptr[0]), .A0(ififoRdata[576]), .A1(ififoRdata[640]), .Z(n6739));
Q_MX02 U1669 ( .S(rptr[0]), .A0(ififoRdata[575]), .A1(ififoRdata[639]), .Z(n6738));
Q_MX02 U1670 ( .S(rptr[0]), .A0(ififoRdata[574]), .A1(ififoRdata[638]), .Z(n6737));
Q_MX02 U1671 ( .S(rptr[0]), .A0(ififoRdata[573]), .A1(ififoRdata[637]), .Z(n6736));
Q_MX02 U1672 ( .S(rptr[0]), .A0(ififoRdata[572]), .A1(ififoRdata[636]), .Z(n6735));
Q_MX02 U1673 ( .S(rptr[0]), .A0(ififoRdata[571]), .A1(ififoRdata[635]), .Z(n6734));
Q_MX02 U1674 ( .S(rptr[0]), .A0(ififoRdata[570]), .A1(ififoRdata[634]), .Z(n6733));
Q_MX02 U1675 ( .S(rptr[0]), .A0(ififoRdata[569]), .A1(ififoRdata[633]), .Z(n6732));
Q_MX02 U1676 ( .S(rptr[0]), .A0(ififoRdata[568]), .A1(ififoRdata[632]), .Z(n6731));
Q_MX02 U1677 ( .S(rptr[0]), .A0(ififoRdata[567]), .A1(ififoRdata[631]), .Z(n6730));
Q_MX02 U1678 ( .S(rptr[0]), .A0(ififoRdata[566]), .A1(ififoRdata[630]), .Z(n6729));
Q_MX02 U1679 ( .S(rptr[0]), .A0(ififoRdata[565]), .A1(ififoRdata[629]), .Z(n6728));
Q_MX02 U1680 ( .S(rptr[0]), .A0(ififoRdata[564]), .A1(ififoRdata[628]), .Z(n6727));
Q_MX02 U1681 ( .S(rptr[0]), .A0(ififoRdata[563]), .A1(ififoRdata[627]), .Z(n6726));
Q_MX02 U1682 ( .S(rptr[0]), .A0(ififoRdata[562]), .A1(ififoRdata[626]), .Z(n6725));
Q_MX02 U1683 ( .S(rptr[0]), .A0(ififoRdata[561]), .A1(ififoRdata[625]), .Z(n6724));
Q_MX02 U1684 ( .S(rptr[0]), .A0(ififoRdata[560]), .A1(ififoRdata[624]), .Z(n6723));
Q_MX02 U1685 ( .S(rptr[0]), .A0(ififoRdata[559]), .A1(ififoRdata[623]), .Z(n6722));
Q_MX02 U1686 ( .S(rptr[0]), .A0(ififoRdata[558]), .A1(ififoRdata[622]), .Z(n6721));
Q_MX02 U1687 ( .S(rptr[0]), .A0(ififoRdata[557]), .A1(ififoRdata[621]), .Z(n6720));
Q_MX02 U1688 ( .S(rptr[0]), .A0(ififoRdata[556]), .A1(ififoRdata[620]), .Z(n6719));
Q_MX02 U1689 ( .S(rptr[0]), .A0(ififoRdata[555]), .A1(ififoRdata[619]), .Z(n6718));
Q_MX02 U1690 ( .S(rptr[0]), .A0(ififoRdata[554]), .A1(ififoRdata[618]), .Z(n6717));
Q_MX02 U1691 ( .S(rptr[0]), .A0(ififoRdata[553]), .A1(ififoRdata[617]), .Z(n6716));
Q_MX02 U1692 ( .S(rptr[0]), .A0(ififoRdata[552]), .A1(ififoRdata[616]), .Z(n6715));
Q_MX02 U1693 ( .S(rptr[0]), .A0(ififoRdata[551]), .A1(ififoRdata[615]), .Z(n6714));
Q_MX02 U1694 ( .S(rptr[0]), .A0(ififoRdata[550]), .A1(ififoRdata[614]), .Z(n6713));
Q_MX02 U1695 ( .S(rptr[0]), .A0(ififoRdata[549]), .A1(ififoRdata[613]), .Z(n6712));
Q_MX02 U1696 ( .S(rptr[0]), .A0(ififoRdata[548]), .A1(ififoRdata[612]), .Z(n6711));
Q_MX02 U1697 ( .S(rptr[0]), .A0(ififoRdata[547]), .A1(ififoRdata[611]), .Z(n6710));
Q_MX02 U1698 ( .S(rptr[0]), .A0(ififoRdata[546]), .A1(ififoRdata[610]), .Z(n6709));
Q_MX02 U1699 ( .S(rptr[0]), .A0(ififoRdata[545]), .A1(ififoRdata[609]), .Z(n6708));
Q_MX02 U1700 ( .S(rptr[0]), .A0(ififoRdata[544]), .A1(ififoRdata[608]), .Z(n6707));
Q_MX02 U1701 ( .S(rptr[0]), .A0(ififoRdata[543]), .A1(ififoRdata[607]), .Z(n6706));
Q_MX02 U1702 ( .S(rptr[0]), .A0(ififoRdata[542]), .A1(ififoRdata[606]), .Z(n6705));
Q_MX02 U1703 ( .S(rptr[0]), .A0(ififoRdata[541]), .A1(ififoRdata[605]), .Z(n6704));
Q_MX02 U1704 ( .S(rptr[0]), .A0(ififoRdata[540]), .A1(ififoRdata[604]), .Z(n6703));
Q_MX02 U1705 ( .S(rptr[0]), .A0(ififoRdata[539]), .A1(ififoRdata[603]), .Z(n6702));
Q_MX02 U1706 ( .S(rptr[0]), .A0(ififoRdata[538]), .A1(ififoRdata[602]), .Z(n6701));
Q_MX02 U1707 ( .S(rptr[0]), .A0(ififoRdata[537]), .A1(ififoRdata[601]), .Z(n6700));
Q_MX02 U1708 ( .S(rptr[0]), .A0(ififoRdata[536]), .A1(ififoRdata[600]), .Z(n6699));
Q_MX02 U1709 ( .S(rptr[0]), .A0(ififoRdata[535]), .A1(ififoRdata[599]), .Z(n6698));
Q_MX02 U1710 ( .S(rptr[0]), .A0(ififoRdata[534]), .A1(ififoRdata[598]), .Z(n6697));
Q_MX02 U1711 ( .S(rptr[0]), .A0(ififoRdata[533]), .A1(ififoRdata[597]), .Z(n6696));
Q_MX02 U1712 ( .S(rptr[0]), .A0(ififoRdata[532]), .A1(ififoRdata[596]), .Z(n6695));
Q_MX02 U1713 ( .S(rptr[0]), .A0(ififoRdata[531]), .A1(ififoRdata[595]), .Z(n6694));
Q_MX02 U1714 ( .S(rptr[0]), .A0(ififoRdata[530]), .A1(ififoRdata[594]), .Z(n6693));
Q_MX02 U1715 ( .S(rptr[0]), .A0(ififoRdata[529]), .A1(ififoRdata[593]), .Z(n6692));
Q_MX02 U1716 ( .S(rptr[0]), .A0(ififoRdata[528]), .A1(ififoRdata[592]), .Z(n6691));
Q_MX02 U1717 ( .S(rptr[0]), .A0(ififoRdata[527]), .A1(ififoRdata[591]), .Z(n6690));
Q_MX02 U1718 ( .S(rptr[0]), .A0(ififoRdata[526]), .A1(ififoRdata[590]), .Z(n6689));
Q_MX02 U1719 ( .S(rptr[0]), .A0(ififoRdata[525]), .A1(ififoRdata[589]), .Z(n6688));
Q_MX02 U1720 ( .S(rptr[0]), .A0(ififoRdata[524]), .A1(ififoRdata[588]), .Z(n6687));
Q_MX02 U1721 ( .S(rptr[0]), .A0(ififoRdata[523]), .A1(ififoRdata[587]), .Z(n6686));
Q_MX02 U1722 ( .S(rptr[0]), .A0(ififoRdata[522]), .A1(ififoRdata[586]), .Z(n6685));
Q_MX02 U1723 ( .S(rptr[0]), .A0(ififoRdata[521]), .A1(ififoRdata[585]), .Z(n6684));
Q_MX02 U1724 ( .S(rptr[0]), .A0(ififoRdata[520]), .A1(ififoRdata[584]), .Z(n6683));
Q_MX02 U1725 ( .S(rptr[0]), .A0(ififoRdata[519]), .A1(ififoRdata[583]), .Z(n6682));
Q_MX02 U1726 ( .S(rptr[0]), .A0(ififoRdata[518]), .A1(ififoRdata[582]), .Z(n6681));
Q_MX02 U1727 ( .S(rptr[0]), .A0(ififoRdata[517]), .A1(ififoRdata[581]), .Z(n6680));
Q_MX02 U1728 ( .S(rptr[0]), .A0(ififoRdata[516]), .A1(ififoRdata[580]), .Z(n6679));
Q_MX02 U1729 ( .S(rptr[0]), .A0(ififoRdata[515]), .A1(ififoRdata[579]), .Z(n6678));
Q_MX02 U1730 ( .S(rptr[0]), .A0(ififoRdata[514]), .A1(ififoRdata[578]), .Z(n6677));
Q_MX02 U1731 ( .S(rptr[0]), .A0(ififoRdata[513]), .A1(ififoRdata[577]), .Z(n6676));
Q_MX02 U1732 ( .S(rptr[0]), .A0(ififoRdata[512]), .A1(ififoRdata[576]), .Z(n6675));
Q_MX02 U1733 ( .S(rptr[0]), .A0(ififoRdata[511]), .A1(ififoRdata[575]), .Z(n6674));
Q_MX02 U1734 ( .S(rptr[0]), .A0(ififoRdata[510]), .A1(ififoRdata[574]), .Z(n6673));
Q_MX02 U1735 ( .S(rptr[0]), .A0(ififoRdata[509]), .A1(ififoRdata[573]), .Z(n6672));
Q_MX02 U1736 ( .S(rptr[0]), .A0(ififoRdata[508]), .A1(ififoRdata[572]), .Z(n6671));
Q_MX02 U1737 ( .S(rptr[0]), .A0(ififoRdata[507]), .A1(ififoRdata[571]), .Z(n6670));
Q_MX02 U1738 ( .S(rptr[0]), .A0(ififoRdata[506]), .A1(ififoRdata[570]), .Z(n6669));
Q_MX02 U1739 ( .S(rptr[0]), .A0(ififoRdata[505]), .A1(ififoRdata[569]), .Z(n6668));
Q_MX02 U1740 ( .S(rptr[0]), .A0(ififoRdata[504]), .A1(ififoRdata[568]), .Z(n6667));
Q_MX02 U1741 ( .S(rptr[0]), .A0(ififoRdata[503]), .A1(ififoRdata[567]), .Z(n6666));
Q_MX02 U1742 ( .S(rptr[0]), .A0(ififoRdata[502]), .A1(ififoRdata[566]), .Z(n6665));
Q_MX02 U1743 ( .S(rptr[0]), .A0(ififoRdata[501]), .A1(ififoRdata[565]), .Z(n6664));
Q_MX02 U1744 ( .S(rptr[0]), .A0(ififoRdata[500]), .A1(ififoRdata[564]), .Z(n6663));
Q_MX02 U1745 ( .S(rptr[0]), .A0(ififoRdata[499]), .A1(ififoRdata[563]), .Z(n6662));
Q_MX02 U1746 ( .S(rptr[0]), .A0(ififoRdata[498]), .A1(ififoRdata[562]), .Z(n6661));
Q_MX02 U1747 ( .S(rptr[0]), .A0(ififoRdata[497]), .A1(ififoRdata[561]), .Z(n6660));
Q_MX02 U1748 ( .S(rptr[0]), .A0(ififoRdata[496]), .A1(ififoRdata[560]), .Z(n6659));
Q_MX02 U1749 ( .S(rptr[0]), .A0(ififoRdata[495]), .A1(ififoRdata[559]), .Z(n6658));
Q_MX02 U1750 ( .S(rptr[0]), .A0(ififoRdata[494]), .A1(ififoRdata[558]), .Z(n6657));
Q_MX02 U1751 ( .S(rptr[0]), .A0(ififoRdata[493]), .A1(ififoRdata[557]), .Z(n6656));
Q_MX02 U1752 ( .S(rptr[0]), .A0(ififoRdata[492]), .A1(ififoRdata[556]), .Z(n6655));
Q_MX02 U1753 ( .S(rptr[0]), .A0(ififoRdata[491]), .A1(ififoRdata[555]), .Z(n6654));
Q_MX02 U1754 ( .S(rptr[0]), .A0(ififoRdata[490]), .A1(ififoRdata[554]), .Z(n6653));
Q_MX02 U1755 ( .S(rptr[0]), .A0(ififoRdata[489]), .A1(ififoRdata[553]), .Z(n6652));
Q_MX02 U1756 ( .S(rptr[0]), .A0(ififoRdata[488]), .A1(ififoRdata[552]), .Z(n6651));
Q_MX02 U1757 ( .S(rptr[0]), .A0(ififoRdata[487]), .A1(ififoRdata[551]), .Z(n6650));
Q_MX02 U1758 ( .S(rptr[0]), .A0(ififoRdata[486]), .A1(ififoRdata[550]), .Z(n6649));
Q_MX02 U1759 ( .S(rptr[0]), .A0(ififoRdata[485]), .A1(ififoRdata[549]), .Z(n6648));
Q_MX02 U1760 ( .S(rptr[0]), .A0(ififoRdata[484]), .A1(ififoRdata[548]), .Z(n6647));
Q_MX02 U1761 ( .S(rptr[0]), .A0(ififoRdata[483]), .A1(ififoRdata[547]), .Z(n6646));
Q_MX02 U1762 ( .S(rptr[0]), .A0(ififoRdata[482]), .A1(ififoRdata[546]), .Z(n6645));
Q_MX02 U1763 ( .S(rptr[0]), .A0(ififoRdata[481]), .A1(ififoRdata[545]), .Z(n6644));
Q_MX02 U1764 ( .S(rptr[0]), .A0(ififoRdata[480]), .A1(ififoRdata[544]), .Z(n6643));
Q_MX02 U1765 ( .S(rptr[0]), .A0(ififoRdata[479]), .A1(ififoRdata[543]), .Z(n6642));
Q_MX02 U1766 ( .S(rptr[0]), .A0(ififoRdata[478]), .A1(ififoRdata[542]), .Z(n6641));
Q_MX02 U1767 ( .S(rptr[0]), .A0(ififoRdata[477]), .A1(ififoRdata[541]), .Z(n6640));
Q_MX02 U1768 ( .S(rptr[0]), .A0(ififoRdata[476]), .A1(ififoRdata[540]), .Z(n6639));
Q_MX02 U1769 ( .S(rptr[0]), .A0(ififoRdata[475]), .A1(ififoRdata[539]), .Z(n6638));
Q_MX02 U1770 ( .S(rptr[0]), .A0(ififoRdata[474]), .A1(ififoRdata[538]), .Z(n6637));
Q_MX02 U1771 ( .S(rptr[0]), .A0(ififoRdata[473]), .A1(ififoRdata[537]), .Z(n6636));
Q_MX02 U1772 ( .S(rptr[0]), .A0(ififoRdata[472]), .A1(ififoRdata[536]), .Z(n6635));
Q_MX02 U1773 ( .S(rptr[0]), .A0(ififoRdata[471]), .A1(ififoRdata[535]), .Z(n6634));
Q_MX02 U1774 ( .S(rptr[0]), .A0(ififoRdata[470]), .A1(ififoRdata[534]), .Z(n6633));
Q_MX02 U1775 ( .S(rptr[0]), .A0(ififoRdata[469]), .A1(ififoRdata[533]), .Z(n6632));
Q_MX02 U1776 ( .S(rptr[0]), .A0(ififoRdata[468]), .A1(ififoRdata[532]), .Z(n6631));
Q_MX02 U1777 ( .S(rptr[0]), .A0(ififoRdata[467]), .A1(ififoRdata[531]), .Z(n6630));
Q_MX02 U1778 ( .S(rptr[0]), .A0(ififoRdata[466]), .A1(ififoRdata[530]), .Z(n6629));
Q_MX02 U1779 ( .S(rptr[0]), .A0(ififoRdata[465]), .A1(ififoRdata[529]), .Z(n6628));
Q_MX02 U1780 ( .S(rptr[0]), .A0(ififoRdata[464]), .A1(ififoRdata[528]), .Z(n6627));
Q_MX02 U1781 ( .S(rptr[0]), .A0(ififoRdata[463]), .A1(ififoRdata[527]), .Z(n6626));
Q_MX02 U1782 ( .S(rptr[0]), .A0(ififoRdata[462]), .A1(ififoRdata[526]), .Z(n6625));
Q_MX02 U1783 ( .S(rptr[0]), .A0(ififoRdata[461]), .A1(ififoRdata[525]), .Z(n6624));
Q_MX02 U1784 ( .S(rptr[0]), .A0(ififoRdata[460]), .A1(ififoRdata[524]), .Z(n6623));
Q_MX02 U1785 ( .S(rptr[0]), .A0(ififoRdata[459]), .A1(ififoRdata[523]), .Z(n6622));
Q_MX02 U1786 ( .S(rptr[0]), .A0(ififoRdata[458]), .A1(ififoRdata[522]), .Z(n6621));
Q_MX02 U1787 ( .S(rptr[0]), .A0(ififoRdata[457]), .A1(ififoRdata[521]), .Z(n6620));
Q_MX02 U1788 ( .S(rptr[0]), .A0(ififoRdata[456]), .A1(ififoRdata[520]), .Z(n6619));
Q_MX02 U1789 ( .S(rptr[0]), .A0(ififoRdata[455]), .A1(ififoRdata[519]), .Z(n6618));
Q_MX02 U1790 ( .S(rptr[0]), .A0(ififoRdata[454]), .A1(ififoRdata[518]), .Z(n6617));
Q_MX02 U1791 ( .S(rptr[0]), .A0(ififoRdata[453]), .A1(ififoRdata[517]), .Z(n6616));
Q_MX02 U1792 ( .S(rptr[0]), .A0(ififoRdata[452]), .A1(ififoRdata[516]), .Z(n6615));
Q_MX02 U1793 ( .S(rptr[0]), .A0(ififoRdata[451]), .A1(ififoRdata[515]), .Z(n6614));
Q_MX02 U1794 ( .S(rptr[0]), .A0(ififoRdata[450]), .A1(ififoRdata[514]), .Z(n6613));
Q_MX02 U1795 ( .S(rptr[0]), .A0(ififoRdata[449]), .A1(ififoRdata[513]), .Z(n6612));
Q_MX02 U1796 ( .S(rptr[0]), .A0(ififoRdata[448]), .A1(ififoRdata[512]), .Z(n6611));
Q_MX02 U1797 ( .S(rptr[0]), .A0(ififoRdata[447]), .A1(ififoRdata[511]), .Z(n6610));
Q_MX02 U1798 ( .S(rptr[0]), .A0(ififoRdata[446]), .A1(ififoRdata[510]), .Z(n6609));
Q_MX02 U1799 ( .S(rptr[0]), .A0(ififoRdata[445]), .A1(ififoRdata[509]), .Z(n6608));
Q_MX02 U1800 ( .S(rptr[0]), .A0(ififoRdata[444]), .A1(ififoRdata[508]), .Z(n6607));
Q_MX02 U1801 ( .S(rptr[0]), .A0(ififoRdata[443]), .A1(ififoRdata[507]), .Z(n6606));
Q_MX02 U1802 ( .S(rptr[0]), .A0(ififoRdata[442]), .A1(ififoRdata[506]), .Z(n6605));
Q_MX02 U1803 ( .S(rptr[0]), .A0(ififoRdata[441]), .A1(ififoRdata[505]), .Z(n6604));
Q_MX02 U1804 ( .S(rptr[0]), .A0(ififoRdata[440]), .A1(ififoRdata[504]), .Z(n6603));
Q_MX02 U1805 ( .S(rptr[0]), .A0(ififoRdata[439]), .A1(ififoRdata[503]), .Z(n6602));
Q_MX02 U1806 ( .S(rptr[0]), .A0(ififoRdata[438]), .A1(ififoRdata[502]), .Z(n6601));
Q_MX02 U1807 ( .S(rptr[0]), .A0(ififoRdata[437]), .A1(ififoRdata[501]), .Z(n6600));
Q_MX02 U1808 ( .S(rptr[0]), .A0(ififoRdata[436]), .A1(ififoRdata[500]), .Z(n6599));
Q_MX02 U1809 ( .S(rptr[0]), .A0(ififoRdata[435]), .A1(ififoRdata[499]), .Z(n6598));
Q_MX02 U1810 ( .S(rptr[0]), .A0(ififoRdata[434]), .A1(ififoRdata[498]), .Z(n6597));
Q_MX02 U1811 ( .S(rptr[0]), .A0(ififoRdata[433]), .A1(ififoRdata[497]), .Z(n6596));
Q_MX02 U1812 ( .S(rptr[0]), .A0(ififoRdata[432]), .A1(ififoRdata[496]), .Z(n6595));
Q_MX02 U1813 ( .S(rptr[0]), .A0(ififoRdata[431]), .A1(ififoRdata[495]), .Z(n6594));
Q_MX02 U1814 ( .S(rptr[0]), .A0(ififoRdata[430]), .A1(ififoRdata[494]), .Z(n6593));
Q_MX02 U1815 ( .S(rptr[0]), .A0(ififoRdata[429]), .A1(ififoRdata[493]), .Z(n6592));
Q_MX02 U1816 ( .S(rptr[0]), .A0(ififoRdata[428]), .A1(ififoRdata[492]), .Z(n6591));
Q_MX02 U1817 ( .S(rptr[0]), .A0(ififoRdata[427]), .A1(ififoRdata[491]), .Z(n6590));
Q_MX02 U1818 ( .S(rptr[0]), .A0(ififoRdata[426]), .A1(ififoRdata[490]), .Z(n6589));
Q_MX02 U1819 ( .S(rptr[0]), .A0(ififoRdata[425]), .A1(ififoRdata[489]), .Z(n6588));
Q_MX02 U1820 ( .S(rptr[0]), .A0(ififoRdata[424]), .A1(ififoRdata[488]), .Z(n6587));
Q_MX02 U1821 ( .S(rptr[0]), .A0(ififoRdata[423]), .A1(ififoRdata[487]), .Z(n6586));
Q_MX02 U1822 ( .S(rptr[0]), .A0(ififoRdata[422]), .A1(ififoRdata[486]), .Z(n6585));
Q_MX02 U1823 ( .S(rptr[0]), .A0(ififoRdata[421]), .A1(ififoRdata[485]), .Z(n6584));
Q_MX02 U1824 ( .S(rptr[0]), .A0(ififoRdata[420]), .A1(ififoRdata[484]), .Z(n6583));
Q_MX02 U1825 ( .S(rptr[0]), .A0(ififoRdata[419]), .A1(ififoRdata[483]), .Z(n6582));
Q_MX02 U1826 ( .S(rptr[0]), .A0(ififoRdata[418]), .A1(ififoRdata[482]), .Z(n6581));
Q_MX02 U1827 ( .S(rptr[0]), .A0(ififoRdata[417]), .A1(ififoRdata[481]), .Z(n6580));
Q_MX02 U1828 ( .S(rptr[0]), .A0(ififoRdata[416]), .A1(ififoRdata[480]), .Z(n6579));
Q_MX02 U1829 ( .S(rptr[0]), .A0(ififoRdata[415]), .A1(ififoRdata[479]), .Z(n6578));
Q_MX02 U1830 ( .S(rptr[0]), .A0(ififoRdata[414]), .A1(ififoRdata[478]), .Z(n6577));
Q_MX02 U1831 ( .S(rptr[0]), .A0(ififoRdata[413]), .A1(ififoRdata[477]), .Z(n6576));
Q_MX02 U1832 ( .S(rptr[0]), .A0(ififoRdata[412]), .A1(ififoRdata[476]), .Z(n6575));
Q_MX02 U1833 ( .S(rptr[0]), .A0(ififoRdata[411]), .A1(ififoRdata[475]), .Z(n6574));
Q_MX02 U1834 ( .S(rptr[0]), .A0(ififoRdata[410]), .A1(ififoRdata[474]), .Z(n6573));
Q_MX02 U1835 ( .S(rptr[0]), .A0(ififoRdata[409]), .A1(ififoRdata[473]), .Z(n6572));
Q_MX02 U1836 ( .S(rptr[0]), .A0(ififoRdata[408]), .A1(ififoRdata[472]), .Z(n6571));
Q_MX02 U1837 ( .S(rptr[0]), .A0(ififoRdata[407]), .A1(ififoRdata[471]), .Z(n6570));
Q_MX02 U1838 ( .S(rptr[0]), .A0(ififoRdata[406]), .A1(ififoRdata[470]), .Z(n6569));
Q_MX02 U1839 ( .S(rptr[0]), .A0(ififoRdata[405]), .A1(ififoRdata[469]), .Z(n6568));
Q_MX02 U1840 ( .S(rptr[0]), .A0(ififoRdata[404]), .A1(ififoRdata[468]), .Z(n6567));
Q_MX02 U1841 ( .S(rptr[0]), .A0(ififoRdata[403]), .A1(ififoRdata[467]), .Z(n6566));
Q_MX02 U1842 ( .S(rptr[0]), .A0(ififoRdata[402]), .A1(ififoRdata[466]), .Z(n6565));
Q_MX02 U1843 ( .S(rptr[0]), .A0(ififoRdata[401]), .A1(ififoRdata[465]), .Z(n6564));
Q_MX02 U1844 ( .S(rptr[0]), .A0(ififoRdata[400]), .A1(ififoRdata[464]), .Z(n6563));
Q_MX02 U1845 ( .S(rptr[0]), .A0(ififoRdata[399]), .A1(ififoRdata[463]), .Z(n6562));
Q_MX02 U1846 ( .S(rptr[0]), .A0(ififoRdata[398]), .A1(ififoRdata[462]), .Z(n6561));
Q_MX02 U1847 ( .S(rptr[0]), .A0(ififoRdata[397]), .A1(ififoRdata[461]), .Z(n6560));
Q_MX02 U1848 ( .S(rptr[0]), .A0(ififoRdata[396]), .A1(ififoRdata[460]), .Z(n6559));
Q_MX02 U1849 ( .S(rptr[0]), .A0(ififoRdata[395]), .A1(ififoRdata[459]), .Z(n6558));
Q_MX02 U1850 ( .S(rptr[0]), .A0(ififoRdata[394]), .A1(ififoRdata[458]), .Z(n6557));
Q_MX02 U1851 ( .S(rptr[0]), .A0(ififoRdata[393]), .A1(ififoRdata[457]), .Z(n6556));
Q_MX02 U1852 ( .S(rptr[0]), .A0(ififoRdata[392]), .A1(ififoRdata[456]), .Z(n6555));
Q_MX02 U1853 ( .S(rptr[0]), .A0(ififoRdata[391]), .A1(ififoRdata[455]), .Z(n6554));
Q_MX02 U1854 ( .S(rptr[0]), .A0(ififoRdata[390]), .A1(ififoRdata[454]), .Z(n6553));
Q_MX02 U1855 ( .S(rptr[0]), .A0(ififoRdata[389]), .A1(ififoRdata[453]), .Z(n6552));
Q_MX02 U1856 ( .S(rptr[0]), .A0(ififoRdata[388]), .A1(ififoRdata[452]), .Z(n6551));
Q_MX02 U1857 ( .S(rptr[0]), .A0(ififoRdata[387]), .A1(ififoRdata[451]), .Z(n6550));
Q_MX02 U1858 ( .S(rptr[0]), .A0(ififoRdata[386]), .A1(ififoRdata[450]), .Z(n6549));
Q_MX02 U1859 ( .S(rptr[0]), .A0(ififoRdata[385]), .A1(ififoRdata[449]), .Z(n6548));
Q_MX02 U1860 ( .S(rptr[0]), .A0(ififoRdata[384]), .A1(ififoRdata[448]), .Z(n6547));
Q_MX02 U1861 ( .S(rptr[0]), .A0(ififoRdata[383]), .A1(ififoRdata[447]), .Z(n6546));
Q_MX02 U1862 ( .S(rptr[0]), .A0(ififoRdata[382]), .A1(ififoRdata[446]), .Z(n6545));
Q_MX02 U1863 ( .S(rptr[0]), .A0(ififoRdata[381]), .A1(ififoRdata[445]), .Z(n6544));
Q_MX02 U1864 ( .S(rptr[0]), .A0(ififoRdata[380]), .A1(ififoRdata[444]), .Z(n6543));
Q_MX02 U1865 ( .S(rptr[0]), .A0(ififoRdata[379]), .A1(ififoRdata[443]), .Z(n6542));
Q_MX02 U1866 ( .S(rptr[0]), .A0(ififoRdata[378]), .A1(ififoRdata[442]), .Z(n6541));
Q_MX02 U1867 ( .S(rptr[0]), .A0(ififoRdata[377]), .A1(ififoRdata[441]), .Z(n6540));
Q_MX02 U1868 ( .S(rptr[0]), .A0(ififoRdata[376]), .A1(ififoRdata[440]), .Z(n6539));
Q_MX02 U1869 ( .S(rptr[0]), .A0(ififoRdata[375]), .A1(ififoRdata[439]), .Z(n6538));
Q_MX02 U1870 ( .S(rptr[0]), .A0(ififoRdata[374]), .A1(ififoRdata[438]), .Z(n6537));
Q_MX02 U1871 ( .S(rptr[0]), .A0(ififoRdata[373]), .A1(ififoRdata[437]), .Z(n6536));
Q_MX02 U1872 ( .S(rptr[0]), .A0(ififoRdata[372]), .A1(ififoRdata[436]), .Z(n6535));
Q_MX02 U1873 ( .S(rptr[0]), .A0(ififoRdata[371]), .A1(ififoRdata[435]), .Z(n6534));
Q_MX02 U1874 ( .S(rptr[0]), .A0(ififoRdata[370]), .A1(ififoRdata[434]), .Z(n6533));
Q_MX02 U1875 ( .S(rptr[0]), .A0(ififoRdata[369]), .A1(ififoRdata[433]), .Z(n6532));
Q_MX02 U1876 ( .S(rptr[0]), .A0(ififoRdata[368]), .A1(ififoRdata[432]), .Z(n6531));
Q_MX02 U1877 ( .S(rptr[0]), .A0(ififoRdata[367]), .A1(ififoRdata[431]), .Z(n6530));
Q_MX02 U1878 ( .S(rptr[0]), .A0(ififoRdata[366]), .A1(ififoRdata[430]), .Z(n6529));
Q_MX02 U1879 ( .S(rptr[0]), .A0(ififoRdata[365]), .A1(ififoRdata[429]), .Z(n6528));
Q_MX02 U1880 ( .S(rptr[0]), .A0(ififoRdata[364]), .A1(ififoRdata[428]), .Z(n6527));
Q_MX02 U1881 ( .S(rptr[0]), .A0(ififoRdata[363]), .A1(ififoRdata[427]), .Z(n6526));
Q_MX02 U1882 ( .S(rptr[0]), .A0(ififoRdata[362]), .A1(ififoRdata[426]), .Z(n6525));
Q_MX02 U1883 ( .S(rptr[0]), .A0(ififoRdata[361]), .A1(ififoRdata[425]), .Z(n6524));
Q_MX02 U1884 ( .S(rptr[0]), .A0(ififoRdata[360]), .A1(ififoRdata[424]), .Z(n6523));
Q_MX02 U1885 ( .S(rptr[0]), .A0(ififoRdata[359]), .A1(ififoRdata[423]), .Z(n6522));
Q_MX02 U1886 ( .S(rptr[0]), .A0(ififoRdata[358]), .A1(ififoRdata[422]), .Z(n6521));
Q_MX02 U1887 ( .S(rptr[0]), .A0(ififoRdata[357]), .A1(ififoRdata[421]), .Z(n6520));
Q_MX02 U1888 ( .S(rptr[0]), .A0(ififoRdata[356]), .A1(ififoRdata[420]), .Z(n6519));
Q_MX02 U1889 ( .S(rptr[0]), .A0(ififoRdata[355]), .A1(ififoRdata[419]), .Z(n6518));
Q_MX02 U1890 ( .S(rptr[0]), .A0(ififoRdata[354]), .A1(ififoRdata[418]), .Z(n6517));
Q_MX02 U1891 ( .S(rptr[0]), .A0(ififoRdata[353]), .A1(ififoRdata[417]), .Z(n6516));
Q_MX02 U1892 ( .S(rptr[0]), .A0(ififoRdata[352]), .A1(ififoRdata[416]), .Z(n6515));
Q_MX02 U1893 ( .S(rptr[0]), .A0(ififoRdata[351]), .A1(ififoRdata[415]), .Z(n6514));
Q_MX02 U1894 ( .S(rptr[0]), .A0(ififoRdata[350]), .A1(ififoRdata[414]), .Z(n6513));
Q_MX02 U1895 ( .S(rptr[0]), .A0(ififoRdata[349]), .A1(ififoRdata[413]), .Z(n6512));
Q_MX02 U1896 ( .S(rptr[0]), .A0(ififoRdata[348]), .A1(ififoRdata[412]), .Z(n6511));
Q_MX02 U1897 ( .S(rptr[0]), .A0(ififoRdata[347]), .A1(ififoRdata[411]), .Z(n6510));
Q_MX02 U1898 ( .S(rptr[0]), .A0(ififoRdata[346]), .A1(ififoRdata[410]), .Z(n6509));
Q_MX02 U1899 ( .S(rptr[0]), .A0(ififoRdata[345]), .A1(ififoRdata[409]), .Z(n6508));
Q_MX02 U1900 ( .S(rptr[0]), .A0(ififoRdata[344]), .A1(ififoRdata[408]), .Z(n6507));
Q_MX02 U1901 ( .S(rptr[0]), .A0(ififoRdata[343]), .A1(ififoRdata[407]), .Z(n6506));
Q_MX02 U1902 ( .S(rptr[0]), .A0(ififoRdata[342]), .A1(ififoRdata[406]), .Z(n6505));
Q_MX02 U1903 ( .S(rptr[0]), .A0(ififoRdata[341]), .A1(ififoRdata[405]), .Z(n6504));
Q_MX02 U1904 ( .S(rptr[0]), .A0(ififoRdata[340]), .A1(ififoRdata[404]), .Z(n6503));
Q_MX02 U1905 ( .S(rptr[0]), .A0(ififoRdata[339]), .A1(ififoRdata[403]), .Z(n6502));
Q_MX02 U1906 ( .S(rptr[0]), .A0(ififoRdata[338]), .A1(ififoRdata[402]), .Z(n6501));
Q_MX02 U1907 ( .S(rptr[0]), .A0(ififoRdata[337]), .A1(ififoRdata[401]), .Z(n6500));
Q_MX02 U1908 ( .S(rptr[0]), .A0(ififoRdata[336]), .A1(ififoRdata[400]), .Z(n6499));
Q_MX02 U1909 ( .S(rptr[0]), .A0(ififoRdata[335]), .A1(ififoRdata[399]), .Z(n6498));
Q_MX02 U1910 ( .S(rptr[0]), .A0(ififoRdata[334]), .A1(ififoRdata[398]), .Z(n6497));
Q_MX02 U1911 ( .S(rptr[0]), .A0(ififoRdata[333]), .A1(ififoRdata[397]), .Z(n6496));
Q_MX02 U1912 ( .S(rptr[0]), .A0(ififoRdata[332]), .A1(ififoRdata[396]), .Z(n6495));
Q_MX02 U1913 ( .S(rptr[0]), .A0(ififoRdata[331]), .A1(ififoRdata[395]), .Z(n6494));
Q_MX02 U1914 ( .S(rptr[0]), .A0(ififoRdata[330]), .A1(ififoRdata[394]), .Z(n6493));
Q_MX02 U1915 ( .S(rptr[0]), .A0(ififoRdata[329]), .A1(ififoRdata[393]), .Z(n6492));
Q_MX02 U1916 ( .S(rptr[0]), .A0(ififoRdata[328]), .A1(ififoRdata[392]), .Z(n6491));
Q_MX02 U1917 ( .S(rptr[0]), .A0(ififoRdata[327]), .A1(ififoRdata[391]), .Z(n6490));
Q_MX02 U1918 ( .S(rptr[0]), .A0(ififoRdata[326]), .A1(ififoRdata[390]), .Z(n6489));
Q_MX02 U1919 ( .S(rptr[0]), .A0(ififoRdata[325]), .A1(ififoRdata[389]), .Z(n6488));
Q_MX02 U1920 ( .S(rptr[0]), .A0(ififoRdata[324]), .A1(ififoRdata[388]), .Z(n6487));
Q_MX02 U1921 ( .S(rptr[0]), .A0(ififoRdata[323]), .A1(ififoRdata[387]), .Z(n6486));
Q_MX02 U1922 ( .S(rptr[0]), .A0(ififoRdata[322]), .A1(ififoRdata[386]), .Z(n6485));
Q_MX02 U1923 ( .S(rptr[0]), .A0(ififoRdata[321]), .A1(ififoRdata[385]), .Z(n6484));
Q_MX02 U1924 ( .S(rptr[0]), .A0(ififoRdata[320]), .A1(ififoRdata[384]), .Z(n6483));
Q_MX02 U1925 ( .S(rptr[0]), .A0(ififoRdata[319]), .A1(ififoRdata[383]), .Z(n6482));
Q_MX02 U1926 ( .S(rptr[0]), .A0(ififoRdata[318]), .A1(ififoRdata[382]), .Z(n6481));
Q_MX02 U1927 ( .S(rptr[0]), .A0(ififoRdata[317]), .A1(ififoRdata[381]), .Z(n6480));
Q_MX02 U1928 ( .S(rptr[0]), .A0(ififoRdata[316]), .A1(ififoRdata[380]), .Z(n6479));
Q_MX02 U1929 ( .S(rptr[0]), .A0(ififoRdata[315]), .A1(ififoRdata[379]), .Z(n6478));
Q_MX02 U1930 ( .S(rptr[0]), .A0(ififoRdata[314]), .A1(ififoRdata[378]), .Z(n6477));
Q_MX02 U1931 ( .S(rptr[0]), .A0(ififoRdata[313]), .A1(ififoRdata[377]), .Z(n6476));
Q_MX02 U1932 ( .S(rptr[0]), .A0(ififoRdata[312]), .A1(ififoRdata[376]), .Z(n6475));
Q_MX02 U1933 ( .S(rptr[0]), .A0(ififoRdata[311]), .A1(ififoRdata[375]), .Z(n6474));
Q_MX02 U1934 ( .S(rptr[0]), .A0(ififoRdata[310]), .A1(ififoRdata[374]), .Z(n6473));
Q_MX02 U1935 ( .S(rptr[0]), .A0(ififoRdata[309]), .A1(ififoRdata[373]), .Z(n6472));
Q_MX02 U1936 ( .S(rptr[0]), .A0(ififoRdata[308]), .A1(ififoRdata[372]), .Z(n6471));
Q_MX02 U1937 ( .S(rptr[0]), .A0(ififoRdata[307]), .A1(ififoRdata[371]), .Z(n6470));
Q_MX02 U1938 ( .S(rptr[0]), .A0(ififoRdata[306]), .A1(ififoRdata[370]), .Z(n6469));
Q_MX02 U1939 ( .S(rptr[0]), .A0(ififoRdata[305]), .A1(ififoRdata[369]), .Z(n6468));
Q_MX02 U1940 ( .S(rptr[0]), .A0(ififoRdata[304]), .A1(ififoRdata[368]), .Z(n6467));
Q_MX02 U1941 ( .S(rptr[0]), .A0(ififoRdata[303]), .A1(ififoRdata[367]), .Z(n6466));
Q_MX02 U1942 ( .S(rptr[0]), .A0(ififoRdata[302]), .A1(ififoRdata[366]), .Z(n6465));
Q_MX02 U1943 ( .S(rptr[0]), .A0(ififoRdata[301]), .A1(ififoRdata[365]), .Z(n6464));
Q_MX02 U1944 ( .S(rptr[0]), .A0(ififoRdata[300]), .A1(ififoRdata[364]), .Z(n6463));
Q_MX02 U1945 ( .S(rptr[0]), .A0(ififoRdata[299]), .A1(ififoRdata[363]), .Z(n6462));
Q_MX02 U1946 ( .S(rptr[0]), .A0(ififoRdata[298]), .A1(ififoRdata[362]), .Z(n6461));
Q_MX02 U1947 ( .S(rptr[0]), .A0(ififoRdata[297]), .A1(ififoRdata[361]), .Z(n6460));
Q_MX02 U1948 ( .S(rptr[0]), .A0(ififoRdata[296]), .A1(ififoRdata[360]), .Z(n6459));
Q_MX02 U1949 ( .S(rptr[0]), .A0(ififoRdata[295]), .A1(ififoRdata[359]), .Z(n6458));
Q_MX02 U1950 ( .S(rptr[0]), .A0(ififoRdata[294]), .A1(ififoRdata[358]), .Z(n6457));
Q_MX02 U1951 ( .S(rptr[0]), .A0(ififoRdata[293]), .A1(ififoRdata[357]), .Z(n6456));
Q_MX02 U1952 ( .S(rptr[0]), .A0(ififoRdata[292]), .A1(ififoRdata[356]), .Z(n6455));
Q_MX02 U1953 ( .S(rptr[0]), .A0(ififoRdata[291]), .A1(ififoRdata[355]), .Z(n6454));
Q_MX02 U1954 ( .S(rptr[0]), .A0(ififoRdata[290]), .A1(ififoRdata[354]), .Z(n6453));
Q_MX02 U1955 ( .S(rptr[0]), .A0(ififoRdata[289]), .A1(ififoRdata[353]), .Z(n6452));
Q_MX02 U1956 ( .S(rptr[0]), .A0(ififoRdata[288]), .A1(ififoRdata[352]), .Z(n6451));
Q_MX02 U1957 ( .S(rptr[0]), .A0(ififoRdata[287]), .A1(ififoRdata[351]), .Z(n6450));
Q_MX02 U1958 ( .S(rptr[0]), .A0(ififoRdata[286]), .A1(ififoRdata[350]), .Z(n6449));
Q_MX02 U1959 ( .S(rptr[0]), .A0(ififoRdata[285]), .A1(ififoRdata[349]), .Z(n6448));
Q_MX02 U1960 ( .S(rptr[0]), .A0(ififoRdata[284]), .A1(ififoRdata[348]), .Z(n6447));
Q_MX02 U1961 ( .S(rptr[0]), .A0(ififoRdata[283]), .A1(ififoRdata[347]), .Z(n6446));
Q_MX02 U1962 ( .S(rptr[0]), .A0(ififoRdata[282]), .A1(ififoRdata[346]), .Z(n6445));
Q_MX02 U1963 ( .S(rptr[0]), .A0(ififoRdata[281]), .A1(ififoRdata[345]), .Z(n6444));
Q_MX02 U1964 ( .S(rptr[0]), .A0(ififoRdata[280]), .A1(ififoRdata[344]), .Z(n6443));
Q_MX02 U1965 ( .S(rptr[0]), .A0(ififoRdata[279]), .A1(ififoRdata[343]), .Z(n6442));
Q_MX02 U1966 ( .S(rptr[0]), .A0(ififoRdata[278]), .A1(ififoRdata[342]), .Z(n6441));
Q_MX02 U1967 ( .S(rptr[0]), .A0(ififoRdata[277]), .A1(ififoRdata[341]), .Z(n6440));
Q_MX02 U1968 ( .S(rptr[0]), .A0(ififoRdata[276]), .A1(ififoRdata[340]), .Z(n6439));
Q_MX02 U1969 ( .S(rptr[0]), .A0(ififoRdata[275]), .A1(ififoRdata[339]), .Z(n6438));
Q_MX02 U1970 ( .S(rptr[0]), .A0(ififoRdata[274]), .A1(ififoRdata[338]), .Z(n6437));
Q_MX02 U1971 ( .S(rptr[0]), .A0(ififoRdata[273]), .A1(ififoRdata[337]), .Z(n6436));
Q_MX02 U1972 ( .S(rptr[0]), .A0(ififoRdata[272]), .A1(ififoRdata[336]), .Z(n6435));
Q_MX02 U1973 ( .S(rptr[0]), .A0(ififoRdata[271]), .A1(ififoRdata[335]), .Z(n6434));
Q_MX02 U1974 ( .S(rptr[0]), .A0(ififoRdata[270]), .A1(ififoRdata[334]), .Z(n6433));
Q_MX02 U1975 ( .S(rptr[0]), .A0(ififoRdata[269]), .A1(ififoRdata[333]), .Z(n6432));
Q_MX02 U1976 ( .S(rptr[0]), .A0(ififoRdata[268]), .A1(ififoRdata[332]), .Z(n6431));
Q_MX02 U1977 ( .S(rptr[0]), .A0(ififoRdata[267]), .A1(ififoRdata[331]), .Z(n6430));
Q_MX02 U1978 ( .S(rptr[0]), .A0(ififoRdata[266]), .A1(ififoRdata[330]), .Z(n6429));
Q_MX02 U1979 ( .S(rptr[0]), .A0(ififoRdata[265]), .A1(ififoRdata[329]), .Z(n6428));
Q_MX02 U1980 ( .S(rptr[0]), .A0(ififoRdata[264]), .A1(ififoRdata[328]), .Z(n6427));
Q_MX02 U1981 ( .S(rptr[0]), .A0(ififoRdata[263]), .A1(ififoRdata[327]), .Z(n6426));
Q_MX02 U1982 ( .S(rptr[0]), .A0(ififoRdata[262]), .A1(ififoRdata[326]), .Z(n6425));
Q_MX02 U1983 ( .S(rptr[0]), .A0(ififoRdata[261]), .A1(ififoRdata[325]), .Z(n6424));
Q_MX02 U1984 ( .S(rptr[0]), .A0(ififoRdata[260]), .A1(ififoRdata[324]), .Z(n6423));
Q_MX02 U1985 ( .S(rptr[0]), .A0(ififoRdata[259]), .A1(ififoRdata[323]), .Z(n6422));
Q_MX02 U1986 ( .S(rptr[0]), .A0(ififoRdata[258]), .A1(ififoRdata[322]), .Z(n6421));
Q_MX02 U1987 ( .S(rptr[0]), .A0(ififoRdata[257]), .A1(ififoRdata[321]), .Z(n6420));
Q_MX02 U1988 ( .S(rptr[0]), .A0(ififoRdata[256]), .A1(ififoRdata[320]), .Z(n6419));
Q_MX02 U1989 ( .S(rptr[0]), .A0(ififoRdata[255]), .A1(ififoRdata[319]), .Z(n6418));
Q_MX02 U1990 ( .S(rptr[0]), .A0(ififoRdata[254]), .A1(ififoRdata[318]), .Z(n6417));
Q_MX02 U1991 ( .S(rptr[0]), .A0(ififoRdata[253]), .A1(ififoRdata[317]), .Z(n6416));
Q_MX02 U1992 ( .S(rptr[0]), .A0(ififoRdata[252]), .A1(ififoRdata[316]), .Z(n6415));
Q_MX02 U1993 ( .S(rptr[0]), .A0(ififoRdata[251]), .A1(ififoRdata[315]), .Z(n6414));
Q_MX02 U1994 ( .S(rptr[0]), .A0(ififoRdata[250]), .A1(ififoRdata[314]), .Z(n6413));
Q_MX02 U1995 ( .S(rptr[0]), .A0(ififoRdata[249]), .A1(ififoRdata[313]), .Z(n6412));
Q_MX02 U1996 ( .S(rptr[0]), .A0(ififoRdata[248]), .A1(ififoRdata[312]), .Z(n6411));
Q_MX02 U1997 ( .S(rptr[0]), .A0(ififoRdata[247]), .A1(ififoRdata[311]), .Z(n6410));
Q_MX02 U1998 ( .S(rptr[0]), .A0(ififoRdata[246]), .A1(ififoRdata[310]), .Z(n6409));
Q_MX02 U1999 ( .S(rptr[0]), .A0(ififoRdata[245]), .A1(ififoRdata[309]), .Z(n6408));
Q_MX02 U2000 ( .S(rptr[0]), .A0(ififoRdata[244]), .A1(ififoRdata[308]), .Z(n6407));
Q_MX02 U2001 ( .S(rptr[0]), .A0(ififoRdata[243]), .A1(ififoRdata[307]), .Z(n6406));
Q_MX02 U2002 ( .S(rptr[0]), .A0(ififoRdata[242]), .A1(ififoRdata[306]), .Z(n6405));
Q_MX02 U2003 ( .S(rptr[0]), .A0(ififoRdata[241]), .A1(ififoRdata[305]), .Z(n6404));
Q_MX02 U2004 ( .S(rptr[0]), .A0(ififoRdata[240]), .A1(ififoRdata[304]), .Z(n6403));
Q_MX02 U2005 ( .S(rptr[0]), .A0(ififoRdata[239]), .A1(ififoRdata[303]), .Z(n6402));
Q_MX02 U2006 ( .S(rptr[0]), .A0(ififoRdata[238]), .A1(ififoRdata[302]), .Z(n6401));
Q_MX02 U2007 ( .S(rptr[0]), .A0(ififoRdata[237]), .A1(ififoRdata[301]), .Z(n6400));
Q_MX02 U2008 ( .S(rptr[0]), .A0(ififoRdata[236]), .A1(ififoRdata[300]), .Z(n6399));
Q_MX02 U2009 ( .S(rptr[0]), .A0(ififoRdata[235]), .A1(ififoRdata[299]), .Z(n6398));
Q_MX02 U2010 ( .S(rptr[0]), .A0(ififoRdata[234]), .A1(ififoRdata[298]), .Z(n6397));
Q_MX02 U2011 ( .S(rptr[0]), .A0(ififoRdata[233]), .A1(ififoRdata[297]), .Z(n6396));
Q_MX02 U2012 ( .S(rptr[0]), .A0(ififoRdata[232]), .A1(ififoRdata[296]), .Z(n6395));
Q_MX02 U2013 ( .S(rptr[0]), .A0(ififoRdata[231]), .A1(ififoRdata[295]), .Z(n6394));
Q_MX02 U2014 ( .S(rptr[0]), .A0(ififoRdata[230]), .A1(ififoRdata[294]), .Z(n6393));
Q_MX02 U2015 ( .S(rptr[0]), .A0(ififoRdata[229]), .A1(ififoRdata[293]), .Z(n6392));
Q_MX02 U2016 ( .S(rptr[0]), .A0(ififoRdata[228]), .A1(ififoRdata[292]), .Z(n6391));
Q_MX02 U2017 ( .S(rptr[0]), .A0(ififoRdata[227]), .A1(ififoRdata[291]), .Z(n6390));
Q_MX02 U2018 ( .S(rptr[0]), .A0(ififoRdata[226]), .A1(ififoRdata[290]), .Z(n6389));
Q_MX02 U2019 ( .S(rptr[0]), .A0(ififoRdata[225]), .A1(ififoRdata[289]), .Z(n6388));
Q_MX02 U2020 ( .S(rptr[0]), .A0(ififoRdata[224]), .A1(ififoRdata[288]), .Z(n6387));
Q_MX02 U2021 ( .S(rptr[0]), .A0(ififoRdata[223]), .A1(ififoRdata[287]), .Z(n6386));
Q_MX02 U2022 ( .S(rptr[0]), .A0(ififoRdata[222]), .A1(ififoRdata[286]), .Z(n6385));
Q_MX02 U2023 ( .S(rptr[0]), .A0(ififoRdata[221]), .A1(ififoRdata[285]), .Z(n6384));
Q_MX02 U2024 ( .S(rptr[0]), .A0(ififoRdata[220]), .A1(ififoRdata[284]), .Z(n6383));
Q_MX02 U2025 ( .S(rptr[0]), .A0(ififoRdata[219]), .A1(ififoRdata[283]), .Z(n6382));
Q_MX02 U2026 ( .S(rptr[0]), .A0(ififoRdata[218]), .A1(ififoRdata[282]), .Z(n6381));
Q_MX02 U2027 ( .S(rptr[0]), .A0(ififoRdata[217]), .A1(ififoRdata[281]), .Z(n6380));
Q_MX02 U2028 ( .S(rptr[0]), .A0(ififoRdata[216]), .A1(ififoRdata[280]), .Z(n6379));
Q_MX02 U2029 ( .S(rptr[0]), .A0(ififoRdata[215]), .A1(ififoRdata[279]), .Z(n6378));
Q_MX02 U2030 ( .S(rptr[0]), .A0(ififoRdata[214]), .A1(ififoRdata[278]), .Z(n6377));
Q_MX02 U2031 ( .S(rptr[0]), .A0(ififoRdata[213]), .A1(ififoRdata[277]), .Z(n6376));
Q_MX02 U2032 ( .S(rptr[0]), .A0(ififoRdata[212]), .A1(ififoRdata[276]), .Z(n6375));
Q_MX02 U2033 ( .S(rptr[0]), .A0(ififoRdata[211]), .A1(ififoRdata[275]), .Z(n6374));
Q_MX02 U2034 ( .S(rptr[0]), .A0(ififoRdata[210]), .A1(ififoRdata[274]), .Z(n6373));
Q_MX02 U2035 ( .S(rptr[0]), .A0(ififoRdata[209]), .A1(ififoRdata[273]), .Z(n6372));
Q_MX02 U2036 ( .S(rptr[0]), .A0(ififoRdata[208]), .A1(ififoRdata[272]), .Z(n6371));
Q_MX02 U2037 ( .S(rptr[0]), .A0(ififoRdata[207]), .A1(ififoRdata[271]), .Z(n6370));
Q_MX02 U2038 ( .S(rptr[0]), .A0(ififoRdata[206]), .A1(ififoRdata[270]), .Z(n6369));
Q_MX02 U2039 ( .S(rptr[0]), .A0(ififoRdata[205]), .A1(ififoRdata[269]), .Z(n6368));
Q_MX02 U2040 ( .S(rptr[0]), .A0(ififoRdata[204]), .A1(ififoRdata[268]), .Z(n6367));
Q_MX02 U2041 ( .S(rptr[0]), .A0(ififoRdata[203]), .A1(ififoRdata[267]), .Z(n6366));
Q_MX02 U2042 ( .S(rptr[0]), .A0(ififoRdata[202]), .A1(ififoRdata[266]), .Z(n6365));
Q_MX02 U2043 ( .S(rptr[0]), .A0(ififoRdata[201]), .A1(ififoRdata[265]), .Z(n6364));
Q_MX02 U2044 ( .S(rptr[0]), .A0(ififoRdata[200]), .A1(ififoRdata[264]), .Z(n6363));
Q_MX02 U2045 ( .S(rptr[0]), .A0(ififoRdata[199]), .A1(ififoRdata[263]), .Z(n6362));
Q_MX02 U2046 ( .S(rptr[0]), .A0(ififoRdata[198]), .A1(ififoRdata[262]), .Z(n6361));
Q_MX02 U2047 ( .S(rptr[0]), .A0(ififoRdata[197]), .A1(ififoRdata[261]), .Z(n6360));
Q_MX02 U2048 ( .S(rptr[0]), .A0(ififoRdata[196]), .A1(ififoRdata[260]), .Z(n6359));
Q_MX02 U2049 ( .S(rptr[0]), .A0(ififoRdata[195]), .A1(ififoRdata[259]), .Z(n6358));
Q_MX02 U2050 ( .S(rptr[0]), .A0(ififoRdata[194]), .A1(ififoRdata[258]), .Z(n6357));
Q_MX02 U2051 ( .S(rptr[0]), .A0(ififoRdata[193]), .A1(ififoRdata[257]), .Z(n6356));
Q_MX02 U2052 ( .S(rptr[0]), .A0(ififoRdata[192]), .A1(ififoRdata[256]), .Z(n6355));
Q_MX02 U2053 ( .S(rptr[0]), .A0(ififoRdata[191]), .A1(ififoRdata[255]), .Z(n6354));
Q_MX02 U2054 ( .S(rptr[0]), .A0(ififoRdata[190]), .A1(ififoRdata[254]), .Z(n6353));
Q_MX02 U2055 ( .S(rptr[0]), .A0(ififoRdata[189]), .A1(ififoRdata[253]), .Z(n6352));
Q_MX02 U2056 ( .S(rptr[0]), .A0(ififoRdata[188]), .A1(ififoRdata[252]), .Z(n6351));
Q_MX02 U2057 ( .S(rptr[0]), .A0(ififoRdata[187]), .A1(ififoRdata[251]), .Z(n6350));
Q_MX02 U2058 ( .S(rptr[0]), .A0(ififoRdata[186]), .A1(ififoRdata[250]), .Z(n6349));
Q_MX02 U2059 ( .S(rptr[0]), .A0(ififoRdata[185]), .A1(ififoRdata[249]), .Z(n6348));
Q_MX02 U2060 ( .S(rptr[0]), .A0(ififoRdata[184]), .A1(ififoRdata[248]), .Z(n6347));
Q_MX02 U2061 ( .S(rptr[0]), .A0(ififoRdata[183]), .A1(ififoRdata[247]), .Z(n6346));
Q_MX02 U2062 ( .S(rptr[0]), .A0(ififoRdata[182]), .A1(ififoRdata[246]), .Z(n6345));
Q_MX02 U2063 ( .S(rptr[0]), .A0(ififoRdata[181]), .A1(ififoRdata[245]), .Z(n6344));
Q_MX02 U2064 ( .S(rptr[0]), .A0(ififoRdata[180]), .A1(ififoRdata[244]), .Z(n6343));
Q_MX02 U2065 ( .S(rptr[0]), .A0(ififoRdata[179]), .A1(ififoRdata[243]), .Z(n6342));
Q_MX02 U2066 ( .S(rptr[0]), .A0(ififoRdata[178]), .A1(ififoRdata[242]), .Z(n6341));
Q_MX02 U2067 ( .S(rptr[0]), .A0(ififoRdata[177]), .A1(ififoRdata[241]), .Z(n6340));
Q_MX02 U2068 ( .S(rptr[0]), .A0(ififoRdata[176]), .A1(ififoRdata[240]), .Z(n6339));
Q_MX02 U2069 ( .S(rptr[0]), .A0(ififoRdata[175]), .A1(ififoRdata[239]), .Z(n6338));
Q_MX02 U2070 ( .S(rptr[0]), .A0(ififoRdata[174]), .A1(ififoRdata[238]), .Z(n6337));
Q_MX02 U2071 ( .S(rptr[0]), .A0(ififoRdata[173]), .A1(ififoRdata[237]), .Z(n6336));
Q_MX02 U2072 ( .S(rptr[0]), .A0(ififoRdata[172]), .A1(ififoRdata[236]), .Z(n6335));
Q_MX02 U2073 ( .S(rptr[0]), .A0(ififoRdata[171]), .A1(ififoRdata[235]), .Z(n6334));
Q_MX02 U2074 ( .S(rptr[0]), .A0(ififoRdata[170]), .A1(ififoRdata[234]), .Z(n6333));
Q_MX02 U2075 ( .S(rptr[0]), .A0(ififoRdata[169]), .A1(ififoRdata[233]), .Z(n6332));
Q_MX02 U2076 ( .S(rptr[0]), .A0(ififoRdata[168]), .A1(ififoRdata[232]), .Z(n6331));
Q_MX02 U2077 ( .S(rptr[0]), .A0(ififoRdata[167]), .A1(ififoRdata[231]), .Z(n6330));
Q_MX02 U2078 ( .S(rptr[0]), .A0(ififoRdata[166]), .A1(ififoRdata[230]), .Z(n6329));
Q_MX02 U2079 ( .S(rptr[0]), .A0(ififoRdata[165]), .A1(ififoRdata[229]), .Z(n6328));
Q_MX02 U2080 ( .S(rptr[0]), .A0(ififoRdata[164]), .A1(ififoRdata[228]), .Z(n6327));
Q_MX02 U2081 ( .S(rptr[0]), .A0(ififoRdata[163]), .A1(ififoRdata[227]), .Z(n6326));
Q_MX02 U2082 ( .S(rptr[0]), .A0(ififoRdata[162]), .A1(ififoRdata[226]), .Z(n6325));
Q_MX02 U2083 ( .S(rptr[0]), .A0(ififoRdata[161]), .A1(ififoRdata[225]), .Z(n6324));
Q_MX02 U2084 ( .S(rptr[0]), .A0(ififoRdata[160]), .A1(ififoRdata[224]), .Z(n6323));
Q_MX02 U2085 ( .S(rptr[0]), .A0(ififoRdata[159]), .A1(ififoRdata[223]), .Z(n6322));
Q_MX02 U2086 ( .S(rptr[0]), .A0(ififoRdata[158]), .A1(ififoRdata[222]), .Z(n6321));
Q_MX02 U2087 ( .S(rptr[0]), .A0(ififoRdata[157]), .A1(ififoRdata[221]), .Z(n6320));
Q_MX02 U2088 ( .S(rptr[0]), .A0(ififoRdata[156]), .A1(ififoRdata[220]), .Z(n6319));
Q_MX02 U2089 ( .S(rptr[0]), .A0(ififoRdata[155]), .A1(ififoRdata[219]), .Z(n6318));
Q_MX02 U2090 ( .S(rptr[0]), .A0(ififoRdata[154]), .A1(ififoRdata[218]), .Z(n6317));
Q_MX02 U2091 ( .S(rptr[0]), .A0(ififoRdata[153]), .A1(ififoRdata[217]), .Z(n6316));
Q_MX02 U2092 ( .S(rptr[0]), .A0(ififoRdata[152]), .A1(ififoRdata[216]), .Z(n6315));
Q_MX02 U2093 ( .S(rptr[0]), .A0(ififoRdata[151]), .A1(ififoRdata[215]), .Z(n6314));
Q_MX02 U2094 ( .S(rptr[0]), .A0(ififoRdata[150]), .A1(ififoRdata[214]), .Z(n6313));
Q_MX02 U2095 ( .S(rptr[0]), .A0(ififoRdata[149]), .A1(ififoRdata[213]), .Z(n6312));
Q_MX02 U2096 ( .S(rptr[0]), .A0(ififoRdata[148]), .A1(ififoRdata[212]), .Z(n6311));
Q_MX02 U2097 ( .S(rptr[0]), .A0(ififoRdata[147]), .A1(ififoRdata[211]), .Z(n6310));
Q_MX02 U2098 ( .S(rptr[0]), .A0(ififoRdata[146]), .A1(ififoRdata[210]), .Z(n6309));
Q_MX02 U2099 ( .S(rptr[0]), .A0(ififoRdata[145]), .A1(ififoRdata[209]), .Z(n6308));
Q_MX02 U2100 ( .S(rptr[0]), .A0(ififoRdata[144]), .A1(ififoRdata[208]), .Z(n6307));
Q_MX02 U2101 ( .S(rptr[0]), .A0(ififoRdata[143]), .A1(ififoRdata[207]), .Z(n6306));
Q_MX02 U2102 ( .S(rptr[0]), .A0(ififoRdata[142]), .A1(ififoRdata[206]), .Z(n6305));
Q_MX02 U2103 ( .S(rptr[0]), .A0(ififoRdata[141]), .A1(ififoRdata[205]), .Z(n6304));
Q_MX02 U2104 ( .S(rptr[0]), .A0(ififoRdata[140]), .A1(ififoRdata[204]), .Z(n6303));
Q_MX02 U2105 ( .S(rptr[0]), .A0(ififoRdata[139]), .A1(ififoRdata[203]), .Z(n6302));
Q_MX02 U2106 ( .S(rptr[0]), .A0(ififoRdata[138]), .A1(ififoRdata[202]), .Z(n6301));
Q_MX02 U2107 ( .S(rptr[0]), .A0(ififoRdata[137]), .A1(ififoRdata[201]), .Z(n6300));
Q_MX02 U2108 ( .S(rptr[0]), .A0(ififoRdata[136]), .A1(ififoRdata[200]), .Z(n6299));
Q_MX02 U2109 ( .S(rptr[0]), .A0(ififoRdata[135]), .A1(ififoRdata[199]), .Z(n6298));
Q_MX02 U2110 ( .S(rptr[0]), .A0(ififoRdata[134]), .A1(ififoRdata[198]), .Z(n6297));
Q_MX02 U2111 ( .S(rptr[0]), .A0(ififoRdata[133]), .A1(ififoRdata[197]), .Z(n6296));
Q_MX02 U2112 ( .S(rptr[0]), .A0(ififoRdata[132]), .A1(ififoRdata[196]), .Z(n6295));
Q_MX02 U2113 ( .S(rptr[0]), .A0(ififoRdata[131]), .A1(ififoRdata[195]), .Z(n6294));
Q_MX02 U2114 ( .S(rptr[0]), .A0(ififoRdata[130]), .A1(ififoRdata[194]), .Z(n6293));
Q_MX02 U2115 ( .S(rptr[0]), .A0(ififoRdata[129]), .A1(ififoRdata[193]), .Z(n6292));
Q_MX02 U2116 ( .S(rptr[0]), .A0(ififoRdata[128]), .A1(ififoRdata[192]), .Z(n6291));
Q_OR02 U2117 ( .A0(n6257), .A1(n6256), .Z(n6290));
Q_OR02 U2118 ( .A0(n6252), .A1(n6251), .Z(n6289));
Q_INV U2119 ( .A(n6289), .Z(n6288));
Q_NR03 U2120 ( .A0(n6290), .A1(n6289), .A2(scgGFreq), .Z(n5640));
Q_XNR2 U2121 ( .A0(wptr[0]), .A1(rptr[0]), .Z(n6287));
Q_XNR2 U2122 ( .A0(wptr[1]), .A1(rptr[1]), .Z(n6286));
Q_XNR2 U2123 ( .A0(wptr[2]), .A1(rptr[2]), .Z(n6285));
Q_XNR2 U2124 ( .A0(wptr[3]), .A1(rptr[3]), .Z(n6284));
Q_XNR2 U2125 ( .A0(wptr[4]), .A1(rptr[4]), .Z(n6283));
Q_XNR2 U2126 ( .A0(wptr[5]), .A1(rptr[5]), .Z(n6282));
Q_XNR2 U2127 ( .A0(wptr[6]), .A1(rptr[6]), .Z(n6281));
Q_XNR2 U2128 ( .A0(wptr[7]), .A1(rptr[7]), .Z(n6280));
Q_XNR2 U2129 ( .A0(wptr[8]), .A1(rptr[8]), .Z(n6279));
Q_XNR2 U2130 ( .A0(wptr[9]), .A1(rptr[9]), .Z(n6278));
Q_XNR2 U2131 ( .A0(wptr[10]), .A1(rptr[10]), .Z(n6277));
Q_XNR2 U2132 ( .A0(wptr[11]), .A1(rptr[11]), .Z(n6276));
Q_XNR2 U2133 ( .A0(wptr[12]), .A1(rptr[12]), .Z(n6275));
Q_XNR2 U2134 ( .A0(wptr[13]), .A1(rptr[13]), .Z(n6274));
Q_XNR2 U2135 ( .A0(wptr[14]), .A1(rptr[14]), .Z(n6273));
Q_XNR2 U2136 ( .A0(wptr[15]), .A1(rptr[15]), .Z(n6272));
Q_XNR2 U2137 ( .A0(wptr[16]), .A1(rptr[16]), .Z(n6271));
Q_AN03 U2138 ( .A0(n6271), .A1(n6272), .A2(n6273), .Z(n6270));
Q_AN03 U2139 ( .A0(n6274), .A1(n6275), .A2(n6276), .Z(n6269));
Q_AN03 U2140 ( .A0(n6277), .A1(n6278), .A2(n6279), .Z(n6268));
Q_AN03 U2141 ( .A0(n6280), .A1(n6281), .A2(n6282), .Z(n6267));
Q_AN03 U2142 ( .A0(n6283), .A1(n6284), .A2(n6285), .Z(n6266));
Q_AN03 U2143 ( .A0(n6286), .A1(n6287), .A2(n6270), .Z(n6265));
Q_AN03 U2144 ( .A0(n6269), .A1(n6268), .A2(n6267), .Z(n6264));
Q_AN03 U2145 ( .A0(n6266), .A1(n6265), .A2(n6264), .Z(n6263));
Q_INV U2146 ( .A(n6263), .Z(n5636));
Q_OR03 U2147 ( .A0(pktl[15]), .A1(pktl[14]), .A2(pktl[13]), .Z(n6262));
Q_OR03 U2148 ( .A0(pktl[12]), .A1(pktl[11]), .A2(pktl[10]), .Z(n6261));
Q_OR03 U2149 ( .A0(pktl[9]), .A1(pktl[8]), .A2(pktl[7]), .Z(n6260));
Q_OR03 U2150 ( .A0(pktl[6]), .A1(pktl[5]), .A2(pktl[4]), .Z(n6259));
Q_OR03 U2151 ( .A0(pktl[3]), .A1(pktl[2]), .A2(pktl[1]), .Z(n6258));
Q_OR03 U2152 ( .A0(pktl[0]), .A1(n6262), .A2(n6261), .Z(n6257));
Q_OR03 U2153 ( .A0(n6260), .A1(n6259), .A2(n6258), .Z(n6256));
Q_OR03 U2154 ( .A0(odly[11]), .A1(odly[10]), .A2(odly[9]), .Z(n6255));
Q_OR03 U2155 ( .A0(odly[8]), .A1(odly[7]), .A2(odly[6]), .Z(n6254));
Q_OR03 U2156 ( .A0(odly[5]), .A1(odly[4]), .A2(odly[3]), .Z(n6253));
Q_OR03 U2157 ( .A0(odly[2]), .A1(odly[1]), .A2(odly[0]), .Z(n6252));
Q_OR03 U2158 ( .A0(n6255), .A1(n6254), .A2(n6253), .Z(n6251));
Q_OR02 U2159 ( .A0(n6289), .A1(scgGFreq), .Z(n6250));
Q_INV U2160 ( .A(xc_top.GFLock1), .Z(n6249));
Q_ND02 U2161 ( .A0(n6250), .A1(n6249), .Z(n5639));
Q_OR02 U2162 ( .A0(pktl[13]), .A1(pktl[12]), .Z(n6248));
Q_OR03 U2163 ( .A0(pktl[15]), .A1(pktl[14]), .A2(n6248), .Z(n6247));
Q_OR02 U2164 ( .A0(pktl[9]), .A1(pktl[8]), .Z(n6246));
Q_OR03 U2165 ( .A0(pktl[11]), .A1(pktl[10]), .A2(n6246), .Z(n6245));
Q_OR02 U2166 ( .A0(pktl[5]), .A1(pktl[4]), .Z(n6244));
Q_OR03 U2167 ( .A0(pktl[7]), .A1(pktl[6]), .A2(n6244), .Z(n6243));
Q_OA21 U2168 ( .A0(pktl[1]), .A1(pktl[0]), .B0(pktl[3]), .Z(n6242));
Q_AN02 U2169 ( .A0(pktl[3]), .A1(pktl[2]), .Z(n6241));
Q_OR03 U2170 ( .A0(n6241), .A1(n6242), .A2(n6243), .Z(n6240));
Q_OR03 U2171 ( .A0(n6247), .A1(n6245), .A2(n6240), .Z(n5634));
Q_OR03 U2172 ( .A0(vlen[9]), .A1(vlen[8]), .A2(vlen[7]), .Z(n6239));
Q_OR03 U2173 ( .A0(vlen[6]), .A1(vlen[5]), .A2(vlen[4]), .Z(n6238));
Q_OR03 U2174 ( .A0(vlen[3]), .A1(vlen[2]), .A2(vlen[1]), .Z(n6237));
Q_OR03 U2175 ( .A0(vlen[0]), .A1(n6239), .A2(n6238), .Z(n6236));
Q_OR02 U2176 ( .A0(n6237), .A1(n6236), .Z(vmode));
Q_INV U2177 ( .A(rptr[3]), .Z(n6235));
Q_AD01HF U2178 ( .A0(rptr[4]), .B0(rptr[3]), .S(n6234), .CO(n6233));
Q_AD01HF U2179 ( .A0(rptr[5]), .B0(n6233), .S(n6232), .CO(n6231));
Q_AD01HF U2180 ( .A0(rptr[6]), .B0(n6231), .S(n6230), .CO(n6229));
Q_AD01HF U2181 ( .A0(rptr[7]), .B0(n6229), .S(n6228), .CO(n6227));
Q_AD01HF U2182 ( .A0(rptr[8]), .B0(n6227), .S(n6226), .CO(n6225));
Q_AD01HF U2183 ( .A0(rptr[9]), .B0(n6225), .S(n6224), .CO(n6223));
Q_AD01HF U2184 ( .A0(rptr[10]), .B0(n6223), .S(n6222), .CO(n6221));
Q_AD01HF U2185 ( .A0(rptr[11]), .B0(n6221), .S(n6220), .CO(n6219));
Q_AD01HF U2186 ( .A0(rptr[12]), .B0(n6219), .S(n6218), .CO(n6217));
Q_AD01HF U2187 ( .A0(rptr[13]), .B0(n6217), .S(n6216), .CO(n6215));
Q_AD01HF U2188 ( .A0(rptr[14]), .B0(n6215), .S(n6214), .CO(n6213));
Q_AD01HF U2189 ( .A0(rptr[15]), .B0(n6213), .S(n6212), .CO(n6211));
Q_XOR2 U2190 ( .A0(rptr[16]), .A1(n6211), .Z(n6210));
Q_INV U2191 ( .A(rptr[0]), .Z(n6209));
Q_AD01HF U2192 ( .A0(rptr[1]), .B0(rptr[0]), .S(n6208), .CO(n6207));
Q_AD01HF U2193 ( .A0(rptr[2]), .B0(n6207), .S(n6206), .CO(n6205));
Q_AD01HF U2194 ( .A0(rptr[3]), .B0(n6205), .S(n6204), .CO(n6203));
Q_AD01HF U2195 ( .A0(rptr[4]), .B0(n6203), .S(n6202), .CO(n6201));
Q_AD01HF U2196 ( .A0(rptr[5]), .B0(n6201), .S(n6200), .CO(n6199));
Q_AD01HF U2197 ( .A0(rptr[6]), .B0(n6199), .S(n6198), .CO(n6197));
Q_AD01HF U2198 ( .A0(rptr[7]), .B0(n6197), .S(n6196), .CO(n6195));
Q_AD01HF U2199 ( .A0(rptr[8]), .B0(n6195), .S(n6194), .CO(n6193));
Q_AD01HF U2200 ( .A0(rptr[9]), .B0(n6193), .S(n6192), .CO(n6191));
Q_AD01HF U2201 ( .A0(rptr[10]), .B0(n6191), .S(n6190), .CO(n6189));
Q_AD01HF U2202 ( .A0(rptr[11]), .B0(n6189), .S(n6188), .CO(n6187));
Q_AD01HF U2203 ( .A0(rptr[12]), .B0(n6187), .S(n6186), .CO(n6185));
Q_AD01HF U2204 ( .A0(rptr[13]), .B0(n6185), .S(n6184), .CO(n6183));
Q_AD01HF U2205 ( .A0(rptr[14]), .B0(n6183), .S(n6182), .CO(n6181));
Q_AD01HF U2206 ( .A0(rptr[15]), .B0(n6181), .S(n6180), .CO(n6179));
Q_XOR2 U2207 ( .A0(n6178), .A1(rptr[16]), .Z(n5899));
Q_INV U2208 ( .A(pktl[3]), .Z(n6177));
Q_XNR2 U2209 ( .A0(pktl[4]), .A1(pktl[3]), .Z(n6176));
Q_OR02 U2210 ( .A0(pktl[4]), .A1(pktl[3]), .Z(n6175));
Q_XNR2 U2211 ( .A0(pktl[5]), .A1(n6175), .Z(n6174));
Q_OR02 U2212 ( .A0(pktl[5]), .A1(n6175), .Z(n6173));
Q_XNR2 U2213 ( .A0(pktl[6]), .A1(n6173), .Z(n6172));
Q_OR02 U2214 ( .A0(pktl[6]), .A1(n6173), .Z(n6171));
Q_XNR2 U2215 ( .A0(pktl[7]), .A1(n6171), .Z(n6170));
Q_OR02 U2216 ( .A0(pktl[7]), .A1(n6171), .Z(n6169));
Q_XNR2 U2217 ( .A0(pktl[8]), .A1(n6169), .Z(n6168));
Q_OR02 U2218 ( .A0(pktl[8]), .A1(n6169), .Z(n6167));
Q_XNR2 U2219 ( .A0(pktl[9]), .A1(n6167), .Z(n6166));
Q_OR02 U2220 ( .A0(pktl[9]), .A1(n6167), .Z(n6165));
Q_XNR2 U2221 ( .A0(pktl[10]), .A1(n6165), .Z(n6164));
Q_OR02 U2222 ( .A0(pktl[10]), .A1(n6165), .Z(n6163));
Q_XNR2 U2223 ( .A0(pktl[11]), .A1(n6163), .Z(n6162));
Q_OR02 U2224 ( .A0(pktl[11]), .A1(n6163), .Z(n6161));
Q_XNR2 U2225 ( .A0(pktl[12]), .A1(n6161), .Z(n6160));
Q_OR02 U2226 ( .A0(pktl[12]), .A1(n6161), .Z(n6159));
Q_XNR2 U2227 ( .A0(pktl[13]), .A1(n6159), .Z(n6158));
Q_OR02 U2228 ( .A0(pktl[13]), .A1(n6159), .Z(n6157));
Q_XNR2 U2229 ( .A0(pktl[14]), .A1(n6157), .Z(n6156));
Q_OR02 U2230 ( .A0(pktl[14]), .A1(n6157), .Z(n6155));
Q_XNR2 U2231 ( .A0(pktl[15]), .A1(n6155), .Z(n6154));
Q_INV U2232 ( .A(pktl[0]), .Z(n6153));
Q_INV U2233 ( .A(pktl[1]), .Z(n6152));
Q_INV U2234 ( .A(pktl[2]), .Z(n6151));
Q_INV U2235 ( .A(pktl[4]), .Z(n6150));
Q_INV U2236 ( .A(pktl[5]), .Z(n6149));
Q_INV U2237 ( .A(pktl[6]), .Z(n6148));
Q_INV U2238 ( .A(pktl[7]), .Z(n6147));
Q_INV U2239 ( .A(pktl[8]), .Z(n6146));
Q_XNR2 U2240 ( .A0(vlen[0]), .A1(n6153), .Z(n6145));
Q_OR02 U2241 ( .A0(vlen[0]), .A1(n6153), .Z(n6144));
Q_AD01 U2242 ( .CI(n6144), .A0(vlen[1]), .B0(n6152), .S(n6143), .CO(n6142));
Q_AD02 U2243 ( .CI(n6142), .A0(vlen[2]), .A1(vlen[3]), .B0(n6151), .B1(n6177), .S0(n6141), .S1(n6140), .CO(n6139));
Q_AD02 U2244 ( .CI(n6139), .A0(vlen[4]), .A1(vlen[5]), .B0(n6150), .B1(n6149), .S0(n6138), .S1(n6137), .CO(n6136));
Q_AD02 U2245 ( .CI(n6136), .A0(vlen[6]), .A1(vlen[7]), .B0(n6148), .B1(n6147), .S0(n6135), .S1(n6134), .CO(n6133));
Q_OR03 U2246 ( .A0(n6145), .A1(n6143), .A2(n6141), .Z(n6130));
Q_OR03 U2247 ( .A0(n6140), .A1(n6130), .A2(n6138), .Z(n6129));
Q_OR03 U2248 ( .A0(n6137), .A1(n6129), .A2(n6135), .Z(n6128));
Q_OR03 U2249 ( .A0(n6134), .A1(n6128), .A2(n6132), .Z(n6127));
Q_NR02 U2250 ( .A0(n6131), .A1(n6127), .Z(n6126));
Q_AD02 U2251 ( .CI(n6126), .A0(rptr[0]), .A1(rptr[1]), .B0(pktl[0]), .B1(pktl[1]), .S0(n6125), .S1(n6124), .CO(n6123));
Q_AD02 U2252 ( .CI(n6123), .A0(rptr[2]), .A1(rptr[3]), .B0(pktl[2]), .B1(pktl[3]), .S0(n6122), .S1(n6121), .CO(n6120));
Q_AD02 U2253 ( .CI(n6120), .A0(rptr[4]), .A1(rptr[5]), .B0(pktl[4]), .B1(pktl[5]), .S0(n6119), .S1(n6118), .CO(n6117));
Q_AD02 U2254 ( .CI(n6117), .A0(rptr[6]), .A1(rptr[7]), .B0(pktl[6]), .B1(pktl[7]), .S0(n6116), .S1(n6115), .CO(n6114));
Q_AD02 U2255 ( .CI(n6114), .A0(rptr[8]), .A1(rptr[9]), .B0(pktl[8]), .B1(pktl[9]), .S0(n6113), .S1(n6112), .CO(n6111));
Q_AD02 U2256 ( .CI(n6111), .A0(rptr[10]), .A1(rptr[11]), .B0(pktl[10]), .B1(pktl[11]), .S0(n6110), .S1(n6109), .CO(n6108));
Q_AD02 U2257 ( .CI(n6108), .A0(rptr[12]), .A1(rptr[13]), .B0(pktl[12]), .B1(pktl[13]), .S0(n6107), .S1(n6106), .CO(n6105));
Q_AD02 U2258 ( .CI(n6105), .A0(rptr[14]), .A1(rptr[15]), .B0(pktl[14]), .B1(pktl[15]), .S0(n6104), .S1(n6103), .CO(n6102));
Q_XOR2 U2259 ( .A0(rptr[16]), .A1(n6102), .Z(n6101));
Q_INV U2260 ( .A(odly[0]), .Z(n6100));
Q_XNR2 U2261 ( .A0(odly[1]), .A1(odly[0]), .Z(n6099));
Q_OR02 U2262 ( .A0(odly[1]), .A1(odly[0]), .Z(n6098));
Q_XNR2 U2263 ( .A0(odly[2]), .A1(n6098), .Z(n6097));
Q_OR02 U2264 ( .A0(odly[2]), .A1(n6098), .Z(n6096));
Q_XNR2 U2265 ( .A0(odly[3]), .A1(n6096), .Z(n6095));
Q_OR02 U2266 ( .A0(odly[3]), .A1(n6096), .Z(n6094));
Q_XNR2 U2267 ( .A0(odly[4]), .A1(n6094), .Z(n6093));
Q_OR02 U2268 ( .A0(odly[4]), .A1(n6094), .Z(n6092));
Q_XNR2 U2269 ( .A0(odly[5]), .A1(n6092), .Z(n6091));
Q_OR02 U2270 ( .A0(odly[5]), .A1(n6092), .Z(n6090));
Q_XNR2 U2271 ( .A0(odly[6]), .A1(n6090), .Z(n6089));
Q_OR02 U2272 ( .A0(odly[6]), .A1(n6090), .Z(n6088));
Q_XNR2 U2273 ( .A0(odly[7]), .A1(n6088), .Z(n6087));
Q_OR02 U2274 ( .A0(odly[7]), .A1(n6088), .Z(n6086));
Q_XNR2 U2275 ( .A0(odly[8]), .A1(n6086), .Z(n6085));
Q_OR02 U2276 ( .A0(odly[8]), .A1(n6086), .Z(n6084));
Q_XNR2 U2277 ( .A0(odly[9]), .A1(n6084), .Z(n6083));
Q_OR02 U2278 ( .A0(odly[9]), .A1(n6084), .Z(n6082));
Q_XNR2 U2279 ( .A0(odly[10]), .A1(n6082), .Z(n6081));
Q_OR02 U2280 ( .A0(odly[10]), .A1(n6082), .Z(n6080));
Q_XNR2 U2281 ( .A0(odly[11]), .A1(n6080), .Z(n6079));
Q_MX02 U2282 ( .S(vmode), .A0(tmpData[0]), .A1(vhead[0]), .Z(head[0]));
Q_MX02 U2283 ( .S(vmode), .A0(tmpData[1]), .A1(vhead[1]), .Z(head[1]));
Q_MX02 U2284 ( .S(vmode), .A0(tmpData[2]), .A1(vhead[2]), .Z(head[2]));
Q_MX02 U2285 ( .S(vmode), .A0(tmpData[3]), .A1(vhead[3]), .Z(head[3]));
Q_MX02 U2286 ( .S(vmode), .A0(tmpData[4]), .A1(vhead[4]), .Z(head[4]));
Q_MX02 U2287 ( .S(vmode), .A0(tmpData[5]), .A1(vhead[5]), .Z(head[5]));
Q_MX02 U2288 ( .S(vmode), .A0(tmpData[6]), .A1(vhead[6]), .Z(head[6]));
Q_MX02 U2289 ( .S(vmode), .A0(tmpData[7]), .A1(vhead[7]), .Z(head[7]));
Q_MX02 U2290 ( .S(vmode), .A0(tmpData[8]), .A1(vhead[8]), .Z(head[8]));
Q_MX02 U2291 ( .S(vmode), .A0(tmpData[9]), .A1(vhead[9]), .Z(head[9]));
Q_MX02 U2292 ( .S(vmode), .A0(tmpData[10]), .A1(vhead[10]), .Z(head[10]));
Q_MX02 U2293 ( .S(vmode), .A0(tmpData[11]), .A1(vhead[11]), .Z(head[11]));
Q_MX02 U2294 ( .S(vmode), .A0(tmpData[12]), .A1(vhead[12]), .Z(head[12]));
Q_MX02 U2295 ( .S(vmode), .A0(tmpData[13]), .A1(vhead[13]), .Z(head[13]));
Q_MX02 U2296 ( .S(vmode), .A0(tmpData[14]), .A1(vhead[14]), .Z(head[14]));
Q_MX02 U2297 ( .S(vmode), .A0(tmpData[15]), .A1(vhead[15]), .Z(head[15]));
Q_MX02 U2298 ( .S(vmode), .A0(tmpData[16]), .A1(vhead[16]), .Z(head[16]));
Q_MX02 U2299 ( .S(vmode), .A0(tmpData[17]), .A1(vhead[17]), .Z(head[17]));
Q_MX02 U2300 ( .S(vmode), .A0(tmpData[18]), .A1(vhead[18]), .Z(head[18]));
Q_MX02 U2301 ( .S(vmode), .A0(tmpData[19]), .A1(vhead[19]), .Z(head[19]));
Q_MX02 U2302 ( .S(vmode), .A0(tmpData[20]), .A1(vhead[20]), .Z(head[20]));
Q_MX02 U2303 ( .S(vmode), .A0(tmpData[21]), .A1(vhead[21]), .Z(head[21]));
Q_MX02 U2304 ( .S(vmode), .A0(tmpData[22]), .A1(vhead[22]), .Z(head[22]));
Q_MX02 U2305 ( .S(vmode), .A0(tmpData[23]), .A1(vhead[23]), .Z(head[23]));
Q_MX02 U2306 ( .S(vmode), .A0(tmpData[24]), .A1(vhead[24]), .Z(head[24]));
Q_MX02 U2307 ( .S(vmode), .A0(tmpData[25]), .A1(vhead[25]), .Z(head[25]));
Q_MX02 U2308 ( .S(vmode), .A0(tmpData[26]), .A1(vhead[26]), .Z(head[26]));
Q_MX02 U2309 ( .S(vmode), .A0(tmpData[27]), .A1(vhead[27]), .Z(head[27]));
Q_MX02 U2310 ( .S(vmode), .A0(tmpData[28]), .A1(vhead[28]), .Z(head[28]));
Q_MX02 U2311 ( .S(vmode), .A0(tmpData[29]), .A1(vhead[29]), .Z(head[29]));
Q_MX02 U2312 ( .S(vmode), .A0(tmpData[30]), .A1(vhead[30]), .Z(head[30]));
Q_MX02 U2313 ( .S(vmode), .A0(tmpData[31]), .A1(vhead[31]), .Z(head[31]));
Q_MX02 U2314 ( .S(vmode), .A0(tmpData[32]), .A1(vhead[32]), .Z(head[32]));
Q_MX02 U2315 ( .S(vmode), .A0(tmpData[33]), .A1(vhead[33]), .Z(head[33]));
Q_MX02 U2316 ( .S(vmode), .A0(tmpData[34]), .A1(vhead[34]), .Z(head[34]));
Q_MX02 U2317 ( .S(vmode), .A0(tmpData[35]), .A1(vhead[35]), .Z(head[35]));
Q_MX02 U2318 ( .S(vmode), .A0(tmpData[36]), .A1(vhead[36]), .Z(head[36]));
Q_MX02 U2319 ( .S(vmode), .A0(tmpData[37]), .A1(vhead[37]), .Z(head[37]));
Q_MX02 U2320 ( .S(vmode), .A0(tmpData[38]), .A1(vhead[38]), .Z(head[38]));
Q_MX02 U2321 ( .S(vmode), .A0(tmpData[39]), .A1(vhead[39]), .Z(head[39]));
Q_MX02 U2322 ( .S(vmode), .A0(tmpData[40]), .A1(vhead[40]), .Z(head[40]));
Q_MX02 U2323 ( .S(vmode), .A0(tmpData[41]), .A1(vhead[41]), .Z(head[41]));
Q_MX02 U2324 ( .S(vmode), .A0(tmpData[42]), .A1(vhead[42]), .Z(head[42]));
Q_MX02 U2325 ( .S(vmode), .A0(tmpData[43]), .A1(vhead[43]), .Z(head[43]));
Q_MX02 U2326 ( .S(vmode), .A0(tmpData[44]), .A1(vhead[44]), .Z(head[44]));
Q_MX02 U2327 ( .S(vmode), .A0(tmpData[45]), .A1(vhead[45]), .Z(head[45]));
Q_MX02 U2328 ( .S(vmode), .A0(tmpData[46]), .A1(vhead[46]), .Z(head[46]));
Q_MX02 U2329 ( .S(vmode), .A0(tmpData[47]), .A1(vhead[47]), .Z(head[47]));
Q_MX02 U2330 ( .S(vmode), .A0(tmpData[48]), .A1(vhead[48]), .Z(head[48]));
Q_MX02 U2331 ( .S(vmode), .A0(tmpData[49]), .A1(vhead[49]), .Z(head[49]));
Q_MX02 U2332 ( .S(vmode), .A0(tmpData[50]), .A1(vhead[50]), .Z(head[50]));
Q_MX02 U2333 ( .S(vmode), .A0(tmpData[51]), .A1(vhead[51]), .Z(head[51]));
Q_MX02 U2334 ( .S(vmode), .A0(tmpData[52]), .A1(vhead[52]), .Z(head[52]));
Q_MX02 U2335 ( .S(vmode), .A0(tmpData[53]), .A1(vhead[53]), .Z(head[53]));
Q_MX02 U2336 ( .S(vmode), .A0(tmpData[54]), .A1(vhead[54]), .Z(head[54]));
Q_MX02 U2337 ( .S(vmode), .A0(tmpData[55]), .A1(vhead[55]), .Z(head[55]));
Q_MX02 U2338 ( .S(vmode), .A0(tmpData[56]), .A1(vhead[56]), .Z(head[56]));
Q_MX02 U2339 ( .S(vmode), .A0(tmpData[57]), .A1(vhead[57]), .Z(head[57]));
Q_MX02 U2340 ( .S(vmode), .A0(tmpData[58]), .A1(vhead[58]), .Z(head[58]));
Q_MX02 U2341 ( .S(vmode), .A0(tmpData[59]), .A1(vhead[59]), .Z(head[59]));
Q_MX02 U2342 ( .S(vmode), .A0(tmpData[60]), .A1(vhead[60]), .Z(head[60]));
Q_MX02 U2343 ( .S(vmode), .A0(tmpData[61]), .A1(vhead[61]), .Z(head[61]));
Q_MX02 U2344 ( .S(vmode), .A0(tmpData[62]), .A1(vhead[62]), .Z(head[62]));
Q_MX02 U2345 ( .S(vmode), .A0(tmpData[63]), .A1(vhead[63]), .Z(head[63]));
Q_INV U2346 ( .A(head[10]), .Z(n6078));
Q_AN03 U2347 ( .A0(n6078), .A1(n6075), .A2(n6074), .Z(n6077));
Q_AN03 U2348 ( .A0(n6070), .A1(n6069), .A2(n6077), .Z(n6076));
Q_AN02 U2349 ( .A0(n6067), .A1(n6076), .Z(n5638));
Q_AN03 U2350 ( .A0(head[31]), .A1(head[30]), .A2(head[29]), .Z(n6075));
Q_AN03 U2351 ( .A0(head[28]), .A1(head[27]), .A2(head[26]), .Z(n6074));
Q_AN03 U2352 ( .A0(head[25]), .A1(head[24]), .A2(head[23]), .Z(n6073));
Q_AN03 U2353 ( .A0(head[22]), .A1(head[21]), .A2(head[20]), .Z(n6072));
Q_AN03 U2354 ( .A0(head[19]), .A1(head[18]), .A2(head[17]), .Z(n6071));
Q_AN03 U2355 ( .A0(head[16]), .A1(head[15]), .A2(head[14]), .Z(n6070));
Q_AN03 U2356 ( .A0(head[13]), .A1(head[12]), .A2(head[11]), .Z(n6069));
Q_AN03 U2357 ( .A0(head[10]), .A1(n6075), .A2(n6074), .Z(n6068));
Q_AN03 U2358 ( .A0(n6073), .A1(n6072), .A2(n6071), .Z(n6067));
Q_AN03 U2359 ( .A0(n6070), .A1(n6069), .A2(n6068), .Z(n6066));
Q_AN02 U2360 ( .A0(n6067), .A1(n6066), .Z(n5637));
Q_OR02 U2361 ( .A0(head[39]), .A1(head[38]), .Z(n6065));
Q_OR03 U2362 ( .A0(head[41]), .A1(head[40]), .A2(n6065), .Z(n6064));
Q_AN02 U2363 ( .A0(head[35]), .A1(head[34]), .Z(n6063));
Q_OR03 U2364 ( .A0(head[37]), .A1(head[36]), .A2(n6063), .Z(n6062));
Q_OR03 U2365 ( .A0(n6064), .A1(n6062), .A2(n6061), .Z(n5635));
Q_INV U2366 ( .A(head[35]), .Z(n6060));
Q_XNR2 U2367 ( .A0(head[36]), .A1(head[35]), .Z(n6059));
Q_OR02 U2368 ( .A0(head[36]), .A1(head[35]), .Z(n6058));
Q_XNR2 U2369 ( .A0(head[37]), .A1(n6058), .Z(n6057));
Q_OR02 U2370 ( .A0(head[37]), .A1(n6058), .Z(n6056));
Q_XNR2 U2371 ( .A0(head[38]), .A1(n6056), .Z(n6055));
Q_OR02 U2372 ( .A0(head[38]), .A1(n6056), .Z(n6054));
Q_XNR2 U2373 ( .A0(head[39]), .A1(n6054), .Z(n6053));
Q_OR02 U2374 ( .A0(head[39]), .A1(n6054), .Z(n6052));
Q_XNR2 U2375 ( .A0(head[40]), .A1(n6052), .Z(n6051));
Q_OR02 U2376 ( .A0(head[40]), .A1(n6052), .Z(n6050));
Q_XNR2 U2377 ( .A0(head[41]), .A1(n6050), .Z(n6049));
Q_NR03 U2378 ( .A0(head[41]), .A1(n6050), .A2(n5655), .Z(n5796));
Q_XNR2 U2379 ( .A0(rptr[0]), .A1(head[0]), .Z(n6048));
Q_OR02 U2380 ( .A0(rptr[0]), .A1(head[0]), .Z(n6047));
Q_AD01 U2381 ( .CI(n6047), .A0(rptr[1]), .B0(head[1]), .S(n6046), .CO(n6045));
Q_AD02 U2382 ( .CI(n6045), .A0(rptr[2]), .A1(rptr[3]), .B0(head[2]), .B1(head[3]), .S0(n6044), .S1(n6043), .CO(n6042));
Q_AD02 U2383 ( .CI(n6042), .A0(rptr[4]), .A1(rptr[5]), .B0(head[4]), .B1(head[5]), .S0(n6041), .S1(n6040), .CO(n6039));
Q_AD02 U2384 ( .CI(n6039), .A0(rptr[6]), .A1(rptr[7]), .B0(head[6]), .B1(head[7]), .S0(n6038), .S1(n6037), .CO(n6036));
Q_AD02 U2385 ( .CI(n6036), .A0(rptr[8]), .A1(rptr[9]), .B0(head[8]), .B1(head[9]), .S0(n6035), .S1(n6034), .CO(n6033));
Q_AD01HF U2386 ( .A0(rptr[10]), .B0(n6033), .S(n6032), .CO(n6031));
Q_AD01HF U2387 ( .A0(rptr[11]), .B0(n6031), .S(n6030), .CO(n6029));
Q_AD01HF U2388 ( .A0(rptr[12]), .B0(n6029), .S(n6028), .CO(n6027));
Q_AD01HF U2389 ( .A0(rptr[13]), .B0(n6027), .S(n6026), .CO(n6025));
Q_AD01HF U2390 ( .A0(rptr[14]), .B0(n6025), .S(n6024), .CO(n6023));
Q_AD01HF U2391 ( .A0(rptr[15]), .B0(n6023), .S(n6022), .CO(n6021));
Q_XNR2 U2392 ( .A0(n6005), .A1(n6006), .Z(n6020));
Q_OR02 U2393 ( .A0(n6005), .A1(n6006), .Z(n6019));
Q_XNR2 U2394 ( .A0(n6004), .A1(n6019), .Z(n6018));
Q_OR02 U2395 ( .A0(n6004), .A1(n6019), .Z(n6017));
Q_XNR2 U2396 ( .A0(n6003), .A1(n6017), .Z(n6016));
Q_OR02 U2397 ( .A0(n6003), .A1(n6017), .Z(n6015));
Q_XNR2 U2398 ( .A0(n6002), .A1(n6015), .Z(n6014));
Q_OR02 U2399 ( .A0(n6002), .A1(n6015), .Z(n6013));
Q_XNR2 U2400 ( .A0(n6001), .A1(n6013), .Z(n6012));
Q_OR02 U2401 ( .A0(n6001), .A1(n6013), .Z(n6011));
Q_XNR2 U2402 ( .A0(n6000), .A1(n6011), .Z(n6010));
Q_MX02 U2403 ( .S(vmode), .A0(head[0]), .A1(vlen[0]), .Z(n6009));
Q_MX02 U2404 ( .S(vmode), .A0(head[1]), .A1(vlen[1]), .Z(n6008));
Q_MX02 U2405 ( .S(vmode), .A0(head[2]), .A1(vlen[2]), .Z(n6007));
Q_MX02 U2406 ( .S(vmode), .A0(head[3]), .A1(vlen[3]), .Z(n6006));
Q_MX02 U2407 ( .S(vmode), .A0(head[4]), .A1(vlen[4]), .Z(n6005));
Q_MX02 U2408 ( .S(vmode), .A0(head[5]), .A1(vlen[5]), .Z(n6004));
Q_MX02 U2409 ( .S(vmode), .A0(head[6]), .A1(vlen[6]), .Z(n6003));
Q_MX02 U2410 ( .S(vmode), .A0(head[7]), .A1(vlen[7]), .Z(n6002));
Q_MX02 U2411 ( .S(vmode), .A0(head[8]), .A1(vlen[8]), .Z(n6001));
Q_MX02 U2412 ( .S(vmode), .A0(head[9]), .A1(vlen[9]), .Z(n6000));
Q_OR02 U2413 ( .A0(n284), .A1(head[10]), .Z(tId[0]));
Q_OR02 U2414 ( .A0(n284), .A1(head[11]), .Z(tId[1]));
Q_OR02 U2415 ( .A0(n284), .A1(head[12]), .Z(tId[2]));
Q_OR02 U2416 ( .A0(n284), .A1(head[13]), .Z(tId[3]));
Q_OR02 U2417 ( .A0(n284), .A1(head[14]), .Z(tId[4]));
Q_OR02 U2418 ( .A0(n284), .A1(head[15]), .Z(tId[5]));
Q_OR02 U2419 ( .A0(n284), .A1(head[16]), .Z(tId[6]));
Q_OR02 U2420 ( .A0(n284), .A1(head[17]), .Z(tId[7]));
Q_OR02 U2421 ( .A0(n284), .A1(head[18]), .Z(tId[8]));
Q_OR02 U2422 ( .A0(n284), .A1(head[19]), .Z(tId[9]));
Q_OR02 U2423 ( .A0(n284), .A1(head[20]), .Z(tId[10]));
Q_OR02 U2424 ( .A0(n284), .A1(head[21]), .Z(tId[11]));
Q_OR02 U2425 ( .A0(n284), .A1(head[22]), .Z(tId[12]));
Q_OR02 U2426 ( .A0(n284), .A1(head[23]), .Z(tId[13]));
Q_OR02 U2427 ( .A0(n284), .A1(head[24]), .Z(tId[14]));
Q_OR02 U2428 ( .A0(n284), .A1(head[25]), .Z(tId[15]));
Q_OR02 U2429 ( .A0(n284), .A1(head[26]), .Z(tId[16]));
Q_OR02 U2430 ( .A0(n284), .A1(head[27]), .Z(tId[17]));
Q_OR02 U2431 ( .A0(n284), .A1(head[28]), .Z(tId[18]));
Q_OR02 U2432 ( .A0(n284), .A1(head[29]), .Z(tId[19]));
Q_OR02 U2433 ( .A0(n284), .A1(head[30]), .Z(tId[20]));
Q_OR02 U2434 ( .A0(n284), .A1(head[31]), .Z(tId[21]));
Q_INV U2435 ( .A(n5999), .Z(n5699));
Q_XNR2 U2436 ( .A0(vlen[4]), .A1(vlen[3]), .Z(n5998));
Q_OR02 U2437 ( .A0(vlen[4]), .A1(vlen[3]), .Z(n5997));
Q_XNR2 U2438 ( .A0(vlen[5]), .A1(n5997), .Z(n5996));
Q_OR02 U2439 ( .A0(vlen[5]), .A1(n5997), .Z(n5995));
Q_XNR2 U2440 ( .A0(vlen[6]), .A1(n5995), .Z(n5994));
Q_OR02 U2441 ( .A0(vlen[6]), .A1(n5995), .Z(n5993));
Q_XNR2 U2442 ( .A0(vlen[7]), .A1(n5993), .Z(n5992));
Q_OR02 U2443 ( .A0(vlen[7]), .A1(n5993), .Z(n5991));
Q_XNR2 U2444 ( .A0(vlen[8]), .A1(n5991), .Z(n5990));
Q_OR02 U2445 ( .A0(vlen[8]), .A1(n5991), .Z(n5989));
Q_XNR2 U2446 ( .A0(vlen[9]), .A1(n5989), .Z(n5988));
Q_INV U2447 ( .A(head[32]), .Z(n5987));
Q_INV U2448 ( .A(head[33]), .Z(n5986));
Q_INV U2449 ( .A(head[34]), .Z(n5985));
Q_INV U2450 ( .A(head[36]), .Z(n5984));
Q_INV U2451 ( .A(head[37]), .Z(n5983));
Q_INV U2452 ( .A(head[38]), .Z(n5982));
Q_INV U2453 ( .A(head[39]), .Z(n5981));
Q_INV U2454 ( .A(head[40]), .Z(n5980));
Q_XNR3 U2455 ( .A0(head[41]), .A1(n6000), .A2(n5966), .Z(n5965));
Q_XNR2 U2456 ( .A0(n5987), .A1(n6009), .Z(n5979));
Q_OR02 U2457 ( .A0(n5987), .A1(n6009), .Z(n5978));
Q_AD02 U2458 ( .CI(n5978), .A0(n5986), .A1(n5985), .B0(n6008), .B1(n6007), .S0(n5977), .S1(n5976), .CO(n5975));
Q_AD02 U2459 ( .CI(n5975), .A0(n6060), .A1(n5984), .B0(n6006), .B1(n6005), .S0(n5974), .S1(n5973), .CO(n5972));
Q_AD02 U2460 ( .CI(n5972), .A0(n5983), .A1(n5982), .B0(n6004), .B1(n6003), .S0(n5971), .S1(n5970), .CO(n5969));
Q_AD02 U2461 ( .CI(n5969), .A0(n5981), .A1(n5980), .B0(n6002), .B1(n6001), .S0(n5968), .S1(n5967), .CO(n5966));
Q_OR03 U2462 ( .A0(n5979), .A1(n5977), .A2(n5976), .Z(n5964));
Q_OR03 U2463 ( .A0(n5974), .A1(n5964), .A2(n5973), .Z(n5963));
Q_OR03 U2464 ( .A0(n5971), .A1(n5963), .A2(n5970), .Z(n5962));
Q_OR03 U2465 ( .A0(n5968), .A1(n5962), .A2(n5967), .Z(n5961));
Q_NR02 U2466 ( .A0(n5965), .A1(n5961), .Z(n5960));
Q_AD02 U2467 ( .CI(n5960), .A0(rptr[0]), .A1(rptr[1]), .B0(head[32]), .B1(head[33]), .S0(n5959), .S1(n5958), .CO(n5957));
Q_AD02 U2468 ( .CI(n5957), .A0(rptr[2]), .A1(rptr[3]), .B0(head[34]), .B1(head[35]), .S0(n5956), .S1(n5955), .CO(n5954));
Q_AD02 U2469 ( .CI(n5954), .A0(rptr[4]), .A1(rptr[5]), .B0(head[36]), .B1(head[37]), .S0(n5953), .S1(n5952), .CO(n5951));
Q_AD02 U2470 ( .CI(n5951), .A0(rptr[6]), .A1(rptr[7]), .B0(head[38]), .B1(head[39]), .S0(n5950), .S1(n5949), .CO(n5948));
Q_AD02 U2471 ( .CI(n5948), .A0(rptr[8]), .A1(rptr[9]), .B0(head[40]), .B1(head[41]), .S0(n5947), .S1(n5946), .CO(n5945));
Q_AD01HF U2472 ( .A0(rptr[10]), .B0(n5945), .S(n5944), .CO(n5943));
Q_AD01HF U2473 ( .A0(rptr[11]), .B0(n5943), .S(n5942), .CO(n5941));
Q_AD01HF U2474 ( .A0(rptr[12]), .B0(n5941), .S(n5940), .CO(n5939));
Q_AD01HF U2475 ( .A0(rptr[13]), .B0(n5939), .S(n5938), .CO(n5937));
Q_AD01HF U2476 ( .A0(rptr[14]), .B0(n5937), .S(n5936), .CO(n5935));
Q_AD01HF U2477 ( .A0(rptr[15]), .B0(n5935), .S(n5934), .CO(n5933));
Q_XOR2 U2478 ( .A0(rptr[16]), .A1(n5933), .Z(n5932));
Q_MX02 U2479 ( .S(n5648), .A0(n6048), .A1(n6209), .Z(n5931));
Q_MX04 U2480 ( .S0(n5648), .S1(n5647), .A0(rptr[0]), .A1(n6125), .A2(n5959), .A3(rptr[0]), .Z(n5930));
Q_MX02 U2481 ( .S(n5646), .A0(n5930), .A1(n5931), .Z(rptrN[0]));
Q_MX02 U2482 ( .S(n5648), .A0(n6046), .A1(n6208), .Z(n5929));
Q_MX04 U2483 ( .S0(n5648), .S1(n5647), .A0(rptr[1]), .A1(n6124), .A2(n5958), .A3(rptr[1]), .Z(n5928));
Q_MX02 U2484 ( .S(n5646), .A0(n5928), .A1(n5929), .Z(rptrN[1]));
Q_MX02 U2485 ( .S(n5648), .A0(n6044), .A1(n6206), .Z(n5927));
Q_MX04 U2486 ( .S0(n5648), .S1(n5647), .A0(rptr[2]), .A1(n6122), .A2(n5956), .A3(rptr[2]), .Z(n5926));
Q_MX02 U2487 ( .S(n5646), .A0(n5926), .A1(n5927), .Z(rptrN[2]));
Q_MX02 U2488 ( .S(n5648), .A0(n6043), .A1(n6204), .Z(n5925));
Q_MX04 U2489 ( .S0(n5648), .S1(n5647), .A0(rptr[3]), .A1(n6121), .A2(n5955), .A3(n6235), .Z(n5924));
Q_MX02 U2490 ( .S(n5646), .A0(n5924), .A1(n5925), .Z(rptrN[3]));
Q_MX02 U2491 ( .S(n5648), .A0(n6041), .A1(n6202), .Z(n5923));
Q_MX04 U2492 ( .S0(n5648), .S1(n5647), .A0(rptr[4]), .A1(n6119), .A2(n5953), .A3(n6234), .Z(n5922));
Q_MX02 U2493 ( .S(n5646), .A0(n5922), .A1(n5923), .Z(rptrN[4]));
Q_MX02 U2494 ( .S(n5648), .A0(n6040), .A1(n6200), .Z(n5921));
Q_MX04 U2495 ( .S0(n5648), .S1(n5647), .A0(rptr[5]), .A1(n6118), .A2(n5952), .A3(n6232), .Z(n5920));
Q_MX02 U2496 ( .S(n5646), .A0(n5920), .A1(n5921), .Z(rptrN[5]));
Q_MX02 U2497 ( .S(n5648), .A0(n6038), .A1(n6198), .Z(n5919));
Q_MX04 U2498 ( .S0(n5648), .S1(n5647), .A0(rptr[6]), .A1(n6116), .A2(n5950), .A3(n6230), .Z(n5918));
Q_MX02 U2499 ( .S(n5646), .A0(n5918), .A1(n5919), .Z(rptrN[6]));
Q_MX02 U2500 ( .S(n5648), .A0(n6037), .A1(n6196), .Z(n5917));
Q_MX04 U2501 ( .S0(n5648), .S1(n5647), .A0(rptr[7]), .A1(n6115), .A2(n5949), .A3(n6228), .Z(n5916));
Q_MX02 U2502 ( .S(n5646), .A0(n5916), .A1(n5917), .Z(rptrN[7]));
Q_MX02 U2503 ( .S(n5648), .A0(n6035), .A1(n6194), .Z(n5915));
Q_MX04 U2504 ( .S0(n5648), .S1(n5647), .A0(rptr[8]), .A1(n6113), .A2(n5947), .A3(n6226), .Z(n5914));
Q_MX02 U2505 ( .S(n5646), .A0(n5914), .A1(n5915), .Z(rptrN[8]));
Q_MX02 U2506 ( .S(n5648), .A0(n6034), .A1(n6192), .Z(n5913));
Q_MX04 U2507 ( .S0(n5648), .S1(n5647), .A0(rptr[9]), .A1(n6112), .A2(n5946), .A3(n6224), .Z(n5912));
Q_MX02 U2508 ( .S(n5646), .A0(n5912), .A1(n5913), .Z(rptrN[9]));
Q_MX02 U2509 ( .S(n5648), .A0(n6032), .A1(n6190), .Z(n5911));
Q_MX04 U2510 ( .S0(n5648), .S1(n5647), .A0(rptr[10]), .A1(n6110), .A2(n5944), .A3(n6222), .Z(n5910));
Q_MX02 U2511 ( .S(n5646), .A0(n5910), .A1(n5911), .Z(rptrN[10]));
Q_MX02 U2512 ( .S(n5648), .A0(n6030), .A1(n6188), .Z(n5909));
Q_MX04 U2513 ( .S0(n5648), .S1(n5647), .A0(rptr[11]), .A1(n6109), .A2(n5942), .A3(n6220), .Z(n5908));
Q_MX02 U2514 ( .S(n5646), .A0(n5908), .A1(n5909), .Z(rptrN[11]));
Q_MX02 U2515 ( .S(n5648), .A0(n6028), .A1(n6186), .Z(n5907));
Q_MX04 U2516 ( .S0(n5648), .S1(n5647), .A0(rptr[12]), .A1(n6107), .A2(n5940), .A3(n6218), .Z(n5906));
Q_MX02 U2517 ( .S(n5646), .A0(n5906), .A1(n5907), .Z(rptrN[12]));
Q_MX02 U2518 ( .S(n5648), .A0(n6026), .A1(n6184), .Z(n5905));
Q_MX04 U2519 ( .S0(n5648), .S1(n5647), .A0(rptr[13]), .A1(n6106), .A2(n5938), .A3(n6216), .Z(n5904));
Q_MX02 U2520 ( .S(n5646), .A0(n5904), .A1(n5905), .Z(rptrN[13]));
Q_MX02 U2521 ( .S(n5648), .A0(n6024), .A1(n6182), .Z(n5903));
Q_MX04 U2522 ( .S0(n5648), .S1(n5647), .A0(rptr[14]), .A1(n6104), .A2(n5936), .A3(n6214), .Z(n5902));
Q_MX02 U2523 ( .S(n5646), .A0(n5902), .A1(n5903), .Z(rptrN[14]));
Q_MX02 U2524 ( .S(n5648), .A0(n6022), .A1(n6180), .Z(n5901));
Q_MX04 U2525 ( .S0(n5648), .S1(n5647), .A0(rptr[15]), .A1(n6103), .A2(n5934), .A3(n6212), .Z(n5900));
Q_MX02 U2526 ( .S(n5646), .A0(n5900), .A1(n5901), .Z(rptrN[15]));
Q_MX02 U2527 ( .S(n5648), .A0(n6021), .A1(n6179), .Z(n6178));
Q_MX04 U2528 ( .S0(n5648), .S1(n5647), .A0(rptr[16]), .A1(n6101), .A2(n5932), .A3(n6210), .Z(n5898));
Q_MX02 U2529 ( .S(n5646), .A0(n5898), .A1(n5899), .Z(rptrN[16]));
Q_INV U2530 ( .A(rptrN[16]), .Z(n5897));
Q_AN02 U2531 ( .A0(rptr[16]), .A1(n5897), .Z(n5896));
Q_OR02 U2532 ( .A0(rptr[16]), .A1(n5897), .Z(n5895));
Q_INV U2533 ( .A(rptrN[15]), .Z(n5894));
Q_AN03 U2534 ( .A0(rptr[15]), .A1(n5894), .A2(n5895), .Z(n5886));
Q_OA21 U2535 ( .A0(rptr[15]), .A1(n5894), .B0(n5895), .Z(n5890));
Q_INV U2536 ( .A(rptrN[14]), .Z(n5893));
Q_AN02 U2537 ( .A0(rptr[14]), .A1(n5893), .Z(n5892));
Q_OA21 U2538 ( .A0(rptr[14]), .A1(n5893), .B0(n5890), .Z(n5889));
Q_INV U2539 ( .A(rptrN[13]), .Z(n5891));
Q_AN03 U2540 ( .A0(rptr[13]), .A1(n5891), .A2(n5889), .Z(n5888));
Q_OA21 U2541 ( .A0(rptr[13]), .A1(n5891), .B0(n5889), .Z(n5884));
Q_AO21 U2542 ( .A0(n5890), .A1(n5892), .B0(n5888), .Z(n5887));
Q_OR03 U2543 ( .A0(n5896), .A1(n5886), .A2(n5887), .Z(n5885));
Q_INV U2544 ( .A(rptrN[12]), .Z(n5883));
Q_AN02 U2545 ( .A0(rptr[12]), .A1(n5883), .Z(n5882));
Q_OR02 U2546 ( .A0(rptr[12]), .A1(n5883), .Z(n5881));
Q_INV U2547 ( .A(rptrN[11]), .Z(n5880));
Q_AN02 U2548 ( .A0(rptr[11]), .A1(n5880), .Z(n5879));
Q_OA21 U2549 ( .A0(rptr[11]), .A1(n5880), .B0(n5881), .Z(n5874));
Q_INV U2550 ( .A(rptrN[10]), .Z(n5878));
Q_AN02 U2551 ( .A0(rptr[10]), .A1(n5878), .Z(n5877));
Q_OA21 U2552 ( .A0(rptr[10]), .A1(n5878), .B0(n5874), .Z(n5873));
Q_INV U2553 ( .A(rptrN[9]), .Z(n5876));
Q_AN03 U2554 ( .A0(rptr[9]), .A1(n5876), .A2(n5873), .Z(n5872));
Q_OR02 U2555 ( .A0(rptr[9]), .A1(n5876), .Z(n5875));
Q_AO21 U2556 ( .A0(n5874), .A1(n5877), .B0(n5872), .Z(n5871));
Q_AO21 U2557 ( .A0(n5881), .A1(n5879), .B0(n5882), .Z(n5870));
Q_OA21 U2558 ( .A0(n5870), .A1(n5871), .B0(n5884), .Z(n5837));
Q_AN03 U2559 ( .A0(n5873), .A1(n5875), .A2(n5884), .Z(n5841));
Q_INV U2560 ( .A(rptrN[8]), .Z(n5869));
Q_AN02 U2561 ( .A0(rptr[8]), .A1(n5869), .Z(n5868));
Q_OR02 U2562 ( .A0(rptr[8]), .A1(n5869), .Z(n5867));
Q_INV U2563 ( .A(rptrN[7]), .Z(n5866));
Q_AN03 U2564 ( .A0(rptr[7]), .A1(n5866), .A2(n5867), .Z(n5857));
Q_OA21 U2565 ( .A0(rptr[7]), .A1(n5866), .B0(n5867), .Z(n5861));
Q_INV U2566 ( .A(rptrN[6]), .Z(n5865));
Q_AN02 U2567 ( .A0(rptr[6]), .A1(n5865), .Z(n5864));
Q_OA21 U2568 ( .A0(rptr[6]), .A1(n5865), .B0(n5861), .Z(n5860));
Q_INV U2569 ( .A(rptrN[5]), .Z(n5863));
Q_AN03 U2570 ( .A0(rptr[5]), .A1(n5863), .A2(n5860), .Z(n5859));
Q_OR02 U2571 ( .A0(rptr[5]), .A1(n5863), .Z(n5862));
Q_AO21 U2572 ( .A0(n5861), .A1(n5864), .B0(n5859), .Z(n5858));
Q_OR03 U2573 ( .A0(n5868), .A1(n5857), .A2(n5858), .Z(n5856));
Q_AN03 U2574 ( .A0(n5860), .A1(n5862), .A2(n5841), .Z(n5840));
Q_INV U2575 ( .A(rptrN[4]), .Z(n5855));
Q_AN02 U2576 ( .A0(rptr[4]), .A1(n5855), .Z(n5854));
Q_OR02 U2577 ( .A0(rptr[4]), .A1(n5855), .Z(n5853));
Q_AN02 U2578 ( .A0(rptr[3]), .A1(n5374), .Z(n5852));
Q_OA21 U2579 ( .A0(rptr[3]), .A1(n5374), .B0(n5853), .Z(n5848));
Q_AN02 U2580 ( .A0(rptr[2]), .A1(n5402), .Z(n5851));
Q_OA21 U2581 ( .A0(rptr[2]), .A1(n5402), .B0(n5848), .Z(n5847));
Q_INV U2582 ( .A(rptrN[1]), .Z(n5850));
Q_AN03 U2583 ( .A0(rptr[1]), .A1(n5850), .A2(n5847), .Z(n5846));
Q_OR02 U2584 ( .A0(rptr[1]), .A1(n5850), .Z(n5849));
Q_AO21 U2585 ( .A0(n5848), .A1(n5851), .B0(n5846), .Z(n5845));
Q_AO21 U2586 ( .A0(n5853), .A1(n5852), .B0(n5854), .Z(n5844));
Q_OA21 U2587 ( .A0(n5844), .A1(n5845), .B0(n5840), .Z(n5839));
Q_AN03 U2588 ( .A0(n5847), .A1(n5849), .A2(n5840), .Z(n5835));
Q_INV U2589 ( .A(rptrN[0]), .Z(n5843));
Q_AN02 U2590 ( .A0(rptr[0]), .A1(n5843), .Z(n5842));
Q_AO21 U2591 ( .A0(n5841), .A1(n5856), .B0(n5839), .Z(n5838));
Q_OR03 U2592 ( .A0(n5885), .A1(n5837), .A2(n5838), .Z(n5836));
Q_AO21 U2593 ( .A0(n5835), .A1(n5842), .B0(n5836), .Z(n5834));
Q_INV U2594 ( .A(n5834), .Z(n5641));
Q_AN02 U2595 ( .A0(n5643), .A1(odly[0]), .Z(n5833));
Q_MX03 U2596 ( .S0(n5643), .S1(n5658), .A0(n6100), .A1(head[48]), .A2(n5833), .Z(odlyN[0]));
Q_AN02 U2597 ( .A0(n5643), .A1(odly[1]), .Z(n5832));
Q_MX03 U2598 ( .S0(n5643), .S1(n5658), .A0(n6099), .A1(head[49]), .A2(n5832), .Z(odlyN[1]));
Q_AN02 U2599 ( .A0(n5643), .A1(odly[2]), .Z(n5831));
Q_MX03 U2600 ( .S0(n5643), .S1(n5658), .A0(n6097), .A1(head[50]), .A2(n5831), .Z(odlyN[2]));
Q_AN02 U2601 ( .A0(n5643), .A1(odly[3]), .Z(n5830));
Q_MX03 U2602 ( .S0(n5643), .S1(n5658), .A0(n6095), .A1(head[51]), .A2(n5830), .Z(odlyN[3]));
Q_AN02 U2603 ( .A0(n5643), .A1(odly[4]), .Z(n5829));
Q_MX03 U2604 ( .S0(n5643), .S1(n5658), .A0(n6093), .A1(head[52]), .A2(n5829), .Z(odlyN[4]));
Q_AN02 U2605 ( .A0(n5643), .A1(odly[5]), .Z(n5828));
Q_MX03 U2606 ( .S0(n5643), .S1(n5658), .A0(n6091), .A1(head[53]), .A2(n5828), .Z(odlyN[5]));
Q_AN02 U2607 ( .A0(n5643), .A1(odly[6]), .Z(n5827));
Q_MX03 U2608 ( .S0(n5643), .S1(n5658), .A0(n6089), .A1(head[54]), .A2(n5827), .Z(odlyN[6]));
Q_AN02 U2609 ( .A0(n5643), .A1(odly[7]), .Z(n5826));
Q_MX03 U2610 ( .S0(n5643), .S1(n5658), .A0(n6087), .A1(head[55]), .A2(n5826), .Z(odlyN[7]));
Q_AN02 U2611 ( .A0(n5643), .A1(odly[8]), .Z(n5825));
Q_MX03 U2612 ( .S0(n5643), .S1(n5658), .A0(n6085), .A1(head[56]), .A2(n5825), .Z(odlyN[8]));
Q_AN02 U2613 ( .A0(n5643), .A1(odly[9]), .Z(n5824));
Q_MX03 U2614 ( .S0(n5643), .S1(n5658), .A0(n6083), .A1(head[57]), .A2(n5824), .Z(odlyN[9]));
Q_AN02 U2615 ( .A0(n5643), .A1(odly[10]), .Z(n5823));
Q_MX03 U2616 ( .S0(n5643), .S1(n5658), .A0(n6081), .A1(head[58]), .A2(n5823), .Z(odlyN[10]));
Q_AN02 U2617 ( .A0(n5643), .A1(odly[11]), .Z(n5822));
Q_MX03 U2618 ( .S0(n5643), .S1(n5658), .A0(n6079), .A1(head[59]), .A2(n5822), .Z(odlyN[11]));
Q_AN02 U2619 ( .A0(eob), .A1(head[61]), .Z(rstDone));
Q_AN02 U2620 ( .A0(n5642), .A1(head[32]), .Z(n5821));
Q_MX02 U2621 ( .S(n5653), .A0(pktl[0]), .A1(n5821), .Z(n5820));
Q_AN02 U2622 ( .A0(n5642), .A1(head[33]), .Z(n5819));
Q_MX02 U2623 ( .S(n5653), .A0(pktl[1]), .A1(n5819), .Z(n5818));
Q_AN02 U2624 ( .A0(n5642), .A1(head[34]), .Z(n5817));
Q_MX02 U2625 ( .S(n5653), .A0(pktl[2]), .A1(n5817), .Z(n5816));
Q_NR02 U2626 ( .A0(n5655), .A1(head[35]), .Z(n5815));
Q_MX02 U2627 ( .S(n5653), .A0(n6177), .A1(n5815), .Z(n5814));
Q_AN02 U2628 ( .A0(n5642), .A1(n6059), .Z(n5813));
Q_MX02 U2629 ( .S(n5653), .A0(n6176), .A1(n5813), .Z(n5812));
Q_AN02 U2630 ( .A0(n5642), .A1(n6057), .Z(n5811));
Q_MX02 U2631 ( .S(n5653), .A0(n6174), .A1(n5811), .Z(n5810));
Q_AN02 U2632 ( .A0(n5642), .A1(n6055), .Z(n5809));
Q_MX02 U2633 ( .S(n5653), .A0(n6172), .A1(n5809), .Z(n5808));
Q_AN02 U2634 ( .A0(n5642), .A1(n6053), .Z(n5807));
Q_MX02 U2635 ( .S(n5653), .A0(n6170), .A1(n5807), .Z(n5806));
Q_AN02 U2636 ( .A0(n5642), .A1(n6051), .Z(n5805));
Q_MX02 U2637 ( .S(n5653), .A0(n6168), .A1(n5805), .Z(n5804));
Q_AN02 U2638 ( .A0(n5642), .A1(n6049), .Z(n5803));
Q_MX02 U2639 ( .S(n5653), .A0(n6166), .A1(n5803), .Z(n5802));
Q_MX02 U2640 ( .S(n5653), .A0(n6164), .A1(n5796), .Z(n5801));
Q_MX02 U2641 ( .S(n5653), .A0(n6162), .A1(n5796), .Z(n5800));
Q_MX02 U2642 ( .S(n5653), .A0(n6160), .A1(n5796), .Z(n5799));
Q_MX02 U2643 ( .S(n5653), .A0(n6158), .A1(n5796), .Z(n5798));
Q_MX02 U2644 ( .S(n5653), .A0(n6156), .A1(n5796), .Z(n5797));
Q_MX02 U2645 ( .S(n5653), .A0(n6154), .A1(n5796), .Z(n5795));
Q_LDP0 \pktlN_REG[15] ( .G(n5649), .D(n5795), .Q(pktlN[15]), .QN( ));
Q_LDP0 \pktlN_REG[14] ( .G(n5649), .D(n5797), .Q(pktlN[14]), .QN( ));
Q_LDP0 \pktlN_REG[13] ( .G(n5649), .D(n5798), .Q(pktlN[13]), .QN( ));
Q_LDP0 \pktlN_REG[12] ( .G(n5649), .D(n5799), .Q(pktlN[12]), .QN( ));
Q_LDP0 \pktlN_REG[11] ( .G(n5649), .D(n5800), .Q(pktlN[11]), .QN( ));
Q_LDP0 \pktlN_REG[10] ( .G(n5649), .D(n5801), .Q(pktlN[10]), .QN( ));
Q_LDP0 \pktlN_REG[9] ( .G(n5649), .D(n5802), .Q(pktlN[9]), .QN( ));
Q_LDP0 \pktlN_REG[8] ( .G(n5649), .D(n5804), .Q(pktlN[8]), .QN( ));
Q_LDP0 \pktlN_REG[7] ( .G(n5649), .D(n5806), .Q(pktlN[7]), .QN( ));
Q_LDP0 \pktlN_REG[6] ( .G(n5649), .D(n5808), .Q(pktlN[6]), .QN( ));
Q_LDP0 \pktlN_REG[5] ( .G(n5649), .D(n5810), .Q(pktlN[5]), .QN( ));
Q_LDP0 \pktlN_REG[4] ( .G(n5649), .D(n5812), .Q(pktlN[4]), .QN( ));
Q_LDP0 \pktlN_REG[3] ( .G(n5649), .D(n5814), .Q(pktlN[3]), .QN( ));
Q_LDP0 \pktlN_REG[2] ( .G(n5649), .D(n5816), .Q(pktlN[2]), .QN( ));
Q_LDP0 \pktlN_REG[1] ( .G(n5649), .D(n5818), .Q(pktlN[1]), .QN( ));
Q_LDP0 \pktlN_REG[0] ( .G(n5649), .D(n5820), .Q(pktlN[0]), .QN( ));
Q_AN02 U2662 ( .A0(n5641), .A1(rptrN[0]), .Z(n5794));
Q_AN02 U2663 ( .A0(n5641), .A1(rptrN[1]), .Z(n5793));
Q_AN02 U2664 ( .A0(n5641), .A1(rptrN[2]), .Z(n5792));
Q_AN02 U2665 ( .A0(n5641), .A1(rptrN[3]), .Z(n5791));
Q_AN02 U2666 ( .A0(n5641), .A1(rptrN[4]), .Z(n5790));
Q_AN02 U2667 ( .A0(n5641), .A1(rptrN[5]), .Z(n5789));
Q_AN02 U2668 ( .A0(n5641), .A1(rptrN[6]), .Z(n5788));
Q_AN02 U2669 ( .A0(n5641), .A1(rptrN[7]), .Z(n5787));
Q_AN02 U2670 ( .A0(n5641), .A1(rptrN[8]), .Z(n5786));
Q_AN02 U2671 ( .A0(n5641), .A1(rptrN[9]), .Z(n5785));
Q_AN02 U2672 ( .A0(n5641), .A1(rptrN[10]), .Z(n5784));
Q_AN02 U2673 ( .A0(n5641), .A1(rptrN[11]), .Z(n5783));
Q_AN02 U2674 ( .A0(n5641), .A1(rptrN[12]), .Z(n5782));
Q_AN02 U2675 ( .A0(n5641), .A1(rptrN[13]), .Z(n5781));
Q_AN02 U2676 ( .A0(n5641), .A1(rptrN[14]), .Z(n5780));
Q_AN02 U2677 ( .A0(n5641), .A1(rptrN[15]), .Z(n5779));
Q_AN02 U2678 ( .A0(n5641), .A1(rptrN[16]), .Z(n5778));
Q_INV U2679 ( .A(rptr[1]), .Z(n5777));
Q_INV U2680 ( .A(rptr[2]), .Z(n5776));
Q_INV U2681 ( .A(rptr[4]), .Z(n5775));
Q_INV U2682 ( .A(rptr[5]), .Z(n5774));
Q_INV U2683 ( .A(rptr[6]), .Z(n5773));
Q_INV U2684 ( .A(rptr[7]), .Z(n5772));
Q_INV U2685 ( .A(rptr[8]), .Z(n5771));
Q_INV U2686 ( .A(rptr[9]), .Z(n5770));
Q_INV U2687 ( .A(rptr[10]), .Z(n5769));
Q_INV U2688 ( .A(rptr[11]), .Z(n5768));
Q_INV U2689 ( .A(rptr[12]), .Z(n5767));
Q_INV U2690 ( .A(rptr[13]), .Z(n5766));
Q_INV U2691 ( .A(rptr[14]), .Z(n5765));
Q_INV U2692 ( .A(rptr[15]), .Z(n5764));
Q_INV U2693 ( .A(rptr[16]), .Z(n5763));
Q_XNR2 U2694 ( .A0(n6209), .A1(n5794), .Z(n5762));
Q_OR02 U2695 ( .A0(n6209), .A1(n5794), .Z(n5761));
Q_AD01 U2696 ( .CI(n5793), .A0(n5777), .B0(n5761), .S(n5760), .CO(n5759));
Q_AD02 U2697 ( .CI(n5759), .A0(n5776), .A1(n6235), .B0(n5792), .B1(n5791), .S0(n5758), .S1(n5757), .CO(n5756));
Q_AD02 U2698 ( .CI(n5756), .A0(n5775), .A1(n5774), .B0(n5790), .B1(n5789), .S0(n5755), .S1(n5754), .CO(n5753));
Q_AD02 U2699 ( .CI(n5753), .A0(n5773), .A1(n5772), .B0(n5788), .B1(n5787), .S0(n5752), .S1(n5751), .CO(n5750));
Q_AD02 U2700 ( .CI(n5750), .A0(n5771), .A1(n5770), .B0(n5786), .B1(n5785), .S0(n5749), .S1(n5748), .CO(n5747));
Q_AD02 U2701 ( .CI(n5747), .A0(n5769), .A1(n5768), .B0(n5784), .B1(n5783), .S0(n5746), .S1(n5745), .CO(n5744));
Q_AD02 U2702 ( .CI(n5744), .A0(n5767), .A1(n5766), .B0(n5782), .B1(n5781), .S0(n5743), .S1(n5742), .CO(n5741));
Q_AD02 U2703 ( .CI(n5741), .A0(n5765), .A1(n5764), .B0(n5780), .B1(n5779), .S0(n5740), .S1(n5739), .CO(n5738));
Q_AD01 U2704 ( .CI(n5738), .A0(n5763), .B0(n5778), .S(n5737), .CO(n5736));
Q_XNR3 U2705 ( .A0(n5834), .A1(n5736), .A2(n1), .Z(rdDelta[17]));
Q_AD01HF U2706 ( .A0(rptrN[0]), .B0(n5762), .S(n5735), .CO(n5734));
Q_AD02 U2707 ( .CI(n5760), .A0(n5734), .A1(rptrN[2]), .B0(rptrN[1]), .B1(n5758), .S0(n5733), .S1(n5732), .CO(n5731));
Q_AD02 U2708 ( .CI(n5731), .A0(rptrN[3]), .A1(rptrN[4]), .B0(n5757), .B1(n5755), .S0(n5730), .S1(n5729), .CO(n5728));
Q_AD02 U2709 ( .CI(n5728), .A0(rptrN[5]), .A1(rptrN[6]), .B0(n5754), .B1(n5752), .S0(n5727), .S1(n5726), .CO(n5725));
Q_AD02 U2710 ( .CI(n5725), .A0(rptrN[7]), .A1(rptrN[8]), .B0(n5751), .B1(n5749), .S0(n5724), .S1(n5723), .CO(n5722));
Q_AD02 U2711 ( .CI(n5722), .A0(rptrN[9]), .A1(rptrN[10]), .B0(n5748), .B1(n5746), .S0(n5721), .S1(n5720), .CO(n5719));
Q_AD02 U2712 ( .CI(n5719), .A0(rptrN[11]), .A1(rptrN[12]), .B0(n5745), .B1(n5743), .S0(n5718), .S1(n5717), .CO(n5716));
Q_AD02 U2713 ( .CI(n5716), .A0(rptrN[13]), .A1(rptrN[14]), .B0(n5742), .B1(n5740), .S0(n5715), .S1(n5714), .CO(n5713));
Q_AD02 U2714 ( .CI(n5713), .A0(rptrN[15]), .A1(rptrN[16]), .B0(n5739), .B1(n5737), .S0(n5712), .S1(n5711), .CO(n5710));
Q_MX02 U2715 ( .S(n5834), .A0(n5762), .A1(n5735), .Z(rdDelta[0]));
Q_MX02 U2716 ( .S(n5834), .A0(n5760), .A1(n5733), .Z(rdDelta[1]));
Q_MX02 U2717 ( .S(n5834), .A0(n5758), .A1(n5732), .Z(rdDelta[2]));
Q_MX02 U2718 ( .S(n5834), .A0(n5757), .A1(n5730), .Z(rdDelta[3]));
Q_MX02 U2719 ( .S(n5834), .A0(n5755), .A1(n5729), .Z(rdDelta[4]));
Q_MX02 U2720 ( .S(n5834), .A0(n5754), .A1(n5727), .Z(rdDelta[5]));
Q_MX02 U2721 ( .S(n5834), .A0(n5752), .A1(n5726), .Z(rdDelta[6]));
Q_MX02 U2722 ( .S(n5834), .A0(n5751), .A1(n5724), .Z(rdDelta[7]));
Q_MX02 U2723 ( .S(n5834), .A0(n5749), .A1(n5723), .Z(rdDelta[8]));
Q_MX02 U2724 ( .S(n5834), .A0(n5748), .A1(n5721), .Z(rdDelta[9]));
Q_MX02 U2725 ( .S(n5834), .A0(n5746), .A1(n5720), .Z(rdDelta[10]));
Q_MX02 U2726 ( .S(n5834), .A0(n5745), .A1(n5718), .Z(rdDelta[11]));
Q_MX02 U2727 ( .S(n5834), .A0(n5743), .A1(n5717), .Z(rdDelta[12]));
Q_MX02 U2728 ( .S(n5834), .A0(n5742), .A1(n5715), .Z(rdDelta[13]));
Q_MX02 U2729 ( .S(n5834), .A0(n5740), .A1(n5714), .Z(rdDelta[14]));
Q_MX02 U2730 ( .S(n5834), .A0(n5739), .A1(n5712), .Z(rdDelta[15]));
Q_MX02 U2731 ( .S(n5834), .A0(n5737), .A1(n5711), .Z(rdDelta[16]));
Q_ND03 U2732 ( .A0(n5645), .A1(n5644), .A2(n5665), .Z(n5709));
Q_MX02 U2733 ( .S(n5645), .A0(n6009), .A1(vlen[0]), .Z(n5708));
Q_AN02 U2734 ( .A0(n5645), .A1(vlen[0]), .Z(n5707));
Q_MX04 U2735 ( .S0(n5644), .S1(n5647), .A0(n5707), .A1(n6145), .A2(n5708), .A3(n5979), .Z(n5706));
Q_MX02 U2736 ( .S(n5645), .A0(n6008), .A1(vlen[1]), .Z(n5705));
Q_AN02 U2737 ( .A0(n5645), .A1(vlen[1]), .Z(n5704));
Q_MX04 U2738 ( .S0(n5644), .S1(n5647), .A0(n5704), .A1(n6143), .A2(n5705), .A3(n5977), .Z(n5703));
Q_MX02 U2739 ( .S(n5645), .A0(n6007), .A1(vlen[2]), .Z(n5702));
Q_AN02 U2740 ( .A0(n5645), .A1(vlen[2]), .Z(n5701));
Q_MX04 U2741 ( .S0(n5644), .S1(n5647), .A0(n5701), .A1(n6141), .A2(n5702), .A3(n5976), .Z(n5700));
Q_MX02 U2742 ( .S(n5645), .A0(n6006), .A1(vlen[3]), .Z(n5999));
Q_AN02 U2743 ( .A0(n5645), .A1(vlen[3]), .Z(n5698));
Q_MX04 U2744 ( .S0(n5644), .S1(n5647), .A0(n5698), .A1(n6140), .A2(n5699), .A3(n5974), .Z(n5697));
Q_MX02 U2745 ( .S(n5645), .A0(n6020), .A1(n5998), .Z(n5696));
Q_AN02 U2746 ( .A0(n5645), .A1(vlen[4]), .Z(n5695));
Q_MX04 U2747 ( .S0(n5644), .S1(n5647), .A0(n5695), .A1(n6138), .A2(n5696), .A3(n5973), .Z(n5694));
Q_MX02 U2748 ( .S(n5645), .A0(n6018), .A1(n5996), .Z(n5693));
Q_AN02 U2749 ( .A0(n5645), .A1(vlen[5]), .Z(n5692));
Q_MX04 U2750 ( .S0(n5644), .S1(n5647), .A0(n5692), .A1(n6137), .A2(n5693), .A3(n5971), .Z(n5691));
Q_MX02 U2751 ( .S(n5645), .A0(n6016), .A1(n5994), .Z(n5690));
Q_AN02 U2752 ( .A0(n5645), .A1(vlen[6]), .Z(n5689));
Q_MX04 U2753 ( .S0(n5644), .S1(n5647), .A0(n5689), .A1(n6135), .A2(n5690), .A3(n5970), .Z(n5688));
Q_MX02 U2754 ( .S(n5645), .A0(n6014), .A1(n5992), .Z(n5687));
Q_AN02 U2755 ( .A0(n5645), .A1(vlen[7]), .Z(n5686));
Q_MX04 U2756 ( .S0(n5644), .S1(n5647), .A0(n5686), .A1(n6134), .A2(n5687), .A3(n5968), .Z(n5685));
Q_MX02 U2757 ( .S(n5645), .A0(n6012), .A1(n5990), .Z(n5684));
Q_AN02 U2758 ( .A0(n5645), .A1(vlen[8]), .Z(n5683));
Q_MX04 U2759 ( .S0(n5644), .S1(n5647), .A0(n5683), .A1(n6132), .A2(n5684), .A3(n5967), .Z(n5682));
Q_MX02 U2760 ( .S(n5645), .A0(n6010), .A1(n5988), .Z(n5681));
Q_AN02 U2761 ( .A0(n5645), .A1(vlen[9]), .Z(n5680));
Q_MX04 U2762 ( .S0(n5644), .S1(n5647), .A0(n5680), .A1(n6131), .A2(n5681), .A3(n5965), .Z(n5679));
Q_LDP0 \vlenN_REG[9] ( .G(n5709), .D(n5679), .Q(vlenN[9]), .QN( ));
Q_LDP0 \vlenN_REG[8] ( .G(n5709), .D(n5682), .Q(vlenN[8]), .QN( ));
Q_LDP0 \vlenN_REG[7] ( .G(n5709), .D(n5685), .Q(vlenN[7]), .QN( ));
Q_LDP0 \vlenN_REG[6] ( .G(n5709), .D(n5688), .Q(vlenN[6]), .QN( ));
Q_LDP0 \vlenN_REG[5] ( .G(n5709), .D(n5691), .Q(vlenN[5]), .QN( ));
Q_LDP0 \vlenN_REG[4] ( .G(n5709), .D(n5694), .Q(vlenN[4]), .QN( ));
Q_LDP0 \vlenN_REG[3] ( .G(n5709), .D(n5697), .Q(vlenN[3]), .QN( ));
Q_LDP0 \vlenN_REG[2] ( .G(n5709), .D(n5700), .Q(vlenN[2]), .QN( ));
Q_LDP0 \vlenN_REG[1] ( .G(n5709), .D(n5703), .Q(vlenN[1]), .QN( ));
Q_LDP0 \vlenN_REG[0] ( .G(n5709), .D(n5706), .Q(vlenN[0]), .QN( ));
Q_AN02 U2773 ( .A0(n5636), .A1(n5678), .Z(n5648));
Q_MX02 U2774 ( .S(n5640), .A0(n6290), .A1(n5677), .Z(n5678));
Q_OR02 U2775 ( .A0(n5638), .A1(n5675), .Z(n5677));
Q_INV U2776 ( .A(n5674), .Z(n5675));
Q_AN02 U2777 ( .A0(nps), .A1(n5673), .Z(n5646));
Q_AN02 U2778 ( .A0(n5636), .A1(n5640), .Z(nps));
Q_AN02 U2779 ( .A0(n5636), .A1(n5672), .Z(n5645));
Q_MX02 U2780 ( .S(n5640), .A0(n5671), .A1(n5638), .Z(n5672));
Q_AN02 U2781 ( .A0(n5636), .A1(n5670), .Z(n5644));
Q_MX02 U2782 ( .S(n5640), .A0(n5669), .A1(n5667), .Z(n5670));
Q_INV U2783 ( .A(n5671), .Z(n5669));
Q_OR02 U2784 ( .A0(n5668), .A1(n5634), .Z(n5671));
Q_INV U2785 ( .A(n6290), .Z(n5668));
Q_OR02 U2786 ( .A0(n5638), .A1(n5666), .Z(n5667));
Q_NR02 U2787 ( .A0(n5637), .A1(n5635), .Z(n5666));
Q_INV U2788 ( .A(n5665), .Z(n5647));
Q_OR03 U2789 ( .A0(n5664), .A1(n5663), .A2(n6263), .Z(n5665));
Q_NR02 U2790 ( .A0(n5652), .A1(n5640), .Z(n5663));
Q_AN02 U2791 ( .A0(n5673), .A1(n5640), .Z(n5664));
Q_ND02 U2792 ( .A0(n6289), .A1(n6263), .Z(n5661));
Q_OA21 U2793 ( .A0(n5660), .A1(n6263), .B0(n5661), .Z(n5643));
Q_MX02 U2794 ( .S(n5640), .A0(n6290), .A1(n5659), .Z(n5660));
Q_AN02 U2795 ( .A0(n5657), .A1(n5661), .Z(n5658));
Q_OR03 U2796 ( .A0(n5664), .A1(n5656), .A2(n6263), .Z(n5657));
Q_OA21 U2797 ( .A0(n6290), .A1(n6288), .B0(n5676), .Z(n5656));
Q_OR02 U2798 ( .A0(n5638), .A1(n5637), .Z(n5673));
Q_INV U2799 ( .A(n5655), .Z(n5642));
Q_OR02 U2800 ( .A0(n284), .A1(n5674), .Z(n5655));
Q_OR02 U2801 ( .A0(n5637), .A1(n5654), .Z(n5674));
Q_INV U2802 ( .A(n5635), .Z(n5654));
Q_OR03 U2803 ( .A0(n6263), .A1(n5640), .A2(n5662), .Z(n5653));
Q_INV U2804 ( .A(n5652), .Z(n5662));
Q_AN02 U2805 ( .A0(n6290), .A1(n5634), .Z(n5652));
Q_NR02 U2806 ( .A0(n284), .A1(n5659), .Z(eob));
Q_INV U2807 ( .A(n5640), .Z(n5676));
Q_OR02 U2808 ( .A0(n5638), .A1(n5651), .Z(n5659));
Q_INV U2809 ( .A(n5637), .Z(n5651));
Q_INV U2810 ( .A(n5650), .Z(active));
Q_MX02 U2811 ( .S(n6263), .A0(xc_top.GFLock1), .A1(n5639), .Z(n5650));
Q_ND03 U2812 ( .A0(n5640), .A1(n5638), .A2(n5636), .Z(n5649));
Q_INV U2813 ( .A(ofifoAddr2[15]), .Z(n5633));
Q_INV U2814 ( .A(ofifoAddr1[15]), .Z(n5632));
Q_NR02 U2815 ( .A0(xc_top.GFReset), .A1(n5650), .Z(n5629));
Q_AN02 U2816 ( .A0(n279), .A1(newMarkBits[0]), .Z(n5628));
Q_AN02 U2817 ( .A0(n279), .A1(newMarkBits[1]), .Z(n5627));
Q_AN02 U2818 ( .A0(n279), .A1(newMarkBits[2]), .Z(n5626));
Q_AN02 U2819 ( .A0(n279), .A1(newMarkBits[3]), .Z(n5625));
Q_AN02 U2820 ( .A0(n279), .A1(markBitsN[0]), .Z(n5624));
Q_AN02 U2821 ( .A0(n279), .A1(markBitsN[1]), .Z(n5623));
Q_AN02 U2822 ( .A0(n279), .A1(markBitsN[2]), .Z(n5622));
Q_AN02 U2823 ( .A0(n279), .A1(markBitsN[3]), .Z(n5621));
Q_AN02 U2824 ( .A0(n279), .A1(xptrN[0]), .Z(n5620));
Q_AN02 U2825 ( .A0(n279), .A1(xptrN[1]), .Z(n5619));
Q_AN02 U2826 ( .A0(n279), .A1(xptrN[2]), .Z(n5618));
Q_AN02 U2827 ( .A0(n279), .A1(xptrN[3]), .Z(n5617));
Q_AN02 U2828 ( .A0(n279), .A1(xptrN[4]), .Z(n5616));
Q_AN02 U2829 ( .A0(n279), .A1(xptrN[5]), .Z(n5615));
Q_AN02 U2830 ( .A0(n279), .A1(xptrN[6]), .Z(n5614));
Q_AN02 U2831 ( .A0(n279), .A1(xptrN[7]), .Z(n5613));
Q_AN02 U2832 ( .A0(n279), .A1(xptrN[8]), .Z(n5612));
Q_AN02 U2833 ( .A0(n279), .A1(xptrN[9]), .Z(n5611));
Q_AN02 U2834 ( .A0(n279), .A1(xptrN[10]), .Z(n5610));
Q_AN02 U2835 ( .A0(n279), .A1(xptrN[11]), .Z(n5609));
Q_AN02 U2836 ( .A0(n279), .A1(xptrN[12]), .Z(n5608));
Q_AN02 U2837 ( .A0(n279), .A1(xptrN[13]), .Z(n5607));
Q_AN02 U2838 ( .A0(n279), .A1(xptrN[14]), .Z(n5606));
Q_AN02 U2839 ( .A0(n279), .A1(xptrN[15]), .Z(n5605));
Q_AN02 U2840 ( .A0(n279), .A1(xptrN[16]), .Z(n5604));
Q_AN02 U2841 ( .A0(n279), .A1(wptrN[0]), .Z(n5603));
Q_AN02 U2842 ( .A0(n279), .A1(wptrN[1]), .Z(n5602));
Q_AN02 U2843 ( .A0(n279), .A1(wptrN[2]), .Z(n5601));
Q_AN02 U2844 ( .A0(n279), .A1(wptrN[3]), .Z(n5600));
Q_AN02 U2845 ( .A0(n279), .A1(wptrN[4]), .Z(n5599));
Q_AN02 U2846 ( .A0(n279), .A1(wptrN[5]), .Z(n5598));
Q_AN02 U2847 ( .A0(n279), .A1(wptrN[6]), .Z(n5597));
Q_AN02 U2848 ( .A0(n279), .A1(wptrN[7]), .Z(n5596));
Q_AN02 U2849 ( .A0(n279), .A1(wptrN[8]), .Z(n5595));
Q_AN02 U2850 ( .A0(n279), .A1(wptrN[9]), .Z(n5594));
Q_AN02 U2851 ( .A0(n279), .A1(wptrN[10]), .Z(n5593));
Q_AN02 U2852 ( .A0(n279), .A1(wptrN[11]), .Z(n5592));
Q_AN02 U2853 ( .A0(n279), .A1(wptrN[12]), .Z(n5591));
Q_AN02 U2854 ( .A0(n279), .A1(wptrN[13]), .Z(n5590));
Q_AN02 U2855 ( .A0(n279), .A1(wptrN[14]), .Z(n5589));
Q_AN02 U2856 ( .A0(n279), .A1(wptrN[15]), .Z(n5588));
Q_AN02 U2857 ( .A0(n279), .A1(wptrN[16]), .Z(n5587));
Q_FDP0UA U2858 ( .D(n5587), .QTFCLK( ), .Q(wptr[16]));
Q_FDP0UA U2859 ( .D(n5588), .QTFCLK( ), .Q(wptr[15]));
Q_FDP0UA U2860 ( .D(n5589), .QTFCLK( ), .Q(wptr[14]));
Q_FDP0UA U2861 ( .D(n5590), .QTFCLK( ), .Q(wptr[13]));
Q_FDP0UA U2862 ( .D(n5591), .QTFCLK( ), .Q(wptr[12]));
Q_FDP0UA U2863 ( .D(n5592), .QTFCLK( ), .Q(wptr[11]));
Q_FDP0UA U2864 ( .D(n5593), .QTFCLK( ), .Q(wptr[10]));
Q_FDP0UA U2865 ( .D(n5594), .QTFCLK( ), .Q(wptr[9]));
Q_FDP0UA U2866 ( .D(n5595), .QTFCLK( ), .Q(wptr[8]));
Q_FDP0UA U2867 ( .D(n5596), .QTFCLK( ), .Q(wptr[7]));
Q_FDP0UA U2868 ( .D(n5597), .QTFCLK( ), .Q(wptr[6]));
Q_FDP0UA U2869 ( .D(n5598), .QTFCLK( ), .Q(wptr[5]));
Q_FDP0UA U2870 ( .D(n5599), .QTFCLK( ), .Q(wptr[4]));
Q_FDP0UA U2871 ( .D(n5600), .QTFCLK( ), .Q(wptr[3]));
Q_FDP0UA U2872 ( .D(n5601), .QTFCLK( ), .Q(wptr[2]));
Q_FDP0UA U2873 ( .D(n5602), .QTFCLK( ), .Q(wptr[1]));
Q_FDP0UA U2874 ( .D(n5603), .QTFCLK( ), .Q(wptr[0]));
Q_FDP0UA U2875 ( .D(n5604), .QTFCLK( ), .Q(xptr[16]));
Q_FDP0UA U2876 ( .D(n5605), .QTFCLK( ), .Q(xptr[15]));
Q_FDP0UA U2877 ( .D(n5606), .QTFCLK( ), .Q(xptr[14]));
Q_FDP0UA U2878 ( .D(n5607), .QTFCLK( ), .Q(xptr[13]));
Q_FDP0UA U2879 ( .D(n5608), .QTFCLK( ), .Q(xptr[12]));
Q_FDP0UA U2880 ( .D(n5609), .QTFCLK( ), .Q(xptr[11]));
Q_FDP0UA U2881 ( .D(n5610), .QTFCLK( ), .Q(xptr[10]));
Q_FDP0UA U2882 ( .D(n5611), .QTFCLK( ), .Q(xptr[9]));
Q_FDP0UA U2883 ( .D(n5612), .QTFCLK( ), .Q(xptr[8]));
Q_FDP0UA U2884 ( .D(n5613), .QTFCLK( ), .Q(xptr[7]));
Q_FDP0UA U2885 ( .D(n5614), .QTFCLK( ), .Q(xptr[6]));
Q_FDP0UA U2886 ( .D(n5615), .QTFCLK( ), .Q(xptr[5]));
Q_FDP0UA U2887 ( .D(n5616), .QTFCLK( ), .Q(xptr[4]));
Q_FDP0UA U2888 ( .D(n5617), .QTFCLK( ), .Q(xptr[3]));
Q_FDP0UA U2889 ( .D(n5618), .QTFCLK( ), .Q(xptr[2]));
Q_FDP0UA U2890 ( .D(n5619), .QTFCLK( ), .Q(xptr[1]));
Q_FDP0UA U2891 ( .D(n5620), .QTFCLK( ), .Q(xptr[0]));
Q_FDP0UA U2892 ( .D(n5621), .QTFCLK( ), .Q(markBits[3]));
Q_FDP0UA U2893 ( .D(n5622), .QTFCLK( ), .Q(markBits[2]));
Q_FDP0UA U2894 ( .D(n5623), .QTFCLK( ), .Q(markBits[1]));
Q_FDP0UA U2895 ( .D(n5624), .QTFCLK( ), .Q(markBits[0]));
Q_FDP0UA U2896 ( .D(n5625), .QTFCLK( ), .Q(newMarkBitsD[3]));
Q_FDP0UA U2897 ( .D(n5626), .QTFCLK( ), .Q(newMarkBitsD[2]));
Q_FDP0UA U2898 ( .D(n5627), .QTFCLK( ), .Q(newMarkBitsD[1]));
Q_FDP0UA U2899 ( .D(n5628), .QTFCLK( ), .Q(newMarkBitsD[0]));
Q_FDP0UA U2900 ( .D(n5586), .QTFCLK( ), .Q(moveForward));
Q_FDP0UA U2901 ( .D(n5629), .QTFCLK( ), .Q(activeD));
Q_AN02 U2902 ( .A0(n279), .A1(moveForwardN), .Z(n5586));
Q_AD01HF U2903 ( .A0(rdCnt[0]), .B0(rdDelta[0]), .S(n5585), .CO(n5584));
Q_AD01 U2904 ( .CI(n5584), .A0(rdCnt[1]), .B0(rdDelta[1]), .S(n5583), .CO(n5582));
Q_AD02 U2905 ( .CI(n5582), .A0(rdCnt[2]), .A1(rdCnt[3]), .B0(rdDelta[2]), .B1(rdDelta[3]), .S0(n5581), .S1(n5580), .CO(n5579));
Q_AD02 U2906 ( .CI(n5579), .A0(rdCnt[4]), .A1(rdCnt[5]), .B0(rdDelta[4]), .B1(rdDelta[5]), .S0(n5578), .S1(n5577), .CO(n5576));
Q_AD02 U2907 ( .CI(n5576), .A0(rdCnt[6]), .A1(rdCnt[7]), .B0(rdDelta[6]), .B1(rdDelta[7]), .S0(n5575), .S1(n5574), .CO(n5573));
Q_AD02 U2908 ( .CI(n5573), .A0(rdCnt[8]), .A1(rdCnt[9]), .B0(rdDelta[8]), .B1(rdDelta[9]), .S0(n5572), .S1(n5571), .CO(n5570));
Q_AD02 U2909 ( .CI(n5570), .A0(rdCnt[10]), .A1(rdCnt[11]), .B0(rdDelta[10]), .B1(rdDelta[11]), .S0(n5569), .S1(n5568), .CO(n5567));
Q_AD02 U2910 ( .CI(n5567), .A0(rdCnt[12]), .A1(rdCnt[13]), .B0(rdDelta[12]), .B1(rdDelta[13]), .S0(n5566), .S1(n5565), .CO(n5564));
Q_AD02 U2911 ( .CI(n5564), .A0(rdCnt[14]), .A1(rdCnt[15]), .B0(rdDelta[14]), .B1(rdDelta[15]), .S0(n5563), .S1(n5562), .CO(n5561));
Q_AD02 U2912 ( .CI(n5561), .A0(rdCnt[16]), .A1(rdCnt[17]), .B0(rdDelta[16]), .B1(rdDelta[17]), .S0(n5560), .S1(n5559), .CO(n5558));
Q_AD01HF U2913 ( .A0(rdCnt[18]), .B0(n5558), .S(n5557), .CO(n5556));
Q_AD01HF U2914 ( .A0(rdCnt[19]), .B0(n5556), .S(n5555), .CO(n5554));
Q_AD01HF U2915 ( .A0(rdCnt[20]), .B0(n5554), .S(n5553), .CO(n5552));
Q_AD01HF U2916 ( .A0(rdCnt[21]), .B0(n5552), .S(n5551), .CO(n5550));
Q_AD01HF U2917 ( .A0(rdCnt[22]), .B0(n5550), .S(n5549), .CO(n5548));
Q_AD01HF U2918 ( .A0(rdCnt[23]), .B0(n5548), .S(n5547), .CO(n5546));
Q_AD01HF U2919 ( .A0(rdCnt[24]), .B0(n5546), .S(n5545), .CO(n5544));
Q_AD01HF U2920 ( .A0(rdCnt[25]), .B0(n5544), .S(n5543), .CO(n5542));
Q_AD01HF U2921 ( .A0(rdCnt[26]), .B0(n5542), .S(n5541), .CO(n5540));
Q_AD01HF U2922 ( .A0(rdCnt[27]), .B0(n5540), .S(n5539), .CO(n5538));
Q_AD01HF U2923 ( .A0(rdCnt[28]), .B0(n5538), .S(n5537), .CO(n5536));
Q_AD01HF U2924 ( .A0(rdCnt[29]), .B0(n5536), .S(n5535), .CO(n5534));
Q_AD01HF U2925 ( .A0(rdCnt[30]), .B0(n5534), .S(n5533), .CO(n5532));
Q_AD01HF U2926 ( .A0(rdCnt[31]), .B0(n5532), .S(n5531), .CO(n5530));
Q_AD01HF U2927 ( .A0(rdCnt[32]), .B0(n5530), .S(n5529), .CO(n5528));
Q_AD01HF U2928 ( .A0(rdCnt[33]), .B0(n5528), .S(n5527), .CO(n5526));
Q_AD01HF U2929 ( .A0(rdCnt[34]), .B0(n5526), .S(n5525), .CO(n5524));
Q_AD01HF U2930 ( .A0(rdCnt[35]), .B0(n5524), .S(n5523), .CO(n5522));
Q_AD01HF U2931 ( .A0(rdCnt[36]), .B0(n5522), .S(n5521), .CO(n5520));
Q_AD01HF U2932 ( .A0(rdCnt[37]), .B0(n5520), .S(n5519), .CO(n5518));
Q_AD01HF U2933 ( .A0(rdCnt[38]), .B0(n5518), .S(n5517), .CO(n5516));
Q_AD01HF U2934 ( .A0(rdCnt[39]), .B0(n5516), .S(n5515), .CO(n5514));
Q_AD01HF U2935 ( .A0(rdCnt[40]), .B0(n5514), .S(n5513), .CO(n5512));
Q_AD01HF U2936 ( .A0(rdCnt[41]), .B0(n5512), .S(n5511), .CO(n5510));
Q_AD01HF U2937 ( .A0(rdCnt[42]), .B0(n5510), .S(n5509), .CO(n5508));
Q_AD01HF U2938 ( .A0(rdCnt[43]), .B0(n5508), .S(n5507), .CO(n5506));
Q_AD01HF U2939 ( .A0(rdCnt[44]), .B0(n5506), .S(n5505), .CO(n5504));
Q_AD01HF U2940 ( .A0(rdCnt[45]), .B0(n5504), .S(n5503), .CO(n5502));
Q_AD01HF U2941 ( .A0(rdCnt[46]), .B0(n5502), .S(n5501), .CO(n5500));
Q_AD01HF U2942 ( .A0(rdCnt[47]), .B0(n5500), .S(n5499), .CO(n5498));
Q_AD01HF U2943 ( .A0(rdCnt[48]), .B0(n5498), .S(n5497), .CO(n5496));
Q_AD01HF U2944 ( .A0(rdCnt[49]), .B0(n5496), .S(n5495), .CO(n5494));
Q_AD01HF U2945 ( .A0(rdCnt[50]), .B0(n5494), .S(n5493), .CO(n5492));
Q_AD01HF U2946 ( .A0(rdCnt[51]), .B0(n5492), .S(n5491), .CO(n5490));
Q_AD01HF U2947 ( .A0(rdCnt[52]), .B0(n5490), .S(n5489), .CO(n5488));
Q_AD01HF U2948 ( .A0(rdCnt[53]), .B0(n5488), .S(n5487), .CO(n5486));
Q_AD01HF U2949 ( .A0(rdCnt[54]), .B0(n5486), .S(n5485), .CO(n5484));
Q_AD01HF U2950 ( .A0(rdCnt[55]), .B0(n5484), .S(n5483), .CO(n5482));
Q_AD01HF U2951 ( .A0(rdCnt[56]), .B0(n5482), .S(n5481), .CO(n5480));
Q_AD01HF U2952 ( .A0(rdCnt[57]), .B0(n5480), .S(n5479), .CO(n5478));
Q_AD01HF U2953 ( .A0(rdCnt[58]), .B0(n5478), .S(n5477), .CO(n5476));
Q_AD01HF U2954 ( .A0(rdCnt[59]), .B0(n5476), .S(n5475), .CO(n5474));
Q_AD01HF U2955 ( .A0(rdCnt[60]), .B0(n5474), .S(n5473), .CO(n5472));
Q_AD01HF U2956 ( .A0(rdCnt[61]), .B0(n5472), .S(n5471), .CO(n5470));
Q_AD01HF U2957 ( .A0(rdCnt[62]), .B0(n5470), .S(n5469), .CO(n5468));
Q_XOR2 U2958 ( .A0(rdCnt[63]), .A1(n5468), .Z(n5467));
Q_AN02 U2959 ( .A0(n279), .A1(n5585), .Z(n5466));
Q_AN02 U2960 ( .A0(n279), .A1(n5583), .Z(n5465));
Q_AN02 U2961 ( .A0(n279), .A1(n5581), .Z(n5464));
Q_AN02 U2962 ( .A0(n279), .A1(n5580), .Z(n5463));
Q_AN02 U2963 ( .A0(n279), .A1(n5578), .Z(n5462));
Q_AN02 U2964 ( .A0(n279), .A1(n5577), .Z(n5461));
Q_AN02 U2965 ( .A0(n279), .A1(n5575), .Z(n5460));
Q_AN02 U2966 ( .A0(n279), .A1(n5574), .Z(n5459));
Q_AN02 U2967 ( .A0(n279), .A1(n5572), .Z(n5458));
Q_AN02 U2968 ( .A0(n279), .A1(n5571), .Z(n5457));
Q_AN02 U2969 ( .A0(n279), .A1(n5569), .Z(n5456));
Q_AN02 U2970 ( .A0(n279), .A1(n5568), .Z(n5455));
Q_AN02 U2971 ( .A0(n279), .A1(n5566), .Z(n5454));
Q_AN02 U2972 ( .A0(n279), .A1(n5565), .Z(n5453));
Q_AN02 U2973 ( .A0(n279), .A1(n5563), .Z(n5452));
Q_AN02 U2974 ( .A0(n279), .A1(n5562), .Z(n5451));
Q_AN02 U2975 ( .A0(n279), .A1(n5560), .Z(n5450));
Q_AN02 U2976 ( .A0(n279), .A1(n5559), .Z(n5449));
Q_AN02 U2977 ( .A0(n279), .A1(n5557), .Z(n5448));
Q_AN02 U2978 ( .A0(n279), .A1(n5555), .Z(n5447));
Q_AN02 U2979 ( .A0(n279), .A1(n5553), .Z(n5446));
Q_AN02 U2980 ( .A0(n279), .A1(n5551), .Z(n5445));
Q_AN02 U2981 ( .A0(n279), .A1(n5549), .Z(n5444));
Q_AN02 U2982 ( .A0(n279), .A1(n5547), .Z(n5443));
Q_AN02 U2983 ( .A0(n279), .A1(n5545), .Z(n5442));
Q_AN02 U2984 ( .A0(n279), .A1(n5543), .Z(n5441));
Q_AN02 U2985 ( .A0(n279), .A1(n5541), .Z(n5440));
Q_AN02 U2986 ( .A0(n279), .A1(n5539), .Z(n5439));
Q_AN02 U2987 ( .A0(n279), .A1(n5537), .Z(n5438));
Q_AN02 U2988 ( .A0(n279), .A1(n5535), .Z(n5437));
Q_AN02 U2989 ( .A0(n279), .A1(n5533), .Z(n5436));
Q_AN02 U2990 ( .A0(n279), .A1(n5531), .Z(n5435));
Q_AN02 U2991 ( .A0(n279), .A1(n5529), .Z(n5434));
Q_AN02 U2992 ( .A0(n279), .A1(n5527), .Z(n5433));
Q_AN02 U2993 ( .A0(n279), .A1(n5525), .Z(n5432));
Q_AN02 U2994 ( .A0(n279), .A1(n5523), .Z(n5431));
Q_AN02 U2995 ( .A0(n279), .A1(n5521), .Z(n5430));
Q_AN02 U2996 ( .A0(n279), .A1(n5519), .Z(n5429));
Q_AN02 U2997 ( .A0(n279), .A1(n5517), .Z(n5428));
Q_AN02 U2998 ( .A0(n279), .A1(n5515), .Z(n5427));
Q_AN02 U2999 ( .A0(n279), .A1(n5513), .Z(n5426));
Q_AN02 U3000 ( .A0(n279), .A1(n5511), .Z(n5425));
Q_AN02 U3001 ( .A0(n279), .A1(n5509), .Z(n5424));
Q_AN02 U3002 ( .A0(n279), .A1(n5507), .Z(n5423));
Q_AN02 U3003 ( .A0(n279), .A1(n5505), .Z(n5422));
Q_AN02 U3004 ( .A0(n279), .A1(n5503), .Z(n5421));
Q_AN02 U3005 ( .A0(n279), .A1(n5501), .Z(n5420));
Q_AN02 U3006 ( .A0(n279), .A1(n5499), .Z(n5419));
Q_AN02 U3007 ( .A0(n279), .A1(n5497), .Z(n5418));
Q_AN02 U3008 ( .A0(n279), .A1(n5495), .Z(n5417));
Q_AN02 U3009 ( .A0(n279), .A1(n5493), .Z(n5416));
Q_AN02 U3010 ( .A0(n279), .A1(n5491), .Z(n5415));
Q_AN02 U3011 ( .A0(n279), .A1(n5489), .Z(n5414));
Q_AN02 U3012 ( .A0(n279), .A1(n5487), .Z(n5413));
Q_AN02 U3013 ( .A0(n279), .A1(n5485), .Z(n5412));
Q_AN02 U3014 ( .A0(n279), .A1(n5483), .Z(n5411));
Q_AN02 U3015 ( .A0(n279), .A1(n5481), .Z(n5410));
Q_AN02 U3016 ( .A0(n279), .A1(n5479), .Z(n5409));
Q_AN02 U3017 ( .A0(n279), .A1(n5477), .Z(n5408));
Q_AN02 U3018 ( .A0(n279), .A1(n5475), .Z(n5407));
Q_AN02 U3019 ( .A0(n279), .A1(n5473), .Z(n5406));
Q_AN02 U3020 ( .A0(n279), .A1(n5471), .Z(n5405));
Q_AN02 U3021 ( .A0(n279), .A1(n5469), .Z(n5404));
Q_AN02 U3022 ( .A0(n279), .A1(n5467), .Z(n5403));
Q_FDP0UA U3023 ( .D(n5403), .QTFCLK( ), .Q(rdCnt[63]));
Q_FDP0UA U3024 ( .D(n5404), .QTFCLK( ), .Q(rdCnt[62]));
Q_FDP0UA U3025 ( .D(n5405), .QTFCLK( ), .Q(rdCnt[61]));
Q_FDP0UA U3026 ( .D(n5406), .QTFCLK( ), .Q(rdCnt[60]));
Q_FDP0UA U3027 ( .D(n5407), .QTFCLK( ), .Q(rdCnt[59]));
Q_FDP0UA U3028 ( .D(n5408), .QTFCLK( ), .Q(rdCnt[58]));
Q_FDP0UA U3029 ( .D(n5409), .QTFCLK( ), .Q(rdCnt[57]));
Q_FDP0UA U3030 ( .D(n5410), .QTFCLK( ), .Q(rdCnt[56]));
Q_FDP0UA U3031 ( .D(n5411), .QTFCLK( ), .Q(rdCnt[55]));
Q_FDP0UA U3032 ( .D(n5412), .QTFCLK( ), .Q(rdCnt[54]));
Q_FDP0UA U3033 ( .D(n5413), .QTFCLK( ), .Q(rdCnt[53]));
Q_FDP0UA U3034 ( .D(n5414), .QTFCLK( ), .Q(rdCnt[52]));
Q_FDP0UA U3035 ( .D(n5415), .QTFCLK( ), .Q(rdCnt[51]));
Q_FDP0UA U3036 ( .D(n5416), .QTFCLK( ), .Q(rdCnt[50]));
Q_FDP0UA U3037 ( .D(n5417), .QTFCLK( ), .Q(rdCnt[49]));
Q_FDP0UA U3038 ( .D(n5418), .QTFCLK( ), .Q(rdCnt[48]));
Q_FDP0UA U3039 ( .D(n5419), .QTFCLK( ), .Q(rdCnt[47]));
Q_FDP0UA U3040 ( .D(n5420), .QTFCLK( ), .Q(rdCnt[46]));
Q_FDP0UA U3041 ( .D(n5421), .QTFCLK( ), .Q(rdCnt[45]));
Q_FDP0UA U3042 ( .D(n5422), .QTFCLK( ), .Q(rdCnt[44]));
Q_FDP0UA U3043 ( .D(n5423), .QTFCLK( ), .Q(rdCnt[43]));
Q_FDP0UA U3044 ( .D(n5424), .QTFCLK( ), .Q(rdCnt[42]));
Q_FDP0UA U3045 ( .D(n5425), .QTFCLK( ), .Q(rdCnt[41]));
Q_FDP0UA U3046 ( .D(n5426), .QTFCLK( ), .Q(rdCnt[40]));
Q_FDP0UA U3047 ( .D(n5427), .QTFCLK( ), .Q(rdCnt[39]));
Q_FDP0UA U3048 ( .D(n5428), .QTFCLK( ), .Q(rdCnt[38]));
Q_FDP0UA U3049 ( .D(n5429), .QTFCLK( ), .Q(rdCnt[37]));
Q_FDP0UA U3050 ( .D(n5430), .QTFCLK( ), .Q(rdCnt[36]));
Q_FDP0UA U3051 ( .D(n5431), .QTFCLK( ), .Q(rdCnt[35]));
Q_FDP0UA U3052 ( .D(n5432), .QTFCLK( ), .Q(rdCnt[34]));
Q_FDP0UA U3053 ( .D(n5433), .QTFCLK( ), .Q(rdCnt[33]));
Q_FDP0UA U3054 ( .D(n5434), .QTFCLK( ), .Q(rdCnt[32]));
Q_FDP0UA U3055 ( .D(n5435), .QTFCLK( ), .Q(rdCnt[31]));
Q_FDP0UA U3056 ( .D(n5436), .QTFCLK( ), .Q(rdCnt[30]));
Q_FDP0UA U3057 ( .D(n5437), .QTFCLK( ), .Q(rdCnt[29]));
Q_FDP0UA U3058 ( .D(n5438), .QTFCLK( ), .Q(rdCnt[28]));
Q_FDP0UA U3059 ( .D(n5439), .QTFCLK( ), .Q(rdCnt[27]));
Q_FDP0UA U3060 ( .D(n5440), .QTFCLK( ), .Q(rdCnt[26]));
Q_FDP0UA U3061 ( .D(n5441), .QTFCLK( ), .Q(rdCnt[25]));
Q_FDP0UA U3062 ( .D(n5442), .QTFCLK( ), .Q(rdCnt[24]));
Q_FDP0UA U3063 ( .D(n5443), .QTFCLK( ), .Q(rdCnt[23]));
Q_FDP0UA U3064 ( .D(n5444), .QTFCLK( ), .Q(rdCnt[22]));
Q_FDP0UA U3065 ( .D(n5445), .QTFCLK( ), .Q(rdCnt[21]));
Q_FDP0UA U3066 ( .D(n5446), .QTFCLK( ), .Q(rdCnt[20]));
Q_FDP0UA U3067 ( .D(n5447), .QTFCLK( ), .Q(rdCnt[19]));
Q_FDP0UA U3068 ( .D(n5448), .QTFCLK( ), .Q(rdCnt[18]));
Q_FDP0UA U3069 ( .D(n5449), .QTFCLK( ), .Q(rdCnt[17]));
Q_FDP0UA U3070 ( .D(n5450), .QTFCLK( ), .Q(rdCnt[16]));
Q_FDP0UA U3071 ( .D(n5451), .QTFCLK( ), .Q(rdCnt[15]));
Q_FDP0UA U3072 ( .D(n5452), .QTFCLK( ), .Q(rdCnt[14]));
Q_FDP0UA U3073 ( .D(n5453), .QTFCLK( ), .Q(rdCnt[13]));
Q_FDP0UA U3074 ( .D(n5454), .QTFCLK( ), .Q(rdCnt[12]));
Q_FDP0UA U3075 ( .D(n5455), .QTFCLK( ), .Q(rdCnt[11]));
Q_FDP0UA U3076 ( .D(n5456), .QTFCLK( ), .Q(rdCnt[10]));
Q_FDP0UA U3077 ( .D(n5457), .QTFCLK( ), .Q(rdCnt[9]));
Q_FDP0UA U3078 ( .D(n5458), .QTFCLK( ), .Q(rdCnt[8]));
Q_FDP0UA U3079 ( .D(n5459), .QTFCLK( ), .Q(rdCnt[7]));
Q_FDP0UA U3080 ( .D(n5460), .QTFCLK( ), .Q(rdCnt[6]));
Q_FDP0UA U3081 ( .D(n5461), .QTFCLK( ), .Q(rdCnt[5]));
Q_FDP0UA U3082 ( .D(n5462), .QTFCLK( ), .Q(rdCnt[4]));
Q_FDP0UA U3083 ( .D(n5463), .QTFCLK( ), .Q(rdCnt[3]));
Q_FDP0UA U3084 ( .D(n5464), .QTFCLK( ), .Q(rdCnt[2]));
Q_FDP0UA U3085 ( .D(n5465), .QTFCLK( ), .Q(rdCnt[1]));
Q_FDP0UA U3086 ( .D(n5466), .QTFCLK( ), .Q(rdCnt[0]));
Q_INV U3087 ( .A(rptrN[2]), .Z(n5402));
Q_AD01HF U3088 ( .A0(rptrN[3]), .B0(rptrN[2]), .S(n5401), .CO(n5400));
Q_AD01HF U3089 ( .A0(rptrN[4]), .B0(n5400), .S(n5399), .CO(n5398));
Q_AD01HF U3090 ( .A0(rptrN[5]), .B0(n5398), .S(n5397), .CO(n5396));
Q_AD01HF U3091 ( .A0(rptrN[6]), .B0(n5396), .S(n5395), .CO(n5394));
Q_AD01HF U3092 ( .A0(rptrN[7]), .B0(n5394), .S(n5393), .CO(n5392));
Q_AD01HF U3093 ( .A0(rptrN[8]), .B0(n5392), .S(n5391), .CO(n5390));
Q_AD01HF U3094 ( .A0(rptrN[9]), .B0(n5390), .S(n5389), .CO(n5388));
Q_AD01HF U3095 ( .A0(rptrN[10]), .B0(n5388), .S(n5387), .CO(n5386));
Q_AD01HF U3096 ( .A0(rptrN[11]), .B0(n5386), .S(n5385), .CO(n5384));
Q_AD01HF U3097 ( .A0(rptrN[12]), .B0(n5384), .S(n5383), .CO(n5382));
Q_AD01HF U3098 ( .A0(rptrN[13]), .B0(n5382), .S(n5381), .CO(n5380));
Q_AD01HF U3099 ( .A0(rptrN[14]), .B0(n5380), .S(n5379), .CO(n5378));
Q_AD01HF U3100 ( .A0(rptrN[15]), .B0(n5378), .S(n5377), .CO(n5376));
Q_XOR2 U3101 ( .A0(rptrN[16]), .A1(n5376), .Z(n5375));
Q_INV U3102 ( .A(rptrN[3]), .Z(n5374));
Q_AD01HF U3103 ( .A0(rptrN[4]), .B0(rptrN[3]), .S(n5373), .CO(n5372));
Q_AD01HF U3104 ( .A0(rptrN[5]), .B0(n5372), .S(n5371), .CO(n5370));
Q_AD01HF U3105 ( .A0(rptrN[6]), .B0(n5370), .S(n5369), .CO(n5368));
Q_AD01HF U3106 ( .A0(rptrN[7]), .B0(n5368), .S(n5367), .CO(n5366));
Q_AD01HF U3107 ( .A0(rptrN[8]), .B0(n5366), .S(n5365), .CO(n5364));
Q_AD01HF U3108 ( .A0(rptrN[9]), .B0(n5364), .S(n5363), .CO(n5362));
Q_AD01HF U3109 ( .A0(rptrN[10]), .B0(n5362), .S(n5361), .CO(n5360));
Q_AD01HF U3110 ( .A0(rptrN[11]), .B0(n5360), .S(n5359), .CO(n5358));
Q_AD01HF U3111 ( .A0(rptrN[12]), .B0(n5358), .S(n5357), .CO(n5356));
Q_AD01HF U3112 ( .A0(rptrN[13]), .B0(n5356), .S(n5355), .CO(n5354));
Q_AD01HF U3113 ( .A0(rptrN[14]), .B0(n5354), .S(n5353), .CO(n5352));
Q_AD01HF U3114 ( .A0(rptrN[15]), .B0(n5352), .S(n5351), .CO(n5350));
Q_XOR2 U3115 ( .A0(rptrN[16]), .A1(n5350), .Z(n5349));
Q_AN02 U3116 ( .A0(n279), .A1(odlyN[0]), .Z(n5348));
Q_AN02 U3117 ( .A0(n279), .A1(odlyN[1]), .Z(n5347));
Q_AN02 U3118 ( .A0(n279), .A1(odlyN[2]), .Z(n5346));
Q_AN02 U3119 ( .A0(n279), .A1(odlyN[3]), .Z(n5345));
Q_AN02 U3120 ( .A0(n279), .A1(odlyN[4]), .Z(n5344));
Q_AN02 U3121 ( .A0(n279), .A1(odlyN[5]), .Z(n5343));
Q_AN02 U3122 ( .A0(n279), .A1(odlyN[6]), .Z(n5342));
Q_AN02 U3123 ( .A0(n279), .A1(odlyN[7]), .Z(n5341));
Q_AN02 U3124 ( .A0(n279), .A1(odlyN[8]), .Z(n5340));
Q_AN02 U3125 ( .A0(n279), .A1(odlyN[9]), .Z(n5339));
Q_AN02 U3126 ( .A0(n279), .A1(odlyN[10]), .Z(n5338));
Q_AN02 U3127 ( .A0(n279), .A1(odlyN[11]), .Z(n5337));
Q_AN02 U3128 ( .A0(n279), .A1(vlenN[0]), .Z(n5336));
Q_AN02 U3129 ( .A0(n279), .A1(vlenN[1]), .Z(n5335));
Q_AN02 U3130 ( .A0(n279), .A1(vlenN[2]), .Z(n5334));
Q_AN02 U3131 ( .A0(n279), .A1(vlenN[3]), .Z(n5333));
Q_AN02 U3132 ( .A0(n279), .A1(vlenN[4]), .Z(n5332));
Q_AN02 U3133 ( .A0(n279), .A1(vlenN[5]), .Z(n5331));
Q_AN02 U3134 ( .A0(n279), .A1(vlenN[6]), .Z(n5330));
Q_AN02 U3135 ( .A0(n279), .A1(vlenN[7]), .Z(n5329));
Q_AN02 U3136 ( .A0(n279), .A1(vlenN[8]), .Z(n5328));
Q_AN02 U3137 ( .A0(n279), .A1(vlenN[9]), .Z(n5327));
Q_AN02 U3138 ( .A0(n279), .A1(pktlN[0]), .Z(n5326));
Q_AN02 U3139 ( .A0(n279), .A1(pktlN[1]), .Z(n5325));
Q_AN02 U3140 ( .A0(n279), .A1(pktlN[2]), .Z(n5324));
Q_AN02 U3141 ( .A0(n279), .A1(pktlN[3]), .Z(n5323));
Q_AN02 U3142 ( .A0(n279), .A1(pktlN[4]), .Z(n5322));
Q_AN02 U3143 ( .A0(n279), .A1(pktlN[5]), .Z(n5321));
Q_AN02 U3144 ( .A0(n279), .A1(pktlN[6]), .Z(n5320));
Q_AN02 U3145 ( .A0(n279), .A1(pktlN[7]), .Z(n5319));
Q_AN02 U3146 ( .A0(n279), .A1(pktlN[8]), .Z(n5318));
Q_AN02 U3147 ( .A0(n279), .A1(pktlN[9]), .Z(n5317));
Q_AN02 U3148 ( .A0(n279), .A1(pktlN[10]), .Z(n5316));
Q_AN02 U3149 ( .A0(n279), .A1(pktlN[11]), .Z(n5315));
Q_AN02 U3150 ( .A0(n279), .A1(pktlN[12]), .Z(n5314));
Q_AN02 U3151 ( .A0(n279), .A1(pktlN[13]), .Z(n5313));
Q_AN02 U3152 ( .A0(n279), .A1(pktlN[14]), .Z(n5312));
Q_AN02 U3153 ( .A0(n279), .A1(pktlN[15]), .Z(n5311));
Q_AN02 U3154 ( .A0(n279), .A1(head[0]), .Z(n5310));
Q_AN02 U3155 ( .A0(n279), .A1(head[1]), .Z(n5309));
Q_AN02 U3156 ( .A0(n279), .A1(head[2]), .Z(n5308));
Q_AN02 U3157 ( .A0(n279), .A1(head[3]), .Z(n5307));
Q_AN02 U3158 ( .A0(n279), .A1(head[4]), .Z(n5306));
Q_AN02 U3159 ( .A0(n279), .A1(head[5]), .Z(n5305));
Q_AN02 U3160 ( .A0(n279), .A1(head[6]), .Z(n5304));
Q_AN02 U3161 ( .A0(n279), .A1(head[7]), .Z(n5303));
Q_AN02 U3162 ( .A0(n279), .A1(head[8]), .Z(n5302));
Q_AN02 U3163 ( .A0(n279), .A1(head[9]), .Z(n5301));
Q_AN02 U3164 ( .A0(n279), .A1(head[10]), .Z(n5300));
Q_AN02 U3165 ( .A0(n279), .A1(head[11]), .Z(n5299));
Q_AN02 U3166 ( .A0(n279), .A1(head[12]), .Z(n5298));
Q_AN02 U3167 ( .A0(n279), .A1(head[13]), .Z(n5297));
Q_AN02 U3168 ( .A0(n279), .A1(head[14]), .Z(n5296));
Q_AN02 U3169 ( .A0(n279), .A1(head[15]), .Z(n5295));
Q_AN02 U3170 ( .A0(n279), .A1(head[16]), .Z(n5294));
Q_AN02 U3171 ( .A0(n279), .A1(head[17]), .Z(n5293));
Q_AN02 U3172 ( .A0(n279), .A1(head[18]), .Z(n5292));
Q_AN02 U3173 ( .A0(n279), .A1(head[19]), .Z(n5291));
Q_AN02 U3174 ( .A0(n279), .A1(head[20]), .Z(n5290));
Q_AN02 U3175 ( .A0(n279), .A1(head[21]), .Z(n5289));
Q_AN02 U3176 ( .A0(n279), .A1(head[22]), .Z(n5288));
Q_AN02 U3177 ( .A0(n279), .A1(head[23]), .Z(n5287));
Q_AN02 U3178 ( .A0(n279), .A1(head[24]), .Z(n5286));
Q_AN02 U3179 ( .A0(n279), .A1(head[25]), .Z(n5285));
Q_AN02 U3180 ( .A0(n279), .A1(head[26]), .Z(n5284));
Q_AN02 U3181 ( .A0(n279), .A1(head[27]), .Z(n5283));
Q_AN02 U3182 ( .A0(n279), .A1(head[28]), .Z(n5282));
Q_AN02 U3183 ( .A0(n279), .A1(head[29]), .Z(n5281));
Q_AN02 U3184 ( .A0(n279), .A1(head[30]), .Z(n5280));
Q_AN02 U3185 ( .A0(n279), .A1(head[31]), .Z(n5279));
Q_AN02 U3186 ( .A0(n279), .A1(head[32]), .Z(n5278));
Q_AN02 U3187 ( .A0(n279), .A1(head[33]), .Z(n5277));
Q_AN02 U3188 ( .A0(n279), .A1(head[34]), .Z(n5276));
Q_AN02 U3189 ( .A0(n279), .A1(head[35]), .Z(n5275));
Q_AN02 U3190 ( .A0(n279), .A1(head[36]), .Z(n5274));
Q_AN02 U3191 ( .A0(n279), .A1(head[37]), .Z(n5273));
Q_AN02 U3192 ( .A0(n279), .A1(head[38]), .Z(n5272));
Q_AN02 U3193 ( .A0(n279), .A1(head[39]), .Z(n5271));
Q_AN02 U3194 ( .A0(n279), .A1(head[40]), .Z(n5270));
Q_AN02 U3195 ( .A0(n279), .A1(head[41]), .Z(n5269));
Q_AN02 U3196 ( .A0(n279), .A1(head[42]), .Z(n5268));
Q_AN02 U3197 ( .A0(n279), .A1(head[43]), .Z(n5267));
Q_AN02 U3198 ( .A0(n279), .A1(head[44]), .Z(n5266));
Q_AN02 U3199 ( .A0(n279), .A1(head[45]), .Z(n5265));
Q_AN02 U3200 ( .A0(n279), .A1(head[46]), .Z(n5264));
Q_AN02 U3201 ( .A0(n279), .A1(head[47]), .Z(n5263));
Q_AN02 U3202 ( .A0(n279), .A1(head[48]), .Z(n5262));
Q_AN02 U3203 ( .A0(n279), .A1(head[49]), .Z(n5261));
Q_AN02 U3204 ( .A0(n279), .A1(head[50]), .Z(n5260));
Q_AN02 U3205 ( .A0(n279), .A1(head[51]), .Z(n5259));
Q_AN02 U3206 ( .A0(n279), .A1(head[52]), .Z(n5258));
Q_AN02 U3207 ( .A0(n279), .A1(head[53]), .Z(n5257));
Q_AN02 U3208 ( .A0(n279), .A1(head[54]), .Z(n5256));
Q_AN02 U3209 ( .A0(n279), .A1(head[55]), .Z(n5255));
Q_AN02 U3210 ( .A0(n279), .A1(head[56]), .Z(n5254));
Q_AN02 U3211 ( .A0(n279), .A1(head[57]), .Z(n5253));
Q_AN02 U3212 ( .A0(n279), .A1(head[58]), .Z(n5252));
Q_AN02 U3213 ( .A0(n279), .A1(head[59]), .Z(n5251));
Q_AN02 U3214 ( .A0(n279), .A1(head[60]), .Z(n5250));
Q_AN02 U3215 ( .A0(n279), .A1(head[61]), .Z(n5249));
Q_AN02 U3216 ( .A0(n279), .A1(head[62]), .Z(n5248));
Q_AN02 U3217 ( .A0(n279), .A1(head[63]), .Z(n5247));
Q_AN02 U3218 ( .A0(n279), .A1(n5373), .Z(n5246));
Q_AN02 U3219 ( .A0(n279), .A1(n5371), .Z(n5245));
Q_AN02 U3220 ( .A0(n279), .A1(n5369), .Z(n5244));
Q_AN02 U3221 ( .A0(n279), .A1(n5367), .Z(n5243));
Q_AN02 U3222 ( .A0(n279), .A1(n5365), .Z(n5242));
Q_AN02 U3223 ( .A0(n279), .A1(n5363), .Z(n5241));
Q_AN02 U3224 ( .A0(n279), .A1(n5361), .Z(n5240));
Q_AN02 U3225 ( .A0(n279), .A1(n5359), .Z(n5239));
Q_AN02 U3226 ( .A0(n279), .A1(n5357), .Z(n5238));
Q_AN02 U3227 ( .A0(n279), .A1(n5355), .Z(n5237));
Q_AN02 U3228 ( .A0(n279), .A1(n5353), .Z(n5236));
Q_AN02 U3229 ( .A0(n279), .A1(n5351), .Z(n5235));
Q_AN02 U3230 ( .A0(n279), .A1(n5349), .Z(n5234));
Q_AN02 U3231 ( .A0(n279), .A1(n5401), .Z(n5233));
Q_AN02 U3232 ( .A0(n279), .A1(n5399), .Z(n5232));
Q_AN02 U3233 ( .A0(n279), .A1(n5397), .Z(n5231));
Q_AN02 U3234 ( .A0(n279), .A1(n5395), .Z(n5230));
Q_AN02 U3235 ( .A0(n279), .A1(n5393), .Z(n5229));
Q_AN02 U3236 ( .A0(n279), .A1(n5391), .Z(n5228));
Q_AN02 U3237 ( .A0(n279), .A1(n5389), .Z(n5227));
Q_AN02 U3238 ( .A0(n279), .A1(n5387), .Z(n5226));
Q_AN02 U3239 ( .A0(n279), .A1(n5385), .Z(n5225));
Q_AN02 U3240 ( .A0(n279), .A1(n5383), .Z(n5224));
Q_AN02 U3241 ( .A0(n279), .A1(n5381), .Z(n5223));
Q_AN02 U3242 ( .A0(n279), .A1(n5379), .Z(n5222));
Q_AN02 U3243 ( .A0(n279), .A1(n5377), .Z(n5221));
Q_AN02 U3244 ( .A0(n279), .A1(n5375), .Z(n5220));
Q_AN02 U3245 ( .A0(n279), .A1(rptrN[0]), .Z(n5219));
Q_AN02 U3246 ( .A0(n279), .A1(rptrN[1]), .Z(n5218));
Q_AN02 U3247 ( .A0(n279), .A1(rptrN[2]), .Z(n5217));
Q_AN02 U3248 ( .A0(n279), .A1(rptrN[3]), .Z(n5216));
Q_AN02 U3249 ( .A0(n279), .A1(rptrN[4]), .Z(n5215));
Q_AN02 U3250 ( .A0(n279), .A1(rptrN[5]), .Z(n5214));
Q_AN02 U3251 ( .A0(n279), .A1(rptrN[6]), .Z(n5213));
Q_AN02 U3252 ( .A0(n279), .A1(rptrN[7]), .Z(n5212));
Q_AN02 U3253 ( .A0(n279), .A1(rptrN[8]), .Z(n5211));
Q_AN02 U3254 ( .A0(n279), .A1(rptrN[9]), .Z(n5210));
Q_AN02 U3255 ( .A0(n279), .A1(rptrN[10]), .Z(n5209));
Q_AN02 U3256 ( .A0(n279), .A1(rptrN[11]), .Z(n5208));
Q_AN02 U3257 ( .A0(n279), .A1(rptrN[12]), .Z(n5207));
Q_AN02 U3258 ( .A0(n279), .A1(rptrN[13]), .Z(n5206));
Q_AN02 U3259 ( .A0(n279), .A1(rptrN[14]), .Z(n5205));
Q_AN02 U3260 ( .A0(n279), .A1(rptrN[15]), .Z(n5204));
Q_AN02 U3261 ( .A0(n279), .A1(rptrN[16]), .Z(n5203));
Q_FDP0UA U3262 ( .D(n5203), .QTFCLK( ), .Q(rptr[16]));
Q_FDP0UA U3263 ( .D(n5204), .QTFCLK( ), .Q(rptr[15]));
Q_FDP0UA U3264 ( .D(n5205), .QTFCLK( ), .Q(rptr[14]));
Q_FDP0UA U3265 ( .D(n5206), .QTFCLK( ), .Q(rptr[13]));
Q_FDP0UA U3266 ( .D(n5207), .QTFCLK( ), .Q(rptr[12]));
Q_FDP0UA U3267 ( .D(n5208), .QTFCLK( ), .Q(rptr[11]));
Q_FDP0UA U3268 ( .D(n5209), .QTFCLK( ), .Q(rptr[10]));
Q_FDP0UA U3269 ( .D(n5210), .QTFCLK( ), .Q(rptr[9]));
Q_FDP0UA U3270 ( .D(n5211), .QTFCLK( ), .Q(rptr[8]));
Q_FDP0UA U3271 ( .D(n5212), .QTFCLK( ), .Q(rptr[7]));
Q_FDP0UA U3272 ( .D(n5213), .QTFCLK( ), .Q(rptr[6]));
Q_FDP0UA U3273 ( .D(n5214), .QTFCLK( ), .Q(rptr[5]));
Q_FDP0UA U3274 ( .D(n5215), .QTFCLK( ), .Q(rptr[4]));
Q_FDP0UA U3275 ( .D(n5216), .QTFCLK( ), .Q(rptr[3]));
Q_FDP0UA U3276 ( .D(n5217), .QTFCLK( ), .Q(rptr[2]));
Q_FDP0UA U3277 ( .D(n5218), .QTFCLK( ), .Q(rptr[1]));
Q_FDP0UA U3278 ( .D(n5219), .QTFCLK( ), .Q(rptr[0]));
Q_FDP0UA U3279 ( .D(n5203), .QTFCLK( ), .Q(ififoRaddr0[14]));
Q_FDP0UA U3280 ( .D(n5204), .QTFCLK( ), .Q(ififoRaddr0[13]));
Q_FDP0UA U3281 ( .D(n5205), .QTFCLK( ), .Q(ififoRaddr0[12]));
Q_FDP0UA U3282 ( .D(n5206), .QTFCLK( ), .Q(ififoRaddr0[11]));
Q_FDP0UA U3283 ( .D(n5207), .QTFCLK( ), .Q(ififoRaddr0[10]));
Q_FDP0UA U3284 ( .D(n5208), .QTFCLK( ), .Q(ififoRaddr0[9]));
Q_FDP0UA U3285 ( .D(n5209), .QTFCLK( ), .Q(ififoRaddr0[8]));
Q_FDP0UA U3286 ( .D(n5210), .QTFCLK( ), .Q(ififoRaddr0[7]));
Q_FDP0UA U3287 ( .D(n5211), .QTFCLK( ), .Q(ififoRaddr0[6]));
Q_FDP0UA U3288 ( .D(n5212), .QTFCLK( ), .Q(ififoRaddr0[5]));
Q_FDP0UA U3289 ( .D(n5213), .QTFCLK( ), .Q(ififoRaddr0[4]));
Q_FDP0UA U3290 ( .D(n5214), .QTFCLK( ), .Q(ififoRaddr0[3]));
Q_FDP0UA U3291 ( .D(n5215), .QTFCLK( ), .Q(ififoRaddr0[2]));
Q_FDP0UA U3292 ( .D(n5216), .QTFCLK( ), .Q(ififoRaddr0[1]));
Q_FDP0UA U3293 ( .D(n5217), .QTFCLK( ), .Q(ififoRaddr0[0]));
Q_FDP0UA U3294 ( .D(n5220), .QTFCLK( ), .Q(ififoRaddr1[14]));
Q_FDP0UA U3295 ( .D(n5221), .QTFCLK( ), .Q(ififoRaddr1[13]));
Q_FDP0UA U3296 ( .D(n5222), .QTFCLK( ), .Q(ififoRaddr1[12]));
Q_FDP0UA U3297 ( .D(n5223), .QTFCLK( ), .Q(ififoRaddr1[11]));
Q_FDP0UA U3298 ( .D(n5224), .QTFCLK( ), .Q(ififoRaddr1[10]));
Q_FDP0UA U3299 ( .D(n5225), .QTFCLK( ), .Q(ififoRaddr1[9]));
Q_FDP0UA U3300 ( .D(n5226), .QTFCLK( ), .Q(ififoRaddr1[8]));
Q_FDP0UA U3301 ( .D(n5227), .QTFCLK( ), .Q(ififoRaddr1[7]));
Q_FDP0UA U3302 ( .D(n5228), .QTFCLK( ), .Q(ififoRaddr1[6]));
Q_FDP0UA U3303 ( .D(n5229), .QTFCLK( ), .Q(ififoRaddr1[5]));
Q_FDP0UA U3304 ( .D(n5230), .QTFCLK( ), .Q(ififoRaddr1[4]));
Q_FDP0UA U3305 ( .D(n5231), .QTFCLK( ), .Q(ififoRaddr1[3]));
Q_FDP0UA U3306 ( .D(n5232), .QTFCLK( ), .Q(ififoRaddr1[2]));
Q_FDP0UA U3307 ( .D(n5233), .QTFCLK( ), .Q(ififoRaddr1[1]));
Q_FDP0UA U3308 ( .D(n6885), .QTFCLK( ), .Q(ififoRaddr1[0]));
Q_FDP0UA U3309 ( .D(n5234), .QTFCLK( ), .Q(ififoRaddr2[14]));
Q_FDP0UA U3310 ( .D(n5235), .QTFCLK( ), .Q(ififoRaddr2[13]));
Q_FDP0UA U3311 ( .D(n5236), .QTFCLK( ), .Q(ififoRaddr2[12]));
Q_FDP0UA U3312 ( .D(n5237), .QTFCLK( ), .Q(ififoRaddr2[11]));
Q_FDP0UA U3313 ( .D(n5238), .QTFCLK( ), .Q(ififoRaddr2[10]));
Q_FDP0UA U3314 ( .D(n5239), .QTFCLK( ), .Q(ififoRaddr2[9]));
Q_FDP0UA U3315 ( .D(n5240), .QTFCLK( ), .Q(ififoRaddr2[8]));
Q_FDP0UA U3316 ( .D(n5241), .QTFCLK( ), .Q(ififoRaddr2[7]));
Q_FDP0UA U3317 ( .D(n5242), .QTFCLK( ), .Q(ififoRaddr2[6]));
Q_FDP0UA U3318 ( .D(n5243), .QTFCLK( ), .Q(ififoRaddr2[5]));
Q_FDP0UA U3319 ( .D(n5244), .QTFCLK( ), .Q(ififoRaddr2[4]));
Q_FDP0UA U3320 ( .D(n5245), .QTFCLK( ), .Q(ififoRaddr2[3]));
Q_FDP0UA U3321 ( .D(n5246), .QTFCLK( ), .Q(ififoRaddr2[2]));
Q_FDP0UA U3322 ( .D(n6886), .QTFCLK( ), .Q(ififoRaddr2[1]));
Q_FDP0UA U3323 ( .D(n5217), .QTFCLK( ), .Q(ififoRaddr2[0]));
Q_FDP0UA U3324 ( .D(n5247), .QTFCLK( ), .Q(vhead[63]));
Q_FDP0UA U3325 ( .D(n5248), .QTFCLK( ), .Q(vhead[62]));
Q_FDP0UA U3326 ( .D(n5249), .QTFCLK( ), .Q(vhead[61]));
Q_FDP0UA U3327 ( .D(n5250), .QTFCLK( ), .Q(vhead[60]));
Q_FDP0UA U3328 ( .D(n5251), .QTFCLK( ), .Q(vhead[59]));
Q_FDP0UA U3329 ( .D(n5252), .QTFCLK( ), .Q(vhead[58]));
Q_FDP0UA U3330 ( .D(n5253), .QTFCLK( ), .Q(vhead[57]));
Q_FDP0UA U3331 ( .D(n5254), .QTFCLK( ), .Q(vhead[56]));
Q_FDP0UA U3332 ( .D(n5255), .QTFCLK( ), .Q(vhead[55]));
Q_FDP0UA U3333 ( .D(n5256), .QTFCLK( ), .Q(vhead[54]));
Q_FDP0UA U3334 ( .D(n5257), .QTFCLK( ), .Q(vhead[53]));
Q_FDP0UA U3335 ( .D(n5258), .QTFCLK( ), .Q(vhead[52]));
Q_FDP0UA U3336 ( .D(n5259), .QTFCLK( ), .Q(vhead[51]));
Q_FDP0UA U3337 ( .D(n5260), .QTFCLK( ), .Q(vhead[50]));
Q_FDP0UA U3338 ( .D(n5261), .QTFCLK( ), .Q(vhead[49]));
Q_FDP0UA U3339 ( .D(n5262), .QTFCLK( ), .Q(vhead[48]));
Q_FDP0UA U3340 ( .D(n5263), .QTFCLK( ), .Q(vhead[47]));
Q_FDP0UA U3341 ( .D(n5264), .QTFCLK( ), .Q(vhead[46]));
Q_FDP0UA U3342 ( .D(n5265), .QTFCLK( ), .Q(vhead[45]));
Q_FDP0UA U3343 ( .D(n5266), .QTFCLK( ), .Q(vhead[44]));
Q_FDP0UA U3344 ( .D(n5267), .QTFCLK( ), .Q(vhead[43]));
Q_FDP0UA U3345 ( .D(n5268), .QTFCLK( ), .Q(vhead[42]));
Q_FDP0UA U3346 ( .D(n5269), .QTFCLK( ), .Q(vhead[41]));
Q_FDP0UA U3347 ( .D(n5270), .QTFCLK( ), .Q(vhead[40]));
Q_FDP0UA U3348 ( .D(n5271), .QTFCLK( ), .Q(vhead[39]));
Q_FDP0UA U3349 ( .D(n5272), .QTFCLK( ), .Q(vhead[38]));
Q_FDP0UA U3350 ( .D(n5273), .QTFCLK( ), .Q(vhead[37]));
Q_FDP0UA U3351 ( .D(n5274), .QTFCLK( ), .Q(vhead[36]));
Q_FDP0UA U3352 ( .D(n5275), .QTFCLK( ), .Q(vhead[35]));
Q_FDP0UA U3353 ( .D(n5276), .QTFCLK( ), .Q(vhead[34]));
Q_FDP0UA U3354 ( .D(n5277), .QTFCLK( ), .Q(vhead[33]));
Q_FDP0UA U3355 ( .D(n5278), .QTFCLK( ), .Q(vhead[32]));
Q_FDP0UA U3356 ( .D(n5279), .QTFCLK( ), .Q(vhead[31]));
Q_FDP0UA U3357 ( .D(n5280), .QTFCLK( ), .Q(vhead[30]));
Q_FDP0UA U3358 ( .D(n5281), .QTFCLK( ), .Q(vhead[29]));
Q_FDP0UA U3359 ( .D(n5282), .QTFCLK( ), .Q(vhead[28]));
Q_FDP0UA U3360 ( .D(n5283), .QTFCLK( ), .Q(vhead[27]));
Q_FDP0UA U3361 ( .D(n5284), .QTFCLK( ), .Q(vhead[26]));
Q_FDP0UA U3362 ( .D(n5285), .QTFCLK( ), .Q(vhead[25]));
Q_FDP0UA U3363 ( .D(n5286), .QTFCLK( ), .Q(vhead[24]));
Q_FDP0UA U3364 ( .D(n5287), .QTFCLK( ), .Q(vhead[23]));
Q_FDP0UA U3365 ( .D(n5288), .QTFCLK( ), .Q(vhead[22]));
Q_FDP0UA U3366 ( .D(n5289), .QTFCLK( ), .Q(vhead[21]));
Q_FDP0UA U3367 ( .D(n5290), .QTFCLK( ), .Q(vhead[20]));
Q_FDP0UA U3368 ( .D(n5291), .QTFCLK( ), .Q(vhead[19]));
Q_FDP0UA U3369 ( .D(n5292), .QTFCLK( ), .Q(vhead[18]));
Q_FDP0UA U3370 ( .D(n5293), .QTFCLK( ), .Q(vhead[17]));
Q_FDP0UA U3371 ( .D(n5294), .QTFCLK( ), .Q(vhead[16]));
Q_FDP0UA U3372 ( .D(n5295), .QTFCLK( ), .Q(vhead[15]));
Q_FDP0UA U3373 ( .D(n5296), .QTFCLK( ), .Q(vhead[14]));
Q_FDP0UA U3374 ( .D(n5297), .QTFCLK( ), .Q(vhead[13]));
Q_FDP0UA U3375 ( .D(n5298), .QTFCLK( ), .Q(vhead[12]));
Q_FDP0UA U3376 ( .D(n5299), .QTFCLK( ), .Q(vhead[11]));
Q_FDP0UA U3377 ( .D(n5300), .QTFCLK( ), .Q(vhead[10]));
Q_FDP0UA U3378 ( .D(n5301), .QTFCLK( ), .Q(vhead[9]));
Q_FDP0UA U3379 ( .D(n5302), .QTFCLK( ), .Q(vhead[8]));
Q_FDP0UA U3380 ( .D(n5303), .QTFCLK( ), .Q(vhead[7]));
Q_FDP0UA U3381 ( .D(n5304), .QTFCLK( ), .Q(vhead[6]));
Q_FDP0UA U3382 ( .D(n5305), .QTFCLK( ), .Q(vhead[5]));
Q_FDP0UA U3383 ( .D(n5306), .QTFCLK( ), .Q(vhead[4]));
Q_FDP0UA U3384 ( .D(n5307), .QTFCLK( ), .Q(vhead[3]));
Q_FDP0UA U3385 ( .D(n5308), .QTFCLK( ), .Q(vhead[2]));
Q_FDP0UA U3386 ( .D(n5309), .QTFCLK( ), .Q(vhead[1]));
Q_FDP0UA U3387 ( .D(n5310), .QTFCLK( ), .Q(vhead[0]));
Q_FDP0UA U3388 ( .D(n5311), .QTFCLK( ), .Q(pktl[15]));
Q_FDP0UA U3389 ( .D(n5312), .QTFCLK( ), .Q(pktl[14]));
Q_FDP0UA U3390 ( .D(n5313), .QTFCLK( ), .Q(pktl[13]));
Q_FDP0UA U3391 ( .D(n5314), .QTFCLK( ), .Q(pktl[12]));
Q_FDP0UA U3392 ( .D(n5315), .QTFCLK( ), .Q(pktl[11]));
Q_FDP0UA U3393 ( .D(n5316), .QTFCLK( ), .Q(pktl[10]));
Q_FDP0UA U3394 ( .D(n5317), .QTFCLK( ), .Q(pktl[9]));
Q_FDP0UA U3395 ( .D(n5318), .QTFCLK( ), .Q(pktl[8]));
Q_FDP0UA U3396 ( .D(n5319), .QTFCLK( ), .Q(pktl[7]));
Q_FDP0UA U3397 ( .D(n5320), .QTFCLK( ), .Q(pktl[6]));
Q_FDP0UA U3398 ( .D(n5321), .QTFCLK( ), .Q(pktl[5]));
Q_FDP0UA U3399 ( .D(n5322), .QTFCLK( ), .Q(pktl[4]));
Q_FDP0UA U3400 ( .D(n5323), .QTFCLK( ), .Q(pktl[3]));
Q_FDP0UA U3401 ( .D(n5324), .QTFCLK( ), .Q(pktl[2]));
Q_FDP0UA U3402 ( .D(n5325), .QTFCLK( ), .Q(pktl[1]));
Q_FDP0UA U3403 ( .D(n5326), .QTFCLK( ), .Q(pktl[0]));
Q_FDP0UA U3404 ( .D(n5327), .QTFCLK( ), .Q(vlen[9]));
Q_FDP0UA U3405 ( .D(n5328), .QTFCLK( ), .Q(vlen[8]));
Q_FDP0UA U3406 ( .D(n5329), .QTFCLK( ), .Q(vlen[7]));
Q_FDP0UA U3407 ( .D(n5330), .QTFCLK( ), .Q(vlen[6]));
Q_FDP0UA U3408 ( .D(n5331), .QTFCLK( ), .Q(vlen[5]));
Q_FDP0UA U3409 ( .D(n5332), .QTFCLK( ), .Q(vlen[4]));
Q_FDP0UA U3410 ( .D(n5333), .QTFCLK( ), .Q(vlen[3]));
Q_FDP0UA U3411 ( .D(n5334), .QTFCLK( ), .Q(vlen[2]));
Q_FDP0UA U3412 ( .D(n5335), .QTFCLK( ), .Q(vlen[1]));
Q_FDP0UA U3413 ( .D(n5336), .QTFCLK( ), .Q(vlen[0]));
Q_FDP0UA U3414 ( .D(n5337), .QTFCLK( ), .Q(odly[11]));
Q_FDP0UA U3415 ( .D(n5338), .QTFCLK( ), .Q(odly[10]));
Q_FDP0UA U3416 ( .D(n5339), .QTFCLK( ), .Q(odly[9]));
Q_FDP0UA U3417 ( .D(n5340), .QTFCLK( ), .Q(odly[8]));
Q_FDP0UA U3418 ( .D(n5341), .QTFCLK( ), .Q(odly[7]));
Q_FDP0UA U3419 ( .D(n5342), .QTFCLK( ), .Q(odly[6]));
Q_FDP0UA U3420 ( .D(n5343), .QTFCLK( ), .Q(odly[5]));
Q_FDP0UA U3421 ( .D(n5344), .QTFCLK( ), .Q(odly[4]));
Q_FDP0UA U3422 ( .D(n5345), .QTFCLK( ), .Q(odly[3]));
Q_FDP0UA U3423 ( .D(n5346), .QTFCLK( ), .Q(odly[2]));
Q_FDP0UA U3424 ( .D(n5347), .QTFCLK( ), .Q(odly[1]));
Q_FDP0UA U3425 ( .D(n5348), .QTFCLK( ), .Q(odly[0]));
Q_AN02 U3426 ( .A0(n279), .A1(rstDoneD), .Z(n5202));
Q_AN02 U3427 ( .A0(n279), .A1(rstDone), .Z(n5201));
Q_FDP0UA U3428 ( .D(n5201), .QTFCLK( ), .Q(rstDoneD));
Q_FDP0UA U3429 ( .D(n5202), .QTFCLK( ), .Q(rstDoneD2));
Q_FDP0UA U3430 ( .D(n5200), .QTFCLK( ), .Q(oMark[254]));
Q_AN02 U3431 ( .A0(n279), .A1(oMark[254]), .Z(n5200));
Q_FDP0UA U3432 ( .D(n5199), .QTFCLK( ), .Q(oMark[253]));
Q_AN02 U3433 ( .A0(n279), .A1(oMark[253]), .Z(n5199));
Q_FDP0UA U3434 ( .D(n5198), .QTFCLK( ), .Q(oMark[252]));
Q_AN02 U3435 ( .A0(n279), .A1(oMark[252]), .Z(n5198));
Q_FDP0UA U3436 ( .D(n5197), .QTFCLK( ), .Q(oMark[251]));
Q_AN02 U3437 ( .A0(n279), .A1(oMark[251]), .Z(n5197));
Q_FDP0UA U3438 ( .D(n5196), .QTFCLK( ), .Q(oMark[250]));
Q_AN02 U3439 ( .A0(n279), .A1(oMark[250]), .Z(n5196));
Q_FDP0UA U3440 ( .D(n5195), .QTFCLK( ), .Q(oMark[249]));
Q_AN02 U3441 ( .A0(n279), .A1(oMark[249]), .Z(n5195));
Q_FDP0UA U3442 ( .D(n5194), .QTFCLK( ), .Q(oMark[248]));
Q_AN02 U3443 ( .A0(n279), .A1(oMark[248]), .Z(n5194));
Q_FDP0UA U3444 ( .D(n5193), .QTFCLK( ), .Q(oMark[247]));
Q_AN02 U3445 ( .A0(n279), .A1(oMark[247]), .Z(n5193));
Q_FDP0UA U3446 ( .D(n5192), .QTFCLK( ), .Q(oMark[246]));
Q_AN02 U3447 ( .A0(n279), .A1(oMark[246]), .Z(n5192));
Q_FDP0UA U3448 ( .D(n5191), .QTFCLK( ), .Q(oMark[245]));
Q_AN02 U3449 ( .A0(n279), .A1(oMark[245]), .Z(n5191));
Q_FDP0UA U3450 ( .D(n5190), .QTFCLK( ), .Q(oMark[244]));
Q_AN02 U3451 ( .A0(n279), .A1(oMark[244]), .Z(n5190));
Q_FDP0UA U3452 ( .D(n5189), .QTFCLK( ), .Q(oMark[243]));
Q_AN02 U3453 ( .A0(n279), .A1(oMark[243]), .Z(n5189));
Q_FDP0UA U3454 ( .D(n5188), .QTFCLK( ), .Q(oMark[242]));
Q_AN02 U3455 ( .A0(n279), .A1(oMark[242]), .Z(n5188));
Q_FDP0UA U3456 ( .D(n5187), .QTFCLK( ), .Q(oMark[241]));
Q_AN02 U3457 ( .A0(n279), .A1(oMark[241]), .Z(n5187));
Q_FDP0UA U3458 ( .D(n5186), .QTFCLK( ), .Q(oMark[240]));
Q_AN02 U3459 ( .A0(n279), .A1(oMark[240]), .Z(n5186));
Q_FDP0UA U3460 ( .D(n5185), .QTFCLK( ), .Q(oMark[239]));
Q_AN02 U3461 ( .A0(n279), .A1(oMark[239]), .Z(n5185));
Q_FDP0UA U3462 ( .D(n5184), .QTFCLK( ), .Q(oMark[238]));
Q_AN02 U3463 ( .A0(n279), .A1(oMark[238]), .Z(n5184));
Q_FDP0UA U3464 ( .D(n5183), .QTFCLK( ), .Q(oMark[237]));
Q_AN02 U3465 ( .A0(n279), .A1(oMark[237]), .Z(n5183));
Q_FDP0UA U3466 ( .D(n5182), .QTFCLK( ), .Q(oMark[236]));
Q_AN02 U3467 ( .A0(n279), .A1(oMark[236]), .Z(n5182));
Q_FDP0UA U3468 ( .D(n5181), .QTFCLK( ), .Q(oMark[235]));
Q_AN02 U3469 ( .A0(n279), .A1(oMark[235]), .Z(n5181));
Q_FDP0UA U3470 ( .D(n5180), .QTFCLK( ), .Q(oMark[234]));
Q_AN02 U3471 ( .A0(n279), .A1(oMark[234]), .Z(n5180));
Q_FDP0UA U3472 ( .D(n5179), .QTFCLK( ), .Q(oMark[233]));
Q_AN02 U3473 ( .A0(n279), .A1(oMark[233]), .Z(n5179));
Q_FDP0UA U3474 ( .D(n5178), .QTFCLK( ), .Q(oMark[232]));
Q_AN02 U3475 ( .A0(n279), .A1(oMark[232]), .Z(n5178));
Q_FDP0UA U3476 ( .D(n5177), .QTFCLK( ), .Q(oMark[231]));
Q_AN02 U3477 ( .A0(n279), .A1(oMark[231]), .Z(n5177));
Q_FDP0UA U3478 ( .D(n5176), .QTFCLK( ), .Q(oMark[230]));
Q_AN02 U3479 ( .A0(n279), .A1(oMark[230]), .Z(n5176));
Q_FDP0UA U3480 ( .D(n5175), .QTFCLK( ), .Q(oMark[229]));
Q_AN02 U3481 ( .A0(n279), .A1(oMark[229]), .Z(n5175));
Q_FDP0UA U3482 ( .D(n5174), .QTFCLK( ), .Q(oMark[228]));
Q_AN02 U3483 ( .A0(n279), .A1(oMark[228]), .Z(n5174));
Q_FDP0UA U3484 ( .D(n5173), .QTFCLK( ), .Q(oMark[227]));
Q_AN02 U3485 ( .A0(n279), .A1(oMark[227]), .Z(n5173));
Q_FDP0UA U3486 ( .D(n5172), .QTFCLK( ), .Q(oMark[226]));
Q_AN02 U3487 ( .A0(n279), .A1(oMark[226]), .Z(n5172));
Q_FDP0UA U3488 ( .D(n5171), .QTFCLK( ), .Q(oMark[225]));
Q_AN02 U3489 ( .A0(n279), .A1(oMark[225]), .Z(n5171));
Q_FDP0UA U3490 ( .D(n5170), .QTFCLK( ), .Q(oMark[224]));
Q_AN02 U3491 ( .A0(n279), .A1(oMark[224]), .Z(n5170));
Q_FDP0UA U3492 ( .D(n5169), .QTFCLK( ), .Q(oMark[223]));
Q_AN02 U3493 ( .A0(n279), .A1(oMark[223]), .Z(n5169));
Q_FDP0UA U3494 ( .D(n5168), .QTFCLK( ), .Q(oMark[222]));
Q_AN02 U3495 ( .A0(n279), .A1(oMark[222]), .Z(n5168));
Q_FDP0UA U3496 ( .D(n5167), .QTFCLK( ), .Q(oMark[221]));
Q_AN02 U3497 ( .A0(n279), .A1(oMark[221]), .Z(n5167));
Q_FDP0UA U3498 ( .D(n5166), .QTFCLK( ), .Q(oMark[220]));
Q_AN02 U3499 ( .A0(n279), .A1(oMark[220]), .Z(n5166));
Q_FDP0UA U3500 ( .D(n5165), .QTFCLK( ), .Q(oMark[219]));
Q_AN02 U3501 ( .A0(n279), .A1(oMark[219]), .Z(n5165));
Q_FDP0UA U3502 ( .D(n5164), .QTFCLK( ), .Q(oMark[218]));
Q_AN02 U3503 ( .A0(n279), .A1(oMark[218]), .Z(n5164));
Q_FDP0UA U3504 ( .D(n5163), .QTFCLK( ), .Q(oMark[217]));
Q_AN02 U3505 ( .A0(n279), .A1(oMark[217]), .Z(n5163));
Q_FDP0UA U3506 ( .D(n5162), .QTFCLK( ), .Q(oMark[216]));
Q_AN02 U3507 ( .A0(n279), .A1(oMark[216]), .Z(n5162));
Q_FDP0UA U3508 ( .D(n5161), .QTFCLK( ), .Q(oMark[215]));
Q_AN02 U3509 ( .A0(n279), .A1(oMark[215]), .Z(n5161));
Q_FDP0UA U3510 ( .D(n5160), .QTFCLK( ), .Q(oMark[214]));
Q_AN02 U3511 ( .A0(n279), .A1(oMark[214]), .Z(n5160));
Q_FDP0UA U3512 ( .D(n5159), .QTFCLK( ), .Q(oMark[213]));
Q_AN02 U3513 ( .A0(n279), .A1(oMark[213]), .Z(n5159));
Q_FDP0UA U3514 ( .D(n5158), .QTFCLK( ), .Q(oMark[212]));
Q_AN02 U3515 ( .A0(n279), .A1(oMark[212]), .Z(n5158));
Q_FDP0UA U3516 ( .D(n5157), .QTFCLK( ), .Q(oMark[211]));
Q_AN02 U3517 ( .A0(n279), .A1(oMark[211]), .Z(n5157));
Q_FDP0UA U3518 ( .D(n5156), .QTFCLK( ), .Q(oMark[210]));
Q_AN02 U3519 ( .A0(n279), .A1(oMark[210]), .Z(n5156));
Q_FDP0UA U3520 ( .D(n5155), .QTFCLK( ), .Q(oMark[209]));
Q_AN02 U3521 ( .A0(n279), .A1(oMark[209]), .Z(n5155));
Q_FDP0UA U3522 ( .D(n5154), .QTFCLK( ), .Q(oMark[208]));
Q_AN02 U3523 ( .A0(n279), .A1(oMark[208]), .Z(n5154));
Q_FDP0UA U3524 ( .D(n5153), .QTFCLK( ), .Q(oMark[207]));
Q_AN02 U3525 ( .A0(n279), .A1(oMark[207]), .Z(n5153));
Q_FDP0UA U3526 ( .D(n5152), .QTFCLK( ), .Q(oMark[206]));
Q_AN02 U3527 ( .A0(n279), .A1(oMark[206]), .Z(n5152));
Q_FDP0UA U3528 ( .D(n5151), .QTFCLK( ), .Q(oMark[205]));
Q_AN02 U3529 ( .A0(n279), .A1(oMark[205]), .Z(n5151));
Q_FDP0UA U3530 ( .D(n5150), .QTFCLK( ), .Q(oMark[204]));
Q_AN02 U3531 ( .A0(n279), .A1(oMark[204]), .Z(n5150));
Q_FDP0UA U3532 ( .D(n5149), .QTFCLK( ), .Q(oMark[203]));
Q_AN02 U3533 ( .A0(n279), .A1(oMark[203]), .Z(n5149));
Q_FDP0UA U3534 ( .D(n5148), .QTFCLK( ), .Q(oMark[202]));
Q_AN02 U3535 ( .A0(n279), .A1(oMark[202]), .Z(n5148));
Q_FDP0UA U3536 ( .D(n5147), .QTFCLK( ), .Q(oMark[201]));
Q_AN02 U3537 ( .A0(n279), .A1(oMark[201]), .Z(n5147));
Q_FDP0UA U3538 ( .D(n5146), .QTFCLK( ), .Q(oMark[200]));
Q_AN02 U3539 ( .A0(n279), .A1(oMark[200]), .Z(n5146));
Q_FDP0UA U3540 ( .D(n5145), .QTFCLK( ), .Q(oMark[199]));
Q_AN02 U3541 ( .A0(n279), .A1(oMark[199]), .Z(n5145));
Q_FDP0UA U3542 ( .D(n5144), .QTFCLK( ), .Q(oMark[198]));
Q_AN02 U3543 ( .A0(n279), .A1(oMark[198]), .Z(n5144));
Q_FDP0UA U3544 ( .D(n5143), .QTFCLK( ), .Q(oMark[197]));
Q_AN02 U3545 ( .A0(n279), .A1(oMark[197]), .Z(n5143));
Q_FDP0UA U3546 ( .D(n5142), .QTFCLK( ), .Q(oMark[196]));
Q_AN02 U3547 ( .A0(n279), .A1(oMark[196]), .Z(n5142));
Q_FDP0UA U3548 ( .D(n5141), .QTFCLK( ), .Q(oMark[195]));
Q_AN02 U3549 ( .A0(n279), .A1(oMark[195]), .Z(n5141));
Q_FDP0UA U3550 ( .D(n5140), .QTFCLK( ), .Q(oMark[194]));
Q_AN02 U3551 ( .A0(n279), .A1(oMark[194]), .Z(n5140));
Q_FDP0UA U3552 ( .D(n5139), .QTFCLK( ), .Q(oMark[193]));
Q_AN02 U3553 ( .A0(n279), .A1(oMark[193]), .Z(n5139));
Q_FDP0UA U3554 ( .D(n5138), .QTFCLK( ), .Q(oMark[192]));
Q_AN02 U3555 ( .A0(n279), .A1(oMark[192]), .Z(n5138));
Q_FDP0UA U3556 ( .D(n5137), .QTFCLK( ), .Q(oMark[190]));
Q_AN02 U3557 ( .A0(n279), .A1(oMark[190]), .Z(n5137));
Q_FDP0UA U3558 ( .D(n5136), .QTFCLK( ), .Q(oMark[189]));
Q_AN02 U3559 ( .A0(n279), .A1(oMark[189]), .Z(n5136));
Q_FDP0UA U3560 ( .D(n5135), .QTFCLK( ), .Q(oMark[188]));
Q_AN02 U3561 ( .A0(n279), .A1(oMark[188]), .Z(n5135));
Q_FDP0UA U3562 ( .D(n5134), .QTFCLK( ), .Q(oMark[187]));
Q_AN02 U3563 ( .A0(n279), .A1(oMark[187]), .Z(n5134));
Q_FDP0UA U3564 ( .D(n5133), .QTFCLK( ), .Q(oMark[186]));
Q_AN02 U3565 ( .A0(n279), .A1(oMark[186]), .Z(n5133));
Q_FDP0UA U3566 ( .D(n5132), .QTFCLK( ), .Q(oMark[185]));
Q_AN02 U3567 ( .A0(n279), .A1(oMark[185]), .Z(n5132));
Q_FDP0UA U3568 ( .D(n5131), .QTFCLK( ), .Q(oMark[184]));
Q_AN02 U3569 ( .A0(n279), .A1(oMark[184]), .Z(n5131));
Q_FDP0UA U3570 ( .D(n5130), .QTFCLK( ), .Q(oMark[183]));
Q_AN02 U3571 ( .A0(n279), .A1(oMark[183]), .Z(n5130));
Q_FDP0UA U3572 ( .D(n5129), .QTFCLK( ), .Q(oMark[182]));
Q_AN02 U3573 ( .A0(n279), .A1(oMark[182]), .Z(n5129));
Q_FDP0UA U3574 ( .D(n5128), .QTFCLK( ), .Q(oMark[181]));
Q_AN02 U3575 ( .A0(n279), .A1(oMark[181]), .Z(n5128));
Q_FDP0UA U3576 ( .D(n5127), .QTFCLK( ), .Q(oMark[180]));
Q_AN02 U3577 ( .A0(n279), .A1(oMark[180]), .Z(n5127));
Q_FDP0UA U3578 ( .D(n5126), .QTFCLK( ), .Q(oMark[179]));
Q_AN02 U3579 ( .A0(n279), .A1(oMark[179]), .Z(n5126));
Q_FDP0UA U3580 ( .D(n5125), .QTFCLK( ), .Q(oMark[178]));
Q_AN02 U3581 ( .A0(n279), .A1(oMark[178]), .Z(n5125));
Q_FDP0UA U3582 ( .D(n5124), .QTFCLK( ), .Q(oMark[177]));
Q_AN02 U3583 ( .A0(n279), .A1(oMark[177]), .Z(n5124));
Q_FDP0UA U3584 ( .D(n5123), .QTFCLK( ), .Q(oMark[176]));
Q_AN02 U3585 ( .A0(n279), .A1(oMark[176]), .Z(n5123));
Q_FDP0UA U3586 ( .D(n5122), .QTFCLK( ), .Q(oMark[175]));
Q_AN02 U3587 ( .A0(n279), .A1(oMark[175]), .Z(n5122));
Q_FDP0UA U3588 ( .D(n5121), .QTFCLK( ), .Q(oMark[174]));
Q_AN02 U3589 ( .A0(n279), .A1(oMark[174]), .Z(n5121));
Q_FDP0UA U3590 ( .D(n5120), .QTFCLK( ), .Q(oMark[173]));
Q_AN02 U3591 ( .A0(n279), .A1(oMark[173]), .Z(n5120));
Q_FDP0UA U3592 ( .D(n5119), .QTFCLK( ), .Q(oMark[172]));
Q_AN02 U3593 ( .A0(n279), .A1(oMark[172]), .Z(n5119));
Q_FDP0UA U3594 ( .D(n5118), .QTFCLK( ), .Q(oMark[171]));
Q_AN02 U3595 ( .A0(n279), .A1(oMark[171]), .Z(n5118));
Q_FDP0UA U3596 ( .D(n5117), .QTFCLK( ), .Q(oMark[170]));
Q_AN02 U3597 ( .A0(n279), .A1(oMark[170]), .Z(n5117));
Q_FDP0UA U3598 ( .D(n5116), .QTFCLK( ), .Q(oMark[169]));
Q_AN02 U3599 ( .A0(n279), .A1(oMark[169]), .Z(n5116));
Q_FDP0UA U3600 ( .D(n5115), .QTFCLK( ), .Q(oMark[168]));
Q_AN02 U3601 ( .A0(n279), .A1(oMark[168]), .Z(n5115));
Q_FDP0UA U3602 ( .D(n5114), .QTFCLK( ), .Q(oMark[167]));
Q_AN02 U3603 ( .A0(n279), .A1(oMark[167]), .Z(n5114));
Q_FDP0UA U3604 ( .D(n5113), .QTFCLK( ), .Q(oMark[166]));
Q_AN02 U3605 ( .A0(n279), .A1(oMark[166]), .Z(n5113));
Q_FDP0UA U3606 ( .D(n5112), .QTFCLK( ), .Q(oMark[165]));
Q_AN02 U3607 ( .A0(n279), .A1(oMark[165]), .Z(n5112));
Q_FDP0UA U3608 ( .D(n5111), .QTFCLK( ), .Q(oMark[164]));
Q_AN02 U3609 ( .A0(n279), .A1(oMark[164]), .Z(n5111));
Q_FDP0UA U3610 ( .D(n5110), .QTFCLK( ), .Q(oMark[163]));
Q_AN02 U3611 ( .A0(n279), .A1(oMark[163]), .Z(n5110));
Q_FDP0UA U3612 ( .D(n5109), .QTFCLK( ), .Q(oMark[162]));
Q_AN02 U3613 ( .A0(n279), .A1(oMark[162]), .Z(n5109));
Q_FDP0UA U3614 ( .D(n5108), .QTFCLK( ), .Q(oMark[161]));
Q_AN02 U3615 ( .A0(n279), .A1(oMark[161]), .Z(n5108));
Q_FDP0UA U3616 ( .D(n5107), .QTFCLK( ), .Q(oMark[160]));
Q_AN02 U3617 ( .A0(n279), .A1(oMark[160]), .Z(n5107));
Q_FDP0UA U3618 ( .D(n5106), .QTFCLK( ), .Q(oMark[159]));
Q_AN02 U3619 ( .A0(n279), .A1(oMark[159]), .Z(n5106));
Q_FDP0UA U3620 ( .D(n5105), .QTFCLK( ), .Q(oMark[158]));
Q_AN02 U3621 ( .A0(n279), .A1(oMark[158]), .Z(n5105));
Q_FDP0UA U3622 ( .D(n5104), .QTFCLK( ), .Q(oMark[157]));
Q_AN02 U3623 ( .A0(n279), .A1(oMark[157]), .Z(n5104));
Q_FDP0UA U3624 ( .D(n5103), .QTFCLK( ), .Q(oMark[156]));
Q_AN02 U3625 ( .A0(n279), .A1(oMark[156]), .Z(n5103));
Q_FDP0UA U3626 ( .D(n5102), .QTFCLK( ), .Q(oMark[155]));
Q_AN02 U3627 ( .A0(n279), .A1(oMark[155]), .Z(n5102));
Q_FDP0UA U3628 ( .D(n5101), .QTFCLK( ), .Q(oMark[154]));
Q_AN02 U3629 ( .A0(n279), .A1(oMark[154]), .Z(n5101));
Q_FDP0UA U3630 ( .D(n5100), .QTFCLK( ), .Q(oMark[153]));
Q_AN02 U3631 ( .A0(n279), .A1(oMark[153]), .Z(n5100));
Q_FDP0UA U3632 ( .D(n5099), .QTFCLK( ), .Q(oMark[152]));
Q_AN02 U3633 ( .A0(n279), .A1(oMark[152]), .Z(n5099));
Q_FDP0UA U3634 ( .D(n5098), .QTFCLK( ), .Q(oMark[151]));
Q_AN02 U3635 ( .A0(n279), .A1(oMark[151]), .Z(n5098));
Q_FDP0UA U3636 ( .D(n5097), .QTFCLK( ), .Q(oMark[150]));
Q_AN02 U3637 ( .A0(n279), .A1(oMark[150]), .Z(n5097));
Q_FDP0UA U3638 ( .D(n5096), .QTFCLK( ), .Q(oMark[149]));
Q_AN02 U3639 ( .A0(n279), .A1(oMark[149]), .Z(n5096));
Q_FDP0UA U3640 ( .D(n5095), .QTFCLK( ), .Q(oMark[148]));
Q_AN02 U3641 ( .A0(n279), .A1(oMark[148]), .Z(n5095));
Q_FDP0UA U3642 ( .D(n5094), .QTFCLK( ), .Q(oMark[147]));
Q_AN02 U3643 ( .A0(n279), .A1(oMark[147]), .Z(n5094));
Q_FDP0UA U3644 ( .D(n5093), .QTFCLK( ), .Q(oMark[146]));
Q_AN02 U3645 ( .A0(n279), .A1(oMark[146]), .Z(n5093));
Q_FDP0UA U3646 ( .D(n5092), .QTFCLK( ), .Q(oMark[145]));
Q_AN02 U3647 ( .A0(n279), .A1(oMark[145]), .Z(n5092));
Q_FDP0UA U3648 ( .D(n5091), .QTFCLK( ), .Q(oMark[144]));
Q_AN02 U3649 ( .A0(n279), .A1(oMark[144]), .Z(n5091));
Q_FDP0UA U3650 ( .D(n5090), .QTFCLK( ), .Q(oMark[143]));
Q_AN02 U3651 ( .A0(n279), .A1(oMark[143]), .Z(n5090));
Q_FDP0UA U3652 ( .D(n5089), .QTFCLK( ), .Q(oMark[142]));
Q_AN02 U3653 ( .A0(n279), .A1(oMark[142]), .Z(n5089));
Q_FDP0UA U3654 ( .D(n5088), .QTFCLK( ), .Q(oMark[141]));
Q_AN02 U3655 ( .A0(n279), .A1(oMark[141]), .Z(n5088));
Q_FDP0UA U3656 ( .D(n5087), .QTFCLK( ), .Q(oMark[140]));
Q_AN02 U3657 ( .A0(n279), .A1(oMark[140]), .Z(n5087));
Q_FDP0UA U3658 ( .D(n5086), .QTFCLK( ), .Q(oMark[139]));
Q_AN02 U3659 ( .A0(n279), .A1(oMark[139]), .Z(n5086));
Q_FDP0UA U3660 ( .D(n5085), .QTFCLK( ), .Q(oMark[138]));
Q_AN02 U3661 ( .A0(n279), .A1(oMark[138]), .Z(n5085));
Q_FDP0UA U3662 ( .D(n5084), .QTFCLK( ), .Q(oMark[137]));
Q_AN02 U3663 ( .A0(n279), .A1(oMark[137]), .Z(n5084));
Q_FDP0UA U3664 ( .D(n5083), .QTFCLK( ), .Q(oMark[136]));
Q_AN02 U3665 ( .A0(n279), .A1(oMark[136]), .Z(n5083));
Q_FDP0UA U3666 ( .D(n5082), .QTFCLK( ), .Q(oMark[135]));
Q_AN02 U3667 ( .A0(n279), .A1(oMark[135]), .Z(n5082));
Q_FDP0UA U3668 ( .D(n5081), .QTFCLK( ), .Q(oMark[134]));
Q_AN02 U3669 ( .A0(n279), .A1(oMark[134]), .Z(n5081));
Q_FDP0UA U3670 ( .D(n5080), .QTFCLK( ), .Q(oMark[133]));
Q_AN02 U3671 ( .A0(n279), .A1(oMark[133]), .Z(n5080));
Q_FDP0UA U3672 ( .D(n5079), .QTFCLK( ), .Q(oMark[132]));
Q_AN02 U3673 ( .A0(n279), .A1(oMark[132]), .Z(n5079));
Q_FDP0UA U3674 ( .D(n5078), .QTFCLK( ), .Q(oMark[131]));
Q_AN02 U3675 ( .A0(n279), .A1(oMark[131]), .Z(n5078));
Q_FDP0UA U3676 ( .D(n5077), .QTFCLK( ), .Q(oMark[130]));
Q_AN02 U3677 ( .A0(n279), .A1(oMark[130]), .Z(n5077));
Q_FDP0UA U3678 ( .D(n5076), .QTFCLK( ), .Q(oMark[129]));
Q_AN02 U3679 ( .A0(n279), .A1(oMark[129]), .Z(n5076));
Q_FDP0UA U3680 ( .D(n5075), .QTFCLK( ), .Q(oMark[128]));
Q_AN02 U3681 ( .A0(n279), .A1(oMark[128]), .Z(n5075));
Q_FDP0UA U3682 ( .D(n5074), .QTFCLK( ), .Q(oMark[126]));
Q_AN02 U3683 ( .A0(n279), .A1(oMark[126]), .Z(n5074));
Q_FDP0UA U3684 ( .D(n5073), .QTFCLK( ), .Q(oMark[125]));
Q_AN02 U3685 ( .A0(n279), .A1(oMark[125]), .Z(n5073));
Q_FDP0UA U3686 ( .D(n5072), .QTFCLK( ), .Q(oMark[124]));
Q_AN02 U3687 ( .A0(n279), .A1(oMark[124]), .Z(n5072));
Q_FDP0UA U3688 ( .D(n5071), .QTFCLK( ), .Q(oMark[123]));
Q_AN02 U3689 ( .A0(n279), .A1(oMark[123]), .Z(n5071));
Q_FDP0UA U3690 ( .D(n5070), .QTFCLK( ), .Q(oMark[122]));
Q_AN02 U3691 ( .A0(n279), .A1(oMark[122]), .Z(n5070));
Q_FDP0UA U3692 ( .D(n5069), .QTFCLK( ), .Q(oMark[121]));
Q_AN02 U3693 ( .A0(n279), .A1(oMark[121]), .Z(n5069));
Q_FDP0UA U3694 ( .D(n5068), .QTFCLK( ), .Q(oMark[120]));
Q_AN02 U3695 ( .A0(n279), .A1(oMark[120]), .Z(n5068));
Q_FDP0UA U3696 ( .D(n5067), .QTFCLK( ), .Q(oMark[119]));
Q_AN02 U3697 ( .A0(n279), .A1(oMark[119]), .Z(n5067));
Q_FDP0UA U3698 ( .D(n5066), .QTFCLK( ), .Q(oMark[118]));
Q_AN02 U3699 ( .A0(n279), .A1(oMark[118]), .Z(n5066));
Q_FDP0UA U3700 ( .D(n5065), .QTFCLK( ), .Q(oMark[117]));
Q_AN02 U3701 ( .A0(n279), .A1(oMark[117]), .Z(n5065));
Q_FDP0UA U3702 ( .D(n5064), .QTFCLK( ), .Q(oMark[116]));
Q_AN02 U3703 ( .A0(n279), .A1(oMark[116]), .Z(n5064));
Q_FDP0UA U3704 ( .D(n5063), .QTFCLK( ), .Q(oMark[115]));
Q_AN02 U3705 ( .A0(n279), .A1(oMark[115]), .Z(n5063));
Q_FDP0UA U3706 ( .D(n5062), .QTFCLK( ), .Q(oMark[114]));
Q_AN02 U3707 ( .A0(n279), .A1(oMark[114]), .Z(n5062));
Q_FDP0UA U3708 ( .D(n5061), .QTFCLK( ), .Q(oMark[113]));
Q_AN02 U3709 ( .A0(n279), .A1(oMark[113]), .Z(n5061));
Q_FDP0UA U3710 ( .D(n5060), .QTFCLK( ), .Q(oMark[112]));
Q_AN02 U3711 ( .A0(n279), .A1(oMark[112]), .Z(n5060));
Q_FDP0UA U3712 ( .D(n5059), .QTFCLK( ), .Q(oMark[111]));
Q_AN02 U3713 ( .A0(n279), .A1(oMark[111]), .Z(n5059));
Q_FDP0UA U3714 ( .D(n5058), .QTFCLK( ), .Q(oMark[110]));
Q_AN02 U3715 ( .A0(n279), .A1(oMark[110]), .Z(n5058));
Q_FDP0UA U3716 ( .D(n5057), .QTFCLK( ), .Q(oMark[109]));
Q_AN02 U3717 ( .A0(n279), .A1(oMark[109]), .Z(n5057));
Q_FDP0UA U3718 ( .D(n5056), .QTFCLK( ), .Q(oMark[108]));
Q_AN02 U3719 ( .A0(n279), .A1(oMark[108]), .Z(n5056));
Q_FDP0UA U3720 ( .D(n5055), .QTFCLK( ), .Q(oMark[107]));
Q_AN02 U3721 ( .A0(n279), .A1(oMark[107]), .Z(n5055));
Q_FDP0UA U3722 ( .D(n5054), .QTFCLK( ), .Q(oMark[106]));
Q_AN02 U3723 ( .A0(n279), .A1(oMark[106]), .Z(n5054));
Q_FDP0UA U3724 ( .D(n5053), .QTFCLK( ), .Q(oMark[105]));
Q_AN02 U3725 ( .A0(n279), .A1(oMark[105]), .Z(n5053));
Q_FDP0UA U3726 ( .D(n5052), .QTFCLK( ), .Q(oMark[104]));
Q_AN02 U3727 ( .A0(n279), .A1(oMark[104]), .Z(n5052));
Q_FDP0UA U3728 ( .D(n5051), .QTFCLK( ), .Q(oMark[103]));
Q_AN02 U3729 ( .A0(n279), .A1(oMark[103]), .Z(n5051));
Q_FDP0UA U3730 ( .D(n5050), .QTFCLK( ), .Q(oMark[102]));
Q_AN02 U3731 ( .A0(n279), .A1(oMark[102]), .Z(n5050));
Q_FDP0UA U3732 ( .D(n5049), .QTFCLK( ), .Q(oMark[101]));
Q_AN02 U3733 ( .A0(n279), .A1(oMark[101]), .Z(n5049));
Q_FDP0UA U3734 ( .D(n5048), .QTFCLK( ), .Q(oMark[100]));
Q_AN02 U3735 ( .A0(n279), .A1(oMark[100]), .Z(n5048));
Q_FDP0UA U3736 ( .D(n5047), .QTFCLK( ), .Q(oMark[99]));
Q_AN02 U3737 ( .A0(n279), .A1(oMark[99]), .Z(n5047));
Q_FDP0UA U3738 ( .D(n5046), .QTFCLK( ), .Q(oMark[98]));
Q_AN02 U3739 ( .A0(n279), .A1(oMark[98]), .Z(n5046));
Q_FDP0UA U3740 ( .D(n5045), .QTFCLK( ), .Q(oMark[97]));
Q_AN02 U3741 ( .A0(n279), .A1(oMark[97]), .Z(n5045));
Q_FDP0UA U3742 ( .D(n5044), .QTFCLK( ), .Q(oMark[96]));
Q_AN02 U3743 ( .A0(n279), .A1(oMark[96]), .Z(n5044));
Q_FDP0UA U3744 ( .D(n5043), .QTFCLK( ), .Q(oMark[95]));
Q_AN02 U3745 ( .A0(n279), .A1(oMark[95]), .Z(n5043));
Q_FDP0UA U3746 ( .D(n5042), .QTFCLK( ), .Q(oMark[94]));
Q_AN02 U3747 ( .A0(n279), .A1(oMark[94]), .Z(n5042));
Q_FDP0UA U3748 ( .D(n5041), .QTFCLK( ), .Q(oMark[93]));
Q_AN02 U3749 ( .A0(n279), .A1(oMark[93]), .Z(n5041));
Q_FDP0UA U3750 ( .D(n5040), .QTFCLK( ), .Q(oMark[92]));
Q_AN02 U3751 ( .A0(n279), .A1(oMark[92]), .Z(n5040));
Q_FDP0UA U3752 ( .D(n5039), .QTFCLK( ), .Q(oMark[91]));
Q_AN02 U3753 ( .A0(n279), .A1(oMark[91]), .Z(n5039));
Q_FDP0UA U3754 ( .D(n5038), .QTFCLK( ), .Q(oMark[90]));
Q_AN02 U3755 ( .A0(n279), .A1(oMark[90]), .Z(n5038));
Q_FDP0UA U3756 ( .D(n5037), .QTFCLK( ), .Q(oMark[89]));
Q_AN02 U3757 ( .A0(n279), .A1(oMark[89]), .Z(n5037));
Q_FDP0UA U3758 ( .D(n5036), .QTFCLK( ), .Q(oMark[88]));
Q_AN02 U3759 ( .A0(n279), .A1(oMark[88]), .Z(n5036));
Q_FDP0UA U3760 ( .D(n5035), .QTFCLK( ), .Q(oMark[87]));
Q_AN02 U3761 ( .A0(n279), .A1(oMark[87]), .Z(n5035));
Q_FDP0UA U3762 ( .D(n5034), .QTFCLK( ), .Q(oMark[86]));
Q_AN02 U3763 ( .A0(n279), .A1(oMark[86]), .Z(n5034));
Q_FDP0UA U3764 ( .D(n5033), .QTFCLK( ), .Q(oMark[85]));
Q_AN02 U3765 ( .A0(n279), .A1(oMark[85]), .Z(n5033));
Q_FDP0UA U3766 ( .D(n5032), .QTFCLK( ), .Q(oMark[84]));
Q_AN02 U3767 ( .A0(n279), .A1(oMark[84]), .Z(n5032));
Q_FDP0UA U3768 ( .D(n5031), .QTFCLK( ), .Q(oMark[83]));
Q_AN02 U3769 ( .A0(n279), .A1(oMark[83]), .Z(n5031));
Q_FDP0UA U3770 ( .D(n5030), .QTFCLK( ), .Q(oMark[82]));
Q_AN02 U3771 ( .A0(n279), .A1(oMark[82]), .Z(n5030));
Q_FDP0UA U3772 ( .D(n5029), .QTFCLK( ), .Q(oMark[81]));
Q_AN02 U3773 ( .A0(n279), .A1(oMark[81]), .Z(n5029));
Q_FDP0UA U3774 ( .D(n5028), .QTFCLK( ), .Q(oMark[80]));
Q_AN02 U3775 ( .A0(n279), .A1(oMark[80]), .Z(n5028));
Q_FDP0UA U3776 ( .D(n5027), .QTFCLK( ), .Q(oMark[79]));
Q_AN02 U3777 ( .A0(n279), .A1(oMark[79]), .Z(n5027));
Q_FDP0UA U3778 ( .D(n5026), .QTFCLK( ), .Q(oMark[78]));
Q_AN02 U3779 ( .A0(n279), .A1(oMark[78]), .Z(n5026));
Q_FDP0UA U3780 ( .D(n5025), .QTFCLK( ), .Q(oMark[77]));
Q_AN02 U3781 ( .A0(n279), .A1(oMark[77]), .Z(n5025));
Q_FDP0UA U3782 ( .D(n5024), .QTFCLK( ), .Q(oMark[76]));
Q_AN02 U3783 ( .A0(n279), .A1(oMark[76]), .Z(n5024));
Q_FDP0UA U3784 ( .D(n5023), .QTFCLK( ), .Q(oMark[75]));
Q_AN02 U3785 ( .A0(n279), .A1(oMark[75]), .Z(n5023));
Q_FDP0UA U3786 ( .D(n5022), .QTFCLK( ), .Q(oMark[74]));
Q_AN02 U3787 ( .A0(n279), .A1(oMark[74]), .Z(n5022));
Q_FDP0UA U3788 ( .D(n5021), .QTFCLK( ), .Q(oMark[73]));
Q_AN02 U3789 ( .A0(n279), .A1(oMark[73]), .Z(n5021));
Q_FDP0UA U3790 ( .D(n5020), .QTFCLK( ), .Q(oMark[72]));
Q_AN02 U3791 ( .A0(n279), .A1(oMark[72]), .Z(n5020));
Q_FDP0UA U3792 ( .D(n5019), .QTFCLK( ), .Q(oMark[71]));
Q_AN02 U3793 ( .A0(n279), .A1(oMark[71]), .Z(n5019));
Q_FDP0UA U3794 ( .D(n5018), .QTFCLK( ), .Q(oMark[70]));
Q_AN02 U3795 ( .A0(n279), .A1(oMark[70]), .Z(n5018));
Q_FDP0UA U3796 ( .D(n5017), .QTFCLK( ), .Q(oMark[69]));
Q_AN02 U3797 ( .A0(n279), .A1(oMark[69]), .Z(n5017));
Q_FDP0UA U3798 ( .D(n5016), .QTFCLK( ), .Q(oMark[68]));
Q_AN02 U3799 ( .A0(n279), .A1(oMark[68]), .Z(n5016));
Q_FDP0UA U3800 ( .D(n5015), .QTFCLK( ), .Q(oMark[67]));
Q_AN02 U3801 ( .A0(n279), .A1(oMark[67]), .Z(n5015));
Q_FDP0UA U3802 ( .D(n5014), .QTFCLK( ), .Q(oMark[66]));
Q_AN02 U3803 ( .A0(n279), .A1(oMark[66]), .Z(n5014));
Q_FDP0UA U3804 ( .D(n5013), .QTFCLK( ), .Q(oMark[65]));
Q_AN02 U3805 ( .A0(n279), .A1(oMark[65]), .Z(n5013));
Q_FDP0UA U3806 ( .D(n5012), .QTFCLK( ), .Q(oMark[64]));
Q_AN02 U3807 ( .A0(n279), .A1(oMark[64]), .Z(n5012));
Q_AN02 U3808 ( .A0(oFill[0]), .A1(oData[511]), .Z(n5011));
Q_AN02 U3809 ( .A0(oFill[0]), .A1(oData[510]), .Z(n5010));
Q_AN02 U3810 ( .A0(oFill[0]), .A1(oData[509]), .Z(n5009));
Q_AN02 U3811 ( .A0(oFill[0]), .A1(oData[508]), .Z(n5008));
Q_AN02 U3812 ( .A0(oFill[0]), .A1(oData[507]), .Z(n5007));
Q_AN02 U3813 ( .A0(oFill[0]), .A1(oData[506]), .Z(n5006));
Q_AN02 U3814 ( .A0(oFill[0]), .A1(oData[505]), .Z(n5005));
Q_AN02 U3815 ( .A0(oFill[0]), .A1(oData[504]), .Z(n5004));
Q_AN02 U3816 ( .A0(oFill[0]), .A1(oData[503]), .Z(n5003));
Q_AN02 U3817 ( .A0(oFill[0]), .A1(oData[502]), .Z(n5002));
Q_AN02 U3818 ( .A0(oFill[0]), .A1(oData[501]), .Z(n5001));
Q_AN02 U3819 ( .A0(oFill[0]), .A1(oData[500]), .Z(n5000));
Q_AN02 U3820 ( .A0(oFill[0]), .A1(oData[499]), .Z(n4999));
Q_AN02 U3821 ( .A0(oFill[0]), .A1(oData[498]), .Z(n4998));
Q_AN02 U3822 ( .A0(oFill[0]), .A1(oData[497]), .Z(n4997));
Q_AN02 U3823 ( .A0(oFill[0]), .A1(oData[496]), .Z(n4996));
Q_AN02 U3824 ( .A0(oFill[0]), .A1(oData[495]), .Z(n4995));
Q_AN02 U3825 ( .A0(oFill[0]), .A1(oData[494]), .Z(n4994));
Q_AN02 U3826 ( .A0(oFill[0]), .A1(oData[493]), .Z(n4993));
Q_AN02 U3827 ( .A0(oFill[0]), .A1(oData[492]), .Z(n4992));
Q_AN02 U3828 ( .A0(oFill[0]), .A1(oData[491]), .Z(n4991));
Q_AN02 U3829 ( .A0(oFill[0]), .A1(oData[490]), .Z(n4990));
Q_AN02 U3830 ( .A0(oFill[0]), .A1(oData[489]), .Z(n4989));
Q_AN02 U3831 ( .A0(oFill[0]), .A1(oData[488]), .Z(n4988));
Q_AN02 U3832 ( .A0(oFill[0]), .A1(oData[487]), .Z(n4987));
Q_AN02 U3833 ( .A0(oFill[0]), .A1(oData[486]), .Z(n4986));
Q_AN02 U3834 ( .A0(oFill[0]), .A1(oData[485]), .Z(n4985));
Q_AN02 U3835 ( .A0(oFill[0]), .A1(oData[484]), .Z(n4984));
Q_AN02 U3836 ( .A0(oFill[0]), .A1(oData[483]), .Z(n4983));
Q_AN02 U3837 ( .A0(oFill[0]), .A1(oData[482]), .Z(n4982));
Q_AN02 U3838 ( .A0(oFill[0]), .A1(oData[481]), .Z(n4981));
Q_AN02 U3839 ( .A0(oFill[0]), .A1(oData[480]), .Z(n4980));
Q_AN02 U3840 ( .A0(oFill[0]), .A1(oData[479]), .Z(n4979));
Q_AN02 U3841 ( .A0(oFill[0]), .A1(oData[478]), .Z(n4978));
Q_AN02 U3842 ( .A0(oFill[0]), .A1(oData[477]), .Z(n4977));
Q_AN02 U3843 ( .A0(oFill[0]), .A1(oData[476]), .Z(n4976));
Q_AN02 U3844 ( .A0(oFill[0]), .A1(oData[475]), .Z(n4975));
Q_AN02 U3845 ( .A0(oFill[0]), .A1(oData[474]), .Z(n4974));
Q_AN02 U3846 ( .A0(oFill[0]), .A1(oData[473]), .Z(n4973));
Q_AN02 U3847 ( .A0(oFill[0]), .A1(oData[472]), .Z(n4972));
Q_AN02 U3848 ( .A0(oFill[0]), .A1(oData[471]), .Z(n4971));
Q_AN02 U3849 ( .A0(oFill[0]), .A1(oData[470]), .Z(n4970));
Q_AN02 U3850 ( .A0(oFill[0]), .A1(oData[469]), .Z(n4969));
Q_AN02 U3851 ( .A0(oFill[0]), .A1(oData[468]), .Z(n4968));
Q_AN02 U3852 ( .A0(oFill[0]), .A1(oData[467]), .Z(n4967));
Q_AN02 U3853 ( .A0(oFill[0]), .A1(oData[466]), .Z(n4966));
Q_AN02 U3854 ( .A0(oFill[0]), .A1(oData[465]), .Z(n4965));
Q_AN02 U3855 ( .A0(oFill[0]), .A1(oData[464]), .Z(n4964));
Q_AN02 U3856 ( .A0(oFill[0]), .A1(oData[463]), .Z(n4963));
Q_AN02 U3857 ( .A0(oFill[0]), .A1(oData[462]), .Z(n4962));
Q_AN02 U3858 ( .A0(oFill[0]), .A1(oData[461]), .Z(n4961));
Q_AN02 U3859 ( .A0(oFill[0]), .A1(oData[460]), .Z(n4960));
Q_AN02 U3860 ( .A0(oFill[0]), .A1(oData[459]), .Z(n4959));
Q_AN02 U3861 ( .A0(oFill[0]), .A1(oData[458]), .Z(n4958));
Q_AN02 U3862 ( .A0(oFill[0]), .A1(oData[457]), .Z(n4957));
Q_AN02 U3863 ( .A0(oFill[0]), .A1(oData[456]), .Z(n4956));
Q_AN02 U3864 ( .A0(oFill[0]), .A1(oData[455]), .Z(n4955));
Q_AN02 U3865 ( .A0(oFill[0]), .A1(oData[454]), .Z(n4954));
Q_AN02 U3866 ( .A0(oFill[0]), .A1(oData[453]), .Z(n4953));
Q_AN02 U3867 ( .A0(oFill[0]), .A1(oData[452]), .Z(n4952));
Q_AN02 U3868 ( .A0(oFill[0]), .A1(oData[451]), .Z(n4951));
Q_AN02 U3869 ( .A0(oFill[0]), .A1(oData[450]), .Z(n4950));
Q_AN02 U3870 ( .A0(oFill[0]), .A1(oData[449]), .Z(n4949));
Q_AN02 U3871 ( .A0(oFill[0]), .A1(oData[448]), .Z(n4948));
Q_MX02 U3872 ( .S(oFill[0]), .A0(oData[511]), .A1(oData[447]), .Z(n4947));
Q_MX02 U3873 ( .S(oFill[0]), .A0(oData[510]), .A1(oData[446]), .Z(n4946));
Q_MX02 U3874 ( .S(oFill[0]), .A0(oData[509]), .A1(oData[445]), .Z(n4945));
Q_MX02 U3875 ( .S(oFill[0]), .A0(oData[508]), .A1(oData[444]), .Z(n4944));
Q_MX02 U3876 ( .S(oFill[0]), .A0(oData[507]), .A1(oData[443]), .Z(n4943));
Q_MX02 U3877 ( .S(oFill[0]), .A0(oData[506]), .A1(oData[442]), .Z(n4942));
Q_MX02 U3878 ( .S(oFill[0]), .A0(oData[505]), .A1(oData[441]), .Z(n4941));
Q_MX02 U3879 ( .S(oFill[0]), .A0(oData[504]), .A1(oData[440]), .Z(n4940));
Q_MX02 U3880 ( .S(oFill[0]), .A0(oData[503]), .A1(oData[439]), .Z(n4939));
Q_MX02 U3881 ( .S(oFill[0]), .A0(oData[502]), .A1(oData[438]), .Z(n4938));
Q_MX02 U3882 ( .S(oFill[0]), .A0(oData[501]), .A1(oData[437]), .Z(n4937));
Q_MX02 U3883 ( .S(oFill[0]), .A0(oData[500]), .A1(oData[436]), .Z(n4936));
Q_MX02 U3884 ( .S(oFill[0]), .A0(oData[499]), .A1(oData[435]), .Z(n4935));
Q_MX02 U3885 ( .S(oFill[0]), .A0(oData[498]), .A1(oData[434]), .Z(n4934));
Q_MX02 U3886 ( .S(oFill[0]), .A0(oData[497]), .A1(oData[433]), .Z(n4933));
Q_MX02 U3887 ( .S(oFill[0]), .A0(oData[496]), .A1(oData[432]), .Z(n4932));
Q_MX02 U3888 ( .S(oFill[0]), .A0(oData[495]), .A1(oData[431]), .Z(n4931));
Q_MX02 U3889 ( .S(oFill[0]), .A0(oData[494]), .A1(oData[430]), .Z(n4930));
Q_MX02 U3890 ( .S(oFill[0]), .A0(oData[493]), .A1(oData[429]), .Z(n4929));
Q_MX02 U3891 ( .S(oFill[0]), .A0(oData[492]), .A1(oData[428]), .Z(n4928));
Q_MX02 U3892 ( .S(oFill[0]), .A0(oData[491]), .A1(oData[427]), .Z(n4927));
Q_MX02 U3893 ( .S(oFill[0]), .A0(oData[490]), .A1(oData[426]), .Z(n4926));
Q_MX02 U3894 ( .S(oFill[0]), .A0(oData[489]), .A1(oData[425]), .Z(n4925));
Q_MX02 U3895 ( .S(oFill[0]), .A0(oData[488]), .A1(oData[424]), .Z(n4924));
Q_MX02 U3896 ( .S(oFill[0]), .A0(oData[487]), .A1(oData[423]), .Z(n4923));
Q_MX02 U3897 ( .S(oFill[0]), .A0(oData[486]), .A1(oData[422]), .Z(n4922));
Q_MX02 U3898 ( .S(oFill[0]), .A0(oData[485]), .A1(oData[421]), .Z(n4921));
Q_MX02 U3899 ( .S(oFill[0]), .A0(oData[484]), .A1(oData[420]), .Z(n4920));
Q_MX02 U3900 ( .S(oFill[0]), .A0(oData[483]), .A1(oData[419]), .Z(n4919));
Q_MX02 U3901 ( .S(oFill[0]), .A0(oData[482]), .A1(oData[418]), .Z(n4918));
Q_MX02 U3902 ( .S(oFill[0]), .A0(oData[481]), .A1(oData[417]), .Z(n4917));
Q_MX02 U3903 ( .S(oFill[0]), .A0(oData[480]), .A1(oData[416]), .Z(n4916));
Q_MX02 U3904 ( .S(oFill[0]), .A0(oData[479]), .A1(oData[415]), .Z(n4915));
Q_MX02 U3905 ( .S(oFill[0]), .A0(oData[478]), .A1(oData[414]), .Z(n4914));
Q_MX02 U3906 ( .S(oFill[0]), .A0(oData[477]), .A1(oData[413]), .Z(n4913));
Q_MX02 U3907 ( .S(oFill[0]), .A0(oData[476]), .A1(oData[412]), .Z(n4912));
Q_MX02 U3908 ( .S(oFill[0]), .A0(oData[475]), .A1(oData[411]), .Z(n4911));
Q_MX02 U3909 ( .S(oFill[0]), .A0(oData[474]), .A1(oData[410]), .Z(n4910));
Q_MX02 U3910 ( .S(oFill[0]), .A0(oData[473]), .A1(oData[409]), .Z(n4909));
Q_MX02 U3911 ( .S(oFill[0]), .A0(oData[472]), .A1(oData[408]), .Z(n4908));
Q_MX02 U3912 ( .S(oFill[0]), .A0(oData[471]), .A1(oData[407]), .Z(n4907));
Q_MX02 U3913 ( .S(oFill[0]), .A0(oData[470]), .A1(oData[406]), .Z(n4906));
Q_MX02 U3914 ( .S(oFill[0]), .A0(oData[469]), .A1(oData[405]), .Z(n4905));
Q_MX02 U3915 ( .S(oFill[0]), .A0(oData[468]), .A1(oData[404]), .Z(n4904));
Q_MX02 U3916 ( .S(oFill[0]), .A0(oData[467]), .A1(oData[403]), .Z(n4903));
Q_MX02 U3917 ( .S(oFill[0]), .A0(oData[466]), .A1(oData[402]), .Z(n4902));
Q_MX02 U3918 ( .S(oFill[0]), .A0(oData[465]), .A1(oData[401]), .Z(n4901));
Q_MX02 U3919 ( .S(oFill[0]), .A0(oData[464]), .A1(oData[400]), .Z(n4900));
Q_MX02 U3920 ( .S(oFill[0]), .A0(oData[463]), .A1(oData[399]), .Z(n4899));
Q_MX02 U3921 ( .S(oFill[0]), .A0(oData[462]), .A1(oData[398]), .Z(n4898));
Q_MX02 U3922 ( .S(oFill[0]), .A0(oData[461]), .A1(oData[397]), .Z(n4897));
Q_MX02 U3923 ( .S(oFill[0]), .A0(oData[460]), .A1(oData[396]), .Z(n4896));
Q_MX02 U3924 ( .S(oFill[0]), .A0(oData[459]), .A1(oData[395]), .Z(n4895));
Q_MX02 U3925 ( .S(oFill[0]), .A0(oData[458]), .A1(oData[394]), .Z(n4894));
Q_MX02 U3926 ( .S(oFill[0]), .A0(oData[457]), .A1(oData[393]), .Z(n4893));
Q_MX02 U3927 ( .S(oFill[0]), .A0(oData[456]), .A1(oData[392]), .Z(n4892));
Q_MX02 U3928 ( .S(oFill[0]), .A0(oData[455]), .A1(oData[391]), .Z(n4891));
Q_MX02 U3929 ( .S(oFill[0]), .A0(oData[454]), .A1(oData[390]), .Z(n4890));
Q_MX02 U3930 ( .S(oFill[0]), .A0(oData[453]), .A1(oData[389]), .Z(n4889));
Q_MX02 U3931 ( .S(oFill[0]), .A0(oData[452]), .A1(oData[388]), .Z(n4888));
Q_MX02 U3932 ( .S(oFill[0]), .A0(oData[451]), .A1(oData[387]), .Z(n4887));
Q_MX02 U3933 ( .S(oFill[0]), .A0(oData[450]), .A1(oData[386]), .Z(n4886));
Q_MX02 U3934 ( .S(oFill[0]), .A0(oData[449]), .A1(oData[385]), .Z(n4885));
Q_MX02 U3935 ( .S(oFill[0]), .A0(oData[448]), .A1(oData[384]), .Z(n4884));
Q_MX02 U3936 ( .S(oFill[0]), .A0(oData[447]), .A1(oData[383]), .Z(n4883));
Q_MX02 U3937 ( .S(oFill[0]), .A0(oData[446]), .A1(oData[382]), .Z(n4882));
Q_MX02 U3938 ( .S(oFill[0]), .A0(oData[445]), .A1(oData[381]), .Z(n4881));
Q_MX02 U3939 ( .S(oFill[0]), .A0(oData[444]), .A1(oData[380]), .Z(n4880));
Q_MX02 U3940 ( .S(oFill[0]), .A0(oData[443]), .A1(oData[379]), .Z(n4879));
Q_MX02 U3941 ( .S(oFill[0]), .A0(oData[442]), .A1(oData[378]), .Z(n4878));
Q_MX02 U3942 ( .S(oFill[0]), .A0(oData[441]), .A1(oData[377]), .Z(n4877));
Q_MX02 U3943 ( .S(oFill[0]), .A0(oData[440]), .A1(oData[376]), .Z(n4876));
Q_MX02 U3944 ( .S(oFill[0]), .A0(oData[439]), .A1(oData[375]), .Z(n4875));
Q_MX02 U3945 ( .S(oFill[0]), .A0(oData[438]), .A1(oData[374]), .Z(n4874));
Q_MX02 U3946 ( .S(oFill[0]), .A0(oData[437]), .A1(oData[373]), .Z(n4873));
Q_MX02 U3947 ( .S(oFill[0]), .A0(oData[436]), .A1(oData[372]), .Z(n4872));
Q_MX02 U3948 ( .S(oFill[0]), .A0(oData[435]), .A1(oData[371]), .Z(n4871));
Q_MX02 U3949 ( .S(oFill[0]), .A0(oData[434]), .A1(oData[370]), .Z(n4870));
Q_MX02 U3950 ( .S(oFill[0]), .A0(oData[433]), .A1(oData[369]), .Z(n4869));
Q_MX02 U3951 ( .S(oFill[0]), .A0(oData[432]), .A1(oData[368]), .Z(n4868));
Q_MX02 U3952 ( .S(oFill[0]), .A0(oData[431]), .A1(oData[367]), .Z(n4867));
Q_MX02 U3953 ( .S(oFill[0]), .A0(oData[430]), .A1(oData[366]), .Z(n4866));
Q_MX02 U3954 ( .S(oFill[0]), .A0(oData[429]), .A1(oData[365]), .Z(n4865));
Q_MX02 U3955 ( .S(oFill[0]), .A0(oData[428]), .A1(oData[364]), .Z(n4864));
Q_MX02 U3956 ( .S(oFill[0]), .A0(oData[427]), .A1(oData[363]), .Z(n4863));
Q_MX02 U3957 ( .S(oFill[0]), .A0(oData[426]), .A1(oData[362]), .Z(n4862));
Q_MX02 U3958 ( .S(oFill[0]), .A0(oData[425]), .A1(oData[361]), .Z(n4861));
Q_MX02 U3959 ( .S(oFill[0]), .A0(oData[424]), .A1(oData[360]), .Z(n4860));
Q_MX02 U3960 ( .S(oFill[0]), .A0(oData[423]), .A1(oData[359]), .Z(n4859));
Q_MX02 U3961 ( .S(oFill[0]), .A0(oData[422]), .A1(oData[358]), .Z(n4858));
Q_MX02 U3962 ( .S(oFill[0]), .A0(oData[421]), .A1(oData[357]), .Z(n4857));
Q_MX02 U3963 ( .S(oFill[0]), .A0(oData[420]), .A1(oData[356]), .Z(n4856));
Q_MX02 U3964 ( .S(oFill[0]), .A0(oData[419]), .A1(oData[355]), .Z(n4855));
Q_MX02 U3965 ( .S(oFill[0]), .A0(oData[418]), .A1(oData[354]), .Z(n4854));
Q_MX02 U3966 ( .S(oFill[0]), .A0(oData[417]), .A1(oData[353]), .Z(n4853));
Q_MX02 U3967 ( .S(oFill[0]), .A0(oData[416]), .A1(oData[352]), .Z(n4852));
Q_MX02 U3968 ( .S(oFill[0]), .A0(oData[415]), .A1(oData[351]), .Z(n4851));
Q_MX02 U3969 ( .S(oFill[0]), .A0(oData[414]), .A1(oData[350]), .Z(n4850));
Q_MX02 U3970 ( .S(oFill[0]), .A0(oData[413]), .A1(oData[349]), .Z(n4849));
Q_MX02 U3971 ( .S(oFill[0]), .A0(oData[412]), .A1(oData[348]), .Z(n4848));
Q_MX02 U3972 ( .S(oFill[0]), .A0(oData[411]), .A1(oData[347]), .Z(n4847));
Q_MX02 U3973 ( .S(oFill[0]), .A0(oData[410]), .A1(oData[346]), .Z(n4846));
Q_MX02 U3974 ( .S(oFill[0]), .A0(oData[409]), .A1(oData[345]), .Z(n4845));
Q_MX02 U3975 ( .S(oFill[0]), .A0(oData[408]), .A1(oData[344]), .Z(n4844));
Q_MX02 U3976 ( .S(oFill[0]), .A0(oData[407]), .A1(oData[343]), .Z(n4843));
Q_MX02 U3977 ( .S(oFill[0]), .A0(oData[406]), .A1(oData[342]), .Z(n4842));
Q_MX02 U3978 ( .S(oFill[0]), .A0(oData[405]), .A1(oData[341]), .Z(n4841));
Q_MX02 U3979 ( .S(oFill[0]), .A0(oData[404]), .A1(oData[340]), .Z(n4840));
Q_MX02 U3980 ( .S(oFill[0]), .A0(oData[403]), .A1(oData[339]), .Z(n4839));
Q_MX02 U3981 ( .S(oFill[0]), .A0(oData[402]), .A1(oData[338]), .Z(n4838));
Q_MX02 U3982 ( .S(oFill[0]), .A0(oData[401]), .A1(oData[337]), .Z(n4837));
Q_MX02 U3983 ( .S(oFill[0]), .A0(oData[400]), .A1(oData[336]), .Z(n4836));
Q_MX02 U3984 ( .S(oFill[0]), .A0(oData[399]), .A1(oData[335]), .Z(n4835));
Q_MX02 U3985 ( .S(oFill[0]), .A0(oData[398]), .A1(oData[334]), .Z(n4834));
Q_MX02 U3986 ( .S(oFill[0]), .A0(oData[397]), .A1(oData[333]), .Z(n4833));
Q_MX02 U3987 ( .S(oFill[0]), .A0(oData[396]), .A1(oData[332]), .Z(n4832));
Q_MX02 U3988 ( .S(oFill[0]), .A0(oData[395]), .A1(oData[331]), .Z(n4831));
Q_MX02 U3989 ( .S(oFill[0]), .A0(oData[394]), .A1(oData[330]), .Z(n4830));
Q_MX02 U3990 ( .S(oFill[0]), .A0(oData[393]), .A1(oData[329]), .Z(n4829));
Q_MX02 U3991 ( .S(oFill[0]), .A0(oData[392]), .A1(oData[328]), .Z(n4828));
Q_MX02 U3992 ( .S(oFill[0]), .A0(oData[391]), .A1(oData[327]), .Z(n4827));
Q_MX02 U3993 ( .S(oFill[0]), .A0(oData[390]), .A1(oData[326]), .Z(n4826));
Q_MX02 U3994 ( .S(oFill[0]), .A0(oData[389]), .A1(oData[325]), .Z(n4825));
Q_MX02 U3995 ( .S(oFill[0]), .A0(oData[388]), .A1(oData[324]), .Z(n4824));
Q_MX02 U3996 ( .S(oFill[0]), .A0(oData[387]), .A1(oData[323]), .Z(n4823));
Q_MX02 U3997 ( .S(oFill[0]), .A0(oData[386]), .A1(oData[322]), .Z(n4822));
Q_MX02 U3998 ( .S(oFill[0]), .A0(oData[385]), .A1(oData[321]), .Z(n4821));
Q_MX02 U3999 ( .S(oFill[0]), .A0(oData[384]), .A1(oData[320]), .Z(n4820));
Q_MX02 U4000 ( .S(oFill[0]), .A0(oData[383]), .A1(oData[319]), .Z(n4819));
Q_MX02 U4001 ( .S(oFill[0]), .A0(oData[382]), .A1(oData[318]), .Z(n4818));
Q_MX02 U4002 ( .S(oFill[0]), .A0(oData[381]), .A1(oData[317]), .Z(n4817));
Q_MX02 U4003 ( .S(oFill[0]), .A0(oData[380]), .A1(oData[316]), .Z(n4816));
Q_MX02 U4004 ( .S(oFill[0]), .A0(oData[379]), .A1(oData[315]), .Z(n4815));
Q_MX02 U4005 ( .S(oFill[0]), .A0(oData[378]), .A1(oData[314]), .Z(n4814));
Q_MX02 U4006 ( .S(oFill[0]), .A0(oData[377]), .A1(oData[313]), .Z(n4813));
Q_MX02 U4007 ( .S(oFill[0]), .A0(oData[376]), .A1(oData[312]), .Z(n4812));
Q_MX02 U4008 ( .S(oFill[0]), .A0(oData[375]), .A1(oData[311]), .Z(n4811));
Q_MX02 U4009 ( .S(oFill[0]), .A0(oData[374]), .A1(oData[310]), .Z(n4810));
Q_MX02 U4010 ( .S(oFill[0]), .A0(oData[373]), .A1(oData[309]), .Z(n4809));
Q_MX02 U4011 ( .S(oFill[0]), .A0(oData[372]), .A1(oData[308]), .Z(n4808));
Q_MX02 U4012 ( .S(oFill[0]), .A0(oData[371]), .A1(oData[307]), .Z(n4807));
Q_MX02 U4013 ( .S(oFill[0]), .A0(oData[370]), .A1(oData[306]), .Z(n4806));
Q_MX02 U4014 ( .S(oFill[0]), .A0(oData[369]), .A1(oData[305]), .Z(n4805));
Q_MX02 U4015 ( .S(oFill[0]), .A0(oData[368]), .A1(oData[304]), .Z(n4804));
Q_MX02 U4016 ( .S(oFill[0]), .A0(oData[367]), .A1(oData[303]), .Z(n4803));
Q_MX02 U4017 ( .S(oFill[0]), .A0(oData[366]), .A1(oData[302]), .Z(n4802));
Q_MX02 U4018 ( .S(oFill[0]), .A0(oData[365]), .A1(oData[301]), .Z(n4801));
Q_MX02 U4019 ( .S(oFill[0]), .A0(oData[364]), .A1(oData[300]), .Z(n4800));
Q_MX02 U4020 ( .S(oFill[0]), .A0(oData[363]), .A1(oData[299]), .Z(n4799));
Q_MX02 U4021 ( .S(oFill[0]), .A0(oData[362]), .A1(oData[298]), .Z(n4798));
Q_MX02 U4022 ( .S(oFill[0]), .A0(oData[361]), .A1(oData[297]), .Z(n4797));
Q_MX02 U4023 ( .S(oFill[0]), .A0(oData[360]), .A1(oData[296]), .Z(n4796));
Q_MX02 U4024 ( .S(oFill[0]), .A0(oData[359]), .A1(oData[295]), .Z(n4795));
Q_MX02 U4025 ( .S(oFill[0]), .A0(oData[358]), .A1(oData[294]), .Z(n4794));
Q_MX02 U4026 ( .S(oFill[0]), .A0(oData[357]), .A1(oData[293]), .Z(n4793));
Q_MX02 U4027 ( .S(oFill[0]), .A0(oData[356]), .A1(oData[292]), .Z(n4792));
Q_MX02 U4028 ( .S(oFill[0]), .A0(oData[355]), .A1(oData[291]), .Z(n4791));
Q_MX02 U4029 ( .S(oFill[0]), .A0(oData[354]), .A1(oData[290]), .Z(n4790));
Q_MX02 U4030 ( .S(oFill[0]), .A0(oData[353]), .A1(oData[289]), .Z(n4789));
Q_MX02 U4031 ( .S(oFill[0]), .A0(oData[352]), .A1(oData[288]), .Z(n4788));
Q_MX02 U4032 ( .S(oFill[0]), .A0(oData[351]), .A1(oData[287]), .Z(n4787));
Q_MX02 U4033 ( .S(oFill[0]), .A0(oData[350]), .A1(oData[286]), .Z(n4786));
Q_MX02 U4034 ( .S(oFill[0]), .A0(oData[349]), .A1(oData[285]), .Z(n4785));
Q_MX02 U4035 ( .S(oFill[0]), .A0(oData[348]), .A1(oData[284]), .Z(n4784));
Q_MX02 U4036 ( .S(oFill[0]), .A0(oData[347]), .A1(oData[283]), .Z(n4783));
Q_MX02 U4037 ( .S(oFill[0]), .A0(oData[346]), .A1(oData[282]), .Z(n4782));
Q_MX02 U4038 ( .S(oFill[0]), .A0(oData[345]), .A1(oData[281]), .Z(n4781));
Q_MX02 U4039 ( .S(oFill[0]), .A0(oData[344]), .A1(oData[280]), .Z(n4780));
Q_MX02 U4040 ( .S(oFill[0]), .A0(oData[343]), .A1(oData[279]), .Z(n4779));
Q_MX02 U4041 ( .S(oFill[0]), .A0(oData[342]), .A1(oData[278]), .Z(n4778));
Q_MX02 U4042 ( .S(oFill[0]), .A0(oData[341]), .A1(oData[277]), .Z(n4777));
Q_MX02 U4043 ( .S(oFill[0]), .A0(oData[340]), .A1(oData[276]), .Z(n4776));
Q_MX02 U4044 ( .S(oFill[0]), .A0(oData[339]), .A1(oData[275]), .Z(n4775));
Q_MX02 U4045 ( .S(oFill[0]), .A0(oData[338]), .A1(oData[274]), .Z(n4774));
Q_MX02 U4046 ( .S(oFill[0]), .A0(oData[337]), .A1(oData[273]), .Z(n4773));
Q_MX02 U4047 ( .S(oFill[0]), .A0(oData[336]), .A1(oData[272]), .Z(n4772));
Q_MX02 U4048 ( .S(oFill[0]), .A0(oData[335]), .A1(oData[271]), .Z(n4771));
Q_MX02 U4049 ( .S(oFill[0]), .A0(oData[334]), .A1(oData[270]), .Z(n4770));
Q_MX02 U4050 ( .S(oFill[0]), .A0(oData[333]), .A1(oData[269]), .Z(n4769));
Q_MX02 U4051 ( .S(oFill[0]), .A0(oData[332]), .A1(oData[268]), .Z(n4768));
Q_MX02 U4052 ( .S(oFill[0]), .A0(oData[331]), .A1(oData[267]), .Z(n4767));
Q_MX02 U4053 ( .S(oFill[0]), .A0(oData[330]), .A1(oData[266]), .Z(n4766));
Q_MX02 U4054 ( .S(oFill[0]), .A0(oData[329]), .A1(oData[265]), .Z(n4765));
Q_MX02 U4055 ( .S(oFill[0]), .A0(oData[328]), .A1(oData[264]), .Z(n4764));
Q_MX02 U4056 ( .S(oFill[0]), .A0(oData[327]), .A1(oData[263]), .Z(n4763));
Q_MX02 U4057 ( .S(oFill[0]), .A0(oData[326]), .A1(oData[262]), .Z(n4762));
Q_MX02 U4058 ( .S(oFill[0]), .A0(oData[325]), .A1(oData[261]), .Z(n4761));
Q_MX02 U4059 ( .S(oFill[0]), .A0(oData[324]), .A1(oData[260]), .Z(n4760));
Q_MX02 U4060 ( .S(oFill[0]), .A0(oData[323]), .A1(oData[259]), .Z(n4759));
Q_MX02 U4061 ( .S(oFill[0]), .A0(oData[322]), .A1(oData[258]), .Z(n4758));
Q_MX02 U4062 ( .S(oFill[0]), .A0(oData[321]), .A1(oData[257]), .Z(n4757));
Q_MX02 U4063 ( .S(oFill[0]), .A0(oData[320]), .A1(oData[256]), .Z(n4756));
Q_MX02 U4064 ( .S(oFill[0]), .A0(oData[319]), .A1(oData[255]), .Z(n4755));
Q_MX02 U4065 ( .S(oFill[0]), .A0(oData[318]), .A1(oData[254]), .Z(n4754));
Q_MX02 U4066 ( .S(oFill[0]), .A0(oData[317]), .A1(oData[253]), .Z(n4753));
Q_MX02 U4067 ( .S(oFill[0]), .A0(oData[316]), .A1(oData[252]), .Z(n4752));
Q_MX02 U4068 ( .S(oFill[0]), .A0(oData[315]), .A1(oData[251]), .Z(n4751));
Q_MX02 U4069 ( .S(oFill[0]), .A0(oData[314]), .A1(oData[250]), .Z(n4750));
Q_MX02 U4070 ( .S(oFill[0]), .A0(oData[313]), .A1(oData[249]), .Z(n4749));
Q_MX02 U4071 ( .S(oFill[0]), .A0(oData[312]), .A1(oData[248]), .Z(n4748));
Q_MX02 U4072 ( .S(oFill[0]), .A0(oData[311]), .A1(oData[247]), .Z(n4747));
Q_MX02 U4073 ( .S(oFill[0]), .A0(oData[310]), .A1(oData[246]), .Z(n4746));
Q_MX02 U4074 ( .S(oFill[0]), .A0(oData[309]), .A1(oData[245]), .Z(n4745));
Q_MX02 U4075 ( .S(oFill[0]), .A0(oData[308]), .A1(oData[244]), .Z(n4744));
Q_MX02 U4076 ( .S(oFill[0]), .A0(oData[307]), .A1(oData[243]), .Z(n4743));
Q_MX02 U4077 ( .S(oFill[0]), .A0(oData[306]), .A1(oData[242]), .Z(n4742));
Q_MX02 U4078 ( .S(oFill[0]), .A0(oData[305]), .A1(oData[241]), .Z(n4741));
Q_MX02 U4079 ( .S(oFill[0]), .A0(oData[304]), .A1(oData[240]), .Z(n4740));
Q_MX02 U4080 ( .S(oFill[0]), .A0(oData[303]), .A1(oData[239]), .Z(n4739));
Q_MX02 U4081 ( .S(oFill[0]), .A0(oData[302]), .A1(oData[238]), .Z(n4738));
Q_MX02 U4082 ( .S(oFill[0]), .A0(oData[301]), .A1(oData[237]), .Z(n4737));
Q_MX02 U4083 ( .S(oFill[0]), .A0(oData[300]), .A1(oData[236]), .Z(n4736));
Q_MX02 U4084 ( .S(oFill[0]), .A0(oData[299]), .A1(oData[235]), .Z(n4735));
Q_MX02 U4085 ( .S(oFill[0]), .A0(oData[298]), .A1(oData[234]), .Z(n4734));
Q_MX02 U4086 ( .S(oFill[0]), .A0(oData[297]), .A1(oData[233]), .Z(n4733));
Q_MX02 U4087 ( .S(oFill[0]), .A0(oData[296]), .A1(oData[232]), .Z(n4732));
Q_MX02 U4088 ( .S(oFill[0]), .A0(oData[295]), .A1(oData[231]), .Z(n4731));
Q_MX02 U4089 ( .S(oFill[0]), .A0(oData[294]), .A1(oData[230]), .Z(n4730));
Q_MX02 U4090 ( .S(oFill[0]), .A0(oData[293]), .A1(oData[229]), .Z(n4729));
Q_MX02 U4091 ( .S(oFill[0]), .A0(oData[292]), .A1(oData[228]), .Z(n4728));
Q_MX02 U4092 ( .S(oFill[0]), .A0(oData[291]), .A1(oData[227]), .Z(n4727));
Q_MX02 U4093 ( .S(oFill[0]), .A0(oData[290]), .A1(oData[226]), .Z(n4726));
Q_MX02 U4094 ( .S(oFill[0]), .A0(oData[289]), .A1(oData[225]), .Z(n4725));
Q_MX02 U4095 ( .S(oFill[0]), .A0(oData[288]), .A1(oData[224]), .Z(n4724));
Q_MX02 U4096 ( .S(oFill[0]), .A0(oData[287]), .A1(oData[223]), .Z(n4723));
Q_MX02 U4097 ( .S(oFill[0]), .A0(oData[286]), .A1(oData[222]), .Z(n4722));
Q_MX02 U4098 ( .S(oFill[0]), .A0(oData[285]), .A1(oData[221]), .Z(n4721));
Q_MX02 U4099 ( .S(oFill[0]), .A0(oData[284]), .A1(oData[220]), .Z(n4720));
Q_MX02 U4100 ( .S(oFill[0]), .A0(oData[283]), .A1(oData[219]), .Z(n4719));
Q_MX02 U4101 ( .S(oFill[0]), .A0(oData[282]), .A1(oData[218]), .Z(n4718));
Q_MX02 U4102 ( .S(oFill[0]), .A0(oData[281]), .A1(oData[217]), .Z(n4717));
Q_MX02 U4103 ( .S(oFill[0]), .A0(oData[280]), .A1(oData[216]), .Z(n4716));
Q_MX02 U4104 ( .S(oFill[0]), .A0(oData[279]), .A1(oData[215]), .Z(n4715));
Q_MX02 U4105 ( .S(oFill[0]), .A0(oData[278]), .A1(oData[214]), .Z(n4714));
Q_MX02 U4106 ( .S(oFill[0]), .A0(oData[277]), .A1(oData[213]), .Z(n4713));
Q_MX02 U4107 ( .S(oFill[0]), .A0(oData[276]), .A1(oData[212]), .Z(n4712));
Q_MX02 U4108 ( .S(oFill[0]), .A0(oData[275]), .A1(oData[211]), .Z(n4711));
Q_MX02 U4109 ( .S(oFill[0]), .A0(oData[274]), .A1(oData[210]), .Z(n4710));
Q_MX02 U4110 ( .S(oFill[0]), .A0(oData[273]), .A1(oData[209]), .Z(n4709));
Q_MX02 U4111 ( .S(oFill[0]), .A0(oData[272]), .A1(oData[208]), .Z(n4708));
Q_MX02 U4112 ( .S(oFill[0]), .A0(oData[271]), .A1(oData[207]), .Z(n4707));
Q_MX02 U4113 ( .S(oFill[0]), .A0(oData[270]), .A1(oData[206]), .Z(n4706));
Q_MX02 U4114 ( .S(oFill[0]), .A0(oData[269]), .A1(oData[205]), .Z(n4705));
Q_MX02 U4115 ( .S(oFill[0]), .A0(oData[268]), .A1(oData[204]), .Z(n4704));
Q_MX02 U4116 ( .S(oFill[0]), .A0(oData[267]), .A1(oData[203]), .Z(n4703));
Q_MX02 U4117 ( .S(oFill[0]), .A0(oData[266]), .A1(oData[202]), .Z(n4702));
Q_MX02 U4118 ( .S(oFill[0]), .A0(oData[265]), .A1(oData[201]), .Z(n4701));
Q_MX02 U4119 ( .S(oFill[0]), .A0(oData[264]), .A1(oData[200]), .Z(n4700));
Q_MX02 U4120 ( .S(oFill[0]), .A0(oData[263]), .A1(oData[199]), .Z(n4699));
Q_MX02 U4121 ( .S(oFill[0]), .A0(oData[262]), .A1(oData[198]), .Z(n4698));
Q_MX02 U4122 ( .S(oFill[0]), .A0(oData[261]), .A1(oData[197]), .Z(n4697));
Q_MX02 U4123 ( .S(oFill[0]), .A0(oData[260]), .A1(oData[196]), .Z(n4696));
Q_MX02 U4124 ( .S(oFill[0]), .A0(oData[259]), .A1(oData[195]), .Z(n4695));
Q_MX02 U4125 ( .S(oFill[0]), .A0(oData[258]), .A1(oData[194]), .Z(n4694));
Q_MX02 U4126 ( .S(oFill[0]), .A0(oData[257]), .A1(oData[193]), .Z(n4693));
Q_MX02 U4127 ( .S(oFill[0]), .A0(oData[256]), .A1(oData[192]), .Z(n4692));
Q_MX02 U4128 ( .S(oFill[0]), .A0(oData[255]), .A1(oData[191]), .Z(n4691));
Q_MX02 U4129 ( .S(oFill[0]), .A0(oData[254]), .A1(oData[190]), .Z(n4690));
Q_MX02 U4130 ( .S(oFill[0]), .A0(oData[253]), .A1(oData[189]), .Z(n4689));
Q_MX02 U4131 ( .S(oFill[0]), .A0(oData[252]), .A1(oData[188]), .Z(n4688));
Q_MX02 U4132 ( .S(oFill[0]), .A0(oData[251]), .A1(oData[187]), .Z(n4687));
Q_MX02 U4133 ( .S(oFill[0]), .A0(oData[250]), .A1(oData[186]), .Z(n4686));
Q_MX02 U4134 ( .S(oFill[0]), .A0(oData[249]), .A1(oData[185]), .Z(n4685));
Q_MX02 U4135 ( .S(oFill[0]), .A0(oData[248]), .A1(oData[184]), .Z(n4684));
Q_MX02 U4136 ( .S(oFill[0]), .A0(oData[247]), .A1(oData[183]), .Z(n4683));
Q_MX02 U4137 ( .S(oFill[0]), .A0(oData[246]), .A1(oData[182]), .Z(n4682));
Q_MX02 U4138 ( .S(oFill[0]), .A0(oData[245]), .A1(oData[181]), .Z(n4681));
Q_MX02 U4139 ( .S(oFill[0]), .A0(oData[244]), .A1(oData[180]), .Z(n4680));
Q_MX02 U4140 ( .S(oFill[0]), .A0(oData[243]), .A1(oData[179]), .Z(n4679));
Q_MX02 U4141 ( .S(oFill[0]), .A0(oData[242]), .A1(oData[178]), .Z(n4678));
Q_MX02 U4142 ( .S(oFill[0]), .A0(oData[241]), .A1(oData[177]), .Z(n4677));
Q_MX02 U4143 ( .S(oFill[0]), .A0(oData[240]), .A1(oData[176]), .Z(n4676));
Q_MX02 U4144 ( .S(oFill[0]), .A0(oData[239]), .A1(oData[175]), .Z(n4675));
Q_MX02 U4145 ( .S(oFill[0]), .A0(oData[238]), .A1(oData[174]), .Z(n4674));
Q_MX02 U4146 ( .S(oFill[0]), .A0(oData[237]), .A1(oData[173]), .Z(n4673));
Q_MX02 U4147 ( .S(oFill[0]), .A0(oData[236]), .A1(oData[172]), .Z(n4672));
Q_MX02 U4148 ( .S(oFill[0]), .A0(oData[235]), .A1(oData[171]), .Z(n4671));
Q_MX02 U4149 ( .S(oFill[0]), .A0(oData[234]), .A1(oData[170]), .Z(n4670));
Q_MX02 U4150 ( .S(oFill[0]), .A0(oData[233]), .A1(oData[169]), .Z(n4669));
Q_MX02 U4151 ( .S(oFill[0]), .A0(oData[232]), .A1(oData[168]), .Z(n4668));
Q_MX02 U4152 ( .S(oFill[0]), .A0(oData[231]), .A1(oData[167]), .Z(n4667));
Q_MX02 U4153 ( .S(oFill[0]), .A0(oData[230]), .A1(oData[166]), .Z(n4666));
Q_MX02 U4154 ( .S(oFill[0]), .A0(oData[229]), .A1(oData[165]), .Z(n4665));
Q_MX02 U4155 ( .S(oFill[0]), .A0(oData[228]), .A1(oData[164]), .Z(n4664));
Q_MX02 U4156 ( .S(oFill[0]), .A0(oData[227]), .A1(oData[163]), .Z(n4663));
Q_MX02 U4157 ( .S(oFill[0]), .A0(oData[226]), .A1(oData[162]), .Z(n4662));
Q_MX02 U4158 ( .S(oFill[0]), .A0(oData[225]), .A1(oData[161]), .Z(n4661));
Q_MX02 U4159 ( .S(oFill[0]), .A0(oData[224]), .A1(oData[160]), .Z(n4660));
Q_MX02 U4160 ( .S(oFill[0]), .A0(oData[223]), .A1(oData[159]), .Z(n4659));
Q_MX02 U4161 ( .S(oFill[0]), .A0(oData[222]), .A1(oData[158]), .Z(n4658));
Q_MX02 U4162 ( .S(oFill[0]), .A0(oData[221]), .A1(oData[157]), .Z(n4657));
Q_MX02 U4163 ( .S(oFill[0]), .A0(oData[220]), .A1(oData[156]), .Z(n4656));
Q_MX02 U4164 ( .S(oFill[0]), .A0(oData[219]), .A1(oData[155]), .Z(n4655));
Q_MX02 U4165 ( .S(oFill[0]), .A0(oData[218]), .A1(oData[154]), .Z(n4654));
Q_MX02 U4166 ( .S(oFill[0]), .A0(oData[217]), .A1(oData[153]), .Z(n4653));
Q_MX02 U4167 ( .S(oFill[0]), .A0(oData[216]), .A1(oData[152]), .Z(n4652));
Q_MX02 U4168 ( .S(oFill[0]), .A0(oData[215]), .A1(oData[151]), .Z(n4651));
Q_MX02 U4169 ( .S(oFill[0]), .A0(oData[214]), .A1(oData[150]), .Z(n4650));
Q_MX02 U4170 ( .S(oFill[0]), .A0(oData[213]), .A1(oData[149]), .Z(n4649));
Q_MX02 U4171 ( .S(oFill[0]), .A0(oData[212]), .A1(oData[148]), .Z(n4648));
Q_MX02 U4172 ( .S(oFill[0]), .A0(oData[211]), .A1(oData[147]), .Z(n4647));
Q_MX02 U4173 ( .S(oFill[0]), .A0(oData[210]), .A1(oData[146]), .Z(n4646));
Q_MX02 U4174 ( .S(oFill[0]), .A0(oData[209]), .A1(oData[145]), .Z(n4645));
Q_MX02 U4175 ( .S(oFill[0]), .A0(oData[208]), .A1(oData[144]), .Z(n4644));
Q_MX02 U4176 ( .S(oFill[0]), .A0(oData[207]), .A1(oData[143]), .Z(n4643));
Q_MX02 U4177 ( .S(oFill[0]), .A0(oData[206]), .A1(oData[142]), .Z(n4642));
Q_MX02 U4178 ( .S(oFill[0]), .A0(oData[205]), .A1(oData[141]), .Z(n4641));
Q_MX02 U4179 ( .S(oFill[0]), .A0(oData[204]), .A1(oData[140]), .Z(n4640));
Q_MX02 U4180 ( .S(oFill[0]), .A0(oData[203]), .A1(oData[139]), .Z(n4639));
Q_MX02 U4181 ( .S(oFill[0]), .A0(oData[202]), .A1(oData[138]), .Z(n4638));
Q_MX02 U4182 ( .S(oFill[0]), .A0(oData[201]), .A1(oData[137]), .Z(n4637));
Q_MX02 U4183 ( .S(oFill[0]), .A0(oData[200]), .A1(oData[136]), .Z(n4636));
Q_MX02 U4184 ( .S(oFill[0]), .A0(oData[199]), .A1(oData[135]), .Z(n4635));
Q_MX02 U4185 ( .S(oFill[0]), .A0(oData[198]), .A1(oData[134]), .Z(n4634));
Q_MX02 U4186 ( .S(oFill[0]), .A0(oData[197]), .A1(oData[133]), .Z(n4633));
Q_MX02 U4187 ( .S(oFill[0]), .A0(oData[196]), .A1(oData[132]), .Z(n4632));
Q_MX02 U4188 ( .S(oFill[0]), .A0(oData[195]), .A1(oData[131]), .Z(n4631));
Q_MX02 U4189 ( .S(oFill[0]), .A0(oData[194]), .A1(oData[130]), .Z(n4630));
Q_MX02 U4190 ( .S(oFill[0]), .A0(oData[193]), .A1(oData[129]), .Z(n4629));
Q_MX02 U4191 ( .S(oFill[0]), .A0(oData[192]), .A1(oData[128]), .Z(n4628));
Q_MX02 U4192 ( .S(oFill[0]), .A0(oData[191]), .A1(oData[127]), .Z(n4627));
Q_MX02 U4193 ( .S(oFill[0]), .A0(oData[190]), .A1(oData[126]), .Z(n4626));
Q_MX02 U4194 ( .S(oFill[0]), .A0(oData[189]), .A1(oData[125]), .Z(n4625));
Q_MX02 U4195 ( .S(oFill[0]), .A0(oData[188]), .A1(oData[124]), .Z(n4624));
Q_MX02 U4196 ( .S(oFill[0]), .A0(oData[187]), .A1(oData[123]), .Z(n4623));
Q_MX02 U4197 ( .S(oFill[0]), .A0(oData[186]), .A1(oData[122]), .Z(n4622));
Q_MX02 U4198 ( .S(oFill[0]), .A0(oData[185]), .A1(oData[121]), .Z(n4621));
Q_MX02 U4199 ( .S(oFill[0]), .A0(oData[184]), .A1(oData[120]), .Z(n4620));
Q_MX02 U4200 ( .S(oFill[0]), .A0(oData[183]), .A1(oData[119]), .Z(n4619));
Q_MX02 U4201 ( .S(oFill[0]), .A0(oData[182]), .A1(oData[118]), .Z(n4618));
Q_MX02 U4202 ( .S(oFill[0]), .A0(oData[181]), .A1(oData[117]), .Z(n4617));
Q_MX02 U4203 ( .S(oFill[0]), .A0(oData[180]), .A1(oData[116]), .Z(n4616));
Q_MX02 U4204 ( .S(oFill[0]), .A0(oData[179]), .A1(oData[115]), .Z(n4615));
Q_MX02 U4205 ( .S(oFill[0]), .A0(oData[178]), .A1(oData[114]), .Z(n4614));
Q_MX02 U4206 ( .S(oFill[0]), .A0(oData[177]), .A1(oData[113]), .Z(n4613));
Q_MX02 U4207 ( .S(oFill[0]), .A0(oData[176]), .A1(oData[112]), .Z(n4612));
Q_MX02 U4208 ( .S(oFill[0]), .A0(oData[175]), .A1(oData[111]), .Z(n4611));
Q_MX02 U4209 ( .S(oFill[0]), .A0(oData[174]), .A1(oData[110]), .Z(n4610));
Q_MX02 U4210 ( .S(oFill[0]), .A0(oData[173]), .A1(oData[109]), .Z(n4609));
Q_MX02 U4211 ( .S(oFill[0]), .A0(oData[172]), .A1(oData[108]), .Z(n4608));
Q_MX02 U4212 ( .S(oFill[0]), .A0(oData[171]), .A1(oData[107]), .Z(n4607));
Q_MX02 U4213 ( .S(oFill[0]), .A0(oData[170]), .A1(oData[106]), .Z(n4606));
Q_MX02 U4214 ( .S(oFill[0]), .A0(oData[169]), .A1(oData[105]), .Z(n4605));
Q_MX02 U4215 ( .S(oFill[0]), .A0(oData[168]), .A1(oData[104]), .Z(n4604));
Q_MX02 U4216 ( .S(oFill[0]), .A0(oData[167]), .A1(oData[103]), .Z(n4603));
Q_MX02 U4217 ( .S(oFill[0]), .A0(oData[166]), .A1(oData[102]), .Z(n4602));
Q_MX02 U4218 ( .S(oFill[0]), .A0(oData[165]), .A1(oData[101]), .Z(n4601));
Q_MX02 U4219 ( .S(oFill[0]), .A0(oData[164]), .A1(oData[100]), .Z(n4600));
Q_MX02 U4220 ( .S(oFill[0]), .A0(oData[163]), .A1(oData[99]), .Z(n4599));
Q_MX02 U4221 ( .S(oFill[0]), .A0(oData[162]), .A1(oData[98]), .Z(n4598));
Q_MX02 U4222 ( .S(oFill[0]), .A0(oData[161]), .A1(oData[97]), .Z(n4597));
Q_MX02 U4223 ( .S(oFill[0]), .A0(oData[160]), .A1(oData[96]), .Z(n4596));
Q_MX02 U4224 ( .S(oFill[0]), .A0(oData[159]), .A1(oData[95]), .Z(n4595));
Q_MX02 U4225 ( .S(oFill[0]), .A0(oData[158]), .A1(oData[94]), .Z(n4594));
Q_MX02 U4226 ( .S(oFill[0]), .A0(oData[157]), .A1(oData[93]), .Z(n4593));
Q_MX02 U4227 ( .S(oFill[0]), .A0(oData[156]), .A1(oData[92]), .Z(n4592));
Q_MX02 U4228 ( .S(oFill[0]), .A0(oData[155]), .A1(oData[91]), .Z(n4591));
Q_MX02 U4229 ( .S(oFill[0]), .A0(oData[154]), .A1(oData[90]), .Z(n4590));
Q_MX02 U4230 ( .S(oFill[0]), .A0(oData[153]), .A1(oData[89]), .Z(n4589));
Q_MX02 U4231 ( .S(oFill[0]), .A0(oData[152]), .A1(oData[88]), .Z(n4588));
Q_MX02 U4232 ( .S(oFill[0]), .A0(oData[151]), .A1(oData[87]), .Z(n4587));
Q_MX02 U4233 ( .S(oFill[0]), .A0(oData[150]), .A1(oData[86]), .Z(n4586));
Q_MX02 U4234 ( .S(oFill[0]), .A0(oData[149]), .A1(oData[85]), .Z(n4585));
Q_MX02 U4235 ( .S(oFill[0]), .A0(oData[148]), .A1(oData[84]), .Z(n4584));
Q_MX02 U4236 ( .S(oFill[0]), .A0(oData[147]), .A1(oData[83]), .Z(n4583));
Q_MX02 U4237 ( .S(oFill[0]), .A0(oData[146]), .A1(oData[82]), .Z(n4582));
Q_MX02 U4238 ( .S(oFill[0]), .A0(oData[145]), .A1(oData[81]), .Z(n4581));
Q_MX02 U4239 ( .S(oFill[0]), .A0(oData[144]), .A1(oData[80]), .Z(n4580));
Q_MX02 U4240 ( .S(oFill[0]), .A0(oData[143]), .A1(oData[79]), .Z(n4579));
Q_MX02 U4241 ( .S(oFill[0]), .A0(oData[142]), .A1(oData[78]), .Z(n4578));
Q_MX02 U4242 ( .S(oFill[0]), .A0(oData[141]), .A1(oData[77]), .Z(n4577));
Q_MX02 U4243 ( .S(oFill[0]), .A0(oData[140]), .A1(oData[76]), .Z(n4576));
Q_MX02 U4244 ( .S(oFill[0]), .A0(oData[139]), .A1(oData[75]), .Z(n4575));
Q_MX02 U4245 ( .S(oFill[0]), .A0(oData[138]), .A1(oData[74]), .Z(n4574));
Q_MX02 U4246 ( .S(oFill[0]), .A0(oData[137]), .A1(oData[73]), .Z(n4573));
Q_MX02 U4247 ( .S(oFill[0]), .A0(oData[136]), .A1(oData[72]), .Z(n4572));
Q_MX02 U4248 ( .S(oFill[0]), .A0(oData[135]), .A1(oData[71]), .Z(n4571));
Q_MX02 U4249 ( .S(oFill[0]), .A0(oData[134]), .A1(oData[70]), .Z(n4570));
Q_MX02 U4250 ( .S(oFill[0]), .A0(oData[133]), .A1(oData[69]), .Z(n4569));
Q_MX02 U4251 ( .S(oFill[0]), .A0(oData[132]), .A1(oData[68]), .Z(n4568));
Q_MX02 U4252 ( .S(oFill[0]), .A0(oData[131]), .A1(oData[67]), .Z(n4567));
Q_MX02 U4253 ( .S(oFill[0]), .A0(oData[130]), .A1(oData[66]), .Z(n4566));
Q_MX02 U4254 ( .S(oFill[0]), .A0(oData[129]), .A1(oData[65]), .Z(n4565));
Q_MX02 U4255 ( .S(oFill[0]), .A0(oData[128]), .A1(oData[64]), .Z(n4564));
Q_MX02 U4256 ( .S(oFill[0]), .A0(oData[127]), .A1(oData[63]), .Z(n4563));
Q_MX02 U4257 ( .S(oFill[0]), .A0(oData[126]), .A1(oData[62]), .Z(n4562));
Q_MX02 U4258 ( .S(oFill[0]), .A0(oData[125]), .A1(oData[61]), .Z(n4561));
Q_MX02 U4259 ( .S(oFill[0]), .A0(oData[124]), .A1(oData[60]), .Z(n4560));
Q_MX02 U4260 ( .S(oFill[0]), .A0(oData[123]), .A1(oData[59]), .Z(n4559));
Q_MX02 U4261 ( .S(oFill[0]), .A0(oData[122]), .A1(oData[58]), .Z(n4558));
Q_MX02 U4262 ( .S(oFill[0]), .A0(oData[121]), .A1(oData[57]), .Z(n4557));
Q_MX02 U4263 ( .S(oFill[0]), .A0(oData[120]), .A1(oData[56]), .Z(n4556));
Q_MX02 U4264 ( .S(oFill[0]), .A0(oData[119]), .A1(oData[55]), .Z(n4555));
Q_MX02 U4265 ( .S(oFill[0]), .A0(oData[118]), .A1(oData[54]), .Z(n4554));
Q_MX02 U4266 ( .S(oFill[0]), .A0(oData[117]), .A1(oData[53]), .Z(n4553));
Q_MX02 U4267 ( .S(oFill[0]), .A0(oData[116]), .A1(oData[52]), .Z(n4552));
Q_MX02 U4268 ( .S(oFill[0]), .A0(oData[115]), .A1(oData[51]), .Z(n4551));
Q_MX02 U4269 ( .S(oFill[0]), .A0(oData[114]), .A1(oData[50]), .Z(n4550));
Q_MX02 U4270 ( .S(oFill[0]), .A0(oData[113]), .A1(oData[49]), .Z(n4549));
Q_MX02 U4271 ( .S(oFill[0]), .A0(oData[112]), .A1(oData[48]), .Z(n4548));
Q_MX02 U4272 ( .S(oFill[0]), .A0(oData[111]), .A1(oData[47]), .Z(n4547));
Q_MX02 U4273 ( .S(oFill[0]), .A0(oData[110]), .A1(oData[46]), .Z(n4546));
Q_MX02 U4274 ( .S(oFill[0]), .A0(oData[109]), .A1(oData[45]), .Z(n4545));
Q_MX02 U4275 ( .S(oFill[0]), .A0(oData[108]), .A1(oData[44]), .Z(n4544));
Q_MX02 U4276 ( .S(oFill[0]), .A0(oData[107]), .A1(oData[43]), .Z(n4543));
Q_MX02 U4277 ( .S(oFill[0]), .A0(oData[106]), .A1(oData[42]), .Z(n4542));
Q_MX02 U4278 ( .S(oFill[0]), .A0(oData[105]), .A1(oData[41]), .Z(n4541));
Q_MX02 U4279 ( .S(oFill[0]), .A0(oData[104]), .A1(oData[40]), .Z(n4540));
Q_MX02 U4280 ( .S(oFill[0]), .A0(oData[103]), .A1(oData[39]), .Z(n4539));
Q_MX02 U4281 ( .S(oFill[0]), .A0(oData[102]), .A1(oData[38]), .Z(n4538));
Q_MX02 U4282 ( .S(oFill[0]), .A0(oData[101]), .A1(oData[37]), .Z(n4537));
Q_MX02 U4283 ( .S(oFill[0]), .A0(oData[100]), .A1(oData[36]), .Z(n4536));
Q_MX02 U4284 ( .S(oFill[0]), .A0(oData[99]), .A1(oData[35]), .Z(n4535));
Q_MX02 U4285 ( .S(oFill[0]), .A0(oData[98]), .A1(oData[34]), .Z(n4534));
Q_MX02 U4286 ( .S(oFill[0]), .A0(oData[97]), .A1(oData[33]), .Z(n4533));
Q_MX02 U4287 ( .S(oFill[0]), .A0(oData[96]), .A1(oData[32]), .Z(n4532));
Q_MX02 U4288 ( .S(oFill[0]), .A0(oData[95]), .A1(oData[31]), .Z(n4531));
Q_MX02 U4289 ( .S(oFill[0]), .A0(oData[94]), .A1(oData[30]), .Z(n4530));
Q_MX02 U4290 ( .S(oFill[0]), .A0(oData[93]), .A1(oData[29]), .Z(n4529));
Q_MX02 U4291 ( .S(oFill[0]), .A0(oData[92]), .A1(oData[28]), .Z(n4528));
Q_MX02 U4292 ( .S(oFill[0]), .A0(oData[91]), .A1(oData[27]), .Z(n4527));
Q_MX02 U4293 ( .S(oFill[0]), .A0(oData[90]), .A1(oData[26]), .Z(n4526));
Q_MX02 U4294 ( .S(oFill[0]), .A0(oData[89]), .A1(oData[25]), .Z(n4525));
Q_MX02 U4295 ( .S(oFill[0]), .A0(oData[88]), .A1(oData[24]), .Z(n4524));
Q_MX02 U4296 ( .S(oFill[0]), .A0(oData[87]), .A1(oData[23]), .Z(n4523));
Q_MX02 U4297 ( .S(oFill[0]), .A0(oData[86]), .A1(oData[22]), .Z(n4522));
Q_MX02 U4298 ( .S(oFill[0]), .A0(oData[85]), .A1(oData[21]), .Z(n4521));
Q_MX02 U4299 ( .S(oFill[0]), .A0(oData[84]), .A1(oData[20]), .Z(n4520));
Q_MX02 U4300 ( .S(oFill[0]), .A0(oData[83]), .A1(oData[19]), .Z(n4519));
Q_MX02 U4301 ( .S(oFill[0]), .A0(oData[82]), .A1(oData[18]), .Z(n4518));
Q_MX02 U4302 ( .S(oFill[0]), .A0(oData[81]), .A1(oData[17]), .Z(n4517));
Q_MX02 U4303 ( .S(oFill[0]), .A0(oData[80]), .A1(oData[16]), .Z(n4516));
Q_MX02 U4304 ( .S(oFill[0]), .A0(oData[79]), .A1(oData[15]), .Z(n4515));
Q_MX02 U4305 ( .S(oFill[0]), .A0(oData[78]), .A1(oData[14]), .Z(n4514));
Q_MX02 U4306 ( .S(oFill[0]), .A0(oData[77]), .A1(oData[13]), .Z(n4513));
Q_MX02 U4307 ( .S(oFill[0]), .A0(oData[76]), .A1(oData[12]), .Z(n4512));
Q_MX02 U4308 ( .S(oFill[0]), .A0(oData[75]), .A1(oData[11]), .Z(n4511));
Q_MX02 U4309 ( .S(oFill[0]), .A0(oData[74]), .A1(oData[10]), .Z(n4510));
Q_MX02 U4310 ( .S(oFill[0]), .A0(oData[73]), .A1(oData[9]), .Z(n4509));
Q_MX02 U4311 ( .S(oFill[0]), .A0(oData[72]), .A1(oData[8]), .Z(n4508));
Q_MX02 U4312 ( .S(oFill[0]), .A0(oData[71]), .A1(oData[7]), .Z(n4507));
Q_MX02 U4313 ( .S(oFill[0]), .A0(oData[70]), .A1(oData[6]), .Z(n4506));
Q_MX02 U4314 ( .S(oFill[0]), .A0(oData[69]), .A1(oData[5]), .Z(n4505));
Q_MX02 U4315 ( .S(oFill[0]), .A0(oData[68]), .A1(oData[4]), .Z(n4504));
Q_MX02 U4316 ( .S(oFill[0]), .A0(oData[67]), .A1(oData[3]), .Z(n4503));
Q_MX02 U4317 ( .S(oFill[0]), .A0(oData[66]), .A1(oData[2]), .Z(n4502));
Q_MX02 U4318 ( .S(oFill[0]), .A0(oData[65]), .A1(oData[1]), .Z(n4501));
Q_MX02 U4319 ( .S(oFill[0]), .A0(oData[64]), .A1(oData[0]), .Z(n4500));
Q_INV U4320 ( .A(oFill[0]), .Z(n4499));
Q_AN02 U4321 ( .A0(n4499), .A1(oData[63]), .Z(n4498));
Q_AN02 U4322 ( .A0(n4499), .A1(oData[62]), .Z(n4497));
Q_AN02 U4323 ( .A0(n4499), .A1(oData[61]), .Z(n4496));
Q_AN02 U4324 ( .A0(n4499), .A1(oData[60]), .Z(n4495));
Q_AN02 U4325 ( .A0(n4499), .A1(oData[59]), .Z(n4494));
Q_AN02 U4326 ( .A0(n4499), .A1(oData[58]), .Z(n4493));
Q_AN02 U4327 ( .A0(n4499), .A1(oData[57]), .Z(n4492));
Q_AN02 U4328 ( .A0(n4499), .A1(oData[56]), .Z(n4491));
Q_AN02 U4329 ( .A0(n4499), .A1(oData[55]), .Z(n4490));
Q_AN02 U4330 ( .A0(n4499), .A1(oData[54]), .Z(n4489));
Q_AN02 U4331 ( .A0(n4499), .A1(oData[53]), .Z(n4488));
Q_AN02 U4332 ( .A0(n4499), .A1(oData[52]), .Z(n4487));
Q_AN02 U4333 ( .A0(n4499), .A1(oData[51]), .Z(n4486));
Q_AN02 U4334 ( .A0(n4499), .A1(oData[50]), .Z(n4485));
Q_AN02 U4335 ( .A0(n4499), .A1(oData[49]), .Z(n4484));
Q_AN02 U4336 ( .A0(n4499), .A1(oData[48]), .Z(n4483));
Q_AN02 U4337 ( .A0(n4499), .A1(oData[47]), .Z(n4482));
Q_AN02 U4338 ( .A0(n4499), .A1(oData[46]), .Z(n4481));
Q_AN02 U4339 ( .A0(n4499), .A1(oData[45]), .Z(n4480));
Q_AN02 U4340 ( .A0(n4499), .A1(oData[44]), .Z(n4479));
Q_AN02 U4341 ( .A0(n4499), .A1(oData[43]), .Z(n4478));
Q_AN02 U4342 ( .A0(n4499), .A1(oData[42]), .Z(n4477));
Q_AN02 U4343 ( .A0(n4499), .A1(oData[41]), .Z(n4476));
Q_AN02 U4344 ( .A0(n4499), .A1(oData[40]), .Z(n4475));
Q_AN02 U4345 ( .A0(n4499), .A1(oData[39]), .Z(n4474));
Q_AN02 U4346 ( .A0(n4499), .A1(oData[38]), .Z(n4473));
Q_AN02 U4347 ( .A0(n4499), .A1(oData[37]), .Z(n4472));
Q_AN02 U4348 ( .A0(n4499), .A1(oData[36]), .Z(n4471));
Q_AN02 U4349 ( .A0(n4499), .A1(oData[35]), .Z(n4470));
Q_AN02 U4350 ( .A0(n4499), .A1(oData[34]), .Z(n4469));
Q_AN02 U4351 ( .A0(n4499), .A1(oData[33]), .Z(n4468));
Q_AN02 U4352 ( .A0(n4499), .A1(oData[32]), .Z(n4467));
Q_AN02 U4353 ( .A0(n4499), .A1(oData[31]), .Z(n4466));
Q_AN02 U4354 ( .A0(n4499), .A1(oData[30]), .Z(n4465));
Q_AN02 U4355 ( .A0(n4499), .A1(oData[29]), .Z(n4464));
Q_AN02 U4356 ( .A0(n4499), .A1(oData[28]), .Z(n4463));
Q_AN02 U4357 ( .A0(n4499), .A1(oData[27]), .Z(n4462));
Q_AN02 U4358 ( .A0(n4499), .A1(oData[26]), .Z(n4461));
Q_AN02 U4359 ( .A0(n4499), .A1(oData[25]), .Z(n4460));
Q_AN02 U4360 ( .A0(n4499), .A1(oData[24]), .Z(n4459));
Q_AN02 U4361 ( .A0(n4499), .A1(oData[23]), .Z(n4458));
Q_AN02 U4362 ( .A0(n4499), .A1(oData[22]), .Z(n4457));
Q_AN02 U4363 ( .A0(n4499), .A1(oData[21]), .Z(n4456));
Q_AN02 U4364 ( .A0(n4499), .A1(oData[20]), .Z(n4455));
Q_AN02 U4365 ( .A0(n4499), .A1(oData[19]), .Z(n4454));
Q_AN02 U4366 ( .A0(n4499), .A1(oData[18]), .Z(n4453));
Q_AN02 U4367 ( .A0(n4499), .A1(oData[17]), .Z(n4452));
Q_AN02 U4368 ( .A0(n4499), .A1(oData[16]), .Z(n4451));
Q_AN02 U4369 ( .A0(n4499), .A1(oData[15]), .Z(n4450));
Q_AN02 U4370 ( .A0(n4499), .A1(oData[14]), .Z(n4449));
Q_AN02 U4371 ( .A0(n4499), .A1(oData[13]), .Z(n4448));
Q_AN02 U4372 ( .A0(n4499), .A1(oData[12]), .Z(n4447));
Q_AN02 U4373 ( .A0(n4499), .A1(oData[11]), .Z(n4446));
Q_AN02 U4374 ( .A0(n4499), .A1(oData[10]), .Z(n4445));
Q_AN02 U4375 ( .A0(n4499), .A1(oData[9]), .Z(n4444));
Q_AN02 U4376 ( .A0(n4499), .A1(oData[8]), .Z(n4443));
Q_AN02 U4377 ( .A0(n4499), .A1(oData[7]), .Z(n4442));
Q_AN02 U4378 ( .A0(n4499), .A1(oData[6]), .Z(n4441));
Q_AN02 U4379 ( .A0(n4499), .A1(oData[5]), .Z(n4440));
Q_AN02 U4380 ( .A0(n4499), .A1(oData[4]), .Z(n4439));
Q_AN02 U4381 ( .A0(n4499), .A1(oData[3]), .Z(n4438));
Q_AN02 U4382 ( .A0(n4499), .A1(oData[2]), .Z(n4437));
Q_AN02 U4383 ( .A0(n4499), .A1(oData[1]), .Z(n4436));
Q_AN02 U4384 ( .A0(n4499), .A1(oData[0]), .Z(n4435));
Q_AN02 U4385 ( .A0(oFill[1]), .A1(n5011), .Z(n4434));
Q_AN02 U4386 ( .A0(oFill[1]), .A1(n5010), .Z(n4433));
Q_AN02 U4387 ( .A0(oFill[1]), .A1(n5009), .Z(n4432));
Q_AN02 U4388 ( .A0(oFill[1]), .A1(n5008), .Z(n4431));
Q_AN02 U4389 ( .A0(oFill[1]), .A1(n5007), .Z(n4430));
Q_AN02 U4390 ( .A0(oFill[1]), .A1(n5006), .Z(n4429));
Q_AN02 U4391 ( .A0(oFill[1]), .A1(n5005), .Z(n4428));
Q_AN02 U4392 ( .A0(oFill[1]), .A1(n5004), .Z(n4427));
Q_AN02 U4393 ( .A0(oFill[1]), .A1(n5003), .Z(n4426));
Q_AN02 U4394 ( .A0(oFill[1]), .A1(n5002), .Z(n4425));
Q_AN02 U4395 ( .A0(oFill[1]), .A1(n5001), .Z(n4424));
Q_AN02 U4396 ( .A0(oFill[1]), .A1(n5000), .Z(n4423));
Q_AN02 U4397 ( .A0(oFill[1]), .A1(n4999), .Z(n4422));
Q_AN02 U4398 ( .A0(oFill[1]), .A1(n4998), .Z(n4421));
Q_AN02 U4399 ( .A0(oFill[1]), .A1(n4997), .Z(n4420));
Q_AN02 U4400 ( .A0(oFill[1]), .A1(n4996), .Z(n4419));
Q_AN02 U4401 ( .A0(oFill[1]), .A1(n4995), .Z(n4418));
Q_AN02 U4402 ( .A0(oFill[1]), .A1(n4994), .Z(n4417));
Q_AN02 U4403 ( .A0(oFill[1]), .A1(n4993), .Z(n4416));
Q_AN02 U4404 ( .A0(oFill[1]), .A1(n4992), .Z(n4415));
Q_AN02 U4405 ( .A0(oFill[1]), .A1(n4991), .Z(n4414));
Q_AN02 U4406 ( .A0(oFill[1]), .A1(n4990), .Z(n4413));
Q_AN02 U4407 ( .A0(oFill[1]), .A1(n4989), .Z(n4412));
Q_AN02 U4408 ( .A0(oFill[1]), .A1(n4988), .Z(n4411));
Q_AN02 U4409 ( .A0(oFill[1]), .A1(n4987), .Z(n4410));
Q_AN02 U4410 ( .A0(oFill[1]), .A1(n4986), .Z(n4409));
Q_AN02 U4411 ( .A0(oFill[1]), .A1(n4985), .Z(n4408));
Q_AN02 U4412 ( .A0(oFill[1]), .A1(n4984), .Z(n4407));
Q_AN02 U4413 ( .A0(oFill[1]), .A1(n4983), .Z(n4406));
Q_AN02 U4414 ( .A0(oFill[1]), .A1(n4982), .Z(n4405));
Q_AN02 U4415 ( .A0(oFill[1]), .A1(n4981), .Z(n4404));
Q_AN02 U4416 ( .A0(oFill[1]), .A1(n4980), .Z(n4403));
Q_AN02 U4417 ( .A0(oFill[1]), .A1(n4979), .Z(n4402));
Q_AN02 U4418 ( .A0(oFill[1]), .A1(n4978), .Z(n4401));
Q_AN02 U4419 ( .A0(oFill[1]), .A1(n4977), .Z(n4400));
Q_AN02 U4420 ( .A0(oFill[1]), .A1(n4976), .Z(n4399));
Q_AN02 U4421 ( .A0(oFill[1]), .A1(n4975), .Z(n4398));
Q_AN02 U4422 ( .A0(oFill[1]), .A1(n4974), .Z(n4397));
Q_AN02 U4423 ( .A0(oFill[1]), .A1(n4973), .Z(n4396));
Q_AN02 U4424 ( .A0(oFill[1]), .A1(n4972), .Z(n4395));
Q_AN02 U4425 ( .A0(oFill[1]), .A1(n4971), .Z(n4394));
Q_AN02 U4426 ( .A0(oFill[1]), .A1(n4970), .Z(n4393));
Q_AN02 U4427 ( .A0(oFill[1]), .A1(n4969), .Z(n4392));
Q_AN02 U4428 ( .A0(oFill[1]), .A1(n4968), .Z(n4391));
Q_AN02 U4429 ( .A0(oFill[1]), .A1(n4967), .Z(n4390));
Q_AN02 U4430 ( .A0(oFill[1]), .A1(n4966), .Z(n4389));
Q_AN02 U4431 ( .A0(oFill[1]), .A1(n4965), .Z(n4388));
Q_AN02 U4432 ( .A0(oFill[1]), .A1(n4964), .Z(n4387));
Q_AN02 U4433 ( .A0(oFill[1]), .A1(n4963), .Z(n4386));
Q_AN02 U4434 ( .A0(oFill[1]), .A1(n4962), .Z(n4385));
Q_AN02 U4435 ( .A0(oFill[1]), .A1(n4961), .Z(n4384));
Q_AN02 U4436 ( .A0(oFill[1]), .A1(n4960), .Z(n4383));
Q_AN02 U4437 ( .A0(oFill[1]), .A1(n4959), .Z(n4382));
Q_AN02 U4438 ( .A0(oFill[1]), .A1(n4958), .Z(n4381));
Q_AN02 U4439 ( .A0(oFill[1]), .A1(n4957), .Z(n4380));
Q_AN02 U4440 ( .A0(oFill[1]), .A1(n4956), .Z(n4379));
Q_AN02 U4441 ( .A0(oFill[1]), .A1(n4955), .Z(n4378));
Q_AN02 U4442 ( .A0(oFill[1]), .A1(n4954), .Z(n4377));
Q_AN02 U4443 ( .A0(oFill[1]), .A1(n4953), .Z(n4376));
Q_AN02 U4444 ( .A0(oFill[1]), .A1(n4952), .Z(n4375));
Q_AN02 U4445 ( .A0(oFill[1]), .A1(n4951), .Z(n4374));
Q_AN02 U4446 ( .A0(oFill[1]), .A1(n4950), .Z(n4373));
Q_AN02 U4447 ( .A0(oFill[1]), .A1(n4949), .Z(n4372));
Q_AN02 U4448 ( .A0(oFill[1]), .A1(n4948), .Z(n4371));
Q_AN02 U4449 ( .A0(oFill[1]), .A1(n4947), .Z(n4370));
Q_AN02 U4450 ( .A0(oFill[1]), .A1(n4946), .Z(n4369));
Q_AN02 U4451 ( .A0(oFill[1]), .A1(n4945), .Z(n4368));
Q_AN02 U4452 ( .A0(oFill[1]), .A1(n4944), .Z(n4367));
Q_AN02 U4453 ( .A0(oFill[1]), .A1(n4943), .Z(n4366));
Q_AN02 U4454 ( .A0(oFill[1]), .A1(n4942), .Z(n4365));
Q_AN02 U4455 ( .A0(oFill[1]), .A1(n4941), .Z(n4364));
Q_AN02 U4456 ( .A0(oFill[1]), .A1(n4940), .Z(n4363));
Q_AN02 U4457 ( .A0(oFill[1]), .A1(n4939), .Z(n4362));
Q_AN02 U4458 ( .A0(oFill[1]), .A1(n4938), .Z(n4361));
Q_AN02 U4459 ( .A0(oFill[1]), .A1(n4937), .Z(n4360));
Q_AN02 U4460 ( .A0(oFill[1]), .A1(n4936), .Z(n4359));
Q_AN02 U4461 ( .A0(oFill[1]), .A1(n4935), .Z(n4358));
Q_AN02 U4462 ( .A0(oFill[1]), .A1(n4934), .Z(n4357));
Q_AN02 U4463 ( .A0(oFill[1]), .A1(n4933), .Z(n4356));
Q_AN02 U4464 ( .A0(oFill[1]), .A1(n4932), .Z(n4355));
Q_AN02 U4465 ( .A0(oFill[1]), .A1(n4931), .Z(n4354));
Q_AN02 U4466 ( .A0(oFill[1]), .A1(n4930), .Z(n4353));
Q_AN02 U4467 ( .A0(oFill[1]), .A1(n4929), .Z(n4352));
Q_AN02 U4468 ( .A0(oFill[1]), .A1(n4928), .Z(n4351));
Q_AN02 U4469 ( .A0(oFill[1]), .A1(n4927), .Z(n4350));
Q_AN02 U4470 ( .A0(oFill[1]), .A1(n4926), .Z(n4349));
Q_AN02 U4471 ( .A0(oFill[1]), .A1(n4925), .Z(n4348));
Q_AN02 U4472 ( .A0(oFill[1]), .A1(n4924), .Z(n4347));
Q_AN02 U4473 ( .A0(oFill[1]), .A1(n4923), .Z(n4346));
Q_AN02 U4474 ( .A0(oFill[1]), .A1(n4922), .Z(n4345));
Q_AN02 U4475 ( .A0(oFill[1]), .A1(n4921), .Z(n4344));
Q_AN02 U4476 ( .A0(oFill[1]), .A1(n4920), .Z(n4343));
Q_AN02 U4477 ( .A0(oFill[1]), .A1(n4919), .Z(n4342));
Q_AN02 U4478 ( .A0(oFill[1]), .A1(n4918), .Z(n4341));
Q_AN02 U4479 ( .A0(oFill[1]), .A1(n4917), .Z(n4340));
Q_AN02 U4480 ( .A0(oFill[1]), .A1(n4916), .Z(n4339));
Q_AN02 U4481 ( .A0(oFill[1]), .A1(n4915), .Z(n4338));
Q_AN02 U4482 ( .A0(oFill[1]), .A1(n4914), .Z(n4337));
Q_AN02 U4483 ( .A0(oFill[1]), .A1(n4913), .Z(n4336));
Q_AN02 U4484 ( .A0(oFill[1]), .A1(n4912), .Z(n4335));
Q_AN02 U4485 ( .A0(oFill[1]), .A1(n4911), .Z(n4334));
Q_AN02 U4486 ( .A0(oFill[1]), .A1(n4910), .Z(n4333));
Q_AN02 U4487 ( .A0(oFill[1]), .A1(n4909), .Z(n4332));
Q_AN02 U4488 ( .A0(oFill[1]), .A1(n4908), .Z(n4331));
Q_AN02 U4489 ( .A0(oFill[1]), .A1(n4907), .Z(n4330));
Q_AN02 U4490 ( .A0(oFill[1]), .A1(n4906), .Z(n4329));
Q_AN02 U4491 ( .A0(oFill[1]), .A1(n4905), .Z(n4328));
Q_AN02 U4492 ( .A0(oFill[1]), .A1(n4904), .Z(n4327));
Q_AN02 U4493 ( .A0(oFill[1]), .A1(n4903), .Z(n4326));
Q_AN02 U4494 ( .A0(oFill[1]), .A1(n4902), .Z(n4325));
Q_AN02 U4495 ( .A0(oFill[1]), .A1(n4901), .Z(n4324));
Q_AN02 U4496 ( .A0(oFill[1]), .A1(n4900), .Z(n4323));
Q_AN02 U4497 ( .A0(oFill[1]), .A1(n4899), .Z(n4322));
Q_AN02 U4498 ( .A0(oFill[1]), .A1(n4898), .Z(n4321));
Q_AN02 U4499 ( .A0(oFill[1]), .A1(n4897), .Z(n4320));
Q_AN02 U4500 ( .A0(oFill[1]), .A1(n4896), .Z(n4319));
Q_AN02 U4501 ( .A0(oFill[1]), .A1(n4895), .Z(n4318));
Q_AN02 U4502 ( .A0(oFill[1]), .A1(n4894), .Z(n4317));
Q_AN02 U4503 ( .A0(oFill[1]), .A1(n4893), .Z(n4316));
Q_AN02 U4504 ( .A0(oFill[1]), .A1(n4892), .Z(n4315));
Q_AN02 U4505 ( .A0(oFill[1]), .A1(n4891), .Z(n4314));
Q_AN02 U4506 ( .A0(oFill[1]), .A1(n4890), .Z(n4313));
Q_AN02 U4507 ( .A0(oFill[1]), .A1(n4889), .Z(n4312));
Q_AN02 U4508 ( .A0(oFill[1]), .A1(n4888), .Z(n4311));
Q_AN02 U4509 ( .A0(oFill[1]), .A1(n4887), .Z(n4310));
Q_AN02 U4510 ( .A0(oFill[1]), .A1(n4886), .Z(n4309));
Q_AN02 U4511 ( .A0(oFill[1]), .A1(n4885), .Z(n4308));
Q_AN02 U4512 ( .A0(oFill[1]), .A1(n4884), .Z(n4307));
Q_MX02 U4513 ( .S(oFill[1]), .A0(n5011), .A1(n4883), .Z(n4306));
Q_MX02 U4514 ( .S(oFill[1]), .A0(n5010), .A1(n4882), .Z(n4305));
Q_MX02 U4515 ( .S(oFill[1]), .A0(n5009), .A1(n4881), .Z(n4304));
Q_MX02 U4516 ( .S(oFill[1]), .A0(n5008), .A1(n4880), .Z(n4303));
Q_MX02 U4517 ( .S(oFill[1]), .A0(n5007), .A1(n4879), .Z(n4302));
Q_MX02 U4518 ( .S(oFill[1]), .A0(n5006), .A1(n4878), .Z(n4301));
Q_MX02 U4519 ( .S(oFill[1]), .A0(n5005), .A1(n4877), .Z(n4300));
Q_MX02 U4520 ( .S(oFill[1]), .A0(n5004), .A1(n4876), .Z(n4299));
Q_MX02 U4521 ( .S(oFill[1]), .A0(n5003), .A1(n4875), .Z(n4298));
Q_MX02 U4522 ( .S(oFill[1]), .A0(n5002), .A1(n4874), .Z(n4297));
Q_MX02 U4523 ( .S(oFill[1]), .A0(n5001), .A1(n4873), .Z(n4296));
Q_MX02 U4524 ( .S(oFill[1]), .A0(n5000), .A1(n4872), .Z(n4295));
Q_MX02 U4525 ( .S(oFill[1]), .A0(n4999), .A1(n4871), .Z(n4294));
Q_MX02 U4526 ( .S(oFill[1]), .A0(n4998), .A1(n4870), .Z(n4293));
Q_MX02 U4527 ( .S(oFill[1]), .A0(n4997), .A1(n4869), .Z(n4292));
Q_MX02 U4528 ( .S(oFill[1]), .A0(n4996), .A1(n4868), .Z(n4291));
Q_MX02 U4529 ( .S(oFill[1]), .A0(n4995), .A1(n4867), .Z(n4290));
Q_MX02 U4530 ( .S(oFill[1]), .A0(n4994), .A1(n4866), .Z(n4289));
Q_MX02 U4531 ( .S(oFill[1]), .A0(n4993), .A1(n4865), .Z(n4288));
Q_MX02 U4532 ( .S(oFill[1]), .A0(n4992), .A1(n4864), .Z(n4287));
Q_MX02 U4533 ( .S(oFill[1]), .A0(n4991), .A1(n4863), .Z(n4286));
Q_MX02 U4534 ( .S(oFill[1]), .A0(n4990), .A1(n4862), .Z(n4285));
Q_MX02 U4535 ( .S(oFill[1]), .A0(n4989), .A1(n4861), .Z(n4284));
Q_MX02 U4536 ( .S(oFill[1]), .A0(n4988), .A1(n4860), .Z(n4283));
Q_MX02 U4537 ( .S(oFill[1]), .A0(n4987), .A1(n4859), .Z(n4282));
Q_MX02 U4538 ( .S(oFill[1]), .A0(n4986), .A1(n4858), .Z(n4281));
Q_MX02 U4539 ( .S(oFill[1]), .A0(n4985), .A1(n4857), .Z(n4280));
Q_MX02 U4540 ( .S(oFill[1]), .A0(n4984), .A1(n4856), .Z(n4279));
Q_MX02 U4541 ( .S(oFill[1]), .A0(n4983), .A1(n4855), .Z(n4278));
Q_MX02 U4542 ( .S(oFill[1]), .A0(n4982), .A1(n4854), .Z(n4277));
Q_MX02 U4543 ( .S(oFill[1]), .A0(n4981), .A1(n4853), .Z(n4276));
Q_MX02 U4544 ( .S(oFill[1]), .A0(n4980), .A1(n4852), .Z(n4275));
Q_MX02 U4545 ( .S(oFill[1]), .A0(n4979), .A1(n4851), .Z(n4274));
Q_MX02 U4546 ( .S(oFill[1]), .A0(n4978), .A1(n4850), .Z(n4273));
Q_MX02 U4547 ( .S(oFill[1]), .A0(n4977), .A1(n4849), .Z(n4272));
Q_MX02 U4548 ( .S(oFill[1]), .A0(n4976), .A1(n4848), .Z(n4271));
Q_MX02 U4549 ( .S(oFill[1]), .A0(n4975), .A1(n4847), .Z(n4270));
Q_MX02 U4550 ( .S(oFill[1]), .A0(n4974), .A1(n4846), .Z(n4269));
Q_MX02 U4551 ( .S(oFill[1]), .A0(n4973), .A1(n4845), .Z(n4268));
Q_MX02 U4552 ( .S(oFill[1]), .A0(n4972), .A1(n4844), .Z(n4267));
Q_MX02 U4553 ( .S(oFill[1]), .A0(n4971), .A1(n4843), .Z(n4266));
Q_MX02 U4554 ( .S(oFill[1]), .A0(n4970), .A1(n4842), .Z(n4265));
Q_MX02 U4555 ( .S(oFill[1]), .A0(n4969), .A1(n4841), .Z(n4264));
Q_MX02 U4556 ( .S(oFill[1]), .A0(n4968), .A1(n4840), .Z(n4263));
Q_MX02 U4557 ( .S(oFill[1]), .A0(n4967), .A1(n4839), .Z(n4262));
Q_MX02 U4558 ( .S(oFill[1]), .A0(n4966), .A1(n4838), .Z(n4261));
Q_MX02 U4559 ( .S(oFill[1]), .A0(n4965), .A1(n4837), .Z(n4260));
Q_MX02 U4560 ( .S(oFill[1]), .A0(n4964), .A1(n4836), .Z(n4259));
Q_MX02 U4561 ( .S(oFill[1]), .A0(n4963), .A1(n4835), .Z(n4258));
Q_MX02 U4562 ( .S(oFill[1]), .A0(n4962), .A1(n4834), .Z(n4257));
Q_MX02 U4563 ( .S(oFill[1]), .A0(n4961), .A1(n4833), .Z(n4256));
Q_MX02 U4564 ( .S(oFill[1]), .A0(n4960), .A1(n4832), .Z(n4255));
Q_MX02 U4565 ( .S(oFill[1]), .A0(n4959), .A1(n4831), .Z(n4254));
Q_MX02 U4566 ( .S(oFill[1]), .A0(n4958), .A1(n4830), .Z(n4253));
Q_MX02 U4567 ( .S(oFill[1]), .A0(n4957), .A1(n4829), .Z(n4252));
Q_MX02 U4568 ( .S(oFill[1]), .A0(n4956), .A1(n4828), .Z(n4251));
Q_MX02 U4569 ( .S(oFill[1]), .A0(n4955), .A1(n4827), .Z(n4250));
Q_MX02 U4570 ( .S(oFill[1]), .A0(n4954), .A1(n4826), .Z(n4249));
Q_MX02 U4571 ( .S(oFill[1]), .A0(n4953), .A1(n4825), .Z(n4248));
Q_MX02 U4572 ( .S(oFill[1]), .A0(n4952), .A1(n4824), .Z(n4247));
Q_MX02 U4573 ( .S(oFill[1]), .A0(n4951), .A1(n4823), .Z(n4246));
Q_MX02 U4574 ( .S(oFill[1]), .A0(n4950), .A1(n4822), .Z(n4245));
Q_MX02 U4575 ( .S(oFill[1]), .A0(n4949), .A1(n4821), .Z(n4244));
Q_MX02 U4576 ( .S(oFill[1]), .A0(n4948), .A1(n4820), .Z(n4243));
Q_MX02 U4577 ( .S(oFill[1]), .A0(n4947), .A1(n4819), .Z(n4242));
Q_MX02 U4578 ( .S(oFill[1]), .A0(n4946), .A1(n4818), .Z(n4241));
Q_MX02 U4579 ( .S(oFill[1]), .A0(n4945), .A1(n4817), .Z(n4240));
Q_MX02 U4580 ( .S(oFill[1]), .A0(n4944), .A1(n4816), .Z(n4239));
Q_MX02 U4581 ( .S(oFill[1]), .A0(n4943), .A1(n4815), .Z(n4238));
Q_MX02 U4582 ( .S(oFill[1]), .A0(n4942), .A1(n4814), .Z(n4237));
Q_MX02 U4583 ( .S(oFill[1]), .A0(n4941), .A1(n4813), .Z(n4236));
Q_MX02 U4584 ( .S(oFill[1]), .A0(n4940), .A1(n4812), .Z(n4235));
Q_MX02 U4585 ( .S(oFill[1]), .A0(n4939), .A1(n4811), .Z(n4234));
Q_MX02 U4586 ( .S(oFill[1]), .A0(n4938), .A1(n4810), .Z(n4233));
Q_MX02 U4587 ( .S(oFill[1]), .A0(n4937), .A1(n4809), .Z(n4232));
Q_MX02 U4588 ( .S(oFill[1]), .A0(n4936), .A1(n4808), .Z(n4231));
Q_MX02 U4589 ( .S(oFill[1]), .A0(n4935), .A1(n4807), .Z(n4230));
Q_MX02 U4590 ( .S(oFill[1]), .A0(n4934), .A1(n4806), .Z(n4229));
Q_MX02 U4591 ( .S(oFill[1]), .A0(n4933), .A1(n4805), .Z(n4228));
Q_MX02 U4592 ( .S(oFill[1]), .A0(n4932), .A1(n4804), .Z(n4227));
Q_MX02 U4593 ( .S(oFill[1]), .A0(n4931), .A1(n4803), .Z(n4226));
Q_MX02 U4594 ( .S(oFill[1]), .A0(n4930), .A1(n4802), .Z(n4225));
Q_MX02 U4595 ( .S(oFill[1]), .A0(n4929), .A1(n4801), .Z(n4224));
Q_MX02 U4596 ( .S(oFill[1]), .A0(n4928), .A1(n4800), .Z(n4223));
Q_MX02 U4597 ( .S(oFill[1]), .A0(n4927), .A1(n4799), .Z(n4222));
Q_MX02 U4598 ( .S(oFill[1]), .A0(n4926), .A1(n4798), .Z(n4221));
Q_MX02 U4599 ( .S(oFill[1]), .A0(n4925), .A1(n4797), .Z(n4220));
Q_MX02 U4600 ( .S(oFill[1]), .A0(n4924), .A1(n4796), .Z(n4219));
Q_MX02 U4601 ( .S(oFill[1]), .A0(n4923), .A1(n4795), .Z(n4218));
Q_MX02 U4602 ( .S(oFill[1]), .A0(n4922), .A1(n4794), .Z(n4217));
Q_MX02 U4603 ( .S(oFill[1]), .A0(n4921), .A1(n4793), .Z(n4216));
Q_MX02 U4604 ( .S(oFill[1]), .A0(n4920), .A1(n4792), .Z(n4215));
Q_MX02 U4605 ( .S(oFill[1]), .A0(n4919), .A1(n4791), .Z(n4214));
Q_MX02 U4606 ( .S(oFill[1]), .A0(n4918), .A1(n4790), .Z(n4213));
Q_MX02 U4607 ( .S(oFill[1]), .A0(n4917), .A1(n4789), .Z(n4212));
Q_MX02 U4608 ( .S(oFill[1]), .A0(n4916), .A1(n4788), .Z(n4211));
Q_MX02 U4609 ( .S(oFill[1]), .A0(n4915), .A1(n4787), .Z(n4210));
Q_MX02 U4610 ( .S(oFill[1]), .A0(n4914), .A1(n4786), .Z(n4209));
Q_MX02 U4611 ( .S(oFill[1]), .A0(n4913), .A1(n4785), .Z(n4208));
Q_MX02 U4612 ( .S(oFill[1]), .A0(n4912), .A1(n4784), .Z(n4207));
Q_MX02 U4613 ( .S(oFill[1]), .A0(n4911), .A1(n4783), .Z(n4206));
Q_MX02 U4614 ( .S(oFill[1]), .A0(n4910), .A1(n4782), .Z(n4205));
Q_MX02 U4615 ( .S(oFill[1]), .A0(n4909), .A1(n4781), .Z(n4204));
Q_MX02 U4616 ( .S(oFill[1]), .A0(n4908), .A1(n4780), .Z(n4203));
Q_MX02 U4617 ( .S(oFill[1]), .A0(n4907), .A1(n4779), .Z(n4202));
Q_MX02 U4618 ( .S(oFill[1]), .A0(n4906), .A1(n4778), .Z(n4201));
Q_MX02 U4619 ( .S(oFill[1]), .A0(n4905), .A1(n4777), .Z(n4200));
Q_MX02 U4620 ( .S(oFill[1]), .A0(n4904), .A1(n4776), .Z(n4199));
Q_MX02 U4621 ( .S(oFill[1]), .A0(n4903), .A1(n4775), .Z(n4198));
Q_MX02 U4622 ( .S(oFill[1]), .A0(n4902), .A1(n4774), .Z(n4197));
Q_MX02 U4623 ( .S(oFill[1]), .A0(n4901), .A1(n4773), .Z(n4196));
Q_MX02 U4624 ( .S(oFill[1]), .A0(n4900), .A1(n4772), .Z(n4195));
Q_MX02 U4625 ( .S(oFill[1]), .A0(n4899), .A1(n4771), .Z(n4194));
Q_MX02 U4626 ( .S(oFill[1]), .A0(n4898), .A1(n4770), .Z(n4193));
Q_MX02 U4627 ( .S(oFill[1]), .A0(n4897), .A1(n4769), .Z(n4192));
Q_MX02 U4628 ( .S(oFill[1]), .A0(n4896), .A1(n4768), .Z(n4191));
Q_MX02 U4629 ( .S(oFill[1]), .A0(n4895), .A1(n4767), .Z(n4190));
Q_MX02 U4630 ( .S(oFill[1]), .A0(n4894), .A1(n4766), .Z(n4189));
Q_MX02 U4631 ( .S(oFill[1]), .A0(n4893), .A1(n4765), .Z(n4188));
Q_MX02 U4632 ( .S(oFill[1]), .A0(n4892), .A1(n4764), .Z(n4187));
Q_MX02 U4633 ( .S(oFill[1]), .A0(n4891), .A1(n4763), .Z(n4186));
Q_MX02 U4634 ( .S(oFill[1]), .A0(n4890), .A1(n4762), .Z(n4185));
Q_MX02 U4635 ( .S(oFill[1]), .A0(n4889), .A1(n4761), .Z(n4184));
Q_MX02 U4636 ( .S(oFill[1]), .A0(n4888), .A1(n4760), .Z(n4183));
Q_MX02 U4637 ( .S(oFill[1]), .A0(n4887), .A1(n4759), .Z(n4182));
Q_MX02 U4638 ( .S(oFill[1]), .A0(n4886), .A1(n4758), .Z(n4181));
Q_MX02 U4639 ( .S(oFill[1]), .A0(n4885), .A1(n4757), .Z(n4180));
Q_MX02 U4640 ( .S(oFill[1]), .A0(n4884), .A1(n4756), .Z(n4179));
Q_MX02 U4641 ( .S(oFill[1]), .A0(n4883), .A1(n4755), .Z(n4178));
Q_MX02 U4642 ( .S(oFill[1]), .A0(n4882), .A1(n4754), .Z(n4177));
Q_MX02 U4643 ( .S(oFill[1]), .A0(n4881), .A1(n4753), .Z(n4176));
Q_MX02 U4644 ( .S(oFill[1]), .A0(n4880), .A1(n4752), .Z(n4175));
Q_MX02 U4645 ( .S(oFill[1]), .A0(n4879), .A1(n4751), .Z(n4174));
Q_MX02 U4646 ( .S(oFill[1]), .A0(n4878), .A1(n4750), .Z(n4173));
Q_MX02 U4647 ( .S(oFill[1]), .A0(n4877), .A1(n4749), .Z(n4172));
Q_MX02 U4648 ( .S(oFill[1]), .A0(n4876), .A1(n4748), .Z(n4171));
Q_MX02 U4649 ( .S(oFill[1]), .A0(n4875), .A1(n4747), .Z(n4170));
Q_MX02 U4650 ( .S(oFill[1]), .A0(n4874), .A1(n4746), .Z(n4169));
Q_MX02 U4651 ( .S(oFill[1]), .A0(n4873), .A1(n4745), .Z(n4168));
Q_MX02 U4652 ( .S(oFill[1]), .A0(n4872), .A1(n4744), .Z(n4167));
Q_MX02 U4653 ( .S(oFill[1]), .A0(n4871), .A1(n4743), .Z(n4166));
Q_MX02 U4654 ( .S(oFill[1]), .A0(n4870), .A1(n4742), .Z(n4165));
Q_MX02 U4655 ( .S(oFill[1]), .A0(n4869), .A1(n4741), .Z(n4164));
Q_MX02 U4656 ( .S(oFill[1]), .A0(n4868), .A1(n4740), .Z(n4163));
Q_MX02 U4657 ( .S(oFill[1]), .A0(n4867), .A1(n4739), .Z(n4162));
Q_MX02 U4658 ( .S(oFill[1]), .A0(n4866), .A1(n4738), .Z(n4161));
Q_MX02 U4659 ( .S(oFill[1]), .A0(n4865), .A1(n4737), .Z(n4160));
Q_MX02 U4660 ( .S(oFill[1]), .A0(n4864), .A1(n4736), .Z(n4159));
Q_MX02 U4661 ( .S(oFill[1]), .A0(n4863), .A1(n4735), .Z(n4158));
Q_MX02 U4662 ( .S(oFill[1]), .A0(n4862), .A1(n4734), .Z(n4157));
Q_MX02 U4663 ( .S(oFill[1]), .A0(n4861), .A1(n4733), .Z(n4156));
Q_MX02 U4664 ( .S(oFill[1]), .A0(n4860), .A1(n4732), .Z(n4155));
Q_MX02 U4665 ( .S(oFill[1]), .A0(n4859), .A1(n4731), .Z(n4154));
Q_MX02 U4666 ( .S(oFill[1]), .A0(n4858), .A1(n4730), .Z(n4153));
Q_MX02 U4667 ( .S(oFill[1]), .A0(n4857), .A1(n4729), .Z(n4152));
Q_MX02 U4668 ( .S(oFill[1]), .A0(n4856), .A1(n4728), .Z(n4151));
Q_MX02 U4669 ( .S(oFill[1]), .A0(n4855), .A1(n4727), .Z(n4150));
Q_MX02 U4670 ( .S(oFill[1]), .A0(n4854), .A1(n4726), .Z(n4149));
Q_MX02 U4671 ( .S(oFill[1]), .A0(n4853), .A1(n4725), .Z(n4148));
Q_MX02 U4672 ( .S(oFill[1]), .A0(n4852), .A1(n4724), .Z(n4147));
Q_MX02 U4673 ( .S(oFill[1]), .A0(n4851), .A1(n4723), .Z(n4146));
Q_MX02 U4674 ( .S(oFill[1]), .A0(n4850), .A1(n4722), .Z(n4145));
Q_MX02 U4675 ( .S(oFill[1]), .A0(n4849), .A1(n4721), .Z(n4144));
Q_MX02 U4676 ( .S(oFill[1]), .A0(n4848), .A1(n4720), .Z(n4143));
Q_MX02 U4677 ( .S(oFill[1]), .A0(n4847), .A1(n4719), .Z(n4142));
Q_MX02 U4678 ( .S(oFill[1]), .A0(n4846), .A1(n4718), .Z(n4141));
Q_MX02 U4679 ( .S(oFill[1]), .A0(n4845), .A1(n4717), .Z(n4140));
Q_MX02 U4680 ( .S(oFill[1]), .A0(n4844), .A1(n4716), .Z(n4139));
Q_MX02 U4681 ( .S(oFill[1]), .A0(n4843), .A1(n4715), .Z(n4138));
Q_MX02 U4682 ( .S(oFill[1]), .A0(n4842), .A1(n4714), .Z(n4137));
Q_MX02 U4683 ( .S(oFill[1]), .A0(n4841), .A1(n4713), .Z(n4136));
Q_MX02 U4684 ( .S(oFill[1]), .A0(n4840), .A1(n4712), .Z(n4135));
Q_MX02 U4685 ( .S(oFill[1]), .A0(n4839), .A1(n4711), .Z(n4134));
Q_MX02 U4686 ( .S(oFill[1]), .A0(n4838), .A1(n4710), .Z(n4133));
Q_MX02 U4687 ( .S(oFill[1]), .A0(n4837), .A1(n4709), .Z(n4132));
Q_MX02 U4688 ( .S(oFill[1]), .A0(n4836), .A1(n4708), .Z(n4131));
Q_MX02 U4689 ( .S(oFill[1]), .A0(n4835), .A1(n4707), .Z(n4130));
Q_MX02 U4690 ( .S(oFill[1]), .A0(n4834), .A1(n4706), .Z(n4129));
Q_MX02 U4691 ( .S(oFill[1]), .A0(n4833), .A1(n4705), .Z(n4128));
Q_MX02 U4692 ( .S(oFill[1]), .A0(n4832), .A1(n4704), .Z(n4127));
Q_MX02 U4693 ( .S(oFill[1]), .A0(n4831), .A1(n4703), .Z(n4126));
Q_MX02 U4694 ( .S(oFill[1]), .A0(n4830), .A1(n4702), .Z(n4125));
Q_MX02 U4695 ( .S(oFill[1]), .A0(n4829), .A1(n4701), .Z(n4124));
Q_MX02 U4696 ( .S(oFill[1]), .A0(n4828), .A1(n4700), .Z(n4123));
Q_MX02 U4697 ( .S(oFill[1]), .A0(n4827), .A1(n4699), .Z(n4122));
Q_MX02 U4698 ( .S(oFill[1]), .A0(n4826), .A1(n4698), .Z(n4121));
Q_MX02 U4699 ( .S(oFill[1]), .A0(n4825), .A1(n4697), .Z(n4120));
Q_MX02 U4700 ( .S(oFill[1]), .A0(n4824), .A1(n4696), .Z(n4119));
Q_MX02 U4701 ( .S(oFill[1]), .A0(n4823), .A1(n4695), .Z(n4118));
Q_MX02 U4702 ( .S(oFill[1]), .A0(n4822), .A1(n4694), .Z(n4117));
Q_MX02 U4703 ( .S(oFill[1]), .A0(n4821), .A1(n4693), .Z(n4116));
Q_MX02 U4704 ( .S(oFill[1]), .A0(n4820), .A1(n4692), .Z(n4115));
Q_MX02 U4705 ( .S(oFill[1]), .A0(n4819), .A1(n4691), .Z(n4114));
Q_MX02 U4706 ( .S(oFill[1]), .A0(n4818), .A1(n4690), .Z(n4113));
Q_MX02 U4707 ( .S(oFill[1]), .A0(n4817), .A1(n4689), .Z(n4112));
Q_MX02 U4708 ( .S(oFill[1]), .A0(n4816), .A1(n4688), .Z(n4111));
Q_MX02 U4709 ( .S(oFill[1]), .A0(n4815), .A1(n4687), .Z(n4110));
Q_MX02 U4710 ( .S(oFill[1]), .A0(n4814), .A1(n4686), .Z(n4109));
Q_MX02 U4711 ( .S(oFill[1]), .A0(n4813), .A1(n4685), .Z(n4108));
Q_MX02 U4712 ( .S(oFill[1]), .A0(n4812), .A1(n4684), .Z(n4107));
Q_MX02 U4713 ( .S(oFill[1]), .A0(n4811), .A1(n4683), .Z(n4106));
Q_MX02 U4714 ( .S(oFill[1]), .A0(n4810), .A1(n4682), .Z(n4105));
Q_MX02 U4715 ( .S(oFill[1]), .A0(n4809), .A1(n4681), .Z(n4104));
Q_MX02 U4716 ( .S(oFill[1]), .A0(n4808), .A1(n4680), .Z(n4103));
Q_MX02 U4717 ( .S(oFill[1]), .A0(n4807), .A1(n4679), .Z(n4102));
Q_MX02 U4718 ( .S(oFill[1]), .A0(n4806), .A1(n4678), .Z(n4101));
Q_MX02 U4719 ( .S(oFill[1]), .A0(n4805), .A1(n4677), .Z(n4100));
Q_MX02 U4720 ( .S(oFill[1]), .A0(n4804), .A1(n4676), .Z(n4099));
Q_MX02 U4721 ( .S(oFill[1]), .A0(n4803), .A1(n4675), .Z(n4098));
Q_MX02 U4722 ( .S(oFill[1]), .A0(n4802), .A1(n4674), .Z(n4097));
Q_MX02 U4723 ( .S(oFill[1]), .A0(n4801), .A1(n4673), .Z(n4096));
Q_MX02 U4724 ( .S(oFill[1]), .A0(n4800), .A1(n4672), .Z(n4095));
Q_MX02 U4725 ( .S(oFill[1]), .A0(n4799), .A1(n4671), .Z(n4094));
Q_MX02 U4726 ( .S(oFill[1]), .A0(n4798), .A1(n4670), .Z(n4093));
Q_MX02 U4727 ( .S(oFill[1]), .A0(n4797), .A1(n4669), .Z(n4092));
Q_MX02 U4728 ( .S(oFill[1]), .A0(n4796), .A1(n4668), .Z(n4091));
Q_MX02 U4729 ( .S(oFill[1]), .A0(n4795), .A1(n4667), .Z(n4090));
Q_MX02 U4730 ( .S(oFill[1]), .A0(n4794), .A1(n4666), .Z(n4089));
Q_MX02 U4731 ( .S(oFill[1]), .A0(n4793), .A1(n4665), .Z(n4088));
Q_MX02 U4732 ( .S(oFill[1]), .A0(n4792), .A1(n4664), .Z(n4087));
Q_MX02 U4733 ( .S(oFill[1]), .A0(n4791), .A1(n4663), .Z(n4086));
Q_MX02 U4734 ( .S(oFill[1]), .A0(n4790), .A1(n4662), .Z(n4085));
Q_MX02 U4735 ( .S(oFill[1]), .A0(n4789), .A1(n4661), .Z(n4084));
Q_MX02 U4736 ( .S(oFill[1]), .A0(n4788), .A1(n4660), .Z(n4083));
Q_MX02 U4737 ( .S(oFill[1]), .A0(n4787), .A1(n4659), .Z(n4082));
Q_MX02 U4738 ( .S(oFill[1]), .A0(n4786), .A1(n4658), .Z(n4081));
Q_MX02 U4739 ( .S(oFill[1]), .A0(n4785), .A1(n4657), .Z(n4080));
Q_MX02 U4740 ( .S(oFill[1]), .A0(n4784), .A1(n4656), .Z(n4079));
Q_MX02 U4741 ( .S(oFill[1]), .A0(n4783), .A1(n4655), .Z(n4078));
Q_MX02 U4742 ( .S(oFill[1]), .A0(n4782), .A1(n4654), .Z(n4077));
Q_MX02 U4743 ( .S(oFill[1]), .A0(n4781), .A1(n4653), .Z(n4076));
Q_MX02 U4744 ( .S(oFill[1]), .A0(n4780), .A1(n4652), .Z(n4075));
Q_MX02 U4745 ( .S(oFill[1]), .A0(n4779), .A1(n4651), .Z(n4074));
Q_MX02 U4746 ( .S(oFill[1]), .A0(n4778), .A1(n4650), .Z(n4073));
Q_MX02 U4747 ( .S(oFill[1]), .A0(n4777), .A1(n4649), .Z(n4072));
Q_MX02 U4748 ( .S(oFill[1]), .A0(n4776), .A1(n4648), .Z(n4071));
Q_MX02 U4749 ( .S(oFill[1]), .A0(n4775), .A1(n4647), .Z(n4070));
Q_MX02 U4750 ( .S(oFill[1]), .A0(n4774), .A1(n4646), .Z(n4069));
Q_MX02 U4751 ( .S(oFill[1]), .A0(n4773), .A1(n4645), .Z(n4068));
Q_MX02 U4752 ( .S(oFill[1]), .A0(n4772), .A1(n4644), .Z(n4067));
Q_MX02 U4753 ( .S(oFill[1]), .A0(n4771), .A1(n4643), .Z(n4066));
Q_MX02 U4754 ( .S(oFill[1]), .A0(n4770), .A1(n4642), .Z(n4065));
Q_MX02 U4755 ( .S(oFill[1]), .A0(n4769), .A1(n4641), .Z(n4064));
Q_MX02 U4756 ( .S(oFill[1]), .A0(n4768), .A1(n4640), .Z(n4063));
Q_MX02 U4757 ( .S(oFill[1]), .A0(n4767), .A1(n4639), .Z(n4062));
Q_MX02 U4758 ( .S(oFill[1]), .A0(n4766), .A1(n4638), .Z(n4061));
Q_MX02 U4759 ( .S(oFill[1]), .A0(n4765), .A1(n4637), .Z(n4060));
Q_MX02 U4760 ( .S(oFill[1]), .A0(n4764), .A1(n4636), .Z(n4059));
Q_MX02 U4761 ( .S(oFill[1]), .A0(n4763), .A1(n4635), .Z(n4058));
Q_MX02 U4762 ( .S(oFill[1]), .A0(n4762), .A1(n4634), .Z(n4057));
Q_MX02 U4763 ( .S(oFill[1]), .A0(n4761), .A1(n4633), .Z(n4056));
Q_MX02 U4764 ( .S(oFill[1]), .A0(n4760), .A1(n4632), .Z(n4055));
Q_MX02 U4765 ( .S(oFill[1]), .A0(n4759), .A1(n4631), .Z(n4054));
Q_MX02 U4766 ( .S(oFill[1]), .A0(n4758), .A1(n4630), .Z(n4053));
Q_MX02 U4767 ( .S(oFill[1]), .A0(n4757), .A1(n4629), .Z(n4052));
Q_MX02 U4768 ( .S(oFill[1]), .A0(n4756), .A1(n4628), .Z(n4051));
Q_MX02 U4769 ( .S(oFill[1]), .A0(n4755), .A1(n4627), .Z(n4050));
Q_MX02 U4770 ( .S(oFill[1]), .A0(n4754), .A1(n4626), .Z(n4049));
Q_MX02 U4771 ( .S(oFill[1]), .A0(n4753), .A1(n4625), .Z(n4048));
Q_MX02 U4772 ( .S(oFill[1]), .A0(n4752), .A1(n4624), .Z(n4047));
Q_MX02 U4773 ( .S(oFill[1]), .A0(n4751), .A1(n4623), .Z(n4046));
Q_MX02 U4774 ( .S(oFill[1]), .A0(n4750), .A1(n4622), .Z(n4045));
Q_MX02 U4775 ( .S(oFill[1]), .A0(n4749), .A1(n4621), .Z(n4044));
Q_MX02 U4776 ( .S(oFill[1]), .A0(n4748), .A1(n4620), .Z(n4043));
Q_MX02 U4777 ( .S(oFill[1]), .A0(n4747), .A1(n4619), .Z(n4042));
Q_MX02 U4778 ( .S(oFill[1]), .A0(n4746), .A1(n4618), .Z(n4041));
Q_MX02 U4779 ( .S(oFill[1]), .A0(n4745), .A1(n4617), .Z(n4040));
Q_MX02 U4780 ( .S(oFill[1]), .A0(n4744), .A1(n4616), .Z(n4039));
Q_MX02 U4781 ( .S(oFill[1]), .A0(n4743), .A1(n4615), .Z(n4038));
Q_MX02 U4782 ( .S(oFill[1]), .A0(n4742), .A1(n4614), .Z(n4037));
Q_MX02 U4783 ( .S(oFill[1]), .A0(n4741), .A1(n4613), .Z(n4036));
Q_MX02 U4784 ( .S(oFill[1]), .A0(n4740), .A1(n4612), .Z(n4035));
Q_MX02 U4785 ( .S(oFill[1]), .A0(n4739), .A1(n4611), .Z(n4034));
Q_MX02 U4786 ( .S(oFill[1]), .A0(n4738), .A1(n4610), .Z(n4033));
Q_MX02 U4787 ( .S(oFill[1]), .A0(n4737), .A1(n4609), .Z(n4032));
Q_MX02 U4788 ( .S(oFill[1]), .A0(n4736), .A1(n4608), .Z(n4031));
Q_MX02 U4789 ( .S(oFill[1]), .A0(n4735), .A1(n4607), .Z(n4030));
Q_MX02 U4790 ( .S(oFill[1]), .A0(n4734), .A1(n4606), .Z(n4029));
Q_MX02 U4791 ( .S(oFill[1]), .A0(n4733), .A1(n4605), .Z(n4028));
Q_MX02 U4792 ( .S(oFill[1]), .A0(n4732), .A1(n4604), .Z(n4027));
Q_MX02 U4793 ( .S(oFill[1]), .A0(n4731), .A1(n4603), .Z(n4026));
Q_MX02 U4794 ( .S(oFill[1]), .A0(n4730), .A1(n4602), .Z(n4025));
Q_MX02 U4795 ( .S(oFill[1]), .A0(n4729), .A1(n4601), .Z(n4024));
Q_MX02 U4796 ( .S(oFill[1]), .A0(n4728), .A1(n4600), .Z(n4023));
Q_MX02 U4797 ( .S(oFill[1]), .A0(n4727), .A1(n4599), .Z(n4022));
Q_MX02 U4798 ( .S(oFill[1]), .A0(n4726), .A1(n4598), .Z(n4021));
Q_MX02 U4799 ( .S(oFill[1]), .A0(n4725), .A1(n4597), .Z(n4020));
Q_MX02 U4800 ( .S(oFill[1]), .A0(n4724), .A1(n4596), .Z(n4019));
Q_MX02 U4801 ( .S(oFill[1]), .A0(n4723), .A1(n4595), .Z(n4018));
Q_MX02 U4802 ( .S(oFill[1]), .A0(n4722), .A1(n4594), .Z(n4017));
Q_MX02 U4803 ( .S(oFill[1]), .A0(n4721), .A1(n4593), .Z(n4016));
Q_MX02 U4804 ( .S(oFill[1]), .A0(n4720), .A1(n4592), .Z(n4015));
Q_MX02 U4805 ( .S(oFill[1]), .A0(n4719), .A1(n4591), .Z(n4014));
Q_MX02 U4806 ( .S(oFill[1]), .A0(n4718), .A1(n4590), .Z(n4013));
Q_MX02 U4807 ( .S(oFill[1]), .A0(n4717), .A1(n4589), .Z(n4012));
Q_MX02 U4808 ( .S(oFill[1]), .A0(n4716), .A1(n4588), .Z(n4011));
Q_MX02 U4809 ( .S(oFill[1]), .A0(n4715), .A1(n4587), .Z(n4010));
Q_MX02 U4810 ( .S(oFill[1]), .A0(n4714), .A1(n4586), .Z(n4009));
Q_MX02 U4811 ( .S(oFill[1]), .A0(n4713), .A1(n4585), .Z(n4008));
Q_MX02 U4812 ( .S(oFill[1]), .A0(n4712), .A1(n4584), .Z(n4007));
Q_MX02 U4813 ( .S(oFill[1]), .A0(n4711), .A1(n4583), .Z(n4006));
Q_MX02 U4814 ( .S(oFill[1]), .A0(n4710), .A1(n4582), .Z(n4005));
Q_MX02 U4815 ( .S(oFill[1]), .A0(n4709), .A1(n4581), .Z(n4004));
Q_MX02 U4816 ( .S(oFill[1]), .A0(n4708), .A1(n4580), .Z(n4003));
Q_MX02 U4817 ( .S(oFill[1]), .A0(n4707), .A1(n4579), .Z(n4002));
Q_MX02 U4818 ( .S(oFill[1]), .A0(n4706), .A1(n4578), .Z(n4001));
Q_MX02 U4819 ( .S(oFill[1]), .A0(n4705), .A1(n4577), .Z(n4000));
Q_MX02 U4820 ( .S(oFill[1]), .A0(n4704), .A1(n4576), .Z(n3999));
Q_MX02 U4821 ( .S(oFill[1]), .A0(n4703), .A1(n4575), .Z(n3998));
Q_MX02 U4822 ( .S(oFill[1]), .A0(n4702), .A1(n4574), .Z(n3997));
Q_MX02 U4823 ( .S(oFill[1]), .A0(n4701), .A1(n4573), .Z(n3996));
Q_MX02 U4824 ( .S(oFill[1]), .A0(n4700), .A1(n4572), .Z(n3995));
Q_MX02 U4825 ( .S(oFill[1]), .A0(n4699), .A1(n4571), .Z(n3994));
Q_MX02 U4826 ( .S(oFill[1]), .A0(n4698), .A1(n4570), .Z(n3993));
Q_MX02 U4827 ( .S(oFill[1]), .A0(n4697), .A1(n4569), .Z(n3992));
Q_MX02 U4828 ( .S(oFill[1]), .A0(n4696), .A1(n4568), .Z(n3991));
Q_MX02 U4829 ( .S(oFill[1]), .A0(n4695), .A1(n4567), .Z(n3990));
Q_MX02 U4830 ( .S(oFill[1]), .A0(n4694), .A1(n4566), .Z(n3989));
Q_MX02 U4831 ( .S(oFill[1]), .A0(n4693), .A1(n4565), .Z(n3988));
Q_MX02 U4832 ( .S(oFill[1]), .A0(n4692), .A1(n4564), .Z(n3987));
Q_MX02 U4833 ( .S(oFill[1]), .A0(n4691), .A1(n4563), .Z(n3986));
Q_MX02 U4834 ( .S(oFill[1]), .A0(n4690), .A1(n4562), .Z(n3985));
Q_MX02 U4835 ( .S(oFill[1]), .A0(n4689), .A1(n4561), .Z(n3984));
Q_MX02 U4836 ( .S(oFill[1]), .A0(n4688), .A1(n4560), .Z(n3983));
Q_MX02 U4837 ( .S(oFill[1]), .A0(n4687), .A1(n4559), .Z(n3982));
Q_MX02 U4838 ( .S(oFill[1]), .A0(n4686), .A1(n4558), .Z(n3981));
Q_MX02 U4839 ( .S(oFill[1]), .A0(n4685), .A1(n4557), .Z(n3980));
Q_MX02 U4840 ( .S(oFill[1]), .A0(n4684), .A1(n4556), .Z(n3979));
Q_MX02 U4841 ( .S(oFill[1]), .A0(n4683), .A1(n4555), .Z(n3978));
Q_MX02 U4842 ( .S(oFill[1]), .A0(n4682), .A1(n4554), .Z(n3977));
Q_MX02 U4843 ( .S(oFill[1]), .A0(n4681), .A1(n4553), .Z(n3976));
Q_MX02 U4844 ( .S(oFill[1]), .A0(n4680), .A1(n4552), .Z(n3975));
Q_MX02 U4845 ( .S(oFill[1]), .A0(n4679), .A1(n4551), .Z(n3974));
Q_MX02 U4846 ( .S(oFill[1]), .A0(n4678), .A1(n4550), .Z(n3973));
Q_MX02 U4847 ( .S(oFill[1]), .A0(n4677), .A1(n4549), .Z(n3972));
Q_MX02 U4848 ( .S(oFill[1]), .A0(n4676), .A1(n4548), .Z(n3971));
Q_MX02 U4849 ( .S(oFill[1]), .A0(n4675), .A1(n4547), .Z(n3970));
Q_MX02 U4850 ( .S(oFill[1]), .A0(n4674), .A1(n4546), .Z(n3969));
Q_MX02 U4851 ( .S(oFill[1]), .A0(n4673), .A1(n4545), .Z(n3968));
Q_MX02 U4852 ( .S(oFill[1]), .A0(n4672), .A1(n4544), .Z(n3967));
Q_MX02 U4853 ( .S(oFill[1]), .A0(n4671), .A1(n4543), .Z(n3966));
Q_MX02 U4854 ( .S(oFill[1]), .A0(n4670), .A1(n4542), .Z(n3965));
Q_MX02 U4855 ( .S(oFill[1]), .A0(n4669), .A1(n4541), .Z(n3964));
Q_MX02 U4856 ( .S(oFill[1]), .A0(n4668), .A1(n4540), .Z(n3963));
Q_MX02 U4857 ( .S(oFill[1]), .A0(n4667), .A1(n4539), .Z(n3962));
Q_MX02 U4858 ( .S(oFill[1]), .A0(n4666), .A1(n4538), .Z(n3961));
Q_MX02 U4859 ( .S(oFill[1]), .A0(n4665), .A1(n4537), .Z(n3960));
Q_MX02 U4860 ( .S(oFill[1]), .A0(n4664), .A1(n4536), .Z(n3959));
Q_MX02 U4861 ( .S(oFill[1]), .A0(n4663), .A1(n4535), .Z(n3958));
Q_MX02 U4862 ( .S(oFill[1]), .A0(n4662), .A1(n4534), .Z(n3957));
Q_MX02 U4863 ( .S(oFill[1]), .A0(n4661), .A1(n4533), .Z(n3956));
Q_MX02 U4864 ( .S(oFill[1]), .A0(n4660), .A1(n4532), .Z(n3955));
Q_MX02 U4865 ( .S(oFill[1]), .A0(n4659), .A1(n4531), .Z(n3954));
Q_MX02 U4866 ( .S(oFill[1]), .A0(n4658), .A1(n4530), .Z(n3953));
Q_MX02 U4867 ( .S(oFill[1]), .A0(n4657), .A1(n4529), .Z(n3952));
Q_MX02 U4868 ( .S(oFill[1]), .A0(n4656), .A1(n4528), .Z(n3951));
Q_MX02 U4869 ( .S(oFill[1]), .A0(n4655), .A1(n4527), .Z(n3950));
Q_MX02 U4870 ( .S(oFill[1]), .A0(n4654), .A1(n4526), .Z(n3949));
Q_MX02 U4871 ( .S(oFill[1]), .A0(n4653), .A1(n4525), .Z(n3948));
Q_MX02 U4872 ( .S(oFill[1]), .A0(n4652), .A1(n4524), .Z(n3947));
Q_MX02 U4873 ( .S(oFill[1]), .A0(n4651), .A1(n4523), .Z(n3946));
Q_MX02 U4874 ( .S(oFill[1]), .A0(n4650), .A1(n4522), .Z(n3945));
Q_MX02 U4875 ( .S(oFill[1]), .A0(n4649), .A1(n4521), .Z(n3944));
Q_MX02 U4876 ( .S(oFill[1]), .A0(n4648), .A1(n4520), .Z(n3943));
Q_MX02 U4877 ( .S(oFill[1]), .A0(n4647), .A1(n4519), .Z(n3942));
Q_MX02 U4878 ( .S(oFill[1]), .A0(n4646), .A1(n4518), .Z(n3941));
Q_MX02 U4879 ( .S(oFill[1]), .A0(n4645), .A1(n4517), .Z(n3940));
Q_MX02 U4880 ( .S(oFill[1]), .A0(n4644), .A1(n4516), .Z(n3939));
Q_MX02 U4881 ( .S(oFill[1]), .A0(n4643), .A1(n4515), .Z(n3938));
Q_MX02 U4882 ( .S(oFill[1]), .A0(n4642), .A1(n4514), .Z(n3937));
Q_MX02 U4883 ( .S(oFill[1]), .A0(n4641), .A1(n4513), .Z(n3936));
Q_MX02 U4884 ( .S(oFill[1]), .A0(n4640), .A1(n4512), .Z(n3935));
Q_MX02 U4885 ( .S(oFill[1]), .A0(n4639), .A1(n4511), .Z(n3934));
Q_MX02 U4886 ( .S(oFill[1]), .A0(n4638), .A1(n4510), .Z(n3933));
Q_MX02 U4887 ( .S(oFill[1]), .A0(n4637), .A1(n4509), .Z(n3932));
Q_MX02 U4888 ( .S(oFill[1]), .A0(n4636), .A1(n4508), .Z(n3931));
Q_MX02 U4889 ( .S(oFill[1]), .A0(n4635), .A1(n4507), .Z(n3930));
Q_MX02 U4890 ( .S(oFill[1]), .A0(n4634), .A1(n4506), .Z(n3929));
Q_MX02 U4891 ( .S(oFill[1]), .A0(n4633), .A1(n4505), .Z(n3928));
Q_MX02 U4892 ( .S(oFill[1]), .A0(n4632), .A1(n4504), .Z(n3927));
Q_MX02 U4893 ( .S(oFill[1]), .A0(n4631), .A1(n4503), .Z(n3926));
Q_MX02 U4894 ( .S(oFill[1]), .A0(n4630), .A1(n4502), .Z(n3925));
Q_MX02 U4895 ( .S(oFill[1]), .A0(n4629), .A1(n4501), .Z(n3924));
Q_MX02 U4896 ( .S(oFill[1]), .A0(n4628), .A1(n4500), .Z(n3923));
Q_MX02 U4897 ( .S(oFill[1]), .A0(n4627), .A1(n4498), .Z(n3922));
Q_MX02 U4898 ( .S(oFill[1]), .A0(n4626), .A1(n4497), .Z(n3921));
Q_MX02 U4899 ( .S(oFill[1]), .A0(n4625), .A1(n4496), .Z(n3920));
Q_MX02 U4900 ( .S(oFill[1]), .A0(n4624), .A1(n4495), .Z(n3919));
Q_MX02 U4901 ( .S(oFill[1]), .A0(n4623), .A1(n4494), .Z(n3918));
Q_MX02 U4902 ( .S(oFill[1]), .A0(n4622), .A1(n4493), .Z(n3917));
Q_MX02 U4903 ( .S(oFill[1]), .A0(n4621), .A1(n4492), .Z(n3916));
Q_MX02 U4904 ( .S(oFill[1]), .A0(n4620), .A1(n4491), .Z(n3915));
Q_MX02 U4905 ( .S(oFill[1]), .A0(n4619), .A1(n4490), .Z(n3914));
Q_MX02 U4906 ( .S(oFill[1]), .A0(n4618), .A1(n4489), .Z(n3913));
Q_MX02 U4907 ( .S(oFill[1]), .A0(n4617), .A1(n4488), .Z(n3912));
Q_MX02 U4908 ( .S(oFill[1]), .A0(n4616), .A1(n4487), .Z(n3911));
Q_MX02 U4909 ( .S(oFill[1]), .A0(n4615), .A1(n4486), .Z(n3910));
Q_MX02 U4910 ( .S(oFill[1]), .A0(n4614), .A1(n4485), .Z(n3909));
Q_MX02 U4911 ( .S(oFill[1]), .A0(n4613), .A1(n4484), .Z(n3908));
Q_MX02 U4912 ( .S(oFill[1]), .A0(n4612), .A1(n4483), .Z(n3907));
Q_MX02 U4913 ( .S(oFill[1]), .A0(n4611), .A1(n4482), .Z(n3906));
Q_MX02 U4914 ( .S(oFill[1]), .A0(n4610), .A1(n4481), .Z(n3905));
Q_MX02 U4915 ( .S(oFill[1]), .A0(n4609), .A1(n4480), .Z(n3904));
Q_MX02 U4916 ( .S(oFill[1]), .A0(n4608), .A1(n4479), .Z(n3903));
Q_MX02 U4917 ( .S(oFill[1]), .A0(n4607), .A1(n4478), .Z(n3902));
Q_MX02 U4918 ( .S(oFill[1]), .A0(n4606), .A1(n4477), .Z(n3901));
Q_MX02 U4919 ( .S(oFill[1]), .A0(n4605), .A1(n4476), .Z(n3900));
Q_MX02 U4920 ( .S(oFill[1]), .A0(n4604), .A1(n4475), .Z(n3899));
Q_MX02 U4921 ( .S(oFill[1]), .A0(n4603), .A1(n4474), .Z(n3898));
Q_MX02 U4922 ( .S(oFill[1]), .A0(n4602), .A1(n4473), .Z(n3897));
Q_MX02 U4923 ( .S(oFill[1]), .A0(n4601), .A1(n4472), .Z(n3896));
Q_MX02 U4924 ( .S(oFill[1]), .A0(n4600), .A1(n4471), .Z(n3895));
Q_MX02 U4925 ( .S(oFill[1]), .A0(n4599), .A1(n4470), .Z(n3894));
Q_MX02 U4926 ( .S(oFill[1]), .A0(n4598), .A1(n4469), .Z(n3893));
Q_MX02 U4927 ( .S(oFill[1]), .A0(n4597), .A1(n4468), .Z(n3892));
Q_MX02 U4928 ( .S(oFill[1]), .A0(n4596), .A1(n4467), .Z(n3891));
Q_MX02 U4929 ( .S(oFill[1]), .A0(n4595), .A1(n4466), .Z(n3890));
Q_MX02 U4930 ( .S(oFill[1]), .A0(n4594), .A1(n4465), .Z(n3889));
Q_MX02 U4931 ( .S(oFill[1]), .A0(n4593), .A1(n4464), .Z(n3888));
Q_MX02 U4932 ( .S(oFill[1]), .A0(n4592), .A1(n4463), .Z(n3887));
Q_MX02 U4933 ( .S(oFill[1]), .A0(n4591), .A1(n4462), .Z(n3886));
Q_MX02 U4934 ( .S(oFill[1]), .A0(n4590), .A1(n4461), .Z(n3885));
Q_MX02 U4935 ( .S(oFill[1]), .A0(n4589), .A1(n4460), .Z(n3884));
Q_MX02 U4936 ( .S(oFill[1]), .A0(n4588), .A1(n4459), .Z(n3883));
Q_MX02 U4937 ( .S(oFill[1]), .A0(n4587), .A1(n4458), .Z(n3882));
Q_MX02 U4938 ( .S(oFill[1]), .A0(n4586), .A1(n4457), .Z(n3881));
Q_MX02 U4939 ( .S(oFill[1]), .A0(n4585), .A1(n4456), .Z(n3880));
Q_MX02 U4940 ( .S(oFill[1]), .A0(n4584), .A1(n4455), .Z(n3879));
Q_MX02 U4941 ( .S(oFill[1]), .A0(n4583), .A1(n4454), .Z(n3878));
Q_MX02 U4942 ( .S(oFill[1]), .A0(n4582), .A1(n4453), .Z(n3877));
Q_MX02 U4943 ( .S(oFill[1]), .A0(n4581), .A1(n4452), .Z(n3876));
Q_MX02 U4944 ( .S(oFill[1]), .A0(n4580), .A1(n4451), .Z(n3875));
Q_MX02 U4945 ( .S(oFill[1]), .A0(n4579), .A1(n4450), .Z(n3874));
Q_MX02 U4946 ( .S(oFill[1]), .A0(n4578), .A1(n4449), .Z(n3873));
Q_MX02 U4947 ( .S(oFill[1]), .A0(n4577), .A1(n4448), .Z(n3872));
Q_MX02 U4948 ( .S(oFill[1]), .A0(n4576), .A1(n4447), .Z(n3871));
Q_MX02 U4949 ( .S(oFill[1]), .A0(n4575), .A1(n4446), .Z(n3870));
Q_MX02 U4950 ( .S(oFill[1]), .A0(n4574), .A1(n4445), .Z(n3869));
Q_MX02 U4951 ( .S(oFill[1]), .A0(n4573), .A1(n4444), .Z(n3868));
Q_MX02 U4952 ( .S(oFill[1]), .A0(n4572), .A1(n4443), .Z(n3867));
Q_MX02 U4953 ( .S(oFill[1]), .A0(n4571), .A1(n4442), .Z(n3866));
Q_MX02 U4954 ( .S(oFill[1]), .A0(n4570), .A1(n4441), .Z(n3865));
Q_MX02 U4955 ( .S(oFill[1]), .A0(n4569), .A1(n4440), .Z(n3864));
Q_MX02 U4956 ( .S(oFill[1]), .A0(n4568), .A1(n4439), .Z(n3863));
Q_MX02 U4957 ( .S(oFill[1]), .A0(n4567), .A1(n4438), .Z(n3862));
Q_MX02 U4958 ( .S(oFill[1]), .A0(n4566), .A1(n4437), .Z(n3861));
Q_MX02 U4959 ( .S(oFill[1]), .A0(n4565), .A1(n4436), .Z(n3860));
Q_MX02 U4960 ( .S(oFill[1]), .A0(n4564), .A1(n4435), .Z(n3859));
Q_INV U4961 ( .A(oFill[1]), .Z(n3858));
Q_AN02 U4962 ( .A0(n3858), .A1(n4563), .Z(n3857));
Q_AN02 U4963 ( .A0(n3858), .A1(n4562), .Z(n3856));
Q_AN02 U4964 ( .A0(n3858), .A1(n4561), .Z(n3855));
Q_AN02 U4965 ( .A0(n3858), .A1(n4560), .Z(n3854));
Q_AN02 U4966 ( .A0(n3858), .A1(n4559), .Z(n3853));
Q_AN02 U4967 ( .A0(n3858), .A1(n4558), .Z(n3852));
Q_AN02 U4968 ( .A0(n3858), .A1(n4557), .Z(n3851));
Q_AN02 U4969 ( .A0(n3858), .A1(n4556), .Z(n3850));
Q_AN02 U4970 ( .A0(n3858), .A1(n4555), .Z(n3849));
Q_AN02 U4971 ( .A0(n3858), .A1(n4554), .Z(n3848));
Q_AN02 U4972 ( .A0(n3858), .A1(n4553), .Z(n3847));
Q_AN02 U4973 ( .A0(n3858), .A1(n4552), .Z(n3846));
Q_AN02 U4974 ( .A0(n3858), .A1(n4551), .Z(n3845));
Q_AN02 U4975 ( .A0(n3858), .A1(n4550), .Z(n3844));
Q_AN02 U4976 ( .A0(n3858), .A1(n4549), .Z(n3843));
Q_AN02 U4977 ( .A0(n3858), .A1(n4548), .Z(n3842));
Q_AN02 U4978 ( .A0(n3858), .A1(n4547), .Z(n3841));
Q_AN02 U4979 ( .A0(n3858), .A1(n4546), .Z(n3840));
Q_AN02 U4980 ( .A0(n3858), .A1(n4545), .Z(n3839));
Q_AN02 U4981 ( .A0(n3858), .A1(n4544), .Z(n3838));
Q_AN02 U4982 ( .A0(n3858), .A1(n4543), .Z(n3837));
Q_AN02 U4983 ( .A0(n3858), .A1(n4542), .Z(n3836));
Q_AN02 U4984 ( .A0(n3858), .A1(n4541), .Z(n3835));
Q_AN02 U4985 ( .A0(n3858), .A1(n4540), .Z(n3834));
Q_AN02 U4986 ( .A0(n3858), .A1(n4539), .Z(n3833));
Q_AN02 U4987 ( .A0(n3858), .A1(n4538), .Z(n3832));
Q_AN02 U4988 ( .A0(n3858), .A1(n4537), .Z(n3831));
Q_AN02 U4989 ( .A0(n3858), .A1(n4536), .Z(n3830));
Q_AN02 U4990 ( .A0(n3858), .A1(n4535), .Z(n3829));
Q_AN02 U4991 ( .A0(n3858), .A1(n4534), .Z(n3828));
Q_AN02 U4992 ( .A0(n3858), .A1(n4533), .Z(n3827));
Q_AN02 U4993 ( .A0(n3858), .A1(n4532), .Z(n3826));
Q_AN02 U4994 ( .A0(n3858), .A1(n4531), .Z(n3825));
Q_AN02 U4995 ( .A0(n3858), .A1(n4530), .Z(n3824));
Q_AN02 U4996 ( .A0(n3858), .A1(n4529), .Z(n3823));
Q_AN02 U4997 ( .A0(n3858), .A1(n4528), .Z(n3822));
Q_AN02 U4998 ( .A0(n3858), .A1(n4527), .Z(n3821));
Q_AN02 U4999 ( .A0(n3858), .A1(n4526), .Z(n3820));
Q_AN02 U5000 ( .A0(n3858), .A1(n4525), .Z(n3819));
Q_AN02 U5001 ( .A0(n3858), .A1(n4524), .Z(n3818));
Q_AN02 U5002 ( .A0(n3858), .A1(n4523), .Z(n3817));
Q_AN02 U5003 ( .A0(n3858), .A1(n4522), .Z(n3816));
Q_AN02 U5004 ( .A0(n3858), .A1(n4521), .Z(n3815));
Q_AN02 U5005 ( .A0(n3858), .A1(n4520), .Z(n3814));
Q_AN02 U5006 ( .A0(n3858), .A1(n4519), .Z(n3813));
Q_AN02 U5007 ( .A0(n3858), .A1(n4518), .Z(n3812));
Q_AN02 U5008 ( .A0(n3858), .A1(n4517), .Z(n3811));
Q_AN02 U5009 ( .A0(n3858), .A1(n4516), .Z(n3810));
Q_AN02 U5010 ( .A0(n3858), .A1(n4515), .Z(n3809));
Q_AN02 U5011 ( .A0(n3858), .A1(n4514), .Z(n3808));
Q_AN02 U5012 ( .A0(n3858), .A1(n4513), .Z(n3807));
Q_AN02 U5013 ( .A0(n3858), .A1(n4512), .Z(n3806));
Q_AN02 U5014 ( .A0(n3858), .A1(n4511), .Z(n3805));
Q_AN02 U5015 ( .A0(n3858), .A1(n4510), .Z(n3804));
Q_AN02 U5016 ( .A0(n3858), .A1(n4509), .Z(n3803));
Q_AN02 U5017 ( .A0(n3858), .A1(n4508), .Z(n3802));
Q_AN02 U5018 ( .A0(n3858), .A1(n4507), .Z(n3801));
Q_AN02 U5019 ( .A0(n3858), .A1(n4506), .Z(n3800));
Q_AN02 U5020 ( .A0(n3858), .A1(n4505), .Z(n3799));
Q_AN02 U5021 ( .A0(n3858), .A1(n4504), .Z(n3798));
Q_AN02 U5022 ( .A0(n3858), .A1(n4503), .Z(n3797));
Q_AN02 U5023 ( .A0(n3858), .A1(n4502), .Z(n3796));
Q_AN02 U5024 ( .A0(n3858), .A1(n4501), .Z(n3795));
Q_AN02 U5025 ( .A0(n3858), .A1(n4500), .Z(n3794));
Q_AN02 U5026 ( .A0(n3858), .A1(n4498), .Z(n3793));
Q_AN02 U5027 ( .A0(n3858), .A1(n4497), .Z(n3792));
Q_AN02 U5028 ( .A0(n3858), .A1(n4496), .Z(n3791));
Q_AN02 U5029 ( .A0(n3858), .A1(n4495), .Z(n3790));
Q_AN02 U5030 ( .A0(n3858), .A1(n4494), .Z(n3789));
Q_AN02 U5031 ( .A0(n3858), .A1(n4493), .Z(n3788));
Q_AN02 U5032 ( .A0(n3858), .A1(n4492), .Z(n3787));
Q_AN02 U5033 ( .A0(n3858), .A1(n4491), .Z(n3786));
Q_AN02 U5034 ( .A0(n3858), .A1(n4490), .Z(n3785));
Q_AN02 U5035 ( .A0(n3858), .A1(n4489), .Z(n3784));
Q_AN02 U5036 ( .A0(n3858), .A1(n4488), .Z(n3783));
Q_AN02 U5037 ( .A0(n3858), .A1(n4487), .Z(n3782));
Q_AN02 U5038 ( .A0(n3858), .A1(n4486), .Z(n3781));
Q_AN02 U5039 ( .A0(n3858), .A1(n4485), .Z(n3780));
Q_AN02 U5040 ( .A0(n3858), .A1(n4484), .Z(n3779));
Q_AN02 U5041 ( .A0(n3858), .A1(n4483), .Z(n3778));
Q_AN02 U5042 ( .A0(n3858), .A1(n4482), .Z(n3777));
Q_AN02 U5043 ( .A0(n3858), .A1(n4481), .Z(n3776));
Q_AN02 U5044 ( .A0(n3858), .A1(n4480), .Z(n3775));
Q_AN02 U5045 ( .A0(n3858), .A1(n4479), .Z(n3774));
Q_AN02 U5046 ( .A0(n3858), .A1(n4478), .Z(n3773));
Q_AN02 U5047 ( .A0(n3858), .A1(n4477), .Z(n3772));
Q_AN02 U5048 ( .A0(n3858), .A1(n4476), .Z(n3771));
Q_AN02 U5049 ( .A0(n3858), .A1(n4475), .Z(n3770));
Q_AN02 U5050 ( .A0(n3858), .A1(n4474), .Z(n3769));
Q_AN02 U5051 ( .A0(n3858), .A1(n4473), .Z(n3768));
Q_AN02 U5052 ( .A0(n3858), .A1(n4472), .Z(n3767));
Q_AN02 U5053 ( .A0(n3858), .A1(n4471), .Z(n3766));
Q_AN02 U5054 ( .A0(n3858), .A1(n4470), .Z(n3765));
Q_AN02 U5055 ( .A0(n3858), .A1(n4469), .Z(n3764));
Q_AN02 U5056 ( .A0(n3858), .A1(n4468), .Z(n3763));
Q_AN02 U5057 ( .A0(n3858), .A1(n4467), .Z(n3762));
Q_AN02 U5058 ( .A0(n3858), .A1(n4466), .Z(n3761));
Q_AN02 U5059 ( .A0(n3858), .A1(n4465), .Z(n3760));
Q_AN02 U5060 ( .A0(n3858), .A1(n4464), .Z(n3759));
Q_AN02 U5061 ( .A0(n3858), .A1(n4463), .Z(n3758));
Q_AN02 U5062 ( .A0(n3858), .A1(n4462), .Z(n3757));
Q_AN02 U5063 ( .A0(n3858), .A1(n4461), .Z(n3756));
Q_AN02 U5064 ( .A0(n3858), .A1(n4460), .Z(n3755));
Q_AN02 U5065 ( .A0(n3858), .A1(n4459), .Z(n3754));
Q_AN02 U5066 ( .A0(n3858), .A1(n4458), .Z(n3753));
Q_AN02 U5067 ( .A0(n3858), .A1(n4457), .Z(n3752));
Q_AN02 U5068 ( .A0(n3858), .A1(n4456), .Z(n3751));
Q_AN02 U5069 ( .A0(n3858), .A1(n4455), .Z(n3750));
Q_AN02 U5070 ( .A0(n3858), .A1(n4454), .Z(n3749));
Q_AN02 U5071 ( .A0(n3858), .A1(n4453), .Z(n3748));
Q_AN02 U5072 ( .A0(n3858), .A1(n4452), .Z(n3747));
Q_AN02 U5073 ( .A0(n3858), .A1(n4451), .Z(n3746));
Q_AN02 U5074 ( .A0(n3858), .A1(n4450), .Z(n3745));
Q_AN02 U5075 ( .A0(n3858), .A1(n4449), .Z(n3744));
Q_AN02 U5076 ( .A0(n3858), .A1(n4448), .Z(n3743));
Q_AN02 U5077 ( .A0(n3858), .A1(n4447), .Z(n3742));
Q_AN02 U5078 ( .A0(n3858), .A1(n4446), .Z(n3741));
Q_AN02 U5079 ( .A0(n3858), .A1(n4445), .Z(n3740));
Q_AN02 U5080 ( .A0(n3858), .A1(n4444), .Z(n3739));
Q_AN02 U5081 ( .A0(n3858), .A1(n4443), .Z(n3738));
Q_AN02 U5082 ( .A0(n3858), .A1(n4442), .Z(n3737));
Q_AN02 U5083 ( .A0(n3858), .A1(n4441), .Z(n3736));
Q_AN02 U5084 ( .A0(n3858), .A1(n4440), .Z(n3735));
Q_AN02 U5085 ( .A0(n3858), .A1(n4439), .Z(n3734));
Q_AN02 U5086 ( .A0(n3858), .A1(n4438), .Z(n3733));
Q_AN02 U5087 ( .A0(n3858), .A1(n4437), .Z(n3732));
Q_AN02 U5088 ( .A0(n3858), .A1(n4436), .Z(n3731));
Q_AN02 U5089 ( .A0(n3858), .A1(n4435), .Z(n3730));
Q_OR02 U5090 ( .A0(n3729), .A1(n3730), .Z(n3256));
Q_OR02 U5091 ( .A0(n3728), .A1(n3731), .Z(n3253));
Q_OR02 U5092 ( .A0(n3727), .A1(n3732), .Z(n3250));
Q_OR02 U5093 ( .A0(n3726), .A1(n3733), .Z(n3247));
Q_OR02 U5094 ( .A0(n3725), .A1(n3734), .Z(n3244));
Q_OR02 U5095 ( .A0(n3724), .A1(n3735), .Z(n3241));
Q_OR02 U5096 ( .A0(n3723), .A1(n3736), .Z(n3238));
Q_OR02 U5097 ( .A0(n3722), .A1(n3737), .Z(n3235));
Q_OR02 U5098 ( .A0(n3721), .A1(n3738), .Z(n3232));
Q_OR02 U5099 ( .A0(n3720), .A1(n3739), .Z(n3229));
Q_OR02 U5100 ( .A0(n3719), .A1(n3740), .Z(n3226));
Q_OR02 U5101 ( .A0(n3718), .A1(n3741), .Z(n3223));
Q_OR02 U5102 ( .A0(n3717), .A1(n3742), .Z(n3220));
Q_OR02 U5103 ( .A0(n3716), .A1(n3743), .Z(n3217));
Q_OR02 U5104 ( .A0(n3715), .A1(n3744), .Z(n3214));
Q_OR02 U5105 ( .A0(n3714), .A1(n3745), .Z(n3211));
Q_OR02 U5106 ( .A0(n3713), .A1(n3746), .Z(n3208));
Q_OR02 U5107 ( .A0(n3712), .A1(n3747), .Z(n3205));
Q_OR02 U5108 ( .A0(n3711), .A1(n3748), .Z(n3202));
Q_OR02 U5109 ( .A0(n3710), .A1(n3749), .Z(n3199));
Q_OR02 U5110 ( .A0(n3709), .A1(n3750), .Z(n3196));
Q_OR02 U5111 ( .A0(n3708), .A1(n3751), .Z(n3193));
Q_OR02 U5112 ( .A0(n3707), .A1(n3752), .Z(n3190));
Q_OR02 U5113 ( .A0(n3706), .A1(n3753), .Z(n3187));
Q_OR02 U5114 ( .A0(n3705), .A1(n3754), .Z(n3184));
Q_OR02 U5115 ( .A0(n3704), .A1(n3755), .Z(n3181));
Q_OR02 U5116 ( .A0(n3703), .A1(n3756), .Z(n3178));
Q_OR02 U5117 ( .A0(n3702), .A1(n3757), .Z(n3175));
Q_OR02 U5118 ( .A0(n3701), .A1(n3758), .Z(n3172));
Q_OR02 U5119 ( .A0(n3700), .A1(n3759), .Z(n3169));
Q_OR02 U5120 ( .A0(n3699), .A1(n3760), .Z(n3166));
Q_OR02 U5121 ( .A0(n3698), .A1(n3761), .Z(n3163));
Q_OR02 U5122 ( .A0(n3697), .A1(n3762), .Z(n3160));
Q_OR02 U5123 ( .A0(n3696), .A1(n3763), .Z(n3157));
Q_OR02 U5124 ( .A0(n3695), .A1(n3764), .Z(n3154));
Q_OR02 U5125 ( .A0(n3694), .A1(n3765), .Z(n3151));
Q_OR02 U5126 ( .A0(n3693), .A1(n3766), .Z(n3148));
Q_OR02 U5127 ( .A0(n3692), .A1(n3767), .Z(n3145));
Q_OR02 U5128 ( .A0(n3691), .A1(n3768), .Z(n3142));
Q_OR02 U5129 ( .A0(n3690), .A1(n3769), .Z(n3139));
Q_OR02 U5130 ( .A0(n3689), .A1(n3770), .Z(n3136));
Q_OR02 U5131 ( .A0(n3688), .A1(n3771), .Z(n3133));
Q_OR02 U5132 ( .A0(n3687), .A1(n3772), .Z(n3130));
Q_OR02 U5133 ( .A0(n3686), .A1(n3773), .Z(n3127));
Q_OR02 U5134 ( .A0(n3685), .A1(n3774), .Z(n3124));
Q_OR02 U5135 ( .A0(n3684), .A1(n3775), .Z(n3121));
Q_OR02 U5136 ( .A0(n3683), .A1(n3776), .Z(n3118));
Q_OR02 U5137 ( .A0(n3682), .A1(n3777), .Z(n3115));
Q_OR02 U5138 ( .A0(n3681), .A1(n3778), .Z(n3112));
Q_OR02 U5139 ( .A0(n3680), .A1(n3779), .Z(n3109));
Q_OR02 U5140 ( .A0(n3679), .A1(n3780), .Z(n3106));
Q_OR02 U5141 ( .A0(n3678), .A1(n3781), .Z(n3103));
Q_OR02 U5142 ( .A0(n3677), .A1(n3782), .Z(n3100));
Q_OR02 U5143 ( .A0(n3676), .A1(n3783), .Z(n3097));
Q_OR02 U5144 ( .A0(n3675), .A1(n3784), .Z(n3094));
Q_OR02 U5145 ( .A0(n3674), .A1(n3785), .Z(n3091));
Q_OR02 U5146 ( .A0(n3673), .A1(n3786), .Z(n3088));
Q_OR02 U5147 ( .A0(n3672), .A1(n3787), .Z(n3085));
Q_OR02 U5148 ( .A0(n3671), .A1(n3788), .Z(n3082));
Q_OR02 U5149 ( .A0(n3670), .A1(n3789), .Z(n3079));
Q_OR02 U5150 ( .A0(n3669), .A1(n3790), .Z(n3076));
Q_OR02 U5151 ( .A0(n3668), .A1(n3791), .Z(n3073));
Q_OR02 U5152 ( .A0(n3667), .A1(n3792), .Z(n3070));
Q_OR02 U5153 ( .A0(n3666), .A1(n3793), .Z(n3067));
Q_OR02 U5154 ( .A0(n3665), .A1(n3794), .Z(n3064));
Q_OR02 U5155 ( .A0(n3664), .A1(n3795), .Z(n3061));
Q_OR02 U5156 ( .A0(n3663), .A1(n3796), .Z(n3058));
Q_OR02 U5157 ( .A0(n3662), .A1(n3797), .Z(n3055));
Q_OR02 U5158 ( .A0(n3661), .A1(n3798), .Z(n3052));
Q_OR02 U5159 ( .A0(n3660), .A1(n3799), .Z(n3049));
Q_OR02 U5160 ( .A0(n3659), .A1(n3800), .Z(n3046));
Q_OR02 U5161 ( .A0(n3658), .A1(n3801), .Z(n3043));
Q_OR02 U5162 ( .A0(n3657), .A1(n3802), .Z(n3040));
Q_OR02 U5163 ( .A0(n3656), .A1(n3803), .Z(n3037));
Q_OR02 U5164 ( .A0(n3655), .A1(n3804), .Z(n3034));
Q_OR02 U5165 ( .A0(n3654), .A1(n3805), .Z(n3031));
Q_OR02 U5166 ( .A0(n3653), .A1(n3806), .Z(n3028));
Q_OR02 U5167 ( .A0(n3652), .A1(n3807), .Z(n3025));
Q_OR02 U5168 ( .A0(n3651), .A1(n3808), .Z(n3022));
Q_OR02 U5169 ( .A0(n3650), .A1(n3809), .Z(n3019));
Q_OR02 U5170 ( .A0(n3649), .A1(n3810), .Z(n3016));
Q_OR02 U5171 ( .A0(n3648), .A1(n3811), .Z(n3013));
Q_OR02 U5172 ( .A0(n3647), .A1(n3812), .Z(n3010));
Q_OR02 U5173 ( .A0(n3646), .A1(n3813), .Z(n3007));
Q_OR02 U5174 ( .A0(n3645), .A1(n3814), .Z(n3004));
Q_OR02 U5175 ( .A0(n3644), .A1(n3815), .Z(n3001));
Q_OR02 U5176 ( .A0(n3643), .A1(n3816), .Z(n2998));
Q_OR02 U5177 ( .A0(n3642), .A1(n3817), .Z(n2995));
Q_OR02 U5178 ( .A0(n3641), .A1(n3818), .Z(n2992));
Q_OR02 U5179 ( .A0(n3640), .A1(n3819), .Z(n2989));
Q_OR02 U5180 ( .A0(n3639), .A1(n3820), .Z(n2986));
Q_OR02 U5181 ( .A0(n3638), .A1(n3821), .Z(n2983));
Q_OR02 U5182 ( .A0(n3637), .A1(n3822), .Z(n2980));
Q_OR02 U5183 ( .A0(n3636), .A1(n3823), .Z(n2977));
Q_OR02 U5184 ( .A0(n3635), .A1(n3824), .Z(n2974));
Q_OR02 U5185 ( .A0(n3634), .A1(n3825), .Z(n2971));
Q_OR02 U5186 ( .A0(n3633), .A1(n3826), .Z(n2968));
Q_OR02 U5187 ( .A0(n3632), .A1(n3827), .Z(n2965));
Q_OR02 U5188 ( .A0(n3631), .A1(n3828), .Z(n2962));
Q_OR02 U5189 ( .A0(n3630), .A1(n3829), .Z(n2959));
Q_OR02 U5190 ( .A0(n3629), .A1(n3830), .Z(n2956));
Q_OR02 U5191 ( .A0(n3628), .A1(n3831), .Z(n2953));
Q_OR02 U5192 ( .A0(n3627), .A1(n3832), .Z(n2950));
Q_OR02 U5193 ( .A0(n3626), .A1(n3833), .Z(n2947));
Q_OR02 U5194 ( .A0(n3625), .A1(n3834), .Z(n2944));
Q_OR02 U5195 ( .A0(n3624), .A1(n3835), .Z(n2941));
Q_OR02 U5196 ( .A0(n3623), .A1(n3836), .Z(n2938));
Q_OR02 U5197 ( .A0(n3622), .A1(n3837), .Z(n2935));
Q_OR02 U5198 ( .A0(n3621), .A1(n3838), .Z(n2932));
Q_OR02 U5199 ( .A0(n3620), .A1(n3839), .Z(n2929));
Q_OR02 U5200 ( .A0(n3619), .A1(n3840), .Z(n2926));
Q_OR02 U5201 ( .A0(n3618), .A1(n3841), .Z(n2923));
Q_OR02 U5202 ( .A0(n3617), .A1(n3842), .Z(n2920));
Q_OR02 U5203 ( .A0(n3616), .A1(n3843), .Z(n2917));
Q_OR02 U5204 ( .A0(n3615), .A1(n3844), .Z(n2914));
Q_OR02 U5205 ( .A0(n3614), .A1(n3845), .Z(n2911));
Q_OR02 U5206 ( .A0(n3613), .A1(n3846), .Z(n2908));
Q_OR02 U5207 ( .A0(n3612), .A1(n3847), .Z(n2905));
Q_OR02 U5208 ( .A0(n3611), .A1(n3848), .Z(n2902));
Q_OR02 U5209 ( .A0(n3610), .A1(n3849), .Z(n2899));
Q_OR02 U5210 ( .A0(n3609), .A1(n3850), .Z(n2896));
Q_OR02 U5211 ( .A0(n3608), .A1(n3851), .Z(n2893));
Q_OR02 U5212 ( .A0(n3607), .A1(n3852), .Z(n2890));
Q_OR02 U5213 ( .A0(n3606), .A1(n3853), .Z(n2887));
Q_OR02 U5214 ( .A0(n3605), .A1(n3854), .Z(n2884));
Q_OR02 U5215 ( .A0(n3604), .A1(n3855), .Z(n2881));
Q_OR02 U5216 ( .A0(n3603), .A1(n3856), .Z(n2878));
Q_OR02 U5217 ( .A0(n3602), .A1(n3857), .Z(n2875));
Q_OR02 U5218 ( .A0(n3601), .A1(n3859), .Z(n2872));
Q_OR02 U5219 ( .A0(n3600), .A1(n3860), .Z(n2869));
Q_OR02 U5220 ( .A0(n3599), .A1(n3861), .Z(n2866));
Q_OR02 U5221 ( .A0(n3598), .A1(n3862), .Z(n2863));
Q_OR02 U5222 ( .A0(n3597), .A1(n3863), .Z(n2860));
Q_OR02 U5223 ( .A0(n3596), .A1(n3864), .Z(n2857));
Q_OR02 U5224 ( .A0(n3595), .A1(n3865), .Z(n2854));
Q_OR02 U5225 ( .A0(n3594), .A1(n3866), .Z(n2851));
Q_OR02 U5226 ( .A0(n3593), .A1(n3867), .Z(n2848));
Q_OR02 U5227 ( .A0(n3592), .A1(n3868), .Z(n2845));
Q_OR02 U5228 ( .A0(n3591), .A1(n3869), .Z(n2842));
Q_OR02 U5229 ( .A0(n3590), .A1(n3870), .Z(n2839));
Q_OR02 U5230 ( .A0(n3589), .A1(n3871), .Z(n2836));
Q_OR02 U5231 ( .A0(n3588), .A1(n3872), .Z(n2833));
Q_OR02 U5232 ( .A0(n3587), .A1(n3873), .Z(n2830));
Q_OR02 U5233 ( .A0(n3586), .A1(n3874), .Z(n2827));
Q_OR02 U5234 ( .A0(n3585), .A1(n3875), .Z(n2824));
Q_OR02 U5235 ( .A0(n3584), .A1(n3876), .Z(n2821));
Q_OR02 U5236 ( .A0(n3583), .A1(n3877), .Z(n2818));
Q_OR02 U5237 ( .A0(n3582), .A1(n3878), .Z(n2815));
Q_OR02 U5238 ( .A0(n3581), .A1(n3879), .Z(n2812));
Q_OR02 U5239 ( .A0(n3580), .A1(n3880), .Z(n2809));
Q_OR02 U5240 ( .A0(n3579), .A1(n3881), .Z(n2806));
Q_OR02 U5241 ( .A0(n3578), .A1(n3882), .Z(n2803));
Q_OR02 U5242 ( .A0(n3577), .A1(n3883), .Z(n2800));
Q_OR02 U5243 ( .A0(n3576), .A1(n3884), .Z(n2797));
Q_OR02 U5244 ( .A0(n3575), .A1(n3885), .Z(n2794));
Q_OR02 U5245 ( .A0(n3574), .A1(n3886), .Z(n2791));
Q_OR02 U5246 ( .A0(n3573), .A1(n3887), .Z(n2788));
Q_OR02 U5247 ( .A0(n3572), .A1(n3888), .Z(n2785));
Q_OR02 U5248 ( .A0(n3571), .A1(n3889), .Z(n2782));
Q_OR02 U5249 ( .A0(n3570), .A1(n3890), .Z(n2779));
Q_OR02 U5250 ( .A0(n3569), .A1(n3891), .Z(n2776));
Q_OR02 U5251 ( .A0(n3568), .A1(n3892), .Z(n2773));
Q_OR02 U5252 ( .A0(n3567), .A1(n3893), .Z(n2770));
Q_OR02 U5253 ( .A0(n3566), .A1(n3894), .Z(n2767));
Q_OR02 U5254 ( .A0(n3565), .A1(n3895), .Z(n2764));
Q_OR02 U5255 ( .A0(n3564), .A1(n3896), .Z(n2761));
Q_OR02 U5256 ( .A0(n3563), .A1(n3897), .Z(n2758));
Q_OR02 U5257 ( .A0(n3562), .A1(n3898), .Z(n2755));
Q_OR02 U5258 ( .A0(n3561), .A1(n3899), .Z(n2752));
Q_OR02 U5259 ( .A0(n3560), .A1(n3900), .Z(n2749));
Q_OR02 U5260 ( .A0(n3559), .A1(n3901), .Z(n2746));
Q_OR02 U5261 ( .A0(n3558), .A1(n3902), .Z(n2743));
Q_OR02 U5262 ( .A0(n3557), .A1(n3903), .Z(n2740));
Q_OR02 U5263 ( .A0(n3556), .A1(n3904), .Z(n2737));
Q_OR02 U5264 ( .A0(n3555), .A1(n3905), .Z(n2734));
Q_OR02 U5265 ( .A0(n3554), .A1(n3906), .Z(n2731));
Q_OR02 U5266 ( .A0(n3553), .A1(n3907), .Z(n2728));
Q_OR02 U5267 ( .A0(n3552), .A1(n3908), .Z(n2725));
Q_OR02 U5268 ( .A0(n3551), .A1(n3909), .Z(n2722));
Q_OR02 U5269 ( .A0(n3550), .A1(n3910), .Z(n2719));
Q_OR02 U5270 ( .A0(n3549), .A1(n3911), .Z(n2716));
Q_OR02 U5271 ( .A0(n3548), .A1(n3912), .Z(n2713));
Q_OR02 U5272 ( .A0(n3547), .A1(n3913), .Z(n2710));
Q_OR02 U5273 ( .A0(n3546), .A1(n3914), .Z(n2707));
Q_OR02 U5274 ( .A0(n3545), .A1(n3915), .Z(n2704));
Q_OR02 U5275 ( .A0(n3544), .A1(n3916), .Z(n2701));
Q_OR02 U5276 ( .A0(n3543), .A1(n3917), .Z(n2698));
Q_OR02 U5277 ( .A0(n3542), .A1(n3918), .Z(n2695));
Q_OR02 U5278 ( .A0(n3541), .A1(n3919), .Z(n2692));
Q_OR02 U5279 ( .A0(n3540), .A1(n3920), .Z(n2689));
Q_OR02 U5280 ( .A0(n3539), .A1(n3921), .Z(n2686));
Q_OR02 U5281 ( .A0(n3538), .A1(n3922), .Z(n2683));
Q_OR02 U5282 ( .A0(n3537), .A1(n3923), .Z(n2680));
Q_OR02 U5283 ( .A0(n3536), .A1(n3924), .Z(n2677));
Q_OR02 U5284 ( .A0(n3535), .A1(n3925), .Z(n2674));
Q_OR02 U5285 ( .A0(n3534), .A1(n3926), .Z(n2671));
Q_OR02 U5286 ( .A0(n3533), .A1(n3927), .Z(n2668));
Q_OR02 U5287 ( .A0(n3532), .A1(n3928), .Z(n2665));
Q_OR02 U5288 ( .A0(n3531), .A1(n3929), .Z(n2662));
Q_OR02 U5289 ( .A0(n3530), .A1(n3930), .Z(n2659));
Q_OR02 U5290 ( .A0(n3529), .A1(n3931), .Z(n2656));
Q_OR02 U5291 ( .A0(n3528), .A1(n3932), .Z(n2653));
Q_OR02 U5292 ( .A0(n3527), .A1(n3933), .Z(n2650));
Q_OR02 U5293 ( .A0(n3526), .A1(n3934), .Z(n2647));
Q_OR02 U5294 ( .A0(n3525), .A1(n3935), .Z(n2644));
Q_OR02 U5295 ( .A0(n3524), .A1(n3936), .Z(n2641));
Q_OR02 U5296 ( .A0(n3523), .A1(n3937), .Z(n2638));
Q_OR02 U5297 ( .A0(n3522), .A1(n3938), .Z(n2635));
Q_OR02 U5298 ( .A0(n3521), .A1(n3939), .Z(n2632));
Q_OR02 U5299 ( .A0(n3520), .A1(n3940), .Z(n2629));
Q_OR02 U5300 ( .A0(n3519), .A1(n3941), .Z(n2626));
Q_OR02 U5301 ( .A0(n3518), .A1(n3942), .Z(n2623));
Q_OR02 U5302 ( .A0(n3517), .A1(n3943), .Z(n2620));
Q_OR02 U5303 ( .A0(n3516), .A1(n3944), .Z(n2617));
Q_OR02 U5304 ( .A0(n3515), .A1(n3945), .Z(n2614));
Q_OR02 U5305 ( .A0(n3514), .A1(n3946), .Z(n2611));
Q_OR02 U5306 ( .A0(n3513), .A1(n3947), .Z(n2608));
Q_OR02 U5307 ( .A0(n3512), .A1(n3948), .Z(n2605));
Q_OR02 U5308 ( .A0(n3511), .A1(n3949), .Z(n2602));
Q_OR02 U5309 ( .A0(n3510), .A1(n3950), .Z(n2599));
Q_OR02 U5310 ( .A0(n3509), .A1(n3951), .Z(n2596));
Q_OR02 U5311 ( .A0(n3508), .A1(n3952), .Z(n2593));
Q_OR02 U5312 ( .A0(n3507), .A1(n3953), .Z(n2590));
Q_OR02 U5313 ( .A0(n3506), .A1(n3954), .Z(n2587));
Q_OR02 U5314 ( .A0(n3505), .A1(n3955), .Z(n2584));
Q_OR02 U5315 ( .A0(n3504), .A1(n3956), .Z(n2581));
Q_OR02 U5316 ( .A0(n3503), .A1(n3957), .Z(n2578));
Q_OR02 U5317 ( .A0(n3502), .A1(n3958), .Z(n2575));
Q_OR02 U5318 ( .A0(n3501), .A1(n3959), .Z(n2572));
Q_OR02 U5319 ( .A0(n3500), .A1(n3960), .Z(n2569));
Q_OR02 U5320 ( .A0(n3499), .A1(n3961), .Z(n2566));
Q_OR02 U5321 ( .A0(n3498), .A1(n3962), .Z(n2563));
Q_OR02 U5322 ( .A0(n3497), .A1(n3963), .Z(n2560));
Q_OR02 U5323 ( .A0(n3496), .A1(n3964), .Z(n2557));
Q_OR02 U5324 ( .A0(n3495), .A1(n3965), .Z(n2554));
Q_OR02 U5325 ( .A0(n3494), .A1(n3966), .Z(n2551));
Q_OR02 U5326 ( .A0(n3493), .A1(n3967), .Z(n2548));
Q_OR02 U5327 ( .A0(n3492), .A1(n3968), .Z(n2545));
Q_OR02 U5328 ( .A0(n3491), .A1(n3969), .Z(n2542));
Q_OR02 U5329 ( .A0(n3490), .A1(n3970), .Z(n2539));
Q_OR02 U5330 ( .A0(n3489), .A1(n3971), .Z(n2536));
Q_OR02 U5331 ( .A0(n3488), .A1(n3972), .Z(n2533));
Q_OR02 U5332 ( .A0(n3487), .A1(n3973), .Z(n2530));
Q_OR02 U5333 ( .A0(n3486), .A1(n3974), .Z(n2527));
Q_OR02 U5334 ( .A0(n3485), .A1(n3975), .Z(n2524));
Q_OR02 U5335 ( .A0(n3484), .A1(n3976), .Z(n2521));
Q_OR02 U5336 ( .A0(n3483), .A1(n3977), .Z(n2518));
Q_OR02 U5337 ( .A0(n3482), .A1(n3978), .Z(n2515));
Q_OR02 U5338 ( .A0(n3481), .A1(n3979), .Z(n2512));
Q_OR02 U5339 ( .A0(n3480), .A1(n3980), .Z(n2509));
Q_OR02 U5340 ( .A0(n3479), .A1(n3981), .Z(n2506));
Q_OR02 U5341 ( .A0(n3478), .A1(n3982), .Z(n2503));
Q_OR02 U5342 ( .A0(n3477), .A1(n3983), .Z(n2500));
Q_OR02 U5343 ( .A0(n3476), .A1(n3984), .Z(n2497));
Q_OR02 U5344 ( .A0(n3475), .A1(n3985), .Z(n2494));
Q_OR02 U5345 ( .A0(n3474), .A1(n3986), .Z(n2491));
Q_OA21 U5346 ( .A0(n3730), .A1(ofifoData[0]), .B0(n278), .Z(n3255));
Q_OA21 U5347 ( .A0(n3731), .A1(ofifoData[1]), .B0(n278), .Z(n3252));
Q_OA21 U5348 ( .A0(n3732), .A1(ofifoData[2]), .B0(n278), .Z(n3249));
Q_OA21 U5349 ( .A0(n3733), .A1(ofifoData[3]), .B0(n278), .Z(n3246));
Q_OA21 U5350 ( .A0(n3734), .A1(ofifoData[4]), .B0(n278), .Z(n3243));
Q_OA21 U5351 ( .A0(n3735), .A1(ofifoData[5]), .B0(n278), .Z(n3240));
Q_OA21 U5352 ( .A0(n3736), .A1(ofifoData[6]), .B0(n278), .Z(n3237));
Q_OA21 U5353 ( .A0(n3737), .A1(ofifoData[7]), .B0(n278), .Z(n3234));
Q_OA21 U5354 ( .A0(n3738), .A1(ofifoData[8]), .B0(n278), .Z(n3231));
Q_OA21 U5355 ( .A0(n3739), .A1(ofifoData[9]), .B0(n278), .Z(n3228));
Q_OA21 U5356 ( .A0(n3740), .A1(ofifoData[10]), .B0(n278), .Z(n3225));
Q_OA21 U5357 ( .A0(n3741), .A1(ofifoData[11]), .B0(n278), .Z(n3222));
Q_OA21 U5358 ( .A0(n3742), .A1(ofifoData[12]), .B0(n278), .Z(n3219));
Q_OA21 U5359 ( .A0(n3743), .A1(ofifoData[13]), .B0(n278), .Z(n3216));
Q_OA21 U5360 ( .A0(n3744), .A1(ofifoData[14]), .B0(n278), .Z(n3213));
Q_OA21 U5361 ( .A0(n3745), .A1(ofifoData[15]), .B0(n278), .Z(n3210));
Q_OA21 U5362 ( .A0(n3746), .A1(ofifoData[16]), .B0(n278), .Z(n3207));
Q_OA21 U5363 ( .A0(n3747), .A1(ofifoData[17]), .B0(n278), .Z(n3204));
Q_OA21 U5364 ( .A0(n3748), .A1(ofifoData[18]), .B0(n278), .Z(n3201));
Q_OA21 U5365 ( .A0(n3749), .A1(ofifoData[19]), .B0(n278), .Z(n3198));
Q_OA21 U5366 ( .A0(n3750), .A1(ofifoData[20]), .B0(n278), .Z(n3195));
Q_OA21 U5367 ( .A0(n3751), .A1(ofifoData[21]), .B0(n278), .Z(n3192));
Q_OA21 U5368 ( .A0(n3752), .A1(ofifoData[22]), .B0(n278), .Z(n3189));
Q_OA21 U5369 ( .A0(n3753), .A1(ofifoData[23]), .B0(n278), .Z(n3186));
Q_OA21 U5370 ( .A0(n3754), .A1(ofifoData[24]), .B0(n278), .Z(n3183));
Q_OA21 U5371 ( .A0(n3755), .A1(ofifoData[25]), .B0(n278), .Z(n3180));
Q_OA21 U5372 ( .A0(n3756), .A1(ofifoData[26]), .B0(n278), .Z(n3177));
Q_OA21 U5373 ( .A0(n3757), .A1(ofifoData[27]), .B0(n278), .Z(n3174));
Q_OA21 U5374 ( .A0(n3758), .A1(ofifoData[28]), .B0(n278), .Z(n3171));
Q_OA21 U5375 ( .A0(n3759), .A1(ofifoData[29]), .B0(n278), .Z(n3168));
Q_OA21 U5376 ( .A0(n3760), .A1(ofifoData[30]), .B0(n278), .Z(n3165));
Q_OA21 U5377 ( .A0(n3761), .A1(ofifoData[31]), .B0(n278), .Z(n3162));
Q_OA21 U5378 ( .A0(n3762), .A1(ofifoData[32]), .B0(n278), .Z(n3159));
Q_OA21 U5379 ( .A0(n3763), .A1(ofifoData[33]), .B0(n278), .Z(n3156));
Q_OA21 U5380 ( .A0(n3764), .A1(ofifoData[34]), .B0(n278), .Z(n3153));
Q_OA21 U5381 ( .A0(n3765), .A1(ofifoData[35]), .B0(n278), .Z(n3150));
Q_OA21 U5382 ( .A0(n3766), .A1(ofifoData[36]), .B0(n278), .Z(n3147));
Q_OA21 U5383 ( .A0(n3767), .A1(ofifoData[37]), .B0(n278), .Z(n3144));
Q_OA21 U5384 ( .A0(n3768), .A1(ofifoData[38]), .B0(n278), .Z(n3141));
Q_OA21 U5385 ( .A0(n3769), .A1(ofifoData[39]), .B0(n278), .Z(n3138));
Q_OA21 U5386 ( .A0(n3770), .A1(ofifoData[40]), .B0(n278), .Z(n3135));
Q_OA21 U5387 ( .A0(n3771), .A1(ofifoData[41]), .B0(n278), .Z(n3132));
Q_OA21 U5388 ( .A0(n3772), .A1(ofifoData[42]), .B0(n278), .Z(n3129));
Q_OA21 U5389 ( .A0(n3773), .A1(ofifoData[43]), .B0(n278), .Z(n3126));
Q_OA21 U5390 ( .A0(n3774), .A1(ofifoData[44]), .B0(n278), .Z(n3123));
Q_OA21 U5391 ( .A0(n3775), .A1(ofifoData[45]), .B0(n278), .Z(n3120));
Q_OA21 U5392 ( .A0(n3776), .A1(ofifoData[46]), .B0(n278), .Z(n3117));
Q_OA21 U5393 ( .A0(n3777), .A1(ofifoData[47]), .B0(n278), .Z(n3114));
Q_OA21 U5394 ( .A0(n3778), .A1(ofifoData[48]), .B0(n278), .Z(n3111));
Q_OA21 U5395 ( .A0(n3779), .A1(ofifoData[49]), .B0(n278), .Z(n3108));
Q_OA21 U5396 ( .A0(n3780), .A1(ofifoData[50]), .B0(n278), .Z(n3105));
Q_OA21 U5397 ( .A0(n3781), .A1(ofifoData[51]), .B0(n278), .Z(n3102));
Q_OA21 U5398 ( .A0(n3782), .A1(ofifoData[52]), .B0(n278), .Z(n3099));
Q_OA21 U5399 ( .A0(n3783), .A1(ofifoData[53]), .B0(n278), .Z(n3096));
Q_OA21 U5400 ( .A0(n3784), .A1(ofifoData[54]), .B0(n278), .Z(n3093));
Q_OA21 U5401 ( .A0(n3785), .A1(ofifoData[55]), .B0(n278), .Z(n3090));
Q_OA21 U5402 ( .A0(n3786), .A1(ofifoData[56]), .B0(n278), .Z(n3087));
Q_OA21 U5403 ( .A0(n3787), .A1(ofifoData[57]), .B0(n278), .Z(n3084));
Q_OA21 U5404 ( .A0(n3788), .A1(ofifoData[58]), .B0(n278), .Z(n3081));
Q_OA21 U5405 ( .A0(n3789), .A1(ofifoData[59]), .B0(n278), .Z(n3078));
Q_OA21 U5406 ( .A0(n3790), .A1(ofifoData[60]), .B0(n278), .Z(n3075));
Q_OA21 U5407 ( .A0(n3791), .A1(ofifoData[61]), .B0(n278), .Z(n3072));
Q_OA21 U5408 ( .A0(n3792), .A1(ofifoData[62]), .B0(n278), .Z(n3069));
Q_OA21 U5409 ( .A0(n3793), .A1(ofifoData[63]), .B0(n278), .Z(n3066));
Q_OA21 U5410 ( .A0(n3794), .A1(ofifoData[64]), .B0(n278), .Z(n3063));
Q_OA21 U5411 ( .A0(n3795), .A1(ofifoData[65]), .B0(n278), .Z(n3060));
Q_OA21 U5412 ( .A0(n3796), .A1(ofifoData[66]), .B0(n278), .Z(n3057));
Q_OA21 U5413 ( .A0(n3797), .A1(ofifoData[67]), .B0(n278), .Z(n3054));
Q_OA21 U5414 ( .A0(n3798), .A1(ofifoData[68]), .B0(n278), .Z(n3051));
Q_OA21 U5415 ( .A0(n3799), .A1(ofifoData[69]), .B0(n278), .Z(n3048));
Q_OA21 U5416 ( .A0(n3800), .A1(ofifoData[70]), .B0(n278), .Z(n3045));
Q_OA21 U5417 ( .A0(n3801), .A1(ofifoData[71]), .B0(n278), .Z(n3042));
Q_OA21 U5418 ( .A0(n3802), .A1(ofifoData[72]), .B0(n278), .Z(n3039));
Q_OA21 U5419 ( .A0(n3803), .A1(ofifoData[73]), .B0(n278), .Z(n3036));
Q_OA21 U5420 ( .A0(n3804), .A1(ofifoData[74]), .B0(n278), .Z(n3033));
Q_OA21 U5421 ( .A0(n3805), .A1(ofifoData[75]), .B0(n278), .Z(n3030));
Q_OA21 U5422 ( .A0(n3806), .A1(ofifoData[76]), .B0(n278), .Z(n3027));
Q_OA21 U5423 ( .A0(n3807), .A1(ofifoData[77]), .B0(n278), .Z(n3024));
Q_OA21 U5424 ( .A0(n3808), .A1(ofifoData[78]), .B0(n278), .Z(n3021));
Q_OA21 U5425 ( .A0(n3809), .A1(ofifoData[79]), .B0(n278), .Z(n3018));
Q_OA21 U5426 ( .A0(n3810), .A1(ofifoData[80]), .B0(n278), .Z(n3015));
Q_OA21 U5427 ( .A0(n3811), .A1(ofifoData[81]), .B0(n278), .Z(n3012));
Q_OA21 U5428 ( .A0(n3812), .A1(ofifoData[82]), .B0(n278), .Z(n3009));
Q_OA21 U5429 ( .A0(n3813), .A1(ofifoData[83]), .B0(n278), .Z(n3006));
Q_OA21 U5430 ( .A0(n3814), .A1(ofifoData[84]), .B0(n278), .Z(n3003));
Q_OA21 U5431 ( .A0(n3815), .A1(ofifoData[85]), .B0(n278), .Z(n3000));
Q_OA21 U5432 ( .A0(n3816), .A1(ofifoData[86]), .B0(n278), .Z(n2997));
Q_OA21 U5433 ( .A0(n3817), .A1(ofifoData[87]), .B0(n278), .Z(n2994));
Q_OA21 U5434 ( .A0(n3818), .A1(ofifoData[88]), .B0(n278), .Z(n2991));
Q_OA21 U5435 ( .A0(n3819), .A1(ofifoData[89]), .B0(n278), .Z(n2988));
Q_OA21 U5436 ( .A0(n3820), .A1(ofifoData[90]), .B0(n278), .Z(n2985));
Q_OA21 U5437 ( .A0(n3821), .A1(ofifoData[91]), .B0(n278), .Z(n2982));
Q_OA21 U5438 ( .A0(n3822), .A1(ofifoData[92]), .B0(n278), .Z(n2979));
Q_OA21 U5439 ( .A0(n3823), .A1(ofifoData[93]), .B0(n278), .Z(n2976));
Q_OA21 U5440 ( .A0(n3824), .A1(ofifoData[94]), .B0(n278), .Z(n2973));
Q_OA21 U5441 ( .A0(n3825), .A1(ofifoData[95]), .B0(n278), .Z(n2970));
Q_OA21 U5442 ( .A0(n3826), .A1(ofifoData[96]), .B0(n278), .Z(n2967));
Q_OA21 U5443 ( .A0(n3827), .A1(ofifoData[97]), .B0(n278), .Z(n2964));
Q_OA21 U5444 ( .A0(n3828), .A1(ofifoData[98]), .B0(n278), .Z(n2961));
Q_OA21 U5445 ( .A0(n3829), .A1(ofifoData[99]), .B0(n278), .Z(n2958));
Q_OA21 U5446 ( .A0(n3830), .A1(ofifoData[100]), .B0(n278), .Z(n2955));
Q_OA21 U5447 ( .A0(n3831), .A1(ofifoData[101]), .B0(n278), .Z(n2952));
Q_OA21 U5448 ( .A0(n3832), .A1(ofifoData[102]), .B0(n278), .Z(n2949));
Q_OA21 U5449 ( .A0(n3833), .A1(ofifoData[103]), .B0(n278), .Z(n2946));
Q_OA21 U5450 ( .A0(n3834), .A1(ofifoData[104]), .B0(n278), .Z(n2943));
Q_OA21 U5451 ( .A0(n3835), .A1(ofifoData[105]), .B0(n278), .Z(n2940));
Q_OA21 U5452 ( .A0(n3836), .A1(ofifoData[106]), .B0(n278), .Z(n2937));
Q_OA21 U5453 ( .A0(n3837), .A1(ofifoData[107]), .B0(n278), .Z(n2934));
Q_OA21 U5454 ( .A0(n3838), .A1(ofifoData[108]), .B0(n278), .Z(n2931));
Q_OA21 U5455 ( .A0(n3839), .A1(ofifoData[109]), .B0(n278), .Z(n2928));
Q_OA21 U5456 ( .A0(n3840), .A1(ofifoData[110]), .B0(n278), .Z(n2925));
Q_OA21 U5457 ( .A0(n3841), .A1(ofifoData[111]), .B0(n278), .Z(n2922));
Q_OA21 U5458 ( .A0(n3842), .A1(ofifoData[112]), .B0(n278), .Z(n2919));
Q_OA21 U5459 ( .A0(n3843), .A1(ofifoData[113]), .B0(n278), .Z(n2916));
Q_OA21 U5460 ( .A0(n3844), .A1(ofifoData[114]), .B0(n278), .Z(n2913));
Q_OA21 U5461 ( .A0(n3845), .A1(ofifoData[115]), .B0(n278), .Z(n2910));
Q_OA21 U5462 ( .A0(n3846), .A1(ofifoData[116]), .B0(n278), .Z(n2907));
Q_OA21 U5463 ( .A0(n3847), .A1(ofifoData[117]), .B0(n278), .Z(n2904));
Q_OA21 U5464 ( .A0(n3848), .A1(ofifoData[118]), .B0(n278), .Z(n2901));
Q_OA21 U5465 ( .A0(n3849), .A1(ofifoData[119]), .B0(n278), .Z(n2898));
Q_OA21 U5466 ( .A0(n3850), .A1(ofifoData[120]), .B0(n278), .Z(n2895));
Q_OA21 U5467 ( .A0(n3851), .A1(ofifoData[121]), .B0(n278), .Z(n2892));
Q_OA21 U5468 ( .A0(n3852), .A1(ofifoData[122]), .B0(n278), .Z(n2889));
Q_OA21 U5469 ( .A0(n3853), .A1(ofifoData[123]), .B0(n278), .Z(n2886));
Q_OA21 U5470 ( .A0(n3854), .A1(ofifoData[124]), .B0(n278), .Z(n2883));
Q_OA21 U5471 ( .A0(n3855), .A1(ofifoData[125]), .B0(n278), .Z(n2880));
Q_OA21 U5472 ( .A0(n3856), .A1(ofifoData[126]), .B0(n278), .Z(n2877));
Q_OA21 U5473 ( .A0(n3857), .A1(ofifoData[127]), .B0(n278), .Z(n2874));
Q_OA21 U5474 ( .A0(n3859), .A1(ofifoData[128]), .B0(n278), .Z(n2871));
Q_OA21 U5475 ( .A0(n3860), .A1(ofifoData[129]), .B0(n278), .Z(n2868));
Q_OA21 U5476 ( .A0(n3861), .A1(ofifoData[130]), .B0(n278), .Z(n2865));
Q_OA21 U5477 ( .A0(n3862), .A1(ofifoData[131]), .B0(n278), .Z(n2862));
Q_OA21 U5478 ( .A0(n3863), .A1(ofifoData[132]), .B0(n278), .Z(n2859));
Q_OA21 U5479 ( .A0(n3864), .A1(ofifoData[133]), .B0(n278), .Z(n2856));
Q_OA21 U5480 ( .A0(n3865), .A1(ofifoData[134]), .B0(n278), .Z(n2853));
Q_OA21 U5481 ( .A0(n3866), .A1(ofifoData[135]), .B0(n278), .Z(n2850));
Q_OA21 U5482 ( .A0(n3867), .A1(ofifoData[136]), .B0(n278), .Z(n2847));
Q_OA21 U5483 ( .A0(n3868), .A1(ofifoData[137]), .B0(n278), .Z(n2844));
Q_OA21 U5484 ( .A0(n3869), .A1(ofifoData[138]), .B0(n278), .Z(n2841));
Q_OA21 U5485 ( .A0(n3870), .A1(ofifoData[139]), .B0(n278), .Z(n2838));
Q_OA21 U5486 ( .A0(n3871), .A1(ofifoData[140]), .B0(n278), .Z(n2835));
Q_OA21 U5487 ( .A0(n3872), .A1(ofifoData[141]), .B0(n278), .Z(n2832));
Q_OA21 U5488 ( .A0(n3873), .A1(ofifoData[142]), .B0(n278), .Z(n2829));
Q_OA21 U5489 ( .A0(n3874), .A1(ofifoData[143]), .B0(n278), .Z(n2826));
Q_OA21 U5490 ( .A0(n3875), .A1(ofifoData[144]), .B0(n278), .Z(n2823));
Q_OA21 U5491 ( .A0(n3876), .A1(ofifoData[145]), .B0(n278), .Z(n2820));
Q_OA21 U5492 ( .A0(n3877), .A1(ofifoData[146]), .B0(n278), .Z(n2817));
Q_OA21 U5493 ( .A0(n3878), .A1(ofifoData[147]), .B0(n278), .Z(n2814));
Q_OA21 U5494 ( .A0(n3879), .A1(ofifoData[148]), .B0(n278), .Z(n2811));
Q_OA21 U5495 ( .A0(n3880), .A1(ofifoData[149]), .B0(n278), .Z(n2808));
Q_OA21 U5496 ( .A0(n3881), .A1(ofifoData[150]), .B0(n278), .Z(n2805));
Q_OA21 U5497 ( .A0(n3882), .A1(ofifoData[151]), .B0(n278), .Z(n2802));
Q_OA21 U5498 ( .A0(n3883), .A1(ofifoData[152]), .B0(n278), .Z(n2799));
Q_OA21 U5499 ( .A0(n3884), .A1(ofifoData[153]), .B0(n278), .Z(n2796));
Q_OA21 U5500 ( .A0(n3885), .A1(ofifoData[154]), .B0(n278), .Z(n2793));
Q_OA21 U5501 ( .A0(n3886), .A1(ofifoData[155]), .B0(n278), .Z(n2790));
Q_OA21 U5502 ( .A0(n3887), .A1(ofifoData[156]), .B0(n278), .Z(n2787));
Q_OA21 U5503 ( .A0(n3888), .A1(ofifoData[157]), .B0(n278), .Z(n2784));
Q_OA21 U5504 ( .A0(n3889), .A1(ofifoData[158]), .B0(n278), .Z(n2781));
Q_OA21 U5505 ( .A0(n3890), .A1(ofifoData[159]), .B0(n278), .Z(n2778));
Q_OA21 U5506 ( .A0(n3891), .A1(ofifoData[160]), .B0(n278), .Z(n2775));
Q_OA21 U5507 ( .A0(n3892), .A1(ofifoData[161]), .B0(n278), .Z(n2772));
Q_OA21 U5508 ( .A0(n3893), .A1(ofifoData[162]), .B0(n278), .Z(n2769));
Q_OA21 U5509 ( .A0(n3894), .A1(ofifoData[163]), .B0(n278), .Z(n2766));
Q_OA21 U5510 ( .A0(n3895), .A1(ofifoData[164]), .B0(n278), .Z(n2763));
Q_OA21 U5511 ( .A0(n3896), .A1(ofifoData[165]), .B0(n278), .Z(n2760));
Q_OA21 U5512 ( .A0(n3897), .A1(ofifoData[166]), .B0(n278), .Z(n2757));
Q_OA21 U5513 ( .A0(n3898), .A1(ofifoData[167]), .B0(n278), .Z(n2754));
Q_OA21 U5514 ( .A0(n3899), .A1(ofifoData[168]), .B0(n278), .Z(n2751));
Q_OA21 U5515 ( .A0(n3900), .A1(ofifoData[169]), .B0(n278), .Z(n2748));
Q_OA21 U5516 ( .A0(n3901), .A1(ofifoData[170]), .B0(n278), .Z(n2745));
Q_OA21 U5517 ( .A0(n3902), .A1(ofifoData[171]), .B0(n278), .Z(n2742));
Q_OA21 U5518 ( .A0(n3903), .A1(ofifoData[172]), .B0(n278), .Z(n2739));
Q_OA21 U5519 ( .A0(n3904), .A1(ofifoData[173]), .B0(n278), .Z(n2736));
Q_OA21 U5520 ( .A0(n3905), .A1(ofifoData[174]), .B0(n278), .Z(n2733));
Q_OA21 U5521 ( .A0(n3906), .A1(ofifoData[175]), .B0(n278), .Z(n2730));
Q_OA21 U5522 ( .A0(n3907), .A1(ofifoData[176]), .B0(n278), .Z(n2727));
Q_OA21 U5523 ( .A0(n3908), .A1(ofifoData[177]), .B0(n278), .Z(n2724));
Q_OA21 U5524 ( .A0(n3909), .A1(ofifoData[178]), .B0(n278), .Z(n2721));
Q_OA21 U5525 ( .A0(n3910), .A1(ofifoData[179]), .B0(n278), .Z(n2718));
Q_OA21 U5526 ( .A0(n3911), .A1(ofifoData[180]), .B0(n278), .Z(n2715));
Q_OA21 U5527 ( .A0(n3912), .A1(ofifoData[181]), .B0(n278), .Z(n2712));
Q_OA21 U5528 ( .A0(n3913), .A1(ofifoData[182]), .B0(n278), .Z(n2709));
Q_OA21 U5529 ( .A0(n3914), .A1(ofifoData[183]), .B0(n278), .Z(n2706));
Q_OA21 U5530 ( .A0(n3915), .A1(ofifoData[184]), .B0(n278), .Z(n2703));
Q_OA21 U5531 ( .A0(n3916), .A1(ofifoData[185]), .B0(n278), .Z(n2700));
Q_OA21 U5532 ( .A0(n3917), .A1(ofifoData[186]), .B0(n278), .Z(n2697));
Q_OA21 U5533 ( .A0(n3918), .A1(ofifoData[187]), .B0(n278), .Z(n2694));
Q_OA21 U5534 ( .A0(n3919), .A1(ofifoData[188]), .B0(n278), .Z(n2691));
Q_OA21 U5535 ( .A0(n3920), .A1(ofifoData[189]), .B0(n278), .Z(n2688));
Q_OA21 U5536 ( .A0(n3921), .A1(ofifoData[190]), .B0(n278), .Z(n2685));
Q_OA21 U5537 ( .A0(n3922), .A1(ofifoData[191]), .B0(n278), .Z(n2682));
Q_OA21 U5538 ( .A0(n3923), .A1(ofifoData[192]), .B0(n278), .Z(n2679));
Q_OA21 U5539 ( .A0(n3924), .A1(ofifoData[193]), .B0(n278), .Z(n2676));
Q_OA21 U5540 ( .A0(n3925), .A1(ofifoData[194]), .B0(n278), .Z(n2673));
Q_OA21 U5541 ( .A0(n3926), .A1(ofifoData[195]), .B0(n278), .Z(n2670));
Q_OA21 U5542 ( .A0(n3927), .A1(ofifoData[196]), .B0(n278), .Z(n2667));
Q_OA21 U5543 ( .A0(n3928), .A1(ofifoData[197]), .B0(n278), .Z(n2664));
Q_OA21 U5544 ( .A0(n3929), .A1(ofifoData[198]), .B0(n278), .Z(n2661));
Q_OA21 U5545 ( .A0(n3930), .A1(ofifoData[199]), .B0(n278), .Z(n2658));
Q_OA21 U5546 ( .A0(n3931), .A1(ofifoData[200]), .B0(n278), .Z(n2655));
Q_OA21 U5547 ( .A0(n3932), .A1(ofifoData[201]), .B0(n278), .Z(n2652));
Q_OA21 U5548 ( .A0(n3933), .A1(ofifoData[202]), .B0(n278), .Z(n2649));
Q_OA21 U5549 ( .A0(n3934), .A1(ofifoData[203]), .B0(n278), .Z(n2646));
Q_OA21 U5550 ( .A0(n3935), .A1(ofifoData[204]), .B0(n278), .Z(n2643));
Q_OA21 U5551 ( .A0(n3936), .A1(ofifoData[205]), .B0(n278), .Z(n2640));
Q_OA21 U5552 ( .A0(n3937), .A1(ofifoData[206]), .B0(n278), .Z(n2637));
Q_OA21 U5553 ( .A0(n3938), .A1(ofifoData[207]), .B0(n278), .Z(n2634));
Q_OA21 U5554 ( .A0(n3939), .A1(ofifoData[208]), .B0(n278), .Z(n2631));
Q_OA21 U5555 ( .A0(n3940), .A1(ofifoData[209]), .B0(n278), .Z(n2628));
Q_OA21 U5556 ( .A0(n3941), .A1(ofifoData[210]), .B0(n278), .Z(n2625));
Q_OA21 U5557 ( .A0(n3942), .A1(ofifoData[211]), .B0(n278), .Z(n2622));
Q_OA21 U5558 ( .A0(n3943), .A1(ofifoData[212]), .B0(n278), .Z(n2619));
Q_OA21 U5559 ( .A0(n3944), .A1(ofifoData[213]), .B0(n278), .Z(n2616));
Q_OA21 U5560 ( .A0(n3945), .A1(ofifoData[214]), .B0(n278), .Z(n2613));
Q_OA21 U5561 ( .A0(n3946), .A1(ofifoData[215]), .B0(n278), .Z(n2610));
Q_OA21 U5562 ( .A0(n3947), .A1(ofifoData[216]), .B0(n278), .Z(n2607));
Q_OA21 U5563 ( .A0(n3948), .A1(ofifoData[217]), .B0(n278), .Z(n2604));
Q_OA21 U5564 ( .A0(n3949), .A1(ofifoData[218]), .B0(n278), .Z(n2601));
Q_OA21 U5565 ( .A0(n3950), .A1(ofifoData[219]), .B0(n278), .Z(n2598));
Q_OA21 U5566 ( .A0(n3951), .A1(ofifoData[220]), .B0(n278), .Z(n2595));
Q_OA21 U5567 ( .A0(n3952), .A1(ofifoData[221]), .B0(n278), .Z(n2592));
Q_OA21 U5568 ( .A0(n3953), .A1(ofifoData[222]), .B0(n278), .Z(n2589));
Q_OA21 U5569 ( .A0(n3954), .A1(ofifoData[223]), .B0(n278), .Z(n2586));
Q_OA21 U5570 ( .A0(n3955), .A1(ofifoData[224]), .B0(n278), .Z(n2583));
Q_OA21 U5571 ( .A0(n3956), .A1(ofifoData[225]), .B0(n278), .Z(n2580));
Q_OA21 U5572 ( .A0(n3957), .A1(ofifoData[226]), .B0(n278), .Z(n2577));
Q_OA21 U5573 ( .A0(n3958), .A1(ofifoData[227]), .B0(n278), .Z(n2574));
Q_OA21 U5574 ( .A0(n3959), .A1(ofifoData[228]), .B0(n278), .Z(n2571));
Q_OA21 U5575 ( .A0(n3960), .A1(ofifoData[229]), .B0(n278), .Z(n2568));
Q_OA21 U5576 ( .A0(n3961), .A1(ofifoData[230]), .B0(n278), .Z(n2565));
Q_OA21 U5577 ( .A0(n3962), .A1(ofifoData[231]), .B0(n278), .Z(n2562));
Q_OA21 U5578 ( .A0(n3963), .A1(ofifoData[232]), .B0(n278), .Z(n2559));
Q_OA21 U5579 ( .A0(n3964), .A1(ofifoData[233]), .B0(n278), .Z(n2556));
Q_OA21 U5580 ( .A0(n3965), .A1(ofifoData[234]), .B0(n278), .Z(n2553));
Q_OA21 U5581 ( .A0(n3966), .A1(ofifoData[235]), .B0(n278), .Z(n2550));
Q_OA21 U5582 ( .A0(n3967), .A1(ofifoData[236]), .B0(n278), .Z(n2547));
Q_OA21 U5583 ( .A0(n3968), .A1(ofifoData[237]), .B0(n278), .Z(n2544));
Q_OA21 U5584 ( .A0(n3969), .A1(ofifoData[238]), .B0(n278), .Z(n2541));
Q_OA21 U5585 ( .A0(n3970), .A1(ofifoData[239]), .B0(n278), .Z(n2538));
Q_OA21 U5586 ( .A0(n3971), .A1(ofifoData[240]), .B0(n278), .Z(n2535));
Q_OA21 U5587 ( .A0(n3972), .A1(ofifoData[241]), .B0(n278), .Z(n2532));
Q_OA21 U5588 ( .A0(n3973), .A1(ofifoData[242]), .B0(n278), .Z(n2529));
Q_OA21 U5589 ( .A0(n3974), .A1(ofifoData[243]), .B0(n278), .Z(n2526));
Q_OA21 U5590 ( .A0(n3975), .A1(ofifoData[244]), .B0(n278), .Z(n2523));
Q_OA21 U5591 ( .A0(n3976), .A1(ofifoData[245]), .B0(n278), .Z(n2520));
Q_OA21 U5592 ( .A0(n3977), .A1(ofifoData[246]), .B0(n278), .Z(n2517));
Q_OA21 U5593 ( .A0(n3978), .A1(ofifoData[247]), .B0(n278), .Z(n2514));
Q_OA21 U5594 ( .A0(n3979), .A1(ofifoData[248]), .B0(n278), .Z(n2511));
Q_OA21 U5595 ( .A0(n3980), .A1(ofifoData[249]), .B0(n278), .Z(n2508));
Q_OA21 U5596 ( .A0(n3981), .A1(ofifoData[250]), .B0(n278), .Z(n2505));
Q_OA21 U5597 ( .A0(n3982), .A1(ofifoData[251]), .B0(n278), .Z(n2502));
Q_OA21 U5598 ( .A0(n3983), .A1(ofifoData[252]), .B0(n278), .Z(n2499));
Q_OA21 U5599 ( .A0(n3984), .A1(ofifoData[253]), .B0(n278), .Z(n2496));
Q_OA21 U5600 ( .A0(n3985), .A1(ofifoData[254]), .B0(n278), .Z(n2493));
Q_OA21 U5601 ( .A0(n3986), .A1(ofifoData[255]), .B0(n278), .Z(n2490));
Q_AN02 U5602 ( .A0(oDataEn), .A1(oDataLen[0]), .Z(n3473));
Q_AN02 U5603 ( .A0(oDataEn), .A1(oDataLen[1]), .Z(n3472));
Q_AN02 U5604 ( .A0(oDataEn), .A1(oDataLen[2]), .Z(n3471));
Q_AN02 U5605 ( .A0(oDataEn), .A1(oDataLen[3]), .Z(n3470));
Q_INV U5606 ( .A(numRsts[0]), .Z(n3469));
Q_AD01HF U5607 ( .A0(numRsts[1]), .B0(numRsts[0]), .S(n3468), .CO(n3467));
Q_AD01HF U5608 ( .A0(numRsts[2]), .B0(n3467), .S(n3466), .CO(n3465));
Q_AD01HF U5609 ( .A0(numRsts[3]), .B0(n3465), .S(n3464), .CO(n3463));
Q_AD01HF U5610 ( .A0(numRsts[4]), .B0(n3463), .S(n3462), .CO(n3461));
Q_AD01HF U5611 ( .A0(numRsts[5]), .B0(n3461), .S(n3460), .CO(n3459));
Q_AD01HF U5612 ( .A0(numRsts[6]), .B0(n3459), .S(n3458), .CO(n3457));
Q_AD01HF U5613 ( .A0(numRsts[7]), .B0(n3457), .S(n3456), .CO(n3455));
Q_AD01HF U5614 ( .A0(numRsts[8]), .B0(n3455), .S(n3454), .CO(n3453));
Q_AD01HF U5615 ( .A0(numRsts[9]), .B0(n3453), .S(n3452), .CO(n3451));
Q_AD01HF U5616 ( .A0(numRsts[10]), .B0(n3451), .S(n3450), .CO(n3449));
Q_AD01HF U5617 ( .A0(numRsts[11]), .B0(n3449), .S(n3448), .CO(n3447));
Q_AD01HF U5618 ( .A0(numRsts[12]), .B0(n3447), .S(n3446), .CO(n3445));
Q_AD01HF U5619 ( .A0(numRsts[13]), .B0(n3445), .S(n3444), .CO(n3443));
Q_AD01HF U5620 ( .A0(numRsts[14]), .B0(n3443), .S(n3442), .CO(n3441));
Q_AD01HF U5621 ( .A0(numRsts[15]), .B0(n3441), .S(n3440), .CO(n3439));
Q_AD01HF U5622 ( .A0(numRsts[16]), .B0(n3439), .S(n3438), .CO(n3437));
Q_AD01HF U5623 ( .A0(numRsts[17]), .B0(n3437), .S(n3436), .CO(n3435));
Q_AD01HF U5624 ( .A0(numRsts[18]), .B0(n3435), .S(n3434), .CO(n3433));
Q_AD01HF U5625 ( .A0(numRsts[19]), .B0(n3433), .S(n3432), .CO(n3431));
Q_AD01HF U5626 ( .A0(numRsts[20]), .B0(n3431), .S(n3430), .CO(n3429));
Q_AD01HF U5627 ( .A0(numRsts[21]), .B0(n3429), .S(n3428), .CO(n3427));
Q_AD01HF U5628 ( .A0(numRsts[22]), .B0(n3427), .S(n3426), .CO(n3425));
Q_AD01HF U5629 ( .A0(numRsts[23]), .B0(n3425), .S(n3424), .CO(n3423));
Q_AD01HF U5630 ( .A0(numRsts[24]), .B0(n3423), .S(n3422), .CO(n3421));
Q_AD01HF U5631 ( .A0(numRsts[25]), .B0(n3421), .S(n3420), .CO(n3419));
Q_AD01HF U5632 ( .A0(numRsts[26]), .B0(n3419), .S(n3418), .CO(n3417));
Q_AD01HF U5633 ( .A0(numRsts[27]), .B0(n3417), .S(n3416), .CO(n3415));
Q_AD01HF U5634 ( .A0(numRsts[28]), .B0(n3415), .S(n3414), .CO(n3413));
Q_AD01HF U5635 ( .A0(numRsts[29]), .B0(n3413), .S(n3412), .CO(n3411));
Q_AD01HF U5636 ( .A0(numRsts[30]), .B0(n3411), .S(n3410), .CO(n3409));
Q_XOR2 U5637 ( .A0(numRsts[31]), .A1(n3409), .Z(n3408));
Q_AD01HF U5638 ( .A0(ofifoWptr[1]), .B0(ofifoWptr[0]), .S(n3407), .CO(n3406));
Q_AD01HF U5639 ( .A0(ofifoWptr[2]), .B0(n3406), .S(n3405), .CO(n3404));
Q_AD01HF U5640 ( .A0(ofifoWptr[3]), .B0(n3404), .S(n3403), .CO(n3402));
Q_AD01HF U5641 ( .A0(ofifoWptr[4]), .B0(n3402), .S(n3401), .CO(n3400));
Q_AD01HF U5642 ( .A0(ofifoWptr[5]), .B0(n3400), .S(n3399), .CO(n3398));
Q_AD01HF U5643 ( .A0(ofifoWptr[6]), .B0(n3398), .S(n3397), .CO(n3396));
Q_AD01HF U5644 ( .A0(ofifoWptr[7]), .B0(n3396), .S(n3395), .CO(n3394));
Q_AD01HF U5645 ( .A0(ofifoWptr[8]), .B0(n3394), .S(n3393), .CO(n3392));
Q_AD01HF U5646 ( .A0(ofifoWptr[9]), .B0(n3392), .S(n3391), .CO(n3390));
Q_AD01HF U5647 ( .A0(ofifoWptr[10]), .B0(n3390), .S(n3389), .CO(n3388));
Q_AD01HF U5648 ( .A0(ofifoWptr[11]), .B0(n3388), .S(n3387), .CO(n3386));
Q_AD01HF U5649 ( .A0(ofifoWptr[12]), .B0(n3386), .S(n3385), .CO(n3384));
Q_AD01HF U5650 ( .A0(ofifoWptr[13]), .B0(n3384), .S(n3383), .CO(n3382));
Q_AD01HF U5651 ( .A0(ofifoWptr[14]), .B0(n3382), .S(n3381), .CO(n3380));
Q_INV U5652 ( .A(ofifoWptr[1]), .Z(n3379));
Q_AD01HF U5653 ( .A0(ofifoWptr[2]), .B0(ofifoWptr[1]), .S(n3378), .CO(n3377));
Q_AD01HF U5654 ( .A0(ofifoWptr[3]), .B0(n3377), .S(n3376), .CO(n3375));
Q_AD01HF U5655 ( .A0(ofifoWptr[4]), .B0(n3375), .S(n3374), .CO(n3373));
Q_AD01HF U5656 ( .A0(ofifoWptr[5]), .B0(n3373), .S(n3372), .CO(n3371));
Q_AD01HF U5657 ( .A0(ofifoWptr[6]), .B0(n3371), .S(n3370), .CO(n3369));
Q_AD01HF U5658 ( .A0(ofifoWptr[7]), .B0(n3369), .S(n3368), .CO(n3367));
Q_AD01HF U5659 ( .A0(ofifoWptr[8]), .B0(n3367), .S(n3366), .CO(n3365));
Q_AD01HF U5660 ( .A0(ofifoWptr[9]), .B0(n3365), .S(n3364), .CO(n3363));
Q_AD01HF U5661 ( .A0(ofifoWptr[10]), .B0(n3363), .S(n3362), .CO(n3361));
Q_AD01HF U5662 ( .A0(ofifoWptr[11]), .B0(n3361), .S(n3360), .CO(n3359));
Q_AD01HF U5663 ( .A0(ofifoWptr[12]), .B0(n3359), .S(n3358), .CO(n3357));
Q_AD01HF U5664 ( .A0(ofifoWptr[13]), .B0(n3357), .S(n3356), .CO(n3355));
Q_AD01HF U5665 ( .A0(ofifoWptr[14]), .B0(n3355), .S(n3354), .CO(n3353));
Q_AD01HF U5666 ( .A0(oFill[0]), .B0(n3473), .S(n3352), .CO(n3351));
Q_AD01 U5667 ( .CI(n3472), .A0(oFill[1]), .B0(n3351), .S(n3350), .CO(n3349));
Q_AD01HF U5668 ( .A0(n3471), .B0(n3349), .S(n3348), .CO(n3347));
Q_AD01HF U5669 ( .A0(ofifoWptr[0]), .B0(n3348), .S(n3345), .CO(n3344));
Q_AD01 U5670 ( .CI(n3346), .A0(ofifoWptr[1]), .B0(n3344), .S(n3343), .CO(n3342));
Q_AD01HF U5671 ( .A0(ofifoWptr[2]), .B0(n3342), .S(n3341), .CO(n3340));
Q_AD01HF U5672 ( .A0(ofifoWptr[3]), .B0(n3340), .S(n3339), .CO(n3338));
Q_AD01HF U5673 ( .A0(ofifoWptr[4]), .B0(n3338), .S(n3337), .CO(n3336));
Q_AD01HF U5674 ( .A0(ofifoWptr[5]), .B0(n3336), .S(n3335), .CO(n3334));
Q_AD01HF U5675 ( .A0(ofifoWptr[6]), .B0(n3334), .S(n3333), .CO(n3332));
Q_AD01HF U5676 ( .A0(ofifoWptr[7]), .B0(n3332), .S(n3331), .CO(n3330));
Q_AD01HF U5677 ( .A0(ofifoWptr[8]), .B0(n3330), .S(n3329), .CO(n3328));
Q_AD01HF U5678 ( .A0(ofifoWptr[9]), .B0(n3328), .S(n3327), .CO(n3326));
Q_AD01HF U5679 ( .A0(ofifoWptr[10]), .B0(n3326), .S(n3325), .CO(n3324));
Q_AD01HF U5680 ( .A0(ofifoWptr[11]), .B0(n3324), .S(n3323), .CO(n3322));
Q_AD01HF U5681 ( .A0(ofifoWptr[12]), .B0(n3322), .S(n3321), .CO(n3320));
Q_AD01HF U5682 ( .A0(ofifoWptr[13]), .B0(n3320), .S(n3319), .CO(n3318));
Q_XOR2 U5683 ( .A0(ofifoWptr[14]), .A1(n3318), .Z(n3317));
Q_OR02 U5684 ( .A0(n301), .A1(n3345), .Z(n3316));
Q_AN02 U5685 ( .A0(n280), .A1(n3343), .Z(n3315));
Q_AN02 U5686 ( .A0(n280), .A1(n3341), .Z(n3314));
Q_AN02 U5687 ( .A0(n280), .A1(n3339), .Z(n3313));
Q_AN02 U5688 ( .A0(n280), .A1(n3337), .Z(n3312));
Q_AN02 U5689 ( .A0(n280), .A1(n3335), .Z(n3311));
Q_AN02 U5690 ( .A0(n280), .A1(n3333), .Z(n3310));
Q_AN02 U5691 ( .A0(n280), .A1(n3331), .Z(n3309));
Q_AN02 U5692 ( .A0(n280), .A1(n3329), .Z(n3308));
Q_AN02 U5693 ( .A0(n280), .A1(n3327), .Z(n3307));
Q_AN02 U5694 ( .A0(n280), .A1(n3325), .Z(n3306));
Q_AN02 U5695 ( .A0(n280), .A1(n3323), .Z(n3305));
Q_AN02 U5696 ( .A0(n280), .A1(n3321), .Z(n3304));
Q_AN02 U5697 ( .A0(n280), .A1(n3319), .Z(n3303));
Q_AN02 U5698 ( .A0(n280), .A1(n3317), .Z(n3302));
Q_OR02 U5699 ( .A0(xc_top.GFReset), .A1(n3379), .Z(n3301));
Q_AN02 U5700 ( .A0(n279), .A1(n3378), .Z(n3300));
Q_AN02 U5701 ( .A0(n279), .A1(n3376), .Z(n3299));
Q_AN02 U5702 ( .A0(n279), .A1(n3374), .Z(n3298));
Q_AN02 U5703 ( .A0(n279), .A1(n3372), .Z(n3297));
Q_AN02 U5704 ( .A0(n279), .A1(n3370), .Z(n3296));
Q_AN02 U5705 ( .A0(n279), .A1(n3368), .Z(n3295));
Q_AN02 U5706 ( .A0(n279), .A1(n3366), .Z(n3294));
Q_AN02 U5707 ( .A0(n279), .A1(n3364), .Z(n3293));
Q_AN02 U5708 ( .A0(n279), .A1(n3362), .Z(n3292));
Q_AN02 U5709 ( .A0(n279), .A1(n3360), .Z(n3291));
Q_AN02 U5710 ( .A0(n279), .A1(n3358), .Z(n3290));
Q_AN02 U5711 ( .A0(n279), .A1(n3356), .Z(n3289));
Q_AN02 U5712 ( .A0(n279), .A1(n3354), .Z(n3288));
Q_AN02 U5713 ( .A0(n279), .A1(n3353), .Z(n3287));
Q_OR02 U5714 ( .A0(xc_top.GFReset), .A1(n3407), .Z(n3286));
Q_AN02 U5715 ( .A0(n279), .A1(n3405), .Z(n3285));
Q_AN02 U5716 ( .A0(n279), .A1(n3403), .Z(n3284));
Q_AN02 U5717 ( .A0(n279), .A1(n3401), .Z(n3283));
Q_AN02 U5718 ( .A0(n279), .A1(n3399), .Z(n3282));
Q_AN02 U5719 ( .A0(n279), .A1(n3397), .Z(n3281));
Q_AN02 U5720 ( .A0(n279), .A1(n3395), .Z(n3280));
Q_AN02 U5721 ( .A0(n279), .A1(n3393), .Z(n3279));
Q_AN02 U5722 ( .A0(n279), .A1(n3391), .Z(n3278));
Q_AN02 U5723 ( .A0(n279), .A1(n3389), .Z(n3277));
Q_AN02 U5724 ( .A0(n279), .A1(n3387), .Z(n3276));
Q_AN02 U5725 ( .A0(n279), .A1(n3385), .Z(n3275));
Q_AN02 U5726 ( .A0(n279), .A1(n3383), .Z(n3274));
Q_AN02 U5727 ( .A0(n279), .A1(n3381), .Z(n3273));
Q_AN02 U5728 ( .A0(n279), .A1(n3380), .Z(n3272));
Q_OR02 U5729 ( .A0(xc_top.GFReset), .A1(ofifoWptr[0]), .Z(n3271));
Q_AN02 U5730 ( .A0(n279), .A1(ofifoWptr[1]), .Z(n3270));
Q_AN02 U5731 ( .A0(n279), .A1(ofifoWptr[2]), .Z(n3269));
Q_AN02 U5732 ( .A0(n279), .A1(ofifoWptr[3]), .Z(n3268));
Q_AN02 U5733 ( .A0(n279), .A1(ofifoWptr[4]), .Z(n3267));
Q_AN02 U5734 ( .A0(n279), .A1(ofifoWptr[5]), .Z(n3266));
Q_AN02 U5735 ( .A0(n279), .A1(ofifoWptr[6]), .Z(n3265));
Q_AN02 U5736 ( .A0(n279), .A1(ofifoWptr[7]), .Z(n3264));
Q_AN02 U5737 ( .A0(n279), .A1(ofifoWptr[8]), .Z(n3263));
Q_AN02 U5738 ( .A0(n279), .A1(ofifoWptr[9]), .Z(n3262));
Q_AN02 U5739 ( .A0(n279), .A1(ofifoWptr[10]), .Z(n3261));
Q_AN02 U5740 ( .A0(n279), .A1(ofifoWptr[11]), .Z(n3260));
Q_AN02 U5741 ( .A0(n279), .A1(ofifoWptr[12]), .Z(n3259));
Q_AN02 U5742 ( .A0(n279), .A1(ofifoWptr[13]), .Z(n3258));
Q_AN02 U5743 ( .A0(n279), .A1(ofifoWptr[14]), .Z(n3257));
Q_MX02 U5744 ( .S(n278), .A0(ofifoData[256]), .A1(ofifoData[512]), .Z(n3729));
Q_MX03 U5745 ( .S0(n277), .S1(n276), .A0(n3255), .A1(n3256), .A2(n3730), .Z(n3254));
Q_MX02 U5746 ( .S(n278), .A0(ofifoData[257]), .A1(ofifoData[513]), .Z(n3728));
Q_MX03 U5747 ( .S0(n277), .S1(n276), .A0(n3252), .A1(n3253), .A2(n3731), .Z(n3251));
Q_MX02 U5748 ( .S(n278), .A0(ofifoData[258]), .A1(ofifoData[514]), .Z(n3727));
Q_MX03 U5749 ( .S0(n277), .S1(n276), .A0(n3249), .A1(n3250), .A2(n3732), .Z(n3248));
Q_MX02 U5750 ( .S(n278), .A0(ofifoData[259]), .A1(ofifoData[515]), .Z(n3726));
Q_MX03 U5751 ( .S0(n277), .S1(n276), .A0(n3246), .A1(n3247), .A2(n3733), .Z(n3245));
Q_MX02 U5752 ( .S(n278), .A0(ofifoData[260]), .A1(ofifoData[516]), .Z(n3725));
Q_MX03 U5753 ( .S0(n277), .S1(n276), .A0(n3243), .A1(n3244), .A2(n3734), .Z(n3242));
Q_MX02 U5754 ( .S(n278), .A0(ofifoData[261]), .A1(ofifoData[517]), .Z(n3724));
Q_MX03 U5755 ( .S0(n277), .S1(n276), .A0(n3240), .A1(n3241), .A2(n3735), .Z(n3239));
Q_MX02 U5756 ( .S(n278), .A0(ofifoData[262]), .A1(ofifoData[518]), .Z(n3723));
Q_MX03 U5757 ( .S0(n277), .S1(n276), .A0(n3237), .A1(n3238), .A2(n3736), .Z(n3236));
Q_MX02 U5758 ( .S(n278), .A0(ofifoData[263]), .A1(ofifoData[519]), .Z(n3722));
Q_MX03 U5759 ( .S0(n277), .S1(n276), .A0(n3234), .A1(n3235), .A2(n3737), .Z(n3233));
Q_MX02 U5760 ( .S(n278), .A0(ofifoData[264]), .A1(ofifoData[520]), .Z(n3721));
Q_MX03 U5761 ( .S0(n277), .S1(n276), .A0(n3231), .A1(n3232), .A2(n3738), .Z(n3230));
Q_MX02 U5762 ( .S(n278), .A0(ofifoData[265]), .A1(ofifoData[521]), .Z(n3720));
Q_MX03 U5763 ( .S0(n277), .S1(n276), .A0(n3228), .A1(n3229), .A2(n3739), .Z(n3227));
Q_MX02 U5764 ( .S(n278), .A0(ofifoData[266]), .A1(ofifoData[522]), .Z(n3719));
Q_MX03 U5765 ( .S0(n277), .S1(n276), .A0(n3225), .A1(n3226), .A2(n3740), .Z(n3224));
Q_MX02 U5766 ( .S(n278), .A0(ofifoData[267]), .A1(ofifoData[523]), .Z(n3718));
Q_MX03 U5767 ( .S0(n277), .S1(n276), .A0(n3222), .A1(n3223), .A2(n3741), .Z(n3221));
Q_MX02 U5768 ( .S(n278), .A0(ofifoData[268]), .A1(ofifoData[524]), .Z(n3717));
Q_MX03 U5769 ( .S0(n277), .S1(n276), .A0(n3219), .A1(n3220), .A2(n3742), .Z(n3218));
Q_MX02 U5770 ( .S(n278), .A0(ofifoData[269]), .A1(ofifoData[525]), .Z(n3716));
Q_MX03 U5771 ( .S0(n277), .S1(n276), .A0(n3216), .A1(n3217), .A2(n3743), .Z(n3215));
Q_MX02 U5772 ( .S(n278), .A0(ofifoData[270]), .A1(ofifoData[526]), .Z(n3715));
Q_MX03 U5773 ( .S0(n277), .S1(n276), .A0(n3213), .A1(n3214), .A2(n3744), .Z(n3212));
Q_MX02 U5774 ( .S(n278), .A0(ofifoData[271]), .A1(ofifoData[527]), .Z(n3714));
Q_MX03 U5775 ( .S0(n277), .S1(n276), .A0(n3210), .A1(n3211), .A2(n3745), .Z(n3209));
Q_MX02 U5776 ( .S(n278), .A0(ofifoData[272]), .A1(ofifoData[528]), .Z(n3713));
Q_MX03 U5777 ( .S0(n277), .S1(n276), .A0(n3207), .A1(n3208), .A2(n3746), .Z(n3206));
Q_MX02 U5778 ( .S(n278), .A0(ofifoData[273]), .A1(ofifoData[529]), .Z(n3712));
Q_MX03 U5779 ( .S0(n277), .S1(n276), .A0(n3204), .A1(n3205), .A2(n3747), .Z(n3203));
Q_MX02 U5780 ( .S(n278), .A0(ofifoData[274]), .A1(ofifoData[530]), .Z(n3711));
Q_MX03 U5781 ( .S0(n277), .S1(n276), .A0(n3201), .A1(n3202), .A2(n3748), .Z(n3200));
Q_MX02 U5782 ( .S(n278), .A0(ofifoData[275]), .A1(ofifoData[531]), .Z(n3710));
Q_MX03 U5783 ( .S0(n277), .S1(n276), .A0(n3198), .A1(n3199), .A2(n3749), .Z(n3197));
Q_MX02 U5784 ( .S(n278), .A0(ofifoData[276]), .A1(ofifoData[532]), .Z(n3709));
Q_MX03 U5785 ( .S0(n277), .S1(n276), .A0(n3195), .A1(n3196), .A2(n3750), .Z(n3194));
Q_MX02 U5786 ( .S(n278), .A0(ofifoData[277]), .A1(ofifoData[533]), .Z(n3708));
Q_MX03 U5787 ( .S0(n277), .S1(n276), .A0(n3192), .A1(n3193), .A2(n3751), .Z(n3191));
Q_MX02 U5788 ( .S(n278), .A0(ofifoData[278]), .A1(ofifoData[534]), .Z(n3707));
Q_MX03 U5789 ( .S0(n277), .S1(n276), .A0(n3189), .A1(n3190), .A2(n3752), .Z(n3188));
Q_MX02 U5790 ( .S(n278), .A0(ofifoData[279]), .A1(ofifoData[535]), .Z(n3706));
Q_MX03 U5791 ( .S0(n277), .S1(n276), .A0(n3186), .A1(n3187), .A2(n3753), .Z(n3185));
Q_MX02 U5792 ( .S(n278), .A0(ofifoData[280]), .A1(ofifoData[536]), .Z(n3705));
Q_MX03 U5793 ( .S0(n277), .S1(n276), .A0(n3183), .A1(n3184), .A2(n3754), .Z(n3182));
Q_MX02 U5794 ( .S(n278), .A0(ofifoData[281]), .A1(ofifoData[537]), .Z(n3704));
Q_MX03 U5795 ( .S0(n277), .S1(n276), .A0(n3180), .A1(n3181), .A2(n3755), .Z(n3179));
Q_MX02 U5796 ( .S(n278), .A0(ofifoData[282]), .A1(ofifoData[538]), .Z(n3703));
Q_MX03 U5797 ( .S0(n277), .S1(n276), .A0(n3177), .A1(n3178), .A2(n3756), .Z(n3176));
Q_MX02 U5798 ( .S(n278), .A0(ofifoData[283]), .A1(ofifoData[539]), .Z(n3702));
Q_MX03 U5799 ( .S0(n277), .S1(n276), .A0(n3174), .A1(n3175), .A2(n3757), .Z(n3173));
Q_MX02 U5800 ( .S(n278), .A0(ofifoData[284]), .A1(ofifoData[540]), .Z(n3701));
Q_MX03 U5801 ( .S0(n277), .S1(n276), .A0(n3171), .A1(n3172), .A2(n3758), .Z(n3170));
Q_MX02 U5802 ( .S(n278), .A0(ofifoData[285]), .A1(ofifoData[541]), .Z(n3700));
Q_MX03 U5803 ( .S0(n277), .S1(n276), .A0(n3168), .A1(n3169), .A2(n3759), .Z(n3167));
Q_MX02 U5804 ( .S(n278), .A0(ofifoData[286]), .A1(ofifoData[542]), .Z(n3699));
Q_MX03 U5805 ( .S0(n277), .S1(n276), .A0(n3165), .A1(n3166), .A2(n3760), .Z(n3164));
Q_MX02 U5806 ( .S(n278), .A0(ofifoData[287]), .A1(ofifoData[543]), .Z(n3698));
Q_MX03 U5807 ( .S0(n277), .S1(n276), .A0(n3162), .A1(n3163), .A2(n3761), .Z(n3161));
Q_MX02 U5808 ( .S(n278), .A0(ofifoData[288]), .A1(ofifoData[544]), .Z(n3697));
Q_MX03 U5809 ( .S0(n277), .S1(n276), .A0(n3159), .A1(n3160), .A2(n3762), .Z(n3158));
Q_MX02 U5810 ( .S(n278), .A0(ofifoData[289]), .A1(ofifoData[545]), .Z(n3696));
Q_MX03 U5811 ( .S0(n277), .S1(n276), .A0(n3156), .A1(n3157), .A2(n3763), .Z(n3155));
Q_MX02 U5812 ( .S(n278), .A0(ofifoData[290]), .A1(ofifoData[546]), .Z(n3695));
Q_MX03 U5813 ( .S0(n277), .S1(n276), .A0(n3153), .A1(n3154), .A2(n3764), .Z(n3152));
Q_MX02 U5814 ( .S(n278), .A0(ofifoData[291]), .A1(ofifoData[547]), .Z(n3694));
Q_MX03 U5815 ( .S0(n277), .S1(n276), .A0(n3150), .A1(n3151), .A2(n3765), .Z(n3149));
Q_MX02 U5816 ( .S(n278), .A0(ofifoData[292]), .A1(ofifoData[548]), .Z(n3693));
Q_MX03 U5817 ( .S0(n277), .S1(n276), .A0(n3147), .A1(n3148), .A2(n3766), .Z(n3146));
Q_MX02 U5818 ( .S(n278), .A0(ofifoData[293]), .A1(ofifoData[549]), .Z(n3692));
Q_MX03 U5819 ( .S0(n277), .S1(n276), .A0(n3144), .A1(n3145), .A2(n3767), .Z(n3143));
Q_MX02 U5820 ( .S(n278), .A0(ofifoData[294]), .A1(ofifoData[550]), .Z(n3691));
Q_MX03 U5821 ( .S0(n277), .S1(n276), .A0(n3141), .A1(n3142), .A2(n3768), .Z(n3140));
Q_MX02 U5822 ( .S(n278), .A0(ofifoData[295]), .A1(ofifoData[551]), .Z(n3690));
Q_MX03 U5823 ( .S0(n277), .S1(n276), .A0(n3138), .A1(n3139), .A2(n3769), .Z(n3137));
Q_MX02 U5824 ( .S(n278), .A0(ofifoData[296]), .A1(ofifoData[552]), .Z(n3689));
Q_MX03 U5825 ( .S0(n277), .S1(n276), .A0(n3135), .A1(n3136), .A2(n3770), .Z(n3134));
Q_MX02 U5826 ( .S(n278), .A0(ofifoData[297]), .A1(ofifoData[553]), .Z(n3688));
Q_MX03 U5827 ( .S0(n277), .S1(n276), .A0(n3132), .A1(n3133), .A2(n3771), .Z(n3131));
Q_MX02 U5828 ( .S(n278), .A0(ofifoData[298]), .A1(ofifoData[554]), .Z(n3687));
Q_MX03 U5829 ( .S0(n277), .S1(n276), .A0(n3129), .A1(n3130), .A2(n3772), .Z(n3128));
Q_MX02 U5830 ( .S(n278), .A0(ofifoData[299]), .A1(ofifoData[555]), .Z(n3686));
Q_MX03 U5831 ( .S0(n277), .S1(n276), .A0(n3126), .A1(n3127), .A2(n3773), .Z(n3125));
Q_MX02 U5832 ( .S(n278), .A0(ofifoData[300]), .A1(ofifoData[556]), .Z(n3685));
Q_MX03 U5833 ( .S0(n277), .S1(n276), .A0(n3123), .A1(n3124), .A2(n3774), .Z(n3122));
Q_MX02 U5834 ( .S(n278), .A0(ofifoData[301]), .A1(ofifoData[557]), .Z(n3684));
Q_MX03 U5835 ( .S0(n277), .S1(n276), .A0(n3120), .A1(n3121), .A2(n3775), .Z(n3119));
Q_MX02 U5836 ( .S(n278), .A0(ofifoData[302]), .A1(ofifoData[558]), .Z(n3683));
Q_MX03 U5837 ( .S0(n277), .S1(n276), .A0(n3117), .A1(n3118), .A2(n3776), .Z(n3116));
Q_MX02 U5838 ( .S(n278), .A0(ofifoData[303]), .A1(ofifoData[559]), .Z(n3682));
Q_MX03 U5839 ( .S0(n277), .S1(n276), .A0(n3114), .A1(n3115), .A2(n3777), .Z(n3113));
Q_MX02 U5840 ( .S(n278), .A0(ofifoData[304]), .A1(ofifoData[560]), .Z(n3681));
Q_MX03 U5841 ( .S0(n277), .S1(n276), .A0(n3111), .A1(n3112), .A2(n3778), .Z(n3110));
Q_MX02 U5842 ( .S(n278), .A0(ofifoData[305]), .A1(ofifoData[561]), .Z(n3680));
Q_MX03 U5843 ( .S0(n277), .S1(n276), .A0(n3108), .A1(n3109), .A2(n3779), .Z(n3107));
Q_MX02 U5844 ( .S(n278), .A0(ofifoData[306]), .A1(ofifoData[562]), .Z(n3679));
Q_MX03 U5845 ( .S0(n277), .S1(n276), .A0(n3105), .A1(n3106), .A2(n3780), .Z(n3104));
Q_MX02 U5846 ( .S(n278), .A0(ofifoData[307]), .A1(ofifoData[563]), .Z(n3678));
Q_MX03 U5847 ( .S0(n277), .S1(n276), .A0(n3102), .A1(n3103), .A2(n3781), .Z(n3101));
Q_MX02 U5848 ( .S(n278), .A0(ofifoData[308]), .A1(ofifoData[564]), .Z(n3677));
Q_MX03 U5849 ( .S0(n277), .S1(n276), .A0(n3099), .A1(n3100), .A2(n3782), .Z(n3098));
Q_MX02 U5850 ( .S(n278), .A0(ofifoData[309]), .A1(ofifoData[565]), .Z(n3676));
Q_MX03 U5851 ( .S0(n277), .S1(n276), .A0(n3096), .A1(n3097), .A2(n3783), .Z(n3095));
Q_MX02 U5852 ( .S(n278), .A0(ofifoData[310]), .A1(ofifoData[566]), .Z(n3675));
Q_MX03 U5853 ( .S0(n277), .S1(n276), .A0(n3093), .A1(n3094), .A2(n3784), .Z(n3092));
Q_MX02 U5854 ( .S(n278), .A0(ofifoData[311]), .A1(ofifoData[567]), .Z(n3674));
Q_MX03 U5855 ( .S0(n277), .S1(n276), .A0(n3090), .A1(n3091), .A2(n3785), .Z(n3089));
Q_MX02 U5856 ( .S(n278), .A0(ofifoData[312]), .A1(ofifoData[568]), .Z(n3673));
Q_MX03 U5857 ( .S0(n277), .S1(n276), .A0(n3087), .A1(n3088), .A2(n3786), .Z(n3086));
Q_MX02 U5858 ( .S(n278), .A0(ofifoData[313]), .A1(ofifoData[569]), .Z(n3672));
Q_MX03 U5859 ( .S0(n277), .S1(n276), .A0(n3084), .A1(n3085), .A2(n3787), .Z(n3083));
Q_MX02 U5860 ( .S(n278), .A0(ofifoData[314]), .A1(ofifoData[570]), .Z(n3671));
Q_MX03 U5861 ( .S0(n277), .S1(n276), .A0(n3081), .A1(n3082), .A2(n3788), .Z(n3080));
Q_MX02 U5862 ( .S(n278), .A0(ofifoData[315]), .A1(ofifoData[571]), .Z(n3670));
Q_MX03 U5863 ( .S0(n277), .S1(n276), .A0(n3078), .A1(n3079), .A2(n3789), .Z(n3077));
Q_MX02 U5864 ( .S(n278), .A0(ofifoData[316]), .A1(ofifoData[572]), .Z(n3669));
Q_MX03 U5865 ( .S0(n277), .S1(n276), .A0(n3075), .A1(n3076), .A2(n3790), .Z(n3074));
Q_MX02 U5866 ( .S(n278), .A0(ofifoData[317]), .A1(ofifoData[573]), .Z(n3668));
Q_MX03 U5867 ( .S0(n277), .S1(n276), .A0(n3072), .A1(n3073), .A2(n3791), .Z(n3071));
Q_MX02 U5868 ( .S(n278), .A0(ofifoData[318]), .A1(ofifoData[574]), .Z(n3667));
Q_MX03 U5869 ( .S0(n277), .S1(n276), .A0(n3069), .A1(n3070), .A2(n3792), .Z(n3068));
Q_MX02 U5870 ( .S(n278), .A0(ofifoData[319]), .A1(ofifoData[575]), .Z(n3666));
Q_MX03 U5871 ( .S0(n277), .S1(n276), .A0(n3066), .A1(n3067), .A2(n3793), .Z(n3065));
Q_MX02 U5872 ( .S(n278), .A0(ofifoData[320]), .A1(ofifoData[576]), .Z(n3665));
Q_MX03 U5873 ( .S0(n277), .S1(n276), .A0(n3063), .A1(n3064), .A2(n3794), .Z(n3062));
Q_MX02 U5874 ( .S(n278), .A0(ofifoData[321]), .A1(ofifoData[577]), .Z(n3664));
Q_MX03 U5875 ( .S0(n277), .S1(n276), .A0(n3060), .A1(n3061), .A2(n3795), .Z(n3059));
Q_MX02 U5876 ( .S(n278), .A0(ofifoData[322]), .A1(ofifoData[578]), .Z(n3663));
Q_MX03 U5877 ( .S0(n277), .S1(n276), .A0(n3057), .A1(n3058), .A2(n3796), .Z(n3056));
Q_MX02 U5878 ( .S(n278), .A0(ofifoData[323]), .A1(ofifoData[579]), .Z(n3662));
Q_MX03 U5879 ( .S0(n277), .S1(n276), .A0(n3054), .A1(n3055), .A2(n3797), .Z(n3053));
Q_MX02 U5880 ( .S(n278), .A0(ofifoData[324]), .A1(ofifoData[580]), .Z(n3661));
Q_MX03 U5881 ( .S0(n277), .S1(n276), .A0(n3051), .A1(n3052), .A2(n3798), .Z(n3050));
Q_MX02 U5882 ( .S(n278), .A0(ofifoData[325]), .A1(ofifoData[581]), .Z(n3660));
Q_MX03 U5883 ( .S0(n277), .S1(n276), .A0(n3048), .A1(n3049), .A2(n3799), .Z(n3047));
Q_MX02 U5884 ( .S(n278), .A0(ofifoData[326]), .A1(ofifoData[582]), .Z(n3659));
Q_MX03 U5885 ( .S0(n277), .S1(n276), .A0(n3045), .A1(n3046), .A2(n3800), .Z(n3044));
Q_MX02 U5886 ( .S(n278), .A0(ofifoData[327]), .A1(ofifoData[583]), .Z(n3658));
Q_MX03 U5887 ( .S0(n277), .S1(n276), .A0(n3042), .A1(n3043), .A2(n3801), .Z(n3041));
Q_MX02 U5888 ( .S(n278), .A0(ofifoData[328]), .A1(ofifoData[584]), .Z(n3657));
Q_MX03 U5889 ( .S0(n277), .S1(n276), .A0(n3039), .A1(n3040), .A2(n3802), .Z(n3038));
Q_MX02 U5890 ( .S(n278), .A0(ofifoData[329]), .A1(ofifoData[585]), .Z(n3656));
Q_MX03 U5891 ( .S0(n277), .S1(n276), .A0(n3036), .A1(n3037), .A2(n3803), .Z(n3035));
Q_MX02 U5892 ( .S(n278), .A0(ofifoData[330]), .A1(ofifoData[586]), .Z(n3655));
Q_MX03 U5893 ( .S0(n277), .S1(n276), .A0(n3033), .A1(n3034), .A2(n3804), .Z(n3032));
Q_MX02 U5894 ( .S(n278), .A0(ofifoData[331]), .A1(ofifoData[587]), .Z(n3654));
Q_MX03 U5895 ( .S0(n277), .S1(n276), .A0(n3030), .A1(n3031), .A2(n3805), .Z(n3029));
Q_MX02 U5896 ( .S(n278), .A0(ofifoData[332]), .A1(ofifoData[588]), .Z(n3653));
Q_MX03 U5897 ( .S0(n277), .S1(n276), .A0(n3027), .A1(n3028), .A2(n3806), .Z(n3026));
Q_MX02 U5898 ( .S(n278), .A0(ofifoData[333]), .A1(ofifoData[589]), .Z(n3652));
Q_MX03 U5899 ( .S0(n277), .S1(n276), .A0(n3024), .A1(n3025), .A2(n3807), .Z(n3023));
Q_MX02 U5900 ( .S(n278), .A0(ofifoData[334]), .A1(ofifoData[590]), .Z(n3651));
Q_MX03 U5901 ( .S0(n277), .S1(n276), .A0(n3021), .A1(n3022), .A2(n3808), .Z(n3020));
Q_MX02 U5902 ( .S(n278), .A0(ofifoData[335]), .A1(ofifoData[591]), .Z(n3650));
Q_MX03 U5903 ( .S0(n277), .S1(n276), .A0(n3018), .A1(n3019), .A2(n3809), .Z(n3017));
Q_MX02 U5904 ( .S(n278), .A0(ofifoData[336]), .A1(ofifoData[592]), .Z(n3649));
Q_MX03 U5905 ( .S0(n277), .S1(n276), .A0(n3015), .A1(n3016), .A2(n3810), .Z(n3014));
Q_MX02 U5906 ( .S(n278), .A0(ofifoData[337]), .A1(ofifoData[593]), .Z(n3648));
Q_MX03 U5907 ( .S0(n277), .S1(n276), .A0(n3012), .A1(n3013), .A2(n3811), .Z(n3011));
Q_MX02 U5908 ( .S(n278), .A0(ofifoData[338]), .A1(ofifoData[594]), .Z(n3647));
Q_MX03 U5909 ( .S0(n277), .S1(n276), .A0(n3009), .A1(n3010), .A2(n3812), .Z(n3008));
Q_MX02 U5910 ( .S(n278), .A0(ofifoData[339]), .A1(ofifoData[595]), .Z(n3646));
Q_MX03 U5911 ( .S0(n277), .S1(n276), .A0(n3006), .A1(n3007), .A2(n3813), .Z(n3005));
Q_MX02 U5912 ( .S(n278), .A0(ofifoData[340]), .A1(ofifoData[596]), .Z(n3645));
Q_MX03 U5913 ( .S0(n277), .S1(n276), .A0(n3003), .A1(n3004), .A2(n3814), .Z(n3002));
Q_MX02 U5914 ( .S(n278), .A0(ofifoData[341]), .A1(ofifoData[597]), .Z(n3644));
Q_MX03 U5915 ( .S0(n277), .S1(n276), .A0(n3000), .A1(n3001), .A2(n3815), .Z(n2999));
Q_MX02 U5916 ( .S(n278), .A0(ofifoData[342]), .A1(ofifoData[598]), .Z(n3643));
Q_MX03 U5917 ( .S0(n277), .S1(n276), .A0(n2997), .A1(n2998), .A2(n3816), .Z(n2996));
Q_MX02 U5918 ( .S(n278), .A0(ofifoData[343]), .A1(ofifoData[599]), .Z(n3642));
Q_MX03 U5919 ( .S0(n277), .S1(n276), .A0(n2994), .A1(n2995), .A2(n3817), .Z(n2993));
Q_MX02 U5920 ( .S(n278), .A0(ofifoData[344]), .A1(ofifoData[600]), .Z(n3641));
Q_MX03 U5921 ( .S0(n277), .S1(n276), .A0(n2991), .A1(n2992), .A2(n3818), .Z(n2990));
Q_MX02 U5922 ( .S(n278), .A0(ofifoData[345]), .A1(ofifoData[601]), .Z(n3640));
Q_MX03 U5923 ( .S0(n277), .S1(n276), .A0(n2988), .A1(n2989), .A2(n3819), .Z(n2987));
Q_MX02 U5924 ( .S(n278), .A0(ofifoData[346]), .A1(ofifoData[602]), .Z(n3639));
Q_MX03 U5925 ( .S0(n277), .S1(n276), .A0(n2985), .A1(n2986), .A2(n3820), .Z(n2984));
Q_MX02 U5926 ( .S(n278), .A0(ofifoData[347]), .A1(ofifoData[603]), .Z(n3638));
Q_MX03 U5927 ( .S0(n277), .S1(n276), .A0(n2982), .A1(n2983), .A2(n3821), .Z(n2981));
Q_MX02 U5928 ( .S(n278), .A0(ofifoData[348]), .A1(ofifoData[604]), .Z(n3637));
Q_MX03 U5929 ( .S0(n277), .S1(n276), .A0(n2979), .A1(n2980), .A2(n3822), .Z(n2978));
Q_MX02 U5930 ( .S(n278), .A0(ofifoData[349]), .A1(ofifoData[605]), .Z(n3636));
Q_MX03 U5931 ( .S0(n277), .S1(n276), .A0(n2976), .A1(n2977), .A2(n3823), .Z(n2975));
Q_MX02 U5932 ( .S(n278), .A0(ofifoData[350]), .A1(ofifoData[606]), .Z(n3635));
Q_MX03 U5933 ( .S0(n277), .S1(n276), .A0(n2973), .A1(n2974), .A2(n3824), .Z(n2972));
Q_MX02 U5934 ( .S(n278), .A0(ofifoData[351]), .A1(ofifoData[607]), .Z(n3634));
Q_MX03 U5935 ( .S0(n277), .S1(n276), .A0(n2970), .A1(n2971), .A2(n3825), .Z(n2969));
Q_MX02 U5936 ( .S(n278), .A0(ofifoData[352]), .A1(ofifoData[608]), .Z(n3633));
Q_MX03 U5937 ( .S0(n277), .S1(n276), .A0(n2967), .A1(n2968), .A2(n3826), .Z(n2966));
Q_MX02 U5938 ( .S(n278), .A0(ofifoData[353]), .A1(ofifoData[609]), .Z(n3632));
Q_MX03 U5939 ( .S0(n277), .S1(n276), .A0(n2964), .A1(n2965), .A2(n3827), .Z(n2963));
Q_MX02 U5940 ( .S(n278), .A0(ofifoData[354]), .A1(ofifoData[610]), .Z(n3631));
Q_MX03 U5941 ( .S0(n277), .S1(n276), .A0(n2961), .A1(n2962), .A2(n3828), .Z(n2960));
Q_MX02 U5942 ( .S(n278), .A0(ofifoData[355]), .A1(ofifoData[611]), .Z(n3630));
Q_MX03 U5943 ( .S0(n277), .S1(n276), .A0(n2958), .A1(n2959), .A2(n3829), .Z(n2957));
Q_MX02 U5944 ( .S(n278), .A0(ofifoData[356]), .A1(ofifoData[612]), .Z(n3629));
Q_MX03 U5945 ( .S0(n277), .S1(n276), .A0(n2955), .A1(n2956), .A2(n3830), .Z(n2954));
Q_MX02 U5946 ( .S(n278), .A0(ofifoData[357]), .A1(ofifoData[613]), .Z(n3628));
Q_MX03 U5947 ( .S0(n277), .S1(n276), .A0(n2952), .A1(n2953), .A2(n3831), .Z(n2951));
Q_MX02 U5948 ( .S(n278), .A0(ofifoData[358]), .A1(ofifoData[614]), .Z(n3627));
Q_MX03 U5949 ( .S0(n277), .S1(n276), .A0(n2949), .A1(n2950), .A2(n3832), .Z(n2948));
Q_MX02 U5950 ( .S(n278), .A0(ofifoData[359]), .A1(ofifoData[615]), .Z(n3626));
Q_MX03 U5951 ( .S0(n277), .S1(n276), .A0(n2946), .A1(n2947), .A2(n3833), .Z(n2945));
Q_MX02 U5952 ( .S(n278), .A0(ofifoData[360]), .A1(ofifoData[616]), .Z(n3625));
Q_MX03 U5953 ( .S0(n277), .S1(n276), .A0(n2943), .A1(n2944), .A2(n3834), .Z(n2942));
Q_MX02 U5954 ( .S(n278), .A0(ofifoData[361]), .A1(ofifoData[617]), .Z(n3624));
Q_MX03 U5955 ( .S0(n277), .S1(n276), .A0(n2940), .A1(n2941), .A2(n3835), .Z(n2939));
Q_MX02 U5956 ( .S(n278), .A0(ofifoData[362]), .A1(ofifoData[618]), .Z(n3623));
Q_MX03 U5957 ( .S0(n277), .S1(n276), .A0(n2937), .A1(n2938), .A2(n3836), .Z(n2936));
Q_MX02 U5958 ( .S(n278), .A0(ofifoData[363]), .A1(ofifoData[619]), .Z(n3622));
Q_MX03 U5959 ( .S0(n277), .S1(n276), .A0(n2934), .A1(n2935), .A2(n3837), .Z(n2933));
Q_MX02 U5960 ( .S(n278), .A0(ofifoData[364]), .A1(ofifoData[620]), .Z(n3621));
Q_MX03 U5961 ( .S0(n277), .S1(n276), .A0(n2931), .A1(n2932), .A2(n3838), .Z(n2930));
Q_MX02 U5962 ( .S(n278), .A0(ofifoData[365]), .A1(ofifoData[621]), .Z(n3620));
Q_MX03 U5963 ( .S0(n277), .S1(n276), .A0(n2928), .A1(n2929), .A2(n3839), .Z(n2927));
Q_MX02 U5964 ( .S(n278), .A0(ofifoData[366]), .A1(ofifoData[622]), .Z(n3619));
Q_MX03 U5965 ( .S0(n277), .S1(n276), .A0(n2925), .A1(n2926), .A2(n3840), .Z(n2924));
Q_MX02 U5966 ( .S(n278), .A0(ofifoData[367]), .A1(ofifoData[623]), .Z(n3618));
Q_MX03 U5967 ( .S0(n277), .S1(n276), .A0(n2922), .A1(n2923), .A2(n3841), .Z(n2921));
Q_MX02 U5968 ( .S(n278), .A0(ofifoData[368]), .A1(ofifoData[624]), .Z(n3617));
Q_MX03 U5969 ( .S0(n277), .S1(n276), .A0(n2919), .A1(n2920), .A2(n3842), .Z(n2918));
Q_MX02 U5970 ( .S(n278), .A0(ofifoData[369]), .A1(ofifoData[625]), .Z(n3616));
Q_MX03 U5971 ( .S0(n277), .S1(n276), .A0(n2916), .A1(n2917), .A2(n3843), .Z(n2915));
Q_MX02 U5972 ( .S(n278), .A0(ofifoData[370]), .A1(ofifoData[626]), .Z(n3615));
Q_MX03 U5973 ( .S0(n277), .S1(n276), .A0(n2913), .A1(n2914), .A2(n3844), .Z(n2912));
Q_MX02 U5974 ( .S(n278), .A0(ofifoData[371]), .A1(ofifoData[627]), .Z(n3614));
Q_MX03 U5975 ( .S0(n277), .S1(n276), .A0(n2910), .A1(n2911), .A2(n3845), .Z(n2909));
Q_MX02 U5976 ( .S(n278), .A0(ofifoData[372]), .A1(ofifoData[628]), .Z(n3613));
Q_MX03 U5977 ( .S0(n277), .S1(n276), .A0(n2907), .A1(n2908), .A2(n3846), .Z(n2906));
Q_MX02 U5978 ( .S(n278), .A0(ofifoData[373]), .A1(ofifoData[629]), .Z(n3612));
Q_MX03 U5979 ( .S0(n277), .S1(n276), .A0(n2904), .A1(n2905), .A2(n3847), .Z(n2903));
Q_MX02 U5980 ( .S(n278), .A0(ofifoData[374]), .A1(ofifoData[630]), .Z(n3611));
Q_MX03 U5981 ( .S0(n277), .S1(n276), .A0(n2901), .A1(n2902), .A2(n3848), .Z(n2900));
Q_MX02 U5982 ( .S(n278), .A0(ofifoData[375]), .A1(ofifoData[631]), .Z(n3610));
Q_MX03 U5983 ( .S0(n277), .S1(n276), .A0(n2898), .A1(n2899), .A2(n3849), .Z(n2897));
Q_MX02 U5984 ( .S(n278), .A0(ofifoData[376]), .A1(ofifoData[632]), .Z(n3609));
Q_MX03 U5985 ( .S0(n277), .S1(n276), .A0(n2895), .A1(n2896), .A2(n3850), .Z(n2894));
Q_MX02 U5986 ( .S(n278), .A0(ofifoData[377]), .A1(ofifoData[633]), .Z(n3608));
Q_MX03 U5987 ( .S0(n277), .S1(n276), .A0(n2892), .A1(n2893), .A2(n3851), .Z(n2891));
Q_MX02 U5988 ( .S(n278), .A0(ofifoData[378]), .A1(ofifoData[634]), .Z(n3607));
Q_MX03 U5989 ( .S0(n277), .S1(n276), .A0(n2889), .A1(n2890), .A2(n3852), .Z(n2888));
Q_MX02 U5990 ( .S(n278), .A0(ofifoData[379]), .A1(ofifoData[635]), .Z(n3606));
Q_MX03 U5991 ( .S0(n277), .S1(n276), .A0(n2886), .A1(n2887), .A2(n3853), .Z(n2885));
Q_MX02 U5992 ( .S(n278), .A0(ofifoData[380]), .A1(ofifoData[636]), .Z(n3605));
Q_MX03 U5993 ( .S0(n277), .S1(n276), .A0(n2883), .A1(n2884), .A2(n3854), .Z(n2882));
Q_MX02 U5994 ( .S(n278), .A0(ofifoData[381]), .A1(ofifoData[637]), .Z(n3604));
Q_MX03 U5995 ( .S0(n277), .S1(n276), .A0(n2880), .A1(n2881), .A2(n3855), .Z(n2879));
Q_MX02 U5996 ( .S(n278), .A0(ofifoData[382]), .A1(ofifoData[638]), .Z(n3603));
Q_MX03 U5997 ( .S0(n277), .S1(n276), .A0(n2877), .A1(n2878), .A2(n3856), .Z(n2876));
Q_MX02 U5998 ( .S(n278), .A0(ofifoData[383]), .A1(ofifoData[639]), .Z(n3602));
Q_MX03 U5999 ( .S0(n277), .S1(n276), .A0(n2874), .A1(n2875), .A2(n3857), .Z(n2873));
Q_MX02 U6000 ( .S(n278), .A0(ofifoData[384]), .A1(ofifoData[640]), .Z(n3601));
Q_MX03 U6001 ( .S0(n277), .S1(n276), .A0(n2871), .A1(n2872), .A2(n3859), .Z(n2870));
Q_MX02 U6002 ( .S(n278), .A0(ofifoData[385]), .A1(ofifoData[641]), .Z(n3600));
Q_MX03 U6003 ( .S0(n277), .S1(n276), .A0(n2868), .A1(n2869), .A2(n3860), .Z(n2867));
Q_MX02 U6004 ( .S(n278), .A0(ofifoData[386]), .A1(ofifoData[642]), .Z(n3599));
Q_MX03 U6005 ( .S0(n277), .S1(n276), .A0(n2865), .A1(n2866), .A2(n3861), .Z(n2864));
Q_MX02 U6006 ( .S(n278), .A0(ofifoData[387]), .A1(ofifoData[643]), .Z(n3598));
Q_MX03 U6007 ( .S0(n277), .S1(n276), .A0(n2862), .A1(n2863), .A2(n3862), .Z(n2861));
Q_MX02 U6008 ( .S(n278), .A0(ofifoData[388]), .A1(ofifoData[644]), .Z(n3597));
Q_MX03 U6009 ( .S0(n277), .S1(n276), .A0(n2859), .A1(n2860), .A2(n3863), .Z(n2858));
Q_MX02 U6010 ( .S(n278), .A0(ofifoData[389]), .A1(ofifoData[645]), .Z(n3596));
Q_MX03 U6011 ( .S0(n277), .S1(n276), .A0(n2856), .A1(n2857), .A2(n3864), .Z(n2855));
Q_MX02 U6012 ( .S(n278), .A0(ofifoData[390]), .A1(ofifoData[646]), .Z(n3595));
Q_MX03 U6013 ( .S0(n277), .S1(n276), .A0(n2853), .A1(n2854), .A2(n3865), .Z(n2852));
Q_MX02 U6014 ( .S(n278), .A0(ofifoData[391]), .A1(ofifoData[647]), .Z(n3594));
Q_MX03 U6015 ( .S0(n277), .S1(n276), .A0(n2850), .A1(n2851), .A2(n3866), .Z(n2849));
Q_MX02 U6016 ( .S(n278), .A0(ofifoData[392]), .A1(ofifoData[648]), .Z(n3593));
Q_MX03 U6017 ( .S0(n277), .S1(n276), .A0(n2847), .A1(n2848), .A2(n3867), .Z(n2846));
Q_MX02 U6018 ( .S(n278), .A0(ofifoData[393]), .A1(ofifoData[649]), .Z(n3592));
Q_MX03 U6019 ( .S0(n277), .S1(n276), .A0(n2844), .A1(n2845), .A2(n3868), .Z(n2843));
Q_MX02 U6020 ( .S(n278), .A0(ofifoData[394]), .A1(ofifoData[650]), .Z(n3591));
Q_MX03 U6021 ( .S0(n277), .S1(n276), .A0(n2841), .A1(n2842), .A2(n3869), .Z(n2840));
Q_MX02 U6022 ( .S(n278), .A0(ofifoData[395]), .A1(ofifoData[651]), .Z(n3590));
Q_MX03 U6023 ( .S0(n277), .S1(n276), .A0(n2838), .A1(n2839), .A2(n3870), .Z(n2837));
Q_MX02 U6024 ( .S(n278), .A0(ofifoData[396]), .A1(ofifoData[652]), .Z(n3589));
Q_MX03 U6025 ( .S0(n277), .S1(n276), .A0(n2835), .A1(n2836), .A2(n3871), .Z(n2834));
Q_MX02 U6026 ( .S(n278), .A0(ofifoData[397]), .A1(ofifoData[653]), .Z(n3588));
Q_MX03 U6027 ( .S0(n277), .S1(n276), .A0(n2832), .A1(n2833), .A2(n3872), .Z(n2831));
Q_MX02 U6028 ( .S(n278), .A0(ofifoData[398]), .A1(ofifoData[654]), .Z(n3587));
Q_MX03 U6029 ( .S0(n277), .S1(n276), .A0(n2829), .A1(n2830), .A2(n3873), .Z(n2828));
Q_MX02 U6030 ( .S(n278), .A0(ofifoData[399]), .A1(ofifoData[655]), .Z(n3586));
Q_MX03 U6031 ( .S0(n277), .S1(n276), .A0(n2826), .A1(n2827), .A2(n3874), .Z(n2825));
Q_MX02 U6032 ( .S(n278), .A0(ofifoData[400]), .A1(ofifoData[656]), .Z(n3585));
Q_MX03 U6033 ( .S0(n277), .S1(n276), .A0(n2823), .A1(n2824), .A2(n3875), .Z(n2822));
Q_MX02 U6034 ( .S(n278), .A0(ofifoData[401]), .A1(ofifoData[657]), .Z(n3584));
Q_MX03 U6035 ( .S0(n277), .S1(n276), .A0(n2820), .A1(n2821), .A2(n3876), .Z(n2819));
Q_MX02 U6036 ( .S(n278), .A0(ofifoData[402]), .A1(ofifoData[658]), .Z(n3583));
Q_MX03 U6037 ( .S0(n277), .S1(n276), .A0(n2817), .A1(n2818), .A2(n3877), .Z(n2816));
Q_MX02 U6038 ( .S(n278), .A0(ofifoData[403]), .A1(ofifoData[659]), .Z(n3582));
Q_MX03 U6039 ( .S0(n277), .S1(n276), .A0(n2814), .A1(n2815), .A2(n3878), .Z(n2813));
Q_MX02 U6040 ( .S(n278), .A0(ofifoData[404]), .A1(ofifoData[660]), .Z(n3581));
Q_MX03 U6041 ( .S0(n277), .S1(n276), .A0(n2811), .A1(n2812), .A2(n3879), .Z(n2810));
Q_MX02 U6042 ( .S(n278), .A0(ofifoData[405]), .A1(ofifoData[661]), .Z(n3580));
Q_MX03 U6043 ( .S0(n277), .S1(n276), .A0(n2808), .A1(n2809), .A2(n3880), .Z(n2807));
Q_MX02 U6044 ( .S(n278), .A0(ofifoData[406]), .A1(ofifoData[662]), .Z(n3579));
Q_MX03 U6045 ( .S0(n277), .S1(n276), .A0(n2805), .A1(n2806), .A2(n3881), .Z(n2804));
Q_MX02 U6046 ( .S(n278), .A0(ofifoData[407]), .A1(ofifoData[663]), .Z(n3578));
Q_MX03 U6047 ( .S0(n277), .S1(n276), .A0(n2802), .A1(n2803), .A2(n3882), .Z(n2801));
Q_MX02 U6048 ( .S(n278), .A0(ofifoData[408]), .A1(ofifoData[664]), .Z(n3577));
Q_MX03 U6049 ( .S0(n277), .S1(n276), .A0(n2799), .A1(n2800), .A2(n3883), .Z(n2798));
Q_MX02 U6050 ( .S(n278), .A0(ofifoData[409]), .A1(ofifoData[665]), .Z(n3576));
Q_MX03 U6051 ( .S0(n277), .S1(n276), .A0(n2796), .A1(n2797), .A2(n3884), .Z(n2795));
Q_MX02 U6052 ( .S(n278), .A0(ofifoData[410]), .A1(ofifoData[666]), .Z(n3575));
Q_MX03 U6053 ( .S0(n277), .S1(n276), .A0(n2793), .A1(n2794), .A2(n3885), .Z(n2792));
Q_MX02 U6054 ( .S(n278), .A0(ofifoData[411]), .A1(ofifoData[667]), .Z(n3574));
Q_MX03 U6055 ( .S0(n277), .S1(n276), .A0(n2790), .A1(n2791), .A2(n3886), .Z(n2789));
Q_MX02 U6056 ( .S(n278), .A0(ofifoData[412]), .A1(ofifoData[668]), .Z(n3573));
Q_MX03 U6057 ( .S0(n277), .S1(n276), .A0(n2787), .A1(n2788), .A2(n3887), .Z(n2786));
Q_MX02 U6058 ( .S(n278), .A0(ofifoData[413]), .A1(ofifoData[669]), .Z(n3572));
Q_MX03 U6059 ( .S0(n277), .S1(n276), .A0(n2784), .A1(n2785), .A2(n3888), .Z(n2783));
Q_MX02 U6060 ( .S(n278), .A0(ofifoData[414]), .A1(ofifoData[670]), .Z(n3571));
Q_MX03 U6061 ( .S0(n277), .S1(n276), .A0(n2781), .A1(n2782), .A2(n3889), .Z(n2780));
Q_MX02 U6062 ( .S(n278), .A0(ofifoData[415]), .A1(ofifoData[671]), .Z(n3570));
Q_MX03 U6063 ( .S0(n277), .S1(n276), .A0(n2778), .A1(n2779), .A2(n3890), .Z(n2777));
Q_MX02 U6064 ( .S(n278), .A0(ofifoData[416]), .A1(ofifoData[672]), .Z(n3569));
Q_MX03 U6065 ( .S0(n277), .S1(n276), .A0(n2775), .A1(n2776), .A2(n3891), .Z(n2774));
Q_MX02 U6066 ( .S(n278), .A0(ofifoData[417]), .A1(ofifoData[673]), .Z(n3568));
Q_MX03 U6067 ( .S0(n277), .S1(n276), .A0(n2772), .A1(n2773), .A2(n3892), .Z(n2771));
Q_MX02 U6068 ( .S(n278), .A0(ofifoData[418]), .A1(ofifoData[674]), .Z(n3567));
Q_MX03 U6069 ( .S0(n277), .S1(n276), .A0(n2769), .A1(n2770), .A2(n3893), .Z(n2768));
Q_MX02 U6070 ( .S(n278), .A0(ofifoData[419]), .A1(ofifoData[675]), .Z(n3566));
Q_MX03 U6071 ( .S0(n277), .S1(n276), .A0(n2766), .A1(n2767), .A2(n3894), .Z(n2765));
Q_MX02 U6072 ( .S(n278), .A0(ofifoData[420]), .A1(ofifoData[676]), .Z(n3565));
Q_MX03 U6073 ( .S0(n277), .S1(n276), .A0(n2763), .A1(n2764), .A2(n3895), .Z(n2762));
Q_MX02 U6074 ( .S(n278), .A0(ofifoData[421]), .A1(ofifoData[677]), .Z(n3564));
Q_MX03 U6075 ( .S0(n277), .S1(n276), .A0(n2760), .A1(n2761), .A2(n3896), .Z(n2759));
Q_MX02 U6076 ( .S(n278), .A0(ofifoData[422]), .A1(ofifoData[678]), .Z(n3563));
Q_MX03 U6077 ( .S0(n277), .S1(n276), .A0(n2757), .A1(n2758), .A2(n3897), .Z(n2756));
Q_MX02 U6078 ( .S(n278), .A0(ofifoData[423]), .A1(ofifoData[679]), .Z(n3562));
Q_MX03 U6079 ( .S0(n277), .S1(n276), .A0(n2754), .A1(n2755), .A2(n3898), .Z(n2753));
Q_MX02 U6080 ( .S(n278), .A0(ofifoData[424]), .A1(ofifoData[680]), .Z(n3561));
Q_MX03 U6081 ( .S0(n277), .S1(n276), .A0(n2751), .A1(n2752), .A2(n3899), .Z(n2750));
Q_MX02 U6082 ( .S(n278), .A0(ofifoData[425]), .A1(ofifoData[681]), .Z(n3560));
Q_MX03 U6083 ( .S0(n277), .S1(n276), .A0(n2748), .A1(n2749), .A2(n3900), .Z(n2747));
Q_MX02 U6084 ( .S(n278), .A0(ofifoData[426]), .A1(ofifoData[682]), .Z(n3559));
Q_MX03 U6085 ( .S0(n277), .S1(n276), .A0(n2745), .A1(n2746), .A2(n3901), .Z(n2744));
Q_MX02 U6086 ( .S(n278), .A0(ofifoData[427]), .A1(ofifoData[683]), .Z(n3558));
Q_MX03 U6087 ( .S0(n277), .S1(n276), .A0(n2742), .A1(n2743), .A2(n3902), .Z(n2741));
Q_MX02 U6088 ( .S(n278), .A0(ofifoData[428]), .A1(ofifoData[684]), .Z(n3557));
Q_MX03 U6089 ( .S0(n277), .S1(n276), .A0(n2739), .A1(n2740), .A2(n3903), .Z(n2738));
Q_MX02 U6090 ( .S(n278), .A0(ofifoData[429]), .A1(ofifoData[685]), .Z(n3556));
Q_MX03 U6091 ( .S0(n277), .S1(n276), .A0(n2736), .A1(n2737), .A2(n3904), .Z(n2735));
Q_MX02 U6092 ( .S(n278), .A0(ofifoData[430]), .A1(ofifoData[686]), .Z(n3555));
Q_MX03 U6093 ( .S0(n277), .S1(n276), .A0(n2733), .A1(n2734), .A2(n3905), .Z(n2732));
Q_MX02 U6094 ( .S(n278), .A0(ofifoData[431]), .A1(ofifoData[687]), .Z(n3554));
Q_MX03 U6095 ( .S0(n277), .S1(n276), .A0(n2730), .A1(n2731), .A2(n3906), .Z(n2729));
Q_MX02 U6096 ( .S(n278), .A0(ofifoData[432]), .A1(ofifoData[688]), .Z(n3553));
Q_MX03 U6097 ( .S0(n277), .S1(n276), .A0(n2727), .A1(n2728), .A2(n3907), .Z(n2726));
Q_MX02 U6098 ( .S(n278), .A0(ofifoData[433]), .A1(ofifoData[689]), .Z(n3552));
Q_MX03 U6099 ( .S0(n277), .S1(n276), .A0(n2724), .A1(n2725), .A2(n3908), .Z(n2723));
Q_MX02 U6100 ( .S(n278), .A0(ofifoData[434]), .A1(ofifoData[690]), .Z(n3551));
Q_MX03 U6101 ( .S0(n277), .S1(n276), .A0(n2721), .A1(n2722), .A2(n3909), .Z(n2720));
Q_MX02 U6102 ( .S(n278), .A0(ofifoData[435]), .A1(ofifoData[691]), .Z(n3550));
Q_MX03 U6103 ( .S0(n277), .S1(n276), .A0(n2718), .A1(n2719), .A2(n3910), .Z(n2717));
Q_MX02 U6104 ( .S(n278), .A0(ofifoData[436]), .A1(ofifoData[692]), .Z(n3549));
Q_MX03 U6105 ( .S0(n277), .S1(n276), .A0(n2715), .A1(n2716), .A2(n3911), .Z(n2714));
Q_MX02 U6106 ( .S(n278), .A0(ofifoData[437]), .A1(ofifoData[693]), .Z(n3548));
Q_MX03 U6107 ( .S0(n277), .S1(n276), .A0(n2712), .A1(n2713), .A2(n3912), .Z(n2711));
Q_MX02 U6108 ( .S(n278), .A0(ofifoData[438]), .A1(ofifoData[694]), .Z(n3547));
Q_MX03 U6109 ( .S0(n277), .S1(n276), .A0(n2709), .A1(n2710), .A2(n3913), .Z(n2708));
Q_MX02 U6110 ( .S(n278), .A0(ofifoData[439]), .A1(ofifoData[695]), .Z(n3546));
Q_MX03 U6111 ( .S0(n277), .S1(n276), .A0(n2706), .A1(n2707), .A2(n3914), .Z(n2705));
Q_MX02 U6112 ( .S(n278), .A0(ofifoData[440]), .A1(ofifoData[696]), .Z(n3545));
Q_MX03 U6113 ( .S0(n277), .S1(n276), .A0(n2703), .A1(n2704), .A2(n3915), .Z(n2702));
Q_MX02 U6114 ( .S(n278), .A0(ofifoData[441]), .A1(ofifoData[697]), .Z(n3544));
Q_MX03 U6115 ( .S0(n277), .S1(n276), .A0(n2700), .A1(n2701), .A2(n3916), .Z(n2699));
Q_MX02 U6116 ( .S(n278), .A0(ofifoData[442]), .A1(ofifoData[698]), .Z(n3543));
Q_MX03 U6117 ( .S0(n277), .S1(n276), .A0(n2697), .A1(n2698), .A2(n3917), .Z(n2696));
Q_MX02 U6118 ( .S(n278), .A0(ofifoData[443]), .A1(ofifoData[699]), .Z(n3542));
Q_MX03 U6119 ( .S0(n277), .S1(n276), .A0(n2694), .A1(n2695), .A2(n3918), .Z(n2693));
Q_MX02 U6120 ( .S(n278), .A0(ofifoData[444]), .A1(ofifoData[700]), .Z(n3541));
Q_MX03 U6121 ( .S0(n277), .S1(n276), .A0(n2691), .A1(n2692), .A2(n3919), .Z(n2690));
Q_MX02 U6122 ( .S(n278), .A0(ofifoData[445]), .A1(ofifoData[701]), .Z(n3540));
Q_MX03 U6123 ( .S0(n277), .S1(n276), .A0(n2688), .A1(n2689), .A2(n3920), .Z(n2687));
Q_MX02 U6124 ( .S(n278), .A0(ofifoData[446]), .A1(ofifoData[702]), .Z(n3539));
Q_MX03 U6125 ( .S0(n277), .S1(n276), .A0(n2685), .A1(n2686), .A2(n3921), .Z(n2684));
Q_MX02 U6126 ( .S(n278), .A0(ofifoData[447]), .A1(ofifoData[703]), .Z(n3538));
Q_MX03 U6127 ( .S0(n277), .S1(n276), .A0(n2682), .A1(n2683), .A2(n3922), .Z(n2681));
Q_MX02 U6128 ( .S(n278), .A0(ofifoData[448]), .A1(ofifoData[704]), .Z(n3537));
Q_MX03 U6129 ( .S0(n277), .S1(n276), .A0(n2679), .A1(n2680), .A2(n3923), .Z(n2678));
Q_MX02 U6130 ( .S(n278), .A0(ofifoData[449]), .A1(ofifoData[705]), .Z(n3536));
Q_MX03 U6131 ( .S0(n277), .S1(n276), .A0(n2676), .A1(n2677), .A2(n3924), .Z(n2675));
Q_MX02 U6132 ( .S(n278), .A0(ofifoData[450]), .A1(ofifoData[706]), .Z(n3535));
Q_MX03 U6133 ( .S0(n277), .S1(n276), .A0(n2673), .A1(n2674), .A2(n3925), .Z(n2672));
Q_MX02 U6134 ( .S(n278), .A0(ofifoData[451]), .A1(ofifoData[707]), .Z(n3534));
Q_MX03 U6135 ( .S0(n277), .S1(n276), .A0(n2670), .A1(n2671), .A2(n3926), .Z(n2669));
Q_MX02 U6136 ( .S(n278), .A0(ofifoData[452]), .A1(ofifoData[708]), .Z(n3533));
Q_MX03 U6137 ( .S0(n277), .S1(n276), .A0(n2667), .A1(n2668), .A2(n3927), .Z(n2666));
Q_MX02 U6138 ( .S(n278), .A0(ofifoData[453]), .A1(ofifoData[709]), .Z(n3532));
Q_MX03 U6139 ( .S0(n277), .S1(n276), .A0(n2664), .A1(n2665), .A2(n3928), .Z(n2663));
Q_MX02 U6140 ( .S(n278), .A0(ofifoData[454]), .A1(ofifoData[710]), .Z(n3531));
Q_MX03 U6141 ( .S0(n277), .S1(n276), .A0(n2661), .A1(n2662), .A2(n3929), .Z(n2660));
Q_MX02 U6142 ( .S(n278), .A0(ofifoData[455]), .A1(ofifoData[711]), .Z(n3530));
Q_MX03 U6143 ( .S0(n277), .S1(n276), .A0(n2658), .A1(n2659), .A2(n3930), .Z(n2657));
Q_MX02 U6144 ( .S(n278), .A0(ofifoData[456]), .A1(ofifoData[712]), .Z(n3529));
Q_MX03 U6145 ( .S0(n277), .S1(n276), .A0(n2655), .A1(n2656), .A2(n3931), .Z(n2654));
Q_MX02 U6146 ( .S(n278), .A0(ofifoData[457]), .A1(ofifoData[713]), .Z(n3528));
Q_MX03 U6147 ( .S0(n277), .S1(n276), .A0(n2652), .A1(n2653), .A2(n3932), .Z(n2651));
Q_MX02 U6148 ( .S(n278), .A0(ofifoData[458]), .A1(ofifoData[714]), .Z(n3527));
Q_MX03 U6149 ( .S0(n277), .S1(n276), .A0(n2649), .A1(n2650), .A2(n3933), .Z(n2648));
Q_MX02 U6150 ( .S(n278), .A0(ofifoData[459]), .A1(ofifoData[715]), .Z(n3526));
Q_MX03 U6151 ( .S0(n277), .S1(n276), .A0(n2646), .A1(n2647), .A2(n3934), .Z(n2645));
Q_MX02 U6152 ( .S(n278), .A0(ofifoData[460]), .A1(ofifoData[716]), .Z(n3525));
Q_MX03 U6153 ( .S0(n277), .S1(n276), .A0(n2643), .A1(n2644), .A2(n3935), .Z(n2642));
Q_MX02 U6154 ( .S(n278), .A0(ofifoData[461]), .A1(ofifoData[717]), .Z(n3524));
Q_MX03 U6155 ( .S0(n277), .S1(n276), .A0(n2640), .A1(n2641), .A2(n3936), .Z(n2639));
Q_MX02 U6156 ( .S(n278), .A0(ofifoData[462]), .A1(ofifoData[718]), .Z(n3523));
Q_MX03 U6157 ( .S0(n277), .S1(n276), .A0(n2637), .A1(n2638), .A2(n3937), .Z(n2636));
Q_MX02 U6158 ( .S(n278), .A0(ofifoData[463]), .A1(ofifoData[719]), .Z(n3522));
Q_MX03 U6159 ( .S0(n277), .S1(n276), .A0(n2634), .A1(n2635), .A2(n3938), .Z(n2633));
Q_MX02 U6160 ( .S(n278), .A0(ofifoData[464]), .A1(ofifoData[720]), .Z(n3521));
Q_MX03 U6161 ( .S0(n277), .S1(n276), .A0(n2631), .A1(n2632), .A2(n3939), .Z(n2630));
Q_MX02 U6162 ( .S(n278), .A0(ofifoData[465]), .A1(ofifoData[721]), .Z(n3520));
Q_MX03 U6163 ( .S0(n277), .S1(n276), .A0(n2628), .A1(n2629), .A2(n3940), .Z(n2627));
Q_MX02 U6164 ( .S(n278), .A0(ofifoData[466]), .A1(ofifoData[722]), .Z(n3519));
Q_MX03 U6165 ( .S0(n277), .S1(n276), .A0(n2625), .A1(n2626), .A2(n3941), .Z(n2624));
Q_MX02 U6166 ( .S(n278), .A0(ofifoData[467]), .A1(ofifoData[723]), .Z(n3518));
Q_MX03 U6167 ( .S0(n277), .S1(n276), .A0(n2622), .A1(n2623), .A2(n3942), .Z(n2621));
Q_MX02 U6168 ( .S(n278), .A0(ofifoData[468]), .A1(ofifoData[724]), .Z(n3517));
Q_MX03 U6169 ( .S0(n277), .S1(n276), .A0(n2619), .A1(n2620), .A2(n3943), .Z(n2618));
Q_MX02 U6170 ( .S(n278), .A0(ofifoData[469]), .A1(ofifoData[725]), .Z(n3516));
Q_MX03 U6171 ( .S0(n277), .S1(n276), .A0(n2616), .A1(n2617), .A2(n3944), .Z(n2615));
Q_MX02 U6172 ( .S(n278), .A0(ofifoData[470]), .A1(ofifoData[726]), .Z(n3515));
Q_MX03 U6173 ( .S0(n277), .S1(n276), .A0(n2613), .A1(n2614), .A2(n3945), .Z(n2612));
Q_MX02 U6174 ( .S(n278), .A0(ofifoData[471]), .A1(ofifoData[727]), .Z(n3514));
Q_MX03 U6175 ( .S0(n277), .S1(n276), .A0(n2610), .A1(n2611), .A2(n3946), .Z(n2609));
Q_MX02 U6176 ( .S(n278), .A0(ofifoData[472]), .A1(ofifoData[728]), .Z(n3513));
Q_MX03 U6177 ( .S0(n277), .S1(n276), .A0(n2607), .A1(n2608), .A2(n3947), .Z(n2606));
Q_MX02 U6178 ( .S(n278), .A0(ofifoData[473]), .A1(ofifoData[729]), .Z(n3512));
Q_MX03 U6179 ( .S0(n277), .S1(n276), .A0(n2604), .A1(n2605), .A2(n3948), .Z(n2603));
Q_MX02 U6180 ( .S(n278), .A0(ofifoData[474]), .A1(ofifoData[730]), .Z(n3511));
Q_MX03 U6181 ( .S0(n277), .S1(n276), .A0(n2601), .A1(n2602), .A2(n3949), .Z(n2600));
Q_MX02 U6182 ( .S(n278), .A0(ofifoData[475]), .A1(ofifoData[731]), .Z(n3510));
Q_MX03 U6183 ( .S0(n277), .S1(n276), .A0(n2598), .A1(n2599), .A2(n3950), .Z(n2597));
Q_MX02 U6184 ( .S(n278), .A0(ofifoData[476]), .A1(ofifoData[732]), .Z(n3509));
Q_MX03 U6185 ( .S0(n277), .S1(n276), .A0(n2595), .A1(n2596), .A2(n3951), .Z(n2594));
Q_MX02 U6186 ( .S(n278), .A0(ofifoData[477]), .A1(ofifoData[733]), .Z(n3508));
Q_MX03 U6187 ( .S0(n277), .S1(n276), .A0(n2592), .A1(n2593), .A2(n3952), .Z(n2591));
Q_MX02 U6188 ( .S(n278), .A0(ofifoData[478]), .A1(ofifoData[734]), .Z(n3507));
Q_MX03 U6189 ( .S0(n277), .S1(n276), .A0(n2589), .A1(n2590), .A2(n3953), .Z(n2588));
Q_MX02 U6190 ( .S(n278), .A0(ofifoData[479]), .A1(ofifoData[735]), .Z(n3506));
Q_MX03 U6191 ( .S0(n277), .S1(n276), .A0(n2586), .A1(n2587), .A2(n3954), .Z(n2585));
Q_MX02 U6192 ( .S(n278), .A0(ofifoData[480]), .A1(ofifoData[736]), .Z(n3505));
Q_MX03 U6193 ( .S0(n277), .S1(n276), .A0(n2583), .A1(n2584), .A2(n3955), .Z(n2582));
Q_MX02 U6194 ( .S(n278), .A0(ofifoData[481]), .A1(ofifoData[737]), .Z(n3504));
Q_MX03 U6195 ( .S0(n277), .S1(n276), .A0(n2580), .A1(n2581), .A2(n3956), .Z(n2579));
Q_MX02 U6196 ( .S(n278), .A0(ofifoData[482]), .A1(ofifoData[738]), .Z(n3503));
Q_MX03 U6197 ( .S0(n277), .S1(n276), .A0(n2577), .A1(n2578), .A2(n3957), .Z(n2576));
Q_MX02 U6198 ( .S(n278), .A0(ofifoData[483]), .A1(ofifoData[739]), .Z(n3502));
Q_MX03 U6199 ( .S0(n277), .S1(n276), .A0(n2574), .A1(n2575), .A2(n3958), .Z(n2573));
Q_MX02 U6200 ( .S(n278), .A0(ofifoData[484]), .A1(ofifoData[740]), .Z(n3501));
Q_MX03 U6201 ( .S0(n277), .S1(n276), .A0(n2571), .A1(n2572), .A2(n3959), .Z(n2570));
Q_MX02 U6202 ( .S(n278), .A0(ofifoData[485]), .A1(ofifoData[741]), .Z(n3500));
Q_MX03 U6203 ( .S0(n277), .S1(n276), .A0(n2568), .A1(n2569), .A2(n3960), .Z(n2567));
Q_MX02 U6204 ( .S(n278), .A0(ofifoData[486]), .A1(ofifoData[742]), .Z(n3499));
Q_MX03 U6205 ( .S0(n277), .S1(n276), .A0(n2565), .A1(n2566), .A2(n3961), .Z(n2564));
Q_MX02 U6206 ( .S(n278), .A0(ofifoData[487]), .A1(ofifoData[743]), .Z(n3498));
Q_MX03 U6207 ( .S0(n277), .S1(n276), .A0(n2562), .A1(n2563), .A2(n3962), .Z(n2561));
Q_MX02 U6208 ( .S(n278), .A0(ofifoData[488]), .A1(ofifoData[744]), .Z(n3497));
Q_MX03 U6209 ( .S0(n277), .S1(n276), .A0(n2559), .A1(n2560), .A2(n3963), .Z(n2558));
Q_MX02 U6210 ( .S(n278), .A0(ofifoData[489]), .A1(ofifoData[745]), .Z(n3496));
Q_MX03 U6211 ( .S0(n277), .S1(n276), .A0(n2556), .A1(n2557), .A2(n3964), .Z(n2555));
Q_MX02 U6212 ( .S(n278), .A0(ofifoData[490]), .A1(ofifoData[746]), .Z(n3495));
Q_MX03 U6213 ( .S0(n277), .S1(n276), .A0(n2553), .A1(n2554), .A2(n3965), .Z(n2552));
Q_MX02 U6214 ( .S(n278), .A0(ofifoData[491]), .A1(ofifoData[747]), .Z(n3494));
Q_MX03 U6215 ( .S0(n277), .S1(n276), .A0(n2550), .A1(n2551), .A2(n3966), .Z(n2549));
Q_MX02 U6216 ( .S(n278), .A0(ofifoData[492]), .A1(ofifoData[748]), .Z(n3493));
Q_MX03 U6217 ( .S0(n277), .S1(n276), .A0(n2547), .A1(n2548), .A2(n3967), .Z(n2546));
Q_MX02 U6218 ( .S(n278), .A0(ofifoData[493]), .A1(ofifoData[749]), .Z(n3492));
Q_MX03 U6219 ( .S0(n277), .S1(n276), .A0(n2544), .A1(n2545), .A2(n3968), .Z(n2543));
Q_MX02 U6220 ( .S(n278), .A0(ofifoData[494]), .A1(ofifoData[750]), .Z(n3491));
Q_MX03 U6221 ( .S0(n277), .S1(n276), .A0(n2541), .A1(n2542), .A2(n3969), .Z(n2540));
Q_MX02 U6222 ( .S(n278), .A0(ofifoData[495]), .A1(ofifoData[751]), .Z(n3490));
Q_MX03 U6223 ( .S0(n277), .S1(n276), .A0(n2538), .A1(n2539), .A2(n3970), .Z(n2537));
Q_MX02 U6224 ( .S(n278), .A0(ofifoData[496]), .A1(ofifoData[752]), .Z(n3489));
Q_MX03 U6225 ( .S0(n277), .S1(n276), .A0(n2535), .A1(n2536), .A2(n3971), .Z(n2534));
Q_MX02 U6226 ( .S(n278), .A0(ofifoData[497]), .A1(ofifoData[753]), .Z(n3488));
Q_MX03 U6227 ( .S0(n277), .S1(n276), .A0(n2532), .A1(n2533), .A2(n3972), .Z(n2531));
Q_MX02 U6228 ( .S(n278), .A0(ofifoData[498]), .A1(ofifoData[754]), .Z(n3487));
Q_MX03 U6229 ( .S0(n277), .S1(n276), .A0(n2529), .A1(n2530), .A2(n3973), .Z(n2528));
Q_MX02 U6230 ( .S(n278), .A0(ofifoData[499]), .A1(ofifoData[755]), .Z(n3486));
Q_MX03 U6231 ( .S0(n277), .S1(n276), .A0(n2526), .A1(n2527), .A2(n3974), .Z(n2525));
Q_MX02 U6232 ( .S(n278), .A0(ofifoData[500]), .A1(ofifoData[756]), .Z(n3485));
Q_MX03 U6233 ( .S0(n277), .S1(n276), .A0(n2523), .A1(n2524), .A2(n3975), .Z(n2522));
Q_MX02 U6234 ( .S(n278), .A0(ofifoData[501]), .A1(ofifoData[757]), .Z(n3484));
Q_MX03 U6235 ( .S0(n277), .S1(n276), .A0(n2520), .A1(n2521), .A2(n3976), .Z(n2519));
Q_MX02 U6236 ( .S(n278), .A0(ofifoData[502]), .A1(ofifoData[758]), .Z(n3483));
Q_MX03 U6237 ( .S0(n277), .S1(n276), .A0(n2517), .A1(n2518), .A2(n3977), .Z(n2516));
Q_MX02 U6238 ( .S(n278), .A0(ofifoData[503]), .A1(ofifoData[759]), .Z(n3482));
Q_MX03 U6239 ( .S0(n277), .S1(n276), .A0(n2514), .A1(n2515), .A2(n3978), .Z(n2513));
Q_MX02 U6240 ( .S(n278), .A0(ofifoData[504]), .A1(ofifoData[760]), .Z(n3481));
Q_MX03 U6241 ( .S0(n277), .S1(n276), .A0(n2511), .A1(n2512), .A2(n3979), .Z(n2510));
Q_MX02 U6242 ( .S(n278), .A0(ofifoData[505]), .A1(ofifoData[761]), .Z(n3480));
Q_MX03 U6243 ( .S0(n277), .S1(n276), .A0(n2508), .A1(n2509), .A2(n3980), .Z(n2507));
Q_MX02 U6244 ( .S(n278), .A0(ofifoData[506]), .A1(ofifoData[762]), .Z(n3479));
Q_MX03 U6245 ( .S0(n277), .S1(n276), .A0(n2505), .A1(n2506), .A2(n3981), .Z(n2504));
Q_MX02 U6246 ( .S(n278), .A0(ofifoData[507]), .A1(ofifoData[763]), .Z(n3478));
Q_MX03 U6247 ( .S0(n277), .S1(n276), .A0(n2502), .A1(n2503), .A2(n3982), .Z(n2501));
Q_MX02 U6248 ( .S(n278), .A0(ofifoData[508]), .A1(ofifoData[764]), .Z(n3477));
Q_MX03 U6249 ( .S0(n277), .S1(n276), .A0(n2499), .A1(n2500), .A2(n3983), .Z(n2498));
Q_MX02 U6250 ( .S(n278), .A0(ofifoData[509]), .A1(ofifoData[765]), .Z(n3476));
Q_MX03 U6251 ( .S0(n277), .S1(n276), .A0(n2496), .A1(n2497), .A2(n3984), .Z(n2495));
Q_MX02 U6252 ( .S(n278), .A0(ofifoData[510]), .A1(ofifoData[766]), .Z(n3475));
Q_MX03 U6253 ( .S0(n277), .S1(n276), .A0(n2493), .A1(n2494), .A2(n3985), .Z(n2492));
Q_MX02 U6254 ( .S(n278), .A0(ofifoData[511]), .A1(ofifoData[767]), .Z(n3474));
Q_MX03 U6255 ( .S0(n277), .S1(n276), .A0(n2490), .A1(n2491), .A2(n3986), .Z(n2489));
Q_AN02 U6256 ( .A0(n9332), .A1(n3987), .Z(n2488));
Q_AN02 U6257 ( .A0(n9332), .A1(n3988), .Z(n2487));
Q_AN02 U6258 ( .A0(n9332), .A1(n3989), .Z(n2486));
Q_AN02 U6259 ( .A0(n9332), .A1(n3990), .Z(n2485));
Q_AN02 U6260 ( .A0(n9332), .A1(n3991), .Z(n2484));
Q_AN02 U6261 ( .A0(n9332), .A1(n3992), .Z(n2483));
Q_AN02 U6262 ( .A0(n9332), .A1(n3993), .Z(n2482));
Q_AN02 U6263 ( .A0(n9332), .A1(n3994), .Z(n2481));
Q_AN02 U6264 ( .A0(n9332), .A1(n3995), .Z(n2480));
Q_AN02 U6265 ( .A0(n9332), .A1(n3996), .Z(n2479));
Q_AN02 U6266 ( .A0(n9332), .A1(n3997), .Z(n2478));
Q_AN02 U6267 ( .A0(n9332), .A1(n3998), .Z(n2477));
Q_AN02 U6268 ( .A0(n9332), .A1(n3999), .Z(n2476));
Q_AN02 U6269 ( .A0(n9332), .A1(n4000), .Z(n2475));
Q_AN02 U6270 ( .A0(n9332), .A1(n4001), .Z(n2474));
Q_AN02 U6271 ( .A0(n9332), .A1(n4002), .Z(n2473));
Q_AN02 U6272 ( .A0(n9332), .A1(n4003), .Z(n2472));
Q_AN02 U6273 ( .A0(n9332), .A1(n4004), .Z(n2471));
Q_AN02 U6274 ( .A0(n9332), .A1(n4005), .Z(n2470));
Q_AN02 U6275 ( .A0(n9332), .A1(n4006), .Z(n2469));
Q_AN02 U6276 ( .A0(n9332), .A1(n4007), .Z(n2468));
Q_AN02 U6277 ( .A0(n9332), .A1(n4008), .Z(n2467));
Q_AN02 U6278 ( .A0(n9332), .A1(n4009), .Z(n2466));
Q_AN02 U6279 ( .A0(n9332), .A1(n4010), .Z(n2465));
Q_AN02 U6280 ( .A0(n9332), .A1(n4011), .Z(n2464));
Q_AN02 U6281 ( .A0(n9332), .A1(n4012), .Z(n2463));
Q_AN02 U6282 ( .A0(n9332), .A1(n4013), .Z(n2462));
Q_AN02 U6283 ( .A0(n9332), .A1(n4014), .Z(n2461));
Q_AN02 U6284 ( .A0(n9332), .A1(n4015), .Z(n2460));
Q_AN02 U6285 ( .A0(n9332), .A1(n4016), .Z(n2459));
Q_AN02 U6286 ( .A0(n9332), .A1(n4017), .Z(n2458));
Q_AN02 U6287 ( .A0(n9332), .A1(n4018), .Z(n2457));
Q_AN02 U6288 ( .A0(n9332), .A1(n4019), .Z(n2456));
Q_AN02 U6289 ( .A0(n9332), .A1(n4020), .Z(n2455));
Q_AN02 U6290 ( .A0(n9332), .A1(n4021), .Z(n2454));
Q_AN02 U6291 ( .A0(n9332), .A1(n4022), .Z(n2453));
Q_AN02 U6292 ( .A0(n9332), .A1(n4023), .Z(n2452));
Q_AN02 U6293 ( .A0(n9332), .A1(n4024), .Z(n2451));
Q_AN02 U6294 ( .A0(n9332), .A1(n4025), .Z(n2450));
Q_AN02 U6295 ( .A0(n9332), .A1(n4026), .Z(n2449));
Q_AN02 U6296 ( .A0(n9332), .A1(n4027), .Z(n2448));
Q_AN02 U6297 ( .A0(n9332), .A1(n4028), .Z(n2447));
Q_AN02 U6298 ( .A0(n9332), .A1(n4029), .Z(n2446));
Q_AN02 U6299 ( .A0(n9332), .A1(n4030), .Z(n2445));
Q_AN02 U6300 ( .A0(n9332), .A1(n4031), .Z(n2444));
Q_AN02 U6301 ( .A0(n9332), .A1(n4032), .Z(n2443));
Q_AN02 U6302 ( .A0(n9332), .A1(n4033), .Z(n2442));
Q_AN02 U6303 ( .A0(n9332), .A1(n4034), .Z(n2441));
Q_AN02 U6304 ( .A0(n9332), .A1(n4035), .Z(n2440));
Q_AN02 U6305 ( .A0(n9332), .A1(n4036), .Z(n2439));
Q_AN02 U6306 ( .A0(n9332), .A1(n4037), .Z(n2438));
Q_AN02 U6307 ( .A0(n9332), .A1(n4038), .Z(n2437));
Q_AN02 U6308 ( .A0(n9332), .A1(n4039), .Z(n2436));
Q_AN02 U6309 ( .A0(n9332), .A1(n4040), .Z(n2435));
Q_AN02 U6310 ( .A0(n9332), .A1(n4041), .Z(n2434));
Q_AN02 U6311 ( .A0(n9332), .A1(n4042), .Z(n2433));
Q_AN02 U6312 ( .A0(n9332), .A1(n4043), .Z(n2432));
Q_AN02 U6313 ( .A0(n9332), .A1(n4044), .Z(n2431));
Q_AN02 U6314 ( .A0(n9332), .A1(n4045), .Z(n2430));
Q_AN02 U6315 ( .A0(n9332), .A1(n4046), .Z(n2429));
Q_AN02 U6316 ( .A0(n9332), .A1(n4047), .Z(n2428));
Q_AN02 U6317 ( .A0(n9332), .A1(n4048), .Z(n2427));
Q_AN02 U6318 ( .A0(n9332), .A1(n4049), .Z(n2426));
Q_AN02 U6319 ( .A0(n9332), .A1(n4050), .Z(n2425));
Q_AN02 U6320 ( .A0(n9332), .A1(n4051), .Z(n2424));
Q_AN02 U6321 ( .A0(n9332), .A1(n4052), .Z(n2423));
Q_AN02 U6322 ( .A0(n9332), .A1(n4053), .Z(n2422));
Q_AN02 U6323 ( .A0(n9332), .A1(n4054), .Z(n2421));
Q_AN02 U6324 ( .A0(n9332), .A1(n4055), .Z(n2420));
Q_AN02 U6325 ( .A0(n9332), .A1(n4056), .Z(n2419));
Q_AN02 U6326 ( .A0(n9332), .A1(n4057), .Z(n2418));
Q_AN02 U6327 ( .A0(n9332), .A1(n4058), .Z(n2417));
Q_AN02 U6328 ( .A0(n9332), .A1(n4059), .Z(n2416));
Q_AN02 U6329 ( .A0(n9332), .A1(n4060), .Z(n2415));
Q_AN02 U6330 ( .A0(n9332), .A1(n4061), .Z(n2414));
Q_AN02 U6331 ( .A0(n9332), .A1(n4062), .Z(n2413));
Q_AN02 U6332 ( .A0(n9332), .A1(n4063), .Z(n2412));
Q_AN02 U6333 ( .A0(n9332), .A1(n4064), .Z(n2411));
Q_AN02 U6334 ( .A0(n9332), .A1(n4065), .Z(n2410));
Q_AN02 U6335 ( .A0(n9332), .A1(n4066), .Z(n2409));
Q_AN02 U6336 ( .A0(n9332), .A1(n4067), .Z(n2408));
Q_AN02 U6337 ( .A0(n9332), .A1(n4068), .Z(n2407));
Q_AN02 U6338 ( .A0(n9332), .A1(n4069), .Z(n2406));
Q_AN02 U6339 ( .A0(n9332), .A1(n4070), .Z(n2405));
Q_AN02 U6340 ( .A0(n9332), .A1(n4071), .Z(n2404));
Q_AN02 U6341 ( .A0(n9332), .A1(n4072), .Z(n2403));
Q_AN02 U6342 ( .A0(n9332), .A1(n4073), .Z(n2402));
Q_AN02 U6343 ( .A0(n9332), .A1(n4074), .Z(n2401));
Q_AN02 U6344 ( .A0(n9332), .A1(n4075), .Z(n2400));
Q_AN02 U6345 ( .A0(n9332), .A1(n4076), .Z(n2399));
Q_AN02 U6346 ( .A0(n9332), .A1(n4077), .Z(n2398));
Q_AN02 U6347 ( .A0(n9332), .A1(n4078), .Z(n2397));
Q_AN02 U6348 ( .A0(n9332), .A1(n4079), .Z(n2396));
Q_AN02 U6349 ( .A0(n9332), .A1(n4080), .Z(n2395));
Q_AN02 U6350 ( .A0(n9332), .A1(n4081), .Z(n2394));
Q_AN02 U6351 ( .A0(n9332), .A1(n4082), .Z(n2393));
Q_AN02 U6352 ( .A0(n9332), .A1(n4083), .Z(n2392));
Q_AN02 U6353 ( .A0(n9332), .A1(n4084), .Z(n2391));
Q_AN02 U6354 ( .A0(n9332), .A1(n4085), .Z(n2390));
Q_AN02 U6355 ( .A0(n9332), .A1(n4086), .Z(n2389));
Q_AN02 U6356 ( .A0(n9332), .A1(n4087), .Z(n2388));
Q_AN02 U6357 ( .A0(n9332), .A1(n4088), .Z(n2387));
Q_AN02 U6358 ( .A0(n9332), .A1(n4089), .Z(n2386));
Q_AN02 U6359 ( .A0(n9332), .A1(n4090), .Z(n2385));
Q_AN02 U6360 ( .A0(n9332), .A1(n4091), .Z(n2384));
Q_AN02 U6361 ( .A0(n9332), .A1(n4092), .Z(n2383));
Q_AN02 U6362 ( .A0(n9332), .A1(n4093), .Z(n2382));
Q_AN02 U6363 ( .A0(n9332), .A1(n4094), .Z(n2381));
Q_AN02 U6364 ( .A0(n9332), .A1(n4095), .Z(n2380));
Q_AN02 U6365 ( .A0(n9332), .A1(n4096), .Z(n2379));
Q_AN02 U6366 ( .A0(n9332), .A1(n4097), .Z(n2378));
Q_AN02 U6367 ( .A0(n9332), .A1(n4098), .Z(n2377));
Q_AN02 U6368 ( .A0(n9332), .A1(n4099), .Z(n2376));
Q_AN02 U6369 ( .A0(n9332), .A1(n4100), .Z(n2375));
Q_AN02 U6370 ( .A0(n9332), .A1(n4101), .Z(n2374));
Q_AN02 U6371 ( .A0(n9332), .A1(n4102), .Z(n2373));
Q_AN02 U6372 ( .A0(n9332), .A1(n4103), .Z(n2372));
Q_AN02 U6373 ( .A0(n9332), .A1(n4104), .Z(n2371));
Q_AN02 U6374 ( .A0(n9332), .A1(n4105), .Z(n2370));
Q_AN02 U6375 ( .A0(n9332), .A1(n4106), .Z(n2369));
Q_AN02 U6376 ( .A0(n9332), .A1(n4107), .Z(n2368));
Q_AN02 U6377 ( .A0(n9332), .A1(n4108), .Z(n2367));
Q_AN02 U6378 ( .A0(n9332), .A1(n4109), .Z(n2366));
Q_AN02 U6379 ( .A0(n9332), .A1(n4110), .Z(n2365));
Q_AN02 U6380 ( .A0(n9332), .A1(n4111), .Z(n2364));
Q_AN02 U6381 ( .A0(n9332), .A1(n4112), .Z(n2363));
Q_AN02 U6382 ( .A0(n9332), .A1(n4113), .Z(n2362));
Q_AN02 U6383 ( .A0(n9332), .A1(n4114), .Z(n2361));
Q_AN02 U6384 ( .A0(n9332), .A1(n4115), .Z(n2360));
Q_AN02 U6385 ( .A0(n9332), .A1(n4116), .Z(n2359));
Q_AN02 U6386 ( .A0(n9332), .A1(n4117), .Z(n2358));
Q_AN02 U6387 ( .A0(n9332), .A1(n4118), .Z(n2357));
Q_AN02 U6388 ( .A0(n9332), .A1(n4119), .Z(n2356));
Q_AN02 U6389 ( .A0(n9332), .A1(n4120), .Z(n2355));
Q_AN02 U6390 ( .A0(n9332), .A1(n4121), .Z(n2354));
Q_AN02 U6391 ( .A0(n9332), .A1(n4122), .Z(n2353));
Q_AN02 U6392 ( .A0(n9332), .A1(n4123), .Z(n2352));
Q_AN02 U6393 ( .A0(n9332), .A1(n4124), .Z(n2351));
Q_AN02 U6394 ( .A0(n9332), .A1(n4125), .Z(n2350));
Q_AN02 U6395 ( .A0(n9332), .A1(n4126), .Z(n2349));
Q_AN02 U6396 ( .A0(n9332), .A1(n4127), .Z(n2348));
Q_AN02 U6397 ( .A0(n9332), .A1(n4128), .Z(n2347));
Q_AN02 U6398 ( .A0(n9332), .A1(n4129), .Z(n2346));
Q_AN02 U6399 ( .A0(n9332), .A1(n4130), .Z(n2345));
Q_AN02 U6400 ( .A0(n9332), .A1(n4131), .Z(n2344));
Q_AN02 U6401 ( .A0(n9332), .A1(n4132), .Z(n2343));
Q_AN02 U6402 ( .A0(n9332), .A1(n4133), .Z(n2342));
Q_AN02 U6403 ( .A0(n9332), .A1(n4134), .Z(n2341));
Q_AN02 U6404 ( .A0(n9332), .A1(n4135), .Z(n2340));
Q_AN02 U6405 ( .A0(n9332), .A1(n4136), .Z(n2339));
Q_AN02 U6406 ( .A0(n9332), .A1(n4137), .Z(n2338));
Q_AN02 U6407 ( .A0(n9332), .A1(n4138), .Z(n2337));
Q_AN02 U6408 ( .A0(n9332), .A1(n4139), .Z(n2336));
Q_AN02 U6409 ( .A0(n9332), .A1(n4140), .Z(n2335));
Q_AN02 U6410 ( .A0(n9332), .A1(n4141), .Z(n2334));
Q_AN02 U6411 ( .A0(n9332), .A1(n4142), .Z(n2333));
Q_AN02 U6412 ( .A0(n9332), .A1(n4143), .Z(n2332));
Q_AN02 U6413 ( .A0(n9332), .A1(n4144), .Z(n2331));
Q_AN02 U6414 ( .A0(n9332), .A1(n4145), .Z(n2330));
Q_AN02 U6415 ( .A0(n9332), .A1(n4146), .Z(n2329));
Q_AN02 U6416 ( .A0(n9332), .A1(n4147), .Z(n2328));
Q_AN02 U6417 ( .A0(n9332), .A1(n4148), .Z(n2327));
Q_AN02 U6418 ( .A0(n9332), .A1(n4149), .Z(n2326));
Q_AN02 U6419 ( .A0(n9332), .A1(n4150), .Z(n2325));
Q_AN02 U6420 ( .A0(n9332), .A1(n4151), .Z(n2324));
Q_AN02 U6421 ( .A0(n9332), .A1(n4152), .Z(n2323));
Q_AN02 U6422 ( .A0(n9332), .A1(n4153), .Z(n2322));
Q_AN02 U6423 ( .A0(n9332), .A1(n4154), .Z(n2321));
Q_AN02 U6424 ( .A0(n9332), .A1(n4155), .Z(n2320));
Q_AN02 U6425 ( .A0(n9332), .A1(n4156), .Z(n2319));
Q_AN02 U6426 ( .A0(n9332), .A1(n4157), .Z(n2318));
Q_AN02 U6427 ( .A0(n9332), .A1(n4158), .Z(n2317));
Q_AN02 U6428 ( .A0(n9332), .A1(n4159), .Z(n2316));
Q_AN02 U6429 ( .A0(n9332), .A1(n4160), .Z(n2315));
Q_AN02 U6430 ( .A0(n9332), .A1(n4161), .Z(n2314));
Q_AN02 U6431 ( .A0(n9332), .A1(n4162), .Z(n2313));
Q_AN02 U6432 ( .A0(n9332), .A1(n4163), .Z(n2312));
Q_AN02 U6433 ( .A0(n9332), .A1(n4164), .Z(n2311));
Q_AN02 U6434 ( .A0(n9332), .A1(n4165), .Z(n2310));
Q_AN02 U6435 ( .A0(n9332), .A1(n4166), .Z(n2309));
Q_AN02 U6436 ( .A0(n9332), .A1(n4167), .Z(n2308));
Q_AN02 U6437 ( .A0(n9332), .A1(n4168), .Z(n2307));
Q_AN02 U6438 ( .A0(n9332), .A1(n4169), .Z(n2306));
Q_AN02 U6439 ( .A0(n9332), .A1(n4170), .Z(n2305));
Q_AN02 U6440 ( .A0(n9332), .A1(n4171), .Z(n2304));
Q_AN02 U6441 ( .A0(n9332), .A1(n4172), .Z(n2303));
Q_AN02 U6442 ( .A0(n9332), .A1(n4173), .Z(n2302));
Q_AN02 U6443 ( .A0(n9332), .A1(n4174), .Z(n2301));
Q_AN02 U6444 ( .A0(n9332), .A1(n4175), .Z(n2300));
Q_AN02 U6445 ( .A0(n9332), .A1(n4176), .Z(n2299));
Q_AN02 U6446 ( .A0(n9332), .A1(n4177), .Z(n2298));
Q_AN02 U6447 ( .A0(n9332), .A1(n4178), .Z(n2297));
Q_AN02 U6448 ( .A0(n9332), .A1(n4179), .Z(n2296));
Q_AN02 U6449 ( .A0(n9332), .A1(n4180), .Z(n2295));
Q_AN02 U6450 ( .A0(n9332), .A1(n4181), .Z(n2294));
Q_AN02 U6451 ( .A0(n9332), .A1(n4182), .Z(n2293));
Q_AN02 U6452 ( .A0(n9332), .A1(n4183), .Z(n2292));
Q_AN02 U6453 ( .A0(n9332), .A1(n4184), .Z(n2291));
Q_AN02 U6454 ( .A0(n9332), .A1(n4185), .Z(n2290));
Q_AN02 U6455 ( .A0(n9332), .A1(n4186), .Z(n2289));
Q_AN02 U6456 ( .A0(n9332), .A1(n4187), .Z(n2288));
Q_AN02 U6457 ( .A0(n9332), .A1(n4188), .Z(n2287));
Q_AN02 U6458 ( .A0(n9332), .A1(n4189), .Z(n2286));
Q_AN02 U6459 ( .A0(n9332), .A1(n4190), .Z(n2285));
Q_AN02 U6460 ( .A0(n9332), .A1(n4191), .Z(n2284));
Q_AN02 U6461 ( .A0(n9332), .A1(n4192), .Z(n2283));
Q_AN02 U6462 ( .A0(n9332), .A1(n4193), .Z(n2282));
Q_AN02 U6463 ( .A0(n9332), .A1(n4194), .Z(n2281));
Q_AN02 U6464 ( .A0(n9332), .A1(n4195), .Z(n2280));
Q_AN02 U6465 ( .A0(n9332), .A1(n4196), .Z(n2279));
Q_AN02 U6466 ( .A0(n9332), .A1(n4197), .Z(n2278));
Q_AN02 U6467 ( .A0(n9332), .A1(n4198), .Z(n2277));
Q_AN02 U6468 ( .A0(n9332), .A1(n4199), .Z(n2276));
Q_AN02 U6469 ( .A0(n9332), .A1(n4200), .Z(n2275));
Q_AN02 U6470 ( .A0(n9332), .A1(n4201), .Z(n2274));
Q_AN02 U6471 ( .A0(n9332), .A1(n4202), .Z(n2273));
Q_AN02 U6472 ( .A0(n9332), .A1(n4203), .Z(n2272));
Q_AN02 U6473 ( .A0(n9332), .A1(n4204), .Z(n2271));
Q_AN02 U6474 ( .A0(n9332), .A1(n4205), .Z(n2270));
Q_AN02 U6475 ( .A0(n9332), .A1(n4206), .Z(n2269));
Q_AN02 U6476 ( .A0(n9332), .A1(n4207), .Z(n2268));
Q_AN02 U6477 ( .A0(n9332), .A1(n4208), .Z(n2267));
Q_AN02 U6478 ( .A0(n9332), .A1(n4209), .Z(n2266));
Q_AN02 U6479 ( .A0(n9332), .A1(n4210), .Z(n2265));
Q_AN02 U6480 ( .A0(n9332), .A1(n4211), .Z(n2264));
Q_AN02 U6481 ( .A0(n9332), .A1(n4212), .Z(n2263));
Q_AN02 U6482 ( .A0(n9332), .A1(n4213), .Z(n2262));
Q_AN02 U6483 ( .A0(n9332), .A1(n4214), .Z(n2261));
Q_AN02 U6484 ( .A0(n9332), .A1(n4215), .Z(n2260));
Q_AN02 U6485 ( .A0(n9332), .A1(n4216), .Z(n2259));
Q_AN02 U6486 ( .A0(n9332), .A1(n4217), .Z(n2258));
Q_AN02 U6487 ( .A0(n9332), .A1(n4218), .Z(n2257));
Q_AN02 U6488 ( .A0(n9332), .A1(n4219), .Z(n2256));
Q_AN02 U6489 ( .A0(n9332), .A1(n4220), .Z(n2255));
Q_AN02 U6490 ( .A0(n9332), .A1(n4221), .Z(n2254));
Q_AN02 U6491 ( .A0(n9332), .A1(n4222), .Z(n2253));
Q_AN02 U6492 ( .A0(n9332), .A1(n4223), .Z(n2252));
Q_AN02 U6493 ( .A0(n9332), .A1(n4224), .Z(n2251));
Q_AN02 U6494 ( .A0(n9332), .A1(n4225), .Z(n2250));
Q_AN02 U6495 ( .A0(n9332), .A1(n4226), .Z(n2249));
Q_AN02 U6496 ( .A0(n9332), .A1(n4227), .Z(n2248));
Q_AN02 U6497 ( .A0(n9332), .A1(n4228), .Z(n2247));
Q_AN02 U6498 ( .A0(n9332), .A1(n4229), .Z(n2246));
Q_AN02 U6499 ( .A0(n9332), .A1(n4230), .Z(n2245));
Q_AN02 U6500 ( .A0(n9332), .A1(n4231), .Z(n2244));
Q_AN02 U6501 ( .A0(n9332), .A1(n4232), .Z(n2243));
Q_AN02 U6502 ( .A0(n9332), .A1(n4233), .Z(n2242));
Q_AN02 U6503 ( .A0(n9332), .A1(n4234), .Z(n2241));
Q_AN02 U6504 ( .A0(n9332), .A1(n4235), .Z(n2240));
Q_AN02 U6505 ( .A0(n9332), .A1(n4236), .Z(n2239));
Q_AN02 U6506 ( .A0(n9332), .A1(n4237), .Z(n2238));
Q_AN02 U6507 ( .A0(n9332), .A1(n4238), .Z(n2237));
Q_AN02 U6508 ( .A0(n9332), .A1(n4239), .Z(n2236));
Q_AN02 U6509 ( .A0(n9332), .A1(n4240), .Z(n2235));
Q_AN02 U6510 ( .A0(n9332), .A1(n4241), .Z(n2234));
Q_AN02 U6511 ( .A0(n9332), .A1(n4242), .Z(n2233));
Q_AN02 U6512 ( .A0(n9332), .A1(n4243), .Z(n2232));
Q_AN02 U6513 ( .A0(n9332), .A1(n4244), .Z(n2231));
Q_AN02 U6514 ( .A0(n9332), .A1(n4245), .Z(n2230));
Q_AN02 U6515 ( .A0(n9332), .A1(n4246), .Z(n2229));
Q_AN02 U6516 ( .A0(n9332), .A1(n4247), .Z(n2228));
Q_AN02 U6517 ( .A0(n9332), .A1(n4248), .Z(n2227));
Q_AN02 U6518 ( .A0(n9332), .A1(n4249), .Z(n2226));
Q_AN02 U6519 ( .A0(n9332), .A1(n4250), .Z(n2225));
Q_AN02 U6520 ( .A0(n9332), .A1(n4251), .Z(n2224));
Q_AN02 U6521 ( .A0(n9332), .A1(n4252), .Z(n2223));
Q_AN02 U6522 ( .A0(n9332), .A1(n4253), .Z(n2222));
Q_AN02 U6523 ( .A0(n9332), .A1(n4254), .Z(n2221));
Q_AN02 U6524 ( .A0(n9332), .A1(n4255), .Z(n2220));
Q_AN02 U6525 ( .A0(n9332), .A1(n4256), .Z(n2219));
Q_AN02 U6526 ( .A0(n9332), .A1(n4257), .Z(n2218));
Q_AN02 U6527 ( .A0(n9332), .A1(n4258), .Z(n2217));
Q_AN02 U6528 ( .A0(n9332), .A1(n4259), .Z(n2216));
Q_AN02 U6529 ( .A0(n9332), .A1(n4260), .Z(n2215));
Q_AN02 U6530 ( .A0(n9332), .A1(n4261), .Z(n2214));
Q_AN02 U6531 ( .A0(n9332), .A1(n4262), .Z(n2213));
Q_AN02 U6532 ( .A0(n9332), .A1(n4263), .Z(n2212));
Q_AN02 U6533 ( .A0(n9332), .A1(n4264), .Z(n2211));
Q_AN02 U6534 ( .A0(n9332), .A1(n4265), .Z(n2210));
Q_AN02 U6535 ( .A0(n9332), .A1(n4266), .Z(n2209));
Q_AN02 U6536 ( .A0(n9332), .A1(n4267), .Z(n2208));
Q_AN02 U6537 ( .A0(n9332), .A1(n4268), .Z(n2207));
Q_AN02 U6538 ( .A0(n9332), .A1(n4269), .Z(n2206));
Q_AN02 U6539 ( .A0(n9332), .A1(n4270), .Z(n2205));
Q_AN02 U6540 ( .A0(n9332), .A1(n4271), .Z(n2204));
Q_AN02 U6541 ( .A0(n9332), .A1(n4272), .Z(n2203));
Q_AN02 U6542 ( .A0(n9332), .A1(n4273), .Z(n2202));
Q_AN02 U6543 ( .A0(n9332), .A1(n4274), .Z(n2201));
Q_AN02 U6544 ( .A0(n9332), .A1(n4275), .Z(n2200));
Q_AN02 U6545 ( .A0(n9332), .A1(n4276), .Z(n2199));
Q_AN02 U6546 ( .A0(n9332), .A1(n4277), .Z(n2198));
Q_AN02 U6547 ( .A0(n9332), .A1(n4278), .Z(n2197));
Q_AN02 U6548 ( .A0(n9332), .A1(n4279), .Z(n2196));
Q_AN02 U6549 ( .A0(n9332), .A1(n4280), .Z(n2195));
Q_AN02 U6550 ( .A0(n9332), .A1(n4281), .Z(n2194));
Q_AN02 U6551 ( .A0(n9332), .A1(n4282), .Z(n2193));
Q_AN02 U6552 ( .A0(n9332), .A1(n4283), .Z(n2192));
Q_AN02 U6553 ( .A0(n9332), .A1(n4284), .Z(n2191));
Q_AN02 U6554 ( .A0(n9332), .A1(n4285), .Z(n2190));
Q_AN02 U6555 ( .A0(n9332), .A1(n4286), .Z(n2189));
Q_AN02 U6556 ( .A0(n9332), .A1(n4287), .Z(n2188));
Q_AN02 U6557 ( .A0(n9332), .A1(n4288), .Z(n2187));
Q_AN02 U6558 ( .A0(n9332), .A1(n4289), .Z(n2186));
Q_AN02 U6559 ( .A0(n9332), .A1(n4290), .Z(n2185));
Q_AN02 U6560 ( .A0(n9332), .A1(n4291), .Z(n2184));
Q_AN02 U6561 ( .A0(n9332), .A1(n4292), .Z(n2183));
Q_AN02 U6562 ( .A0(n9332), .A1(n4293), .Z(n2182));
Q_AN02 U6563 ( .A0(n9332), .A1(n4294), .Z(n2181));
Q_AN02 U6564 ( .A0(n9332), .A1(n4295), .Z(n2180));
Q_AN02 U6565 ( .A0(n9332), .A1(n4296), .Z(n2179));
Q_AN02 U6566 ( .A0(n9332), .A1(n4297), .Z(n2178));
Q_AN02 U6567 ( .A0(n9332), .A1(n4298), .Z(n2177));
Q_AN02 U6568 ( .A0(n9332), .A1(n4299), .Z(n2176));
Q_AN02 U6569 ( .A0(n9332), .A1(n4300), .Z(n2175));
Q_AN02 U6570 ( .A0(n9332), .A1(n4301), .Z(n2174));
Q_AN02 U6571 ( .A0(n9332), .A1(n4302), .Z(n2173));
Q_AN02 U6572 ( .A0(n9332), .A1(n4303), .Z(n2172));
Q_AN02 U6573 ( .A0(n9332), .A1(n4304), .Z(n2171));
Q_AN02 U6574 ( .A0(n9332), .A1(n4305), .Z(n2170));
Q_AN02 U6575 ( .A0(n9332), .A1(n4306), .Z(n2169));
Q_AN02 U6576 ( .A0(n9332), .A1(n4307), .Z(n2168));
Q_AN02 U6577 ( .A0(n9332), .A1(n4308), .Z(n2167));
Q_AN02 U6578 ( .A0(n9332), .A1(n4309), .Z(n2166));
Q_AN02 U6579 ( .A0(n9332), .A1(n4310), .Z(n2165));
Q_AN02 U6580 ( .A0(n9332), .A1(n4311), .Z(n2164));
Q_AN02 U6581 ( .A0(n9332), .A1(n4312), .Z(n2163));
Q_AN02 U6582 ( .A0(n9332), .A1(n4313), .Z(n2162));
Q_AN02 U6583 ( .A0(n9332), .A1(n4314), .Z(n2161));
Q_AN02 U6584 ( .A0(n9332), .A1(n4315), .Z(n2160));
Q_AN02 U6585 ( .A0(n9332), .A1(n4316), .Z(n2159));
Q_AN02 U6586 ( .A0(n9332), .A1(n4317), .Z(n2158));
Q_AN02 U6587 ( .A0(n9332), .A1(n4318), .Z(n2157));
Q_AN02 U6588 ( .A0(n9332), .A1(n4319), .Z(n2156));
Q_AN02 U6589 ( .A0(n9332), .A1(n4320), .Z(n2155));
Q_AN02 U6590 ( .A0(n9332), .A1(n4321), .Z(n2154));
Q_AN02 U6591 ( .A0(n9332), .A1(n4322), .Z(n2153));
Q_AN02 U6592 ( .A0(n9332), .A1(n4323), .Z(n2152));
Q_AN02 U6593 ( .A0(n9332), .A1(n4324), .Z(n2151));
Q_AN02 U6594 ( .A0(n9332), .A1(n4325), .Z(n2150));
Q_AN02 U6595 ( .A0(n9332), .A1(n4326), .Z(n2149));
Q_AN02 U6596 ( .A0(n9332), .A1(n4327), .Z(n2148));
Q_AN02 U6597 ( .A0(n9332), .A1(n4328), .Z(n2147));
Q_AN02 U6598 ( .A0(n9332), .A1(n4329), .Z(n2146));
Q_AN02 U6599 ( .A0(n9332), .A1(n4330), .Z(n2145));
Q_AN02 U6600 ( .A0(n9332), .A1(n4331), .Z(n2144));
Q_AN02 U6601 ( .A0(n9332), .A1(n4332), .Z(n2143));
Q_AN02 U6602 ( .A0(n9332), .A1(n4333), .Z(n2142));
Q_AN02 U6603 ( .A0(n9332), .A1(n4334), .Z(n2141));
Q_AN02 U6604 ( .A0(n9332), .A1(n4335), .Z(n2140));
Q_AN02 U6605 ( .A0(n9332), .A1(n4336), .Z(n2139));
Q_AN02 U6606 ( .A0(n9332), .A1(n4337), .Z(n2138));
Q_AN02 U6607 ( .A0(n9332), .A1(n4338), .Z(n2137));
Q_AN02 U6608 ( .A0(n9332), .A1(n4339), .Z(n2136));
Q_AN02 U6609 ( .A0(n9332), .A1(n4340), .Z(n2135));
Q_AN02 U6610 ( .A0(n9332), .A1(n4341), .Z(n2134));
Q_AN02 U6611 ( .A0(n9332), .A1(n4342), .Z(n2133));
Q_AN02 U6612 ( .A0(n9332), .A1(n4343), .Z(n2132));
Q_AN02 U6613 ( .A0(n9332), .A1(n4344), .Z(n2131));
Q_AN02 U6614 ( .A0(n9332), .A1(n4345), .Z(n2130));
Q_AN02 U6615 ( .A0(n9332), .A1(n4346), .Z(n2129));
Q_AN02 U6616 ( .A0(n9332), .A1(n4347), .Z(n2128));
Q_AN02 U6617 ( .A0(n9332), .A1(n4348), .Z(n2127));
Q_AN02 U6618 ( .A0(n9332), .A1(n4349), .Z(n2126));
Q_AN02 U6619 ( .A0(n9332), .A1(n4350), .Z(n2125));
Q_AN02 U6620 ( .A0(n9332), .A1(n4351), .Z(n2124));
Q_AN02 U6621 ( .A0(n9332), .A1(n4352), .Z(n2123));
Q_AN02 U6622 ( .A0(n9332), .A1(n4353), .Z(n2122));
Q_AN02 U6623 ( .A0(n9332), .A1(n4354), .Z(n2121));
Q_AN02 U6624 ( .A0(n9332), .A1(n4355), .Z(n2120));
Q_AN02 U6625 ( .A0(n9332), .A1(n4356), .Z(n2119));
Q_AN02 U6626 ( .A0(n9332), .A1(n4357), .Z(n2118));
Q_AN02 U6627 ( .A0(n9332), .A1(n4358), .Z(n2117));
Q_AN02 U6628 ( .A0(n9332), .A1(n4359), .Z(n2116));
Q_AN02 U6629 ( .A0(n9332), .A1(n4360), .Z(n2115));
Q_AN02 U6630 ( .A0(n9332), .A1(n4361), .Z(n2114));
Q_AN02 U6631 ( .A0(n9332), .A1(n4362), .Z(n2113));
Q_AN02 U6632 ( .A0(n9332), .A1(n4363), .Z(n2112));
Q_AN02 U6633 ( .A0(n9332), .A1(n4364), .Z(n2111));
Q_AN02 U6634 ( .A0(n9332), .A1(n4365), .Z(n2110));
Q_AN02 U6635 ( .A0(n9332), .A1(n4366), .Z(n2109));
Q_AN02 U6636 ( .A0(n9332), .A1(n4367), .Z(n2108));
Q_AN02 U6637 ( .A0(n9332), .A1(n4368), .Z(n2107));
Q_AN02 U6638 ( .A0(n9332), .A1(n4369), .Z(n2106));
Q_AN02 U6639 ( .A0(n9332), .A1(n4370), .Z(n2105));
Q_AN02 U6640 ( .A0(n9332), .A1(n4371), .Z(n2104));
Q_AN02 U6641 ( .A0(n9332), .A1(n4372), .Z(n2103));
Q_AN02 U6642 ( .A0(n9332), .A1(n4373), .Z(n2102));
Q_AN02 U6643 ( .A0(n9332), .A1(n4374), .Z(n2101));
Q_AN02 U6644 ( .A0(n9332), .A1(n4375), .Z(n2100));
Q_AN02 U6645 ( .A0(n9332), .A1(n4376), .Z(n2099));
Q_AN02 U6646 ( .A0(n9332), .A1(n4377), .Z(n2098));
Q_AN02 U6647 ( .A0(n9332), .A1(n4378), .Z(n2097));
Q_AN02 U6648 ( .A0(n9332), .A1(n4379), .Z(n2096));
Q_AN02 U6649 ( .A0(n9332), .A1(n4380), .Z(n2095));
Q_AN02 U6650 ( .A0(n9332), .A1(n4381), .Z(n2094));
Q_AN02 U6651 ( .A0(n9332), .A1(n4382), .Z(n2093));
Q_AN02 U6652 ( .A0(n9332), .A1(n4383), .Z(n2092));
Q_AN02 U6653 ( .A0(n9332), .A1(n4384), .Z(n2091));
Q_AN02 U6654 ( .A0(n9332), .A1(n4385), .Z(n2090));
Q_AN02 U6655 ( .A0(n9332), .A1(n4386), .Z(n2089));
Q_AN02 U6656 ( .A0(n9332), .A1(n4387), .Z(n2088));
Q_AN02 U6657 ( .A0(n9332), .A1(n4388), .Z(n2087));
Q_AN02 U6658 ( .A0(n9332), .A1(n4389), .Z(n2086));
Q_AN02 U6659 ( .A0(n9332), .A1(n4390), .Z(n2085));
Q_AN02 U6660 ( .A0(n9332), .A1(n4391), .Z(n2084));
Q_AN02 U6661 ( .A0(n9332), .A1(n4392), .Z(n2083));
Q_AN02 U6662 ( .A0(n9332), .A1(n4393), .Z(n2082));
Q_AN02 U6663 ( .A0(n9332), .A1(n4394), .Z(n2081));
Q_AN02 U6664 ( .A0(n9332), .A1(n4395), .Z(n2080));
Q_AN02 U6665 ( .A0(n9332), .A1(n4396), .Z(n2079));
Q_AN02 U6666 ( .A0(n9332), .A1(n4397), .Z(n2078));
Q_AN02 U6667 ( .A0(n9332), .A1(n4398), .Z(n2077));
Q_AN02 U6668 ( .A0(n9332), .A1(n4399), .Z(n2076));
Q_AN02 U6669 ( .A0(n9332), .A1(n4400), .Z(n2075));
Q_AN02 U6670 ( .A0(n9332), .A1(n4401), .Z(n2074));
Q_AN02 U6671 ( .A0(n9332), .A1(n4402), .Z(n2073));
Q_AN02 U6672 ( .A0(n9332), .A1(n4403), .Z(n2072));
Q_AN02 U6673 ( .A0(n9332), .A1(n4404), .Z(n2071));
Q_AN02 U6674 ( .A0(n9332), .A1(n4405), .Z(n2070));
Q_AN02 U6675 ( .A0(n9332), .A1(n4406), .Z(n2069));
Q_AN02 U6676 ( .A0(n9332), .A1(n4407), .Z(n2068));
Q_AN02 U6677 ( .A0(n9332), .A1(n4408), .Z(n2067));
Q_AN02 U6678 ( .A0(n9332), .A1(n4409), .Z(n2066));
Q_AN02 U6679 ( .A0(n9332), .A1(n4410), .Z(n2065));
Q_AN02 U6680 ( .A0(n9332), .A1(n4411), .Z(n2064));
Q_AN02 U6681 ( .A0(n9332), .A1(n4412), .Z(n2063));
Q_AN02 U6682 ( .A0(n9332), .A1(n4413), .Z(n2062));
Q_AN02 U6683 ( .A0(n9332), .A1(n4414), .Z(n2061));
Q_AN02 U6684 ( .A0(n9332), .A1(n4415), .Z(n2060));
Q_AN02 U6685 ( .A0(n9332), .A1(n4416), .Z(n2059));
Q_AN02 U6686 ( .A0(n9332), .A1(n4417), .Z(n2058));
Q_AN02 U6687 ( .A0(n9332), .A1(n4418), .Z(n2057));
Q_AN02 U6688 ( .A0(n9332), .A1(n4419), .Z(n2056));
Q_AN02 U6689 ( .A0(n9332), .A1(n4420), .Z(n2055));
Q_AN02 U6690 ( .A0(n9332), .A1(n4421), .Z(n2054));
Q_AN02 U6691 ( .A0(n9332), .A1(n4422), .Z(n2053));
Q_AN02 U6692 ( .A0(n9332), .A1(n4423), .Z(n2052));
Q_AN02 U6693 ( .A0(n9332), .A1(n4424), .Z(n2051));
Q_AN02 U6694 ( .A0(n9332), .A1(n4425), .Z(n2050));
Q_AN02 U6695 ( .A0(n9332), .A1(n4426), .Z(n2049));
Q_AN02 U6696 ( .A0(n9332), .A1(n4427), .Z(n2048));
Q_AN02 U6697 ( .A0(n9332), .A1(n4428), .Z(n2047));
Q_AN02 U6698 ( .A0(n9332), .A1(n4429), .Z(n2046));
Q_AN02 U6699 ( .A0(n9332), .A1(n4430), .Z(n2045));
Q_AN02 U6700 ( .A0(n9332), .A1(n4431), .Z(n2044));
Q_AN02 U6701 ( .A0(n9332), .A1(n4432), .Z(n2043));
Q_AN02 U6702 ( .A0(n9332), .A1(n4433), .Z(n2042));
Q_AN02 U6703 ( .A0(n9332), .A1(n4434), .Z(n2041));
Q_AN02 U6704 ( .A0(n279), .A1(n3469), .Z(n2040));
Q_AN02 U6705 ( .A0(n279), .A1(n3468), .Z(n2039));
Q_AN02 U6706 ( .A0(n279), .A1(n3466), .Z(n2038));
Q_AN02 U6707 ( .A0(n279), .A1(n3464), .Z(n2037));
Q_AN02 U6708 ( .A0(n279), .A1(n3462), .Z(n2036));
Q_AN02 U6709 ( .A0(n279), .A1(n3460), .Z(n2035));
Q_AN02 U6710 ( .A0(n279), .A1(n3458), .Z(n2034));
Q_AN02 U6711 ( .A0(n279), .A1(n3456), .Z(n2033));
Q_AN02 U6712 ( .A0(n279), .A1(n3454), .Z(n2032));
Q_AN02 U6713 ( .A0(n279), .A1(n3452), .Z(n2031));
Q_AN02 U6714 ( .A0(n279), .A1(n3450), .Z(n2030));
Q_AN02 U6715 ( .A0(n279), .A1(n3448), .Z(n2029));
Q_AN02 U6716 ( .A0(n279), .A1(n3446), .Z(n2028));
Q_AN02 U6717 ( .A0(n279), .A1(n3444), .Z(n2027));
Q_AN02 U6718 ( .A0(n279), .A1(n3442), .Z(n2026));
Q_AN02 U6719 ( .A0(n279), .A1(n3440), .Z(n2025));
Q_AN02 U6720 ( .A0(n279), .A1(n3438), .Z(n2024));
Q_AN02 U6721 ( .A0(n279), .A1(n3436), .Z(n2023));
Q_AN02 U6722 ( .A0(n279), .A1(n3434), .Z(n2022));
Q_AN02 U6723 ( .A0(n279), .A1(n3432), .Z(n2021));
Q_AN02 U6724 ( .A0(n279), .A1(n3430), .Z(n2020));
Q_AN02 U6725 ( .A0(n279), .A1(n3428), .Z(n2019));
Q_AN02 U6726 ( .A0(n279), .A1(n3426), .Z(n2018));
Q_AN02 U6727 ( .A0(n279), .A1(n3424), .Z(n2017));
Q_AN02 U6728 ( .A0(n279), .A1(n3422), .Z(n2016));
Q_AN02 U6729 ( .A0(n279), .A1(n3420), .Z(n2015));
Q_AN02 U6730 ( .A0(n279), .A1(n3418), .Z(n2014));
Q_AN02 U6731 ( .A0(n279), .A1(n3416), .Z(n2013));
Q_AN02 U6732 ( .A0(n279), .A1(n3414), .Z(n2012));
Q_AN02 U6733 ( .A0(n279), .A1(n3412), .Z(n2011));
Q_AN02 U6734 ( .A0(n279), .A1(n3410), .Z(n2010));
Q_AN02 U6735 ( .A0(n279), .A1(n3408), .Z(n2009));
Q_AN02 U6736 ( .A0(n279), .A1(rdCnt[0]), .Z(n2008));
Q_AN02 U6737 ( .A0(n279), .A1(rdCnt[1]), .Z(n2007));
Q_AN02 U6738 ( .A0(n279), .A1(rdCnt[2]), .Z(n2006));
Q_AN02 U6739 ( .A0(n279), .A1(rdCnt[3]), .Z(n2005));
Q_AN02 U6740 ( .A0(n279), .A1(rdCnt[4]), .Z(n2004));
Q_AN02 U6741 ( .A0(n279), .A1(rdCnt[5]), .Z(n2003));
Q_AN02 U6742 ( .A0(n279), .A1(rdCnt[6]), .Z(n2002));
Q_AN02 U6743 ( .A0(n279), .A1(rdCnt[7]), .Z(n2001));
Q_AN02 U6744 ( .A0(n279), .A1(rdCnt[8]), .Z(n2000));
Q_AN02 U6745 ( .A0(n279), .A1(rdCnt[9]), .Z(n1999));
Q_AN02 U6746 ( .A0(n279), .A1(rdCnt[10]), .Z(n1998));
Q_AN02 U6747 ( .A0(n279), .A1(rdCnt[11]), .Z(n1997));
Q_AN02 U6748 ( .A0(n279), .A1(rdCnt[12]), .Z(n1996));
Q_AN02 U6749 ( .A0(n279), .A1(rdCnt[13]), .Z(n1995));
Q_AN02 U6750 ( .A0(n279), .A1(rdCnt[14]), .Z(n1994));
Q_AN02 U6751 ( .A0(n279), .A1(rdCnt[15]), .Z(n1993));
Q_AN02 U6752 ( .A0(n279), .A1(rdCnt[16]), .Z(n1992));
Q_AN02 U6753 ( .A0(n279), .A1(rdCnt[17]), .Z(n1991));
Q_AN02 U6754 ( .A0(n279), .A1(rdCnt[18]), .Z(n1990));
Q_AN02 U6755 ( .A0(n279), .A1(rdCnt[19]), .Z(n1989));
Q_AN02 U6756 ( .A0(n279), .A1(rdCnt[20]), .Z(n1988));
Q_AN02 U6757 ( .A0(n279), .A1(rdCnt[21]), .Z(n1987));
Q_AN02 U6758 ( .A0(n279), .A1(rdCnt[22]), .Z(n1986));
Q_AN02 U6759 ( .A0(n279), .A1(rdCnt[23]), .Z(n1985));
Q_AN02 U6760 ( .A0(n279), .A1(rdCnt[24]), .Z(n1984));
Q_AN02 U6761 ( .A0(n279), .A1(rdCnt[25]), .Z(n1983));
Q_AN02 U6762 ( .A0(n279), .A1(rdCnt[26]), .Z(n1982));
Q_AN02 U6763 ( .A0(n279), .A1(rdCnt[27]), .Z(n1981));
Q_AN02 U6764 ( .A0(n279), .A1(rdCnt[28]), .Z(n1980));
Q_AN02 U6765 ( .A0(n279), .A1(rdCnt[29]), .Z(n1979));
Q_AN02 U6766 ( .A0(n279), .A1(rdCnt[30]), .Z(n1978));
Q_AN02 U6767 ( .A0(n279), .A1(rdCnt[31]), .Z(n1977));
Q_AN02 U6768 ( .A0(n279), .A1(rdCnt[32]), .Z(n1976));
Q_AN02 U6769 ( .A0(n279), .A1(rdCnt[33]), .Z(n1975));
Q_AN02 U6770 ( .A0(n279), .A1(rdCnt[34]), .Z(n1974));
Q_AN02 U6771 ( .A0(n279), .A1(rdCnt[35]), .Z(n1973));
Q_AN02 U6772 ( .A0(n279), .A1(rdCnt[36]), .Z(n1972));
Q_AN02 U6773 ( .A0(n279), .A1(rdCnt[37]), .Z(n1971));
Q_AN02 U6774 ( .A0(n279), .A1(rdCnt[38]), .Z(n1970));
Q_AN02 U6775 ( .A0(n279), .A1(rdCnt[39]), .Z(n1969));
Q_AN02 U6776 ( .A0(n279), .A1(rdCnt[40]), .Z(n1968));
Q_AN02 U6777 ( .A0(n279), .A1(rdCnt[41]), .Z(n1967));
Q_AN02 U6778 ( .A0(n279), .A1(rdCnt[42]), .Z(n1966));
Q_AN02 U6779 ( .A0(n279), .A1(rdCnt[43]), .Z(n1965));
Q_AN02 U6780 ( .A0(n279), .A1(rdCnt[44]), .Z(n1964));
Q_AN02 U6781 ( .A0(n279), .A1(rdCnt[45]), .Z(n1963));
Q_AN02 U6782 ( .A0(n279), .A1(rdCnt[46]), .Z(n1962));
Q_AN02 U6783 ( .A0(n279), .A1(rdCnt[47]), .Z(n1961));
Q_AN02 U6784 ( .A0(n279), .A1(rdCnt[48]), .Z(n1960));
Q_AN02 U6785 ( .A0(n279), .A1(rdCnt[49]), .Z(n1959));
Q_AN02 U6786 ( .A0(n279), .A1(rdCnt[50]), .Z(n1958));
Q_AN02 U6787 ( .A0(n279), .A1(rdCnt[51]), .Z(n1957));
Q_AN02 U6788 ( .A0(n279), .A1(rdCnt[52]), .Z(n1956));
Q_AN02 U6789 ( .A0(n279), .A1(rdCnt[53]), .Z(n1955));
Q_AN02 U6790 ( .A0(n279), .A1(rdCnt[54]), .Z(n1954));
Q_AN02 U6791 ( .A0(n279), .A1(rdCnt[55]), .Z(n1953));
Q_AN02 U6792 ( .A0(n279), .A1(rdCnt[56]), .Z(n1952));
Q_AN02 U6793 ( .A0(n279), .A1(rdCnt[57]), .Z(n1951));
Q_AN02 U6794 ( .A0(n279), .A1(rdCnt[58]), .Z(n1950));
Q_AN02 U6795 ( .A0(n279), .A1(rdCnt[59]), .Z(n1949));
Q_AN02 U6796 ( .A0(n279), .A1(rdCnt[60]), .Z(n1948));
Q_AN02 U6797 ( .A0(n279), .A1(rdCnt[61]), .Z(n1947));
Q_AN02 U6798 ( .A0(n279), .A1(rdCnt[62]), .Z(n1946));
Q_NR02 U6799 ( .A0(xc_top.GFReset), .A1(oMark[63]), .Z(n1945));
Q_NR02 U6800 ( .A0(xc_top.GFReset), .A1(oMark[127]), .Z(n1944));
Q_NR02 U6801 ( .A0(xc_top.GFReset), .A1(oMark[191]), .Z(n1943));
Q_NR02 U6802 ( .A0(xc_top.GFReset), .A1(oMark[255]), .Z(n1942));
Q_AN02 U6803 ( .A0(n280), .A1(n3352), .Z(n1941));
Q_AN02 U6804 ( .A0(n280), .A1(n3350), .Z(n1940));
Q_AN02 U6805 ( .A0(n280), .A1(n3348), .Z(n1939));
Q_AN02 U6806 ( .A0(n280), .A1(n3346), .Z(n1938));
Q_FDP0UA U6807 ( .D(n1937), .QTFCLK( ), .Q(oMark[255]));
Q_MX02 U6808 ( .S(n283), .A0(n1942), .A1(oMark[255]), .Z(n1937));
Q_FDP0UA U6809 ( .D(n1936), .QTFCLK( ), .Q(oMark[191]));
Q_MX02 U6810 ( .S(n283), .A0(n1943), .A1(oMark[191]), .Z(n1936));
Q_FDP0UA U6811 ( .D(n1935), .QTFCLK( ), .Q(oMark[127]));
Q_MX02 U6812 ( .S(n283), .A0(n1944), .A1(oMark[127]), .Z(n1935));
Q_FDP0UA U6813 ( .D(n1934), .QTFCLK( ), .Q(oMark[63]));
Q_MX02 U6814 ( .S(n283), .A0(n1945), .A1(oMark[63]), .Z(n1934));
Q_FDP0UA U6815 ( .D(n1946), .QTFCLK( ), .Q(oMark[62]));
Q_FDP0UA U6816 ( .D(n1947), .QTFCLK( ), .Q(oMark[61]));
Q_FDP0UA U6817 ( .D(n1948), .QTFCLK( ), .Q(oMark[60]));
Q_FDP0UA U6818 ( .D(n1949), .QTFCLK( ), .Q(oMark[59]));
Q_FDP0UA U6819 ( .D(n1950), .QTFCLK( ), .Q(oMark[58]));
Q_FDP0UA U6820 ( .D(n1951), .QTFCLK( ), .Q(oMark[57]));
Q_FDP0UA U6821 ( .D(n1952), .QTFCLK( ), .Q(oMark[56]));
Q_FDP0UA U6822 ( .D(n1953), .QTFCLK( ), .Q(oMark[55]));
Q_FDP0UA U6823 ( .D(n1954), .QTFCLK( ), .Q(oMark[54]));
Q_FDP0UA U6824 ( .D(n1955), .QTFCLK( ), .Q(oMark[53]));
Q_FDP0UA U6825 ( .D(n1956), .QTFCLK( ), .Q(oMark[52]));
Q_FDP0UA U6826 ( .D(n1957), .QTFCLK( ), .Q(oMark[51]));
Q_FDP0UA U6827 ( .D(n1958), .QTFCLK( ), .Q(oMark[50]));
Q_FDP0UA U6828 ( .D(n1959), .QTFCLK( ), .Q(oMark[49]));
Q_FDP0UA U6829 ( .D(n1960), .QTFCLK( ), .Q(oMark[48]));
Q_FDP0UA U6830 ( .D(n1961), .QTFCLK( ), .Q(oMark[47]));
Q_FDP0UA U6831 ( .D(n1962), .QTFCLK( ), .Q(oMark[46]));
Q_FDP0UA U6832 ( .D(n1963), .QTFCLK( ), .Q(oMark[45]));
Q_FDP0UA U6833 ( .D(n1964), .QTFCLK( ), .Q(oMark[44]));
Q_FDP0UA U6834 ( .D(n1965), .QTFCLK( ), .Q(oMark[43]));
Q_FDP0UA U6835 ( .D(n1966), .QTFCLK( ), .Q(oMark[42]));
Q_FDP0UA U6836 ( .D(n1967), .QTFCLK( ), .Q(oMark[41]));
Q_FDP0UA U6837 ( .D(n1968), .QTFCLK( ), .Q(oMark[40]));
Q_FDP0UA U6838 ( .D(n1969), .QTFCLK( ), .Q(oMark[39]));
Q_FDP0UA U6839 ( .D(n1970), .QTFCLK( ), .Q(oMark[38]));
Q_FDP0UA U6840 ( .D(n1971), .QTFCLK( ), .Q(oMark[37]));
Q_FDP0UA U6841 ( .D(n1972), .QTFCLK( ), .Q(oMark[36]));
Q_FDP0UA U6842 ( .D(n1973), .QTFCLK( ), .Q(oMark[35]));
Q_FDP0UA U6843 ( .D(n1974), .QTFCLK( ), .Q(oMark[34]));
Q_FDP0UA U6844 ( .D(n1975), .QTFCLK( ), .Q(oMark[33]));
Q_FDP0UA U6845 ( .D(n1976), .QTFCLK( ), .Q(oMark[32]));
Q_FDP0UA U6846 ( .D(n1977), .QTFCLK( ), .Q(oMark[31]));
Q_FDP0UA U6847 ( .D(n1978), .QTFCLK( ), .Q(oMark[30]));
Q_FDP0UA U6848 ( .D(n1979), .QTFCLK( ), .Q(oMark[29]));
Q_FDP0UA U6849 ( .D(n1980), .QTFCLK( ), .Q(oMark[28]));
Q_FDP0UA U6850 ( .D(n1981), .QTFCLK( ), .Q(oMark[27]));
Q_FDP0UA U6851 ( .D(n1982), .QTFCLK( ), .Q(oMark[26]));
Q_FDP0UA U6852 ( .D(n1983), .QTFCLK( ), .Q(oMark[25]));
Q_FDP0UA U6853 ( .D(n1984), .QTFCLK( ), .Q(oMark[24]));
Q_FDP0UA U6854 ( .D(n1985), .QTFCLK( ), .Q(oMark[23]));
Q_FDP0UA U6855 ( .D(n1986), .QTFCLK( ), .Q(oMark[22]));
Q_FDP0UA U6856 ( .D(n1987), .QTFCLK( ), .Q(oMark[21]));
Q_FDP0UA U6857 ( .D(n1988), .QTFCLK( ), .Q(oMark[20]));
Q_FDP0UA U6858 ( .D(n1989), .QTFCLK( ), .Q(oMark[19]));
Q_FDP0UA U6859 ( .D(n1990), .QTFCLK( ), .Q(oMark[18]));
Q_FDP0UA U6860 ( .D(n1991), .QTFCLK( ), .Q(oMark[17]));
Q_FDP0UA U6861 ( .D(n1992), .QTFCLK( ), .Q(oMark[16]));
Q_FDP0UA U6862 ( .D(n1993), .QTFCLK( ), .Q(oMark[15]));
Q_FDP0UA U6863 ( .D(n1994), .QTFCLK( ), .Q(oMark[14]));
Q_FDP0UA U6864 ( .D(n1995), .QTFCLK( ), .Q(oMark[13]));
Q_FDP0UA U6865 ( .D(n1996), .QTFCLK( ), .Q(oMark[12]));
Q_FDP0UA U6866 ( .D(n1997), .QTFCLK( ), .Q(oMark[11]));
Q_FDP0UA U6867 ( .D(n1998), .QTFCLK( ), .Q(oMark[10]));
Q_FDP0UA U6868 ( .D(n1999), .QTFCLK( ), .Q(oMark[9]));
Q_FDP0UA U6869 ( .D(n2000), .QTFCLK( ), .Q(oMark[8]));
Q_FDP0UA U6870 ( .D(n2001), .QTFCLK( ), .Q(oMark[7]));
Q_FDP0UA U6871 ( .D(n2002), .QTFCLK( ), .Q(oMark[6]));
Q_FDP0UA U6872 ( .D(n2003), .QTFCLK( ), .Q(oMark[5]));
Q_FDP0UA U6873 ( .D(n2004), .QTFCLK( ), .Q(oMark[4]));
Q_FDP0UA U6874 ( .D(n2005), .QTFCLK( ), .Q(oMark[3]));
Q_FDP0UA U6875 ( .D(n2006), .QTFCLK( ), .Q(oMark[2]));
Q_FDP0UA U6876 ( .D(n2007), .QTFCLK( ), .Q(oMark[1]));
Q_FDP0UA U6877 ( .D(n2008), .QTFCLK( ), .Q(oMark[0]));
Q_FDP0UA U6878 ( .D(n1933), .QTFCLK( ), .Q(numRsts[31]));
Q_MX02 U6879 ( .S(n283), .A0(n2009), .A1(numRsts[31]), .Z(n1933));
Q_FDP0UA U6880 ( .D(n1932), .QTFCLK( ), .Q(numRsts[30]));
Q_MX02 U6881 ( .S(n283), .A0(n2010), .A1(numRsts[30]), .Z(n1932));
Q_FDP0UA U6882 ( .D(n1931), .QTFCLK( ), .Q(numRsts[29]));
Q_MX02 U6883 ( .S(n283), .A0(n2011), .A1(numRsts[29]), .Z(n1931));
Q_FDP0UA U6884 ( .D(n1930), .QTFCLK( ), .Q(numRsts[28]));
Q_MX02 U6885 ( .S(n283), .A0(n2012), .A1(numRsts[28]), .Z(n1930));
Q_FDP0UA U6886 ( .D(n1929), .QTFCLK( ), .Q(numRsts[27]));
Q_MX02 U6887 ( .S(n283), .A0(n2013), .A1(numRsts[27]), .Z(n1929));
Q_FDP0UA U6888 ( .D(n1928), .QTFCLK( ), .Q(numRsts[26]));
Q_MX02 U6889 ( .S(n283), .A0(n2014), .A1(numRsts[26]), .Z(n1928));
Q_FDP0UA U6890 ( .D(n1927), .QTFCLK( ), .Q(numRsts[25]));
Q_MX02 U6891 ( .S(n283), .A0(n2015), .A1(numRsts[25]), .Z(n1927));
Q_FDP0UA U6892 ( .D(n1926), .QTFCLK( ), .Q(numRsts[24]));
Q_MX02 U6893 ( .S(n283), .A0(n2016), .A1(numRsts[24]), .Z(n1926));
Q_FDP0UA U6894 ( .D(n1925), .QTFCLK( ), .Q(numRsts[23]));
Q_MX02 U6895 ( .S(n283), .A0(n2017), .A1(numRsts[23]), .Z(n1925));
Q_FDP0UA U6896 ( .D(n1924), .QTFCLK( ), .Q(numRsts[22]));
Q_MX02 U6897 ( .S(n283), .A0(n2018), .A1(numRsts[22]), .Z(n1924));
Q_FDP0UA U6898 ( .D(n1923), .QTFCLK( ), .Q(numRsts[21]));
Q_MX02 U6899 ( .S(n283), .A0(n2019), .A1(numRsts[21]), .Z(n1923));
Q_FDP0UA U6900 ( .D(n1922), .QTFCLK( ), .Q(numRsts[20]));
Q_MX02 U6901 ( .S(n283), .A0(n2020), .A1(numRsts[20]), .Z(n1922));
Q_FDP0UA U6902 ( .D(n1921), .QTFCLK( ), .Q(numRsts[19]));
Q_MX02 U6903 ( .S(n283), .A0(n2021), .A1(numRsts[19]), .Z(n1921));
Q_FDP0UA U6904 ( .D(n1920), .QTFCLK( ), .Q(numRsts[18]));
Q_MX02 U6905 ( .S(n283), .A0(n2022), .A1(numRsts[18]), .Z(n1920));
Q_FDP0UA U6906 ( .D(n1919), .QTFCLK( ), .Q(numRsts[17]));
Q_MX02 U6907 ( .S(n283), .A0(n2023), .A1(numRsts[17]), .Z(n1919));
Q_FDP0UA U6908 ( .D(n1918), .QTFCLK( ), .Q(numRsts[16]));
Q_MX02 U6909 ( .S(n283), .A0(n2024), .A1(numRsts[16]), .Z(n1918));
Q_FDP0UA U6910 ( .D(n1917), .QTFCLK( ), .Q(numRsts[15]));
Q_MX02 U6911 ( .S(n283), .A0(n2025), .A1(numRsts[15]), .Z(n1917));
Q_FDP0UA U6912 ( .D(n1916), .QTFCLK( ), .Q(numRsts[14]));
Q_MX02 U6913 ( .S(n283), .A0(n2026), .A1(numRsts[14]), .Z(n1916));
Q_FDP0UA U6914 ( .D(n1915), .QTFCLK( ), .Q(numRsts[13]));
Q_MX02 U6915 ( .S(n283), .A0(n2027), .A1(numRsts[13]), .Z(n1915));
Q_FDP0UA U6916 ( .D(n1914), .QTFCLK( ), .Q(numRsts[12]));
Q_MX02 U6917 ( .S(n283), .A0(n2028), .A1(numRsts[12]), .Z(n1914));
Q_FDP0UA U6918 ( .D(n1913), .QTFCLK( ), .Q(numRsts[11]));
Q_MX02 U6919 ( .S(n283), .A0(n2029), .A1(numRsts[11]), .Z(n1913));
Q_FDP0UA U6920 ( .D(n1912), .QTFCLK( ), .Q(numRsts[10]));
Q_MX02 U6921 ( .S(n283), .A0(n2030), .A1(numRsts[10]), .Z(n1912));
Q_FDP0UA U6922 ( .D(n1911), .QTFCLK( ), .Q(numRsts[9]));
Q_MX02 U6923 ( .S(n283), .A0(n2031), .A1(numRsts[9]), .Z(n1911));
Q_FDP0UA U6924 ( .D(n1910), .QTFCLK( ), .Q(numRsts[8]));
Q_MX02 U6925 ( .S(n283), .A0(n2032), .A1(numRsts[8]), .Z(n1910));
Q_FDP0UA U6926 ( .D(n1909), .QTFCLK( ), .Q(numRsts[7]));
Q_MX02 U6927 ( .S(n283), .A0(n2033), .A1(numRsts[7]), .Z(n1909));
Q_FDP0UA U6928 ( .D(n1908), .QTFCLK( ), .Q(numRsts[6]));
Q_MX02 U6929 ( .S(n283), .A0(n2034), .A1(numRsts[6]), .Z(n1908));
Q_FDP0UA U6930 ( .D(n1907), .QTFCLK( ), .Q(numRsts[5]));
Q_MX02 U6931 ( .S(n283), .A0(n2035), .A1(numRsts[5]), .Z(n1907));
Q_FDP0UA U6932 ( .D(n1906), .QTFCLK( ), .Q(numRsts[4]));
Q_MX02 U6933 ( .S(n283), .A0(n2036), .A1(numRsts[4]), .Z(n1906));
Q_FDP0UA U6934 ( .D(n1905), .QTFCLK( ), .Q(numRsts[3]));
Q_MX02 U6935 ( .S(n283), .A0(n2037), .A1(numRsts[3]), .Z(n1905));
Q_FDP0UA U6936 ( .D(n1904), .QTFCLK( ), .Q(numRsts[2]));
Q_MX02 U6937 ( .S(n283), .A0(n2038), .A1(numRsts[2]), .Z(n1904));
Q_FDP0UA U6938 ( .D(n1903), .QTFCLK( ), .Q(numRsts[1]));
Q_MX02 U6939 ( .S(n283), .A0(n2039), .A1(numRsts[1]), .Z(n1903));
Q_FDP0UA U6940 ( .D(n1902), .QTFCLK( ), .Q(numRsts[0]));
Q_MX02 U6941 ( .S(n283), .A0(n2040), .A1(numRsts[0]), .Z(n1902));
Q_FDP0UA U6942 ( .D(n1901), .QTFCLK( ), .Q(ofifoData[767]));
Q_AN02 U6943 ( .A0(n281), .A1(ofifoData[767]), .Z(n1901));
Q_FDP0UA U6944 ( .D(n1900), .QTFCLK( ), .Q(ofifoData[766]));
Q_AN02 U6945 ( .A0(n281), .A1(ofifoData[766]), .Z(n1900));
Q_FDP0UA U6946 ( .D(n1899), .QTFCLK( ), .Q(ofifoData[765]));
Q_AN02 U6947 ( .A0(n281), .A1(ofifoData[765]), .Z(n1899));
Q_FDP0UA U6948 ( .D(n1898), .QTFCLK( ), .Q(ofifoData[764]));
Q_AN02 U6949 ( .A0(n281), .A1(ofifoData[764]), .Z(n1898));
Q_FDP0UA U6950 ( .D(n1897), .QTFCLK( ), .Q(ofifoData[763]));
Q_AN02 U6951 ( .A0(n281), .A1(ofifoData[763]), .Z(n1897));
Q_FDP0UA U6952 ( .D(n1896), .QTFCLK( ), .Q(ofifoData[762]));
Q_AN02 U6953 ( .A0(n281), .A1(ofifoData[762]), .Z(n1896));
Q_FDP0UA U6954 ( .D(n1895), .QTFCLK( ), .Q(ofifoData[761]));
Q_AN02 U6955 ( .A0(n281), .A1(ofifoData[761]), .Z(n1895));
Q_FDP0UA U6956 ( .D(n1894), .QTFCLK( ), .Q(ofifoData[760]));
Q_AN02 U6957 ( .A0(n281), .A1(ofifoData[760]), .Z(n1894));
Q_FDP0UA U6958 ( .D(n1893), .QTFCLK( ), .Q(ofifoData[759]));
Q_AN02 U6959 ( .A0(n281), .A1(ofifoData[759]), .Z(n1893));
Q_FDP0UA U6960 ( .D(n1892), .QTFCLK( ), .Q(ofifoData[758]));
Q_AN02 U6961 ( .A0(n281), .A1(ofifoData[758]), .Z(n1892));
Q_FDP0UA U6962 ( .D(n1891), .QTFCLK( ), .Q(ofifoData[757]));
Q_AN02 U6963 ( .A0(n281), .A1(ofifoData[757]), .Z(n1891));
Q_FDP0UA U6964 ( .D(n1890), .QTFCLK( ), .Q(ofifoData[756]));
Q_AN02 U6965 ( .A0(n281), .A1(ofifoData[756]), .Z(n1890));
Q_FDP0UA U6966 ( .D(n1889), .QTFCLK( ), .Q(ofifoData[755]));
Q_AN02 U6967 ( .A0(n281), .A1(ofifoData[755]), .Z(n1889));
Q_FDP0UA U6968 ( .D(n1888), .QTFCLK( ), .Q(ofifoData[754]));
Q_AN02 U6969 ( .A0(n281), .A1(ofifoData[754]), .Z(n1888));
Q_FDP0UA U6970 ( .D(n1887), .QTFCLK( ), .Q(ofifoData[753]));
Q_AN02 U6971 ( .A0(n281), .A1(ofifoData[753]), .Z(n1887));
Q_FDP0UA U6972 ( .D(n1886), .QTFCLK( ), .Q(ofifoData[752]));
Q_AN02 U6973 ( .A0(n281), .A1(ofifoData[752]), .Z(n1886));
Q_FDP0UA U6974 ( .D(n1885), .QTFCLK( ), .Q(ofifoData[751]));
Q_AN02 U6975 ( .A0(n281), .A1(ofifoData[751]), .Z(n1885));
Q_FDP0UA U6976 ( .D(n1884), .QTFCLK( ), .Q(ofifoData[750]));
Q_AN02 U6977 ( .A0(n281), .A1(ofifoData[750]), .Z(n1884));
Q_FDP0UA U6978 ( .D(n1883), .QTFCLK( ), .Q(ofifoData[749]));
Q_AN02 U6979 ( .A0(n281), .A1(ofifoData[749]), .Z(n1883));
Q_FDP0UA U6980 ( .D(n1882), .QTFCLK( ), .Q(ofifoData[748]));
Q_AN02 U6981 ( .A0(n281), .A1(ofifoData[748]), .Z(n1882));
Q_FDP0UA U6982 ( .D(n1881), .QTFCLK( ), .Q(ofifoData[747]));
Q_AN02 U6983 ( .A0(n281), .A1(ofifoData[747]), .Z(n1881));
Q_FDP0UA U6984 ( .D(n1880), .QTFCLK( ), .Q(ofifoData[746]));
Q_AN02 U6985 ( .A0(n281), .A1(ofifoData[746]), .Z(n1880));
Q_FDP0UA U6986 ( .D(n1879), .QTFCLK( ), .Q(ofifoData[745]));
Q_AN02 U6987 ( .A0(n281), .A1(ofifoData[745]), .Z(n1879));
Q_FDP0UA U6988 ( .D(n1878), .QTFCLK( ), .Q(ofifoData[744]));
Q_AN02 U6989 ( .A0(n281), .A1(ofifoData[744]), .Z(n1878));
Q_FDP0UA U6990 ( .D(n1877), .QTFCLK( ), .Q(ofifoData[743]));
Q_AN02 U6991 ( .A0(n281), .A1(ofifoData[743]), .Z(n1877));
Q_FDP0UA U6992 ( .D(n1876), .QTFCLK( ), .Q(ofifoData[742]));
Q_AN02 U6993 ( .A0(n281), .A1(ofifoData[742]), .Z(n1876));
Q_FDP0UA U6994 ( .D(n1875), .QTFCLK( ), .Q(ofifoData[741]));
Q_AN02 U6995 ( .A0(n281), .A1(ofifoData[741]), .Z(n1875));
Q_FDP0UA U6996 ( .D(n1874), .QTFCLK( ), .Q(ofifoData[740]));
Q_AN02 U6997 ( .A0(n281), .A1(ofifoData[740]), .Z(n1874));
Q_FDP0UA U6998 ( .D(n1873), .QTFCLK( ), .Q(ofifoData[739]));
Q_AN02 U6999 ( .A0(n281), .A1(ofifoData[739]), .Z(n1873));
Q_FDP0UA U7000 ( .D(n1872), .QTFCLK( ), .Q(ofifoData[738]));
Q_AN02 U7001 ( .A0(n281), .A1(ofifoData[738]), .Z(n1872));
Q_FDP0UA U7002 ( .D(n1871), .QTFCLK( ), .Q(ofifoData[737]));
Q_AN02 U7003 ( .A0(n281), .A1(ofifoData[737]), .Z(n1871));
Q_FDP0UA U7004 ( .D(n1870), .QTFCLK( ), .Q(ofifoData[736]));
Q_AN02 U7005 ( .A0(n281), .A1(ofifoData[736]), .Z(n1870));
Q_FDP0UA U7006 ( .D(n1869), .QTFCLK( ), .Q(ofifoData[735]));
Q_AN02 U7007 ( .A0(n281), .A1(ofifoData[735]), .Z(n1869));
Q_FDP0UA U7008 ( .D(n1868), .QTFCLK( ), .Q(ofifoData[734]));
Q_AN02 U7009 ( .A0(n281), .A1(ofifoData[734]), .Z(n1868));
Q_FDP0UA U7010 ( .D(n1867), .QTFCLK( ), .Q(ofifoData[733]));
Q_AN02 U7011 ( .A0(n281), .A1(ofifoData[733]), .Z(n1867));
Q_FDP0UA U7012 ( .D(n1866), .QTFCLK( ), .Q(ofifoData[732]));
Q_AN02 U7013 ( .A0(n281), .A1(ofifoData[732]), .Z(n1866));
Q_FDP0UA U7014 ( .D(n1865), .QTFCLK( ), .Q(ofifoData[731]));
Q_AN02 U7015 ( .A0(n281), .A1(ofifoData[731]), .Z(n1865));
Q_FDP0UA U7016 ( .D(n1864), .QTFCLK( ), .Q(ofifoData[730]));
Q_AN02 U7017 ( .A0(n281), .A1(ofifoData[730]), .Z(n1864));
Q_FDP0UA U7018 ( .D(n1863), .QTFCLK( ), .Q(ofifoData[729]));
Q_AN02 U7019 ( .A0(n281), .A1(ofifoData[729]), .Z(n1863));
Q_FDP0UA U7020 ( .D(n1862), .QTFCLK( ), .Q(ofifoData[728]));
Q_AN02 U7021 ( .A0(n281), .A1(ofifoData[728]), .Z(n1862));
Q_FDP0UA U7022 ( .D(n1861), .QTFCLK( ), .Q(ofifoData[727]));
Q_AN02 U7023 ( .A0(n281), .A1(ofifoData[727]), .Z(n1861));
Q_FDP0UA U7024 ( .D(n1860), .QTFCLK( ), .Q(ofifoData[726]));
Q_AN02 U7025 ( .A0(n281), .A1(ofifoData[726]), .Z(n1860));
Q_FDP0UA U7026 ( .D(n1859), .QTFCLK( ), .Q(ofifoData[725]));
Q_AN02 U7027 ( .A0(n281), .A1(ofifoData[725]), .Z(n1859));
Q_FDP0UA U7028 ( .D(n1858), .QTFCLK( ), .Q(ofifoData[724]));
Q_AN02 U7029 ( .A0(n281), .A1(ofifoData[724]), .Z(n1858));
Q_FDP0UA U7030 ( .D(n1857), .QTFCLK( ), .Q(ofifoData[723]));
Q_AN02 U7031 ( .A0(n281), .A1(ofifoData[723]), .Z(n1857));
Q_FDP0UA U7032 ( .D(n1856), .QTFCLK( ), .Q(ofifoData[722]));
Q_AN02 U7033 ( .A0(n281), .A1(ofifoData[722]), .Z(n1856));
Q_FDP0UA U7034 ( .D(n1855), .QTFCLK( ), .Q(ofifoData[721]));
Q_AN02 U7035 ( .A0(n281), .A1(ofifoData[721]), .Z(n1855));
Q_FDP0UA U7036 ( .D(n1854), .QTFCLK( ), .Q(ofifoData[720]));
Q_AN02 U7037 ( .A0(n281), .A1(ofifoData[720]), .Z(n1854));
Q_FDP0UA U7038 ( .D(n1853), .QTFCLK( ), .Q(ofifoData[719]));
Q_AN02 U7039 ( .A0(n281), .A1(ofifoData[719]), .Z(n1853));
Q_FDP0UA U7040 ( .D(n1852), .QTFCLK( ), .Q(ofifoData[718]));
Q_AN02 U7041 ( .A0(n281), .A1(ofifoData[718]), .Z(n1852));
Q_FDP0UA U7042 ( .D(n1851), .QTFCLK( ), .Q(ofifoData[717]));
Q_AN02 U7043 ( .A0(n281), .A1(ofifoData[717]), .Z(n1851));
Q_FDP0UA U7044 ( .D(n1850), .QTFCLK( ), .Q(ofifoData[716]));
Q_AN02 U7045 ( .A0(n281), .A1(ofifoData[716]), .Z(n1850));
Q_FDP0UA U7046 ( .D(n1849), .QTFCLK( ), .Q(ofifoData[715]));
Q_AN02 U7047 ( .A0(n281), .A1(ofifoData[715]), .Z(n1849));
Q_FDP0UA U7048 ( .D(n1848), .QTFCLK( ), .Q(ofifoData[714]));
Q_AN02 U7049 ( .A0(n281), .A1(ofifoData[714]), .Z(n1848));
Q_FDP0UA U7050 ( .D(n1847), .QTFCLK( ), .Q(ofifoData[713]));
Q_AN02 U7051 ( .A0(n281), .A1(ofifoData[713]), .Z(n1847));
Q_FDP0UA U7052 ( .D(n1846), .QTFCLK( ), .Q(ofifoData[712]));
Q_AN02 U7053 ( .A0(n281), .A1(ofifoData[712]), .Z(n1846));
Q_FDP0UA U7054 ( .D(n1845), .QTFCLK( ), .Q(ofifoData[711]));
Q_AN02 U7055 ( .A0(n281), .A1(ofifoData[711]), .Z(n1845));
Q_FDP0UA U7056 ( .D(n1844), .QTFCLK( ), .Q(ofifoData[710]));
Q_AN02 U7057 ( .A0(n281), .A1(ofifoData[710]), .Z(n1844));
Q_FDP0UA U7058 ( .D(n1843), .QTFCLK( ), .Q(ofifoData[709]));
Q_AN02 U7059 ( .A0(n281), .A1(ofifoData[709]), .Z(n1843));
Q_FDP0UA U7060 ( .D(n1842), .QTFCLK( ), .Q(ofifoData[708]));
Q_AN02 U7061 ( .A0(n281), .A1(ofifoData[708]), .Z(n1842));
Q_FDP0UA U7062 ( .D(n1841), .QTFCLK( ), .Q(ofifoData[707]));
Q_AN02 U7063 ( .A0(n281), .A1(ofifoData[707]), .Z(n1841));
Q_FDP0UA U7064 ( .D(n1840), .QTFCLK( ), .Q(ofifoData[706]));
Q_AN02 U7065 ( .A0(n281), .A1(ofifoData[706]), .Z(n1840));
Q_FDP0UA U7066 ( .D(n1839), .QTFCLK( ), .Q(ofifoData[705]));
Q_AN02 U7067 ( .A0(n281), .A1(ofifoData[705]), .Z(n1839));
Q_FDP0UA U7068 ( .D(n1838), .QTFCLK( ), .Q(ofifoData[704]));
Q_AN02 U7069 ( .A0(n281), .A1(ofifoData[704]), .Z(n1838));
Q_FDP0UA U7070 ( .D(n1837), .QTFCLK( ), .Q(ofifoData[703]));
Q_MX02 U7071 ( .S(n281), .A0(n2041), .A1(ofifoData[703]), .Z(n1837));
Q_FDP0UA U7072 ( .D(n1836), .QTFCLK( ), .Q(ofifoData[702]));
Q_MX02 U7073 ( .S(n281), .A0(n2042), .A1(ofifoData[702]), .Z(n1836));
Q_FDP0UA U7074 ( .D(n1835), .QTFCLK( ), .Q(ofifoData[701]));
Q_MX02 U7075 ( .S(n281), .A0(n2043), .A1(ofifoData[701]), .Z(n1835));
Q_FDP0UA U7076 ( .D(n1834), .QTFCLK( ), .Q(ofifoData[700]));
Q_MX02 U7077 ( .S(n281), .A0(n2044), .A1(ofifoData[700]), .Z(n1834));
Q_FDP0UA U7078 ( .D(n1833), .QTFCLK( ), .Q(ofifoData[699]));
Q_MX02 U7079 ( .S(n281), .A0(n2045), .A1(ofifoData[699]), .Z(n1833));
Q_FDP0UA U7080 ( .D(n1832), .QTFCLK( ), .Q(ofifoData[698]));
Q_MX02 U7081 ( .S(n281), .A0(n2046), .A1(ofifoData[698]), .Z(n1832));
Q_FDP0UA U7082 ( .D(n1831), .QTFCLK( ), .Q(ofifoData[697]));
Q_MX02 U7083 ( .S(n281), .A0(n2047), .A1(ofifoData[697]), .Z(n1831));
Q_FDP0UA U7084 ( .D(n1830), .QTFCLK( ), .Q(ofifoData[696]));
Q_MX02 U7085 ( .S(n281), .A0(n2048), .A1(ofifoData[696]), .Z(n1830));
Q_FDP0UA U7086 ( .D(n1829), .QTFCLK( ), .Q(ofifoData[695]));
Q_MX02 U7087 ( .S(n281), .A0(n2049), .A1(ofifoData[695]), .Z(n1829));
Q_FDP0UA U7088 ( .D(n1828), .QTFCLK( ), .Q(ofifoData[694]));
Q_MX02 U7089 ( .S(n281), .A0(n2050), .A1(ofifoData[694]), .Z(n1828));
Q_FDP0UA U7090 ( .D(n1827), .QTFCLK( ), .Q(ofifoData[693]));
Q_MX02 U7091 ( .S(n281), .A0(n2051), .A1(ofifoData[693]), .Z(n1827));
Q_FDP0UA U7092 ( .D(n1826), .QTFCLK( ), .Q(ofifoData[692]));
Q_MX02 U7093 ( .S(n281), .A0(n2052), .A1(ofifoData[692]), .Z(n1826));
Q_FDP0UA U7094 ( .D(n1825), .QTFCLK( ), .Q(ofifoData[691]));
Q_MX02 U7095 ( .S(n281), .A0(n2053), .A1(ofifoData[691]), .Z(n1825));
Q_FDP0UA U7096 ( .D(n1824), .QTFCLK( ), .Q(ofifoData[690]));
Q_MX02 U7097 ( .S(n281), .A0(n2054), .A1(ofifoData[690]), .Z(n1824));
Q_FDP0UA U7098 ( .D(n1823), .QTFCLK( ), .Q(ofifoData[689]));
Q_MX02 U7099 ( .S(n281), .A0(n2055), .A1(ofifoData[689]), .Z(n1823));
Q_FDP0UA U7100 ( .D(n1822), .QTFCLK( ), .Q(ofifoData[688]));
Q_MX02 U7101 ( .S(n281), .A0(n2056), .A1(ofifoData[688]), .Z(n1822));
Q_FDP0UA U7102 ( .D(n1821), .QTFCLK( ), .Q(ofifoData[687]));
Q_MX02 U7103 ( .S(n281), .A0(n2057), .A1(ofifoData[687]), .Z(n1821));
Q_FDP0UA U7104 ( .D(n1820), .QTFCLK( ), .Q(ofifoData[686]));
Q_MX02 U7105 ( .S(n281), .A0(n2058), .A1(ofifoData[686]), .Z(n1820));
Q_FDP0UA U7106 ( .D(n1819), .QTFCLK( ), .Q(ofifoData[685]));
Q_MX02 U7107 ( .S(n281), .A0(n2059), .A1(ofifoData[685]), .Z(n1819));
Q_FDP0UA U7108 ( .D(n1818), .QTFCLK( ), .Q(ofifoData[684]));
Q_MX02 U7109 ( .S(n281), .A0(n2060), .A1(ofifoData[684]), .Z(n1818));
Q_FDP0UA U7110 ( .D(n1817), .QTFCLK( ), .Q(ofifoData[683]));
Q_MX02 U7111 ( .S(n281), .A0(n2061), .A1(ofifoData[683]), .Z(n1817));
Q_FDP0UA U7112 ( .D(n1816), .QTFCLK( ), .Q(ofifoData[682]));
Q_MX02 U7113 ( .S(n281), .A0(n2062), .A1(ofifoData[682]), .Z(n1816));
Q_FDP0UA U7114 ( .D(n1815), .QTFCLK( ), .Q(ofifoData[681]));
Q_MX02 U7115 ( .S(n281), .A0(n2063), .A1(ofifoData[681]), .Z(n1815));
Q_FDP0UA U7116 ( .D(n1814), .QTFCLK( ), .Q(ofifoData[680]));
Q_MX02 U7117 ( .S(n281), .A0(n2064), .A1(ofifoData[680]), .Z(n1814));
Q_FDP0UA U7118 ( .D(n1813), .QTFCLK( ), .Q(ofifoData[679]));
Q_MX02 U7119 ( .S(n281), .A0(n2065), .A1(ofifoData[679]), .Z(n1813));
Q_FDP0UA U7120 ( .D(n1812), .QTFCLK( ), .Q(ofifoData[678]));
Q_MX02 U7121 ( .S(n281), .A0(n2066), .A1(ofifoData[678]), .Z(n1812));
Q_FDP0UA U7122 ( .D(n1811), .QTFCLK( ), .Q(ofifoData[677]));
Q_MX02 U7123 ( .S(n281), .A0(n2067), .A1(ofifoData[677]), .Z(n1811));
Q_FDP0UA U7124 ( .D(n1810), .QTFCLK( ), .Q(ofifoData[676]));
Q_MX02 U7125 ( .S(n281), .A0(n2068), .A1(ofifoData[676]), .Z(n1810));
Q_FDP0UA U7126 ( .D(n1809), .QTFCLK( ), .Q(ofifoData[675]));
Q_MX02 U7127 ( .S(n281), .A0(n2069), .A1(ofifoData[675]), .Z(n1809));
Q_FDP0UA U7128 ( .D(n1808), .QTFCLK( ), .Q(ofifoData[674]));
Q_MX02 U7129 ( .S(n281), .A0(n2070), .A1(ofifoData[674]), .Z(n1808));
Q_FDP0UA U7130 ( .D(n1807), .QTFCLK( ), .Q(ofifoData[673]));
Q_MX02 U7131 ( .S(n281), .A0(n2071), .A1(ofifoData[673]), .Z(n1807));
Q_FDP0UA U7132 ( .D(n1806), .QTFCLK( ), .Q(ofifoData[672]));
Q_MX02 U7133 ( .S(n281), .A0(n2072), .A1(ofifoData[672]), .Z(n1806));
Q_FDP0UA U7134 ( .D(n1805), .QTFCLK( ), .Q(ofifoData[671]));
Q_MX02 U7135 ( .S(n281), .A0(n2073), .A1(ofifoData[671]), .Z(n1805));
Q_FDP0UA U7136 ( .D(n1804), .QTFCLK( ), .Q(ofifoData[670]));
Q_MX02 U7137 ( .S(n281), .A0(n2074), .A1(ofifoData[670]), .Z(n1804));
Q_FDP0UA U7138 ( .D(n1803), .QTFCLK( ), .Q(ofifoData[669]));
Q_MX02 U7139 ( .S(n281), .A0(n2075), .A1(ofifoData[669]), .Z(n1803));
Q_FDP0UA U7140 ( .D(n1802), .QTFCLK( ), .Q(ofifoData[668]));
Q_MX02 U7141 ( .S(n281), .A0(n2076), .A1(ofifoData[668]), .Z(n1802));
Q_FDP0UA U7142 ( .D(n1801), .QTFCLK( ), .Q(ofifoData[667]));
Q_MX02 U7143 ( .S(n281), .A0(n2077), .A1(ofifoData[667]), .Z(n1801));
Q_FDP0UA U7144 ( .D(n1800), .QTFCLK( ), .Q(ofifoData[666]));
Q_MX02 U7145 ( .S(n281), .A0(n2078), .A1(ofifoData[666]), .Z(n1800));
Q_FDP0UA U7146 ( .D(n1799), .QTFCLK( ), .Q(ofifoData[665]));
Q_MX02 U7147 ( .S(n281), .A0(n2079), .A1(ofifoData[665]), .Z(n1799));
Q_FDP0UA U7148 ( .D(n1798), .QTFCLK( ), .Q(ofifoData[664]));
Q_MX02 U7149 ( .S(n281), .A0(n2080), .A1(ofifoData[664]), .Z(n1798));
Q_FDP0UA U7150 ( .D(n1797), .QTFCLK( ), .Q(ofifoData[663]));
Q_MX02 U7151 ( .S(n281), .A0(n2081), .A1(ofifoData[663]), .Z(n1797));
Q_FDP0UA U7152 ( .D(n1796), .QTFCLK( ), .Q(ofifoData[662]));
Q_MX02 U7153 ( .S(n281), .A0(n2082), .A1(ofifoData[662]), .Z(n1796));
Q_FDP0UA U7154 ( .D(n1795), .QTFCLK( ), .Q(ofifoData[661]));
Q_MX02 U7155 ( .S(n281), .A0(n2083), .A1(ofifoData[661]), .Z(n1795));
Q_FDP0UA U7156 ( .D(n1794), .QTFCLK( ), .Q(ofifoData[660]));
Q_MX02 U7157 ( .S(n281), .A0(n2084), .A1(ofifoData[660]), .Z(n1794));
Q_FDP0UA U7158 ( .D(n1793), .QTFCLK( ), .Q(ofifoData[659]));
Q_MX02 U7159 ( .S(n281), .A0(n2085), .A1(ofifoData[659]), .Z(n1793));
Q_FDP0UA U7160 ( .D(n1792), .QTFCLK( ), .Q(ofifoData[658]));
Q_MX02 U7161 ( .S(n281), .A0(n2086), .A1(ofifoData[658]), .Z(n1792));
Q_FDP0UA U7162 ( .D(n1791), .QTFCLK( ), .Q(ofifoData[657]));
Q_MX02 U7163 ( .S(n281), .A0(n2087), .A1(ofifoData[657]), .Z(n1791));
Q_FDP0UA U7164 ( .D(n1790), .QTFCLK( ), .Q(ofifoData[656]));
Q_MX02 U7165 ( .S(n281), .A0(n2088), .A1(ofifoData[656]), .Z(n1790));
Q_FDP0UA U7166 ( .D(n1789), .QTFCLK( ), .Q(ofifoData[655]));
Q_MX02 U7167 ( .S(n281), .A0(n2089), .A1(ofifoData[655]), .Z(n1789));
Q_FDP0UA U7168 ( .D(n1788), .QTFCLK( ), .Q(ofifoData[654]));
Q_MX02 U7169 ( .S(n281), .A0(n2090), .A1(ofifoData[654]), .Z(n1788));
Q_FDP0UA U7170 ( .D(n1787), .QTFCLK( ), .Q(ofifoData[653]));
Q_MX02 U7171 ( .S(n281), .A0(n2091), .A1(ofifoData[653]), .Z(n1787));
Q_FDP0UA U7172 ( .D(n1786), .QTFCLK( ), .Q(ofifoData[652]));
Q_MX02 U7173 ( .S(n281), .A0(n2092), .A1(ofifoData[652]), .Z(n1786));
Q_FDP0UA U7174 ( .D(n1785), .QTFCLK( ), .Q(ofifoData[651]));
Q_MX02 U7175 ( .S(n281), .A0(n2093), .A1(ofifoData[651]), .Z(n1785));
Q_FDP0UA U7176 ( .D(n1784), .QTFCLK( ), .Q(ofifoData[650]));
Q_MX02 U7177 ( .S(n281), .A0(n2094), .A1(ofifoData[650]), .Z(n1784));
Q_FDP0UA U7178 ( .D(n1783), .QTFCLK( ), .Q(ofifoData[649]));
Q_MX02 U7179 ( .S(n281), .A0(n2095), .A1(ofifoData[649]), .Z(n1783));
Q_FDP0UA U7180 ( .D(n1782), .QTFCLK( ), .Q(ofifoData[648]));
Q_MX02 U7181 ( .S(n281), .A0(n2096), .A1(ofifoData[648]), .Z(n1782));
Q_FDP0UA U7182 ( .D(n1781), .QTFCLK( ), .Q(ofifoData[647]));
Q_MX02 U7183 ( .S(n281), .A0(n2097), .A1(ofifoData[647]), .Z(n1781));
Q_FDP0UA U7184 ( .D(n1780), .QTFCLK( ), .Q(ofifoData[646]));
Q_MX02 U7185 ( .S(n281), .A0(n2098), .A1(ofifoData[646]), .Z(n1780));
Q_FDP0UA U7186 ( .D(n1779), .QTFCLK( ), .Q(ofifoData[645]));
Q_MX02 U7187 ( .S(n281), .A0(n2099), .A1(ofifoData[645]), .Z(n1779));
Q_FDP0UA U7188 ( .D(n1778), .QTFCLK( ), .Q(ofifoData[644]));
Q_MX02 U7189 ( .S(n281), .A0(n2100), .A1(ofifoData[644]), .Z(n1778));
Q_FDP0UA U7190 ( .D(n1777), .QTFCLK( ), .Q(ofifoData[643]));
Q_MX02 U7191 ( .S(n281), .A0(n2101), .A1(ofifoData[643]), .Z(n1777));
Q_FDP0UA U7192 ( .D(n1776), .QTFCLK( ), .Q(ofifoData[642]));
Q_MX02 U7193 ( .S(n281), .A0(n2102), .A1(ofifoData[642]), .Z(n1776));
Q_FDP0UA U7194 ( .D(n1775), .QTFCLK( ), .Q(ofifoData[641]));
Q_MX02 U7195 ( .S(n281), .A0(n2103), .A1(ofifoData[641]), .Z(n1775));
Q_FDP0UA U7196 ( .D(n1774), .QTFCLK( ), .Q(ofifoData[640]));
Q_MX02 U7197 ( .S(n281), .A0(n2104), .A1(ofifoData[640]), .Z(n1774));
Q_FDP0UA U7198 ( .D(n1773), .QTFCLK( ), .Q(ofifoData[639]));
Q_MX02 U7199 ( .S(n281), .A0(n2105), .A1(ofifoData[639]), .Z(n1773));
Q_FDP0UA U7200 ( .D(n1772), .QTFCLK( ), .Q(ofifoData[638]));
Q_MX02 U7201 ( .S(n281), .A0(n2106), .A1(ofifoData[638]), .Z(n1772));
Q_FDP0UA U7202 ( .D(n1771), .QTFCLK( ), .Q(ofifoData[637]));
Q_MX02 U7203 ( .S(n281), .A0(n2107), .A1(ofifoData[637]), .Z(n1771));
Q_FDP0UA U7204 ( .D(n1770), .QTFCLK( ), .Q(ofifoData[636]));
Q_MX02 U7205 ( .S(n281), .A0(n2108), .A1(ofifoData[636]), .Z(n1770));
Q_FDP0UA U7206 ( .D(n1769), .QTFCLK( ), .Q(ofifoData[635]));
Q_MX02 U7207 ( .S(n281), .A0(n2109), .A1(ofifoData[635]), .Z(n1769));
Q_FDP0UA U7208 ( .D(n1768), .QTFCLK( ), .Q(ofifoData[634]));
Q_MX02 U7209 ( .S(n281), .A0(n2110), .A1(ofifoData[634]), .Z(n1768));
Q_FDP0UA U7210 ( .D(n1767), .QTFCLK( ), .Q(ofifoData[633]));
Q_MX02 U7211 ( .S(n281), .A0(n2111), .A1(ofifoData[633]), .Z(n1767));
Q_FDP0UA U7212 ( .D(n1766), .QTFCLK( ), .Q(ofifoData[632]));
Q_MX02 U7213 ( .S(n281), .A0(n2112), .A1(ofifoData[632]), .Z(n1766));
Q_FDP0UA U7214 ( .D(n1765), .QTFCLK( ), .Q(ofifoData[631]));
Q_MX02 U7215 ( .S(n281), .A0(n2113), .A1(ofifoData[631]), .Z(n1765));
Q_FDP0UA U7216 ( .D(n1764), .QTFCLK( ), .Q(ofifoData[630]));
Q_MX02 U7217 ( .S(n281), .A0(n2114), .A1(ofifoData[630]), .Z(n1764));
Q_FDP0UA U7218 ( .D(n1763), .QTFCLK( ), .Q(ofifoData[629]));
Q_MX02 U7219 ( .S(n281), .A0(n2115), .A1(ofifoData[629]), .Z(n1763));
Q_FDP0UA U7220 ( .D(n1762), .QTFCLK( ), .Q(ofifoData[628]));
Q_MX02 U7221 ( .S(n281), .A0(n2116), .A1(ofifoData[628]), .Z(n1762));
Q_FDP0UA U7222 ( .D(n1761), .QTFCLK( ), .Q(ofifoData[627]));
Q_MX02 U7223 ( .S(n281), .A0(n2117), .A1(ofifoData[627]), .Z(n1761));
Q_FDP0UA U7224 ( .D(n1760), .QTFCLK( ), .Q(ofifoData[626]));
Q_MX02 U7225 ( .S(n281), .A0(n2118), .A1(ofifoData[626]), .Z(n1760));
Q_FDP0UA U7226 ( .D(n1759), .QTFCLK( ), .Q(ofifoData[625]));
Q_MX02 U7227 ( .S(n281), .A0(n2119), .A1(ofifoData[625]), .Z(n1759));
Q_FDP0UA U7228 ( .D(n1758), .QTFCLK( ), .Q(ofifoData[624]));
Q_MX02 U7229 ( .S(n281), .A0(n2120), .A1(ofifoData[624]), .Z(n1758));
Q_FDP0UA U7230 ( .D(n1757), .QTFCLK( ), .Q(ofifoData[623]));
Q_MX02 U7231 ( .S(n281), .A0(n2121), .A1(ofifoData[623]), .Z(n1757));
Q_FDP0UA U7232 ( .D(n1756), .QTFCLK( ), .Q(ofifoData[622]));
Q_MX02 U7233 ( .S(n281), .A0(n2122), .A1(ofifoData[622]), .Z(n1756));
Q_FDP0UA U7234 ( .D(n1755), .QTFCLK( ), .Q(ofifoData[621]));
Q_MX02 U7235 ( .S(n281), .A0(n2123), .A1(ofifoData[621]), .Z(n1755));
Q_FDP0UA U7236 ( .D(n1754), .QTFCLK( ), .Q(ofifoData[620]));
Q_MX02 U7237 ( .S(n281), .A0(n2124), .A1(ofifoData[620]), .Z(n1754));
Q_FDP0UA U7238 ( .D(n1753), .QTFCLK( ), .Q(ofifoData[619]));
Q_MX02 U7239 ( .S(n281), .A0(n2125), .A1(ofifoData[619]), .Z(n1753));
Q_FDP0UA U7240 ( .D(n1752), .QTFCLK( ), .Q(ofifoData[618]));
Q_MX02 U7241 ( .S(n281), .A0(n2126), .A1(ofifoData[618]), .Z(n1752));
Q_FDP0UA U7242 ( .D(n1751), .QTFCLK( ), .Q(ofifoData[617]));
Q_MX02 U7243 ( .S(n281), .A0(n2127), .A1(ofifoData[617]), .Z(n1751));
Q_FDP0UA U7244 ( .D(n1750), .QTFCLK( ), .Q(ofifoData[616]));
Q_MX02 U7245 ( .S(n281), .A0(n2128), .A1(ofifoData[616]), .Z(n1750));
Q_FDP0UA U7246 ( .D(n1749), .QTFCLK( ), .Q(ofifoData[615]));
Q_MX02 U7247 ( .S(n281), .A0(n2129), .A1(ofifoData[615]), .Z(n1749));
Q_FDP0UA U7248 ( .D(n1748), .QTFCLK( ), .Q(ofifoData[614]));
Q_MX02 U7249 ( .S(n281), .A0(n2130), .A1(ofifoData[614]), .Z(n1748));
Q_FDP0UA U7250 ( .D(n1747), .QTFCLK( ), .Q(ofifoData[613]));
Q_MX02 U7251 ( .S(n281), .A0(n2131), .A1(ofifoData[613]), .Z(n1747));
Q_FDP0UA U7252 ( .D(n1746), .QTFCLK( ), .Q(ofifoData[612]));
Q_MX02 U7253 ( .S(n281), .A0(n2132), .A1(ofifoData[612]), .Z(n1746));
Q_FDP0UA U7254 ( .D(n1745), .QTFCLK( ), .Q(ofifoData[611]));
Q_MX02 U7255 ( .S(n281), .A0(n2133), .A1(ofifoData[611]), .Z(n1745));
Q_FDP0UA U7256 ( .D(n1744), .QTFCLK( ), .Q(ofifoData[610]));
Q_MX02 U7257 ( .S(n281), .A0(n2134), .A1(ofifoData[610]), .Z(n1744));
Q_FDP0UA U7258 ( .D(n1743), .QTFCLK( ), .Q(ofifoData[609]));
Q_MX02 U7259 ( .S(n281), .A0(n2135), .A1(ofifoData[609]), .Z(n1743));
Q_FDP0UA U7260 ( .D(n1742), .QTFCLK( ), .Q(ofifoData[608]));
Q_MX02 U7261 ( .S(n281), .A0(n2136), .A1(ofifoData[608]), .Z(n1742));
Q_FDP0UA U7262 ( .D(n1741), .QTFCLK( ), .Q(ofifoData[607]));
Q_MX02 U7263 ( .S(n281), .A0(n2137), .A1(ofifoData[607]), .Z(n1741));
Q_FDP0UA U7264 ( .D(n1740), .QTFCLK( ), .Q(ofifoData[606]));
Q_MX02 U7265 ( .S(n281), .A0(n2138), .A1(ofifoData[606]), .Z(n1740));
Q_FDP0UA U7266 ( .D(n1739), .QTFCLK( ), .Q(ofifoData[605]));
Q_MX02 U7267 ( .S(n281), .A0(n2139), .A1(ofifoData[605]), .Z(n1739));
Q_FDP0UA U7268 ( .D(n1738), .QTFCLK( ), .Q(ofifoData[604]));
Q_MX02 U7269 ( .S(n281), .A0(n2140), .A1(ofifoData[604]), .Z(n1738));
Q_FDP0UA U7270 ( .D(n1737), .QTFCLK( ), .Q(ofifoData[603]));
Q_MX02 U7271 ( .S(n281), .A0(n2141), .A1(ofifoData[603]), .Z(n1737));
Q_FDP0UA U7272 ( .D(n1736), .QTFCLK( ), .Q(ofifoData[602]));
Q_MX02 U7273 ( .S(n281), .A0(n2142), .A1(ofifoData[602]), .Z(n1736));
Q_FDP0UA U7274 ( .D(n1735), .QTFCLK( ), .Q(ofifoData[601]));
Q_MX02 U7275 ( .S(n281), .A0(n2143), .A1(ofifoData[601]), .Z(n1735));
Q_FDP0UA U7276 ( .D(n1734), .QTFCLK( ), .Q(ofifoData[600]));
Q_MX02 U7277 ( .S(n281), .A0(n2144), .A1(ofifoData[600]), .Z(n1734));
Q_FDP0UA U7278 ( .D(n1733), .QTFCLK( ), .Q(ofifoData[599]));
Q_MX02 U7279 ( .S(n281), .A0(n2145), .A1(ofifoData[599]), .Z(n1733));
Q_FDP0UA U7280 ( .D(n1732), .QTFCLK( ), .Q(ofifoData[598]));
Q_MX02 U7281 ( .S(n281), .A0(n2146), .A1(ofifoData[598]), .Z(n1732));
Q_FDP0UA U7282 ( .D(n1731), .QTFCLK( ), .Q(ofifoData[597]));
Q_MX02 U7283 ( .S(n281), .A0(n2147), .A1(ofifoData[597]), .Z(n1731));
Q_FDP0UA U7284 ( .D(n1730), .QTFCLK( ), .Q(ofifoData[596]));
Q_MX02 U7285 ( .S(n281), .A0(n2148), .A1(ofifoData[596]), .Z(n1730));
Q_FDP0UA U7286 ( .D(n1729), .QTFCLK( ), .Q(ofifoData[595]));
Q_MX02 U7287 ( .S(n281), .A0(n2149), .A1(ofifoData[595]), .Z(n1729));
Q_FDP0UA U7288 ( .D(n1728), .QTFCLK( ), .Q(ofifoData[594]));
Q_MX02 U7289 ( .S(n281), .A0(n2150), .A1(ofifoData[594]), .Z(n1728));
Q_FDP0UA U7290 ( .D(n1727), .QTFCLK( ), .Q(ofifoData[593]));
Q_MX02 U7291 ( .S(n281), .A0(n2151), .A1(ofifoData[593]), .Z(n1727));
Q_FDP0UA U7292 ( .D(n1726), .QTFCLK( ), .Q(ofifoData[592]));
Q_MX02 U7293 ( .S(n281), .A0(n2152), .A1(ofifoData[592]), .Z(n1726));
Q_FDP0UA U7294 ( .D(n1725), .QTFCLK( ), .Q(ofifoData[591]));
Q_MX02 U7295 ( .S(n281), .A0(n2153), .A1(ofifoData[591]), .Z(n1725));
Q_FDP0UA U7296 ( .D(n1724), .QTFCLK( ), .Q(ofifoData[590]));
Q_MX02 U7297 ( .S(n281), .A0(n2154), .A1(ofifoData[590]), .Z(n1724));
Q_FDP0UA U7298 ( .D(n1723), .QTFCLK( ), .Q(ofifoData[589]));
Q_MX02 U7299 ( .S(n281), .A0(n2155), .A1(ofifoData[589]), .Z(n1723));
Q_FDP0UA U7300 ( .D(n1722), .QTFCLK( ), .Q(ofifoData[588]));
Q_MX02 U7301 ( .S(n281), .A0(n2156), .A1(ofifoData[588]), .Z(n1722));
Q_FDP0UA U7302 ( .D(n1721), .QTFCLK( ), .Q(ofifoData[587]));
Q_MX02 U7303 ( .S(n281), .A0(n2157), .A1(ofifoData[587]), .Z(n1721));
Q_FDP0UA U7304 ( .D(n1720), .QTFCLK( ), .Q(ofifoData[586]));
Q_MX02 U7305 ( .S(n281), .A0(n2158), .A1(ofifoData[586]), .Z(n1720));
Q_FDP0UA U7306 ( .D(n1719), .QTFCLK( ), .Q(ofifoData[585]));
Q_MX02 U7307 ( .S(n281), .A0(n2159), .A1(ofifoData[585]), .Z(n1719));
Q_FDP0UA U7308 ( .D(n1718), .QTFCLK( ), .Q(ofifoData[584]));
Q_MX02 U7309 ( .S(n281), .A0(n2160), .A1(ofifoData[584]), .Z(n1718));
Q_FDP0UA U7310 ( .D(n1717), .QTFCLK( ), .Q(ofifoData[583]));
Q_MX02 U7311 ( .S(n281), .A0(n2161), .A1(ofifoData[583]), .Z(n1717));
Q_FDP0UA U7312 ( .D(n1716), .QTFCLK( ), .Q(ofifoData[582]));
Q_MX02 U7313 ( .S(n281), .A0(n2162), .A1(ofifoData[582]), .Z(n1716));
Q_FDP0UA U7314 ( .D(n1715), .QTFCLK( ), .Q(ofifoData[581]));
Q_MX02 U7315 ( .S(n281), .A0(n2163), .A1(ofifoData[581]), .Z(n1715));
Q_FDP0UA U7316 ( .D(n1714), .QTFCLK( ), .Q(ofifoData[580]));
Q_MX02 U7317 ( .S(n281), .A0(n2164), .A1(ofifoData[580]), .Z(n1714));
Q_FDP0UA U7318 ( .D(n1713), .QTFCLK( ), .Q(ofifoData[579]));
Q_MX02 U7319 ( .S(n281), .A0(n2165), .A1(ofifoData[579]), .Z(n1713));
Q_FDP0UA U7320 ( .D(n1712), .QTFCLK( ), .Q(ofifoData[578]));
Q_MX02 U7321 ( .S(n281), .A0(n2166), .A1(ofifoData[578]), .Z(n1712));
Q_FDP0UA U7322 ( .D(n1711), .QTFCLK( ), .Q(ofifoData[577]));
Q_MX02 U7323 ( .S(n281), .A0(n2167), .A1(ofifoData[577]), .Z(n1711));
Q_FDP0UA U7324 ( .D(n1710), .QTFCLK( ), .Q(ofifoData[576]));
Q_MX02 U7325 ( .S(n281), .A0(n2168), .A1(ofifoData[576]), .Z(n1710));
Q_FDP0UA U7326 ( .D(n1709), .QTFCLK( ), .Q(ofifoData[575]));
Q_MX02 U7327 ( .S(n281), .A0(n2169), .A1(ofifoData[575]), .Z(n1709));
Q_FDP0UA U7328 ( .D(n1708), .QTFCLK( ), .Q(ofifoData[574]));
Q_MX02 U7329 ( .S(n281), .A0(n2170), .A1(ofifoData[574]), .Z(n1708));
Q_FDP0UA U7330 ( .D(n1707), .QTFCLK( ), .Q(ofifoData[573]));
Q_MX02 U7331 ( .S(n281), .A0(n2171), .A1(ofifoData[573]), .Z(n1707));
Q_FDP0UA U7332 ( .D(n1706), .QTFCLK( ), .Q(ofifoData[572]));
Q_MX02 U7333 ( .S(n281), .A0(n2172), .A1(ofifoData[572]), .Z(n1706));
Q_FDP0UA U7334 ( .D(n1705), .QTFCLK( ), .Q(ofifoData[571]));
Q_MX02 U7335 ( .S(n281), .A0(n2173), .A1(ofifoData[571]), .Z(n1705));
Q_FDP0UA U7336 ( .D(n1704), .QTFCLK( ), .Q(ofifoData[570]));
Q_MX02 U7337 ( .S(n281), .A0(n2174), .A1(ofifoData[570]), .Z(n1704));
Q_FDP0UA U7338 ( .D(n1703), .QTFCLK( ), .Q(ofifoData[569]));
Q_MX02 U7339 ( .S(n281), .A0(n2175), .A1(ofifoData[569]), .Z(n1703));
Q_FDP0UA U7340 ( .D(n1702), .QTFCLK( ), .Q(ofifoData[568]));
Q_MX02 U7341 ( .S(n281), .A0(n2176), .A1(ofifoData[568]), .Z(n1702));
Q_FDP0UA U7342 ( .D(n1701), .QTFCLK( ), .Q(ofifoData[567]));
Q_MX02 U7343 ( .S(n281), .A0(n2177), .A1(ofifoData[567]), .Z(n1701));
Q_FDP0UA U7344 ( .D(n1700), .QTFCLK( ), .Q(ofifoData[566]));
Q_MX02 U7345 ( .S(n281), .A0(n2178), .A1(ofifoData[566]), .Z(n1700));
Q_FDP0UA U7346 ( .D(n1699), .QTFCLK( ), .Q(ofifoData[565]));
Q_MX02 U7347 ( .S(n281), .A0(n2179), .A1(ofifoData[565]), .Z(n1699));
Q_FDP0UA U7348 ( .D(n1698), .QTFCLK( ), .Q(ofifoData[564]));
Q_MX02 U7349 ( .S(n281), .A0(n2180), .A1(ofifoData[564]), .Z(n1698));
Q_FDP0UA U7350 ( .D(n1697), .QTFCLK( ), .Q(ofifoData[563]));
Q_MX02 U7351 ( .S(n281), .A0(n2181), .A1(ofifoData[563]), .Z(n1697));
Q_FDP0UA U7352 ( .D(n1696), .QTFCLK( ), .Q(ofifoData[562]));
Q_MX02 U7353 ( .S(n281), .A0(n2182), .A1(ofifoData[562]), .Z(n1696));
Q_FDP0UA U7354 ( .D(n1695), .QTFCLK( ), .Q(ofifoData[561]));
Q_MX02 U7355 ( .S(n281), .A0(n2183), .A1(ofifoData[561]), .Z(n1695));
Q_FDP0UA U7356 ( .D(n1694), .QTFCLK( ), .Q(ofifoData[560]));
Q_MX02 U7357 ( .S(n281), .A0(n2184), .A1(ofifoData[560]), .Z(n1694));
Q_FDP0UA U7358 ( .D(n1693), .QTFCLK( ), .Q(ofifoData[559]));
Q_MX02 U7359 ( .S(n281), .A0(n2185), .A1(ofifoData[559]), .Z(n1693));
Q_FDP0UA U7360 ( .D(n1692), .QTFCLK( ), .Q(ofifoData[558]));
Q_MX02 U7361 ( .S(n281), .A0(n2186), .A1(ofifoData[558]), .Z(n1692));
Q_FDP0UA U7362 ( .D(n1691), .QTFCLK( ), .Q(ofifoData[557]));
Q_MX02 U7363 ( .S(n281), .A0(n2187), .A1(ofifoData[557]), .Z(n1691));
Q_FDP0UA U7364 ( .D(n1690), .QTFCLK( ), .Q(ofifoData[556]));
Q_MX02 U7365 ( .S(n281), .A0(n2188), .A1(ofifoData[556]), .Z(n1690));
Q_FDP0UA U7366 ( .D(n1689), .QTFCLK( ), .Q(ofifoData[555]));
Q_MX02 U7367 ( .S(n281), .A0(n2189), .A1(ofifoData[555]), .Z(n1689));
Q_FDP0UA U7368 ( .D(n1688), .QTFCLK( ), .Q(ofifoData[554]));
Q_MX02 U7369 ( .S(n281), .A0(n2190), .A1(ofifoData[554]), .Z(n1688));
Q_FDP0UA U7370 ( .D(n1687), .QTFCLK( ), .Q(ofifoData[553]));
Q_MX02 U7371 ( .S(n281), .A0(n2191), .A1(ofifoData[553]), .Z(n1687));
Q_FDP0UA U7372 ( .D(n1686), .QTFCLK( ), .Q(ofifoData[552]));
Q_MX02 U7373 ( .S(n281), .A0(n2192), .A1(ofifoData[552]), .Z(n1686));
Q_FDP0UA U7374 ( .D(n1685), .QTFCLK( ), .Q(ofifoData[551]));
Q_MX02 U7375 ( .S(n281), .A0(n2193), .A1(ofifoData[551]), .Z(n1685));
Q_FDP0UA U7376 ( .D(n1684), .QTFCLK( ), .Q(ofifoData[550]));
Q_MX02 U7377 ( .S(n281), .A0(n2194), .A1(ofifoData[550]), .Z(n1684));
Q_FDP0UA U7378 ( .D(n1683), .QTFCLK( ), .Q(ofifoData[549]));
Q_MX02 U7379 ( .S(n281), .A0(n2195), .A1(ofifoData[549]), .Z(n1683));
Q_FDP0UA U7380 ( .D(n1682), .QTFCLK( ), .Q(ofifoData[548]));
Q_MX02 U7381 ( .S(n281), .A0(n2196), .A1(ofifoData[548]), .Z(n1682));
Q_FDP0UA U7382 ( .D(n1681), .QTFCLK( ), .Q(ofifoData[547]));
Q_MX02 U7383 ( .S(n281), .A0(n2197), .A1(ofifoData[547]), .Z(n1681));
Q_FDP0UA U7384 ( .D(n1680), .QTFCLK( ), .Q(ofifoData[546]));
Q_MX02 U7385 ( .S(n281), .A0(n2198), .A1(ofifoData[546]), .Z(n1680));
Q_FDP0UA U7386 ( .D(n1679), .QTFCLK( ), .Q(ofifoData[545]));
Q_MX02 U7387 ( .S(n281), .A0(n2199), .A1(ofifoData[545]), .Z(n1679));
Q_FDP0UA U7388 ( .D(n1678), .QTFCLK( ), .Q(ofifoData[544]));
Q_MX02 U7389 ( .S(n281), .A0(n2200), .A1(ofifoData[544]), .Z(n1678));
Q_FDP0UA U7390 ( .D(n1677), .QTFCLK( ), .Q(ofifoData[543]));
Q_MX02 U7391 ( .S(n281), .A0(n2201), .A1(ofifoData[543]), .Z(n1677));
Q_FDP0UA U7392 ( .D(n1676), .QTFCLK( ), .Q(ofifoData[542]));
Q_MX02 U7393 ( .S(n281), .A0(n2202), .A1(ofifoData[542]), .Z(n1676));
Q_FDP0UA U7394 ( .D(n1675), .QTFCLK( ), .Q(ofifoData[541]));
Q_MX02 U7395 ( .S(n281), .A0(n2203), .A1(ofifoData[541]), .Z(n1675));
Q_FDP0UA U7396 ( .D(n1674), .QTFCLK( ), .Q(ofifoData[540]));
Q_MX02 U7397 ( .S(n281), .A0(n2204), .A1(ofifoData[540]), .Z(n1674));
Q_FDP0UA U7398 ( .D(n1673), .QTFCLK( ), .Q(ofifoData[539]));
Q_MX02 U7399 ( .S(n281), .A0(n2205), .A1(ofifoData[539]), .Z(n1673));
Q_FDP0UA U7400 ( .D(n1672), .QTFCLK( ), .Q(ofifoData[538]));
Q_MX02 U7401 ( .S(n281), .A0(n2206), .A1(ofifoData[538]), .Z(n1672));
Q_FDP0UA U7402 ( .D(n1671), .QTFCLK( ), .Q(ofifoData[537]));
Q_MX02 U7403 ( .S(n281), .A0(n2207), .A1(ofifoData[537]), .Z(n1671));
Q_FDP0UA U7404 ( .D(n1670), .QTFCLK( ), .Q(ofifoData[536]));
Q_MX02 U7405 ( .S(n281), .A0(n2208), .A1(ofifoData[536]), .Z(n1670));
Q_FDP0UA U7406 ( .D(n1669), .QTFCLK( ), .Q(ofifoData[535]));
Q_MX02 U7407 ( .S(n281), .A0(n2209), .A1(ofifoData[535]), .Z(n1669));
Q_FDP0UA U7408 ( .D(n1668), .QTFCLK( ), .Q(ofifoData[534]));
Q_MX02 U7409 ( .S(n281), .A0(n2210), .A1(ofifoData[534]), .Z(n1668));
Q_FDP0UA U7410 ( .D(n1667), .QTFCLK( ), .Q(ofifoData[533]));
Q_MX02 U7411 ( .S(n281), .A0(n2211), .A1(ofifoData[533]), .Z(n1667));
Q_FDP0UA U7412 ( .D(n1666), .QTFCLK( ), .Q(ofifoData[532]));
Q_MX02 U7413 ( .S(n281), .A0(n2212), .A1(ofifoData[532]), .Z(n1666));
Q_FDP0UA U7414 ( .D(n1665), .QTFCLK( ), .Q(ofifoData[531]));
Q_MX02 U7415 ( .S(n281), .A0(n2213), .A1(ofifoData[531]), .Z(n1665));
Q_FDP0UA U7416 ( .D(n1664), .QTFCLK( ), .Q(ofifoData[530]));
Q_MX02 U7417 ( .S(n281), .A0(n2214), .A1(ofifoData[530]), .Z(n1664));
Q_FDP0UA U7418 ( .D(n1663), .QTFCLK( ), .Q(ofifoData[529]));
Q_MX02 U7419 ( .S(n281), .A0(n2215), .A1(ofifoData[529]), .Z(n1663));
Q_FDP0UA U7420 ( .D(n1662), .QTFCLK( ), .Q(ofifoData[528]));
Q_MX02 U7421 ( .S(n281), .A0(n2216), .A1(ofifoData[528]), .Z(n1662));
Q_FDP0UA U7422 ( .D(n1661), .QTFCLK( ), .Q(ofifoData[527]));
Q_MX02 U7423 ( .S(n281), .A0(n2217), .A1(ofifoData[527]), .Z(n1661));
Q_FDP0UA U7424 ( .D(n1660), .QTFCLK( ), .Q(ofifoData[526]));
Q_MX02 U7425 ( .S(n281), .A0(n2218), .A1(ofifoData[526]), .Z(n1660));
Q_FDP0UA U7426 ( .D(n1659), .QTFCLK( ), .Q(ofifoData[525]));
Q_MX02 U7427 ( .S(n281), .A0(n2219), .A1(ofifoData[525]), .Z(n1659));
Q_FDP0UA U7428 ( .D(n1658), .QTFCLK( ), .Q(ofifoData[524]));
Q_MX02 U7429 ( .S(n281), .A0(n2220), .A1(ofifoData[524]), .Z(n1658));
Q_FDP0UA U7430 ( .D(n1657), .QTFCLK( ), .Q(ofifoData[523]));
Q_MX02 U7431 ( .S(n281), .A0(n2221), .A1(ofifoData[523]), .Z(n1657));
Q_FDP0UA U7432 ( .D(n1656), .QTFCLK( ), .Q(ofifoData[522]));
Q_MX02 U7433 ( .S(n281), .A0(n2222), .A1(ofifoData[522]), .Z(n1656));
Q_FDP0UA U7434 ( .D(n1655), .QTFCLK( ), .Q(ofifoData[521]));
Q_MX02 U7435 ( .S(n281), .A0(n2223), .A1(ofifoData[521]), .Z(n1655));
Q_FDP0UA U7436 ( .D(n1654), .QTFCLK( ), .Q(ofifoData[520]));
Q_MX02 U7437 ( .S(n281), .A0(n2224), .A1(ofifoData[520]), .Z(n1654));
Q_FDP0UA U7438 ( .D(n1653), .QTFCLK( ), .Q(ofifoData[519]));
Q_MX02 U7439 ( .S(n281), .A0(n2225), .A1(ofifoData[519]), .Z(n1653));
Q_FDP0UA U7440 ( .D(n1652), .QTFCLK( ), .Q(ofifoData[518]));
Q_MX02 U7441 ( .S(n281), .A0(n2226), .A1(ofifoData[518]), .Z(n1652));
Q_FDP0UA U7442 ( .D(n1651), .QTFCLK( ), .Q(ofifoData[517]));
Q_MX02 U7443 ( .S(n281), .A0(n2227), .A1(ofifoData[517]), .Z(n1651));
Q_FDP0UA U7444 ( .D(n1650), .QTFCLK( ), .Q(ofifoData[516]));
Q_MX02 U7445 ( .S(n281), .A0(n2228), .A1(ofifoData[516]), .Z(n1650));
Q_FDP0UA U7446 ( .D(n1649), .QTFCLK( ), .Q(ofifoData[515]));
Q_MX02 U7447 ( .S(n281), .A0(n2229), .A1(ofifoData[515]), .Z(n1649));
Q_FDP0UA U7448 ( .D(n1648), .QTFCLK( ), .Q(ofifoData[514]));
Q_MX02 U7449 ( .S(n281), .A0(n2230), .A1(ofifoData[514]), .Z(n1648));
Q_FDP0UA U7450 ( .D(n1647), .QTFCLK( ), .Q(ofifoData[513]));
Q_MX02 U7451 ( .S(n281), .A0(n2231), .A1(ofifoData[513]), .Z(n1647));
Q_FDP0UA U7452 ( .D(n1646), .QTFCLK( ), .Q(ofifoData[512]));
Q_MX02 U7453 ( .S(n281), .A0(n2232), .A1(ofifoData[512]), .Z(n1646));
Q_FDP0UA U7454 ( .D(n1645), .QTFCLK( ), .Q(ofifoData[511]));
Q_MX02 U7455 ( .S(n281), .A0(n2233), .A1(ofifoData[511]), .Z(n1645));
Q_FDP0UA U7456 ( .D(n1644), .QTFCLK( ), .Q(ofifoData[510]));
Q_MX02 U7457 ( .S(n281), .A0(n2234), .A1(ofifoData[510]), .Z(n1644));
Q_FDP0UA U7458 ( .D(n1643), .QTFCLK( ), .Q(ofifoData[509]));
Q_MX02 U7459 ( .S(n281), .A0(n2235), .A1(ofifoData[509]), .Z(n1643));
Q_FDP0UA U7460 ( .D(n1642), .QTFCLK( ), .Q(ofifoData[508]));
Q_MX02 U7461 ( .S(n281), .A0(n2236), .A1(ofifoData[508]), .Z(n1642));
Q_FDP0UA U7462 ( .D(n1641), .QTFCLK( ), .Q(ofifoData[507]));
Q_MX02 U7463 ( .S(n281), .A0(n2237), .A1(ofifoData[507]), .Z(n1641));
Q_FDP0UA U7464 ( .D(n1640), .QTFCLK( ), .Q(ofifoData[506]));
Q_MX02 U7465 ( .S(n281), .A0(n2238), .A1(ofifoData[506]), .Z(n1640));
Q_FDP0UA U7466 ( .D(n1639), .QTFCLK( ), .Q(ofifoData[505]));
Q_MX02 U7467 ( .S(n281), .A0(n2239), .A1(ofifoData[505]), .Z(n1639));
Q_FDP0UA U7468 ( .D(n1638), .QTFCLK( ), .Q(ofifoData[504]));
Q_MX02 U7469 ( .S(n281), .A0(n2240), .A1(ofifoData[504]), .Z(n1638));
Q_FDP0UA U7470 ( .D(n1637), .QTFCLK( ), .Q(ofifoData[503]));
Q_MX02 U7471 ( .S(n281), .A0(n2241), .A1(ofifoData[503]), .Z(n1637));
Q_FDP0UA U7472 ( .D(n1636), .QTFCLK( ), .Q(ofifoData[502]));
Q_MX02 U7473 ( .S(n281), .A0(n2242), .A1(ofifoData[502]), .Z(n1636));
Q_FDP0UA U7474 ( .D(n1635), .QTFCLK( ), .Q(ofifoData[501]));
Q_MX02 U7475 ( .S(n281), .A0(n2243), .A1(ofifoData[501]), .Z(n1635));
Q_FDP0UA U7476 ( .D(n1634), .QTFCLK( ), .Q(ofifoData[500]));
Q_MX02 U7477 ( .S(n281), .A0(n2244), .A1(ofifoData[500]), .Z(n1634));
Q_FDP0UA U7478 ( .D(n1633), .QTFCLK( ), .Q(ofifoData[499]));
Q_MX02 U7479 ( .S(n281), .A0(n2245), .A1(ofifoData[499]), .Z(n1633));
Q_FDP0UA U7480 ( .D(n1632), .QTFCLK( ), .Q(ofifoData[498]));
Q_MX02 U7481 ( .S(n281), .A0(n2246), .A1(ofifoData[498]), .Z(n1632));
Q_FDP0UA U7482 ( .D(n1631), .QTFCLK( ), .Q(ofifoData[497]));
Q_MX02 U7483 ( .S(n281), .A0(n2247), .A1(ofifoData[497]), .Z(n1631));
Q_FDP0UA U7484 ( .D(n1630), .QTFCLK( ), .Q(ofifoData[496]));
Q_MX02 U7485 ( .S(n281), .A0(n2248), .A1(ofifoData[496]), .Z(n1630));
Q_FDP0UA U7486 ( .D(n1629), .QTFCLK( ), .Q(ofifoData[495]));
Q_MX02 U7487 ( .S(n281), .A0(n2249), .A1(ofifoData[495]), .Z(n1629));
Q_FDP0UA U7488 ( .D(n1628), .QTFCLK( ), .Q(ofifoData[494]));
Q_MX02 U7489 ( .S(n281), .A0(n2250), .A1(ofifoData[494]), .Z(n1628));
Q_FDP0UA U7490 ( .D(n1627), .QTFCLK( ), .Q(ofifoData[493]));
Q_MX02 U7491 ( .S(n281), .A0(n2251), .A1(ofifoData[493]), .Z(n1627));
Q_FDP0UA U7492 ( .D(n1626), .QTFCLK( ), .Q(ofifoData[492]));
Q_MX02 U7493 ( .S(n281), .A0(n2252), .A1(ofifoData[492]), .Z(n1626));
Q_FDP0UA U7494 ( .D(n1625), .QTFCLK( ), .Q(ofifoData[491]));
Q_MX02 U7495 ( .S(n281), .A0(n2253), .A1(ofifoData[491]), .Z(n1625));
Q_FDP0UA U7496 ( .D(n1624), .QTFCLK( ), .Q(ofifoData[490]));
Q_MX02 U7497 ( .S(n281), .A0(n2254), .A1(ofifoData[490]), .Z(n1624));
Q_FDP0UA U7498 ( .D(n1623), .QTFCLK( ), .Q(ofifoData[489]));
Q_MX02 U7499 ( .S(n281), .A0(n2255), .A1(ofifoData[489]), .Z(n1623));
Q_FDP0UA U7500 ( .D(n1622), .QTFCLK( ), .Q(ofifoData[488]));
Q_MX02 U7501 ( .S(n281), .A0(n2256), .A1(ofifoData[488]), .Z(n1622));
Q_FDP0UA U7502 ( .D(n1621), .QTFCLK( ), .Q(ofifoData[487]));
Q_MX02 U7503 ( .S(n281), .A0(n2257), .A1(ofifoData[487]), .Z(n1621));
Q_FDP0UA U7504 ( .D(n1620), .QTFCLK( ), .Q(ofifoData[486]));
Q_MX02 U7505 ( .S(n281), .A0(n2258), .A1(ofifoData[486]), .Z(n1620));
Q_FDP0UA U7506 ( .D(n1619), .QTFCLK( ), .Q(ofifoData[485]));
Q_MX02 U7507 ( .S(n281), .A0(n2259), .A1(ofifoData[485]), .Z(n1619));
Q_FDP0UA U7508 ( .D(n1618), .QTFCLK( ), .Q(ofifoData[484]));
Q_MX02 U7509 ( .S(n281), .A0(n2260), .A1(ofifoData[484]), .Z(n1618));
Q_FDP0UA U7510 ( .D(n1617), .QTFCLK( ), .Q(ofifoData[483]));
Q_MX02 U7511 ( .S(n281), .A0(n2261), .A1(ofifoData[483]), .Z(n1617));
Q_FDP0UA U7512 ( .D(n1616), .QTFCLK( ), .Q(ofifoData[482]));
Q_MX02 U7513 ( .S(n281), .A0(n2262), .A1(ofifoData[482]), .Z(n1616));
Q_FDP0UA U7514 ( .D(n1615), .QTFCLK( ), .Q(ofifoData[481]));
Q_MX02 U7515 ( .S(n281), .A0(n2263), .A1(ofifoData[481]), .Z(n1615));
Q_FDP0UA U7516 ( .D(n1614), .QTFCLK( ), .Q(ofifoData[480]));
Q_MX02 U7517 ( .S(n281), .A0(n2264), .A1(ofifoData[480]), .Z(n1614));
Q_FDP0UA U7518 ( .D(n1613), .QTFCLK( ), .Q(ofifoData[479]));
Q_MX02 U7519 ( .S(n281), .A0(n2265), .A1(ofifoData[479]), .Z(n1613));
Q_FDP0UA U7520 ( .D(n1612), .QTFCLK( ), .Q(ofifoData[478]));
Q_MX02 U7521 ( .S(n281), .A0(n2266), .A1(ofifoData[478]), .Z(n1612));
Q_FDP0UA U7522 ( .D(n1611), .QTFCLK( ), .Q(ofifoData[477]));
Q_MX02 U7523 ( .S(n281), .A0(n2267), .A1(ofifoData[477]), .Z(n1611));
Q_FDP0UA U7524 ( .D(n1610), .QTFCLK( ), .Q(ofifoData[476]));
Q_MX02 U7525 ( .S(n281), .A0(n2268), .A1(ofifoData[476]), .Z(n1610));
Q_FDP0UA U7526 ( .D(n1609), .QTFCLK( ), .Q(ofifoData[475]));
Q_MX02 U7527 ( .S(n281), .A0(n2269), .A1(ofifoData[475]), .Z(n1609));
Q_FDP0UA U7528 ( .D(n1608), .QTFCLK( ), .Q(ofifoData[474]));
Q_MX02 U7529 ( .S(n281), .A0(n2270), .A1(ofifoData[474]), .Z(n1608));
Q_FDP0UA U7530 ( .D(n1607), .QTFCLK( ), .Q(ofifoData[473]));
Q_MX02 U7531 ( .S(n281), .A0(n2271), .A1(ofifoData[473]), .Z(n1607));
Q_FDP0UA U7532 ( .D(n1606), .QTFCLK( ), .Q(ofifoData[472]));
Q_MX02 U7533 ( .S(n281), .A0(n2272), .A1(ofifoData[472]), .Z(n1606));
Q_FDP0UA U7534 ( .D(n1605), .QTFCLK( ), .Q(ofifoData[471]));
Q_MX02 U7535 ( .S(n281), .A0(n2273), .A1(ofifoData[471]), .Z(n1605));
Q_FDP0UA U7536 ( .D(n1604), .QTFCLK( ), .Q(ofifoData[470]));
Q_MX02 U7537 ( .S(n281), .A0(n2274), .A1(ofifoData[470]), .Z(n1604));
Q_FDP0UA U7538 ( .D(n1603), .QTFCLK( ), .Q(ofifoData[469]));
Q_MX02 U7539 ( .S(n281), .A0(n2275), .A1(ofifoData[469]), .Z(n1603));
Q_FDP0UA U7540 ( .D(n1602), .QTFCLK( ), .Q(ofifoData[468]));
Q_MX02 U7541 ( .S(n281), .A0(n2276), .A1(ofifoData[468]), .Z(n1602));
Q_FDP0UA U7542 ( .D(n1601), .QTFCLK( ), .Q(ofifoData[467]));
Q_MX02 U7543 ( .S(n281), .A0(n2277), .A1(ofifoData[467]), .Z(n1601));
Q_FDP0UA U7544 ( .D(n1600), .QTFCLK( ), .Q(ofifoData[466]));
Q_MX02 U7545 ( .S(n281), .A0(n2278), .A1(ofifoData[466]), .Z(n1600));
Q_FDP0UA U7546 ( .D(n1599), .QTFCLK( ), .Q(ofifoData[465]));
Q_MX02 U7547 ( .S(n281), .A0(n2279), .A1(ofifoData[465]), .Z(n1599));
Q_FDP0UA U7548 ( .D(n1598), .QTFCLK( ), .Q(ofifoData[464]));
Q_MX02 U7549 ( .S(n281), .A0(n2280), .A1(ofifoData[464]), .Z(n1598));
Q_FDP0UA U7550 ( .D(n1597), .QTFCLK( ), .Q(ofifoData[463]));
Q_MX02 U7551 ( .S(n281), .A0(n2281), .A1(ofifoData[463]), .Z(n1597));
Q_FDP0UA U7552 ( .D(n1596), .QTFCLK( ), .Q(ofifoData[462]));
Q_MX02 U7553 ( .S(n281), .A0(n2282), .A1(ofifoData[462]), .Z(n1596));
Q_FDP0UA U7554 ( .D(n1595), .QTFCLK( ), .Q(ofifoData[461]));
Q_MX02 U7555 ( .S(n281), .A0(n2283), .A1(ofifoData[461]), .Z(n1595));
Q_FDP0UA U7556 ( .D(n1594), .QTFCLK( ), .Q(ofifoData[460]));
Q_MX02 U7557 ( .S(n281), .A0(n2284), .A1(ofifoData[460]), .Z(n1594));
Q_FDP0UA U7558 ( .D(n1593), .QTFCLK( ), .Q(ofifoData[459]));
Q_MX02 U7559 ( .S(n281), .A0(n2285), .A1(ofifoData[459]), .Z(n1593));
Q_FDP0UA U7560 ( .D(n1592), .QTFCLK( ), .Q(ofifoData[458]));
Q_MX02 U7561 ( .S(n281), .A0(n2286), .A1(ofifoData[458]), .Z(n1592));
Q_FDP0UA U7562 ( .D(n1591), .QTFCLK( ), .Q(ofifoData[457]));
Q_MX02 U7563 ( .S(n281), .A0(n2287), .A1(ofifoData[457]), .Z(n1591));
Q_FDP0UA U7564 ( .D(n1590), .QTFCLK( ), .Q(ofifoData[456]));
Q_MX02 U7565 ( .S(n281), .A0(n2288), .A1(ofifoData[456]), .Z(n1590));
Q_FDP0UA U7566 ( .D(n1589), .QTFCLK( ), .Q(ofifoData[455]));
Q_MX02 U7567 ( .S(n281), .A0(n2289), .A1(ofifoData[455]), .Z(n1589));
Q_FDP0UA U7568 ( .D(n1588), .QTFCLK( ), .Q(ofifoData[454]));
Q_MX02 U7569 ( .S(n281), .A0(n2290), .A1(ofifoData[454]), .Z(n1588));
Q_FDP0UA U7570 ( .D(n1587), .QTFCLK( ), .Q(ofifoData[453]));
Q_MX02 U7571 ( .S(n281), .A0(n2291), .A1(ofifoData[453]), .Z(n1587));
Q_FDP0UA U7572 ( .D(n1586), .QTFCLK( ), .Q(ofifoData[452]));
Q_MX02 U7573 ( .S(n281), .A0(n2292), .A1(ofifoData[452]), .Z(n1586));
Q_FDP0UA U7574 ( .D(n1585), .QTFCLK( ), .Q(ofifoData[451]));
Q_MX02 U7575 ( .S(n281), .A0(n2293), .A1(ofifoData[451]), .Z(n1585));
Q_FDP0UA U7576 ( .D(n1584), .QTFCLK( ), .Q(ofifoData[450]));
Q_MX02 U7577 ( .S(n281), .A0(n2294), .A1(ofifoData[450]), .Z(n1584));
Q_FDP0UA U7578 ( .D(n1583), .QTFCLK( ), .Q(ofifoData[449]));
Q_MX02 U7579 ( .S(n281), .A0(n2295), .A1(ofifoData[449]), .Z(n1583));
Q_FDP0UA U7580 ( .D(n1582), .QTFCLK( ), .Q(ofifoData[448]));
Q_MX02 U7581 ( .S(n281), .A0(n2296), .A1(ofifoData[448]), .Z(n1582));
Q_FDP0UA U7582 ( .D(n1581), .QTFCLK( ), .Q(ofifoData[447]));
Q_MX02 U7583 ( .S(n281), .A0(n2297), .A1(ofifoData[447]), .Z(n1581));
Q_FDP0UA U7584 ( .D(n1580), .QTFCLK( ), .Q(ofifoData[446]));
Q_MX02 U7585 ( .S(n281), .A0(n2298), .A1(ofifoData[446]), .Z(n1580));
Q_FDP0UA U7586 ( .D(n1579), .QTFCLK( ), .Q(ofifoData[445]));
Q_MX02 U7587 ( .S(n281), .A0(n2299), .A1(ofifoData[445]), .Z(n1579));
Q_FDP0UA U7588 ( .D(n1578), .QTFCLK( ), .Q(ofifoData[444]));
Q_MX02 U7589 ( .S(n281), .A0(n2300), .A1(ofifoData[444]), .Z(n1578));
Q_FDP0UA U7590 ( .D(n1577), .QTFCLK( ), .Q(ofifoData[443]));
Q_MX02 U7591 ( .S(n281), .A0(n2301), .A1(ofifoData[443]), .Z(n1577));
Q_FDP0UA U7592 ( .D(n1576), .QTFCLK( ), .Q(ofifoData[442]));
Q_MX02 U7593 ( .S(n281), .A0(n2302), .A1(ofifoData[442]), .Z(n1576));
Q_FDP0UA U7594 ( .D(n1575), .QTFCLK( ), .Q(ofifoData[441]));
Q_MX02 U7595 ( .S(n281), .A0(n2303), .A1(ofifoData[441]), .Z(n1575));
Q_FDP0UA U7596 ( .D(n1574), .QTFCLK( ), .Q(ofifoData[440]));
Q_MX02 U7597 ( .S(n281), .A0(n2304), .A1(ofifoData[440]), .Z(n1574));
Q_FDP0UA U7598 ( .D(n1573), .QTFCLK( ), .Q(ofifoData[439]));
Q_MX02 U7599 ( .S(n281), .A0(n2305), .A1(ofifoData[439]), .Z(n1573));
Q_FDP0UA U7600 ( .D(n1572), .QTFCLK( ), .Q(ofifoData[438]));
Q_MX02 U7601 ( .S(n281), .A0(n2306), .A1(ofifoData[438]), .Z(n1572));
Q_FDP0UA U7602 ( .D(n1571), .QTFCLK( ), .Q(ofifoData[437]));
Q_MX02 U7603 ( .S(n281), .A0(n2307), .A1(ofifoData[437]), .Z(n1571));
Q_FDP0UA U7604 ( .D(n1570), .QTFCLK( ), .Q(ofifoData[436]));
Q_MX02 U7605 ( .S(n281), .A0(n2308), .A1(ofifoData[436]), .Z(n1570));
Q_FDP0UA U7606 ( .D(n1569), .QTFCLK( ), .Q(ofifoData[435]));
Q_MX02 U7607 ( .S(n281), .A0(n2309), .A1(ofifoData[435]), .Z(n1569));
Q_FDP0UA U7608 ( .D(n1568), .QTFCLK( ), .Q(ofifoData[434]));
Q_MX02 U7609 ( .S(n281), .A0(n2310), .A1(ofifoData[434]), .Z(n1568));
Q_FDP0UA U7610 ( .D(n1567), .QTFCLK( ), .Q(ofifoData[433]));
Q_MX02 U7611 ( .S(n281), .A0(n2311), .A1(ofifoData[433]), .Z(n1567));
Q_FDP0UA U7612 ( .D(n1566), .QTFCLK( ), .Q(ofifoData[432]));
Q_MX02 U7613 ( .S(n281), .A0(n2312), .A1(ofifoData[432]), .Z(n1566));
Q_FDP0UA U7614 ( .D(n1565), .QTFCLK( ), .Q(ofifoData[431]));
Q_MX02 U7615 ( .S(n281), .A0(n2313), .A1(ofifoData[431]), .Z(n1565));
Q_FDP0UA U7616 ( .D(n1564), .QTFCLK( ), .Q(ofifoData[430]));
Q_MX02 U7617 ( .S(n281), .A0(n2314), .A1(ofifoData[430]), .Z(n1564));
Q_FDP0UA U7618 ( .D(n1563), .QTFCLK( ), .Q(ofifoData[429]));
Q_MX02 U7619 ( .S(n281), .A0(n2315), .A1(ofifoData[429]), .Z(n1563));
Q_FDP0UA U7620 ( .D(n1562), .QTFCLK( ), .Q(ofifoData[428]));
Q_MX02 U7621 ( .S(n281), .A0(n2316), .A1(ofifoData[428]), .Z(n1562));
Q_FDP0UA U7622 ( .D(n1561), .QTFCLK( ), .Q(ofifoData[427]));
Q_MX02 U7623 ( .S(n281), .A0(n2317), .A1(ofifoData[427]), .Z(n1561));
Q_FDP0UA U7624 ( .D(n1560), .QTFCLK( ), .Q(ofifoData[426]));
Q_MX02 U7625 ( .S(n281), .A0(n2318), .A1(ofifoData[426]), .Z(n1560));
Q_FDP0UA U7626 ( .D(n1559), .QTFCLK( ), .Q(ofifoData[425]));
Q_MX02 U7627 ( .S(n281), .A0(n2319), .A1(ofifoData[425]), .Z(n1559));
Q_FDP0UA U7628 ( .D(n1558), .QTFCLK( ), .Q(ofifoData[424]));
Q_MX02 U7629 ( .S(n281), .A0(n2320), .A1(ofifoData[424]), .Z(n1558));
Q_FDP0UA U7630 ( .D(n1557), .QTFCLK( ), .Q(ofifoData[423]));
Q_MX02 U7631 ( .S(n281), .A0(n2321), .A1(ofifoData[423]), .Z(n1557));
Q_FDP0UA U7632 ( .D(n1556), .QTFCLK( ), .Q(ofifoData[422]));
Q_MX02 U7633 ( .S(n281), .A0(n2322), .A1(ofifoData[422]), .Z(n1556));
Q_FDP0UA U7634 ( .D(n1555), .QTFCLK( ), .Q(ofifoData[421]));
Q_MX02 U7635 ( .S(n281), .A0(n2323), .A1(ofifoData[421]), .Z(n1555));
Q_FDP0UA U7636 ( .D(n1554), .QTFCLK( ), .Q(ofifoData[420]));
Q_MX02 U7637 ( .S(n281), .A0(n2324), .A1(ofifoData[420]), .Z(n1554));
Q_FDP0UA U7638 ( .D(n1553), .QTFCLK( ), .Q(ofifoData[419]));
Q_MX02 U7639 ( .S(n281), .A0(n2325), .A1(ofifoData[419]), .Z(n1553));
Q_FDP0UA U7640 ( .D(n1552), .QTFCLK( ), .Q(ofifoData[418]));
Q_MX02 U7641 ( .S(n281), .A0(n2326), .A1(ofifoData[418]), .Z(n1552));
Q_FDP0UA U7642 ( .D(n1551), .QTFCLK( ), .Q(ofifoData[417]));
Q_MX02 U7643 ( .S(n281), .A0(n2327), .A1(ofifoData[417]), .Z(n1551));
Q_FDP0UA U7644 ( .D(n1550), .QTFCLK( ), .Q(ofifoData[416]));
Q_MX02 U7645 ( .S(n281), .A0(n2328), .A1(ofifoData[416]), .Z(n1550));
Q_FDP0UA U7646 ( .D(n1549), .QTFCLK( ), .Q(ofifoData[415]));
Q_MX02 U7647 ( .S(n281), .A0(n2329), .A1(ofifoData[415]), .Z(n1549));
Q_FDP0UA U7648 ( .D(n1548), .QTFCLK( ), .Q(ofifoData[414]));
Q_MX02 U7649 ( .S(n281), .A0(n2330), .A1(ofifoData[414]), .Z(n1548));
Q_FDP0UA U7650 ( .D(n1547), .QTFCLK( ), .Q(ofifoData[413]));
Q_MX02 U7651 ( .S(n281), .A0(n2331), .A1(ofifoData[413]), .Z(n1547));
Q_FDP0UA U7652 ( .D(n1546), .QTFCLK( ), .Q(ofifoData[412]));
Q_MX02 U7653 ( .S(n281), .A0(n2332), .A1(ofifoData[412]), .Z(n1546));
Q_FDP0UA U7654 ( .D(n1545), .QTFCLK( ), .Q(ofifoData[411]));
Q_MX02 U7655 ( .S(n281), .A0(n2333), .A1(ofifoData[411]), .Z(n1545));
Q_FDP0UA U7656 ( .D(n1544), .QTFCLK( ), .Q(ofifoData[410]));
Q_MX02 U7657 ( .S(n281), .A0(n2334), .A1(ofifoData[410]), .Z(n1544));
Q_FDP0UA U7658 ( .D(n1543), .QTFCLK( ), .Q(ofifoData[409]));
Q_MX02 U7659 ( .S(n281), .A0(n2335), .A1(ofifoData[409]), .Z(n1543));
Q_FDP0UA U7660 ( .D(n1542), .QTFCLK( ), .Q(ofifoData[408]));
Q_MX02 U7661 ( .S(n281), .A0(n2336), .A1(ofifoData[408]), .Z(n1542));
Q_FDP0UA U7662 ( .D(n1541), .QTFCLK( ), .Q(ofifoData[407]));
Q_MX02 U7663 ( .S(n281), .A0(n2337), .A1(ofifoData[407]), .Z(n1541));
Q_FDP0UA U7664 ( .D(n1540), .QTFCLK( ), .Q(ofifoData[406]));
Q_MX02 U7665 ( .S(n281), .A0(n2338), .A1(ofifoData[406]), .Z(n1540));
Q_FDP0UA U7666 ( .D(n1539), .QTFCLK( ), .Q(ofifoData[405]));
Q_MX02 U7667 ( .S(n281), .A0(n2339), .A1(ofifoData[405]), .Z(n1539));
Q_FDP0UA U7668 ( .D(n1538), .QTFCLK( ), .Q(ofifoData[404]));
Q_MX02 U7669 ( .S(n281), .A0(n2340), .A1(ofifoData[404]), .Z(n1538));
Q_FDP0UA U7670 ( .D(n1537), .QTFCLK( ), .Q(ofifoData[403]));
Q_MX02 U7671 ( .S(n281), .A0(n2341), .A1(ofifoData[403]), .Z(n1537));
Q_FDP0UA U7672 ( .D(n1536), .QTFCLK( ), .Q(ofifoData[402]));
Q_MX02 U7673 ( .S(n281), .A0(n2342), .A1(ofifoData[402]), .Z(n1536));
Q_FDP0UA U7674 ( .D(n1535), .QTFCLK( ), .Q(ofifoData[401]));
Q_MX02 U7675 ( .S(n281), .A0(n2343), .A1(ofifoData[401]), .Z(n1535));
Q_FDP0UA U7676 ( .D(n1534), .QTFCLK( ), .Q(ofifoData[400]));
Q_MX02 U7677 ( .S(n281), .A0(n2344), .A1(ofifoData[400]), .Z(n1534));
Q_FDP0UA U7678 ( .D(n1533), .QTFCLK( ), .Q(ofifoData[399]));
Q_MX02 U7679 ( .S(n281), .A0(n2345), .A1(ofifoData[399]), .Z(n1533));
Q_FDP0UA U7680 ( .D(n1532), .QTFCLK( ), .Q(ofifoData[398]));
Q_MX02 U7681 ( .S(n281), .A0(n2346), .A1(ofifoData[398]), .Z(n1532));
Q_FDP0UA U7682 ( .D(n1531), .QTFCLK( ), .Q(ofifoData[397]));
Q_MX02 U7683 ( .S(n281), .A0(n2347), .A1(ofifoData[397]), .Z(n1531));
Q_FDP0UA U7684 ( .D(n1530), .QTFCLK( ), .Q(ofifoData[396]));
Q_MX02 U7685 ( .S(n281), .A0(n2348), .A1(ofifoData[396]), .Z(n1530));
Q_FDP0UA U7686 ( .D(n1529), .QTFCLK( ), .Q(ofifoData[395]));
Q_MX02 U7687 ( .S(n281), .A0(n2349), .A1(ofifoData[395]), .Z(n1529));
Q_FDP0UA U7688 ( .D(n1528), .QTFCLK( ), .Q(ofifoData[394]));
Q_MX02 U7689 ( .S(n281), .A0(n2350), .A1(ofifoData[394]), .Z(n1528));
Q_FDP0UA U7690 ( .D(n1527), .QTFCLK( ), .Q(ofifoData[393]));
Q_MX02 U7691 ( .S(n281), .A0(n2351), .A1(ofifoData[393]), .Z(n1527));
Q_FDP0UA U7692 ( .D(n1526), .QTFCLK( ), .Q(ofifoData[392]));
Q_MX02 U7693 ( .S(n281), .A0(n2352), .A1(ofifoData[392]), .Z(n1526));
Q_FDP0UA U7694 ( .D(n1525), .QTFCLK( ), .Q(ofifoData[391]));
Q_MX02 U7695 ( .S(n281), .A0(n2353), .A1(ofifoData[391]), .Z(n1525));
Q_FDP0UA U7696 ( .D(n1524), .QTFCLK( ), .Q(ofifoData[390]));
Q_MX02 U7697 ( .S(n281), .A0(n2354), .A1(ofifoData[390]), .Z(n1524));
Q_FDP0UA U7698 ( .D(n1523), .QTFCLK( ), .Q(ofifoData[389]));
Q_MX02 U7699 ( .S(n281), .A0(n2355), .A1(ofifoData[389]), .Z(n1523));
Q_FDP0UA U7700 ( .D(n1522), .QTFCLK( ), .Q(ofifoData[388]));
Q_MX02 U7701 ( .S(n281), .A0(n2356), .A1(ofifoData[388]), .Z(n1522));
Q_FDP0UA U7702 ( .D(n1521), .QTFCLK( ), .Q(ofifoData[387]));
Q_MX02 U7703 ( .S(n281), .A0(n2357), .A1(ofifoData[387]), .Z(n1521));
Q_FDP0UA U7704 ( .D(n1520), .QTFCLK( ), .Q(ofifoData[386]));
Q_MX02 U7705 ( .S(n281), .A0(n2358), .A1(ofifoData[386]), .Z(n1520));
Q_FDP0UA U7706 ( .D(n1519), .QTFCLK( ), .Q(ofifoData[385]));
Q_MX02 U7707 ( .S(n281), .A0(n2359), .A1(ofifoData[385]), .Z(n1519));
Q_FDP0UA U7708 ( .D(n1518), .QTFCLK( ), .Q(ofifoData[384]));
Q_MX02 U7709 ( .S(n281), .A0(n2360), .A1(ofifoData[384]), .Z(n1518));
Q_FDP0UA U7710 ( .D(n1517), .QTFCLK( ), .Q(ofifoData[383]));
Q_MX02 U7711 ( .S(n281), .A0(n2361), .A1(ofifoData[383]), .Z(n1517));
Q_FDP0UA U7712 ( .D(n1516), .QTFCLK( ), .Q(ofifoData[382]));
Q_MX02 U7713 ( .S(n281), .A0(n2362), .A1(ofifoData[382]), .Z(n1516));
Q_FDP0UA U7714 ( .D(n1515), .QTFCLK( ), .Q(ofifoData[381]));
Q_MX02 U7715 ( .S(n281), .A0(n2363), .A1(ofifoData[381]), .Z(n1515));
Q_FDP0UA U7716 ( .D(n1514), .QTFCLK( ), .Q(ofifoData[380]));
Q_MX02 U7717 ( .S(n281), .A0(n2364), .A1(ofifoData[380]), .Z(n1514));
Q_FDP0UA U7718 ( .D(n1513), .QTFCLK( ), .Q(ofifoData[379]));
Q_MX02 U7719 ( .S(n281), .A0(n2365), .A1(ofifoData[379]), .Z(n1513));
Q_FDP0UA U7720 ( .D(n1512), .QTFCLK( ), .Q(ofifoData[378]));
Q_MX02 U7721 ( .S(n281), .A0(n2366), .A1(ofifoData[378]), .Z(n1512));
Q_FDP0UA U7722 ( .D(n1511), .QTFCLK( ), .Q(ofifoData[377]));
Q_MX02 U7723 ( .S(n281), .A0(n2367), .A1(ofifoData[377]), .Z(n1511));
Q_FDP0UA U7724 ( .D(n1510), .QTFCLK( ), .Q(ofifoData[376]));
Q_MX02 U7725 ( .S(n281), .A0(n2368), .A1(ofifoData[376]), .Z(n1510));
Q_FDP0UA U7726 ( .D(n1509), .QTFCLK( ), .Q(ofifoData[375]));
Q_MX02 U7727 ( .S(n281), .A0(n2369), .A1(ofifoData[375]), .Z(n1509));
Q_FDP0UA U7728 ( .D(n1508), .QTFCLK( ), .Q(ofifoData[374]));
Q_MX02 U7729 ( .S(n281), .A0(n2370), .A1(ofifoData[374]), .Z(n1508));
Q_FDP0UA U7730 ( .D(n1507), .QTFCLK( ), .Q(ofifoData[373]));
Q_MX02 U7731 ( .S(n281), .A0(n2371), .A1(ofifoData[373]), .Z(n1507));
Q_FDP0UA U7732 ( .D(n1506), .QTFCLK( ), .Q(ofifoData[372]));
Q_MX02 U7733 ( .S(n281), .A0(n2372), .A1(ofifoData[372]), .Z(n1506));
Q_FDP0UA U7734 ( .D(n1505), .QTFCLK( ), .Q(ofifoData[371]));
Q_MX02 U7735 ( .S(n281), .A0(n2373), .A1(ofifoData[371]), .Z(n1505));
Q_FDP0UA U7736 ( .D(n1504), .QTFCLK( ), .Q(ofifoData[370]));
Q_MX02 U7737 ( .S(n281), .A0(n2374), .A1(ofifoData[370]), .Z(n1504));
Q_FDP0UA U7738 ( .D(n1503), .QTFCLK( ), .Q(ofifoData[369]));
Q_MX02 U7739 ( .S(n281), .A0(n2375), .A1(ofifoData[369]), .Z(n1503));
Q_FDP0UA U7740 ( .D(n1502), .QTFCLK( ), .Q(ofifoData[368]));
Q_MX02 U7741 ( .S(n281), .A0(n2376), .A1(ofifoData[368]), .Z(n1502));
Q_FDP0UA U7742 ( .D(n1501), .QTFCLK( ), .Q(ofifoData[367]));
Q_MX02 U7743 ( .S(n281), .A0(n2377), .A1(ofifoData[367]), .Z(n1501));
Q_FDP0UA U7744 ( .D(n1500), .QTFCLK( ), .Q(ofifoData[366]));
Q_MX02 U7745 ( .S(n281), .A0(n2378), .A1(ofifoData[366]), .Z(n1500));
Q_FDP0UA U7746 ( .D(n1499), .QTFCLK( ), .Q(ofifoData[365]));
Q_MX02 U7747 ( .S(n281), .A0(n2379), .A1(ofifoData[365]), .Z(n1499));
Q_FDP0UA U7748 ( .D(n1498), .QTFCLK( ), .Q(ofifoData[364]));
Q_MX02 U7749 ( .S(n281), .A0(n2380), .A1(ofifoData[364]), .Z(n1498));
Q_FDP0UA U7750 ( .D(n1497), .QTFCLK( ), .Q(ofifoData[363]));
Q_MX02 U7751 ( .S(n281), .A0(n2381), .A1(ofifoData[363]), .Z(n1497));
Q_FDP0UA U7752 ( .D(n1496), .QTFCLK( ), .Q(ofifoData[362]));
Q_MX02 U7753 ( .S(n281), .A0(n2382), .A1(ofifoData[362]), .Z(n1496));
Q_FDP0UA U7754 ( .D(n1495), .QTFCLK( ), .Q(ofifoData[361]));
Q_MX02 U7755 ( .S(n281), .A0(n2383), .A1(ofifoData[361]), .Z(n1495));
Q_FDP0UA U7756 ( .D(n1494), .QTFCLK( ), .Q(ofifoData[360]));
Q_MX02 U7757 ( .S(n281), .A0(n2384), .A1(ofifoData[360]), .Z(n1494));
Q_FDP0UA U7758 ( .D(n1493), .QTFCLK( ), .Q(ofifoData[359]));
Q_MX02 U7759 ( .S(n281), .A0(n2385), .A1(ofifoData[359]), .Z(n1493));
Q_FDP0UA U7760 ( .D(n1492), .QTFCLK( ), .Q(ofifoData[358]));
Q_MX02 U7761 ( .S(n281), .A0(n2386), .A1(ofifoData[358]), .Z(n1492));
Q_FDP0UA U7762 ( .D(n1491), .QTFCLK( ), .Q(ofifoData[357]));
Q_MX02 U7763 ( .S(n281), .A0(n2387), .A1(ofifoData[357]), .Z(n1491));
Q_FDP0UA U7764 ( .D(n1490), .QTFCLK( ), .Q(ofifoData[356]));
Q_MX02 U7765 ( .S(n281), .A0(n2388), .A1(ofifoData[356]), .Z(n1490));
Q_FDP0UA U7766 ( .D(n1489), .QTFCLK( ), .Q(ofifoData[355]));
Q_MX02 U7767 ( .S(n281), .A0(n2389), .A1(ofifoData[355]), .Z(n1489));
Q_FDP0UA U7768 ( .D(n1488), .QTFCLK( ), .Q(ofifoData[354]));
Q_MX02 U7769 ( .S(n281), .A0(n2390), .A1(ofifoData[354]), .Z(n1488));
Q_FDP0UA U7770 ( .D(n1487), .QTFCLK( ), .Q(ofifoData[353]));
Q_MX02 U7771 ( .S(n281), .A0(n2391), .A1(ofifoData[353]), .Z(n1487));
Q_FDP0UA U7772 ( .D(n1486), .QTFCLK( ), .Q(ofifoData[352]));
Q_MX02 U7773 ( .S(n281), .A0(n2392), .A1(ofifoData[352]), .Z(n1486));
Q_FDP0UA U7774 ( .D(n1485), .QTFCLK( ), .Q(ofifoData[351]));
Q_MX02 U7775 ( .S(n281), .A0(n2393), .A1(ofifoData[351]), .Z(n1485));
Q_FDP0UA U7776 ( .D(n1484), .QTFCLK( ), .Q(ofifoData[350]));
Q_MX02 U7777 ( .S(n281), .A0(n2394), .A1(ofifoData[350]), .Z(n1484));
Q_FDP0UA U7778 ( .D(n1483), .QTFCLK( ), .Q(ofifoData[349]));
Q_MX02 U7779 ( .S(n281), .A0(n2395), .A1(ofifoData[349]), .Z(n1483));
Q_FDP0UA U7780 ( .D(n1482), .QTFCLK( ), .Q(ofifoData[348]));
Q_MX02 U7781 ( .S(n281), .A0(n2396), .A1(ofifoData[348]), .Z(n1482));
Q_FDP0UA U7782 ( .D(n1481), .QTFCLK( ), .Q(ofifoData[347]));
Q_MX02 U7783 ( .S(n281), .A0(n2397), .A1(ofifoData[347]), .Z(n1481));
Q_FDP0UA U7784 ( .D(n1480), .QTFCLK( ), .Q(ofifoData[346]));
Q_MX02 U7785 ( .S(n281), .A0(n2398), .A1(ofifoData[346]), .Z(n1480));
Q_FDP0UA U7786 ( .D(n1479), .QTFCLK( ), .Q(ofifoData[345]));
Q_MX02 U7787 ( .S(n281), .A0(n2399), .A1(ofifoData[345]), .Z(n1479));
Q_FDP0UA U7788 ( .D(n1478), .QTFCLK( ), .Q(ofifoData[344]));
Q_MX02 U7789 ( .S(n281), .A0(n2400), .A1(ofifoData[344]), .Z(n1478));
Q_FDP0UA U7790 ( .D(n1477), .QTFCLK( ), .Q(ofifoData[343]));
Q_MX02 U7791 ( .S(n281), .A0(n2401), .A1(ofifoData[343]), .Z(n1477));
Q_FDP0UA U7792 ( .D(n1476), .QTFCLK( ), .Q(ofifoData[342]));
Q_MX02 U7793 ( .S(n281), .A0(n2402), .A1(ofifoData[342]), .Z(n1476));
Q_FDP0UA U7794 ( .D(n1475), .QTFCLK( ), .Q(ofifoData[341]));
Q_MX02 U7795 ( .S(n281), .A0(n2403), .A1(ofifoData[341]), .Z(n1475));
Q_FDP0UA U7796 ( .D(n1474), .QTFCLK( ), .Q(ofifoData[340]));
Q_MX02 U7797 ( .S(n281), .A0(n2404), .A1(ofifoData[340]), .Z(n1474));
Q_FDP0UA U7798 ( .D(n1473), .QTFCLK( ), .Q(ofifoData[339]));
Q_MX02 U7799 ( .S(n281), .A0(n2405), .A1(ofifoData[339]), .Z(n1473));
Q_FDP0UA U7800 ( .D(n1472), .QTFCLK( ), .Q(ofifoData[338]));
Q_MX02 U7801 ( .S(n281), .A0(n2406), .A1(ofifoData[338]), .Z(n1472));
Q_FDP0UA U7802 ( .D(n1471), .QTFCLK( ), .Q(ofifoData[337]));
Q_MX02 U7803 ( .S(n281), .A0(n2407), .A1(ofifoData[337]), .Z(n1471));
Q_FDP0UA U7804 ( .D(n1470), .QTFCLK( ), .Q(ofifoData[336]));
Q_MX02 U7805 ( .S(n281), .A0(n2408), .A1(ofifoData[336]), .Z(n1470));
Q_FDP0UA U7806 ( .D(n1469), .QTFCLK( ), .Q(ofifoData[335]));
Q_MX02 U7807 ( .S(n281), .A0(n2409), .A1(ofifoData[335]), .Z(n1469));
Q_FDP0UA U7808 ( .D(n1468), .QTFCLK( ), .Q(ofifoData[334]));
Q_MX02 U7809 ( .S(n281), .A0(n2410), .A1(ofifoData[334]), .Z(n1468));
Q_FDP0UA U7810 ( .D(n1467), .QTFCLK( ), .Q(ofifoData[333]));
Q_MX02 U7811 ( .S(n281), .A0(n2411), .A1(ofifoData[333]), .Z(n1467));
Q_FDP0UA U7812 ( .D(n1466), .QTFCLK( ), .Q(ofifoData[332]));
Q_MX02 U7813 ( .S(n281), .A0(n2412), .A1(ofifoData[332]), .Z(n1466));
Q_FDP0UA U7814 ( .D(n1465), .QTFCLK( ), .Q(ofifoData[331]));
Q_MX02 U7815 ( .S(n281), .A0(n2413), .A1(ofifoData[331]), .Z(n1465));
Q_FDP0UA U7816 ( .D(n1464), .QTFCLK( ), .Q(ofifoData[330]));
Q_MX02 U7817 ( .S(n281), .A0(n2414), .A1(ofifoData[330]), .Z(n1464));
Q_FDP0UA U7818 ( .D(n1463), .QTFCLK( ), .Q(ofifoData[329]));
Q_MX02 U7819 ( .S(n281), .A0(n2415), .A1(ofifoData[329]), .Z(n1463));
Q_FDP0UA U7820 ( .D(n1462), .QTFCLK( ), .Q(ofifoData[328]));
Q_MX02 U7821 ( .S(n281), .A0(n2416), .A1(ofifoData[328]), .Z(n1462));
Q_FDP0UA U7822 ( .D(n1461), .QTFCLK( ), .Q(ofifoData[327]));
Q_MX02 U7823 ( .S(n281), .A0(n2417), .A1(ofifoData[327]), .Z(n1461));
Q_FDP0UA U7824 ( .D(n1460), .QTFCLK( ), .Q(ofifoData[326]));
Q_MX02 U7825 ( .S(n281), .A0(n2418), .A1(ofifoData[326]), .Z(n1460));
Q_FDP0UA U7826 ( .D(n1459), .QTFCLK( ), .Q(ofifoData[325]));
Q_MX02 U7827 ( .S(n281), .A0(n2419), .A1(ofifoData[325]), .Z(n1459));
Q_FDP0UA U7828 ( .D(n1458), .QTFCLK( ), .Q(ofifoData[324]));
Q_MX02 U7829 ( .S(n281), .A0(n2420), .A1(ofifoData[324]), .Z(n1458));
Q_FDP0UA U7830 ( .D(n1457), .QTFCLK( ), .Q(ofifoData[323]));
Q_MX02 U7831 ( .S(n281), .A0(n2421), .A1(ofifoData[323]), .Z(n1457));
Q_FDP0UA U7832 ( .D(n1456), .QTFCLK( ), .Q(ofifoData[322]));
Q_MX02 U7833 ( .S(n281), .A0(n2422), .A1(ofifoData[322]), .Z(n1456));
Q_FDP0UA U7834 ( .D(n1455), .QTFCLK( ), .Q(ofifoData[321]));
Q_MX02 U7835 ( .S(n281), .A0(n2423), .A1(ofifoData[321]), .Z(n1455));
Q_FDP0UA U7836 ( .D(n1454), .QTFCLK( ), .Q(ofifoData[320]));
Q_MX02 U7837 ( .S(n281), .A0(n2424), .A1(ofifoData[320]), .Z(n1454));
Q_FDP0UA U7838 ( .D(n1453), .QTFCLK( ), .Q(ofifoData[319]));
Q_MX02 U7839 ( .S(n281), .A0(n2425), .A1(ofifoData[319]), .Z(n1453));
Q_FDP0UA U7840 ( .D(n1452), .QTFCLK( ), .Q(ofifoData[318]));
Q_MX02 U7841 ( .S(n281), .A0(n2426), .A1(ofifoData[318]), .Z(n1452));
Q_FDP0UA U7842 ( .D(n1451), .QTFCLK( ), .Q(ofifoData[317]));
Q_MX02 U7843 ( .S(n281), .A0(n2427), .A1(ofifoData[317]), .Z(n1451));
Q_FDP0UA U7844 ( .D(n1450), .QTFCLK( ), .Q(ofifoData[316]));
Q_MX02 U7845 ( .S(n281), .A0(n2428), .A1(ofifoData[316]), .Z(n1450));
Q_FDP0UA U7846 ( .D(n1449), .QTFCLK( ), .Q(ofifoData[315]));
Q_MX02 U7847 ( .S(n281), .A0(n2429), .A1(ofifoData[315]), .Z(n1449));
Q_FDP0UA U7848 ( .D(n1448), .QTFCLK( ), .Q(ofifoData[314]));
Q_MX02 U7849 ( .S(n281), .A0(n2430), .A1(ofifoData[314]), .Z(n1448));
Q_FDP0UA U7850 ( .D(n1447), .QTFCLK( ), .Q(ofifoData[313]));
Q_MX02 U7851 ( .S(n281), .A0(n2431), .A1(ofifoData[313]), .Z(n1447));
Q_FDP0UA U7852 ( .D(n1446), .QTFCLK( ), .Q(ofifoData[312]));
Q_MX02 U7853 ( .S(n281), .A0(n2432), .A1(ofifoData[312]), .Z(n1446));
Q_FDP0UA U7854 ( .D(n1445), .QTFCLK( ), .Q(ofifoData[311]));
Q_MX02 U7855 ( .S(n281), .A0(n2433), .A1(ofifoData[311]), .Z(n1445));
Q_FDP0UA U7856 ( .D(n1444), .QTFCLK( ), .Q(ofifoData[310]));
Q_MX02 U7857 ( .S(n281), .A0(n2434), .A1(ofifoData[310]), .Z(n1444));
Q_FDP0UA U7858 ( .D(n1443), .QTFCLK( ), .Q(ofifoData[309]));
Q_MX02 U7859 ( .S(n281), .A0(n2435), .A1(ofifoData[309]), .Z(n1443));
Q_FDP0UA U7860 ( .D(n1442), .QTFCLK( ), .Q(ofifoData[308]));
Q_MX02 U7861 ( .S(n281), .A0(n2436), .A1(ofifoData[308]), .Z(n1442));
Q_FDP0UA U7862 ( .D(n1441), .QTFCLK( ), .Q(ofifoData[307]));
Q_MX02 U7863 ( .S(n281), .A0(n2437), .A1(ofifoData[307]), .Z(n1441));
Q_FDP0UA U7864 ( .D(n1440), .QTFCLK( ), .Q(ofifoData[306]));
Q_MX02 U7865 ( .S(n281), .A0(n2438), .A1(ofifoData[306]), .Z(n1440));
Q_FDP0UA U7866 ( .D(n1439), .QTFCLK( ), .Q(ofifoData[305]));
Q_MX02 U7867 ( .S(n281), .A0(n2439), .A1(ofifoData[305]), .Z(n1439));
Q_FDP0UA U7868 ( .D(n1438), .QTFCLK( ), .Q(ofifoData[304]));
Q_MX02 U7869 ( .S(n281), .A0(n2440), .A1(ofifoData[304]), .Z(n1438));
Q_FDP0UA U7870 ( .D(n1437), .QTFCLK( ), .Q(ofifoData[303]));
Q_MX02 U7871 ( .S(n281), .A0(n2441), .A1(ofifoData[303]), .Z(n1437));
Q_FDP0UA U7872 ( .D(n1436), .QTFCLK( ), .Q(ofifoData[302]));
Q_MX02 U7873 ( .S(n281), .A0(n2442), .A1(ofifoData[302]), .Z(n1436));
Q_FDP0UA U7874 ( .D(n1435), .QTFCLK( ), .Q(ofifoData[301]));
Q_MX02 U7875 ( .S(n281), .A0(n2443), .A1(ofifoData[301]), .Z(n1435));
Q_FDP0UA U7876 ( .D(n1434), .QTFCLK( ), .Q(ofifoData[300]));
Q_MX02 U7877 ( .S(n281), .A0(n2444), .A1(ofifoData[300]), .Z(n1434));
Q_FDP0UA U7878 ( .D(n1433), .QTFCLK( ), .Q(ofifoData[299]));
Q_MX02 U7879 ( .S(n281), .A0(n2445), .A1(ofifoData[299]), .Z(n1433));
Q_FDP0UA U7880 ( .D(n1432), .QTFCLK( ), .Q(ofifoData[298]));
Q_MX02 U7881 ( .S(n281), .A0(n2446), .A1(ofifoData[298]), .Z(n1432));
Q_FDP0UA U7882 ( .D(n1431), .QTFCLK( ), .Q(ofifoData[297]));
Q_MX02 U7883 ( .S(n281), .A0(n2447), .A1(ofifoData[297]), .Z(n1431));
Q_FDP0UA U7884 ( .D(n1430), .QTFCLK( ), .Q(ofifoData[296]));
Q_MX02 U7885 ( .S(n281), .A0(n2448), .A1(ofifoData[296]), .Z(n1430));
Q_FDP0UA U7886 ( .D(n1429), .QTFCLK( ), .Q(ofifoData[295]));
Q_MX02 U7887 ( .S(n281), .A0(n2449), .A1(ofifoData[295]), .Z(n1429));
Q_FDP0UA U7888 ( .D(n1428), .QTFCLK( ), .Q(ofifoData[294]));
Q_MX02 U7889 ( .S(n281), .A0(n2450), .A1(ofifoData[294]), .Z(n1428));
Q_FDP0UA U7890 ( .D(n1427), .QTFCLK( ), .Q(ofifoData[293]));
Q_MX02 U7891 ( .S(n281), .A0(n2451), .A1(ofifoData[293]), .Z(n1427));
Q_FDP0UA U7892 ( .D(n1426), .QTFCLK( ), .Q(ofifoData[292]));
Q_MX02 U7893 ( .S(n281), .A0(n2452), .A1(ofifoData[292]), .Z(n1426));
Q_FDP0UA U7894 ( .D(n1425), .QTFCLK( ), .Q(ofifoData[291]));
Q_MX02 U7895 ( .S(n281), .A0(n2453), .A1(ofifoData[291]), .Z(n1425));
Q_FDP0UA U7896 ( .D(n1424), .QTFCLK( ), .Q(ofifoData[290]));
Q_MX02 U7897 ( .S(n281), .A0(n2454), .A1(ofifoData[290]), .Z(n1424));
Q_FDP0UA U7898 ( .D(n1423), .QTFCLK( ), .Q(ofifoData[289]));
Q_MX02 U7899 ( .S(n281), .A0(n2455), .A1(ofifoData[289]), .Z(n1423));
Q_FDP0UA U7900 ( .D(n1422), .QTFCLK( ), .Q(ofifoData[288]));
Q_MX02 U7901 ( .S(n281), .A0(n2456), .A1(ofifoData[288]), .Z(n1422));
Q_FDP0UA U7902 ( .D(n1421), .QTFCLK( ), .Q(ofifoData[287]));
Q_MX02 U7903 ( .S(n281), .A0(n2457), .A1(ofifoData[287]), .Z(n1421));
Q_FDP0UA U7904 ( .D(n1420), .QTFCLK( ), .Q(ofifoData[286]));
Q_MX02 U7905 ( .S(n281), .A0(n2458), .A1(ofifoData[286]), .Z(n1420));
Q_FDP0UA U7906 ( .D(n1419), .QTFCLK( ), .Q(ofifoData[285]));
Q_MX02 U7907 ( .S(n281), .A0(n2459), .A1(ofifoData[285]), .Z(n1419));
Q_FDP0UA U7908 ( .D(n1418), .QTFCLK( ), .Q(ofifoData[284]));
Q_MX02 U7909 ( .S(n281), .A0(n2460), .A1(ofifoData[284]), .Z(n1418));
Q_FDP0UA U7910 ( .D(n1417), .QTFCLK( ), .Q(ofifoData[283]));
Q_MX02 U7911 ( .S(n281), .A0(n2461), .A1(ofifoData[283]), .Z(n1417));
Q_FDP0UA U7912 ( .D(n1416), .QTFCLK( ), .Q(ofifoData[282]));
Q_MX02 U7913 ( .S(n281), .A0(n2462), .A1(ofifoData[282]), .Z(n1416));
Q_FDP0UA U7914 ( .D(n1415), .QTFCLK( ), .Q(ofifoData[281]));
Q_MX02 U7915 ( .S(n281), .A0(n2463), .A1(ofifoData[281]), .Z(n1415));
Q_FDP0UA U7916 ( .D(n1414), .QTFCLK( ), .Q(ofifoData[280]));
Q_MX02 U7917 ( .S(n281), .A0(n2464), .A1(ofifoData[280]), .Z(n1414));
Q_FDP0UA U7918 ( .D(n1413), .QTFCLK( ), .Q(ofifoData[279]));
Q_MX02 U7919 ( .S(n281), .A0(n2465), .A1(ofifoData[279]), .Z(n1413));
Q_FDP0UA U7920 ( .D(n1412), .QTFCLK( ), .Q(ofifoData[278]));
Q_MX02 U7921 ( .S(n281), .A0(n2466), .A1(ofifoData[278]), .Z(n1412));
Q_FDP0UA U7922 ( .D(n1411), .QTFCLK( ), .Q(ofifoData[277]));
Q_MX02 U7923 ( .S(n281), .A0(n2467), .A1(ofifoData[277]), .Z(n1411));
Q_FDP0UA U7924 ( .D(n1410), .QTFCLK( ), .Q(ofifoData[276]));
Q_MX02 U7925 ( .S(n281), .A0(n2468), .A1(ofifoData[276]), .Z(n1410));
Q_FDP0UA U7926 ( .D(n1409), .QTFCLK( ), .Q(ofifoData[275]));
Q_MX02 U7927 ( .S(n281), .A0(n2469), .A1(ofifoData[275]), .Z(n1409));
Q_FDP0UA U7928 ( .D(n1408), .QTFCLK( ), .Q(ofifoData[274]));
Q_MX02 U7929 ( .S(n281), .A0(n2470), .A1(ofifoData[274]), .Z(n1408));
Q_FDP0UA U7930 ( .D(n1407), .QTFCLK( ), .Q(ofifoData[273]));
Q_MX02 U7931 ( .S(n281), .A0(n2471), .A1(ofifoData[273]), .Z(n1407));
Q_FDP0UA U7932 ( .D(n1406), .QTFCLK( ), .Q(ofifoData[272]));
Q_MX02 U7933 ( .S(n281), .A0(n2472), .A1(ofifoData[272]), .Z(n1406));
Q_FDP0UA U7934 ( .D(n1405), .QTFCLK( ), .Q(ofifoData[271]));
Q_MX02 U7935 ( .S(n281), .A0(n2473), .A1(ofifoData[271]), .Z(n1405));
Q_FDP0UA U7936 ( .D(n1404), .QTFCLK( ), .Q(ofifoData[270]));
Q_MX02 U7937 ( .S(n281), .A0(n2474), .A1(ofifoData[270]), .Z(n1404));
Q_FDP0UA U7938 ( .D(n1403), .QTFCLK( ), .Q(ofifoData[269]));
Q_MX02 U7939 ( .S(n281), .A0(n2475), .A1(ofifoData[269]), .Z(n1403));
Q_FDP0UA U7940 ( .D(n1402), .QTFCLK( ), .Q(ofifoData[268]));
Q_MX02 U7941 ( .S(n281), .A0(n2476), .A1(ofifoData[268]), .Z(n1402));
Q_FDP0UA U7942 ( .D(n1401), .QTFCLK( ), .Q(ofifoData[267]));
Q_MX02 U7943 ( .S(n281), .A0(n2477), .A1(ofifoData[267]), .Z(n1401));
Q_FDP0UA U7944 ( .D(n1400), .QTFCLK( ), .Q(ofifoData[266]));
Q_MX02 U7945 ( .S(n281), .A0(n2478), .A1(ofifoData[266]), .Z(n1400));
Q_FDP0UA U7946 ( .D(n1399), .QTFCLK( ), .Q(ofifoData[265]));
Q_MX02 U7947 ( .S(n281), .A0(n2479), .A1(ofifoData[265]), .Z(n1399));
Q_FDP0UA U7948 ( .D(n1398), .QTFCLK( ), .Q(ofifoData[264]));
Q_MX02 U7949 ( .S(n281), .A0(n2480), .A1(ofifoData[264]), .Z(n1398));
Q_FDP0UA U7950 ( .D(n1397), .QTFCLK( ), .Q(ofifoData[263]));
Q_MX02 U7951 ( .S(n281), .A0(n2481), .A1(ofifoData[263]), .Z(n1397));
Q_FDP0UA U7952 ( .D(n1396), .QTFCLK( ), .Q(ofifoData[262]));
Q_MX02 U7953 ( .S(n281), .A0(n2482), .A1(ofifoData[262]), .Z(n1396));
Q_FDP0UA U7954 ( .D(n1395), .QTFCLK( ), .Q(ofifoData[261]));
Q_MX02 U7955 ( .S(n281), .A0(n2483), .A1(ofifoData[261]), .Z(n1395));
Q_FDP0UA U7956 ( .D(n1394), .QTFCLK( ), .Q(ofifoData[260]));
Q_MX02 U7957 ( .S(n281), .A0(n2484), .A1(ofifoData[260]), .Z(n1394));
Q_FDP0UA U7958 ( .D(n1393), .QTFCLK( ), .Q(ofifoData[259]));
Q_MX02 U7959 ( .S(n281), .A0(n2485), .A1(ofifoData[259]), .Z(n1393));
Q_FDP0UA U7960 ( .D(n1392), .QTFCLK( ), .Q(ofifoData[258]));
Q_MX02 U7961 ( .S(n281), .A0(n2486), .A1(ofifoData[258]), .Z(n1392));
Q_FDP0UA U7962 ( .D(n1391), .QTFCLK( ), .Q(ofifoData[257]));
Q_MX02 U7963 ( .S(n281), .A0(n2487), .A1(ofifoData[257]), .Z(n1391));
Q_FDP0UA U7964 ( .D(n1390), .QTFCLK( ), .Q(ofifoData[256]));
Q_MX02 U7965 ( .S(n281), .A0(n2488), .A1(ofifoData[256]), .Z(n1390));
Q_FDP0UA U7966 ( .D(n1389), .QTFCLK( ), .Q(ofifoData[255]));
Q_MX02 U7967 ( .S(n281), .A0(n2489), .A1(ofifoData[255]), .Z(n1389));
Q_FDP0UA U7968 ( .D(n1388), .QTFCLK( ), .Q(ofifoData[254]));
Q_MX02 U7969 ( .S(n281), .A0(n2492), .A1(ofifoData[254]), .Z(n1388));
Q_FDP0UA U7970 ( .D(n1387), .QTFCLK( ), .Q(ofifoData[253]));
Q_MX02 U7971 ( .S(n281), .A0(n2495), .A1(ofifoData[253]), .Z(n1387));
Q_FDP0UA U7972 ( .D(n1386), .QTFCLK( ), .Q(ofifoData[252]));
Q_MX02 U7973 ( .S(n281), .A0(n2498), .A1(ofifoData[252]), .Z(n1386));
Q_FDP0UA U7974 ( .D(n1385), .QTFCLK( ), .Q(ofifoData[251]));
Q_MX02 U7975 ( .S(n281), .A0(n2501), .A1(ofifoData[251]), .Z(n1385));
Q_FDP0UA U7976 ( .D(n1384), .QTFCLK( ), .Q(ofifoData[250]));
Q_MX02 U7977 ( .S(n281), .A0(n2504), .A1(ofifoData[250]), .Z(n1384));
Q_FDP0UA U7978 ( .D(n1383), .QTFCLK( ), .Q(ofifoData[249]));
Q_MX02 U7979 ( .S(n281), .A0(n2507), .A1(ofifoData[249]), .Z(n1383));
Q_FDP0UA U7980 ( .D(n1382), .QTFCLK( ), .Q(ofifoData[248]));
Q_MX02 U7981 ( .S(n281), .A0(n2510), .A1(ofifoData[248]), .Z(n1382));
Q_FDP0UA U7982 ( .D(n1381), .QTFCLK( ), .Q(ofifoData[247]));
Q_MX02 U7983 ( .S(n281), .A0(n2513), .A1(ofifoData[247]), .Z(n1381));
Q_FDP0UA U7984 ( .D(n1380), .QTFCLK( ), .Q(ofifoData[246]));
Q_MX02 U7985 ( .S(n281), .A0(n2516), .A1(ofifoData[246]), .Z(n1380));
Q_FDP0UA U7986 ( .D(n1379), .QTFCLK( ), .Q(ofifoData[245]));
Q_MX02 U7987 ( .S(n281), .A0(n2519), .A1(ofifoData[245]), .Z(n1379));
Q_FDP0UA U7988 ( .D(n1378), .QTFCLK( ), .Q(ofifoData[244]));
Q_MX02 U7989 ( .S(n281), .A0(n2522), .A1(ofifoData[244]), .Z(n1378));
Q_FDP0UA U7990 ( .D(n1377), .QTFCLK( ), .Q(ofifoData[243]));
Q_MX02 U7991 ( .S(n281), .A0(n2525), .A1(ofifoData[243]), .Z(n1377));
Q_FDP0UA U7992 ( .D(n1376), .QTFCLK( ), .Q(ofifoData[242]));
Q_MX02 U7993 ( .S(n281), .A0(n2528), .A1(ofifoData[242]), .Z(n1376));
Q_FDP0UA U7994 ( .D(n1375), .QTFCLK( ), .Q(ofifoData[241]));
Q_MX02 U7995 ( .S(n281), .A0(n2531), .A1(ofifoData[241]), .Z(n1375));
Q_FDP0UA U7996 ( .D(n1374), .QTFCLK( ), .Q(ofifoData[240]));
Q_MX02 U7997 ( .S(n281), .A0(n2534), .A1(ofifoData[240]), .Z(n1374));
Q_FDP0UA U7998 ( .D(n1373), .QTFCLK( ), .Q(ofifoData[239]));
Q_MX02 U7999 ( .S(n281), .A0(n2537), .A1(ofifoData[239]), .Z(n1373));
Q_FDP0UA U8000 ( .D(n1372), .QTFCLK( ), .Q(ofifoData[238]));
Q_MX02 U8001 ( .S(n281), .A0(n2540), .A1(ofifoData[238]), .Z(n1372));
Q_FDP0UA U8002 ( .D(n1371), .QTFCLK( ), .Q(ofifoData[237]));
Q_MX02 U8003 ( .S(n281), .A0(n2543), .A1(ofifoData[237]), .Z(n1371));
Q_FDP0UA U8004 ( .D(n1370), .QTFCLK( ), .Q(ofifoData[236]));
Q_MX02 U8005 ( .S(n281), .A0(n2546), .A1(ofifoData[236]), .Z(n1370));
Q_FDP0UA U8006 ( .D(n1369), .QTFCLK( ), .Q(ofifoData[235]));
Q_MX02 U8007 ( .S(n281), .A0(n2549), .A1(ofifoData[235]), .Z(n1369));
Q_FDP0UA U8008 ( .D(n1368), .QTFCLK( ), .Q(ofifoData[234]));
Q_MX02 U8009 ( .S(n281), .A0(n2552), .A1(ofifoData[234]), .Z(n1368));
Q_FDP0UA U8010 ( .D(n1367), .QTFCLK( ), .Q(ofifoData[233]));
Q_MX02 U8011 ( .S(n281), .A0(n2555), .A1(ofifoData[233]), .Z(n1367));
Q_FDP0UA U8012 ( .D(n1366), .QTFCLK( ), .Q(ofifoData[232]));
Q_MX02 U8013 ( .S(n281), .A0(n2558), .A1(ofifoData[232]), .Z(n1366));
Q_FDP0UA U8014 ( .D(n1365), .QTFCLK( ), .Q(ofifoData[231]));
Q_MX02 U8015 ( .S(n281), .A0(n2561), .A1(ofifoData[231]), .Z(n1365));
Q_FDP0UA U8016 ( .D(n1364), .QTFCLK( ), .Q(ofifoData[230]));
Q_MX02 U8017 ( .S(n281), .A0(n2564), .A1(ofifoData[230]), .Z(n1364));
Q_FDP0UA U8018 ( .D(n1363), .QTFCLK( ), .Q(ofifoData[229]));
Q_MX02 U8019 ( .S(n281), .A0(n2567), .A1(ofifoData[229]), .Z(n1363));
Q_FDP0UA U8020 ( .D(n1362), .QTFCLK( ), .Q(ofifoData[228]));
Q_MX02 U8021 ( .S(n281), .A0(n2570), .A1(ofifoData[228]), .Z(n1362));
Q_FDP0UA U8022 ( .D(n1361), .QTFCLK( ), .Q(ofifoData[227]));
Q_MX02 U8023 ( .S(n281), .A0(n2573), .A1(ofifoData[227]), .Z(n1361));
Q_FDP0UA U8024 ( .D(n1360), .QTFCLK( ), .Q(ofifoData[226]));
Q_MX02 U8025 ( .S(n281), .A0(n2576), .A1(ofifoData[226]), .Z(n1360));
Q_FDP0UA U8026 ( .D(n1359), .QTFCLK( ), .Q(ofifoData[225]));
Q_MX02 U8027 ( .S(n281), .A0(n2579), .A1(ofifoData[225]), .Z(n1359));
Q_FDP0UA U8028 ( .D(n1358), .QTFCLK( ), .Q(ofifoData[224]));
Q_MX02 U8029 ( .S(n281), .A0(n2582), .A1(ofifoData[224]), .Z(n1358));
Q_FDP0UA U8030 ( .D(n1357), .QTFCLK( ), .Q(ofifoData[223]));
Q_MX02 U8031 ( .S(n281), .A0(n2585), .A1(ofifoData[223]), .Z(n1357));
Q_FDP0UA U8032 ( .D(n1356), .QTFCLK( ), .Q(ofifoData[222]));
Q_MX02 U8033 ( .S(n281), .A0(n2588), .A1(ofifoData[222]), .Z(n1356));
Q_FDP0UA U8034 ( .D(n1355), .QTFCLK( ), .Q(ofifoData[221]));
Q_MX02 U8035 ( .S(n281), .A0(n2591), .A1(ofifoData[221]), .Z(n1355));
Q_FDP0UA U8036 ( .D(n1354), .QTFCLK( ), .Q(ofifoData[220]));
Q_MX02 U8037 ( .S(n281), .A0(n2594), .A1(ofifoData[220]), .Z(n1354));
Q_FDP0UA U8038 ( .D(n1353), .QTFCLK( ), .Q(ofifoData[219]));
Q_MX02 U8039 ( .S(n281), .A0(n2597), .A1(ofifoData[219]), .Z(n1353));
Q_FDP0UA U8040 ( .D(n1352), .QTFCLK( ), .Q(ofifoData[218]));
Q_MX02 U8041 ( .S(n281), .A0(n2600), .A1(ofifoData[218]), .Z(n1352));
Q_FDP0UA U8042 ( .D(n1351), .QTFCLK( ), .Q(ofifoData[217]));
Q_MX02 U8043 ( .S(n281), .A0(n2603), .A1(ofifoData[217]), .Z(n1351));
Q_FDP0UA U8044 ( .D(n1350), .QTFCLK( ), .Q(ofifoData[216]));
Q_MX02 U8045 ( .S(n281), .A0(n2606), .A1(ofifoData[216]), .Z(n1350));
Q_FDP0UA U8046 ( .D(n1349), .QTFCLK( ), .Q(ofifoData[215]));
Q_MX02 U8047 ( .S(n281), .A0(n2609), .A1(ofifoData[215]), .Z(n1349));
Q_FDP0UA U8048 ( .D(n1348), .QTFCLK( ), .Q(ofifoData[214]));
Q_MX02 U8049 ( .S(n281), .A0(n2612), .A1(ofifoData[214]), .Z(n1348));
Q_FDP0UA U8050 ( .D(n1347), .QTFCLK( ), .Q(ofifoData[213]));
Q_MX02 U8051 ( .S(n281), .A0(n2615), .A1(ofifoData[213]), .Z(n1347));
Q_FDP0UA U8052 ( .D(n1346), .QTFCLK( ), .Q(ofifoData[212]));
Q_MX02 U8053 ( .S(n281), .A0(n2618), .A1(ofifoData[212]), .Z(n1346));
Q_FDP0UA U8054 ( .D(n1345), .QTFCLK( ), .Q(ofifoData[211]));
Q_MX02 U8055 ( .S(n281), .A0(n2621), .A1(ofifoData[211]), .Z(n1345));
Q_FDP0UA U8056 ( .D(n1344), .QTFCLK( ), .Q(ofifoData[210]));
Q_MX02 U8057 ( .S(n281), .A0(n2624), .A1(ofifoData[210]), .Z(n1344));
Q_FDP0UA U8058 ( .D(n1343), .QTFCLK( ), .Q(ofifoData[209]));
Q_MX02 U8059 ( .S(n281), .A0(n2627), .A1(ofifoData[209]), .Z(n1343));
Q_FDP0UA U8060 ( .D(n1342), .QTFCLK( ), .Q(ofifoData[208]));
Q_MX02 U8061 ( .S(n281), .A0(n2630), .A1(ofifoData[208]), .Z(n1342));
Q_FDP0UA U8062 ( .D(n1341), .QTFCLK( ), .Q(ofifoData[207]));
Q_MX02 U8063 ( .S(n281), .A0(n2633), .A1(ofifoData[207]), .Z(n1341));
Q_FDP0UA U8064 ( .D(n1340), .QTFCLK( ), .Q(ofifoData[206]));
Q_MX02 U8065 ( .S(n281), .A0(n2636), .A1(ofifoData[206]), .Z(n1340));
Q_FDP0UA U8066 ( .D(n1339), .QTFCLK( ), .Q(ofifoData[205]));
Q_MX02 U8067 ( .S(n281), .A0(n2639), .A1(ofifoData[205]), .Z(n1339));
Q_FDP0UA U8068 ( .D(n1338), .QTFCLK( ), .Q(ofifoData[204]));
Q_MX02 U8069 ( .S(n281), .A0(n2642), .A1(ofifoData[204]), .Z(n1338));
Q_FDP0UA U8070 ( .D(n1337), .QTFCLK( ), .Q(ofifoData[203]));
Q_MX02 U8071 ( .S(n281), .A0(n2645), .A1(ofifoData[203]), .Z(n1337));
Q_FDP0UA U8072 ( .D(n1336), .QTFCLK( ), .Q(ofifoData[202]));
Q_MX02 U8073 ( .S(n281), .A0(n2648), .A1(ofifoData[202]), .Z(n1336));
Q_FDP0UA U8074 ( .D(n1335), .QTFCLK( ), .Q(ofifoData[201]));
Q_MX02 U8075 ( .S(n281), .A0(n2651), .A1(ofifoData[201]), .Z(n1335));
Q_FDP0UA U8076 ( .D(n1334), .QTFCLK( ), .Q(ofifoData[200]));
Q_MX02 U8077 ( .S(n281), .A0(n2654), .A1(ofifoData[200]), .Z(n1334));
Q_FDP0UA U8078 ( .D(n1333), .QTFCLK( ), .Q(ofifoData[199]));
Q_MX02 U8079 ( .S(n281), .A0(n2657), .A1(ofifoData[199]), .Z(n1333));
Q_FDP0UA U8080 ( .D(n1332), .QTFCLK( ), .Q(ofifoData[198]));
Q_MX02 U8081 ( .S(n281), .A0(n2660), .A1(ofifoData[198]), .Z(n1332));
Q_FDP0UA U8082 ( .D(n1331), .QTFCLK( ), .Q(ofifoData[197]));
Q_MX02 U8083 ( .S(n281), .A0(n2663), .A1(ofifoData[197]), .Z(n1331));
Q_FDP0UA U8084 ( .D(n1330), .QTFCLK( ), .Q(ofifoData[196]));
Q_MX02 U8085 ( .S(n281), .A0(n2666), .A1(ofifoData[196]), .Z(n1330));
Q_FDP0UA U8086 ( .D(n1329), .QTFCLK( ), .Q(ofifoData[195]));
Q_MX02 U8087 ( .S(n281), .A0(n2669), .A1(ofifoData[195]), .Z(n1329));
Q_FDP0UA U8088 ( .D(n1328), .QTFCLK( ), .Q(ofifoData[194]));
Q_MX02 U8089 ( .S(n281), .A0(n2672), .A1(ofifoData[194]), .Z(n1328));
Q_FDP0UA U8090 ( .D(n1327), .QTFCLK( ), .Q(ofifoData[193]));
Q_MX02 U8091 ( .S(n281), .A0(n2675), .A1(ofifoData[193]), .Z(n1327));
Q_FDP0UA U8092 ( .D(n1326), .QTFCLK( ), .Q(ofifoData[192]));
Q_MX02 U8093 ( .S(n281), .A0(n2678), .A1(ofifoData[192]), .Z(n1326));
Q_FDP0UA U8094 ( .D(n1325), .QTFCLK( ), .Q(ofifoData[191]));
Q_MX02 U8095 ( .S(n281), .A0(n2681), .A1(ofifoData[191]), .Z(n1325));
Q_FDP0UA U8096 ( .D(n1324), .QTFCLK( ), .Q(ofifoData[190]));
Q_MX02 U8097 ( .S(n281), .A0(n2684), .A1(ofifoData[190]), .Z(n1324));
Q_FDP0UA U8098 ( .D(n1323), .QTFCLK( ), .Q(ofifoData[189]));
Q_MX02 U8099 ( .S(n281), .A0(n2687), .A1(ofifoData[189]), .Z(n1323));
Q_FDP0UA U8100 ( .D(n1322), .QTFCLK( ), .Q(ofifoData[188]));
Q_MX02 U8101 ( .S(n281), .A0(n2690), .A1(ofifoData[188]), .Z(n1322));
Q_FDP0UA U8102 ( .D(n1321), .QTFCLK( ), .Q(ofifoData[187]));
Q_MX02 U8103 ( .S(n281), .A0(n2693), .A1(ofifoData[187]), .Z(n1321));
Q_FDP0UA U8104 ( .D(n1320), .QTFCLK( ), .Q(ofifoData[186]));
Q_MX02 U8105 ( .S(n281), .A0(n2696), .A1(ofifoData[186]), .Z(n1320));
Q_FDP0UA U8106 ( .D(n1319), .QTFCLK( ), .Q(ofifoData[185]));
Q_MX02 U8107 ( .S(n281), .A0(n2699), .A1(ofifoData[185]), .Z(n1319));
Q_FDP0UA U8108 ( .D(n1318), .QTFCLK( ), .Q(ofifoData[184]));
Q_MX02 U8109 ( .S(n281), .A0(n2702), .A1(ofifoData[184]), .Z(n1318));
Q_FDP0UA U8110 ( .D(n1317), .QTFCLK( ), .Q(ofifoData[183]));
Q_MX02 U8111 ( .S(n281), .A0(n2705), .A1(ofifoData[183]), .Z(n1317));
Q_FDP0UA U8112 ( .D(n1316), .QTFCLK( ), .Q(ofifoData[182]));
Q_MX02 U8113 ( .S(n281), .A0(n2708), .A1(ofifoData[182]), .Z(n1316));
Q_FDP0UA U8114 ( .D(n1315), .QTFCLK( ), .Q(ofifoData[181]));
Q_MX02 U8115 ( .S(n281), .A0(n2711), .A1(ofifoData[181]), .Z(n1315));
Q_FDP0UA U8116 ( .D(n1314), .QTFCLK( ), .Q(ofifoData[180]));
Q_MX02 U8117 ( .S(n281), .A0(n2714), .A1(ofifoData[180]), .Z(n1314));
Q_FDP0UA U8118 ( .D(n1313), .QTFCLK( ), .Q(ofifoData[179]));
Q_MX02 U8119 ( .S(n281), .A0(n2717), .A1(ofifoData[179]), .Z(n1313));
Q_FDP0UA U8120 ( .D(n1312), .QTFCLK( ), .Q(ofifoData[178]));
Q_MX02 U8121 ( .S(n281), .A0(n2720), .A1(ofifoData[178]), .Z(n1312));
Q_FDP0UA U8122 ( .D(n1311), .QTFCLK( ), .Q(ofifoData[177]));
Q_MX02 U8123 ( .S(n281), .A0(n2723), .A1(ofifoData[177]), .Z(n1311));
Q_FDP0UA U8124 ( .D(n1310), .QTFCLK( ), .Q(ofifoData[176]));
Q_MX02 U8125 ( .S(n281), .A0(n2726), .A1(ofifoData[176]), .Z(n1310));
Q_FDP0UA U8126 ( .D(n1309), .QTFCLK( ), .Q(ofifoData[175]));
Q_MX02 U8127 ( .S(n281), .A0(n2729), .A1(ofifoData[175]), .Z(n1309));
Q_FDP0UA U8128 ( .D(n1308), .QTFCLK( ), .Q(ofifoData[174]));
Q_MX02 U8129 ( .S(n281), .A0(n2732), .A1(ofifoData[174]), .Z(n1308));
Q_FDP0UA U8130 ( .D(n1307), .QTFCLK( ), .Q(ofifoData[173]));
Q_MX02 U8131 ( .S(n281), .A0(n2735), .A1(ofifoData[173]), .Z(n1307));
Q_FDP0UA U8132 ( .D(n1306), .QTFCLK( ), .Q(ofifoData[172]));
Q_MX02 U8133 ( .S(n281), .A0(n2738), .A1(ofifoData[172]), .Z(n1306));
Q_FDP0UA U8134 ( .D(n1305), .QTFCLK( ), .Q(ofifoData[171]));
Q_MX02 U8135 ( .S(n281), .A0(n2741), .A1(ofifoData[171]), .Z(n1305));
Q_FDP0UA U8136 ( .D(n1304), .QTFCLK( ), .Q(ofifoData[170]));
Q_MX02 U8137 ( .S(n281), .A0(n2744), .A1(ofifoData[170]), .Z(n1304));
Q_FDP0UA U8138 ( .D(n1303), .QTFCLK( ), .Q(ofifoData[169]));
Q_MX02 U8139 ( .S(n281), .A0(n2747), .A1(ofifoData[169]), .Z(n1303));
Q_FDP0UA U8140 ( .D(n1302), .QTFCLK( ), .Q(ofifoData[168]));
Q_MX02 U8141 ( .S(n281), .A0(n2750), .A1(ofifoData[168]), .Z(n1302));
Q_FDP0UA U8142 ( .D(n1301), .QTFCLK( ), .Q(ofifoData[167]));
Q_MX02 U8143 ( .S(n281), .A0(n2753), .A1(ofifoData[167]), .Z(n1301));
Q_FDP0UA U8144 ( .D(n1300), .QTFCLK( ), .Q(ofifoData[166]));
Q_MX02 U8145 ( .S(n281), .A0(n2756), .A1(ofifoData[166]), .Z(n1300));
Q_FDP0UA U8146 ( .D(n1299), .QTFCLK( ), .Q(ofifoData[165]));
Q_MX02 U8147 ( .S(n281), .A0(n2759), .A1(ofifoData[165]), .Z(n1299));
Q_FDP0UA U8148 ( .D(n1298), .QTFCLK( ), .Q(ofifoData[164]));
Q_MX02 U8149 ( .S(n281), .A0(n2762), .A1(ofifoData[164]), .Z(n1298));
Q_FDP0UA U8150 ( .D(n1297), .QTFCLK( ), .Q(ofifoData[163]));
Q_MX02 U8151 ( .S(n281), .A0(n2765), .A1(ofifoData[163]), .Z(n1297));
Q_FDP0UA U8152 ( .D(n1296), .QTFCLK( ), .Q(ofifoData[162]));
Q_MX02 U8153 ( .S(n281), .A0(n2768), .A1(ofifoData[162]), .Z(n1296));
Q_FDP0UA U8154 ( .D(n1295), .QTFCLK( ), .Q(ofifoData[161]));
Q_MX02 U8155 ( .S(n281), .A0(n2771), .A1(ofifoData[161]), .Z(n1295));
Q_FDP0UA U8156 ( .D(n1294), .QTFCLK( ), .Q(ofifoData[160]));
Q_MX02 U8157 ( .S(n281), .A0(n2774), .A1(ofifoData[160]), .Z(n1294));
Q_FDP0UA U8158 ( .D(n1293), .QTFCLK( ), .Q(ofifoData[159]));
Q_MX02 U8159 ( .S(n281), .A0(n2777), .A1(ofifoData[159]), .Z(n1293));
Q_FDP0UA U8160 ( .D(n1292), .QTFCLK( ), .Q(ofifoData[158]));
Q_MX02 U8161 ( .S(n281), .A0(n2780), .A1(ofifoData[158]), .Z(n1292));
Q_FDP0UA U8162 ( .D(n1291), .QTFCLK( ), .Q(ofifoData[157]));
Q_MX02 U8163 ( .S(n281), .A0(n2783), .A1(ofifoData[157]), .Z(n1291));
Q_FDP0UA U8164 ( .D(n1290), .QTFCLK( ), .Q(ofifoData[156]));
Q_MX02 U8165 ( .S(n281), .A0(n2786), .A1(ofifoData[156]), .Z(n1290));
Q_FDP0UA U8166 ( .D(n1289), .QTFCLK( ), .Q(ofifoData[155]));
Q_MX02 U8167 ( .S(n281), .A0(n2789), .A1(ofifoData[155]), .Z(n1289));
Q_FDP0UA U8168 ( .D(n1288), .QTFCLK( ), .Q(ofifoData[154]));
Q_MX02 U8169 ( .S(n281), .A0(n2792), .A1(ofifoData[154]), .Z(n1288));
Q_FDP0UA U8170 ( .D(n1287), .QTFCLK( ), .Q(ofifoData[153]));
Q_MX02 U8171 ( .S(n281), .A0(n2795), .A1(ofifoData[153]), .Z(n1287));
Q_FDP0UA U8172 ( .D(n1286), .QTFCLK( ), .Q(ofifoData[152]));
Q_MX02 U8173 ( .S(n281), .A0(n2798), .A1(ofifoData[152]), .Z(n1286));
Q_FDP0UA U8174 ( .D(n1285), .QTFCLK( ), .Q(ofifoData[151]));
Q_MX02 U8175 ( .S(n281), .A0(n2801), .A1(ofifoData[151]), .Z(n1285));
Q_FDP0UA U8176 ( .D(n1284), .QTFCLK( ), .Q(ofifoData[150]));
Q_MX02 U8177 ( .S(n281), .A0(n2804), .A1(ofifoData[150]), .Z(n1284));
Q_FDP0UA U8178 ( .D(n1283), .QTFCLK( ), .Q(ofifoData[149]));
Q_MX02 U8179 ( .S(n281), .A0(n2807), .A1(ofifoData[149]), .Z(n1283));
Q_FDP0UA U8180 ( .D(n1282), .QTFCLK( ), .Q(ofifoData[148]));
Q_MX02 U8181 ( .S(n281), .A0(n2810), .A1(ofifoData[148]), .Z(n1282));
Q_FDP0UA U8182 ( .D(n1281), .QTFCLK( ), .Q(ofifoData[147]));
Q_MX02 U8183 ( .S(n281), .A0(n2813), .A1(ofifoData[147]), .Z(n1281));
Q_FDP0UA U8184 ( .D(n1280), .QTFCLK( ), .Q(ofifoData[146]));
Q_MX02 U8185 ( .S(n281), .A0(n2816), .A1(ofifoData[146]), .Z(n1280));
Q_FDP0UA U8186 ( .D(n1279), .QTFCLK( ), .Q(ofifoData[145]));
Q_MX02 U8187 ( .S(n281), .A0(n2819), .A1(ofifoData[145]), .Z(n1279));
Q_FDP0UA U8188 ( .D(n1278), .QTFCLK( ), .Q(ofifoData[144]));
Q_MX02 U8189 ( .S(n281), .A0(n2822), .A1(ofifoData[144]), .Z(n1278));
Q_FDP0UA U8190 ( .D(n1277), .QTFCLK( ), .Q(ofifoData[143]));
Q_MX02 U8191 ( .S(n281), .A0(n2825), .A1(ofifoData[143]), .Z(n1277));
Q_FDP0UA U8192 ( .D(n1276), .QTFCLK( ), .Q(ofifoData[142]));
Q_MX02 U8193 ( .S(n281), .A0(n2828), .A1(ofifoData[142]), .Z(n1276));
Q_FDP0UA U8194 ( .D(n1275), .QTFCLK( ), .Q(ofifoData[141]));
Q_MX02 U8195 ( .S(n281), .A0(n2831), .A1(ofifoData[141]), .Z(n1275));
Q_FDP0UA U8196 ( .D(n1274), .QTFCLK( ), .Q(ofifoData[140]));
Q_MX02 U8197 ( .S(n281), .A0(n2834), .A1(ofifoData[140]), .Z(n1274));
Q_FDP0UA U8198 ( .D(n1273), .QTFCLK( ), .Q(ofifoData[139]));
Q_MX02 U8199 ( .S(n281), .A0(n2837), .A1(ofifoData[139]), .Z(n1273));
Q_FDP0UA U8200 ( .D(n1272), .QTFCLK( ), .Q(ofifoData[138]));
Q_MX02 U8201 ( .S(n281), .A0(n2840), .A1(ofifoData[138]), .Z(n1272));
Q_FDP0UA U8202 ( .D(n1271), .QTFCLK( ), .Q(ofifoData[137]));
Q_MX02 U8203 ( .S(n281), .A0(n2843), .A1(ofifoData[137]), .Z(n1271));
Q_FDP0UA U8204 ( .D(n1270), .QTFCLK( ), .Q(ofifoData[136]));
Q_MX02 U8205 ( .S(n281), .A0(n2846), .A1(ofifoData[136]), .Z(n1270));
Q_FDP0UA U8206 ( .D(n1269), .QTFCLK( ), .Q(ofifoData[135]));
Q_MX02 U8207 ( .S(n281), .A0(n2849), .A1(ofifoData[135]), .Z(n1269));
Q_FDP0UA U8208 ( .D(n1268), .QTFCLK( ), .Q(ofifoData[134]));
Q_MX02 U8209 ( .S(n281), .A0(n2852), .A1(ofifoData[134]), .Z(n1268));
Q_FDP0UA U8210 ( .D(n1267), .QTFCLK( ), .Q(ofifoData[133]));
Q_MX02 U8211 ( .S(n281), .A0(n2855), .A1(ofifoData[133]), .Z(n1267));
Q_FDP0UA U8212 ( .D(n1266), .QTFCLK( ), .Q(ofifoData[132]));
Q_MX02 U8213 ( .S(n281), .A0(n2858), .A1(ofifoData[132]), .Z(n1266));
Q_FDP0UA U8214 ( .D(n1265), .QTFCLK( ), .Q(ofifoData[131]));
Q_MX02 U8215 ( .S(n281), .A0(n2861), .A1(ofifoData[131]), .Z(n1265));
Q_FDP0UA U8216 ( .D(n1264), .QTFCLK( ), .Q(ofifoData[130]));
Q_MX02 U8217 ( .S(n281), .A0(n2864), .A1(ofifoData[130]), .Z(n1264));
Q_FDP0UA U8218 ( .D(n1263), .QTFCLK( ), .Q(ofifoData[129]));
Q_MX02 U8219 ( .S(n281), .A0(n2867), .A1(ofifoData[129]), .Z(n1263));
Q_FDP0UA U8220 ( .D(n1262), .QTFCLK( ), .Q(ofifoData[128]));
Q_MX02 U8221 ( .S(n281), .A0(n2870), .A1(ofifoData[128]), .Z(n1262));
Q_FDP0UA U8222 ( .D(n1261), .QTFCLK( ), .Q(ofifoData[127]));
Q_MX02 U8223 ( .S(n281), .A0(n2873), .A1(ofifoData[127]), .Z(n1261));
Q_FDP0UA U8224 ( .D(n1260), .QTFCLK( ), .Q(ofifoData[126]));
Q_MX02 U8225 ( .S(n281), .A0(n2876), .A1(ofifoData[126]), .Z(n1260));
Q_FDP0UA U8226 ( .D(n1259), .QTFCLK( ), .Q(ofifoData[125]));
Q_MX02 U8227 ( .S(n281), .A0(n2879), .A1(ofifoData[125]), .Z(n1259));
Q_FDP0UA U8228 ( .D(n1258), .QTFCLK( ), .Q(ofifoData[124]));
Q_MX02 U8229 ( .S(n281), .A0(n2882), .A1(ofifoData[124]), .Z(n1258));
Q_FDP0UA U8230 ( .D(n1257), .QTFCLK( ), .Q(ofifoData[123]));
Q_MX02 U8231 ( .S(n281), .A0(n2885), .A1(ofifoData[123]), .Z(n1257));
Q_FDP0UA U8232 ( .D(n1256), .QTFCLK( ), .Q(ofifoData[122]));
Q_MX02 U8233 ( .S(n281), .A0(n2888), .A1(ofifoData[122]), .Z(n1256));
Q_FDP0UA U8234 ( .D(n1255), .QTFCLK( ), .Q(ofifoData[121]));
Q_MX02 U8235 ( .S(n281), .A0(n2891), .A1(ofifoData[121]), .Z(n1255));
Q_FDP0UA U8236 ( .D(n1254), .QTFCLK( ), .Q(ofifoData[120]));
Q_MX02 U8237 ( .S(n281), .A0(n2894), .A1(ofifoData[120]), .Z(n1254));
Q_FDP0UA U8238 ( .D(n1253), .QTFCLK( ), .Q(ofifoData[119]));
Q_MX02 U8239 ( .S(n281), .A0(n2897), .A1(ofifoData[119]), .Z(n1253));
Q_FDP0UA U8240 ( .D(n1252), .QTFCLK( ), .Q(ofifoData[118]));
Q_MX02 U8241 ( .S(n281), .A0(n2900), .A1(ofifoData[118]), .Z(n1252));
Q_FDP0UA U8242 ( .D(n1251), .QTFCLK( ), .Q(ofifoData[117]));
Q_MX02 U8243 ( .S(n281), .A0(n2903), .A1(ofifoData[117]), .Z(n1251));
Q_FDP0UA U8244 ( .D(n1250), .QTFCLK( ), .Q(ofifoData[116]));
Q_MX02 U8245 ( .S(n281), .A0(n2906), .A1(ofifoData[116]), .Z(n1250));
Q_FDP0UA U8246 ( .D(n1249), .QTFCLK( ), .Q(ofifoData[115]));
Q_MX02 U8247 ( .S(n281), .A0(n2909), .A1(ofifoData[115]), .Z(n1249));
Q_FDP0UA U8248 ( .D(n1248), .QTFCLK( ), .Q(ofifoData[114]));
Q_MX02 U8249 ( .S(n281), .A0(n2912), .A1(ofifoData[114]), .Z(n1248));
Q_FDP0UA U8250 ( .D(n1247), .QTFCLK( ), .Q(ofifoData[113]));
Q_MX02 U8251 ( .S(n281), .A0(n2915), .A1(ofifoData[113]), .Z(n1247));
Q_FDP0UA U8252 ( .D(n1246), .QTFCLK( ), .Q(ofifoData[112]));
Q_MX02 U8253 ( .S(n281), .A0(n2918), .A1(ofifoData[112]), .Z(n1246));
Q_FDP0UA U8254 ( .D(n1245), .QTFCLK( ), .Q(ofifoData[111]));
Q_MX02 U8255 ( .S(n281), .A0(n2921), .A1(ofifoData[111]), .Z(n1245));
Q_FDP0UA U8256 ( .D(n1244), .QTFCLK( ), .Q(ofifoData[110]));
Q_MX02 U8257 ( .S(n281), .A0(n2924), .A1(ofifoData[110]), .Z(n1244));
Q_FDP0UA U8258 ( .D(n1243), .QTFCLK( ), .Q(ofifoData[109]));
Q_MX02 U8259 ( .S(n281), .A0(n2927), .A1(ofifoData[109]), .Z(n1243));
Q_FDP0UA U8260 ( .D(n1242), .QTFCLK( ), .Q(ofifoData[108]));
Q_MX02 U8261 ( .S(n281), .A0(n2930), .A1(ofifoData[108]), .Z(n1242));
Q_FDP0UA U8262 ( .D(n1241), .QTFCLK( ), .Q(ofifoData[107]));
Q_MX02 U8263 ( .S(n281), .A0(n2933), .A1(ofifoData[107]), .Z(n1241));
Q_FDP0UA U8264 ( .D(n1240), .QTFCLK( ), .Q(ofifoData[106]));
Q_MX02 U8265 ( .S(n281), .A0(n2936), .A1(ofifoData[106]), .Z(n1240));
Q_FDP0UA U8266 ( .D(n1239), .QTFCLK( ), .Q(ofifoData[105]));
Q_MX02 U8267 ( .S(n281), .A0(n2939), .A1(ofifoData[105]), .Z(n1239));
Q_FDP0UA U8268 ( .D(n1238), .QTFCLK( ), .Q(ofifoData[104]));
Q_MX02 U8269 ( .S(n281), .A0(n2942), .A1(ofifoData[104]), .Z(n1238));
Q_FDP0UA U8270 ( .D(n1237), .QTFCLK( ), .Q(ofifoData[103]));
Q_MX02 U8271 ( .S(n281), .A0(n2945), .A1(ofifoData[103]), .Z(n1237));
Q_FDP0UA U8272 ( .D(n1236), .QTFCLK( ), .Q(ofifoData[102]));
Q_MX02 U8273 ( .S(n281), .A0(n2948), .A1(ofifoData[102]), .Z(n1236));
Q_FDP0UA U8274 ( .D(n1235), .QTFCLK( ), .Q(ofifoData[101]));
Q_MX02 U8275 ( .S(n281), .A0(n2951), .A1(ofifoData[101]), .Z(n1235));
Q_FDP0UA U8276 ( .D(n1234), .QTFCLK( ), .Q(ofifoData[100]));
Q_MX02 U8277 ( .S(n281), .A0(n2954), .A1(ofifoData[100]), .Z(n1234));
Q_FDP0UA U8278 ( .D(n1233), .QTFCLK( ), .Q(ofifoData[99]));
Q_MX02 U8279 ( .S(n281), .A0(n2957), .A1(ofifoData[99]), .Z(n1233));
Q_FDP0UA U8280 ( .D(n1232), .QTFCLK( ), .Q(ofifoData[98]));
Q_MX02 U8281 ( .S(n281), .A0(n2960), .A1(ofifoData[98]), .Z(n1232));
Q_FDP0UA U8282 ( .D(n1231), .QTFCLK( ), .Q(ofifoData[97]));
Q_MX02 U8283 ( .S(n281), .A0(n2963), .A1(ofifoData[97]), .Z(n1231));
Q_FDP0UA U8284 ( .D(n1230), .QTFCLK( ), .Q(ofifoData[96]));
Q_MX02 U8285 ( .S(n281), .A0(n2966), .A1(ofifoData[96]), .Z(n1230));
Q_FDP0UA U8286 ( .D(n1229), .QTFCLK( ), .Q(ofifoData[95]));
Q_MX02 U8287 ( .S(n281), .A0(n2969), .A1(ofifoData[95]), .Z(n1229));
Q_FDP0UA U8288 ( .D(n1228), .QTFCLK( ), .Q(ofifoData[94]));
Q_MX02 U8289 ( .S(n281), .A0(n2972), .A1(ofifoData[94]), .Z(n1228));
Q_FDP0UA U8290 ( .D(n1227), .QTFCLK( ), .Q(ofifoData[93]));
Q_MX02 U8291 ( .S(n281), .A0(n2975), .A1(ofifoData[93]), .Z(n1227));
Q_FDP0UA U8292 ( .D(n1226), .QTFCLK( ), .Q(ofifoData[92]));
Q_MX02 U8293 ( .S(n281), .A0(n2978), .A1(ofifoData[92]), .Z(n1226));
Q_FDP0UA U8294 ( .D(n1225), .QTFCLK( ), .Q(ofifoData[91]));
Q_MX02 U8295 ( .S(n281), .A0(n2981), .A1(ofifoData[91]), .Z(n1225));
Q_FDP0UA U8296 ( .D(n1224), .QTFCLK( ), .Q(ofifoData[90]));
Q_MX02 U8297 ( .S(n281), .A0(n2984), .A1(ofifoData[90]), .Z(n1224));
Q_FDP0UA U8298 ( .D(n1223), .QTFCLK( ), .Q(ofifoData[89]));
Q_MX02 U8299 ( .S(n281), .A0(n2987), .A1(ofifoData[89]), .Z(n1223));
Q_FDP0UA U8300 ( .D(n1222), .QTFCLK( ), .Q(ofifoData[88]));
Q_MX02 U8301 ( .S(n281), .A0(n2990), .A1(ofifoData[88]), .Z(n1222));
Q_FDP0UA U8302 ( .D(n1221), .QTFCLK( ), .Q(ofifoData[87]));
Q_MX02 U8303 ( .S(n281), .A0(n2993), .A1(ofifoData[87]), .Z(n1221));
Q_FDP0UA U8304 ( .D(n1220), .QTFCLK( ), .Q(ofifoData[86]));
Q_MX02 U8305 ( .S(n281), .A0(n2996), .A1(ofifoData[86]), .Z(n1220));
Q_FDP0UA U8306 ( .D(n1219), .QTFCLK( ), .Q(ofifoData[85]));
Q_MX02 U8307 ( .S(n281), .A0(n2999), .A1(ofifoData[85]), .Z(n1219));
Q_FDP0UA U8308 ( .D(n1218), .QTFCLK( ), .Q(ofifoData[84]));
Q_MX02 U8309 ( .S(n281), .A0(n3002), .A1(ofifoData[84]), .Z(n1218));
Q_FDP0UA U8310 ( .D(n1217), .QTFCLK( ), .Q(ofifoData[83]));
Q_MX02 U8311 ( .S(n281), .A0(n3005), .A1(ofifoData[83]), .Z(n1217));
Q_FDP0UA U8312 ( .D(n1216), .QTFCLK( ), .Q(ofifoData[82]));
Q_MX02 U8313 ( .S(n281), .A0(n3008), .A1(ofifoData[82]), .Z(n1216));
Q_FDP0UA U8314 ( .D(n1215), .QTFCLK( ), .Q(ofifoData[81]));
Q_MX02 U8315 ( .S(n281), .A0(n3011), .A1(ofifoData[81]), .Z(n1215));
Q_FDP0UA U8316 ( .D(n1214), .QTFCLK( ), .Q(ofifoData[80]));
Q_MX02 U8317 ( .S(n281), .A0(n3014), .A1(ofifoData[80]), .Z(n1214));
Q_FDP0UA U8318 ( .D(n1213), .QTFCLK( ), .Q(ofifoData[79]));
Q_MX02 U8319 ( .S(n281), .A0(n3017), .A1(ofifoData[79]), .Z(n1213));
Q_FDP0UA U8320 ( .D(n1212), .QTFCLK( ), .Q(ofifoData[78]));
Q_MX02 U8321 ( .S(n281), .A0(n3020), .A1(ofifoData[78]), .Z(n1212));
Q_FDP0UA U8322 ( .D(n1211), .QTFCLK( ), .Q(ofifoData[77]));
Q_MX02 U8323 ( .S(n281), .A0(n3023), .A1(ofifoData[77]), .Z(n1211));
Q_FDP0UA U8324 ( .D(n1210), .QTFCLK( ), .Q(ofifoData[76]));
Q_MX02 U8325 ( .S(n281), .A0(n3026), .A1(ofifoData[76]), .Z(n1210));
Q_FDP0UA U8326 ( .D(n1209), .QTFCLK( ), .Q(ofifoData[75]));
Q_MX02 U8327 ( .S(n281), .A0(n3029), .A1(ofifoData[75]), .Z(n1209));
Q_FDP0UA U8328 ( .D(n1208), .QTFCLK( ), .Q(ofifoData[74]));
Q_MX02 U8329 ( .S(n281), .A0(n3032), .A1(ofifoData[74]), .Z(n1208));
Q_FDP0UA U8330 ( .D(n1207), .QTFCLK( ), .Q(ofifoData[73]));
Q_MX02 U8331 ( .S(n281), .A0(n3035), .A1(ofifoData[73]), .Z(n1207));
Q_FDP0UA U8332 ( .D(n1206), .QTFCLK( ), .Q(ofifoData[72]));
Q_MX02 U8333 ( .S(n281), .A0(n3038), .A1(ofifoData[72]), .Z(n1206));
Q_FDP0UA U8334 ( .D(n1205), .QTFCLK( ), .Q(ofifoData[71]));
Q_MX02 U8335 ( .S(n281), .A0(n3041), .A1(ofifoData[71]), .Z(n1205));
Q_FDP0UA U8336 ( .D(n1204), .QTFCLK( ), .Q(ofifoData[70]));
Q_MX02 U8337 ( .S(n281), .A0(n3044), .A1(ofifoData[70]), .Z(n1204));
Q_FDP0UA U8338 ( .D(n1203), .QTFCLK( ), .Q(ofifoData[69]));
Q_MX02 U8339 ( .S(n281), .A0(n3047), .A1(ofifoData[69]), .Z(n1203));
Q_FDP0UA U8340 ( .D(n1202), .QTFCLK( ), .Q(ofifoData[68]));
Q_MX02 U8341 ( .S(n281), .A0(n3050), .A1(ofifoData[68]), .Z(n1202));
Q_FDP0UA U8342 ( .D(n1201), .QTFCLK( ), .Q(ofifoData[67]));
Q_MX02 U8343 ( .S(n281), .A0(n3053), .A1(ofifoData[67]), .Z(n1201));
Q_FDP0UA U8344 ( .D(n1200), .QTFCLK( ), .Q(ofifoData[66]));
Q_MX02 U8345 ( .S(n281), .A0(n3056), .A1(ofifoData[66]), .Z(n1200));
Q_FDP0UA U8346 ( .D(n1199), .QTFCLK( ), .Q(ofifoData[65]));
Q_MX02 U8347 ( .S(n281), .A0(n3059), .A1(ofifoData[65]), .Z(n1199));
Q_FDP0UA U8348 ( .D(n1198), .QTFCLK( ), .Q(ofifoData[64]));
Q_MX02 U8349 ( .S(n281), .A0(n3062), .A1(ofifoData[64]), .Z(n1198));
Q_FDP0UA U8350 ( .D(n1197), .QTFCLK( ), .Q(ofifoData[63]));
Q_MX02 U8351 ( .S(n281), .A0(n3065), .A1(ofifoData[63]), .Z(n1197));
Q_FDP0UA U8352 ( .D(n1196), .QTFCLK( ), .Q(ofifoData[62]));
Q_MX02 U8353 ( .S(n281), .A0(n3068), .A1(ofifoData[62]), .Z(n1196));
Q_FDP0UA U8354 ( .D(n1195), .QTFCLK( ), .Q(ofifoData[61]));
Q_MX02 U8355 ( .S(n281), .A0(n3071), .A1(ofifoData[61]), .Z(n1195));
Q_FDP0UA U8356 ( .D(n1194), .QTFCLK( ), .Q(ofifoData[60]));
Q_MX02 U8357 ( .S(n281), .A0(n3074), .A1(ofifoData[60]), .Z(n1194));
Q_FDP0UA U8358 ( .D(n1193), .QTFCLK( ), .Q(ofifoData[59]));
Q_MX02 U8359 ( .S(n281), .A0(n3077), .A1(ofifoData[59]), .Z(n1193));
Q_FDP0UA U8360 ( .D(n1192), .QTFCLK( ), .Q(ofifoData[58]));
Q_MX02 U8361 ( .S(n281), .A0(n3080), .A1(ofifoData[58]), .Z(n1192));
Q_FDP0UA U8362 ( .D(n1191), .QTFCLK( ), .Q(ofifoData[57]));
Q_MX02 U8363 ( .S(n281), .A0(n3083), .A1(ofifoData[57]), .Z(n1191));
Q_FDP0UA U8364 ( .D(n1190), .QTFCLK( ), .Q(ofifoData[56]));
Q_MX02 U8365 ( .S(n281), .A0(n3086), .A1(ofifoData[56]), .Z(n1190));
Q_FDP0UA U8366 ( .D(n1189), .QTFCLK( ), .Q(ofifoData[55]));
Q_MX02 U8367 ( .S(n281), .A0(n3089), .A1(ofifoData[55]), .Z(n1189));
Q_FDP0UA U8368 ( .D(n1188), .QTFCLK( ), .Q(ofifoData[54]));
Q_MX02 U8369 ( .S(n281), .A0(n3092), .A1(ofifoData[54]), .Z(n1188));
Q_FDP0UA U8370 ( .D(n1187), .QTFCLK( ), .Q(ofifoData[53]));
Q_MX02 U8371 ( .S(n281), .A0(n3095), .A1(ofifoData[53]), .Z(n1187));
Q_FDP0UA U8372 ( .D(n1186), .QTFCLK( ), .Q(ofifoData[52]));
Q_MX02 U8373 ( .S(n281), .A0(n3098), .A1(ofifoData[52]), .Z(n1186));
Q_FDP0UA U8374 ( .D(n1185), .QTFCLK( ), .Q(ofifoData[51]));
Q_MX02 U8375 ( .S(n281), .A0(n3101), .A1(ofifoData[51]), .Z(n1185));
Q_FDP0UA U8376 ( .D(n1184), .QTFCLK( ), .Q(ofifoData[50]));
Q_MX02 U8377 ( .S(n281), .A0(n3104), .A1(ofifoData[50]), .Z(n1184));
Q_FDP0UA U8378 ( .D(n1183), .QTFCLK( ), .Q(ofifoData[49]));
Q_MX02 U8379 ( .S(n281), .A0(n3107), .A1(ofifoData[49]), .Z(n1183));
Q_FDP0UA U8380 ( .D(n1182), .QTFCLK( ), .Q(ofifoData[48]));
Q_MX02 U8381 ( .S(n281), .A0(n3110), .A1(ofifoData[48]), .Z(n1182));
Q_FDP0UA U8382 ( .D(n1181), .QTFCLK( ), .Q(ofifoData[47]));
Q_MX02 U8383 ( .S(n281), .A0(n3113), .A1(ofifoData[47]), .Z(n1181));
Q_FDP0UA U8384 ( .D(n1180), .QTFCLK( ), .Q(ofifoData[46]));
Q_MX02 U8385 ( .S(n281), .A0(n3116), .A1(ofifoData[46]), .Z(n1180));
Q_FDP0UA U8386 ( .D(n1179), .QTFCLK( ), .Q(ofifoData[45]));
Q_MX02 U8387 ( .S(n281), .A0(n3119), .A1(ofifoData[45]), .Z(n1179));
Q_FDP0UA U8388 ( .D(n1178), .QTFCLK( ), .Q(ofifoData[44]));
Q_MX02 U8389 ( .S(n281), .A0(n3122), .A1(ofifoData[44]), .Z(n1178));
Q_FDP0UA U8390 ( .D(n1177), .QTFCLK( ), .Q(ofifoData[43]));
Q_MX02 U8391 ( .S(n281), .A0(n3125), .A1(ofifoData[43]), .Z(n1177));
Q_FDP0UA U8392 ( .D(n1176), .QTFCLK( ), .Q(ofifoData[42]));
Q_MX02 U8393 ( .S(n281), .A0(n3128), .A1(ofifoData[42]), .Z(n1176));
Q_FDP0UA U8394 ( .D(n1175), .QTFCLK( ), .Q(ofifoData[41]));
Q_MX02 U8395 ( .S(n281), .A0(n3131), .A1(ofifoData[41]), .Z(n1175));
Q_FDP0UA U8396 ( .D(n1174), .QTFCLK( ), .Q(ofifoData[40]));
Q_MX02 U8397 ( .S(n281), .A0(n3134), .A1(ofifoData[40]), .Z(n1174));
Q_FDP0UA U8398 ( .D(n1173), .QTFCLK( ), .Q(ofifoData[39]));
Q_MX02 U8399 ( .S(n281), .A0(n3137), .A1(ofifoData[39]), .Z(n1173));
Q_FDP0UA U8400 ( .D(n1172), .QTFCLK( ), .Q(ofifoData[38]));
Q_MX02 U8401 ( .S(n281), .A0(n3140), .A1(ofifoData[38]), .Z(n1172));
Q_FDP0UA U8402 ( .D(n1171), .QTFCLK( ), .Q(ofifoData[37]));
Q_MX02 U8403 ( .S(n281), .A0(n3143), .A1(ofifoData[37]), .Z(n1171));
Q_FDP0UA U8404 ( .D(n1170), .QTFCLK( ), .Q(ofifoData[36]));
Q_MX02 U8405 ( .S(n281), .A0(n3146), .A1(ofifoData[36]), .Z(n1170));
Q_FDP0UA U8406 ( .D(n1169), .QTFCLK( ), .Q(ofifoData[35]));
Q_MX02 U8407 ( .S(n281), .A0(n3149), .A1(ofifoData[35]), .Z(n1169));
Q_FDP0UA U8408 ( .D(n1168), .QTFCLK( ), .Q(ofifoData[34]));
Q_MX02 U8409 ( .S(n281), .A0(n3152), .A1(ofifoData[34]), .Z(n1168));
Q_FDP0UA U8410 ( .D(n1167), .QTFCLK( ), .Q(ofifoData[33]));
Q_MX02 U8411 ( .S(n281), .A0(n3155), .A1(ofifoData[33]), .Z(n1167));
Q_FDP0UA U8412 ( .D(n1166), .QTFCLK( ), .Q(ofifoData[32]));
Q_MX02 U8413 ( .S(n281), .A0(n3158), .A1(ofifoData[32]), .Z(n1166));
Q_FDP0UA U8414 ( .D(n1165), .QTFCLK( ), .Q(ofifoData[31]));
Q_MX02 U8415 ( .S(n281), .A0(n3161), .A1(ofifoData[31]), .Z(n1165));
Q_FDP0UA U8416 ( .D(n1164), .QTFCLK( ), .Q(ofifoData[30]));
Q_MX02 U8417 ( .S(n281), .A0(n3164), .A1(ofifoData[30]), .Z(n1164));
Q_FDP0UA U8418 ( .D(n1163), .QTFCLK( ), .Q(ofifoData[29]));
Q_MX02 U8419 ( .S(n281), .A0(n3167), .A1(ofifoData[29]), .Z(n1163));
Q_FDP0UA U8420 ( .D(n1162), .QTFCLK( ), .Q(ofifoData[28]));
Q_MX02 U8421 ( .S(n281), .A0(n3170), .A1(ofifoData[28]), .Z(n1162));
Q_FDP0UA U8422 ( .D(n1161), .QTFCLK( ), .Q(ofifoData[27]));
Q_MX02 U8423 ( .S(n281), .A0(n3173), .A1(ofifoData[27]), .Z(n1161));
Q_FDP0UA U8424 ( .D(n1160), .QTFCLK( ), .Q(ofifoData[26]));
Q_MX02 U8425 ( .S(n281), .A0(n3176), .A1(ofifoData[26]), .Z(n1160));
Q_FDP0UA U8426 ( .D(n1159), .QTFCLK( ), .Q(ofifoData[25]));
Q_MX02 U8427 ( .S(n281), .A0(n3179), .A1(ofifoData[25]), .Z(n1159));
Q_FDP0UA U8428 ( .D(n1158), .QTFCLK( ), .Q(ofifoData[24]));
Q_MX02 U8429 ( .S(n281), .A0(n3182), .A1(ofifoData[24]), .Z(n1158));
Q_FDP0UA U8430 ( .D(n1157), .QTFCLK( ), .Q(ofifoData[23]));
Q_MX02 U8431 ( .S(n281), .A0(n3185), .A1(ofifoData[23]), .Z(n1157));
Q_FDP0UA U8432 ( .D(n1156), .QTFCLK( ), .Q(ofifoData[22]));
Q_MX02 U8433 ( .S(n281), .A0(n3188), .A1(ofifoData[22]), .Z(n1156));
Q_FDP0UA U8434 ( .D(n1155), .QTFCLK( ), .Q(ofifoData[21]));
Q_MX02 U8435 ( .S(n281), .A0(n3191), .A1(ofifoData[21]), .Z(n1155));
Q_FDP0UA U8436 ( .D(n1154), .QTFCLK( ), .Q(ofifoData[20]));
Q_MX02 U8437 ( .S(n281), .A0(n3194), .A1(ofifoData[20]), .Z(n1154));
Q_FDP0UA U8438 ( .D(n1153), .QTFCLK( ), .Q(ofifoData[19]));
Q_MX02 U8439 ( .S(n281), .A0(n3197), .A1(ofifoData[19]), .Z(n1153));
Q_FDP0UA U8440 ( .D(n1152), .QTFCLK( ), .Q(ofifoData[18]));
Q_MX02 U8441 ( .S(n281), .A0(n3200), .A1(ofifoData[18]), .Z(n1152));
Q_FDP0UA U8442 ( .D(n1151), .QTFCLK( ), .Q(ofifoData[17]));
Q_MX02 U8443 ( .S(n281), .A0(n3203), .A1(ofifoData[17]), .Z(n1151));
Q_FDP0UA U8444 ( .D(n1150), .QTFCLK( ), .Q(ofifoData[16]));
Q_MX02 U8445 ( .S(n281), .A0(n3206), .A1(ofifoData[16]), .Z(n1150));
Q_FDP0UA U8446 ( .D(n1149), .QTFCLK( ), .Q(ofifoData[15]));
Q_MX02 U8447 ( .S(n281), .A0(n3209), .A1(ofifoData[15]), .Z(n1149));
Q_FDP0UA U8448 ( .D(n1148), .QTFCLK( ), .Q(ofifoData[14]));
Q_MX02 U8449 ( .S(n281), .A0(n3212), .A1(ofifoData[14]), .Z(n1148));
Q_FDP0UA U8450 ( .D(n1147), .QTFCLK( ), .Q(ofifoData[13]));
Q_MX02 U8451 ( .S(n281), .A0(n3215), .A1(ofifoData[13]), .Z(n1147));
Q_FDP0UA U8452 ( .D(n1146), .QTFCLK( ), .Q(ofifoData[12]));
Q_MX02 U8453 ( .S(n281), .A0(n3218), .A1(ofifoData[12]), .Z(n1146));
Q_FDP0UA U8454 ( .D(n1145), .QTFCLK( ), .Q(ofifoData[11]));
Q_MX02 U8455 ( .S(n281), .A0(n3221), .A1(ofifoData[11]), .Z(n1145));
Q_FDP0UA U8456 ( .D(n1144), .QTFCLK( ), .Q(ofifoData[10]));
Q_MX02 U8457 ( .S(n281), .A0(n3224), .A1(ofifoData[10]), .Z(n1144));
Q_FDP0UA U8458 ( .D(n1143), .QTFCLK( ), .Q(ofifoData[9]));
Q_MX02 U8459 ( .S(n281), .A0(n3227), .A1(ofifoData[9]), .Z(n1143));
Q_FDP0UA U8460 ( .D(n1142), .QTFCLK( ), .Q(ofifoData[8]));
Q_MX02 U8461 ( .S(n281), .A0(n3230), .A1(ofifoData[8]), .Z(n1142));
Q_FDP0UA U8462 ( .D(n1141), .QTFCLK( ), .Q(ofifoData[7]));
Q_MX02 U8463 ( .S(n281), .A0(n3233), .A1(ofifoData[7]), .Z(n1141));
Q_FDP0UA U8464 ( .D(n1140), .QTFCLK( ), .Q(ofifoData[6]));
Q_MX02 U8465 ( .S(n281), .A0(n3236), .A1(ofifoData[6]), .Z(n1140));
Q_FDP0UA U8466 ( .D(n1139), .QTFCLK( ), .Q(ofifoData[5]));
Q_MX02 U8467 ( .S(n281), .A0(n3239), .A1(ofifoData[5]), .Z(n1139));
Q_FDP0UA U8468 ( .D(n1138), .QTFCLK( ), .Q(ofifoData[4]));
Q_MX02 U8469 ( .S(n281), .A0(n3242), .A1(ofifoData[4]), .Z(n1138));
Q_FDP0UA U8470 ( .D(n1137), .QTFCLK( ), .Q(ofifoData[3]));
Q_MX02 U8471 ( .S(n281), .A0(n3245), .A1(ofifoData[3]), .Z(n1137));
Q_FDP0UA U8472 ( .D(n1136), .QTFCLK( ), .Q(ofifoData[2]));
Q_MX02 U8473 ( .S(n281), .A0(n3248), .A1(ofifoData[2]), .Z(n1136));
Q_FDP0UA U8474 ( .D(n1135), .QTFCLK( ), .Q(ofifoData[1]));
Q_MX02 U8475 ( .S(n281), .A0(n3251), .A1(ofifoData[1]), .Z(n1135));
Q_FDP0UA U8476 ( .D(n1134), .QTFCLK( ), .Q(ofifoData[0]));
Q_MX02 U8477 ( .S(n281), .A0(n3254), .A1(ofifoData[0]), .Z(n1134));
Q_FDP0UA U8478 ( .D(n1133), .QTFCLK( ), .Q(ofifoAddr0[14]));
Q_MX02 U8479 ( .S(n275), .A0(n3257), .A1(ofifoAddr0[14]), .Z(n1133));
Q_FDP0UA U8480 ( .D(n1132), .QTFCLK( ), .Q(ofifoAddr0[13]));
Q_MX02 U8481 ( .S(n275), .A0(n3258), .A1(ofifoAddr0[13]), .Z(n1132));
Q_FDP0UA U8482 ( .D(n1131), .QTFCLK( ), .Q(ofifoAddr0[12]));
Q_MX02 U8483 ( .S(n275), .A0(n3259), .A1(ofifoAddr0[12]), .Z(n1131));
Q_FDP0UA U8484 ( .D(n1130), .QTFCLK( ), .Q(ofifoAddr0[11]));
Q_MX02 U8485 ( .S(n275), .A0(n3260), .A1(ofifoAddr0[11]), .Z(n1130));
Q_FDP0UA U8486 ( .D(n1129), .QTFCLK( ), .Q(ofifoAddr0[10]));
Q_MX02 U8487 ( .S(n275), .A0(n3261), .A1(ofifoAddr0[10]), .Z(n1129));
Q_FDP0UA U8488 ( .D(n1128), .QTFCLK( ), .Q(ofifoAddr0[9]));
Q_MX02 U8489 ( .S(n275), .A0(n3262), .A1(ofifoAddr0[9]), .Z(n1128));
Q_FDP0UA U8490 ( .D(n1127), .QTFCLK( ), .Q(ofifoAddr0[8]));
Q_MX02 U8491 ( .S(n275), .A0(n3263), .A1(ofifoAddr0[8]), .Z(n1127));
Q_FDP0UA U8492 ( .D(n1126), .QTFCLK( ), .Q(ofifoAddr0[7]));
Q_MX02 U8493 ( .S(n275), .A0(n3264), .A1(ofifoAddr0[7]), .Z(n1126));
Q_FDP0UA U8494 ( .D(n1125), .QTFCLK( ), .Q(ofifoAddr0[6]));
Q_MX02 U8495 ( .S(n275), .A0(n3265), .A1(ofifoAddr0[6]), .Z(n1125));
Q_FDP0UA U8496 ( .D(n1124), .QTFCLK( ), .Q(ofifoAddr0[5]));
Q_MX02 U8497 ( .S(n275), .A0(n3266), .A1(ofifoAddr0[5]), .Z(n1124));
Q_FDP0UA U8498 ( .D(n1123), .QTFCLK( ), .Q(ofifoAddr0[4]));
Q_MX02 U8499 ( .S(n275), .A0(n3267), .A1(ofifoAddr0[4]), .Z(n1123));
Q_FDP0UA U8500 ( .D(n1122), .QTFCLK( ), .Q(ofifoAddr0[3]));
Q_MX02 U8501 ( .S(n275), .A0(n3268), .A1(ofifoAddr0[3]), .Z(n1122));
Q_FDP0UA U8502 ( .D(n1121), .QTFCLK( ), .Q(ofifoAddr0[2]));
Q_MX02 U8503 ( .S(n275), .A0(n3269), .A1(ofifoAddr0[2]), .Z(n1121));
Q_FDP0UA U8504 ( .D(n1120), .QTFCLK( ), .Q(ofifoAddr0[1]));
Q_MX02 U8505 ( .S(n275), .A0(n3270), .A1(ofifoAddr0[1]), .Z(n1120));
Q_FDP0UA U8506 ( .D(n1119), .QTFCLK( ), .Q(ofifoAddr0[0]));
Q_MX02 U8507 ( .S(n275), .A0(n3271), .A1(ofifoAddr0[0]), .Z(n1119));
Q_FDP0UA U8508 ( .D(n1118), .QTFCLK( ), .Q(ofifoAddr1[15]));
Q_MX02 U8509 ( .S(n275), .A0(n3272), .A1(ofifoAddr1[15]), .Z(n1118));
Q_FDP0UA U8510 ( .D(n1117), .QTFCLK( ), .Q(ofifoAddr1[14]));
Q_MX02 U8511 ( .S(n275), .A0(n3273), .A1(ofifoAddr1[14]), .Z(n1117));
Q_FDP0UA U8512 ( .D(n1116), .QTFCLK( ), .Q(ofifoAddr1[13]));
Q_MX02 U8513 ( .S(n275), .A0(n3274), .A1(ofifoAddr1[13]), .Z(n1116));
Q_FDP0UA U8514 ( .D(n1115), .QTFCLK( ), .Q(ofifoAddr1[12]));
Q_MX02 U8515 ( .S(n275), .A0(n3275), .A1(ofifoAddr1[12]), .Z(n1115));
Q_FDP0UA U8516 ( .D(n1114), .QTFCLK( ), .Q(ofifoAddr1[11]));
Q_MX02 U8517 ( .S(n275), .A0(n3276), .A1(ofifoAddr1[11]), .Z(n1114));
Q_FDP0UA U8518 ( .D(n1113), .QTFCLK( ), .Q(ofifoAddr1[10]));
Q_MX02 U8519 ( .S(n275), .A0(n3277), .A1(ofifoAddr1[10]), .Z(n1113));
Q_FDP0UA U8520 ( .D(n1112), .QTFCLK( ), .Q(ofifoAddr1[9]));
Q_MX02 U8521 ( .S(n275), .A0(n3278), .A1(ofifoAddr1[9]), .Z(n1112));
Q_FDP0UA U8522 ( .D(n1111), .QTFCLK( ), .Q(ofifoAddr1[8]));
Q_MX02 U8523 ( .S(n275), .A0(n3279), .A1(ofifoAddr1[8]), .Z(n1111));
Q_FDP0UA U8524 ( .D(n1110), .QTFCLK( ), .Q(ofifoAddr1[7]));
Q_MX02 U8525 ( .S(n275), .A0(n3280), .A1(ofifoAddr1[7]), .Z(n1110));
Q_FDP0UA U8526 ( .D(n1109), .QTFCLK( ), .Q(ofifoAddr1[6]));
Q_MX02 U8527 ( .S(n275), .A0(n3281), .A1(ofifoAddr1[6]), .Z(n1109));
Q_FDP0UA U8528 ( .D(n1108), .QTFCLK( ), .Q(ofifoAddr1[5]));
Q_MX02 U8529 ( .S(n275), .A0(n3282), .A1(ofifoAddr1[5]), .Z(n1108));
Q_FDP0UA U8530 ( .D(n1107), .QTFCLK( ), .Q(ofifoAddr1[4]));
Q_MX02 U8531 ( .S(n275), .A0(n3283), .A1(ofifoAddr1[4]), .Z(n1107));
Q_FDP0UA U8532 ( .D(n1106), .QTFCLK( ), .Q(ofifoAddr1[3]));
Q_MX02 U8533 ( .S(n275), .A0(n3284), .A1(ofifoAddr1[3]), .Z(n1106));
Q_FDP0UA U8534 ( .D(n1105), .QTFCLK( ), .Q(ofifoAddr1[2]));
Q_MX02 U8535 ( .S(n275), .A0(n3285), .A1(ofifoAddr1[2]), .Z(n1105));
Q_FDP0UA U8536 ( .D(n1104), .QTFCLK( ), .Q(ofifoAddr1[1]));
Q_MX02 U8537 ( .S(n275), .A0(n3286), .A1(ofifoAddr1[1]), .Z(n1104));
Q_FDP0UA U8538 ( .D(n1103), .QTFCLK( ), .Q(ofifoAddr1[0]));
Q_MX02 U8539 ( .S(n275), .A0(n6887), .A1(ofifoAddr1[0]), .Z(n1103));
Q_FDP0UA U8540 ( .D(n1102), .QTFCLK( ), .Q(ofifoAddr2[15]));
Q_MX02 U8541 ( .S(n275), .A0(n3287), .A1(ofifoAddr2[15]), .Z(n1102));
Q_FDP0UA U8542 ( .D(n1101), .QTFCLK( ), .Q(ofifoAddr2[14]));
Q_MX02 U8543 ( .S(n275), .A0(n3288), .A1(ofifoAddr2[14]), .Z(n1101));
Q_FDP0UA U8544 ( .D(n1100), .QTFCLK( ), .Q(ofifoAddr2[13]));
Q_MX02 U8545 ( .S(n275), .A0(n3289), .A1(ofifoAddr2[13]), .Z(n1100));
Q_FDP0UA U8546 ( .D(n1099), .QTFCLK( ), .Q(ofifoAddr2[12]));
Q_MX02 U8547 ( .S(n275), .A0(n3290), .A1(ofifoAddr2[12]), .Z(n1099));
Q_FDP0UA U8548 ( .D(n1098), .QTFCLK( ), .Q(ofifoAddr2[11]));
Q_MX02 U8549 ( .S(n275), .A0(n3291), .A1(ofifoAddr2[11]), .Z(n1098));
Q_FDP0UA U8550 ( .D(n1097), .QTFCLK( ), .Q(ofifoAddr2[10]));
Q_MX02 U8551 ( .S(n275), .A0(n3292), .A1(ofifoAddr2[10]), .Z(n1097));
Q_FDP0UA U8552 ( .D(n1096), .QTFCLK( ), .Q(ofifoAddr2[9]));
Q_MX02 U8553 ( .S(n275), .A0(n3293), .A1(ofifoAddr2[9]), .Z(n1096));
Q_FDP0UA U8554 ( .D(n1095), .QTFCLK( ), .Q(ofifoAddr2[8]));
Q_MX02 U8555 ( .S(n275), .A0(n3294), .A1(ofifoAddr2[8]), .Z(n1095));
Q_FDP0UA U8556 ( .D(n1094), .QTFCLK( ), .Q(ofifoAddr2[7]));
Q_MX02 U8557 ( .S(n275), .A0(n3295), .A1(ofifoAddr2[7]), .Z(n1094));
Q_FDP0UA U8558 ( .D(n1093), .QTFCLK( ), .Q(ofifoAddr2[6]));
Q_MX02 U8559 ( .S(n275), .A0(n3296), .A1(ofifoAddr2[6]), .Z(n1093));
Q_FDP0UA U8560 ( .D(n1092), .QTFCLK( ), .Q(ofifoAddr2[5]));
Q_MX02 U8561 ( .S(n275), .A0(n3297), .A1(ofifoAddr2[5]), .Z(n1092));
Q_FDP0UA U8562 ( .D(n1091), .QTFCLK( ), .Q(ofifoAddr2[4]));
Q_MX02 U8563 ( .S(n275), .A0(n3298), .A1(ofifoAddr2[4]), .Z(n1091));
Q_FDP0UA U8564 ( .D(n1090), .QTFCLK( ), .Q(ofifoAddr2[3]));
Q_MX02 U8565 ( .S(n275), .A0(n3299), .A1(ofifoAddr2[3]), .Z(n1090));
Q_FDP0UA U8566 ( .D(n1089), .QTFCLK( ), .Q(ofifoAddr2[2]));
Q_MX02 U8567 ( .S(n275), .A0(n3300), .A1(ofifoAddr2[2]), .Z(n1089));
Q_FDP0UA U8568 ( .D(n1088), .QTFCLK( ), .Q(ofifoAddr2[1]));
Q_MX02 U8569 ( .S(n275), .A0(n3301), .A1(ofifoAddr2[1]), .Z(n1088));
Q_FDP0UA U8570 ( .D(n1087), .QTFCLK( ), .Q(ofifoAddr2[0]));
Q_MX02 U8571 ( .S(n275), .A0(n3271), .A1(ofifoAddr2[0]), .Z(n1087));
Q_FDP0UA U8572 ( .D(n1086), .QTFCLK( ), .Q(ofifoWptr[14]));
Q_MX02 U8573 ( .S(n281), .A0(n3302), .A1(ofifoWptr[14]), .Z(n1086));
Q_FDP0UA U8574 ( .D(n1085), .QTFCLK( ), .Q(ofifoWptr[13]));
Q_MX02 U8575 ( .S(n281), .A0(n3303), .A1(ofifoWptr[13]), .Z(n1085));
Q_FDP0UA U8576 ( .D(n1084), .QTFCLK( ), .Q(ofifoWptr[12]));
Q_MX02 U8577 ( .S(n281), .A0(n3304), .A1(ofifoWptr[12]), .Z(n1084));
Q_FDP0UA U8578 ( .D(n1083), .QTFCLK( ), .Q(ofifoWptr[11]));
Q_MX02 U8579 ( .S(n281), .A0(n3305), .A1(ofifoWptr[11]), .Z(n1083));
Q_FDP0UA U8580 ( .D(n1082), .QTFCLK( ), .Q(ofifoWptr[10]));
Q_MX02 U8581 ( .S(n281), .A0(n3306), .A1(ofifoWptr[10]), .Z(n1082));
Q_FDP0UA U8582 ( .D(n1081), .QTFCLK( ), .Q(ofifoWptr[9]));
Q_MX02 U8583 ( .S(n281), .A0(n3307), .A1(ofifoWptr[9]), .Z(n1081));
Q_FDP0UA U8584 ( .D(n1080), .QTFCLK( ), .Q(ofifoWptr[8]));
Q_MX02 U8585 ( .S(n281), .A0(n3308), .A1(ofifoWptr[8]), .Z(n1080));
Q_FDP0UA U8586 ( .D(n1079), .QTFCLK( ), .Q(ofifoWptr[7]));
Q_MX02 U8587 ( .S(n281), .A0(n3309), .A1(ofifoWptr[7]), .Z(n1079));
Q_FDP0UA U8588 ( .D(n1078), .QTFCLK( ), .Q(ofifoWptr[6]));
Q_MX02 U8589 ( .S(n281), .A0(n3310), .A1(ofifoWptr[6]), .Z(n1078));
Q_FDP0UA U8590 ( .D(n1077), .QTFCLK( ), .Q(ofifoWptr[5]));
Q_MX02 U8591 ( .S(n281), .A0(n3311), .A1(ofifoWptr[5]), .Z(n1077));
Q_FDP0UA U8592 ( .D(n1076), .QTFCLK( ), .Q(ofifoWptr[4]));
Q_MX02 U8593 ( .S(n281), .A0(n3312), .A1(ofifoWptr[4]), .Z(n1076));
Q_FDP0UA U8594 ( .D(n1075), .QTFCLK( ), .Q(ofifoWptr[3]));
Q_MX02 U8595 ( .S(n281), .A0(n3313), .A1(ofifoWptr[3]), .Z(n1075));
Q_FDP0UA U8596 ( .D(n1074), .QTFCLK( ), .Q(ofifoWptr[2]));
Q_MX02 U8597 ( .S(n281), .A0(n3314), .A1(ofifoWptr[2]), .Z(n1074));
Q_FDP0UA U8598 ( .D(n1073), .QTFCLK( ), .Q(ofifoWptr[1]));
Q_MX02 U8599 ( .S(n281), .A0(n3315), .A1(ofifoWptr[1]), .Z(n1073));
Q_FDP0UA U8600 ( .D(n1072), .QTFCLK( ), .Q(ofifoWptr[0]));
Q_MX02 U8601 ( .S(n281), .A0(n3316), .A1(ofifoWptr[0]), .Z(n1072));
Q_FDP0UA U8602 ( .D(n1071), .QTFCLK( ), .Q(shiftedOData[767]));
Q_AN02 U8603 ( .A0(n301), .A1(shiftedOData[767]), .Z(n1071));
Q_FDP0UA U8604 ( .D(n1070), .QTFCLK( ), .Q(shiftedOData[766]));
Q_AN02 U8605 ( .A0(n301), .A1(shiftedOData[766]), .Z(n1070));
Q_FDP0UA U8606 ( .D(n1069), .QTFCLK( ), .Q(shiftedOData[765]));
Q_AN02 U8607 ( .A0(n301), .A1(shiftedOData[765]), .Z(n1069));
Q_FDP0UA U8608 ( .D(n1068), .QTFCLK( ), .Q(shiftedOData[764]));
Q_AN02 U8609 ( .A0(n301), .A1(shiftedOData[764]), .Z(n1068));
Q_FDP0UA U8610 ( .D(n1067), .QTFCLK( ), .Q(shiftedOData[763]));
Q_AN02 U8611 ( .A0(n301), .A1(shiftedOData[763]), .Z(n1067));
Q_FDP0UA U8612 ( .D(n1066), .QTFCLK( ), .Q(shiftedOData[762]));
Q_AN02 U8613 ( .A0(n301), .A1(shiftedOData[762]), .Z(n1066));
Q_FDP0UA U8614 ( .D(n1065), .QTFCLK( ), .Q(shiftedOData[761]));
Q_AN02 U8615 ( .A0(n301), .A1(shiftedOData[761]), .Z(n1065));
Q_FDP0UA U8616 ( .D(n1064), .QTFCLK( ), .Q(shiftedOData[760]));
Q_AN02 U8617 ( .A0(n301), .A1(shiftedOData[760]), .Z(n1064));
Q_FDP0UA U8618 ( .D(n1063), .QTFCLK( ), .Q(shiftedOData[759]));
Q_AN02 U8619 ( .A0(n301), .A1(shiftedOData[759]), .Z(n1063));
Q_FDP0UA U8620 ( .D(n1062), .QTFCLK( ), .Q(shiftedOData[758]));
Q_AN02 U8621 ( .A0(n301), .A1(shiftedOData[758]), .Z(n1062));
Q_FDP0UA U8622 ( .D(n1061), .QTFCLK( ), .Q(shiftedOData[757]));
Q_AN02 U8623 ( .A0(n301), .A1(shiftedOData[757]), .Z(n1061));
Q_FDP0UA U8624 ( .D(n1060), .QTFCLK( ), .Q(shiftedOData[756]));
Q_AN02 U8625 ( .A0(n301), .A1(shiftedOData[756]), .Z(n1060));
Q_FDP0UA U8626 ( .D(n1059), .QTFCLK( ), .Q(shiftedOData[755]));
Q_AN02 U8627 ( .A0(n301), .A1(shiftedOData[755]), .Z(n1059));
Q_FDP0UA U8628 ( .D(n1058), .QTFCLK( ), .Q(shiftedOData[754]));
Q_AN02 U8629 ( .A0(n301), .A1(shiftedOData[754]), .Z(n1058));
Q_FDP0UA U8630 ( .D(n1057), .QTFCLK( ), .Q(shiftedOData[753]));
Q_AN02 U8631 ( .A0(n301), .A1(shiftedOData[753]), .Z(n1057));
Q_FDP0UA U8632 ( .D(n1056), .QTFCLK( ), .Q(shiftedOData[752]));
Q_AN02 U8633 ( .A0(n301), .A1(shiftedOData[752]), .Z(n1056));
Q_FDP0UA U8634 ( .D(n1055), .QTFCLK( ), .Q(shiftedOData[751]));
Q_AN02 U8635 ( .A0(n301), .A1(shiftedOData[751]), .Z(n1055));
Q_FDP0UA U8636 ( .D(n1054), .QTFCLK( ), .Q(shiftedOData[750]));
Q_AN02 U8637 ( .A0(n301), .A1(shiftedOData[750]), .Z(n1054));
Q_FDP0UA U8638 ( .D(n1053), .QTFCLK( ), .Q(shiftedOData[749]));
Q_AN02 U8639 ( .A0(n301), .A1(shiftedOData[749]), .Z(n1053));
Q_FDP0UA U8640 ( .D(n1052), .QTFCLK( ), .Q(shiftedOData[748]));
Q_AN02 U8641 ( .A0(n301), .A1(shiftedOData[748]), .Z(n1052));
Q_FDP0UA U8642 ( .D(n1051), .QTFCLK( ), .Q(shiftedOData[747]));
Q_AN02 U8643 ( .A0(n301), .A1(shiftedOData[747]), .Z(n1051));
Q_FDP0UA U8644 ( .D(n1050), .QTFCLK( ), .Q(shiftedOData[746]));
Q_AN02 U8645 ( .A0(n301), .A1(shiftedOData[746]), .Z(n1050));
Q_FDP0UA U8646 ( .D(n1049), .QTFCLK( ), .Q(shiftedOData[745]));
Q_AN02 U8647 ( .A0(n301), .A1(shiftedOData[745]), .Z(n1049));
Q_FDP0UA U8648 ( .D(n1048), .QTFCLK( ), .Q(shiftedOData[744]));
Q_AN02 U8649 ( .A0(n301), .A1(shiftedOData[744]), .Z(n1048));
Q_FDP0UA U8650 ( .D(n1047), .QTFCLK( ), .Q(shiftedOData[743]));
Q_AN02 U8651 ( .A0(n301), .A1(shiftedOData[743]), .Z(n1047));
Q_FDP0UA U8652 ( .D(n1046), .QTFCLK( ), .Q(shiftedOData[742]));
Q_AN02 U8653 ( .A0(n301), .A1(shiftedOData[742]), .Z(n1046));
Q_FDP0UA U8654 ( .D(n1045), .QTFCLK( ), .Q(shiftedOData[741]));
Q_AN02 U8655 ( .A0(n301), .A1(shiftedOData[741]), .Z(n1045));
Q_FDP0UA U8656 ( .D(n1044), .QTFCLK( ), .Q(shiftedOData[740]));
Q_AN02 U8657 ( .A0(n301), .A1(shiftedOData[740]), .Z(n1044));
Q_FDP0UA U8658 ( .D(n1043), .QTFCLK( ), .Q(shiftedOData[739]));
Q_AN02 U8659 ( .A0(n301), .A1(shiftedOData[739]), .Z(n1043));
Q_FDP0UA U8660 ( .D(n1042), .QTFCLK( ), .Q(shiftedOData[738]));
Q_AN02 U8661 ( .A0(n301), .A1(shiftedOData[738]), .Z(n1042));
Q_FDP0UA U8662 ( .D(n1041), .QTFCLK( ), .Q(shiftedOData[737]));
Q_AN02 U8663 ( .A0(n301), .A1(shiftedOData[737]), .Z(n1041));
Q_FDP0UA U8664 ( .D(n1040), .QTFCLK( ), .Q(shiftedOData[736]));
Q_AN02 U8665 ( .A0(n301), .A1(shiftedOData[736]), .Z(n1040));
Q_FDP0UA U8666 ( .D(n1039), .QTFCLK( ), .Q(shiftedOData[735]));
Q_AN02 U8667 ( .A0(n301), .A1(shiftedOData[735]), .Z(n1039));
Q_FDP0UA U8668 ( .D(n1038), .QTFCLK( ), .Q(shiftedOData[734]));
Q_AN02 U8669 ( .A0(n301), .A1(shiftedOData[734]), .Z(n1038));
Q_FDP0UA U8670 ( .D(n1037), .QTFCLK( ), .Q(shiftedOData[733]));
Q_AN02 U8671 ( .A0(n301), .A1(shiftedOData[733]), .Z(n1037));
Q_FDP0UA U8672 ( .D(n1036), .QTFCLK( ), .Q(shiftedOData[732]));
Q_AN02 U8673 ( .A0(n301), .A1(shiftedOData[732]), .Z(n1036));
Q_FDP0UA U8674 ( .D(n1035), .QTFCLK( ), .Q(shiftedOData[731]));
Q_AN02 U8675 ( .A0(n301), .A1(shiftedOData[731]), .Z(n1035));
Q_FDP0UA U8676 ( .D(n1034), .QTFCLK( ), .Q(shiftedOData[730]));
Q_AN02 U8677 ( .A0(n301), .A1(shiftedOData[730]), .Z(n1034));
Q_FDP0UA U8678 ( .D(n1033), .QTFCLK( ), .Q(shiftedOData[729]));
Q_AN02 U8679 ( .A0(n301), .A1(shiftedOData[729]), .Z(n1033));
Q_FDP0UA U8680 ( .D(n1032), .QTFCLK( ), .Q(shiftedOData[728]));
Q_AN02 U8681 ( .A0(n301), .A1(shiftedOData[728]), .Z(n1032));
Q_FDP0UA U8682 ( .D(n1031), .QTFCLK( ), .Q(shiftedOData[727]));
Q_AN02 U8683 ( .A0(n301), .A1(shiftedOData[727]), .Z(n1031));
Q_FDP0UA U8684 ( .D(n1030), .QTFCLK( ), .Q(shiftedOData[726]));
Q_AN02 U8685 ( .A0(n301), .A1(shiftedOData[726]), .Z(n1030));
Q_FDP0UA U8686 ( .D(n1029), .QTFCLK( ), .Q(shiftedOData[725]));
Q_AN02 U8687 ( .A0(n301), .A1(shiftedOData[725]), .Z(n1029));
Q_FDP0UA U8688 ( .D(n1028), .QTFCLK( ), .Q(shiftedOData[724]));
Q_AN02 U8689 ( .A0(n301), .A1(shiftedOData[724]), .Z(n1028));
Q_FDP0UA U8690 ( .D(n1027), .QTFCLK( ), .Q(shiftedOData[723]));
Q_AN02 U8691 ( .A0(n301), .A1(shiftedOData[723]), .Z(n1027));
Q_FDP0UA U8692 ( .D(n1026), .QTFCLK( ), .Q(shiftedOData[722]));
Q_AN02 U8693 ( .A0(n301), .A1(shiftedOData[722]), .Z(n1026));
Q_FDP0UA U8694 ( .D(n1025), .QTFCLK( ), .Q(shiftedOData[721]));
Q_AN02 U8695 ( .A0(n301), .A1(shiftedOData[721]), .Z(n1025));
Q_FDP0UA U8696 ( .D(n1024), .QTFCLK( ), .Q(shiftedOData[720]));
Q_AN02 U8697 ( .A0(n301), .A1(shiftedOData[720]), .Z(n1024));
Q_FDP0UA U8698 ( .D(n1023), .QTFCLK( ), .Q(shiftedOData[719]));
Q_AN02 U8699 ( .A0(n301), .A1(shiftedOData[719]), .Z(n1023));
Q_FDP0UA U8700 ( .D(n1022), .QTFCLK( ), .Q(shiftedOData[718]));
Q_AN02 U8701 ( .A0(n301), .A1(shiftedOData[718]), .Z(n1022));
Q_FDP0UA U8702 ( .D(n1021), .QTFCLK( ), .Q(shiftedOData[717]));
Q_AN02 U8703 ( .A0(n301), .A1(shiftedOData[717]), .Z(n1021));
Q_FDP0UA U8704 ( .D(n1020), .QTFCLK( ), .Q(shiftedOData[716]));
Q_AN02 U8705 ( .A0(n301), .A1(shiftedOData[716]), .Z(n1020));
Q_FDP0UA U8706 ( .D(n1019), .QTFCLK( ), .Q(shiftedOData[715]));
Q_AN02 U8707 ( .A0(n301), .A1(shiftedOData[715]), .Z(n1019));
Q_FDP0UA U8708 ( .D(n1018), .QTFCLK( ), .Q(shiftedOData[714]));
Q_AN02 U8709 ( .A0(n301), .A1(shiftedOData[714]), .Z(n1018));
Q_FDP0UA U8710 ( .D(n1017), .QTFCLK( ), .Q(shiftedOData[713]));
Q_AN02 U8711 ( .A0(n301), .A1(shiftedOData[713]), .Z(n1017));
Q_FDP0UA U8712 ( .D(n1016), .QTFCLK( ), .Q(shiftedOData[712]));
Q_AN02 U8713 ( .A0(n301), .A1(shiftedOData[712]), .Z(n1016));
Q_FDP0UA U8714 ( .D(n1015), .QTFCLK( ), .Q(shiftedOData[711]));
Q_AN02 U8715 ( .A0(n301), .A1(shiftedOData[711]), .Z(n1015));
Q_FDP0UA U8716 ( .D(n1014), .QTFCLK( ), .Q(shiftedOData[710]));
Q_AN02 U8717 ( .A0(n301), .A1(shiftedOData[710]), .Z(n1014));
Q_FDP0UA U8718 ( .D(n1013), .QTFCLK( ), .Q(shiftedOData[709]));
Q_AN02 U8719 ( .A0(n301), .A1(shiftedOData[709]), .Z(n1013));
Q_FDP0UA U8720 ( .D(n1012), .QTFCLK( ), .Q(shiftedOData[708]));
Q_AN02 U8721 ( .A0(n301), .A1(shiftedOData[708]), .Z(n1012));
Q_FDP0UA U8722 ( .D(n1011), .QTFCLK( ), .Q(shiftedOData[707]));
Q_AN02 U8723 ( .A0(n301), .A1(shiftedOData[707]), .Z(n1011));
Q_FDP0UA U8724 ( .D(n1010), .QTFCLK( ), .Q(shiftedOData[706]));
Q_AN02 U8725 ( .A0(n301), .A1(shiftedOData[706]), .Z(n1010));
Q_FDP0UA U8726 ( .D(n1009), .QTFCLK( ), .Q(shiftedOData[705]));
Q_AN02 U8727 ( .A0(n301), .A1(shiftedOData[705]), .Z(n1009));
Q_FDP0UA U8728 ( .D(n1008), .QTFCLK( ), .Q(shiftedOData[704]));
Q_AN02 U8729 ( .A0(n301), .A1(shiftedOData[704]), .Z(n1008));
Q_FDP0UA U8730 ( .D(n1007), .QTFCLK( ), .Q(shiftedOData[703]));
Q_MX02 U8731 ( .S(n280), .A0(shiftedOData[703]), .A1(n4434), .Z(n1007));
Q_FDP0UA U8732 ( .D(n1006), .QTFCLK( ), .Q(shiftedOData[702]));
Q_MX02 U8733 ( .S(n280), .A0(shiftedOData[702]), .A1(n4433), .Z(n1006));
Q_FDP0UA U8734 ( .D(n1005), .QTFCLK( ), .Q(shiftedOData[701]));
Q_MX02 U8735 ( .S(n280), .A0(shiftedOData[701]), .A1(n4432), .Z(n1005));
Q_FDP0UA U8736 ( .D(n1004), .QTFCLK( ), .Q(shiftedOData[700]));
Q_MX02 U8737 ( .S(n280), .A0(shiftedOData[700]), .A1(n4431), .Z(n1004));
Q_FDP0UA U8738 ( .D(n1003), .QTFCLK( ), .Q(shiftedOData[699]));
Q_MX02 U8739 ( .S(n280), .A0(shiftedOData[699]), .A1(n4430), .Z(n1003));
Q_FDP0UA U8740 ( .D(n1002), .QTFCLK( ), .Q(shiftedOData[698]));
Q_MX02 U8741 ( .S(n280), .A0(shiftedOData[698]), .A1(n4429), .Z(n1002));
Q_FDP0UA U8742 ( .D(n1001), .QTFCLK( ), .Q(shiftedOData[697]));
Q_MX02 U8743 ( .S(n280), .A0(shiftedOData[697]), .A1(n4428), .Z(n1001));
Q_FDP0UA U8744 ( .D(n1000), .QTFCLK( ), .Q(shiftedOData[696]));
Q_MX02 U8745 ( .S(n280), .A0(shiftedOData[696]), .A1(n4427), .Z(n1000));
Q_FDP0UA U8746 ( .D(n999), .QTFCLK( ), .Q(shiftedOData[695]));
Q_MX02 U8747 ( .S(n280), .A0(shiftedOData[695]), .A1(n4426), .Z(n999));
Q_FDP0UA U8748 ( .D(n998), .QTFCLK( ), .Q(shiftedOData[694]));
Q_MX02 U8749 ( .S(n280), .A0(shiftedOData[694]), .A1(n4425), .Z(n998));
Q_FDP0UA U8750 ( .D(n997), .QTFCLK( ), .Q(shiftedOData[693]));
Q_MX02 U8751 ( .S(n280), .A0(shiftedOData[693]), .A1(n4424), .Z(n997));
Q_FDP0UA U8752 ( .D(n996), .QTFCLK( ), .Q(shiftedOData[692]));
Q_MX02 U8753 ( .S(n280), .A0(shiftedOData[692]), .A1(n4423), .Z(n996));
Q_FDP0UA U8754 ( .D(n995), .QTFCLK( ), .Q(shiftedOData[691]));
Q_MX02 U8755 ( .S(n280), .A0(shiftedOData[691]), .A1(n4422), .Z(n995));
Q_FDP0UA U8756 ( .D(n994), .QTFCLK( ), .Q(shiftedOData[690]));
Q_MX02 U8757 ( .S(n280), .A0(shiftedOData[690]), .A1(n4421), .Z(n994));
Q_FDP0UA U8758 ( .D(n993), .QTFCLK( ), .Q(shiftedOData[689]));
Q_MX02 U8759 ( .S(n280), .A0(shiftedOData[689]), .A1(n4420), .Z(n993));
Q_FDP0UA U8760 ( .D(n992), .QTFCLK( ), .Q(shiftedOData[688]));
Q_MX02 U8761 ( .S(n280), .A0(shiftedOData[688]), .A1(n4419), .Z(n992));
Q_FDP0UA U8762 ( .D(n991), .QTFCLK( ), .Q(shiftedOData[687]));
Q_MX02 U8763 ( .S(n280), .A0(shiftedOData[687]), .A1(n4418), .Z(n991));
Q_FDP0UA U8764 ( .D(n990), .QTFCLK( ), .Q(shiftedOData[686]));
Q_MX02 U8765 ( .S(n280), .A0(shiftedOData[686]), .A1(n4417), .Z(n990));
Q_FDP0UA U8766 ( .D(n989), .QTFCLK( ), .Q(shiftedOData[685]));
Q_MX02 U8767 ( .S(n280), .A0(shiftedOData[685]), .A1(n4416), .Z(n989));
Q_FDP0UA U8768 ( .D(n988), .QTFCLK( ), .Q(shiftedOData[684]));
Q_MX02 U8769 ( .S(n280), .A0(shiftedOData[684]), .A1(n4415), .Z(n988));
Q_FDP0UA U8770 ( .D(n987), .QTFCLK( ), .Q(shiftedOData[683]));
Q_MX02 U8771 ( .S(n280), .A0(shiftedOData[683]), .A1(n4414), .Z(n987));
Q_FDP0UA U8772 ( .D(n986), .QTFCLK( ), .Q(shiftedOData[682]));
Q_MX02 U8773 ( .S(n280), .A0(shiftedOData[682]), .A1(n4413), .Z(n986));
Q_FDP0UA U8774 ( .D(n985), .QTFCLK( ), .Q(shiftedOData[681]));
Q_MX02 U8775 ( .S(n280), .A0(shiftedOData[681]), .A1(n4412), .Z(n985));
Q_FDP0UA U8776 ( .D(n984), .QTFCLK( ), .Q(shiftedOData[680]));
Q_MX02 U8777 ( .S(n280), .A0(shiftedOData[680]), .A1(n4411), .Z(n984));
Q_FDP0UA U8778 ( .D(n983), .QTFCLK( ), .Q(shiftedOData[679]));
Q_MX02 U8779 ( .S(n280), .A0(shiftedOData[679]), .A1(n4410), .Z(n983));
Q_FDP0UA U8780 ( .D(n982), .QTFCLK( ), .Q(shiftedOData[678]));
Q_MX02 U8781 ( .S(n280), .A0(shiftedOData[678]), .A1(n4409), .Z(n982));
Q_FDP0UA U8782 ( .D(n981), .QTFCLK( ), .Q(shiftedOData[677]));
Q_MX02 U8783 ( .S(n280), .A0(shiftedOData[677]), .A1(n4408), .Z(n981));
Q_FDP0UA U8784 ( .D(n980), .QTFCLK( ), .Q(shiftedOData[676]));
Q_MX02 U8785 ( .S(n280), .A0(shiftedOData[676]), .A1(n4407), .Z(n980));
Q_FDP0UA U8786 ( .D(n979), .QTFCLK( ), .Q(shiftedOData[675]));
Q_MX02 U8787 ( .S(n280), .A0(shiftedOData[675]), .A1(n4406), .Z(n979));
Q_FDP0UA U8788 ( .D(n978), .QTFCLK( ), .Q(shiftedOData[674]));
Q_MX02 U8789 ( .S(n280), .A0(shiftedOData[674]), .A1(n4405), .Z(n978));
Q_FDP0UA U8790 ( .D(n977), .QTFCLK( ), .Q(shiftedOData[673]));
Q_MX02 U8791 ( .S(n280), .A0(shiftedOData[673]), .A1(n4404), .Z(n977));
Q_FDP0UA U8792 ( .D(n976), .QTFCLK( ), .Q(shiftedOData[672]));
Q_MX02 U8793 ( .S(n280), .A0(shiftedOData[672]), .A1(n4403), .Z(n976));
Q_FDP0UA U8794 ( .D(n975), .QTFCLK( ), .Q(shiftedOData[671]));
Q_MX02 U8795 ( .S(n280), .A0(shiftedOData[671]), .A1(n4402), .Z(n975));
Q_FDP0UA U8796 ( .D(n974), .QTFCLK( ), .Q(shiftedOData[670]));
Q_MX02 U8797 ( .S(n280), .A0(shiftedOData[670]), .A1(n4401), .Z(n974));
Q_FDP0UA U8798 ( .D(n973), .QTFCLK( ), .Q(shiftedOData[669]));
Q_MX02 U8799 ( .S(n280), .A0(shiftedOData[669]), .A1(n4400), .Z(n973));
Q_FDP0UA U8800 ( .D(n972), .QTFCLK( ), .Q(shiftedOData[668]));
Q_MX02 U8801 ( .S(n280), .A0(shiftedOData[668]), .A1(n4399), .Z(n972));
Q_FDP0UA U8802 ( .D(n971), .QTFCLK( ), .Q(shiftedOData[667]));
Q_MX02 U8803 ( .S(n280), .A0(shiftedOData[667]), .A1(n4398), .Z(n971));
Q_FDP0UA U8804 ( .D(n970), .QTFCLK( ), .Q(shiftedOData[666]));
Q_MX02 U8805 ( .S(n280), .A0(shiftedOData[666]), .A1(n4397), .Z(n970));
Q_FDP0UA U8806 ( .D(n969), .QTFCLK( ), .Q(shiftedOData[665]));
Q_MX02 U8807 ( .S(n280), .A0(shiftedOData[665]), .A1(n4396), .Z(n969));
Q_FDP0UA U8808 ( .D(n968), .QTFCLK( ), .Q(shiftedOData[664]));
Q_MX02 U8809 ( .S(n280), .A0(shiftedOData[664]), .A1(n4395), .Z(n968));
Q_FDP0UA U8810 ( .D(n967), .QTFCLK( ), .Q(shiftedOData[663]));
Q_MX02 U8811 ( .S(n280), .A0(shiftedOData[663]), .A1(n4394), .Z(n967));
Q_FDP0UA U8812 ( .D(n966), .QTFCLK( ), .Q(shiftedOData[662]));
Q_MX02 U8813 ( .S(n280), .A0(shiftedOData[662]), .A1(n4393), .Z(n966));
Q_FDP0UA U8814 ( .D(n965), .QTFCLK( ), .Q(shiftedOData[661]));
Q_MX02 U8815 ( .S(n280), .A0(shiftedOData[661]), .A1(n4392), .Z(n965));
Q_FDP0UA U8816 ( .D(n964), .QTFCLK( ), .Q(shiftedOData[660]));
Q_MX02 U8817 ( .S(n280), .A0(shiftedOData[660]), .A1(n4391), .Z(n964));
Q_FDP0UA U8818 ( .D(n963), .QTFCLK( ), .Q(shiftedOData[659]));
Q_MX02 U8819 ( .S(n280), .A0(shiftedOData[659]), .A1(n4390), .Z(n963));
Q_FDP0UA U8820 ( .D(n962), .QTFCLK( ), .Q(shiftedOData[658]));
Q_MX02 U8821 ( .S(n280), .A0(shiftedOData[658]), .A1(n4389), .Z(n962));
Q_FDP0UA U8822 ( .D(n961), .QTFCLK( ), .Q(shiftedOData[657]));
Q_MX02 U8823 ( .S(n280), .A0(shiftedOData[657]), .A1(n4388), .Z(n961));
Q_FDP0UA U8824 ( .D(n960), .QTFCLK( ), .Q(shiftedOData[656]));
Q_MX02 U8825 ( .S(n280), .A0(shiftedOData[656]), .A1(n4387), .Z(n960));
Q_FDP0UA U8826 ( .D(n959), .QTFCLK( ), .Q(shiftedOData[655]));
Q_MX02 U8827 ( .S(n280), .A0(shiftedOData[655]), .A1(n4386), .Z(n959));
Q_FDP0UA U8828 ( .D(n958), .QTFCLK( ), .Q(shiftedOData[654]));
Q_MX02 U8829 ( .S(n280), .A0(shiftedOData[654]), .A1(n4385), .Z(n958));
Q_FDP0UA U8830 ( .D(n957), .QTFCLK( ), .Q(shiftedOData[653]));
Q_MX02 U8831 ( .S(n280), .A0(shiftedOData[653]), .A1(n4384), .Z(n957));
Q_FDP0UA U8832 ( .D(n956), .QTFCLK( ), .Q(shiftedOData[652]));
Q_MX02 U8833 ( .S(n280), .A0(shiftedOData[652]), .A1(n4383), .Z(n956));
Q_FDP0UA U8834 ( .D(n955), .QTFCLK( ), .Q(shiftedOData[651]));
Q_MX02 U8835 ( .S(n280), .A0(shiftedOData[651]), .A1(n4382), .Z(n955));
Q_FDP0UA U8836 ( .D(n954), .QTFCLK( ), .Q(shiftedOData[650]));
Q_MX02 U8837 ( .S(n280), .A0(shiftedOData[650]), .A1(n4381), .Z(n954));
Q_FDP0UA U8838 ( .D(n953), .QTFCLK( ), .Q(shiftedOData[649]));
Q_MX02 U8839 ( .S(n280), .A0(shiftedOData[649]), .A1(n4380), .Z(n953));
Q_FDP0UA U8840 ( .D(n952), .QTFCLK( ), .Q(shiftedOData[648]));
Q_MX02 U8841 ( .S(n280), .A0(shiftedOData[648]), .A1(n4379), .Z(n952));
Q_FDP0UA U8842 ( .D(n951), .QTFCLK( ), .Q(shiftedOData[647]));
Q_MX02 U8843 ( .S(n280), .A0(shiftedOData[647]), .A1(n4378), .Z(n951));
Q_FDP0UA U8844 ( .D(n950), .QTFCLK( ), .Q(shiftedOData[646]));
Q_MX02 U8845 ( .S(n280), .A0(shiftedOData[646]), .A1(n4377), .Z(n950));
Q_FDP0UA U8846 ( .D(n949), .QTFCLK( ), .Q(shiftedOData[645]));
Q_MX02 U8847 ( .S(n280), .A0(shiftedOData[645]), .A1(n4376), .Z(n949));
Q_FDP0UA U8848 ( .D(n948), .QTFCLK( ), .Q(shiftedOData[644]));
Q_MX02 U8849 ( .S(n280), .A0(shiftedOData[644]), .A1(n4375), .Z(n948));
Q_FDP0UA U8850 ( .D(n947), .QTFCLK( ), .Q(shiftedOData[643]));
Q_MX02 U8851 ( .S(n280), .A0(shiftedOData[643]), .A1(n4374), .Z(n947));
Q_FDP0UA U8852 ( .D(n946), .QTFCLK( ), .Q(shiftedOData[642]));
Q_MX02 U8853 ( .S(n280), .A0(shiftedOData[642]), .A1(n4373), .Z(n946));
Q_FDP0UA U8854 ( .D(n945), .QTFCLK( ), .Q(shiftedOData[641]));
Q_MX02 U8855 ( .S(n280), .A0(shiftedOData[641]), .A1(n4372), .Z(n945));
Q_FDP0UA U8856 ( .D(n944), .QTFCLK( ), .Q(shiftedOData[640]));
Q_MX02 U8857 ( .S(n280), .A0(shiftedOData[640]), .A1(n4371), .Z(n944));
Q_FDP0UA U8858 ( .D(n943), .QTFCLK( ), .Q(shiftedOData[639]));
Q_MX02 U8859 ( .S(n280), .A0(shiftedOData[639]), .A1(n4370), .Z(n943));
Q_FDP0UA U8860 ( .D(n942), .QTFCLK( ), .Q(shiftedOData[638]));
Q_MX02 U8861 ( .S(n280), .A0(shiftedOData[638]), .A1(n4369), .Z(n942));
Q_FDP0UA U8862 ( .D(n941), .QTFCLK( ), .Q(shiftedOData[637]));
Q_MX02 U8863 ( .S(n280), .A0(shiftedOData[637]), .A1(n4368), .Z(n941));
Q_FDP0UA U8864 ( .D(n940), .QTFCLK( ), .Q(shiftedOData[636]));
Q_MX02 U8865 ( .S(n280), .A0(shiftedOData[636]), .A1(n4367), .Z(n940));
Q_FDP0UA U8866 ( .D(n939), .QTFCLK( ), .Q(shiftedOData[635]));
Q_MX02 U8867 ( .S(n280), .A0(shiftedOData[635]), .A1(n4366), .Z(n939));
Q_FDP0UA U8868 ( .D(n938), .QTFCLK( ), .Q(shiftedOData[634]));
Q_MX02 U8869 ( .S(n280), .A0(shiftedOData[634]), .A1(n4365), .Z(n938));
Q_FDP0UA U8870 ( .D(n937), .QTFCLK( ), .Q(shiftedOData[633]));
Q_MX02 U8871 ( .S(n280), .A0(shiftedOData[633]), .A1(n4364), .Z(n937));
Q_FDP0UA U8872 ( .D(n936), .QTFCLK( ), .Q(shiftedOData[632]));
Q_MX02 U8873 ( .S(n280), .A0(shiftedOData[632]), .A1(n4363), .Z(n936));
Q_FDP0UA U8874 ( .D(n935), .QTFCLK( ), .Q(shiftedOData[631]));
Q_MX02 U8875 ( .S(n280), .A0(shiftedOData[631]), .A1(n4362), .Z(n935));
Q_FDP0UA U8876 ( .D(n934), .QTFCLK( ), .Q(shiftedOData[630]));
Q_MX02 U8877 ( .S(n280), .A0(shiftedOData[630]), .A1(n4361), .Z(n934));
Q_FDP0UA U8878 ( .D(n933), .QTFCLK( ), .Q(shiftedOData[629]));
Q_MX02 U8879 ( .S(n280), .A0(shiftedOData[629]), .A1(n4360), .Z(n933));
Q_FDP0UA U8880 ( .D(n932), .QTFCLK( ), .Q(shiftedOData[628]));
Q_MX02 U8881 ( .S(n280), .A0(shiftedOData[628]), .A1(n4359), .Z(n932));
Q_FDP0UA U8882 ( .D(n931), .QTFCLK( ), .Q(shiftedOData[627]));
Q_MX02 U8883 ( .S(n280), .A0(shiftedOData[627]), .A1(n4358), .Z(n931));
Q_FDP0UA U8884 ( .D(n930), .QTFCLK( ), .Q(shiftedOData[626]));
Q_MX02 U8885 ( .S(n280), .A0(shiftedOData[626]), .A1(n4357), .Z(n930));
Q_FDP0UA U8886 ( .D(n929), .QTFCLK( ), .Q(shiftedOData[625]));
Q_MX02 U8887 ( .S(n280), .A0(shiftedOData[625]), .A1(n4356), .Z(n929));
Q_FDP0UA U8888 ( .D(n928), .QTFCLK( ), .Q(shiftedOData[624]));
Q_MX02 U8889 ( .S(n280), .A0(shiftedOData[624]), .A1(n4355), .Z(n928));
Q_FDP0UA U8890 ( .D(n927), .QTFCLK( ), .Q(shiftedOData[623]));
Q_MX02 U8891 ( .S(n280), .A0(shiftedOData[623]), .A1(n4354), .Z(n927));
Q_FDP0UA U8892 ( .D(n926), .QTFCLK( ), .Q(shiftedOData[622]));
Q_MX02 U8893 ( .S(n280), .A0(shiftedOData[622]), .A1(n4353), .Z(n926));
Q_FDP0UA U8894 ( .D(n925), .QTFCLK( ), .Q(shiftedOData[621]));
Q_MX02 U8895 ( .S(n280), .A0(shiftedOData[621]), .A1(n4352), .Z(n925));
Q_FDP0UA U8896 ( .D(n924), .QTFCLK( ), .Q(shiftedOData[620]));
Q_MX02 U8897 ( .S(n280), .A0(shiftedOData[620]), .A1(n4351), .Z(n924));
Q_FDP0UA U8898 ( .D(n923), .QTFCLK( ), .Q(shiftedOData[619]));
Q_MX02 U8899 ( .S(n280), .A0(shiftedOData[619]), .A1(n4350), .Z(n923));
Q_FDP0UA U8900 ( .D(n922), .QTFCLK( ), .Q(shiftedOData[618]));
Q_MX02 U8901 ( .S(n280), .A0(shiftedOData[618]), .A1(n4349), .Z(n922));
Q_FDP0UA U8902 ( .D(n921), .QTFCLK( ), .Q(shiftedOData[617]));
Q_MX02 U8903 ( .S(n280), .A0(shiftedOData[617]), .A1(n4348), .Z(n921));
Q_FDP0UA U8904 ( .D(n920), .QTFCLK( ), .Q(shiftedOData[616]));
Q_MX02 U8905 ( .S(n280), .A0(shiftedOData[616]), .A1(n4347), .Z(n920));
Q_FDP0UA U8906 ( .D(n919), .QTFCLK( ), .Q(shiftedOData[615]));
Q_MX02 U8907 ( .S(n280), .A0(shiftedOData[615]), .A1(n4346), .Z(n919));
Q_FDP0UA U8908 ( .D(n918), .QTFCLK( ), .Q(shiftedOData[614]));
Q_MX02 U8909 ( .S(n280), .A0(shiftedOData[614]), .A1(n4345), .Z(n918));
Q_FDP0UA U8910 ( .D(n917), .QTFCLK( ), .Q(shiftedOData[613]));
Q_MX02 U8911 ( .S(n280), .A0(shiftedOData[613]), .A1(n4344), .Z(n917));
Q_FDP0UA U8912 ( .D(n916), .QTFCLK( ), .Q(shiftedOData[612]));
Q_MX02 U8913 ( .S(n280), .A0(shiftedOData[612]), .A1(n4343), .Z(n916));
Q_FDP0UA U8914 ( .D(n915), .QTFCLK( ), .Q(shiftedOData[611]));
Q_MX02 U8915 ( .S(n280), .A0(shiftedOData[611]), .A1(n4342), .Z(n915));
Q_FDP0UA U8916 ( .D(n914), .QTFCLK( ), .Q(shiftedOData[610]));
Q_MX02 U8917 ( .S(n280), .A0(shiftedOData[610]), .A1(n4341), .Z(n914));
Q_FDP0UA U8918 ( .D(n913), .QTFCLK( ), .Q(shiftedOData[609]));
Q_MX02 U8919 ( .S(n280), .A0(shiftedOData[609]), .A1(n4340), .Z(n913));
Q_FDP0UA U8920 ( .D(n912), .QTFCLK( ), .Q(shiftedOData[608]));
Q_MX02 U8921 ( .S(n280), .A0(shiftedOData[608]), .A1(n4339), .Z(n912));
Q_FDP0UA U8922 ( .D(n911), .QTFCLK( ), .Q(shiftedOData[607]));
Q_MX02 U8923 ( .S(n280), .A0(shiftedOData[607]), .A1(n4338), .Z(n911));
Q_FDP0UA U8924 ( .D(n910), .QTFCLK( ), .Q(shiftedOData[606]));
Q_MX02 U8925 ( .S(n280), .A0(shiftedOData[606]), .A1(n4337), .Z(n910));
Q_FDP0UA U8926 ( .D(n909), .QTFCLK( ), .Q(shiftedOData[605]));
Q_MX02 U8927 ( .S(n280), .A0(shiftedOData[605]), .A1(n4336), .Z(n909));
Q_FDP0UA U8928 ( .D(n908), .QTFCLK( ), .Q(shiftedOData[604]));
Q_MX02 U8929 ( .S(n280), .A0(shiftedOData[604]), .A1(n4335), .Z(n908));
Q_FDP0UA U8930 ( .D(n907), .QTFCLK( ), .Q(shiftedOData[603]));
Q_MX02 U8931 ( .S(n280), .A0(shiftedOData[603]), .A1(n4334), .Z(n907));
Q_FDP0UA U8932 ( .D(n906), .QTFCLK( ), .Q(shiftedOData[602]));
Q_MX02 U8933 ( .S(n280), .A0(shiftedOData[602]), .A1(n4333), .Z(n906));
Q_FDP0UA U8934 ( .D(n905), .QTFCLK( ), .Q(shiftedOData[601]));
Q_MX02 U8935 ( .S(n280), .A0(shiftedOData[601]), .A1(n4332), .Z(n905));
Q_FDP0UA U8936 ( .D(n904), .QTFCLK( ), .Q(shiftedOData[600]));
Q_MX02 U8937 ( .S(n280), .A0(shiftedOData[600]), .A1(n4331), .Z(n904));
Q_FDP0UA U8938 ( .D(n903), .QTFCLK( ), .Q(shiftedOData[599]));
Q_MX02 U8939 ( .S(n280), .A0(shiftedOData[599]), .A1(n4330), .Z(n903));
Q_FDP0UA U8940 ( .D(n902), .QTFCLK( ), .Q(shiftedOData[598]));
Q_MX02 U8941 ( .S(n280), .A0(shiftedOData[598]), .A1(n4329), .Z(n902));
Q_FDP0UA U8942 ( .D(n901), .QTFCLK( ), .Q(shiftedOData[597]));
Q_MX02 U8943 ( .S(n280), .A0(shiftedOData[597]), .A1(n4328), .Z(n901));
Q_FDP0UA U8944 ( .D(n900), .QTFCLK( ), .Q(shiftedOData[596]));
Q_MX02 U8945 ( .S(n280), .A0(shiftedOData[596]), .A1(n4327), .Z(n900));
Q_FDP0UA U8946 ( .D(n899), .QTFCLK( ), .Q(shiftedOData[595]));
Q_MX02 U8947 ( .S(n280), .A0(shiftedOData[595]), .A1(n4326), .Z(n899));
Q_FDP0UA U8948 ( .D(n898), .QTFCLK( ), .Q(shiftedOData[594]));
Q_MX02 U8949 ( .S(n280), .A0(shiftedOData[594]), .A1(n4325), .Z(n898));
Q_FDP0UA U8950 ( .D(n897), .QTFCLK( ), .Q(shiftedOData[593]));
Q_MX02 U8951 ( .S(n280), .A0(shiftedOData[593]), .A1(n4324), .Z(n897));
Q_FDP0UA U8952 ( .D(n896), .QTFCLK( ), .Q(shiftedOData[592]));
Q_MX02 U8953 ( .S(n280), .A0(shiftedOData[592]), .A1(n4323), .Z(n896));
Q_FDP0UA U8954 ( .D(n895), .QTFCLK( ), .Q(shiftedOData[591]));
Q_MX02 U8955 ( .S(n280), .A0(shiftedOData[591]), .A1(n4322), .Z(n895));
Q_FDP0UA U8956 ( .D(n894), .QTFCLK( ), .Q(shiftedOData[590]));
Q_MX02 U8957 ( .S(n280), .A0(shiftedOData[590]), .A1(n4321), .Z(n894));
Q_FDP0UA U8958 ( .D(n893), .QTFCLK( ), .Q(shiftedOData[589]));
Q_MX02 U8959 ( .S(n280), .A0(shiftedOData[589]), .A1(n4320), .Z(n893));
Q_FDP0UA U8960 ( .D(n892), .QTFCLK( ), .Q(shiftedOData[588]));
Q_MX02 U8961 ( .S(n280), .A0(shiftedOData[588]), .A1(n4319), .Z(n892));
Q_FDP0UA U8962 ( .D(n891), .QTFCLK( ), .Q(shiftedOData[587]));
Q_MX02 U8963 ( .S(n280), .A0(shiftedOData[587]), .A1(n4318), .Z(n891));
Q_FDP0UA U8964 ( .D(n890), .QTFCLK( ), .Q(shiftedOData[586]));
Q_MX02 U8965 ( .S(n280), .A0(shiftedOData[586]), .A1(n4317), .Z(n890));
Q_FDP0UA U8966 ( .D(n889), .QTFCLK( ), .Q(shiftedOData[585]));
Q_MX02 U8967 ( .S(n280), .A0(shiftedOData[585]), .A1(n4316), .Z(n889));
Q_FDP0UA U8968 ( .D(n888), .QTFCLK( ), .Q(shiftedOData[584]));
Q_MX02 U8969 ( .S(n280), .A0(shiftedOData[584]), .A1(n4315), .Z(n888));
Q_FDP0UA U8970 ( .D(n887), .QTFCLK( ), .Q(shiftedOData[583]));
Q_MX02 U8971 ( .S(n280), .A0(shiftedOData[583]), .A1(n4314), .Z(n887));
Q_FDP0UA U8972 ( .D(n886), .QTFCLK( ), .Q(shiftedOData[582]));
Q_MX02 U8973 ( .S(n280), .A0(shiftedOData[582]), .A1(n4313), .Z(n886));
Q_FDP0UA U8974 ( .D(n885), .QTFCLK( ), .Q(shiftedOData[581]));
Q_MX02 U8975 ( .S(n280), .A0(shiftedOData[581]), .A1(n4312), .Z(n885));
Q_FDP0UA U8976 ( .D(n884), .QTFCLK( ), .Q(shiftedOData[580]));
Q_MX02 U8977 ( .S(n280), .A0(shiftedOData[580]), .A1(n4311), .Z(n884));
Q_FDP0UA U8978 ( .D(n883), .QTFCLK( ), .Q(shiftedOData[579]));
Q_MX02 U8979 ( .S(n280), .A0(shiftedOData[579]), .A1(n4310), .Z(n883));
Q_FDP0UA U8980 ( .D(n882), .QTFCLK( ), .Q(shiftedOData[578]));
Q_MX02 U8981 ( .S(n280), .A0(shiftedOData[578]), .A1(n4309), .Z(n882));
Q_FDP0UA U8982 ( .D(n881), .QTFCLK( ), .Q(shiftedOData[577]));
Q_MX02 U8983 ( .S(n280), .A0(shiftedOData[577]), .A1(n4308), .Z(n881));
Q_FDP0UA U8984 ( .D(n880), .QTFCLK( ), .Q(shiftedOData[576]));
Q_MX02 U8985 ( .S(n280), .A0(shiftedOData[576]), .A1(n4307), .Z(n880));
Q_FDP0UA U8986 ( .D(n879), .QTFCLK( ), .Q(shiftedOData[575]));
Q_MX02 U8987 ( .S(n280), .A0(shiftedOData[575]), .A1(n4306), .Z(n879));
Q_FDP0UA U8988 ( .D(n878), .QTFCLK( ), .Q(shiftedOData[574]));
Q_MX02 U8989 ( .S(n280), .A0(shiftedOData[574]), .A1(n4305), .Z(n878));
Q_FDP0UA U8990 ( .D(n877), .QTFCLK( ), .Q(shiftedOData[573]));
Q_MX02 U8991 ( .S(n280), .A0(shiftedOData[573]), .A1(n4304), .Z(n877));
Q_FDP0UA U8992 ( .D(n876), .QTFCLK( ), .Q(shiftedOData[572]));
Q_MX02 U8993 ( .S(n280), .A0(shiftedOData[572]), .A1(n4303), .Z(n876));
Q_FDP0UA U8994 ( .D(n875), .QTFCLK( ), .Q(shiftedOData[571]));
Q_MX02 U8995 ( .S(n280), .A0(shiftedOData[571]), .A1(n4302), .Z(n875));
Q_FDP0UA U8996 ( .D(n874), .QTFCLK( ), .Q(shiftedOData[570]));
Q_MX02 U8997 ( .S(n280), .A0(shiftedOData[570]), .A1(n4301), .Z(n874));
Q_FDP0UA U8998 ( .D(n873), .QTFCLK( ), .Q(shiftedOData[569]));
Q_MX02 U8999 ( .S(n280), .A0(shiftedOData[569]), .A1(n4300), .Z(n873));
Q_FDP0UA U9000 ( .D(n872), .QTFCLK( ), .Q(shiftedOData[568]));
Q_MX02 U9001 ( .S(n280), .A0(shiftedOData[568]), .A1(n4299), .Z(n872));
Q_FDP0UA U9002 ( .D(n871), .QTFCLK( ), .Q(shiftedOData[567]));
Q_MX02 U9003 ( .S(n280), .A0(shiftedOData[567]), .A1(n4298), .Z(n871));
Q_FDP0UA U9004 ( .D(n870), .QTFCLK( ), .Q(shiftedOData[566]));
Q_MX02 U9005 ( .S(n280), .A0(shiftedOData[566]), .A1(n4297), .Z(n870));
Q_FDP0UA U9006 ( .D(n869), .QTFCLK( ), .Q(shiftedOData[565]));
Q_MX02 U9007 ( .S(n280), .A0(shiftedOData[565]), .A1(n4296), .Z(n869));
Q_FDP0UA U9008 ( .D(n868), .QTFCLK( ), .Q(shiftedOData[564]));
Q_MX02 U9009 ( .S(n280), .A0(shiftedOData[564]), .A1(n4295), .Z(n868));
Q_FDP0UA U9010 ( .D(n867), .QTFCLK( ), .Q(shiftedOData[563]));
Q_MX02 U9011 ( .S(n280), .A0(shiftedOData[563]), .A1(n4294), .Z(n867));
Q_FDP0UA U9012 ( .D(n866), .QTFCLK( ), .Q(shiftedOData[562]));
Q_MX02 U9013 ( .S(n280), .A0(shiftedOData[562]), .A1(n4293), .Z(n866));
Q_FDP0UA U9014 ( .D(n865), .QTFCLK( ), .Q(shiftedOData[561]));
Q_MX02 U9015 ( .S(n280), .A0(shiftedOData[561]), .A1(n4292), .Z(n865));
Q_FDP0UA U9016 ( .D(n864), .QTFCLK( ), .Q(shiftedOData[560]));
Q_MX02 U9017 ( .S(n280), .A0(shiftedOData[560]), .A1(n4291), .Z(n864));
Q_FDP0UA U9018 ( .D(n863), .QTFCLK( ), .Q(shiftedOData[559]));
Q_MX02 U9019 ( .S(n280), .A0(shiftedOData[559]), .A1(n4290), .Z(n863));
Q_FDP0UA U9020 ( .D(n862), .QTFCLK( ), .Q(shiftedOData[558]));
Q_MX02 U9021 ( .S(n280), .A0(shiftedOData[558]), .A1(n4289), .Z(n862));
Q_FDP0UA U9022 ( .D(n861), .QTFCLK( ), .Q(shiftedOData[557]));
Q_MX02 U9023 ( .S(n280), .A0(shiftedOData[557]), .A1(n4288), .Z(n861));
Q_FDP0UA U9024 ( .D(n860), .QTFCLK( ), .Q(shiftedOData[556]));
Q_MX02 U9025 ( .S(n280), .A0(shiftedOData[556]), .A1(n4287), .Z(n860));
Q_FDP0UA U9026 ( .D(n859), .QTFCLK( ), .Q(shiftedOData[555]));
Q_MX02 U9027 ( .S(n280), .A0(shiftedOData[555]), .A1(n4286), .Z(n859));
Q_FDP0UA U9028 ( .D(n858), .QTFCLK( ), .Q(shiftedOData[554]));
Q_MX02 U9029 ( .S(n280), .A0(shiftedOData[554]), .A1(n4285), .Z(n858));
Q_FDP0UA U9030 ( .D(n857), .QTFCLK( ), .Q(shiftedOData[553]));
Q_MX02 U9031 ( .S(n280), .A0(shiftedOData[553]), .A1(n4284), .Z(n857));
Q_FDP0UA U9032 ( .D(n856), .QTFCLK( ), .Q(shiftedOData[552]));
Q_MX02 U9033 ( .S(n280), .A0(shiftedOData[552]), .A1(n4283), .Z(n856));
Q_FDP0UA U9034 ( .D(n855), .QTFCLK( ), .Q(shiftedOData[551]));
Q_MX02 U9035 ( .S(n280), .A0(shiftedOData[551]), .A1(n4282), .Z(n855));
Q_FDP0UA U9036 ( .D(n854), .QTFCLK( ), .Q(shiftedOData[550]));
Q_MX02 U9037 ( .S(n280), .A0(shiftedOData[550]), .A1(n4281), .Z(n854));
Q_FDP0UA U9038 ( .D(n853), .QTFCLK( ), .Q(shiftedOData[549]));
Q_MX02 U9039 ( .S(n280), .A0(shiftedOData[549]), .A1(n4280), .Z(n853));
Q_FDP0UA U9040 ( .D(n852), .QTFCLK( ), .Q(shiftedOData[548]));
Q_MX02 U9041 ( .S(n280), .A0(shiftedOData[548]), .A1(n4279), .Z(n852));
Q_FDP0UA U9042 ( .D(n851), .QTFCLK( ), .Q(shiftedOData[547]));
Q_MX02 U9043 ( .S(n280), .A0(shiftedOData[547]), .A1(n4278), .Z(n851));
Q_FDP0UA U9044 ( .D(n850), .QTFCLK( ), .Q(shiftedOData[546]));
Q_MX02 U9045 ( .S(n280), .A0(shiftedOData[546]), .A1(n4277), .Z(n850));
Q_FDP0UA U9046 ( .D(n849), .QTFCLK( ), .Q(shiftedOData[545]));
Q_MX02 U9047 ( .S(n280), .A0(shiftedOData[545]), .A1(n4276), .Z(n849));
Q_FDP0UA U9048 ( .D(n848), .QTFCLK( ), .Q(shiftedOData[544]));
Q_MX02 U9049 ( .S(n280), .A0(shiftedOData[544]), .A1(n4275), .Z(n848));
Q_FDP0UA U9050 ( .D(n847), .QTFCLK( ), .Q(shiftedOData[543]));
Q_MX02 U9051 ( .S(n280), .A0(shiftedOData[543]), .A1(n4274), .Z(n847));
Q_FDP0UA U9052 ( .D(n846), .QTFCLK( ), .Q(shiftedOData[542]));
Q_MX02 U9053 ( .S(n280), .A0(shiftedOData[542]), .A1(n4273), .Z(n846));
Q_FDP0UA U9054 ( .D(n845), .QTFCLK( ), .Q(shiftedOData[541]));
Q_MX02 U9055 ( .S(n280), .A0(shiftedOData[541]), .A1(n4272), .Z(n845));
Q_FDP0UA U9056 ( .D(n844), .QTFCLK( ), .Q(shiftedOData[540]));
Q_MX02 U9057 ( .S(n280), .A0(shiftedOData[540]), .A1(n4271), .Z(n844));
Q_FDP0UA U9058 ( .D(n843), .QTFCLK( ), .Q(shiftedOData[539]));
Q_MX02 U9059 ( .S(n280), .A0(shiftedOData[539]), .A1(n4270), .Z(n843));
Q_FDP0UA U9060 ( .D(n842), .QTFCLK( ), .Q(shiftedOData[538]));
Q_MX02 U9061 ( .S(n280), .A0(shiftedOData[538]), .A1(n4269), .Z(n842));
Q_FDP0UA U9062 ( .D(n841), .QTFCLK( ), .Q(shiftedOData[537]));
Q_MX02 U9063 ( .S(n280), .A0(shiftedOData[537]), .A1(n4268), .Z(n841));
Q_FDP0UA U9064 ( .D(n840), .QTFCLK( ), .Q(shiftedOData[536]));
Q_MX02 U9065 ( .S(n280), .A0(shiftedOData[536]), .A1(n4267), .Z(n840));
Q_FDP0UA U9066 ( .D(n839), .QTFCLK( ), .Q(shiftedOData[535]));
Q_MX02 U9067 ( .S(n280), .A0(shiftedOData[535]), .A1(n4266), .Z(n839));
Q_FDP0UA U9068 ( .D(n838), .QTFCLK( ), .Q(shiftedOData[534]));
Q_MX02 U9069 ( .S(n280), .A0(shiftedOData[534]), .A1(n4265), .Z(n838));
Q_FDP0UA U9070 ( .D(n837), .QTFCLK( ), .Q(shiftedOData[533]));
Q_MX02 U9071 ( .S(n280), .A0(shiftedOData[533]), .A1(n4264), .Z(n837));
Q_FDP0UA U9072 ( .D(n836), .QTFCLK( ), .Q(shiftedOData[532]));
Q_MX02 U9073 ( .S(n280), .A0(shiftedOData[532]), .A1(n4263), .Z(n836));
Q_FDP0UA U9074 ( .D(n835), .QTFCLK( ), .Q(shiftedOData[531]));
Q_MX02 U9075 ( .S(n280), .A0(shiftedOData[531]), .A1(n4262), .Z(n835));
Q_FDP0UA U9076 ( .D(n834), .QTFCLK( ), .Q(shiftedOData[530]));
Q_MX02 U9077 ( .S(n280), .A0(shiftedOData[530]), .A1(n4261), .Z(n834));
Q_FDP0UA U9078 ( .D(n833), .QTFCLK( ), .Q(shiftedOData[529]));
Q_MX02 U9079 ( .S(n280), .A0(shiftedOData[529]), .A1(n4260), .Z(n833));
Q_FDP0UA U9080 ( .D(n832), .QTFCLK( ), .Q(shiftedOData[528]));
Q_MX02 U9081 ( .S(n280), .A0(shiftedOData[528]), .A1(n4259), .Z(n832));
Q_FDP0UA U9082 ( .D(n831), .QTFCLK( ), .Q(shiftedOData[527]));
Q_MX02 U9083 ( .S(n280), .A0(shiftedOData[527]), .A1(n4258), .Z(n831));
Q_FDP0UA U9084 ( .D(n830), .QTFCLK( ), .Q(shiftedOData[526]));
Q_MX02 U9085 ( .S(n280), .A0(shiftedOData[526]), .A1(n4257), .Z(n830));
Q_FDP0UA U9086 ( .D(n829), .QTFCLK( ), .Q(shiftedOData[525]));
Q_MX02 U9087 ( .S(n280), .A0(shiftedOData[525]), .A1(n4256), .Z(n829));
Q_FDP0UA U9088 ( .D(n828), .QTFCLK( ), .Q(shiftedOData[524]));
Q_MX02 U9089 ( .S(n280), .A0(shiftedOData[524]), .A1(n4255), .Z(n828));
Q_FDP0UA U9090 ( .D(n827), .QTFCLK( ), .Q(shiftedOData[523]));
Q_MX02 U9091 ( .S(n280), .A0(shiftedOData[523]), .A1(n4254), .Z(n827));
Q_FDP0UA U9092 ( .D(n826), .QTFCLK( ), .Q(shiftedOData[522]));
Q_MX02 U9093 ( .S(n280), .A0(shiftedOData[522]), .A1(n4253), .Z(n826));
Q_FDP0UA U9094 ( .D(n825), .QTFCLK( ), .Q(shiftedOData[521]));
Q_MX02 U9095 ( .S(n280), .A0(shiftedOData[521]), .A1(n4252), .Z(n825));
Q_FDP0UA U9096 ( .D(n824), .QTFCLK( ), .Q(shiftedOData[520]));
Q_MX02 U9097 ( .S(n280), .A0(shiftedOData[520]), .A1(n4251), .Z(n824));
Q_FDP0UA U9098 ( .D(n823), .QTFCLK( ), .Q(shiftedOData[519]));
Q_MX02 U9099 ( .S(n280), .A0(shiftedOData[519]), .A1(n4250), .Z(n823));
Q_FDP0UA U9100 ( .D(n822), .QTFCLK( ), .Q(shiftedOData[518]));
Q_MX02 U9101 ( .S(n280), .A0(shiftedOData[518]), .A1(n4249), .Z(n822));
Q_FDP0UA U9102 ( .D(n821), .QTFCLK( ), .Q(shiftedOData[517]));
Q_MX02 U9103 ( .S(n280), .A0(shiftedOData[517]), .A1(n4248), .Z(n821));
Q_FDP0UA U9104 ( .D(n820), .QTFCLK( ), .Q(shiftedOData[516]));
Q_MX02 U9105 ( .S(n280), .A0(shiftedOData[516]), .A1(n4247), .Z(n820));
Q_FDP0UA U9106 ( .D(n819), .QTFCLK( ), .Q(shiftedOData[515]));
Q_MX02 U9107 ( .S(n280), .A0(shiftedOData[515]), .A1(n4246), .Z(n819));
Q_FDP0UA U9108 ( .D(n818), .QTFCLK( ), .Q(shiftedOData[514]));
Q_MX02 U9109 ( .S(n280), .A0(shiftedOData[514]), .A1(n4245), .Z(n818));
Q_FDP0UA U9110 ( .D(n817), .QTFCLK( ), .Q(shiftedOData[513]));
Q_MX02 U9111 ( .S(n280), .A0(shiftedOData[513]), .A1(n4244), .Z(n817));
Q_FDP0UA U9112 ( .D(n816), .QTFCLK( ), .Q(shiftedOData[512]));
Q_MX02 U9113 ( .S(n280), .A0(shiftedOData[512]), .A1(n4243), .Z(n816));
Q_FDP0UA U9114 ( .D(n815), .QTFCLK( ), .Q(shiftedOData[511]));
Q_MX02 U9115 ( .S(n280), .A0(shiftedOData[511]), .A1(n4242), .Z(n815));
Q_FDP0UA U9116 ( .D(n814), .QTFCLK( ), .Q(shiftedOData[510]));
Q_MX02 U9117 ( .S(n280), .A0(shiftedOData[510]), .A1(n4241), .Z(n814));
Q_FDP0UA U9118 ( .D(n813), .QTFCLK( ), .Q(shiftedOData[509]));
Q_MX02 U9119 ( .S(n280), .A0(shiftedOData[509]), .A1(n4240), .Z(n813));
Q_FDP0UA U9120 ( .D(n812), .QTFCLK( ), .Q(shiftedOData[508]));
Q_MX02 U9121 ( .S(n280), .A0(shiftedOData[508]), .A1(n4239), .Z(n812));
Q_FDP0UA U9122 ( .D(n811), .QTFCLK( ), .Q(shiftedOData[507]));
Q_MX02 U9123 ( .S(n280), .A0(shiftedOData[507]), .A1(n4238), .Z(n811));
Q_FDP0UA U9124 ( .D(n810), .QTFCLK( ), .Q(shiftedOData[506]));
Q_MX02 U9125 ( .S(n280), .A0(shiftedOData[506]), .A1(n4237), .Z(n810));
Q_FDP0UA U9126 ( .D(n809), .QTFCLK( ), .Q(shiftedOData[505]));
Q_MX02 U9127 ( .S(n280), .A0(shiftedOData[505]), .A1(n4236), .Z(n809));
Q_FDP0UA U9128 ( .D(n808), .QTFCLK( ), .Q(shiftedOData[504]));
Q_MX02 U9129 ( .S(n280), .A0(shiftedOData[504]), .A1(n4235), .Z(n808));
Q_FDP0UA U9130 ( .D(n807), .QTFCLK( ), .Q(shiftedOData[503]));
Q_MX02 U9131 ( .S(n280), .A0(shiftedOData[503]), .A1(n4234), .Z(n807));
Q_FDP0UA U9132 ( .D(n806), .QTFCLK( ), .Q(shiftedOData[502]));
Q_MX02 U9133 ( .S(n280), .A0(shiftedOData[502]), .A1(n4233), .Z(n806));
Q_FDP0UA U9134 ( .D(n805), .QTFCLK( ), .Q(shiftedOData[501]));
Q_MX02 U9135 ( .S(n280), .A0(shiftedOData[501]), .A1(n4232), .Z(n805));
Q_FDP0UA U9136 ( .D(n804), .QTFCLK( ), .Q(shiftedOData[500]));
Q_MX02 U9137 ( .S(n280), .A0(shiftedOData[500]), .A1(n4231), .Z(n804));
Q_FDP0UA U9138 ( .D(n803), .QTFCLK( ), .Q(shiftedOData[499]));
Q_MX02 U9139 ( .S(n280), .A0(shiftedOData[499]), .A1(n4230), .Z(n803));
Q_FDP0UA U9140 ( .D(n802), .QTFCLK( ), .Q(shiftedOData[498]));
Q_MX02 U9141 ( .S(n280), .A0(shiftedOData[498]), .A1(n4229), .Z(n802));
Q_FDP0UA U9142 ( .D(n801), .QTFCLK( ), .Q(shiftedOData[497]));
Q_MX02 U9143 ( .S(n280), .A0(shiftedOData[497]), .A1(n4228), .Z(n801));
Q_FDP0UA U9144 ( .D(n800), .QTFCLK( ), .Q(shiftedOData[496]));
Q_MX02 U9145 ( .S(n280), .A0(shiftedOData[496]), .A1(n4227), .Z(n800));
Q_FDP0UA U9146 ( .D(n799), .QTFCLK( ), .Q(shiftedOData[495]));
Q_MX02 U9147 ( .S(n280), .A0(shiftedOData[495]), .A1(n4226), .Z(n799));
Q_FDP0UA U9148 ( .D(n798), .QTFCLK( ), .Q(shiftedOData[494]));
Q_MX02 U9149 ( .S(n280), .A0(shiftedOData[494]), .A1(n4225), .Z(n798));
Q_FDP0UA U9150 ( .D(n797), .QTFCLK( ), .Q(shiftedOData[493]));
Q_MX02 U9151 ( .S(n280), .A0(shiftedOData[493]), .A1(n4224), .Z(n797));
Q_FDP0UA U9152 ( .D(n796), .QTFCLK( ), .Q(shiftedOData[492]));
Q_MX02 U9153 ( .S(n280), .A0(shiftedOData[492]), .A1(n4223), .Z(n796));
Q_FDP0UA U9154 ( .D(n795), .QTFCLK( ), .Q(shiftedOData[491]));
Q_MX02 U9155 ( .S(n280), .A0(shiftedOData[491]), .A1(n4222), .Z(n795));
Q_FDP0UA U9156 ( .D(n794), .QTFCLK( ), .Q(shiftedOData[490]));
Q_MX02 U9157 ( .S(n280), .A0(shiftedOData[490]), .A1(n4221), .Z(n794));
Q_FDP0UA U9158 ( .D(n793), .QTFCLK( ), .Q(shiftedOData[489]));
Q_MX02 U9159 ( .S(n280), .A0(shiftedOData[489]), .A1(n4220), .Z(n793));
Q_FDP0UA U9160 ( .D(n792), .QTFCLK( ), .Q(shiftedOData[488]));
Q_MX02 U9161 ( .S(n280), .A0(shiftedOData[488]), .A1(n4219), .Z(n792));
Q_FDP0UA U9162 ( .D(n791), .QTFCLK( ), .Q(shiftedOData[487]));
Q_MX02 U9163 ( .S(n280), .A0(shiftedOData[487]), .A1(n4218), .Z(n791));
Q_FDP0UA U9164 ( .D(n790), .QTFCLK( ), .Q(shiftedOData[486]));
Q_MX02 U9165 ( .S(n280), .A0(shiftedOData[486]), .A1(n4217), .Z(n790));
Q_FDP0UA U9166 ( .D(n789), .QTFCLK( ), .Q(shiftedOData[485]));
Q_MX02 U9167 ( .S(n280), .A0(shiftedOData[485]), .A1(n4216), .Z(n789));
Q_FDP0UA U9168 ( .D(n788), .QTFCLK( ), .Q(shiftedOData[484]));
Q_MX02 U9169 ( .S(n280), .A0(shiftedOData[484]), .A1(n4215), .Z(n788));
Q_FDP0UA U9170 ( .D(n787), .QTFCLK( ), .Q(shiftedOData[483]));
Q_MX02 U9171 ( .S(n280), .A0(shiftedOData[483]), .A1(n4214), .Z(n787));
Q_FDP0UA U9172 ( .D(n786), .QTFCLK( ), .Q(shiftedOData[482]));
Q_MX02 U9173 ( .S(n280), .A0(shiftedOData[482]), .A1(n4213), .Z(n786));
Q_FDP0UA U9174 ( .D(n785), .QTFCLK( ), .Q(shiftedOData[481]));
Q_MX02 U9175 ( .S(n280), .A0(shiftedOData[481]), .A1(n4212), .Z(n785));
Q_FDP0UA U9176 ( .D(n784), .QTFCLK( ), .Q(shiftedOData[480]));
Q_MX02 U9177 ( .S(n280), .A0(shiftedOData[480]), .A1(n4211), .Z(n784));
Q_FDP0UA U9178 ( .D(n783), .QTFCLK( ), .Q(shiftedOData[479]));
Q_MX02 U9179 ( .S(n280), .A0(shiftedOData[479]), .A1(n4210), .Z(n783));
Q_FDP0UA U9180 ( .D(n782), .QTFCLK( ), .Q(shiftedOData[478]));
Q_MX02 U9181 ( .S(n280), .A0(shiftedOData[478]), .A1(n4209), .Z(n782));
Q_FDP0UA U9182 ( .D(n781), .QTFCLK( ), .Q(shiftedOData[477]));
Q_MX02 U9183 ( .S(n280), .A0(shiftedOData[477]), .A1(n4208), .Z(n781));
Q_FDP0UA U9184 ( .D(n780), .QTFCLK( ), .Q(shiftedOData[476]));
Q_MX02 U9185 ( .S(n280), .A0(shiftedOData[476]), .A1(n4207), .Z(n780));
Q_FDP0UA U9186 ( .D(n779), .QTFCLK( ), .Q(shiftedOData[475]));
Q_MX02 U9187 ( .S(n280), .A0(shiftedOData[475]), .A1(n4206), .Z(n779));
Q_FDP0UA U9188 ( .D(n778), .QTFCLK( ), .Q(shiftedOData[474]));
Q_MX02 U9189 ( .S(n280), .A0(shiftedOData[474]), .A1(n4205), .Z(n778));
Q_FDP0UA U9190 ( .D(n777), .QTFCLK( ), .Q(shiftedOData[473]));
Q_MX02 U9191 ( .S(n280), .A0(shiftedOData[473]), .A1(n4204), .Z(n777));
Q_FDP0UA U9192 ( .D(n776), .QTFCLK( ), .Q(shiftedOData[472]));
Q_MX02 U9193 ( .S(n280), .A0(shiftedOData[472]), .A1(n4203), .Z(n776));
Q_FDP0UA U9194 ( .D(n775), .QTFCLK( ), .Q(shiftedOData[471]));
Q_MX02 U9195 ( .S(n280), .A0(shiftedOData[471]), .A1(n4202), .Z(n775));
Q_FDP0UA U9196 ( .D(n774), .QTFCLK( ), .Q(shiftedOData[470]));
Q_MX02 U9197 ( .S(n280), .A0(shiftedOData[470]), .A1(n4201), .Z(n774));
Q_FDP0UA U9198 ( .D(n773), .QTFCLK( ), .Q(shiftedOData[469]));
Q_MX02 U9199 ( .S(n280), .A0(shiftedOData[469]), .A1(n4200), .Z(n773));
Q_FDP0UA U9200 ( .D(n772), .QTFCLK( ), .Q(shiftedOData[468]));
Q_MX02 U9201 ( .S(n280), .A0(shiftedOData[468]), .A1(n4199), .Z(n772));
Q_FDP0UA U9202 ( .D(n771), .QTFCLK( ), .Q(shiftedOData[467]));
Q_MX02 U9203 ( .S(n280), .A0(shiftedOData[467]), .A1(n4198), .Z(n771));
Q_FDP0UA U9204 ( .D(n770), .QTFCLK( ), .Q(shiftedOData[466]));
Q_MX02 U9205 ( .S(n280), .A0(shiftedOData[466]), .A1(n4197), .Z(n770));
Q_FDP0UA U9206 ( .D(n769), .QTFCLK( ), .Q(shiftedOData[465]));
Q_MX02 U9207 ( .S(n280), .A0(shiftedOData[465]), .A1(n4196), .Z(n769));
Q_FDP0UA U9208 ( .D(n768), .QTFCLK( ), .Q(shiftedOData[464]));
Q_MX02 U9209 ( .S(n280), .A0(shiftedOData[464]), .A1(n4195), .Z(n768));
Q_FDP0UA U9210 ( .D(n767), .QTFCLK( ), .Q(shiftedOData[463]));
Q_MX02 U9211 ( .S(n280), .A0(shiftedOData[463]), .A1(n4194), .Z(n767));
Q_FDP0UA U9212 ( .D(n766), .QTFCLK( ), .Q(shiftedOData[462]));
Q_MX02 U9213 ( .S(n280), .A0(shiftedOData[462]), .A1(n4193), .Z(n766));
Q_FDP0UA U9214 ( .D(n765), .QTFCLK( ), .Q(shiftedOData[461]));
Q_MX02 U9215 ( .S(n280), .A0(shiftedOData[461]), .A1(n4192), .Z(n765));
Q_FDP0UA U9216 ( .D(n764), .QTFCLK( ), .Q(shiftedOData[460]));
Q_MX02 U9217 ( .S(n280), .A0(shiftedOData[460]), .A1(n4191), .Z(n764));
Q_FDP0UA U9218 ( .D(n763), .QTFCLK( ), .Q(shiftedOData[459]));
Q_MX02 U9219 ( .S(n280), .A0(shiftedOData[459]), .A1(n4190), .Z(n763));
Q_FDP0UA U9220 ( .D(n762), .QTFCLK( ), .Q(shiftedOData[458]));
Q_MX02 U9221 ( .S(n280), .A0(shiftedOData[458]), .A1(n4189), .Z(n762));
Q_FDP0UA U9222 ( .D(n761), .QTFCLK( ), .Q(shiftedOData[457]));
Q_MX02 U9223 ( .S(n280), .A0(shiftedOData[457]), .A1(n4188), .Z(n761));
Q_FDP0UA U9224 ( .D(n760), .QTFCLK( ), .Q(shiftedOData[456]));
Q_MX02 U9225 ( .S(n280), .A0(shiftedOData[456]), .A1(n4187), .Z(n760));
Q_FDP0UA U9226 ( .D(n759), .QTFCLK( ), .Q(shiftedOData[455]));
Q_MX02 U9227 ( .S(n280), .A0(shiftedOData[455]), .A1(n4186), .Z(n759));
Q_FDP0UA U9228 ( .D(n758), .QTFCLK( ), .Q(shiftedOData[454]));
Q_MX02 U9229 ( .S(n280), .A0(shiftedOData[454]), .A1(n4185), .Z(n758));
Q_FDP0UA U9230 ( .D(n757), .QTFCLK( ), .Q(shiftedOData[453]));
Q_MX02 U9231 ( .S(n280), .A0(shiftedOData[453]), .A1(n4184), .Z(n757));
Q_FDP0UA U9232 ( .D(n756), .QTFCLK( ), .Q(shiftedOData[452]));
Q_MX02 U9233 ( .S(n280), .A0(shiftedOData[452]), .A1(n4183), .Z(n756));
Q_FDP0UA U9234 ( .D(n755), .QTFCLK( ), .Q(shiftedOData[451]));
Q_MX02 U9235 ( .S(n280), .A0(shiftedOData[451]), .A1(n4182), .Z(n755));
Q_FDP0UA U9236 ( .D(n754), .QTFCLK( ), .Q(shiftedOData[450]));
Q_MX02 U9237 ( .S(n280), .A0(shiftedOData[450]), .A1(n4181), .Z(n754));
Q_FDP0UA U9238 ( .D(n753), .QTFCLK( ), .Q(shiftedOData[449]));
Q_MX02 U9239 ( .S(n280), .A0(shiftedOData[449]), .A1(n4180), .Z(n753));
Q_FDP0UA U9240 ( .D(n752), .QTFCLK( ), .Q(shiftedOData[448]));
Q_MX02 U9241 ( .S(n280), .A0(shiftedOData[448]), .A1(n4179), .Z(n752));
Q_FDP0UA U9242 ( .D(n751), .QTFCLK( ), .Q(shiftedOData[447]));
Q_MX02 U9243 ( .S(n280), .A0(shiftedOData[447]), .A1(n4178), .Z(n751));
Q_FDP0UA U9244 ( .D(n750), .QTFCLK( ), .Q(shiftedOData[446]));
Q_MX02 U9245 ( .S(n280), .A0(shiftedOData[446]), .A1(n4177), .Z(n750));
Q_FDP0UA U9246 ( .D(n749), .QTFCLK( ), .Q(shiftedOData[445]));
Q_MX02 U9247 ( .S(n280), .A0(shiftedOData[445]), .A1(n4176), .Z(n749));
Q_FDP0UA U9248 ( .D(n748), .QTFCLK( ), .Q(shiftedOData[444]));
Q_MX02 U9249 ( .S(n280), .A0(shiftedOData[444]), .A1(n4175), .Z(n748));
Q_FDP0UA U9250 ( .D(n747), .QTFCLK( ), .Q(shiftedOData[443]));
Q_MX02 U9251 ( .S(n280), .A0(shiftedOData[443]), .A1(n4174), .Z(n747));
Q_FDP0UA U9252 ( .D(n746), .QTFCLK( ), .Q(shiftedOData[442]));
Q_MX02 U9253 ( .S(n280), .A0(shiftedOData[442]), .A1(n4173), .Z(n746));
Q_FDP0UA U9254 ( .D(n745), .QTFCLK( ), .Q(shiftedOData[441]));
Q_MX02 U9255 ( .S(n280), .A0(shiftedOData[441]), .A1(n4172), .Z(n745));
Q_FDP0UA U9256 ( .D(n744), .QTFCLK( ), .Q(shiftedOData[440]));
Q_MX02 U9257 ( .S(n280), .A0(shiftedOData[440]), .A1(n4171), .Z(n744));
Q_FDP0UA U9258 ( .D(n743), .QTFCLK( ), .Q(shiftedOData[439]));
Q_MX02 U9259 ( .S(n280), .A0(shiftedOData[439]), .A1(n4170), .Z(n743));
Q_FDP0UA U9260 ( .D(n742), .QTFCLK( ), .Q(shiftedOData[438]));
Q_MX02 U9261 ( .S(n280), .A0(shiftedOData[438]), .A1(n4169), .Z(n742));
Q_FDP0UA U9262 ( .D(n741), .QTFCLK( ), .Q(shiftedOData[437]));
Q_MX02 U9263 ( .S(n280), .A0(shiftedOData[437]), .A1(n4168), .Z(n741));
Q_FDP0UA U9264 ( .D(n740), .QTFCLK( ), .Q(shiftedOData[436]));
Q_MX02 U9265 ( .S(n280), .A0(shiftedOData[436]), .A1(n4167), .Z(n740));
Q_FDP0UA U9266 ( .D(n739), .QTFCLK( ), .Q(shiftedOData[435]));
Q_MX02 U9267 ( .S(n280), .A0(shiftedOData[435]), .A1(n4166), .Z(n739));
Q_FDP0UA U9268 ( .D(n738), .QTFCLK( ), .Q(shiftedOData[434]));
Q_MX02 U9269 ( .S(n280), .A0(shiftedOData[434]), .A1(n4165), .Z(n738));
Q_FDP0UA U9270 ( .D(n737), .QTFCLK( ), .Q(shiftedOData[433]));
Q_MX02 U9271 ( .S(n280), .A0(shiftedOData[433]), .A1(n4164), .Z(n737));
Q_FDP0UA U9272 ( .D(n736), .QTFCLK( ), .Q(shiftedOData[432]));
Q_MX02 U9273 ( .S(n280), .A0(shiftedOData[432]), .A1(n4163), .Z(n736));
Q_FDP0UA U9274 ( .D(n735), .QTFCLK( ), .Q(shiftedOData[431]));
Q_MX02 U9275 ( .S(n280), .A0(shiftedOData[431]), .A1(n4162), .Z(n735));
Q_FDP0UA U9276 ( .D(n734), .QTFCLK( ), .Q(shiftedOData[430]));
Q_MX02 U9277 ( .S(n280), .A0(shiftedOData[430]), .A1(n4161), .Z(n734));
Q_FDP0UA U9278 ( .D(n733), .QTFCLK( ), .Q(shiftedOData[429]));
Q_MX02 U9279 ( .S(n280), .A0(shiftedOData[429]), .A1(n4160), .Z(n733));
Q_FDP0UA U9280 ( .D(n732), .QTFCLK( ), .Q(shiftedOData[428]));
Q_MX02 U9281 ( .S(n280), .A0(shiftedOData[428]), .A1(n4159), .Z(n732));
Q_FDP0UA U9282 ( .D(n731), .QTFCLK( ), .Q(shiftedOData[427]));
Q_MX02 U9283 ( .S(n280), .A0(shiftedOData[427]), .A1(n4158), .Z(n731));
Q_FDP0UA U9284 ( .D(n730), .QTFCLK( ), .Q(shiftedOData[426]));
Q_MX02 U9285 ( .S(n280), .A0(shiftedOData[426]), .A1(n4157), .Z(n730));
Q_FDP0UA U9286 ( .D(n729), .QTFCLK( ), .Q(shiftedOData[425]));
Q_MX02 U9287 ( .S(n280), .A0(shiftedOData[425]), .A1(n4156), .Z(n729));
Q_FDP0UA U9288 ( .D(n728), .QTFCLK( ), .Q(shiftedOData[424]));
Q_MX02 U9289 ( .S(n280), .A0(shiftedOData[424]), .A1(n4155), .Z(n728));
Q_FDP0UA U9290 ( .D(n727), .QTFCLK( ), .Q(shiftedOData[423]));
Q_MX02 U9291 ( .S(n280), .A0(shiftedOData[423]), .A1(n4154), .Z(n727));
Q_FDP0UA U9292 ( .D(n726), .QTFCLK( ), .Q(shiftedOData[422]));
Q_MX02 U9293 ( .S(n280), .A0(shiftedOData[422]), .A1(n4153), .Z(n726));
Q_FDP0UA U9294 ( .D(n725), .QTFCLK( ), .Q(shiftedOData[421]));
Q_MX02 U9295 ( .S(n280), .A0(shiftedOData[421]), .A1(n4152), .Z(n725));
Q_FDP0UA U9296 ( .D(n724), .QTFCLK( ), .Q(shiftedOData[420]));
Q_MX02 U9297 ( .S(n280), .A0(shiftedOData[420]), .A1(n4151), .Z(n724));
Q_FDP0UA U9298 ( .D(n723), .QTFCLK( ), .Q(shiftedOData[419]));
Q_MX02 U9299 ( .S(n280), .A0(shiftedOData[419]), .A1(n4150), .Z(n723));
Q_FDP0UA U9300 ( .D(n722), .QTFCLK( ), .Q(shiftedOData[418]));
Q_MX02 U9301 ( .S(n280), .A0(shiftedOData[418]), .A1(n4149), .Z(n722));
Q_FDP0UA U9302 ( .D(n721), .QTFCLK( ), .Q(shiftedOData[417]));
Q_MX02 U9303 ( .S(n280), .A0(shiftedOData[417]), .A1(n4148), .Z(n721));
Q_FDP0UA U9304 ( .D(n720), .QTFCLK( ), .Q(shiftedOData[416]));
Q_MX02 U9305 ( .S(n280), .A0(shiftedOData[416]), .A1(n4147), .Z(n720));
Q_FDP0UA U9306 ( .D(n719), .QTFCLK( ), .Q(shiftedOData[415]));
Q_MX02 U9307 ( .S(n280), .A0(shiftedOData[415]), .A1(n4146), .Z(n719));
Q_FDP0UA U9308 ( .D(n718), .QTFCLK( ), .Q(shiftedOData[414]));
Q_MX02 U9309 ( .S(n280), .A0(shiftedOData[414]), .A1(n4145), .Z(n718));
Q_FDP0UA U9310 ( .D(n717), .QTFCLK( ), .Q(shiftedOData[413]));
Q_MX02 U9311 ( .S(n280), .A0(shiftedOData[413]), .A1(n4144), .Z(n717));
Q_FDP0UA U9312 ( .D(n716), .QTFCLK( ), .Q(shiftedOData[412]));
Q_MX02 U9313 ( .S(n280), .A0(shiftedOData[412]), .A1(n4143), .Z(n716));
Q_FDP0UA U9314 ( .D(n715), .QTFCLK( ), .Q(shiftedOData[411]));
Q_MX02 U9315 ( .S(n280), .A0(shiftedOData[411]), .A1(n4142), .Z(n715));
Q_FDP0UA U9316 ( .D(n714), .QTFCLK( ), .Q(shiftedOData[410]));
Q_MX02 U9317 ( .S(n280), .A0(shiftedOData[410]), .A1(n4141), .Z(n714));
Q_FDP0UA U9318 ( .D(n713), .QTFCLK( ), .Q(shiftedOData[409]));
Q_MX02 U9319 ( .S(n280), .A0(shiftedOData[409]), .A1(n4140), .Z(n713));
Q_FDP0UA U9320 ( .D(n712), .QTFCLK( ), .Q(shiftedOData[408]));
Q_MX02 U9321 ( .S(n280), .A0(shiftedOData[408]), .A1(n4139), .Z(n712));
Q_FDP0UA U9322 ( .D(n711), .QTFCLK( ), .Q(shiftedOData[407]));
Q_MX02 U9323 ( .S(n280), .A0(shiftedOData[407]), .A1(n4138), .Z(n711));
Q_FDP0UA U9324 ( .D(n710), .QTFCLK( ), .Q(shiftedOData[406]));
Q_MX02 U9325 ( .S(n280), .A0(shiftedOData[406]), .A1(n4137), .Z(n710));
Q_FDP0UA U9326 ( .D(n709), .QTFCLK( ), .Q(shiftedOData[405]));
Q_MX02 U9327 ( .S(n280), .A0(shiftedOData[405]), .A1(n4136), .Z(n709));
Q_FDP0UA U9328 ( .D(n708), .QTFCLK( ), .Q(shiftedOData[404]));
Q_MX02 U9329 ( .S(n280), .A0(shiftedOData[404]), .A1(n4135), .Z(n708));
Q_FDP0UA U9330 ( .D(n707), .QTFCLK( ), .Q(shiftedOData[403]));
Q_MX02 U9331 ( .S(n280), .A0(shiftedOData[403]), .A1(n4134), .Z(n707));
Q_FDP0UA U9332 ( .D(n706), .QTFCLK( ), .Q(shiftedOData[402]));
Q_MX02 U9333 ( .S(n280), .A0(shiftedOData[402]), .A1(n4133), .Z(n706));
Q_FDP0UA U9334 ( .D(n705), .QTFCLK( ), .Q(shiftedOData[401]));
Q_MX02 U9335 ( .S(n280), .A0(shiftedOData[401]), .A1(n4132), .Z(n705));
Q_FDP0UA U9336 ( .D(n704), .QTFCLK( ), .Q(shiftedOData[400]));
Q_MX02 U9337 ( .S(n280), .A0(shiftedOData[400]), .A1(n4131), .Z(n704));
Q_FDP0UA U9338 ( .D(n703), .QTFCLK( ), .Q(shiftedOData[399]));
Q_MX02 U9339 ( .S(n280), .A0(shiftedOData[399]), .A1(n4130), .Z(n703));
Q_FDP0UA U9340 ( .D(n702), .QTFCLK( ), .Q(shiftedOData[398]));
Q_MX02 U9341 ( .S(n280), .A0(shiftedOData[398]), .A1(n4129), .Z(n702));
Q_FDP0UA U9342 ( .D(n701), .QTFCLK( ), .Q(shiftedOData[397]));
Q_MX02 U9343 ( .S(n280), .A0(shiftedOData[397]), .A1(n4128), .Z(n701));
Q_FDP0UA U9344 ( .D(n700), .QTFCLK( ), .Q(shiftedOData[396]));
Q_MX02 U9345 ( .S(n280), .A0(shiftedOData[396]), .A1(n4127), .Z(n700));
Q_FDP0UA U9346 ( .D(n699), .QTFCLK( ), .Q(shiftedOData[395]));
Q_MX02 U9347 ( .S(n280), .A0(shiftedOData[395]), .A1(n4126), .Z(n699));
Q_FDP0UA U9348 ( .D(n698), .QTFCLK( ), .Q(shiftedOData[394]));
Q_MX02 U9349 ( .S(n280), .A0(shiftedOData[394]), .A1(n4125), .Z(n698));
Q_FDP0UA U9350 ( .D(n697), .QTFCLK( ), .Q(shiftedOData[393]));
Q_MX02 U9351 ( .S(n280), .A0(shiftedOData[393]), .A1(n4124), .Z(n697));
Q_FDP0UA U9352 ( .D(n696), .QTFCLK( ), .Q(shiftedOData[392]));
Q_MX02 U9353 ( .S(n280), .A0(shiftedOData[392]), .A1(n4123), .Z(n696));
Q_FDP0UA U9354 ( .D(n695), .QTFCLK( ), .Q(shiftedOData[391]));
Q_MX02 U9355 ( .S(n280), .A0(shiftedOData[391]), .A1(n4122), .Z(n695));
Q_FDP0UA U9356 ( .D(n694), .QTFCLK( ), .Q(shiftedOData[390]));
Q_MX02 U9357 ( .S(n280), .A0(shiftedOData[390]), .A1(n4121), .Z(n694));
Q_FDP0UA U9358 ( .D(n693), .QTFCLK( ), .Q(shiftedOData[389]));
Q_MX02 U9359 ( .S(n280), .A0(shiftedOData[389]), .A1(n4120), .Z(n693));
Q_FDP0UA U9360 ( .D(n692), .QTFCLK( ), .Q(shiftedOData[388]));
Q_MX02 U9361 ( .S(n280), .A0(shiftedOData[388]), .A1(n4119), .Z(n692));
Q_FDP0UA U9362 ( .D(n691), .QTFCLK( ), .Q(shiftedOData[387]));
Q_MX02 U9363 ( .S(n280), .A0(shiftedOData[387]), .A1(n4118), .Z(n691));
Q_FDP0UA U9364 ( .D(n690), .QTFCLK( ), .Q(shiftedOData[386]));
Q_MX02 U9365 ( .S(n280), .A0(shiftedOData[386]), .A1(n4117), .Z(n690));
Q_FDP0UA U9366 ( .D(n689), .QTFCLK( ), .Q(shiftedOData[385]));
Q_MX02 U9367 ( .S(n280), .A0(shiftedOData[385]), .A1(n4116), .Z(n689));
Q_FDP0UA U9368 ( .D(n688), .QTFCLK( ), .Q(shiftedOData[384]));
Q_MX02 U9369 ( .S(n280), .A0(shiftedOData[384]), .A1(n4115), .Z(n688));
Q_FDP0UA U9370 ( .D(n687), .QTFCLK( ), .Q(shiftedOData[383]));
Q_MX02 U9371 ( .S(n280), .A0(shiftedOData[383]), .A1(n4114), .Z(n687));
Q_FDP0UA U9372 ( .D(n686), .QTFCLK( ), .Q(shiftedOData[382]));
Q_MX02 U9373 ( .S(n280), .A0(shiftedOData[382]), .A1(n4113), .Z(n686));
Q_FDP0UA U9374 ( .D(n685), .QTFCLK( ), .Q(shiftedOData[381]));
Q_MX02 U9375 ( .S(n280), .A0(shiftedOData[381]), .A1(n4112), .Z(n685));
Q_FDP0UA U9376 ( .D(n684), .QTFCLK( ), .Q(shiftedOData[380]));
Q_MX02 U9377 ( .S(n280), .A0(shiftedOData[380]), .A1(n4111), .Z(n684));
Q_FDP0UA U9378 ( .D(n683), .QTFCLK( ), .Q(shiftedOData[379]));
Q_MX02 U9379 ( .S(n280), .A0(shiftedOData[379]), .A1(n4110), .Z(n683));
Q_FDP0UA U9380 ( .D(n682), .QTFCLK( ), .Q(shiftedOData[378]));
Q_MX02 U9381 ( .S(n280), .A0(shiftedOData[378]), .A1(n4109), .Z(n682));
Q_FDP0UA U9382 ( .D(n681), .QTFCLK( ), .Q(shiftedOData[377]));
Q_MX02 U9383 ( .S(n280), .A0(shiftedOData[377]), .A1(n4108), .Z(n681));
Q_FDP0UA U9384 ( .D(n680), .QTFCLK( ), .Q(shiftedOData[376]));
Q_MX02 U9385 ( .S(n280), .A0(shiftedOData[376]), .A1(n4107), .Z(n680));
Q_FDP0UA U9386 ( .D(n679), .QTFCLK( ), .Q(shiftedOData[375]));
Q_MX02 U9387 ( .S(n280), .A0(shiftedOData[375]), .A1(n4106), .Z(n679));
Q_FDP0UA U9388 ( .D(n678), .QTFCLK( ), .Q(shiftedOData[374]));
Q_MX02 U9389 ( .S(n280), .A0(shiftedOData[374]), .A1(n4105), .Z(n678));
Q_FDP0UA U9390 ( .D(n677), .QTFCLK( ), .Q(shiftedOData[373]));
Q_MX02 U9391 ( .S(n280), .A0(shiftedOData[373]), .A1(n4104), .Z(n677));
Q_FDP0UA U9392 ( .D(n676), .QTFCLK( ), .Q(shiftedOData[372]));
Q_MX02 U9393 ( .S(n280), .A0(shiftedOData[372]), .A1(n4103), .Z(n676));
Q_FDP0UA U9394 ( .D(n675), .QTFCLK( ), .Q(shiftedOData[371]));
Q_MX02 U9395 ( .S(n280), .A0(shiftedOData[371]), .A1(n4102), .Z(n675));
Q_FDP0UA U9396 ( .D(n674), .QTFCLK( ), .Q(shiftedOData[370]));
Q_MX02 U9397 ( .S(n280), .A0(shiftedOData[370]), .A1(n4101), .Z(n674));
Q_FDP0UA U9398 ( .D(n673), .QTFCLK( ), .Q(shiftedOData[369]));
Q_MX02 U9399 ( .S(n280), .A0(shiftedOData[369]), .A1(n4100), .Z(n673));
Q_FDP0UA U9400 ( .D(n672), .QTFCLK( ), .Q(shiftedOData[368]));
Q_MX02 U9401 ( .S(n280), .A0(shiftedOData[368]), .A1(n4099), .Z(n672));
Q_FDP0UA U9402 ( .D(n671), .QTFCLK( ), .Q(shiftedOData[367]));
Q_MX02 U9403 ( .S(n280), .A0(shiftedOData[367]), .A1(n4098), .Z(n671));
Q_FDP0UA U9404 ( .D(n670), .QTFCLK( ), .Q(shiftedOData[366]));
Q_MX02 U9405 ( .S(n280), .A0(shiftedOData[366]), .A1(n4097), .Z(n670));
Q_FDP0UA U9406 ( .D(n669), .QTFCLK( ), .Q(shiftedOData[365]));
Q_MX02 U9407 ( .S(n280), .A0(shiftedOData[365]), .A1(n4096), .Z(n669));
Q_FDP0UA U9408 ( .D(n668), .QTFCLK( ), .Q(shiftedOData[364]));
Q_MX02 U9409 ( .S(n280), .A0(shiftedOData[364]), .A1(n4095), .Z(n668));
Q_FDP0UA U9410 ( .D(n667), .QTFCLK( ), .Q(shiftedOData[363]));
Q_MX02 U9411 ( .S(n280), .A0(shiftedOData[363]), .A1(n4094), .Z(n667));
Q_FDP0UA U9412 ( .D(n666), .QTFCLK( ), .Q(shiftedOData[362]));
Q_MX02 U9413 ( .S(n280), .A0(shiftedOData[362]), .A1(n4093), .Z(n666));
Q_FDP0UA U9414 ( .D(n665), .QTFCLK( ), .Q(shiftedOData[361]));
Q_MX02 U9415 ( .S(n280), .A0(shiftedOData[361]), .A1(n4092), .Z(n665));
Q_FDP0UA U9416 ( .D(n664), .QTFCLK( ), .Q(shiftedOData[360]));
Q_MX02 U9417 ( .S(n280), .A0(shiftedOData[360]), .A1(n4091), .Z(n664));
Q_FDP0UA U9418 ( .D(n663), .QTFCLK( ), .Q(shiftedOData[359]));
Q_MX02 U9419 ( .S(n280), .A0(shiftedOData[359]), .A1(n4090), .Z(n663));
Q_FDP0UA U9420 ( .D(n662), .QTFCLK( ), .Q(shiftedOData[358]));
Q_MX02 U9421 ( .S(n280), .A0(shiftedOData[358]), .A1(n4089), .Z(n662));
Q_FDP0UA U9422 ( .D(n661), .QTFCLK( ), .Q(shiftedOData[357]));
Q_MX02 U9423 ( .S(n280), .A0(shiftedOData[357]), .A1(n4088), .Z(n661));
Q_FDP0UA U9424 ( .D(n660), .QTFCLK( ), .Q(shiftedOData[356]));
Q_MX02 U9425 ( .S(n280), .A0(shiftedOData[356]), .A1(n4087), .Z(n660));
Q_FDP0UA U9426 ( .D(n659), .QTFCLK( ), .Q(shiftedOData[355]));
Q_MX02 U9427 ( .S(n280), .A0(shiftedOData[355]), .A1(n4086), .Z(n659));
Q_FDP0UA U9428 ( .D(n658), .QTFCLK( ), .Q(shiftedOData[354]));
Q_MX02 U9429 ( .S(n280), .A0(shiftedOData[354]), .A1(n4085), .Z(n658));
Q_FDP0UA U9430 ( .D(n657), .QTFCLK( ), .Q(shiftedOData[353]));
Q_MX02 U9431 ( .S(n280), .A0(shiftedOData[353]), .A1(n4084), .Z(n657));
Q_FDP0UA U9432 ( .D(n656), .QTFCLK( ), .Q(shiftedOData[352]));
Q_MX02 U9433 ( .S(n280), .A0(shiftedOData[352]), .A1(n4083), .Z(n656));
Q_FDP0UA U9434 ( .D(n655), .QTFCLK( ), .Q(shiftedOData[351]));
Q_MX02 U9435 ( .S(n280), .A0(shiftedOData[351]), .A1(n4082), .Z(n655));
Q_FDP0UA U9436 ( .D(n654), .QTFCLK( ), .Q(shiftedOData[350]));
Q_MX02 U9437 ( .S(n280), .A0(shiftedOData[350]), .A1(n4081), .Z(n654));
Q_FDP0UA U9438 ( .D(n653), .QTFCLK( ), .Q(shiftedOData[349]));
Q_MX02 U9439 ( .S(n280), .A0(shiftedOData[349]), .A1(n4080), .Z(n653));
Q_FDP0UA U9440 ( .D(n652), .QTFCLK( ), .Q(shiftedOData[348]));
Q_MX02 U9441 ( .S(n280), .A0(shiftedOData[348]), .A1(n4079), .Z(n652));
Q_FDP0UA U9442 ( .D(n651), .QTFCLK( ), .Q(shiftedOData[347]));
Q_MX02 U9443 ( .S(n280), .A0(shiftedOData[347]), .A1(n4078), .Z(n651));
Q_FDP0UA U9444 ( .D(n650), .QTFCLK( ), .Q(shiftedOData[346]));
Q_MX02 U9445 ( .S(n280), .A0(shiftedOData[346]), .A1(n4077), .Z(n650));
Q_FDP0UA U9446 ( .D(n649), .QTFCLK( ), .Q(shiftedOData[345]));
Q_MX02 U9447 ( .S(n280), .A0(shiftedOData[345]), .A1(n4076), .Z(n649));
Q_FDP0UA U9448 ( .D(n648), .QTFCLK( ), .Q(shiftedOData[344]));
Q_MX02 U9449 ( .S(n280), .A0(shiftedOData[344]), .A1(n4075), .Z(n648));
Q_FDP0UA U9450 ( .D(n647), .QTFCLK( ), .Q(shiftedOData[343]));
Q_MX02 U9451 ( .S(n280), .A0(shiftedOData[343]), .A1(n4074), .Z(n647));
Q_FDP0UA U9452 ( .D(n646), .QTFCLK( ), .Q(shiftedOData[342]));
Q_MX02 U9453 ( .S(n280), .A0(shiftedOData[342]), .A1(n4073), .Z(n646));
Q_FDP0UA U9454 ( .D(n645), .QTFCLK( ), .Q(shiftedOData[341]));
Q_MX02 U9455 ( .S(n280), .A0(shiftedOData[341]), .A1(n4072), .Z(n645));
Q_FDP0UA U9456 ( .D(n644), .QTFCLK( ), .Q(shiftedOData[340]));
Q_MX02 U9457 ( .S(n280), .A0(shiftedOData[340]), .A1(n4071), .Z(n644));
Q_FDP0UA U9458 ( .D(n643), .QTFCLK( ), .Q(shiftedOData[339]));
Q_MX02 U9459 ( .S(n280), .A0(shiftedOData[339]), .A1(n4070), .Z(n643));
Q_FDP0UA U9460 ( .D(n642), .QTFCLK( ), .Q(shiftedOData[338]));
Q_MX02 U9461 ( .S(n280), .A0(shiftedOData[338]), .A1(n4069), .Z(n642));
Q_FDP0UA U9462 ( .D(n641), .QTFCLK( ), .Q(shiftedOData[337]));
Q_MX02 U9463 ( .S(n280), .A0(shiftedOData[337]), .A1(n4068), .Z(n641));
Q_FDP0UA U9464 ( .D(n640), .QTFCLK( ), .Q(shiftedOData[336]));
Q_MX02 U9465 ( .S(n280), .A0(shiftedOData[336]), .A1(n4067), .Z(n640));
Q_FDP0UA U9466 ( .D(n639), .QTFCLK( ), .Q(shiftedOData[335]));
Q_MX02 U9467 ( .S(n280), .A0(shiftedOData[335]), .A1(n4066), .Z(n639));
Q_FDP0UA U9468 ( .D(n638), .QTFCLK( ), .Q(shiftedOData[334]));
Q_MX02 U9469 ( .S(n280), .A0(shiftedOData[334]), .A1(n4065), .Z(n638));
Q_FDP0UA U9470 ( .D(n637), .QTFCLK( ), .Q(shiftedOData[333]));
Q_MX02 U9471 ( .S(n280), .A0(shiftedOData[333]), .A1(n4064), .Z(n637));
Q_FDP0UA U9472 ( .D(n636), .QTFCLK( ), .Q(shiftedOData[332]));
Q_MX02 U9473 ( .S(n280), .A0(shiftedOData[332]), .A1(n4063), .Z(n636));
Q_FDP0UA U9474 ( .D(n635), .QTFCLK( ), .Q(shiftedOData[331]));
Q_MX02 U9475 ( .S(n280), .A0(shiftedOData[331]), .A1(n4062), .Z(n635));
Q_FDP0UA U9476 ( .D(n634), .QTFCLK( ), .Q(shiftedOData[330]));
Q_MX02 U9477 ( .S(n280), .A0(shiftedOData[330]), .A1(n4061), .Z(n634));
Q_FDP0UA U9478 ( .D(n633), .QTFCLK( ), .Q(shiftedOData[329]));
Q_MX02 U9479 ( .S(n280), .A0(shiftedOData[329]), .A1(n4060), .Z(n633));
Q_FDP0UA U9480 ( .D(n632), .QTFCLK( ), .Q(shiftedOData[328]));
Q_MX02 U9481 ( .S(n280), .A0(shiftedOData[328]), .A1(n4059), .Z(n632));
Q_FDP0UA U9482 ( .D(n631), .QTFCLK( ), .Q(shiftedOData[327]));
Q_MX02 U9483 ( .S(n280), .A0(shiftedOData[327]), .A1(n4058), .Z(n631));
Q_FDP0UA U9484 ( .D(n630), .QTFCLK( ), .Q(shiftedOData[326]));
Q_MX02 U9485 ( .S(n280), .A0(shiftedOData[326]), .A1(n4057), .Z(n630));
Q_FDP0UA U9486 ( .D(n629), .QTFCLK( ), .Q(shiftedOData[325]));
Q_MX02 U9487 ( .S(n280), .A0(shiftedOData[325]), .A1(n4056), .Z(n629));
Q_FDP0UA U9488 ( .D(n628), .QTFCLK( ), .Q(shiftedOData[324]));
Q_MX02 U9489 ( .S(n280), .A0(shiftedOData[324]), .A1(n4055), .Z(n628));
Q_FDP0UA U9490 ( .D(n627), .QTFCLK( ), .Q(shiftedOData[323]));
Q_MX02 U9491 ( .S(n280), .A0(shiftedOData[323]), .A1(n4054), .Z(n627));
Q_FDP0UA U9492 ( .D(n626), .QTFCLK( ), .Q(shiftedOData[322]));
Q_MX02 U9493 ( .S(n280), .A0(shiftedOData[322]), .A1(n4053), .Z(n626));
Q_FDP0UA U9494 ( .D(n625), .QTFCLK( ), .Q(shiftedOData[321]));
Q_MX02 U9495 ( .S(n280), .A0(shiftedOData[321]), .A1(n4052), .Z(n625));
Q_FDP0UA U9496 ( .D(n624), .QTFCLK( ), .Q(shiftedOData[320]));
Q_MX02 U9497 ( .S(n280), .A0(shiftedOData[320]), .A1(n4051), .Z(n624));
Q_FDP0UA U9498 ( .D(n623), .QTFCLK( ), .Q(shiftedOData[319]));
Q_MX02 U9499 ( .S(n280), .A0(shiftedOData[319]), .A1(n4050), .Z(n623));
Q_FDP0UA U9500 ( .D(n622), .QTFCLK( ), .Q(shiftedOData[318]));
Q_MX02 U9501 ( .S(n280), .A0(shiftedOData[318]), .A1(n4049), .Z(n622));
Q_FDP0UA U9502 ( .D(n621), .QTFCLK( ), .Q(shiftedOData[317]));
Q_MX02 U9503 ( .S(n280), .A0(shiftedOData[317]), .A1(n4048), .Z(n621));
Q_FDP0UA U9504 ( .D(n620), .QTFCLK( ), .Q(shiftedOData[316]));
Q_MX02 U9505 ( .S(n280), .A0(shiftedOData[316]), .A1(n4047), .Z(n620));
Q_FDP0UA U9506 ( .D(n619), .QTFCLK( ), .Q(shiftedOData[315]));
Q_MX02 U9507 ( .S(n280), .A0(shiftedOData[315]), .A1(n4046), .Z(n619));
Q_FDP0UA U9508 ( .D(n618), .QTFCLK( ), .Q(shiftedOData[314]));
Q_MX02 U9509 ( .S(n280), .A0(shiftedOData[314]), .A1(n4045), .Z(n618));
Q_FDP0UA U9510 ( .D(n617), .QTFCLK( ), .Q(shiftedOData[313]));
Q_MX02 U9511 ( .S(n280), .A0(shiftedOData[313]), .A1(n4044), .Z(n617));
Q_FDP0UA U9512 ( .D(n616), .QTFCLK( ), .Q(shiftedOData[312]));
Q_MX02 U9513 ( .S(n280), .A0(shiftedOData[312]), .A1(n4043), .Z(n616));
Q_FDP0UA U9514 ( .D(n615), .QTFCLK( ), .Q(shiftedOData[311]));
Q_MX02 U9515 ( .S(n280), .A0(shiftedOData[311]), .A1(n4042), .Z(n615));
Q_FDP0UA U9516 ( .D(n614), .QTFCLK( ), .Q(shiftedOData[310]));
Q_MX02 U9517 ( .S(n280), .A0(shiftedOData[310]), .A1(n4041), .Z(n614));
Q_FDP0UA U9518 ( .D(n613), .QTFCLK( ), .Q(shiftedOData[309]));
Q_MX02 U9519 ( .S(n280), .A0(shiftedOData[309]), .A1(n4040), .Z(n613));
Q_FDP0UA U9520 ( .D(n612), .QTFCLK( ), .Q(shiftedOData[308]));
Q_MX02 U9521 ( .S(n280), .A0(shiftedOData[308]), .A1(n4039), .Z(n612));
Q_FDP0UA U9522 ( .D(n611), .QTFCLK( ), .Q(shiftedOData[307]));
Q_MX02 U9523 ( .S(n280), .A0(shiftedOData[307]), .A1(n4038), .Z(n611));
Q_FDP0UA U9524 ( .D(n610), .QTFCLK( ), .Q(shiftedOData[306]));
Q_MX02 U9525 ( .S(n280), .A0(shiftedOData[306]), .A1(n4037), .Z(n610));
Q_FDP0UA U9526 ( .D(n609), .QTFCLK( ), .Q(shiftedOData[305]));
Q_MX02 U9527 ( .S(n280), .A0(shiftedOData[305]), .A1(n4036), .Z(n609));
Q_FDP0UA U9528 ( .D(n608), .QTFCLK( ), .Q(shiftedOData[304]));
Q_MX02 U9529 ( .S(n280), .A0(shiftedOData[304]), .A1(n4035), .Z(n608));
Q_FDP0UA U9530 ( .D(n607), .QTFCLK( ), .Q(shiftedOData[303]));
Q_MX02 U9531 ( .S(n280), .A0(shiftedOData[303]), .A1(n4034), .Z(n607));
Q_FDP0UA U9532 ( .D(n606), .QTFCLK( ), .Q(shiftedOData[302]));
Q_MX02 U9533 ( .S(n280), .A0(shiftedOData[302]), .A1(n4033), .Z(n606));
Q_FDP0UA U9534 ( .D(n605), .QTFCLK( ), .Q(shiftedOData[301]));
Q_MX02 U9535 ( .S(n280), .A0(shiftedOData[301]), .A1(n4032), .Z(n605));
Q_FDP0UA U9536 ( .D(n604), .QTFCLK( ), .Q(shiftedOData[300]));
Q_MX02 U9537 ( .S(n280), .A0(shiftedOData[300]), .A1(n4031), .Z(n604));
Q_FDP0UA U9538 ( .D(n603), .QTFCLK( ), .Q(shiftedOData[299]));
Q_MX02 U9539 ( .S(n280), .A0(shiftedOData[299]), .A1(n4030), .Z(n603));
Q_FDP0UA U9540 ( .D(n602), .QTFCLK( ), .Q(shiftedOData[298]));
Q_MX02 U9541 ( .S(n280), .A0(shiftedOData[298]), .A1(n4029), .Z(n602));
Q_FDP0UA U9542 ( .D(n601), .QTFCLK( ), .Q(shiftedOData[297]));
Q_MX02 U9543 ( .S(n280), .A0(shiftedOData[297]), .A1(n4028), .Z(n601));
Q_FDP0UA U9544 ( .D(n600), .QTFCLK( ), .Q(shiftedOData[296]));
Q_MX02 U9545 ( .S(n280), .A0(shiftedOData[296]), .A1(n4027), .Z(n600));
Q_FDP0UA U9546 ( .D(n599), .QTFCLK( ), .Q(shiftedOData[295]));
Q_MX02 U9547 ( .S(n280), .A0(shiftedOData[295]), .A1(n4026), .Z(n599));
Q_FDP0UA U9548 ( .D(n598), .QTFCLK( ), .Q(shiftedOData[294]));
Q_MX02 U9549 ( .S(n280), .A0(shiftedOData[294]), .A1(n4025), .Z(n598));
Q_FDP0UA U9550 ( .D(n597), .QTFCLK( ), .Q(shiftedOData[293]));
Q_MX02 U9551 ( .S(n280), .A0(shiftedOData[293]), .A1(n4024), .Z(n597));
Q_FDP0UA U9552 ( .D(n596), .QTFCLK( ), .Q(shiftedOData[292]));
Q_MX02 U9553 ( .S(n280), .A0(shiftedOData[292]), .A1(n4023), .Z(n596));
Q_FDP0UA U9554 ( .D(n595), .QTFCLK( ), .Q(shiftedOData[291]));
Q_MX02 U9555 ( .S(n280), .A0(shiftedOData[291]), .A1(n4022), .Z(n595));
Q_FDP0UA U9556 ( .D(n594), .QTFCLK( ), .Q(shiftedOData[290]));
Q_MX02 U9557 ( .S(n280), .A0(shiftedOData[290]), .A1(n4021), .Z(n594));
Q_FDP0UA U9558 ( .D(n593), .QTFCLK( ), .Q(shiftedOData[289]));
Q_MX02 U9559 ( .S(n280), .A0(shiftedOData[289]), .A1(n4020), .Z(n593));
Q_FDP0UA U9560 ( .D(n592), .QTFCLK( ), .Q(shiftedOData[288]));
Q_MX02 U9561 ( .S(n280), .A0(shiftedOData[288]), .A1(n4019), .Z(n592));
Q_FDP0UA U9562 ( .D(n591), .QTFCLK( ), .Q(shiftedOData[287]));
Q_MX02 U9563 ( .S(n280), .A0(shiftedOData[287]), .A1(n4018), .Z(n591));
Q_FDP0UA U9564 ( .D(n590), .QTFCLK( ), .Q(shiftedOData[286]));
Q_MX02 U9565 ( .S(n280), .A0(shiftedOData[286]), .A1(n4017), .Z(n590));
Q_FDP0UA U9566 ( .D(n589), .QTFCLK( ), .Q(shiftedOData[285]));
Q_MX02 U9567 ( .S(n280), .A0(shiftedOData[285]), .A1(n4016), .Z(n589));
Q_FDP0UA U9568 ( .D(n588), .QTFCLK( ), .Q(shiftedOData[284]));
Q_MX02 U9569 ( .S(n280), .A0(shiftedOData[284]), .A1(n4015), .Z(n588));
Q_FDP0UA U9570 ( .D(n587), .QTFCLK( ), .Q(shiftedOData[283]));
Q_MX02 U9571 ( .S(n280), .A0(shiftedOData[283]), .A1(n4014), .Z(n587));
Q_FDP0UA U9572 ( .D(n586), .QTFCLK( ), .Q(shiftedOData[282]));
Q_MX02 U9573 ( .S(n280), .A0(shiftedOData[282]), .A1(n4013), .Z(n586));
Q_FDP0UA U9574 ( .D(n585), .QTFCLK( ), .Q(shiftedOData[281]));
Q_MX02 U9575 ( .S(n280), .A0(shiftedOData[281]), .A1(n4012), .Z(n585));
Q_FDP0UA U9576 ( .D(n584), .QTFCLK( ), .Q(shiftedOData[280]));
Q_MX02 U9577 ( .S(n280), .A0(shiftedOData[280]), .A1(n4011), .Z(n584));
Q_FDP0UA U9578 ( .D(n583), .QTFCLK( ), .Q(shiftedOData[279]));
Q_MX02 U9579 ( .S(n280), .A0(shiftedOData[279]), .A1(n4010), .Z(n583));
Q_FDP0UA U9580 ( .D(n582), .QTFCLK( ), .Q(shiftedOData[278]));
Q_MX02 U9581 ( .S(n280), .A0(shiftedOData[278]), .A1(n4009), .Z(n582));
Q_FDP0UA U9582 ( .D(n581), .QTFCLK( ), .Q(shiftedOData[277]));
Q_MX02 U9583 ( .S(n280), .A0(shiftedOData[277]), .A1(n4008), .Z(n581));
Q_FDP0UA U9584 ( .D(n580), .QTFCLK( ), .Q(shiftedOData[276]));
Q_MX02 U9585 ( .S(n280), .A0(shiftedOData[276]), .A1(n4007), .Z(n580));
Q_FDP0UA U9586 ( .D(n579), .QTFCLK( ), .Q(shiftedOData[275]));
Q_MX02 U9587 ( .S(n280), .A0(shiftedOData[275]), .A1(n4006), .Z(n579));
Q_FDP0UA U9588 ( .D(n578), .QTFCLK( ), .Q(shiftedOData[274]));
Q_MX02 U9589 ( .S(n280), .A0(shiftedOData[274]), .A1(n4005), .Z(n578));
Q_FDP0UA U9590 ( .D(n577), .QTFCLK( ), .Q(shiftedOData[273]));
Q_MX02 U9591 ( .S(n280), .A0(shiftedOData[273]), .A1(n4004), .Z(n577));
Q_FDP0UA U9592 ( .D(n576), .QTFCLK( ), .Q(shiftedOData[272]));
Q_MX02 U9593 ( .S(n280), .A0(shiftedOData[272]), .A1(n4003), .Z(n576));
Q_FDP0UA U9594 ( .D(n575), .QTFCLK( ), .Q(shiftedOData[271]));
Q_MX02 U9595 ( .S(n280), .A0(shiftedOData[271]), .A1(n4002), .Z(n575));
Q_FDP0UA U9596 ( .D(n574), .QTFCLK( ), .Q(shiftedOData[270]));
Q_MX02 U9597 ( .S(n280), .A0(shiftedOData[270]), .A1(n4001), .Z(n574));
Q_FDP0UA U9598 ( .D(n573), .QTFCLK( ), .Q(shiftedOData[269]));
Q_MX02 U9599 ( .S(n280), .A0(shiftedOData[269]), .A1(n4000), .Z(n573));
Q_FDP0UA U9600 ( .D(n572), .QTFCLK( ), .Q(shiftedOData[268]));
Q_MX02 U9601 ( .S(n280), .A0(shiftedOData[268]), .A1(n3999), .Z(n572));
Q_FDP0UA U9602 ( .D(n571), .QTFCLK( ), .Q(shiftedOData[267]));
Q_MX02 U9603 ( .S(n280), .A0(shiftedOData[267]), .A1(n3998), .Z(n571));
Q_FDP0UA U9604 ( .D(n570), .QTFCLK( ), .Q(shiftedOData[266]));
Q_MX02 U9605 ( .S(n280), .A0(shiftedOData[266]), .A1(n3997), .Z(n570));
Q_FDP0UA U9606 ( .D(n569), .QTFCLK( ), .Q(shiftedOData[265]));
Q_MX02 U9607 ( .S(n280), .A0(shiftedOData[265]), .A1(n3996), .Z(n569));
Q_FDP0UA U9608 ( .D(n568), .QTFCLK( ), .Q(shiftedOData[264]));
Q_MX02 U9609 ( .S(n280), .A0(shiftedOData[264]), .A1(n3995), .Z(n568));
Q_FDP0UA U9610 ( .D(n567), .QTFCLK( ), .Q(shiftedOData[263]));
Q_MX02 U9611 ( .S(n280), .A0(shiftedOData[263]), .A1(n3994), .Z(n567));
Q_FDP0UA U9612 ( .D(n566), .QTFCLK( ), .Q(shiftedOData[262]));
Q_MX02 U9613 ( .S(n280), .A0(shiftedOData[262]), .A1(n3993), .Z(n566));
Q_FDP0UA U9614 ( .D(n565), .QTFCLK( ), .Q(shiftedOData[261]));
Q_MX02 U9615 ( .S(n280), .A0(shiftedOData[261]), .A1(n3992), .Z(n565));
Q_FDP0UA U9616 ( .D(n564), .QTFCLK( ), .Q(shiftedOData[260]));
Q_MX02 U9617 ( .S(n280), .A0(shiftedOData[260]), .A1(n3991), .Z(n564));
Q_FDP0UA U9618 ( .D(n563), .QTFCLK( ), .Q(shiftedOData[259]));
Q_MX02 U9619 ( .S(n280), .A0(shiftedOData[259]), .A1(n3990), .Z(n563));
Q_FDP0UA U9620 ( .D(n562), .QTFCLK( ), .Q(shiftedOData[258]));
Q_MX02 U9621 ( .S(n280), .A0(shiftedOData[258]), .A1(n3989), .Z(n562));
Q_FDP0UA U9622 ( .D(n561), .QTFCLK( ), .Q(shiftedOData[257]));
Q_MX02 U9623 ( .S(n280), .A0(shiftedOData[257]), .A1(n3988), .Z(n561));
Q_FDP0UA U9624 ( .D(n560), .QTFCLK( ), .Q(shiftedOData[256]));
Q_MX02 U9625 ( .S(n280), .A0(shiftedOData[256]), .A1(n3987), .Z(n560));
Q_FDP0UA U9626 ( .D(n559), .QTFCLK( ), .Q(shiftedOData[255]));
Q_MX02 U9627 ( .S(n280), .A0(shiftedOData[255]), .A1(n3986), .Z(n559));
Q_FDP0UA U9628 ( .D(n558), .QTFCLK( ), .Q(shiftedOData[254]));
Q_MX02 U9629 ( .S(n280), .A0(shiftedOData[254]), .A1(n3985), .Z(n558));
Q_FDP0UA U9630 ( .D(n557), .QTFCLK( ), .Q(shiftedOData[253]));
Q_MX02 U9631 ( .S(n280), .A0(shiftedOData[253]), .A1(n3984), .Z(n557));
Q_FDP0UA U9632 ( .D(n556), .QTFCLK( ), .Q(shiftedOData[252]));
Q_MX02 U9633 ( .S(n280), .A0(shiftedOData[252]), .A1(n3983), .Z(n556));
Q_FDP0UA U9634 ( .D(n555), .QTFCLK( ), .Q(shiftedOData[251]));
Q_MX02 U9635 ( .S(n280), .A0(shiftedOData[251]), .A1(n3982), .Z(n555));
Q_FDP0UA U9636 ( .D(n554), .QTFCLK( ), .Q(shiftedOData[250]));
Q_MX02 U9637 ( .S(n280), .A0(shiftedOData[250]), .A1(n3981), .Z(n554));
Q_FDP0UA U9638 ( .D(n553), .QTFCLK( ), .Q(shiftedOData[249]));
Q_MX02 U9639 ( .S(n280), .A0(shiftedOData[249]), .A1(n3980), .Z(n553));
Q_FDP0UA U9640 ( .D(n552), .QTFCLK( ), .Q(shiftedOData[248]));
Q_MX02 U9641 ( .S(n280), .A0(shiftedOData[248]), .A1(n3979), .Z(n552));
Q_FDP0UA U9642 ( .D(n551), .QTFCLK( ), .Q(shiftedOData[247]));
Q_MX02 U9643 ( .S(n280), .A0(shiftedOData[247]), .A1(n3978), .Z(n551));
Q_FDP0UA U9644 ( .D(n550), .QTFCLK( ), .Q(shiftedOData[246]));
Q_MX02 U9645 ( .S(n280), .A0(shiftedOData[246]), .A1(n3977), .Z(n550));
Q_FDP0UA U9646 ( .D(n549), .QTFCLK( ), .Q(shiftedOData[245]));
Q_MX02 U9647 ( .S(n280), .A0(shiftedOData[245]), .A1(n3976), .Z(n549));
Q_FDP0UA U9648 ( .D(n548), .QTFCLK( ), .Q(shiftedOData[244]));
Q_MX02 U9649 ( .S(n280), .A0(shiftedOData[244]), .A1(n3975), .Z(n548));
Q_FDP0UA U9650 ( .D(n547), .QTFCLK( ), .Q(shiftedOData[243]));
Q_MX02 U9651 ( .S(n280), .A0(shiftedOData[243]), .A1(n3974), .Z(n547));
Q_FDP0UA U9652 ( .D(n546), .QTFCLK( ), .Q(shiftedOData[242]));
Q_MX02 U9653 ( .S(n280), .A0(shiftedOData[242]), .A1(n3973), .Z(n546));
Q_FDP0UA U9654 ( .D(n545), .QTFCLK( ), .Q(shiftedOData[241]));
Q_MX02 U9655 ( .S(n280), .A0(shiftedOData[241]), .A1(n3972), .Z(n545));
Q_FDP0UA U9656 ( .D(n544), .QTFCLK( ), .Q(shiftedOData[240]));
Q_MX02 U9657 ( .S(n280), .A0(shiftedOData[240]), .A1(n3971), .Z(n544));
Q_FDP0UA U9658 ( .D(n543), .QTFCLK( ), .Q(shiftedOData[239]));
Q_MX02 U9659 ( .S(n280), .A0(shiftedOData[239]), .A1(n3970), .Z(n543));
Q_FDP0UA U9660 ( .D(n542), .QTFCLK( ), .Q(shiftedOData[238]));
Q_MX02 U9661 ( .S(n280), .A0(shiftedOData[238]), .A1(n3969), .Z(n542));
Q_FDP0UA U9662 ( .D(n541), .QTFCLK( ), .Q(shiftedOData[237]));
Q_MX02 U9663 ( .S(n280), .A0(shiftedOData[237]), .A1(n3968), .Z(n541));
Q_FDP0UA U9664 ( .D(n540), .QTFCLK( ), .Q(shiftedOData[236]));
Q_MX02 U9665 ( .S(n280), .A0(shiftedOData[236]), .A1(n3967), .Z(n540));
Q_FDP0UA U9666 ( .D(n539), .QTFCLK( ), .Q(shiftedOData[235]));
Q_MX02 U9667 ( .S(n280), .A0(shiftedOData[235]), .A1(n3966), .Z(n539));
Q_FDP0UA U9668 ( .D(n538), .QTFCLK( ), .Q(shiftedOData[234]));
Q_MX02 U9669 ( .S(n280), .A0(shiftedOData[234]), .A1(n3965), .Z(n538));
Q_FDP0UA U9670 ( .D(n537), .QTFCLK( ), .Q(shiftedOData[233]));
Q_MX02 U9671 ( .S(n280), .A0(shiftedOData[233]), .A1(n3964), .Z(n537));
Q_FDP0UA U9672 ( .D(n536), .QTFCLK( ), .Q(shiftedOData[232]));
Q_MX02 U9673 ( .S(n280), .A0(shiftedOData[232]), .A1(n3963), .Z(n536));
Q_FDP0UA U9674 ( .D(n535), .QTFCLK( ), .Q(shiftedOData[231]));
Q_MX02 U9675 ( .S(n280), .A0(shiftedOData[231]), .A1(n3962), .Z(n535));
Q_FDP0UA U9676 ( .D(n534), .QTFCLK( ), .Q(shiftedOData[230]));
Q_MX02 U9677 ( .S(n280), .A0(shiftedOData[230]), .A1(n3961), .Z(n534));
Q_FDP0UA U9678 ( .D(n533), .QTFCLK( ), .Q(shiftedOData[229]));
Q_MX02 U9679 ( .S(n280), .A0(shiftedOData[229]), .A1(n3960), .Z(n533));
Q_FDP0UA U9680 ( .D(n532), .QTFCLK( ), .Q(shiftedOData[228]));
Q_MX02 U9681 ( .S(n280), .A0(shiftedOData[228]), .A1(n3959), .Z(n532));
Q_FDP0UA U9682 ( .D(n531), .QTFCLK( ), .Q(shiftedOData[227]));
Q_MX02 U9683 ( .S(n280), .A0(shiftedOData[227]), .A1(n3958), .Z(n531));
Q_FDP0UA U9684 ( .D(n530), .QTFCLK( ), .Q(shiftedOData[226]));
Q_MX02 U9685 ( .S(n280), .A0(shiftedOData[226]), .A1(n3957), .Z(n530));
Q_FDP0UA U9686 ( .D(n529), .QTFCLK( ), .Q(shiftedOData[225]));
Q_MX02 U9687 ( .S(n280), .A0(shiftedOData[225]), .A1(n3956), .Z(n529));
Q_FDP0UA U9688 ( .D(n528), .QTFCLK( ), .Q(shiftedOData[224]));
Q_MX02 U9689 ( .S(n280), .A0(shiftedOData[224]), .A1(n3955), .Z(n528));
Q_FDP0UA U9690 ( .D(n527), .QTFCLK( ), .Q(shiftedOData[223]));
Q_MX02 U9691 ( .S(n280), .A0(shiftedOData[223]), .A1(n3954), .Z(n527));
Q_FDP0UA U9692 ( .D(n526), .QTFCLK( ), .Q(shiftedOData[222]));
Q_MX02 U9693 ( .S(n280), .A0(shiftedOData[222]), .A1(n3953), .Z(n526));
Q_FDP0UA U9694 ( .D(n525), .QTFCLK( ), .Q(shiftedOData[221]));
Q_MX02 U9695 ( .S(n280), .A0(shiftedOData[221]), .A1(n3952), .Z(n525));
Q_FDP0UA U9696 ( .D(n524), .QTFCLK( ), .Q(shiftedOData[220]));
Q_MX02 U9697 ( .S(n280), .A0(shiftedOData[220]), .A1(n3951), .Z(n524));
Q_FDP0UA U9698 ( .D(n523), .QTFCLK( ), .Q(shiftedOData[219]));
Q_MX02 U9699 ( .S(n280), .A0(shiftedOData[219]), .A1(n3950), .Z(n523));
Q_FDP0UA U9700 ( .D(n522), .QTFCLK( ), .Q(shiftedOData[218]));
Q_MX02 U9701 ( .S(n280), .A0(shiftedOData[218]), .A1(n3949), .Z(n522));
Q_FDP0UA U9702 ( .D(n521), .QTFCLK( ), .Q(shiftedOData[217]));
Q_MX02 U9703 ( .S(n280), .A0(shiftedOData[217]), .A1(n3948), .Z(n521));
Q_FDP0UA U9704 ( .D(n520), .QTFCLK( ), .Q(shiftedOData[216]));
Q_MX02 U9705 ( .S(n280), .A0(shiftedOData[216]), .A1(n3947), .Z(n520));
Q_FDP0UA U9706 ( .D(n519), .QTFCLK( ), .Q(shiftedOData[215]));
Q_MX02 U9707 ( .S(n280), .A0(shiftedOData[215]), .A1(n3946), .Z(n519));
Q_FDP0UA U9708 ( .D(n518), .QTFCLK( ), .Q(shiftedOData[214]));
Q_MX02 U9709 ( .S(n280), .A0(shiftedOData[214]), .A1(n3945), .Z(n518));
Q_FDP0UA U9710 ( .D(n517), .QTFCLK( ), .Q(shiftedOData[213]));
Q_MX02 U9711 ( .S(n280), .A0(shiftedOData[213]), .A1(n3944), .Z(n517));
Q_FDP0UA U9712 ( .D(n516), .QTFCLK( ), .Q(shiftedOData[212]));
Q_MX02 U9713 ( .S(n280), .A0(shiftedOData[212]), .A1(n3943), .Z(n516));
Q_FDP0UA U9714 ( .D(n515), .QTFCLK( ), .Q(shiftedOData[211]));
Q_MX02 U9715 ( .S(n280), .A0(shiftedOData[211]), .A1(n3942), .Z(n515));
Q_FDP0UA U9716 ( .D(n514), .QTFCLK( ), .Q(shiftedOData[210]));
Q_MX02 U9717 ( .S(n280), .A0(shiftedOData[210]), .A1(n3941), .Z(n514));
Q_FDP0UA U9718 ( .D(n513), .QTFCLK( ), .Q(shiftedOData[209]));
Q_MX02 U9719 ( .S(n280), .A0(shiftedOData[209]), .A1(n3940), .Z(n513));
Q_FDP0UA U9720 ( .D(n512), .QTFCLK( ), .Q(shiftedOData[208]));
Q_MX02 U9721 ( .S(n280), .A0(shiftedOData[208]), .A1(n3939), .Z(n512));
Q_FDP0UA U9722 ( .D(n511), .QTFCLK( ), .Q(shiftedOData[207]));
Q_MX02 U9723 ( .S(n280), .A0(shiftedOData[207]), .A1(n3938), .Z(n511));
Q_FDP0UA U9724 ( .D(n510), .QTFCLK( ), .Q(shiftedOData[206]));
Q_MX02 U9725 ( .S(n280), .A0(shiftedOData[206]), .A1(n3937), .Z(n510));
Q_FDP0UA U9726 ( .D(n509), .QTFCLK( ), .Q(shiftedOData[205]));
Q_MX02 U9727 ( .S(n280), .A0(shiftedOData[205]), .A1(n3936), .Z(n509));
Q_FDP0UA U9728 ( .D(n508), .QTFCLK( ), .Q(shiftedOData[204]));
Q_MX02 U9729 ( .S(n280), .A0(shiftedOData[204]), .A1(n3935), .Z(n508));
Q_FDP0UA U9730 ( .D(n507), .QTFCLK( ), .Q(shiftedOData[203]));
Q_MX02 U9731 ( .S(n280), .A0(shiftedOData[203]), .A1(n3934), .Z(n507));
Q_FDP0UA U9732 ( .D(n506), .QTFCLK( ), .Q(shiftedOData[202]));
Q_MX02 U9733 ( .S(n280), .A0(shiftedOData[202]), .A1(n3933), .Z(n506));
Q_FDP0UA U9734 ( .D(n505), .QTFCLK( ), .Q(shiftedOData[201]));
Q_MX02 U9735 ( .S(n280), .A0(shiftedOData[201]), .A1(n3932), .Z(n505));
Q_FDP0UA U9736 ( .D(n504), .QTFCLK( ), .Q(shiftedOData[200]));
Q_MX02 U9737 ( .S(n280), .A0(shiftedOData[200]), .A1(n3931), .Z(n504));
Q_FDP0UA U9738 ( .D(n503), .QTFCLK( ), .Q(shiftedOData[199]));
Q_MX02 U9739 ( .S(n280), .A0(shiftedOData[199]), .A1(n3930), .Z(n503));
Q_FDP0UA U9740 ( .D(n502), .QTFCLK( ), .Q(shiftedOData[198]));
Q_MX02 U9741 ( .S(n280), .A0(shiftedOData[198]), .A1(n3929), .Z(n502));
Q_FDP0UA U9742 ( .D(n501), .QTFCLK( ), .Q(shiftedOData[197]));
Q_MX02 U9743 ( .S(n280), .A0(shiftedOData[197]), .A1(n3928), .Z(n501));
Q_FDP0UA U9744 ( .D(n500), .QTFCLK( ), .Q(shiftedOData[196]));
Q_MX02 U9745 ( .S(n280), .A0(shiftedOData[196]), .A1(n3927), .Z(n500));
Q_FDP0UA U9746 ( .D(n499), .QTFCLK( ), .Q(shiftedOData[195]));
Q_MX02 U9747 ( .S(n280), .A0(shiftedOData[195]), .A1(n3926), .Z(n499));
Q_FDP0UA U9748 ( .D(n498), .QTFCLK( ), .Q(shiftedOData[194]));
Q_MX02 U9749 ( .S(n280), .A0(shiftedOData[194]), .A1(n3925), .Z(n498));
Q_FDP0UA U9750 ( .D(n497), .QTFCLK( ), .Q(shiftedOData[193]));
Q_MX02 U9751 ( .S(n280), .A0(shiftedOData[193]), .A1(n3924), .Z(n497));
Q_FDP0UA U9752 ( .D(n496), .QTFCLK( ), .Q(shiftedOData[192]));
Q_MX02 U9753 ( .S(n280), .A0(shiftedOData[192]), .A1(n3923), .Z(n496));
Q_FDP0UA U9754 ( .D(n495), .QTFCLK( ), .Q(shiftedOData[191]));
Q_MX02 U9755 ( .S(n280), .A0(shiftedOData[191]), .A1(n3922), .Z(n495));
Q_FDP0UA U9756 ( .D(n494), .QTFCLK( ), .Q(shiftedOData[190]));
Q_MX02 U9757 ( .S(n280), .A0(shiftedOData[190]), .A1(n3921), .Z(n494));
Q_FDP0UA U9758 ( .D(n493), .QTFCLK( ), .Q(shiftedOData[189]));
Q_MX02 U9759 ( .S(n280), .A0(shiftedOData[189]), .A1(n3920), .Z(n493));
Q_FDP0UA U9760 ( .D(n492), .QTFCLK( ), .Q(shiftedOData[188]));
Q_MX02 U9761 ( .S(n280), .A0(shiftedOData[188]), .A1(n3919), .Z(n492));
Q_FDP0UA U9762 ( .D(n491), .QTFCLK( ), .Q(shiftedOData[187]));
Q_MX02 U9763 ( .S(n280), .A0(shiftedOData[187]), .A1(n3918), .Z(n491));
Q_FDP0UA U9764 ( .D(n490), .QTFCLK( ), .Q(shiftedOData[186]));
Q_MX02 U9765 ( .S(n280), .A0(shiftedOData[186]), .A1(n3917), .Z(n490));
Q_FDP0UA U9766 ( .D(n489), .QTFCLK( ), .Q(shiftedOData[185]));
Q_MX02 U9767 ( .S(n280), .A0(shiftedOData[185]), .A1(n3916), .Z(n489));
Q_FDP0UA U9768 ( .D(n488), .QTFCLK( ), .Q(shiftedOData[184]));
Q_MX02 U9769 ( .S(n280), .A0(shiftedOData[184]), .A1(n3915), .Z(n488));
Q_FDP0UA U9770 ( .D(n487), .QTFCLK( ), .Q(shiftedOData[183]));
Q_MX02 U9771 ( .S(n280), .A0(shiftedOData[183]), .A1(n3914), .Z(n487));
Q_FDP0UA U9772 ( .D(n486), .QTFCLK( ), .Q(shiftedOData[182]));
Q_MX02 U9773 ( .S(n280), .A0(shiftedOData[182]), .A1(n3913), .Z(n486));
Q_FDP0UA U9774 ( .D(n485), .QTFCLK( ), .Q(shiftedOData[181]));
Q_MX02 U9775 ( .S(n280), .A0(shiftedOData[181]), .A1(n3912), .Z(n485));
Q_FDP0UA U9776 ( .D(n484), .QTFCLK( ), .Q(shiftedOData[180]));
Q_MX02 U9777 ( .S(n280), .A0(shiftedOData[180]), .A1(n3911), .Z(n484));
Q_FDP0UA U9778 ( .D(n483), .QTFCLK( ), .Q(shiftedOData[179]));
Q_MX02 U9779 ( .S(n280), .A0(shiftedOData[179]), .A1(n3910), .Z(n483));
Q_FDP0UA U9780 ( .D(n482), .QTFCLK( ), .Q(shiftedOData[178]));
Q_MX02 U9781 ( .S(n280), .A0(shiftedOData[178]), .A1(n3909), .Z(n482));
Q_FDP0UA U9782 ( .D(n481), .QTFCLK( ), .Q(shiftedOData[177]));
Q_MX02 U9783 ( .S(n280), .A0(shiftedOData[177]), .A1(n3908), .Z(n481));
Q_FDP0UA U9784 ( .D(n480), .QTFCLK( ), .Q(shiftedOData[176]));
Q_MX02 U9785 ( .S(n280), .A0(shiftedOData[176]), .A1(n3907), .Z(n480));
Q_FDP0UA U9786 ( .D(n479), .QTFCLK( ), .Q(shiftedOData[175]));
Q_MX02 U9787 ( .S(n280), .A0(shiftedOData[175]), .A1(n3906), .Z(n479));
Q_FDP0UA U9788 ( .D(n478), .QTFCLK( ), .Q(shiftedOData[174]));
Q_MX02 U9789 ( .S(n280), .A0(shiftedOData[174]), .A1(n3905), .Z(n478));
Q_FDP0UA U9790 ( .D(n477), .QTFCLK( ), .Q(shiftedOData[173]));
Q_MX02 U9791 ( .S(n280), .A0(shiftedOData[173]), .A1(n3904), .Z(n477));
Q_FDP0UA U9792 ( .D(n476), .QTFCLK( ), .Q(shiftedOData[172]));
Q_MX02 U9793 ( .S(n280), .A0(shiftedOData[172]), .A1(n3903), .Z(n476));
Q_FDP0UA U9794 ( .D(n475), .QTFCLK( ), .Q(shiftedOData[171]));
Q_MX02 U9795 ( .S(n280), .A0(shiftedOData[171]), .A1(n3902), .Z(n475));
Q_FDP0UA U9796 ( .D(n474), .QTFCLK( ), .Q(shiftedOData[170]));
Q_MX02 U9797 ( .S(n280), .A0(shiftedOData[170]), .A1(n3901), .Z(n474));
Q_FDP0UA U9798 ( .D(n473), .QTFCLK( ), .Q(shiftedOData[169]));
Q_MX02 U9799 ( .S(n280), .A0(shiftedOData[169]), .A1(n3900), .Z(n473));
Q_FDP0UA U9800 ( .D(n472), .QTFCLK( ), .Q(shiftedOData[168]));
Q_MX02 U9801 ( .S(n280), .A0(shiftedOData[168]), .A1(n3899), .Z(n472));
Q_FDP0UA U9802 ( .D(n471), .QTFCLK( ), .Q(shiftedOData[167]));
Q_MX02 U9803 ( .S(n280), .A0(shiftedOData[167]), .A1(n3898), .Z(n471));
Q_FDP0UA U9804 ( .D(n470), .QTFCLK( ), .Q(shiftedOData[166]));
Q_MX02 U9805 ( .S(n280), .A0(shiftedOData[166]), .A1(n3897), .Z(n470));
Q_FDP0UA U9806 ( .D(n469), .QTFCLK( ), .Q(shiftedOData[165]));
Q_MX02 U9807 ( .S(n280), .A0(shiftedOData[165]), .A1(n3896), .Z(n469));
Q_FDP0UA U9808 ( .D(n468), .QTFCLK( ), .Q(shiftedOData[164]));
Q_MX02 U9809 ( .S(n280), .A0(shiftedOData[164]), .A1(n3895), .Z(n468));
Q_FDP0UA U9810 ( .D(n467), .QTFCLK( ), .Q(shiftedOData[163]));
Q_MX02 U9811 ( .S(n280), .A0(shiftedOData[163]), .A1(n3894), .Z(n467));
Q_FDP0UA U9812 ( .D(n466), .QTFCLK( ), .Q(shiftedOData[162]));
Q_MX02 U9813 ( .S(n280), .A0(shiftedOData[162]), .A1(n3893), .Z(n466));
Q_FDP0UA U9814 ( .D(n465), .QTFCLK( ), .Q(shiftedOData[161]));
Q_MX02 U9815 ( .S(n280), .A0(shiftedOData[161]), .A1(n3892), .Z(n465));
Q_FDP0UA U9816 ( .D(n464), .QTFCLK( ), .Q(shiftedOData[160]));
Q_MX02 U9817 ( .S(n280), .A0(shiftedOData[160]), .A1(n3891), .Z(n464));
Q_FDP0UA U9818 ( .D(n463), .QTFCLK( ), .Q(shiftedOData[159]));
Q_MX02 U9819 ( .S(n280), .A0(shiftedOData[159]), .A1(n3890), .Z(n463));
Q_FDP0UA U9820 ( .D(n462), .QTFCLK( ), .Q(shiftedOData[158]));
Q_MX02 U9821 ( .S(n280), .A0(shiftedOData[158]), .A1(n3889), .Z(n462));
Q_FDP0UA U9822 ( .D(n461), .QTFCLK( ), .Q(shiftedOData[157]));
Q_MX02 U9823 ( .S(n280), .A0(shiftedOData[157]), .A1(n3888), .Z(n461));
Q_FDP0UA U9824 ( .D(n460), .QTFCLK( ), .Q(shiftedOData[156]));
Q_MX02 U9825 ( .S(n280), .A0(shiftedOData[156]), .A1(n3887), .Z(n460));
Q_FDP0UA U9826 ( .D(n459), .QTFCLK( ), .Q(shiftedOData[155]));
Q_MX02 U9827 ( .S(n280), .A0(shiftedOData[155]), .A1(n3886), .Z(n459));
Q_FDP0UA U9828 ( .D(n458), .QTFCLK( ), .Q(shiftedOData[154]));
Q_MX02 U9829 ( .S(n280), .A0(shiftedOData[154]), .A1(n3885), .Z(n458));
Q_FDP0UA U9830 ( .D(n457), .QTFCLK( ), .Q(shiftedOData[153]));
Q_MX02 U9831 ( .S(n280), .A0(shiftedOData[153]), .A1(n3884), .Z(n457));
Q_FDP0UA U9832 ( .D(n456), .QTFCLK( ), .Q(shiftedOData[152]));
Q_MX02 U9833 ( .S(n280), .A0(shiftedOData[152]), .A1(n3883), .Z(n456));
Q_FDP0UA U9834 ( .D(n455), .QTFCLK( ), .Q(shiftedOData[151]));
Q_MX02 U9835 ( .S(n280), .A0(shiftedOData[151]), .A1(n3882), .Z(n455));
Q_FDP0UA U9836 ( .D(n454), .QTFCLK( ), .Q(shiftedOData[150]));
Q_MX02 U9837 ( .S(n280), .A0(shiftedOData[150]), .A1(n3881), .Z(n454));
Q_FDP0UA U9838 ( .D(n453), .QTFCLK( ), .Q(shiftedOData[149]));
Q_MX02 U9839 ( .S(n280), .A0(shiftedOData[149]), .A1(n3880), .Z(n453));
Q_FDP0UA U9840 ( .D(n452), .QTFCLK( ), .Q(shiftedOData[148]));
Q_MX02 U9841 ( .S(n280), .A0(shiftedOData[148]), .A1(n3879), .Z(n452));
Q_FDP0UA U9842 ( .D(n451), .QTFCLK( ), .Q(shiftedOData[147]));
Q_MX02 U9843 ( .S(n280), .A0(shiftedOData[147]), .A1(n3878), .Z(n451));
Q_FDP0UA U9844 ( .D(n450), .QTFCLK( ), .Q(shiftedOData[146]));
Q_MX02 U9845 ( .S(n280), .A0(shiftedOData[146]), .A1(n3877), .Z(n450));
Q_FDP0UA U9846 ( .D(n449), .QTFCLK( ), .Q(shiftedOData[145]));
Q_MX02 U9847 ( .S(n280), .A0(shiftedOData[145]), .A1(n3876), .Z(n449));
Q_FDP0UA U9848 ( .D(n448), .QTFCLK( ), .Q(shiftedOData[144]));
Q_MX02 U9849 ( .S(n280), .A0(shiftedOData[144]), .A1(n3875), .Z(n448));
Q_FDP0UA U9850 ( .D(n447), .QTFCLK( ), .Q(shiftedOData[143]));
Q_MX02 U9851 ( .S(n280), .A0(shiftedOData[143]), .A1(n3874), .Z(n447));
Q_FDP0UA U9852 ( .D(n446), .QTFCLK( ), .Q(shiftedOData[142]));
Q_MX02 U9853 ( .S(n280), .A0(shiftedOData[142]), .A1(n3873), .Z(n446));
Q_FDP0UA U9854 ( .D(n445), .QTFCLK( ), .Q(shiftedOData[141]));
Q_MX02 U9855 ( .S(n280), .A0(shiftedOData[141]), .A1(n3872), .Z(n445));
Q_FDP0UA U9856 ( .D(n444), .QTFCLK( ), .Q(shiftedOData[140]));
Q_MX02 U9857 ( .S(n280), .A0(shiftedOData[140]), .A1(n3871), .Z(n444));
Q_FDP0UA U9858 ( .D(n443), .QTFCLK( ), .Q(shiftedOData[139]));
Q_MX02 U9859 ( .S(n280), .A0(shiftedOData[139]), .A1(n3870), .Z(n443));
Q_FDP0UA U9860 ( .D(n442), .QTFCLK( ), .Q(shiftedOData[138]));
Q_MX02 U9861 ( .S(n280), .A0(shiftedOData[138]), .A1(n3869), .Z(n442));
Q_FDP0UA U9862 ( .D(n441), .QTFCLK( ), .Q(shiftedOData[137]));
Q_MX02 U9863 ( .S(n280), .A0(shiftedOData[137]), .A1(n3868), .Z(n441));
Q_FDP0UA U9864 ( .D(n440), .QTFCLK( ), .Q(shiftedOData[136]));
Q_MX02 U9865 ( .S(n280), .A0(shiftedOData[136]), .A1(n3867), .Z(n440));
Q_FDP0UA U9866 ( .D(n439), .QTFCLK( ), .Q(shiftedOData[135]));
Q_MX02 U9867 ( .S(n280), .A0(shiftedOData[135]), .A1(n3866), .Z(n439));
Q_FDP0UA U9868 ( .D(n438), .QTFCLK( ), .Q(shiftedOData[134]));
Q_MX02 U9869 ( .S(n280), .A0(shiftedOData[134]), .A1(n3865), .Z(n438));
Q_FDP0UA U9870 ( .D(n437), .QTFCLK( ), .Q(shiftedOData[133]));
Q_MX02 U9871 ( .S(n280), .A0(shiftedOData[133]), .A1(n3864), .Z(n437));
Q_FDP0UA U9872 ( .D(n436), .QTFCLK( ), .Q(shiftedOData[132]));
Q_MX02 U9873 ( .S(n280), .A0(shiftedOData[132]), .A1(n3863), .Z(n436));
Q_FDP0UA U9874 ( .D(n435), .QTFCLK( ), .Q(shiftedOData[131]));
Q_MX02 U9875 ( .S(n280), .A0(shiftedOData[131]), .A1(n3862), .Z(n435));
Q_FDP0UA U9876 ( .D(n434), .QTFCLK( ), .Q(shiftedOData[130]));
Q_MX02 U9877 ( .S(n280), .A0(shiftedOData[130]), .A1(n3861), .Z(n434));
Q_FDP0UA U9878 ( .D(n433), .QTFCLK( ), .Q(shiftedOData[129]));
Q_MX02 U9879 ( .S(n280), .A0(shiftedOData[129]), .A1(n3860), .Z(n433));
Q_FDP0UA U9880 ( .D(n432), .QTFCLK( ), .Q(shiftedOData[128]));
Q_MX02 U9881 ( .S(n280), .A0(shiftedOData[128]), .A1(n3859), .Z(n432));
Q_FDP0UA U9882 ( .D(n431), .QTFCLK( ), .Q(shiftedOData[127]));
Q_MX02 U9883 ( .S(n280), .A0(shiftedOData[127]), .A1(n3857), .Z(n431));
Q_FDP0UA U9884 ( .D(n430), .QTFCLK( ), .Q(shiftedOData[126]));
Q_MX02 U9885 ( .S(n280), .A0(shiftedOData[126]), .A1(n3856), .Z(n430));
Q_FDP0UA U9886 ( .D(n429), .QTFCLK( ), .Q(shiftedOData[125]));
Q_MX02 U9887 ( .S(n280), .A0(shiftedOData[125]), .A1(n3855), .Z(n429));
Q_FDP0UA U9888 ( .D(n428), .QTFCLK( ), .Q(shiftedOData[124]));
Q_MX02 U9889 ( .S(n280), .A0(shiftedOData[124]), .A1(n3854), .Z(n428));
Q_FDP0UA U9890 ( .D(n427), .QTFCLK( ), .Q(shiftedOData[123]));
Q_MX02 U9891 ( .S(n280), .A0(shiftedOData[123]), .A1(n3853), .Z(n427));
Q_FDP0UA U9892 ( .D(n426), .QTFCLK( ), .Q(shiftedOData[122]));
Q_MX02 U9893 ( .S(n280), .A0(shiftedOData[122]), .A1(n3852), .Z(n426));
Q_FDP0UA U9894 ( .D(n425), .QTFCLK( ), .Q(shiftedOData[121]));
Q_MX02 U9895 ( .S(n280), .A0(shiftedOData[121]), .A1(n3851), .Z(n425));
Q_FDP0UA U9896 ( .D(n424), .QTFCLK( ), .Q(shiftedOData[120]));
Q_MX02 U9897 ( .S(n280), .A0(shiftedOData[120]), .A1(n3850), .Z(n424));
Q_FDP0UA U9898 ( .D(n423), .QTFCLK( ), .Q(shiftedOData[119]));
Q_MX02 U9899 ( .S(n280), .A0(shiftedOData[119]), .A1(n3849), .Z(n423));
Q_FDP0UA U9900 ( .D(n422), .QTFCLK( ), .Q(shiftedOData[118]));
Q_MX02 U9901 ( .S(n280), .A0(shiftedOData[118]), .A1(n3848), .Z(n422));
Q_FDP0UA U9902 ( .D(n421), .QTFCLK( ), .Q(shiftedOData[117]));
Q_MX02 U9903 ( .S(n280), .A0(shiftedOData[117]), .A1(n3847), .Z(n421));
Q_FDP0UA U9904 ( .D(n420), .QTFCLK( ), .Q(shiftedOData[116]));
Q_MX02 U9905 ( .S(n280), .A0(shiftedOData[116]), .A1(n3846), .Z(n420));
Q_FDP0UA U9906 ( .D(n419), .QTFCLK( ), .Q(shiftedOData[115]));
Q_MX02 U9907 ( .S(n280), .A0(shiftedOData[115]), .A1(n3845), .Z(n419));
Q_FDP0UA U9908 ( .D(n418), .QTFCLK( ), .Q(shiftedOData[114]));
Q_MX02 U9909 ( .S(n280), .A0(shiftedOData[114]), .A1(n3844), .Z(n418));
Q_FDP0UA U9910 ( .D(n417), .QTFCLK( ), .Q(shiftedOData[113]));
Q_MX02 U9911 ( .S(n280), .A0(shiftedOData[113]), .A1(n3843), .Z(n417));
Q_FDP0UA U9912 ( .D(n416), .QTFCLK( ), .Q(shiftedOData[112]));
Q_MX02 U9913 ( .S(n280), .A0(shiftedOData[112]), .A1(n3842), .Z(n416));
Q_FDP0UA U9914 ( .D(n415), .QTFCLK( ), .Q(shiftedOData[111]));
Q_MX02 U9915 ( .S(n280), .A0(shiftedOData[111]), .A1(n3841), .Z(n415));
Q_FDP0UA U9916 ( .D(n414), .QTFCLK( ), .Q(shiftedOData[110]));
Q_MX02 U9917 ( .S(n280), .A0(shiftedOData[110]), .A1(n3840), .Z(n414));
Q_FDP0UA U9918 ( .D(n413), .QTFCLK( ), .Q(shiftedOData[109]));
Q_MX02 U9919 ( .S(n280), .A0(shiftedOData[109]), .A1(n3839), .Z(n413));
Q_FDP0UA U9920 ( .D(n412), .QTFCLK( ), .Q(shiftedOData[108]));
Q_MX02 U9921 ( .S(n280), .A0(shiftedOData[108]), .A1(n3838), .Z(n412));
Q_FDP0UA U9922 ( .D(n411), .QTFCLK( ), .Q(shiftedOData[107]));
Q_MX02 U9923 ( .S(n280), .A0(shiftedOData[107]), .A1(n3837), .Z(n411));
Q_FDP0UA U9924 ( .D(n410), .QTFCLK( ), .Q(shiftedOData[106]));
Q_MX02 U9925 ( .S(n280), .A0(shiftedOData[106]), .A1(n3836), .Z(n410));
Q_FDP0UA U9926 ( .D(n409), .QTFCLK( ), .Q(shiftedOData[105]));
Q_MX02 U9927 ( .S(n280), .A0(shiftedOData[105]), .A1(n3835), .Z(n409));
Q_FDP0UA U9928 ( .D(n408), .QTFCLK( ), .Q(shiftedOData[104]));
Q_MX02 U9929 ( .S(n280), .A0(shiftedOData[104]), .A1(n3834), .Z(n408));
Q_FDP0UA U9930 ( .D(n407), .QTFCLK( ), .Q(shiftedOData[103]));
Q_MX02 U9931 ( .S(n280), .A0(shiftedOData[103]), .A1(n3833), .Z(n407));
Q_FDP0UA U9932 ( .D(n406), .QTFCLK( ), .Q(shiftedOData[102]));
Q_MX02 U9933 ( .S(n280), .A0(shiftedOData[102]), .A1(n3832), .Z(n406));
Q_FDP0UA U9934 ( .D(n405), .QTFCLK( ), .Q(shiftedOData[101]));
Q_MX02 U9935 ( .S(n280), .A0(shiftedOData[101]), .A1(n3831), .Z(n405));
Q_FDP0UA U9936 ( .D(n404), .QTFCLK( ), .Q(shiftedOData[100]));
Q_MX02 U9937 ( .S(n280), .A0(shiftedOData[100]), .A1(n3830), .Z(n404));
Q_FDP0UA U9938 ( .D(n403), .QTFCLK( ), .Q(shiftedOData[99]));
Q_MX02 U9939 ( .S(n280), .A0(shiftedOData[99]), .A1(n3829), .Z(n403));
Q_FDP0UA U9940 ( .D(n402), .QTFCLK( ), .Q(shiftedOData[98]));
Q_MX02 U9941 ( .S(n280), .A0(shiftedOData[98]), .A1(n3828), .Z(n402));
Q_FDP0UA U9942 ( .D(n401), .QTFCLK( ), .Q(shiftedOData[97]));
Q_MX02 U9943 ( .S(n280), .A0(shiftedOData[97]), .A1(n3827), .Z(n401));
Q_FDP0UA U9944 ( .D(n400), .QTFCLK( ), .Q(shiftedOData[96]));
Q_MX02 U9945 ( .S(n280), .A0(shiftedOData[96]), .A1(n3826), .Z(n400));
Q_FDP0UA U9946 ( .D(n399), .QTFCLK( ), .Q(shiftedOData[95]));
Q_MX02 U9947 ( .S(n280), .A0(shiftedOData[95]), .A1(n3825), .Z(n399));
Q_FDP0UA U9948 ( .D(n398), .QTFCLK( ), .Q(shiftedOData[94]));
Q_MX02 U9949 ( .S(n280), .A0(shiftedOData[94]), .A1(n3824), .Z(n398));
Q_FDP0UA U9950 ( .D(n397), .QTFCLK( ), .Q(shiftedOData[93]));
Q_MX02 U9951 ( .S(n280), .A0(shiftedOData[93]), .A1(n3823), .Z(n397));
Q_FDP0UA U9952 ( .D(n396), .QTFCLK( ), .Q(shiftedOData[92]));
Q_MX02 U9953 ( .S(n280), .A0(shiftedOData[92]), .A1(n3822), .Z(n396));
Q_FDP0UA U9954 ( .D(n395), .QTFCLK( ), .Q(shiftedOData[91]));
Q_MX02 U9955 ( .S(n280), .A0(shiftedOData[91]), .A1(n3821), .Z(n395));
Q_FDP0UA U9956 ( .D(n394), .QTFCLK( ), .Q(shiftedOData[90]));
Q_MX02 U9957 ( .S(n280), .A0(shiftedOData[90]), .A1(n3820), .Z(n394));
Q_FDP0UA U9958 ( .D(n393), .QTFCLK( ), .Q(shiftedOData[89]));
Q_MX02 U9959 ( .S(n280), .A0(shiftedOData[89]), .A1(n3819), .Z(n393));
Q_FDP0UA U9960 ( .D(n392), .QTFCLK( ), .Q(shiftedOData[88]));
Q_MX02 U9961 ( .S(n280), .A0(shiftedOData[88]), .A1(n3818), .Z(n392));
Q_FDP0UA U9962 ( .D(n391), .QTFCLK( ), .Q(shiftedOData[87]));
Q_MX02 U9963 ( .S(n280), .A0(shiftedOData[87]), .A1(n3817), .Z(n391));
Q_FDP0UA U9964 ( .D(n390), .QTFCLK( ), .Q(shiftedOData[86]));
Q_MX02 U9965 ( .S(n280), .A0(shiftedOData[86]), .A1(n3816), .Z(n390));
Q_FDP0UA U9966 ( .D(n389), .QTFCLK( ), .Q(shiftedOData[85]));
Q_MX02 U9967 ( .S(n280), .A0(shiftedOData[85]), .A1(n3815), .Z(n389));
Q_FDP0UA U9968 ( .D(n388), .QTFCLK( ), .Q(shiftedOData[84]));
Q_MX02 U9969 ( .S(n280), .A0(shiftedOData[84]), .A1(n3814), .Z(n388));
Q_FDP0UA U9970 ( .D(n387), .QTFCLK( ), .Q(shiftedOData[83]));
Q_MX02 U9971 ( .S(n280), .A0(shiftedOData[83]), .A1(n3813), .Z(n387));
Q_FDP0UA U9972 ( .D(n386), .QTFCLK( ), .Q(shiftedOData[82]));
Q_MX02 U9973 ( .S(n280), .A0(shiftedOData[82]), .A1(n3812), .Z(n386));
Q_FDP0UA U9974 ( .D(n385), .QTFCLK( ), .Q(shiftedOData[81]));
Q_MX02 U9975 ( .S(n280), .A0(shiftedOData[81]), .A1(n3811), .Z(n385));
Q_FDP0UA U9976 ( .D(n384), .QTFCLK( ), .Q(shiftedOData[80]));
Q_MX02 U9977 ( .S(n280), .A0(shiftedOData[80]), .A1(n3810), .Z(n384));
Q_FDP0UA U9978 ( .D(n383), .QTFCLK( ), .Q(shiftedOData[79]));
Q_MX02 U9979 ( .S(n280), .A0(shiftedOData[79]), .A1(n3809), .Z(n383));
Q_FDP0UA U9980 ( .D(n382), .QTFCLK( ), .Q(shiftedOData[78]));
Q_MX02 U9981 ( .S(n280), .A0(shiftedOData[78]), .A1(n3808), .Z(n382));
Q_FDP0UA U9982 ( .D(n381), .QTFCLK( ), .Q(shiftedOData[77]));
Q_MX02 U9983 ( .S(n280), .A0(shiftedOData[77]), .A1(n3807), .Z(n381));
Q_FDP0UA U9984 ( .D(n380), .QTFCLK( ), .Q(shiftedOData[76]));
Q_MX02 U9985 ( .S(n280), .A0(shiftedOData[76]), .A1(n3806), .Z(n380));
Q_FDP0UA U9986 ( .D(n379), .QTFCLK( ), .Q(shiftedOData[75]));
Q_MX02 U9987 ( .S(n280), .A0(shiftedOData[75]), .A1(n3805), .Z(n379));
Q_FDP0UA U9988 ( .D(n378), .QTFCLK( ), .Q(shiftedOData[74]));
Q_MX02 U9989 ( .S(n280), .A0(shiftedOData[74]), .A1(n3804), .Z(n378));
Q_FDP0UA U9990 ( .D(n377), .QTFCLK( ), .Q(shiftedOData[73]));
Q_MX02 U9991 ( .S(n280), .A0(shiftedOData[73]), .A1(n3803), .Z(n377));
Q_FDP0UA U9992 ( .D(n376), .QTFCLK( ), .Q(shiftedOData[72]));
Q_MX02 U9993 ( .S(n280), .A0(shiftedOData[72]), .A1(n3802), .Z(n376));
Q_FDP0UA U9994 ( .D(n375), .QTFCLK( ), .Q(shiftedOData[71]));
Q_MX02 U9995 ( .S(n280), .A0(shiftedOData[71]), .A1(n3801), .Z(n375));
Q_FDP0UA U9996 ( .D(n374), .QTFCLK( ), .Q(shiftedOData[70]));
Q_MX02 U9997 ( .S(n280), .A0(shiftedOData[70]), .A1(n3800), .Z(n374));
Q_FDP0UA U9998 ( .D(n373), .QTFCLK( ), .Q(shiftedOData[69]));
Q_MX02 U9999 ( .S(n280), .A0(shiftedOData[69]), .A1(n3799), .Z(n373));
Q_FDP0UA U10000 ( .D(n372), .QTFCLK( ), .Q(shiftedOData[68]));
Q_MX02 U10001 ( .S(n280), .A0(shiftedOData[68]), .A1(n3798), .Z(n372));
Q_FDP0UA U10002 ( .D(n371), .QTFCLK( ), .Q(shiftedOData[67]));
Q_MX02 U10003 ( .S(n280), .A0(shiftedOData[67]), .A1(n3797), .Z(n371));
Q_FDP0UA U10004 ( .D(n370), .QTFCLK( ), .Q(shiftedOData[66]));
Q_MX02 U10005 ( .S(n280), .A0(shiftedOData[66]), .A1(n3796), .Z(n370));
Q_FDP0UA U10006 ( .D(n369), .QTFCLK( ), .Q(shiftedOData[65]));
Q_MX02 U10007 ( .S(n280), .A0(shiftedOData[65]), .A1(n3795), .Z(n369));
Q_FDP0UA U10008 ( .D(n368), .QTFCLK( ), .Q(shiftedOData[64]));
Q_MX02 U10009 ( .S(n280), .A0(shiftedOData[64]), .A1(n3794), .Z(n368));
Q_FDP0UA U10010 ( .D(n367), .QTFCLK( ), .Q(shiftedOData[63]));
Q_MX02 U10011 ( .S(n280), .A0(shiftedOData[63]), .A1(n3793), .Z(n367));
Q_FDP0UA U10012 ( .D(n366), .QTFCLK( ), .Q(shiftedOData[62]));
Q_MX02 U10013 ( .S(n280), .A0(shiftedOData[62]), .A1(n3792), .Z(n366));
Q_FDP0UA U10014 ( .D(n365), .QTFCLK( ), .Q(shiftedOData[61]));
Q_MX02 U10015 ( .S(n280), .A0(shiftedOData[61]), .A1(n3791), .Z(n365));
Q_FDP0UA U10016 ( .D(n364), .QTFCLK( ), .Q(shiftedOData[60]));
Q_MX02 U10017 ( .S(n280), .A0(shiftedOData[60]), .A1(n3790), .Z(n364));
Q_FDP0UA U10018 ( .D(n363), .QTFCLK( ), .Q(shiftedOData[59]));
Q_MX02 U10019 ( .S(n280), .A0(shiftedOData[59]), .A1(n3789), .Z(n363));
Q_FDP0UA U10020 ( .D(n362), .QTFCLK( ), .Q(shiftedOData[58]));
Q_MX02 U10021 ( .S(n280), .A0(shiftedOData[58]), .A1(n3788), .Z(n362));
Q_FDP0UA U10022 ( .D(n361), .QTFCLK( ), .Q(shiftedOData[57]));
Q_MX02 U10023 ( .S(n280), .A0(shiftedOData[57]), .A1(n3787), .Z(n361));
Q_FDP0UA U10024 ( .D(n360), .QTFCLK( ), .Q(shiftedOData[56]));
Q_MX02 U10025 ( .S(n280), .A0(shiftedOData[56]), .A1(n3786), .Z(n360));
Q_FDP0UA U10026 ( .D(n359), .QTFCLK( ), .Q(shiftedOData[55]));
Q_MX02 U10027 ( .S(n280), .A0(shiftedOData[55]), .A1(n3785), .Z(n359));
Q_FDP0UA U10028 ( .D(n358), .QTFCLK( ), .Q(shiftedOData[54]));
Q_MX02 U10029 ( .S(n280), .A0(shiftedOData[54]), .A1(n3784), .Z(n358));
Q_FDP0UA U10030 ( .D(n357), .QTFCLK( ), .Q(shiftedOData[53]));
Q_MX02 U10031 ( .S(n280), .A0(shiftedOData[53]), .A1(n3783), .Z(n357));
Q_FDP0UA U10032 ( .D(n356), .QTFCLK( ), .Q(shiftedOData[52]));
Q_MX02 U10033 ( .S(n280), .A0(shiftedOData[52]), .A1(n3782), .Z(n356));
Q_FDP0UA U10034 ( .D(n355), .QTFCLK( ), .Q(shiftedOData[51]));
Q_MX02 U10035 ( .S(n280), .A0(shiftedOData[51]), .A1(n3781), .Z(n355));
Q_FDP0UA U10036 ( .D(n354), .QTFCLK( ), .Q(shiftedOData[50]));
Q_MX02 U10037 ( .S(n280), .A0(shiftedOData[50]), .A1(n3780), .Z(n354));
Q_FDP0UA U10038 ( .D(n353), .QTFCLK( ), .Q(shiftedOData[49]));
Q_MX02 U10039 ( .S(n280), .A0(shiftedOData[49]), .A1(n3779), .Z(n353));
Q_FDP0UA U10040 ( .D(n352), .QTFCLK( ), .Q(shiftedOData[48]));
Q_MX02 U10041 ( .S(n280), .A0(shiftedOData[48]), .A1(n3778), .Z(n352));
Q_FDP0UA U10042 ( .D(n351), .QTFCLK( ), .Q(shiftedOData[47]));
Q_MX02 U10043 ( .S(n280), .A0(shiftedOData[47]), .A1(n3777), .Z(n351));
Q_FDP0UA U10044 ( .D(n350), .QTFCLK( ), .Q(shiftedOData[46]));
Q_MX02 U10045 ( .S(n280), .A0(shiftedOData[46]), .A1(n3776), .Z(n350));
Q_FDP0UA U10046 ( .D(n349), .QTFCLK( ), .Q(shiftedOData[45]));
Q_MX02 U10047 ( .S(n280), .A0(shiftedOData[45]), .A1(n3775), .Z(n349));
Q_FDP0UA U10048 ( .D(n348), .QTFCLK( ), .Q(shiftedOData[44]));
Q_MX02 U10049 ( .S(n280), .A0(shiftedOData[44]), .A1(n3774), .Z(n348));
Q_FDP0UA U10050 ( .D(n347), .QTFCLK( ), .Q(shiftedOData[43]));
Q_MX02 U10051 ( .S(n280), .A0(shiftedOData[43]), .A1(n3773), .Z(n347));
Q_FDP0UA U10052 ( .D(n346), .QTFCLK( ), .Q(shiftedOData[42]));
Q_MX02 U10053 ( .S(n280), .A0(shiftedOData[42]), .A1(n3772), .Z(n346));
Q_FDP0UA U10054 ( .D(n345), .QTFCLK( ), .Q(shiftedOData[41]));
Q_MX02 U10055 ( .S(n280), .A0(shiftedOData[41]), .A1(n3771), .Z(n345));
Q_FDP0UA U10056 ( .D(n344), .QTFCLK( ), .Q(shiftedOData[40]));
Q_MX02 U10057 ( .S(n280), .A0(shiftedOData[40]), .A1(n3770), .Z(n344));
Q_FDP0UA U10058 ( .D(n343), .QTFCLK( ), .Q(shiftedOData[39]));
Q_MX02 U10059 ( .S(n280), .A0(shiftedOData[39]), .A1(n3769), .Z(n343));
Q_FDP0UA U10060 ( .D(n342), .QTFCLK( ), .Q(shiftedOData[38]));
Q_MX02 U10061 ( .S(n280), .A0(shiftedOData[38]), .A1(n3768), .Z(n342));
Q_FDP0UA U10062 ( .D(n341), .QTFCLK( ), .Q(shiftedOData[37]));
Q_MX02 U10063 ( .S(n280), .A0(shiftedOData[37]), .A1(n3767), .Z(n341));
Q_FDP0UA U10064 ( .D(n340), .QTFCLK( ), .Q(shiftedOData[36]));
Q_MX02 U10065 ( .S(n280), .A0(shiftedOData[36]), .A1(n3766), .Z(n340));
Q_FDP0UA U10066 ( .D(n339), .QTFCLK( ), .Q(shiftedOData[35]));
Q_MX02 U10067 ( .S(n280), .A0(shiftedOData[35]), .A1(n3765), .Z(n339));
Q_FDP0UA U10068 ( .D(n338), .QTFCLK( ), .Q(shiftedOData[34]));
Q_MX02 U10069 ( .S(n280), .A0(shiftedOData[34]), .A1(n3764), .Z(n338));
Q_FDP0UA U10070 ( .D(n337), .QTFCLK( ), .Q(shiftedOData[33]));
Q_MX02 U10071 ( .S(n280), .A0(shiftedOData[33]), .A1(n3763), .Z(n337));
Q_FDP0UA U10072 ( .D(n336), .QTFCLK( ), .Q(shiftedOData[32]));
Q_MX02 U10073 ( .S(n280), .A0(shiftedOData[32]), .A1(n3762), .Z(n336));
Q_FDP0UA U10074 ( .D(n335), .QTFCLK( ), .Q(shiftedOData[31]));
Q_MX02 U10075 ( .S(n280), .A0(shiftedOData[31]), .A1(n3761), .Z(n335));
Q_FDP0UA U10076 ( .D(n334), .QTFCLK( ), .Q(shiftedOData[30]));
Q_MX02 U10077 ( .S(n280), .A0(shiftedOData[30]), .A1(n3760), .Z(n334));
Q_FDP0UA U10078 ( .D(n333), .QTFCLK( ), .Q(shiftedOData[29]));
Q_MX02 U10079 ( .S(n280), .A0(shiftedOData[29]), .A1(n3759), .Z(n333));
Q_FDP0UA U10080 ( .D(n332), .QTFCLK( ), .Q(shiftedOData[28]));
Q_MX02 U10081 ( .S(n280), .A0(shiftedOData[28]), .A1(n3758), .Z(n332));
Q_FDP0UA U10082 ( .D(n331), .QTFCLK( ), .Q(shiftedOData[27]));
Q_MX02 U10083 ( .S(n280), .A0(shiftedOData[27]), .A1(n3757), .Z(n331));
Q_FDP0UA U10084 ( .D(n330), .QTFCLK( ), .Q(shiftedOData[26]));
Q_MX02 U10085 ( .S(n280), .A0(shiftedOData[26]), .A1(n3756), .Z(n330));
Q_FDP0UA U10086 ( .D(n329), .QTFCLK( ), .Q(shiftedOData[25]));
Q_MX02 U10087 ( .S(n280), .A0(shiftedOData[25]), .A1(n3755), .Z(n329));
Q_FDP0UA U10088 ( .D(n328), .QTFCLK( ), .Q(shiftedOData[24]));
Q_MX02 U10089 ( .S(n280), .A0(shiftedOData[24]), .A1(n3754), .Z(n328));
Q_FDP0UA U10090 ( .D(n327), .QTFCLK( ), .Q(shiftedOData[23]));
Q_MX02 U10091 ( .S(n280), .A0(shiftedOData[23]), .A1(n3753), .Z(n327));
Q_FDP0UA U10092 ( .D(n326), .QTFCLK( ), .Q(shiftedOData[22]));
Q_MX02 U10093 ( .S(n280), .A0(shiftedOData[22]), .A1(n3752), .Z(n326));
Q_FDP0UA U10094 ( .D(n325), .QTFCLK( ), .Q(shiftedOData[21]));
Q_MX02 U10095 ( .S(n280), .A0(shiftedOData[21]), .A1(n3751), .Z(n325));
Q_FDP0UA U10096 ( .D(n324), .QTFCLK( ), .Q(shiftedOData[20]));
Q_MX02 U10097 ( .S(n280), .A0(shiftedOData[20]), .A1(n3750), .Z(n324));
Q_FDP0UA U10098 ( .D(n323), .QTFCLK( ), .Q(shiftedOData[19]));
Q_MX02 U10099 ( .S(n280), .A0(shiftedOData[19]), .A1(n3749), .Z(n323));
Q_FDP0UA U10100 ( .D(n322), .QTFCLK( ), .Q(shiftedOData[18]));
Q_MX02 U10101 ( .S(n280), .A0(shiftedOData[18]), .A1(n3748), .Z(n322));
Q_FDP0UA U10102 ( .D(n321), .QTFCLK( ), .Q(shiftedOData[17]));
Q_MX02 U10103 ( .S(n280), .A0(shiftedOData[17]), .A1(n3747), .Z(n321));
Q_FDP0UA U10104 ( .D(n320), .QTFCLK( ), .Q(shiftedOData[16]));
Q_MX02 U10105 ( .S(n280), .A0(shiftedOData[16]), .A1(n3746), .Z(n320));
Q_FDP0UA U10106 ( .D(n319), .QTFCLK( ), .Q(shiftedOData[15]));
Q_MX02 U10107 ( .S(n280), .A0(shiftedOData[15]), .A1(n3745), .Z(n319));
Q_FDP0UA U10108 ( .D(n318), .QTFCLK( ), .Q(shiftedOData[14]));
Q_MX02 U10109 ( .S(n280), .A0(shiftedOData[14]), .A1(n3744), .Z(n318));
Q_FDP0UA U10110 ( .D(n317), .QTFCLK( ), .Q(shiftedOData[13]));
Q_MX02 U10111 ( .S(n280), .A0(shiftedOData[13]), .A1(n3743), .Z(n317));
Q_FDP0UA U10112 ( .D(n316), .QTFCLK( ), .Q(shiftedOData[12]));
Q_MX02 U10113 ( .S(n280), .A0(shiftedOData[12]), .A1(n3742), .Z(n316));
Q_FDP0UA U10114 ( .D(n315), .QTFCLK( ), .Q(shiftedOData[11]));
Q_MX02 U10115 ( .S(n280), .A0(shiftedOData[11]), .A1(n3741), .Z(n315));
Q_FDP0UA U10116 ( .D(n314), .QTFCLK( ), .Q(shiftedOData[10]));
Q_MX02 U10117 ( .S(n280), .A0(shiftedOData[10]), .A1(n3740), .Z(n314));
Q_FDP0UA U10118 ( .D(n313), .QTFCLK( ), .Q(shiftedOData[9]));
Q_MX02 U10119 ( .S(n280), .A0(shiftedOData[9]), .A1(n3739), .Z(n313));
Q_FDP0UA U10120 ( .D(n312), .QTFCLK( ), .Q(shiftedOData[8]));
Q_MX02 U10121 ( .S(n280), .A0(shiftedOData[8]), .A1(n3738), .Z(n312));
Q_FDP0UA U10122 ( .D(n311), .QTFCLK( ), .Q(shiftedOData[7]));
Q_MX02 U10123 ( .S(n280), .A0(shiftedOData[7]), .A1(n3737), .Z(n311));
Q_FDP0UA U10124 ( .D(n310), .QTFCLK( ), .Q(shiftedOData[6]));
Q_MX02 U10125 ( .S(n280), .A0(shiftedOData[6]), .A1(n3736), .Z(n310));
Q_FDP0UA U10126 ( .D(n309), .QTFCLK( ), .Q(shiftedOData[5]));
Q_MX02 U10127 ( .S(n280), .A0(shiftedOData[5]), .A1(n3735), .Z(n309));
Q_FDP0UA U10128 ( .D(n308), .QTFCLK( ), .Q(shiftedOData[4]));
Q_MX02 U10129 ( .S(n280), .A0(shiftedOData[4]), .A1(n3734), .Z(n308));
Q_FDP0UA U10130 ( .D(n307), .QTFCLK( ), .Q(shiftedOData[3]));
Q_MX02 U10131 ( .S(n280), .A0(shiftedOData[3]), .A1(n3733), .Z(n307));
Q_FDP0UA U10132 ( .D(n306), .QTFCLK( ), .Q(shiftedOData[2]));
Q_MX02 U10133 ( .S(n280), .A0(shiftedOData[2]), .A1(n3732), .Z(n306));
Q_FDP0UA U10134 ( .D(n305), .QTFCLK( ), .Q(shiftedOData[1]));
Q_MX02 U10135 ( .S(n280), .A0(shiftedOData[1]), .A1(n3731), .Z(n305));
Q_FDP0UA U10136 ( .D(n304), .QTFCLK( ), .Q(shiftedOData[0]));
Q_MX02 U10137 ( .S(n280), .A0(shiftedOData[0]), .A1(n3730), .Z(n304));
Q_FDP0UA U10138 ( .D(n303), .QTFCLK( ), .Q(shiftCount[7]));
Q_MX02 U10139 ( .S(n280), .A0(shiftCount[7]), .A1(oFill[1]), .Z(n303));
Q_FDP0UA U10140 ( .D(n302), .QTFCLK( ), .Q(shiftCount[6]));
Q_MX02 U10141 ( .S(n280), .A0(shiftCount[6]), .A1(oFill[0]), .Z(n302));
Q_FDP0UA U10142 ( .D(n300), .QTFCLK( ), .Q(shiftCount[5]));
Q_INV U10143 ( .A(n280), .Z(n301));
Q_AN02 U10144 ( .A0(n301), .A1(shiftCount[5]), .Z(n300));
Q_FDP0UA U10145 ( .D(n299), .QTFCLK( ), .Q(shiftCount[4]));
Q_AN02 U10146 ( .A0(n301), .A1(shiftCount[4]), .Z(n299));
Q_FDP0UA U10147 ( .D(n298), .QTFCLK( ), .Q(shiftCount[3]));
Q_AN02 U10148 ( .A0(n301), .A1(shiftCount[3]), .Z(n298));
Q_FDP0UA U10149 ( .D(n297), .QTFCLK( ), .Q(shiftCount[2]));
Q_AN02 U10150 ( .A0(n301), .A1(shiftCount[2]), .Z(n297));
Q_FDP0UA U10151 ( .D(n296), .QTFCLK( ), .Q(shiftCount[1]));
Q_AN02 U10152 ( .A0(n301), .A1(shiftCount[1]), .Z(n296));
Q_FDP0UA U10153 ( .D(n295), .QTFCLK( ), .Q(shiftCount[0]));
Q_AN02 U10154 ( .A0(n301), .A1(shiftCount[0]), .Z(n295));
Q_FDP0UA U10155 ( .D(n294), .QTFCLK( ), .Q(oFill[3]));
Q_MX02 U10156 ( .S(n281), .A0(n1938), .A1(oFill[3]), .Z(n294));
Q_FDP0UA U10157 ( .D(n293), .QTFCLK( ), .Q(oFill[2]));
Q_MX02 U10158 ( .S(n281), .A0(n1939), .A1(oFill[2]), .Z(n293));
Q_FDP0UA U10159 ( .D(n292), .QTFCLK( ), .Q(oFill[1]));
Q_MX02 U10160 ( .S(n281), .A0(n1940), .A1(oFill[1]), .Z(n292));
Q_FDP0UA U10161 ( .D(n291), .QTFCLK( ), .Q(oFill[0]));
Q_MX02 U10162 ( .S(n281), .A0(n1941), .A1(oFill[0]), .Z(n291));
Q_FDP0UA U10163 ( .D(n290), .QTFCLK( ), .Q(oSt));
Q_MX02 U10164 ( .S(n287), .A0(n275), .A1(oSt), .Z(n290));
Q_AN02 U10165 ( .A0(n280), .A1(n289), .Z(n278));
Q_AN02 U10166 ( .A0(n280), .A1(n288), .Z(n277));
Q_INV U10167 ( .A(oFill[2]), .Z(n289));
Q_AN03 U10168 ( .A0(oFill[3]), .A1(oFill[2]), .A2(n280), .Z(n276));
Q_AN02 U10169 ( .A0(n279), .A1(oSt), .Z(n280));
Q_AN02 U10170 ( .A0(n279), .A1(n286), .Z(n287));
Q_MX02 U10171 ( .S(oSt), .A0(n284), .A1(n285), .Z(n286));
Q_AN02 U10172 ( .A0(n279), .A1(n282), .Z(n283));
Q_ND02 U10173 ( .A0(oSt), .A1(rstDoneD2), .Z(n282));
Q_INV U10174 ( .A(rstDoneD2), .Z(n285));
Q_AN02 U10175 ( .A0(n275), .A1(n284), .Z(n281));
Q_INV U10176 ( .A(nps), .Z(n284));
Q_NR02 U10177 ( .A0(xc_top.GFReset), .A1(oSt), .Z(n275));
Q_INV U10178 ( .A(xc_top.GFReset), .Z(n279));
Q_FDP0B U10179 ( .D(n5586), .QTFCLK( ), .Q(n274));
Q_FDP0UA U10180 ( .D(xptrN[2]), .QTFCLK( ), .Q(n273));
Q_FDP0UA U10181 ( .D(xptrN[3]), .QTFCLK( ), .Q(n272));
Q_FDP0UA U10182 ( .D(xptrN[4]), .QTFCLK( ), .Q(n271));
Q_FDP0UA U10183 ( .D(xptrN[5]), .QTFCLK( ), .Q(n270));
Q_FDP0UA U10184 ( .D(xptrN[6]), .QTFCLK( ), .Q(n269));
Q_FDP0UA U10185 ( .D(xptrN[7]), .QTFCLK( ), .Q(n268));
Q_FDP0UA U10186 ( .D(xptrN[8]), .QTFCLK( ), .Q(n267));
Q_FDP0UA U10187 ( .D(xptrN[9]), .QTFCLK( ), .Q(n266));
Q_FDP0UA U10188 ( .D(xptrN[10]), .QTFCLK( ), .Q(n265));
Q_FDP0UA U10189 ( .D(xptrN[11]), .QTFCLK( ), .Q(n264));
Q_FDP0UA U10190 ( .D(xptrN[12]), .QTFCLK( ), .Q(n263));
Q_FDP0UA U10191 ( .D(xptrN[13]), .QTFCLK( ), .Q(n262));
Q_FDP0UA U10192 ( .D(xptrN[14]), .QTFCLK( ), .Q(n261));
Q_FDP0UA U10193 ( .D(xptrN[15]), .QTFCLK( ), .Q(n260));
Q_FDP0UA U10194 ( .D(xptrN[16]), .QTFCLK( ), .Q(n259));
Q_FDP0UA U10195 ( .D(ififoXdataFinal[0]), .QTFCLK( ), .Q(n258));
Q_FDP0UA U10196 ( .D(ififoXdataFinal[1]), .QTFCLK( ), .Q(n257));
Q_FDP0UA U10197 ( .D(ififoXdataFinal[2]), .QTFCLK( ), .Q(n256));
Q_FDP0UA U10198 ( .D(ififoXdataFinal[3]), .QTFCLK( ), .Q(n255));
Q_FDP0UA U10199 ( .D(ififoXdataFinal[4]), .QTFCLK( ), .Q(n254));
Q_FDP0UA U10200 ( .D(ififoXdataFinal[5]), .QTFCLK( ), .Q(n253));
Q_FDP0UA U10201 ( .D(ififoXdataFinal[6]), .QTFCLK( ), .Q(n252));
Q_FDP0UA U10202 ( .D(ififoXdataFinal[7]), .QTFCLK( ), .Q(n251));
Q_FDP0UA U10203 ( .D(ififoXdataFinal[8]), .QTFCLK( ), .Q(n250));
Q_FDP0UA U10204 ( .D(ififoXdataFinal[9]), .QTFCLK( ), .Q(n249));
Q_FDP0UA U10205 ( .D(ififoXdataFinal[10]), .QTFCLK( ), .Q(n248));
Q_FDP0UA U10206 ( .D(ififoXdataFinal[11]), .QTFCLK( ), .Q(n247));
Q_FDP0UA U10207 ( .D(ififoXdataFinal[12]), .QTFCLK( ), .Q(n246));
Q_FDP0UA U10208 ( .D(ififoXdataFinal[13]), .QTFCLK( ), .Q(n245));
Q_FDP0UA U10209 ( .D(ififoXdataFinal[14]), .QTFCLK( ), .Q(n244));
Q_FDP0UA U10210 ( .D(ififoXdataFinal[15]), .QTFCLK( ), .Q(n243));
Q_FDP0UA U10211 ( .D(ififoXdataFinal[16]), .QTFCLK( ), .Q(n242));
Q_FDP0UA U10212 ( .D(ififoXdataFinal[17]), .QTFCLK( ), .Q(n241));
Q_FDP0UA U10213 ( .D(ififoXdataFinal[18]), .QTFCLK( ), .Q(n240));
Q_FDP0UA U10214 ( .D(ififoXdataFinal[19]), .QTFCLK( ), .Q(n239));
Q_FDP0UA U10215 ( .D(ififoXdataFinal[20]), .QTFCLK( ), .Q(n238));
Q_FDP0UA U10216 ( .D(ififoXdataFinal[21]), .QTFCLK( ), .Q(n237));
Q_FDP0UA U10217 ( .D(ififoXdataFinal[22]), .QTFCLK( ), .Q(n236));
Q_FDP0UA U10218 ( .D(ififoXdataFinal[23]), .QTFCLK( ), .Q(n235));
Q_FDP0UA U10219 ( .D(ififoXdataFinal[24]), .QTFCLK( ), .Q(n234));
Q_FDP0UA U10220 ( .D(ififoXdataFinal[25]), .QTFCLK( ), .Q(n233));
Q_FDP0UA U10221 ( .D(ififoXdataFinal[26]), .QTFCLK( ), .Q(n232));
Q_FDP0UA U10222 ( .D(ififoXdataFinal[27]), .QTFCLK( ), .Q(n231));
Q_FDP0UA U10223 ( .D(ififoXdataFinal[28]), .QTFCLK( ), .Q(n230));
Q_FDP0UA U10224 ( .D(ififoXdataFinal[29]), .QTFCLK( ), .Q(n229));
Q_FDP0UA U10225 ( .D(ififoXdataFinal[30]), .QTFCLK( ), .Q(n228));
Q_FDP0UA U10226 ( .D(ififoXdataFinal[31]), .QTFCLK( ), .Q(n227));
Q_FDP0UA U10227 ( .D(ififoXdataFinal[32]), .QTFCLK( ), .Q(n226));
Q_FDP0UA U10228 ( .D(ififoXdataFinal[33]), .QTFCLK( ), .Q(n225));
Q_FDP0UA U10229 ( .D(ififoXdataFinal[34]), .QTFCLK( ), .Q(n224));
Q_FDP0UA U10230 ( .D(ififoXdataFinal[35]), .QTFCLK( ), .Q(n223));
Q_FDP0UA U10231 ( .D(ififoXdataFinal[36]), .QTFCLK( ), .Q(n222));
Q_FDP0UA U10232 ( .D(ififoXdataFinal[37]), .QTFCLK( ), .Q(n221));
Q_FDP0UA U10233 ( .D(ififoXdataFinal[38]), .QTFCLK( ), .Q(n220));
Q_FDP0UA U10234 ( .D(ififoXdataFinal[39]), .QTFCLK( ), .Q(n219));
Q_FDP0UA U10235 ( .D(ififoXdataFinal[40]), .QTFCLK( ), .Q(n218));
Q_FDP0UA U10236 ( .D(ififoXdataFinal[41]), .QTFCLK( ), .Q(n217));
Q_FDP0UA U10237 ( .D(ififoXdataFinal[42]), .QTFCLK( ), .Q(n216));
Q_FDP0UA U10238 ( .D(ififoXdataFinal[43]), .QTFCLK( ), .Q(n215));
Q_FDP0UA U10239 ( .D(ififoXdataFinal[44]), .QTFCLK( ), .Q(n214));
Q_FDP0UA U10240 ( .D(ififoXdataFinal[45]), .QTFCLK( ), .Q(n213));
Q_FDP0UA U10241 ( .D(ififoXdataFinal[46]), .QTFCLK( ), .Q(n212));
Q_FDP0UA U10242 ( .D(ififoXdataFinal[47]), .QTFCLK( ), .Q(n211));
Q_FDP0UA U10243 ( .D(ififoXdataFinal[48]), .QTFCLK( ), .Q(n210));
Q_FDP0UA U10244 ( .D(ififoXdataFinal[49]), .QTFCLK( ), .Q(n209));
Q_FDP0UA U10245 ( .D(ififoXdataFinal[50]), .QTFCLK( ), .Q(n208));
Q_FDP0UA U10246 ( .D(ififoXdataFinal[51]), .QTFCLK( ), .Q(n207));
Q_FDP0UA U10247 ( .D(ififoXdataFinal[52]), .QTFCLK( ), .Q(n206));
Q_FDP0UA U10248 ( .D(ififoXdataFinal[53]), .QTFCLK( ), .Q(n205));
Q_FDP0UA U10249 ( .D(ififoXdataFinal[54]), .QTFCLK( ), .Q(n204));
Q_FDP0UA U10250 ( .D(ififoXdataFinal[55]), .QTFCLK( ), .Q(n203));
Q_FDP0UA U10251 ( .D(ififoXdataFinal[56]), .QTFCLK( ), .Q(n202));
Q_FDP0UA U10252 ( .D(ififoXdataFinal[57]), .QTFCLK( ), .Q(n201));
Q_FDP0UA U10253 ( .D(ififoXdataFinal[58]), .QTFCLK( ), .Q(n200));
Q_FDP0UA U10254 ( .D(ififoXdataFinal[59]), .QTFCLK( ), .Q(n199));
Q_FDP0UA U10255 ( .D(ififoXdataFinal[60]), .QTFCLK( ), .Q(n198));
Q_FDP0UA U10256 ( .D(ififoXdataFinal[61]), .QTFCLK( ), .Q(n197));
Q_FDP0UA U10257 ( .D(ififoXdataFinal[62]), .QTFCLK( ), .Q(n196));
Q_FDP0UA U10258 ( .D(ififoXdataFinal[63]), .QTFCLK( ), .Q(n195));
Q_FDP0UA U10259 ( .D(ififoXdataFinal[64]), .QTFCLK( ), .Q(n194));
Q_FDP0UA U10260 ( .D(ififoXdataFinal[65]), .QTFCLK( ), .Q(n193));
Q_FDP0UA U10261 ( .D(ififoXdataFinal[66]), .QTFCLK( ), .Q(n192));
Q_FDP0UA U10262 ( .D(ififoXdataFinal[67]), .QTFCLK( ), .Q(n191));
Q_FDP0UA U10263 ( .D(ififoXdataFinal[68]), .QTFCLK( ), .Q(n190));
Q_FDP0UA U10264 ( .D(ififoXdataFinal[69]), .QTFCLK( ), .Q(n189));
Q_FDP0UA U10265 ( .D(ififoXdataFinal[70]), .QTFCLK( ), .Q(n188));
Q_FDP0UA U10266 ( .D(ififoXdataFinal[71]), .QTFCLK( ), .Q(n187));
Q_FDP0UA U10267 ( .D(ififoXdataFinal[72]), .QTFCLK( ), .Q(n186));
Q_FDP0UA U10268 ( .D(ififoXdataFinal[73]), .QTFCLK( ), .Q(n185));
Q_FDP0UA U10269 ( .D(ififoXdataFinal[74]), .QTFCLK( ), .Q(n184));
Q_FDP0UA U10270 ( .D(ififoXdataFinal[75]), .QTFCLK( ), .Q(n183));
Q_FDP0UA U10271 ( .D(ififoXdataFinal[76]), .QTFCLK( ), .Q(n182));
Q_FDP0UA U10272 ( .D(ififoXdataFinal[77]), .QTFCLK( ), .Q(n181));
Q_FDP0UA U10273 ( .D(ififoXdataFinal[78]), .QTFCLK( ), .Q(n180));
Q_FDP0UA U10274 ( .D(ififoXdataFinal[79]), .QTFCLK( ), .Q(n179));
Q_FDP0UA U10275 ( .D(ififoXdataFinal[80]), .QTFCLK( ), .Q(n178));
Q_FDP0UA U10276 ( .D(ififoXdataFinal[81]), .QTFCLK( ), .Q(n177));
Q_FDP0UA U10277 ( .D(ififoXdataFinal[82]), .QTFCLK( ), .Q(n176));
Q_FDP0UA U10278 ( .D(ififoXdataFinal[83]), .QTFCLK( ), .Q(n175));
Q_FDP0UA U10279 ( .D(ififoXdataFinal[84]), .QTFCLK( ), .Q(n174));
Q_FDP0UA U10280 ( .D(ififoXdataFinal[85]), .QTFCLK( ), .Q(n173));
Q_FDP0UA U10281 ( .D(ififoXdataFinal[86]), .QTFCLK( ), .Q(n172));
Q_FDP0UA U10282 ( .D(ififoXdataFinal[87]), .QTFCLK( ), .Q(n171));
Q_FDP0UA U10283 ( .D(ififoXdataFinal[88]), .QTFCLK( ), .Q(n170));
Q_FDP0UA U10284 ( .D(ififoXdataFinal[89]), .QTFCLK( ), .Q(n169));
Q_FDP0UA U10285 ( .D(ififoXdataFinal[90]), .QTFCLK( ), .Q(n168));
Q_FDP0UA U10286 ( .D(ififoXdataFinal[91]), .QTFCLK( ), .Q(n167));
Q_FDP0UA U10287 ( .D(ififoXdataFinal[92]), .QTFCLK( ), .Q(n166));
Q_FDP0UA U10288 ( .D(ififoXdataFinal[93]), .QTFCLK( ), .Q(n165));
Q_FDP0UA U10289 ( .D(ififoXdataFinal[94]), .QTFCLK( ), .Q(n164));
Q_FDP0UA U10290 ( .D(ififoXdataFinal[95]), .QTFCLK( ), .Q(n163));
Q_FDP0UA U10291 ( .D(ififoXdataFinal[96]), .QTFCLK( ), .Q(n162));
Q_FDP0UA U10292 ( .D(ififoXdataFinal[97]), .QTFCLK( ), .Q(n161));
Q_FDP0UA U10293 ( .D(ififoXdataFinal[98]), .QTFCLK( ), .Q(n160));
Q_FDP0UA U10294 ( .D(ififoXdataFinal[99]), .QTFCLK( ), .Q(n159));
Q_FDP0UA U10295 ( .D(ififoXdataFinal[100]), .QTFCLK( ), .Q(n158));
Q_FDP0UA U10296 ( .D(ififoXdataFinal[101]), .QTFCLK( ), .Q(n157));
Q_FDP0UA U10297 ( .D(ififoXdataFinal[102]), .QTFCLK( ), .Q(n156));
Q_FDP0UA U10298 ( .D(ififoXdataFinal[103]), .QTFCLK( ), .Q(n155));
Q_FDP0UA U10299 ( .D(ififoXdataFinal[104]), .QTFCLK( ), .Q(n154));
Q_FDP0UA U10300 ( .D(ififoXdataFinal[105]), .QTFCLK( ), .Q(n153));
Q_FDP0UA U10301 ( .D(ififoXdataFinal[106]), .QTFCLK( ), .Q(n152));
Q_FDP0UA U10302 ( .D(ififoXdataFinal[107]), .QTFCLK( ), .Q(n151));
Q_FDP0UA U10303 ( .D(ififoXdataFinal[108]), .QTFCLK( ), .Q(n150));
Q_FDP0UA U10304 ( .D(ififoXdataFinal[109]), .QTFCLK( ), .Q(n149));
Q_FDP0UA U10305 ( .D(ififoXdataFinal[110]), .QTFCLK( ), .Q(n148));
Q_FDP0UA U10306 ( .D(ififoXdataFinal[111]), .QTFCLK( ), .Q(n147));
Q_FDP0UA U10307 ( .D(ififoXdataFinal[112]), .QTFCLK( ), .Q(n146));
Q_FDP0UA U10308 ( .D(ififoXdataFinal[113]), .QTFCLK( ), .Q(n145));
Q_FDP0UA U10309 ( .D(ififoXdataFinal[114]), .QTFCLK( ), .Q(n144));
Q_FDP0UA U10310 ( .D(ififoXdataFinal[115]), .QTFCLK( ), .Q(n143));
Q_FDP0UA U10311 ( .D(ififoXdataFinal[116]), .QTFCLK( ), .Q(n142));
Q_FDP0UA U10312 ( .D(ififoXdataFinal[117]), .QTFCLK( ), .Q(n141));
Q_FDP0UA U10313 ( .D(ififoXdataFinal[118]), .QTFCLK( ), .Q(n140));
Q_FDP0UA U10314 ( .D(ififoXdataFinal[119]), .QTFCLK( ), .Q(n139));
Q_FDP0UA U10315 ( .D(ififoXdataFinal[120]), .QTFCLK( ), .Q(n138));
Q_FDP0UA U10316 ( .D(ififoXdataFinal[121]), .QTFCLK( ), .Q(n137));
Q_FDP0UA U10317 ( .D(ififoXdataFinal[122]), .QTFCLK( ), .Q(n136));
Q_FDP0UA U10318 ( .D(ififoXdataFinal[123]), .QTFCLK( ), .Q(n135));
Q_FDP0UA U10319 ( .D(ififoXdataFinal[124]), .QTFCLK( ), .Q(n134));
Q_FDP0UA U10320 ( .D(ififoXdataFinal[125]), .QTFCLK( ), .Q(n133));
Q_FDP0UA U10321 ( .D(ififoXdataFinal[126]), .QTFCLK( ), .Q(n132));
Q_FDP0UA U10322 ( .D(ififoXdataFinal[127]), .QTFCLK( ), .Q(n131));
Q_FDP0UA U10323 ( .D(ififoXdataFinal[128]), .QTFCLK( ), .Q(n130));
Q_FDP0UA U10324 ( .D(ififoXdataFinal[129]), .QTFCLK( ), .Q(n129));
Q_FDP0UA U10325 ( .D(ififoXdataFinal[130]), .QTFCLK( ), .Q(n128));
Q_FDP0UA U10326 ( .D(ififoXdataFinal[131]), .QTFCLK( ), .Q(n127));
Q_FDP0UA U10327 ( .D(ififoXdataFinal[132]), .QTFCLK( ), .Q(n126));
Q_FDP0UA U10328 ( .D(ififoXdataFinal[133]), .QTFCLK( ), .Q(n125));
Q_FDP0UA U10329 ( .D(ififoXdataFinal[134]), .QTFCLK( ), .Q(n124));
Q_FDP0UA U10330 ( .D(ififoXdataFinal[135]), .QTFCLK( ), .Q(n123));
Q_FDP0UA U10331 ( .D(ififoXdataFinal[136]), .QTFCLK( ), .Q(n122));
Q_FDP0UA U10332 ( .D(ififoXdataFinal[137]), .QTFCLK( ), .Q(n121));
Q_FDP0UA U10333 ( .D(ififoXdataFinal[138]), .QTFCLK( ), .Q(n120));
Q_FDP0UA U10334 ( .D(ififoXdataFinal[139]), .QTFCLK( ), .Q(n119));
Q_FDP0UA U10335 ( .D(ififoXdataFinal[140]), .QTFCLK( ), .Q(n118));
Q_FDP0UA U10336 ( .D(ififoXdataFinal[141]), .QTFCLK( ), .Q(n117));
Q_FDP0UA U10337 ( .D(ififoXdataFinal[142]), .QTFCLK( ), .Q(n116));
Q_FDP0UA U10338 ( .D(ififoXdataFinal[143]), .QTFCLK( ), .Q(n115));
Q_FDP0UA U10339 ( .D(ififoXdataFinal[144]), .QTFCLK( ), .Q(n114));
Q_FDP0UA U10340 ( .D(ififoXdataFinal[145]), .QTFCLK( ), .Q(n113));
Q_FDP0UA U10341 ( .D(ififoXdataFinal[146]), .QTFCLK( ), .Q(n112));
Q_FDP0UA U10342 ( .D(ififoXdataFinal[147]), .QTFCLK( ), .Q(n111));
Q_FDP0UA U10343 ( .D(ififoXdataFinal[148]), .QTFCLK( ), .Q(n110));
Q_FDP0UA U10344 ( .D(ififoXdataFinal[149]), .QTFCLK( ), .Q(n109));
Q_FDP0UA U10345 ( .D(ififoXdataFinal[150]), .QTFCLK( ), .Q(n108));
Q_FDP0UA U10346 ( .D(ififoXdataFinal[151]), .QTFCLK( ), .Q(n107));
Q_FDP0UA U10347 ( .D(ififoXdataFinal[152]), .QTFCLK( ), .Q(n106));
Q_FDP0UA U10348 ( .D(ififoXdataFinal[153]), .QTFCLK( ), .Q(n105));
Q_FDP0UA U10349 ( .D(ififoXdataFinal[154]), .QTFCLK( ), .Q(n104));
Q_FDP0UA U10350 ( .D(ififoXdataFinal[155]), .QTFCLK( ), .Q(n103));
Q_FDP0UA U10351 ( .D(ififoXdataFinal[156]), .QTFCLK( ), .Q(n102));
Q_FDP0UA U10352 ( .D(ififoXdataFinal[157]), .QTFCLK( ), .Q(n101));
Q_FDP0UA U10353 ( .D(ififoXdataFinal[158]), .QTFCLK( ), .Q(n100));
Q_FDP0UA U10354 ( .D(ififoXdataFinal[159]), .QTFCLK( ), .Q(n99));
Q_FDP0UA U10355 ( .D(ififoXdataFinal[160]), .QTFCLK( ), .Q(n98));
Q_FDP0UA U10356 ( .D(ififoXdataFinal[161]), .QTFCLK( ), .Q(n97));
Q_FDP0UA U10357 ( .D(ififoXdataFinal[162]), .QTFCLK( ), .Q(n96));
Q_FDP0UA U10358 ( .D(ififoXdataFinal[163]), .QTFCLK( ), .Q(n95));
Q_FDP0UA U10359 ( .D(ififoXdataFinal[164]), .QTFCLK( ), .Q(n94));
Q_FDP0UA U10360 ( .D(ififoXdataFinal[165]), .QTFCLK( ), .Q(n93));
Q_FDP0UA U10361 ( .D(ififoXdataFinal[166]), .QTFCLK( ), .Q(n92));
Q_FDP0UA U10362 ( .D(ififoXdataFinal[167]), .QTFCLK( ), .Q(n91));
Q_FDP0UA U10363 ( .D(ififoXdataFinal[168]), .QTFCLK( ), .Q(n90));
Q_FDP0UA U10364 ( .D(ififoXdataFinal[169]), .QTFCLK( ), .Q(n89));
Q_FDP0UA U10365 ( .D(ififoXdataFinal[170]), .QTFCLK( ), .Q(n88));
Q_FDP0UA U10366 ( .D(ififoXdataFinal[171]), .QTFCLK( ), .Q(n87));
Q_FDP0UA U10367 ( .D(ififoXdataFinal[172]), .QTFCLK( ), .Q(n86));
Q_FDP0UA U10368 ( .D(ififoXdataFinal[173]), .QTFCLK( ), .Q(n85));
Q_FDP0UA U10369 ( .D(ififoXdataFinal[174]), .QTFCLK( ), .Q(n84));
Q_FDP0UA U10370 ( .D(ififoXdataFinal[175]), .QTFCLK( ), .Q(n83));
Q_FDP0UA U10371 ( .D(ififoXdataFinal[176]), .QTFCLK( ), .Q(n82));
Q_FDP0UA U10372 ( .D(ififoXdataFinal[177]), .QTFCLK( ), .Q(n81));
Q_FDP0UA U10373 ( .D(ififoXdataFinal[178]), .QTFCLK( ), .Q(n80));
Q_FDP0UA U10374 ( .D(ififoXdataFinal[179]), .QTFCLK( ), .Q(n79));
Q_FDP0UA U10375 ( .D(ififoXdataFinal[180]), .QTFCLK( ), .Q(n78));
Q_FDP0UA U10376 ( .D(ififoXdataFinal[181]), .QTFCLK( ), .Q(n77));
Q_FDP0UA U10377 ( .D(ififoXdataFinal[182]), .QTFCLK( ), .Q(n76));
Q_FDP0UA U10378 ( .D(ififoXdataFinal[183]), .QTFCLK( ), .Q(n75));
Q_FDP0UA U10379 ( .D(ififoXdataFinal[184]), .QTFCLK( ), .Q(n74));
Q_FDP0UA U10380 ( .D(ififoXdataFinal[185]), .QTFCLK( ), .Q(n73));
Q_FDP0UA U10381 ( .D(ififoXdataFinal[186]), .QTFCLK( ), .Q(n72));
Q_FDP0UA U10382 ( .D(ififoXdataFinal[187]), .QTFCLK( ), .Q(n71));
Q_FDP0UA U10383 ( .D(ififoXdataFinal[188]), .QTFCLK( ), .Q(n70));
Q_FDP0UA U10384 ( .D(ififoXdataFinal[189]), .QTFCLK( ), .Q(n69));
Q_FDP0UA U10385 ( .D(ififoXdataFinal[190]), .QTFCLK( ), .Q(n68));
Q_FDP0UA U10386 ( .D(ififoXdataFinal[191]), .QTFCLK( ), .Q(n67));
Q_FDP0UA U10387 ( .D(ififoXdataFinal[192]), .QTFCLK( ), .Q(n66));
Q_FDP0UA U10388 ( .D(ififoXdataFinal[193]), .QTFCLK( ), .Q(n65));
Q_FDP0UA U10389 ( .D(ififoXdataFinal[194]), .QTFCLK( ), .Q(n64));
Q_FDP0UA U10390 ( .D(ififoXdataFinal[195]), .QTFCLK( ), .Q(n63));
Q_FDP0UA U10391 ( .D(ififoXdataFinal[196]), .QTFCLK( ), .Q(n62));
Q_FDP0UA U10392 ( .D(ififoXdataFinal[197]), .QTFCLK( ), .Q(n61));
Q_FDP0UA U10393 ( .D(ififoXdataFinal[198]), .QTFCLK( ), .Q(n60));
Q_FDP0UA U10394 ( .D(ififoXdataFinal[199]), .QTFCLK( ), .Q(n59));
Q_FDP0UA U10395 ( .D(ififoXdataFinal[200]), .QTFCLK( ), .Q(n58));
Q_FDP0UA U10396 ( .D(ififoXdataFinal[201]), .QTFCLK( ), .Q(n57));
Q_FDP0UA U10397 ( .D(ififoXdataFinal[202]), .QTFCLK( ), .Q(n56));
Q_FDP0UA U10398 ( .D(ififoXdataFinal[203]), .QTFCLK( ), .Q(n55));
Q_FDP0UA U10399 ( .D(ififoXdataFinal[204]), .QTFCLK( ), .Q(n54));
Q_FDP0UA U10400 ( .D(ififoXdataFinal[205]), .QTFCLK( ), .Q(n53));
Q_FDP0UA U10401 ( .D(ififoXdataFinal[206]), .QTFCLK( ), .Q(n52));
Q_FDP0UA U10402 ( .D(ififoXdataFinal[207]), .QTFCLK( ), .Q(n51));
Q_FDP0UA U10403 ( .D(ififoXdataFinal[208]), .QTFCLK( ), .Q(n50));
Q_FDP0UA U10404 ( .D(ififoXdataFinal[209]), .QTFCLK( ), .Q(n49));
Q_FDP0UA U10405 ( .D(ififoXdataFinal[210]), .QTFCLK( ), .Q(n48));
Q_FDP0UA U10406 ( .D(ififoXdataFinal[211]), .QTFCLK( ), .Q(n47));
Q_FDP0UA U10407 ( .D(ififoXdataFinal[212]), .QTFCLK( ), .Q(n46));
Q_FDP0UA U10408 ( .D(ififoXdataFinal[213]), .QTFCLK( ), .Q(n45));
Q_FDP0UA U10409 ( .D(ififoXdataFinal[214]), .QTFCLK( ), .Q(n44));
Q_FDP0UA U10410 ( .D(ififoXdataFinal[215]), .QTFCLK( ), .Q(n43));
Q_FDP0UA U10411 ( .D(ififoXdataFinal[216]), .QTFCLK( ), .Q(n42));
Q_FDP0UA U10412 ( .D(ififoXdataFinal[217]), .QTFCLK( ), .Q(n41));
Q_FDP0UA U10413 ( .D(ififoXdataFinal[218]), .QTFCLK( ), .Q(n40));
Q_FDP0UA U10414 ( .D(ififoXdataFinal[219]), .QTFCLK( ), .Q(n39));
Q_FDP0UA U10415 ( .D(ififoXdataFinal[220]), .QTFCLK( ), .Q(n38));
Q_FDP0UA U10416 ( .D(ififoXdataFinal[221]), .QTFCLK( ), .Q(n37));
Q_FDP0UA U10417 ( .D(ififoXdataFinal[222]), .QTFCLK( ), .Q(n36));
Q_FDP0UA U10418 ( .D(ififoXdataFinal[223]), .QTFCLK( ), .Q(n35));
Q_FDP0UA U10419 ( .D(ififoXdataFinal[224]), .QTFCLK( ), .Q(n34));
Q_FDP0UA U10420 ( .D(ififoXdataFinal[225]), .QTFCLK( ), .Q(n33));
Q_FDP0UA U10421 ( .D(ififoXdataFinal[226]), .QTFCLK( ), .Q(n32));
Q_FDP0UA U10422 ( .D(ififoXdataFinal[227]), .QTFCLK( ), .Q(n31));
Q_FDP0UA U10423 ( .D(ififoXdataFinal[228]), .QTFCLK( ), .Q(n30));
Q_FDP0UA U10424 ( .D(ififoXdataFinal[229]), .QTFCLK( ), .Q(n29));
Q_FDP0UA U10425 ( .D(ififoXdataFinal[230]), .QTFCLK( ), .Q(n28));
Q_FDP0UA U10426 ( .D(ififoXdataFinal[231]), .QTFCLK( ), .Q(n27));
Q_FDP0UA U10427 ( .D(ififoXdataFinal[232]), .QTFCLK( ), .Q(n26));
Q_FDP0UA U10428 ( .D(ififoXdataFinal[233]), .QTFCLK( ), .Q(n25));
Q_FDP0UA U10429 ( .D(ififoXdataFinal[234]), .QTFCLK( ), .Q(n24));
Q_FDP0UA U10430 ( .D(ififoXdataFinal[235]), .QTFCLK( ), .Q(n23));
Q_FDP0UA U10431 ( .D(ififoXdataFinal[236]), .QTFCLK( ), .Q(n22));
Q_FDP0UA U10432 ( .D(ififoXdataFinal[237]), .QTFCLK( ), .Q(n21));
Q_FDP0UA U10433 ( .D(ififoXdataFinal[238]), .QTFCLK( ), .Q(n20));
Q_FDP0UA U10434 ( .D(ififoXdataFinal[239]), .QTFCLK( ), .Q(n19));
Q_FDP0UA U10435 ( .D(ififoXdataFinal[240]), .QTFCLK( ), .Q(n18));
Q_FDP0UA U10436 ( .D(ififoXdataFinal[241]), .QTFCLK( ), .Q(n17));
Q_FDP0UA U10437 ( .D(ififoXdataFinal[242]), .QTFCLK( ), .Q(n16));
Q_FDP0UA U10438 ( .D(ififoXdataFinal[243]), .QTFCLK( ), .Q(n15));
Q_FDP0UA U10439 ( .D(ififoXdataFinal[244]), .QTFCLK( ), .Q(n14));
Q_FDP0UA U10440 ( .D(ififoXdataFinal[245]), .QTFCLK( ), .Q(n13));
Q_FDP0UA U10441 ( .D(ififoXdataFinal[246]), .QTFCLK( ), .Q(n12));
Q_FDP0UA U10442 ( .D(ififoXdataFinal[247]), .QTFCLK( ), .Q(n11));
Q_FDP0UA U10443 ( .D(ififoXdataFinal[248]), .QTFCLK( ), .Q(n10));
Q_FDP0UA U10444 ( .D(ififoXdataFinal[249]), .QTFCLK( ), .Q(n9));
Q_FDP0UA U10445 ( .D(ififoXdataFinal[250]), .QTFCLK( ), .Q(n8));
Q_FDP0UA U10446 ( .D(ififoXdataFinal[251]), .QTFCLK( ), .Q(n7));
Q_FDP0UA U10447 ( .D(ififoXdataFinal[252]), .QTFCLK( ), .Q(n6));
Q_FDP0UA U10448 ( .D(ififoXdataFinal[253]), .QTFCLK( ), .Q(n5));
Q_FDP0UA U10449 ( .D(ififoXdataFinal[254]), .QTFCLK( ), .Q(n4));
Q_FDP0UA U10450 ( .D(ififoXdataFinal[255]), .QTFCLK( ), .Q(n3));
Q_XOR2 U10451 ( .A0(n3347), .A1(n3470), .Z(n3346));
Q_OA21 U10452 ( .A0(head[32]), .A1(head[33]), .B0(head[35]), .Z(n6061));
Q_AD01 U10453 ( .CI(n6133), .A0(vlen[8]), .B0(n6146), .S(n6132), .CO(n2));
Q_XNR3 U10454 ( .A0(n2), .A1(vlen[9]), .A2(pktl[9]), .Z(n6131));
Q_OR03 U10455 ( .A0(n278), .A1(n277), .A2(n276), .Z(n9332));
Q_AN02 U10456 ( .A0(n5710), .A1(n5834), .Z(n1));
Q_XOR2 U10457 ( .A0(oFill[3]), .A1(oFill[2]), .Z(n288));
`ifdef CBV

reg [255:0] ixc_gfm_ofifo [0:32767];
always @(n5631 or oMark[255] or oMark[254] or oMark[253] or oMark[252]
 or oMark[251] or oMark[250] or oMark[249] or oMark[248] or oMark[247] or oMark[246] or oMark[245] or oMark[244]
 or oMark[243] or oMark[242] or oMark[241] or oMark[240] or oMark[239] or oMark[238] or oMark[237] or oMark[236]
 or oMark[235] or oMark[234] or oMark[233] or oMark[232] or oMark[231] or oMark[230] or oMark[229] or oMark[228]
 or oMark[227] or oMark[226] or oMark[225] or oMark[224] or oMark[223] or oMark[222] or oMark[221] or oMark[220]
 or oMark[219] or oMark[218] or oMark[217] or oMark[216] or oMark[215] or oMark[214] or oMark[213] or oMark[212]
 or oMark[211] or oMark[210] or oMark[209] or oMark[208] or oMark[207] or oMark[206] or oMark[205] or oMark[204]
 or oMark[203] or oMark[202] or oMark[201] or oMark[200] or oMark[199] or oMark[198] or oMark[197] or oMark[196]
 or oMark[195] or oMark[194] or oMark[193] or oMark[192] or oMark[191] or oMark[190] or oMark[189] or oMark[188]
 or oMark[187] or oMark[186] or oMark[185] or oMark[184] or oMark[183] or oMark[182] or oMark[181] or oMark[180]
 or oMark[179] or oMark[178] or oMark[177] or oMark[176] or oMark[175] or oMark[174] or oMark[173] or oMark[172]
 or oMark[171] or oMark[170] or oMark[169] or oMark[168] or oMark[167] or oMark[166] or oMark[165] or oMark[164]
 or oMark[163] or oMark[162] or oMark[161] or oMark[160] or oMark[159] or oMark[158] or oMark[157] or oMark[156]
 or oMark[155] or oMark[154] or oMark[153] or oMark[152] or oMark[151] or oMark[150] or oMark[149] or oMark[148]
 or oMark[147] or oMark[146] or oMark[145] or oMark[144] or oMark[143] or oMark[142] or oMark[141] or oMark[140]
 or oMark[139] or oMark[138] or oMark[137] or oMark[136] or oMark[135] or oMark[134] or oMark[133] or oMark[132]
 or oMark[131] or oMark[130] or oMark[129] or oMark[128] or oMark[127] or oMark[126] or oMark[125] or oMark[124]
 or oMark[123] or oMark[122] or oMark[121] or oMark[120] or oMark[119] or oMark[118] or oMark[117] or oMark[116]
 or oMark[115] or oMark[114] or oMark[113] or oMark[112] or oMark[111] or oMark[110] or oMark[109] or oMark[108]
 or oMark[107] or oMark[106] or oMark[105] or oMark[104] or oMark[103] or oMark[102] or oMark[101] or oMark[100]
 or oMark[99] or oMark[98] or oMark[97] or oMark[96] or oMark[95] or oMark[94] or oMark[93] or oMark[92]
 or oMark[91] or oMark[90] or oMark[89] or oMark[88] or oMark[87] or oMark[86] or oMark[85] or oMark[84]
 or oMark[83] or oMark[82] or oMark[81] or oMark[80] or oMark[79] or oMark[78] or oMark[77] or oMark[76]
 or oMark[75] or oMark[74] or oMark[73] or oMark[72] or oMark[71] or oMark[70] or oMark[69] or oMark[68]
 or oMark[67] or oMark[66] or oMark[65] or oMark[64] or oMark[63] or oMark[62] or oMark[61] or oMark[60]
 or oMark[59] or oMark[58] or oMark[57] or oMark[56] or oMark[55] or oMark[54] or oMark[53] or oMark[52]
 or oMark[51] or oMark[50] or oMark[49] or oMark[48] or oMark[47] or oMark[46] or oMark[45] or oMark[44]
 or oMark[43] or oMark[42] or oMark[41] or oMark[40] or oMark[39] or oMark[38] or oMark[37] or oMark[36]
 or oMark[35] or oMark[34] or oMark[33] or oMark[32] or oMark[31] or oMark[30] or oMark[29] or oMark[28]
 or oMark[27] or oMark[26] or oMark[25] or oMark[24] or oMark[23] or oMark[22] or oMark[21] or oMark[20]
 or oMark[19] or oMark[18] or oMark[17] or oMark[16] or oMark[15] or oMark[14] or oMark[13] or oMark[12]
 or oMark[11] or oMark[10] or oMark[9] or oMark[8] or oMark[7] or oMark[6] or oMark[5] or oMark[4]
 or oMark[3] or oMark[2] or oMark[1] or oMark[0] or n6882 or ofifoAddr0[14] or ofifoAddr0[13] or ofifoAddr0[12]
 or ofifoAddr0[11] or ofifoAddr0[10] or ofifoAddr0[9] or ofifoAddr0[8] or ofifoAddr0[7] or ofifoAddr0[6] or ofifoAddr0[5] or ofifoAddr0[4]
 or ofifoAddr0[3] or ofifoAddr0[2] or ofifoAddr0[1] or ofifoAddr0[0] or ofifoData[255] or ofifoData[254] or ofifoData[253] or ofifoData[252]
 or ofifoData[251] or ofifoData[250] or ofifoData[249] or ofifoData[248] or ofifoData[247] or ofifoData[246] or ofifoData[245] or ofifoData[244]
 or ofifoData[243] or ofifoData[242] or ofifoData[241] or ofifoData[240] or ofifoData[239] or ofifoData[238] or ofifoData[237] or ofifoData[236]
 or ofifoData[235] or ofifoData[234] or ofifoData[233] or ofifoData[232] or ofifoData[231] or ofifoData[230] or ofifoData[229] or ofifoData[228]
 or ofifoData[227] or ofifoData[226] or ofifoData[225] or ofifoData[224] or ofifoData[223] or ofifoData[222] or ofifoData[221] or ofifoData[220]
 or ofifoData[219] or ofifoData[218] or ofifoData[217] or ofifoData[216] or ofifoData[215] or ofifoData[214] or ofifoData[213] or ofifoData[212]
 or ofifoData[211] or ofifoData[210] or ofifoData[209] or ofifoData[208] or ofifoData[207] or ofifoData[206] or ofifoData[205] or ofifoData[204]
 or ofifoData[203] or ofifoData[202] or ofifoData[201] or ofifoData[200] or ofifoData[199] or ofifoData[198] or ofifoData[197] or ofifoData[196]
 or ofifoData[195] or ofifoData[194] or ofifoData[193] or ofifoData[192] or ofifoData[191] or ofifoData[190] or ofifoData[189] or ofifoData[188]
 or ofifoData[187] or ofifoData[186] or ofifoData[185] or ofifoData[184] or ofifoData[183] or ofifoData[182] or ofifoData[181] or ofifoData[180]
 or ofifoData[179] or ofifoData[178] or ofifoData[177] or ofifoData[176] or ofifoData[175] or ofifoData[174] or ofifoData[173] or ofifoData[172]
 or ofifoData[171] or ofifoData[170] or ofifoData[169] or ofifoData[168] or ofifoData[167] or ofifoData[166] or ofifoData[165] or ofifoData[164]
 or ofifoData[163] or ofifoData[162] or ofifoData[161] or ofifoData[160] or ofifoData[159] or ofifoData[158] or ofifoData[157] or ofifoData[156]
 or ofifoData[155] or ofifoData[154] or ofifoData[153] or ofifoData[152] or ofifoData[151] or ofifoData[150] or ofifoData[149] or ofifoData[148]
 or ofifoData[147] or ofifoData[146] or ofifoData[145] or ofifoData[144] or ofifoData[143] or ofifoData[142] or ofifoData[141] or ofifoData[140]
 or ofifoData[139] or ofifoData[138] or ofifoData[137] or ofifoData[136] or ofifoData[135] or ofifoData[134] or ofifoData[133] or ofifoData[132]
 or ofifoData[131] or ofifoData[130] or ofifoData[129] or ofifoData[128] or ofifoData[127] or ofifoData[126] or ofifoData[125] or ofifoData[124]
 or ofifoData[123] or ofifoData[122] or ofifoData[121] or ofifoData[120] or ofifoData[119] or ofifoData[118] or ofifoData[117] or ofifoData[116]
 or ofifoData[115] or ofifoData[114] or ofifoData[113] or ofifoData[112] or ofifoData[111] or ofifoData[110] or ofifoData[109] or ofifoData[108]
 or ofifoData[107] or ofifoData[106] or ofifoData[105] or ofifoData[104] or ofifoData[103] or ofifoData[102] or ofifoData[101] or ofifoData[100]
 or ofifoData[99] or ofifoData[98] or ofifoData[97] or ofifoData[96] or ofifoData[95] or ofifoData[94] or ofifoData[93] or ofifoData[92]
 or ofifoData[91] or ofifoData[90] or ofifoData[89] or ofifoData[88] or ofifoData[87] or ofifoData[86] or ofifoData[85] or ofifoData[84]
 or ofifoData[83] or ofifoData[82] or ofifoData[81] or ofifoData[80] or ofifoData[79] or ofifoData[78] or ofifoData[77] or ofifoData[76]
 or ofifoData[75] or ofifoData[74] or ofifoData[73] or ofifoData[72] or ofifoData[71] or ofifoData[70] or ofifoData[69] or ofifoData[68]
 or ofifoData[67] or ofifoData[66] or ofifoData[65] or ofifoData[64] or ofifoData[63] or ofifoData[62] or ofifoData[61] or ofifoData[60]
 or ofifoData[59] or ofifoData[58] or ofifoData[57] or ofifoData[56] or ofifoData[55] or ofifoData[54] or ofifoData[53] or ofifoData[52]
 or ofifoData[51] or ofifoData[50] or ofifoData[49] or ofifoData[48] or ofifoData[47] or ofifoData[46] or ofifoData[45] or ofifoData[44]
 or ofifoData[43] or ofifoData[42] or ofifoData[41] or ofifoData[40] or ofifoData[39] or ofifoData[38] or ofifoData[37] or ofifoData[36]
 or ofifoData[35] or ofifoData[34] or ofifoData[33] or ofifoData[32] or ofifoData[31] or ofifoData[30] or ofifoData[29] or ofifoData[28]
 or ofifoData[27] or ofifoData[26] or ofifoData[25] or ofifoData[24] or ofifoData[23] or ofifoData[22] or ofifoData[21] or ofifoData[20]
 or ofifoData[19] or ofifoData[18] or ofifoData[17] or ofifoData[16] or ofifoData[15] or ofifoData[14] or ofifoData[13] or ofifoData[12]
 or ofifoData[11] or ofifoData[10] or ofifoData[9] or ofifoData[8] or ofifoData[7] or ofifoData[6] or ofifoData[5] or ofifoData[4]
 or ofifoData[3] or ofifoData[2] or ofifoData[1] or ofifoData[0] or ofifoAddr1[14] or ofifoAddr1[13] or ofifoAddr1[12] or ofifoAddr1[11]
 or ofifoAddr1[10] or ofifoAddr1[9] or ofifoAddr1[8] or ofifoAddr1[7] or ofifoAddr1[6] or ofifoAddr1[5] or ofifoAddr1[4] or ofifoAddr1[3]
 or ofifoAddr1[2] or ofifoAddr1[1] or ofifoAddr1[0] or ofifoData[511] or ofifoData[510] or ofifoData[509] or ofifoData[508] or ofifoData[507]
 or ofifoData[506] or ofifoData[505] or ofifoData[504] or ofifoData[503] or ofifoData[502] or ofifoData[501] or ofifoData[500] or ofifoData[499]
 or ofifoData[498] or ofifoData[497] or ofifoData[496] or ofifoData[495] or ofifoData[494] or ofifoData[493] or ofifoData[492] or ofifoData[491]
 or ofifoData[490] or ofifoData[489] or ofifoData[488] or ofifoData[487] or ofifoData[486] or ofifoData[485] or ofifoData[484] or ofifoData[483]
 or ofifoData[482] or ofifoData[481] or ofifoData[480] or ofifoData[479] or ofifoData[478] or ofifoData[477] or ofifoData[476] or ofifoData[475]
 or ofifoData[474] or ofifoData[473] or ofifoData[472] or ofifoData[471] or ofifoData[470] or ofifoData[469] or ofifoData[468] or ofifoData[467]
 or ofifoData[466] or ofifoData[465] or ofifoData[464] or ofifoData[463] or ofifoData[462] or ofifoData[461] or ofifoData[460] or ofifoData[459]
 or ofifoData[458] or ofifoData[457] or ofifoData[456] or ofifoData[455] or ofifoData[454] or ofifoData[453] or ofifoData[452] or ofifoData[451]
 or ofifoData[450] or ofifoData[449] or ofifoData[448] or ofifoData[447] or ofifoData[446] or ofifoData[445] or ofifoData[444] or ofifoData[443]
 or ofifoData[442] or ofifoData[441] or ofifoData[440] or ofifoData[439] or ofifoData[438] or ofifoData[437] or ofifoData[436] or ofifoData[435]
 or ofifoData[434] or ofifoData[433] or ofifoData[432] or ofifoData[431] or ofifoData[430] or ofifoData[429] or ofifoData[428] or ofifoData[427]
 or ofifoData[426] or ofifoData[425] or ofifoData[424] or ofifoData[423] or ofifoData[422] or ofifoData[421] or ofifoData[420] or ofifoData[419]
 or ofifoData[418] or ofifoData[417] or ofifoData[416] or ofifoData[415] or ofifoData[414] or ofifoData[413] or ofifoData[412] or ofifoData[411]
 or ofifoData[410] or ofifoData[409] or ofifoData[408] or ofifoData[407] or ofifoData[406] or ofifoData[405] or ofifoData[404] or ofifoData[403]
 or ofifoData[402] or ofifoData[401] or ofifoData[400] or ofifoData[399] or ofifoData[398] or ofifoData[397] or ofifoData[396] or ofifoData[395]
 or ofifoData[394] or ofifoData[393] or ofifoData[392] or ofifoData[391] or ofifoData[390] or ofifoData[389] or ofifoData[388] or ofifoData[387]
 or ofifoData[386] or ofifoData[385] or ofifoData[384] or ofifoData[383] or ofifoData[382] or ofifoData[381] or ofifoData[380] or ofifoData[379]
 or ofifoData[378] or ofifoData[377] or ofifoData[376] or ofifoData[375] or ofifoData[374] or ofifoData[373] or ofifoData[372] or ofifoData[371]
 or ofifoData[370] or ofifoData[369] or ofifoData[368] or ofifoData[367] or ofifoData[366] or ofifoData[365] or ofifoData[364] or ofifoData[363]
 or ofifoData[362] or ofifoData[361] or ofifoData[360] or ofifoData[359] or ofifoData[358] or ofifoData[357] or ofifoData[356] or ofifoData[355]
 or ofifoData[354] or ofifoData[353] or ofifoData[352] or ofifoData[351] or ofifoData[350] or ofifoData[349] or ofifoData[348] or ofifoData[347]
 or ofifoData[346] or ofifoData[345] or ofifoData[344] or ofifoData[343] or ofifoData[342] or ofifoData[341] or ofifoData[340] or ofifoData[339]
 or ofifoData[338] or ofifoData[337] or ofifoData[336] or ofifoData[335] or ofifoData[334] or ofifoData[333] or ofifoData[332] or ofifoData[331]
 or ofifoData[330] or ofifoData[329] or ofifoData[328] or ofifoData[327] or ofifoData[326] or ofifoData[325] or ofifoData[324] or ofifoData[323]
 or ofifoData[322] or ofifoData[321] or ofifoData[320] or ofifoData[319] or ofifoData[318] or ofifoData[317] or ofifoData[316] or ofifoData[315]
 or ofifoData[314] or ofifoData[313] or ofifoData[312] or ofifoData[311] or ofifoData[310] or ofifoData[309] or ofifoData[308] or ofifoData[307]
 or ofifoData[306] or ofifoData[305] or ofifoData[304] or ofifoData[303] or ofifoData[302] or ofifoData[301] or ofifoData[300] or ofifoData[299]
 or ofifoData[298] or ofifoData[297] or ofifoData[296] or ofifoData[295] or ofifoData[294] or ofifoData[293] or ofifoData[292] or ofifoData[291]
 or ofifoData[290] or ofifoData[289] or ofifoData[288] or ofifoData[287] or ofifoData[286] or ofifoData[285] or ofifoData[284] or ofifoData[283]
 or ofifoData[282] or ofifoData[281] or ofifoData[280] or ofifoData[279] or ofifoData[278] or ofifoData[277] or ofifoData[276] or ofifoData[275]
 or ofifoData[274] or ofifoData[273] or ofifoData[272] or ofifoData[271] or ofifoData[270] or ofifoData[269] or ofifoData[268] or ofifoData[267]
 or ofifoData[266] or ofifoData[265] or ofifoData[264] or ofifoData[263] or ofifoData[262] or ofifoData[261] or ofifoData[260] or ofifoData[259]
 or ofifoData[258] or ofifoData[257] or ofifoData[256] or n5632 or ofifoAddr2[14] or ofifoAddr2[13] or ofifoAddr2[12] or ofifoAddr2[11]
 or ofifoAddr2[10] or ofifoAddr2[9] or ofifoAddr2[8] or ofifoAddr2[7] or ofifoAddr2[6] or ofifoAddr2[5] or ofifoAddr2[4] or ofifoAddr2[3]
 or ofifoAddr2[2] or ofifoAddr2[1] or ofifoAddr2[0] or ofifoData[767] or ofifoData[766] or ofifoData[765] or ofifoData[764] or ofifoData[763]
 or ofifoData[762] or ofifoData[761] or ofifoData[760] or ofifoData[759] or ofifoData[758] or ofifoData[757] or ofifoData[756] or ofifoData[755]
 or ofifoData[754] or ofifoData[753] or ofifoData[752] or ofifoData[751] or ofifoData[750] or ofifoData[749] or ofifoData[748] or ofifoData[747]
 or ofifoData[746] or ofifoData[745] or ofifoData[744] or ofifoData[743] or ofifoData[742] or ofifoData[741] or ofifoData[740] or ofifoData[739]
 or ofifoData[738] or ofifoData[737] or ofifoData[736] or ofifoData[735] or ofifoData[734] or ofifoData[733] or ofifoData[732] or ofifoData[731]
 or ofifoData[730] or ofifoData[729] or ofifoData[728] or ofifoData[727] or ofifoData[726] or ofifoData[725] or ofifoData[724] or ofifoData[723]
 or ofifoData[722] or ofifoData[721] or ofifoData[720] or ofifoData[719] or ofifoData[718] or ofifoData[717] or ofifoData[716] or ofifoData[715]
 or ofifoData[714] or ofifoData[713] or ofifoData[712] or ofifoData[711] or ofifoData[710] or ofifoData[709] or ofifoData[708] or ofifoData[707]
 or ofifoData[706] or ofifoData[705] or ofifoData[704] or ofifoData[703] or ofifoData[702] or ofifoData[701] or ofifoData[700] or ofifoData[699]
 or ofifoData[698] or ofifoData[697] or ofifoData[696] or ofifoData[695] or ofifoData[694] or ofifoData[693] or ofifoData[692] or ofifoData[691]
 or ofifoData[690] or ofifoData[689] or ofifoData[688] or ofifoData[687] or ofifoData[686] or ofifoData[685] or ofifoData[684] or ofifoData[683]
 or ofifoData[682] or ofifoData[681] or ofifoData[680] or ofifoData[679] or ofifoData[678] or ofifoData[677] or ofifoData[676] or ofifoData[675]
 or ofifoData[674] or ofifoData[673] or ofifoData[672] or ofifoData[671] or ofifoData[670] or ofifoData[669] or ofifoData[668] or ofifoData[667]
 or ofifoData[666] or ofifoData[665] or ofifoData[664] or ofifoData[663] or ofifoData[662] or ofifoData[661] or ofifoData[660] or ofifoData[659]
 or ofifoData[658] or ofifoData[657] or ofifoData[656] or ofifoData[655] or ofifoData[654] or ofifoData[653] or ofifoData[652] or ofifoData[651]
 or ofifoData[650] or ofifoData[649] or ofifoData[648] or ofifoData[647] or ofifoData[646] or ofifoData[645] or ofifoData[644] or ofifoData[643]
 or ofifoData[642] or ofifoData[641] or ofifoData[640] or ofifoData[639] or ofifoData[638] or ofifoData[637] or ofifoData[636] or ofifoData[635]
 or ofifoData[634] or ofifoData[633] or ofifoData[632] or ofifoData[631] or ofifoData[630] or ofifoData[629] or ofifoData[628] or ofifoData[627]
 or ofifoData[626] or ofifoData[625] or ofifoData[624] or ofifoData[623] or ofifoData[622] or ofifoData[621] or ofifoData[620] or ofifoData[619]
 or ofifoData[618] or ofifoData[617] or ofifoData[616] or ofifoData[615] or ofifoData[614] or ofifoData[613] or ofifoData[612] or ofifoData[611]
 or ofifoData[610] or ofifoData[609] or ofifoData[608] or ofifoData[607] or ofifoData[606] or ofifoData[605] or ofifoData[604] or ofifoData[603]
 or ofifoData[602] or ofifoData[601] or ofifoData[600] or ofifoData[599] or ofifoData[598] or ofifoData[597] or ofifoData[596] or ofifoData[595]
 or ofifoData[594] or ofifoData[593] or ofifoData[592] or ofifoData[591] or ofifoData[590] or ofifoData[589] or ofifoData[588] or ofifoData[587]
 or ofifoData[586] or ofifoData[585] or ofifoData[584] or ofifoData[583] or ofifoData[582] or ofifoData[581] or ofifoData[580] or ofifoData[579]
 or ofifoData[578] or ofifoData[577] or ofifoData[576] or ofifoData[575] or ofifoData[574] or ofifoData[573] or ofifoData[572] or ofifoData[571]
 or ofifoData[570] or ofifoData[569] or ofifoData[568] or ofifoData[567] or ofifoData[566] or ofifoData[565] or ofifoData[564] or ofifoData[563]
 or ofifoData[562] or ofifoData[561] or ofifoData[560] or ofifoData[559] or ofifoData[558] or ofifoData[557] or ofifoData[556] or ofifoData[555]
 or ofifoData[554] or ofifoData[553] or ofifoData[552] or ofifoData[551] or ofifoData[550] or ofifoData[549] or ofifoData[548] or ofifoData[547]
 or ofifoData[546] or ofifoData[545] or ofifoData[544] or ofifoData[543] or ofifoData[542] or ofifoData[541] or ofifoData[540] or ofifoData[539]
 or ofifoData[538] or ofifoData[537] or ofifoData[536] or ofifoData[535] or ofifoData[534] or ofifoData[533] or ofifoData[532] or ofifoData[531]
 or ofifoData[530] or ofifoData[529] or ofifoData[528] or ofifoData[527] or ofifoData[526] or ofifoData[525] or ofifoData[524] or ofifoData[523]
 or ofifoData[522] or ofifoData[521] or ofifoData[520] or ofifoData[519] or ofifoData[518] or ofifoData[517] or ofifoData[516] or ofifoData[515]
 or ofifoData[514] or ofifoData[513] or ofifoData[512] or n5633)
#0 begin
if (n6882)
ixc_gfm_ofifo[{n5631, n5631, n5631, n5631, n5631,
 n5631, n5631, n5631, n5631, n5631, n5631, n5631, n5631,
 n5631, n5631}] =
{oMark[255], oMark[254], oMark[253], oMark[252], oMark[251],
 oMark[250], oMark[249], oMark[248], oMark[247], oMark[246], oMark[245], oMark[244], oMark[243],
 oMark[242], oMark[241], oMark[240], oMark[239], oMark[238], oMark[237], oMark[236], oMark[235],
 oMark[234], oMark[233], oMark[232], oMark[231], oMark[230], oMark[229], oMark[228], oMark[227],
 oMark[226], oMark[225], oMark[224], oMark[223], oMark[222], oMark[221], oMark[220], oMark[219],
 oMark[218], oMark[217], oMark[216], oMark[215], oMark[214], oMark[213], oMark[212], oMark[211],
 oMark[210], oMark[209], oMark[208], oMark[207], oMark[206], oMark[205], oMark[204], oMark[203],
 oMark[202], oMark[201], oMark[200], oMark[199], oMark[198], oMark[197], oMark[196], oMark[195],
 oMark[194], oMark[193], oMark[192], oMark[191], oMark[190], oMark[189], oMark[188], oMark[187],
 oMark[186], oMark[185], oMark[184], oMark[183], oMark[182], oMark[181], oMark[180], oMark[179],
 oMark[178], oMark[177], oMark[176], oMark[175], oMark[174], oMark[173], oMark[172], oMark[171],
 oMark[170], oMark[169], oMark[168], oMark[167], oMark[166], oMark[165], oMark[164], oMark[163],
 oMark[162], oMark[161], oMark[160], oMark[159], oMark[158], oMark[157], oMark[156], oMark[155],
 oMark[154], oMark[153], oMark[152], oMark[151], oMark[150], oMark[149], oMark[148], oMark[147],
 oMark[146], oMark[145], oMark[144], oMark[143], oMark[142], oMark[141], oMark[140], oMark[139],
 oMark[138], oMark[137], oMark[136], oMark[135], oMark[134], oMark[133], oMark[132], oMark[131],
 oMark[130], oMark[129], oMark[128], oMark[127], oMark[126], oMark[125], oMark[124], oMark[123],
 oMark[122], oMark[121], oMark[120], oMark[119], oMark[118], oMark[117], oMark[116], oMark[115],
 oMark[114], oMark[113], oMark[112], oMark[111], oMark[110], oMark[109], oMark[108], oMark[107],
 oMark[106], oMark[105], oMark[104], oMark[103], oMark[102], oMark[101], oMark[100], oMark[99],
 oMark[98], oMark[97], oMark[96], oMark[95], oMark[94], oMark[93], oMark[92], oMark[91],
 oMark[90], oMark[89], oMark[88], oMark[87], oMark[86], oMark[85], oMark[84], oMark[83],
 oMark[82], oMark[81], oMark[80], oMark[79], oMark[78], oMark[77], oMark[76], oMark[75],
 oMark[74], oMark[73], oMark[72], oMark[71], oMark[70], oMark[69], oMark[68], oMark[67],
 oMark[66], oMark[65], oMark[64], oMark[63], oMark[62], oMark[61], oMark[60], oMark[59],
 oMark[58], oMark[57], oMark[56], oMark[55], oMark[54], oMark[53], oMark[52], oMark[51],
 oMark[50], oMark[49], oMark[48], oMark[47], oMark[46], oMark[45], oMark[44], oMark[43],
 oMark[42], oMark[41], oMark[40], oMark[39], oMark[38], oMark[37], oMark[36], oMark[35],
 oMark[34], oMark[33], oMark[32], oMark[31], oMark[30], oMark[29], oMark[28], oMark[27],
 oMark[26], oMark[25], oMark[24], oMark[23], oMark[22], oMark[21], oMark[20], oMark[19],
 oMark[18], oMark[17], oMark[16], oMark[15], oMark[14], oMark[13], oMark[12], oMark[11],
 oMark[10], oMark[9], oMark[8], oMark[7], oMark[6], oMark[5], oMark[4], oMark[3],
 oMark[2], oMark[1], oMark[0]};
if (n6882)
ixc_gfm_ofifo[{ofifoAddr0[14], ofifoAddr0[13], ofifoAddr0[12], ofifoAddr0[11], ofifoAddr0[10],
 ofifoAddr0[9], ofifoAddr0[8], ofifoAddr0[7], ofifoAddr0[6], ofifoAddr0[5], ofifoAddr0[4], ofifoAddr0[3], ofifoAddr0[2],
 ofifoAddr0[1], ofifoAddr0[0]}] =
{ofifoData[255], ofifoData[254], ofifoData[253], ofifoData[252], ofifoData[251],
 ofifoData[250], ofifoData[249], ofifoData[248], ofifoData[247], ofifoData[246], ofifoData[245], ofifoData[244], ofifoData[243],
 ofifoData[242], ofifoData[241], ofifoData[240], ofifoData[239], ofifoData[238], ofifoData[237], ofifoData[236], ofifoData[235],
 ofifoData[234], ofifoData[233], ofifoData[232], ofifoData[231], ofifoData[230], ofifoData[229], ofifoData[228], ofifoData[227],
 ofifoData[226], ofifoData[225], ofifoData[224], ofifoData[223], ofifoData[222], ofifoData[221], ofifoData[220], ofifoData[219],
 ofifoData[218], ofifoData[217], ofifoData[216], ofifoData[215], ofifoData[214], ofifoData[213], ofifoData[212], ofifoData[211],
 ofifoData[210], ofifoData[209], ofifoData[208], ofifoData[207], ofifoData[206], ofifoData[205], ofifoData[204], ofifoData[203],
 ofifoData[202], ofifoData[201], ofifoData[200], ofifoData[199], ofifoData[198], ofifoData[197], ofifoData[196], ofifoData[195],
 ofifoData[194], ofifoData[193], ofifoData[192], ofifoData[191], ofifoData[190], ofifoData[189], ofifoData[188], ofifoData[187],
 ofifoData[186], ofifoData[185], ofifoData[184], ofifoData[183], ofifoData[182], ofifoData[181], ofifoData[180], ofifoData[179],
 ofifoData[178], ofifoData[177], ofifoData[176], ofifoData[175], ofifoData[174], ofifoData[173], ofifoData[172], ofifoData[171],
 ofifoData[170], ofifoData[169], ofifoData[168], ofifoData[167], ofifoData[166], ofifoData[165], ofifoData[164], ofifoData[163],
 ofifoData[162], ofifoData[161], ofifoData[160], ofifoData[159], ofifoData[158], ofifoData[157], ofifoData[156], ofifoData[155],
 ofifoData[154], ofifoData[153], ofifoData[152], ofifoData[151], ofifoData[150], ofifoData[149], ofifoData[148], ofifoData[147],
 ofifoData[146], ofifoData[145], ofifoData[144], ofifoData[143], ofifoData[142], ofifoData[141], ofifoData[140], ofifoData[139],
 ofifoData[138], ofifoData[137], ofifoData[136], ofifoData[135], ofifoData[134], ofifoData[133], ofifoData[132], ofifoData[131],
 ofifoData[130], ofifoData[129], ofifoData[128], ofifoData[127], ofifoData[126], ofifoData[125], ofifoData[124], ofifoData[123],
 ofifoData[122], ofifoData[121], ofifoData[120], ofifoData[119], ofifoData[118], ofifoData[117], ofifoData[116], ofifoData[115],
 ofifoData[114], ofifoData[113], ofifoData[112], ofifoData[111], ofifoData[110], ofifoData[109], ofifoData[108], ofifoData[107],
 ofifoData[106], ofifoData[105], ofifoData[104], ofifoData[103], ofifoData[102], ofifoData[101], ofifoData[100], ofifoData[99],
 ofifoData[98], ofifoData[97], ofifoData[96], ofifoData[95], ofifoData[94], ofifoData[93], ofifoData[92], ofifoData[91],
 ofifoData[90], ofifoData[89], ofifoData[88], ofifoData[87], ofifoData[86], ofifoData[85], ofifoData[84], ofifoData[83],
 ofifoData[82], ofifoData[81], ofifoData[80], ofifoData[79], ofifoData[78], ofifoData[77], ofifoData[76], ofifoData[75],
 ofifoData[74], ofifoData[73], ofifoData[72], ofifoData[71], ofifoData[70], ofifoData[69], ofifoData[68], ofifoData[67],
 ofifoData[66], ofifoData[65], ofifoData[64], ofifoData[63], ofifoData[62], ofifoData[61], ofifoData[60], ofifoData[59],
 ofifoData[58], ofifoData[57], ofifoData[56], ofifoData[55], ofifoData[54], ofifoData[53], ofifoData[52], ofifoData[51],
 ofifoData[50], ofifoData[49], ofifoData[48], ofifoData[47], ofifoData[46], ofifoData[45], ofifoData[44], ofifoData[43],
 ofifoData[42], ofifoData[41], ofifoData[40], ofifoData[39], ofifoData[38], ofifoData[37], ofifoData[36], ofifoData[35],
 ofifoData[34], ofifoData[33], ofifoData[32], ofifoData[31], ofifoData[30], ofifoData[29], ofifoData[28], ofifoData[27],
 ofifoData[26], ofifoData[25], ofifoData[24], ofifoData[23], ofifoData[22], ofifoData[21], ofifoData[20], ofifoData[19],
 ofifoData[18], ofifoData[17], ofifoData[16], ofifoData[15], ofifoData[14], ofifoData[13], ofifoData[12], ofifoData[11],
 ofifoData[10], ofifoData[9], ofifoData[8], ofifoData[7], ofifoData[6], ofifoData[5], ofifoData[4], ofifoData[3],
 ofifoData[2], ofifoData[1], ofifoData[0]};
if (n5632)
ixc_gfm_ofifo[{ofifoAddr1[14], ofifoAddr1[13], ofifoAddr1[12], ofifoAddr1[11], ofifoAddr1[10],
 ofifoAddr1[9], ofifoAddr1[8], ofifoAddr1[7], ofifoAddr1[6], ofifoAddr1[5], ofifoAddr1[4], ofifoAddr1[3], ofifoAddr1[2],
 ofifoAddr1[1], ofifoAddr1[0]}] =
{ofifoData[511], ofifoData[510], ofifoData[509], ofifoData[508], ofifoData[507],
 ofifoData[506], ofifoData[505], ofifoData[504], ofifoData[503], ofifoData[502], ofifoData[501], ofifoData[500], ofifoData[499],
 ofifoData[498], ofifoData[497], ofifoData[496], ofifoData[495], ofifoData[494], ofifoData[493], ofifoData[492], ofifoData[491],
 ofifoData[490], ofifoData[489], ofifoData[488], ofifoData[487], ofifoData[486], ofifoData[485], ofifoData[484], ofifoData[483],
 ofifoData[482], ofifoData[481], ofifoData[480], ofifoData[479], ofifoData[478], ofifoData[477], ofifoData[476], ofifoData[475],
 ofifoData[474], ofifoData[473], ofifoData[472], ofifoData[471], ofifoData[470], ofifoData[469], ofifoData[468], ofifoData[467],
 ofifoData[466], ofifoData[465], ofifoData[464], ofifoData[463], ofifoData[462], ofifoData[461], ofifoData[460], ofifoData[459],
 ofifoData[458], ofifoData[457], ofifoData[456], ofifoData[455], ofifoData[454], ofifoData[453], ofifoData[452], ofifoData[451],
 ofifoData[450], ofifoData[449], ofifoData[448], ofifoData[447], ofifoData[446], ofifoData[445], ofifoData[444], ofifoData[443],
 ofifoData[442], ofifoData[441], ofifoData[440], ofifoData[439], ofifoData[438], ofifoData[437], ofifoData[436], ofifoData[435],
 ofifoData[434], ofifoData[433], ofifoData[432], ofifoData[431], ofifoData[430], ofifoData[429], ofifoData[428], ofifoData[427],
 ofifoData[426], ofifoData[425], ofifoData[424], ofifoData[423], ofifoData[422], ofifoData[421], ofifoData[420], ofifoData[419],
 ofifoData[418], ofifoData[417], ofifoData[416], ofifoData[415], ofifoData[414], ofifoData[413], ofifoData[412], ofifoData[411],
 ofifoData[410], ofifoData[409], ofifoData[408], ofifoData[407], ofifoData[406], ofifoData[405], ofifoData[404], ofifoData[403],
 ofifoData[402], ofifoData[401], ofifoData[400], ofifoData[399], ofifoData[398], ofifoData[397], ofifoData[396], ofifoData[395],
 ofifoData[394], ofifoData[393], ofifoData[392], ofifoData[391], ofifoData[390], ofifoData[389], ofifoData[388], ofifoData[387],
 ofifoData[386], ofifoData[385], ofifoData[384], ofifoData[383], ofifoData[382], ofifoData[381], ofifoData[380], ofifoData[379],
 ofifoData[378], ofifoData[377], ofifoData[376], ofifoData[375], ofifoData[374], ofifoData[373], ofifoData[372], ofifoData[371],
 ofifoData[370], ofifoData[369], ofifoData[368], ofifoData[367], ofifoData[366], ofifoData[365], ofifoData[364], ofifoData[363],
 ofifoData[362], ofifoData[361], ofifoData[360], ofifoData[359], ofifoData[358], ofifoData[357], ofifoData[356], ofifoData[355],
 ofifoData[354], ofifoData[353], ofifoData[352], ofifoData[351], ofifoData[350], ofifoData[349], ofifoData[348], ofifoData[347],
 ofifoData[346], ofifoData[345], ofifoData[344], ofifoData[343], ofifoData[342], ofifoData[341], ofifoData[340], ofifoData[339],
 ofifoData[338], ofifoData[337], ofifoData[336], ofifoData[335], ofifoData[334], ofifoData[333], ofifoData[332], ofifoData[331],
 ofifoData[330], ofifoData[329], ofifoData[328], ofifoData[327], ofifoData[326], ofifoData[325], ofifoData[324], ofifoData[323],
 ofifoData[322], ofifoData[321], ofifoData[320], ofifoData[319], ofifoData[318], ofifoData[317], ofifoData[316], ofifoData[315],
 ofifoData[314], ofifoData[313], ofifoData[312], ofifoData[311], ofifoData[310], ofifoData[309], ofifoData[308], ofifoData[307],
 ofifoData[306], ofifoData[305], ofifoData[304], ofifoData[303], ofifoData[302], ofifoData[301], ofifoData[300], ofifoData[299],
 ofifoData[298], ofifoData[297], ofifoData[296], ofifoData[295], ofifoData[294], ofifoData[293], ofifoData[292], ofifoData[291],
 ofifoData[290], ofifoData[289], ofifoData[288], ofifoData[287], ofifoData[286], ofifoData[285], ofifoData[284], ofifoData[283],
 ofifoData[282], ofifoData[281], ofifoData[280], ofifoData[279], ofifoData[278], ofifoData[277], ofifoData[276], ofifoData[275],
 ofifoData[274], ofifoData[273], ofifoData[272], ofifoData[271], ofifoData[270], ofifoData[269], ofifoData[268], ofifoData[267],
 ofifoData[266], ofifoData[265], ofifoData[264], ofifoData[263], ofifoData[262], ofifoData[261], ofifoData[260], ofifoData[259],
 ofifoData[258], ofifoData[257], ofifoData[256]};
if (n5633)
ixc_gfm_ofifo[{ofifoAddr2[14], ofifoAddr2[13], ofifoAddr2[12], ofifoAddr2[11], ofifoAddr2[10],
 ofifoAddr2[9], ofifoAddr2[8], ofifoAddr2[7], ofifoAddr2[6], ofifoAddr2[5], ofifoAddr2[4], ofifoAddr2[3], ofifoAddr2[2],
 ofifoAddr2[1], ofifoAddr2[0]}] =
{ofifoData[767], ofifoData[766], ofifoData[765], ofifoData[764], ofifoData[763],
 ofifoData[762], ofifoData[761], ofifoData[760], ofifoData[759], ofifoData[758], ofifoData[757], ofifoData[756], ofifoData[755],
 ofifoData[754], ofifoData[753], ofifoData[752], ofifoData[751], ofifoData[750], ofifoData[749], ofifoData[748], ofifoData[747],
 ofifoData[746], ofifoData[745], ofifoData[744], ofifoData[743], ofifoData[742], ofifoData[741], ofifoData[740], ofifoData[739],
 ofifoData[738], ofifoData[737], ofifoData[736], ofifoData[735], ofifoData[734], ofifoData[733], ofifoData[732], ofifoData[731],
 ofifoData[730], ofifoData[729], ofifoData[728], ofifoData[727], ofifoData[726], ofifoData[725], ofifoData[724], ofifoData[723],
 ofifoData[722], ofifoData[721], ofifoData[720], ofifoData[719], ofifoData[718], ofifoData[717], ofifoData[716], ofifoData[715],
 ofifoData[714], ofifoData[713], ofifoData[712], ofifoData[711], ofifoData[710], ofifoData[709], ofifoData[708], ofifoData[707],
 ofifoData[706], ofifoData[705], ofifoData[704], ofifoData[703], ofifoData[702], ofifoData[701], ofifoData[700], ofifoData[699],
 ofifoData[698], ofifoData[697], ofifoData[696], ofifoData[695], ofifoData[694], ofifoData[693], ofifoData[692], ofifoData[691],
 ofifoData[690], ofifoData[689], ofifoData[688], ofifoData[687], ofifoData[686], ofifoData[685], ofifoData[684], ofifoData[683],
 ofifoData[682], ofifoData[681], ofifoData[680], ofifoData[679], ofifoData[678], ofifoData[677], ofifoData[676], ofifoData[675],
 ofifoData[674], ofifoData[673], ofifoData[672], ofifoData[671], ofifoData[670], ofifoData[669], ofifoData[668], ofifoData[667],
 ofifoData[666], ofifoData[665], ofifoData[664], ofifoData[663], ofifoData[662], ofifoData[661], ofifoData[660], ofifoData[659],
 ofifoData[658], ofifoData[657], ofifoData[656], ofifoData[655], ofifoData[654], ofifoData[653], ofifoData[652], ofifoData[651],
 ofifoData[650], ofifoData[649], ofifoData[648], ofifoData[647], ofifoData[646], ofifoData[645], ofifoData[644], ofifoData[643],
 ofifoData[642], ofifoData[641], ofifoData[640], ofifoData[639], ofifoData[638], ofifoData[637], ofifoData[636], ofifoData[635],
 ofifoData[634], ofifoData[633], ofifoData[632], ofifoData[631], ofifoData[630], ofifoData[629], ofifoData[628], ofifoData[627],
 ofifoData[626], ofifoData[625], ofifoData[624], ofifoData[623], ofifoData[622], ofifoData[621], ofifoData[620], ofifoData[619],
 ofifoData[618], ofifoData[617], ofifoData[616], ofifoData[615], ofifoData[614], ofifoData[613], ofifoData[612], ofifoData[611],
 ofifoData[610], ofifoData[609], ofifoData[608], ofifoData[607], ofifoData[606], ofifoData[605], ofifoData[604], ofifoData[603],
 ofifoData[602], ofifoData[601], ofifoData[600], ofifoData[599], ofifoData[598], ofifoData[597], ofifoData[596], ofifoData[595],
 ofifoData[594], ofifoData[593], ofifoData[592], ofifoData[591], ofifoData[590], ofifoData[589], ofifoData[588], ofifoData[587],
 ofifoData[586], ofifoData[585], ofifoData[584], ofifoData[583], ofifoData[582], ofifoData[581], ofifoData[580], ofifoData[579],
 ofifoData[578], ofifoData[577], ofifoData[576], ofifoData[575], ofifoData[574], ofifoData[573], ofifoData[572], ofifoData[571],
 ofifoData[570], ofifoData[569], ofifoData[568], ofifoData[567], ofifoData[566], ofifoData[565], ofifoData[564], ofifoData[563],
 ofifoData[562], ofifoData[561], ofifoData[560], ofifoData[559], ofifoData[558], ofifoData[557], ofifoData[556], ofifoData[555],
 ofifoData[554], ofifoData[553], ofifoData[552], ofifoData[551], ofifoData[550], ofifoData[549], ofifoData[548], ofifoData[547],
 ofifoData[546], ofifoData[545], ofifoData[544], ofifoData[543], ofifoData[542], ofifoData[541], ofifoData[540], ofifoData[539],
 ofifoData[538], ofifoData[537], ofifoData[536], ofifoData[535], ofifoData[534], ofifoData[533], ofifoData[532], ofifoData[531],
 ofifoData[530], ofifoData[529], ofifoData[528], ofifoData[527], ofifoData[526], ofifoData[525], ofifoData[524], ofifoData[523],
 ofifoData[522], ofifoData[521], ofifoData[520], ofifoData[519], ofifoData[518], ofifoData[517], ofifoData[516], ofifoData[515],
 ofifoData[514], ofifoData[513], ofifoData[512]};
end
`else

MPW32KX256 ixc_gfm_ofifo ( .A14(n5631), .A13(n5631), .A12(n5631), .A11(n5631), .A10(n5631), .A9(n5631),
 .A8(n5631), .A7(n5631), .A6(n5631), .A5(n5631), .A4(n5631), .A3(n5631), .A2(n5631), .A1(n5631),
 .A0(n5631), .DI255(oMark[255]), .DI254(oMark[254]), .DI253(oMark[253]), .DI252(oMark[252]), .DI251(oMark[251]), .DI250(oMark[250]), .DI249(oMark[249]),
 .DI248(oMark[248]), .DI247(oMark[247]), .DI246(oMark[246]), .DI245(oMark[245]), .DI244(oMark[244]), .DI243(oMark[243]), .DI242(oMark[242]), .DI241(oMark[241]),
 .DI240(oMark[240]), .DI239(oMark[239]), .DI238(oMark[238]), .DI237(oMark[237]), .DI236(oMark[236]), .DI235(oMark[235]), .DI234(oMark[234]), .DI233(oMark[233]),
 .DI232(oMark[232]), .DI231(oMark[231]), .DI230(oMark[230]), .DI229(oMark[229]), .DI228(oMark[228]), .DI227(oMark[227]), .DI226(oMark[226]), .DI225(oMark[225]),
 .DI224(oMark[224]), .DI223(oMark[223]), .DI222(oMark[222]), .DI221(oMark[221]), .DI220(oMark[220]), .DI219(oMark[219]), .DI218(oMark[218]), .DI217(oMark[217]),
 .DI216(oMark[216]), .DI215(oMark[215]), .DI214(oMark[214]), .DI213(oMark[213]), .DI212(oMark[212]), .DI211(oMark[211]), .DI210(oMark[210]), .DI209(oMark[209]),
 .DI208(oMark[208]), .DI207(oMark[207]), .DI206(oMark[206]), .DI205(oMark[205]), .DI204(oMark[204]), .DI203(oMark[203]), .DI202(oMark[202]), .DI201(oMark[201]),
 .DI200(oMark[200]), .DI199(oMark[199]), .DI198(oMark[198]), .DI197(oMark[197]), .DI196(oMark[196]), .DI195(oMark[195]), .DI194(oMark[194]), .DI193(oMark[193]),
 .DI192(oMark[192]), .DI191(oMark[191]), .DI190(oMark[190]), .DI189(oMark[189]), .DI188(oMark[188]), .DI187(oMark[187]), .DI186(oMark[186]), .DI185(oMark[185]),
 .DI184(oMark[184]), .DI183(oMark[183]), .DI182(oMark[182]), .DI181(oMark[181]), .DI180(oMark[180]), .DI179(oMark[179]), .DI178(oMark[178]), .DI177(oMark[177]),
 .DI176(oMark[176]), .DI175(oMark[175]), .DI174(oMark[174]), .DI173(oMark[173]), .DI172(oMark[172]), .DI171(oMark[171]), .DI170(oMark[170]), .DI169(oMark[169]),
 .DI168(oMark[168]), .DI167(oMark[167]), .DI166(oMark[166]), .DI165(oMark[165]), .DI164(oMark[164]), .DI163(oMark[163]), .DI162(oMark[162]), .DI161(oMark[161]),
 .DI160(oMark[160]), .DI159(oMark[159]), .DI158(oMark[158]), .DI157(oMark[157]), .DI156(oMark[156]), .DI155(oMark[155]), .DI154(oMark[154]), .DI153(oMark[153]),
 .DI152(oMark[152]), .DI151(oMark[151]), .DI150(oMark[150]), .DI149(oMark[149]), .DI148(oMark[148]), .DI147(oMark[147]), .DI146(oMark[146]), .DI145(oMark[145]),
 .DI144(oMark[144]), .DI143(oMark[143]), .DI142(oMark[142]), .DI141(oMark[141]), .DI140(oMark[140]), .DI139(oMark[139]), .DI138(oMark[138]), .DI137(oMark[137]),
 .DI136(oMark[136]), .DI135(oMark[135]), .DI134(oMark[134]), .DI133(oMark[133]), .DI132(oMark[132]), .DI131(oMark[131]), .DI130(oMark[130]), .DI129(oMark[129]),
 .DI128(oMark[128]), .DI127(oMark[127]), .DI126(oMark[126]), .DI125(oMark[125]), .DI124(oMark[124]), .DI123(oMark[123]), .DI122(oMark[122]), .DI121(oMark[121]),
 .DI120(oMark[120]), .DI119(oMark[119]), .DI118(oMark[118]), .DI117(oMark[117]), .DI116(oMark[116]), .DI115(oMark[115]), .DI114(oMark[114]), .DI113(oMark[113]),
 .DI112(oMark[112]), .DI111(oMark[111]), .DI110(oMark[110]), .DI109(oMark[109]), .DI108(oMark[108]), .DI107(oMark[107]), .DI106(oMark[106]), .DI105(oMark[105]),
 .DI104(oMark[104]), .DI103(oMark[103]), .DI102(oMark[102]), .DI101(oMark[101]), .DI100(oMark[100]), .DI99(oMark[99]), .DI98(oMark[98]), .DI97(oMark[97]),
 .DI96(oMark[96]), .DI95(oMark[95]), .DI94(oMark[94]), .DI93(oMark[93]), .DI92(oMark[92]), .DI91(oMark[91]), .DI90(oMark[90]), .DI89(oMark[89]),
 .DI88(oMark[88]), .DI87(oMark[87]), .DI86(oMark[86]), .DI85(oMark[85]), .DI84(oMark[84]), .DI83(oMark[83]), .DI82(oMark[82]), .DI81(oMark[81]),
 .DI80(oMark[80]), .DI79(oMark[79]), .DI78(oMark[78]), .DI77(oMark[77]), .DI76(oMark[76]), .DI75(oMark[75]), .DI74(oMark[74]), .DI73(oMark[73]),
 .DI72(oMark[72]), .DI71(oMark[71]), .DI70(oMark[70]), .DI69(oMark[69]), .DI68(oMark[68]), .DI67(oMark[67]), .DI66(oMark[66]), .DI65(oMark[65]),
 .DI64(oMark[64]), .DI63(oMark[63]), .DI62(oMark[62]), .DI61(oMark[61]), .DI60(oMark[60]), .DI59(oMark[59]), .DI58(oMark[58]), .DI57(oMark[57]),
 .DI56(oMark[56]), .DI55(oMark[55]), .DI54(oMark[54]), .DI53(oMark[53]), .DI52(oMark[52]), .DI51(oMark[51]), .DI50(oMark[50]), .DI49(oMark[49]),
 .DI48(oMark[48]), .DI47(oMark[47]), .DI46(oMark[46]), .DI45(oMark[45]), .DI44(oMark[44]), .DI43(oMark[43]), .DI42(oMark[42]), .DI41(oMark[41]),
 .DI40(oMark[40]), .DI39(oMark[39]), .DI38(oMark[38]), .DI37(oMark[37]), .DI36(oMark[36]), .DI35(oMark[35]), .DI34(oMark[34]), .DI33(oMark[33]),
 .DI32(oMark[32]), .DI31(oMark[31]), .DI30(oMark[30]), .DI29(oMark[29]), .DI28(oMark[28]), .DI27(oMark[27]), .DI26(oMark[26]), .DI25(oMark[25]),
 .DI24(oMark[24]), .DI23(oMark[23]), .DI22(oMark[22]), .DI21(oMark[21]), .DI20(oMark[20]), .DI19(oMark[19]), .DI18(oMark[18]), .DI17(oMark[17]),
 .DI16(oMark[16]), .DI15(oMark[15]), .DI14(oMark[14]), .DI13(oMark[13]), .DI12(oMark[12]), .DI11(oMark[11]), .DI10(oMark[10]), .DI9(oMark[9]),
 .DI8(oMark[8]), .DI7(oMark[7]), .DI6(oMark[6]), .DI5(oMark[5]), .DI4(oMark[4]), .DI3(oMark[3]), .DI2(oMark[2]), .DI1(oMark[1]),
 .DI0(oMark[0]), .WE(n6882), .SYNC_IN(n5631), .SYNC_OUT(n9333));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ofifo" HDL_MEMORY_DECL "1 255 0 0 32767"
MPW32KX256 U10459 ( .A14(ofifoAddr0[14]), .A13(ofifoAddr0[13]), .A12(ofifoAddr0[12]), .A11(ofifoAddr0[11]), .A10(ofifoAddr0[10]), .A9(ofifoAddr0[9]),
 .A8(ofifoAddr0[8]), .A7(ofifoAddr0[7]), .A6(ofifoAddr0[6]), .A5(ofifoAddr0[5]), .A4(ofifoAddr0[4]), .A3(ofifoAddr0[3]), .A2(ofifoAddr0[2]), .A1(ofifoAddr0[1]),
 .A0(ofifoAddr0[0]), .DI255(ofifoData[255]), .DI254(ofifoData[254]), .DI253(ofifoData[253]), .DI252(ofifoData[252]), .DI251(ofifoData[251]), .DI250(ofifoData[250]), .DI249(ofifoData[249]),
 .DI248(ofifoData[248]), .DI247(ofifoData[247]), .DI246(ofifoData[246]), .DI245(ofifoData[245]), .DI244(ofifoData[244]), .DI243(ofifoData[243]), .DI242(ofifoData[242]), .DI241(ofifoData[241]),
 .DI240(ofifoData[240]), .DI239(ofifoData[239]), .DI238(ofifoData[238]), .DI237(ofifoData[237]), .DI236(ofifoData[236]), .DI235(ofifoData[235]), .DI234(ofifoData[234]), .DI233(ofifoData[233]),
 .DI232(ofifoData[232]), .DI231(ofifoData[231]), .DI230(ofifoData[230]), .DI229(ofifoData[229]), .DI228(ofifoData[228]), .DI227(ofifoData[227]), .DI226(ofifoData[226]), .DI225(ofifoData[225]),
 .DI224(ofifoData[224]), .DI223(ofifoData[223]), .DI222(ofifoData[222]), .DI221(ofifoData[221]), .DI220(ofifoData[220]), .DI219(ofifoData[219]), .DI218(ofifoData[218]), .DI217(ofifoData[217]),
 .DI216(ofifoData[216]), .DI215(ofifoData[215]), .DI214(ofifoData[214]), .DI213(ofifoData[213]), .DI212(ofifoData[212]), .DI211(ofifoData[211]), .DI210(ofifoData[210]), .DI209(ofifoData[209]),
 .DI208(ofifoData[208]), .DI207(ofifoData[207]), .DI206(ofifoData[206]), .DI205(ofifoData[205]), .DI204(ofifoData[204]), .DI203(ofifoData[203]), .DI202(ofifoData[202]), .DI201(ofifoData[201]),
 .DI200(ofifoData[200]), .DI199(ofifoData[199]), .DI198(ofifoData[198]), .DI197(ofifoData[197]), .DI196(ofifoData[196]), .DI195(ofifoData[195]), .DI194(ofifoData[194]), .DI193(ofifoData[193]),
 .DI192(ofifoData[192]), .DI191(ofifoData[191]), .DI190(ofifoData[190]), .DI189(ofifoData[189]), .DI188(ofifoData[188]), .DI187(ofifoData[187]), .DI186(ofifoData[186]), .DI185(ofifoData[185]),
 .DI184(ofifoData[184]), .DI183(ofifoData[183]), .DI182(ofifoData[182]), .DI181(ofifoData[181]), .DI180(ofifoData[180]), .DI179(ofifoData[179]), .DI178(ofifoData[178]), .DI177(ofifoData[177]),
 .DI176(ofifoData[176]), .DI175(ofifoData[175]), .DI174(ofifoData[174]), .DI173(ofifoData[173]), .DI172(ofifoData[172]), .DI171(ofifoData[171]), .DI170(ofifoData[170]), .DI169(ofifoData[169]),
 .DI168(ofifoData[168]), .DI167(ofifoData[167]), .DI166(ofifoData[166]), .DI165(ofifoData[165]), .DI164(ofifoData[164]), .DI163(ofifoData[163]), .DI162(ofifoData[162]), .DI161(ofifoData[161]),
 .DI160(ofifoData[160]), .DI159(ofifoData[159]), .DI158(ofifoData[158]), .DI157(ofifoData[157]), .DI156(ofifoData[156]), .DI155(ofifoData[155]), .DI154(ofifoData[154]), .DI153(ofifoData[153]),
 .DI152(ofifoData[152]), .DI151(ofifoData[151]), .DI150(ofifoData[150]), .DI149(ofifoData[149]), .DI148(ofifoData[148]), .DI147(ofifoData[147]), .DI146(ofifoData[146]), .DI145(ofifoData[145]),
 .DI144(ofifoData[144]), .DI143(ofifoData[143]), .DI142(ofifoData[142]), .DI141(ofifoData[141]), .DI140(ofifoData[140]), .DI139(ofifoData[139]), .DI138(ofifoData[138]), .DI137(ofifoData[137]),
 .DI136(ofifoData[136]), .DI135(ofifoData[135]), .DI134(ofifoData[134]), .DI133(ofifoData[133]), .DI132(ofifoData[132]), .DI131(ofifoData[131]), .DI130(ofifoData[130]), .DI129(ofifoData[129]),
 .DI128(ofifoData[128]), .DI127(ofifoData[127]), .DI126(ofifoData[126]), .DI125(ofifoData[125]), .DI124(ofifoData[124]), .DI123(ofifoData[123]), .DI122(ofifoData[122]), .DI121(ofifoData[121]),
 .DI120(ofifoData[120]), .DI119(ofifoData[119]), .DI118(ofifoData[118]), .DI117(ofifoData[117]), .DI116(ofifoData[116]), .DI115(ofifoData[115]), .DI114(ofifoData[114]), .DI113(ofifoData[113]),
 .DI112(ofifoData[112]), .DI111(ofifoData[111]), .DI110(ofifoData[110]), .DI109(ofifoData[109]), .DI108(ofifoData[108]), .DI107(ofifoData[107]), .DI106(ofifoData[106]), .DI105(ofifoData[105]),
 .DI104(ofifoData[104]), .DI103(ofifoData[103]), .DI102(ofifoData[102]), .DI101(ofifoData[101]), .DI100(ofifoData[100]), .DI99(ofifoData[99]), .DI98(ofifoData[98]), .DI97(ofifoData[97]),
 .DI96(ofifoData[96]), .DI95(ofifoData[95]), .DI94(ofifoData[94]), .DI93(ofifoData[93]), .DI92(ofifoData[92]), .DI91(ofifoData[91]), .DI90(ofifoData[90]), .DI89(ofifoData[89]),
 .DI88(ofifoData[88]), .DI87(ofifoData[87]), .DI86(ofifoData[86]), .DI85(ofifoData[85]), .DI84(ofifoData[84]), .DI83(ofifoData[83]), .DI82(ofifoData[82]), .DI81(ofifoData[81]),
 .DI80(ofifoData[80]), .DI79(ofifoData[79]), .DI78(ofifoData[78]), .DI77(ofifoData[77]), .DI76(ofifoData[76]), .DI75(ofifoData[75]), .DI74(ofifoData[74]), .DI73(ofifoData[73]),
 .DI72(ofifoData[72]), .DI71(ofifoData[71]), .DI70(ofifoData[70]), .DI69(ofifoData[69]), .DI68(ofifoData[68]), .DI67(ofifoData[67]), .DI66(ofifoData[66]), .DI65(ofifoData[65]),
 .DI64(ofifoData[64]), .DI63(ofifoData[63]), .DI62(ofifoData[62]), .DI61(ofifoData[61]), .DI60(ofifoData[60]), .DI59(ofifoData[59]), .DI58(ofifoData[58]), .DI57(ofifoData[57]),
 .DI56(ofifoData[56]), .DI55(ofifoData[55]), .DI54(ofifoData[54]), .DI53(ofifoData[53]), .DI52(ofifoData[52]), .DI51(ofifoData[51]), .DI50(ofifoData[50]), .DI49(ofifoData[49]),
 .DI48(ofifoData[48]), .DI47(ofifoData[47]), .DI46(ofifoData[46]), .DI45(ofifoData[45]), .DI44(ofifoData[44]), .DI43(ofifoData[43]), .DI42(ofifoData[42]), .DI41(ofifoData[41]),
 .DI40(ofifoData[40]), .DI39(ofifoData[39]), .DI38(ofifoData[38]), .DI37(ofifoData[37]), .DI36(ofifoData[36]), .DI35(ofifoData[35]), .DI34(ofifoData[34]), .DI33(ofifoData[33]),
 .DI32(ofifoData[32]), .DI31(ofifoData[31]), .DI30(ofifoData[30]), .DI29(ofifoData[29]), .DI28(ofifoData[28]), .DI27(ofifoData[27]), .DI26(ofifoData[26]), .DI25(ofifoData[25]),
 .DI24(ofifoData[24]), .DI23(ofifoData[23]), .DI22(ofifoData[22]), .DI21(ofifoData[21]), .DI20(ofifoData[20]), .DI19(ofifoData[19]), .DI18(ofifoData[18]), .DI17(ofifoData[17]),
 .DI16(ofifoData[16]), .DI15(ofifoData[15]), .DI14(ofifoData[14]), .DI13(ofifoData[13]), .DI12(ofifoData[12]), .DI11(ofifoData[11]), .DI10(ofifoData[10]), .DI9(ofifoData[9]),
 .DI8(ofifoData[8]), .DI7(ofifoData[7]), .DI6(ofifoData[6]), .DI5(ofifoData[5]), .DI4(ofifoData[4]), .DI3(ofifoData[3]), .DI2(ofifoData[2]), .DI1(ofifoData[1]),
 .DI0(ofifoData[0]), .WE(n6882), .SYNC_IN(n9333), .SYNC_OUT(n9334));
MPW32KX256 U10460 ( .A14(ofifoAddr1[14]), .A13(ofifoAddr1[13]), .A12(ofifoAddr1[12]), .A11(ofifoAddr1[11]), .A10(ofifoAddr1[10]), .A9(ofifoAddr1[9]),
 .A8(ofifoAddr1[8]), .A7(ofifoAddr1[7]), .A6(ofifoAddr1[6]), .A5(ofifoAddr1[5]), .A4(ofifoAddr1[4]), .A3(ofifoAddr1[3]), .A2(ofifoAddr1[2]), .A1(ofifoAddr1[1]),
 .A0(ofifoAddr1[0]), .DI255(ofifoData[511]), .DI254(ofifoData[510]), .DI253(ofifoData[509]), .DI252(ofifoData[508]), .DI251(ofifoData[507]), .DI250(ofifoData[506]), .DI249(ofifoData[505]),
 .DI248(ofifoData[504]), .DI247(ofifoData[503]), .DI246(ofifoData[502]), .DI245(ofifoData[501]), .DI244(ofifoData[500]), .DI243(ofifoData[499]), .DI242(ofifoData[498]), .DI241(ofifoData[497]),
 .DI240(ofifoData[496]), .DI239(ofifoData[495]), .DI238(ofifoData[494]), .DI237(ofifoData[493]), .DI236(ofifoData[492]), .DI235(ofifoData[491]), .DI234(ofifoData[490]), .DI233(ofifoData[489]),
 .DI232(ofifoData[488]), .DI231(ofifoData[487]), .DI230(ofifoData[486]), .DI229(ofifoData[485]), .DI228(ofifoData[484]), .DI227(ofifoData[483]), .DI226(ofifoData[482]), .DI225(ofifoData[481]),
 .DI224(ofifoData[480]), .DI223(ofifoData[479]), .DI222(ofifoData[478]), .DI221(ofifoData[477]), .DI220(ofifoData[476]), .DI219(ofifoData[475]), .DI218(ofifoData[474]), .DI217(ofifoData[473]),
 .DI216(ofifoData[472]), .DI215(ofifoData[471]), .DI214(ofifoData[470]), .DI213(ofifoData[469]), .DI212(ofifoData[468]), .DI211(ofifoData[467]), .DI210(ofifoData[466]), .DI209(ofifoData[465]),
 .DI208(ofifoData[464]), .DI207(ofifoData[463]), .DI206(ofifoData[462]), .DI205(ofifoData[461]), .DI204(ofifoData[460]), .DI203(ofifoData[459]), .DI202(ofifoData[458]), .DI201(ofifoData[457]),
 .DI200(ofifoData[456]), .DI199(ofifoData[455]), .DI198(ofifoData[454]), .DI197(ofifoData[453]), .DI196(ofifoData[452]), .DI195(ofifoData[451]), .DI194(ofifoData[450]), .DI193(ofifoData[449]),
 .DI192(ofifoData[448]), .DI191(ofifoData[447]), .DI190(ofifoData[446]), .DI189(ofifoData[445]), .DI188(ofifoData[444]), .DI187(ofifoData[443]), .DI186(ofifoData[442]), .DI185(ofifoData[441]),
 .DI184(ofifoData[440]), .DI183(ofifoData[439]), .DI182(ofifoData[438]), .DI181(ofifoData[437]), .DI180(ofifoData[436]), .DI179(ofifoData[435]), .DI178(ofifoData[434]), .DI177(ofifoData[433]),
 .DI176(ofifoData[432]), .DI175(ofifoData[431]), .DI174(ofifoData[430]), .DI173(ofifoData[429]), .DI172(ofifoData[428]), .DI171(ofifoData[427]), .DI170(ofifoData[426]), .DI169(ofifoData[425]),
 .DI168(ofifoData[424]), .DI167(ofifoData[423]), .DI166(ofifoData[422]), .DI165(ofifoData[421]), .DI164(ofifoData[420]), .DI163(ofifoData[419]), .DI162(ofifoData[418]), .DI161(ofifoData[417]),
 .DI160(ofifoData[416]), .DI159(ofifoData[415]), .DI158(ofifoData[414]), .DI157(ofifoData[413]), .DI156(ofifoData[412]), .DI155(ofifoData[411]), .DI154(ofifoData[410]), .DI153(ofifoData[409]),
 .DI152(ofifoData[408]), .DI151(ofifoData[407]), .DI150(ofifoData[406]), .DI149(ofifoData[405]), .DI148(ofifoData[404]), .DI147(ofifoData[403]), .DI146(ofifoData[402]), .DI145(ofifoData[401]),
 .DI144(ofifoData[400]), .DI143(ofifoData[399]), .DI142(ofifoData[398]), .DI141(ofifoData[397]), .DI140(ofifoData[396]), .DI139(ofifoData[395]), .DI138(ofifoData[394]), .DI137(ofifoData[393]),
 .DI136(ofifoData[392]), .DI135(ofifoData[391]), .DI134(ofifoData[390]), .DI133(ofifoData[389]), .DI132(ofifoData[388]), .DI131(ofifoData[387]), .DI130(ofifoData[386]), .DI129(ofifoData[385]),
 .DI128(ofifoData[384]), .DI127(ofifoData[383]), .DI126(ofifoData[382]), .DI125(ofifoData[381]), .DI124(ofifoData[380]), .DI123(ofifoData[379]), .DI122(ofifoData[378]), .DI121(ofifoData[377]),
 .DI120(ofifoData[376]), .DI119(ofifoData[375]), .DI118(ofifoData[374]), .DI117(ofifoData[373]), .DI116(ofifoData[372]), .DI115(ofifoData[371]), .DI114(ofifoData[370]), .DI113(ofifoData[369]),
 .DI112(ofifoData[368]), .DI111(ofifoData[367]), .DI110(ofifoData[366]), .DI109(ofifoData[365]), .DI108(ofifoData[364]), .DI107(ofifoData[363]), .DI106(ofifoData[362]), .DI105(ofifoData[361]),
 .DI104(ofifoData[360]), .DI103(ofifoData[359]), .DI102(ofifoData[358]), .DI101(ofifoData[357]), .DI100(ofifoData[356]), .DI99(ofifoData[355]), .DI98(ofifoData[354]), .DI97(ofifoData[353]),
 .DI96(ofifoData[352]), .DI95(ofifoData[351]), .DI94(ofifoData[350]), .DI93(ofifoData[349]), .DI92(ofifoData[348]), .DI91(ofifoData[347]), .DI90(ofifoData[346]), .DI89(ofifoData[345]),
 .DI88(ofifoData[344]), .DI87(ofifoData[343]), .DI86(ofifoData[342]), .DI85(ofifoData[341]), .DI84(ofifoData[340]), .DI83(ofifoData[339]), .DI82(ofifoData[338]), .DI81(ofifoData[337]),
 .DI80(ofifoData[336]), .DI79(ofifoData[335]), .DI78(ofifoData[334]), .DI77(ofifoData[333]), .DI76(ofifoData[332]), .DI75(ofifoData[331]), .DI74(ofifoData[330]), .DI73(ofifoData[329]),
 .DI72(ofifoData[328]), .DI71(ofifoData[327]), .DI70(ofifoData[326]), .DI69(ofifoData[325]), .DI68(ofifoData[324]), .DI67(ofifoData[323]), .DI66(ofifoData[322]), .DI65(ofifoData[321]),
 .DI64(ofifoData[320]), .DI63(ofifoData[319]), .DI62(ofifoData[318]), .DI61(ofifoData[317]), .DI60(ofifoData[316]), .DI59(ofifoData[315]), .DI58(ofifoData[314]), .DI57(ofifoData[313]),
 .DI56(ofifoData[312]), .DI55(ofifoData[311]), .DI54(ofifoData[310]), .DI53(ofifoData[309]), .DI52(ofifoData[308]), .DI51(ofifoData[307]), .DI50(ofifoData[306]), .DI49(ofifoData[305]),
 .DI48(ofifoData[304]), .DI47(ofifoData[303]), .DI46(ofifoData[302]), .DI45(ofifoData[301]), .DI44(ofifoData[300]), .DI43(ofifoData[299]), .DI42(ofifoData[298]), .DI41(ofifoData[297]),
 .DI40(ofifoData[296]), .DI39(ofifoData[295]), .DI38(ofifoData[294]), .DI37(ofifoData[293]), .DI36(ofifoData[292]), .DI35(ofifoData[291]), .DI34(ofifoData[290]), .DI33(ofifoData[289]),
 .DI32(ofifoData[288]), .DI31(ofifoData[287]), .DI30(ofifoData[286]), .DI29(ofifoData[285]), .DI28(ofifoData[284]), .DI27(ofifoData[283]), .DI26(ofifoData[282]), .DI25(ofifoData[281]),
 .DI24(ofifoData[280]), .DI23(ofifoData[279]), .DI22(ofifoData[278]), .DI21(ofifoData[277]), .DI20(ofifoData[276]), .DI19(ofifoData[275]), .DI18(ofifoData[274]), .DI17(ofifoData[273]),
 .DI16(ofifoData[272]), .DI15(ofifoData[271]), .DI14(ofifoData[270]), .DI13(ofifoData[269]), .DI12(ofifoData[268]), .DI11(ofifoData[267]), .DI10(ofifoData[266]), .DI9(ofifoData[265]),
 .DI8(ofifoData[264]), .DI7(ofifoData[263]), .DI6(ofifoData[262]), .DI5(ofifoData[261]), .DI4(ofifoData[260]), .DI3(ofifoData[259]), .DI2(ofifoData[258]), .DI1(ofifoData[257]),
 .DI0(ofifoData[256]), .WE(n5632), .SYNC_IN(n9334), .SYNC_OUT(n9335));
MPW32KX256 U10461 ( .A14(ofifoAddr2[14]), .A13(ofifoAddr2[13]), .A12(ofifoAddr2[12]), .A11(ofifoAddr2[11]), .A10(ofifoAddr2[10]), .A9(ofifoAddr2[9]),
 .A8(ofifoAddr2[8]), .A7(ofifoAddr2[7]), .A6(ofifoAddr2[6]), .A5(ofifoAddr2[5]), .A4(ofifoAddr2[4]), .A3(ofifoAddr2[3]), .A2(ofifoAddr2[2]), .A1(ofifoAddr2[1]),
 .A0(ofifoAddr2[0]), .DI255(ofifoData[767]), .DI254(ofifoData[766]), .DI253(ofifoData[765]), .DI252(ofifoData[764]), .DI251(ofifoData[763]), .DI250(ofifoData[762]), .DI249(ofifoData[761]),
 .DI248(ofifoData[760]), .DI247(ofifoData[759]), .DI246(ofifoData[758]), .DI245(ofifoData[757]), .DI244(ofifoData[756]), .DI243(ofifoData[755]), .DI242(ofifoData[754]), .DI241(ofifoData[753]),
 .DI240(ofifoData[752]), .DI239(ofifoData[751]), .DI238(ofifoData[750]), .DI237(ofifoData[749]), .DI236(ofifoData[748]), .DI235(ofifoData[747]), .DI234(ofifoData[746]), .DI233(ofifoData[745]),
 .DI232(ofifoData[744]), .DI231(ofifoData[743]), .DI230(ofifoData[742]), .DI229(ofifoData[741]), .DI228(ofifoData[740]), .DI227(ofifoData[739]), .DI226(ofifoData[738]), .DI225(ofifoData[737]),
 .DI224(ofifoData[736]), .DI223(ofifoData[735]), .DI222(ofifoData[734]), .DI221(ofifoData[733]), .DI220(ofifoData[732]), .DI219(ofifoData[731]), .DI218(ofifoData[730]), .DI217(ofifoData[729]),
 .DI216(ofifoData[728]), .DI215(ofifoData[727]), .DI214(ofifoData[726]), .DI213(ofifoData[725]), .DI212(ofifoData[724]), .DI211(ofifoData[723]), .DI210(ofifoData[722]), .DI209(ofifoData[721]),
 .DI208(ofifoData[720]), .DI207(ofifoData[719]), .DI206(ofifoData[718]), .DI205(ofifoData[717]), .DI204(ofifoData[716]), .DI203(ofifoData[715]), .DI202(ofifoData[714]), .DI201(ofifoData[713]),
 .DI200(ofifoData[712]), .DI199(ofifoData[711]), .DI198(ofifoData[710]), .DI197(ofifoData[709]), .DI196(ofifoData[708]), .DI195(ofifoData[707]), .DI194(ofifoData[706]), .DI193(ofifoData[705]),
 .DI192(ofifoData[704]), .DI191(ofifoData[703]), .DI190(ofifoData[702]), .DI189(ofifoData[701]), .DI188(ofifoData[700]), .DI187(ofifoData[699]), .DI186(ofifoData[698]), .DI185(ofifoData[697]),
 .DI184(ofifoData[696]), .DI183(ofifoData[695]), .DI182(ofifoData[694]), .DI181(ofifoData[693]), .DI180(ofifoData[692]), .DI179(ofifoData[691]), .DI178(ofifoData[690]), .DI177(ofifoData[689]),
 .DI176(ofifoData[688]), .DI175(ofifoData[687]), .DI174(ofifoData[686]), .DI173(ofifoData[685]), .DI172(ofifoData[684]), .DI171(ofifoData[683]), .DI170(ofifoData[682]), .DI169(ofifoData[681]),
 .DI168(ofifoData[680]), .DI167(ofifoData[679]), .DI166(ofifoData[678]), .DI165(ofifoData[677]), .DI164(ofifoData[676]), .DI163(ofifoData[675]), .DI162(ofifoData[674]), .DI161(ofifoData[673]),
 .DI160(ofifoData[672]), .DI159(ofifoData[671]), .DI158(ofifoData[670]), .DI157(ofifoData[669]), .DI156(ofifoData[668]), .DI155(ofifoData[667]), .DI154(ofifoData[666]), .DI153(ofifoData[665]),
 .DI152(ofifoData[664]), .DI151(ofifoData[663]), .DI150(ofifoData[662]), .DI149(ofifoData[661]), .DI148(ofifoData[660]), .DI147(ofifoData[659]), .DI146(ofifoData[658]), .DI145(ofifoData[657]),
 .DI144(ofifoData[656]), .DI143(ofifoData[655]), .DI142(ofifoData[654]), .DI141(ofifoData[653]), .DI140(ofifoData[652]), .DI139(ofifoData[651]), .DI138(ofifoData[650]), .DI137(ofifoData[649]),
 .DI136(ofifoData[648]), .DI135(ofifoData[647]), .DI134(ofifoData[646]), .DI133(ofifoData[645]), .DI132(ofifoData[644]), .DI131(ofifoData[643]), .DI130(ofifoData[642]), .DI129(ofifoData[641]),
 .DI128(ofifoData[640]), .DI127(ofifoData[639]), .DI126(ofifoData[638]), .DI125(ofifoData[637]), .DI124(ofifoData[636]), .DI123(ofifoData[635]), .DI122(ofifoData[634]), .DI121(ofifoData[633]),
 .DI120(ofifoData[632]), .DI119(ofifoData[631]), .DI118(ofifoData[630]), .DI117(ofifoData[629]), .DI116(ofifoData[628]), .DI115(ofifoData[627]), .DI114(ofifoData[626]), .DI113(ofifoData[625]),
 .DI112(ofifoData[624]), .DI111(ofifoData[623]), .DI110(ofifoData[622]), .DI109(ofifoData[621]), .DI108(ofifoData[620]), .DI107(ofifoData[619]), .DI106(ofifoData[618]), .DI105(ofifoData[617]),
 .DI104(ofifoData[616]), .DI103(ofifoData[615]), .DI102(ofifoData[614]), .DI101(ofifoData[613]), .DI100(ofifoData[612]), .DI99(ofifoData[611]), .DI98(ofifoData[610]), .DI97(ofifoData[609]),
 .DI96(ofifoData[608]), .DI95(ofifoData[607]), .DI94(ofifoData[606]), .DI93(ofifoData[605]), .DI92(ofifoData[604]), .DI91(ofifoData[603]), .DI90(ofifoData[602]), .DI89(ofifoData[601]),
 .DI88(ofifoData[600]), .DI87(ofifoData[599]), .DI86(ofifoData[598]), .DI85(ofifoData[597]), .DI84(ofifoData[596]), .DI83(ofifoData[595]), .DI82(ofifoData[594]), .DI81(ofifoData[593]),
 .DI80(ofifoData[592]), .DI79(ofifoData[591]), .DI78(ofifoData[590]), .DI77(ofifoData[589]), .DI76(ofifoData[588]), .DI75(ofifoData[587]), .DI74(ofifoData[586]), .DI73(ofifoData[585]),
 .DI72(ofifoData[584]), .DI71(ofifoData[583]), .DI70(ofifoData[582]), .DI69(ofifoData[581]), .DI68(ofifoData[580]), .DI67(ofifoData[579]), .DI66(ofifoData[578]), .DI65(ofifoData[577]),
 .DI64(ofifoData[576]), .DI63(ofifoData[575]), .DI62(ofifoData[574]), .DI61(ofifoData[573]), .DI60(ofifoData[572]), .DI59(ofifoData[571]), .DI58(ofifoData[570]), .DI57(ofifoData[569]),
 .DI56(ofifoData[568]), .DI55(ofifoData[567]), .DI54(ofifoData[566]), .DI53(ofifoData[565]), .DI52(ofifoData[564]), .DI51(ofifoData[563]), .DI50(ofifoData[562]), .DI49(ofifoData[561]),
 .DI48(ofifoData[560]), .DI47(ofifoData[559]), .DI46(ofifoData[558]), .DI45(ofifoData[557]), .DI44(ofifoData[556]), .DI43(ofifoData[555]), .DI42(ofifoData[554]), .DI41(ofifoData[553]),
 .DI40(ofifoData[552]), .DI39(ofifoData[551]), .DI38(ofifoData[550]), .DI37(ofifoData[549]), .DI36(ofifoData[548]), .DI35(ofifoData[547]), .DI34(ofifoData[546]), .DI33(ofifoData[545]),
 .DI32(ofifoData[544]), .DI31(ofifoData[543]), .DI30(ofifoData[542]), .DI29(ofifoData[541]), .DI28(ofifoData[540]), .DI27(ofifoData[539]), .DI26(ofifoData[538]), .DI25(ofifoData[537]),
 .DI24(ofifoData[536]), .DI23(ofifoData[535]), .DI22(ofifoData[534]), .DI21(ofifoData[533]), .DI20(ofifoData[532]), .DI19(ofifoData[531]), .DI18(ofifoData[530]), .DI17(ofifoData[529]),
 .DI16(ofifoData[528]), .DI15(ofifoData[527]), .DI14(ofifoData[526]), .DI13(ofifoData[525]), .DI12(ofifoData[524]), .DI11(ofifoData[523]), .DI10(ofifoData[522]), .DI9(ofifoData[521]),
 .DI8(ofifoData[520]), .DI7(ofifoData[519]), .DI6(ofifoData[518]), .DI5(ofifoData[517]), .DI4(ofifoData[516]), .DI3(ofifoData[515]), .DI2(ofifoData[514]), .DI1(ofifoData[513]),
 .DI0(ofifoData[512]), .WE(n5633), .SYNC_IN(n9335), .SYNC_OUT( ));
`endif
`ifdef CBV

reg [255:0] ixc_gfm_ififo [0:32767];
initial begin: U10462
  integer j;
  for (j=0; j<=32767; j=j+1) ixc_gfm_ififo[j] =
`ifdef CBV_MEM_INIT1
  {256{1'b1}};
`else
  256'b0;
`endif
end
reg [255:0] n9336;
assign {ififoXdata[255], ififoXdata[254], ififoXdata[253], ififoXdata[252], ififoXdata[251], ififoXdata[250], ififoXdata[249],
ififoXdata[248], ififoXdata[247], ififoXdata[246], ififoXdata[245], ififoXdata[244], ififoXdata[243], ififoXdata[242], ififoXdata[241],
ififoXdata[240], ififoXdata[239], ififoXdata[238], ififoXdata[237], ififoXdata[236], ififoXdata[235], ififoXdata[234], ififoXdata[233],
ififoXdata[232], ififoXdata[231], ififoXdata[230], ififoXdata[229], ififoXdata[228], ififoXdata[227], ififoXdata[226], ififoXdata[225],
ififoXdata[224], ififoXdata[223], ififoXdata[222], ififoXdata[221], ififoXdata[220], ififoXdata[219], ififoXdata[218], ififoXdata[217],
ififoXdata[216], ififoXdata[215], ififoXdata[214], ififoXdata[213], ififoXdata[212], ififoXdata[211], ififoXdata[210], ififoXdata[209],
ififoXdata[208], ififoXdata[207], ififoXdata[206], ififoXdata[205], ififoXdata[204], ififoXdata[203], ififoXdata[202], ififoXdata[201],
ififoXdata[200], ififoXdata[199], ififoXdata[198], ififoXdata[197], ififoXdata[196], ififoXdata[195], ififoXdata[194], ififoXdata[193],
ififoXdata[192], ififoXdata[191], ififoXdata[190], ififoXdata[189], ififoXdata[188], ififoXdata[187], ififoXdata[186], ififoXdata[185],
ififoXdata[184], ififoXdata[183], ififoXdata[182], ififoXdata[181], ififoXdata[180], ififoXdata[179], ififoXdata[178], ififoXdata[177],
ififoXdata[176], ififoXdata[175], ififoXdata[174], ififoXdata[173], ififoXdata[172], ififoXdata[171], ififoXdata[170], ififoXdata[169],
ififoXdata[168], ififoXdata[167], ififoXdata[166], ififoXdata[165], ififoXdata[164], ififoXdata[163], ififoXdata[162], ififoXdata[161],
ififoXdata[160], ififoXdata[159], ififoXdata[158], ififoXdata[157], ififoXdata[156], ififoXdata[155], ififoXdata[154], ififoXdata[153],
ififoXdata[152], ififoXdata[151], ififoXdata[150], ififoXdata[149], ififoXdata[148], ififoXdata[147], ififoXdata[146], ififoXdata[145],
ififoXdata[144], ififoXdata[143], ififoXdata[142], ififoXdata[141], ififoXdata[140], ififoXdata[139], ififoXdata[138], ififoXdata[137],
ififoXdata[136], ififoXdata[135], ififoXdata[134], ififoXdata[133], ififoXdata[132], ififoXdata[131], ififoXdata[130], ififoXdata[129],
ififoXdata[128], ififoXdata[127], ififoXdata[126], ififoXdata[125], ififoXdata[124], ififoXdata[123], ififoXdata[122], ififoXdata[121],
ififoXdata[120], ififoXdata[119], ififoXdata[118], ififoXdata[117], ififoXdata[116], ififoXdata[115], ififoXdata[114], ififoXdata[113],
ififoXdata[112], ififoXdata[111], ififoXdata[110], ififoXdata[109], ififoXdata[108], ififoXdata[107], ififoXdata[106], ififoXdata[105],
ififoXdata[104], ififoXdata[103], ififoXdata[102], ififoXdata[101], ififoXdata[100], ififoXdata[99], ififoXdata[98], ififoXdata[97],
ififoXdata[96], ififoXdata[95], ififoXdata[94], ififoXdata[93], ififoXdata[92], ififoXdata[91], ififoXdata[90], ififoXdata[89],
ififoXdata[88], ififoXdata[87], ififoXdata[86], ififoXdata[85], ififoXdata[84], ififoXdata[83], ififoXdata[82], ififoXdata[81],
ififoXdata[80], ififoXdata[79], ififoXdata[78], ififoXdata[77], ififoXdata[76], ififoXdata[75], ififoXdata[74], ififoXdata[73],
ififoXdata[72], ififoXdata[71], ififoXdata[70], ififoXdata[69], ififoXdata[68], ififoXdata[67], ififoXdata[66], ififoXdata[65],
ififoXdata[64], ififoXdata[63], ififoXdata[62], ififoXdata[61], ififoXdata[60], ififoXdata[59], ififoXdata[58], ififoXdata[57],
ififoXdata[56], ififoXdata[55], ififoXdata[54], ififoXdata[53], ififoXdata[52], ififoXdata[51], ififoXdata[50], ififoXdata[49],
ififoXdata[48], ififoXdata[47], ififoXdata[46], ififoXdata[45], ififoXdata[44], ififoXdata[43], ififoXdata[42], ififoXdata[41],
ififoXdata[40], ififoXdata[39], ififoXdata[38], ififoXdata[37], ififoXdata[36], ififoXdata[35], ififoXdata[34], ififoXdata[33],
ififoXdata[32], ififoXdata[31], ififoXdata[30], ififoXdata[29], ififoXdata[28], ififoXdata[27], ififoXdata[26], ififoXdata[25],
ififoXdata[24], ififoXdata[23], ififoXdata[22], ififoXdata[21], ififoXdata[20], ififoXdata[19], ififoXdata[18], ififoXdata[17],
ififoXdata[16], ififoXdata[15], ififoXdata[14], ififoXdata[13], ififoXdata[12], ififoXdata[11], ififoXdata[10], ififoXdata[9],
ififoXdata[8], ififoXdata[7], ififoXdata[6], ififoXdata[5], ififoXdata[4], ififoXdata[3], ififoXdata[2], ififoXdata[1],
ififoXdata[0]} = n9336; 
reg [255:0] n9337;
assign {ififoRdata[255], ififoRdata[254], ififoRdata[253], ififoRdata[252], ififoRdata[251], ififoRdata[250], ififoRdata[249],
ififoRdata[248], ififoRdata[247], ififoRdata[246], ififoRdata[245], ififoRdata[244], ififoRdata[243], ififoRdata[242], ififoRdata[241],
ififoRdata[240], ififoRdata[239], ififoRdata[238], ififoRdata[237], ififoRdata[236], ififoRdata[235], ififoRdata[234], ififoRdata[233],
ififoRdata[232], ififoRdata[231], ififoRdata[230], ififoRdata[229], ififoRdata[228], ififoRdata[227], ififoRdata[226], ififoRdata[225],
ififoRdata[224], ififoRdata[223], ififoRdata[222], ififoRdata[221], ififoRdata[220], ififoRdata[219], ififoRdata[218], ififoRdata[217],
ififoRdata[216], ififoRdata[215], ififoRdata[214], ififoRdata[213], ififoRdata[212], ififoRdata[211], ififoRdata[210], ififoRdata[209],
ififoRdata[208], ififoRdata[207], ififoRdata[206], ififoRdata[205], ififoRdata[204], ififoRdata[203], ififoRdata[202], ififoRdata[201],
ififoRdata[200], ififoRdata[199], ififoRdata[198], ififoRdata[197], ififoRdata[196], ififoRdata[195], ififoRdata[194], ififoRdata[193],
ififoRdata[192], ififoRdata[191], ififoRdata[190], ififoRdata[189], ififoRdata[188], ififoRdata[187], ififoRdata[186], ififoRdata[185],
ififoRdata[184], ififoRdata[183], ififoRdata[182], ififoRdata[181], ififoRdata[180], ififoRdata[179], ififoRdata[178], ififoRdata[177],
ififoRdata[176], ififoRdata[175], ififoRdata[174], ififoRdata[173], ififoRdata[172], ififoRdata[171], ififoRdata[170], ififoRdata[169],
ififoRdata[168], ififoRdata[167], ififoRdata[166], ififoRdata[165], ififoRdata[164], ififoRdata[163], ififoRdata[162], ififoRdata[161],
ififoRdata[160], ififoRdata[159], ififoRdata[158], ififoRdata[157], ififoRdata[156], ififoRdata[155], ififoRdata[154], ififoRdata[153],
ififoRdata[152], ififoRdata[151], ififoRdata[150], ififoRdata[149], ififoRdata[148], ififoRdata[147], ififoRdata[146], ififoRdata[145],
ififoRdata[144], ififoRdata[143], ififoRdata[142], ififoRdata[141], ififoRdata[140], ififoRdata[139], ififoRdata[138], ififoRdata[137],
ififoRdata[136], ififoRdata[135], ififoRdata[134], ififoRdata[133], ififoRdata[132], ififoRdata[131], ififoRdata[130], ififoRdata[129],
ififoRdata[128], ififoRdata[127], ififoRdata[126], ififoRdata[125], ififoRdata[124], ififoRdata[123], ififoRdata[122], ififoRdata[121],
ififoRdata[120], ififoRdata[119], ififoRdata[118], ififoRdata[117], ififoRdata[116], ififoRdata[115], ififoRdata[114], ififoRdata[113],
ififoRdata[112], ififoRdata[111], ififoRdata[110], ififoRdata[109], ififoRdata[108], ififoRdata[107], ififoRdata[106], ififoRdata[105],
ififoRdata[104], ififoRdata[103], ififoRdata[102], ififoRdata[101], ififoRdata[100], ififoRdata[99], ififoRdata[98], ififoRdata[97],
ififoRdata[96], ififoRdata[95], ififoRdata[94], ififoRdata[93], ififoRdata[92], ififoRdata[91], ififoRdata[90], ififoRdata[89],
ififoRdata[88], ififoRdata[87], ififoRdata[86], ififoRdata[85], ififoRdata[84], ififoRdata[83], ififoRdata[82], ififoRdata[81],
ififoRdata[80], ififoRdata[79], ififoRdata[78], ififoRdata[77], ififoRdata[76], ififoRdata[75], ififoRdata[74], ififoRdata[73],
ififoRdata[72], ififoRdata[71], ififoRdata[70], ififoRdata[69], ififoRdata[68], ififoRdata[67], ififoRdata[66], ififoRdata[65],
ififoRdata[64], ififoRdata[63], ififoRdata[62], ififoRdata[61], ififoRdata[60], ififoRdata[59], ififoRdata[58], ififoRdata[57],
ififoRdata[56], ififoRdata[55], ififoRdata[54], ififoRdata[53], ififoRdata[52], ififoRdata[51], ififoRdata[50], ififoRdata[49],
ififoRdata[48], ififoRdata[47], ififoRdata[46], ififoRdata[45], ififoRdata[44], ififoRdata[43], ififoRdata[42], ififoRdata[41],
ififoRdata[40], ififoRdata[39], ififoRdata[38], ififoRdata[37], ififoRdata[36], ififoRdata[35], ififoRdata[34], ififoRdata[33],
ififoRdata[32], ififoRdata[31], ififoRdata[30], ififoRdata[29], ififoRdata[28], ififoRdata[27], ififoRdata[26], ififoRdata[25],
ififoRdata[24], ififoRdata[23], ififoRdata[22], ififoRdata[21], ififoRdata[20], ififoRdata[19], ififoRdata[18], ififoRdata[17],
ififoRdata[16], ififoRdata[15], ififoRdata[14], ififoRdata[13], ififoRdata[12], ififoRdata[11], ififoRdata[10], ififoRdata[9],
ififoRdata[8], ififoRdata[7], ififoRdata[6], ififoRdata[5], ififoRdata[4], ififoRdata[3], ififoRdata[2], ififoRdata[1],
ififoRdata[0]} = n9337; 
reg [255:0] n9338;
assign {ififoRdata[511], ififoRdata[510], ififoRdata[509], ififoRdata[508], ififoRdata[507], ififoRdata[506], ififoRdata[505],
ififoRdata[504], ififoRdata[503], ififoRdata[502], ififoRdata[501], ififoRdata[500], ififoRdata[499], ififoRdata[498], ififoRdata[497],
ififoRdata[496], ififoRdata[495], ififoRdata[494], ififoRdata[493], ififoRdata[492], ififoRdata[491], ififoRdata[490], ififoRdata[489],
ififoRdata[488], ififoRdata[487], ififoRdata[486], ififoRdata[485], ififoRdata[484], ififoRdata[483], ififoRdata[482], ififoRdata[481],
ififoRdata[480], ififoRdata[479], ififoRdata[478], ififoRdata[477], ififoRdata[476], ififoRdata[475], ififoRdata[474], ififoRdata[473],
ififoRdata[472], ififoRdata[471], ififoRdata[470], ififoRdata[469], ififoRdata[468], ififoRdata[467], ififoRdata[466], ififoRdata[465],
ififoRdata[464], ififoRdata[463], ififoRdata[462], ififoRdata[461], ififoRdata[460], ififoRdata[459], ififoRdata[458], ififoRdata[457],
ififoRdata[456], ififoRdata[455], ififoRdata[454], ififoRdata[453], ififoRdata[452], ififoRdata[451], ififoRdata[450], ififoRdata[449],
ififoRdata[448], ififoRdata[447], ififoRdata[446], ififoRdata[445], ififoRdata[444], ififoRdata[443], ififoRdata[442], ififoRdata[441],
ififoRdata[440], ififoRdata[439], ififoRdata[438], ififoRdata[437], ififoRdata[436], ififoRdata[435], ififoRdata[434], ififoRdata[433],
ififoRdata[432], ififoRdata[431], ififoRdata[430], ififoRdata[429], ififoRdata[428], ififoRdata[427], ififoRdata[426], ififoRdata[425],
ififoRdata[424], ififoRdata[423], ififoRdata[422], ififoRdata[421], ififoRdata[420], ififoRdata[419], ififoRdata[418], ififoRdata[417],
ififoRdata[416], ififoRdata[415], ififoRdata[414], ififoRdata[413], ififoRdata[412], ififoRdata[411], ififoRdata[410], ififoRdata[409],
ififoRdata[408], ififoRdata[407], ififoRdata[406], ififoRdata[405], ififoRdata[404], ififoRdata[403], ififoRdata[402], ififoRdata[401],
ififoRdata[400], ififoRdata[399], ififoRdata[398], ififoRdata[397], ififoRdata[396], ififoRdata[395], ififoRdata[394], ififoRdata[393],
ififoRdata[392], ififoRdata[391], ififoRdata[390], ififoRdata[389], ififoRdata[388], ififoRdata[387], ififoRdata[386], ififoRdata[385],
ififoRdata[384], ififoRdata[383], ififoRdata[382], ififoRdata[381], ififoRdata[380], ififoRdata[379], ififoRdata[378], ififoRdata[377],
ififoRdata[376], ififoRdata[375], ififoRdata[374], ififoRdata[373], ififoRdata[372], ififoRdata[371], ififoRdata[370], ififoRdata[369],
ififoRdata[368], ififoRdata[367], ififoRdata[366], ififoRdata[365], ififoRdata[364], ififoRdata[363], ififoRdata[362], ififoRdata[361],
ififoRdata[360], ififoRdata[359], ififoRdata[358], ififoRdata[357], ififoRdata[356], ififoRdata[355], ififoRdata[354], ififoRdata[353],
ififoRdata[352], ififoRdata[351], ififoRdata[350], ififoRdata[349], ififoRdata[348], ififoRdata[347], ififoRdata[346], ififoRdata[345],
ififoRdata[344], ififoRdata[343], ififoRdata[342], ififoRdata[341], ififoRdata[340], ififoRdata[339], ififoRdata[338], ififoRdata[337],
ififoRdata[336], ififoRdata[335], ififoRdata[334], ififoRdata[333], ififoRdata[332], ififoRdata[331], ififoRdata[330], ififoRdata[329],
ififoRdata[328], ififoRdata[327], ififoRdata[326], ififoRdata[325], ififoRdata[324], ififoRdata[323], ififoRdata[322], ififoRdata[321],
ififoRdata[320], ififoRdata[319], ififoRdata[318], ififoRdata[317], ififoRdata[316], ififoRdata[315], ififoRdata[314], ififoRdata[313],
ififoRdata[312], ififoRdata[311], ififoRdata[310], ififoRdata[309], ififoRdata[308], ififoRdata[307], ififoRdata[306], ififoRdata[305],
ififoRdata[304], ififoRdata[303], ififoRdata[302], ififoRdata[301], ififoRdata[300], ififoRdata[299], ififoRdata[298], ififoRdata[297],
ififoRdata[296], ififoRdata[295], ififoRdata[294], ififoRdata[293], ififoRdata[292], ififoRdata[291], ififoRdata[290], ififoRdata[289],
ififoRdata[288], ififoRdata[287], ififoRdata[286], ififoRdata[285], ififoRdata[284], ififoRdata[283], ififoRdata[282], ififoRdata[281],
ififoRdata[280], ififoRdata[279], ififoRdata[278], ififoRdata[277], ififoRdata[276], ififoRdata[275], ififoRdata[274], ififoRdata[273],
ififoRdata[272], ififoRdata[271], ififoRdata[270], ififoRdata[269], ififoRdata[268], ififoRdata[267], ififoRdata[266], ififoRdata[265],
ififoRdata[264], ififoRdata[263], ififoRdata[262], ififoRdata[261], ififoRdata[260], ififoRdata[259], ififoRdata[258], ififoRdata[257],
ififoRdata[256]} = n9338; 
reg [255:0] n9339;
assign {ififoRdata[767], ififoRdata[766], ififoRdata[765], ififoRdata[764], ififoRdata[763], ififoRdata[762], ififoRdata[761],
ififoRdata[760], ififoRdata[759], ififoRdata[758], ififoRdata[757], ififoRdata[756], ififoRdata[755], ififoRdata[754], ififoRdata[753],
ififoRdata[752], ififoRdata[751], ififoRdata[750], ififoRdata[749], ififoRdata[748], ififoRdata[747], ififoRdata[746], ififoRdata[745],
ififoRdata[744], ififoRdata[743], ififoRdata[742], ififoRdata[741], ififoRdata[740], ififoRdata[739], ififoRdata[738], ififoRdata[737],
ififoRdata[736], ififoRdata[735], ififoRdata[734], ififoRdata[733], ififoRdata[732], ififoRdata[731], ififoRdata[730], ififoRdata[729],
ififoRdata[728], ififoRdata[727], ififoRdata[726], ififoRdata[725], ififoRdata[724], ififoRdata[723], ififoRdata[722], ififoRdata[721],
ififoRdata[720], ififoRdata[719], ififoRdata[718], ififoRdata[717], ififoRdata[716], ififoRdata[715], ififoRdata[714], ififoRdata[713],
ififoRdata[712], ififoRdata[711], ififoRdata[710], ififoRdata[709], ififoRdata[708], ififoRdata[707], ififoRdata[706], ififoRdata[705],
ififoRdata[704], ififoRdata[703], ififoRdata[702], ififoRdata[701], ififoRdata[700], ififoRdata[699], ififoRdata[698], ififoRdata[697],
ififoRdata[696], ififoRdata[695], ififoRdata[694], ififoRdata[693], ififoRdata[692], ififoRdata[691], ififoRdata[690], ififoRdata[689],
ififoRdata[688], ififoRdata[687], ififoRdata[686], ififoRdata[685], ififoRdata[684], ififoRdata[683], ififoRdata[682], ififoRdata[681],
ififoRdata[680], ififoRdata[679], ififoRdata[678], ififoRdata[677], ififoRdata[676], ififoRdata[675], ififoRdata[674], ififoRdata[673],
ififoRdata[672], ififoRdata[671], ififoRdata[670], ififoRdata[669], ififoRdata[668], ififoRdata[667], ififoRdata[666], ififoRdata[665],
ififoRdata[664], ififoRdata[663], ififoRdata[662], ififoRdata[661], ififoRdata[660], ififoRdata[659], ififoRdata[658], ififoRdata[657],
ififoRdata[656], ififoRdata[655], ififoRdata[654], ififoRdata[653], ififoRdata[652], ififoRdata[651], ififoRdata[650], ififoRdata[649],
ififoRdata[648], ififoRdata[647], ififoRdata[646], ififoRdata[645], ififoRdata[644], ififoRdata[643], ififoRdata[642], ififoRdata[641],
ififoRdata[640], ififoRdata[639], ififoRdata[638], ififoRdata[637], ififoRdata[636], ififoRdata[635], ififoRdata[634], ififoRdata[633],
ififoRdata[632], ififoRdata[631], ififoRdata[630], ififoRdata[629], ififoRdata[628], ififoRdata[627], ififoRdata[626], ififoRdata[625],
ififoRdata[624], ififoRdata[623], ififoRdata[622], ififoRdata[621], ififoRdata[620], ififoRdata[619], ififoRdata[618], ififoRdata[617],
ififoRdata[616], ififoRdata[615], ififoRdata[614], ififoRdata[613], ififoRdata[612], ififoRdata[611], ififoRdata[610], ififoRdata[609],
ififoRdata[608], ififoRdata[607], ififoRdata[606], ififoRdata[605], ififoRdata[604], ififoRdata[603], ififoRdata[602], ififoRdata[601],
ififoRdata[600], ififoRdata[599], ififoRdata[598], ififoRdata[597], ififoRdata[596], ififoRdata[595], ififoRdata[594], ififoRdata[593],
ififoRdata[592], ififoRdata[591], ififoRdata[590], ififoRdata[589], ififoRdata[588], ififoRdata[587], ififoRdata[586], ififoRdata[585],
ififoRdata[584], ififoRdata[583], ififoRdata[582], ififoRdata[581], ififoRdata[580], ififoRdata[579], ififoRdata[578], ififoRdata[577],
ififoRdata[576], ififoRdata[575], ififoRdata[574], ififoRdata[573], ififoRdata[572], ififoRdata[571], ififoRdata[570], ififoRdata[569],
ififoRdata[568], ififoRdata[567], ififoRdata[566], ififoRdata[565], ififoRdata[564], ififoRdata[563], ififoRdata[562], ififoRdata[561],
ififoRdata[560], ififoRdata[559], ififoRdata[558], ififoRdata[557], ififoRdata[556], ififoRdata[555], ififoRdata[554], ififoRdata[553],
ififoRdata[552], ififoRdata[551], ififoRdata[550], ififoRdata[549], ififoRdata[548], ififoRdata[547], ififoRdata[546], ififoRdata[545],
ififoRdata[544], ififoRdata[543], ififoRdata[542], ififoRdata[541], ififoRdata[540], ififoRdata[539], ififoRdata[538], ififoRdata[537],
ififoRdata[536], ififoRdata[535], ififoRdata[534], ififoRdata[533], ififoRdata[532], ififoRdata[531], ififoRdata[530], ififoRdata[529],
ififoRdata[528], ififoRdata[527], ififoRdata[526], ififoRdata[525], ififoRdata[524], ififoRdata[523], ififoRdata[522], ififoRdata[521],
ififoRdata[520], ififoRdata[519], ififoRdata[518], ififoRdata[517], ififoRdata[516], ififoRdata[515], ififoRdata[514], ififoRdata[513],
ififoRdata[512]} = n9339; 
always @(n259 or n260 or n261 or n262 or n263
 or n264 or n265 or n266 or n267 or n268 or n269 or n270 or n271
 or n272 or n273 or n3 or n4 or n5 or n6 or n7 or n8
 or n9 or n10 or n11 or n12 or n13 or n14 or n15 or n16
 or n17 or n18 or n19 or n20 or n21 or n22 or n23 or n24
 or n25 or n26 or n27 or n28 or n29 or n30 or n31 or n32
 or n33 or n34 or n35 or n36 or n37 or n38 or n39 or n40
 or n41 or n42 or n43 or n44 or n45 or n46 or n47 or n48
 or n49 or n50 or n51 or n52 or n53 or n54 or n55 or n56
 or n57 or n58 or n59 or n60 or n61 or n62 or n63 or n64
 or n65 or n66 or n67 or n68 or n69 or n70 or n71 or n72
 or n73 or n74 or n75 or n76 or n77 or n78 or n79 or n80
 or n81 or n82 or n83 or n84 or n85 or n86 or n87 or n88
 or n89 or n90 or n91 or n92 or n93 or n94 or n95 or n96
 or n97 or n98 or n99 or n100 or n101 or n102 or n103 or n104
 or n105 or n106 or n107 or n108 or n109 or n110 or n111 or n112
 or n113 or n114 or n115 or n116 or n117 or n118 or n119 or n120
 or n121 or n122 or n123 or n124 or n125 or n126 or n127 or n128
 or n129 or n130 or n131 or n132 or n133 or n134 or n135 or n136
 or n137 or n138 or n139 or n140 or n141 or n142 or n143 or n144
 or n145 or n146 or n147 or n148 or n149 or n150 or n151 or n152
 or n153 or n154 or n155 or n156 or n157 or n158 or n159 or n160
 or n161 or n162 or n163 or n164 or n165 or n166 or n167 or n168
 or n169 or n170 or n171 or n172 or n173 or n174 or n175 or n176
 or n177 or n178 or n179 or n180 or n181 or n182 or n183 or n184
 or n185 or n186 or n187 or n188 or n189 or n190 or n191 or n192
 or n193 or n194 or n195 or n196 or n197 or n198 or n199 or n200
 or n201 or n202 or n203 or n204 or n205 or n206 or n207 or n208
 or n209 or n210 or n211 or n212 or n213 or n214 or n215 or n216
 or n217 or n218 or n219 or n220 or n221 or n222 or n223 or n224
 or n225 or n226 or n227 or n228 or n229 or n230 or n231 or n232
 or n233 or n234 or n235 or n236 or n237 or n238 or n239 or n240
 or n241 or n242 or n243 or n244 or n245 or n246 or n247 or n248
 or n249 or n250 or n251 or n252 or n253 or n254 or n255 or n256
 or n257 or n258 or n274 or xptr[16] or xptr[15] or xptr[14] or xptr[13] or xptr[12]
 or xptr[11] or xptr[10] or xptr[9] or xptr[8] or xptr[7] or xptr[6] or xptr[5] or xptr[4]
 or xptr[3] or xptr[2] or ififoRaddr0[14] or ififoRaddr0[13] or ififoRaddr0[12] or ififoRaddr0[11] or ififoRaddr0[10] or ififoRaddr0[9]
 or ififoRaddr0[8] or ififoRaddr0[7] or ififoRaddr0[6] or ififoRaddr0[5] or ififoRaddr0[4] or ififoRaddr0[3] or ififoRaddr0[2] or ififoRaddr0[1]
 or ififoRaddr0[0] or ififoRaddr1[14] or ififoRaddr1[13] or ififoRaddr1[12] or ififoRaddr1[11] or ififoRaddr1[10] or ififoRaddr1[9] or ififoRaddr1[8]
 or ififoRaddr1[7] or ififoRaddr1[6] or ififoRaddr1[5] or ififoRaddr1[4] or ififoRaddr1[3] or ififoRaddr1[2] or ififoRaddr1[1] or ififoRaddr1[0]
 or ififoRaddr2[14] or ififoRaddr2[13] or ififoRaddr2[12] or ififoRaddr2[11] or ififoRaddr2[10] or ififoRaddr2[9] or ififoRaddr2[8] or ififoRaddr2[7]
 or ififoRaddr2[6] or ififoRaddr2[5] or ififoRaddr2[4] or ififoRaddr2[3] or ififoRaddr2[2] or ififoRaddr2[1] or ififoRaddr2[0])
#0 begin
if (n274)
ixc_gfm_ififo[{n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273}] =
{n3, n4, n5, n6, n7,
 n8, n9, n10, n11, n12, n13, n14, n15,
 n16, n17, n18, n19, n20, n21, n22, n23,
 n24, n25, n26, n27, n28, n29, n30, n31,
 n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258};
n9336 = ixc_gfm_ififo[{xptr[16], xptr[15], xptr[14], xptr[13], xptr[12],
 xptr[11], xptr[10], xptr[9], xptr[8], xptr[7], xptr[6], xptr[5], xptr[4],
 xptr[3], xptr[2]}];
n9337 = ixc_gfm_ififo[{ififoRaddr0[14], ififoRaddr0[13], ififoRaddr0[12], ififoRaddr0[11], ififoRaddr0[10],
 ififoRaddr0[9], ififoRaddr0[8], ififoRaddr0[7], ififoRaddr0[6], ififoRaddr0[5], ififoRaddr0[4], ififoRaddr0[3], ififoRaddr0[2],
 ififoRaddr0[1], ififoRaddr0[0]}];
n9338 = ixc_gfm_ififo[{ififoRaddr1[14], ififoRaddr1[13], ififoRaddr1[12], ififoRaddr1[11], ififoRaddr1[10],
 ififoRaddr1[9], ififoRaddr1[8], ififoRaddr1[7], ififoRaddr1[6], ififoRaddr1[5], ififoRaddr1[4], ififoRaddr1[3], ififoRaddr1[2],
 ififoRaddr1[1], ififoRaddr1[0]}];
n9339 = ixc_gfm_ififo[{ififoRaddr2[14], ififoRaddr2[13], ififoRaddr2[12], ififoRaddr2[11], ififoRaddr2[10],
 ififoRaddr2[9], ififoRaddr2[8], ififoRaddr2[7], ififoRaddr2[6], ififoRaddr2[5], ififoRaddr2[4], ififoRaddr2[3], ififoRaddr2[2],
 ififoRaddr2[1], ififoRaddr2[0]}];
end
`else

MPW32KX256 ixc_gfm_ififo ( .A14(n259), .A13(n260), .A12(n261), .A11(n262), .A10(n263), .A9(n264),
 .A8(n265), .A7(n266), .A6(n267), .A5(n268), .A4(n269), .A3(n270), .A2(n271), .A1(n272),
 .A0(n273), .DI255(n3), .DI254(n4), .DI253(n5), .DI252(n6), .DI251(n7), .DI250(n8), .DI249(n9),
 .DI248(n10), .DI247(n11), .DI246(n12), .DI245(n13), .DI244(n14), .DI243(n15), .DI242(n16), .DI241(n17),
 .DI240(n18), .DI239(n19), .DI238(n20), .DI237(n21), .DI236(n22), .DI235(n23), .DI234(n24), .DI233(n25),
 .DI232(n26), .DI231(n27), .DI230(n28), .DI229(n29), .DI228(n30), .DI227(n31), .DI226(n32), .DI225(n33),
 .DI224(n34), .DI223(n35), .DI222(n36), .DI221(n37), .DI220(n38), .DI219(n39), .DI218(n40), .DI217(n41),
 .DI216(n42), .DI215(n43), .DI214(n44), .DI213(n45), .DI212(n46), .DI211(n47), .DI210(n48), .DI209(n49),
 .DI208(n50), .DI207(n51), .DI206(n52), .DI205(n53), .DI204(n54), .DI203(n55), .DI202(n56), .DI201(n57),
 .DI200(n58), .DI199(n59), .DI198(n60), .DI197(n61), .DI196(n62), .DI195(n63), .DI194(n64), .DI193(n65),
 .DI192(n66), .DI191(n67), .DI190(n68), .DI189(n69), .DI188(n70), .DI187(n71), .DI186(n72), .DI185(n73),
 .DI184(n74), .DI183(n75), .DI182(n76), .DI181(n77), .DI180(n78), .DI179(n79), .DI178(n80), .DI177(n81),
 .DI176(n82), .DI175(n83), .DI174(n84), .DI173(n85), .DI172(n86), .DI171(n87), .DI170(n88), .DI169(n89),
 .DI168(n90), .DI167(n91), .DI166(n92), .DI165(n93), .DI164(n94), .DI163(n95), .DI162(n96), .DI161(n97),
 .DI160(n98), .DI159(n99), .DI158(n100), .DI157(n101), .DI156(n102), .DI155(n103), .DI154(n104), .DI153(n105),
 .DI152(n106), .DI151(n107), .DI150(n108), .DI149(n109), .DI148(n110), .DI147(n111), .DI146(n112), .DI145(n113),
 .DI144(n114), .DI143(n115), .DI142(n116), .DI141(n117), .DI140(n118), .DI139(n119), .DI138(n120), .DI137(n121),
 .DI136(n122), .DI135(n123), .DI134(n124), .DI133(n125), .DI132(n126), .DI131(n127), .DI130(n128), .DI129(n129),
 .DI128(n130), .DI127(n131), .DI126(n132), .DI125(n133), .DI124(n134), .DI123(n135), .DI122(n136), .DI121(n137),
 .DI120(n138), .DI119(n139), .DI118(n140), .DI117(n141), .DI116(n142), .DI115(n143), .DI114(n144), .DI113(n145),
 .DI112(n146), .DI111(n147), .DI110(n148), .DI109(n149), .DI108(n150), .DI107(n151), .DI106(n152), .DI105(n153),
 .DI104(n154), .DI103(n155), .DI102(n156), .DI101(n157), .DI100(n158), .DI99(n159), .DI98(n160), .DI97(n161),
 .DI96(n162), .DI95(n163), .DI94(n164), .DI93(n165), .DI92(n166), .DI91(n167), .DI90(n168), .DI89(n169),
 .DI88(n170), .DI87(n171), .DI86(n172), .DI85(n173), .DI84(n174), .DI83(n175), .DI82(n176), .DI81(n177),
 .DI80(n178), .DI79(n179), .DI78(n180), .DI77(n181), .DI76(n182), .DI75(n183), .DI74(n184), .DI73(n185),
 .DI72(n186), .DI71(n187), .DI70(n188), .DI69(n189), .DI68(n190), .DI67(n191), .DI66(n192), .DI65(n193),
 .DI64(n194), .DI63(n195), .DI62(n196), .DI61(n197), .DI60(n198), .DI59(n199), .DI58(n200), .DI57(n201),
 .DI56(n202), .DI55(n203), .DI54(n204), .DI53(n205), .DI52(n206), .DI51(n207), .DI50(n208), .DI49(n209),
 .DI48(n210), .DI47(n211), .DI46(n212), .DI45(n213), .DI44(n214), .DI43(n215), .DI42(n216), .DI41(n217),
 .DI40(n218), .DI39(n219), .DI38(n220), .DI37(n221), .DI36(n222), .DI35(n223), .DI34(n224), .DI33(n225),
 .DI32(n226), .DI31(n227), .DI30(n228), .DI29(n229), .DI28(n230), .DI27(n231), .DI26(n232), .DI25(n233),
 .DI24(n234), .DI23(n235), .DI22(n236), .DI21(n237), .DI20(n238), .DI19(n239), .DI18(n240), .DI17(n241),
 .DI16(n242), .DI15(n243), .DI14(n244), .DI13(n245), .DI12(n246), .DI11(n247), .DI10(n248), .DI9(n249),
 .DI8(n250), .DI7(n251), .DI6(n252), .DI5(n253), .DI4(n254), .DI3(n255), .DI2(n256), .DI1(n257),
 .DI0(n258), .WE(n274), .SYNC_IN(n5631), .SYNC_OUT(n9336));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ififo" HDL_MEMORY_DECL "1 255 0 0 32767"
MPR32KX256 U10463 ( .A14(xptr[16]), .A13(xptr[15]), .A12(xptr[14]), .A11(xptr[13]), .A10(xptr[12]), .A9(xptr[11]),
 .A8(xptr[10]), .A7(xptr[9]), .A6(xptr[8]), .A5(xptr[7]), .A4(xptr[6]), .A3(xptr[5]), .A2(xptr[4]), .A1(xptr[3]),
 .A0(xptr[2]), .SYNC_IN(n9336), .DO255(ififoXdata[255]), .DO254(ififoXdata[254]), .DO253(ififoXdata[253]), .DO252(ififoXdata[252]), .DO251(ififoXdata[251]), .DO250(ififoXdata[250]),
 .DO249(ififoXdata[249]), .DO248(ififoXdata[248]), .DO247(ififoXdata[247]), .DO246(ififoXdata[246]), .DO245(ififoXdata[245]), .DO244(ififoXdata[244]), .DO243(ififoXdata[243]), .DO242(ififoXdata[242]),
 .DO241(ififoXdata[241]), .DO240(ififoXdata[240]), .DO239(ififoXdata[239]), .DO238(ififoXdata[238]), .DO237(ififoXdata[237]), .DO236(ififoXdata[236]), .DO235(ififoXdata[235]), .DO234(ififoXdata[234]),
 .DO233(ififoXdata[233]), .DO232(ififoXdata[232]), .DO231(ififoXdata[231]), .DO230(ififoXdata[230]), .DO229(ififoXdata[229]), .DO228(ififoXdata[228]), .DO227(ififoXdata[227]), .DO226(ififoXdata[226]),
 .DO225(ififoXdata[225]), .DO224(ififoXdata[224]), .DO223(ififoXdata[223]), .DO222(ififoXdata[222]), .DO221(ififoXdata[221]), .DO220(ififoXdata[220]), .DO219(ififoXdata[219]), .DO218(ififoXdata[218]),
 .DO217(ififoXdata[217]), .DO216(ififoXdata[216]), .DO215(ififoXdata[215]), .DO214(ififoXdata[214]), .DO213(ififoXdata[213]), .DO212(ififoXdata[212]), .DO211(ififoXdata[211]), .DO210(ififoXdata[210]),
 .DO209(ififoXdata[209]), .DO208(ififoXdata[208]), .DO207(ififoXdata[207]), .DO206(ififoXdata[206]), .DO205(ififoXdata[205]), .DO204(ififoXdata[204]), .DO203(ififoXdata[203]), .DO202(ififoXdata[202]),
 .DO201(ififoXdata[201]), .DO200(ififoXdata[200]), .DO199(ififoXdata[199]), .DO198(ififoXdata[198]), .DO197(ififoXdata[197]), .DO196(ififoXdata[196]), .DO195(ififoXdata[195]), .DO194(ififoXdata[194]),
 .DO193(ififoXdata[193]), .DO192(ififoXdata[192]), .DO191(ififoXdata[191]), .DO190(ififoXdata[190]), .DO189(ififoXdata[189]), .DO188(ififoXdata[188]), .DO187(ififoXdata[187]), .DO186(ififoXdata[186]),
 .DO185(ififoXdata[185]), .DO184(ififoXdata[184]), .DO183(ififoXdata[183]), .DO182(ififoXdata[182]), .DO181(ififoXdata[181]), .DO180(ififoXdata[180]), .DO179(ififoXdata[179]), .DO178(ififoXdata[178]),
 .DO177(ififoXdata[177]), .DO176(ififoXdata[176]), .DO175(ififoXdata[175]), .DO174(ififoXdata[174]), .DO173(ififoXdata[173]), .DO172(ififoXdata[172]), .DO171(ififoXdata[171]), .DO170(ififoXdata[170]),
 .DO169(ififoXdata[169]), .DO168(ififoXdata[168]), .DO167(ififoXdata[167]), .DO166(ififoXdata[166]), .DO165(ififoXdata[165]), .DO164(ififoXdata[164]), .DO163(ififoXdata[163]), .DO162(ififoXdata[162]),
 .DO161(ififoXdata[161]), .DO160(ififoXdata[160]), .DO159(ififoXdata[159]), .DO158(ififoXdata[158]), .DO157(ififoXdata[157]), .DO156(ififoXdata[156]), .DO155(ififoXdata[155]), .DO154(ififoXdata[154]),
 .DO153(ififoXdata[153]), .DO152(ififoXdata[152]), .DO151(ififoXdata[151]), .DO150(ififoXdata[150]), .DO149(ififoXdata[149]), .DO148(ififoXdata[148]), .DO147(ififoXdata[147]), .DO146(ififoXdata[146]),
 .DO145(ififoXdata[145]), .DO144(ififoXdata[144]), .DO143(ififoXdata[143]), .DO142(ififoXdata[142]), .DO141(ififoXdata[141]), .DO140(ififoXdata[140]), .DO139(ififoXdata[139]), .DO138(ififoXdata[138]),
 .DO137(ififoXdata[137]), .DO136(ififoXdata[136]), .DO135(ififoXdata[135]), .DO134(ififoXdata[134]), .DO133(ififoXdata[133]), .DO132(ififoXdata[132]), .DO131(ififoXdata[131]), .DO130(ififoXdata[130]),
 .DO129(ififoXdata[129]), .DO128(ififoXdata[128]), .DO127(ififoXdata[127]), .DO126(ififoXdata[126]), .DO125(ififoXdata[125]), .DO124(ififoXdata[124]), .DO123(ififoXdata[123]), .DO122(ififoXdata[122]),
 .DO121(ififoXdata[121]), .DO120(ififoXdata[120]), .DO119(ififoXdata[119]), .DO118(ififoXdata[118]), .DO117(ififoXdata[117]), .DO116(ififoXdata[116]), .DO115(ififoXdata[115]), .DO114(ififoXdata[114]),
 .DO113(ififoXdata[113]), .DO112(ififoXdata[112]), .DO111(ififoXdata[111]), .DO110(ififoXdata[110]), .DO109(ififoXdata[109]), .DO108(ififoXdata[108]), .DO107(ififoXdata[107]), .DO106(ififoXdata[106]),
 .DO105(ififoXdata[105]), .DO104(ififoXdata[104]), .DO103(ififoXdata[103]), .DO102(ififoXdata[102]), .DO101(ififoXdata[101]), .DO100(ififoXdata[100]), .DO99(ififoXdata[99]), .DO98(ififoXdata[98]),
 .DO97(ififoXdata[97]), .DO96(ififoXdata[96]), .DO95(ififoXdata[95]), .DO94(ififoXdata[94]), .DO93(ififoXdata[93]), .DO92(ififoXdata[92]), .DO91(ififoXdata[91]), .DO90(ififoXdata[90]),
 .DO89(ififoXdata[89]), .DO88(ififoXdata[88]), .DO87(ififoXdata[87]), .DO86(ififoXdata[86]), .DO85(ififoXdata[85]), .DO84(ififoXdata[84]), .DO83(ififoXdata[83]), .DO82(ififoXdata[82]),
 .DO81(ififoXdata[81]), .DO80(ififoXdata[80]), .DO79(ififoXdata[79]), .DO78(ififoXdata[78]), .DO77(ififoXdata[77]), .DO76(ififoXdata[76]), .DO75(ififoXdata[75]), .DO74(ififoXdata[74]),
 .DO73(ififoXdata[73]), .DO72(ififoXdata[72]), .DO71(ififoXdata[71]), .DO70(ififoXdata[70]), .DO69(ififoXdata[69]), .DO68(ififoXdata[68]), .DO67(ififoXdata[67]), .DO66(ififoXdata[66]),
 .DO65(ififoXdata[65]), .DO64(ififoXdata[64]), .DO63(ififoXdata[63]), .DO62(ififoXdata[62]), .DO61(ififoXdata[61]), .DO60(ififoXdata[60]), .DO59(ififoXdata[59]), .DO58(ififoXdata[58]),
 .DO57(ififoXdata[57]), .DO56(ififoXdata[56]), .DO55(ififoXdata[55]), .DO54(ififoXdata[54]), .DO53(ififoXdata[53]), .DO52(ififoXdata[52]), .DO51(ififoXdata[51]), .DO50(ififoXdata[50]),
 .DO49(ififoXdata[49]), .DO48(ififoXdata[48]), .DO47(ififoXdata[47]), .DO46(ififoXdata[46]), .DO45(ififoXdata[45]), .DO44(ififoXdata[44]), .DO43(ififoXdata[43]), .DO42(ififoXdata[42]),
 .DO41(ififoXdata[41]), .DO40(ififoXdata[40]), .DO39(ififoXdata[39]), .DO38(ififoXdata[38]), .DO37(ififoXdata[37]), .DO36(ififoXdata[36]), .DO35(ififoXdata[35]), .DO34(ififoXdata[34]),
 .DO33(ififoXdata[33]), .DO32(ififoXdata[32]), .DO31(ififoXdata[31]), .DO30(ififoXdata[30]), .DO29(ififoXdata[29]), .DO28(ififoXdata[28]), .DO27(ififoXdata[27]), .DO26(ififoXdata[26]),
 .DO25(ififoXdata[25]), .DO24(ififoXdata[24]), .DO23(ififoXdata[23]), .DO22(ififoXdata[22]), .DO21(ififoXdata[21]), .DO20(ififoXdata[20]), .DO19(ififoXdata[19]), .DO18(ififoXdata[18]),
 .DO17(ififoXdata[17]), .DO16(ififoXdata[16]), .DO15(ififoXdata[15]), .DO14(ififoXdata[14]), .DO13(ififoXdata[13]), .DO12(ififoXdata[12]), .DO11(ififoXdata[11]), .DO10(ififoXdata[10]),
 .DO9(ififoXdata[9]), .DO8(ififoXdata[8]), .DO7(ififoXdata[7]), .DO6(ififoXdata[6]), .DO5(ififoXdata[5]), .DO4(ififoXdata[4]), .DO3(ififoXdata[3]), .DO2(ififoXdata[2]),
 .DO1(ififoXdata[1]), .DO0(ififoXdata[0]), .SYNC_OUT(n9337));
MPR32KX256 U10464 ( .A14(ififoRaddr0[14]), .A13(ififoRaddr0[13]), .A12(ififoRaddr0[12]), .A11(ififoRaddr0[11]), .A10(ififoRaddr0[10]), .A9(ififoRaddr0[9]),
 .A8(ififoRaddr0[8]), .A7(ififoRaddr0[7]), .A6(ififoRaddr0[6]), .A5(ififoRaddr0[5]), .A4(ififoRaddr0[4]), .A3(ififoRaddr0[3]), .A2(ififoRaddr0[2]), .A1(ififoRaddr0[1]),
 .A0(ififoRaddr0[0]), .SYNC_IN(n9337), .DO255(ififoRdata[255]), .DO254(ififoRdata[254]), .DO253(ififoRdata[253]), .DO252(ififoRdata[252]), .DO251(ififoRdata[251]), .DO250(ififoRdata[250]),
 .DO249(ififoRdata[249]), .DO248(ififoRdata[248]), .DO247(ififoRdata[247]), .DO246(ififoRdata[246]), .DO245(ififoRdata[245]), .DO244(ififoRdata[244]), .DO243(ififoRdata[243]), .DO242(ififoRdata[242]),
 .DO241(ififoRdata[241]), .DO240(ififoRdata[240]), .DO239(ififoRdata[239]), .DO238(ififoRdata[238]), .DO237(ififoRdata[237]), .DO236(ififoRdata[236]), .DO235(ififoRdata[235]), .DO234(ififoRdata[234]),
 .DO233(ififoRdata[233]), .DO232(ififoRdata[232]), .DO231(ififoRdata[231]), .DO230(ififoRdata[230]), .DO229(ififoRdata[229]), .DO228(ififoRdata[228]), .DO227(ififoRdata[227]), .DO226(ififoRdata[226]),
 .DO225(ififoRdata[225]), .DO224(ififoRdata[224]), .DO223(ififoRdata[223]), .DO222(ififoRdata[222]), .DO221(ififoRdata[221]), .DO220(ififoRdata[220]), .DO219(ififoRdata[219]), .DO218(ififoRdata[218]),
 .DO217(ififoRdata[217]), .DO216(ififoRdata[216]), .DO215(ififoRdata[215]), .DO214(ififoRdata[214]), .DO213(ififoRdata[213]), .DO212(ififoRdata[212]), .DO211(ififoRdata[211]), .DO210(ififoRdata[210]),
 .DO209(ififoRdata[209]), .DO208(ififoRdata[208]), .DO207(ififoRdata[207]), .DO206(ififoRdata[206]), .DO205(ififoRdata[205]), .DO204(ififoRdata[204]), .DO203(ififoRdata[203]), .DO202(ififoRdata[202]),
 .DO201(ififoRdata[201]), .DO200(ififoRdata[200]), .DO199(ififoRdata[199]), .DO198(ififoRdata[198]), .DO197(ififoRdata[197]), .DO196(ififoRdata[196]), .DO195(ififoRdata[195]), .DO194(ififoRdata[194]),
 .DO193(ififoRdata[193]), .DO192(ififoRdata[192]), .DO191(ififoRdata[191]), .DO190(ififoRdata[190]), .DO189(ififoRdata[189]), .DO188(ififoRdata[188]), .DO187(ififoRdata[187]), .DO186(ififoRdata[186]),
 .DO185(ififoRdata[185]), .DO184(ififoRdata[184]), .DO183(ififoRdata[183]), .DO182(ififoRdata[182]), .DO181(ififoRdata[181]), .DO180(ififoRdata[180]), .DO179(ififoRdata[179]), .DO178(ififoRdata[178]),
 .DO177(ififoRdata[177]), .DO176(ififoRdata[176]), .DO175(ififoRdata[175]), .DO174(ififoRdata[174]), .DO173(ififoRdata[173]), .DO172(ififoRdata[172]), .DO171(ififoRdata[171]), .DO170(ififoRdata[170]),
 .DO169(ififoRdata[169]), .DO168(ififoRdata[168]), .DO167(ififoRdata[167]), .DO166(ififoRdata[166]), .DO165(ififoRdata[165]), .DO164(ififoRdata[164]), .DO163(ififoRdata[163]), .DO162(ififoRdata[162]),
 .DO161(ififoRdata[161]), .DO160(ififoRdata[160]), .DO159(ififoRdata[159]), .DO158(ififoRdata[158]), .DO157(ififoRdata[157]), .DO156(ififoRdata[156]), .DO155(ififoRdata[155]), .DO154(ififoRdata[154]),
 .DO153(ififoRdata[153]), .DO152(ififoRdata[152]), .DO151(ififoRdata[151]), .DO150(ififoRdata[150]), .DO149(ififoRdata[149]), .DO148(ififoRdata[148]), .DO147(ififoRdata[147]), .DO146(ififoRdata[146]),
 .DO145(ififoRdata[145]), .DO144(ififoRdata[144]), .DO143(ififoRdata[143]), .DO142(ififoRdata[142]), .DO141(ififoRdata[141]), .DO140(ififoRdata[140]), .DO139(ififoRdata[139]), .DO138(ififoRdata[138]),
 .DO137(ififoRdata[137]), .DO136(ififoRdata[136]), .DO135(ififoRdata[135]), .DO134(ififoRdata[134]), .DO133(ififoRdata[133]), .DO132(ififoRdata[132]), .DO131(ififoRdata[131]), .DO130(ififoRdata[130]),
 .DO129(ififoRdata[129]), .DO128(ififoRdata[128]), .DO127(ififoRdata[127]), .DO126(ififoRdata[126]), .DO125(ififoRdata[125]), .DO124(ififoRdata[124]), .DO123(ififoRdata[123]), .DO122(ififoRdata[122]),
 .DO121(ififoRdata[121]), .DO120(ififoRdata[120]), .DO119(ififoRdata[119]), .DO118(ififoRdata[118]), .DO117(ififoRdata[117]), .DO116(ififoRdata[116]), .DO115(ififoRdata[115]), .DO114(ififoRdata[114]),
 .DO113(ififoRdata[113]), .DO112(ififoRdata[112]), .DO111(ififoRdata[111]), .DO110(ififoRdata[110]), .DO109(ififoRdata[109]), .DO108(ififoRdata[108]), .DO107(ififoRdata[107]), .DO106(ififoRdata[106]),
 .DO105(ififoRdata[105]), .DO104(ififoRdata[104]), .DO103(ififoRdata[103]), .DO102(ififoRdata[102]), .DO101(ififoRdata[101]), .DO100(ififoRdata[100]), .DO99(ififoRdata[99]), .DO98(ififoRdata[98]),
 .DO97(ififoRdata[97]), .DO96(ififoRdata[96]), .DO95(ififoRdata[95]), .DO94(ififoRdata[94]), .DO93(ififoRdata[93]), .DO92(ififoRdata[92]), .DO91(ififoRdata[91]), .DO90(ififoRdata[90]),
 .DO89(ififoRdata[89]), .DO88(ififoRdata[88]), .DO87(ififoRdata[87]), .DO86(ififoRdata[86]), .DO85(ififoRdata[85]), .DO84(ififoRdata[84]), .DO83(ififoRdata[83]), .DO82(ififoRdata[82]),
 .DO81(ififoRdata[81]), .DO80(ififoRdata[80]), .DO79(ififoRdata[79]), .DO78(ififoRdata[78]), .DO77(ififoRdata[77]), .DO76(ififoRdata[76]), .DO75(ififoRdata[75]), .DO74(ififoRdata[74]),
 .DO73(ififoRdata[73]), .DO72(ififoRdata[72]), .DO71(ififoRdata[71]), .DO70(ififoRdata[70]), .DO69(ififoRdata[69]), .DO68(ififoRdata[68]), .DO67(ififoRdata[67]), .DO66(ififoRdata[66]),
 .DO65(ififoRdata[65]), .DO64(ififoRdata[64]), .DO63(ififoRdata[63]), .DO62(ififoRdata[62]), .DO61(ififoRdata[61]), .DO60(ififoRdata[60]), .DO59(ififoRdata[59]), .DO58(ififoRdata[58]),
 .DO57(ififoRdata[57]), .DO56(ififoRdata[56]), .DO55(ififoRdata[55]), .DO54(ififoRdata[54]), .DO53(ififoRdata[53]), .DO52(ififoRdata[52]), .DO51(ififoRdata[51]), .DO50(ififoRdata[50]),
 .DO49(ififoRdata[49]), .DO48(ififoRdata[48]), .DO47(ififoRdata[47]), .DO46(ififoRdata[46]), .DO45(ififoRdata[45]), .DO44(ififoRdata[44]), .DO43(ififoRdata[43]), .DO42(ififoRdata[42]),
 .DO41(ififoRdata[41]), .DO40(ififoRdata[40]), .DO39(ififoRdata[39]), .DO38(ififoRdata[38]), .DO37(ififoRdata[37]), .DO36(ififoRdata[36]), .DO35(ififoRdata[35]), .DO34(ififoRdata[34]),
 .DO33(ififoRdata[33]), .DO32(ififoRdata[32]), .DO31(ififoRdata[31]), .DO30(ififoRdata[30]), .DO29(ififoRdata[29]), .DO28(ififoRdata[28]), .DO27(ififoRdata[27]), .DO26(ififoRdata[26]),
 .DO25(ififoRdata[25]), .DO24(ififoRdata[24]), .DO23(ififoRdata[23]), .DO22(ififoRdata[22]), .DO21(ififoRdata[21]), .DO20(ififoRdata[20]), .DO19(ififoRdata[19]), .DO18(ififoRdata[18]),
 .DO17(ififoRdata[17]), .DO16(ififoRdata[16]), .DO15(ififoRdata[15]), .DO14(ififoRdata[14]), .DO13(ififoRdata[13]), .DO12(ififoRdata[12]), .DO11(ififoRdata[11]), .DO10(ififoRdata[10]),
 .DO9(ififoRdata[9]), .DO8(ififoRdata[8]), .DO7(ififoRdata[7]), .DO6(ififoRdata[6]), .DO5(ififoRdata[5]), .DO4(ififoRdata[4]), .DO3(ififoRdata[3]), .DO2(ififoRdata[2]),
 .DO1(ififoRdata[1]), .DO0(ififoRdata[0]), .SYNC_OUT(n9338));
MPR32KX256 U10465 ( .A14(ififoRaddr1[14]), .A13(ififoRaddr1[13]), .A12(ififoRaddr1[12]), .A11(ififoRaddr1[11]), .A10(ififoRaddr1[10]), .A9(ififoRaddr1[9]),
 .A8(ififoRaddr1[8]), .A7(ififoRaddr1[7]), .A6(ififoRaddr1[6]), .A5(ififoRaddr1[5]), .A4(ififoRaddr1[4]), .A3(ififoRaddr1[3]), .A2(ififoRaddr1[2]), .A1(ififoRaddr1[1]),
 .A0(ififoRaddr1[0]), .SYNC_IN(n9338), .DO255(ififoRdata[511]), .DO254(ififoRdata[510]), .DO253(ififoRdata[509]), .DO252(ififoRdata[508]), .DO251(ififoRdata[507]), .DO250(ififoRdata[506]),
 .DO249(ififoRdata[505]), .DO248(ififoRdata[504]), .DO247(ififoRdata[503]), .DO246(ififoRdata[502]), .DO245(ififoRdata[501]), .DO244(ififoRdata[500]), .DO243(ififoRdata[499]), .DO242(ififoRdata[498]),
 .DO241(ififoRdata[497]), .DO240(ififoRdata[496]), .DO239(ififoRdata[495]), .DO238(ififoRdata[494]), .DO237(ififoRdata[493]), .DO236(ififoRdata[492]), .DO235(ififoRdata[491]), .DO234(ififoRdata[490]),
 .DO233(ififoRdata[489]), .DO232(ififoRdata[488]), .DO231(ififoRdata[487]), .DO230(ififoRdata[486]), .DO229(ififoRdata[485]), .DO228(ififoRdata[484]), .DO227(ififoRdata[483]), .DO226(ififoRdata[482]),
 .DO225(ififoRdata[481]), .DO224(ififoRdata[480]), .DO223(ififoRdata[479]), .DO222(ififoRdata[478]), .DO221(ififoRdata[477]), .DO220(ififoRdata[476]), .DO219(ififoRdata[475]), .DO218(ififoRdata[474]),
 .DO217(ififoRdata[473]), .DO216(ififoRdata[472]), .DO215(ififoRdata[471]), .DO214(ififoRdata[470]), .DO213(ififoRdata[469]), .DO212(ififoRdata[468]), .DO211(ififoRdata[467]), .DO210(ififoRdata[466]),
 .DO209(ififoRdata[465]), .DO208(ififoRdata[464]), .DO207(ififoRdata[463]), .DO206(ififoRdata[462]), .DO205(ififoRdata[461]), .DO204(ififoRdata[460]), .DO203(ififoRdata[459]), .DO202(ififoRdata[458]),
 .DO201(ififoRdata[457]), .DO200(ififoRdata[456]), .DO199(ififoRdata[455]), .DO198(ififoRdata[454]), .DO197(ififoRdata[453]), .DO196(ififoRdata[452]), .DO195(ififoRdata[451]), .DO194(ififoRdata[450]),
 .DO193(ififoRdata[449]), .DO192(ififoRdata[448]), .DO191(ififoRdata[447]), .DO190(ififoRdata[446]), .DO189(ififoRdata[445]), .DO188(ififoRdata[444]), .DO187(ififoRdata[443]), .DO186(ififoRdata[442]),
 .DO185(ififoRdata[441]), .DO184(ififoRdata[440]), .DO183(ififoRdata[439]), .DO182(ififoRdata[438]), .DO181(ififoRdata[437]), .DO180(ififoRdata[436]), .DO179(ififoRdata[435]), .DO178(ififoRdata[434]),
 .DO177(ififoRdata[433]), .DO176(ififoRdata[432]), .DO175(ififoRdata[431]), .DO174(ififoRdata[430]), .DO173(ififoRdata[429]), .DO172(ififoRdata[428]), .DO171(ififoRdata[427]), .DO170(ififoRdata[426]),
 .DO169(ififoRdata[425]), .DO168(ififoRdata[424]), .DO167(ififoRdata[423]), .DO166(ififoRdata[422]), .DO165(ififoRdata[421]), .DO164(ififoRdata[420]), .DO163(ififoRdata[419]), .DO162(ififoRdata[418]),
 .DO161(ififoRdata[417]), .DO160(ififoRdata[416]), .DO159(ififoRdata[415]), .DO158(ififoRdata[414]), .DO157(ififoRdata[413]), .DO156(ififoRdata[412]), .DO155(ififoRdata[411]), .DO154(ififoRdata[410]),
 .DO153(ififoRdata[409]), .DO152(ififoRdata[408]), .DO151(ififoRdata[407]), .DO150(ififoRdata[406]), .DO149(ififoRdata[405]), .DO148(ififoRdata[404]), .DO147(ififoRdata[403]), .DO146(ififoRdata[402]),
 .DO145(ififoRdata[401]), .DO144(ififoRdata[400]), .DO143(ififoRdata[399]), .DO142(ififoRdata[398]), .DO141(ififoRdata[397]), .DO140(ififoRdata[396]), .DO139(ififoRdata[395]), .DO138(ififoRdata[394]),
 .DO137(ififoRdata[393]), .DO136(ififoRdata[392]), .DO135(ififoRdata[391]), .DO134(ififoRdata[390]), .DO133(ififoRdata[389]), .DO132(ififoRdata[388]), .DO131(ififoRdata[387]), .DO130(ififoRdata[386]),
 .DO129(ififoRdata[385]), .DO128(ififoRdata[384]), .DO127(ififoRdata[383]), .DO126(ififoRdata[382]), .DO125(ififoRdata[381]), .DO124(ififoRdata[380]), .DO123(ififoRdata[379]), .DO122(ififoRdata[378]),
 .DO121(ififoRdata[377]), .DO120(ififoRdata[376]), .DO119(ififoRdata[375]), .DO118(ififoRdata[374]), .DO117(ififoRdata[373]), .DO116(ififoRdata[372]), .DO115(ififoRdata[371]), .DO114(ififoRdata[370]),
 .DO113(ififoRdata[369]), .DO112(ififoRdata[368]), .DO111(ififoRdata[367]), .DO110(ififoRdata[366]), .DO109(ififoRdata[365]), .DO108(ififoRdata[364]), .DO107(ififoRdata[363]), .DO106(ififoRdata[362]),
 .DO105(ififoRdata[361]), .DO104(ififoRdata[360]), .DO103(ififoRdata[359]), .DO102(ififoRdata[358]), .DO101(ififoRdata[357]), .DO100(ififoRdata[356]), .DO99(ififoRdata[355]), .DO98(ififoRdata[354]),
 .DO97(ififoRdata[353]), .DO96(ififoRdata[352]), .DO95(ififoRdata[351]), .DO94(ififoRdata[350]), .DO93(ififoRdata[349]), .DO92(ififoRdata[348]), .DO91(ififoRdata[347]), .DO90(ififoRdata[346]),
 .DO89(ififoRdata[345]), .DO88(ififoRdata[344]), .DO87(ififoRdata[343]), .DO86(ififoRdata[342]), .DO85(ififoRdata[341]), .DO84(ififoRdata[340]), .DO83(ififoRdata[339]), .DO82(ififoRdata[338]),
 .DO81(ififoRdata[337]), .DO80(ififoRdata[336]), .DO79(ififoRdata[335]), .DO78(ififoRdata[334]), .DO77(ififoRdata[333]), .DO76(ififoRdata[332]), .DO75(ififoRdata[331]), .DO74(ififoRdata[330]),
 .DO73(ififoRdata[329]), .DO72(ififoRdata[328]), .DO71(ififoRdata[327]), .DO70(ififoRdata[326]), .DO69(ififoRdata[325]), .DO68(ififoRdata[324]), .DO67(ififoRdata[323]), .DO66(ififoRdata[322]),
 .DO65(ififoRdata[321]), .DO64(ififoRdata[320]), .DO63(ififoRdata[319]), .DO62(ififoRdata[318]), .DO61(ififoRdata[317]), .DO60(ififoRdata[316]), .DO59(ififoRdata[315]), .DO58(ififoRdata[314]),
 .DO57(ififoRdata[313]), .DO56(ififoRdata[312]), .DO55(ififoRdata[311]), .DO54(ififoRdata[310]), .DO53(ififoRdata[309]), .DO52(ififoRdata[308]), .DO51(ififoRdata[307]), .DO50(ififoRdata[306]),
 .DO49(ififoRdata[305]), .DO48(ififoRdata[304]), .DO47(ififoRdata[303]), .DO46(ififoRdata[302]), .DO45(ififoRdata[301]), .DO44(ififoRdata[300]), .DO43(ififoRdata[299]), .DO42(ififoRdata[298]),
 .DO41(ififoRdata[297]), .DO40(ififoRdata[296]), .DO39(ififoRdata[295]), .DO38(ififoRdata[294]), .DO37(ififoRdata[293]), .DO36(ififoRdata[292]), .DO35(ififoRdata[291]), .DO34(ififoRdata[290]),
 .DO33(ififoRdata[289]), .DO32(ififoRdata[288]), .DO31(ififoRdata[287]), .DO30(ififoRdata[286]), .DO29(ififoRdata[285]), .DO28(ififoRdata[284]), .DO27(ififoRdata[283]), .DO26(ififoRdata[282]),
 .DO25(ififoRdata[281]), .DO24(ififoRdata[280]), .DO23(ififoRdata[279]), .DO22(ififoRdata[278]), .DO21(ififoRdata[277]), .DO20(ififoRdata[276]), .DO19(ififoRdata[275]), .DO18(ififoRdata[274]),
 .DO17(ififoRdata[273]), .DO16(ififoRdata[272]), .DO15(ififoRdata[271]), .DO14(ififoRdata[270]), .DO13(ififoRdata[269]), .DO12(ififoRdata[268]), .DO11(ififoRdata[267]), .DO10(ififoRdata[266]),
 .DO9(ififoRdata[265]), .DO8(ififoRdata[264]), .DO7(ififoRdata[263]), .DO6(ififoRdata[262]), .DO5(ififoRdata[261]), .DO4(ififoRdata[260]), .DO3(ififoRdata[259]), .DO2(ififoRdata[258]),
 .DO1(ififoRdata[257]), .DO0(ififoRdata[256]), .SYNC_OUT(n9339));
MPR32KX256 U10466 ( .A14(ififoRaddr2[14]), .A13(ififoRaddr2[13]), .A12(ififoRaddr2[12]), .A11(ififoRaddr2[11]), .A10(ififoRaddr2[10]), .A9(ififoRaddr2[9]),
 .A8(ififoRaddr2[8]), .A7(ififoRaddr2[7]), .A6(ififoRaddr2[6]), .A5(ififoRaddr2[5]), .A4(ififoRaddr2[4]), .A3(ififoRaddr2[3]), .A2(ififoRaddr2[2]), .A1(ififoRaddr2[1]),
 .A0(ififoRaddr2[0]), .SYNC_IN(n9339), .DO255(ififoRdata[767]), .DO254(ififoRdata[766]), .DO253(ififoRdata[765]), .DO252(ififoRdata[764]), .DO251(ififoRdata[763]), .DO250(ififoRdata[762]),
 .DO249(ififoRdata[761]), .DO248(ififoRdata[760]), .DO247(ififoRdata[759]), .DO246(ififoRdata[758]), .DO245(ififoRdata[757]), .DO244(ififoRdata[756]), .DO243(ififoRdata[755]), .DO242(ififoRdata[754]),
 .DO241(ififoRdata[753]), .DO240(ififoRdata[752]), .DO239(ififoRdata[751]), .DO238(ififoRdata[750]), .DO237(ififoRdata[749]), .DO236(ififoRdata[748]), .DO235(ififoRdata[747]), .DO234(ififoRdata[746]),
 .DO233(ififoRdata[745]), .DO232(ififoRdata[744]), .DO231(ififoRdata[743]), .DO230(ififoRdata[742]), .DO229(ififoRdata[741]), .DO228(ififoRdata[740]), .DO227(ififoRdata[739]), .DO226(ififoRdata[738]),
 .DO225(ififoRdata[737]), .DO224(ififoRdata[736]), .DO223(ififoRdata[735]), .DO222(ififoRdata[734]), .DO221(ififoRdata[733]), .DO220(ififoRdata[732]), .DO219(ififoRdata[731]), .DO218(ififoRdata[730]),
 .DO217(ififoRdata[729]), .DO216(ififoRdata[728]), .DO215(ififoRdata[727]), .DO214(ififoRdata[726]), .DO213(ififoRdata[725]), .DO212(ififoRdata[724]), .DO211(ififoRdata[723]), .DO210(ififoRdata[722]),
 .DO209(ififoRdata[721]), .DO208(ififoRdata[720]), .DO207(ififoRdata[719]), .DO206(ififoRdata[718]), .DO205(ififoRdata[717]), .DO204(ififoRdata[716]), .DO203(ififoRdata[715]), .DO202(ififoRdata[714]),
 .DO201(ififoRdata[713]), .DO200(ififoRdata[712]), .DO199(ififoRdata[711]), .DO198(ififoRdata[710]), .DO197(ififoRdata[709]), .DO196(ififoRdata[708]), .DO195(ififoRdata[707]), .DO194(ififoRdata[706]),
 .DO193(ififoRdata[705]), .DO192(ififoRdata[704]), .DO191(ififoRdata[703]), .DO190(ififoRdata[702]), .DO189(ififoRdata[701]), .DO188(ififoRdata[700]), .DO187(ififoRdata[699]), .DO186(ififoRdata[698]),
 .DO185(ififoRdata[697]), .DO184(ififoRdata[696]), .DO183(ififoRdata[695]), .DO182(ififoRdata[694]), .DO181(ififoRdata[693]), .DO180(ififoRdata[692]), .DO179(ififoRdata[691]), .DO178(ififoRdata[690]),
 .DO177(ififoRdata[689]), .DO176(ififoRdata[688]), .DO175(ififoRdata[687]), .DO174(ififoRdata[686]), .DO173(ififoRdata[685]), .DO172(ififoRdata[684]), .DO171(ififoRdata[683]), .DO170(ififoRdata[682]),
 .DO169(ififoRdata[681]), .DO168(ififoRdata[680]), .DO167(ififoRdata[679]), .DO166(ififoRdata[678]), .DO165(ififoRdata[677]), .DO164(ififoRdata[676]), .DO163(ififoRdata[675]), .DO162(ififoRdata[674]),
 .DO161(ififoRdata[673]), .DO160(ififoRdata[672]), .DO159(ififoRdata[671]), .DO158(ififoRdata[670]), .DO157(ififoRdata[669]), .DO156(ififoRdata[668]), .DO155(ififoRdata[667]), .DO154(ififoRdata[666]),
 .DO153(ififoRdata[665]), .DO152(ififoRdata[664]), .DO151(ififoRdata[663]), .DO150(ififoRdata[662]), .DO149(ififoRdata[661]), .DO148(ififoRdata[660]), .DO147(ififoRdata[659]), .DO146(ififoRdata[658]),
 .DO145(ififoRdata[657]), .DO144(ififoRdata[656]), .DO143(ififoRdata[655]), .DO142(ififoRdata[654]), .DO141(ififoRdata[653]), .DO140(ififoRdata[652]), .DO139(ififoRdata[651]), .DO138(ififoRdata[650]),
 .DO137(ififoRdata[649]), .DO136(ififoRdata[648]), .DO135(ififoRdata[647]), .DO134(ififoRdata[646]), .DO133(ififoRdata[645]), .DO132(ififoRdata[644]), .DO131(ififoRdata[643]), .DO130(ififoRdata[642]),
 .DO129(ififoRdata[641]), .DO128(ififoRdata[640]), .DO127(ififoRdata[639]), .DO126(ififoRdata[638]), .DO125(ififoRdata[637]), .DO124(ififoRdata[636]), .DO123(ififoRdata[635]), .DO122(ififoRdata[634]),
 .DO121(ififoRdata[633]), .DO120(ififoRdata[632]), .DO119(ififoRdata[631]), .DO118(ififoRdata[630]), .DO117(ififoRdata[629]), .DO116(ififoRdata[628]), .DO115(ififoRdata[627]), .DO114(ififoRdata[626]),
 .DO113(ififoRdata[625]), .DO112(ififoRdata[624]), .DO111(ififoRdata[623]), .DO110(ififoRdata[622]), .DO109(ififoRdata[621]), .DO108(ififoRdata[620]), .DO107(ififoRdata[619]), .DO106(ififoRdata[618]),
 .DO105(ififoRdata[617]), .DO104(ififoRdata[616]), .DO103(ififoRdata[615]), .DO102(ififoRdata[614]), .DO101(ififoRdata[613]), .DO100(ififoRdata[612]), .DO99(ififoRdata[611]), .DO98(ififoRdata[610]),
 .DO97(ififoRdata[609]), .DO96(ififoRdata[608]), .DO95(ififoRdata[607]), .DO94(ififoRdata[606]), .DO93(ififoRdata[605]), .DO92(ififoRdata[604]), .DO91(ififoRdata[603]), .DO90(ififoRdata[602]),
 .DO89(ififoRdata[601]), .DO88(ififoRdata[600]), .DO87(ififoRdata[599]), .DO86(ififoRdata[598]), .DO85(ififoRdata[597]), .DO84(ififoRdata[596]), .DO83(ififoRdata[595]), .DO82(ififoRdata[594]),
 .DO81(ififoRdata[593]), .DO80(ififoRdata[592]), .DO79(ififoRdata[591]), .DO78(ififoRdata[590]), .DO77(ififoRdata[589]), .DO76(ififoRdata[588]), .DO75(ififoRdata[587]), .DO74(ififoRdata[586]),
 .DO73(ififoRdata[585]), .DO72(ififoRdata[584]), .DO71(ififoRdata[583]), .DO70(ififoRdata[582]), .DO69(ififoRdata[581]), .DO68(ififoRdata[580]), .DO67(ififoRdata[579]), .DO66(ififoRdata[578]),
 .DO65(ififoRdata[577]), .DO64(ififoRdata[576]), .DO63(ififoRdata[575]), .DO62(ififoRdata[574]), .DO61(ififoRdata[573]), .DO60(ififoRdata[572]), .DO59(ififoRdata[571]), .DO58(ififoRdata[570]),
 .DO57(ififoRdata[569]), .DO56(ififoRdata[568]), .DO55(ififoRdata[567]), .DO54(ififoRdata[566]), .DO53(ififoRdata[565]), .DO52(ififoRdata[564]), .DO51(ififoRdata[563]), .DO50(ififoRdata[562]),
 .DO49(ififoRdata[561]), .DO48(ififoRdata[560]), .DO47(ififoRdata[559]), .DO46(ififoRdata[558]), .DO45(ififoRdata[557]), .DO44(ififoRdata[556]), .DO43(ififoRdata[555]), .DO42(ififoRdata[554]),
 .DO41(ififoRdata[553]), .DO40(ififoRdata[552]), .DO39(ififoRdata[551]), .DO38(ififoRdata[550]), .DO37(ififoRdata[549]), .DO36(ififoRdata[548]), .DO35(ififoRdata[547]), .DO34(ififoRdata[546]),
 .DO33(ififoRdata[545]), .DO32(ififoRdata[544]), .DO31(ififoRdata[543]), .DO30(ififoRdata[542]), .DO29(ififoRdata[541]), .DO28(ififoRdata[540]), .DO27(ififoRdata[539]), .DO26(ififoRdata[538]),
 .DO25(ififoRdata[537]), .DO24(ififoRdata[536]), .DO23(ififoRdata[535]), .DO22(ififoRdata[534]), .DO21(ififoRdata[533]), .DO20(ififoRdata[532]), .DO19(ififoRdata[531]), .DO18(ififoRdata[530]),
 .DO17(ififoRdata[529]), .DO16(ififoRdata[528]), .DO15(ififoRdata[527]), .DO14(ififoRdata[526]), .DO13(ififoRdata[525]), .DO12(ififoRdata[524]), .DO11(ififoRdata[523]), .DO10(ififoRdata[522]),
 .DO9(ififoRdata[521]), .DO8(ififoRdata[520]), .DO7(ififoRdata[519]), .DO6(ififoRdata[518]), .DO5(ififoRdata[517]), .DO4(ififoRdata[516]), .DO3(ififoRdata[515]), .DO2(ififoRdata[514]),
 .DO1(ififoRdata[513]), .DO0(ififoRdata[512]), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "ixc_gfm_ififo 1 255 0 0 32767"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "ixc_gfm_ofifo 1 255 0 0 32767"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "2"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW32KX256_MPR32KX256
`else
module MPW32KX256( A14, A13, A12, A11, A10, A9, A8,
 A7, A6, A5, A4, A3, A2, A1, A0,
 DI255, DI254, DI253, DI252, DI251, DI250, DI249, DI248,
 DI247, DI246, DI245, DI244, DI243, DI242, DI241, DI240,
 DI239, DI238, DI237, DI236, DI235, DI234, DI233, DI232,
 DI231, DI230, DI229, DI228, DI227, DI226, DI225, DI224,
 DI223, DI222, DI221, DI220, DI219, DI218, DI217, DI216,
 DI215, DI214, DI213, DI212, DI211, DI210, DI209, DI208,
 DI207, DI206, DI205, DI204, DI203, DI202, DI201, DI200,
 DI199, DI198, DI197, DI196, DI195, DI194, DI193, DI192,
 DI191, DI190, DI189, DI188, DI187, DI186, DI185, DI184,
 DI183, DI182, DI181, DI180, DI179, DI178, DI177, DI176,
 DI175, DI174, DI173, DI172, DI171, DI170, DI169, DI168,
 DI167, DI166, DI165, DI164, DI163, DI162, DI161, DI160,
 DI159, DI158, DI157, DI156, DI155, DI154, DI153, DI152,
 DI151, DI150, DI149, DI148, DI147, DI146, DI145, DI144,
 DI143, DI142, DI141, DI140, DI139, DI138, DI137, DI136,
 DI135, DI134, DI133, DI132, DI131, DI130, DI129, DI128,
 DI127, DI126, DI125, DI124, DI123, DI122, DI121, DI120,
 DI119, DI118, DI117, DI116, DI115, DI114, DI113, DI112,
 DI111, DI110, DI109, DI108, DI107, DI106, DI105, DI104,
 DI103, DI102, DI101, DI100, DI99, DI98, DI97, DI96,
 DI95, DI94, DI93, DI92, DI91, DI90, DI89, DI88,
 DI87, DI86, DI85, DI84, DI83, DI82, DI81, DI80,
 DI79, DI78, DI77, DI76, DI75, DI74, DI73, DI72,
 DI71, DI70, DI69, DI68, DI67, DI66, DI65, DI64,
 DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56,
 DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48,
 DI47, DI46, DI45, DI44, DI43, DI42, DI41, DI40,
 DI39, DI38, DI37, DI36, DI35, DI34, DI33, DI32,
 DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24,
 DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16,
 DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8,
 DI7, DI6, DI5, DI4, DI3, DI2, DI1, DI0,
 WE, SYNC_IN, SYNC_OUT);
input  A14, A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, DI255, DI254, DI253,
 DI252, DI251, DI250, DI249, DI248, DI247, DI246, DI245, DI244, DI243,
 DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235, DI234, DI233,
 DI232, DI231, DI230, DI229, DI228, DI227, DI226, DI225, DI224, DI223,
 DI222, DI221, DI220, DI219, DI218, DI217, DI216, DI215, DI214, DI213,
 DI212, DI211, DI210, DI209, DI208, DI207, DI206, DI205, DI204, DI203,
 DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195, DI194, DI193,
 DI192, DI191, DI190, DI189, DI188, DI187, DI186, DI185, DI184, DI183,
 DI182, DI181, DI180, DI179, DI178, DI177, DI176, DI175, DI174, DI173,
 DI172, DI171, DI170, DI169, DI168, DI167, DI166, DI165, DI164, DI163,
 DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155, DI154, DI153,
 DI152, DI151, DI150, DI149, DI148, DI147, DI146, DI145, DI144, DI143,
 DI142, DI141, DI140, DI139, DI138, DI137, DI136, DI135, DI134, DI133,
 DI132, DI131, DI130, DI129, DI128, DI127, DI126, DI125, DI124, DI123,
 DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115, DI114, DI113,
 DI112, DI111, DI110, DI109, DI108, DI107, DI106, DI105, DI104, DI103,
 DI102, DI101, DI100, DI99, DI98, DI97, DI96, DI95, DI94, DI93,
 DI92, DI91, DI90, DI89, DI88, DI87, DI86, DI85, DI84, DI83,
 DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75, DI74, DI73,
 DI72, DI71, DI70, DI69, DI68, DI67, DI66, DI65, DI64, DI63,
 DI62, DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54, DI53,
 DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34, DI33,
 DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24, DI23,
 DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR32KX256_
`else
module MPR32KX256( A14, A13, A12, A11, A10, A9, A8,
 A7, A6, A5, A4, A3, A2, A1, A0,
 SYNC_IN, DO255, DO254, DO253, DO252, DO251, DO250, DO249,
 DO248, DO247, DO246, DO245, DO244, DO243, DO242, DO241,
 DO240, DO239, DO238, DO237, DO236, DO235, DO234, DO233,
 DO232, DO231, DO230, DO229, DO228, DO227, DO226, DO225,
 DO224, DO223, DO222, DO221, DO220, DO219, DO218, DO217,
 DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209,
 DO208, DO207, DO206, DO205, DO204, DO203, DO202, DO201,
 DO200, DO199, DO198, DO197, DO196, DO195, DO194, DO193,
 DO192, DO191, DO190, DO189, DO188, DO187, DO186, DO185,
 DO184, DO183, DO182, DO181, DO180, DO179, DO178, DO177,
 DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169,
 DO168, DO167, DO166, DO165, DO164, DO163, DO162, DO161,
 DO160, DO159, DO158, DO157, DO156, DO155, DO154, DO153,
 DO152, DO151, DO150, DO149, DO148, DO147, DO146, DO145,
 DO144, DO143, DO142, DO141, DO140, DO139, DO138, DO137,
 DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129,
 DO128, DO127, DO126, DO125, DO124, DO123, DO122, DO121,
 DO120, DO119, DO118, DO117, DO116, DO115, DO114, DO113,
 DO112, DO111, DO110, DO109, DO108, DO107, DO106, DO105,
 DO104, DO103, DO102, DO101, DO100, DO99, DO98, DO97,
 DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89,
 DO88, DO87, DO86, DO85, DO84, DO83, DO82, DO81,
 DO80, DO79, DO78, DO77, DO76, DO75, DO74, DO73,
 DO72, DO71, DO70, DO69, DO68, DO67, DO66, DO65,
 DO64, DO63, DO62, DO61, DO60, DO59, DO58, DO57,
 DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49,
 DO48, DO47, DO46, DO45, DO44, DO43, DO42, DO41,
 DO40, DO39, DO38, DO37, DO36, DO35, DO34, DO33,
 DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25,
 DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17,
 DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9,
 DO8, DO7, DO6, DO5, DO4, DO3, DO2, DO1,
 DO0, SYNC_OUT);
input  A14, A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, SYNC_IN;
output  DO255, DO254, DO253, DO252, DO251, DO250, DO249, DO248,
 DO247, DO246, DO245, DO244, DO243, DO242, DO241, DO240, DO239, DO238,
 DO237, DO236, DO235, DO234, DO233, DO232, DO231, DO230, DO229, DO228,
 DO227, DO226, DO225, DO224, DO223, DO222, DO221, DO220, DO219, DO218,
 DO217, DO216, DO215, DO214, DO213, DO212, DO211, DO210, DO209, DO208,
 DO207, DO206, DO205, DO204, DO203, DO202, DO201, DO200, DO199, DO198,
 DO197, DO196, DO195, DO194, DO193, DO192, DO191, DO190, DO189, DO188,
 DO187, DO186, DO185, DO184, DO183, DO182, DO181, DO180, DO179, DO178,
 DO177, DO176, DO175, DO174, DO173, DO172, DO171, DO170, DO169, DO168,
 DO167, DO166, DO165, DO164, DO163, DO162, DO161, DO160, DO159, DO158,
 DO157, DO156, DO155, DO154, DO153, DO152, DO151, DO150, DO149, DO148,
 DO147, DO146, DO145, DO144, DO143, DO142, DO141, DO140, DO139, DO138,
 DO137, DO136, DO135, DO134, DO133, DO132, DO131, DO130, DO129, DO128,
 DO127, DO126, DO125, DO124, DO123, DO122, DO121, DO120, DO119, DO118,
 DO117, DO116, DO115, DO114, DO113, DO112, DO111, DO110, DO109, DO108,
 DO107, DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99, DO98,
 DO97, DO96, DO95, DO94, DO93, DO92, DO91, DO90, DO89, DO88,
 DO87, DO86, DO85, DO84, DO83, DO82, DO81, DO80, DO79, DO78,
 DO77, DO76, DO75, DO74, DO73, DO72, DO71, DO70, DO69, DO68,
 DO67, DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59, DO58,
 DO57, DO56, DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48,
 DO47, DO46, DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28,
 DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18,
 DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8,
 DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR32KX256_
`endif
`define MPW32KX256_MPR32KX256
`endif
`endif
