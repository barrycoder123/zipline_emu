architecture module of ixc_asgn_ecov_rst_pulse is
  -- quickturn CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
  signal DUMMY0 : std_logic ;

begin
  rstsig <= DUMMY0 ;
end module;
