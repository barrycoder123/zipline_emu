
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_credit_manager ( credit_available, .hw_status( {\hw_status.used_err , 
	\hw_status.return_err , \hw_status.credit_issued [9], 
	\hw_status.credit_issued [8], \hw_status.credit_issued [7], 
	\hw_status.credit_issued [6], \hw_status.credit_issued [5], 
	\hw_status.credit_issued [4], \hw_status.credit_issued [3], 
	\hw_status.credit_issued [2], \hw_status.credit_issued [1], 
	\hw_status.credit_issued [0]} ), clk, rst_n, sw_init, credit_return, 
	credit_used, .sw_config( {\sw_config.dis_used , 
	\sw_config.dis_return , \sw_config.credit_limit [9], 
	\sw_config.credit_limit [8], \sw_config.credit_limit [7], 
	\sw_config.credit_limit [6], \sw_config.credit_limit [5], 
	\sw_config.credit_limit [4], \sw_config.credit_limit [3], 
	\sw_config.credit_limit [2], \sw_config.credit_limit [1], 
	\sw_config.credit_limit [0]} ));
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [8:0] credit_available;
output \hw_status.used_err ;
output \hw_status.return_err ;
output [9:0] \hw_status.credit_issued ;
wire [11:0] hw_status;
input clk;
input rst_n;
input sw_init;
input [8:0] credit_return;
input [8:0] credit_used;
input \sw_config.dis_used ;
input \sw_config.dis_return ;
input [9:0] \sw_config.credit_limit ;
wire [11:0] sw_config;
wire [0:8] _zy_simnet_credit_available_0_w$;
wire [0:11] _zy_simnet_hw_status_1_w$;
wire _zy_sva_b0_t;
wire _zy_sva_b1_t;
wire _zy_sva_b2_t;
wire _zyixc_port_1_0_s2hW;
wire _zyixc_port_1_1_s2hW;
wire [9:0] credit_issued_r;
wire used_err_v;
wire return_err_v;
wire [9:0] credit_issued_v;
wire [9:0] remaining_credit_v;
wire [31:0] outstanding;
wire credit_decrease;
wire [9:0] credit_limit;
`_2_ wire _zy_sva_b0;
`_2_ wire _zy_sva_b1;
`_2_ wire [0:0] _zy_sva_credit_return_check_1_0_fail;
`_2_ wire _zy_sva_b2;
`_2_ wire [0:0] _zy_sva_credit_danger_check_2_3_fail;
`_2_ wire _zyixc_port_1_0_req;
`_2_ wire _zyixc_port_1_0_ack;
`_2_ wire _zyixc_port_1_0_isf;
`_2_ wire _zyixc_port_1_0_osf;
`_2_ wire _zyixc_port_1_1_req;
`_2_ wire _zyixc_port_1_1_ack;
`_2_ wire _zyixc_port_1_1_isf;
`_2_ wire _zyixc_port_1_1_osf;
supply0 n234;
supply0 n405;
supply0 n406;
supply0 n407;
supply0 n408;
supply0 n409;
supply0 n410;
tran (hw_status[11], \hw_status.used_err );
tran (hw_status[10], \hw_status.return_err );
tran (hw_status[9], \hw_status.credit_issued [9]);
tran (hw_status[8], \hw_status.credit_issued [8]);
tran (hw_status[7], \hw_status.credit_issued [7]);
tran (hw_status[6], \hw_status.credit_issued [6]);
tran (hw_status[5], \hw_status.credit_issued [5]);
tran (hw_status[4], \hw_status.credit_issued [4]);
tran (hw_status[3], \hw_status.credit_issued [3]);
tran (hw_status[2], \hw_status.credit_issued [2]);
tran (hw_status[1], \hw_status.credit_issued [1]);
tran (hw_status[0], \hw_status.credit_issued [0]);
tran (sw_config[11], \sw_config.dis_used );
tran (sw_config[10], \sw_config.dis_return );
tran (sw_config[9], \sw_config.credit_limit [9]);
tran (sw_config[8], \sw_config.credit_limit [8]);
tran (sw_config[7], \sw_config.credit_limit [7]);
tran (sw_config[6], \sw_config.credit_limit [6]);
tran (sw_config[5], \sw_config.credit_limit [5]);
tran (sw_config[4], \sw_config.credit_limit [4]);
tran (sw_config[3], \sw_config.credit_limit [3]);
tran (sw_config[2], \sw_config.credit_limit [2]);
tran (sw_config[1], \sw_config.credit_limit [1]);
tran (sw_config[0], \sw_config.credit_limit [0]);
Q_OA21 U0 ( .A0(sw_config[0]), .A1(sw_config[1]), .B0(sw_config[9]), .Z(n412));
Q_OA21 U1 ( .A0(remaining_credit_v[0]), .A1(remaining_credit_v[1]), .B0(remaining_credit_v[8]), .Z(n25));
Q_INV U2 ( .A(sw_init), .Z(n1));
Q_FDP1 \credit_issued_r_REG[0] ( .CK(clk), .R(rst_n), .D(n13), .Q(credit_issued_r[0]), .QN(n204));
Q_FDP1 \credit_issued_r_REG[1] ( .CK(clk), .R(rst_n), .D(n12), .Q(credit_issued_r[1]), .QN(n207));
Q_FDP1 \credit_issued_r_REG[2] ( .CK(clk), .R(rst_n), .D(n11), .Q(credit_issued_r[2]), .QN(n214));
Q_FDP1 \credit_issued_r_REG[3] ( .CK(clk), .R(rst_n), .D(n10), .Q(credit_issued_r[3]), .QN(n216));
Q_FDP1 \credit_issued_r_REG[4] ( .CK(clk), .R(rst_n), .D(n9), .Q(credit_issued_r[4]), .QN(n218));
Q_FDP1 \credit_issued_r_REG[5] ( .CK(clk), .R(rst_n), .D(n8), .Q(credit_issued_r[5]), .QN(n221));
Q_FDP1 \credit_issued_r_REG[6] ( .CK(clk), .R(rst_n), .D(n7), .Q(credit_issued_r[6]), .QN(n228));
Q_FDP1 \credit_issued_r_REG[7] ( .CK(clk), .R(rst_n), .D(n6), .Q(credit_issued_r[7]), .QN(n230));
Q_FDP1 \credit_issued_r_REG[8] ( .CK(clk), .R(rst_n), .D(n5), .Q(credit_issued_r[8]), .QN(n232));
Q_FDP1 \credit_issued_r_REG[9] ( .CK(clk), .R(rst_n), .D(n4), .Q(credit_issued_r[9]), .QN(n233));
Q_FDP1 \hw_status_REG[0] ( .CK(clk), .R(rst_n), .D(n13), .Q(hw_status[0]), .QN( ));
Q_FDP1 \hw_status_REG[1] ( .CK(clk), .R(rst_n), .D(n12), .Q(hw_status[1]), .QN( ));
Q_FDP1 \hw_status_REG[2] ( .CK(clk), .R(rst_n), .D(n11), .Q(hw_status[2]), .QN( ));
Q_FDP1 \hw_status_REG[3] ( .CK(clk), .R(rst_n), .D(n10), .Q(hw_status[3]), .QN( ));
Q_FDP1 \hw_status_REG[4] ( .CK(clk), .R(rst_n), .D(n9), .Q(hw_status[4]), .QN( ));
Q_FDP1 \hw_status_REG[5] ( .CK(clk), .R(rst_n), .D(n8), .Q(hw_status[5]), .QN( ));
Q_FDP1 \hw_status_REG[6] ( .CK(clk), .R(rst_n), .D(n7), .Q(hw_status[6]), .QN( ));
Q_FDP1 \hw_status_REG[7] ( .CK(clk), .R(rst_n), .D(n6), .Q(hw_status[7]), .QN( ));
Q_FDP1 \hw_status_REG[8] ( .CK(clk), .R(rst_n), .D(n5), .Q(hw_status[8]), .QN( ));
Q_FDP1 \hw_status_REG[9] ( .CK(clk), .R(rst_n), .D(n4), .Q(hw_status[9]), .QN( ));
Q_FDP1 \hw_status_REG[10] ( .CK(clk), .R(rst_n), .D(n3), .Q(hw_status[10]), .QN( ));
Q_FDP1 \hw_status_REG[11] ( .CK(clk), .R(rst_n), .D(n2), .Q(hw_status[11]), .QN( ));
Q_AN02 U25 ( .A0(n1), .A1(credit_issued_v[9]), .Z(n4));
Q_AN02 U26 ( .A0(n1), .A1(credit_issued_v[8]), .Z(n5));
Q_AN02 U27 ( .A0(n1), .A1(credit_issued_v[7]), .Z(n6));
Q_AN02 U28 ( .A0(n1), .A1(credit_issued_v[6]), .Z(n7));
Q_AN02 U29 ( .A0(n1), .A1(credit_issued_v[5]), .Z(n8));
Q_AN02 U30 ( .A0(n1), .A1(credit_issued_v[4]), .Z(n9));
Q_AN02 U31 ( .A0(n1), .A1(credit_issued_v[3]), .Z(n10));
Q_AN02 U32 ( .A0(n1), .A1(credit_issued_v[2]), .Z(n11));
Q_AN02 U33 ( .A0(n1), .A1(credit_issued_v[1]), .Z(n12));
Q_AN02 U34 ( .A0(n1), .A1(credit_issued_v[0]), .Z(n13));
Q_AN03 U35 ( .A0(n15), .A1(n14), .A2(n1), .Z(n3));
Q_OR02 U36 ( .A0(hw_status[10]), .A1(return_err_v), .Z(n14));
Q_INV U37 ( .A(sw_config[10]), .Z(n15));
Q_AN03 U38 ( .A0(n17), .A1(n16), .A2(n1), .Z(n2));
Q_OR02 U39 ( .A0(hw_status[11]), .A1(used_err_v), .Z(n16));
Q_INV U40 ( .A(sw_config[11]), .Z(n17));
Q_INV U41 ( .A(n18), .Z(n20));
Q_OA21 U42 ( .A0(n18), .A1(remaining_credit_v[8]), .B0(n19), .Z(credit_available[8]));
Q_AN03 U43 ( .A0(n20), .A1(remaining_credit_v[7]), .A2(n19), .Z(credit_available[7]));
Q_AN03 U44 ( .A0(n20), .A1(remaining_credit_v[6]), .A2(n19), .Z(credit_available[6]));
Q_AN03 U45 ( .A0(n20), .A1(remaining_credit_v[5]), .A2(n19), .Z(credit_available[5]));
Q_AN03 U46 ( .A0(n20), .A1(remaining_credit_v[4]), .A2(n19), .Z(credit_available[4]));
Q_AN03 U47 ( .A0(n20), .A1(remaining_credit_v[3]), .A2(n19), .Z(credit_available[3]));
Q_AN03 U48 ( .A0(n20), .A1(remaining_credit_v[2]), .A2(n19), .Z(credit_available[2]));
Q_AN03 U49 ( .A0(n20), .A1(remaining_credit_v[1]), .A2(n19), .Z(credit_available[1]));
Q_AN03 U50 ( .A0(n20), .A1(remaining_credit_v[0]), .A2(n19), .Z(credit_available[0]));
Q_OR03 U51 ( .A0(n28), .A1(n24), .A2(n25), .Z(n18));
Q_OA21 U52 ( .A0(n26), .A1(n27), .B0(remaining_credit_v[8]), .Z(n24));
Q_OR02 U53 ( .A0(remaining_credit_v[5]), .A1(remaining_credit_v[4]), .Z(n26));
Q_OR02 U54 ( .A0(remaining_credit_v[3]), .A1(remaining_credit_v[2]), .Z(n27));
Q_AO21 U55 ( .A0(remaining_credit_v[8]), .A1(n29), .B0(remaining_credit_v[9]), .Z(n28));
Q_OR02 U56 ( .A0(remaining_credit_v[7]), .A1(remaining_credit_v[6]), .Z(n29));
Q_OR02 U57 ( .A0(remaining_credit_v[9]), .A1(n30), .Z(n19));
Q_OR03 U58 ( .A0(remaining_credit_v[7]), .A1(n31), .A2(remaining_credit_v[8]), .Z(n30));
Q_OR03 U59 ( .A0(remaining_credit_v[5]), .A1(n32), .A2(remaining_credit_v[6]), .Z(n31));
Q_OR03 U60 ( .A0(remaining_credit_v[3]), .A1(n33), .A2(remaining_credit_v[4]), .Z(n32));
Q_OR03 U61 ( .A0(remaining_credit_v[0]), .A1(remaining_credit_v[1]), .A2(remaining_credit_v[2]), .Z(n33));
Q_AN02 U62 ( .A0(n21), .A1(n34), .Z(remaining_credit_v[9]));
Q_AN02 U63 ( .A0(n21), .A1(n36), .Z(remaining_credit_v[8]));
Q_AN02 U64 ( .A0(n21), .A1(n37), .Z(remaining_credit_v[7]));
Q_AN02 U65 ( .A0(n21), .A1(n39), .Z(remaining_credit_v[6]));
Q_AN02 U66 ( .A0(n21), .A1(n40), .Z(remaining_credit_v[5]));
Q_AN02 U67 ( .A0(n21), .A1(n42), .Z(remaining_credit_v[4]));
Q_AN02 U68 ( .A0(n21), .A1(n43), .Z(remaining_credit_v[3]));
Q_AN02 U69 ( .A0(n21), .A1(n45), .Z(remaining_credit_v[2]));
Q_AN02 U70 ( .A0(n21), .A1(n46), .Z(remaining_credit_v[1]));
Q_AN02 U71 ( .A0(n21), .A1(n48), .Z(remaining_credit_v[0]));
Q_AD02 U72 ( .CI(n38), .A0(sw_config[7]), .A1(sw_config[8]), .B0(n80), .B1(n81), .S0(n37), .S1(n36), .CO(n35));
Q_AD02 U73 ( .CI(n41), .A0(sw_config[5]), .A1(sw_config[6]), .B0(n70), .B1(n78), .S0(n40), .S1(n39), .CO(n38));
Q_AD02 U74 ( .CI(n44), .A0(sw_config[3]), .A1(sw_config[4]), .B0(n65), .B1(n67), .S0(n43), .S1(n42), .CO(n41));
Q_AD02 U75 ( .CI(n56), .A0(sw_config[1]), .A1(sw_config[2]), .B0(n47), .B1(n63), .S0(n46), .S1(n45), .CO(n44));
Q_OR02 U76 ( .A0(sw_config[0]), .A1(n53), .Z(n47));
Q_XNR2 U77 ( .A0(sw_config[0]), .A1(n53), .Z(n48));
Q_XNR3 U78 ( .A0(sw_config[9]), .A1(n166), .A2(n35), .Z(n34));
Q_OR03 U79 ( .A0(n72), .A1(n49), .A2(n50), .Z(n21));
Q_AN03 U80 ( .A0(n71), .A1(n57), .A2(n51), .Z(n50));
Q_AO21 U81 ( .A0(n54), .A1(n52), .B0(n55), .Z(n51));
Q_AN02 U82 ( .A0(sw_config[0]), .A1(n53), .Z(n52));
Q_INV U83 ( .A(n175), .Z(n53));
Q_OR02 U84 ( .A0(sw_config[1]), .A1(n56), .Z(n54));
Q_AN02 U85 ( .A0(sw_config[1]), .A1(n56), .Z(n55));
Q_INV U86 ( .A(n174), .Z(n56));
Q_OA21 U87 ( .A0(n58), .A1(n59), .B0(n71), .Z(n49));
Q_AO21 U88 ( .A0(n68), .A1(n66), .B0(n69), .Z(n58));
Q_AO21 U89 ( .A0(n62), .A1(n64), .B0(n60), .Z(n59));
Q_OA21 U90 ( .A0(sw_config[2]), .A1(n63), .B0(n61), .Z(n57));
Q_AN03 U91 ( .A0(sw_config[2]), .A1(n63), .A2(n61), .Z(n60));
Q_INV U92 ( .A(n173), .Z(n63));
Q_OA21 U93 ( .A0(sw_config[3]), .A1(n65), .B0(n62), .Z(n61));
Q_AN02 U94 ( .A0(sw_config[3]), .A1(n65), .Z(n64));
Q_INV U95 ( .A(n172), .Z(n65));
Q_OA21 U96 ( .A0(sw_config[4]), .A1(n67), .B0(n68), .Z(n62));
Q_AN02 U97 ( .A0(sw_config[4]), .A1(n67), .Z(n66));
Q_INV U98 ( .A(n171), .Z(n67));
Q_OR02 U99 ( .A0(sw_config[5]), .A1(n70), .Z(n68));
Q_AN02 U100 ( .A0(sw_config[5]), .A1(n70), .Z(n69));
Q_INV U101 ( .A(n170), .Z(n70));
Q_OR03 U102 ( .A0(n83), .A1(n73), .A2(n74), .Z(n72));
Q_AO21 U103 ( .A0(n77), .A1(n79), .B0(n75), .Z(n74));
Q_OA21 U104 ( .A0(sw_config[6]), .A1(n78), .B0(n76), .Z(n71));
Q_AN03 U105 ( .A0(sw_config[6]), .A1(n78), .A2(n76), .Z(n75));
Q_INV U106 ( .A(n169), .Z(n78));
Q_OA21 U107 ( .A0(sw_config[7]), .A1(n80), .B0(n77), .Z(n76));
Q_AN02 U108 ( .A0(sw_config[7]), .A1(n80), .Z(n79));
Q_INV U109 ( .A(n168), .Z(n80));
Q_OA21 U110 ( .A0(sw_config[8]), .A1(n81), .B0(n82), .Z(n77));
Q_AN03 U111 ( .A0(sw_config[8]), .A1(n81), .A2(n82), .Z(n73));
Q_INV U112 ( .A(n167), .Z(n81));
Q_OR02 U113 ( .A0(sw_config[9]), .A1(n84), .Z(n82));
Q_AN02 U114 ( .A0(sw_config[9]), .A1(n84), .Z(n83));
Q_INV U115 ( .A(n166), .Z(n84));
Q_OR03 U116 ( .A0(n117), .A1(n85), .A2(n86), .Z(n22));
Q_AN03 U117 ( .A0(n116), .A1(n98), .A2(n87), .Z(n86));
Q_OR03 U118 ( .A0(n96), .A1(n88), .A2(n89), .Z(n87));
Q_AN02 U119 ( .A0(n95), .A1(n93), .Z(n88));
Q_AN03 U120 ( .A0(n95), .A1(n92), .A2(n90), .Z(n89));
Q_AN02 U121 ( .A0(sw_config[0]), .A1(n91), .Z(n90));
Q_INV U122 ( .A(n147), .Z(n91));
Q_OR02 U123 ( .A0(sw_config[1]), .A1(n94), .Z(n92));
Q_AN02 U124 ( .A0(sw_config[1]), .A1(n94), .Z(n93));
Q_INV U125 ( .A(n145), .Z(n94));
Q_OR02 U126 ( .A0(sw_config[2]), .A1(n97), .Z(n95));
Q_AN02 U127 ( .A0(sw_config[2]), .A1(n97), .Z(n96));
Q_INV U128 ( .A(n144), .Z(n97));
Q_AN02 U129 ( .A0(n102), .A1(n104), .Z(n98));
Q_OA21 U130 ( .A0(n99), .A1(n100), .B0(n116), .Z(n85));
Q_AO21 U131 ( .A0(n113), .A1(n111), .B0(n114), .Z(n99));
Q_AO21 U132 ( .A0(n103), .A1(n108), .B0(n101), .Z(n100));
Q_AN02 U133 ( .A0(n102), .A1(n105), .Z(n101));
Q_AN02 U134 ( .A0(n103), .A1(n107), .Z(n102));
Q_AN02 U135 ( .A0(n113), .A1(n110), .Z(n103));
Q_OR02 U136 ( .A0(sw_config[3]), .A1(n106), .Z(n104));
Q_AN02 U137 ( .A0(sw_config[3]), .A1(n106), .Z(n105));
Q_INV U138 ( .A(n142), .Z(n106));
Q_OR02 U139 ( .A0(sw_config[4]), .A1(n109), .Z(n107));
Q_AN02 U140 ( .A0(sw_config[4]), .A1(n109), .Z(n108));
Q_INV U141 ( .A(n141), .Z(n109));
Q_OR02 U142 ( .A0(sw_config[5]), .A1(n112), .Z(n110));
Q_AN02 U143 ( .A0(sw_config[5]), .A1(n112), .Z(n111));
Q_INV U144 ( .A(n139), .Z(n112));
Q_OR02 U145 ( .A0(sw_config[6]), .A1(n115), .Z(n113));
Q_AN02 U146 ( .A0(sw_config[6]), .A1(n115), .Z(n114));
Q_INV U147 ( .A(n138), .Z(n115));
Q_AN02 U148 ( .A0(n120), .A1(n122), .Z(n116));
Q_AO21 U149 ( .A0(n131), .A1(n129), .B0(n118), .Z(n117));
Q_AO21 U150 ( .A0(n121), .A1(n126), .B0(n119), .Z(n118));
Q_AN02 U151 ( .A0(n120), .A1(n123), .Z(n119));
Q_AN02 U152 ( .A0(n121), .A1(n125), .Z(n120));
Q_AN02 U153 ( .A0(n131), .A1(n128), .Z(n121));
Q_OR02 U154 ( .A0(sw_config[7]), .A1(n124), .Z(n122));
Q_AN02 U155 ( .A0(sw_config[7]), .A1(n124), .Z(n123));
Q_INV U156 ( .A(n136), .Z(n124));
Q_OR02 U157 ( .A0(sw_config[8]), .A1(n127), .Z(n125));
Q_AN02 U158 ( .A0(sw_config[8]), .A1(n127), .Z(n126));
Q_INV U159 ( .A(n135), .Z(n127));
Q_OR02 U160 ( .A0(sw_config[9]), .A1(n130), .Z(n128));
Q_AN02 U161 ( .A0(sw_config[9]), .A1(n130), .Z(n129));
Q_INV U162 ( .A(n133), .Z(n130));
Q_INV U163 ( .A(n132), .Z(n131));
Q_MX02 U164 ( .S(n22), .A0(sw_config[9]), .A1(n133), .Z(credit_issued_v[9]));
Q_MX02 U165 ( .S(n22), .A0(sw_config[8]), .A1(n135), .Z(credit_issued_v[8]));
Q_MX02 U166 ( .S(n22), .A0(sw_config[7]), .A1(n136), .Z(credit_issued_v[7]));
Q_MX02 U167 ( .S(n22), .A0(sw_config[6]), .A1(n138), .Z(credit_issued_v[6]));
Q_MX02 U168 ( .S(n22), .A0(sw_config[5]), .A1(n139), .Z(credit_issued_v[5]));
Q_MX02 U169 ( .S(n22), .A0(sw_config[4]), .A1(n141), .Z(credit_issued_v[4]));
Q_MX02 U170 ( .S(n22), .A0(sw_config[3]), .A1(n142), .Z(credit_issued_v[3]));
Q_MX02 U171 ( .S(n22), .A0(sw_config[2]), .A1(n144), .Z(credit_issued_v[2]));
Q_MX02 U172 ( .S(n22), .A0(sw_config[1]), .A1(n145), .Z(credit_issued_v[1]));
Q_MX02 U173 ( .S(n22), .A0(sw_config[0]), .A1(n147), .Z(credit_issued_v[0]));
Q_AD01HF U174 ( .A0(n166), .B0(n134), .S(n133), .CO(n132));
Q_AD02 U175 ( .CI(n137), .A0(credit_used[7]), .A1(credit_used[8]), .B0(n168), .B1(n167), .S0(n136), .S1(n135), .CO(n134));
Q_AD02 U176 ( .CI(n140), .A0(credit_used[5]), .A1(credit_used[6]), .B0(n170), .B1(n169), .S0(n139), .S1(n138), .CO(n137));
Q_AD02 U177 ( .CI(n143), .A0(credit_used[3]), .A1(credit_used[4]), .B0(n172), .B1(n171), .S0(n142), .S1(n141), .CO(n140));
Q_AD02 U178 ( .CI(n174), .A0(credit_used[1]), .A1(credit_used[2]), .B0(n146), .B1(n173), .S0(n145), .S1(n144), .CO(n143));
Q_AD01HF U179 ( .A0(credit_used[0]), .B0(n175), .S(n147), .CO(n146));
Q_OR03 U180 ( .A0(n148), .A1(n149), .A2(n164), .Z(used_err_v));
Q_AN03 U181 ( .A0(n163), .A1(n156), .A2(n150), .Z(n149));
Q_OR03 U182 ( .A0(n519), .A1(n151), .A2(n152), .Z(n150));
Q_NR02 U183 ( .A0(n105), .A1(n95), .Z(n151));
Q_AO21 U184 ( .A0(n154), .A1(n516), .B0(n153), .Z(n152));
Q_AN03 U185 ( .A0(n154), .A1(n515), .A2(n155), .Z(n153));
Q_NR02 U186 ( .A0(n105), .A1(n96), .Z(n154));
Q_AN02 U187 ( .A0(n147), .A1(n483), .Z(n155));
Q_AN02 U188 ( .A0(n161), .A1(n517), .Z(n156));
Q_OA21 U189 ( .A0(n157), .A1(n159), .B0(n163), .Z(n148));
Q_OR02 U190 ( .A0(n522), .A1(n158), .Z(n157));
Q_NR02 U191 ( .A0(n123), .A1(n113), .Z(n158));
Q_AO21 U192 ( .A0(n162), .A1(n521), .B0(n160), .Z(n159));
Q_AN02 U193 ( .A0(n161), .A1(n518), .Z(n160));
Q_AN02 U194 ( .A0(n162), .A1(n520), .Z(n161));
Q_NR02 U195 ( .A0(n123), .A1(n114), .Z(n162));
Q_NR02 U196 ( .A0(n129), .A1(n126), .Z(n163));
Q_OR03 U197 ( .A0(n523), .A1(n165), .A2(n132), .Z(n164));
Q_NR02 U198 ( .A0(n129), .A1(n125), .Z(n165));
Q_AN02 U199 ( .A0(n23), .A1(n176), .Z(n166));
Q_AN02 U200 ( .A0(n23), .A1(n178), .Z(n167));
Q_AN02 U201 ( .A0(n23), .A1(n179), .Z(n168));
Q_AN02 U202 ( .A0(n23), .A1(n181), .Z(n169));
Q_AN02 U203 ( .A0(n23), .A1(n182), .Z(n170));
Q_AN02 U204 ( .A0(n23), .A1(n184), .Z(n171));
Q_AN02 U205 ( .A0(n23), .A1(n185), .Z(n172));
Q_AN02 U206 ( .A0(n23), .A1(n187), .Z(n173));
Q_AN02 U207 ( .A0(n23), .A1(n188), .Z(n174));
Q_AN02 U208 ( .A0(n23), .A1(n190), .Z(n175));
Q_XOR2 U209 ( .A0(n233), .A1(n177), .Z(n176));
Q_AD02 U210 ( .CI(n180), .A0(credit_issued_r[7]), .A1(credit_issued_r[8]), .B0(n192), .B1(n191), .S0(n179), .S1(n178), .CO(n177));
Q_AD02 U211 ( .CI(n183), .A0(credit_issued_r[5]), .A1(credit_issued_r[6]), .B0(n194), .B1(n193), .S0(n182), .S1(n181), .CO(n180));
Q_AD02 U212 ( .CI(n186), .A0(credit_issued_r[3]), .A1(credit_issued_r[4]), .B0(n196), .B1(n195), .S0(n185), .S1(n184), .CO(n183));
Q_AD02 U213 ( .CI(n189), .A0(credit_issued_r[1]), .A1(credit_issued_r[2]), .B0(n198), .B1(n197), .S0(n188), .S1(n187), .CO(n186));
Q_OR02 U214 ( .A0(credit_issued_r[0]), .A1(n199), .Z(n189));
Q_XNR2 U215 ( .A0(credit_issued_r[0]), .A1(n199), .Z(n190));
Q_INV U216 ( .A(credit_return[8]), .Z(n191));
Q_INV U217 ( .A(credit_return[7]), .Z(n192));
Q_INV U218 ( .A(credit_return[6]), .Z(n193));
Q_INV U219 ( .A(credit_return[5]), .Z(n194));
Q_INV U220 ( .A(credit_return[4]), .Z(n195));
Q_INV U221 ( .A(credit_return[3]), .Z(n196));
Q_INV U222 ( .A(credit_return[2]), .Z(n197));
Q_INV U223 ( .A(credit_return[1]), .Z(n198));
Q_INV U224 ( .A(credit_return[0]), .Z(n199));
Q_INV U225 ( .A(return_err_v), .Z(n23));
Q_OR03 U226 ( .A0(n223), .A1(n200), .A2(n201), .Z(return_err_v));
Q_AN03 U227 ( .A0(n222), .A1(n208), .A2(n202), .Z(n201));
Q_AO21 U228 ( .A0(n205), .A1(n203), .B0(n206), .Z(n202));
Q_AN02 U229 ( .A0(credit_return[0]), .A1(n204), .Z(n203));
Q_OR02 U230 ( .A0(credit_return[1]), .A1(n207), .Z(n205));
Q_AN02 U231 ( .A0(credit_return[1]), .A1(n207), .Z(n206));
Q_OA21 U232 ( .A0(n209), .A1(n210), .B0(n222), .Z(n200));
Q_AO21 U233 ( .A0(n219), .A1(n217), .B0(n220), .Z(n209));
Q_AO21 U234 ( .A0(n213), .A1(n215), .B0(n211), .Z(n210));
Q_OA21 U235 ( .A0(credit_return[2]), .A1(n214), .B0(n212), .Z(n208));
Q_AN03 U236 ( .A0(credit_return[2]), .A1(n214), .A2(n212), .Z(n211));
Q_OA21 U237 ( .A0(credit_return[3]), .A1(n216), .B0(n213), .Z(n212));
Q_AN02 U238 ( .A0(credit_return[3]), .A1(n216), .Z(n215));
Q_OA21 U239 ( .A0(credit_return[4]), .A1(n218), .B0(n219), .Z(n213));
Q_AN02 U240 ( .A0(credit_return[4]), .A1(n218), .Z(n217));
Q_OR02 U241 ( .A0(credit_return[5]), .A1(n221), .Z(n219));
Q_AN02 U242 ( .A0(credit_return[5]), .A1(n221), .Z(n220));
Q_AO21 U243 ( .A0(n233), .A1(n231), .B0(n224), .Z(n223));
Q_AO21 U244 ( .A0(n227), .A1(n229), .B0(n225), .Z(n224));
Q_OA21 U245 ( .A0(credit_return[6]), .A1(n228), .B0(n226), .Z(n222));
Q_AN03 U246 ( .A0(credit_return[6]), .A1(n228), .A2(n226), .Z(n225));
Q_OA21 U247 ( .A0(credit_return[7]), .A1(n230), .B0(n227), .Z(n226));
Q_AN02 U248 ( .A0(credit_return[7]), .A1(n230), .Z(n229));
Q_OA21 U249 ( .A0(credit_return[8]), .A1(n232), .B0(n233), .Z(n227));
Q_AN02 U250 ( .A0(credit_return[8]), .A1(n232), .Z(n231));
Q_FDP1 \credit_limit_REG[0] ( .CK(clk), .R(rst_n), .D(n276), .Q(credit_limit[0]), .QN( ));
Q_FDP1 \credit_limit_REG[1] ( .CK(clk), .R(rst_n), .D(n275), .Q(credit_limit[1]), .QN( ));
Q_FDP1 \credit_limit_REG[2] ( .CK(clk), .R(rst_n), .D(n274), .Q(credit_limit[2]), .QN( ));
Q_FDP1 \credit_limit_REG[3] ( .CK(clk), .R(rst_n), .D(n273), .Q(credit_limit[3]), .QN( ));
Q_FDP1 \credit_limit_REG[4] ( .CK(clk), .R(rst_n), .D(n272), .Q(credit_limit[4]), .QN( ));
Q_FDP1 \credit_limit_REG[5] ( .CK(clk), .R(rst_n), .D(n271), .Q(credit_limit[5]), .QN( ));
Q_FDP1 \credit_limit_REG[6] ( .CK(clk), .R(rst_n), .D(n270), .Q(credit_limit[6]), .QN( ));
Q_FDP1 \credit_limit_REG[7] ( .CK(clk), .R(rst_n), .D(n269), .Q(credit_limit[7]), .QN( ));
Q_FDP1 \credit_limit_REG[8] ( .CK(clk), .R(rst_n), .D(n268), .Q(credit_limit[8]), .QN( ));
Q_FDP2 \credit_limit_REG[9] ( .CK(clk), .S(rst_n), .D(n267), .Q(credit_limit[9]), .QN( ));
Q_FDP1 \outstanding_REG[0] ( .CK(clk), .R(rst_n), .D(n266), .Q(outstanding[0]), .QN(n428));
Q_FDP1 \outstanding_REG[1] ( .CK(clk), .R(rst_n), .D(n265), .Q(outstanding[1]), .QN(n431));
Q_FDP1 \outstanding_REG[2] ( .CK(clk), .R(rst_n), .D(n264), .Q(outstanding[2]), .QN(n432));
Q_FDP1 \outstanding_REG[3] ( .CK(clk), .R(rst_n), .D(n263), .Q(outstanding[3]), .QN(n435));
Q_FDP1 \outstanding_REG[4] ( .CK(clk), .R(rst_n), .D(n262), .Q(outstanding[4]), .QN(n443));
Q_FDP1 \outstanding_REG[5] ( .CK(clk), .R(rst_n), .D(n261), .Q(outstanding[5]), .QN(n445));
Q_FDP1 \outstanding_REG[6] ( .CK(clk), .R(rst_n), .D(n260), .Q(outstanding[6]), .QN(n446));
Q_FDP1 \outstanding_REG[7] ( .CK(clk), .R(rst_n), .D(n259), .Q(outstanding[7]), .QN(n449));
Q_FDP1 \outstanding_REG[8] ( .CK(clk), .R(rst_n), .D(n258), .Q(outstanding[8]), .QN(n454));
Q_FDP1 \outstanding_REG[9] ( .CK(clk), .R(rst_n), .D(n257), .Q(outstanding[9]), .QN(n455));
Q_FDP1 \outstanding_REG[10] ( .CK(clk), .R(rst_n), .D(n256), .Q(outstanding[10]), .QN( ));
Q_FDP1 \outstanding_REG[11] ( .CK(clk), .R(rst_n), .D(n255), .Q(outstanding[11]), .QN( ));
Q_FDP1 \outstanding_REG[12] ( .CK(clk), .R(rst_n), .D(n254), .Q(outstanding[12]), .QN(n458));
Q_FDP1 \outstanding_REG[13] ( .CK(clk), .R(rst_n), .D(n253), .Q(outstanding[13]), .QN(n459));
Q_FDP1 \outstanding_REG[14] ( .CK(clk), .R(rst_n), .D(n252), .Q(outstanding[14]), .QN( ));
Q_FDP1 \outstanding_REG[15] ( .CK(clk), .R(rst_n), .D(n251), .Q(outstanding[15]), .QN( ));
Q_FDP1 \outstanding_REG[16] ( .CK(clk), .R(rst_n), .D(n250), .Q(outstanding[16]), .QN(n462));
Q_FDP1 \outstanding_REG[17] ( .CK(clk), .R(rst_n), .D(n249), .Q(outstanding[17]), .QN(n463));
Q_FDP1 \outstanding_REG[18] ( .CK(clk), .R(rst_n), .D(n248), .Q(outstanding[18]), .QN( ));
Q_FDP1 \outstanding_REG[19] ( .CK(clk), .R(rst_n), .D(n247), .Q(outstanding[19]), .QN( ));
Q_FDP1 \outstanding_REG[20] ( .CK(clk), .R(rst_n), .D(n246), .Q(outstanding[20]), .QN(n466));
Q_FDP1 \outstanding_REG[21] ( .CK(clk), .R(rst_n), .D(n245), .Q(outstanding[21]), .QN(n467));
Q_FDP1 \outstanding_REG[22] ( .CK(clk), .R(rst_n), .D(n244), .Q(outstanding[22]), .QN( ));
Q_FDP1 \outstanding_REG[23] ( .CK(clk), .R(rst_n), .D(n243), .Q(outstanding[23]), .QN( ));
Q_FDP1 \outstanding_REG[24] ( .CK(clk), .R(rst_n), .D(n242), .Q(outstanding[24]), .QN(n470));
Q_FDP1 \outstanding_REG[25] ( .CK(clk), .R(rst_n), .D(n241), .Q(outstanding[25]), .QN(n471));
Q_FDP1 \outstanding_REG[26] ( .CK(clk), .R(rst_n), .D(n240), .Q(outstanding[26]), .QN( ));
Q_FDP1 \outstanding_REG[27] ( .CK(clk), .R(rst_n), .D(n239), .Q(outstanding[27]), .QN( ));
Q_FDP1 \outstanding_REG[28] ( .CK(clk), .R(rst_n), .D(n238), .Q(outstanding[28]), .QN(n474));
Q_FDP1 \outstanding_REG[29] ( .CK(clk), .R(rst_n), .D(n237), .Q(outstanding[29]), .QN(n475));
Q_FDP1 \outstanding_REG[30] ( .CK(clk), .R(rst_n), .D(n236), .Q(outstanding[30]), .QN( ));
Q_FDP1 \outstanding_REG[31] ( .CK(clk), .R(rst_n), .D(n235), .Q(outstanding[31]), .QN( ));
Q_AN02 U293 ( .A0(n1), .A1(n277), .Z(n235));
Q_AN02 U294 ( .A0(n1), .A1(n279), .Z(n236));
Q_AN02 U295 ( .A0(n1), .A1(n281), .Z(n237));
Q_AN02 U296 ( .A0(n1), .A1(n283), .Z(n238));
Q_AN02 U297 ( .A0(n1), .A1(n285), .Z(n239));
Q_AN02 U298 ( .A0(n1), .A1(n287), .Z(n240));
Q_AN02 U299 ( .A0(n1), .A1(n289), .Z(n241));
Q_AN02 U300 ( .A0(n1), .A1(n291), .Z(n242));
Q_AN02 U301 ( .A0(n1), .A1(n293), .Z(n243));
Q_AN02 U302 ( .A0(n1), .A1(n295), .Z(n244));
Q_AN02 U303 ( .A0(n1), .A1(n297), .Z(n245));
Q_AN02 U304 ( .A0(n1), .A1(n299), .Z(n246));
Q_AN02 U305 ( .A0(n1), .A1(n301), .Z(n247));
Q_AN02 U306 ( .A0(n1), .A1(n303), .Z(n248));
Q_AN02 U307 ( .A0(n1), .A1(n305), .Z(n249));
Q_AN02 U308 ( .A0(n1), .A1(n307), .Z(n250));
Q_AN02 U309 ( .A0(n1), .A1(n309), .Z(n251));
Q_AN02 U310 ( .A0(n1), .A1(n311), .Z(n252));
Q_AN02 U311 ( .A0(n1), .A1(n313), .Z(n253));
Q_AN02 U312 ( .A0(n1), .A1(n315), .Z(n254));
Q_AN02 U313 ( .A0(n1), .A1(n317), .Z(n255));
Q_AN02 U314 ( .A0(n1), .A1(n319), .Z(n256));
Q_AN02 U315 ( .A0(n1), .A1(n321), .Z(n257));
Q_AN02 U316 ( .A0(n1), .A1(n323), .Z(n258));
Q_AN02 U317 ( .A0(n1), .A1(n325), .Z(n259));
Q_AN02 U318 ( .A0(n1), .A1(n327), .Z(n260));
Q_AN02 U319 ( .A0(n1), .A1(n329), .Z(n261));
Q_AN02 U320 ( .A0(n1), .A1(n331), .Z(n262));
Q_AN02 U321 ( .A0(n1), .A1(n333), .Z(n263));
Q_AN02 U322 ( .A0(n1), .A1(n335), .Z(n264));
Q_AN02 U323 ( .A0(n1), .A1(n337), .Z(n265));
Q_AN02 U324 ( .A0(n1), .A1(n339), .Z(n266));
Q_OR02 U325 ( .A0(sw_init), .A1(sw_config[9]), .Z(n267));
Q_AN02 U326 ( .A0(n1), .A1(sw_config[8]), .Z(n268));
Q_AN02 U327 ( .A0(n1), .A1(sw_config[7]), .Z(n269));
Q_AN02 U328 ( .A0(n1), .A1(sw_config[6]), .Z(n270));
Q_AN02 U329 ( .A0(n1), .A1(sw_config[5]), .Z(n271));
Q_AN02 U330 ( .A0(n1), .A1(sw_config[4]), .Z(n272));
Q_AN02 U331 ( .A0(n1), .A1(sw_config[3]), .Z(n273));
Q_AN02 U332 ( .A0(n1), .A1(sw_config[2]), .Z(n274));
Q_AN02 U333 ( .A0(n1), .A1(sw_config[1]), .Z(n275));
Q_AN02 U334 ( .A0(n1), .A1(sw_config[0]), .Z(n276));
Q_XNR3 U335 ( .A0(n278), .A1(outstanding[31]), .A2(n340), .Z(n277));
Q_AD01HF U336 ( .A0(n280), .B0(n341), .S(n279), .CO(n278));
Q_AD01HF U337 ( .A0(n282), .B0(n343), .S(n281), .CO(n280));
Q_AD01HF U338 ( .A0(n284), .B0(n345), .S(n283), .CO(n282));
Q_AD01HF U339 ( .A0(n286), .B0(n347), .S(n285), .CO(n284));
Q_AD01HF U340 ( .A0(n288), .B0(n349), .S(n287), .CO(n286));
Q_AD01HF U341 ( .A0(n290), .B0(n351), .S(n289), .CO(n288));
Q_AD01HF U342 ( .A0(n292), .B0(n353), .S(n291), .CO(n290));
Q_AD01HF U343 ( .A0(n294), .B0(n355), .S(n293), .CO(n292));
Q_AD01HF U344 ( .A0(n296), .B0(n357), .S(n295), .CO(n294));
Q_AD01HF U345 ( .A0(n298), .B0(n359), .S(n297), .CO(n296));
Q_AD01HF U346 ( .A0(n300), .B0(n361), .S(n299), .CO(n298));
Q_AD01HF U347 ( .A0(n302), .B0(n363), .S(n301), .CO(n300));
Q_AD01HF U348 ( .A0(n304), .B0(n365), .S(n303), .CO(n302));
Q_AD01HF U349 ( .A0(n306), .B0(n367), .S(n305), .CO(n304));
Q_AD01HF U350 ( .A0(n308), .B0(n369), .S(n307), .CO(n306));
Q_AD01HF U351 ( .A0(n310), .B0(n371), .S(n309), .CO(n308));
Q_AD01HF U352 ( .A0(n312), .B0(n373), .S(n311), .CO(n310));
Q_AD01HF U353 ( .A0(n314), .B0(n375), .S(n313), .CO(n312));
Q_AD01HF U354 ( .A0(n316), .B0(n377), .S(n315), .CO(n314));
Q_AD01HF U355 ( .A0(n318), .B0(n379), .S(n317), .CO(n316));
Q_AD01HF U356 ( .A0(n320), .B0(n381), .S(n319), .CO(n318));
Q_AD01HF U357 ( .A0(n383), .B0(n322), .S(n321), .CO(n320));
Q_AD01 U358 ( .CI(n324), .A0(n385), .B0(n386), .S(n323), .CO(n322));
Q_AD01 U359 ( .CI(n326), .A0(n387), .B0(n388), .S(n325), .CO(n324));
Q_AD01 U360 ( .CI(n328), .A0(n389), .B0(n390), .S(n327), .CO(n326));
Q_AD01 U361 ( .CI(n330), .A0(n391), .B0(n392), .S(n329), .CO(n328));
Q_AD01 U362 ( .CI(n332), .A0(n393), .B0(n394), .S(n331), .CO(n330));
Q_AD01 U363 ( .CI(n334), .A0(n395), .B0(n396), .S(n333), .CO(n332));
Q_AD01 U364 ( .CI(n336), .A0(n397), .B0(n398), .S(n335), .CO(n334));
Q_AD01 U365 ( .CI(n399), .A0(n338), .B0(n400), .S(n337), .CO(n336));
Q_AD01HF U366 ( .A0(n199), .B0(n401), .S(n339), .CO(n338));
Q_OR02 U367 ( .A0(outstanding[30]), .A1(n342), .Z(n340));
Q_XNR2 U368 ( .A0(outstanding[30]), .A1(n342), .Z(n341));
Q_OR02 U369 ( .A0(outstanding[29]), .A1(n344), .Z(n342));
Q_XNR2 U370 ( .A0(outstanding[29]), .A1(n344), .Z(n343));
Q_OR02 U371 ( .A0(outstanding[28]), .A1(n346), .Z(n344));
Q_XNR2 U372 ( .A0(outstanding[28]), .A1(n346), .Z(n345));
Q_OR02 U373 ( .A0(outstanding[27]), .A1(n348), .Z(n346));
Q_XNR2 U374 ( .A0(outstanding[27]), .A1(n348), .Z(n347));
Q_OR02 U375 ( .A0(outstanding[26]), .A1(n350), .Z(n348));
Q_XNR2 U376 ( .A0(outstanding[26]), .A1(n350), .Z(n349));
Q_OR02 U377 ( .A0(outstanding[25]), .A1(n352), .Z(n350));
Q_XNR2 U378 ( .A0(outstanding[25]), .A1(n352), .Z(n351));
Q_OR02 U379 ( .A0(outstanding[24]), .A1(n354), .Z(n352));
Q_XNR2 U380 ( .A0(outstanding[24]), .A1(n354), .Z(n353));
Q_OR02 U381 ( .A0(outstanding[23]), .A1(n356), .Z(n354));
Q_XNR2 U382 ( .A0(outstanding[23]), .A1(n356), .Z(n355));
Q_OR02 U383 ( .A0(outstanding[22]), .A1(n358), .Z(n356));
Q_XNR2 U384 ( .A0(outstanding[22]), .A1(n358), .Z(n357));
Q_OR02 U385 ( .A0(outstanding[21]), .A1(n360), .Z(n358));
Q_XNR2 U386 ( .A0(outstanding[21]), .A1(n360), .Z(n359));
Q_OR02 U387 ( .A0(outstanding[20]), .A1(n362), .Z(n360));
Q_XNR2 U388 ( .A0(outstanding[20]), .A1(n362), .Z(n361));
Q_OR02 U389 ( .A0(outstanding[19]), .A1(n364), .Z(n362));
Q_XNR2 U390 ( .A0(outstanding[19]), .A1(n364), .Z(n363));
Q_OR02 U391 ( .A0(outstanding[18]), .A1(n366), .Z(n364));
Q_XNR2 U392 ( .A0(outstanding[18]), .A1(n366), .Z(n365));
Q_OR02 U393 ( .A0(outstanding[17]), .A1(n368), .Z(n366));
Q_XNR2 U394 ( .A0(outstanding[17]), .A1(n368), .Z(n367));
Q_OR02 U395 ( .A0(outstanding[16]), .A1(n370), .Z(n368));
Q_XNR2 U396 ( .A0(outstanding[16]), .A1(n370), .Z(n369));
Q_OR02 U397 ( .A0(outstanding[15]), .A1(n372), .Z(n370));
Q_XNR2 U398 ( .A0(outstanding[15]), .A1(n372), .Z(n371));
Q_OR02 U399 ( .A0(outstanding[14]), .A1(n374), .Z(n372));
Q_XNR2 U400 ( .A0(outstanding[14]), .A1(n374), .Z(n373));
Q_OR02 U401 ( .A0(outstanding[13]), .A1(n376), .Z(n374));
Q_XNR2 U402 ( .A0(outstanding[13]), .A1(n376), .Z(n375));
Q_OR02 U403 ( .A0(outstanding[12]), .A1(n378), .Z(n376));
Q_XNR2 U404 ( .A0(outstanding[12]), .A1(n378), .Z(n377));
Q_OR02 U405 ( .A0(outstanding[11]), .A1(n380), .Z(n378));
Q_XNR2 U406 ( .A0(outstanding[11]), .A1(n380), .Z(n379));
Q_OR02 U407 ( .A0(outstanding[10]), .A1(n382), .Z(n380));
Q_XNR2 U408 ( .A0(outstanding[10]), .A1(n382), .Z(n381));
Q_OR02 U409 ( .A0(outstanding[9]), .A1(n384), .Z(n382));
Q_XNR2 U410 ( .A0(outstanding[9]), .A1(n384), .Z(n383));
Q_AD01 U411 ( .CI(n191), .A0(outstanding[8]), .B0(credit_used[8]), .S(n385), .CO(n384));
Q_AD01 U412 ( .CI(n192), .A0(outstanding[7]), .B0(credit_used[7]), .S(n387), .CO(n386));
Q_AD01 U413 ( .CI(n193), .A0(outstanding[6]), .B0(credit_used[6]), .S(n389), .CO(n388));
Q_AD01 U414 ( .CI(n194), .A0(outstanding[5]), .B0(credit_used[5]), .S(n391), .CO(n390));
Q_AD01 U415 ( .CI(n195), .A0(outstanding[4]), .B0(credit_used[4]), .S(n393), .CO(n392));
Q_AD01 U416 ( .CI(n196), .A0(outstanding[3]), .B0(credit_used[3]), .S(n395), .CO(n394));
Q_AD01 U417 ( .CI(n197), .A0(outstanding[2]), .B0(credit_used[2]), .S(n397), .CO(n396));
Q_AD01 U418 ( .CI(n198), .A0(outstanding[1]), .B0(credit_used[1]), .S(n399), .CO(n398));
Q_OR02 U419 ( .A0(outstanding[0]), .A1(credit_used[0]), .Z(n400));
Q_XNR2 U420 ( .A0(outstanding[0]), .A1(credit_used[0]), .Z(n401));
Q_INV U421 ( .A(_zy_sva_b2), .Z(n402));
Q_AN02 U422 ( .A0(_zy_sva_b0), .A1(n403), .Z(n404));
Q_ND02 U423 ( .A0(_zy_sva_b0), .A1(_zy_sva_b1), .Z(n403));
Q_INV U424 ( .A(sw_config[9]), .Z(n514));
Q_AN02 U425 ( .A0(credit_limit[9]), .A1(n514), .Z(n513));
Q_OR02 U426 ( .A0(credit_limit[9]), .A1(n514), .Z(n512));
Q_INV U427 ( .A(sw_config[8]), .Z(n511));
Q_AN03 U428 ( .A0(credit_limit[8]), .A1(n511), .A2(n512), .Z(n503));
Q_OA21 U429 ( .A0(credit_limit[8]), .A1(n511), .B0(n512), .Z(n507));
Q_INV U430 ( .A(sw_config[7]), .Z(n510));
Q_AN02 U431 ( .A0(credit_limit[7]), .A1(n510), .Z(n509));
Q_OA21 U432 ( .A0(credit_limit[7]), .A1(n510), .B0(n507), .Z(n506));
Q_INV U433 ( .A(sw_config[6]), .Z(n508));
Q_AN03 U434 ( .A0(credit_limit[6]), .A1(n508), .A2(n506), .Z(n505));
Q_OA21 U435 ( .A0(credit_limit[6]), .A1(n508), .B0(n506), .Z(n501));
Q_AO21 U436 ( .A0(n507), .A1(n509), .B0(n505), .Z(n504));
Q_OR03 U437 ( .A0(n513), .A1(n503), .A2(n504), .Z(n502));
Q_INV U438 ( .A(sw_config[5]), .Z(n500));
Q_AN02 U439 ( .A0(credit_limit[5]), .A1(n500), .Z(n499));
Q_OR02 U440 ( .A0(credit_limit[5]), .A1(n500), .Z(n498));
Q_INV U441 ( .A(sw_config[4]), .Z(n497));
Q_AN02 U442 ( .A0(credit_limit[4]), .A1(n497), .Z(n496));
Q_OA21 U443 ( .A0(credit_limit[4]), .A1(n497), .B0(n498), .Z(n492));
Q_INV U444 ( .A(sw_config[3]), .Z(n495));
Q_AN02 U445 ( .A0(credit_limit[3]), .A1(n495), .Z(n494));
Q_OA21 U446 ( .A0(credit_limit[3]), .A1(n495), .B0(n492), .Z(n491));
Q_INV U447 ( .A(sw_config[2]), .Z(n493));
Q_AN03 U448 ( .A0(credit_limit[2]), .A1(n493), .A2(n491), .Z(n490));
Q_OA21 U449 ( .A0(credit_limit[2]), .A1(n493), .B0(n491), .Z(n487));
Q_AO21 U450 ( .A0(n492), .A1(n494), .B0(n490), .Z(n489));
Q_AO21 U451 ( .A0(n498), .A1(n496), .B0(n499), .Z(n488));
Q_OA21 U452 ( .A0(n488), .A1(n489), .B0(n501), .Z(n479));
Q_INV U453 ( .A(sw_config[1]), .Z(n486));
Q_AN02 U454 ( .A0(credit_limit[1]), .A1(n486), .Z(n485));
Q_OR02 U455 ( .A0(credit_limit[1]), .A1(n486), .Z(n484));
Q_INV U456 ( .A(sw_config[0]), .Z(n483));
Q_AN02 U457 ( .A0(credit_limit[0]), .A1(n483), .Z(n482));
Q_AO21 U458 ( .A0(n484), .A1(n482), .B0(n485), .Z(n481));
Q_AN03 U459 ( .A0(n501), .A1(n487), .A2(n481), .Z(n480));
Q_OR03 U460 ( .A0(n502), .A1(n479), .A2(n480), .Z(credit_decrease));
ixc_assign_9 _zz_strnp_0 ( _zy_simnet_credit_available_0_w$[0:8], 
	credit_available[8:0]);
ixc_assign_12 _zz_strnp_1 ( _zy_simnet_hw_status_1_w$[0:11], hw_status[11:0]);
Q_OR03 U463 ( .A0(credit_return[8]), .A1(credit_return[7]), .A2(credit_return[6]), .Z(n478));
Q_OR03 U464 ( .A0(credit_return[5]), .A1(credit_return[4]), .A2(credit_return[3]), .Z(n477));
Q_OR03 U465 ( .A0(credit_return[2]), .A1(credit_return[1]), .A2(credit_return[0]), .Z(n476));
Q_OR03 U466 ( .A0(n478), .A1(n477), .A2(n476), .Z(_zy_sva_b0_t));
Q_NR02 U467 ( .A0(outstanding[31]), .A1(outstanding[30]), .Z(n473));
Q_AN03 U468 ( .A0(n473), .A1(n475), .A2(n474), .Z(n472));
Q_NR02 U469 ( .A0(outstanding[27]), .A1(outstanding[26]), .Z(n469));
Q_AN03 U470 ( .A0(n469), .A1(n471), .A2(n470), .Z(n468));
Q_NR02 U471 ( .A0(outstanding[23]), .A1(outstanding[22]), .Z(n465));
Q_AN03 U472 ( .A0(n465), .A1(n467), .A2(n466), .Z(n464));
Q_NR02 U473 ( .A0(outstanding[19]), .A1(outstanding[18]), .Z(n461));
Q_AN03 U474 ( .A0(n461), .A1(n463), .A2(n462), .Z(n460));
Q_NR02 U475 ( .A0(outstanding[15]), .A1(outstanding[14]), .Z(n457));
Q_AN03 U476 ( .A0(n457), .A1(n459), .A2(n458), .Z(n456));
Q_AN03 U477 ( .A0(credit_return[8]), .A1(n454), .A2(n451), .Z(n450));
Q_OR02 U478 ( .A0(credit_return[8]), .A1(n454), .Z(n453));
Q_NR02 U479 ( .A0(outstanding[11]), .A1(outstanding[10]), .Z(n452));
Q_AN02 U480 ( .A0(n452), .A1(n455), .Z(n451));
Q_AN03 U481 ( .A0(n451), .A1(n453), .A2(n456), .Z(n420));
Q_AN02 U482 ( .A0(credit_return[7]), .A1(n449), .Z(n448));
Q_OR02 U483 ( .A0(credit_return[7]), .A1(n449), .Z(n447));
Q_AN03 U484 ( .A0(credit_return[6]), .A1(n446), .A2(n447), .Z(n438));
Q_OA21 U485 ( .A0(credit_return[6]), .A1(n446), .B0(n447), .Z(n442));
Q_AN02 U486 ( .A0(credit_return[5]), .A1(n445), .Z(n444));
Q_OA21 U487 ( .A0(credit_return[5]), .A1(n445), .B0(n442), .Z(n441));
Q_AN03 U488 ( .A0(credit_return[4]), .A1(n443), .A2(n441), .Z(n440));
Q_OA21 U489 ( .A0(credit_return[4]), .A1(n443), .B0(n441), .Z(n436));
Q_AO21 U490 ( .A0(n442), .A1(n444), .B0(n440), .Z(n439));
Q_OR03 U491 ( .A0(n448), .A1(n438), .A2(n439), .Z(n437));
Q_AN02 U492 ( .A0(credit_return[3]), .A1(n435), .Z(n434));
Q_OR02 U493 ( .A0(credit_return[3]), .A1(n435), .Z(n433));
Q_AN03 U494 ( .A0(credit_return[2]), .A1(n432), .A2(n433), .Z(n423));
Q_OA21 U495 ( .A0(credit_return[2]), .A1(n432), .B0(n433), .Z(n426));
Q_AN02 U496 ( .A0(credit_return[1]), .A1(n431), .Z(n430));
Q_OR02 U497 ( .A0(credit_return[1]), .A1(n431), .Z(n429));
Q_AN02 U498 ( .A0(credit_return[0]), .A1(n428), .Z(n427));
Q_AN03 U499 ( .A0(n426), .A1(n429), .A2(n427), .Z(n425));
Q_AO21 U500 ( .A0(n426), .A1(n430), .B0(n425), .Z(n424));
Q_OR03 U501 ( .A0(n434), .A1(n423), .A2(n424), .Z(n422));
Q_AN03 U502 ( .A0(n472), .A1(n468), .A2(n464), .Z(n421));
Q_ND03 U503 ( .A0(n421), .A1(n460), .A2(n417), .Z(_zy_sva_b1_t));
Q_AN03 U504 ( .A0(n420), .A1(n436), .A2(n422), .Z(n419));
Q_AO21 U505 ( .A0(n420), .A1(n437), .B0(n419), .Z(n418));
Q_AO21 U506 ( .A0(n456), .A1(n450), .B0(n418), .Z(n417));
Q_OR02 U507 ( .A0(sw_config[7]), .A1(sw_config[6]), .Z(n416));
Q_OA21 U508 ( .A0(sw_config[8]), .A1(n416), .B0(sw_config[9]), .Z(n415));
Q_OR02 U509 ( .A0(sw_config[3]), .A1(sw_config[2]), .Z(n414));
Q_OR02 U510 ( .A0(sw_config[5]), .A1(sw_config[4]), .Z(n413));
Q_OA21 U511 ( .A0(n413), .A1(n414), .B0(sw_config[9]), .Z(n411));
Q_NR03 U512 ( .A0(n415), .A1(n411), .A2(n412), .Z(_zy_sva_b2_t));
ixc_sample_logic_1_3 _zz_zy_sva_b0 ( _zy_sva_b0, _zy_sva_b0_t);
ixc_sample_logic_1_3 _zz_zy_sva_b1 ( _zy_sva_b1, _zy_sva_b1_t);
ixc_sample_logic_1_3 _zz_zy_sva_b2 ( _zy_sva_b2, _zy_sva_b2_t);
ixc_pio_call_0_0_0_0_1 _zzixc_tfport_1_1 ( _zyixc_port_1_1_ack, 
	_zyixc_port_1_1_s2hW, _zyixc_port_1_1_isf, _zyixc_port_1_1_req, n410, 
	_zyixc_port_1_1_osf, n409, n408);
ixc_pio_call_0_0_0_0_1 _zzixc_tfport_1_0 ( _zyixc_port_1_0_ack, 
	_zyixc_port_1_0_s2hW, _zyixc_port_1_0_isf, _zyixc_port_1_0_req, n407, 
	_zyixc_port_1_0_osf, n406, n405);
wire [2:0] n528 = 3'b000;
Q_ASSERT credit_return_check ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT( ), .FAIL_COUNT( ), .CHECK_COUNT( ), .KILL_SIGNAL( ), .SEVERITY(n528[0]));
// pragma CVASTRPROP INSTANCE "credit_return_check" HDL_ASSERT "$"
// pragma CVASTRPROP INSTANCE "credit_return_check" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/common/nx_library/nx_credit_manager.v"
//pragma CVAINTPROP INSTANCE "credit_return_check" ASSERT_LINE 116
wire [2:0] n529 = 3'b000;
Q_ASSERT credit_danger_check ( .PASS( ), .FAIL( ), .ACTIVE( ), .FAIL_LEVEL( ), .PASS_LEVEL( ), .DISABLE( ), .PASS_COUNT( ), .FAIL_COUNT( ), .CHECK_COUNT( ), .KILL_SIGNAL( ), .SEVERITY(n529[0]));
// pragma CVASTRPROP INSTANCE "credit_danger_check" HDL_ASSERT "$"
// pragma CVASTRPROP INSTANCE "credit_danger_check" ASSERT_FILENAME "/home/ibarry/Project-Zipline-master/rtl/common/nx_library/nx_credit_manager.v"
//pragma CVAINTPROP INSTANCE "credit_danger_check" ASSERT_LINE 122
Q_INV U520 ( .A(n93), .Z(n515));
Q_INV U521 ( .A(n92), .Z(n516));
Q_INV U522 ( .A(n108), .Z(n517));
Q_INV U523 ( .A(n107), .Z(n518));
Q_INV U524 ( .A(n104), .Z(n519));
Q_INV U525 ( .A(n111), .Z(n520));
Q_INV U526 ( .A(n110), .Z(n521));
Q_INV U527 ( .A(n122), .Z(n522));
Q_INV U528 ( .A(n128), .Z(n523));
Q_INV U529 ( .A(_zy_sva_credit_return_check_1_0_fail[0]), .Z(n524));
Q_FDP4EP \_zy_sva_credit_return_check_1_0_fail_REG[0] ( .CK(clk), .CE(n404), .R(n234), .D(n524), .Q(_zy_sva_credit_return_check_1_0_fail[0]));
Q_INV U531 ( .A(_zyixc_port_1_0_req), .Z(n525));
Q_FDP4EP _zyixc_port_1_0_req_REG  ( .CK(clk), .CE(n404), .R(n234), .D(n525), .Q(_zyixc_port_1_0_req));
Q_INV U533 ( .A(_zy_sva_credit_danger_check_2_3_fail[0]), .Z(n526));
Q_FDP4EP \_zy_sva_credit_danger_check_2_3_fail_REG[0] ( .CK(clk), .CE(n402), .R(n234), .D(n526), .Q(_zy_sva_credit_danger_check_2_3_fail[0]));
Q_INV U535 ( .A(_zyixc_port_1_1_req), .Z(n527));
Q_FDP4EP _zyixc_port_1_1_req_REG  ( .CK(clk), .CE(n402), .R(n234), .D(n527), .Q(_zyixc_port_1_1_req));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\hw_status.credit_issued  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\sw_config.credit_limit  (1,0) 1 9 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "2"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "hw_status 3 \hw_status.used_err  \hw_status.return_err  \hw_status.credit_issued "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "sw_config 3 \sw_config.dis_used  \sw_config.dis_return  \sw_config.credit_limit "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "2"
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
endmodule
