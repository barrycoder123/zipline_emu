
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_core_glue ( disable_debug_cmd_q, set_gcm_tag_fail_int, 
	set_txc_bp_int, set_rsm_is_backpressuring, .kme_ib_out( {
	\kme_ib_out.tready } ), .sa_snapshot( {
	\sa_snapshot[31].r.part1[31] , \sa_snapshot[31].r.part1[30] , 
	\sa_snapshot[31].r.part1[29] , \sa_snapshot[31].r.part1[28] , 
	\sa_snapshot[31].r.part1[27] , \sa_snapshot[31].r.part1[26] , 
	\sa_snapshot[31].r.part1[25] , \sa_snapshot[31].r.part1[24] , 
	\sa_snapshot[31].r.part1[23] , \sa_snapshot[31].r.part1[22] , 
	\sa_snapshot[31].r.part1[21] , \sa_snapshot[31].r.part1[20] , 
	\sa_snapshot[31].r.part1[19] , \sa_snapshot[31].r.part1[18] , 
	\sa_snapshot[31].r.part1[17] , \sa_snapshot[31].r.part1[16] , 
	\sa_snapshot[31].r.part1[15] , \sa_snapshot[31].r.part1[14] , 
	\sa_snapshot[31].r.part1[13] , \sa_snapshot[31].r.part1[12] , 
	\sa_snapshot[31].r.part1[11] , \sa_snapshot[31].r.part1[10] , 
	\sa_snapshot[31].r.part1[9] , \sa_snapshot[31].r.part1[8] , 
	\sa_snapshot[31].r.part1[7] , \sa_snapshot[31].r.part1[6] , 
	\sa_snapshot[31].r.part1[5] , \sa_snapshot[31].r.part1[4] , 
	\sa_snapshot[31].r.part1[3] , \sa_snapshot[31].r.part1[2] , 
	\sa_snapshot[31].r.part1[1] , \sa_snapshot[31].r.part1[0] , 
	\sa_snapshot[31].r.part0[31] , \sa_snapshot[31].r.part0[30] , 
	\sa_snapshot[31].r.part0[29] , \sa_snapshot[31].r.part0[28] , 
	\sa_snapshot[31].r.part0[27] , \sa_snapshot[31].r.part0[26] , 
	\sa_snapshot[31].r.part0[25] , \sa_snapshot[31].r.part0[24] , 
	\sa_snapshot[31].r.part0[23] , \sa_snapshot[31].r.part0[22] , 
	\sa_snapshot[31].r.part0[21] , \sa_snapshot[31].r.part0[20] , 
	\sa_snapshot[31].r.part0[19] , \sa_snapshot[31].r.part0[18] , 
	\sa_snapshot[31].r.part0[17] , \sa_snapshot[31].r.part0[16] , 
	\sa_snapshot[31].r.part0[15] , \sa_snapshot[31].r.part0[14] , 
	\sa_snapshot[31].r.part0[13] , \sa_snapshot[31].r.part0[12] , 
	\sa_snapshot[31].r.part0[11] , \sa_snapshot[31].r.part0[10] , 
	\sa_snapshot[31].r.part0[9] , \sa_snapshot[31].r.part0[8] , 
	\sa_snapshot[31].r.part0[7] , \sa_snapshot[31].r.part0[6] , 
	\sa_snapshot[31].r.part0[5] , \sa_snapshot[31].r.part0[4] , 
	\sa_snapshot[31].r.part0[3] , \sa_snapshot[31].r.part0[2] , 
	\sa_snapshot[31].r.part0[1] , \sa_snapshot[31].r.part0[0] , 
	\sa_snapshot[30].r.part1[31] , \sa_snapshot[30].r.part1[30] , 
	\sa_snapshot[30].r.part1[29] , \sa_snapshot[30].r.part1[28] , 
	\sa_snapshot[30].r.part1[27] , \sa_snapshot[30].r.part1[26] , 
	\sa_snapshot[30].r.part1[25] , \sa_snapshot[30].r.part1[24] , 
	\sa_snapshot[30].r.part1[23] , \sa_snapshot[30].r.part1[22] , 
	\sa_snapshot[30].r.part1[21] , \sa_snapshot[30].r.part1[20] , 
	\sa_snapshot[30].r.part1[19] , \sa_snapshot[30].r.part1[18] , 
	\sa_snapshot[30].r.part1[17] , \sa_snapshot[30].r.part1[16] , 
	\sa_snapshot[30].r.part1[15] , \sa_snapshot[30].r.part1[14] , 
	\sa_snapshot[30].r.part1[13] , \sa_snapshot[30].r.part1[12] , 
	\sa_snapshot[30].r.part1[11] , \sa_snapshot[30].r.part1[10] , 
	\sa_snapshot[30].r.part1[9] , \sa_snapshot[30].r.part1[8] , 
	\sa_snapshot[30].r.part1[7] , \sa_snapshot[30].r.part1[6] , 
	\sa_snapshot[30].r.part1[5] , \sa_snapshot[30].r.part1[4] , 
	\sa_snapshot[30].r.part1[3] , \sa_snapshot[30].r.part1[2] , 
	\sa_snapshot[30].r.part1[1] , \sa_snapshot[30].r.part1[0] , 
	\sa_snapshot[30].r.part0[31] , \sa_snapshot[30].r.part0[30] , 
	\sa_snapshot[30].r.part0[29] , \sa_snapshot[30].r.part0[28] , 
	\sa_snapshot[30].r.part0[27] , \sa_snapshot[30].r.part0[26] , 
	\sa_snapshot[30].r.part0[25] , \sa_snapshot[30].r.part0[24] , 
	\sa_snapshot[30].r.part0[23] , \sa_snapshot[30].r.part0[22] , 
	\sa_snapshot[30].r.part0[21] , \sa_snapshot[30].r.part0[20] , 
	\sa_snapshot[30].r.part0[19] , \sa_snapshot[30].r.part0[18] , 
	\sa_snapshot[30].r.part0[17] , \sa_snapshot[30].r.part0[16] , 
	\sa_snapshot[30].r.part0[15] , \sa_snapshot[30].r.part0[14] , 
	\sa_snapshot[30].r.part0[13] , \sa_snapshot[30].r.part0[12] , 
	\sa_snapshot[30].r.part0[11] , \sa_snapshot[30].r.part0[10] , 
	\sa_snapshot[30].r.part0[9] , \sa_snapshot[30].r.part0[8] , 
	\sa_snapshot[30].r.part0[7] , \sa_snapshot[30].r.part0[6] , 
	\sa_snapshot[30].r.part0[5] , \sa_snapshot[30].r.part0[4] , 
	\sa_snapshot[30].r.part0[3] , \sa_snapshot[30].r.part0[2] , 
	\sa_snapshot[30].r.part0[1] , \sa_snapshot[30].r.part0[0] , 
	\sa_snapshot[29].r.part1[31] , \sa_snapshot[29].r.part1[30] , 
	\sa_snapshot[29].r.part1[29] , \sa_snapshot[29].r.part1[28] , 
	\sa_snapshot[29].r.part1[27] , \sa_snapshot[29].r.part1[26] , 
	\sa_snapshot[29].r.part1[25] , \sa_snapshot[29].r.part1[24] , 
	\sa_snapshot[29].r.part1[23] , \sa_snapshot[29].r.part1[22] , 
	\sa_snapshot[29].r.part1[21] , \sa_snapshot[29].r.part1[20] , 
	\sa_snapshot[29].r.part1[19] , \sa_snapshot[29].r.part1[18] , 
	\sa_snapshot[29].r.part1[17] , \sa_snapshot[29].r.part1[16] , 
	\sa_snapshot[29].r.part1[15] , \sa_snapshot[29].r.part1[14] , 
	\sa_snapshot[29].r.part1[13] , \sa_snapshot[29].r.part1[12] , 
	\sa_snapshot[29].r.part1[11] , \sa_snapshot[29].r.part1[10] , 
	\sa_snapshot[29].r.part1[9] , \sa_snapshot[29].r.part1[8] , 
	\sa_snapshot[29].r.part1[7] , \sa_snapshot[29].r.part1[6] , 
	\sa_snapshot[29].r.part1[5] , \sa_snapshot[29].r.part1[4] , 
	\sa_snapshot[29].r.part1[3] , \sa_snapshot[29].r.part1[2] , 
	\sa_snapshot[29].r.part1[1] , \sa_snapshot[29].r.part1[0] , 
	\sa_snapshot[29].r.part0[31] , \sa_snapshot[29].r.part0[30] , 
	\sa_snapshot[29].r.part0[29] , \sa_snapshot[29].r.part0[28] , 
	\sa_snapshot[29].r.part0[27] , \sa_snapshot[29].r.part0[26] , 
	\sa_snapshot[29].r.part0[25] , \sa_snapshot[29].r.part0[24] , 
	\sa_snapshot[29].r.part0[23] , \sa_snapshot[29].r.part0[22] , 
	\sa_snapshot[29].r.part0[21] , \sa_snapshot[29].r.part0[20] , 
	\sa_snapshot[29].r.part0[19] , \sa_snapshot[29].r.part0[18] , 
	\sa_snapshot[29].r.part0[17] , \sa_snapshot[29].r.part0[16] , 
	\sa_snapshot[29].r.part0[15] , \sa_snapshot[29].r.part0[14] , 
	\sa_snapshot[29].r.part0[13] , \sa_snapshot[29].r.part0[12] , 
	\sa_snapshot[29].r.part0[11] , \sa_snapshot[29].r.part0[10] , 
	\sa_snapshot[29].r.part0[9] , \sa_snapshot[29].r.part0[8] , 
	\sa_snapshot[29].r.part0[7] , \sa_snapshot[29].r.part0[6] , 
	\sa_snapshot[29].r.part0[5] , \sa_snapshot[29].r.part0[4] , 
	\sa_snapshot[29].r.part0[3] , \sa_snapshot[29].r.part0[2] , 
	\sa_snapshot[29].r.part0[1] , \sa_snapshot[29].r.part0[0] , 
	\sa_snapshot[28].r.part1[31] , \sa_snapshot[28].r.part1[30] , 
	\sa_snapshot[28].r.part1[29] , \sa_snapshot[28].r.part1[28] , 
	\sa_snapshot[28].r.part1[27] , \sa_snapshot[28].r.part1[26] , 
	\sa_snapshot[28].r.part1[25] , \sa_snapshot[28].r.part1[24] , 
	\sa_snapshot[28].r.part1[23] , \sa_snapshot[28].r.part1[22] , 
	\sa_snapshot[28].r.part1[21] , \sa_snapshot[28].r.part1[20] , 
	\sa_snapshot[28].r.part1[19] , \sa_snapshot[28].r.part1[18] , 
	\sa_snapshot[28].r.part1[17] , \sa_snapshot[28].r.part1[16] , 
	\sa_snapshot[28].r.part1[15] , \sa_snapshot[28].r.part1[14] , 
	\sa_snapshot[28].r.part1[13] , \sa_snapshot[28].r.part1[12] , 
	\sa_snapshot[28].r.part1[11] , \sa_snapshot[28].r.part1[10] , 
	\sa_snapshot[28].r.part1[9] , \sa_snapshot[28].r.part1[8] , 
	\sa_snapshot[28].r.part1[7] , \sa_snapshot[28].r.part1[6] , 
	\sa_snapshot[28].r.part1[5] , \sa_snapshot[28].r.part1[4] , 
	\sa_snapshot[28].r.part1[3] , \sa_snapshot[28].r.part1[2] , 
	\sa_snapshot[28].r.part1[1] , \sa_snapshot[28].r.part1[0] , 
	\sa_snapshot[28].r.part0[31] , \sa_snapshot[28].r.part0[30] , 
	\sa_snapshot[28].r.part0[29] , \sa_snapshot[28].r.part0[28] , 
	\sa_snapshot[28].r.part0[27] , \sa_snapshot[28].r.part0[26] , 
	\sa_snapshot[28].r.part0[25] , \sa_snapshot[28].r.part0[24] , 
	\sa_snapshot[28].r.part0[23] , \sa_snapshot[28].r.part0[22] , 
	\sa_snapshot[28].r.part0[21] , \sa_snapshot[28].r.part0[20] , 
	\sa_snapshot[28].r.part0[19] , \sa_snapshot[28].r.part0[18] , 
	\sa_snapshot[28].r.part0[17] , \sa_snapshot[28].r.part0[16] , 
	\sa_snapshot[28].r.part0[15] , \sa_snapshot[28].r.part0[14] , 
	\sa_snapshot[28].r.part0[13] , \sa_snapshot[28].r.part0[12] , 
	\sa_snapshot[28].r.part0[11] , \sa_snapshot[28].r.part0[10] , 
	\sa_snapshot[28].r.part0[9] , \sa_snapshot[28].r.part0[8] , 
	\sa_snapshot[28].r.part0[7] , \sa_snapshot[28].r.part0[6] , 
	\sa_snapshot[28].r.part0[5] , \sa_snapshot[28].r.part0[4] , 
	\sa_snapshot[28].r.part0[3] , \sa_snapshot[28].r.part0[2] , 
	\sa_snapshot[28].r.part0[1] , \sa_snapshot[28].r.part0[0] , 
	\sa_snapshot[27].r.part1[31] , \sa_snapshot[27].r.part1[30] , 
	\sa_snapshot[27].r.part1[29] , \sa_snapshot[27].r.part1[28] , 
	\sa_snapshot[27].r.part1[27] , \sa_snapshot[27].r.part1[26] , 
	\sa_snapshot[27].r.part1[25] , \sa_snapshot[27].r.part1[24] , 
	\sa_snapshot[27].r.part1[23] , \sa_snapshot[27].r.part1[22] , 
	\sa_snapshot[27].r.part1[21] , \sa_snapshot[27].r.part1[20] , 
	\sa_snapshot[27].r.part1[19] , \sa_snapshot[27].r.part1[18] , 
	\sa_snapshot[27].r.part1[17] , \sa_snapshot[27].r.part1[16] , 
	\sa_snapshot[27].r.part1[15] , \sa_snapshot[27].r.part1[14] , 
	\sa_snapshot[27].r.part1[13] , \sa_snapshot[27].r.part1[12] , 
	\sa_snapshot[27].r.part1[11] , \sa_snapshot[27].r.part1[10] , 
	\sa_snapshot[27].r.part1[9] , \sa_snapshot[27].r.part1[8] , 
	\sa_snapshot[27].r.part1[7] , \sa_snapshot[27].r.part1[6] , 
	\sa_snapshot[27].r.part1[5] , \sa_snapshot[27].r.part1[4] , 
	\sa_snapshot[27].r.part1[3] , \sa_snapshot[27].r.part1[2] , 
	\sa_snapshot[27].r.part1[1] , \sa_snapshot[27].r.part1[0] , 
	\sa_snapshot[27].r.part0[31] , \sa_snapshot[27].r.part0[30] , 
	\sa_snapshot[27].r.part0[29] , \sa_snapshot[27].r.part0[28] , 
	\sa_snapshot[27].r.part0[27] , \sa_snapshot[27].r.part0[26] , 
	\sa_snapshot[27].r.part0[25] , \sa_snapshot[27].r.part0[24] , 
	\sa_snapshot[27].r.part0[23] , \sa_snapshot[27].r.part0[22] , 
	\sa_snapshot[27].r.part0[21] , \sa_snapshot[27].r.part0[20] , 
	\sa_snapshot[27].r.part0[19] , \sa_snapshot[27].r.part0[18] , 
	\sa_snapshot[27].r.part0[17] , \sa_snapshot[27].r.part0[16] , 
	\sa_snapshot[27].r.part0[15] , \sa_snapshot[27].r.part0[14] , 
	\sa_snapshot[27].r.part0[13] , \sa_snapshot[27].r.part0[12] , 
	\sa_snapshot[27].r.part0[11] , \sa_snapshot[27].r.part0[10] , 
	\sa_snapshot[27].r.part0[9] , \sa_snapshot[27].r.part0[8] , 
	\sa_snapshot[27].r.part0[7] , \sa_snapshot[27].r.part0[6] , 
	\sa_snapshot[27].r.part0[5] , \sa_snapshot[27].r.part0[4] , 
	\sa_snapshot[27].r.part0[3] , \sa_snapshot[27].r.part0[2] , 
	\sa_snapshot[27].r.part0[1] , \sa_snapshot[27].r.part0[0] , 
	\sa_snapshot[26].r.part1[31] , \sa_snapshot[26].r.part1[30] , 
	\sa_snapshot[26].r.part1[29] , \sa_snapshot[26].r.part1[28] , 
	\sa_snapshot[26].r.part1[27] , \sa_snapshot[26].r.part1[26] , 
	\sa_snapshot[26].r.part1[25] , \sa_snapshot[26].r.part1[24] , 
	\sa_snapshot[26].r.part1[23] , \sa_snapshot[26].r.part1[22] , 
	\sa_snapshot[26].r.part1[21] , \sa_snapshot[26].r.part1[20] , 
	\sa_snapshot[26].r.part1[19] , \sa_snapshot[26].r.part1[18] , 
	\sa_snapshot[26].r.part1[17] , \sa_snapshot[26].r.part1[16] , 
	\sa_snapshot[26].r.part1[15] , \sa_snapshot[26].r.part1[14] , 
	\sa_snapshot[26].r.part1[13] , \sa_snapshot[26].r.part1[12] , 
	\sa_snapshot[26].r.part1[11] , \sa_snapshot[26].r.part1[10] , 
	\sa_snapshot[26].r.part1[9] , \sa_snapshot[26].r.part1[8] , 
	\sa_snapshot[26].r.part1[7] , \sa_snapshot[26].r.part1[6] , 
	\sa_snapshot[26].r.part1[5] , \sa_snapshot[26].r.part1[4] , 
	\sa_snapshot[26].r.part1[3] , \sa_snapshot[26].r.part1[2] , 
	\sa_snapshot[26].r.part1[1] , \sa_snapshot[26].r.part1[0] , 
	\sa_snapshot[26].r.part0[31] , \sa_snapshot[26].r.part0[30] , 
	\sa_snapshot[26].r.part0[29] , \sa_snapshot[26].r.part0[28] , 
	\sa_snapshot[26].r.part0[27] , \sa_snapshot[26].r.part0[26] , 
	\sa_snapshot[26].r.part0[25] , \sa_snapshot[26].r.part0[24] , 
	\sa_snapshot[26].r.part0[23] , \sa_snapshot[26].r.part0[22] , 
	\sa_snapshot[26].r.part0[21] , \sa_snapshot[26].r.part0[20] , 
	\sa_snapshot[26].r.part0[19] , \sa_snapshot[26].r.part0[18] , 
	\sa_snapshot[26].r.part0[17] , \sa_snapshot[26].r.part0[16] , 
	\sa_snapshot[26].r.part0[15] , \sa_snapshot[26].r.part0[14] , 
	\sa_snapshot[26].r.part0[13] , \sa_snapshot[26].r.part0[12] , 
	\sa_snapshot[26].r.part0[11] , \sa_snapshot[26].r.part0[10] , 
	\sa_snapshot[26].r.part0[9] , \sa_snapshot[26].r.part0[8] , 
	\sa_snapshot[26].r.part0[7] , \sa_snapshot[26].r.part0[6] , 
	\sa_snapshot[26].r.part0[5] , \sa_snapshot[26].r.part0[4] , 
	\sa_snapshot[26].r.part0[3] , \sa_snapshot[26].r.part0[2] , 
	\sa_snapshot[26].r.part0[1] , \sa_snapshot[26].r.part0[0] , 
	\sa_snapshot[25].r.part1[31] , \sa_snapshot[25].r.part1[30] , 
	\sa_snapshot[25].r.part1[29] , \sa_snapshot[25].r.part1[28] , 
	\sa_snapshot[25].r.part1[27] , \sa_snapshot[25].r.part1[26] , 
	\sa_snapshot[25].r.part1[25] , \sa_snapshot[25].r.part1[24] , 
	\sa_snapshot[25].r.part1[23] , \sa_snapshot[25].r.part1[22] , 
	\sa_snapshot[25].r.part1[21] , \sa_snapshot[25].r.part1[20] , 
	\sa_snapshot[25].r.part1[19] , \sa_snapshot[25].r.part1[18] , 
	\sa_snapshot[25].r.part1[17] , \sa_snapshot[25].r.part1[16] , 
	\sa_snapshot[25].r.part1[15] , \sa_snapshot[25].r.part1[14] , 
	\sa_snapshot[25].r.part1[13] , \sa_snapshot[25].r.part1[12] , 
	\sa_snapshot[25].r.part1[11] , \sa_snapshot[25].r.part1[10] , 
	\sa_snapshot[25].r.part1[9] , \sa_snapshot[25].r.part1[8] , 
	\sa_snapshot[25].r.part1[7] , \sa_snapshot[25].r.part1[6] , 
	\sa_snapshot[25].r.part1[5] , \sa_snapshot[25].r.part1[4] , 
	\sa_snapshot[25].r.part1[3] , \sa_snapshot[25].r.part1[2] , 
	\sa_snapshot[25].r.part1[1] , \sa_snapshot[25].r.part1[0] , 
	\sa_snapshot[25].r.part0[31] , \sa_snapshot[25].r.part0[30] , 
	\sa_snapshot[25].r.part0[29] , \sa_snapshot[25].r.part0[28] , 
	\sa_snapshot[25].r.part0[27] , \sa_snapshot[25].r.part0[26] , 
	\sa_snapshot[25].r.part0[25] , \sa_snapshot[25].r.part0[24] , 
	\sa_snapshot[25].r.part0[23] , \sa_snapshot[25].r.part0[22] , 
	\sa_snapshot[25].r.part0[21] , \sa_snapshot[25].r.part0[20] , 
	\sa_snapshot[25].r.part0[19] , \sa_snapshot[25].r.part0[18] , 
	\sa_snapshot[25].r.part0[17] , \sa_snapshot[25].r.part0[16] , 
	\sa_snapshot[25].r.part0[15] , \sa_snapshot[25].r.part0[14] , 
	\sa_snapshot[25].r.part0[13] , \sa_snapshot[25].r.part0[12] , 
	\sa_snapshot[25].r.part0[11] , \sa_snapshot[25].r.part0[10] , 
	\sa_snapshot[25].r.part0[9] , \sa_snapshot[25].r.part0[8] , 
	\sa_snapshot[25].r.part0[7] , \sa_snapshot[25].r.part0[6] , 
	\sa_snapshot[25].r.part0[5] , \sa_snapshot[25].r.part0[4] , 
	\sa_snapshot[25].r.part0[3] , \sa_snapshot[25].r.part0[2] , 
	\sa_snapshot[25].r.part0[1] , \sa_snapshot[25].r.part0[0] , 
	\sa_snapshot[24].r.part1[31] , \sa_snapshot[24].r.part1[30] , 
	\sa_snapshot[24].r.part1[29] , \sa_snapshot[24].r.part1[28] , 
	\sa_snapshot[24].r.part1[27] , \sa_snapshot[24].r.part1[26] , 
	\sa_snapshot[24].r.part1[25] , \sa_snapshot[24].r.part1[24] , 
	\sa_snapshot[24].r.part1[23] , \sa_snapshot[24].r.part1[22] , 
	\sa_snapshot[24].r.part1[21] , \sa_snapshot[24].r.part1[20] , 
	\sa_snapshot[24].r.part1[19] , \sa_snapshot[24].r.part1[18] , 
	\sa_snapshot[24].r.part1[17] , \sa_snapshot[24].r.part1[16] , 
	\sa_snapshot[24].r.part1[15] , \sa_snapshot[24].r.part1[14] , 
	\sa_snapshot[24].r.part1[13] , \sa_snapshot[24].r.part1[12] , 
	\sa_snapshot[24].r.part1[11] , \sa_snapshot[24].r.part1[10] , 
	\sa_snapshot[24].r.part1[9] , \sa_snapshot[24].r.part1[8] , 
	\sa_snapshot[24].r.part1[7] , \sa_snapshot[24].r.part1[6] , 
	\sa_snapshot[24].r.part1[5] , \sa_snapshot[24].r.part1[4] , 
	\sa_snapshot[24].r.part1[3] , \sa_snapshot[24].r.part1[2] , 
	\sa_snapshot[24].r.part1[1] , \sa_snapshot[24].r.part1[0] , 
	\sa_snapshot[24].r.part0[31] , \sa_snapshot[24].r.part0[30] , 
	\sa_snapshot[24].r.part0[29] , \sa_snapshot[24].r.part0[28] , 
	\sa_snapshot[24].r.part0[27] , \sa_snapshot[24].r.part0[26] , 
	\sa_snapshot[24].r.part0[25] , \sa_snapshot[24].r.part0[24] , 
	\sa_snapshot[24].r.part0[23] , \sa_snapshot[24].r.part0[22] , 
	\sa_snapshot[24].r.part0[21] , \sa_snapshot[24].r.part0[20] , 
	\sa_snapshot[24].r.part0[19] , \sa_snapshot[24].r.part0[18] , 
	\sa_snapshot[24].r.part0[17] , \sa_snapshot[24].r.part0[16] , 
	\sa_snapshot[24].r.part0[15] , \sa_snapshot[24].r.part0[14] , 
	\sa_snapshot[24].r.part0[13] , \sa_snapshot[24].r.part0[12] , 
	\sa_snapshot[24].r.part0[11] , \sa_snapshot[24].r.part0[10] , 
	\sa_snapshot[24].r.part0[9] , \sa_snapshot[24].r.part0[8] , 
	\sa_snapshot[24].r.part0[7] , \sa_snapshot[24].r.part0[6] , 
	\sa_snapshot[24].r.part0[5] , \sa_snapshot[24].r.part0[4] , 
	\sa_snapshot[24].r.part0[3] , \sa_snapshot[24].r.part0[2] , 
	\sa_snapshot[24].r.part0[1] , \sa_snapshot[24].r.part0[0] , 
	\sa_snapshot[23].r.part1[31] , \sa_snapshot[23].r.part1[30] , 
	\sa_snapshot[23].r.part1[29] , \sa_snapshot[23].r.part1[28] , 
	\sa_snapshot[23].r.part1[27] , \sa_snapshot[23].r.part1[26] , 
	\sa_snapshot[23].r.part1[25] , \sa_snapshot[23].r.part1[24] , 
	\sa_snapshot[23].r.part1[23] , \sa_snapshot[23].r.part1[22] , 
	\sa_snapshot[23].r.part1[21] , \sa_snapshot[23].r.part1[20] , 
	\sa_snapshot[23].r.part1[19] , \sa_snapshot[23].r.part1[18] , 
	\sa_snapshot[23].r.part1[17] , \sa_snapshot[23].r.part1[16] , 
	\sa_snapshot[23].r.part1[15] , \sa_snapshot[23].r.part1[14] , 
	\sa_snapshot[23].r.part1[13] , \sa_snapshot[23].r.part1[12] , 
	\sa_snapshot[23].r.part1[11] , \sa_snapshot[23].r.part1[10] , 
	\sa_snapshot[23].r.part1[9] , \sa_snapshot[23].r.part1[8] , 
	\sa_snapshot[23].r.part1[7] , \sa_snapshot[23].r.part1[6] , 
	\sa_snapshot[23].r.part1[5] , \sa_snapshot[23].r.part1[4] , 
	\sa_snapshot[23].r.part1[3] , \sa_snapshot[23].r.part1[2] , 
	\sa_snapshot[23].r.part1[1] , \sa_snapshot[23].r.part1[0] , 
	\sa_snapshot[23].r.part0[31] , \sa_snapshot[23].r.part0[30] , 
	\sa_snapshot[23].r.part0[29] , \sa_snapshot[23].r.part0[28] , 
	\sa_snapshot[23].r.part0[27] , \sa_snapshot[23].r.part0[26] , 
	\sa_snapshot[23].r.part0[25] , \sa_snapshot[23].r.part0[24] , 
	\sa_snapshot[23].r.part0[23] , \sa_snapshot[23].r.part0[22] , 
	\sa_snapshot[23].r.part0[21] , \sa_snapshot[23].r.part0[20] , 
	\sa_snapshot[23].r.part0[19] , \sa_snapshot[23].r.part0[18] , 
	\sa_snapshot[23].r.part0[17] , \sa_snapshot[23].r.part0[16] , 
	\sa_snapshot[23].r.part0[15] , \sa_snapshot[23].r.part0[14] , 
	\sa_snapshot[23].r.part0[13] , \sa_snapshot[23].r.part0[12] , 
	\sa_snapshot[23].r.part0[11] , \sa_snapshot[23].r.part0[10] , 
	\sa_snapshot[23].r.part0[9] , \sa_snapshot[23].r.part0[8] , 
	\sa_snapshot[23].r.part0[7] , \sa_snapshot[23].r.part0[6] , 
	\sa_snapshot[23].r.part0[5] , \sa_snapshot[23].r.part0[4] , 
	\sa_snapshot[23].r.part0[3] , \sa_snapshot[23].r.part0[2] , 
	\sa_snapshot[23].r.part0[1] , \sa_snapshot[23].r.part0[0] , 
	\sa_snapshot[22].r.part1[31] , \sa_snapshot[22].r.part1[30] , 
	\sa_snapshot[22].r.part1[29] , \sa_snapshot[22].r.part1[28] , 
	\sa_snapshot[22].r.part1[27] , \sa_snapshot[22].r.part1[26] , 
	\sa_snapshot[22].r.part1[25] , \sa_snapshot[22].r.part1[24] , 
	\sa_snapshot[22].r.part1[23] , \sa_snapshot[22].r.part1[22] , 
	\sa_snapshot[22].r.part1[21] , \sa_snapshot[22].r.part1[20] , 
	\sa_snapshot[22].r.part1[19] , \sa_snapshot[22].r.part1[18] , 
	\sa_snapshot[22].r.part1[17] , \sa_snapshot[22].r.part1[16] , 
	\sa_snapshot[22].r.part1[15] , \sa_snapshot[22].r.part1[14] , 
	\sa_snapshot[22].r.part1[13] , \sa_snapshot[22].r.part1[12] , 
	\sa_snapshot[22].r.part1[11] , \sa_snapshot[22].r.part1[10] , 
	\sa_snapshot[22].r.part1[9] , \sa_snapshot[22].r.part1[8] , 
	\sa_snapshot[22].r.part1[7] , \sa_snapshot[22].r.part1[6] , 
	\sa_snapshot[22].r.part1[5] , \sa_snapshot[22].r.part1[4] , 
	\sa_snapshot[22].r.part1[3] , \sa_snapshot[22].r.part1[2] , 
	\sa_snapshot[22].r.part1[1] , \sa_snapshot[22].r.part1[0] , 
	\sa_snapshot[22].r.part0[31] , \sa_snapshot[22].r.part0[30] , 
	\sa_snapshot[22].r.part0[29] , \sa_snapshot[22].r.part0[28] , 
	\sa_snapshot[22].r.part0[27] , \sa_snapshot[22].r.part0[26] , 
	\sa_snapshot[22].r.part0[25] , \sa_snapshot[22].r.part0[24] , 
	\sa_snapshot[22].r.part0[23] , \sa_snapshot[22].r.part0[22] , 
	\sa_snapshot[22].r.part0[21] , \sa_snapshot[22].r.part0[20] , 
	\sa_snapshot[22].r.part0[19] , \sa_snapshot[22].r.part0[18] , 
	\sa_snapshot[22].r.part0[17] , \sa_snapshot[22].r.part0[16] , 
	\sa_snapshot[22].r.part0[15] , \sa_snapshot[22].r.part0[14] , 
	\sa_snapshot[22].r.part0[13] , \sa_snapshot[22].r.part0[12] , 
	\sa_snapshot[22].r.part0[11] , \sa_snapshot[22].r.part0[10] , 
	\sa_snapshot[22].r.part0[9] , \sa_snapshot[22].r.part0[8] , 
	\sa_snapshot[22].r.part0[7] , \sa_snapshot[22].r.part0[6] , 
	\sa_snapshot[22].r.part0[5] , \sa_snapshot[22].r.part0[4] , 
	\sa_snapshot[22].r.part0[3] , \sa_snapshot[22].r.part0[2] , 
	\sa_snapshot[22].r.part0[1] , \sa_snapshot[22].r.part0[0] , 
	\sa_snapshot[21].r.part1[31] , \sa_snapshot[21].r.part1[30] , 
	\sa_snapshot[21].r.part1[29] , \sa_snapshot[21].r.part1[28] , 
	\sa_snapshot[21].r.part1[27] , \sa_snapshot[21].r.part1[26] , 
	\sa_snapshot[21].r.part1[25] , \sa_snapshot[21].r.part1[24] , 
	\sa_snapshot[21].r.part1[23] , \sa_snapshot[21].r.part1[22] , 
	\sa_snapshot[21].r.part1[21] , \sa_snapshot[21].r.part1[20] , 
	\sa_snapshot[21].r.part1[19] , \sa_snapshot[21].r.part1[18] , 
	\sa_snapshot[21].r.part1[17] , \sa_snapshot[21].r.part1[16] , 
	\sa_snapshot[21].r.part1[15] , \sa_snapshot[21].r.part1[14] , 
	\sa_snapshot[21].r.part1[13] , \sa_snapshot[21].r.part1[12] , 
	\sa_snapshot[21].r.part1[11] , \sa_snapshot[21].r.part1[10] , 
	\sa_snapshot[21].r.part1[9] , \sa_snapshot[21].r.part1[8] , 
	\sa_snapshot[21].r.part1[7] , \sa_snapshot[21].r.part1[6] , 
	\sa_snapshot[21].r.part1[5] , \sa_snapshot[21].r.part1[4] , 
	\sa_snapshot[21].r.part1[3] , \sa_snapshot[21].r.part1[2] , 
	\sa_snapshot[21].r.part1[1] , \sa_snapshot[21].r.part1[0] , 
	\sa_snapshot[21].r.part0[31] , \sa_snapshot[21].r.part0[30] , 
	\sa_snapshot[21].r.part0[29] , \sa_snapshot[21].r.part0[28] , 
	\sa_snapshot[21].r.part0[27] , \sa_snapshot[21].r.part0[26] , 
	\sa_snapshot[21].r.part0[25] , \sa_snapshot[21].r.part0[24] , 
	\sa_snapshot[21].r.part0[23] , \sa_snapshot[21].r.part0[22] , 
	\sa_snapshot[21].r.part0[21] , \sa_snapshot[21].r.part0[20] , 
	\sa_snapshot[21].r.part0[19] , \sa_snapshot[21].r.part0[18] , 
	\sa_snapshot[21].r.part0[17] , \sa_snapshot[21].r.part0[16] , 
	\sa_snapshot[21].r.part0[15] , \sa_snapshot[21].r.part0[14] , 
	\sa_snapshot[21].r.part0[13] , \sa_snapshot[21].r.part0[12] , 
	\sa_snapshot[21].r.part0[11] , \sa_snapshot[21].r.part0[10] , 
	\sa_snapshot[21].r.part0[9] , \sa_snapshot[21].r.part0[8] , 
	\sa_snapshot[21].r.part0[7] , \sa_snapshot[21].r.part0[6] , 
	\sa_snapshot[21].r.part0[5] , \sa_snapshot[21].r.part0[4] , 
	\sa_snapshot[21].r.part0[3] , \sa_snapshot[21].r.part0[2] , 
	\sa_snapshot[21].r.part0[1] , \sa_snapshot[21].r.part0[0] , 
	\sa_snapshot[20].r.part1[31] , \sa_snapshot[20].r.part1[30] , 
	\sa_snapshot[20].r.part1[29] , \sa_snapshot[20].r.part1[28] , 
	\sa_snapshot[20].r.part1[27] , \sa_snapshot[20].r.part1[26] , 
	\sa_snapshot[20].r.part1[25] , \sa_snapshot[20].r.part1[24] , 
	\sa_snapshot[20].r.part1[23] , \sa_snapshot[20].r.part1[22] , 
	\sa_snapshot[20].r.part1[21] , \sa_snapshot[20].r.part1[20] , 
	\sa_snapshot[20].r.part1[19] , \sa_snapshot[20].r.part1[18] , 
	\sa_snapshot[20].r.part1[17] , \sa_snapshot[20].r.part1[16] , 
	\sa_snapshot[20].r.part1[15] , \sa_snapshot[20].r.part1[14] , 
	\sa_snapshot[20].r.part1[13] , \sa_snapshot[20].r.part1[12] , 
	\sa_snapshot[20].r.part1[11] , \sa_snapshot[20].r.part1[10] , 
	\sa_snapshot[20].r.part1[9] , \sa_snapshot[20].r.part1[8] , 
	\sa_snapshot[20].r.part1[7] , \sa_snapshot[20].r.part1[6] , 
	\sa_snapshot[20].r.part1[5] , \sa_snapshot[20].r.part1[4] , 
	\sa_snapshot[20].r.part1[3] , \sa_snapshot[20].r.part1[2] , 
	\sa_snapshot[20].r.part1[1] , \sa_snapshot[20].r.part1[0] , 
	\sa_snapshot[20].r.part0[31] , \sa_snapshot[20].r.part0[30] , 
	\sa_snapshot[20].r.part0[29] , \sa_snapshot[20].r.part0[28] , 
	\sa_snapshot[20].r.part0[27] , \sa_snapshot[20].r.part0[26] , 
	\sa_snapshot[20].r.part0[25] , \sa_snapshot[20].r.part0[24] , 
	\sa_snapshot[20].r.part0[23] , \sa_snapshot[20].r.part0[22] , 
	\sa_snapshot[20].r.part0[21] , \sa_snapshot[20].r.part0[20] , 
	\sa_snapshot[20].r.part0[19] , \sa_snapshot[20].r.part0[18] , 
	\sa_snapshot[20].r.part0[17] , \sa_snapshot[20].r.part0[16] , 
	\sa_snapshot[20].r.part0[15] , \sa_snapshot[20].r.part0[14] , 
	\sa_snapshot[20].r.part0[13] , \sa_snapshot[20].r.part0[12] , 
	\sa_snapshot[20].r.part0[11] , \sa_snapshot[20].r.part0[10] , 
	\sa_snapshot[20].r.part0[9] , \sa_snapshot[20].r.part0[8] , 
	\sa_snapshot[20].r.part0[7] , \sa_snapshot[20].r.part0[6] , 
	\sa_snapshot[20].r.part0[5] , \sa_snapshot[20].r.part0[4] , 
	\sa_snapshot[20].r.part0[3] , \sa_snapshot[20].r.part0[2] , 
	\sa_snapshot[20].r.part0[1] , \sa_snapshot[20].r.part0[0] , 
	\sa_snapshot[19].r.part1[31] , \sa_snapshot[19].r.part1[30] , 
	\sa_snapshot[19].r.part1[29] , \sa_snapshot[19].r.part1[28] , 
	\sa_snapshot[19].r.part1[27] , \sa_snapshot[19].r.part1[26] , 
	\sa_snapshot[19].r.part1[25] , \sa_snapshot[19].r.part1[24] , 
	\sa_snapshot[19].r.part1[23] , \sa_snapshot[19].r.part1[22] , 
	\sa_snapshot[19].r.part1[21] , \sa_snapshot[19].r.part1[20] , 
	\sa_snapshot[19].r.part1[19] , \sa_snapshot[19].r.part1[18] , 
	\sa_snapshot[19].r.part1[17] , \sa_snapshot[19].r.part1[16] , 
	\sa_snapshot[19].r.part1[15] , \sa_snapshot[19].r.part1[14] , 
	\sa_snapshot[19].r.part1[13] , \sa_snapshot[19].r.part1[12] , 
	\sa_snapshot[19].r.part1[11] , \sa_snapshot[19].r.part1[10] , 
	\sa_snapshot[19].r.part1[9] , \sa_snapshot[19].r.part1[8] , 
	\sa_snapshot[19].r.part1[7] , \sa_snapshot[19].r.part1[6] , 
	\sa_snapshot[19].r.part1[5] , \sa_snapshot[19].r.part1[4] , 
	\sa_snapshot[19].r.part1[3] , \sa_snapshot[19].r.part1[2] , 
	\sa_snapshot[19].r.part1[1] , \sa_snapshot[19].r.part1[0] , 
	\sa_snapshot[19].r.part0[31] , \sa_snapshot[19].r.part0[30] , 
	\sa_snapshot[19].r.part0[29] , \sa_snapshot[19].r.part0[28] , 
	\sa_snapshot[19].r.part0[27] , \sa_snapshot[19].r.part0[26] , 
	\sa_snapshot[19].r.part0[25] , \sa_snapshot[19].r.part0[24] , 
	\sa_snapshot[19].r.part0[23] , \sa_snapshot[19].r.part0[22] , 
	\sa_snapshot[19].r.part0[21] , \sa_snapshot[19].r.part0[20] , 
	\sa_snapshot[19].r.part0[19] , \sa_snapshot[19].r.part0[18] , 
	\sa_snapshot[19].r.part0[17] , \sa_snapshot[19].r.part0[16] , 
	\sa_snapshot[19].r.part0[15] , \sa_snapshot[19].r.part0[14] , 
	\sa_snapshot[19].r.part0[13] , \sa_snapshot[19].r.part0[12] , 
	\sa_snapshot[19].r.part0[11] , \sa_snapshot[19].r.part0[10] , 
	\sa_snapshot[19].r.part0[9] , \sa_snapshot[19].r.part0[8] , 
	\sa_snapshot[19].r.part0[7] , \sa_snapshot[19].r.part0[6] , 
	\sa_snapshot[19].r.part0[5] , \sa_snapshot[19].r.part0[4] , 
	\sa_snapshot[19].r.part0[3] , \sa_snapshot[19].r.part0[2] , 
	\sa_snapshot[19].r.part0[1] , \sa_snapshot[19].r.part0[0] , 
	\sa_snapshot[18].r.part1[31] , \sa_snapshot[18].r.part1[30] , 
	\sa_snapshot[18].r.part1[29] , \sa_snapshot[18].r.part1[28] , 
	\sa_snapshot[18].r.part1[27] , \sa_snapshot[18].r.part1[26] , 
	\sa_snapshot[18].r.part1[25] , \sa_snapshot[18].r.part1[24] , 
	\sa_snapshot[18].r.part1[23] , \sa_snapshot[18].r.part1[22] , 
	\sa_snapshot[18].r.part1[21] , \sa_snapshot[18].r.part1[20] , 
	\sa_snapshot[18].r.part1[19] , \sa_snapshot[18].r.part1[18] , 
	\sa_snapshot[18].r.part1[17] , \sa_snapshot[18].r.part1[16] , 
	\sa_snapshot[18].r.part1[15] , \sa_snapshot[18].r.part1[14] , 
	\sa_snapshot[18].r.part1[13] , \sa_snapshot[18].r.part1[12] , 
	\sa_snapshot[18].r.part1[11] , \sa_snapshot[18].r.part1[10] , 
	\sa_snapshot[18].r.part1[9] , \sa_snapshot[18].r.part1[8] , 
	\sa_snapshot[18].r.part1[7] , \sa_snapshot[18].r.part1[6] , 
	\sa_snapshot[18].r.part1[5] , \sa_snapshot[18].r.part1[4] , 
	\sa_snapshot[18].r.part1[3] , \sa_snapshot[18].r.part1[2] , 
	\sa_snapshot[18].r.part1[1] , \sa_snapshot[18].r.part1[0] , 
	\sa_snapshot[18].r.part0[31] , \sa_snapshot[18].r.part0[30] , 
	\sa_snapshot[18].r.part0[29] , \sa_snapshot[18].r.part0[28] , 
	\sa_snapshot[18].r.part0[27] , \sa_snapshot[18].r.part0[26] , 
	\sa_snapshot[18].r.part0[25] , \sa_snapshot[18].r.part0[24] , 
	\sa_snapshot[18].r.part0[23] , \sa_snapshot[18].r.part0[22] , 
	\sa_snapshot[18].r.part0[21] , \sa_snapshot[18].r.part0[20] , 
	\sa_snapshot[18].r.part0[19] , \sa_snapshot[18].r.part0[18] , 
	\sa_snapshot[18].r.part0[17] , \sa_snapshot[18].r.part0[16] , 
	\sa_snapshot[18].r.part0[15] , \sa_snapshot[18].r.part0[14] , 
	\sa_snapshot[18].r.part0[13] , \sa_snapshot[18].r.part0[12] , 
	\sa_snapshot[18].r.part0[11] , \sa_snapshot[18].r.part0[10] , 
	\sa_snapshot[18].r.part0[9] , \sa_snapshot[18].r.part0[8] , 
	\sa_snapshot[18].r.part0[7] , \sa_snapshot[18].r.part0[6] , 
	\sa_snapshot[18].r.part0[5] , \sa_snapshot[18].r.part0[4] , 
	\sa_snapshot[18].r.part0[3] , \sa_snapshot[18].r.part0[2] , 
	\sa_snapshot[18].r.part0[1] , \sa_snapshot[18].r.part0[0] , 
	\sa_snapshot[17].r.part1[31] , \sa_snapshot[17].r.part1[30] , 
	\sa_snapshot[17].r.part1[29] , \sa_snapshot[17].r.part1[28] , 
	\sa_snapshot[17].r.part1[27] , \sa_snapshot[17].r.part1[26] , 
	\sa_snapshot[17].r.part1[25] , \sa_snapshot[17].r.part1[24] , 
	\sa_snapshot[17].r.part1[23] , \sa_snapshot[17].r.part1[22] , 
	\sa_snapshot[17].r.part1[21] , \sa_snapshot[17].r.part1[20] , 
	\sa_snapshot[17].r.part1[19] , \sa_snapshot[17].r.part1[18] , 
	\sa_snapshot[17].r.part1[17] , \sa_snapshot[17].r.part1[16] , 
	\sa_snapshot[17].r.part1[15] , \sa_snapshot[17].r.part1[14] , 
	\sa_snapshot[17].r.part1[13] , \sa_snapshot[17].r.part1[12] , 
	\sa_snapshot[17].r.part1[11] , \sa_snapshot[17].r.part1[10] , 
	\sa_snapshot[17].r.part1[9] , \sa_snapshot[17].r.part1[8] , 
	\sa_snapshot[17].r.part1[7] , \sa_snapshot[17].r.part1[6] , 
	\sa_snapshot[17].r.part1[5] , \sa_snapshot[17].r.part1[4] , 
	\sa_snapshot[17].r.part1[3] , \sa_snapshot[17].r.part1[2] , 
	\sa_snapshot[17].r.part1[1] , \sa_snapshot[17].r.part1[0] , 
	\sa_snapshot[17].r.part0[31] , \sa_snapshot[17].r.part0[30] , 
	\sa_snapshot[17].r.part0[29] , \sa_snapshot[17].r.part0[28] , 
	\sa_snapshot[17].r.part0[27] , \sa_snapshot[17].r.part0[26] , 
	\sa_snapshot[17].r.part0[25] , \sa_snapshot[17].r.part0[24] , 
	\sa_snapshot[17].r.part0[23] , \sa_snapshot[17].r.part0[22] , 
	\sa_snapshot[17].r.part0[21] , \sa_snapshot[17].r.part0[20] , 
	\sa_snapshot[17].r.part0[19] , \sa_snapshot[17].r.part0[18] , 
	\sa_snapshot[17].r.part0[17] , \sa_snapshot[17].r.part0[16] , 
	\sa_snapshot[17].r.part0[15] , \sa_snapshot[17].r.part0[14] , 
	\sa_snapshot[17].r.part0[13] , \sa_snapshot[17].r.part0[12] , 
	\sa_snapshot[17].r.part0[11] , \sa_snapshot[17].r.part0[10] , 
	\sa_snapshot[17].r.part0[9] , \sa_snapshot[17].r.part0[8] , 
	\sa_snapshot[17].r.part0[7] , \sa_snapshot[17].r.part0[6] , 
	\sa_snapshot[17].r.part0[5] , \sa_snapshot[17].r.part0[4] , 
	\sa_snapshot[17].r.part0[3] , \sa_snapshot[17].r.part0[2] , 
	\sa_snapshot[17].r.part0[1] , \sa_snapshot[17].r.part0[0] , 
	\sa_snapshot[16].r.part1[31] , \sa_snapshot[16].r.part1[30] , 
	\sa_snapshot[16].r.part1[29] , \sa_snapshot[16].r.part1[28] , 
	\sa_snapshot[16].r.part1[27] , \sa_snapshot[16].r.part1[26] , 
	\sa_snapshot[16].r.part1[25] , \sa_snapshot[16].r.part1[24] , 
	\sa_snapshot[16].r.part1[23] , \sa_snapshot[16].r.part1[22] , 
	\sa_snapshot[16].r.part1[21] , \sa_snapshot[16].r.part1[20] , 
	\sa_snapshot[16].r.part1[19] , \sa_snapshot[16].r.part1[18] , 
	\sa_snapshot[16].r.part1[17] , \sa_snapshot[16].r.part1[16] , 
	\sa_snapshot[16].r.part1[15] , \sa_snapshot[16].r.part1[14] , 
	\sa_snapshot[16].r.part1[13] , \sa_snapshot[16].r.part1[12] , 
	\sa_snapshot[16].r.part1[11] , \sa_snapshot[16].r.part1[10] , 
	\sa_snapshot[16].r.part1[9] , \sa_snapshot[16].r.part1[8] , 
	\sa_snapshot[16].r.part1[7] , \sa_snapshot[16].r.part1[6] , 
	\sa_snapshot[16].r.part1[5] , \sa_snapshot[16].r.part1[4] , 
	\sa_snapshot[16].r.part1[3] , \sa_snapshot[16].r.part1[2] , 
	\sa_snapshot[16].r.part1[1] , \sa_snapshot[16].r.part1[0] , 
	\sa_snapshot[16].r.part0[31] , \sa_snapshot[16].r.part0[30] , 
	\sa_snapshot[16].r.part0[29] , \sa_snapshot[16].r.part0[28] , 
	\sa_snapshot[16].r.part0[27] , \sa_snapshot[16].r.part0[26] , 
	\sa_snapshot[16].r.part0[25] , \sa_snapshot[16].r.part0[24] , 
	\sa_snapshot[16].r.part0[23] , \sa_snapshot[16].r.part0[22] , 
	\sa_snapshot[16].r.part0[21] , \sa_snapshot[16].r.part0[20] , 
	\sa_snapshot[16].r.part0[19] , \sa_snapshot[16].r.part0[18] , 
	\sa_snapshot[16].r.part0[17] , \sa_snapshot[16].r.part0[16] , 
	\sa_snapshot[16].r.part0[15] , \sa_snapshot[16].r.part0[14] , 
	\sa_snapshot[16].r.part0[13] , \sa_snapshot[16].r.part0[12] , 
	\sa_snapshot[16].r.part0[11] , \sa_snapshot[16].r.part0[10] , 
	\sa_snapshot[16].r.part0[9] , \sa_snapshot[16].r.part0[8] , 
	\sa_snapshot[16].r.part0[7] , \sa_snapshot[16].r.part0[6] , 
	\sa_snapshot[16].r.part0[5] , \sa_snapshot[16].r.part0[4] , 
	\sa_snapshot[16].r.part0[3] , \sa_snapshot[16].r.part0[2] , 
	\sa_snapshot[16].r.part0[1] , \sa_snapshot[16].r.part0[0] , 
	\sa_snapshot[15].r.part1[31] , \sa_snapshot[15].r.part1[30] , 
	\sa_snapshot[15].r.part1[29] , \sa_snapshot[15].r.part1[28] , 
	\sa_snapshot[15].r.part1[27] , \sa_snapshot[15].r.part1[26] , 
	\sa_snapshot[15].r.part1[25] , \sa_snapshot[15].r.part1[24] , 
	\sa_snapshot[15].r.part1[23] , \sa_snapshot[15].r.part1[22] , 
	\sa_snapshot[15].r.part1[21] , \sa_snapshot[15].r.part1[20] , 
	\sa_snapshot[15].r.part1[19] , \sa_snapshot[15].r.part1[18] , 
	\sa_snapshot[15].r.part1[17] , \sa_snapshot[15].r.part1[16] , 
	\sa_snapshot[15].r.part1[15] , \sa_snapshot[15].r.part1[14] , 
	\sa_snapshot[15].r.part1[13] , \sa_snapshot[15].r.part1[12] , 
	\sa_snapshot[15].r.part1[11] , \sa_snapshot[15].r.part1[10] , 
	\sa_snapshot[15].r.part1[9] , \sa_snapshot[15].r.part1[8] , 
	\sa_snapshot[15].r.part1[7] , \sa_snapshot[15].r.part1[6] , 
	\sa_snapshot[15].r.part1[5] , \sa_snapshot[15].r.part1[4] , 
	\sa_snapshot[15].r.part1[3] , \sa_snapshot[15].r.part1[2] , 
	\sa_snapshot[15].r.part1[1] , \sa_snapshot[15].r.part1[0] , 
	\sa_snapshot[15].r.part0[31] , \sa_snapshot[15].r.part0[30] , 
	\sa_snapshot[15].r.part0[29] , \sa_snapshot[15].r.part0[28] , 
	\sa_snapshot[15].r.part0[27] , \sa_snapshot[15].r.part0[26] , 
	\sa_snapshot[15].r.part0[25] , \sa_snapshot[15].r.part0[24] , 
	\sa_snapshot[15].r.part0[23] , \sa_snapshot[15].r.part0[22] , 
	\sa_snapshot[15].r.part0[21] , \sa_snapshot[15].r.part0[20] , 
	\sa_snapshot[15].r.part0[19] , \sa_snapshot[15].r.part0[18] , 
	\sa_snapshot[15].r.part0[17] , \sa_snapshot[15].r.part0[16] , 
	\sa_snapshot[15].r.part0[15] , \sa_snapshot[15].r.part0[14] , 
	\sa_snapshot[15].r.part0[13] , \sa_snapshot[15].r.part0[12] , 
	\sa_snapshot[15].r.part0[11] , \sa_snapshot[15].r.part0[10] , 
	\sa_snapshot[15].r.part0[9] , \sa_snapshot[15].r.part0[8] , 
	\sa_snapshot[15].r.part0[7] , \sa_snapshot[15].r.part0[6] , 
	\sa_snapshot[15].r.part0[5] , \sa_snapshot[15].r.part0[4] , 
	\sa_snapshot[15].r.part0[3] , \sa_snapshot[15].r.part0[2] , 
	\sa_snapshot[15].r.part0[1] , \sa_snapshot[15].r.part0[0] , 
	\sa_snapshot[14].r.part1[31] , \sa_snapshot[14].r.part1[30] , 
	\sa_snapshot[14].r.part1[29] , \sa_snapshot[14].r.part1[28] , 
	\sa_snapshot[14].r.part1[27] , \sa_snapshot[14].r.part1[26] , 
	\sa_snapshot[14].r.part1[25] , \sa_snapshot[14].r.part1[24] , 
	\sa_snapshot[14].r.part1[23] , \sa_snapshot[14].r.part1[22] , 
	\sa_snapshot[14].r.part1[21] , \sa_snapshot[14].r.part1[20] , 
	\sa_snapshot[14].r.part1[19] , \sa_snapshot[14].r.part1[18] , 
	\sa_snapshot[14].r.part1[17] , \sa_snapshot[14].r.part1[16] , 
	\sa_snapshot[14].r.part1[15] , \sa_snapshot[14].r.part1[14] , 
	\sa_snapshot[14].r.part1[13] , \sa_snapshot[14].r.part1[12] , 
	\sa_snapshot[14].r.part1[11] , \sa_snapshot[14].r.part1[10] , 
	\sa_snapshot[14].r.part1[9] , \sa_snapshot[14].r.part1[8] , 
	\sa_snapshot[14].r.part1[7] , \sa_snapshot[14].r.part1[6] , 
	\sa_snapshot[14].r.part1[5] , \sa_snapshot[14].r.part1[4] , 
	\sa_snapshot[14].r.part1[3] , \sa_snapshot[14].r.part1[2] , 
	\sa_snapshot[14].r.part1[1] , \sa_snapshot[14].r.part1[0] , 
	\sa_snapshot[14].r.part0[31] , \sa_snapshot[14].r.part0[30] , 
	\sa_snapshot[14].r.part0[29] , \sa_snapshot[14].r.part0[28] , 
	\sa_snapshot[14].r.part0[27] , \sa_snapshot[14].r.part0[26] , 
	\sa_snapshot[14].r.part0[25] , \sa_snapshot[14].r.part0[24] , 
	\sa_snapshot[14].r.part0[23] , \sa_snapshot[14].r.part0[22] , 
	\sa_snapshot[14].r.part0[21] , \sa_snapshot[14].r.part0[20] , 
	\sa_snapshot[14].r.part0[19] , \sa_snapshot[14].r.part0[18] , 
	\sa_snapshot[14].r.part0[17] , \sa_snapshot[14].r.part0[16] , 
	\sa_snapshot[14].r.part0[15] , \sa_snapshot[14].r.part0[14] , 
	\sa_snapshot[14].r.part0[13] , \sa_snapshot[14].r.part0[12] , 
	\sa_snapshot[14].r.part0[11] , \sa_snapshot[14].r.part0[10] , 
	\sa_snapshot[14].r.part0[9] , \sa_snapshot[14].r.part0[8] , 
	\sa_snapshot[14].r.part0[7] , \sa_snapshot[14].r.part0[6] , 
	\sa_snapshot[14].r.part0[5] , \sa_snapshot[14].r.part0[4] , 
	\sa_snapshot[14].r.part0[3] , \sa_snapshot[14].r.part0[2] , 
	\sa_snapshot[14].r.part0[1] , \sa_snapshot[14].r.part0[0] , 
	\sa_snapshot[13].r.part1[31] , \sa_snapshot[13].r.part1[30] , 
	\sa_snapshot[13].r.part1[29] , \sa_snapshot[13].r.part1[28] , 
	\sa_snapshot[13].r.part1[27] , \sa_snapshot[13].r.part1[26] , 
	\sa_snapshot[13].r.part1[25] , \sa_snapshot[13].r.part1[24] , 
	\sa_snapshot[13].r.part1[23] , \sa_snapshot[13].r.part1[22] , 
	\sa_snapshot[13].r.part1[21] , \sa_snapshot[13].r.part1[20] , 
	\sa_snapshot[13].r.part1[19] , \sa_snapshot[13].r.part1[18] , 
	\sa_snapshot[13].r.part1[17] , \sa_snapshot[13].r.part1[16] , 
	\sa_snapshot[13].r.part1[15] , \sa_snapshot[13].r.part1[14] , 
	\sa_snapshot[13].r.part1[13] , \sa_snapshot[13].r.part1[12] , 
	\sa_snapshot[13].r.part1[11] , \sa_snapshot[13].r.part1[10] , 
	\sa_snapshot[13].r.part1[9] , \sa_snapshot[13].r.part1[8] , 
	\sa_snapshot[13].r.part1[7] , \sa_snapshot[13].r.part1[6] , 
	\sa_snapshot[13].r.part1[5] , \sa_snapshot[13].r.part1[4] , 
	\sa_snapshot[13].r.part1[3] , \sa_snapshot[13].r.part1[2] , 
	\sa_snapshot[13].r.part1[1] , \sa_snapshot[13].r.part1[0] , 
	\sa_snapshot[13].r.part0[31] , \sa_snapshot[13].r.part0[30] , 
	\sa_snapshot[13].r.part0[29] , \sa_snapshot[13].r.part0[28] , 
	\sa_snapshot[13].r.part0[27] , \sa_snapshot[13].r.part0[26] , 
	\sa_snapshot[13].r.part0[25] , \sa_snapshot[13].r.part0[24] , 
	\sa_snapshot[13].r.part0[23] , \sa_snapshot[13].r.part0[22] , 
	\sa_snapshot[13].r.part0[21] , \sa_snapshot[13].r.part0[20] , 
	\sa_snapshot[13].r.part0[19] , \sa_snapshot[13].r.part0[18] , 
	\sa_snapshot[13].r.part0[17] , \sa_snapshot[13].r.part0[16] , 
	\sa_snapshot[13].r.part0[15] , \sa_snapshot[13].r.part0[14] , 
	\sa_snapshot[13].r.part0[13] , \sa_snapshot[13].r.part0[12] , 
	\sa_snapshot[13].r.part0[11] , \sa_snapshot[13].r.part0[10] , 
	\sa_snapshot[13].r.part0[9] , \sa_snapshot[13].r.part0[8] , 
	\sa_snapshot[13].r.part0[7] , \sa_snapshot[13].r.part0[6] , 
	\sa_snapshot[13].r.part0[5] , \sa_snapshot[13].r.part0[4] , 
	\sa_snapshot[13].r.part0[3] , \sa_snapshot[13].r.part0[2] , 
	\sa_snapshot[13].r.part0[1] , \sa_snapshot[13].r.part0[0] , 
	\sa_snapshot[12].r.part1[31] , \sa_snapshot[12].r.part1[30] , 
	\sa_snapshot[12].r.part1[29] , \sa_snapshot[12].r.part1[28] , 
	\sa_snapshot[12].r.part1[27] , \sa_snapshot[12].r.part1[26] , 
	\sa_snapshot[12].r.part1[25] , \sa_snapshot[12].r.part1[24] , 
	\sa_snapshot[12].r.part1[23] , \sa_snapshot[12].r.part1[22] , 
	\sa_snapshot[12].r.part1[21] , \sa_snapshot[12].r.part1[20] , 
	\sa_snapshot[12].r.part1[19] , \sa_snapshot[12].r.part1[18] , 
	\sa_snapshot[12].r.part1[17] , \sa_snapshot[12].r.part1[16] , 
	\sa_snapshot[12].r.part1[15] , \sa_snapshot[12].r.part1[14] , 
	\sa_snapshot[12].r.part1[13] , \sa_snapshot[12].r.part1[12] , 
	\sa_snapshot[12].r.part1[11] , \sa_snapshot[12].r.part1[10] , 
	\sa_snapshot[12].r.part1[9] , \sa_snapshot[12].r.part1[8] , 
	\sa_snapshot[12].r.part1[7] , \sa_snapshot[12].r.part1[6] , 
	\sa_snapshot[12].r.part1[5] , \sa_snapshot[12].r.part1[4] , 
	\sa_snapshot[12].r.part1[3] , \sa_snapshot[12].r.part1[2] , 
	\sa_snapshot[12].r.part1[1] , \sa_snapshot[12].r.part1[0] , 
	\sa_snapshot[12].r.part0[31] , \sa_snapshot[12].r.part0[30] , 
	\sa_snapshot[12].r.part0[29] , \sa_snapshot[12].r.part0[28] , 
	\sa_snapshot[12].r.part0[27] , \sa_snapshot[12].r.part0[26] , 
	\sa_snapshot[12].r.part0[25] , \sa_snapshot[12].r.part0[24] , 
	\sa_snapshot[12].r.part0[23] , \sa_snapshot[12].r.part0[22] , 
	\sa_snapshot[12].r.part0[21] , \sa_snapshot[12].r.part0[20] , 
	\sa_snapshot[12].r.part0[19] , \sa_snapshot[12].r.part0[18] , 
	\sa_snapshot[12].r.part0[17] , \sa_snapshot[12].r.part0[16] , 
	\sa_snapshot[12].r.part0[15] , \sa_snapshot[12].r.part0[14] , 
	\sa_snapshot[12].r.part0[13] , \sa_snapshot[12].r.part0[12] , 
	\sa_snapshot[12].r.part0[11] , \sa_snapshot[12].r.part0[10] , 
	\sa_snapshot[12].r.part0[9] , \sa_snapshot[12].r.part0[8] , 
	\sa_snapshot[12].r.part0[7] , \sa_snapshot[12].r.part0[6] , 
	\sa_snapshot[12].r.part0[5] , \sa_snapshot[12].r.part0[4] , 
	\sa_snapshot[12].r.part0[3] , \sa_snapshot[12].r.part0[2] , 
	\sa_snapshot[12].r.part0[1] , \sa_snapshot[12].r.part0[0] , 
	\sa_snapshot[11].r.part1[31] , \sa_snapshot[11].r.part1[30] , 
	\sa_snapshot[11].r.part1[29] , \sa_snapshot[11].r.part1[28] , 
	\sa_snapshot[11].r.part1[27] , \sa_snapshot[11].r.part1[26] , 
	\sa_snapshot[11].r.part1[25] , \sa_snapshot[11].r.part1[24] , 
	\sa_snapshot[11].r.part1[23] , \sa_snapshot[11].r.part1[22] , 
	\sa_snapshot[11].r.part1[21] , \sa_snapshot[11].r.part1[20] , 
	\sa_snapshot[11].r.part1[19] , \sa_snapshot[11].r.part1[18] , 
	\sa_snapshot[11].r.part1[17] , \sa_snapshot[11].r.part1[16] , 
	\sa_snapshot[11].r.part1[15] , \sa_snapshot[11].r.part1[14] , 
	\sa_snapshot[11].r.part1[13] , \sa_snapshot[11].r.part1[12] , 
	\sa_snapshot[11].r.part1[11] , \sa_snapshot[11].r.part1[10] , 
	\sa_snapshot[11].r.part1[9] , \sa_snapshot[11].r.part1[8] , 
	\sa_snapshot[11].r.part1[7] , \sa_snapshot[11].r.part1[6] , 
	\sa_snapshot[11].r.part1[5] , \sa_snapshot[11].r.part1[4] , 
	\sa_snapshot[11].r.part1[3] , \sa_snapshot[11].r.part1[2] , 
	\sa_snapshot[11].r.part1[1] , \sa_snapshot[11].r.part1[0] , 
	\sa_snapshot[11].r.part0[31] , \sa_snapshot[11].r.part0[30] , 
	\sa_snapshot[11].r.part0[29] , \sa_snapshot[11].r.part0[28] , 
	\sa_snapshot[11].r.part0[27] , \sa_snapshot[11].r.part0[26] , 
	\sa_snapshot[11].r.part0[25] , \sa_snapshot[11].r.part0[24] , 
	\sa_snapshot[11].r.part0[23] , \sa_snapshot[11].r.part0[22] , 
	\sa_snapshot[11].r.part0[21] , \sa_snapshot[11].r.part0[20] , 
	\sa_snapshot[11].r.part0[19] , \sa_snapshot[11].r.part0[18] , 
	\sa_snapshot[11].r.part0[17] , \sa_snapshot[11].r.part0[16] , 
	\sa_snapshot[11].r.part0[15] , \sa_snapshot[11].r.part0[14] , 
	\sa_snapshot[11].r.part0[13] , \sa_snapshot[11].r.part0[12] , 
	\sa_snapshot[11].r.part0[11] , \sa_snapshot[11].r.part0[10] , 
	\sa_snapshot[11].r.part0[9] , \sa_snapshot[11].r.part0[8] , 
	\sa_snapshot[11].r.part0[7] , \sa_snapshot[11].r.part0[6] , 
	\sa_snapshot[11].r.part0[5] , \sa_snapshot[11].r.part0[4] , 
	\sa_snapshot[11].r.part0[3] , \sa_snapshot[11].r.part0[2] , 
	\sa_snapshot[11].r.part0[1] , \sa_snapshot[11].r.part0[0] , 
	\sa_snapshot[10].r.part1[31] , \sa_snapshot[10].r.part1[30] , 
	\sa_snapshot[10].r.part1[29] , \sa_snapshot[10].r.part1[28] , 
	\sa_snapshot[10].r.part1[27] , \sa_snapshot[10].r.part1[26] , 
	\sa_snapshot[10].r.part1[25] , \sa_snapshot[10].r.part1[24] , 
	\sa_snapshot[10].r.part1[23] , \sa_snapshot[10].r.part1[22] , 
	\sa_snapshot[10].r.part1[21] , \sa_snapshot[10].r.part1[20] , 
	\sa_snapshot[10].r.part1[19] , \sa_snapshot[10].r.part1[18] , 
	\sa_snapshot[10].r.part1[17] , \sa_snapshot[10].r.part1[16] , 
	\sa_snapshot[10].r.part1[15] , \sa_snapshot[10].r.part1[14] , 
	\sa_snapshot[10].r.part1[13] , \sa_snapshot[10].r.part1[12] , 
	\sa_snapshot[10].r.part1[11] , \sa_snapshot[10].r.part1[10] , 
	\sa_snapshot[10].r.part1[9] , \sa_snapshot[10].r.part1[8] , 
	\sa_snapshot[10].r.part1[7] , \sa_snapshot[10].r.part1[6] , 
	\sa_snapshot[10].r.part1[5] , \sa_snapshot[10].r.part1[4] , 
	\sa_snapshot[10].r.part1[3] , \sa_snapshot[10].r.part1[2] , 
	\sa_snapshot[10].r.part1[1] , \sa_snapshot[10].r.part1[0] , 
	\sa_snapshot[10].r.part0[31] , \sa_snapshot[10].r.part0[30] , 
	\sa_snapshot[10].r.part0[29] , \sa_snapshot[10].r.part0[28] , 
	\sa_snapshot[10].r.part0[27] , \sa_snapshot[10].r.part0[26] , 
	\sa_snapshot[10].r.part0[25] , \sa_snapshot[10].r.part0[24] , 
	\sa_snapshot[10].r.part0[23] , \sa_snapshot[10].r.part0[22] , 
	\sa_snapshot[10].r.part0[21] , \sa_snapshot[10].r.part0[20] , 
	\sa_snapshot[10].r.part0[19] , \sa_snapshot[10].r.part0[18] , 
	\sa_snapshot[10].r.part0[17] , \sa_snapshot[10].r.part0[16] , 
	\sa_snapshot[10].r.part0[15] , \sa_snapshot[10].r.part0[14] , 
	\sa_snapshot[10].r.part0[13] , \sa_snapshot[10].r.part0[12] , 
	\sa_snapshot[10].r.part0[11] , \sa_snapshot[10].r.part0[10] , 
	\sa_snapshot[10].r.part0[9] , \sa_snapshot[10].r.part0[8] , 
	\sa_snapshot[10].r.part0[7] , \sa_snapshot[10].r.part0[6] , 
	\sa_snapshot[10].r.part0[5] , \sa_snapshot[10].r.part0[4] , 
	\sa_snapshot[10].r.part0[3] , \sa_snapshot[10].r.part0[2] , 
	\sa_snapshot[10].r.part0[1] , \sa_snapshot[10].r.part0[0] , 
	\sa_snapshot[9].r.part1[31] , \sa_snapshot[9].r.part1[30] , 
	\sa_snapshot[9].r.part1[29] , \sa_snapshot[9].r.part1[28] , 
	\sa_snapshot[9].r.part1[27] , \sa_snapshot[9].r.part1[26] , 
	\sa_snapshot[9].r.part1[25] , \sa_snapshot[9].r.part1[24] , 
	\sa_snapshot[9].r.part1[23] , \sa_snapshot[9].r.part1[22] , 
	\sa_snapshot[9].r.part1[21] , \sa_snapshot[9].r.part1[20] , 
	\sa_snapshot[9].r.part1[19] , \sa_snapshot[9].r.part1[18] , 
	\sa_snapshot[9].r.part1[17] , \sa_snapshot[9].r.part1[16] , 
	\sa_snapshot[9].r.part1[15] , \sa_snapshot[9].r.part1[14] , 
	\sa_snapshot[9].r.part1[13] , \sa_snapshot[9].r.part1[12] , 
	\sa_snapshot[9].r.part1[11] , \sa_snapshot[9].r.part1[10] , 
	\sa_snapshot[9].r.part1[9] , \sa_snapshot[9].r.part1[8] , 
	\sa_snapshot[9].r.part1[7] , \sa_snapshot[9].r.part1[6] , 
	\sa_snapshot[9].r.part1[5] , \sa_snapshot[9].r.part1[4] , 
	\sa_snapshot[9].r.part1[3] , \sa_snapshot[9].r.part1[2] , 
	\sa_snapshot[9].r.part1[1] , \sa_snapshot[9].r.part1[0] , 
	\sa_snapshot[9].r.part0[31] , \sa_snapshot[9].r.part0[30] , 
	\sa_snapshot[9].r.part0[29] , \sa_snapshot[9].r.part0[28] , 
	\sa_snapshot[9].r.part0[27] , \sa_snapshot[9].r.part0[26] , 
	\sa_snapshot[9].r.part0[25] , \sa_snapshot[9].r.part0[24] , 
	\sa_snapshot[9].r.part0[23] , \sa_snapshot[9].r.part0[22] , 
	\sa_snapshot[9].r.part0[21] , \sa_snapshot[9].r.part0[20] , 
	\sa_snapshot[9].r.part0[19] , \sa_snapshot[9].r.part0[18] , 
	\sa_snapshot[9].r.part0[17] , \sa_snapshot[9].r.part0[16] , 
	\sa_snapshot[9].r.part0[15] , \sa_snapshot[9].r.part0[14] , 
	\sa_snapshot[9].r.part0[13] , \sa_snapshot[9].r.part0[12] , 
	\sa_snapshot[9].r.part0[11] , \sa_snapshot[9].r.part0[10] , 
	\sa_snapshot[9].r.part0[9] , \sa_snapshot[9].r.part0[8] , 
	\sa_snapshot[9].r.part0[7] , \sa_snapshot[9].r.part0[6] , 
	\sa_snapshot[9].r.part0[5] , \sa_snapshot[9].r.part0[4] , 
	\sa_snapshot[9].r.part0[3] , \sa_snapshot[9].r.part0[2] , 
	\sa_snapshot[9].r.part0[1] , \sa_snapshot[9].r.part0[0] , 
	\sa_snapshot[8].r.part1[31] , \sa_snapshot[8].r.part1[30] , 
	\sa_snapshot[8].r.part1[29] , \sa_snapshot[8].r.part1[28] , 
	\sa_snapshot[8].r.part1[27] , \sa_snapshot[8].r.part1[26] , 
	\sa_snapshot[8].r.part1[25] , \sa_snapshot[8].r.part1[24] , 
	\sa_snapshot[8].r.part1[23] , \sa_snapshot[8].r.part1[22] , 
	\sa_snapshot[8].r.part1[21] , \sa_snapshot[8].r.part1[20] , 
	\sa_snapshot[8].r.part1[19] , \sa_snapshot[8].r.part1[18] , 
	\sa_snapshot[8].r.part1[17] , \sa_snapshot[8].r.part1[16] , 
	\sa_snapshot[8].r.part1[15] , \sa_snapshot[8].r.part1[14] , 
	\sa_snapshot[8].r.part1[13] , \sa_snapshot[8].r.part1[12] , 
	\sa_snapshot[8].r.part1[11] , \sa_snapshot[8].r.part1[10] , 
	\sa_snapshot[8].r.part1[9] , \sa_snapshot[8].r.part1[8] , 
	\sa_snapshot[8].r.part1[7] , \sa_snapshot[8].r.part1[6] , 
	\sa_snapshot[8].r.part1[5] , \sa_snapshot[8].r.part1[4] , 
	\sa_snapshot[8].r.part1[3] , \sa_snapshot[8].r.part1[2] , 
	\sa_snapshot[8].r.part1[1] , \sa_snapshot[8].r.part1[0] , 
	\sa_snapshot[8].r.part0[31] , \sa_snapshot[8].r.part0[30] , 
	\sa_snapshot[8].r.part0[29] , \sa_snapshot[8].r.part0[28] , 
	\sa_snapshot[8].r.part0[27] , \sa_snapshot[8].r.part0[26] , 
	\sa_snapshot[8].r.part0[25] , \sa_snapshot[8].r.part0[24] , 
	\sa_snapshot[8].r.part0[23] , \sa_snapshot[8].r.part0[22] , 
	\sa_snapshot[8].r.part0[21] , \sa_snapshot[8].r.part0[20] , 
	\sa_snapshot[8].r.part0[19] , \sa_snapshot[8].r.part0[18] , 
	\sa_snapshot[8].r.part0[17] , \sa_snapshot[8].r.part0[16] , 
	\sa_snapshot[8].r.part0[15] , \sa_snapshot[8].r.part0[14] , 
	\sa_snapshot[8].r.part0[13] , \sa_snapshot[8].r.part0[12] , 
	\sa_snapshot[8].r.part0[11] , \sa_snapshot[8].r.part0[10] , 
	\sa_snapshot[8].r.part0[9] , \sa_snapshot[8].r.part0[8] , 
	\sa_snapshot[8].r.part0[7] , \sa_snapshot[8].r.part0[6] , 
	\sa_snapshot[8].r.part0[5] , \sa_snapshot[8].r.part0[4] , 
	\sa_snapshot[8].r.part0[3] , \sa_snapshot[8].r.part0[2] , 
	\sa_snapshot[8].r.part0[1] , \sa_snapshot[8].r.part0[0] , 
	\sa_snapshot[7].r.part1[31] , \sa_snapshot[7].r.part1[30] , 
	\sa_snapshot[7].r.part1[29] , \sa_snapshot[7].r.part1[28] , 
	\sa_snapshot[7].r.part1[27] , \sa_snapshot[7].r.part1[26] , 
	\sa_snapshot[7].r.part1[25] , \sa_snapshot[7].r.part1[24] , 
	\sa_snapshot[7].r.part1[23] , \sa_snapshot[7].r.part1[22] , 
	\sa_snapshot[7].r.part1[21] , \sa_snapshot[7].r.part1[20] , 
	\sa_snapshot[7].r.part1[19] , \sa_snapshot[7].r.part1[18] , 
	\sa_snapshot[7].r.part1[17] , \sa_snapshot[7].r.part1[16] , 
	\sa_snapshot[7].r.part1[15] , \sa_snapshot[7].r.part1[14] , 
	\sa_snapshot[7].r.part1[13] , \sa_snapshot[7].r.part1[12] , 
	\sa_snapshot[7].r.part1[11] , \sa_snapshot[7].r.part1[10] , 
	\sa_snapshot[7].r.part1[9] , \sa_snapshot[7].r.part1[8] , 
	\sa_snapshot[7].r.part1[7] , \sa_snapshot[7].r.part1[6] , 
	\sa_snapshot[7].r.part1[5] , \sa_snapshot[7].r.part1[4] , 
	\sa_snapshot[7].r.part1[3] , \sa_snapshot[7].r.part1[2] , 
	\sa_snapshot[7].r.part1[1] , \sa_snapshot[7].r.part1[0] , 
	\sa_snapshot[7].r.part0[31] , \sa_snapshot[7].r.part0[30] , 
	\sa_snapshot[7].r.part0[29] , \sa_snapshot[7].r.part0[28] , 
	\sa_snapshot[7].r.part0[27] , \sa_snapshot[7].r.part0[26] , 
	\sa_snapshot[7].r.part0[25] , \sa_snapshot[7].r.part0[24] , 
	\sa_snapshot[7].r.part0[23] , \sa_snapshot[7].r.part0[22] , 
	\sa_snapshot[7].r.part0[21] , \sa_snapshot[7].r.part0[20] , 
	\sa_snapshot[7].r.part0[19] , \sa_snapshot[7].r.part0[18] , 
	\sa_snapshot[7].r.part0[17] , \sa_snapshot[7].r.part0[16] , 
	\sa_snapshot[7].r.part0[15] , \sa_snapshot[7].r.part0[14] , 
	\sa_snapshot[7].r.part0[13] , \sa_snapshot[7].r.part0[12] , 
	\sa_snapshot[7].r.part0[11] , \sa_snapshot[7].r.part0[10] , 
	\sa_snapshot[7].r.part0[9] , \sa_snapshot[7].r.part0[8] , 
	\sa_snapshot[7].r.part0[7] , \sa_snapshot[7].r.part0[6] , 
	\sa_snapshot[7].r.part0[5] , \sa_snapshot[7].r.part0[4] , 
	\sa_snapshot[7].r.part0[3] , \sa_snapshot[7].r.part0[2] , 
	\sa_snapshot[7].r.part0[1] , \sa_snapshot[7].r.part0[0] , 
	\sa_snapshot[6].r.part1[31] , \sa_snapshot[6].r.part1[30] , 
	\sa_snapshot[6].r.part1[29] , \sa_snapshot[6].r.part1[28] , 
	\sa_snapshot[6].r.part1[27] , \sa_snapshot[6].r.part1[26] , 
	\sa_snapshot[6].r.part1[25] , \sa_snapshot[6].r.part1[24] , 
	\sa_snapshot[6].r.part1[23] , \sa_snapshot[6].r.part1[22] , 
	\sa_snapshot[6].r.part1[21] , \sa_snapshot[6].r.part1[20] , 
	\sa_snapshot[6].r.part1[19] , \sa_snapshot[6].r.part1[18] , 
	\sa_snapshot[6].r.part1[17] , \sa_snapshot[6].r.part1[16] , 
	\sa_snapshot[6].r.part1[15] , \sa_snapshot[6].r.part1[14] , 
	\sa_snapshot[6].r.part1[13] , \sa_snapshot[6].r.part1[12] , 
	\sa_snapshot[6].r.part1[11] , \sa_snapshot[6].r.part1[10] , 
	\sa_snapshot[6].r.part1[9] , \sa_snapshot[6].r.part1[8] , 
	\sa_snapshot[6].r.part1[7] , \sa_snapshot[6].r.part1[6] , 
	\sa_snapshot[6].r.part1[5] , \sa_snapshot[6].r.part1[4] , 
	\sa_snapshot[6].r.part1[3] , \sa_snapshot[6].r.part1[2] , 
	\sa_snapshot[6].r.part1[1] , \sa_snapshot[6].r.part1[0] , 
	\sa_snapshot[6].r.part0[31] , \sa_snapshot[6].r.part0[30] , 
	\sa_snapshot[6].r.part0[29] , \sa_snapshot[6].r.part0[28] , 
	\sa_snapshot[6].r.part0[27] , \sa_snapshot[6].r.part0[26] , 
	\sa_snapshot[6].r.part0[25] , \sa_snapshot[6].r.part0[24] , 
	\sa_snapshot[6].r.part0[23] , \sa_snapshot[6].r.part0[22] , 
	\sa_snapshot[6].r.part0[21] , \sa_snapshot[6].r.part0[20] , 
	\sa_snapshot[6].r.part0[19] , \sa_snapshot[6].r.part0[18] , 
	\sa_snapshot[6].r.part0[17] , \sa_snapshot[6].r.part0[16] , 
	\sa_snapshot[6].r.part0[15] , \sa_snapshot[6].r.part0[14] , 
	\sa_snapshot[6].r.part0[13] , \sa_snapshot[6].r.part0[12] , 
	\sa_snapshot[6].r.part0[11] , \sa_snapshot[6].r.part0[10] , 
	\sa_snapshot[6].r.part0[9] , \sa_snapshot[6].r.part0[8] , 
	\sa_snapshot[6].r.part0[7] , \sa_snapshot[6].r.part0[6] , 
	\sa_snapshot[6].r.part0[5] , \sa_snapshot[6].r.part0[4] , 
	\sa_snapshot[6].r.part0[3] , \sa_snapshot[6].r.part0[2] , 
	\sa_snapshot[6].r.part0[1] , \sa_snapshot[6].r.part0[0] , 
	\sa_snapshot[5].r.part1[31] , \sa_snapshot[5].r.part1[30] , 
	\sa_snapshot[5].r.part1[29] , \sa_snapshot[5].r.part1[28] , 
	\sa_snapshot[5].r.part1[27] , \sa_snapshot[5].r.part1[26] , 
	\sa_snapshot[5].r.part1[25] , \sa_snapshot[5].r.part1[24] , 
	\sa_snapshot[5].r.part1[23] , \sa_snapshot[5].r.part1[22] , 
	\sa_snapshot[5].r.part1[21] , \sa_snapshot[5].r.part1[20] , 
	\sa_snapshot[5].r.part1[19] , \sa_snapshot[5].r.part1[18] , 
	\sa_snapshot[5].r.part1[17] , \sa_snapshot[5].r.part1[16] , 
	\sa_snapshot[5].r.part1[15] , \sa_snapshot[5].r.part1[14] , 
	\sa_snapshot[5].r.part1[13] , \sa_snapshot[5].r.part1[12] , 
	\sa_snapshot[5].r.part1[11] , \sa_snapshot[5].r.part1[10] , 
	\sa_snapshot[5].r.part1[9] , \sa_snapshot[5].r.part1[8] , 
	\sa_snapshot[5].r.part1[7] , \sa_snapshot[5].r.part1[6] , 
	\sa_snapshot[5].r.part1[5] , \sa_snapshot[5].r.part1[4] , 
	\sa_snapshot[5].r.part1[3] , \sa_snapshot[5].r.part1[2] , 
	\sa_snapshot[5].r.part1[1] , \sa_snapshot[5].r.part1[0] , 
	\sa_snapshot[5].r.part0[31] , \sa_snapshot[5].r.part0[30] , 
	\sa_snapshot[5].r.part0[29] , \sa_snapshot[5].r.part0[28] , 
	\sa_snapshot[5].r.part0[27] , \sa_snapshot[5].r.part0[26] , 
	\sa_snapshot[5].r.part0[25] , \sa_snapshot[5].r.part0[24] , 
	\sa_snapshot[5].r.part0[23] , \sa_snapshot[5].r.part0[22] , 
	\sa_snapshot[5].r.part0[21] , \sa_snapshot[5].r.part0[20] , 
	\sa_snapshot[5].r.part0[19] , \sa_snapshot[5].r.part0[18] , 
	\sa_snapshot[5].r.part0[17] , \sa_snapshot[5].r.part0[16] , 
	\sa_snapshot[5].r.part0[15] , \sa_snapshot[5].r.part0[14] , 
	\sa_snapshot[5].r.part0[13] , \sa_snapshot[5].r.part0[12] , 
	\sa_snapshot[5].r.part0[11] , \sa_snapshot[5].r.part0[10] , 
	\sa_snapshot[5].r.part0[9] , \sa_snapshot[5].r.part0[8] , 
	\sa_snapshot[5].r.part0[7] , \sa_snapshot[5].r.part0[6] , 
	\sa_snapshot[5].r.part0[5] , \sa_snapshot[5].r.part0[4] , 
	\sa_snapshot[5].r.part0[3] , \sa_snapshot[5].r.part0[2] , 
	\sa_snapshot[5].r.part0[1] , \sa_snapshot[5].r.part0[0] , 
	\sa_snapshot[4].r.part1[31] , \sa_snapshot[4].r.part1[30] , 
	\sa_snapshot[4].r.part1[29] , \sa_snapshot[4].r.part1[28] , 
	\sa_snapshot[4].r.part1[27] , \sa_snapshot[4].r.part1[26] , 
	\sa_snapshot[4].r.part1[25] , \sa_snapshot[4].r.part1[24] , 
	\sa_snapshot[4].r.part1[23] , \sa_snapshot[4].r.part1[22] , 
	\sa_snapshot[4].r.part1[21] , \sa_snapshot[4].r.part1[20] , 
	\sa_snapshot[4].r.part1[19] , \sa_snapshot[4].r.part1[18] , 
	\sa_snapshot[4].r.part1[17] , \sa_snapshot[4].r.part1[16] , 
	\sa_snapshot[4].r.part1[15] , \sa_snapshot[4].r.part1[14] , 
	\sa_snapshot[4].r.part1[13] , \sa_snapshot[4].r.part1[12] , 
	\sa_snapshot[4].r.part1[11] , \sa_snapshot[4].r.part1[10] , 
	\sa_snapshot[4].r.part1[9] , \sa_snapshot[4].r.part1[8] , 
	\sa_snapshot[4].r.part1[7] , \sa_snapshot[4].r.part1[6] , 
	\sa_snapshot[4].r.part1[5] , \sa_snapshot[4].r.part1[4] , 
	\sa_snapshot[4].r.part1[3] , \sa_snapshot[4].r.part1[2] , 
	\sa_snapshot[4].r.part1[1] , \sa_snapshot[4].r.part1[0] , 
	\sa_snapshot[4].r.part0[31] , \sa_snapshot[4].r.part0[30] , 
	\sa_snapshot[4].r.part0[29] , \sa_snapshot[4].r.part0[28] , 
	\sa_snapshot[4].r.part0[27] , \sa_snapshot[4].r.part0[26] , 
	\sa_snapshot[4].r.part0[25] , \sa_snapshot[4].r.part0[24] , 
	\sa_snapshot[4].r.part0[23] , \sa_snapshot[4].r.part0[22] , 
	\sa_snapshot[4].r.part0[21] , \sa_snapshot[4].r.part0[20] , 
	\sa_snapshot[4].r.part0[19] , \sa_snapshot[4].r.part0[18] , 
	\sa_snapshot[4].r.part0[17] , \sa_snapshot[4].r.part0[16] , 
	\sa_snapshot[4].r.part0[15] , \sa_snapshot[4].r.part0[14] , 
	\sa_snapshot[4].r.part0[13] , \sa_snapshot[4].r.part0[12] , 
	\sa_snapshot[4].r.part0[11] , \sa_snapshot[4].r.part0[10] , 
	\sa_snapshot[4].r.part0[9] , \sa_snapshot[4].r.part0[8] , 
	\sa_snapshot[4].r.part0[7] , \sa_snapshot[4].r.part0[6] , 
	\sa_snapshot[4].r.part0[5] , \sa_snapshot[4].r.part0[4] , 
	\sa_snapshot[4].r.part0[3] , \sa_snapshot[4].r.part0[2] , 
	\sa_snapshot[4].r.part0[1] , \sa_snapshot[4].r.part0[0] , 
	\sa_snapshot[3].r.part1[31] , \sa_snapshot[3].r.part1[30] , 
	\sa_snapshot[3].r.part1[29] , \sa_snapshot[3].r.part1[28] , 
	\sa_snapshot[3].r.part1[27] , \sa_snapshot[3].r.part1[26] , 
	\sa_snapshot[3].r.part1[25] , \sa_snapshot[3].r.part1[24] , 
	\sa_snapshot[3].r.part1[23] , \sa_snapshot[3].r.part1[22] , 
	\sa_snapshot[3].r.part1[21] , \sa_snapshot[3].r.part1[20] , 
	\sa_snapshot[3].r.part1[19] , \sa_snapshot[3].r.part1[18] , 
	\sa_snapshot[3].r.part1[17] , \sa_snapshot[3].r.part1[16] , 
	\sa_snapshot[3].r.part1[15] , \sa_snapshot[3].r.part1[14] , 
	\sa_snapshot[3].r.part1[13] , \sa_snapshot[3].r.part1[12] , 
	\sa_snapshot[3].r.part1[11] , \sa_snapshot[3].r.part1[10] , 
	\sa_snapshot[3].r.part1[9] , \sa_snapshot[3].r.part1[8] , 
	\sa_snapshot[3].r.part1[7] , \sa_snapshot[3].r.part1[6] , 
	\sa_snapshot[3].r.part1[5] , \sa_snapshot[3].r.part1[4] , 
	\sa_snapshot[3].r.part1[3] , \sa_snapshot[3].r.part1[2] , 
	\sa_snapshot[3].r.part1[1] , \sa_snapshot[3].r.part1[0] , 
	\sa_snapshot[3].r.part0[31] , \sa_snapshot[3].r.part0[30] , 
	\sa_snapshot[3].r.part0[29] , \sa_snapshot[3].r.part0[28] , 
	\sa_snapshot[3].r.part0[27] , \sa_snapshot[3].r.part0[26] , 
	\sa_snapshot[3].r.part0[25] , \sa_snapshot[3].r.part0[24] , 
	\sa_snapshot[3].r.part0[23] , \sa_snapshot[3].r.part0[22] , 
	\sa_snapshot[3].r.part0[21] , \sa_snapshot[3].r.part0[20] , 
	\sa_snapshot[3].r.part0[19] , \sa_snapshot[3].r.part0[18] , 
	\sa_snapshot[3].r.part0[17] , \sa_snapshot[3].r.part0[16] , 
	\sa_snapshot[3].r.part0[15] , \sa_snapshot[3].r.part0[14] , 
	\sa_snapshot[3].r.part0[13] , \sa_snapshot[3].r.part0[12] , 
	\sa_snapshot[3].r.part0[11] , \sa_snapshot[3].r.part0[10] , 
	\sa_snapshot[3].r.part0[9] , \sa_snapshot[3].r.part0[8] , 
	\sa_snapshot[3].r.part0[7] , \sa_snapshot[3].r.part0[6] , 
	\sa_snapshot[3].r.part0[5] , \sa_snapshot[3].r.part0[4] , 
	\sa_snapshot[3].r.part0[3] , \sa_snapshot[3].r.part0[2] , 
	\sa_snapshot[3].r.part0[1] , \sa_snapshot[3].r.part0[0] , 
	\sa_snapshot[2].r.part1[31] , \sa_snapshot[2].r.part1[30] , 
	\sa_snapshot[2].r.part1[29] , \sa_snapshot[2].r.part1[28] , 
	\sa_snapshot[2].r.part1[27] , \sa_snapshot[2].r.part1[26] , 
	\sa_snapshot[2].r.part1[25] , \sa_snapshot[2].r.part1[24] , 
	\sa_snapshot[2].r.part1[23] , \sa_snapshot[2].r.part1[22] , 
	\sa_snapshot[2].r.part1[21] , \sa_snapshot[2].r.part1[20] , 
	\sa_snapshot[2].r.part1[19] , \sa_snapshot[2].r.part1[18] , 
	\sa_snapshot[2].r.part1[17] , \sa_snapshot[2].r.part1[16] , 
	\sa_snapshot[2].r.part1[15] , \sa_snapshot[2].r.part1[14] , 
	\sa_snapshot[2].r.part1[13] , \sa_snapshot[2].r.part1[12] , 
	\sa_snapshot[2].r.part1[11] , \sa_snapshot[2].r.part1[10] , 
	\sa_snapshot[2].r.part1[9] , \sa_snapshot[2].r.part1[8] , 
	\sa_snapshot[2].r.part1[7] , \sa_snapshot[2].r.part1[6] , 
	\sa_snapshot[2].r.part1[5] , \sa_snapshot[2].r.part1[4] , 
	\sa_snapshot[2].r.part1[3] , \sa_snapshot[2].r.part1[2] , 
	\sa_snapshot[2].r.part1[1] , \sa_snapshot[2].r.part1[0] , 
	\sa_snapshot[2].r.part0[31] , \sa_snapshot[2].r.part0[30] , 
	\sa_snapshot[2].r.part0[29] , \sa_snapshot[2].r.part0[28] , 
	\sa_snapshot[2].r.part0[27] , \sa_snapshot[2].r.part0[26] , 
	\sa_snapshot[2].r.part0[25] , \sa_snapshot[2].r.part0[24] , 
	\sa_snapshot[2].r.part0[23] , \sa_snapshot[2].r.part0[22] , 
	\sa_snapshot[2].r.part0[21] , \sa_snapshot[2].r.part0[20] , 
	\sa_snapshot[2].r.part0[19] , \sa_snapshot[2].r.part0[18] , 
	\sa_snapshot[2].r.part0[17] , \sa_snapshot[2].r.part0[16] , 
	\sa_snapshot[2].r.part0[15] , \sa_snapshot[2].r.part0[14] , 
	\sa_snapshot[2].r.part0[13] , \sa_snapshot[2].r.part0[12] , 
	\sa_snapshot[2].r.part0[11] , \sa_snapshot[2].r.part0[10] , 
	\sa_snapshot[2].r.part0[9] , \sa_snapshot[2].r.part0[8] , 
	\sa_snapshot[2].r.part0[7] , \sa_snapshot[2].r.part0[6] , 
	\sa_snapshot[2].r.part0[5] , \sa_snapshot[2].r.part0[4] , 
	\sa_snapshot[2].r.part0[3] , \sa_snapshot[2].r.part0[2] , 
	\sa_snapshot[2].r.part0[1] , \sa_snapshot[2].r.part0[0] , 
	\sa_snapshot[1].r.part1[31] , \sa_snapshot[1].r.part1[30] , 
	\sa_snapshot[1].r.part1[29] , \sa_snapshot[1].r.part1[28] , 
	\sa_snapshot[1].r.part1[27] , \sa_snapshot[1].r.part1[26] , 
	\sa_snapshot[1].r.part1[25] , \sa_snapshot[1].r.part1[24] , 
	\sa_snapshot[1].r.part1[23] , \sa_snapshot[1].r.part1[22] , 
	\sa_snapshot[1].r.part1[21] , \sa_snapshot[1].r.part1[20] , 
	\sa_snapshot[1].r.part1[19] , \sa_snapshot[1].r.part1[18] , 
	\sa_snapshot[1].r.part1[17] , \sa_snapshot[1].r.part1[16] , 
	\sa_snapshot[1].r.part1[15] , \sa_snapshot[1].r.part1[14] , 
	\sa_snapshot[1].r.part1[13] , \sa_snapshot[1].r.part1[12] , 
	\sa_snapshot[1].r.part1[11] , \sa_snapshot[1].r.part1[10] , 
	\sa_snapshot[1].r.part1[9] , \sa_snapshot[1].r.part1[8] , 
	\sa_snapshot[1].r.part1[7] , \sa_snapshot[1].r.part1[6] , 
	\sa_snapshot[1].r.part1[5] , \sa_snapshot[1].r.part1[4] , 
	\sa_snapshot[1].r.part1[3] , \sa_snapshot[1].r.part1[2] , 
	\sa_snapshot[1].r.part1[1] , \sa_snapshot[1].r.part1[0] , 
	\sa_snapshot[1].r.part0[31] , \sa_snapshot[1].r.part0[30] , 
	\sa_snapshot[1].r.part0[29] , \sa_snapshot[1].r.part0[28] , 
	\sa_snapshot[1].r.part0[27] , \sa_snapshot[1].r.part0[26] , 
	\sa_snapshot[1].r.part0[25] , \sa_snapshot[1].r.part0[24] , 
	\sa_snapshot[1].r.part0[23] , \sa_snapshot[1].r.part0[22] , 
	\sa_snapshot[1].r.part0[21] , \sa_snapshot[1].r.part0[20] , 
	\sa_snapshot[1].r.part0[19] , \sa_snapshot[1].r.part0[18] , 
	\sa_snapshot[1].r.part0[17] , \sa_snapshot[1].r.part0[16] , 
	\sa_snapshot[1].r.part0[15] , \sa_snapshot[1].r.part0[14] , 
	\sa_snapshot[1].r.part0[13] , \sa_snapshot[1].r.part0[12] , 
	\sa_snapshot[1].r.part0[11] , \sa_snapshot[1].r.part0[10] , 
	\sa_snapshot[1].r.part0[9] , \sa_snapshot[1].r.part0[8] , 
	\sa_snapshot[1].r.part0[7] , \sa_snapshot[1].r.part0[6] , 
	\sa_snapshot[1].r.part0[5] , \sa_snapshot[1].r.part0[4] , 
	\sa_snapshot[1].r.part0[3] , \sa_snapshot[1].r.part0[2] , 
	\sa_snapshot[1].r.part0[1] , \sa_snapshot[1].r.part0[0] , 
	\sa_snapshot[0].r.part1[31] , \sa_snapshot[0].r.part1[30] , 
	\sa_snapshot[0].r.part1[29] , \sa_snapshot[0].r.part1[28] , 
	\sa_snapshot[0].r.part1[27] , \sa_snapshot[0].r.part1[26] , 
	\sa_snapshot[0].r.part1[25] , \sa_snapshot[0].r.part1[24] , 
	\sa_snapshot[0].r.part1[23] , \sa_snapshot[0].r.part1[22] , 
	\sa_snapshot[0].r.part1[21] , \sa_snapshot[0].r.part1[20] , 
	\sa_snapshot[0].r.part1[19] , \sa_snapshot[0].r.part1[18] , 
	\sa_snapshot[0].r.part1[17] , \sa_snapshot[0].r.part1[16] , 
	\sa_snapshot[0].r.part1[15] , \sa_snapshot[0].r.part1[14] , 
	\sa_snapshot[0].r.part1[13] , \sa_snapshot[0].r.part1[12] , 
	\sa_snapshot[0].r.part1[11] , \sa_snapshot[0].r.part1[10] , 
	\sa_snapshot[0].r.part1[9] , \sa_snapshot[0].r.part1[8] , 
	\sa_snapshot[0].r.part1[7] , \sa_snapshot[0].r.part1[6] , 
	\sa_snapshot[0].r.part1[5] , \sa_snapshot[0].r.part1[4] , 
	\sa_snapshot[0].r.part1[3] , \sa_snapshot[0].r.part1[2] , 
	\sa_snapshot[0].r.part1[1] , \sa_snapshot[0].r.part1[0] , 
	\sa_snapshot[0].r.part0[31] , \sa_snapshot[0].r.part0[30] , 
	\sa_snapshot[0].r.part0[29] , \sa_snapshot[0].r.part0[28] , 
	\sa_snapshot[0].r.part0[27] , \sa_snapshot[0].r.part0[26] , 
	\sa_snapshot[0].r.part0[25] , \sa_snapshot[0].r.part0[24] , 
	\sa_snapshot[0].r.part0[23] , \sa_snapshot[0].r.part0[22] , 
	\sa_snapshot[0].r.part0[21] , \sa_snapshot[0].r.part0[20] , 
	\sa_snapshot[0].r.part0[19] , \sa_snapshot[0].r.part0[18] , 
	\sa_snapshot[0].r.part0[17] , \sa_snapshot[0].r.part0[16] , 
	\sa_snapshot[0].r.part0[15] , \sa_snapshot[0].r.part0[14] , 
	\sa_snapshot[0].r.part0[13] , \sa_snapshot[0].r.part0[12] , 
	\sa_snapshot[0].r.part0[11] , \sa_snapshot[0].r.part0[10] , 
	\sa_snapshot[0].r.part0[9] , \sa_snapshot[0].r.part0[8] , 
	\sa_snapshot[0].r.part0[7] , \sa_snapshot[0].r.part0[6] , 
	\sa_snapshot[0].r.part0[5] , \sa_snapshot[0].r.part0[4] , 
	\sa_snapshot[0].r.part0[3] , \sa_snapshot[0].r.part0[2] , 
	\sa_snapshot[0].r.part0[1] , \sa_snapshot[0].r.part0[0] } ), 
	.sa_count( {\sa_count[31].r.part1[31] , \sa_count[31].r.part1[30] , 
	\sa_count[31].r.part1[29] , \sa_count[31].r.part1[28] , 
	\sa_count[31].r.part1[27] , \sa_count[31].r.part1[26] , 
	\sa_count[31].r.part1[25] , \sa_count[31].r.part1[24] , 
	\sa_count[31].r.part1[23] , \sa_count[31].r.part1[22] , 
	\sa_count[31].r.part1[21] , \sa_count[31].r.part1[20] , 
	\sa_count[31].r.part1[19] , \sa_count[31].r.part1[18] , 
	\sa_count[31].r.part1[17] , \sa_count[31].r.part1[16] , 
	\sa_count[31].r.part1[15] , \sa_count[31].r.part1[14] , 
	\sa_count[31].r.part1[13] , \sa_count[31].r.part1[12] , 
	\sa_count[31].r.part1[11] , \sa_count[31].r.part1[10] , 
	\sa_count[31].r.part1[9] , \sa_count[31].r.part1[8] , 
	\sa_count[31].r.part1[7] , \sa_count[31].r.part1[6] , 
	\sa_count[31].r.part1[5] , \sa_count[31].r.part1[4] , 
	\sa_count[31].r.part1[3] , \sa_count[31].r.part1[2] , 
	\sa_count[31].r.part1[1] , \sa_count[31].r.part1[0] , 
	\sa_count[31].r.part0[31] , \sa_count[31].r.part0[30] , 
	\sa_count[31].r.part0[29] , \sa_count[31].r.part0[28] , 
	\sa_count[31].r.part0[27] , \sa_count[31].r.part0[26] , 
	\sa_count[31].r.part0[25] , \sa_count[31].r.part0[24] , 
	\sa_count[31].r.part0[23] , \sa_count[31].r.part0[22] , 
	\sa_count[31].r.part0[21] , \sa_count[31].r.part0[20] , 
	\sa_count[31].r.part0[19] , \sa_count[31].r.part0[18] , 
	\sa_count[31].r.part0[17] , \sa_count[31].r.part0[16] , 
	\sa_count[31].r.part0[15] , \sa_count[31].r.part0[14] , 
	\sa_count[31].r.part0[13] , \sa_count[31].r.part0[12] , 
	\sa_count[31].r.part0[11] , \sa_count[31].r.part0[10] , 
	\sa_count[31].r.part0[9] , \sa_count[31].r.part0[8] , 
	\sa_count[31].r.part0[7] , \sa_count[31].r.part0[6] , 
	\sa_count[31].r.part0[5] , \sa_count[31].r.part0[4] , 
	\sa_count[31].r.part0[3] , \sa_count[31].r.part0[2] , 
	\sa_count[31].r.part0[1] , \sa_count[31].r.part0[0] , 
	\sa_count[30].r.part1[31] , \sa_count[30].r.part1[30] , 
	\sa_count[30].r.part1[29] , \sa_count[30].r.part1[28] , 
	\sa_count[30].r.part1[27] , \sa_count[30].r.part1[26] , 
	\sa_count[30].r.part1[25] , \sa_count[30].r.part1[24] , 
	\sa_count[30].r.part1[23] , \sa_count[30].r.part1[22] , 
	\sa_count[30].r.part1[21] , \sa_count[30].r.part1[20] , 
	\sa_count[30].r.part1[19] , \sa_count[30].r.part1[18] , 
	\sa_count[30].r.part1[17] , \sa_count[30].r.part1[16] , 
	\sa_count[30].r.part1[15] , \sa_count[30].r.part1[14] , 
	\sa_count[30].r.part1[13] , \sa_count[30].r.part1[12] , 
	\sa_count[30].r.part1[11] , \sa_count[30].r.part1[10] , 
	\sa_count[30].r.part1[9] , \sa_count[30].r.part1[8] , 
	\sa_count[30].r.part1[7] , \sa_count[30].r.part1[6] , 
	\sa_count[30].r.part1[5] , \sa_count[30].r.part1[4] , 
	\sa_count[30].r.part1[3] , \sa_count[30].r.part1[2] , 
	\sa_count[30].r.part1[1] , \sa_count[30].r.part1[0] , 
	\sa_count[30].r.part0[31] , \sa_count[30].r.part0[30] , 
	\sa_count[30].r.part0[29] , \sa_count[30].r.part0[28] , 
	\sa_count[30].r.part0[27] , \sa_count[30].r.part0[26] , 
	\sa_count[30].r.part0[25] , \sa_count[30].r.part0[24] , 
	\sa_count[30].r.part0[23] , \sa_count[30].r.part0[22] , 
	\sa_count[30].r.part0[21] , \sa_count[30].r.part0[20] , 
	\sa_count[30].r.part0[19] , \sa_count[30].r.part0[18] , 
	\sa_count[30].r.part0[17] , \sa_count[30].r.part0[16] , 
	\sa_count[30].r.part0[15] , \sa_count[30].r.part0[14] , 
	\sa_count[30].r.part0[13] , \sa_count[30].r.part0[12] , 
	\sa_count[30].r.part0[11] , \sa_count[30].r.part0[10] , 
	\sa_count[30].r.part0[9] , \sa_count[30].r.part0[8] , 
	\sa_count[30].r.part0[7] , \sa_count[30].r.part0[6] , 
	\sa_count[30].r.part0[5] , \sa_count[30].r.part0[4] , 
	\sa_count[30].r.part0[3] , \sa_count[30].r.part0[2] , 
	\sa_count[30].r.part0[1] , \sa_count[30].r.part0[0] , 
	\sa_count[29].r.part1[31] , \sa_count[29].r.part1[30] , 
	\sa_count[29].r.part1[29] , \sa_count[29].r.part1[28] , 
	\sa_count[29].r.part1[27] , \sa_count[29].r.part1[26] , 
	\sa_count[29].r.part1[25] , \sa_count[29].r.part1[24] , 
	\sa_count[29].r.part1[23] , \sa_count[29].r.part1[22] , 
	\sa_count[29].r.part1[21] , \sa_count[29].r.part1[20] , 
	\sa_count[29].r.part1[19] , \sa_count[29].r.part1[18] , 
	\sa_count[29].r.part1[17] , \sa_count[29].r.part1[16] , 
	\sa_count[29].r.part1[15] , \sa_count[29].r.part1[14] , 
	\sa_count[29].r.part1[13] , \sa_count[29].r.part1[12] , 
	\sa_count[29].r.part1[11] , \sa_count[29].r.part1[10] , 
	\sa_count[29].r.part1[9] , \sa_count[29].r.part1[8] , 
	\sa_count[29].r.part1[7] , \sa_count[29].r.part1[6] , 
	\sa_count[29].r.part1[5] , \sa_count[29].r.part1[4] , 
	\sa_count[29].r.part1[3] , \sa_count[29].r.part1[2] , 
	\sa_count[29].r.part1[1] , \sa_count[29].r.part1[0] , 
	\sa_count[29].r.part0[31] , \sa_count[29].r.part0[30] , 
	\sa_count[29].r.part0[29] , \sa_count[29].r.part0[28] , 
	\sa_count[29].r.part0[27] , \sa_count[29].r.part0[26] , 
	\sa_count[29].r.part0[25] , \sa_count[29].r.part0[24] , 
	\sa_count[29].r.part0[23] , \sa_count[29].r.part0[22] , 
	\sa_count[29].r.part0[21] , \sa_count[29].r.part0[20] , 
	\sa_count[29].r.part0[19] , \sa_count[29].r.part0[18] , 
	\sa_count[29].r.part0[17] , \sa_count[29].r.part0[16] , 
	\sa_count[29].r.part0[15] , \sa_count[29].r.part0[14] , 
	\sa_count[29].r.part0[13] , \sa_count[29].r.part0[12] , 
	\sa_count[29].r.part0[11] , \sa_count[29].r.part0[10] , 
	\sa_count[29].r.part0[9] , \sa_count[29].r.part0[8] , 
	\sa_count[29].r.part0[7] , \sa_count[29].r.part0[6] , 
	\sa_count[29].r.part0[5] , \sa_count[29].r.part0[4] , 
	\sa_count[29].r.part0[3] , \sa_count[29].r.part0[2] , 
	\sa_count[29].r.part0[1] , \sa_count[29].r.part0[0] , 
	\sa_count[28].r.part1[31] , \sa_count[28].r.part1[30] , 
	\sa_count[28].r.part1[29] , \sa_count[28].r.part1[28] , 
	\sa_count[28].r.part1[27] , \sa_count[28].r.part1[26] , 
	\sa_count[28].r.part1[25] , \sa_count[28].r.part1[24] , 
	\sa_count[28].r.part1[23] , \sa_count[28].r.part1[22] , 
	\sa_count[28].r.part1[21] , \sa_count[28].r.part1[20] , 
	\sa_count[28].r.part1[19] , \sa_count[28].r.part1[18] , 
	\sa_count[28].r.part1[17] , \sa_count[28].r.part1[16] , 
	\sa_count[28].r.part1[15] , \sa_count[28].r.part1[14] , 
	\sa_count[28].r.part1[13] , \sa_count[28].r.part1[12] , 
	\sa_count[28].r.part1[11] , \sa_count[28].r.part1[10] , 
	\sa_count[28].r.part1[9] , \sa_count[28].r.part1[8] , 
	\sa_count[28].r.part1[7] , \sa_count[28].r.part1[6] , 
	\sa_count[28].r.part1[5] , \sa_count[28].r.part1[4] , 
	\sa_count[28].r.part1[3] , \sa_count[28].r.part1[2] , 
	\sa_count[28].r.part1[1] , \sa_count[28].r.part1[0] , 
	\sa_count[28].r.part0[31] , \sa_count[28].r.part0[30] , 
	\sa_count[28].r.part0[29] , \sa_count[28].r.part0[28] , 
	\sa_count[28].r.part0[27] , \sa_count[28].r.part0[26] , 
	\sa_count[28].r.part0[25] , \sa_count[28].r.part0[24] , 
	\sa_count[28].r.part0[23] , \sa_count[28].r.part0[22] , 
	\sa_count[28].r.part0[21] , \sa_count[28].r.part0[20] , 
	\sa_count[28].r.part0[19] , \sa_count[28].r.part0[18] , 
	\sa_count[28].r.part0[17] , \sa_count[28].r.part0[16] , 
	\sa_count[28].r.part0[15] , \sa_count[28].r.part0[14] , 
	\sa_count[28].r.part0[13] , \sa_count[28].r.part0[12] , 
	\sa_count[28].r.part0[11] , \sa_count[28].r.part0[10] , 
	\sa_count[28].r.part0[9] , \sa_count[28].r.part0[8] , 
	\sa_count[28].r.part0[7] , \sa_count[28].r.part0[6] , 
	\sa_count[28].r.part0[5] , \sa_count[28].r.part0[4] , 
	\sa_count[28].r.part0[3] , \sa_count[28].r.part0[2] , 
	\sa_count[28].r.part0[1] , \sa_count[28].r.part0[0] , 
	\sa_count[27].r.part1[31] , \sa_count[27].r.part1[30] , 
	\sa_count[27].r.part1[29] , \sa_count[27].r.part1[28] , 
	\sa_count[27].r.part1[27] , \sa_count[27].r.part1[26] , 
	\sa_count[27].r.part1[25] , \sa_count[27].r.part1[24] , 
	\sa_count[27].r.part1[23] , \sa_count[27].r.part1[22] , 
	\sa_count[27].r.part1[21] , \sa_count[27].r.part1[20] , 
	\sa_count[27].r.part1[19] , \sa_count[27].r.part1[18] , 
	\sa_count[27].r.part1[17] , \sa_count[27].r.part1[16] , 
	\sa_count[27].r.part1[15] , \sa_count[27].r.part1[14] , 
	\sa_count[27].r.part1[13] , \sa_count[27].r.part1[12] , 
	\sa_count[27].r.part1[11] , \sa_count[27].r.part1[10] , 
	\sa_count[27].r.part1[9] , \sa_count[27].r.part1[8] , 
	\sa_count[27].r.part1[7] , \sa_count[27].r.part1[6] , 
	\sa_count[27].r.part1[5] , \sa_count[27].r.part1[4] , 
	\sa_count[27].r.part1[3] , \sa_count[27].r.part1[2] , 
	\sa_count[27].r.part1[1] , \sa_count[27].r.part1[0] , 
	\sa_count[27].r.part0[31] , \sa_count[27].r.part0[30] , 
	\sa_count[27].r.part0[29] , \sa_count[27].r.part0[28] , 
	\sa_count[27].r.part0[27] , \sa_count[27].r.part0[26] , 
	\sa_count[27].r.part0[25] , \sa_count[27].r.part0[24] , 
	\sa_count[27].r.part0[23] , \sa_count[27].r.part0[22] , 
	\sa_count[27].r.part0[21] , \sa_count[27].r.part0[20] , 
	\sa_count[27].r.part0[19] , \sa_count[27].r.part0[18] , 
	\sa_count[27].r.part0[17] , \sa_count[27].r.part0[16] , 
	\sa_count[27].r.part0[15] , \sa_count[27].r.part0[14] , 
	\sa_count[27].r.part0[13] , \sa_count[27].r.part0[12] , 
	\sa_count[27].r.part0[11] , \sa_count[27].r.part0[10] , 
	\sa_count[27].r.part0[9] , \sa_count[27].r.part0[8] , 
	\sa_count[27].r.part0[7] , \sa_count[27].r.part0[6] , 
	\sa_count[27].r.part0[5] , \sa_count[27].r.part0[4] , 
	\sa_count[27].r.part0[3] , \sa_count[27].r.part0[2] , 
	\sa_count[27].r.part0[1] , \sa_count[27].r.part0[0] , 
	\sa_count[26].r.part1[31] , \sa_count[26].r.part1[30] , 
	\sa_count[26].r.part1[29] , \sa_count[26].r.part1[28] , 
	\sa_count[26].r.part1[27] , \sa_count[26].r.part1[26] , 
	\sa_count[26].r.part1[25] , \sa_count[26].r.part1[24] , 
	\sa_count[26].r.part1[23] , \sa_count[26].r.part1[22] , 
	\sa_count[26].r.part1[21] , \sa_count[26].r.part1[20] , 
	\sa_count[26].r.part1[19] , \sa_count[26].r.part1[18] , 
	\sa_count[26].r.part1[17] , \sa_count[26].r.part1[16] , 
	\sa_count[26].r.part1[15] , \sa_count[26].r.part1[14] , 
	\sa_count[26].r.part1[13] , \sa_count[26].r.part1[12] , 
	\sa_count[26].r.part1[11] , \sa_count[26].r.part1[10] , 
	\sa_count[26].r.part1[9] , \sa_count[26].r.part1[8] , 
	\sa_count[26].r.part1[7] , \sa_count[26].r.part1[6] , 
	\sa_count[26].r.part1[5] , \sa_count[26].r.part1[4] , 
	\sa_count[26].r.part1[3] , \sa_count[26].r.part1[2] , 
	\sa_count[26].r.part1[1] , \sa_count[26].r.part1[0] , 
	\sa_count[26].r.part0[31] , \sa_count[26].r.part0[30] , 
	\sa_count[26].r.part0[29] , \sa_count[26].r.part0[28] , 
	\sa_count[26].r.part0[27] , \sa_count[26].r.part0[26] , 
	\sa_count[26].r.part0[25] , \sa_count[26].r.part0[24] , 
	\sa_count[26].r.part0[23] , \sa_count[26].r.part0[22] , 
	\sa_count[26].r.part0[21] , \sa_count[26].r.part0[20] , 
	\sa_count[26].r.part0[19] , \sa_count[26].r.part0[18] , 
	\sa_count[26].r.part0[17] , \sa_count[26].r.part0[16] , 
	\sa_count[26].r.part0[15] , \sa_count[26].r.part0[14] , 
	\sa_count[26].r.part0[13] , \sa_count[26].r.part0[12] , 
	\sa_count[26].r.part0[11] , \sa_count[26].r.part0[10] , 
	\sa_count[26].r.part0[9] , \sa_count[26].r.part0[8] , 
	\sa_count[26].r.part0[7] , \sa_count[26].r.part0[6] , 
	\sa_count[26].r.part0[5] , \sa_count[26].r.part0[4] , 
	\sa_count[26].r.part0[3] , \sa_count[26].r.part0[2] , 
	\sa_count[26].r.part0[1] , \sa_count[26].r.part0[0] , 
	\sa_count[25].r.part1[31] , \sa_count[25].r.part1[30] , 
	\sa_count[25].r.part1[29] , \sa_count[25].r.part1[28] , 
	\sa_count[25].r.part1[27] , \sa_count[25].r.part1[26] , 
	\sa_count[25].r.part1[25] , \sa_count[25].r.part1[24] , 
	\sa_count[25].r.part1[23] , \sa_count[25].r.part1[22] , 
	\sa_count[25].r.part1[21] , \sa_count[25].r.part1[20] , 
	\sa_count[25].r.part1[19] , \sa_count[25].r.part1[18] , 
	\sa_count[25].r.part1[17] , \sa_count[25].r.part1[16] , 
	\sa_count[25].r.part1[15] , \sa_count[25].r.part1[14] , 
	\sa_count[25].r.part1[13] , \sa_count[25].r.part1[12] , 
	\sa_count[25].r.part1[11] , \sa_count[25].r.part1[10] , 
	\sa_count[25].r.part1[9] , \sa_count[25].r.part1[8] , 
	\sa_count[25].r.part1[7] , \sa_count[25].r.part1[6] , 
	\sa_count[25].r.part1[5] , \sa_count[25].r.part1[4] , 
	\sa_count[25].r.part1[3] , \sa_count[25].r.part1[2] , 
	\sa_count[25].r.part1[1] , \sa_count[25].r.part1[0] , 
	\sa_count[25].r.part0[31] , \sa_count[25].r.part0[30] , 
	\sa_count[25].r.part0[29] , \sa_count[25].r.part0[28] , 
	\sa_count[25].r.part0[27] , \sa_count[25].r.part0[26] , 
	\sa_count[25].r.part0[25] , \sa_count[25].r.part0[24] , 
	\sa_count[25].r.part0[23] , \sa_count[25].r.part0[22] , 
	\sa_count[25].r.part0[21] , \sa_count[25].r.part0[20] , 
	\sa_count[25].r.part0[19] , \sa_count[25].r.part0[18] , 
	\sa_count[25].r.part0[17] , \sa_count[25].r.part0[16] , 
	\sa_count[25].r.part0[15] , \sa_count[25].r.part0[14] , 
	\sa_count[25].r.part0[13] , \sa_count[25].r.part0[12] , 
	\sa_count[25].r.part0[11] , \sa_count[25].r.part0[10] , 
	\sa_count[25].r.part0[9] , \sa_count[25].r.part0[8] , 
	\sa_count[25].r.part0[7] , \sa_count[25].r.part0[6] , 
	\sa_count[25].r.part0[5] , \sa_count[25].r.part0[4] , 
	\sa_count[25].r.part0[3] , \sa_count[25].r.part0[2] , 
	\sa_count[25].r.part0[1] , \sa_count[25].r.part0[0] , 
	\sa_count[24].r.part1[31] , \sa_count[24].r.part1[30] , 
	\sa_count[24].r.part1[29] , \sa_count[24].r.part1[28] , 
	\sa_count[24].r.part1[27] , \sa_count[24].r.part1[26] , 
	\sa_count[24].r.part1[25] , \sa_count[24].r.part1[24] , 
	\sa_count[24].r.part1[23] , \sa_count[24].r.part1[22] , 
	\sa_count[24].r.part1[21] , \sa_count[24].r.part1[20] , 
	\sa_count[24].r.part1[19] , \sa_count[24].r.part1[18] , 
	\sa_count[24].r.part1[17] , \sa_count[24].r.part1[16] , 
	\sa_count[24].r.part1[15] , \sa_count[24].r.part1[14] , 
	\sa_count[24].r.part1[13] , \sa_count[24].r.part1[12] , 
	\sa_count[24].r.part1[11] , \sa_count[24].r.part1[10] , 
	\sa_count[24].r.part1[9] , \sa_count[24].r.part1[8] , 
	\sa_count[24].r.part1[7] , \sa_count[24].r.part1[6] , 
	\sa_count[24].r.part1[5] , \sa_count[24].r.part1[4] , 
	\sa_count[24].r.part1[3] , \sa_count[24].r.part1[2] , 
	\sa_count[24].r.part1[1] , \sa_count[24].r.part1[0] , 
	\sa_count[24].r.part0[31] , \sa_count[24].r.part0[30] , 
	\sa_count[24].r.part0[29] , \sa_count[24].r.part0[28] , 
	\sa_count[24].r.part0[27] , \sa_count[24].r.part0[26] , 
	\sa_count[24].r.part0[25] , \sa_count[24].r.part0[24] , 
	\sa_count[24].r.part0[23] , \sa_count[24].r.part0[22] , 
	\sa_count[24].r.part0[21] , \sa_count[24].r.part0[20] , 
	\sa_count[24].r.part0[19] , \sa_count[24].r.part0[18] , 
	\sa_count[24].r.part0[17] , \sa_count[24].r.part0[16] , 
	\sa_count[24].r.part0[15] , \sa_count[24].r.part0[14] , 
	\sa_count[24].r.part0[13] , \sa_count[24].r.part0[12] , 
	\sa_count[24].r.part0[11] , \sa_count[24].r.part0[10] , 
	\sa_count[24].r.part0[9] , \sa_count[24].r.part0[8] , 
	\sa_count[24].r.part0[7] , \sa_count[24].r.part0[6] , 
	\sa_count[24].r.part0[5] , \sa_count[24].r.part0[4] , 
	\sa_count[24].r.part0[3] , \sa_count[24].r.part0[2] , 
	\sa_count[24].r.part0[1] , \sa_count[24].r.part0[0] , 
	\sa_count[23].r.part1[31] , \sa_count[23].r.part1[30] , 
	\sa_count[23].r.part1[29] , \sa_count[23].r.part1[28] , 
	\sa_count[23].r.part1[27] , \sa_count[23].r.part1[26] , 
	\sa_count[23].r.part1[25] , \sa_count[23].r.part1[24] , 
	\sa_count[23].r.part1[23] , \sa_count[23].r.part1[22] , 
	\sa_count[23].r.part1[21] , \sa_count[23].r.part1[20] , 
	\sa_count[23].r.part1[19] , \sa_count[23].r.part1[18] , 
	\sa_count[23].r.part1[17] , \sa_count[23].r.part1[16] , 
	\sa_count[23].r.part1[15] , \sa_count[23].r.part1[14] , 
	\sa_count[23].r.part1[13] , \sa_count[23].r.part1[12] , 
	\sa_count[23].r.part1[11] , \sa_count[23].r.part1[10] , 
	\sa_count[23].r.part1[9] , \sa_count[23].r.part1[8] , 
	\sa_count[23].r.part1[7] , \sa_count[23].r.part1[6] , 
	\sa_count[23].r.part1[5] , \sa_count[23].r.part1[4] , 
	\sa_count[23].r.part1[3] , \sa_count[23].r.part1[2] , 
	\sa_count[23].r.part1[1] , \sa_count[23].r.part1[0] , 
	\sa_count[23].r.part0[31] , \sa_count[23].r.part0[30] , 
	\sa_count[23].r.part0[29] , \sa_count[23].r.part0[28] , 
	\sa_count[23].r.part0[27] , \sa_count[23].r.part0[26] , 
	\sa_count[23].r.part0[25] , \sa_count[23].r.part0[24] , 
	\sa_count[23].r.part0[23] , \sa_count[23].r.part0[22] , 
	\sa_count[23].r.part0[21] , \sa_count[23].r.part0[20] , 
	\sa_count[23].r.part0[19] , \sa_count[23].r.part0[18] , 
	\sa_count[23].r.part0[17] , \sa_count[23].r.part0[16] , 
	\sa_count[23].r.part0[15] , \sa_count[23].r.part0[14] , 
	\sa_count[23].r.part0[13] , \sa_count[23].r.part0[12] , 
	\sa_count[23].r.part0[11] , \sa_count[23].r.part0[10] , 
	\sa_count[23].r.part0[9] , \sa_count[23].r.part0[8] , 
	\sa_count[23].r.part0[7] , \sa_count[23].r.part0[6] , 
	\sa_count[23].r.part0[5] , \sa_count[23].r.part0[4] , 
	\sa_count[23].r.part0[3] , \sa_count[23].r.part0[2] , 
	\sa_count[23].r.part0[1] , \sa_count[23].r.part0[0] , 
	\sa_count[22].r.part1[31] , \sa_count[22].r.part1[30] , 
	\sa_count[22].r.part1[29] , \sa_count[22].r.part1[28] , 
	\sa_count[22].r.part1[27] , \sa_count[22].r.part1[26] , 
	\sa_count[22].r.part1[25] , \sa_count[22].r.part1[24] , 
	\sa_count[22].r.part1[23] , \sa_count[22].r.part1[22] , 
	\sa_count[22].r.part1[21] , \sa_count[22].r.part1[20] , 
	\sa_count[22].r.part1[19] , \sa_count[22].r.part1[18] , 
	\sa_count[22].r.part1[17] , \sa_count[22].r.part1[16] , 
	\sa_count[22].r.part1[15] , \sa_count[22].r.part1[14] , 
	\sa_count[22].r.part1[13] , \sa_count[22].r.part1[12] , 
	\sa_count[22].r.part1[11] , \sa_count[22].r.part1[10] , 
	\sa_count[22].r.part1[9] , \sa_count[22].r.part1[8] , 
	\sa_count[22].r.part1[7] , \sa_count[22].r.part1[6] , 
	\sa_count[22].r.part1[5] , \sa_count[22].r.part1[4] , 
	\sa_count[22].r.part1[3] , \sa_count[22].r.part1[2] , 
	\sa_count[22].r.part1[1] , \sa_count[22].r.part1[0] , 
	\sa_count[22].r.part0[31] , \sa_count[22].r.part0[30] , 
	\sa_count[22].r.part0[29] , \sa_count[22].r.part0[28] , 
	\sa_count[22].r.part0[27] , \sa_count[22].r.part0[26] , 
	\sa_count[22].r.part0[25] , \sa_count[22].r.part0[24] , 
	\sa_count[22].r.part0[23] , \sa_count[22].r.part0[22] , 
	\sa_count[22].r.part0[21] , \sa_count[22].r.part0[20] , 
	\sa_count[22].r.part0[19] , \sa_count[22].r.part0[18] , 
	\sa_count[22].r.part0[17] , \sa_count[22].r.part0[16] , 
	\sa_count[22].r.part0[15] , \sa_count[22].r.part0[14] , 
	\sa_count[22].r.part0[13] , \sa_count[22].r.part0[12] , 
	\sa_count[22].r.part0[11] , \sa_count[22].r.part0[10] , 
	\sa_count[22].r.part0[9] , \sa_count[22].r.part0[8] , 
	\sa_count[22].r.part0[7] , \sa_count[22].r.part0[6] , 
	\sa_count[22].r.part0[5] , \sa_count[22].r.part0[4] , 
	\sa_count[22].r.part0[3] , \sa_count[22].r.part0[2] , 
	\sa_count[22].r.part0[1] , \sa_count[22].r.part0[0] , 
	\sa_count[21].r.part1[31] , \sa_count[21].r.part1[30] , 
	\sa_count[21].r.part1[29] , \sa_count[21].r.part1[28] , 
	\sa_count[21].r.part1[27] , \sa_count[21].r.part1[26] , 
	\sa_count[21].r.part1[25] , \sa_count[21].r.part1[24] , 
	\sa_count[21].r.part1[23] , \sa_count[21].r.part1[22] , 
	\sa_count[21].r.part1[21] , \sa_count[21].r.part1[20] , 
	\sa_count[21].r.part1[19] , \sa_count[21].r.part1[18] , 
	\sa_count[21].r.part1[17] , \sa_count[21].r.part1[16] , 
	\sa_count[21].r.part1[15] , \sa_count[21].r.part1[14] , 
	\sa_count[21].r.part1[13] , \sa_count[21].r.part1[12] , 
	\sa_count[21].r.part1[11] , \sa_count[21].r.part1[10] , 
	\sa_count[21].r.part1[9] , \sa_count[21].r.part1[8] , 
	\sa_count[21].r.part1[7] , \sa_count[21].r.part1[6] , 
	\sa_count[21].r.part1[5] , \sa_count[21].r.part1[4] , 
	\sa_count[21].r.part1[3] , \sa_count[21].r.part1[2] , 
	\sa_count[21].r.part1[1] , \sa_count[21].r.part1[0] , 
	\sa_count[21].r.part0[31] , \sa_count[21].r.part0[30] , 
	\sa_count[21].r.part0[29] , \sa_count[21].r.part0[28] , 
	\sa_count[21].r.part0[27] , \sa_count[21].r.part0[26] , 
	\sa_count[21].r.part0[25] , \sa_count[21].r.part0[24] , 
	\sa_count[21].r.part0[23] , \sa_count[21].r.part0[22] , 
	\sa_count[21].r.part0[21] , \sa_count[21].r.part0[20] , 
	\sa_count[21].r.part0[19] , \sa_count[21].r.part0[18] , 
	\sa_count[21].r.part0[17] , \sa_count[21].r.part0[16] , 
	\sa_count[21].r.part0[15] , \sa_count[21].r.part0[14] , 
	\sa_count[21].r.part0[13] , \sa_count[21].r.part0[12] , 
	\sa_count[21].r.part0[11] , \sa_count[21].r.part0[10] , 
	\sa_count[21].r.part0[9] , \sa_count[21].r.part0[8] , 
	\sa_count[21].r.part0[7] , \sa_count[21].r.part0[6] , 
	\sa_count[21].r.part0[5] , \sa_count[21].r.part0[4] , 
	\sa_count[21].r.part0[3] , \sa_count[21].r.part0[2] , 
	\sa_count[21].r.part0[1] , \sa_count[21].r.part0[0] , 
	\sa_count[20].r.part1[31] , \sa_count[20].r.part1[30] , 
	\sa_count[20].r.part1[29] , \sa_count[20].r.part1[28] , 
	\sa_count[20].r.part1[27] , \sa_count[20].r.part1[26] , 
	\sa_count[20].r.part1[25] , \sa_count[20].r.part1[24] , 
	\sa_count[20].r.part1[23] , \sa_count[20].r.part1[22] , 
	\sa_count[20].r.part1[21] , \sa_count[20].r.part1[20] , 
	\sa_count[20].r.part1[19] , \sa_count[20].r.part1[18] , 
	\sa_count[20].r.part1[17] , \sa_count[20].r.part1[16] , 
	\sa_count[20].r.part1[15] , \sa_count[20].r.part1[14] , 
	\sa_count[20].r.part1[13] , \sa_count[20].r.part1[12] , 
	\sa_count[20].r.part1[11] , \sa_count[20].r.part1[10] , 
	\sa_count[20].r.part1[9] , \sa_count[20].r.part1[8] , 
	\sa_count[20].r.part1[7] , \sa_count[20].r.part1[6] , 
	\sa_count[20].r.part1[5] , \sa_count[20].r.part1[4] , 
	\sa_count[20].r.part1[3] , \sa_count[20].r.part1[2] , 
	\sa_count[20].r.part1[1] , \sa_count[20].r.part1[0] , 
	\sa_count[20].r.part0[31] , \sa_count[20].r.part0[30] , 
	\sa_count[20].r.part0[29] , \sa_count[20].r.part0[28] , 
	\sa_count[20].r.part0[27] , \sa_count[20].r.part0[26] , 
	\sa_count[20].r.part0[25] , \sa_count[20].r.part0[24] , 
	\sa_count[20].r.part0[23] , \sa_count[20].r.part0[22] , 
	\sa_count[20].r.part0[21] , \sa_count[20].r.part0[20] , 
	\sa_count[20].r.part0[19] , \sa_count[20].r.part0[18] , 
	\sa_count[20].r.part0[17] , \sa_count[20].r.part0[16] , 
	\sa_count[20].r.part0[15] , \sa_count[20].r.part0[14] , 
	\sa_count[20].r.part0[13] , \sa_count[20].r.part0[12] , 
	\sa_count[20].r.part0[11] , \sa_count[20].r.part0[10] , 
	\sa_count[20].r.part0[9] , \sa_count[20].r.part0[8] , 
	\sa_count[20].r.part0[7] , \sa_count[20].r.part0[6] , 
	\sa_count[20].r.part0[5] , \sa_count[20].r.part0[4] , 
	\sa_count[20].r.part0[3] , \sa_count[20].r.part0[2] , 
	\sa_count[20].r.part0[1] , \sa_count[20].r.part0[0] , 
	\sa_count[19].r.part1[31] , \sa_count[19].r.part1[30] , 
	\sa_count[19].r.part1[29] , \sa_count[19].r.part1[28] , 
	\sa_count[19].r.part1[27] , \sa_count[19].r.part1[26] , 
	\sa_count[19].r.part1[25] , \sa_count[19].r.part1[24] , 
	\sa_count[19].r.part1[23] , \sa_count[19].r.part1[22] , 
	\sa_count[19].r.part1[21] , \sa_count[19].r.part1[20] , 
	\sa_count[19].r.part1[19] , \sa_count[19].r.part1[18] , 
	\sa_count[19].r.part1[17] , \sa_count[19].r.part1[16] , 
	\sa_count[19].r.part1[15] , \sa_count[19].r.part1[14] , 
	\sa_count[19].r.part1[13] , \sa_count[19].r.part1[12] , 
	\sa_count[19].r.part1[11] , \sa_count[19].r.part1[10] , 
	\sa_count[19].r.part1[9] , \sa_count[19].r.part1[8] , 
	\sa_count[19].r.part1[7] , \sa_count[19].r.part1[6] , 
	\sa_count[19].r.part1[5] , \sa_count[19].r.part1[4] , 
	\sa_count[19].r.part1[3] , \sa_count[19].r.part1[2] , 
	\sa_count[19].r.part1[1] , \sa_count[19].r.part1[0] , 
	\sa_count[19].r.part0[31] , \sa_count[19].r.part0[30] , 
	\sa_count[19].r.part0[29] , \sa_count[19].r.part0[28] , 
	\sa_count[19].r.part0[27] , \sa_count[19].r.part0[26] , 
	\sa_count[19].r.part0[25] , \sa_count[19].r.part0[24] , 
	\sa_count[19].r.part0[23] , \sa_count[19].r.part0[22] , 
	\sa_count[19].r.part0[21] , \sa_count[19].r.part0[20] , 
	\sa_count[19].r.part0[19] , \sa_count[19].r.part0[18] , 
	\sa_count[19].r.part0[17] , \sa_count[19].r.part0[16] , 
	\sa_count[19].r.part0[15] , \sa_count[19].r.part0[14] , 
	\sa_count[19].r.part0[13] , \sa_count[19].r.part0[12] , 
	\sa_count[19].r.part0[11] , \sa_count[19].r.part0[10] , 
	\sa_count[19].r.part0[9] , \sa_count[19].r.part0[8] , 
	\sa_count[19].r.part0[7] , \sa_count[19].r.part0[6] , 
	\sa_count[19].r.part0[5] , \sa_count[19].r.part0[4] , 
	\sa_count[19].r.part0[3] , \sa_count[19].r.part0[2] , 
	\sa_count[19].r.part0[1] , \sa_count[19].r.part0[0] , 
	\sa_count[18].r.part1[31] , \sa_count[18].r.part1[30] , 
	\sa_count[18].r.part1[29] , \sa_count[18].r.part1[28] , 
	\sa_count[18].r.part1[27] , \sa_count[18].r.part1[26] , 
	\sa_count[18].r.part1[25] , \sa_count[18].r.part1[24] , 
	\sa_count[18].r.part1[23] , \sa_count[18].r.part1[22] , 
	\sa_count[18].r.part1[21] , \sa_count[18].r.part1[20] , 
	\sa_count[18].r.part1[19] , \sa_count[18].r.part1[18] , 
	\sa_count[18].r.part1[17] , \sa_count[18].r.part1[16] , 
	\sa_count[18].r.part1[15] , \sa_count[18].r.part1[14] , 
	\sa_count[18].r.part1[13] , \sa_count[18].r.part1[12] , 
	\sa_count[18].r.part1[11] , \sa_count[18].r.part1[10] , 
	\sa_count[18].r.part1[9] , \sa_count[18].r.part1[8] , 
	\sa_count[18].r.part1[7] , \sa_count[18].r.part1[6] , 
	\sa_count[18].r.part1[5] , \sa_count[18].r.part1[4] , 
	\sa_count[18].r.part1[3] , \sa_count[18].r.part1[2] , 
	\sa_count[18].r.part1[1] , \sa_count[18].r.part1[0] , 
	\sa_count[18].r.part0[31] , \sa_count[18].r.part0[30] , 
	\sa_count[18].r.part0[29] , \sa_count[18].r.part0[28] , 
	\sa_count[18].r.part0[27] , \sa_count[18].r.part0[26] , 
	\sa_count[18].r.part0[25] , \sa_count[18].r.part0[24] , 
	\sa_count[18].r.part0[23] , \sa_count[18].r.part0[22] , 
	\sa_count[18].r.part0[21] , \sa_count[18].r.part0[20] , 
	\sa_count[18].r.part0[19] , \sa_count[18].r.part0[18] , 
	\sa_count[18].r.part0[17] , \sa_count[18].r.part0[16] , 
	\sa_count[18].r.part0[15] , \sa_count[18].r.part0[14] , 
	\sa_count[18].r.part0[13] , \sa_count[18].r.part0[12] , 
	\sa_count[18].r.part0[11] , \sa_count[18].r.part0[10] , 
	\sa_count[18].r.part0[9] , \sa_count[18].r.part0[8] , 
	\sa_count[18].r.part0[7] , \sa_count[18].r.part0[6] , 
	\sa_count[18].r.part0[5] , \sa_count[18].r.part0[4] , 
	\sa_count[18].r.part0[3] , \sa_count[18].r.part0[2] , 
	\sa_count[18].r.part0[1] , \sa_count[18].r.part0[0] , 
	\sa_count[17].r.part1[31] , \sa_count[17].r.part1[30] , 
	\sa_count[17].r.part1[29] , \sa_count[17].r.part1[28] , 
	\sa_count[17].r.part1[27] , \sa_count[17].r.part1[26] , 
	\sa_count[17].r.part1[25] , \sa_count[17].r.part1[24] , 
	\sa_count[17].r.part1[23] , \sa_count[17].r.part1[22] , 
	\sa_count[17].r.part1[21] , \sa_count[17].r.part1[20] , 
	\sa_count[17].r.part1[19] , \sa_count[17].r.part1[18] , 
	\sa_count[17].r.part1[17] , \sa_count[17].r.part1[16] , 
	\sa_count[17].r.part1[15] , \sa_count[17].r.part1[14] , 
	\sa_count[17].r.part1[13] , \sa_count[17].r.part1[12] , 
	\sa_count[17].r.part1[11] , \sa_count[17].r.part1[10] , 
	\sa_count[17].r.part1[9] , \sa_count[17].r.part1[8] , 
	\sa_count[17].r.part1[7] , \sa_count[17].r.part1[6] , 
	\sa_count[17].r.part1[5] , \sa_count[17].r.part1[4] , 
	\sa_count[17].r.part1[3] , \sa_count[17].r.part1[2] , 
	\sa_count[17].r.part1[1] , \sa_count[17].r.part1[0] , 
	\sa_count[17].r.part0[31] , \sa_count[17].r.part0[30] , 
	\sa_count[17].r.part0[29] , \sa_count[17].r.part0[28] , 
	\sa_count[17].r.part0[27] , \sa_count[17].r.part0[26] , 
	\sa_count[17].r.part0[25] , \sa_count[17].r.part0[24] , 
	\sa_count[17].r.part0[23] , \sa_count[17].r.part0[22] , 
	\sa_count[17].r.part0[21] , \sa_count[17].r.part0[20] , 
	\sa_count[17].r.part0[19] , \sa_count[17].r.part0[18] , 
	\sa_count[17].r.part0[17] , \sa_count[17].r.part0[16] , 
	\sa_count[17].r.part0[15] , \sa_count[17].r.part0[14] , 
	\sa_count[17].r.part0[13] , \sa_count[17].r.part0[12] , 
	\sa_count[17].r.part0[11] , \sa_count[17].r.part0[10] , 
	\sa_count[17].r.part0[9] , \sa_count[17].r.part0[8] , 
	\sa_count[17].r.part0[7] , \sa_count[17].r.part0[6] , 
	\sa_count[17].r.part0[5] , \sa_count[17].r.part0[4] , 
	\sa_count[17].r.part0[3] , \sa_count[17].r.part0[2] , 
	\sa_count[17].r.part0[1] , \sa_count[17].r.part0[0] , 
	\sa_count[16].r.part1[31] , \sa_count[16].r.part1[30] , 
	\sa_count[16].r.part1[29] , \sa_count[16].r.part1[28] , 
	\sa_count[16].r.part1[27] , \sa_count[16].r.part1[26] , 
	\sa_count[16].r.part1[25] , \sa_count[16].r.part1[24] , 
	\sa_count[16].r.part1[23] , \sa_count[16].r.part1[22] , 
	\sa_count[16].r.part1[21] , \sa_count[16].r.part1[20] , 
	\sa_count[16].r.part1[19] , \sa_count[16].r.part1[18] , 
	\sa_count[16].r.part1[17] , \sa_count[16].r.part1[16] , 
	\sa_count[16].r.part1[15] , \sa_count[16].r.part1[14] , 
	\sa_count[16].r.part1[13] , \sa_count[16].r.part1[12] , 
	\sa_count[16].r.part1[11] , \sa_count[16].r.part1[10] , 
	\sa_count[16].r.part1[9] , \sa_count[16].r.part1[8] , 
	\sa_count[16].r.part1[7] , \sa_count[16].r.part1[6] , 
	\sa_count[16].r.part1[5] , \sa_count[16].r.part1[4] , 
	\sa_count[16].r.part1[3] , \sa_count[16].r.part1[2] , 
	\sa_count[16].r.part1[1] , \sa_count[16].r.part1[0] , 
	\sa_count[16].r.part0[31] , \sa_count[16].r.part0[30] , 
	\sa_count[16].r.part0[29] , \sa_count[16].r.part0[28] , 
	\sa_count[16].r.part0[27] , \sa_count[16].r.part0[26] , 
	\sa_count[16].r.part0[25] , \sa_count[16].r.part0[24] , 
	\sa_count[16].r.part0[23] , \sa_count[16].r.part0[22] , 
	\sa_count[16].r.part0[21] , \sa_count[16].r.part0[20] , 
	\sa_count[16].r.part0[19] , \sa_count[16].r.part0[18] , 
	\sa_count[16].r.part0[17] , \sa_count[16].r.part0[16] , 
	\sa_count[16].r.part0[15] , \sa_count[16].r.part0[14] , 
	\sa_count[16].r.part0[13] , \sa_count[16].r.part0[12] , 
	\sa_count[16].r.part0[11] , \sa_count[16].r.part0[10] , 
	\sa_count[16].r.part0[9] , \sa_count[16].r.part0[8] , 
	\sa_count[16].r.part0[7] , \sa_count[16].r.part0[6] , 
	\sa_count[16].r.part0[5] , \sa_count[16].r.part0[4] , 
	\sa_count[16].r.part0[3] , \sa_count[16].r.part0[2] , 
	\sa_count[16].r.part0[1] , \sa_count[16].r.part0[0] , 
	\sa_count[15].r.part1[31] , \sa_count[15].r.part1[30] , 
	\sa_count[15].r.part1[29] , \sa_count[15].r.part1[28] , 
	\sa_count[15].r.part1[27] , \sa_count[15].r.part1[26] , 
	\sa_count[15].r.part1[25] , \sa_count[15].r.part1[24] , 
	\sa_count[15].r.part1[23] , \sa_count[15].r.part1[22] , 
	\sa_count[15].r.part1[21] , \sa_count[15].r.part1[20] , 
	\sa_count[15].r.part1[19] , \sa_count[15].r.part1[18] , 
	\sa_count[15].r.part1[17] , \sa_count[15].r.part1[16] , 
	\sa_count[15].r.part1[15] , \sa_count[15].r.part1[14] , 
	\sa_count[15].r.part1[13] , \sa_count[15].r.part1[12] , 
	\sa_count[15].r.part1[11] , \sa_count[15].r.part1[10] , 
	\sa_count[15].r.part1[9] , \sa_count[15].r.part1[8] , 
	\sa_count[15].r.part1[7] , \sa_count[15].r.part1[6] , 
	\sa_count[15].r.part1[5] , \sa_count[15].r.part1[4] , 
	\sa_count[15].r.part1[3] , \sa_count[15].r.part1[2] , 
	\sa_count[15].r.part1[1] , \sa_count[15].r.part1[0] , 
	\sa_count[15].r.part0[31] , \sa_count[15].r.part0[30] , 
	\sa_count[15].r.part0[29] , \sa_count[15].r.part0[28] , 
	\sa_count[15].r.part0[27] , \sa_count[15].r.part0[26] , 
	\sa_count[15].r.part0[25] , \sa_count[15].r.part0[24] , 
	\sa_count[15].r.part0[23] , \sa_count[15].r.part0[22] , 
	\sa_count[15].r.part0[21] , \sa_count[15].r.part0[20] , 
	\sa_count[15].r.part0[19] , \sa_count[15].r.part0[18] , 
	\sa_count[15].r.part0[17] , \sa_count[15].r.part0[16] , 
	\sa_count[15].r.part0[15] , \sa_count[15].r.part0[14] , 
	\sa_count[15].r.part0[13] , \sa_count[15].r.part0[12] , 
	\sa_count[15].r.part0[11] , \sa_count[15].r.part0[10] , 
	\sa_count[15].r.part0[9] , \sa_count[15].r.part0[8] , 
	\sa_count[15].r.part0[7] , \sa_count[15].r.part0[6] , 
	\sa_count[15].r.part0[5] , \sa_count[15].r.part0[4] , 
	\sa_count[15].r.part0[3] , \sa_count[15].r.part0[2] , 
	\sa_count[15].r.part0[1] , \sa_count[15].r.part0[0] , 
	\sa_count[14].r.part1[31] , \sa_count[14].r.part1[30] , 
	\sa_count[14].r.part1[29] , \sa_count[14].r.part1[28] , 
	\sa_count[14].r.part1[27] , \sa_count[14].r.part1[26] , 
	\sa_count[14].r.part1[25] , \sa_count[14].r.part1[24] , 
	\sa_count[14].r.part1[23] , \sa_count[14].r.part1[22] , 
	\sa_count[14].r.part1[21] , \sa_count[14].r.part1[20] , 
	\sa_count[14].r.part1[19] , \sa_count[14].r.part1[18] , 
	\sa_count[14].r.part1[17] , \sa_count[14].r.part1[16] , 
	\sa_count[14].r.part1[15] , \sa_count[14].r.part1[14] , 
	\sa_count[14].r.part1[13] , \sa_count[14].r.part1[12] , 
	\sa_count[14].r.part1[11] , \sa_count[14].r.part1[10] , 
	\sa_count[14].r.part1[9] , \sa_count[14].r.part1[8] , 
	\sa_count[14].r.part1[7] , \sa_count[14].r.part1[6] , 
	\sa_count[14].r.part1[5] , \sa_count[14].r.part1[4] , 
	\sa_count[14].r.part1[3] , \sa_count[14].r.part1[2] , 
	\sa_count[14].r.part1[1] , \sa_count[14].r.part1[0] , 
	\sa_count[14].r.part0[31] , \sa_count[14].r.part0[30] , 
	\sa_count[14].r.part0[29] , \sa_count[14].r.part0[28] , 
	\sa_count[14].r.part0[27] , \sa_count[14].r.part0[26] , 
	\sa_count[14].r.part0[25] , \sa_count[14].r.part0[24] , 
	\sa_count[14].r.part0[23] , \sa_count[14].r.part0[22] , 
	\sa_count[14].r.part0[21] , \sa_count[14].r.part0[20] , 
	\sa_count[14].r.part0[19] , \sa_count[14].r.part0[18] , 
	\sa_count[14].r.part0[17] , \sa_count[14].r.part0[16] , 
	\sa_count[14].r.part0[15] , \sa_count[14].r.part0[14] , 
	\sa_count[14].r.part0[13] , \sa_count[14].r.part0[12] , 
	\sa_count[14].r.part0[11] , \sa_count[14].r.part0[10] , 
	\sa_count[14].r.part0[9] , \sa_count[14].r.part0[8] , 
	\sa_count[14].r.part0[7] , \sa_count[14].r.part0[6] , 
	\sa_count[14].r.part0[5] , \sa_count[14].r.part0[4] , 
	\sa_count[14].r.part0[3] , \sa_count[14].r.part0[2] , 
	\sa_count[14].r.part0[1] , \sa_count[14].r.part0[0] , 
	\sa_count[13].r.part1[31] , \sa_count[13].r.part1[30] , 
	\sa_count[13].r.part1[29] , \sa_count[13].r.part1[28] , 
	\sa_count[13].r.part1[27] , \sa_count[13].r.part1[26] , 
	\sa_count[13].r.part1[25] , \sa_count[13].r.part1[24] , 
	\sa_count[13].r.part1[23] , \sa_count[13].r.part1[22] , 
	\sa_count[13].r.part1[21] , \sa_count[13].r.part1[20] , 
	\sa_count[13].r.part1[19] , \sa_count[13].r.part1[18] , 
	\sa_count[13].r.part1[17] , \sa_count[13].r.part1[16] , 
	\sa_count[13].r.part1[15] , \sa_count[13].r.part1[14] , 
	\sa_count[13].r.part1[13] , \sa_count[13].r.part1[12] , 
	\sa_count[13].r.part1[11] , \sa_count[13].r.part1[10] , 
	\sa_count[13].r.part1[9] , \sa_count[13].r.part1[8] , 
	\sa_count[13].r.part1[7] , \sa_count[13].r.part1[6] , 
	\sa_count[13].r.part1[5] , \sa_count[13].r.part1[4] , 
	\sa_count[13].r.part1[3] , \sa_count[13].r.part1[2] , 
	\sa_count[13].r.part1[1] , \sa_count[13].r.part1[0] , 
	\sa_count[13].r.part0[31] , \sa_count[13].r.part0[30] , 
	\sa_count[13].r.part0[29] , \sa_count[13].r.part0[28] , 
	\sa_count[13].r.part0[27] , \sa_count[13].r.part0[26] , 
	\sa_count[13].r.part0[25] , \sa_count[13].r.part0[24] , 
	\sa_count[13].r.part0[23] , \sa_count[13].r.part0[22] , 
	\sa_count[13].r.part0[21] , \sa_count[13].r.part0[20] , 
	\sa_count[13].r.part0[19] , \sa_count[13].r.part0[18] , 
	\sa_count[13].r.part0[17] , \sa_count[13].r.part0[16] , 
	\sa_count[13].r.part0[15] , \sa_count[13].r.part0[14] , 
	\sa_count[13].r.part0[13] , \sa_count[13].r.part0[12] , 
	\sa_count[13].r.part0[11] , \sa_count[13].r.part0[10] , 
	\sa_count[13].r.part0[9] , \sa_count[13].r.part0[8] , 
	\sa_count[13].r.part0[7] , \sa_count[13].r.part0[6] , 
	\sa_count[13].r.part0[5] , \sa_count[13].r.part0[4] , 
	\sa_count[13].r.part0[3] , \sa_count[13].r.part0[2] , 
	\sa_count[13].r.part0[1] , \sa_count[13].r.part0[0] , 
	\sa_count[12].r.part1[31] , \sa_count[12].r.part1[30] , 
	\sa_count[12].r.part1[29] , \sa_count[12].r.part1[28] , 
	\sa_count[12].r.part1[27] , \sa_count[12].r.part1[26] , 
	\sa_count[12].r.part1[25] , \sa_count[12].r.part1[24] , 
	\sa_count[12].r.part1[23] , \sa_count[12].r.part1[22] , 
	\sa_count[12].r.part1[21] , \sa_count[12].r.part1[20] , 
	\sa_count[12].r.part1[19] , \sa_count[12].r.part1[18] , 
	\sa_count[12].r.part1[17] , \sa_count[12].r.part1[16] , 
	\sa_count[12].r.part1[15] , \sa_count[12].r.part1[14] , 
	\sa_count[12].r.part1[13] , \sa_count[12].r.part1[12] , 
	\sa_count[12].r.part1[11] , \sa_count[12].r.part1[10] , 
	\sa_count[12].r.part1[9] , \sa_count[12].r.part1[8] , 
	\sa_count[12].r.part1[7] , \sa_count[12].r.part1[6] , 
	\sa_count[12].r.part1[5] , \sa_count[12].r.part1[4] , 
	\sa_count[12].r.part1[3] , \sa_count[12].r.part1[2] , 
	\sa_count[12].r.part1[1] , \sa_count[12].r.part1[0] , 
	\sa_count[12].r.part0[31] , \sa_count[12].r.part0[30] , 
	\sa_count[12].r.part0[29] , \sa_count[12].r.part0[28] , 
	\sa_count[12].r.part0[27] , \sa_count[12].r.part0[26] , 
	\sa_count[12].r.part0[25] , \sa_count[12].r.part0[24] , 
	\sa_count[12].r.part0[23] , \sa_count[12].r.part0[22] , 
	\sa_count[12].r.part0[21] , \sa_count[12].r.part0[20] , 
	\sa_count[12].r.part0[19] , \sa_count[12].r.part0[18] , 
	\sa_count[12].r.part0[17] , \sa_count[12].r.part0[16] , 
	\sa_count[12].r.part0[15] , \sa_count[12].r.part0[14] , 
	\sa_count[12].r.part0[13] , \sa_count[12].r.part0[12] , 
	\sa_count[12].r.part0[11] , \sa_count[12].r.part0[10] , 
	\sa_count[12].r.part0[9] , \sa_count[12].r.part0[8] , 
	\sa_count[12].r.part0[7] , \sa_count[12].r.part0[6] , 
	\sa_count[12].r.part0[5] , \sa_count[12].r.part0[4] , 
	\sa_count[12].r.part0[3] , \sa_count[12].r.part0[2] , 
	\sa_count[12].r.part0[1] , \sa_count[12].r.part0[0] , 
	\sa_count[11].r.part1[31] , \sa_count[11].r.part1[30] , 
	\sa_count[11].r.part1[29] , \sa_count[11].r.part1[28] , 
	\sa_count[11].r.part1[27] , \sa_count[11].r.part1[26] , 
	\sa_count[11].r.part1[25] , \sa_count[11].r.part1[24] , 
	\sa_count[11].r.part1[23] , \sa_count[11].r.part1[22] , 
	\sa_count[11].r.part1[21] , \sa_count[11].r.part1[20] , 
	\sa_count[11].r.part1[19] , \sa_count[11].r.part1[18] , 
	\sa_count[11].r.part1[17] , \sa_count[11].r.part1[16] , 
	\sa_count[11].r.part1[15] , \sa_count[11].r.part1[14] , 
	\sa_count[11].r.part1[13] , \sa_count[11].r.part1[12] , 
	\sa_count[11].r.part1[11] , \sa_count[11].r.part1[10] , 
	\sa_count[11].r.part1[9] , \sa_count[11].r.part1[8] , 
	\sa_count[11].r.part1[7] , \sa_count[11].r.part1[6] , 
	\sa_count[11].r.part1[5] , \sa_count[11].r.part1[4] , 
	\sa_count[11].r.part1[3] , \sa_count[11].r.part1[2] , 
	\sa_count[11].r.part1[1] , \sa_count[11].r.part1[0] , 
	\sa_count[11].r.part0[31] , \sa_count[11].r.part0[30] , 
	\sa_count[11].r.part0[29] , \sa_count[11].r.part0[28] , 
	\sa_count[11].r.part0[27] , \sa_count[11].r.part0[26] , 
	\sa_count[11].r.part0[25] , \sa_count[11].r.part0[24] , 
	\sa_count[11].r.part0[23] , \sa_count[11].r.part0[22] , 
	\sa_count[11].r.part0[21] , \sa_count[11].r.part0[20] , 
	\sa_count[11].r.part0[19] , \sa_count[11].r.part0[18] , 
	\sa_count[11].r.part0[17] , \sa_count[11].r.part0[16] , 
	\sa_count[11].r.part0[15] , \sa_count[11].r.part0[14] , 
	\sa_count[11].r.part0[13] , \sa_count[11].r.part0[12] , 
	\sa_count[11].r.part0[11] , \sa_count[11].r.part0[10] , 
	\sa_count[11].r.part0[9] , \sa_count[11].r.part0[8] , 
	\sa_count[11].r.part0[7] , \sa_count[11].r.part0[6] , 
	\sa_count[11].r.part0[5] , \sa_count[11].r.part0[4] , 
	\sa_count[11].r.part0[3] , \sa_count[11].r.part0[2] , 
	\sa_count[11].r.part0[1] , \sa_count[11].r.part0[0] , 
	\sa_count[10].r.part1[31] , \sa_count[10].r.part1[30] , 
	\sa_count[10].r.part1[29] , \sa_count[10].r.part1[28] , 
	\sa_count[10].r.part1[27] , \sa_count[10].r.part1[26] , 
	\sa_count[10].r.part1[25] , \sa_count[10].r.part1[24] , 
	\sa_count[10].r.part1[23] , \sa_count[10].r.part1[22] , 
	\sa_count[10].r.part1[21] , \sa_count[10].r.part1[20] , 
	\sa_count[10].r.part1[19] , \sa_count[10].r.part1[18] , 
	\sa_count[10].r.part1[17] , \sa_count[10].r.part1[16] , 
	\sa_count[10].r.part1[15] , \sa_count[10].r.part1[14] , 
	\sa_count[10].r.part1[13] , \sa_count[10].r.part1[12] , 
	\sa_count[10].r.part1[11] , \sa_count[10].r.part1[10] , 
	\sa_count[10].r.part1[9] , \sa_count[10].r.part1[8] , 
	\sa_count[10].r.part1[7] , \sa_count[10].r.part1[6] , 
	\sa_count[10].r.part1[5] , \sa_count[10].r.part1[4] , 
	\sa_count[10].r.part1[3] , \sa_count[10].r.part1[2] , 
	\sa_count[10].r.part1[1] , \sa_count[10].r.part1[0] , 
	\sa_count[10].r.part0[31] , \sa_count[10].r.part0[30] , 
	\sa_count[10].r.part0[29] , \sa_count[10].r.part0[28] , 
	\sa_count[10].r.part0[27] , \sa_count[10].r.part0[26] , 
	\sa_count[10].r.part0[25] , \sa_count[10].r.part0[24] , 
	\sa_count[10].r.part0[23] , \sa_count[10].r.part0[22] , 
	\sa_count[10].r.part0[21] , \sa_count[10].r.part0[20] , 
	\sa_count[10].r.part0[19] , \sa_count[10].r.part0[18] , 
	\sa_count[10].r.part0[17] , \sa_count[10].r.part0[16] , 
	\sa_count[10].r.part0[15] , \sa_count[10].r.part0[14] , 
	\sa_count[10].r.part0[13] , \sa_count[10].r.part0[12] , 
	\sa_count[10].r.part0[11] , \sa_count[10].r.part0[10] , 
	\sa_count[10].r.part0[9] , \sa_count[10].r.part0[8] , 
	\sa_count[10].r.part0[7] , \sa_count[10].r.part0[6] , 
	\sa_count[10].r.part0[5] , \sa_count[10].r.part0[4] , 
	\sa_count[10].r.part0[3] , \sa_count[10].r.part0[2] , 
	\sa_count[10].r.part0[1] , \sa_count[10].r.part0[0] , 
	\sa_count[9].r.part1[31] , \sa_count[9].r.part1[30] , 
	\sa_count[9].r.part1[29] , \sa_count[9].r.part1[28] , 
	\sa_count[9].r.part1[27] , \sa_count[9].r.part1[26] , 
	\sa_count[9].r.part1[25] , \sa_count[9].r.part1[24] , 
	\sa_count[9].r.part1[23] , \sa_count[9].r.part1[22] , 
	\sa_count[9].r.part1[21] , \sa_count[9].r.part1[20] , 
	\sa_count[9].r.part1[19] , \sa_count[9].r.part1[18] , 
	\sa_count[9].r.part1[17] , \sa_count[9].r.part1[16] , 
	\sa_count[9].r.part1[15] , \sa_count[9].r.part1[14] , 
	\sa_count[9].r.part1[13] , \sa_count[9].r.part1[12] , 
	\sa_count[9].r.part1[11] , \sa_count[9].r.part1[10] , 
	\sa_count[9].r.part1[9] , \sa_count[9].r.part1[8] , 
	\sa_count[9].r.part1[7] , \sa_count[9].r.part1[6] , 
	\sa_count[9].r.part1[5] , \sa_count[9].r.part1[4] , 
	\sa_count[9].r.part1[3] , \sa_count[9].r.part1[2] , 
	\sa_count[9].r.part1[1] , \sa_count[9].r.part1[0] , 
	\sa_count[9].r.part0[31] , \sa_count[9].r.part0[30] , 
	\sa_count[9].r.part0[29] , \sa_count[9].r.part0[28] , 
	\sa_count[9].r.part0[27] , \sa_count[9].r.part0[26] , 
	\sa_count[9].r.part0[25] , \sa_count[9].r.part0[24] , 
	\sa_count[9].r.part0[23] , \sa_count[9].r.part0[22] , 
	\sa_count[9].r.part0[21] , \sa_count[9].r.part0[20] , 
	\sa_count[9].r.part0[19] , \sa_count[9].r.part0[18] , 
	\sa_count[9].r.part0[17] , \sa_count[9].r.part0[16] , 
	\sa_count[9].r.part0[15] , \sa_count[9].r.part0[14] , 
	\sa_count[9].r.part0[13] , \sa_count[9].r.part0[12] , 
	\sa_count[9].r.part0[11] , \sa_count[9].r.part0[10] , 
	\sa_count[9].r.part0[9] , \sa_count[9].r.part0[8] , 
	\sa_count[9].r.part0[7] , \sa_count[9].r.part0[6] , 
	\sa_count[9].r.part0[5] , \sa_count[9].r.part0[4] , 
	\sa_count[9].r.part0[3] , \sa_count[9].r.part0[2] , 
	\sa_count[9].r.part0[1] , \sa_count[9].r.part0[0] , 
	\sa_count[8].r.part1[31] , \sa_count[8].r.part1[30] , 
	\sa_count[8].r.part1[29] , \sa_count[8].r.part1[28] , 
	\sa_count[8].r.part1[27] , \sa_count[8].r.part1[26] , 
	\sa_count[8].r.part1[25] , \sa_count[8].r.part1[24] , 
	\sa_count[8].r.part1[23] , \sa_count[8].r.part1[22] , 
	\sa_count[8].r.part1[21] , \sa_count[8].r.part1[20] , 
	\sa_count[8].r.part1[19] , \sa_count[8].r.part1[18] , 
	\sa_count[8].r.part1[17] , \sa_count[8].r.part1[16] , 
	\sa_count[8].r.part1[15] , \sa_count[8].r.part1[14] , 
	\sa_count[8].r.part1[13] , \sa_count[8].r.part1[12] , 
	\sa_count[8].r.part1[11] , \sa_count[8].r.part1[10] , 
	\sa_count[8].r.part1[9] , \sa_count[8].r.part1[8] , 
	\sa_count[8].r.part1[7] , \sa_count[8].r.part1[6] , 
	\sa_count[8].r.part1[5] , \sa_count[8].r.part1[4] , 
	\sa_count[8].r.part1[3] , \sa_count[8].r.part1[2] , 
	\sa_count[8].r.part1[1] , \sa_count[8].r.part1[0] , 
	\sa_count[8].r.part0[31] , \sa_count[8].r.part0[30] , 
	\sa_count[8].r.part0[29] , \sa_count[8].r.part0[28] , 
	\sa_count[8].r.part0[27] , \sa_count[8].r.part0[26] , 
	\sa_count[8].r.part0[25] , \sa_count[8].r.part0[24] , 
	\sa_count[8].r.part0[23] , \sa_count[8].r.part0[22] , 
	\sa_count[8].r.part0[21] , \sa_count[8].r.part0[20] , 
	\sa_count[8].r.part0[19] , \sa_count[8].r.part0[18] , 
	\sa_count[8].r.part0[17] , \sa_count[8].r.part0[16] , 
	\sa_count[8].r.part0[15] , \sa_count[8].r.part0[14] , 
	\sa_count[8].r.part0[13] , \sa_count[8].r.part0[12] , 
	\sa_count[8].r.part0[11] , \sa_count[8].r.part0[10] , 
	\sa_count[8].r.part0[9] , \sa_count[8].r.part0[8] , 
	\sa_count[8].r.part0[7] , \sa_count[8].r.part0[6] , 
	\sa_count[8].r.part0[5] , \sa_count[8].r.part0[4] , 
	\sa_count[8].r.part0[3] , \sa_count[8].r.part0[2] , 
	\sa_count[8].r.part0[1] , \sa_count[8].r.part0[0] , 
	\sa_count[7].r.part1[31] , \sa_count[7].r.part1[30] , 
	\sa_count[7].r.part1[29] , \sa_count[7].r.part1[28] , 
	\sa_count[7].r.part1[27] , \sa_count[7].r.part1[26] , 
	\sa_count[7].r.part1[25] , \sa_count[7].r.part1[24] , 
	\sa_count[7].r.part1[23] , \sa_count[7].r.part1[22] , 
	\sa_count[7].r.part1[21] , \sa_count[7].r.part1[20] , 
	\sa_count[7].r.part1[19] , \sa_count[7].r.part1[18] , 
	\sa_count[7].r.part1[17] , \sa_count[7].r.part1[16] , 
	\sa_count[7].r.part1[15] , \sa_count[7].r.part1[14] , 
	\sa_count[7].r.part1[13] , \sa_count[7].r.part1[12] , 
	\sa_count[7].r.part1[11] , \sa_count[7].r.part1[10] , 
	\sa_count[7].r.part1[9] , \sa_count[7].r.part1[8] , 
	\sa_count[7].r.part1[7] , \sa_count[7].r.part1[6] , 
	\sa_count[7].r.part1[5] , \sa_count[7].r.part1[4] , 
	\sa_count[7].r.part1[3] , \sa_count[7].r.part1[2] , 
	\sa_count[7].r.part1[1] , \sa_count[7].r.part1[0] , 
	\sa_count[7].r.part0[31] , \sa_count[7].r.part0[30] , 
	\sa_count[7].r.part0[29] , \sa_count[7].r.part0[28] , 
	\sa_count[7].r.part0[27] , \sa_count[7].r.part0[26] , 
	\sa_count[7].r.part0[25] , \sa_count[7].r.part0[24] , 
	\sa_count[7].r.part0[23] , \sa_count[7].r.part0[22] , 
	\sa_count[7].r.part0[21] , \sa_count[7].r.part0[20] , 
	\sa_count[7].r.part0[19] , \sa_count[7].r.part0[18] , 
	\sa_count[7].r.part0[17] , \sa_count[7].r.part0[16] , 
	\sa_count[7].r.part0[15] , \sa_count[7].r.part0[14] , 
	\sa_count[7].r.part0[13] , \sa_count[7].r.part0[12] , 
	\sa_count[7].r.part0[11] , \sa_count[7].r.part0[10] , 
	\sa_count[7].r.part0[9] , \sa_count[7].r.part0[8] , 
	\sa_count[7].r.part0[7] , \sa_count[7].r.part0[6] , 
	\sa_count[7].r.part0[5] , \sa_count[7].r.part0[4] , 
	\sa_count[7].r.part0[3] , \sa_count[7].r.part0[2] , 
	\sa_count[7].r.part0[1] , \sa_count[7].r.part0[0] , 
	\sa_count[6].r.part1[31] , \sa_count[6].r.part1[30] , 
	\sa_count[6].r.part1[29] , \sa_count[6].r.part1[28] , 
	\sa_count[6].r.part1[27] , \sa_count[6].r.part1[26] , 
	\sa_count[6].r.part1[25] , \sa_count[6].r.part1[24] , 
	\sa_count[6].r.part1[23] , \sa_count[6].r.part1[22] , 
	\sa_count[6].r.part1[21] , \sa_count[6].r.part1[20] , 
	\sa_count[6].r.part1[19] , \sa_count[6].r.part1[18] , 
	\sa_count[6].r.part1[17] , \sa_count[6].r.part1[16] , 
	\sa_count[6].r.part1[15] , \sa_count[6].r.part1[14] , 
	\sa_count[6].r.part1[13] , \sa_count[6].r.part1[12] , 
	\sa_count[6].r.part1[11] , \sa_count[6].r.part1[10] , 
	\sa_count[6].r.part1[9] , \sa_count[6].r.part1[8] , 
	\sa_count[6].r.part1[7] , \sa_count[6].r.part1[6] , 
	\sa_count[6].r.part1[5] , \sa_count[6].r.part1[4] , 
	\sa_count[6].r.part1[3] , \sa_count[6].r.part1[2] , 
	\sa_count[6].r.part1[1] , \sa_count[6].r.part1[0] , 
	\sa_count[6].r.part0[31] , \sa_count[6].r.part0[30] , 
	\sa_count[6].r.part0[29] , \sa_count[6].r.part0[28] , 
	\sa_count[6].r.part0[27] , \sa_count[6].r.part0[26] , 
	\sa_count[6].r.part0[25] , \sa_count[6].r.part0[24] , 
	\sa_count[6].r.part0[23] , \sa_count[6].r.part0[22] , 
	\sa_count[6].r.part0[21] , \sa_count[6].r.part0[20] , 
	\sa_count[6].r.part0[19] , \sa_count[6].r.part0[18] , 
	\sa_count[6].r.part0[17] , \sa_count[6].r.part0[16] , 
	\sa_count[6].r.part0[15] , \sa_count[6].r.part0[14] , 
	\sa_count[6].r.part0[13] , \sa_count[6].r.part0[12] , 
	\sa_count[6].r.part0[11] , \sa_count[6].r.part0[10] , 
	\sa_count[6].r.part0[9] , \sa_count[6].r.part0[8] , 
	\sa_count[6].r.part0[7] , \sa_count[6].r.part0[6] , 
	\sa_count[6].r.part0[5] , \sa_count[6].r.part0[4] , 
	\sa_count[6].r.part0[3] , \sa_count[6].r.part0[2] , 
	\sa_count[6].r.part0[1] , \sa_count[6].r.part0[0] , 
	\sa_count[5].r.part1[31] , \sa_count[5].r.part1[30] , 
	\sa_count[5].r.part1[29] , \sa_count[5].r.part1[28] , 
	\sa_count[5].r.part1[27] , \sa_count[5].r.part1[26] , 
	\sa_count[5].r.part1[25] , \sa_count[5].r.part1[24] , 
	\sa_count[5].r.part1[23] , \sa_count[5].r.part1[22] , 
	\sa_count[5].r.part1[21] , \sa_count[5].r.part1[20] , 
	\sa_count[5].r.part1[19] , \sa_count[5].r.part1[18] , 
	\sa_count[5].r.part1[17] , \sa_count[5].r.part1[16] , 
	\sa_count[5].r.part1[15] , \sa_count[5].r.part1[14] , 
	\sa_count[5].r.part1[13] , \sa_count[5].r.part1[12] , 
	\sa_count[5].r.part1[11] , \sa_count[5].r.part1[10] , 
	\sa_count[5].r.part1[9] , \sa_count[5].r.part1[8] , 
	\sa_count[5].r.part1[7] , \sa_count[5].r.part1[6] , 
	\sa_count[5].r.part1[5] , \sa_count[5].r.part1[4] , 
	\sa_count[5].r.part1[3] , \sa_count[5].r.part1[2] , 
	\sa_count[5].r.part1[1] , \sa_count[5].r.part1[0] , 
	\sa_count[5].r.part0[31] , \sa_count[5].r.part0[30] , 
	\sa_count[5].r.part0[29] , \sa_count[5].r.part0[28] , 
	\sa_count[5].r.part0[27] , \sa_count[5].r.part0[26] , 
	\sa_count[5].r.part0[25] , \sa_count[5].r.part0[24] , 
	\sa_count[5].r.part0[23] , \sa_count[5].r.part0[22] , 
	\sa_count[5].r.part0[21] , \sa_count[5].r.part0[20] , 
	\sa_count[5].r.part0[19] , \sa_count[5].r.part0[18] , 
	\sa_count[5].r.part0[17] , \sa_count[5].r.part0[16] , 
	\sa_count[5].r.part0[15] , \sa_count[5].r.part0[14] , 
	\sa_count[5].r.part0[13] , \sa_count[5].r.part0[12] , 
	\sa_count[5].r.part0[11] , \sa_count[5].r.part0[10] , 
	\sa_count[5].r.part0[9] , \sa_count[5].r.part0[8] , 
	\sa_count[5].r.part0[7] , \sa_count[5].r.part0[6] , 
	\sa_count[5].r.part0[5] , \sa_count[5].r.part0[4] , 
	\sa_count[5].r.part0[3] , \sa_count[5].r.part0[2] , 
	\sa_count[5].r.part0[1] , \sa_count[5].r.part0[0] , 
	\sa_count[4].r.part1[31] , \sa_count[4].r.part1[30] , 
	\sa_count[4].r.part1[29] , \sa_count[4].r.part1[28] , 
	\sa_count[4].r.part1[27] , \sa_count[4].r.part1[26] , 
	\sa_count[4].r.part1[25] , \sa_count[4].r.part1[24] , 
	\sa_count[4].r.part1[23] , \sa_count[4].r.part1[22] , 
	\sa_count[4].r.part1[21] , \sa_count[4].r.part1[20] , 
	\sa_count[4].r.part1[19] , \sa_count[4].r.part1[18] , 
	\sa_count[4].r.part1[17] , \sa_count[4].r.part1[16] , 
	\sa_count[4].r.part1[15] , \sa_count[4].r.part1[14] , 
	\sa_count[4].r.part1[13] , \sa_count[4].r.part1[12] , 
	\sa_count[4].r.part1[11] , \sa_count[4].r.part1[10] , 
	\sa_count[4].r.part1[9] , \sa_count[4].r.part1[8] , 
	\sa_count[4].r.part1[7] , \sa_count[4].r.part1[6] , 
	\sa_count[4].r.part1[5] , \sa_count[4].r.part1[4] , 
	\sa_count[4].r.part1[3] , \sa_count[4].r.part1[2] , 
	\sa_count[4].r.part1[1] , \sa_count[4].r.part1[0] , 
	\sa_count[4].r.part0[31] , \sa_count[4].r.part0[30] , 
	\sa_count[4].r.part0[29] , \sa_count[4].r.part0[28] , 
	\sa_count[4].r.part0[27] , \sa_count[4].r.part0[26] , 
	\sa_count[4].r.part0[25] , \sa_count[4].r.part0[24] , 
	\sa_count[4].r.part0[23] , \sa_count[4].r.part0[22] , 
	\sa_count[4].r.part0[21] , \sa_count[4].r.part0[20] , 
	\sa_count[4].r.part0[19] , \sa_count[4].r.part0[18] , 
	\sa_count[4].r.part0[17] , \sa_count[4].r.part0[16] , 
	\sa_count[4].r.part0[15] , \sa_count[4].r.part0[14] , 
	\sa_count[4].r.part0[13] , \sa_count[4].r.part0[12] , 
	\sa_count[4].r.part0[11] , \sa_count[4].r.part0[10] , 
	\sa_count[4].r.part0[9] , \sa_count[4].r.part0[8] , 
	\sa_count[4].r.part0[7] , \sa_count[4].r.part0[6] , 
	\sa_count[4].r.part0[5] , \sa_count[4].r.part0[4] , 
	\sa_count[4].r.part0[3] , \sa_count[4].r.part0[2] , 
	\sa_count[4].r.part0[1] , \sa_count[4].r.part0[0] , 
	\sa_count[3].r.part1[31] , \sa_count[3].r.part1[30] , 
	\sa_count[3].r.part1[29] , \sa_count[3].r.part1[28] , 
	\sa_count[3].r.part1[27] , \sa_count[3].r.part1[26] , 
	\sa_count[3].r.part1[25] , \sa_count[3].r.part1[24] , 
	\sa_count[3].r.part1[23] , \sa_count[3].r.part1[22] , 
	\sa_count[3].r.part1[21] , \sa_count[3].r.part1[20] , 
	\sa_count[3].r.part1[19] , \sa_count[3].r.part1[18] , 
	\sa_count[3].r.part1[17] , \sa_count[3].r.part1[16] , 
	\sa_count[3].r.part1[15] , \sa_count[3].r.part1[14] , 
	\sa_count[3].r.part1[13] , \sa_count[3].r.part1[12] , 
	\sa_count[3].r.part1[11] , \sa_count[3].r.part1[10] , 
	\sa_count[3].r.part1[9] , \sa_count[3].r.part1[8] , 
	\sa_count[3].r.part1[7] , \sa_count[3].r.part1[6] , 
	\sa_count[3].r.part1[5] , \sa_count[3].r.part1[4] , 
	\sa_count[3].r.part1[3] , \sa_count[3].r.part1[2] , 
	\sa_count[3].r.part1[1] , \sa_count[3].r.part1[0] , 
	\sa_count[3].r.part0[31] , \sa_count[3].r.part0[30] , 
	\sa_count[3].r.part0[29] , \sa_count[3].r.part0[28] , 
	\sa_count[3].r.part0[27] , \sa_count[3].r.part0[26] , 
	\sa_count[3].r.part0[25] , \sa_count[3].r.part0[24] , 
	\sa_count[3].r.part0[23] , \sa_count[3].r.part0[22] , 
	\sa_count[3].r.part0[21] , \sa_count[3].r.part0[20] , 
	\sa_count[3].r.part0[19] , \sa_count[3].r.part0[18] , 
	\sa_count[3].r.part0[17] , \sa_count[3].r.part0[16] , 
	\sa_count[3].r.part0[15] , \sa_count[3].r.part0[14] , 
	\sa_count[3].r.part0[13] , \sa_count[3].r.part0[12] , 
	\sa_count[3].r.part0[11] , \sa_count[3].r.part0[10] , 
	\sa_count[3].r.part0[9] , \sa_count[3].r.part0[8] , 
	\sa_count[3].r.part0[7] , \sa_count[3].r.part0[6] , 
	\sa_count[3].r.part0[5] , \sa_count[3].r.part0[4] , 
	\sa_count[3].r.part0[3] , \sa_count[3].r.part0[2] , 
	\sa_count[3].r.part0[1] , \sa_count[3].r.part0[0] , 
	\sa_count[2].r.part1[31] , \sa_count[2].r.part1[30] , 
	\sa_count[2].r.part1[29] , \sa_count[2].r.part1[28] , 
	\sa_count[2].r.part1[27] , \sa_count[2].r.part1[26] , 
	\sa_count[2].r.part1[25] , \sa_count[2].r.part1[24] , 
	\sa_count[2].r.part1[23] , \sa_count[2].r.part1[22] , 
	\sa_count[2].r.part1[21] , \sa_count[2].r.part1[20] , 
	\sa_count[2].r.part1[19] , \sa_count[2].r.part1[18] , 
	\sa_count[2].r.part1[17] , \sa_count[2].r.part1[16] , 
	\sa_count[2].r.part1[15] , \sa_count[2].r.part1[14] , 
	\sa_count[2].r.part1[13] , \sa_count[2].r.part1[12] , 
	\sa_count[2].r.part1[11] , \sa_count[2].r.part1[10] , 
	\sa_count[2].r.part1[9] , \sa_count[2].r.part1[8] , 
	\sa_count[2].r.part1[7] , \sa_count[2].r.part1[6] , 
	\sa_count[2].r.part1[5] , \sa_count[2].r.part1[4] , 
	\sa_count[2].r.part1[3] , \sa_count[2].r.part1[2] , 
	\sa_count[2].r.part1[1] , \sa_count[2].r.part1[0] , 
	\sa_count[2].r.part0[31] , \sa_count[2].r.part0[30] , 
	\sa_count[2].r.part0[29] , \sa_count[2].r.part0[28] , 
	\sa_count[2].r.part0[27] , \sa_count[2].r.part0[26] , 
	\sa_count[2].r.part0[25] , \sa_count[2].r.part0[24] , 
	\sa_count[2].r.part0[23] , \sa_count[2].r.part0[22] , 
	\sa_count[2].r.part0[21] , \sa_count[2].r.part0[20] , 
	\sa_count[2].r.part0[19] , \sa_count[2].r.part0[18] , 
	\sa_count[2].r.part0[17] , \sa_count[2].r.part0[16] , 
	\sa_count[2].r.part0[15] , \sa_count[2].r.part0[14] , 
	\sa_count[2].r.part0[13] , \sa_count[2].r.part0[12] , 
	\sa_count[2].r.part0[11] , \sa_count[2].r.part0[10] , 
	\sa_count[2].r.part0[9] , \sa_count[2].r.part0[8] , 
	\sa_count[2].r.part0[7] , \sa_count[2].r.part0[6] , 
	\sa_count[2].r.part0[5] , \sa_count[2].r.part0[4] , 
	\sa_count[2].r.part0[3] , \sa_count[2].r.part0[2] , 
	\sa_count[2].r.part0[1] , \sa_count[2].r.part0[0] , 
	\sa_count[1].r.part1[31] , \sa_count[1].r.part1[30] , 
	\sa_count[1].r.part1[29] , \sa_count[1].r.part1[28] , 
	\sa_count[1].r.part1[27] , \sa_count[1].r.part1[26] , 
	\sa_count[1].r.part1[25] , \sa_count[1].r.part1[24] , 
	\sa_count[1].r.part1[23] , \sa_count[1].r.part1[22] , 
	\sa_count[1].r.part1[21] , \sa_count[1].r.part1[20] , 
	\sa_count[1].r.part1[19] , \sa_count[1].r.part1[18] , 
	\sa_count[1].r.part1[17] , \sa_count[1].r.part1[16] , 
	\sa_count[1].r.part1[15] , \sa_count[1].r.part1[14] , 
	\sa_count[1].r.part1[13] , \sa_count[1].r.part1[12] , 
	\sa_count[1].r.part1[11] , \sa_count[1].r.part1[10] , 
	\sa_count[1].r.part1[9] , \sa_count[1].r.part1[8] , 
	\sa_count[1].r.part1[7] , \sa_count[1].r.part1[6] , 
	\sa_count[1].r.part1[5] , \sa_count[1].r.part1[4] , 
	\sa_count[1].r.part1[3] , \sa_count[1].r.part1[2] , 
	\sa_count[1].r.part1[1] , \sa_count[1].r.part1[0] , 
	\sa_count[1].r.part0[31] , \sa_count[1].r.part0[30] , 
	\sa_count[1].r.part0[29] , \sa_count[1].r.part0[28] , 
	\sa_count[1].r.part0[27] , \sa_count[1].r.part0[26] , 
	\sa_count[1].r.part0[25] , \sa_count[1].r.part0[24] , 
	\sa_count[1].r.part0[23] , \sa_count[1].r.part0[22] , 
	\sa_count[1].r.part0[21] , \sa_count[1].r.part0[20] , 
	\sa_count[1].r.part0[19] , \sa_count[1].r.part0[18] , 
	\sa_count[1].r.part0[17] , \sa_count[1].r.part0[16] , 
	\sa_count[1].r.part0[15] , \sa_count[1].r.part0[14] , 
	\sa_count[1].r.part0[13] , \sa_count[1].r.part0[12] , 
	\sa_count[1].r.part0[11] , \sa_count[1].r.part0[10] , 
	\sa_count[1].r.part0[9] , \sa_count[1].r.part0[8] , 
	\sa_count[1].r.part0[7] , \sa_count[1].r.part0[6] , 
	\sa_count[1].r.part0[5] , \sa_count[1].r.part0[4] , 
	\sa_count[1].r.part0[3] , \sa_count[1].r.part0[2] , 
	\sa_count[1].r.part0[1] , \sa_count[1].r.part0[0] , 
	\sa_count[0].r.part1[31] , \sa_count[0].r.part1[30] , 
	\sa_count[0].r.part1[29] , \sa_count[0].r.part1[28] , 
	\sa_count[0].r.part1[27] , \sa_count[0].r.part1[26] , 
	\sa_count[0].r.part1[25] , \sa_count[0].r.part1[24] , 
	\sa_count[0].r.part1[23] , \sa_count[0].r.part1[22] , 
	\sa_count[0].r.part1[21] , \sa_count[0].r.part1[20] , 
	\sa_count[0].r.part1[19] , \sa_count[0].r.part1[18] , 
	\sa_count[0].r.part1[17] , \sa_count[0].r.part1[16] , 
	\sa_count[0].r.part1[15] , \sa_count[0].r.part1[14] , 
	\sa_count[0].r.part1[13] , \sa_count[0].r.part1[12] , 
	\sa_count[0].r.part1[11] , \sa_count[0].r.part1[10] , 
	\sa_count[0].r.part1[9] , \sa_count[0].r.part1[8] , 
	\sa_count[0].r.part1[7] , \sa_count[0].r.part1[6] , 
	\sa_count[0].r.part1[5] , \sa_count[0].r.part1[4] , 
	\sa_count[0].r.part1[3] , \sa_count[0].r.part1[2] , 
	\sa_count[0].r.part1[1] , \sa_count[0].r.part1[0] , 
	\sa_count[0].r.part0[31] , \sa_count[0].r.part0[30] , 
	\sa_count[0].r.part0[29] , \sa_count[0].r.part0[28] , 
	\sa_count[0].r.part0[27] , \sa_count[0].r.part0[26] , 
	\sa_count[0].r.part0[25] , \sa_count[0].r.part0[24] , 
	\sa_count[0].r.part0[23] , \sa_count[0].r.part0[22] , 
	\sa_count[0].r.part0[21] , \sa_count[0].r.part0[20] , 
	\sa_count[0].r.part0[19] , \sa_count[0].r.part0[18] , 
	\sa_count[0].r.part0[17] , \sa_count[0].r.part0[16] , 
	\sa_count[0].r.part0[15] , \sa_count[0].r.part0[14] , 
	\sa_count[0].r.part0[13] , \sa_count[0].r.part0[12] , 
	\sa_count[0].r.part0[11] , \sa_count[0].r.part0[10] , 
	\sa_count[0].r.part0[9] , \sa_count[0].r.part0[8] , 
	\sa_count[0].r.part0[7] , \sa_count[0].r.part0[6] , 
	\sa_count[0].r.part0[5] , \sa_count[0].r.part0[4] , 
	\sa_count[0].r.part0[3] , \sa_count[0].r.part0[2] , 
	\sa_count[0].r.part0[1] , \sa_count[0].r.part0[0] } ), kme_idle, 
	.idle_components( {\idle_components.r.part0 [31], 
	\idle_components.r.part0 [30], \idle_components.r.part0 [29], 
	\idle_components.r.part0 [28], \idle_components.r.part0 [27], 
	\idle_components.r.part0 [26], \idle_components.r.part0 [25], 
	\idle_components.r.part0 [24], \idle_components.r.part0 [23], 
	\idle_components.r.part0 [22], \idle_components.r.part0 [21], 
	\idle_components.r.part0 [20], \idle_components.r.part0 [19], 
	\idle_components.r.part0 [18], \idle_components.r.part0 [17], 
	\idle_components.r.part0 [16], \idle_components.r.part0 [15], 
	\idle_components.r.part0 [14], \idle_components.r.part0 [13], 
	\idle_components.r.part0 [12], \idle_components.r.part0 [11], 
	\idle_components.r.part0 [10], \idle_components.r.part0 [9], 
	\idle_components.r.part0 [8], \idle_components.r.part0 [7], 
	\idle_components.r.part0 [6], \idle_components.r.part0 [5], 
	\idle_components.r.part0 [4], \idle_components.r.part0 [3], 
	\idle_components.r.part0 [2], \idle_components.r.part0 [1], 
	\idle_components.r.part0 [0]} ), clk, rst_n, disable_debug_cmd, 
	cceip_encrypt_gcm_tag_fail_int, cceip_validate_gcm_tag_fail_int, 
	cddip_decrypt_gcm_tag_fail_int, cceip_ob_full, cddip_ob_full, 
	.tready_override( {\tready_override.r.part0 [8], 
	\tready_override.r.part0 [7], \tready_override.r.part0 [6], 
	\tready_override.r.part0 [5], \tready_override.r.part0 [4], 
	\tready_override.r.part0 [3], \tready_override.r.part0 [2], 
	\tready_override.r.part0 [1], \tready_override.r.part0 [0]} ), 
	.core_kme_ib_out( {\core_kme_ib_out.tready } ), .sa_global_ctrl( {
	\sa_global_ctrl.r.part0 [31], \sa_global_ctrl.r.part0 [30], 
	\sa_global_ctrl.r.part0 [29], \sa_global_ctrl.r.part0 [28], 
	\sa_global_ctrl.r.part0 [27], \sa_global_ctrl.r.part0 [26], 
	\sa_global_ctrl.r.part0 [25], \sa_global_ctrl.r.part0 [24], 
	\sa_global_ctrl.r.part0 [23], \sa_global_ctrl.r.part0 [22], 
	\sa_global_ctrl.r.part0 [21], \sa_global_ctrl.r.part0 [20], 
	\sa_global_ctrl.r.part0 [19], \sa_global_ctrl.r.part0 [18], 
	\sa_global_ctrl.r.part0 [17], \sa_global_ctrl.r.part0 [16], 
	\sa_global_ctrl.r.part0 [15], \sa_global_ctrl.r.part0 [14], 
	\sa_global_ctrl.r.part0 [13], \sa_global_ctrl.r.part0 [12], 
	\sa_global_ctrl.r.part0 [11], \sa_global_ctrl.r.part0 [10], 
	\sa_global_ctrl.r.part0 [9], \sa_global_ctrl.r.part0 [8], 
	\sa_global_ctrl.r.part0 [7], \sa_global_ctrl.r.part0 [6], 
	\sa_global_ctrl.r.part0 [5], \sa_global_ctrl.r.part0 [4], 
	\sa_global_ctrl.r.part0 [3], \sa_global_ctrl.r.part0 [2], 
	\sa_global_ctrl.r.part0 [1], \sa_global_ctrl.r.part0 [0]} ), .sa_ctrl( {
	\sa_ctrl[31].r.part0[31] , \sa_ctrl[31].r.part0[30] , 
	\sa_ctrl[31].r.part0[29] , \sa_ctrl[31].r.part0[28] , 
	\sa_ctrl[31].r.part0[27] , \sa_ctrl[31].r.part0[26] , 
	\sa_ctrl[31].r.part0[25] , \sa_ctrl[31].r.part0[24] , 
	\sa_ctrl[31].r.part0[23] , \sa_ctrl[31].r.part0[22] , 
	\sa_ctrl[31].r.part0[21] , \sa_ctrl[31].r.part0[20] , 
	\sa_ctrl[31].r.part0[19] , \sa_ctrl[31].r.part0[18] , 
	\sa_ctrl[31].r.part0[17] , \sa_ctrl[31].r.part0[16] , 
	\sa_ctrl[31].r.part0[15] , \sa_ctrl[31].r.part0[14] , 
	\sa_ctrl[31].r.part0[13] , \sa_ctrl[31].r.part0[12] , 
	\sa_ctrl[31].r.part0[11] , \sa_ctrl[31].r.part0[10] , 
	\sa_ctrl[31].r.part0[9] , \sa_ctrl[31].r.part0[8] , 
	\sa_ctrl[31].r.part0[7] , \sa_ctrl[31].r.part0[6] , 
	\sa_ctrl[31].r.part0[5] , \sa_ctrl[31].r.part0[4] , 
	\sa_ctrl[31].r.part0[3] , \sa_ctrl[31].r.part0[2] , 
	\sa_ctrl[31].r.part0[1] , \sa_ctrl[31].r.part0[0] , 
	\sa_ctrl[30].r.part0[31] , \sa_ctrl[30].r.part0[30] , 
	\sa_ctrl[30].r.part0[29] , \sa_ctrl[30].r.part0[28] , 
	\sa_ctrl[30].r.part0[27] , \sa_ctrl[30].r.part0[26] , 
	\sa_ctrl[30].r.part0[25] , \sa_ctrl[30].r.part0[24] , 
	\sa_ctrl[30].r.part0[23] , \sa_ctrl[30].r.part0[22] , 
	\sa_ctrl[30].r.part0[21] , \sa_ctrl[30].r.part0[20] , 
	\sa_ctrl[30].r.part0[19] , \sa_ctrl[30].r.part0[18] , 
	\sa_ctrl[30].r.part0[17] , \sa_ctrl[30].r.part0[16] , 
	\sa_ctrl[30].r.part0[15] , \sa_ctrl[30].r.part0[14] , 
	\sa_ctrl[30].r.part0[13] , \sa_ctrl[30].r.part0[12] , 
	\sa_ctrl[30].r.part0[11] , \sa_ctrl[30].r.part0[10] , 
	\sa_ctrl[30].r.part0[9] , \sa_ctrl[30].r.part0[8] , 
	\sa_ctrl[30].r.part0[7] , \sa_ctrl[30].r.part0[6] , 
	\sa_ctrl[30].r.part0[5] , \sa_ctrl[30].r.part0[4] , 
	\sa_ctrl[30].r.part0[3] , \sa_ctrl[30].r.part0[2] , 
	\sa_ctrl[30].r.part0[1] , \sa_ctrl[30].r.part0[0] , 
	\sa_ctrl[29].r.part0[31] , \sa_ctrl[29].r.part0[30] , 
	\sa_ctrl[29].r.part0[29] , \sa_ctrl[29].r.part0[28] , 
	\sa_ctrl[29].r.part0[27] , \sa_ctrl[29].r.part0[26] , 
	\sa_ctrl[29].r.part0[25] , \sa_ctrl[29].r.part0[24] , 
	\sa_ctrl[29].r.part0[23] , \sa_ctrl[29].r.part0[22] , 
	\sa_ctrl[29].r.part0[21] , \sa_ctrl[29].r.part0[20] , 
	\sa_ctrl[29].r.part0[19] , \sa_ctrl[29].r.part0[18] , 
	\sa_ctrl[29].r.part0[17] , \sa_ctrl[29].r.part0[16] , 
	\sa_ctrl[29].r.part0[15] , \sa_ctrl[29].r.part0[14] , 
	\sa_ctrl[29].r.part0[13] , \sa_ctrl[29].r.part0[12] , 
	\sa_ctrl[29].r.part0[11] , \sa_ctrl[29].r.part0[10] , 
	\sa_ctrl[29].r.part0[9] , \sa_ctrl[29].r.part0[8] , 
	\sa_ctrl[29].r.part0[7] , \sa_ctrl[29].r.part0[6] , 
	\sa_ctrl[29].r.part0[5] , \sa_ctrl[29].r.part0[4] , 
	\sa_ctrl[29].r.part0[3] , \sa_ctrl[29].r.part0[2] , 
	\sa_ctrl[29].r.part0[1] , \sa_ctrl[29].r.part0[0] , 
	\sa_ctrl[28].r.part0[31] , \sa_ctrl[28].r.part0[30] , 
	\sa_ctrl[28].r.part0[29] , \sa_ctrl[28].r.part0[28] , 
	\sa_ctrl[28].r.part0[27] , \sa_ctrl[28].r.part0[26] , 
	\sa_ctrl[28].r.part0[25] , \sa_ctrl[28].r.part0[24] , 
	\sa_ctrl[28].r.part0[23] , \sa_ctrl[28].r.part0[22] , 
	\sa_ctrl[28].r.part0[21] , \sa_ctrl[28].r.part0[20] , 
	\sa_ctrl[28].r.part0[19] , \sa_ctrl[28].r.part0[18] , 
	\sa_ctrl[28].r.part0[17] , \sa_ctrl[28].r.part0[16] , 
	\sa_ctrl[28].r.part0[15] , \sa_ctrl[28].r.part0[14] , 
	\sa_ctrl[28].r.part0[13] , \sa_ctrl[28].r.part0[12] , 
	\sa_ctrl[28].r.part0[11] , \sa_ctrl[28].r.part0[10] , 
	\sa_ctrl[28].r.part0[9] , \sa_ctrl[28].r.part0[8] , 
	\sa_ctrl[28].r.part0[7] , \sa_ctrl[28].r.part0[6] , 
	\sa_ctrl[28].r.part0[5] , \sa_ctrl[28].r.part0[4] , 
	\sa_ctrl[28].r.part0[3] , \sa_ctrl[28].r.part0[2] , 
	\sa_ctrl[28].r.part0[1] , \sa_ctrl[28].r.part0[0] , 
	\sa_ctrl[27].r.part0[31] , \sa_ctrl[27].r.part0[30] , 
	\sa_ctrl[27].r.part0[29] , \sa_ctrl[27].r.part0[28] , 
	\sa_ctrl[27].r.part0[27] , \sa_ctrl[27].r.part0[26] , 
	\sa_ctrl[27].r.part0[25] , \sa_ctrl[27].r.part0[24] , 
	\sa_ctrl[27].r.part0[23] , \sa_ctrl[27].r.part0[22] , 
	\sa_ctrl[27].r.part0[21] , \sa_ctrl[27].r.part0[20] , 
	\sa_ctrl[27].r.part0[19] , \sa_ctrl[27].r.part0[18] , 
	\sa_ctrl[27].r.part0[17] , \sa_ctrl[27].r.part0[16] , 
	\sa_ctrl[27].r.part0[15] , \sa_ctrl[27].r.part0[14] , 
	\sa_ctrl[27].r.part0[13] , \sa_ctrl[27].r.part0[12] , 
	\sa_ctrl[27].r.part0[11] , \sa_ctrl[27].r.part0[10] , 
	\sa_ctrl[27].r.part0[9] , \sa_ctrl[27].r.part0[8] , 
	\sa_ctrl[27].r.part0[7] , \sa_ctrl[27].r.part0[6] , 
	\sa_ctrl[27].r.part0[5] , \sa_ctrl[27].r.part0[4] , 
	\sa_ctrl[27].r.part0[3] , \sa_ctrl[27].r.part0[2] , 
	\sa_ctrl[27].r.part0[1] , \sa_ctrl[27].r.part0[0] , 
	\sa_ctrl[26].r.part0[31] , \sa_ctrl[26].r.part0[30] , 
	\sa_ctrl[26].r.part0[29] , \sa_ctrl[26].r.part0[28] , 
	\sa_ctrl[26].r.part0[27] , \sa_ctrl[26].r.part0[26] , 
	\sa_ctrl[26].r.part0[25] , \sa_ctrl[26].r.part0[24] , 
	\sa_ctrl[26].r.part0[23] , \sa_ctrl[26].r.part0[22] , 
	\sa_ctrl[26].r.part0[21] , \sa_ctrl[26].r.part0[20] , 
	\sa_ctrl[26].r.part0[19] , \sa_ctrl[26].r.part0[18] , 
	\sa_ctrl[26].r.part0[17] , \sa_ctrl[26].r.part0[16] , 
	\sa_ctrl[26].r.part0[15] , \sa_ctrl[26].r.part0[14] , 
	\sa_ctrl[26].r.part0[13] , \sa_ctrl[26].r.part0[12] , 
	\sa_ctrl[26].r.part0[11] , \sa_ctrl[26].r.part0[10] , 
	\sa_ctrl[26].r.part0[9] , \sa_ctrl[26].r.part0[8] , 
	\sa_ctrl[26].r.part0[7] , \sa_ctrl[26].r.part0[6] , 
	\sa_ctrl[26].r.part0[5] , \sa_ctrl[26].r.part0[4] , 
	\sa_ctrl[26].r.part0[3] , \sa_ctrl[26].r.part0[2] , 
	\sa_ctrl[26].r.part0[1] , \sa_ctrl[26].r.part0[0] , 
	\sa_ctrl[25].r.part0[31] , \sa_ctrl[25].r.part0[30] , 
	\sa_ctrl[25].r.part0[29] , \sa_ctrl[25].r.part0[28] , 
	\sa_ctrl[25].r.part0[27] , \sa_ctrl[25].r.part0[26] , 
	\sa_ctrl[25].r.part0[25] , \sa_ctrl[25].r.part0[24] , 
	\sa_ctrl[25].r.part0[23] , \sa_ctrl[25].r.part0[22] , 
	\sa_ctrl[25].r.part0[21] , \sa_ctrl[25].r.part0[20] , 
	\sa_ctrl[25].r.part0[19] , \sa_ctrl[25].r.part0[18] , 
	\sa_ctrl[25].r.part0[17] , \sa_ctrl[25].r.part0[16] , 
	\sa_ctrl[25].r.part0[15] , \sa_ctrl[25].r.part0[14] , 
	\sa_ctrl[25].r.part0[13] , \sa_ctrl[25].r.part0[12] , 
	\sa_ctrl[25].r.part0[11] , \sa_ctrl[25].r.part0[10] , 
	\sa_ctrl[25].r.part0[9] , \sa_ctrl[25].r.part0[8] , 
	\sa_ctrl[25].r.part0[7] , \sa_ctrl[25].r.part0[6] , 
	\sa_ctrl[25].r.part0[5] , \sa_ctrl[25].r.part0[4] , 
	\sa_ctrl[25].r.part0[3] , \sa_ctrl[25].r.part0[2] , 
	\sa_ctrl[25].r.part0[1] , \sa_ctrl[25].r.part0[0] , 
	\sa_ctrl[24].r.part0[31] , \sa_ctrl[24].r.part0[30] , 
	\sa_ctrl[24].r.part0[29] , \sa_ctrl[24].r.part0[28] , 
	\sa_ctrl[24].r.part0[27] , \sa_ctrl[24].r.part0[26] , 
	\sa_ctrl[24].r.part0[25] , \sa_ctrl[24].r.part0[24] , 
	\sa_ctrl[24].r.part0[23] , \sa_ctrl[24].r.part0[22] , 
	\sa_ctrl[24].r.part0[21] , \sa_ctrl[24].r.part0[20] , 
	\sa_ctrl[24].r.part0[19] , \sa_ctrl[24].r.part0[18] , 
	\sa_ctrl[24].r.part0[17] , \sa_ctrl[24].r.part0[16] , 
	\sa_ctrl[24].r.part0[15] , \sa_ctrl[24].r.part0[14] , 
	\sa_ctrl[24].r.part0[13] , \sa_ctrl[24].r.part0[12] , 
	\sa_ctrl[24].r.part0[11] , \sa_ctrl[24].r.part0[10] , 
	\sa_ctrl[24].r.part0[9] , \sa_ctrl[24].r.part0[8] , 
	\sa_ctrl[24].r.part0[7] , \sa_ctrl[24].r.part0[6] , 
	\sa_ctrl[24].r.part0[5] , \sa_ctrl[24].r.part0[4] , 
	\sa_ctrl[24].r.part0[3] , \sa_ctrl[24].r.part0[2] , 
	\sa_ctrl[24].r.part0[1] , \sa_ctrl[24].r.part0[0] , 
	\sa_ctrl[23].r.part0[31] , \sa_ctrl[23].r.part0[30] , 
	\sa_ctrl[23].r.part0[29] , \sa_ctrl[23].r.part0[28] , 
	\sa_ctrl[23].r.part0[27] , \sa_ctrl[23].r.part0[26] , 
	\sa_ctrl[23].r.part0[25] , \sa_ctrl[23].r.part0[24] , 
	\sa_ctrl[23].r.part0[23] , \sa_ctrl[23].r.part0[22] , 
	\sa_ctrl[23].r.part0[21] , \sa_ctrl[23].r.part0[20] , 
	\sa_ctrl[23].r.part0[19] , \sa_ctrl[23].r.part0[18] , 
	\sa_ctrl[23].r.part0[17] , \sa_ctrl[23].r.part0[16] , 
	\sa_ctrl[23].r.part0[15] , \sa_ctrl[23].r.part0[14] , 
	\sa_ctrl[23].r.part0[13] , \sa_ctrl[23].r.part0[12] , 
	\sa_ctrl[23].r.part0[11] , \sa_ctrl[23].r.part0[10] , 
	\sa_ctrl[23].r.part0[9] , \sa_ctrl[23].r.part0[8] , 
	\sa_ctrl[23].r.part0[7] , \sa_ctrl[23].r.part0[6] , 
	\sa_ctrl[23].r.part0[5] , \sa_ctrl[23].r.part0[4] , 
	\sa_ctrl[23].r.part0[3] , \sa_ctrl[23].r.part0[2] , 
	\sa_ctrl[23].r.part0[1] , \sa_ctrl[23].r.part0[0] , 
	\sa_ctrl[22].r.part0[31] , \sa_ctrl[22].r.part0[30] , 
	\sa_ctrl[22].r.part0[29] , \sa_ctrl[22].r.part0[28] , 
	\sa_ctrl[22].r.part0[27] , \sa_ctrl[22].r.part0[26] , 
	\sa_ctrl[22].r.part0[25] , \sa_ctrl[22].r.part0[24] , 
	\sa_ctrl[22].r.part0[23] , \sa_ctrl[22].r.part0[22] , 
	\sa_ctrl[22].r.part0[21] , \sa_ctrl[22].r.part0[20] , 
	\sa_ctrl[22].r.part0[19] , \sa_ctrl[22].r.part0[18] , 
	\sa_ctrl[22].r.part0[17] , \sa_ctrl[22].r.part0[16] , 
	\sa_ctrl[22].r.part0[15] , \sa_ctrl[22].r.part0[14] , 
	\sa_ctrl[22].r.part0[13] , \sa_ctrl[22].r.part0[12] , 
	\sa_ctrl[22].r.part0[11] , \sa_ctrl[22].r.part0[10] , 
	\sa_ctrl[22].r.part0[9] , \sa_ctrl[22].r.part0[8] , 
	\sa_ctrl[22].r.part0[7] , \sa_ctrl[22].r.part0[6] , 
	\sa_ctrl[22].r.part0[5] , \sa_ctrl[22].r.part0[4] , 
	\sa_ctrl[22].r.part0[3] , \sa_ctrl[22].r.part0[2] , 
	\sa_ctrl[22].r.part0[1] , \sa_ctrl[22].r.part0[0] , 
	\sa_ctrl[21].r.part0[31] , \sa_ctrl[21].r.part0[30] , 
	\sa_ctrl[21].r.part0[29] , \sa_ctrl[21].r.part0[28] , 
	\sa_ctrl[21].r.part0[27] , \sa_ctrl[21].r.part0[26] , 
	\sa_ctrl[21].r.part0[25] , \sa_ctrl[21].r.part0[24] , 
	\sa_ctrl[21].r.part0[23] , \sa_ctrl[21].r.part0[22] , 
	\sa_ctrl[21].r.part0[21] , \sa_ctrl[21].r.part0[20] , 
	\sa_ctrl[21].r.part0[19] , \sa_ctrl[21].r.part0[18] , 
	\sa_ctrl[21].r.part0[17] , \sa_ctrl[21].r.part0[16] , 
	\sa_ctrl[21].r.part0[15] , \sa_ctrl[21].r.part0[14] , 
	\sa_ctrl[21].r.part0[13] , \sa_ctrl[21].r.part0[12] , 
	\sa_ctrl[21].r.part0[11] , \sa_ctrl[21].r.part0[10] , 
	\sa_ctrl[21].r.part0[9] , \sa_ctrl[21].r.part0[8] , 
	\sa_ctrl[21].r.part0[7] , \sa_ctrl[21].r.part0[6] , 
	\sa_ctrl[21].r.part0[5] , \sa_ctrl[21].r.part0[4] , 
	\sa_ctrl[21].r.part0[3] , \sa_ctrl[21].r.part0[2] , 
	\sa_ctrl[21].r.part0[1] , \sa_ctrl[21].r.part0[0] , 
	\sa_ctrl[20].r.part0[31] , \sa_ctrl[20].r.part0[30] , 
	\sa_ctrl[20].r.part0[29] , \sa_ctrl[20].r.part0[28] , 
	\sa_ctrl[20].r.part0[27] , \sa_ctrl[20].r.part0[26] , 
	\sa_ctrl[20].r.part0[25] , \sa_ctrl[20].r.part0[24] , 
	\sa_ctrl[20].r.part0[23] , \sa_ctrl[20].r.part0[22] , 
	\sa_ctrl[20].r.part0[21] , \sa_ctrl[20].r.part0[20] , 
	\sa_ctrl[20].r.part0[19] , \sa_ctrl[20].r.part0[18] , 
	\sa_ctrl[20].r.part0[17] , \sa_ctrl[20].r.part0[16] , 
	\sa_ctrl[20].r.part0[15] , \sa_ctrl[20].r.part0[14] , 
	\sa_ctrl[20].r.part0[13] , \sa_ctrl[20].r.part0[12] , 
	\sa_ctrl[20].r.part0[11] , \sa_ctrl[20].r.part0[10] , 
	\sa_ctrl[20].r.part0[9] , \sa_ctrl[20].r.part0[8] , 
	\sa_ctrl[20].r.part0[7] , \sa_ctrl[20].r.part0[6] , 
	\sa_ctrl[20].r.part0[5] , \sa_ctrl[20].r.part0[4] , 
	\sa_ctrl[20].r.part0[3] , \sa_ctrl[20].r.part0[2] , 
	\sa_ctrl[20].r.part0[1] , \sa_ctrl[20].r.part0[0] , 
	\sa_ctrl[19].r.part0[31] , \sa_ctrl[19].r.part0[30] , 
	\sa_ctrl[19].r.part0[29] , \sa_ctrl[19].r.part0[28] , 
	\sa_ctrl[19].r.part0[27] , \sa_ctrl[19].r.part0[26] , 
	\sa_ctrl[19].r.part0[25] , \sa_ctrl[19].r.part0[24] , 
	\sa_ctrl[19].r.part0[23] , \sa_ctrl[19].r.part0[22] , 
	\sa_ctrl[19].r.part0[21] , \sa_ctrl[19].r.part0[20] , 
	\sa_ctrl[19].r.part0[19] , \sa_ctrl[19].r.part0[18] , 
	\sa_ctrl[19].r.part0[17] , \sa_ctrl[19].r.part0[16] , 
	\sa_ctrl[19].r.part0[15] , \sa_ctrl[19].r.part0[14] , 
	\sa_ctrl[19].r.part0[13] , \sa_ctrl[19].r.part0[12] , 
	\sa_ctrl[19].r.part0[11] , \sa_ctrl[19].r.part0[10] , 
	\sa_ctrl[19].r.part0[9] , \sa_ctrl[19].r.part0[8] , 
	\sa_ctrl[19].r.part0[7] , \sa_ctrl[19].r.part0[6] , 
	\sa_ctrl[19].r.part0[5] , \sa_ctrl[19].r.part0[4] , 
	\sa_ctrl[19].r.part0[3] , \sa_ctrl[19].r.part0[2] , 
	\sa_ctrl[19].r.part0[1] , \sa_ctrl[19].r.part0[0] , 
	\sa_ctrl[18].r.part0[31] , \sa_ctrl[18].r.part0[30] , 
	\sa_ctrl[18].r.part0[29] , \sa_ctrl[18].r.part0[28] , 
	\sa_ctrl[18].r.part0[27] , \sa_ctrl[18].r.part0[26] , 
	\sa_ctrl[18].r.part0[25] , \sa_ctrl[18].r.part0[24] , 
	\sa_ctrl[18].r.part0[23] , \sa_ctrl[18].r.part0[22] , 
	\sa_ctrl[18].r.part0[21] , \sa_ctrl[18].r.part0[20] , 
	\sa_ctrl[18].r.part0[19] , \sa_ctrl[18].r.part0[18] , 
	\sa_ctrl[18].r.part0[17] , \sa_ctrl[18].r.part0[16] , 
	\sa_ctrl[18].r.part0[15] , \sa_ctrl[18].r.part0[14] , 
	\sa_ctrl[18].r.part0[13] , \sa_ctrl[18].r.part0[12] , 
	\sa_ctrl[18].r.part0[11] , \sa_ctrl[18].r.part0[10] , 
	\sa_ctrl[18].r.part0[9] , \sa_ctrl[18].r.part0[8] , 
	\sa_ctrl[18].r.part0[7] , \sa_ctrl[18].r.part0[6] , 
	\sa_ctrl[18].r.part0[5] , \sa_ctrl[18].r.part0[4] , 
	\sa_ctrl[18].r.part0[3] , \sa_ctrl[18].r.part0[2] , 
	\sa_ctrl[18].r.part0[1] , \sa_ctrl[18].r.part0[0] , 
	\sa_ctrl[17].r.part0[31] , \sa_ctrl[17].r.part0[30] , 
	\sa_ctrl[17].r.part0[29] , \sa_ctrl[17].r.part0[28] , 
	\sa_ctrl[17].r.part0[27] , \sa_ctrl[17].r.part0[26] , 
	\sa_ctrl[17].r.part0[25] , \sa_ctrl[17].r.part0[24] , 
	\sa_ctrl[17].r.part0[23] , \sa_ctrl[17].r.part0[22] , 
	\sa_ctrl[17].r.part0[21] , \sa_ctrl[17].r.part0[20] , 
	\sa_ctrl[17].r.part0[19] , \sa_ctrl[17].r.part0[18] , 
	\sa_ctrl[17].r.part0[17] , \sa_ctrl[17].r.part0[16] , 
	\sa_ctrl[17].r.part0[15] , \sa_ctrl[17].r.part0[14] , 
	\sa_ctrl[17].r.part0[13] , \sa_ctrl[17].r.part0[12] , 
	\sa_ctrl[17].r.part0[11] , \sa_ctrl[17].r.part0[10] , 
	\sa_ctrl[17].r.part0[9] , \sa_ctrl[17].r.part0[8] , 
	\sa_ctrl[17].r.part0[7] , \sa_ctrl[17].r.part0[6] , 
	\sa_ctrl[17].r.part0[5] , \sa_ctrl[17].r.part0[4] , 
	\sa_ctrl[17].r.part0[3] , \sa_ctrl[17].r.part0[2] , 
	\sa_ctrl[17].r.part0[1] , \sa_ctrl[17].r.part0[0] , 
	\sa_ctrl[16].r.part0[31] , \sa_ctrl[16].r.part0[30] , 
	\sa_ctrl[16].r.part0[29] , \sa_ctrl[16].r.part0[28] , 
	\sa_ctrl[16].r.part0[27] , \sa_ctrl[16].r.part0[26] , 
	\sa_ctrl[16].r.part0[25] , \sa_ctrl[16].r.part0[24] , 
	\sa_ctrl[16].r.part0[23] , \sa_ctrl[16].r.part0[22] , 
	\sa_ctrl[16].r.part0[21] , \sa_ctrl[16].r.part0[20] , 
	\sa_ctrl[16].r.part0[19] , \sa_ctrl[16].r.part0[18] , 
	\sa_ctrl[16].r.part0[17] , \sa_ctrl[16].r.part0[16] , 
	\sa_ctrl[16].r.part0[15] , \sa_ctrl[16].r.part0[14] , 
	\sa_ctrl[16].r.part0[13] , \sa_ctrl[16].r.part0[12] , 
	\sa_ctrl[16].r.part0[11] , \sa_ctrl[16].r.part0[10] , 
	\sa_ctrl[16].r.part0[9] , \sa_ctrl[16].r.part0[8] , 
	\sa_ctrl[16].r.part0[7] , \sa_ctrl[16].r.part0[6] , 
	\sa_ctrl[16].r.part0[5] , \sa_ctrl[16].r.part0[4] , 
	\sa_ctrl[16].r.part0[3] , \sa_ctrl[16].r.part0[2] , 
	\sa_ctrl[16].r.part0[1] , \sa_ctrl[16].r.part0[0] , 
	\sa_ctrl[15].r.part0[31] , \sa_ctrl[15].r.part0[30] , 
	\sa_ctrl[15].r.part0[29] , \sa_ctrl[15].r.part0[28] , 
	\sa_ctrl[15].r.part0[27] , \sa_ctrl[15].r.part0[26] , 
	\sa_ctrl[15].r.part0[25] , \sa_ctrl[15].r.part0[24] , 
	\sa_ctrl[15].r.part0[23] , \sa_ctrl[15].r.part0[22] , 
	\sa_ctrl[15].r.part0[21] , \sa_ctrl[15].r.part0[20] , 
	\sa_ctrl[15].r.part0[19] , \sa_ctrl[15].r.part0[18] , 
	\sa_ctrl[15].r.part0[17] , \sa_ctrl[15].r.part0[16] , 
	\sa_ctrl[15].r.part0[15] , \sa_ctrl[15].r.part0[14] , 
	\sa_ctrl[15].r.part0[13] , \sa_ctrl[15].r.part0[12] , 
	\sa_ctrl[15].r.part0[11] , \sa_ctrl[15].r.part0[10] , 
	\sa_ctrl[15].r.part0[9] , \sa_ctrl[15].r.part0[8] , 
	\sa_ctrl[15].r.part0[7] , \sa_ctrl[15].r.part0[6] , 
	\sa_ctrl[15].r.part0[5] , \sa_ctrl[15].r.part0[4] , 
	\sa_ctrl[15].r.part0[3] , \sa_ctrl[15].r.part0[2] , 
	\sa_ctrl[15].r.part0[1] , \sa_ctrl[15].r.part0[0] , 
	\sa_ctrl[14].r.part0[31] , \sa_ctrl[14].r.part0[30] , 
	\sa_ctrl[14].r.part0[29] , \sa_ctrl[14].r.part0[28] , 
	\sa_ctrl[14].r.part0[27] , \sa_ctrl[14].r.part0[26] , 
	\sa_ctrl[14].r.part0[25] , \sa_ctrl[14].r.part0[24] , 
	\sa_ctrl[14].r.part0[23] , \sa_ctrl[14].r.part0[22] , 
	\sa_ctrl[14].r.part0[21] , \sa_ctrl[14].r.part0[20] , 
	\sa_ctrl[14].r.part0[19] , \sa_ctrl[14].r.part0[18] , 
	\sa_ctrl[14].r.part0[17] , \sa_ctrl[14].r.part0[16] , 
	\sa_ctrl[14].r.part0[15] , \sa_ctrl[14].r.part0[14] , 
	\sa_ctrl[14].r.part0[13] , \sa_ctrl[14].r.part0[12] , 
	\sa_ctrl[14].r.part0[11] , \sa_ctrl[14].r.part0[10] , 
	\sa_ctrl[14].r.part0[9] , \sa_ctrl[14].r.part0[8] , 
	\sa_ctrl[14].r.part0[7] , \sa_ctrl[14].r.part0[6] , 
	\sa_ctrl[14].r.part0[5] , \sa_ctrl[14].r.part0[4] , 
	\sa_ctrl[14].r.part0[3] , \sa_ctrl[14].r.part0[2] , 
	\sa_ctrl[14].r.part0[1] , \sa_ctrl[14].r.part0[0] , 
	\sa_ctrl[13].r.part0[31] , \sa_ctrl[13].r.part0[30] , 
	\sa_ctrl[13].r.part0[29] , \sa_ctrl[13].r.part0[28] , 
	\sa_ctrl[13].r.part0[27] , \sa_ctrl[13].r.part0[26] , 
	\sa_ctrl[13].r.part0[25] , \sa_ctrl[13].r.part0[24] , 
	\sa_ctrl[13].r.part0[23] , \sa_ctrl[13].r.part0[22] , 
	\sa_ctrl[13].r.part0[21] , \sa_ctrl[13].r.part0[20] , 
	\sa_ctrl[13].r.part0[19] , \sa_ctrl[13].r.part0[18] , 
	\sa_ctrl[13].r.part0[17] , \sa_ctrl[13].r.part0[16] , 
	\sa_ctrl[13].r.part0[15] , \sa_ctrl[13].r.part0[14] , 
	\sa_ctrl[13].r.part0[13] , \sa_ctrl[13].r.part0[12] , 
	\sa_ctrl[13].r.part0[11] , \sa_ctrl[13].r.part0[10] , 
	\sa_ctrl[13].r.part0[9] , \sa_ctrl[13].r.part0[8] , 
	\sa_ctrl[13].r.part0[7] , \sa_ctrl[13].r.part0[6] , 
	\sa_ctrl[13].r.part0[5] , \sa_ctrl[13].r.part0[4] , 
	\sa_ctrl[13].r.part0[3] , \sa_ctrl[13].r.part0[2] , 
	\sa_ctrl[13].r.part0[1] , \sa_ctrl[13].r.part0[0] , 
	\sa_ctrl[12].r.part0[31] , \sa_ctrl[12].r.part0[30] , 
	\sa_ctrl[12].r.part0[29] , \sa_ctrl[12].r.part0[28] , 
	\sa_ctrl[12].r.part0[27] , \sa_ctrl[12].r.part0[26] , 
	\sa_ctrl[12].r.part0[25] , \sa_ctrl[12].r.part0[24] , 
	\sa_ctrl[12].r.part0[23] , \sa_ctrl[12].r.part0[22] , 
	\sa_ctrl[12].r.part0[21] , \sa_ctrl[12].r.part0[20] , 
	\sa_ctrl[12].r.part0[19] , \sa_ctrl[12].r.part0[18] , 
	\sa_ctrl[12].r.part0[17] , \sa_ctrl[12].r.part0[16] , 
	\sa_ctrl[12].r.part0[15] , \sa_ctrl[12].r.part0[14] , 
	\sa_ctrl[12].r.part0[13] , \sa_ctrl[12].r.part0[12] , 
	\sa_ctrl[12].r.part0[11] , \sa_ctrl[12].r.part0[10] , 
	\sa_ctrl[12].r.part0[9] , \sa_ctrl[12].r.part0[8] , 
	\sa_ctrl[12].r.part0[7] , \sa_ctrl[12].r.part0[6] , 
	\sa_ctrl[12].r.part0[5] , \sa_ctrl[12].r.part0[4] , 
	\sa_ctrl[12].r.part0[3] , \sa_ctrl[12].r.part0[2] , 
	\sa_ctrl[12].r.part0[1] , \sa_ctrl[12].r.part0[0] , 
	\sa_ctrl[11].r.part0[31] , \sa_ctrl[11].r.part0[30] , 
	\sa_ctrl[11].r.part0[29] , \sa_ctrl[11].r.part0[28] , 
	\sa_ctrl[11].r.part0[27] , \sa_ctrl[11].r.part0[26] , 
	\sa_ctrl[11].r.part0[25] , \sa_ctrl[11].r.part0[24] , 
	\sa_ctrl[11].r.part0[23] , \sa_ctrl[11].r.part0[22] , 
	\sa_ctrl[11].r.part0[21] , \sa_ctrl[11].r.part0[20] , 
	\sa_ctrl[11].r.part0[19] , \sa_ctrl[11].r.part0[18] , 
	\sa_ctrl[11].r.part0[17] , \sa_ctrl[11].r.part0[16] , 
	\sa_ctrl[11].r.part0[15] , \sa_ctrl[11].r.part0[14] , 
	\sa_ctrl[11].r.part0[13] , \sa_ctrl[11].r.part0[12] , 
	\sa_ctrl[11].r.part0[11] , \sa_ctrl[11].r.part0[10] , 
	\sa_ctrl[11].r.part0[9] , \sa_ctrl[11].r.part0[8] , 
	\sa_ctrl[11].r.part0[7] , \sa_ctrl[11].r.part0[6] , 
	\sa_ctrl[11].r.part0[5] , \sa_ctrl[11].r.part0[4] , 
	\sa_ctrl[11].r.part0[3] , \sa_ctrl[11].r.part0[2] , 
	\sa_ctrl[11].r.part0[1] , \sa_ctrl[11].r.part0[0] , 
	\sa_ctrl[10].r.part0[31] , \sa_ctrl[10].r.part0[30] , 
	\sa_ctrl[10].r.part0[29] , \sa_ctrl[10].r.part0[28] , 
	\sa_ctrl[10].r.part0[27] , \sa_ctrl[10].r.part0[26] , 
	\sa_ctrl[10].r.part0[25] , \sa_ctrl[10].r.part0[24] , 
	\sa_ctrl[10].r.part0[23] , \sa_ctrl[10].r.part0[22] , 
	\sa_ctrl[10].r.part0[21] , \sa_ctrl[10].r.part0[20] , 
	\sa_ctrl[10].r.part0[19] , \sa_ctrl[10].r.part0[18] , 
	\sa_ctrl[10].r.part0[17] , \sa_ctrl[10].r.part0[16] , 
	\sa_ctrl[10].r.part0[15] , \sa_ctrl[10].r.part0[14] , 
	\sa_ctrl[10].r.part0[13] , \sa_ctrl[10].r.part0[12] , 
	\sa_ctrl[10].r.part0[11] , \sa_ctrl[10].r.part0[10] , 
	\sa_ctrl[10].r.part0[9] , \sa_ctrl[10].r.part0[8] , 
	\sa_ctrl[10].r.part0[7] , \sa_ctrl[10].r.part0[6] , 
	\sa_ctrl[10].r.part0[5] , \sa_ctrl[10].r.part0[4] , 
	\sa_ctrl[10].r.part0[3] , \sa_ctrl[10].r.part0[2] , 
	\sa_ctrl[10].r.part0[1] , \sa_ctrl[10].r.part0[0] , 
	\sa_ctrl[9].r.part0[31] , \sa_ctrl[9].r.part0[30] , 
	\sa_ctrl[9].r.part0[29] , \sa_ctrl[9].r.part0[28] , 
	\sa_ctrl[9].r.part0[27] , \sa_ctrl[9].r.part0[26] , 
	\sa_ctrl[9].r.part0[25] , \sa_ctrl[9].r.part0[24] , 
	\sa_ctrl[9].r.part0[23] , \sa_ctrl[9].r.part0[22] , 
	\sa_ctrl[9].r.part0[21] , \sa_ctrl[9].r.part0[20] , 
	\sa_ctrl[9].r.part0[19] , \sa_ctrl[9].r.part0[18] , 
	\sa_ctrl[9].r.part0[17] , \sa_ctrl[9].r.part0[16] , 
	\sa_ctrl[9].r.part0[15] , \sa_ctrl[9].r.part0[14] , 
	\sa_ctrl[9].r.part0[13] , \sa_ctrl[9].r.part0[12] , 
	\sa_ctrl[9].r.part0[11] , \sa_ctrl[9].r.part0[10] , 
	\sa_ctrl[9].r.part0[9] , \sa_ctrl[9].r.part0[8] , 
	\sa_ctrl[9].r.part0[7] , \sa_ctrl[9].r.part0[6] , 
	\sa_ctrl[9].r.part0[5] , \sa_ctrl[9].r.part0[4] , 
	\sa_ctrl[9].r.part0[3] , \sa_ctrl[9].r.part0[2] , 
	\sa_ctrl[9].r.part0[1] , \sa_ctrl[9].r.part0[0] , 
	\sa_ctrl[8].r.part0[31] , \sa_ctrl[8].r.part0[30] , 
	\sa_ctrl[8].r.part0[29] , \sa_ctrl[8].r.part0[28] , 
	\sa_ctrl[8].r.part0[27] , \sa_ctrl[8].r.part0[26] , 
	\sa_ctrl[8].r.part0[25] , \sa_ctrl[8].r.part0[24] , 
	\sa_ctrl[8].r.part0[23] , \sa_ctrl[8].r.part0[22] , 
	\sa_ctrl[8].r.part0[21] , \sa_ctrl[8].r.part0[20] , 
	\sa_ctrl[8].r.part0[19] , \sa_ctrl[8].r.part0[18] , 
	\sa_ctrl[8].r.part0[17] , \sa_ctrl[8].r.part0[16] , 
	\sa_ctrl[8].r.part0[15] , \sa_ctrl[8].r.part0[14] , 
	\sa_ctrl[8].r.part0[13] , \sa_ctrl[8].r.part0[12] , 
	\sa_ctrl[8].r.part0[11] , \sa_ctrl[8].r.part0[10] , 
	\sa_ctrl[8].r.part0[9] , \sa_ctrl[8].r.part0[8] , 
	\sa_ctrl[8].r.part0[7] , \sa_ctrl[8].r.part0[6] , 
	\sa_ctrl[8].r.part0[5] , \sa_ctrl[8].r.part0[4] , 
	\sa_ctrl[8].r.part0[3] , \sa_ctrl[8].r.part0[2] , 
	\sa_ctrl[8].r.part0[1] , \sa_ctrl[8].r.part0[0] , 
	\sa_ctrl[7].r.part0[31] , \sa_ctrl[7].r.part0[30] , 
	\sa_ctrl[7].r.part0[29] , \sa_ctrl[7].r.part0[28] , 
	\sa_ctrl[7].r.part0[27] , \sa_ctrl[7].r.part0[26] , 
	\sa_ctrl[7].r.part0[25] , \sa_ctrl[7].r.part0[24] , 
	\sa_ctrl[7].r.part0[23] , \sa_ctrl[7].r.part0[22] , 
	\sa_ctrl[7].r.part0[21] , \sa_ctrl[7].r.part0[20] , 
	\sa_ctrl[7].r.part0[19] , \sa_ctrl[7].r.part0[18] , 
	\sa_ctrl[7].r.part0[17] , \sa_ctrl[7].r.part0[16] , 
	\sa_ctrl[7].r.part0[15] , \sa_ctrl[7].r.part0[14] , 
	\sa_ctrl[7].r.part0[13] , \sa_ctrl[7].r.part0[12] , 
	\sa_ctrl[7].r.part0[11] , \sa_ctrl[7].r.part0[10] , 
	\sa_ctrl[7].r.part0[9] , \sa_ctrl[7].r.part0[8] , 
	\sa_ctrl[7].r.part0[7] , \sa_ctrl[7].r.part0[6] , 
	\sa_ctrl[7].r.part0[5] , \sa_ctrl[7].r.part0[4] , 
	\sa_ctrl[7].r.part0[3] , \sa_ctrl[7].r.part0[2] , 
	\sa_ctrl[7].r.part0[1] , \sa_ctrl[7].r.part0[0] , 
	\sa_ctrl[6].r.part0[31] , \sa_ctrl[6].r.part0[30] , 
	\sa_ctrl[6].r.part0[29] , \sa_ctrl[6].r.part0[28] , 
	\sa_ctrl[6].r.part0[27] , \sa_ctrl[6].r.part0[26] , 
	\sa_ctrl[6].r.part0[25] , \sa_ctrl[6].r.part0[24] , 
	\sa_ctrl[6].r.part0[23] , \sa_ctrl[6].r.part0[22] , 
	\sa_ctrl[6].r.part0[21] , \sa_ctrl[6].r.part0[20] , 
	\sa_ctrl[6].r.part0[19] , \sa_ctrl[6].r.part0[18] , 
	\sa_ctrl[6].r.part0[17] , \sa_ctrl[6].r.part0[16] , 
	\sa_ctrl[6].r.part0[15] , \sa_ctrl[6].r.part0[14] , 
	\sa_ctrl[6].r.part0[13] , \sa_ctrl[6].r.part0[12] , 
	\sa_ctrl[6].r.part0[11] , \sa_ctrl[6].r.part0[10] , 
	\sa_ctrl[6].r.part0[9] , \sa_ctrl[6].r.part0[8] , 
	\sa_ctrl[6].r.part0[7] , \sa_ctrl[6].r.part0[6] , 
	\sa_ctrl[6].r.part0[5] , \sa_ctrl[6].r.part0[4] , 
	\sa_ctrl[6].r.part0[3] , \sa_ctrl[6].r.part0[2] , 
	\sa_ctrl[6].r.part0[1] , \sa_ctrl[6].r.part0[0] , 
	\sa_ctrl[5].r.part0[31] , \sa_ctrl[5].r.part0[30] , 
	\sa_ctrl[5].r.part0[29] , \sa_ctrl[5].r.part0[28] , 
	\sa_ctrl[5].r.part0[27] , \sa_ctrl[5].r.part0[26] , 
	\sa_ctrl[5].r.part0[25] , \sa_ctrl[5].r.part0[24] , 
	\sa_ctrl[5].r.part0[23] , \sa_ctrl[5].r.part0[22] , 
	\sa_ctrl[5].r.part0[21] , \sa_ctrl[5].r.part0[20] , 
	\sa_ctrl[5].r.part0[19] , \sa_ctrl[5].r.part0[18] , 
	\sa_ctrl[5].r.part0[17] , \sa_ctrl[5].r.part0[16] , 
	\sa_ctrl[5].r.part0[15] , \sa_ctrl[5].r.part0[14] , 
	\sa_ctrl[5].r.part0[13] , \sa_ctrl[5].r.part0[12] , 
	\sa_ctrl[5].r.part0[11] , \sa_ctrl[5].r.part0[10] , 
	\sa_ctrl[5].r.part0[9] , \sa_ctrl[5].r.part0[8] , 
	\sa_ctrl[5].r.part0[7] , \sa_ctrl[5].r.part0[6] , 
	\sa_ctrl[5].r.part0[5] , \sa_ctrl[5].r.part0[4] , 
	\sa_ctrl[5].r.part0[3] , \sa_ctrl[5].r.part0[2] , 
	\sa_ctrl[5].r.part0[1] , \sa_ctrl[5].r.part0[0] , 
	\sa_ctrl[4].r.part0[31] , \sa_ctrl[4].r.part0[30] , 
	\sa_ctrl[4].r.part0[29] , \sa_ctrl[4].r.part0[28] , 
	\sa_ctrl[4].r.part0[27] , \sa_ctrl[4].r.part0[26] , 
	\sa_ctrl[4].r.part0[25] , \sa_ctrl[4].r.part0[24] , 
	\sa_ctrl[4].r.part0[23] , \sa_ctrl[4].r.part0[22] , 
	\sa_ctrl[4].r.part0[21] , \sa_ctrl[4].r.part0[20] , 
	\sa_ctrl[4].r.part0[19] , \sa_ctrl[4].r.part0[18] , 
	\sa_ctrl[4].r.part0[17] , \sa_ctrl[4].r.part0[16] , 
	\sa_ctrl[4].r.part0[15] , \sa_ctrl[4].r.part0[14] , 
	\sa_ctrl[4].r.part0[13] , \sa_ctrl[4].r.part0[12] , 
	\sa_ctrl[4].r.part0[11] , \sa_ctrl[4].r.part0[10] , 
	\sa_ctrl[4].r.part0[9] , \sa_ctrl[4].r.part0[8] , 
	\sa_ctrl[4].r.part0[7] , \sa_ctrl[4].r.part0[6] , 
	\sa_ctrl[4].r.part0[5] , \sa_ctrl[4].r.part0[4] , 
	\sa_ctrl[4].r.part0[3] , \sa_ctrl[4].r.part0[2] , 
	\sa_ctrl[4].r.part0[1] , \sa_ctrl[4].r.part0[0] , 
	\sa_ctrl[3].r.part0[31] , \sa_ctrl[3].r.part0[30] , 
	\sa_ctrl[3].r.part0[29] , \sa_ctrl[3].r.part0[28] , 
	\sa_ctrl[3].r.part0[27] , \sa_ctrl[3].r.part0[26] , 
	\sa_ctrl[3].r.part0[25] , \sa_ctrl[3].r.part0[24] , 
	\sa_ctrl[3].r.part0[23] , \sa_ctrl[3].r.part0[22] , 
	\sa_ctrl[3].r.part0[21] , \sa_ctrl[3].r.part0[20] , 
	\sa_ctrl[3].r.part0[19] , \sa_ctrl[3].r.part0[18] , 
	\sa_ctrl[3].r.part0[17] , \sa_ctrl[3].r.part0[16] , 
	\sa_ctrl[3].r.part0[15] , \sa_ctrl[3].r.part0[14] , 
	\sa_ctrl[3].r.part0[13] , \sa_ctrl[3].r.part0[12] , 
	\sa_ctrl[3].r.part0[11] , \sa_ctrl[3].r.part0[10] , 
	\sa_ctrl[3].r.part0[9] , \sa_ctrl[3].r.part0[8] , 
	\sa_ctrl[3].r.part0[7] , \sa_ctrl[3].r.part0[6] , 
	\sa_ctrl[3].r.part0[5] , \sa_ctrl[3].r.part0[4] , 
	\sa_ctrl[3].r.part0[3] , \sa_ctrl[3].r.part0[2] , 
	\sa_ctrl[3].r.part0[1] , \sa_ctrl[3].r.part0[0] , 
	\sa_ctrl[2].r.part0[31] , \sa_ctrl[2].r.part0[30] , 
	\sa_ctrl[2].r.part0[29] , \sa_ctrl[2].r.part0[28] , 
	\sa_ctrl[2].r.part0[27] , \sa_ctrl[2].r.part0[26] , 
	\sa_ctrl[2].r.part0[25] , \sa_ctrl[2].r.part0[24] , 
	\sa_ctrl[2].r.part0[23] , \sa_ctrl[2].r.part0[22] , 
	\sa_ctrl[2].r.part0[21] , \sa_ctrl[2].r.part0[20] , 
	\sa_ctrl[2].r.part0[19] , \sa_ctrl[2].r.part0[18] , 
	\sa_ctrl[2].r.part0[17] , \sa_ctrl[2].r.part0[16] , 
	\sa_ctrl[2].r.part0[15] , \sa_ctrl[2].r.part0[14] , 
	\sa_ctrl[2].r.part0[13] , \sa_ctrl[2].r.part0[12] , 
	\sa_ctrl[2].r.part0[11] , \sa_ctrl[2].r.part0[10] , 
	\sa_ctrl[2].r.part0[9] , \sa_ctrl[2].r.part0[8] , 
	\sa_ctrl[2].r.part0[7] , \sa_ctrl[2].r.part0[6] , 
	\sa_ctrl[2].r.part0[5] , \sa_ctrl[2].r.part0[4] , 
	\sa_ctrl[2].r.part0[3] , \sa_ctrl[2].r.part0[2] , 
	\sa_ctrl[2].r.part0[1] , \sa_ctrl[2].r.part0[0] , 
	\sa_ctrl[1].r.part0[31] , \sa_ctrl[1].r.part0[30] , 
	\sa_ctrl[1].r.part0[29] , \sa_ctrl[1].r.part0[28] , 
	\sa_ctrl[1].r.part0[27] , \sa_ctrl[1].r.part0[26] , 
	\sa_ctrl[1].r.part0[25] , \sa_ctrl[1].r.part0[24] , 
	\sa_ctrl[1].r.part0[23] , \sa_ctrl[1].r.part0[22] , 
	\sa_ctrl[1].r.part0[21] , \sa_ctrl[1].r.part0[20] , 
	\sa_ctrl[1].r.part0[19] , \sa_ctrl[1].r.part0[18] , 
	\sa_ctrl[1].r.part0[17] , \sa_ctrl[1].r.part0[16] , 
	\sa_ctrl[1].r.part0[15] , \sa_ctrl[1].r.part0[14] , 
	\sa_ctrl[1].r.part0[13] , \sa_ctrl[1].r.part0[12] , 
	\sa_ctrl[1].r.part0[11] , \sa_ctrl[1].r.part0[10] , 
	\sa_ctrl[1].r.part0[9] , \sa_ctrl[1].r.part0[8] , 
	\sa_ctrl[1].r.part0[7] , \sa_ctrl[1].r.part0[6] , 
	\sa_ctrl[1].r.part0[5] , \sa_ctrl[1].r.part0[4] , 
	\sa_ctrl[1].r.part0[3] , \sa_ctrl[1].r.part0[2] , 
	\sa_ctrl[1].r.part0[1] , \sa_ctrl[1].r.part0[0] , 
	\sa_ctrl[0].r.part0[31] , \sa_ctrl[0].r.part0[30] , 
	\sa_ctrl[0].r.part0[29] , \sa_ctrl[0].r.part0[28] , 
	\sa_ctrl[0].r.part0[27] , \sa_ctrl[0].r.part0[26] , 
	\sa_ctrl[0].r.part0[25] , \sa_ctrl[0].r.part0[24] , 
	\sa_ctrl[0].r.part0[23] , \sa_ctrl[0].r.part0[22] , 
	\sa_ctrl[0].r.part0[21] , \sa_ctrl[0].r.part0[20] , 
	\sa_ctrl[0].r.part0[19] , \sa_ctrl[0].r.part0[18] , 
	\sa_ctrl[0].r.part0[17] , \sa_ctrl[0].r.part0[16] , 
	\sa_ctrl[0].r.part0[15] , \sa_ctrl[0].r.part0[14] , 
	\sa_ctrl[0].r.part0[13] , \sa_ctrl[0].r.part0[12] , 
	\sa_ctrl[0].r.part0[11] , \sa_ctrl[0].r.part0[10] , 
	\sa_ctrl[0].r.part0[9] , \sa_ctrl[0].r.part0[8] , 
	\sa_ctrl[0].r.part0[7] , \sa_ctrl[0].r.part0[6] , 
	\sa_ctrl[0].r.part0[5] , \sa_ctrl[0].r.part0[4] , 
	\sa_ctrl[0].r.part0[3] , \sa_ctrl[0].r.part0[2] , 
	\sa_ctrl[0].r.part0[1] , \sa_ctrl[0].r.part0[0] } ), 
	stat_drbg_reseed, stat_req_with_expired_seed, stat_aux_key_type_0, 
	stat_aux_key_type_1, stat_aux_key_type_2, stat_aux_key_type_3, 
	stat_aux_key_type_4, stat_aux_key_type_5, stat_aux_key_type_6, 
	stat_aux_key_type_7, stat_aux_key_type_8, stat_aux_key_type_9, 
	stat_aux_key_type_10, stat_aux_key_type_11, stat_aux_key_type_12, 
	stat_aux_key_type_13, stat_cceip0_stall_on_valid_key, 
	stat_cceip1_stall_on_valid_key, stat_cceip2_stall_on_valid_key, 
	stat_cceip3_stall_on_valid_key, stat_cddip0_stall_on_valid_key, 
	stat_cddip1_stall_on_valid_key, stat_cddip2_stall_on_valid_key, 
	stat_cddip3_stall_on_valid_key, stat_aux_cmd_with_vf_pf_fail, 
	kme_slv_empty, drng_idle, tlv_parser_idle, 
	tlv_parser_int_tlv_start_pulse, cceip_key_tlv_rsm_end_pulse, 
	cddip_key_tlv_rsm_end_pulse, cceip_key_tlv_rsm_idle, 
	cddip_key_tlv_rsm_idle);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output disable_debug_cmd_q;
output set_gcm_tag_fail_int;
output set_txc_bp_int;
output [7:0] set_rsm_is_backpressuring;
output \kme_ib_out.tready ;
wire [0:0] kme_ib_out;
output \sa_snapshot[31].r.part1[31] ,\sa_snapshot[31].r.part1[30] 
	,\sa_snapshot[31].r.part1[29] ,\sa_snapshot[31].r.part1[28] 
	,\sa_snapshot[31].r.part1[27] ,\sa_snapshot[31].r.part1[26] 
	,\sa_snapshot[31].r.part1[25] ,\sa_snapshot[31].r.part1[24] 
	,\sa_snapshot[31].r.part1[23] ,\sa_snapshot[31].r.part1[22] 
	,\sa_snapshot[31].r.part1[21] ,\sa_snapshot[31].r.part1[20] 
	,\sa_snapshot[31].r.part1[19] ,\sa_snapshot[31].r.part1[18] 
	,\sa_snapshot[31].r.part1[17] ,\sa_snapshot[31].r.part1[16] 
	,\sa_snapshot[31].r.part1[15] ,\sa_snapshot[31].r.part1[14] 
	,\sa_snapshot[31].r.part1[13] ,\sa_snapshot[31].r.part1[12] 
	,\sa_snapshot[31].r.part1[11] ,\sa_snapshot[31].r.part1[10] 
	,\sa_snapshot[31].r.part1[9] ,\sa_snapshot[31].r.part1[8] 
	,\sa_snapshot[31].r.part1[7] ,\sa_snapshot[31].r.part1[6] 
	,\sa_snapshot[31].r.part1[5] ,\sa_snapshot[31].r.part1[4] 
	,\sa_snapshot[31].r.part1[3] ,\sa_snapshot[31].r.part1[2] 
	,\sa_snapshot[31].r.part1[1] ,\sa_snapshot[31].r.part1[0] 
	,\sa_snapshot[31].r.part0[31] ,\sa_snapshot[31].r.part0[30] 
	,\sa_snapshot[31].r.part0[29] ,\sa_snapshot[31].r.part0[28] 
	,\sa_snapshot[31].r.part0[27] ,\sa_snapshot[31].r.part0[26] 
	,\sa_snapshot[31].r.part0[25] ,\sa_snapshot[31].r.part0[24] 
	,\sa_snapshot[31].r.part0[23] ,\sa_snapshot[31].r.part0[22] 
	,\sa_snapshot[31].r.part0[21] ,\sa_snapshot[31].r.part0[20] 
	,\sa_snapshot[31].r.part0[19] ,\sa_snapshot[31].r.part0[18] 
	,\sa_snapshot[31].r.part0[17] ,\sa_snapshot[31].r.part0[16] 
	,\sa_snapshot[31].r.part0[15] ,\sa_snapshot[31].r.part0[14] 
	,\sa_snapshot[31].r.part0[13] ,\sa_snapshot[31].r.part0[12] 
	,\sa_snapshot[31].r.part0[11] ,\sa_snapshot[31].r.part0[10] 
	,\sa_snapshot[31].r.part0[9] ,\sa_snapshot[31].r.part0[8] 
	,\sa_snapshot[31].r.part0[7] ,\sa_snapshot[31].r.part0[6] 
	,\sa_snapshot[31].r.part0[5] ,\sa_snapshot[31].r.part0[4] 
	,\sa_snapshot[31].r.part0[3] ,\sa_snapshot[31].r.part0[2] 
	,\sa_snapshot[31].r.part0[1] ,\sa_snapshot[31].r.part0[0] 
	,\sa_snapshot[30].r.part1[31] ,\sa_snapshot[30].r.part1[30] 
	,\sa_snapshot[30].r.part1[29] ,\sa_snapshot[30].r.part1[28] 
	,\sa_snapshot[30].r.part1[27] ,\sa_snapshot[30].r.part1[26] 
	,\sa_snapshot[30].r.part1[25] ,\sa_snapshot[30].r.part1[24] 
	,\sa_snapshot[30].r.part1[23] ,\sa_snapshot[30].r.part1[22] 
	,\sa_snapshot[30].r.part1[21] ,\sa_snapshot[30].r.part1[20] 
	,\sa_snapshot[30].r.part1[19] ,\sa_snapshot[30].r.part1[18] 
	,\sa_snapshot[30].r.part1[17] ,\sa_snapshot[30].r.part1[16] 
	,\sa_snapshot[30].r.part1[15] ,\sa_snapshot[30].r.part1[14] 
	,\sa_snapshot[30].r.part1[13] ,\sa_snapshot[30].r.part1[12] 
	,\sa_snapshot[30].r.part1[11] ,\sa_snapshot[30].r.part1[10] 
	,\sa_snapshot[30].r.part1[9] ,\sa_snapshot[30].r.part1[8] 
	,\sa_snapshot[30].r.part1[7] ,\sa_snapshot[30].r.part1[6] 
	,\sa_snapshot[30].r.part1[5] ,\sa_snapshot[30].r.part1[4] 
	,\sa_snapshot[30].r.part1[3] ,\sa_snapshot[30].r.part1[2] 
	,\sa_snapshot[30].r.part1[1] ,\sa_snapshot[30].r.part1[0] 
	,\sa_snapshot[30].r.part0[31] ,\sa_snapshot[30].r.part0[30] 
	,\sa_snapshot[30].r.part0[29] ,\sa_snapshot[30].r.part0[28] 
	,\sa_snapshot[30].r.part0[27] ,\sa_snapshot[30].r.part0[26] 
	,\sa_snapshot[30].r.part0[25] ,\sa_snapshot[30].r.part0[24] 
	,\sa_snapshot[30].r.part0[23] ,\sa_snapshot[30].r.part0[22] 
	,\sa_snapshot[30].r.part0[21] ,\sa_snapshot[30].r.part0[20] 
	,\sa_snapshot[30].r.part0[19] ,\sa_snapshot[30].r.part0[18] 
	,\sa_snapshot[30].r.part0[17] ,\sa_snapshot[30].r.part0[16] 
	,\sa_snapshot[30].r.part0[15] ,\sa_snapshot[30].r.part0[14] 
	,\sa_snapshot[30].r.part0[13] ,\sa_snapshot[30].r.part0[12] 
	,\sa_snapshot[30].r.part0[11] ,\sa_snapshot[30].r.part0[10] 
	,\sa_snapshot[30].r.part0[9] ,\sa_snapshot[30].r.part0[8] 
	,\sa_snapshot[30].r.part0[7] ,\sa_snapshot[30].r.part0[6] 
	,\sa_snapshot[30].r.part0[5] ,\sa_snapshot[30].r.part0[4] 
	,\sa_snapshot[30].r.part0[3] ,\sa_snapshot[30].r.part0[2] 
	,\sa_snapshot[30].r.part0[1] ,\sa_snapshot[30].r.part0[0] 
	,\sa_snapshot[29].r.part1[31] ,\sa_snapshot[29].r.part1[30] 
	,\sa_snapshot[29].r.part1[29] ,\sa_snapshot[29].r.part1[28] 
	,\sa_snapshot[29].r.part1[27] ,\sa_snapshot[29].r.part1[26] 
	,\sa_snapshot[29].r.part1[25] ,\sa_snapshot[29].r.part1[24] 
	,\sa_snapshot[29].r.part1[23] ,\sa_snapshot[29].r.part1[22] 
	,\sa_snapshot[29].r.part1[21] ,\sa_snapshot[29].r.part1[20] 
	,\sa_snapshot[29].r.part1[19] ,\sa_snapshot[29].r.part1[18] 
	,\sa_snapshot[29].r.part1[17] ,\sa_snapshot[29].r.part1[16] 
	,\sa_snapshot[29].r.part1[15] ,\sa_snapshot[29].r.part1[14] 
	,\sa_snapshot[29].r.part1[13] ,\sa_snapshot[29].r.part1[12] 
	,\sa_snapshot[29].r.part1[11] ,\sa_snapshot[29].r.part1[10] 
	,\sa_snapshot[29].r.part1[9] ,\sa_snapshot[29].r.part1[8] 
	,\sa_snapshot[29].r.part1[7] ,\sa_snapshot[29].r.part1[6] 
	,\sa_snapshot[29].r.part1[5] ,\sa_snapshot[29].r.part1[4] 
	,\sa_snapshot[29].r.part1[3] ,\sa_snapshot[29].r.part1[2] 
	,\sa_snapshot[29].r.part1[1] ,\sa_snapshot[29].r.part1[0] 
	,\sa_snapshot[29].r.part0[31] ,\sa_snapshot[29].r.part0[30] 
	,\sa_snapshot[29].r.part0[29] ,\sa_snapshot[29].r.part0[28] 
	,\sa_snapshot[29].r.part0[27] ,\sa_snapshot[29].r.part0[26] 
	,\sa_snapshot[29].r.part0[25] ,\sa_snapshot[29].r.part0[24] 
	,\sa_snapshot[29].r.part0[23] ,\sa_snapshot[29].r.part0[22] 
	,\sa_snapshot[29].r.part0[21] ,\sa_snapshot[29].r.part0[20] 
	,\sa_snapshot[29].r.part0[19] ,\sa_snapshot[29].r.part0[18] 
	,\sa_snapshot[29].r.part0[17] ,\sa_snapshot[29].r.part0[16] 
	,\sa_snapshot[29].r.part0[15] ,\sa_snapshot[29].r.part0[14] 
	,\sa_snapshot[29].r.part0[13] ,\sa_snapshot[29].r.part0[12] 
	,\sa_snapshot[29].r.part0[11] ,\sa_snapshot[29].r.part0[10] 
	,\sa_snapshot[29].r.part0[9] ,\sa_snapshot[29].r.part0[8] 
	,\sa_snapshot[29].r.part0[7] ,\sa_snapshot[29].r.part0[6] 
	,\sa_snapshot[29].r.part0[5] ,\sa_snapshot[29].r.part0[4] 
	,\sa_snapshot[29].r.part0[3] ,\sa_snapshot[29].r.part0[2] 
	,\sa_snapshot[29].r.part0[1] ,\sa_snapshot[29].r.part0[0] 
	,\sa_snapshot[28].r.part1[31] ,\sa_snapshot[28].r.part1[30] 
	,\sa_snapshot[28].r.part1[29] ,\sa_snapshot[28].r.part1[28] 
	,\sa_snapshot[28].r.part1[27] ,\sa_snapshot[28].r.part1[26] 
	,\sa_snapshot[28].r.part1[25] ,\sa_snapshot[28].r.part1[24] 
	,\sa_snapshot[28].r.part1[23] ,\sa_snapshot[28].r.part1[22] 
	,\sa_snapshot[28].r.part1[21] ,\sa_snapshot[28].r.part1[20] 
	,\sa_snapshot[28].r.part1[19] ,\sa_snapshot[28].r.part1[18] 
	,\sa_snapshot[28].r.part1[17] ,\sa_snapshot[28].r.part1[16] 
	,\sa_snapshot[28].r.part1[15] ,\sa_snapshot[28].r.part1[14] 
	,\sa_snapshot[28].r.part1[13] ,\sa_snapshot[28].r.part1[12] 
	,\sa_snapshot[28].r.part1[11] ,\sa_snapshot[28].r.part1[10] 
	,\sa_snapshot[28].r.part1[9] ,\sa_snapshot[28].r.part1[8] 
	,\sa_snapshot[28].r.part1[7] ,\sa_snapshot[28].r.part1[6] 
	,\sa_snapshot[28].r.part1[5] ,\sa_snapshot[28].r.part1[4] 
	,\sa_snapshot[28].r.part1[3] ,\sa_snapshot[28].r.part1[2] 
	,\sa_snapshot[28].r.part1[1] ,\sa_snapshot[28].r.part1[0] 
	,\sa_snapshot[28].r.part0[31] ,\sa_snapshot[28].r.part0[30] 
	,\sa_snapshot[28].r.part0[29] ,\sa_snapshot[28].r.part0[28] 
	,\sa_snapshot[28].r.part0[27] ,\sa_snapshot[28].r.part0[26] 
	,\sa_snapshot[28].r.part0[25] ,\sa_snapshot[28].r.part0[24] 
	,\sa_snapshot[28].r.part0[23] ,\sa_snapshot[28].r.part0[22] 
	,\sa_snapshot[28].r.part0[21] ,\sa_snapshot[28].r.part0[20] 
	,\sa_snapshot[28].r.part0[19] ,\sa_snapshot[28].r.part0[18] 
	,\sa_snapshot[28].r.part0[17] ,\sa_snapshot[28].r.part0[16] 
	,\sa_snapshot[28].r.part0[15] ,\sa_snapshot[28].r.part0[14] 
	,\sa_snapshot[28].r.part0[13] ,\sa_snapshot[28].r.part0[12] 
	,\sa_snapshot[28].r.part0[11] ,\sa_snapshot[28].r.part0[10] 
	,\sa_snapshot[28].r.part0[9] ,\sa_snapshot[28].r.part0[8] 
	,\sa_snapshot[28].r.part0[7] ,\sa_snapshot[28].r.part0[6] 
	,\sa_snapshot[28].r.part0[5] ,\sa_snapshot[28].r.part0[4] 
	,\sa_snapshot[28].r.part0[3] ,\sa_snapshot[28].r.part0[2] 
	,\sa_snapshot[28].r.part0[1] ,\sa_snapshot[28].r.part0[0] 
	,\sa_snapshot[27].r.part1[31] ,\sa_snapshot[27].r.part1[30] 
	,\sa_snapshot[27].r.part1[29] ,\sa_snapshot[27].r.part1[28] 
	,\sa_snapshot[27].r.part1[27] ,\sa_snapshot[27].r.part1[26] 
	,\sa_snapshot[27].r.part1[25] ,\sa_snapshot[27].r.part1[24] 
	,\sa_snapshot[27].r.part1[23] ,\sa_snapshot[27].r.part1[22] 
	,\sa_snapshot[27].r.part1[21] ,\sa_snapshot[27].r.part1[20] 
	,\sa_snapshot[27].r.part1[19] ,\sa_snapshot[27].r.part1[18] 
	,\sa_snapshot[27].r.part1[17] ,\sa_snapshot[27].r.part1[16] 
	,\sa_snapshot[27].r.part1[15] ,\sa_snapshot[27].r.part1[14] 
	,\sa_snapshot[27].r.part1[13] ,\sa_snapshot[27].r.part1[12] 
	,\sa_snapshot[27].r.part1[11] ,\sa_snapshot[27].r.part1[10] 
	,\sa_snapshot[27].r.part1[9] ,\sa_snapshot[27].r.part1[8] 
	,\sa_snapshot[27].r.part1[7] ,\sa_snapshot[27].r.part1[6] 
	,\sa_snapshot[27].r.part1[5] ,\sa_snapshot[27].r.part1[4] 
	,\sa_snapshot[27].r.part1[3] ,\sa_snapshot[27].r.part1[2] 
	,\sa_snapshot[27].r.part1[1] ,\sa_snapshot[27].r.part1[0] 
	,\sa_snapshot[27].r.part0[31] ,\sa_snapshot[27].r.part0[30] 
	,\sa_snapshot[27].r.part0[29] ,\sa_snapshot[27].r.part0[28] 
	,\sa_snapshot[27].r.part0[27] ,\sa_snapshot[27].r.part0[26] 
	,\sa_snapshot[27].r.part0[25] ,\sa_snapshot[27].r.part0[24] 
	,\sa_snapshot[27].r.part0[23] ,\sa_snapshot[27].r.part0[22] 
	,\sa_snapshot[27].r.part0[21] ,\sa_snapshot[27].r.part0[20] 
	,\sa_snapshot[27].r.part0[19] ,\sa_snapshot[27].r.part0[18] 
	,\sa_snapshot[27].r.part0[17] ,\sa_snapshot[27].r.part0[16] 
	,\sa_snapshot[27].r.part0[15] ,\sa_snapshot[27].r.part0[14] 
	,\sa_snapshot[27].r.part0[13] ,\sa_snapshot[27].r.part0[12] 
	,\sa_snapshot[27].r.part0[11] ,\sa_snapshot[27].r.part0[10] 
	,\sa_snapshot[27].r.part0[9] ,\sa_snapshot[27].r.part0[8] 
	,\sa_snapshot[27].r.part0[7] ,\sa_snapshot[27].r.part0[6] 
	,\sa_snapshot[27].r.part0[5] ,\sa_snapshot[27].r.part0[4] 
	,\sa_snapshot[27].r.part0[3] ,\sa_snapshot[27].r.part0[2] 
	,\sa_snapshot[27].r.part0[1] ,\sa_snapshot[27].r.part0[0] 
	,\sa_snapshot[26].r.part1[31] ,\sa_snapshot[26].r.part1[30] 
	,\sa_snapshot[26].r.part1[29] ,\sa_snapshot[26].r.part1[28] 
	,\sa_snapshot[26].r.part1[27] ,\sa_snapshot[26].r.part1[26] 
	,\sa_snapshot[26].r.part1[25] ,\sa_snapshot[26].r.part1[24] 
	,\sa_snapshot[26].r.part1[23] ,\sa_snapshot[26].r.part1[22] 
	,\sa_snapshot[26].r.part1[21] ,\sa_snapshot[26].r.part1[20] 
	,\sa_snapshot[26].r.part1[19] ,\sa_snapshot[26].r.part1[18] 
	,\sa_snapshot[26].r.part1[17] ,\sa_snapshot[26].r.part1[16] 
	,\sa_snapshot[26].r.part1[15] ,\sa_snapshot[26].r.part1[14] 
	,\sa_snapshot[26].r.part1[13] ,\sa_snapshot[26].r.part1[12] 
	,\sa_snapshot[26].r.part1[11] ,\sa_snapshot[26].r.part1[10] 
	,\sa_snapshot[26].r.part1[9] ,\sa_snapshot[26].r.part1[8] 
	,\sa_snapshot[26].r.part1[7] ,\sa_snapshot[26].r.part1[6] 
	,\sa_snapshot[26].r.part1[5] ,\sa_snapshot[26].r.part1[4] 
	,\sa_snapshot[26].r.part1[3] ,\sa_snapshot[26].r.part1[2] 
	,\sa_snapshot[26].r.part1[1] ,\sa_snapshot[26].r.part1[0] 
	,\sa_snapshot[26].r.part0[31] ,\sa_snapshot[26].r.part0[30] 
	,\sa_snapshot[26].r.part0[29] ,\sa_snapshot[26].r.part0[28] 
	,\sa_snapshot[26].r.part0[27] ,\sa_snapshot[26].r.part0[26] 
	,\sa_snapshot[26].r.part0[25] ,\sa_snapshot[26].r.part0[24] 
	,\sa_snapshot[26].r.part0[23] ,\sa_snapshot[26].r.part0[22] 
	,\sa_snapshot[26].r.part0[21] ,\sa_snapshot[26].r.part0[20] 
	,\sa_snapshot[26].r.part0[19] ,\sa_snapshot[26].r.part0[18] 
	,\sa_snapshot[26].r.part0[17] ,\sa_snapshot[26].r.part0[16] 
	,\sa_snapshot[26].r.part0[15] ,\sa_snapshot[26].r.part0[14] 
	,\sa_snapshot[26].r.part0[13] ,\sa_snapshot[26].r.part0[12] 
	,\sa_snapshot[26].r.part0[11] ,\sa_snapshot[26].r.part0[10] 
	,\sa_snapshot[26].r.part0[9] ,\sa_snapshot[26].r.part0[8] 
	,\sa_snapshot[26].r.part0[7] ,\sa_snapshot[26].r.part0[6] 
	,\sa_snapshot[26].r.part0[5] ,\sa_snapshot[26].r.part0[4] 
	,\sa_snapshot[26].r.part0[3] ,\sa_snapshot[26].r.part0[2] 
	,\sa_snapshot[26].r.part0[1] ,\sa_snapshot[26].r.part0[0] 
	,\sa_snapshot[25].r.part1[31] ,\sa_snapshot[25].r.part1[30] 
	,\sa_snapshot[25].r.part1[29] ,\sa_snapshot[25].r.part1[28] 
	,\sa_snapshot[25].r.part1[27] ,\sa_snapshot[25].r.part1[26] 
	,\sa_snapshot[25].r.part1[25] ,\sa_snapshot[25].r.part1[24] 
	,\sa_snapshot[25].r.part1[23] ,\sa_snapshot[25].r.part1[22] 
	,\sa_snapshot[25].r.part1[21] ,\sa_snapshot[25].r.part1[20] 
	,\sa_snapshot[25].r.part1[19] ,\sa_snapshot[25].r.part1[18] 
	,\sa_snapshot[25].r.part1[17] ,\sa_snapshot[25].r.part1[16] 
	,\sa_snapshot[25].r.part1[15] ,\sa_snapshot[25].r.part1[14] 
	,\sa_snapshot[25].r.part1[13] ,\sa_snapshot[25].r.part1[12] 
	,\sa_snapshot[25].r.part1[11] ,\sa_snapshot[25].r.part1[10] 
	,\sa_snapshot[25].r.part1[9] ,\sa_snapshot[25].r.part1[8] 
	,\sa_snapshot[25].r.part1[7] ,\sa_snapshot[25].r.part1[6] 
	,\sa_snapshot[25].r.part1[5] ,\sa_snapshot[25].r.part1[4] 
	,\sa_snapshot[25].r.part1[3] ,\sa_snapshot[25].r.part1[2] 
	,\sa_snapshot[25].r.part1[1] ,\sa_snapshot[25].r.part1[0] 
	,\sa_snapshot[25].r.part0[31] ,\sa_snapshot[25].r.part0[30] 
	,\sa_snapshot[25].r.part0[29] ,\sa_snapshot[25].r.part0[28] 
	,\sa_snapshot[25].r.part0[27] ,\sa_snapshot[25].r.part0[26] 
	,\sa_snapshot[25].r.part0[25] ,\sa_snapshot[25].r.part0[24] 
	,\sa_snapshot[25].r.part0[23] ,\sa_snapshot[25].r.part0[22] 
	,\sa_snapshot[25].r.part0[21] ,\sa_snapshot[25].r.part0[20] 
	,\sa_snapshot[25].r.part0[19] ,\sa_snapshot[25].r.part0[18] 
	,\sa_snapshot[25].r.part0[17] ,\sa_snapshot[25].r.part0[16] 
	,\sa_snapshot[25].r.part0[15] ,\sa_snapshot[25].r.part0[14] 
	,\sa_snapshot[25].r.part0[13] ,\sa_snapshot[25].r.part0[12] 
	,\sa_snapshot[25].r.part0[11] ,\sa_snapshot[25].r.part0[10] 
	,\sa_snapshot[25].r.part0[9] ,\sa_snapshot[25].r.part0[8] 
	,\sa_snapshot[25].r.part0[7] ,\sa_snapshot[25].r.part0[6] 
	,\sa_snapshot[25].r.part0[5] ,\sa_snapshot[25].r.part0[4] 
	,\sa_snapshot[25].r.part0[3] ,\sa_snapshot[25].r.part0[2] 
	,\sa_snapshot[25].r.part0[1] ,\sa_snapshot[25].r.part0[0] 
	,\sa_snapshot[24].r.part1[31] ,\sa_snapshot[24].r.part1[30] 
	,\sa_snapshot[24].r.part1[29] ,\sa_snapshot[24].r.part1[28] 
	,\sa_snapshot[24].r.part1[27] ,\sa_snapshot[24].r.part1[26] 
	,\sa_snapshot[24].r.part1[25] ,\sa_snapshot[24].r.part1[24] 
	,\sa_snapshot[24].r.part1[23] ,\sa_snapshot[24].r.part1[22] 
	,\sa_snapshot[24].r.part1[21] ,\sa_snapshot[24].r.part1[20] 
	,\sa_snapshot[24].r.part1[19] ,\sa_snapshot[24].r.part1[18] 
	,\sa_snapshot[24].r.part1[17] ,\sa_snapshot[24].r.part1[16] 
	,\sa_snapshot[24].r.part1[15] ,\sa_snapshot[24].r.part1[14] 
	,\sa_snapshot[24].r.part1[13] ,\sa_snapshot[24].r.part1[12] 
	,\sa_snapshot[24].r.part1[11] ,\sa_snapshot[24].r.part1[10] 
	,\sa_snapshot[24].r.part1[9] ,\sa_snapshot[24].r.part1[8] 
	,\sa_snapshot[24].r.part1[7] ,\sa_snapshot[24].r.part1[6] 
	,\sa_snapshot[24].r.part1[5] ,\sa_snapshot[24].r.part1[4] 
	,\sa_snapshot[24].r.part1[3] ,\sa_snapshot[24].r.part1[2] 
	,\sa_snapshot[24].r.part1[1] ,\sa_snapshot[24].r.part1[0] 
	,\sa_snapshot[24].r.part0[31] ,\sa_snapshot[24].r.part0[30] 
	,\sa_snapshot[24].r.part0[29] ,\sa_snapshot[24].r.part0[28] 
	,\sa_snapshot[24].r.part0[27] ,\sa_snapshot[24].r.part0[26] 
	,\sa_snapshot[24].r.part0[25] ,\sa_snapshot[24].r.part0[24] 
	,\sa_snapshot[24].r.part0[23] ,\sa_snapshot[24].r.part0[22] 
	,\sa_snapshot[24].r.part0[21] ,\sa_snapshot[24].r.part0[20] 
	,\sa_snapshot[24].r.part0[19] ,\sa_snapshot[24].r.part0[18] 
	,\sa_snapshot[24].r.part0[17] ,\sa_snapshot[24].r.part0[16] 
	,\sa_snapshot[24].r.part0[15] ,\sa_snapshot[24].r.part0[14] 
	,\sa_snapshot[24].r.part0[13] ,\sa_snapshot[24].r.part0[12] 
	,\sa_snapshot[24].r.part0[11] ,\sa_snapshot[24].r.part0[10] 
	,\sa_snapshot[24].r.part0[9] ,\sa_snapshot[24].r.part0[8] 
	,\sa_snapshot[24].r.part0[7] ,\sa_snapshot[24].r.part0[6] 
	,\sa_snapshot[24].r.part0[5] ,\sa_snapshot[24].r.part0[4] 
	,\sa_snapshot[24].r.part0[3] ,\sa_snapshot[24].r.part0[2] 
	,\sa_snapshot[24].r.part0[1] ,\sa_snapshot[24].r.part0[0] 
	,\sa_snapshot[23].r.part1[31] ,\sa_snapshot[23].r.part1[30] 
	,\sa_snapshot[23].r.part1[29] ,\sa_snapshot[23].r.part1[28] 
	,\sa_snapshot[23].r.part1[27] ,\sa_snapshot[23].r.part1[26] 
	,\sa_snapshot[23].r.part1[25] ,\sa_snapshot[23].r.part1[24] 
	,\sa_snapshot[23].r.part1[23] ,\sa_snapshot[23].r.part1[22] 
	,\sa_snapshot[23].r.part1[21] ,\sa_snapshot[23].r.part1[20] 
	,\sa_snapshot[23].r.part1[19] ,\sa_snapshot[23].r.part1[18] 
	,\sa_snapshot[23].r.part1[17] ,\sa_snapshot[23].r.part1[16] 
	,\sa_snapshot[23].r.part1[15] ,\sa_snapshot[23].r.part1[14] 
	,\sa_snapshot[23].r.part1[13] ,\sa_snapshot[23].r.part1[12] 
	,\sa_snapshot[23].r.part1[11] ,\sa_snapshot[23].r.part1[10] 
	,\sa_snapshot[23].r.part1[9] ,\sa_snapshot[23].r.part1[8] 
	,\sa_snapshot[23].r.part1[7] ,\sa_snapshot[23].r.part1[6] 
	,\sa_snapshot[23].r.part1[5] ,\sa_snapshot[23].r.part1[4] 
	,\sa_snapshot[23].r.part1[3] ,\sa_snapshot[23].r.part1[2] 
	,\sa_snapshot[23].r.part1[1] ,\sa_snapshot[23].r.part1[0] 
	,\sa_snapshot[23].r.part0[31] ,\sa_snapshot[23].r.part0[30] 
	,\sa_snapshot[23].r.part0[29] ,\sa_snapshot[23].r.part0[28] 
	,\sa_snapshot[23].r.part0[27] ,\sa_snapshot[23].r.part0[26] 
	,\sa_snapshot[23].r.part0[25] ,\sa_snapshot[23].r.part0[24] 
	,\sa_snapshot[23].r.part0[23] ,\sa_snapshot[23].r.part0[22] 
	,\sa_snapshot[23].r.part0[21] ,\sa_snapshot[23].r.part0[20] 
	,\sa_snapshot[23].r.part0[19] ,\sa_snapshot[23].r.part0[18] 
	,\sa_snapshot[23].r.part0[17] ,\sa_snapshot[23].r.part0[16] 
	,\sa_snapshot[23].r.part0[15] ,\sa_snapshot[23].r.part0[14] 
	,\sa_snapshot[23].r.part0[13] ,\sa_snapshot[23].r.part0[12] 
	,\sa_snapshot[23].r.part0[11] ,\sa_snapshot[23].r.part0[10] 
	,\sa_snapshot[23].r.part0[9] ,\sa_snapshot[23].r.part0[8] 
	,\sa_snapshot[23].r.part0[7] ,\sa_snapshot[23].r.part0[6] 
	,\sa_snapshot[23].r.part0[5] ,\sa_snapshot[23].r.part0[4] 
	,\sa_snapshot[23].r.part0[3] ,\sa_snapshot[23].r.part0[2] 
	,\sa_snapshot[23].r.part0[1] ,\sa_snapshot[23].r.part0[0] 
	,\sa_snapshot[22].r.part1[31] ,\sa_snapshot[22].r.part1[30] 
	,\sa_snapshot[22].r.part1[29] ,\sa_snapshot[22].r.part1[28] 
	,\sa_snapshot[22].r.part1[27] ,\sa_snapshot[22].r.part1[26] 
	,\sa_snapshot[22].r.part1[25] ,\sa_snapshot[22].r.part1[24] 
	,\sa_snapshot[22].r.part1[23] ,\sa_snapshot[22].r.part1[22] 
	,\sa_snapshot[22].r.part1[21] ,\sa_snapshot[22].r.part1[20] 
	,\sa_snapshot[22].r.part1[19] ,\sa_snapshot[22].r.part1[18] 
	,\sa_snapshot[22].r.part1[17] ,\sa_snapshot[22].r.part1[16] 
	,\sa_snapshot[22].r.part1[15] ,\sa_snapshot[22].r.part1[14] 
	,\sa_snapshot[22].r.part1[13] ,\sa_snapshot[22].r.part1[12] 
	,\sa_snapshot[22].r.part1[11] ,\sa_snapshot[22].r.part1[10] 
	,\sa_snapshot[22].r.part1[9] ,\sa_snapshot[22].r.part1[8] 
	,\sa_snapshot[22].r.part1[7] ,\sa_snapshot[22].r.part1[6] 
	,\sa_snapshot[22].r.part1[5] ,\sa_snapshot[22].r.part1[4] 
	,\sa_snapshot[22].r.part1[3] ,\sa_snapshot[22].r.part1[2] 
	,\sa_snapshot[22].r.part1[1] ,\sa_snapshot[22].r.part1[0] 
	,\sa_snapshot[22].r.part0[31] ,\sa_snapshot[22].r.part0[30] 
	,\sa_snapshot[22].r.part0[29] ,\sa_snapshot[22].r.part0[28] 
	,\sa_snapshot[22].r.part0[27] ,\sa_snapshot[22].r.part0[26] 
	,\sa_snapshot[22].r.part0[25] ,\sa_snapshot[22].r.part0[24] 
	,\sa_snapshot[22].r.part0[23] ,\sa_snapshot[22].r.part0[22] 
	,\sa_snapshot[22].r.part0[21] ,\sa_snapshot[22].r.part0[20] 
	,\sa_snapshot[22].r.part0[19] ,\sa_snapshot[22].r.part0[18] 
	,\sa_snapshot[22].r.part0[17] ,\sa_snapshot[22].r.part0[16] 
	,\sa_snapshot[22].r.part0[15] ,\sa_snapshot[22].r.part0[14] 
	,\sa_snapshot[22].r.part0[13] ,\sa_snapshot[22].r.part0[12] 
	,\sa_snapshot[22].r.part0[11] ,\sa_snapshot[22].r.part0[10] 
	,\sa_snapshot[22].r.part0[9] ,\sa_snapshot[22].r.part0[8] 
	,\sa_snapshot[22].r.part0[7] ,\sa_snapshot[22].r.part0[6] 
	,\sa_snapshot[22].r.part0[5] ,\sa_snapshot[22].r.part0[4] 
	,\sa_snapshot[22].r.part0[3] ,\sa_snapshot[22].r.part0[2] 
	,\sa_snapshot[22].r.part0[1] ,\sa_snapshot[22].r.part0[0] 
	,\sa_snapshot[21].r.part1[31] ,\sa_snapshot[21].r.part1[30] 
	,\sa_snapshot[21].r.part1[29] ,\sa_snapshot[21].r.part1[28] 
	,\sa_snapshot[21].r.part1[27] ,\sa_snapshot[21].r.part1[26] 
	,\sa_snapshot[21].r.part1[25] ,\sa_snapshot[21].r.part1[24] 
	,\sa_snapshot[21].r.part1[23] ,\sa_snapshot[21].r.part1[22] 
	,\sa_snapshot[21].r.part1[21] ,\sa_snapshot[21].r.part1[20] 
	,\sa_snapshot[21].r.part1[19] ,\sa_snapshot[21].r.part1[18] 
	,\sa_snapshot[21].r.part1[17] ,\sa_snapshot[21].r.part1[16] 
	,\sa_snapshot[21].r.part1[15] ,\sa_snapshot[21].r.part1[14] 
	,\sa_snapshot[21].r.part1[13] ,\sa_snapshot[21].r.part1[12] 
	,\sa_snapshot[21].r.part1[11] ,\sa_snapshot[21].r.part1[10] 
	,\sa_snapshot[21].r.part1[9] ,\sa_snapshot[21].r.part1[8] 
	,\sa_snapshot[21].r.part1[7] ,\sa_snapshot[21].r.part1[6] 
	,\sa_snapshot[21].r.part1[5] ,\sa_snapshot[21].r.part1[4] 
	,\sa_snapshot[21].r.part1[3] ,\sa_snapshot[21].r.part1[2] 
	,\sa_snapshot[21].r.part1[1] ,\sa_snapshot[21].r.part1[0] 
	,\sa_snapshot[21].r.part0[31] ,\sa_snapshot[21].r.part0[30] 
	,\sa_snapshot[21].r.part0[29] ,\sa_snapshot[21].r.part0[28] 
	,\sa_snapshot[21].r.part0[27] ,\sa_snapshot[21].r.part0[26] 
	,\sa_snapshot[21].r.part0[25] ,\sa_snapshot[21].r.part0[24] 
	,\sa_snapshot[21].r.part0[23] ,\sa_snapshot[21].r.part0[22] 
	,\sa_snapshot[21].r.part0[21] ,\sa_snapshot[21].r.part0[20] 
	,\sa_snapshot[21].r.part0[19] ,\sa_snapshot[21].r.part0[18] 
	,\sa_snapshot[21].r.part0[17] ,\sa_snapshot[21].r.part0[16] 
	,\sa_snapshot[21].r.part0[15] ,\sa_snapshot[21].r.part0[14] 
	,\sa_snapshot[21].r.part0[13] ,\sa_snapshot[21].r.part0[12] 
	,\sa_snapshot[21].r.part0[11] ,\sa_snapshot[21].r.part0[10] 
	,\sa_snapshot[21].r.part0[9] ,\sa_snapshot[21].r.part0[8] 
	,\sa_snapshot[21].r.part0[7] ,\sa_snapshot[21].r.part0[6] 
	,\sa_snapshot[21].r.part0[5] ,\sa_snapshot[21].r.part0[4] 
	,\sa_snapshot[21].r.part0[3] ,\sa_snapshot[21].r.part0[2] 
	,\sa_snapshot[21].r.part0[1] ,\sa_snapshot[21].r.part0[0] 
	,\sa_snapshot[20].r.part1[31] ,\sa_snapshot[20].r.part1[30] 
	,\sa_snapshot[20].r.part1[29] ,\sa_snapshot[20].r.part1[28] 
	,\sa_snapshot[20].r.part1[27] ,\sa_snapshot[20].r.part1[26] 
	,\sa_snapshot[20].r.part1[25] ,\sa_snapshot[20].r.part1[24] 
	,\sa_snapshot[20].r.part1[23] ,\sa_snapshot[20].r.part1[22] 
	,\sa_snapshot[20].r.part1[21] ,\sa_snapshot[20].r.part1[20] 
	,\sa_snapshot[20].r.part1[19] ,\sa_snapshot[20].r.part1[18] 
	,\sa_snapshot[20].r.part1[17] ,\sa_snapshot[20].r.part1[16] 
	,\sa_snapshot[20].r.part1[15] ,\sa_snapshot[20].r.part1[14] 
	,\sa_snapshot[20].r.part1[13] ,\sa_snapshot[20].r.part1[12] 
	,\sa_snapshot[20].r.part1[11] ,\sa_snapshot[20].r.part1[10] 
	,\sa_snapshot[20].r.part1[9] ,\sa_snapshot[20].r.part1[8] 
	,\sa_snapshot[20].r.part1[7] ,\sa_snapshot[20].r.part1[6] 
	,\sa_snapshot[20].r.part1[5] ,\sa_snapshot[20].r.part1[4] 
	,\sa_snapshot[20].r.part1[3] ,\sa_snapshot[20].r.part1[2] 
	,\sa_snapshot[20].r.part1[1] ,\sa_snapshot[20].r.part1[0] 
	,\sa_snapshot[20].r.part0[31] ,\sa_snapshot[20].r.part0[30] 
	,\sa_snapshot[20].r.part0[29] ,\sa_snapshot[20].r.part0[28] 
	,\sa_snapshot[20].r.part0[27] ,\sa_snapshot[20].r.part0[26] 
	,\sa_snapshot[20].r.part0[25] ,\sa_snapshot[20].r.part0[24] 
	,\sa_snapshot[20].r.part0[23] ,\sa_snapshot[20].r.part0[22] 
	,\sa_snapshot[20].r.part0[21] ,\sa_snapshot[20].r.part0[20] 
	,\sa_snapshot[20].r.part0[19] ,\sa_snapshot[20].r.part0[18] 
	,\sa_snapshot[20].r.part0[17] ,\sa_snapshot[20].r.part0[16] 
	,\sa_snapshot[20].r.part0[15] ,\sa_snapshot[20].r.part0[14] 
	,\sa_snapshot[20].r.part0[13] ,\sa_snapshot[20].r.part0[12] 
	,\sa_snapshot[20].r.part0[11] ,\sa_snapshot[20].r.part0[10] 
	,\sa_snapshot[20].r.part0[9] ,\sa_snapshot[20].r.part0[8] 
	,\sa_snapshot[20].r.part0[7] ,\sa_snapshot[20].r.part0[6] 
	,\sa_snapshot[20].r.part0[5] ,\sa_snapshot[20].r.part0[4] 
	,\sa_snapshot[20].r.part0[3] ,\sa_snapshot[20].r.part0[2] 
	,\sa_snapshot[20].r.part0[1] ,\sa_snapshot[20].r.part0[0] 
	,\sa_snapshot[19].r.part1[31] ,\sa_snapshot[19].r.part1[30] 
	,\sa_snapshot[19].r.part1[29] ,\sa_snapshot[19].r.part1[28] 
	,\sa_snapshot[19].r.part1[27] ,\sa_snapshot[19].r.part1[26] 
	,\sa_snapshot[19].r.part1[25] ,\sa_snapshot[19].r.part1[24] 
	,\sa_snapshot[19].r.part1[23] ,\sa_snapshot[19].r.part1[22] 
	,\sa_snapshot[19].r.part1[21] ,\sa_snapshot[19].r.part1[20] 
	,\sa_snapshot[19].r.part1[19] ,\sa_snapshot[19].r.part1[18] 
	,\sa_snapshot[19].r.part1[17] ,\sa_snapshot[19].r.part1[16] 
	,\sa_snapshot[19].r.part1[15] ,\sa_snapshot[19].r.part1[14] 
	,\sa_snapshot[19].r.part1[13] ,\sa_snapshot[19].r.part1[12] 
	,\sa_snapshot[19].r.part1[11] ,\sa_snapshot[19].r.part1[10] 
	,\sa_snapshot[19].r.part1[9] ,\sa_snapshot[19].r.part1[8] 
	,\sa_snapshot[19].r.part1[7] ,\sa_snapshot[19].r.part1[6] 
	,\sa_snapshot[19].r.part1[5] ,\sa_snapshot[19].r.part1[4] 
	,\sa_snapshot[19].r.part1[3] ,\sa_snapshot[19].r.part1[2] 
	,\sa_snapshot[19].r.part1[1] ,\sa_snapshot[19].r.part1[0] 
	,\sa_snapshot[19].r.part0[31] ,\sa_snapshot[19].r.part0[30] 
	,\sa_snapshot[19].r.part0[29] ,\sa_snapshot[19].r.part0[28] 
	,\sa_snapshot[19].r.part0[27] ,\sa_snapshot[19].r.part0[26] 
	,\sa_snapshot[19].r.part0[25] ,\sa_snapshot[19].r.part0[24] 
	,\sa_snapshot[19].r.part0[23] ,\sa_snapshot[19].r.part0[22] 
	,\sa_snapshot[19].r.part0[21] ,\sa_snapshot[19].r.part0[20] 
	,\sa_snapshot[19].r.part0[19] ,\sa_snapshot[19].r.part0[18] 
	,\sa_snapshot[19].r.part0[17] ,\sa_snapshot[19].r.part0[16] 
	,\sa_snapshot[19].r.part0[15] ,\sa_snapshot[19].r.part0[14] 
	,\sa_snapshot[19].r.part0[13] ,\sa_snapshot[19].r.part0[12] 
	,\sa_snapshot[19].r.part0[11] ,\sa_snapshot[19].r.part0[10] 
	,\sa_snapshot[19].r.part0[9] ,\sa_snapshot[19].r.part0[8] 
	,\sa_snapshot[19].r.part0[7] ,\sa_snapshot[19].r.part0[6] 
	,\sa_snapshot[19].r.part0[5] ,\sa_snapshot[19].r.part0[4] 
	,\sa_snapshot[19].r.part0[3] ,\sa_snapshot[19].r.part0[2] 
	,\sa_snapshot[19].r.part0[1] ,\sa_snapshot[19].r.part0[0] 
	,\sa_snapshot[18].r.part1[31] ,\sa_snapshot[18].r.part1[30] 
	,\sa_snapshot[18].r.part1[29] ,\sa_snapshot[18].r.part1[28] 
	,\sa_snapshot[18].r.part1[27] ,\sa_snapshot[18].r.part1[26] 
	,\sa_snapshot[18].r.part1[25] ,\sa_snapshot[18].r.part1[24] 
	,\sa_snapshot[18].r.part1[23] ,\sa_snapshot[18].r.part1[22] 
	,\sa_snapshot[18].r.part1[21] ,\sa_snapshot[18].r.part1[20] 
	,\sa_snapshot[18].r.part1[19] ,\sa_snapshot[18].r.part1[18] 
	,\sa_snapshot[18].r.part1[17] ,\sa_snapshot[18].r.part1[16] 
	,\sa_snapshot[18].r.part1[15] ,\sa_snapshot[18].r.part1[14] 
	,\sa_snapshot[18].r.part1[13] ,\sa_snapshot[18].r.part1[12] 
	,\sa_snapshot[18].r.part1[11] ,\sa_snapshot[18].r.part1[10] 
	,\sa_snapshot[18].r.part1[9] ,\sa_snapshot[18].r.part1[8] 
	,\sa_snapshot[18].r.part1[7] ,\sa_snapshot[18].r.part1[6] 
	,\sa_snapshot[18].r.part1[5] ,\sa_snapshot[18].r.part1[4] 
	,\sa_snapshot[18].r.part1[3] ,\sa_snapshot[18].r.part1[2] 
	,\sa_snapshot[18].r.part1[1] ,\sa_snapshot[18].r.part1[0] 
	,\sa_snapshot[18].r.part0[31] ,\sa_snapshot[18].r.part0[30] 
	,\sa_snapshot[18].r.part0[29] ,\sa_snapshot[18].r.part0[28] 
	,\sa_snapshot[18].r.part0[27] ,\sa_snapshot[18].r.part0[26] 
	,\sa_snapshot[18].r.part0[25] ,\sa_snapshot[18].r.part0[24] 
	,\sa_snapshot[18].r.part0[23] ,\sa_snapshot[18].r.part0[22] 
	,\sa_snapshot[18].r.part0[21] ,\sa_snapshot[18].r.part0[20] 
	,\sa_snapshot[18].r.part0[19] ,\sa_snapshot[18].r.part0[18] 
	,\sa_snapshot[18].r.part0[17] ,\sa_snapshot[18].r.part0[16] 
	,\sa_snapshot[18].r.part0[15] ,\sa_snapshot[18].r.part0[14] 
	,\sa_snapshot[18].r.part0[13] ,\sa_snapshot[18].r.part0[12] 
	,\sa_snapshot[18].r.part0[11] ,\sa_snapshot[18].r.part0[10] 
	,\sa_snapshot[18].r.part0[9] ,\sa_snapshot[18].r.part0[8] 
	,\sa_snapshot[18].r.part0[7] ,\sa_snapshot[18].r.part0[6] 
	,\sa_snapshot[18].r.part0[5] ,\sa_snapshot[18].r.part0[4] 
	,\sa_snapshot[18].r.part0[3] ,\sa_snapshot[18].r.part0[2] 
	,\sa_snapshot[18].r.part0[1] ,\sa_snapshot[18].r.part0[0] 
	,\sa_snapshot[17].r.part1[31] ,\sa_snapshot[17].r.part1[30] 
	,\sa_snapshot[17].r.part1[29] ,\sa_snapshot[17].r.part1[28] 
	,\sa_snapshot[17].r.part1[27] ,\sa_snapshot[17].r.part1[26] 
	,\sa_snapshot[17].r.part1[25] ,\sa_snapshot[17].r.part1[24] 
	,\sa_snapshot[17].r.part1[23] ,\sa_snapshot[17].r.part1[22] 
	,\sa_snapshot[17].r.part1[21] ,\sa_snapshot[17].r.part1[20] 
	,\sa_snapshot[17].r.part1[19] ,\sa_snapshot[17].r.part1[18] 
	,\sa_snapshot[17].r.part1[17] ,\sa_snapshot[17].r.part1[16] 
	,\sa_snapshot[17].r.part1[15] ,\sa_snapshot[17].r.part1[14] 
	,\sa_snapshot[17].r.part1[13] ,\sa_snapshot[17].r.part1[12] 
	,\sa_snapshot[17].r.part1[11] ,\sa_snapshot[17].r.part1[10] 
	,\sa_snapshot[17].r.part1[9] ,\sa_snapshot[17].r.part1[8] 
	,\sa_snapshot[17].r.part1[7] ,\sa_snapshot[17].r.part1[6] 
	,\sa_snapshot[17].r.part1[5] ,\sa_snapshot[17].r.part1[4] 
	,\sa_snapshot[17].r.part1[3] ,\sa_snapshot[17].r.part1[2] 
	,\sa_snapshot[17].r.part1[1] ,\sa_snapshot[17].r.part1[0] 
	,\sa_snapshot[17].r.part0[31] ,\sa_snapshot[17].r.part0[30] 
	,\sa_snapshot[17].r.part0[29] ,\sa_snapshot[17].r.part0[28] 
	,\sa_snapshot[17].r.part0[27] ,\sa_snapshot[17].r.part0[26] 
	,\sa_snapshot[17].r.part0[25] ,\sa_snapshot[17].r.part0[24] 
	,\sa_snapshot[17].r.part0[23] ,\sa_snapshot[17].r.part0[22] 
	,\sa_snapshot[17].r.part0[21] ,\sa_snapshot[17].r.part0[20] 
	,\sa_snapshot[17].r.part0[19] ,\sa_snapshot[17].r.part0[18] 
	,\sa_snapshot[17].r.part0[17] ,\sa_snapshot[17].r.part0[16] 
	,\sa_snapshot[17].r.part0[15] ,\sa_snapshot[17].r.part0[14] 
	,\sa_snapshot[17].r.part0[13] ,\sa_snapshot[17].r.part0[12] 
	,\sa_snapshot[17].r.part0[11] ,\sa_snapshot[17].r.part0[10] 
	,\sa_snapshot[17].r.part0[9] ,\sa_snapshot[17].r.part0[8] 
	,\sa_snapshot[17].r.part0[7] ,\sa_snapshot[17].r.part0[6] 
	,\sa_snapshot[17].r.part0[5] ,\sa_snapshot[17].r.part0[4] 
	,\sa_snapshot[17].r.part0[3] ,\sa_snapshot[17].r.part0[2] 
	,\sa_snapshot[17].r.part0[1] ,\sa_snapshot[17].r.part0[0] 
	,\sa_snapshot[16].r.part1[31] ,\sa_snapshot[16].r.part1[30] 
	,\sa_snapshot[16].r.part1[29] ,\sa_snapshot[16].r.part1[28] 
	,\sa_snapshot[16].r.part1[27] ,\sa_snapshot[16].r.part1[26] 
	,\sa_snapshot[16].r.part1[25] ,\sa_snapshot[16].r.part1[24] 
	,\sa_snapshot[16].r.part1[23] ,\sa_snapshot[16].r.part1[22] 
	,\sa_snapshot[16].r.part1[21] ,\sa_snapshot[16].r.part1[20] 
	,\sa_snapshot[16].r.part1[19] ,\sa_snapshot[16].r.part1[18] 
	,\sa_snapshot[16].r.part1[17] ,\sa_snapshot[16].r.part1[16] 
	,\sa_snapshot[16].r.part1[15] ,\sa_snapshot[16].r.part1[14] 
	,\sa_snapshot[16].r.part1[13] ,\sa_snapshot[16].r.part1[12] 
	,\sa_snapshot[16].r.part1[11] ,\sa_snapshot[16].r.part1[10] 
	,\sa_snapshot[16].r.part1[9] ,\sa_snapshot[16].r.part1[8] 
	,\sa_snapshot[16].r.part1[7] ,\sa_snapshot[16].r.part1[6] 
	,\sa_snapshot[16].r.part1[5] ,\sa_snapshot[16].r.part1[4] 
	,\sa_snapshot[16].r.part1[3] ,\sa_snapshot[16].r.part1[2] 
	,\sa_snapshot[16].r.part1[1] ,\sa_snapshot[16].r.part1[0] 
	,\sa_snapshot[16].r.part0[31] ,\sa_snapshot[16].r.part0[30] 
	,\sa_snapshot[16].r.part0[29] ,\sa_snapshot[16].r.part0[28] 
	,\sa_snapshot[16].r.part0[27] ,\sa_snapshot[16].r.part0[26] 
	,\sa_snapshot[16].r.part0[25] ,\sa_snapshot[16].r.part0[24] 
	,\sa_snapshot[16].r.part0[23] ,\sa_snapshot[16].r.part0[22] 
	,\sa_snapshot[16].r.part0[21] ,\sa_snapshot[16].r.part0[20] 
	,\sa_snapshot[16].r.part0[19] ,\sa_snapshot[16].r.part0[18] 
	,\sa_snapshot[16].r.part0[17] ,\sa_snapshot[16].r.part0[16] 
	,\sa_snapshot[16].r.part0[15] ,\sa_snapshot[16].r.part0[14] 
	,\sa_snapshot[16].r.part0[13] ,\sa_snapshot[16].r.part0[12] 
	,\sa_snapshot[16].r.part0[11] ,\sa_snapshot[16].r.part0[10] 
	,\sa_snapshot[16].r.part0[9] ,\sa_snapshot[16].r.part0[8] 
	,\sa_snapshot[16].r.part0[7] ,\sa_snapshot[16].r.part0[6] 
	,\sa_snapshot[16].r.part0[5] ,\sa_snapshot[16].r.part0[4] 
	,\sa_snapshot[16].r.part0[3] ,\sa_snapshot[16].r.part0[2] 
	,\sa_snapshot[16].r.part0[1] ,\sa_snapshot[16].r.part0[0] 
	,\sa_snapshot[15].r.part1[31] ,\sa_snapshot[15].r.part1[30] 
	,\sa_snapshot[15].r.part1[29] ,\sa_snapshot[15].r.part1[28] 
	,\sa_snapshot[15].r.part1[27] ,\sa_snapshot[15].r.part1[26] 
	,\sa_snapshot[15].r.part1[25] ,\sa_snapshot[15].r.part1[24] 
	,\sa_snapshot[15].r.part1[23] ,\sa_snapshot[15].r.part1[22] 
	,\sa_snapshot[15].r.part1[21] ,\sa_snapshot[15].r.part1[20] 
	,\sa_snapshot[15].r.part1[19] ,\sa_snapshot[15].r.part1[18] 
	,\sa_snapshot[15].r.part1[17] ,\sa_snapshot[15].r.part1[16] 
	,\sa_snapshot[15].r.part1[15] ,\sa_snapshot[15].r.part1[14] 
	,\sa_snapshot[15].r.part1[13] ,\sa_snapshot[15].r.part1[12] 
	,\sa_snapshot[15].r.part1[11] ,\sa_snapshot[15].r.part1[10] 
	,\sa_snapshot[15].r.part1[9] ,\sa_snapshot[15].r.part1[8] 
	,\sa_snapshot[15].r.part1[7] ,\sa_snapshot[15].r.part1[6] 
	,\sa_snapshot[15].r.part1[5] ,\sa_snapshot[15].r.part1[4] 
	,\sa_snapshot[15].r.part1[3] ,\sa_snapshot[15].r.part1[2] 
	,\sa_snapshot[15].r.part1[1] ,\sa_snapshot[15].r.part1[0] 
	,\sa_snapshot[15].r.part0[31] ,\sa_snapshot[15].r.part0[30] 
	,\sa_snapshot[15].r.part0[29] ,\sa_snapshot[15].r.part0[28] 
	,\sa_snapshot[15].r.part0[27] ,\sa_snapshot[15].r.part0[26] 
	,\sa_snapshot[15].r.part0[25] ,\sa_snapshot[15].r.part0[24] 
	,\sa_snapshot[15].r.part0[23] ,\sa_snapshot[15].r.part0[22] 
	,\sa_snapshot[15].r.part0[21] ,\sa_snapshot[15].r.part0[20] 
	,\sa_snapshot[15].r.part0[19] ,\sa_snapshot[15].r.part0[18] 
	,\sa_snapshot[15].r.part0[17] ,\sa_snapshot[15].r.part0[16] 
	,\sa_snapshot[15].r.part0[15] ,\sa_snapshot[15].r.part0[14] 
	,\sa_snapshot[15].r.part0[13] ,\sa_snapshot[15].r.part0[12] 
	,\sa_snapshot[15].r.part0[11] ,\sa_snapshot[15].r.part0[10] 
	,\sa_snapshot[15].r.part0[9] ,\sa_snapshot[15].r.part0[8] 
	,\sa_snapshot[15].r.part0[7] ,\sa_snapshot[15].r.part0[6] 
	,\sa_snapshot[15].r.part0[5] ,\sa_snapshot[15].r.part0[4] 
	,\sa_snapshot[15].r.part0[3] ,\sa_snapshot[15].r.part0[2] 
	,\sa_snapshot[15].r.part0[1] ,\sa_snapshot[15].r.part0[0] 
	,\sa_snapshot[14].r.part1[31] ,\sa_snapshot[14].r.part1[30] 
	,\sa_snapshot[14].r.part1[29] ,\sa_snapshot[14].r.part1[28] 
	,\sa_snapshot[14].r.part1[27] ,\sa_snapshot[14].r.part1[26] 
	,\sa_snapshot[14].r.part1[25] ,\sa_snapshot[14].r.part1[24] 
	,\sa_snapshot[14].r.part1[23] ,\sa_snapshot[14].r.part1[22] 
	,\sa_snapshot[14].r.part1[21] ,\sa_snapshot[14].r.part1[20] 
	,\sa_snapshot[14].r.part1[19] ,\sa_snapshot[14].r.part1[18] 
	,\sa_snapshot[14].r.part1[17] ,\sa_snapshot[14].r.part1[16] 
	,\sa_snapshot[14].r.part1[15] ,\sa_snapshot[14].r.part1[14] 
	,\sa_snapshot[14].r.part1[13] ,\sa_snapshot[14].r.part1[12] 
	,\sa_snapshot[14].r.part1[11] ,\sa_snapshot[14].r.part1[10] 
	,\sa_snapshot[14].r.part1[9] ,\sa_snapshot[14].r.part1[8] 
	,\sa_snapshot[14].r.part1[7] ,\sa_snapshot[14].r.part1[6] 
	,\sa_snapshot[14].r.part1[5] ,\sa_snapshot[14].r.part1[4] 
	,\sa_snapshot[14].r.part1[3] ,\sa_snapshot[14].r.part1[2] 
	,\sa_snapshot[14].r.part1[1] ,\sa_snapshot[14].r.part1[0] 
	,\sa_snapshot[14].r.part0[31] ,\sa_snapshot[14].r.part0[30] 
	,\sa_snapshot[14].r.part0[29] ,\sa_snapshot[14].r.part0[28] 
	,\sa_snapshot[14].r.part0[27] ,\sa_snapshot[14].r.part0[26] 
	,\sa_snapshot[14].r.part0[25] ,\sa_snapshot[14].r.part0[24] 
	,\sa_snapshot[14].r.part0[23] ,\sa_snapshot[14].r.part0[22] 
	,\sa_snapshot[14].r.part0[21] ,\sa_snapshot[14].r.part0[20] 
	,\sa_snapshot[14].r.part0[19] ,\sa_snapshot[14].r.part0[18] 
	,\sa_snapshot[14].r.part0[17] ,\sa_snapshot[14].r.part0[16] 
	,\sa_snapshot[14].r.part0[15] ,\sa_snapshot[14].r.part0[14] 
	,\sa_snapshot[14].r.part0[13] ,\sa_snapshot[14].r.part0[12] 
	,\sa_snapshot[14].r.part0[11] ,\sa_snapshot[14].r.part0[10] 
	,\sa_snapshot[14].r.part0[9] ,\sa_snapshot[14].r.part0[8] 
	,\sa_snapshot[14].r.part0[7] ,\sa_snapshot[14].r.part0[6] 
	,\sa_snapshot[14].r.part0[5] ,\sa_snapshot[14].r.part0[4] 
	,\sa_snapshot[14].r.part0[3] ,\sa_snapshot[14].r.part0[2] 
	,\sa_snapshot[14].r.part0[1] ,\sa_snapshot[14].r.part0[0] 
	,\sa_snapshot[13].r.part1[31] ,\sa_snapshot[13].r.part1[30] 
	,\sa_snapshot[13].r.part1[29] ,\sa_snapshot[13].r.part1[28] 
	,\sa_snapshot[13].r.part1[27] ,\sa_snapshot[13].r.part1[26] 
	,\sa_snapshot[13].r.part1[25] ,\sa_snapshot[13].r.part1[24] 
	,\sa_snapshot[13].r.part1[23] ,\sa_snapshot[13].r.part1[22] 
	,\sa_snapshot[13].r.part1[21] ,\sa_snapshot[13].r.part1[20] 
	,\sa_snapshot[13].r.part1[19] ,\sa_snapshot[13].r.part1[18] 
	,\sa_snapshot[13].r.part1[17] ,\sa_snapshot[13].r.part1[16] 
	,\sa_snapshot[13].r.part1[15] ,\sa_snapshot[13].r.part1[14] 
	,\sa_snapshot[13].r.part1[13] ,\sa_snapshot[13].r.part1[12] 
	,\sa_snapshot[13].r.part1[11] ,\sa_snapshot[13].r.part1[10] 
	,\sa_snapshot[13].r.part1[9] ,\sa_snapshot[13].r.part1[8] 
	,\sa_snapshot[13].r.part1[7] ,\sa_snapshot[13].r.part1[6] 
	,\sa_snapshot[13].r.part1[5] ,\sa_snapshot[13].r.part1[4] 
	,\sa_snapshot[13].r.part1[3] ,\sa_snapshot[13].r.part1[2] 
	,\sa_snapshot[13].r.part1[1] ,\sa_snapshot[13].r.part1[0] 
	,\sa_snapshot[13].r.part0[31] ,\sa_snapshot[13].r.part0[30] 
	,\sa_snapshot[13].r.part0[29] ,\sa_snapshot[13].r.part0[28] 
	,\sa_snapshot[13].r.part0[27] ,\sa_snapshot[13].r.part0[26] 
	,\sa_snapshot[13].r.part0[25] ,\sa_snapshot[13].r.part0[24] 
	,\sa_snapshot[13].r.part0[23] ,\sa_snapshot[13].r.part0[22] 
	,\sa_snapshot[13].r.part0[21] ,\sa_snapshot[13].r.part0[20] 
	,\sa_snapshot[13].r.part0[19] ,\sa_snapshot[13].r.part0[18] 
	,\sa_snapshot[13].r.part0[17] ,\sa_snapshot[13].r.part0[16] 
	,\sa_snapshot[13].r.part0[15] ,\sa_snapshot[13].r.part0[14] 
	,\sa_snapshot[13].r.part0[13] ,\sa_snapshot[13].r.part0[12] 
	,\sa_snapshot[13].r.part0[11] ,\sa_snapshot[13].r.part0[10] 
	,\sa_snapshot[13].r.part0[9] ,\sa_snapshot[13].r.part0[8] 
	,\sa_snapshot[13].r.part0[7] ,\sa_snapshot[13].r.part0[6] 
	,\sa_snapshot[13].r.part0[5] ,\sa_snapshot[13].r.part0[4] 
	,\sa_snapshot[13].r.part0[3] ,\sa_snapshot[13].r.part0[2] 
	,\sa_snapshot[13].r.part0[1] ,\sa_snapshot[13].r.part0[0] 
	,\sa_snapshot[12].r.part1[31] ,\sa_snapshot[12].r.part1[30] 
	,\sa_snapshot[12].r.part1[29] ,\sa_snapshot[12].r.part1[28] 
	,\sa_snapshot[12].r.part1[27] ,\sa_snapshot[12].r.part1[26] 
	,\sa_snapshot[12].r.part1[25] ,\sa_snapshot[12].r.part1[24] 
	,\sa_snapshot[12].r.part1[23] ,\sa_snapshot[12].r.part1[22] 
	,\sa_snapshot[12].r.part1[21] ,\sa_snapshot[12].r.part1[20] 
	,\sa_snapshot[12].r.part1[19] ,\sa_snapshot[12].r.part1[18] 
	,\sa_snapshot[12].r.part1[17] ,\sa_snapshot[12].r.part1[16] 
	,\sa_snapshot[12].r.part1[15] ,\sa_snapshot[12].r.part1[14] 
	,\sa_snapshot[12].r.part1[13] ,\sa_snapshot[12].r.part1[12] 
	,\sa_snapshot[12].r.part1[11] ,\sa_snapshot[12].r.part1[10] 
	,\sa_snapshot[12].r.part1[9] ,\sa_snapshot[12].r.part1[8] 
	,\sa_snapshot[12].r.part1[7] ,\sa_snapshot[12].r.part1[6] 
	,\sa_snapshot[12].r.part1[5] ,\sa_snapshot[12].r.part1[4] 
	,\sa_snapshot[12].r.part1[3] ,\sa_snapshot[12].r.part1[2] 
	,\sa_snapshot[12].r.part1[1] ,\sa_snapshot[12].r.part1[0] 
	,\sa_snapshot[12].r.part0[31] ,\sa_snapshot[12].r.part0[30] 
	,\sa_snapshot[12].r.part0[29] ,\sa_snapshot[12].r.part0[28] 
	,\sa_snapshot[12].r.part0[27] ,\sa_snapshot[12].r.part0[26] 
	,\sa_snapshot[12].r.part0[25] ,\sa_snapshot[12].r.part0[24] 
	,\sa_snapshot[12].r.part0[23] ,\sa_snapshot[12].r.part0[22] 
	,\sa_snapshot[12].r.part0[21] ,\sa_snapshot[12].r.part0[20] 
	,\sa_snapshot[12].r.part0[19] ,\sa_snapshot[12].r.part0[18] 
	,\sa_snapshot[12].r.part0[17] ,\sa_snapshot[12].r.part0[16] 
	,\sa_snapshot[12].r.part0[15] ,\sa_snapshot[12].r.part0[14] 
	,\sa_snapshot[12].r.part0[13] ,\sa_snapshot[12].r.part0[12] 
	,\sa_snapshot[12].r.part0[11] ,\sa_snapshot[12].r.part0[10] 
	,\sa_snapshot[12].r.part0[9] ,\sa_snapshot[12].r.part0[8] 
	,\sa_snapshot[12].r.part0[7] ,\sa_snapshot[12].r.part0[6] 
	,\sa_snapshot[12].r.part0[5] ,\sa_snapshot[12].r.part0[4] 
	,\sa_snapshot[12].r.part0[3] ,\sa_snapshot[12].r.part0[2] 
	,\sa_snapshot[12].r.part0[1] ,\sa_snapshot[12].r.part0[0] 
	,\sa_snapshot[11].r.part1[31] ,\sa_snapshot[11].r.part1[30] 
	,\sa_snapshot[11].r.part1[29] ,\sa_snapshot[11].r.part1[28] 
	,\sa_snapshot[11].r.part1[27] ,\sa_snapshot[11].r.part1[26] 
	,\sa_snapshot[11].r.part1[25] ,\sa_snapshot[11].r.part1[24] 
	,\sa_snapshot[11].r.part1[23] ,\sa_snapshot[11].r.part1[22] 
	,\sa_snapshot[11].r.part1[21] ,\sa_snapshot[11].r.part1[20] 
	,\sa_snapshot[11].r.part1[19] ,\sa_snapshot[11].r.part1[18] 
	,\sa_snapshot[11].r.part1[17] ,\sa_snapshot[11].r.part1[16] 
	,\sa_snapshot[11].r.part1[15] ,\sa_snapshot[11].r.part1[14] 
	,\sa_snapshot[11].r.part1[13] ,\sa_snapshot[11].r.part1[12] 
	,\sa_snapshot[11].r.part1[11] ,\sa_snapshot[11].r.part1[10] 
	,\sa_snapshot[11].r.part1[9] ,\sa_snapshot[11].r.part1[8] 
	,\sa_snapshot[11].r.part1[7] ,\sa_snapshot[11].r.part1[6] 
	,\sa_snapshot[11].r.part1[5] ,\sa_snapshot[11].r.part1[4] 
	,\sa_snapshot[11].r.part1[3] ,\sa_snapshot[11].r.part1[2] 
	,\sa_snapshot[11].r.part1[1] ,\sa_snapshot[11].r.part1[0] 
	,\sa_snapshot[11].r.part0[31] ,\sa_snapshot[11].r.part0[30] 
	,\sa_snapshot[11].r.part0[29] ,\sa_snapshot[11].r.part0[28] 
	,\sa_snapshot[11].r.part0[27] ,\sa_snapshot[11].r.part0[26] 
	,\sa_snapshot[11].r.part0[25] ,\sa_snapshot[11].r.part0[24] 
	,\sa_snapshot[11].r.part0[23] ,\sa_snapshot[11].r.part0[22] 
	,\sa_snapshot[11].r.part0[21] ,\sa_snapshot[11].r.part0[20] 
	,\sa_snapshot[11].r.part0[19] ,\sa_snapshot[11].r.part0[18] 
	,\sa_snapshot[11].r.part0[17] ,\sa_snapshot[11].r.part0[16] 
	,\sa_snapshot[11].r.part0[15] ,\sa_snapshot[11].r.part0[14] 
	,\sa_snapshot[11].r.part0[13] ,\sa_snapshot[11].r.part0[12] 
	,\sa_snapshot[11].r.part0[11] ,\sa_snapshot[11].r.part0[10] 
	,\sa_snapshot[11].r.part0[9] ,\sa_snapshot[11].r.part0[8] 
	,\sa_snapshot[11].r.part0[7] ,\sa_snapshot[11].r.part0[6] 
	,\sa_snapshot[11].r.part0[5] ,\sa_snapshot[11].r.part0[4] 
	,\sa_snapshot[11].r.part0[3] ,\sa_snapshot[11].r.part0[2] 
	,\sa_snapshot[11].r.part0[1] ,\sa_snapshot[11].r.part0[0] 
	,\sa_snapshot[10].r.part1[31] ,\sa_snapshot[10].r.part1[30] 
	,\sa_snapshot[10].r.part1[29] ,\sa_snapshot[10].r.part1[28] 
	,\sa_snapshot[10].r.part1[27] ,\sa_snapshot[10].r.part1[26] 
	,\sa_snapshot[10].r.part1[25] ,\sa_snapshot[10].r.part1[24] 
	,\sa_snapshot[10].r.part1[23] ,\sa_snapshot[10].r.part1[22] 
	,\sa_snapshot[10].r.part1[21] ,\sa_snapshot[10].r.part1[20] 
	,\sa_snapshot[10].r.part1[19] ,\sa_snapshot[10].r.part1[18] 
	,\sa_snapshot[10].r.part1[17] ,\sa_snapshot[10].r.part1[16] 
	,\sa_snapshot[10].r.part1[15] ,\sa_snapshot[10].r.part1[14] 
	,\sa_snapshot[10].r.part1[13] ,\sa_snapshot[10].r.part1[12] 
	,\sa_snapshot[10].r.part1[11] ,\sa_snapshot[10].r.part1[10] 
	,\sa_snapshot[10].r.part1[9] ,\sa_snapshot[10].r.part1[8] 
	,\sa_snapshot[10].r.part1[7] ,\sa_snapshot[10].r.part1[6] 
	,\sa_snapshot[10].r.part1[5] ,\sa_snapshot[10].r.part1[4] 
	,\sa_snapshot[10].r.part1[3] ,\sa_snapshot[10].r.part1[2] 
	,\sa_snapshot[10].r.part1[1] ,\sa_snapshot[10].r.part1[0] 
	,\sa_snapshot[10].r.part0[31] ,\sa_snapshot[10].r.part0[30] 
	,\sa_snapshot[10].r.part0[29] ,\sa_snapshot[10].r.part0[28] 
	,\sa_snapshot[10].r.part0[27] ,\sa_snapshot[10].r.part0[26] 
	,\sa_snapshot[10].r.part0[25] ,\sa_snapshot[10].r.part0[24] 
	,\sa_snapshot[10].r.part0[23] ,\sa_snapshot[10].r.part0[22] 
	,\sa_snapshot[10].r.part0[21] ,\sa_snapshot[10].r.part0[20] 
	,\sa_snapshot[10].r.part0[19] ,\sa_snapshot[10].r.part0[18] 
	,\sa_snapshot[10].r.part0[17] ,\sa_snapshot[10].r.part0[16] 
	,\sa_snapshot[10].r.part0[15] ,\sa_snapshot[10].r.part0[14] 
	,\sa_snapshot[10].r.part0[13] ,\sa_snapshot[10].r.part0[12] 
	,\sa_snapshot[10].r.part0[11] ,\sa_snapshot[10].r.part0[10] 
	,\sa_snapshot[10].r.part0[9] ,\sa_snapshot[10].r.part0[8] 
	,\sa_snapshot[10].r.part0[7] ,\sa_snapshot[10].r.part0[6] 
	,\sa_snapshot[10].r.part0[5] ,\sa_snapshot[10].r.part0[4] 
	,\sa_snapshot[10].r.part0[3] ,\sa_snapshot[10].r.part0[2] 
	,\sa_snapshot[10].r.part0[1] ,\sa_snapshot[10].r.part0[0] 
	,\sa_snapshot[9].r.part1[31] ,\sa_snapshot[9].r.part1[30] 
	,\sa_snapshot[9].r.part1[29] ,\sa_snapshot[9].r.part1[28] 
	,\sa_snapshot[9].r.part1[27] ,\sa_snapshot[9].r.part1[26] 
	,\sa_snapshot[9].r.part1[25] ,\sa_snapshot[9].r.part1[24] 
	,\sa_snapshot[9].r.part1[23] ,\sa_snapshot[9].r.part1[22] 
	,\sa_snapshot[9].r.part1[21] ,\sa_snapshot[9].r.part1[20] 
	,\sa_snapshot[9].r.part1[19] ,\sa_snapshot[9].r.part1[18] 
	,\sa_snapshot[9].r.part1[17] ,\sa_snapshot[9].r.part1[16] 
	,\sa_snapshot[9].r.part1[15] ,\sa_snapshot[9].r.part1[14] 
	,\sa_snapshot[9].r.part1[13] ,\sa_snapshot[9].r.part1[12] 
	,\sa_snapshot[9].r.part1[11] ,\sa_snapshot[9].r.part1[10] 
	,\sa_snapshot[9].r.part1[9] ,\sa_snapshot[9].r.part1[8] 
	,\sa_snapshot[9].r.part1[7] ,\sa_snapshot[9].r.part1[6] 
	,\sa_snapshot[9].r.part1[5] ,\sa_snapshot[9].r.part1[4] 
	,\sa_snapshot[9].r.part1[3] ,\sa_snapshot[9].r.part1[2] 
	,\sa_snapshot[9].r.part1[1] ,\sa_snapshot[9].r.part1[0] 
	,\sa_snapshot[9].r.part0[31] ,\sa_snapshot[9].r.part0[30] 
	,\sa_snapshot[9].r.part0[29] ,\sa_snapshot[9].r.part0[28] 
	,\sa_snapshot[9].r.part0[27] ,\sa_snapshot[9].r.part0[26] 
	,\sa_snapshot[9].r.part0[25] ,\sa_snapshot[9].r.part0[24] 
	,\sa_snapshot[9].r.part0[23] ,\sa_snapshot[9].r.part0[22] 
	,\sa_snapshot[9].r.part0[21] ,\sa_snapshot[9].r.part0[20] 
	,\sa_snapshot[9].r.part0[19] ,\sa_snapshot[9].r.part0[18] 
	,\sa_snapshot[9].r.part0[17] ,\sa_snapshot[9].r.part0[16] 
	,\sa_snapshot[9].r.part0[15] ,\sa_snapshot[9].r.part0[14] 
	,\sa_snapshot[9].r.part0[13] ,\sa_snapshot[9].r.part0[12] 
	,\sa_snapshot[9].r.part0[11] ,\sa_snapshot[9].r.part0[10] 
	,\sa_snapshot[9].r.part0[9] ,\sa_snapshot[9].r.part0[8] 
	,\sa_snapshot[9].r.part0[7] ,\sa_snapshot[9].r.part0[6] 
	,\sa_snapshot[9].r.part0[5] ,\sa_snapshot[9].r.part0[4] 
	,\sa_snapshot[9].r.part0[3] ,\sa_snapshot[9].r.part0[2] 
	,\sa_snapshot[9].r.part0[1] ,\sa_snapshot[9].r.part0[0] 
	,\sa_snapshot[8].r.part1[31] ,\sa_snapshot[8].r.part1[30] 
	,\sa_snapshot[8].r.part1[29] ,\sa_snapshot[8].r.part1[28] 
	,\sa_snapshot[8].r.part1[27] ,\sa_snapshot[8].r.part1[26] 
	,\sa_snapshot[8].r.part1[25] ,\sa_snapshot[8].r.part1[24] 
	,\sa_snapshot[8].r.part1[23] ,\sa_snapshot[8].r.part1[22] 
	,\sa_snapshot[8].r.part1[21] ,\sa_snapshot[8].r.part1[20] 
	,\sa_snapshot[8].r.part1[19] ,\sa_snapshot[8].r.part1[18] 
	,\sa_snapshot[8].r.part1[17] ,\sa_snapshot[8].r.part1[16] 
	,\sa_snapshot[8].r.part1[15] ,\sa_snapshot[8].r.part1[14] 
	,\sa_snapshot[8].r.part1[13] ,\sa_snapshot[8].r.part1[12] 
	,\sa_snapshot[8].r.part1[11] ,\sa_snapshot[8].r.part1[10] 
	,\sa_snapshot[8].r.part1[9] ,\sa_snapshot[8].r.part1[8] 
	,\sa_snapshot[8].r.part1[7] ,\sa_snapshot[8].r.part1[6] 
	,\sa_snapshot[8].r.part1[5] ,\sa_snapshot[8].r.part1[4] 
	,\sa_snapshot[8].r.part1[3] ,\sa_snapshot[8].r.part1[2] 
	,\sa_snapshot[8].r.part1[1] ,\sa_snapshot[8].r.part1[0] 
	,\sa_snapshot[8].r.part0[31] ,\sa_snapshot[8].r.part0[30] 
	,\sa_snapshot[8].r.part0[29] ,\sa_snapshot[8].r.part0[28] 
	,\sa_snapshot[8].r.part0[27] ,\sa_snapshot[8].r.part0[26] 
	,\sa_snapshot[8].r.part0[25] ,\sa_snapshot[8].r.part0[24] 
	,\sa_snapshot[8].r.part0[23] ,\sa_snapshot[8].r.part0[22] 
	,\sa_snapshot[8].r.part0[21] ,\sa_snapshot[8].r.part0[20] 
	,\sa_snapshot[8].r.part0[19] ,\sa_snapshot[8].r.part0[18] 
	,\sa_snapshot[8].r.part0[17] ,\sa_snapshot[8].r.part0[16] 
	,\sa_snapshot[8].r.part0[15] ,\sa_snapshot[8].r.part0[14] 
	,\sa_snapshot[8].r.part0[13] ,\sa_snapshot[8].r.part0[12] 
	,\sa_snapshot[8].r.part0[11] ,\sa_snapshot[8].r.part0[10] 
	,\sa_snapshot[8].r.part0[9] ,\sa_snapshot[8].r.part0[8] 
	,\sa_snapshot[8].r.part0[7] ,\sa_snapshot[8].r.part0[6] 
	,\sa_snapshot[8].r.part0[5] ,\sa_snapshot[8].r.part0[4] 
	,\sa_snapshot[8].r.part0[3] ,\sa_snapshot[8].r.part0[2] 
	,\sa_snapshot[8].r.part0[1] ,\sa_snapshot[8].r.part0[0] 
	,\sa_snapshot[7].r.part1[31] ,\sa_snapshot[7].r.part1[30] 
	,\sa_snapshot[7].r.part1[29] ,\sa_snapshot[7].r.part1[28] 
	,\sa_snapshot[7].r.part1[27] ,\sa_snapshot[7].r.part1[26] 
	,\sa_snapshot[7].r.part1[25] ,\sa_snapshot[7].r.part1[24] 
	,\sa_snapshot[7].r.part1[23] ,\sa_snapshot[7].r.part1[22] 
	,\sa_snapshot[7].r.part1[21] ,\sa_snapshot[7].r.part1[20] 
	,\sa_snapshot[7].r.part1[19] ,\sa_snapshot[7].r.part1[18] 
	,\sa_snapshot[7].r.part1[17] ,\sa_snapshot[7].r.part1[16] 
	,\sa_snapshot[7].r.part1[15] ,\sa_snapshot[7].r.part1[14] 
	,\sa_snapshot[7].r.part1[13] ,\sa_snapshot[7].r.part1[12] 
	,\sa_snapshot[7].r.part1[11] ,\sa_snapshot[7].r.part1[10] 
	,\sa_snapshot[7].r.part1[9] ,\sa_snapshot[7].r.part1[8] 
	,\sa_snapshot[7].r.part1[7] ,\sa_snapshot[7].r.part1[6] 
	,\sa_snapshot[7].r.part1[5] ,\sa_snapshot[7].r.part1[4] 
	,\sa_snapshot[7].r.part1[3] ,\sa_snapshot[7].r.part1[2] 
	,\sa_snapshot[7].r.part1[1] ,\sa_snapshot[7].r.part1[0] 
	,\sa_snapshot[7].r.part0[31] ,\sa_snapshot[7].r.part0[30] 
	,\sa_snapshot[7].r.part0[29] ,\sa_snapshot[7].r.part0[28] 
	,\sa_snapshot[7].r.part0[27] ,\sa_snapshot[7].r.part0[26] 
	,\sa_snapshot[7].r.part0[25] ,\sa_snapshot[7].r.part0[24] 
	,\sa_snapshot[7].r.part0[23] ,\sa_snapshot[7].r.part0[22] 
	,\sa_snapshot[7].r.part0[21] ,\sa_snapshot[7].r.part0[20] 
	,\sa_snapshot[7].r.part0[19] ,\sa_snapshot[7].r.part0[18] 
	,\sa_snapshot[7].r.part0[17] ,\sa_snapshot[7].r.part0[16] 
	,\sa_snapshot[7].r.part0[15] ,\sa_snapshot[7].r.part0[14] 
	,\sa_snapshot[7].r.part0[13] ,\sa_snapshot[7].r.part0[12] 
	,\sa_snapshot[7].r.part0[11] ,\sa_snapshot[7].r.part0[10] 
	,\sa_snapshot[7].r.part0[9] ,\sa_snapshot[7].r.part0[8] 
	,\sa_snapshot[7].r.part0[7] ,\sa_snapshot[7].r.part0[6] 
	,\sa_snapshot[7].r.part0[5] ,\sa_snapshot[7].r.part0[4] 
	,\sa_snapshot[7].r.part0[3] ,\sa_snapshot[7].r.part0[2] 
	,\sa_snapshot[7].r.part0[1] ,\sa_snapshot[7].r.part0[0] 
	,\sa_snapshot[6].r.part1[31] ,\sa_snapshot[6].r.part1[30] 
	,\sa_snapshot[6].r.part1[29] ,\sa_snapshot[6].r.part1[28] 
	,\sa_snapshot[6].r.part1[27] ,\sa_snapshot[6].r.part1[26] 
	,\sa_snapshot[6].r.part1[25] ,\sa_snapshot[6].r.part1[24] 
	,\sa_snapshot[6].r.part1[23] ,\sa_snapshot[6].r.part1[22] 
	,\sa_snapshot[6].r.part1[21] ,\sa_snapshot[6].r.part1[20] 
	,\sa_snapshot[6].r.part1[19] ,\sa_snapshot[6].r.part1[18] 
	,\sa_snapshot[6].r.part1[17] ,\sa_snapshot[6].r.part1[16] 
	,\sa_snapshot[6].r.part1[15] ,\sa_snapshot[6].r.part1[14] 
	,\sa_snapshot[6].r.part1[13] ,\sa_snapshot[6].r.part1[12] 
	,\sa_snapshot[6].r.part1[11] ,\sa_snapshot[6].r.part1[10] 
	,\sa_snapshot[6].r.part1[9] ,\sa_snapshot[6].r.part1[8] 
	,\sa_snapshot[6].r.part1[7] ,\sa_snapshot[6].r.part1[6] 
	,\sa_snapshot[6].r.part1[5] ,\sa_snapshot[6].r.part1[4] 
	,\sa_snapshot[6].r.part1[3] ,\sa_snapshot[6].r.part1[2] 
	,\sa_snapshot[6].r.part1[1] ,\sa_snapshot[6].r.part1[0] 
	,\sa_snapshot[6].r.part0[31] ,\sa_snapshot[6].r.part0[30] 
	,\sa_snapshot[6].r.part0[29] ,\sa_snapshot[6].r.part0[28] 
	,\sa_snapshot[6].r.part0[27] ,\sa_snapshot[6].r.part0[26] 
	,\sa_snapshot[6].r.part0[25] ,\sa_snapshot[6].r.part0[24] 
	,\sa_snapshot[6].r.part0[23] ,\sa_snapshot[6].r.part0[22] 
	,\sa_snapshot[6].r.part0[21] ,\sa_snapshot[6].r.part0[20] 
	,\sa_snapshot[6].r.part0[19] ,\sa_snapshot[6].r.part0[18] 
	,\sa_snapshot[6].r.part0[17] ,\sa_snapshot[6].r.part0[16] 
	,\sa_snapshot[6].r.part0[15] ,\sa_snapshot[6].r.part0[14] 
	,\sa_snapshot[6].r.part0[13] ,\sa_snapshot[6].r.part0[12] 
	,\sa_snapshot[6].r.part0[11] ,\sa_snapshot[6].r.part0[10] 
	,\sa_snapshot[6].r.part0[9] ,\sa_snapshot[6].r.part0[8] 
	,\sa_snapshot[6].r.part0[7] ,\sa_snapshot[6].r.part0[6] 
	,\sa_snapshot[6].r.part0[5] ,\sa_snapshot[6].r.part0[4] 
	,\sa_snapshot[6].r.part0[3] ,\sa_snapshot[6].r.part0[2] 
	,\sa_snapshot[6].r.part0[1] ,\sa_snapshot[6].r.part0[0] 
	,\sa_snapshot[5].r.part1[31] ,\sa_snapshot[5].r.part1[30] 
	,\sa_snapshot[5].r.part1[29] ,\sa_snapshot[5].r.part1[28] 
	,\sa_snapshot[5].r.part1[27] ,\sa_snapshot[5].r.part1[26] 
	,\sa_snapshot[5].r.part1[25] ,\sa_snapshot[5].r.part1[24] 
	,\sa_snapshot[5].r.part1[23] ,\sa_snapshot[5].r.part1[22] 
	,\sa_snapshot[5].r.part1[21] ,\sa_snapshot[5].r.part1[20] 
	,\sa_snapshot[5].r.part1[19] ,\sa_snapshot[5].r.part1[18] 
	,\sa_snapshot[5].r.part1[17] ,\sa_snapshot[5].r.part1[16] 
	,\sa_snapshot[5].r.part1[15] ,\sa_snapshot[5].r.part1[14] 
	,\sa_snapshot[5].r.part1[13] ,\sa_snapshot[5].r.part1[12] 
	,\sa_snapshot[5].r.part1[11] ,\sa_snapshot[5].r.part1[10] 
	,\sa_snapshot[5].r.part1[9] ,\sa_snapshot[5].r.part1[8] 
	,\sa_snapshot[5].r.part1[7] ,\sa_snapshot[5].r.part1[6] 
	,\sa_snapshot[5].r.part1[5] ,\sa_snapshot[5].r.part1[4] 
	,\sa_snapshot[5].r.part1[3] ,\sa_snapshot[5].r.part1[2] 
	,\sa_snapshot[5].r.part1[1] ,\sa_snapshot[5].r.part1[0] 
	,\sa_snapshot[5].r.part0[31] ,\sa_snapshot[5].r.part0[30] 
	,\sa_snapshot[5].r.part0[29] ,\sa_snapshot[5].r.part0[28] 
	,\sa_snapshot[5].r.part0[27] ,\sa_snapshot[5].r.part0[26] 
	,\sa_snapshot[5].r.part0[25] ,\sa_snapshot[5].r.part0[24] 
	,\sa_snapshot[5].r.part0[23] ,\sa_snapshot[5].r.part0[22] 
	,\sa_snapshot[5].r.part0[21] ,\sa_snapshot[5].r.part0[20] 
	,\sa_snapshot[5].r.part0[19] ,\sa_snapshot[5].r.part0[18] 
	,\sa_snapshot[5].r.part0[17] ,\sa_snapshot[5].r.part0[16] 
	,\sa_snapshot[5].r.part0[15] ,\sa_snapshot[5].r.part0[14] 
	,\sa_snapshot[5].r.part0[13] ,\sa_snapshot[5].r.part0[12] 
	,\sa_snapshot[5].r.part0[11] ,\sa_snapshot[5].r.part0[10] 
	,\sa_snapshot[5].r.part0[9] ,\sa_snapshot[5].r.part0[8] 
	,\sa_snapshot[5].r.part0[7] ,\sa_snapshot[5].r.part0[6] 
	,\sa_snapshot[5].r.part0[5] ,\sa_snapshot[5].r.part0[4] 
	,\sa_snapshot[5].r.part0[3] ,\sa_snapshot[5].r.part0[2] 
	,\sa_snapshot[5].r.part0[1] ,\sa_snapshot[5].r.part0[0] 
	,\sa_snapshot[4].r.part1[31] ,\sa_snapshot[4].r.part1[30] 
	,\sa_snapshot[4].r.part1[29] ,\sa_snapshot[4].r.part1[28] 
	,\sa_snapshot[4].r.part1[27] ,\sa_snapshot[4].r.part1[26] 
	,\sa_snapshot[4].r.part1[25] ,\sa_snapshot[4].r.part1[24] 
	,\sa_snapshot[4].r.part1[23] ,\sa_snapshot[4].r.part1[22] 
	,\sa_snapshot[4].r.part1[21] ,\sa_snapshot[4].r.part1[20] 
	,\sa_snapshot[4].r.part1[19] ,\sa_snapshot[4].r.part1[18] 
	,\sa_snapshot[4].r.part1[17] ,\sa_snapshot[4].r.part1[16] 
	,\sa_snapshot[4].r.part1[15] ,\sa_snapshot[4].r.part1[14] 
	,\sa_snapshot[4].r.part1[13] ,\sa_snapshot[4].r.part1[12] 
	,\sa_snapshot[4].r.part1[11] ,\sa_snapshot[4].r.part1[10] 
	,\sa_snapshot[4].r.part1[9] ,\sa_snapshot[4].r.part1[8] 
	,\sa_snapshot[4].r.part1[7] ,\sa_snapshot[4].r.part1[6] 
	,\sa_snapshot[4].r.part1[5] ,\sa_snapshot[4].r.part1[4] 
	,\sa_snapshot[4].r.part1[3] ,\sa_snapshot[4].r.part1[2] 
	,\sa_snapshot[4].r.part1[1] ,\sa_snapshot[4].r.part1[0] 
	,\sa_snapshot[4].r.part0[31] ,\sa_snapshot[4].r.part0[30] 
	,\sa_snapshot[4].r.part0[29] ,\sa_snapshot[4].r.part0[28] 
	,\sa_snapshot[4].r.part0[27] ,\sa_snapshot[4].r.part0[26] 
	,\sa_snapshot[4].r.part0[25] ,\sa_snapshot[4].r.part0[24] 
	,\sa_snapshot[4].r.part0[23] ,\sa_snapshot[4].r.part0[22] 
	,\sa_snapshot[4].r.part0[21] ,\sa_snapshot[4].r.part0[20] 
	,\sa_snapshot[4].r.part0[19] ,\sa_snapshot[4].r.part0[18] 
	,\sa_snapshot[4].r.part0[17] ,\sa_snapshot[4].r.part0[16] 
	,\sa_snapshot[4].r.part0[15] ,\sa_snapshot[4].r.part0[14] 
	,\sa_snapshot[4].r.part0[13] ,\sa_snapshot[4].r.part0[12] 
	,\sa_snapshot[4].r.part0[11] ,\sa_snapshot[4].r.part0[10] 
	,\sa_snapshot[4].r.part0[9] ,\sa_snapshot[4].r.part0[8] 
	,\sa_snapshot[4].r.part0[7] ,\sa_snapshot[4].r.part0[6] 
	,\sa_snapshot[4].r.part0[5] ,\sa_snapshot[4].r.part0[4] 
	,\sa_snapshot[4].r.part0[3] ,\sa_snapshot[4].r.part0[2] 
	,\sa_snapshot[4].r.part0[1] ,\sa_snapshot[4].r.part0[0] 
	,\sa_snapshot[3].r.part1[31] ,\sa_snapshot[3].r.part1[30] 
	,\sa_snapshot[3].r.part1[29] ,\sa_snapshot[3].r.part1[28] 
	,\sa_snapshot[3].r.part1[27] ,\sa_snapshot[3].r.part1[26] 
	,\sa_snapshot[3].r.part1[25] ,\sa_snapshot[3].r.part1[24] 
	,\sa_snapshot[3].r.part1[23] ,\sa_snapshot[3].r.part1[22] 
	,\sa_snapshot[3].r.part1[21] ,\sa_snapshot[3].r.part1[20] 
	,\sa_snapshot[3].r.part1[19] ,\sa_snapshot[3].r.part1[18] 
	,\sa_snapshot[3].r.part1[17] ,\sa_snapshot[3].r.part1[16] 
	,\sa_snapshot[3].r.part1[15] ,\sa_snapshot[3].r.part1[14] 
	,\sa_snapshot[3].r.part1[13] ,\sa_snapshot[3].r.part1[12] 
	,\sa_snapshot[3].r.part1[11] ,\sa_snapshot[3].r.part1[10] 
	,\sa_snapshot[3].r.part1[9] ,\sa_snapshot[3].r.part1[8] 
	,\sa_snapshot[3].r.part1[7] ,\sa_snapshot[3].r.part1[6] 
	,\sa_snapshot[3].r.part1[5] ,\sa_snapshot[3].r.part1[4] 
	,\sa_snapshot[3].r.part1[3] ,\sa_snapshot[3].r.part1[2] 
	,\sa_snapshot[3].r.part1[1] ,\sa_snapshot[3].r.part1[0] 
	,\sa_snapshot[3].r.part0[31] ,\sa_snapshot[3].r.part0[30] 
	,\sa_snapshot[3].r.part0[29] ,\sa_snapshot[3].r.part0[28] 
	,\sa_snapshot[3].r.part0[27] ,\sa_snapshot[3].r.part0[26] 
	,\sa_snapshot[3].r.part0[25] ,\sa_snapshot[3].r.part0[24] 
	,\sa_snapshot[3].r.part0[23] ,\sa_snapshot[3].r.part0[22] 
	,\sa_snapshot[3].r.part0[21] ,\sa_snapshot[3].r.part0[20] 
	,\sa_snapshot[3].r.part0[19] ,\sa_snapshot[3].r.part0[18] 
	,\sa_snapshot[3].r.part0[17] ,\sa_snapshot[3].r.part0[16] 
	,\sa_snapshot[3].r.part0[15] ,\sa_snapshot[3].r.part0[14] 
	,\sa_snapshot[3].r.part0[13] ,\sa_snapshot[3].r.part0[12] 
	,\sa_snapshot[3].r.part0[11] ,\sa_snapshot[3].r.part0[10] 
	,\sa_snapshot[3].r.part0[9] ,\sa_snapshot[3].r.part0[8] 
	,\sa_snapshot[3].r.part0[7] ,\sa_snapshot[3].r.part0[6] 
	,\sa_snapshot[3].r.part0[5] ,\sa_snapshot[3].r.part0[4] 
	,\sa_snapshot[3].r.part0[3] ,\sa_snapshot[3].r.part0[2] 
	,\sa_snapshot[3].r.part0[1] ,\sa_snapshot[3].r.part0[0] 
	,\sa_snapshot[2].r.part1[31] ,\sa_snapshot[2].r.part1[30] 
	,\sa_snapshot[2].r.part1[29] ,\sa_snapshot[2].r.part1[28] 
	,\sa_snapshot[2].r.part1[27] ,\sa_snapshot[2].r.part1[26] 
	,\sa_snapshot[2].r.part1[25] ,\sa_snapshot[2].r.part1[24] 
	,\sa_snapshot[2].r.part1[23] ,\sa_snapshot[2].r.part1[22] 
	,\sa_snapshot[2].r.part1[21] ,\sa_snapshot[2].r.part1[20] 
	,\sa_snapshot[2].r.part1[19] ,\sa_snapshot[2].r.part1[18] 
	,\sa_snapshot[2].r.part1[17] ,\sa_snapshot[2].r.part1[16] 
	,\sa_snapshot[2].r.part1[15] ,\sa_snapshot[2].r.part1[14] 
	,\sa_snapshot[2].r.part1[13] ,\sa_snapshot[2].r.part1[12] 
	,\sa_snapshot[2].r.part1[11] ,\sa_snapshot[2].r.part1[10] 
	,\sa_snapshot[2].r.part1[9] ,\sa_snapshot[2].r.part1[8] 
	,\sa_snapshot[2].r.part1[7] ,\sa_snapshot[2].r.part1[6] 
	,\sa_snapshot[2].r.part1[5] ,\sa_snapshot[2].r.part1[4] 
	,\sa_snapshot[2].r.part1[3] ,\sa_snapshot[2].r.part1[2] 
	,\sa_snapshot[2].r.part1[1] ,\sa_snapshot[2].r.part1[0] 
	,\sa_snapshot[2].r.part0[31] ,\sa_snapshot[2].r.part0[30] 
	,\sa_snapshot[2].r.part0[29] ,\sa_snapshot[2].r.part0[28] 
	,\sa_snapshot[2].r.part0[27] ,\sa_snapshot[2].r.part0[26] 
	,\sa_snapshot[2].r.part0[25] ,\sa_snapshot[2].r.part0[24] 
	,\sa_snapshot[2].r.part0[23] ,\sa_snapshot[2].r.part0[22] 
	,\sa_snapshot[2].r.part0[21] ,\sa_snapshot[2].r.part0[20] 
	,\sa_snapshot[2].r.part0[19] ,\sa_snapshot[2].r.part0[18] 
	,\sa_snapshot[2].r.part0[17] ,\sa_snapshot[2].r.part0[16] 
	,\sa_snapshot[2].r.part0[15] ,\sa_snapshot[2].r.part0[14] 
	,\sa_snapshot[2].r.part0[13] ,\sa_snapshot[2].r.part0[12] 
	,\sa_snapshot[2].r.part0[11] ,\sa_snapshot[2].r.part0[10] 
	,\sa_snapshot[2].r.part0[9] ,\sa_snapshot[2].r.part0[8] 
	,\sa_snapshot[2].r.part0[7] ,\sa_snapshot[2].r.part0[6] 
	,\sa_snapshot[2].r.part0[5] ,\sa_snapshot[2].r.part0[4] 
	,\sa_snapshot[2].r.part0[3] ,\sa_snapshot[2].r.part0[2] 
	,\sa_snapshot[2].r.part0[1] ,\sa_snapshot[2].r.part0[0] 
	,\sa_snapshot[1].r.part1[31] ,\sa_snapshot[1].r.part1[30] 
	,\sa_snapshot[1].r.part1[29] ,\sa_snapshot[1].r.part1[28] 
	,\sa_snapshot[1].r.part1[27] ,\sa_snapshot[1].r.part1[26] 
	,\sa_snapshot[1].r.part1[25] ,\sa_snapshot[1].r.part1[24] 
	,\sa_snapshot[1].r.part1[23] ,\sa_snapshot[1].r.part1[22] 
	,\sa_snapshot[1].r.part1[21] ,\sa_snapshot[1].r.part1[20] 
	,\sa_snapshot[1].r.part1[19] ,\sa_snapshot[1].r.part1[18] 
	,\sa_snapshot[1].r.part1[17] ,\sa_snapshot[1].r.part1[16] 
	,\sa_snapshot[1].r.part1[15] ,\sa_snapshot[1].r.part1[14] 
	,\sa_snapshot[1].r.part1[13] ,\sa_snapshot[1].r.part1[12] 
	,\sa_snapshot[1].r.part1[11] ,\sa_snapshot[1].r.part1[10] 
	,\sa_snapshot[1].r.part1[9] ,\sa_snapshot[1].r.part1[8] 
	,\sa_snapshot[1].r.part1[7] ,\sa_snapshot[1].r.part1[6] 
	,\sa_snapshot[1].r.part1[5] ,\sa_snapshot[1].r.part1[4] 
	,\sa_snapshot[1].r.part1[3] ,\sa_snapshot[1].r.part1[2] 
	,\sa_snapshot[1].r.part1[1] ,\sa_snapshot[1].r.part1[0] 
	,\sa_snapshot[1].r.part0[31] ,\sa_snapshot[1].r.part0[30] 
	,\sa_snapshot[1].r.part0[29] ,\sa_snapshot[1].r.part0[28] 
	,\sa_snapshot[1].r.part0[27] ,\sa_snapshot[1].r.part0[26] 
	,\sa_snapshot[1].r.part0[25] ,\sa_snapshot[1].r.part0[24] 
	,\sa_snapshot[1].r.part0[23] ,\sa_snapshot[1].r.part0[22] 
	,\sa_snapshot[1].r.part0[21] ,\sa_snapshot[1].r.part0[20] 
	,\sa_snapshot[1].r.part0[19] ,\sa_snapshot[1].r.part0[18] 
	,\sa_snapshot[1].r.part0[17] ,\sa_snapshot[1].r.part0[16] 
	,\sa_snapshot[1].r.part0[15] ,\sa_snapshot[1].r.part0[14] 
	,\sa_snapshot[1].r.part0[13] ,\sa_snapshot[1].r.part0[12] 
	,\sa_snapshot[1].r.part0[11] ,\sa_snapshot[1].r.part0[10] 
	,\sa_snapshot[1].r.part0[9] ,\sa_snapshot[1].r.part0[8] 
	,\sa_snapshot[1].r.part0[7] ,\sa_snapshot[1].r.part0[6] 
	,\sa_snapshot[1].r.part0[5] ,\sa_snapshot[1].r.part0[4] 
	,\sa_snapshot[1].r.part0[3] ,\sa_snapshot[1].r.part0[2] 
	,\sa_snapshot[1].r.part0[1] ,\sa_snapshot[1].r.part0[0] 
	,\sa_snapshot[0].r.part1[31] ,\sa_snapshot[0].r.part1[30] 
	,\sa_snapshot[0].r.part1[29] ,\sa_snapshot[0].r.part1[28] 
	,\sa_snapshot[0].r.part1[27] ,\sa_snapshot[0].r.part1[26] 
	,\sa_snapshot[0].r.part1[25] ,\sa_snapshot[0].r.part1[24] 
	,\sa_snapshot[0].r.part1[23] ,\sa_snapshot[0].r.part1[22] 
	,\sa_snapshot[0].r.part1[21] ,\sa_snapshot[0].r.part1[20] 
	,\sa_snapshot[0].r.part1[19] ,\sa_snapshot[0].r.part1[18] 
	,\sa_snapshot[0].r.part1[17] ,\sa_snapshot[0].r.part1[16] 
	,\sa_snapshot[0].r.part1[15] ,\sa_snapshot[0].r.part1[14] 
	,\sa_snapshot[0].r.part1[13] ,\sa_snapshot[0].r.part1[12] 
	,\sa_snapshot[0].r.part1[11] ,\sa_snapshot[0].r.part1[10] 
	,\sa_snapshot[0].r.part1[9] ,\sa_snapshot[0].r.part1[8] 
	,\sa_snapshot[0].r.part1[7] ,\sa_snapshot[0].r.part1[6] 
	,\sa_snapshot[0].r.part1[5] ,\sa_snapshot[0].r.part1[4] 
	,\sa_snapshot[0].r.part1[3] ,\sa_snapshot[0].r.part1[2] 
	,\sa_snapshot[0].r.part1[1] ,\sa_snapshot[0].r.part1[0] 
	,\sa_snapshot[0].r.part0[31] ,\sa_snapshot[0].r.part0[30] 
	,\sa_snapshot[0].r.part0[29] ,\sa_snapshot[0].r.part0[28] 
	,\sa_snapshot[0].r.part0[27] ,\sa_snapshot[0].r.part0[26] 
	,\sa_snapshot[0].r.part0[25] ,\sa_snapshot[0].r.part0[24] 
	,\sa_snapshot[0].r.part0[23] ,\sa_snapshot[0].r.part0[22] 
	,\sa_snapshot[0].r.part0[21] ,\sa_snapshot[0].r.part0[20] 
	,\sa_snapshot[0].r.part0[19] ,\sa_snapshot[0].r.part0[18] 
	,\sa_snapshot[0].r.part0[17] ,\sa_snapshot[0].r.part0[16] 
	,\sa_snapshot[0].r.part0[15] ,\sa_snapshot[0].r.part0[14] 
	,\sa_snapshot[0].r.part0[13] ,\sa_snapshot[0].r.part0[12] 
	,\sa_snapshot[0].r.part0[11] ,\sa_snapshot[0].r.part0[10] 
	,\sa_snapshot[0].r.part0[9] ,\sa_snapshot[0].r.part0[8] 
	,\sa_snapshot[0].r.part0[7] ,\sa_snapshot[0].r.part0[6] 
	,\sa_snapshot[0].r.part0[5] ,\sa_snapshot[0].r.part0[4] 
	,\sa_snapshot[0].r.part0[3] ,\sa_snapshot[0].r.part0[2] 
	,\sa_snapshot[0].r.part0[1] ,\sa_snapshot[0].r.part0[0] ;
output \sa_count[31].r.part1[31] ,\sa_count[31].r.part1[30] 
	,\sa_count[31].r.part1[29] ,\sa_count[31].r.part1[28] 
	,\sa_count[31].r.part1[27] ,\sa_count[31].r.part1[26] 
	,\sa_count[31].r.part1[25] ,\sa_count[31].r.part1[24] 
	,\sa_count[31].r.part1[23] ,\sa_count[31].r.part1[22] 
	,\sa_count[31].r.part1[21] ,\sa_count[31].r.part1[20] 
	,\sa_count[31].r.part1[19] ,\sa_count[31].r.part1[18] 
	,\sa_count[31].r.part1[17] ,\sa_count[31].r.part1[16] 
	,\sa_count[31].r.part1[15] ,\sa_count[31].r.part1[14] 
	,\sa_count[31].r.part1[13] ,\sa_count[31].r.part1[12] 
	,\sa_count[31].r.part1[11] ,\sa_count[31].r.part1[10] 
	,\sa_count[31].r.part1[9] ,\sa_count[31].r.part1[8] 
	,\sa_count[31].r.part1[7] ,\sa_count[31].r.part1[6] 
	,\sa_count[31].r.part1[5] ,\sa_count[31].r.part1[4] 
	,\sa_count[31].r.part1[3] ,\sa_count[31].r.part1[2] 
	,\sa_count[31].r.part1[1] ,\sa_count[31].r.part1[0] 
	,\sa_count[31].r.part0[31] ,\sa_count[31].r.part0[30] 
	,\sa_count[31].r.part0[29] ,\sa_count[31].r.part0[28] 
	,\sa_count[31].r.part0[27] ,\sa_count[31].r.part0[26] 
	,\sa_count[31].r.part0[25] ,\sa_count[31].r.part0[24] 
	,\sa_count[31].r.part0[23] ,\sa_count[31].r.part0[22] 
	,\sa_count[31].r.part0[21] ,\sa_count[31].r.part0[20] 
	,\sa_count[31].r.part0[19] ,\sa_count[31].r.part0[18] 
	,\sa_count[31].r.part0[17] ,\sa_count[31].r.part0[16] 
	,\sa_count[31].r.part0[15] ,\sa_count[31].r.part0[14] 
	,\sa_count[31].r.part0[13] ,\sa_count[31].r.part0[12] 
	,\sa_count[31].r.part0[11] ,\sa_count[31].r.part0[10] 
	,\sa_count[31].r.part0[9] ,\sa_count[31].r.part0[8] 
	,\sa_count[31].r.part0[7] ,\sa_count[31].r.part0[6] 
	,\sa_count[31].r.part0[5] ,\sa_count[31].r.part0[4] 
	,\sa_count[31].r.part0[3] ,\sa_count[31].r.part0[2] 
	,\sa_count[31].r.part0[1] ,\sa_count[31].r.part0[0] 
	,\sa_count[30].r.part1[31] ,\sa_count[30].r.part1[30] 
	,\sa_count[30].r.part1[29] ,\sa_count[30].r.part1[28] 
	,\sa_count[30].r.part1[27] ,\sa_count[30].r.part1[26] 
	,\sa_count[30].r.part1[25] ,\sa_count[30].r.part1[24] 
	,\sa_count[30].r.part1[23] ,\sa_count[30].r.part1[22] 
	,\sa_count[30].r.part1[21] ,\sa_count[30].r.part1[20] 
	,\sa_count[30].r.part1[19] ,\sa_count[30].r.part1[18] 
	,\sa_count[30].r.part1[17] ,\sa_count[30].r.part1[16] 
	,\sa_count[30].r.part1[15] ,\sa_count[30].r.part1[14] 
	,\sa_count[30].r.part1[13] ,\sa_count[30].r.part1[12] 
	,\sa_count[30].r.part1[11] ,\sa_count[30].r.part1[10] 
	,\sa_count[30].r.part1[9] ,\sa_count[30].r.part1[8] 
	,\sa_count[30].r.part1[7] ,\sa_count[30].r.part1[6] 
	,\sa_count[30].r.part1[5] ,\sa_count[30].r.part1[4] 
	,\sa_count[30].r.part1[3] ,\sa_count[30].r.part1[2] 
	,\sa_count[30].r.part1[1] ,\sa_count[30].r.part1[0] 
	,\sa_count[30].r.part0[31] ,\sa_count[30].r.part0[30] 
	,\sa_count[30].r.part0[29] ,\sa_count[30].r.part0[28] 
	,\sa_count[30].r.part0[27] ,\sa_count[30].r.part0[26] 
	,\sa_count[30].r.part0[25] ,\sa_count[30].r.part0[24] 
	,\sa_count[30].r.part0[23] ,\sa_count[30].r.part0[22] 
	,\sa_count[30].r.part0[21] ,\sa_count[30].r.part0[20] 
	,\sa_count[30].r.part0[19] ,\sa_count[30].r.part0[18] 
	,\sa_count[30].r.part0[17] ,\sa_count[30].r.part0[16] 
	,\sa_count[30].r.part0[15] ,\sa_count[30].r.part0[14] 
	,\sa_count[30].r.part0[13] ,\sa_count[30].r.part0[12] 
	,\sa_count[30].r.part0[11] ,\sa_count[30].r.part0[10] 
	,\sa_count[30].r.part0[9] ,\sa_count[30].r.part0[8] 
	,\sa_count[30].r.part0[7] ,\sa_count[30].r.part0[6] 
	,\sa_count[30].r.part0[5] ,\sa_count[30].r.part0[4] 
	,\sa_count[30].r.part0[3] ,\sa_count[30].r.part0[2] 
	,\sa_count[30].r.part0[1] ,\sa_count[30].r.part0[0] 
	,\sa_count[29].r.part1[31] ,\sa_count[29].r.part1[30] 
	,\sa_count[29].r.part1[29] ,\sa_count[29].r.part1[28] 
	,\sa_count[29].r.part1[27] ,\sa_count[29].r.part1[26] 
	,\sa_count[29].r.part1[25] ,\sa_count[29].r.part1[24] 
	,\sa_count[29].r.part1[23] ,\sa_count[29].r.part1[22] 
	,\sa_count[29].r.part1[21] ,\sa_count[29].r.part1[20] 
	,\sa_count[29].r.part1[19] ,\sa_count[29].r.part1[18] 
	,\sa_count[29].r.part1[17] ,\sa_count[29].r.part1[16] 
	,\sa_count[29].r.part1[15] ,\sa_count[29].r.part1[14] 
	,\sa_count[29].r.part1[13] ,\sa_count[29].r.part1[12] 
	,\sa_count[29].r.part1[11] ,\sa_count[29].r.part1[10] 
	,\sa_count[29].r.part1[9] ,\sa_count[29].r.part1[8] 
	,\sa_count[29].r.part1[7] ,\sa_count[29].r.part1[6] 
	,\sa_count[29].r.part1[5] ,\sa_count[29].r.part1[4] 
	,\sa_count[29].r.part1[3] ,\sa_count[29].r.part1[2] 
	,\sa_count[29].r.part1[1] ,\sa_count[29].r.part1[0] 
	,\sa_count[29].r.part0[31] ,\sa_count[29].r.part0[30] 
	,\sa_count[29].r.part0[29] ,\sa_count[29].r.part0[28] 
	,\sa_count[29].r.part0[27] ,\sa_count[29].r.part0[26] 
	,\sa_count[29].r.part0[25] ,\sa_count[29].r.part0[24] 
	,\sa_count[29].r.part0[23] ,\sa_count[29].r.part0[22] 
	,\sa_count[29].r.part0[21] ,\sa_count[29].r.part0[20] 
	,\sa_count[29].r.part0[19] ,\sa_count[29].r.part0[18] 
	,\sa_count[29].r.part0[17] ,\sa_count[29].r.part0[16] 
	,\sa_count[29].r.part0[15] ,\sa_count[29].r.part0[14] 
	,\sa_count[29].r.part0[13] ,\sa_count[29].r.part0[12] 
	,\sa_count[29].r.part0[11] ,\sa_count[29].r.part0[10] 
	,\sa_count[29].r.part0[9] ,\sa_count[29].r.part0[8] 
	,\sa_count[29].r.part0[7] ,\sa_count[29].r.part0[6] 
	,\sa_count[29].r.part0[5] ,\sa_count[29].r.part0[4] 
	,\sa_count[29].r.part0[3] ,\sa_count[29].r.part0[2] 
	,\sa_count[29].r.part0[1] ,\sa_count[29].r.part0[0] 
	,\sa_count[28].r.part1[31] ,\sa_count[28].r.part1[30] 
	,\sa_count[28].r.part1[29] ,\sa_count[28].r.part1[28] 
	,\sa_count[28].r.part1[27] ,\sa_count[28].r.part1[26] 
	,\sa_count[28].r.part1[25] ,\sa_count[28].r.part1[24] 
	,\sa_count[28].r.part1[23] ,\sa_count[28].r.part1[22] 
	,\sa_count[28].r.part1[21] ,\sa_count[28].r.part1[20] 
	,\sa_count[28].r.part1[19] ,\sa_count[28].r.part1[18] 
	,\sa_count[28].r.part1[17] ,\sa_count[28].r.part1[16] 
	,\sa_count[28].r.part1[15] ,\sa_count[28].r.part1[14] 
	,\sa_count[28].r.part1[13] ,\sa_count[28].r.part1[12] 
	,\sa_count[28].r.part1[11] ,\sa_count[28].r.part1[10] 
	,\sa_count[28].r.part1[9] ,\sa_count[28].r.part1[8] 
	,\sa_count[28].r.part1[7] ,\sa_count[28].r.part1[6] 
	,\sa_count[28].r.part1[5] ,\sa_count[28].r.part1[4] 
	,\sa_count[28].r.part1[3] ,\sa_count[28].r.part1[2] 
	,\sa_count[28].r.part1[1] ,\sa_count[28].r.part1[0] 
	,\sa_count[28].r.part0[31] ,\sa_count[28].r.part0[30] 
	,\sa_count[28].r.part0[29] ,\sa_count[28].r.part0[28] 
	,\sa_count[28].r.part0[27] ,\sa_count[28].r.part0[26] 
	,\sa_count[28].r.part0[25] ,\sa_count[28].r.part0[24] 
	,\sa_count[28].r.part0[23] ,\sa_count[28].r.part0[22] 
	,\sa_count[28].r.part0[21] ,\sa_count[28].r.part0[20] 
	,\sa_count[28].r.part0[19] ,\sa_count[28].r.part0[18] 
	,\sa_count[28].r.part0[17] ,\sa_count[28].r.part0[16] 
	,\sa_count[28].r.part0[15] ,\sa_count[28].r.part0[14] 
	,\sa_count[28].r.part0[13] ,\sa_count[28].r.part0[12] 
	,\sa_count[28].r.part0[11] ,\sa_count[28].r.part0[10] 
	,\sa_count[28].r.part0[9] ,\sa_count[28].r.part0[8] 
	,\sa_count[28].r.part0[7] ,\sa_count[28].r.part0[6] 
	,\sa_count[28].r.part0[5] ,\sa_count[28].r.part0[4] 
	,\sa_count[28].r.part0[3] ,\sa_count[28].r.part0[2] 
	,\sa_count[28].r.part0[1] ,\sa_count[28].r.part0[0] 
	,\sa_count[27].r.part1[31] ,\sa_count[27].r.part1[30] 
	,\sa_count[27].r.part1[29] ,\sa_count[27].r.part1[28] 
	,\sa_count[27].r.part1[27] ,\sa_count[27].r.part1[26] 
	,\sa_count[27].r.part1[25] ,\sa_count[27].r.part1[24] 
	,\sa_count[27].r.part1[23] ,\sa_count[27].r.part1[22] 
	,\sa_count[27].r.part1[21] ,\sa_count[27].r.part1[20] 
	,\sa_count[27].r.part1[19] ,\sa_count[27].r.part1[18] 
	,\sa_count[27].r.part1[17] ,\sa_count[27].r.part1[16] 
	,\sa_count[27].r.part1[15] ,\sa_count[27].r.part1[14] 
	,\sa_count[27].r.part1[13] ,\sa_count[27].r.part1[12] 
	,\sa_count[27].r.part1[11] ,\sa_count[27].r.part1[10] 
	,\sa_count[27].r.part1[9] ,\sa_count[27].r.part1[8] 
	,\sa_count[27].r.part1[7] ,\sa_count[27].r.part1[6] 
	,\sa_count[27].r.part1[5] ,\sa_count[27].r.part1[4] 
	,\sa_count[27].r.part1[3] ,\sa_count[27].r.part1[2] 
	,\sa_count[27].r.part1[1] ,\sa_count[27].r.part1[0] 
	,\sa_count[27].r.part0[31] ,\sa_count[27].r.part0[30] 
	,\sa_count[27].r.part0[29] ,\sa_count[27].r.part0[28] 
	,\sa_count[27].r.part0[27] ,\sa_count[27].r.part0[26] 
	,\sa_count[27].r.part0[25] ,\sa_count[27].r.part0[24] 
	,\sa_count[27].r.part0[23] ,\sa_count[27].r.part0[22] 
	,\sa_count[27].r.part0[21] ,\sa_count[27].r.part0[20] 
	,\sa_count[27].r.part0[19] ,\sa_count[27].r.part0[18] 
	,\sa_count[27].r.part0[17] ,\sa_count[27].r.part0[16] 
	,\sa_count[27].r.part0[15] ,\sa_count[27].r.part0[14] 
	,\sa_count[27].r.part0[13] ,\sa_count[27].r.part0[12] 
	,\sa_count[27].r.part0[11] ,\sa_count[27].r.part0[10] 
	,\sa_count[27].r.part0[9] ,\sa_count[27].r.part0[8] 
	,\sa_count[27].r.part0[7] ,\sa_count[27].r.part0[6] 
	,\sa_count[27].r.part0[5] ,\sa_count[27].r.part0[4] 
	,\sa_count[27].r.part0[3] ,\sa_count[27].r.part0[2] 
	,\sa_count[27].r.part0[1] ,\sa_count[27].r.part0[0] 
	,\sa_count[26].r.part1[31] ,\sa_count[26].r.part1[30] 
	,\sa_count[26].r.part1[29] ,\sa_count[26].r.part1[28] 
	,\sa_count[26].r.part1[27] ,\sa_count[26].r.part1[26] 
	,\sa_count[26].r.part1[25] ,\sa_count[26].r.part1[24] 
	,\sa_count[26].r.part1[23] ,\sa_count[26].r.part1[22] 
	,\sa_count[26].r.part1[21] ,\sa_count[26].r.part1[20] 
	,\sa_count[26].r.part1[19] ,\sa_count[26].r.part1[18] 
	,\sa_count[26].r.part1[17] ,\sa_count[26].r.part1[16] 
	,\sa_count[26].r.part1[15] ,\sa_count[26].r.part1[14] 
	,\sa_count[26].r.part1[13] ,\sa_count[26].r.part1[12] 
	,\sa_count[26].r.part1[11] ,\sa_count[26].r.part1[10] 
	,\sa_count[26].r.part1[9] ,\sa_count[26].r.part1[8] 
	,\sa_count[26].r.part1[7] ,\sa_count[26].r.part1[6] 
	,\sa_count[26].r.part1[5] ,\sa_count[26].r.part1[4] 
	,\sa_count[26].r.part1[3] ,\sa_count[26].r.part1[2] 
	,\sa_count[26].r.part1[1] ,\sa_count[26].r.part1[0] 
	,\sa_count[26].r.part0[31] ,\sa_count[26].r.part0[30] 
	,\sa_count[26].r.part0[29] ,\sa_count[26].r.part0[28] 
	,\sa_count[26].r.part0[27] ,\sa_count[26].r.part0[26] 
	,\sa_count[26].r.part0[25] ,\sa_count[26].r.part0[24] 
	,\sa_count[26].r.part0[23] ,\sa_count[26].r.part0[22] 
	,\sa_count[26].r.part0[21] ,\sa_count[26].r.part0[20] 
	,\sa_count[26].r.part0[19] ,\sa_count[26].r.part0[18] 
	,\sa_count[26].r.part0[17] ,\sa_count[26].r.part0[16] 
	,\sa_count[26].r.part0[15] ,\sa_count[26].r.part0[14] 
	,\sa_count[26].r.part0[13] ,\sa_count[26].r.part0[12] 
	,\sa_count[26].r.part0[11] ,\sa_count[26].r.part0[10] 
	,\sa_count[26].r.part0[9] ,\sa_count[26].r.part0[8] 
	,\sa_count[26].r.part0[7] ,\sa_count[26].r.part0[6] 
	,\sa_count[26].r.part0[5] ,\sa_count[26].r.part0[4] 
	,\sa_count[26].r.part0[3] ,\sa_count[26].r.part0[2] 
	,\sa_count[26].r.part0[1] ,\sa_count[26].r.part0[0] 
	,\sa_count[25].r.part1[31] ,\sa_count[25].r.part1[30] 
	,\sa_count[25].r.part1[29] ,\sa_count[25].r.part1[28] 
	,\sa_count[25].r.part1[27] ,\sa_count[25].r.part1[26] 
	,\sa_count[25].r.part1[25] ,\sa_count[25].r.part1[24] 
	,\sa_count[25].r.part1[23] ,\sa_count[25].r.part1[22] 
	,\sa_count[25].r.part1[21] ,\sa_count[25].r.part1[20] 
	,\sa_count[25].r.part1[19] ,\sa_count[25].r.part1[18] 
	,\sa_count[25].r.part1[17] ,\sa_count[25].r.part1[16] 
	,\sa_count[25].r.part1[15] ,\sa_count[25].r.part1[14] 
	,\sa_count[25].r.part1[13] ,\sa_count[25].r.part1[12] 
	,\sa_count[25].r.part1[11] ,\sa_count[25].r.part1[10] 
	,\sa_count[25].r.part1[9] ,\sa_count[25].r.part1[8] 
	,\sa_count[25].r.part1[7] ,\sa_count[25].r.part1[6] 
	,\sa_count[25].r.part1[5] ,\sa_count[25].r.part1[4] 
	,\sa_count[25].r.part1[3] ,\sa_count[25].r.part1[2] 
	,\sa_count[25].r.part1[1] ,\sa_count[25].r.part1[0] 
	,\sa_count[25].r.part0[31] ,\sa_count[25].r.part0[30] 
	,\sa_count[25].r.part0[29] ,\sa_count[25].r.part0[28] 
	,\sa_count[25].r.part0[27] ,\sa_count[25].r.part0[26] 
	,\sa_count[25].r.part0[25] ,\sa_count[25].r.part0[24] 
	,\sa_count[25].r.part0[23] ,\sa_count[25].r.part0[22] 
	,\sa_count[25].r.part0[21] ,\sa_count[25].r.part0[20] 
	,\sa_count[25].r.part0[19] ,\sa_count[25].r.part0[18] 
	,\sa_count[25].r.part0[17] ,\sa_count[25].r.part0[16] 
	,\sa_count[25].r.part0[15] ,\sa_count[25].r.part0[14] 
	,\sa_count[25].r.part0[13] ,\sa_count[25].r.part0[12] 
	,\sa_count[25].r.part0[11] ,\sa_count[25].r.part0[10] 
	,\sa_count[25].r.part0[9] ,\sa_count[25].r.part0[8] 
	,\sa_count[25].r.part0[7] ,\sa_count[25].r.part0[6] 
	,\sa_count[25].r.part0[5] ,\sa_count[25].r.part0[4] 
	,\sa_count[25].r.part0[3] ,\sa_count[25].r.part0[2] 
	,\sa_count[25].r.part0[1] ,\sa_count[25].r.part0[0] 
	,\sa_count[24].r.part1[31] ,\sa_count[24].r.part1[30] 
	,\sa_count[24].r.part1[29] ,\sa_count[24].r.part1[28] 
	,\sa_count[24].r.part1[27] ,\sa_count[24].r.part1[26] 
	,\sa_count[24].r.part1[25] ,\sa_count[24].r.part1[24] 
	,\sa_count[24].r.part1[23] ,\sa_count[24].r.part1[22] 
	,\sa_count[24].r.part1[21] ,\sa_count[24].r.part1[20] 
	,\sa_count[24].r.part1[19] ,\sa_count[24].r.part1[18] 
	,\sa_count[24].r.part1[17] ,\sa_count[24].r.part1[16] 
	,\sa_count[24].r.part1[15] ,\sa_count[24].r.part1[14] 
	,\sa_count[24].r.part1[13] ,\sa_count[24].r.part1[12] 
	,\sa_count[24].r.part1[11] ,\sa_count[24].r.part1[10] 
	,\sa_count[24].r.part1[9] ,\sa_count[24].r.part1[8] 
	,\sa_count[24].r.part1[7] ,\sa_count[24].r.part1[6] 
	,\sa_count[24].r.part1[5] ,\sa_count[24].r.part1[4] 
	,\sa_count[24].r.part1[3] ,\sa_count[24].r.part1[2] 
	,\sa_count[24].r.part1[1] ,\sa_count[24].r.part1[0] 
	,\sa_count[24].r.part0[31] ,\sa_count[24].r.part0[30] 
	,\sa_count[24].r.part0[29] ,\sa_count[24].r.part0[28] 
	,\sa_count[24].r.part0[27] ,\sa_count[24].r.part0[26] 
	,\sa_count[24].r.part0[25] ,\sa_count[24].r.part0[24] 
	,\sa_count[24].r.part0[23] ,\sa_count[24].r.part0[22] 
	,\sa_count[24].r.part0[21] ,\sa_count[24].r.part0[20] 
	,\sa_count[24].r.part0[19] ,\sa_count[24].r.part0[18] 
	,\sa_count[24].r.part0[17] ,\sa_count[24].r.part0[16] 
	,\sa_count[24].r.part0[15] ,\sa_count[24].r.part0[14] 
	,\sa_count[24].r.part0[13] ,\sa_count[24].r.part0[12] 
	,\sa_count[24].r.part0[11] ,\sa_count[24].r.part0[10] 
	,\sa_count[24].r.part0[9] ,\sa_count[24].r.part0[8] 
	,\sa_count[24].r.part0[7] ,\sa_count[24].r.part0[6] 
	,\sa_count[24].r.part0[5] ,\sa_count[24].r.part0[4] 
	,\sa_count[24].r.part0[3] ,\sa_count[24].r.part0[2] 
	,\sa_count[24].r.part0[1] ,\sa_count[24].r.part0[0] 
	,\sa_count[23].r.part1[31] ,\sa_count[23].r.part1[30] 
	,\sa_count[23].r.part1[29] ,\sa_count[23].r.part1[28] 
	,\sa_count[23].r.part1[27] ,\sa_count[23].r.part1[26] 
	,\sa_count[23].r.part1[25] ,\sa_count[23].r.part1[24] 
	,\sa_count[23].r.part1[23] ,\sa_count[23].r.part1[22] 
	,\sa_count[23].r.part1[21] ,\sa_count[23].r.part1[20] 
	,\sa_count[23].r.part1[19] ,\sa_count[23].r.part1[18] 
	,\sa_count[23].r.part1[17] ,\sa_count[23].r.part1[16] 
	,\sa_count[23].r.part1[15] ,\sa_count[23].r.part1[14] 
	,\sa_count[23].r.part1[13] ,\sa_count[23].r.part1[12] 
	,\sa_count[23].r.part1[11] ,\sa_count[23].r.part1[10] 
	,\sa_count[23].r.part1[9] ,\sa_count[23].r.part1[8] 
	,\sa_count[23].r.part1[7] ,\sa_count[23].r.part1[6] 
	,\sa_count[23].r.part1[5] ,\sa_count[23].r.part1[4] 
	,\sa_count[23].r.part1[3] ,\sa_count[23].r.part1[2] 
	,\sa_count[23].r.part1[1] ,\sa_count[23].r.part1[0] 
	,\sa_count[23].r.part0[31] ,\sa_count[23].r.part0[30] 
	,\sa_count[23].r.part0[29] ,\sa_count[23].r.part0[28] 
	,\sa_count[23].r.part0[27] ,\sa_count[23].r.part0[26] 
	,\sa_count[23].r.part0[25] ,\sa_count[23].r.part0[24] 
	,\sa_count[23].r.part0[23] ,\sa_count[23].r.part0[22] 
	,\sa_count[23].r.part0[21] ,\sa_count[23].r.part0[20] 
	,\sa_count[23].r.part0[19] ,\sa_count[23].r.part0[18] 
	,\sa_count[23].r.part0[17] ,\sa_count[23].r.part0[16] 
	,\sa_count[23].r.part0[15] ,\sa_count[23].r.part0[14] 
	,\sa_count[23].r.part0[13] ,\sa_count[23].r.part0[12] 
	,\sa_count[23].r.part0[11] ,\sa_count[23].r.part0[10] 
	,\sa_count[23].r.part0[9] ,\sa_count[23].r.part0[8] 
	,\sa_count[23].r.part0[7] ,\sa_count[23].r.part0[6] 
	,\sa_count[23].r.part0[5] ,\sa_count[23].r.part0[4] 
	,\sa_count[23].r.part0[3] ,\sa_count[23].r.part0[2] 
	,\sa_count[23].r.part0[1] ,\sa_count[23].r.part0[0] 
	,\sa_count[22].r.part1[31] ,\sa_count[22].r.part1[30] 
	,\sa_count[22].r.part1[29] ,\sa_count[22].r.part1[28] 
	,\sa_count[22].r.part1[27] ,\sa_count[22].r.part1[26] 
	,\sa_count[22].r.part1[25] ,\sa_count[22].r.part1[24] 
	,\sa_count[22].r.part1[23] ,\sa_count[22].r.part1[22] 
	,\sa_count[22].r.part1[21] ,\sa_count[22].r.part1[20] 
	,\sa_count[22].r.part1[19] ,\sa_count[22].r.part1[18] 
	,\sa_count[22].r.part1[17] ,\sa_count[22].r.part1[16] 
	,\sa_count[22].r.part1[15] ,\sa_count[22].r.part1[14] 
	,\sa_count[22].r.part1[13] ,\sa_count[22].r.part1[12] 
	,\sa_count[22].r.part1[11] ,\sa_count[22].r.part1[10] 
	,\sa_count[22].r.part1[9] ,\sa_count[22].r.part1[8] 
	,\sa_count[22].r.part1[7] ,\sa_count[22].r.part1[6] 
	,\sa_count[22].r.part1[5] ,\sa_count[22].r.part1[4] 
	,\sa_count[22].r.part1[3] ,\sa_count[22].r.part1[2] 
	,\sa_count[22].r.part1[1] ,\sa_count[22].r.part1[0] 
	,\sa_count[22].r.part0[31] ,\sa_count[22].r.part0[30] 
	,\sa_count[22].r.part0[29] ,\sa_count[22].r.part0[28] 
	,\sa_count[22].r.part0[27] ,\sa_count[22].r.part0[26] 
	,\sa_count[22].r.part0[25] ,\sa_count[22].r.part0[24] 
	,\sa_count[22].r.part0[23] ,\sa_count[22].r.part0[22] 
	,\sa_count[22].r.part0[21] ,\sa_count[22].r.part0[20] 
	,\sa_count[22].r.part0[19] ,\sa_count[22].r.part0[18] 
	,\sa_count[22].r.part0[17] ,\sa_count[22].r.part0[16] 
	,\sa_count[22].r.part0[15] ,\sa_count[22].r.part0[14] 
	,\sa_count[22].r.part0[13] ,\sa_count[22].r.part0[12] 
	,\sa_count[22].r.part0[11] ,\sa_count[22].r.part0[10] 
	,\sa_count[22].r.part0[9] ,\sa_count[22].r.part0[8] 
	,\sa_count[22].r.part0[7] ,\sa_count[22].r.part0[6] 
	,\sa_count[22].r.part0[5] ,\sa_count[22].r.part0[4] 
	,\sa_count[22].r.part0[3] ,\sa_count[22].r.part0[2] 
	,\sa_count[22].r.part0[1] ,\sa_count[22].r.part0[0] 
	,\sa_count[21].r.part1[31] ,\sa_count[21].r.part1[30] 
	,\sa_count[21].r.part1[29] ,\sa_count[21].r.part1[28] 
	,\sa_count[21].r.part1[27] ,\sa_count[21].r.part1[26] 
	,\sa_count[21].r.part1[25] ,\sa_count[21].r.part1[24] 
	,\sa_count[21].r.part1[23] ,\sa_count[21].r.part1[22] 
	,\sa_count[21].r.part1[21] ,\sa_count[21].r.part1[20] 
	,\sa_count[21].r.part1[19] ,\sa_count[21].r.part1[18] 
	,\sa_count[21].r.part1[17] ,\sa_count[21].r.part1[16] 
	,\sa_count[21].r.part1[15] ,\sa_count[21].r.part1[14] 
	,\sa_count[21].r.part1[13] ,\sa_count[21].r.part1[12] 
	,\sa_count[21].r.part1[11] ,\sa_count[21].r.part1[10] 
	,\sa_count[21].r.part1[9] ,\sa_count[21].r.part1[8] 
	,\sa_count[21].r.part1[7] ,\sa_count[21].r.part1[6] 
	,\sa_count[21].r.part1[5] ,\sa_count[21].r.part1[4] 
	,\sa_count[21].r.part1[3] ,\sa_count[21].r.part1[2] 
	,\sa_count[21].r.part1[1] ,\sa_count[21].r.part1[0] 
	,\sa_count[21].r.part0[31] ,\sa_count[21].r.part0[30] 
	,\sa_count[21].r.part0[29] ,\sa_count[21].r.part0[28] 
	,\sa_count[21].r.part0[27] ,\sa_count[21].r.part0[26] 
	,\sa_count[21].r.part0[25] ,\sa_count[21].r.part0[24] 
	,\sa_count[21].r.part0[23] ,\sa_count[21].r.part0[22] 
	,\sa_count[21].r.part0[21] ,\sa_count[21].r.part0[20] 
	,\sa_count[21].r.part0[19] ,\sa_count[21].r.part0[18] 
	,\sa_count[21].r.part0[17] ,\sa_count[21].r.part0[16] 
	,\sa_count[21].r.part0[15] ,\sa_count[21].r.part0[14] 
	,\sa_count[21].r.part0[13] ,\sa_count[21].r.part0[12] 
	,\sa_count[21].r.part0[11] ,\sa_count[21].r.part0[10] 
	,\sa_count[21].r.part0[9] ,\sa_count[21].r.part0[8] 
	,\sa_count[21].r.part0[7] ,\sa_count[21].r.part0[6] 
	,\sa_count[21].r.part0[5] ,\sa_count[21].r.part0[4] 
	,\sa_count[21].r.part0[3] ,\sa_count[21].r.part0[2] 
	,\sa_count[21].r.part0[1] ,\sa_count[21].r.part0[0] 
	,\sa_count[20].r.part1[31] ,\sa_count[20].r.part1[30] 
	,\sa_count[20].r.part1[29] ,\sa_count[20].r.part1[28] 
	,\sa_count[20].r.part1[27] ,\sa_count[20].r.part1[26] 
	,\sa_count[20].r.part1[25] ,\sa_count[20].r.part1[24] 
	,\sa_count[20].r.part1[23] ,\sa_count[20].r.part1[22] 
	,\sa_count[20].r.part1[21] ,\sa_count[20].r.part1[20] 
	,\sa_count[20].r.part1[19] ,\sa_count[20].r.part1[18] 
	,\sa_count[20].r.part1[17] ,\sa_count[20].r.part1[16] 
	,\sa_count[20].r.part1[15] ,\sa_count[20].r.part1[14] 
	,\sa_count[20].r.part1[13] ,\sa_count[20].r.part1[12] 
	,\sa_count[20].r.part1[11] ,\sa_count[20].r.part1[10] 
	,\sa_count[20].r.part1[9] ,\sa_count[20].r.part1[8] 
	,\sa_count[20].r.part1[7] ,\sa_count[20].r.part1[6] 
	,\sa_count[20].r.part1[5] ,\sa_count[20].r.part1[4] 
	,\sa_count[20].r.part1[3] ,\sa_count[20].r.part1[2] 
	,\sa_count[20].r.part1[1] ,\sa_count[20].r.part1[0] 
	,\sa_count[20].r.part0[31] ,\sa_count[20].r.part0[30] 
	,\sa_count[20].r.part0[29] ,\sa_count[20].r.part0[28] 
	,\sa_count[20].r.part0[27] ,\sa_count[20].r.part0[26] 
	,\sa_count[20].r.part0[25] ,\sa_count[20].r.part0[24] 
	,\sa_count[20].r.part0[23] ,\sa_count[20].r.part0[22] 
	,\sa_count[20].r.part0[21] ,\sa_count[20].r.part0[20] 
	,\sa_count[20].r.part0[19] ,\sa_count[20].r.part0[18] 
	,\sa_count[20].r.part0[17] ,\sa_count[20].r.part0[16] 
	,\sa_count[20].r.part0[15] ,\sa_count[20].r.part0[14] 
	,\sa_count[20].r.part0[13] ,\sa_count[20].r.part0[12] 
	,\sa_count[20].r.part0[11] ,\sa_count[20].r.part0[10] 
	,\sa_count[20].r.part0[9] ,\sa_count[20].r.part0[8] 
	,\sa_count[20].r.part0[7] ,\sa_count[20].r.part0[6] 
	,\sa_count[20].r.part0[5] ,\sa_count[20].r.part0[4] 
	,\sa_count[20].r.part0[3] ,\sa_count[20].r.part0[2] 
	,\sa_count[20].r.part0[1] ,\sa_count[20].r.part0[0] 
	,\sa_count[19].r.part1[31] ,\sa_count[19].r.part1[30] 
	,\sa_count[19].r.part1[29] ,\sa_count[19].r.part1[28] 
	,\sa_count[19].r.part1[27] ,\sa_count[19].r.part1[26] 
	,\sa_count[19].r.part1[25] ,\sa_count[19].r.part1[24] 
	,\sa_count[19].r.part1[23] ,\sa_count[19].r.part1[22] 
	,\sa_count[19].r.part1[21] ,\sa_count[19].r.part1[20] 
	,\sa_count[19].r.part1[19] ,\sa_count[19].r.part1[18] 
	,\sa_count[19].r.part1[17] ,\sa_count[19].r.part1[16] 
	,\sa_count[19].r.part1[15] ,\sa_count[19].r.part1[14] 
	,\sa_count[19].r.part1[13] ,\sa_count[19].r.part1[12] 
	,\sa_count[19].r.part1[11] ,\sa_count[19].r.part1[10] 
	,\sa_count[19].r.part1[9] ,\sa_count[19].r.part1[8] 
	,\sa_count[19].r.part1[7] ,\sa_count[19].r.part1[6] 
	,\sa_count[19].r.part1[5] ,\sa_count[19].r.part1[4] 
	,\sa_count[19].r.part1[3] ,\sa_count[19].r.part1[2] 
	,\sa_count[19].r.part1[1] ,\sa_count[19].r.part1[0] 
	,\sa_count[19].r.part0[31] ,\sa_count[19].r.part0[30] 
	,\sa_count[19].r.part0[29] ,\sa_count[19].r.part0[28] 
	,\sa_count[19].r.part0[27] ,\sa_count[19].r.part0[26] 
	,\sa_count[19].r.part0[25] ,\sa_count[19].r.part0[24] 
	,\sa_count[19].r.part0[23] ,\sa_count[19].r.part0[22] 
	,\sa_count[19].r.part0[21] ,\sa_count[19].r.part0[20] 
	,\sa_count[19].r.part0[19] ,\sa_count[19].r.part0[18] 
	,\sa_count[19].r.part0[17] ,\sa_count[19].r.part0[16] 
	,\sa_count[19].r.part0[15] ,\sa_count[19].r.part0[14] 
	,\sa_count[19].r.part0[13] ,\sa_count[19].r.part0[12] 
	,\sa_count[19].r.part0[11] ,\sa_count[19].r.part0[10] 
	,\sa_count[19].r.part0[9] ,\sa_count[19].r.part0[8] 
	,\sa_count[19].r.part0[7] ,\sa_count[19].r.part0[6] 
	,\sa_count[19].r.part0[5] ,\sa_count[19].r.part0[4] 
	,\sa_count[19].r.part0[3] ,\sa_count[19].r.part0[2] 
	,\sa_count[19].r.part0[1] ,\sa_count[19].r.part0[0] 
	,\sa_count[18].r.part1[31] ,\sa_count[18].r.part1[30] 
	,\sa_count[18].r.part1[29] ,\sa_count[18].r.part1[28] 
	,\sa_count[18].r.part1[27] ,\sa_count[18].r.part1[26] 
	,\sa_count[18].r.part1[25] ,\sa_count[18].r.part1[24] 
	,\sa_count[18].r.part1[23] ,\sa_count[18].r.part1[22] 
	,\sa_count[18].r.part1[21] ,\sa_count[18].r.part1[20] 
	,\sa_count[18].r.part1[19] ,\sa_count[18].r.part1[18] 
	,\sa_count[18].r.part1[17] ,\sa_count[18].r.part1[16] 
	,\sa_count[18].r.part1[15] ,\sa_count[18].r.part1[14] 
	,\sa_count[18].r.part1[13] ,\sa_count[18].r.part1[12] 
	,\sa_count[18].r.part1[11] ,\sa_count[18].r.part1[10] 
	,\sa_count[18].r.part1[9] ,\sa_count[18].r.part1[8] 
	,\sa_count[18].r.part1[7] ,\sa_count[18].r.part1[6] 
	,\sa_count[18].r.part1[5] ,\sa_count[18].r.part1[4] 
	,\sa_count[18].r.part1[3] ,\sa_count[18].r.part1[2] 
	,\sa_count[18].r.part1[1] ,\sa_count[18].r.part1[0] 
	,\sa_count[18].r.part0[31] ,\sa_count[18].r.part0[30] 
	,\sa_count[18].r.part0[29] ,\sa_count[18].r.part0[28] 
	,\sa_count[18].r.part0[27] ,\sa_count[18].r.part0[26] 
	,\sa_count[18].r.part0[25] ,\sa_count[18].r.part0[24] 
	,\sa_count[18].r.part0[23] ,\sa_count[18].r.part0[22] 
	,\sa_count[18].r.part0[21] ,\sa_count[18].r.part0[20] 
	,\sa_count[18].r.part0[19] ,\sa_count[18].r.part0[18] 
	,\sa_count[18].r.part0[17] ,\sa_count[18].r.part0[16] 
	,\sa_count[18].r.part0[15] ,\sa_count[18].r.part0[14] 
	,\sa_count[18].r.part0[13] ,\sa_count[18].r.part0[12] 
	,\sa_count[18].r.part0[11] ,\sa_count[18].r.part0[10] 
	,\sa_count[18].r.part0[9] ,\sa_count[18].r.part0[8] 
	,\sa_count[18].r.part0[7] ,\sa_count[18].r.part0[6] 
	,\sa_count[18].r.part0[5] ,\sa_count[18].r.part0[4] 
	,\sa_count[18].r.part0[3] ,\sa_count[18].r.part0[2] 
	,\sa_count[18].r.part0[1] ,\sa_count[18].r.part0[0] 
	,\sa_count[17].r.part1[31] ,\sa_count[17].r.part1[30] 
	,\sa_count[17].r.part1[29] ,\sa_count[17].r.part1[28] 
	,\sa_count[17].r.part1[27] ,\sa_count[17].r.part1[26] 
	,\sa_count[17].r.part1[25] ,\sa_count[17].r.part1[24] 
	,\sa_count[17].r.part1[23] ,\sa_count[17].r.part1[22] 
	,\sa_count[17].r.part1[21] ,\sa_count[17].r.part1[20] 
	,\sa_count[17].r.part1[19] ,\sa_count[17].r.part1[18] 
	,\sa_count[17].r.part1[17] ,\sa_count[17].r.part1[16] 
	,\sa_count[17].r.part1[15] ,\sa_count[17].r.part1[14] 
	,\sa_count[17].r.part1[13] ,\sa_count[17].r.part1[12] 
	,\sa_count[17].r.part1[11] ,\sa_count[17].r.part1[10] 
	,\sa_count[17].r.part1[9] ,\sa_count[17].r.part1[8] 
	,\sa_count[17].r.part1[7] ,\sa_count[17].r.part1[6] 
	,\sa_count[17].r.part1[5] ,\sa_count[17].r.part1[4] 
	,\sa_count[17].r.part1[3] ,\sa_count[17].r.part1[2] 
	,\sa_count[17].r.part1[1] ,\sa_count[17].r.part1[0] 
	,\sa_count[17].r.part0[31] ,\sa_count[17].r.part0[30] 
	,\sa_count[17].r.part0[29] ,\sa_count[17].r.part0[28] 
	,\sa_count[17].r.part0[27] ,\sa_count[17].r.part0[26] 
	,\sa_count[17].r.part0[25] ,\sa_count[17].r.part0[24] 
	,\sa_count[17].r.part0[23] ,\sa_count[17].r.part0[22] 
	,\sa_count[17].r.part0[21] ,\sa_count[17].r.part0[20] 
	,\sa_count[17].r.part0[19] ,\sa_count[17].r.part0[18] 
	,\sa_count[17].r.part0[17] ,\sa_count[17].r.part0[16] 
	,\sa_count[17].r.part0[15] ,\sa_count[17].r.part0[14] 
	,\sa_count[17].r.part0[13] ,\sa_count[17].r.part0[12] 
	,\sa_count[17].r.part0[11] ,\sa_count[17].r.part0[10] 
	,\sa_count[17].r.part0[9] ,\sa_count[17].r.part0[8] 
	,\sa_count[17].r.part0[7] ,\sa_count[17].r.part0[6] 
	,\sa_count[17].r.part0[5] ,\sa_count[17].r.part0[4] 
	,\sa_count[17].r.part0[3] ,\sa_count[17].r.part0[2] 
	,\sa_count[17].r.part0[1] ,\sa_count[17].r.part0[0] 
	,\sa_count[16].r.part1[31] ,\sa_count[16].r.part1[30] 
	,\sa_count[16].r.part1[29] ,\sa_count[16].r.part1[28] 
	,\sa_count[16].r.part1[27] ,\sa_count[16].r.part1[26] 
	,\sa_count[16].r.part1[25] ,\sa_count[16].r.part1[24] 
	,\sa_count[16].r.part1[23] ,\sa_count[16].r.part1[22] 
	,\sa_count[16].r.part1[21] ,\sa_count[16].r.part1[20] 
	,\sa_count[16].r.part1[19] ,\sa_count[16].r.part1[18] 
	,\sa_count[16].r.part1[17] ,\sa_count[16].r.part1[16] 
	,\sa_count[16].r.part1[15] ,\sa_count[16].r.part1[14] 
	,\sa_count[16].r.part1[13] ,\sa_count[16].r.part1[12] 
	,\sa_count[16].r.part1[11] ,\sa_count[16].r.part1[10] 
	,\sa_count[16].r.part1[9] ,\sa_count[16].r.part1[8] 
	,\sa_count[16].r.part1[7] ,\sa_count[16].r.part1[6] 
	,\sa_count[16].r.part1[5] ,\sa_count[16].r.part1[4] 
	,\sa_count[16].r.part1[3] ,\sa_count[16].r.part1[2] 
	,\sa_count[16].r.part1[1] ,\sa_count[16].r.part1[0] 
	,\sa_count[16].r.part0[31] ,\sa_count[16].r.part0[30] 
	,\sa_count[16].r.part0[29] ,\sa_count[16].r.part0[28] 
	,\sa_count[16].r.part0[27] ,\sa_count[16].r.part0[26] 
	,\sa_count[16].r.part0[25] ,\sa_count[16].r.part0[24] 
	,\sa_count[16].r.part0[23] ,\sa_count[16].r.part0[22] 
	,\sa_count[16].r.part0[21] ,\sa_count[16].r.part0[20] 
	,\sa_count[16].r.part0[19] ,\sa_count[16].r.part0[18] 
	,\sa_count[16].r.part0[17] ,\sa_count[16].r.part0[16] 
	,\sa_count[16].r.part0[15] ,\sa_count[16].r.part0[14] 
	,\sa_count[16].r.part0[13] ,\sa_count[16].r.part0[12] 
	,\sa_count[16].r.part0[11] ,\sa_count[16].r.part0[10] 
	,\sa_count[16].r.part0[9] ,\sa_count[16].r.part0[8] 
	,\sa_count[16].r.part0[7] ,\sa_count[16].r.part0[6] 
	,\sa_count[16].r.part0[5] ,\sa_count[16].r.part0[4] 
	,\sa_count[16].r.part0[3] ,\sa_count[16].r.part0[2] 
	,\sa_count[16].r.part0[1] ,\sa_count[16].r.part0[0] 
	,\sa_count[15].r.part1[31] ,\sa_count[15].r.part1[30] 
	,\sa_count[15].r.part1[29] ,\sa_count[15].r.part1[28] 
	,\sa_count[15].r.part1[27] ,\sa_count[15].r.part1[26] 
	,\sa_count[15].r.part1[25] ,\sa_count[15].r.part1[24] 
	,\sa_count[15].r.part1[23] ,\sa_count[15].r.part1[22] 
	,\sa_count[15].r.part1[21] ,\sa_count[15].r.part1[20] 
	,\sa_count[15].r.part1[19] ,\sa_count[15].r.part1[18] 
	,\sa_count[15].r.part1[17] ,\sa_count[15].r.part1[16] 
	,\sa_count[15].r.part1[15] ,\sa_count[15].r.part1[14] 
	,\sa_count[15].r.part1[13] ,\sa_count[15].r.part1[12] 
	,\sa_count[15].r.part1[11] ,\sa_count[15].r.part1[10] 
	,\sa_count[15].r.part1[9] ,\sa_count[15].r.part1[8] 
	,\sa_count[15].r.part1[7] ,\sa_count[15].r.part1[6] 
	,\sa_count[15].r.part1[5] ,\sa_count[15].r.part1[4] 
	,\sa_count[15].r.part1[3] ,\sa_count[15].r.part1[2] 
	,\sa_count[15].r.part1[1] ,\sa_count[15].r.part1[0] 
	,\sa_count[15].r.part0[31] ,\sa_count[15].r.part0[30] 
	,\sa_count[15].r.part0[29] ,\sa_count[15].r.part0[28] 
	,\sa_count[15].r.part0[27] ,\sa_count[15].r.part0[26] 
	,\sa_count[15].r.part0[25] ,\sa_count[15].r.part0[24] 
	,\sa_count[15].r.part0[23] ,\sa_count[15].r.part0[22] 
	,\sa_count[15].r.part0[21] ,\sa_count[15].r.part0[20] 
	,\sa_count[15].r.part0[19] ,\sa_count[15].r.part0[18] 
	,\sa_count[15].r.part0[17] ,\sa_count[15].r.part0[16] 
	,\sa_count[15].r.part0[15] ,\sa_count[15].r.part0[14] 
	,\sa_count[15].r.part0[13] ,\sa_count[15].r.part0[12] 
	,\sa_count[15].r.part0[11] ,\sa_count[15].r.part0[10] 
	,\sa_count[15].r.part0[9] ,\sa_count[15].r.part0[8] 
	,\sa_count[15].r.part0[7] ,\sa_count[15].r.part0[6] 
	,\sa_count[15].r.part0[5] ,\sa_count[15].r.part0[4] 
	,\sa_count[15].r.part0[3] ,\sa_count[15].r.part0[2] 
	,\sa_count[15].r.part0[1] ,\sa_count[15].r.part0[0] 
	,\sa_count[14].r.part1[31] ,\sa_count[14].r.part1[30] 
	,\sa_count[14].r.part1[29] ,\sa_count[14].r.part1[28] 
	,\sa_count[14].r.part1[27] ,\sa_count[14].r.part1[26] 
	,\sa_count[14].r.part1[25] ,\sa_count[14].r.part1[24] 
	,\sa_count[14].r.part1[23] ,\sa_count[14].r.part1[22] 
	,\sa_count[14].r.part1[21] ,\sa_count[14].r.part1[20] 
	,\sa_count[14].r.part1[19] ,\sa_count[14].r.part1[18] 
	,\sa_count[14].r.part1[17] ,\sa_count[14].r.part1[16] 
	,\sa_count[14].r.part1[15] ,\sa_count[14].r.part1[14] 
	,\sa_count[14].r.part1[13] ,\sa_count[14].r.part1[12] 
	,\sa_count[14].r.part1[11] ,\sa_count[14].r.part1[10] 
	,\sa_count[14].r.part1[9] ,\sa_count[14].r.part1[8] 
	,\sa_count[14].r.part1[7] ,\sa_count[14].r.part1[6] 
	,\sa_count[14].r.part1[5] ,\sa_count[14].r.part1[4] 
	,\sa_count[14].r.part1[3] ,\sa_count[14].r.part1[2] 
	,\sa_count[14].r.part1[1] ,\sa_count[14].r.part1[0] 
	,\sa_count[14].r.part0[31] ,\sa_count[14].r.part0[30] 
	,\sa_count[14].r.part0[29] ,\sa_count[14].r.part0[28] 
	,\sa_count[14].r.part0[27] ,\sa_count[14].r.part0[26] 
	,\sa_count[14].r.part0[25] ,\sa_count[14].r.part0[24] 
	,\sa_count[14].r.part0[23] ,\sa_count[14].r.part0[22] 
	,\sa_count[14].r.part0[21] ,\sa_count[14].r.part0[20] 
	,\sa_count[14].r.part0[19] ,\sa_count[14].r.part0[18] 
	,\sa_count[14].r.part0[17] ,\sa_count[14].r.part0[16] 
	,\sa_count[14].r.part0[15] ,\sa_count[14].r.part0[14] 
	,\sa_count[14].r.part0[13] ,\sa_count[14].r.part0[12] 
	,\sa_count[14].r.part0[11] ,\sa_count[14].r.part0[10] 
	,\sa_count[14].r.part0[9] ,\sa_count[14].r.part0[8] 
	,\sa_count[14].r.part0[7] ,\sa_count[14].r.part0[6] 
	,\sa_count[14].r.part0[5] ,\sa_count[14].r.part0[4] 
	,\sa_count[14].r.part0[3] ,\sa_count[14].r.part0[2] 
	,\sa_count[14].r.part0[1] ,\sa_count[14].r.part0[0] 
	,\sa_count[13].r.part1[31] ,\sa_count[13].r.part1[30] 
	,\sa_count[13].r.part1[29] ,\sa_count[13].r.part1[28] 
	,\sa_count[13].r.part1[27] ,\sa_count[13].r.part1[26] 
	,\sa_count[13].r.part1[25] ,\sa_count[13].r.part1[24] 
	,\sa_count[13].r.part1[23] ,\sa_count[13].r.part1[22] 
	,\sa_count[13].r.part1[21] ,\sa_count[13].r.part1[20] 
	,\sa_count[13].r.part1[19] ,\sa_count[13].r.part1[18] 
	,\sa_count[13].r.part1[17] ,\sa_count[13].r.part1[16] 
	,\sa_count[13].r.part1[15] ,\sa_count[13].r.part1[14] 
	,\sa_count[13].r.part1[13] ,\sa_count[13].r.part1[12] 
	,\sa_count[13].r.part1[11] ,\sa_count[13].r.part1[10] 
	,\sa_count[13].r.part1[9] ,\sa_count[13].r.part1[8] 
	,\sa_count[13].r.part1[7] ,\sa_count[13].r.part1[6] 
	,\sa_count[13].r.part1[5] ,\sa_count[13].r.part1[4] 
	,\sa_count[13].r.part1[3] ,\sa_count[13].r.part1[2] 
	,\sa_count[13].r.part1[1] ,\sa_count[13].r.part1[0] 
	,\sa_count[13].r.part0[31] ,\sa_count[13].r.part0[30] 
	,\sa_count[13].r.part0[29] ,\sa_count[13].r.part0[28] 
	,\sa_count[13].r.part0[27] ,\sa_count[13].r.part0[26] 
	,\sa_count[13].r.part0[25] ,\sa_count[13].r.part0[24] 
	,\sa_count[13].r.part0[23] ,\sa_count[13].r.part0[22] 
	,\sa_count[13].r.part0[21] ,\sa_count[13].r.part0[20] 
	,\sa_count[13].r.part0[19] ,\sa_count[13].r.part0[18] 
	,\sa_count[13].r.part0[17] ,\sa_count[13].r.part0[16] 
	,\sa_count[13].r.part0[15] ,\sa_count[13].r.part0[14] 
	,\sa_count[13].r.part0[13] ,\sa_count[13].r.part0[12] 
	,\sa_count[13].r.part0[11] ,\sa_count[13].r.part0[10] 
	,\sa_count[13].r.part0[9] ,\sa_count[13].r.part0[8] 
	,\sa_count[13].r.part0[7] ,\sa_count[13].r.part0[6] 
	,\sa_count[13].r.part0[5] ,\sa_count[13].r.part0[4] 
	,\sa_count[13].r.part0[3] ,\sa_count[13].r.part0[2] 
	,\sa_count[13].r.part0[1] ,\sa_count[13].r.part0[0] 
	,\sa_count[12].r.part1[31] ,\sa_count[12].r.part1[30] 
	,\sa_count[12].r.part1[29] ,\sa_count[12].r.part1[28] 
	,\sa_count[12].r.part1[27] ,\sa_count[12].r.part1[26] 
	,\sa_count[12].r.part1[25] ,\sa_count[12].r.part1[24] 
	,\sa_count[12].r.part1[23] ,\sa_count[12].r.part1[22] 
	,\sa_count[12].r.part1[21] ,\sa_count[12].r.part1[20] 
	,\sa_count[12].r.part1[19] ,\sa_count[12].r.part1[18] 
	,\sa_count[12].r.part1[17] ,\sa_count[12].r.part1[16] 
	,\sa_count[12].r.part1[15] ,\sa_count[12].r.part1[14] 
	,\sa_count[12].r.part1[13] ,\sa_count[12].r.part1[12] 
	,\sa_count[12].r.part1[11] ,\sa_count[12].r.part1[10] 
	,\sa_count[12].r.part1[9] ,\sa_count[12].r.part1[8] 
	,\sa_count[12].r.part1[7] ,\sa_count[12].r.part1[6] 
	,\sa_count[12].r.part1[5] ,\sa_count[12].r.part1[4] 
	,\sa_count[12].r.part1[3] ,\sa_count[12].r.part1[2] 
	,\sa_count[12].r.part1[1] ,\sa_count[12].r.part1[0] 
	,\sa_count[12].r.part0[31] ,\sa_count[12].r.part0[30] 
	,\sa_count[12].r.part0[29] ,\sa_count[12].r.part0[28] 
	,\sa_count[12].r.part0[27] ,\sa_count[12].r.part0[26] 
	,\sa_count[12].r.part0[25] ,\sa_count[12].r.part0[24] 
	,\sa_count[12].r.part0[23] ,\sa_count[12].r.part0[22] 
	,\sa_count[12].r.part0[21] ,\sa_count[12].r.part0[20] 
	,\sa_count[12].r.part0[19] ,\sa_count[12].r.part0[18] 
	,\sa_count[12].r.part0[17] ,\sa_count[12].r.part0[16] 
	,\sa_count[12].r.part0[15] ,\sa_count[12].r.part0[14] 
	,\sa_count[12].r.part0[13] ,\sa_count[12].r.part0[12] 
	,\sa_count[12].r.part0[11] ,\sa_count[12].r.part0[10] 
	,\sa_count[12].r.part0[9] ,\sa_count[12].r.part0[8] 
	,\sa_count[12].r.part0[7] ,\sa_count[12].r.part0[6] 
	,\sa_count[12].r.part0[5] ,\sa_count[12].r.part0[4] 
	,\sa_count[12].r.part0[3] ,\sa_count[12].r.part0[2] 
	,\sa_count[12].r.part0[1] ,\sa_count[12].r.part0[0] 
	,\sa_count[11].r.part1[31] ,\sa_count[11].r.part1[30] 
	,\sa_count[11].r.part1[29] ,\sa_count[11].r.part1[28] 
	,\sa_count[11].r.part1[27] ,\sa_count[11].r.part1[26] 
	,\sa_count[11].r.part1[25] ,\sa_count[11].r.part1[24] 
	,\sa_count[11].r.part1[23] ,\sa_count[11].r.part1[22] 
	,\sa_count[11].r.part1[21] ,\sa_count[11].r.part1[20] 
	,\sa_count[11].r.part1[19] ,\sa_count[11].r.part1[18] 
	,\sa_count[11].r.part1[17] ,\sa_count[11].r.part1[16] 
	,\sa_count[11].r.part1[15] ,\sa_count[11].r.part1[14] 
	,\sa_count[11].r.part1[13] ,\sa_count[11].r.part1[12] 
	,\sa_count[11].r.part1[11] ,\sa_count[11].r.part1[10] 
	,\sa_count[11].r.part1[9] ,\sa_count[11].r.part1[8] 
	,\sa_count[11].r.part1[7] ,\sa_count[11].r.part1[6] 
	,\sa_count[11].r.part1[5] ,\sa_count[11].r.part1[4] 
	,\sa_count[11].r.part1[3] ,\sa_count[11].r.part1[2] 
	,\sa_count[11].r.part1[1] ,\sa_count[11].r.part1[0] 
	,\sa_count[11].r.part0[31] ,\sa_count[11].r.part0[30] 
	,\sa_count[11].r.part0[29] ,\sa_count[11].r.part0[28] 
	,\sa_count[11].r.part0[27] ,\sa_count[11].r.part0[26] 
	,\sa_count[11].r.part0[25] ,\sa_count[11].r.part0[24] 
	,\sa_count[11].r.part0[23] ,\sa_count[11].r.part0[22] 
	,\sa_count[11].r.part0[21] ,\sa_count[11].r.part0[20] 
	,\sa_count[11].r.part0[19] ,\sa_count[11].r.part0[18] 
	,\sa_count[11].r.part0[17] ,\sa_count[11].r.part0[16] 
	,\sa_count[11].r.part0[15] ,\sa_count[11].r.part0[14] 
	,\sa_count[11].r.part0[13] ,\sa_count[11].r.part0[12] 
	,\sa_count[11].r.part0[11] ,\sa_count[11].r.part0[10] 
	,\sa_count[11].r.part0[9] ,\sa_count[11].r.part0[8] 
	,\sa_count[11].r.part0[7] ,\sa_count[11].r.part0[6] 
	,\sa_count[11].r.part0[5] ,\sa_count[11].r.part0[4] 
	,\sa_count[11].r.part0[3] ,\sa_count[11].r.part0[2] 
	,\sa_count[11].r.part0[1] ,\sa_count[11].r.part0[0] 
	,\sa_count[10].r.part1[31] ,\sa_count[10].r.part1[30] 
	,\sa_count[10].r.part1[29] ,\sa_count[10].r.part1[28] 
	,\sa_count[10].r.part1[27] ,\sa_count[10].r.part1[26] 
	,\sa_count[10].r.part1[25] ,\sa_count[10].r.part1[24] 
	,\sa_count[10].r.part1[23] ,\sa_count[10].r.part1[22] 
	,\sa_count[10].r.part1[21] ,\sa_count[10].r.part1[20] 
	,\sa_count[10].r.part1[19] ,\sa_count[10].r.part1[18] 
	,\sa_count[10].r.part1[17] ,\sa_count[10].r.part1[16] 
	,\sa_count[10].r.part1[15] ,\sa_count[10].r.part1[14] 
	,\sa_count[10].r.part1[13] ,\sa_count[10].r.part1[12] 
	,\sa_count[10].r.part1[11] ,\sa_count[10].r.part1[10] 
	,\sa_count[10].r.part1[9] ,\sa_count[10].r.part1[8] 
	,\sa_count[10].r.part1[7] ,\sa_count[10].r.part1[6] 
	,\sa_count[10].r.part1[5] ,\sa_count[10].r.part1[4] 
	,\sa_count[10].r.part1[3] ,\sa_count[10].r.part1[2] 
	,\sa_count[10].r.part1[1] ,\sa_count[10].r.part1[0] 
	,\sa_count[10].r.part0[31] ,\sa_count[10].r.part0[30] 
	,\sa_count[10].r.part0[29] ,\sa_count[10].r.part0[28] 
	,\sa_count[10].r.part0[27] ,\sa_count[10].r.part0[26] 
	,\sa_count[10].r.part0[25] ,\sa_count[10].r.part0[24] 
	,\sa_count[10].r.part0[23] ,\sa_count[10].r.part0[22] 
	,\sa_count[10].r.part0[21] ,\sa_count[10].r.part0[20] 
	,\sa_count[10].r.part0[19] ,\sa_count[10].r.part0[18] 
	,\sa_count[10].r.part0[17] ,\sa_count[10].r.part0[16] 
	,\sa_count[10].r.part0[15] ,\sa_count[10].r.part0[14] 
	,\sa_count[10].r.part0[13] ,\sa_count[10].r.part0[12] 
	,\sa_count[10].r.part0[11] ,\sa_count[10].r.part0[10] 
	,\sa_count[10].r.part0[9] ,\sa_count[10].r.part0[8] 
	,\sa_count[10].r.part0[7] ,\sa_count[10].r.part0[6] 
	,\sa_count[10].r.part0[5] ,\sa_count[10].r.part0[4] 
	,\sa_count[10].r.part0[3] ,\sa_count[10].r.part0[2] 
	,\sa_count[10].r.part0[1] ,\sa_count[10].r.part0[0] 
	,\sa_count[9].r.part1[31] ,\sa_count[9].r.part1[30] 
	,\sa_count[9].r.part1[29] ,\sa_count[9].r.part1[28] 
	,\sa_count[9].r.part1[27] ,\sa_count[9].r.part1[26] 
	,\sa_count[9].r.part1[25] ,\sa_count[9].r.part1[24] 
	,\sa_count[9].r.part1[23] ,\sa_count[9].r.part1[22] 
	,\sa_count[9].r.part1[21] ,\sa_count[9].r.part1[20] 
	,\sa_count[9].r.part1[19] ,\sa_count[9].r.part1[18] 
	,\sa_count[9].r.part1[17] ,\sa_count[9].r.part1[16] 
	,\sa_count[9].r.part1[15] ,\sa_count[9].r.part1[14] 
	,\sa_count[9].r.part1[13] ,\sa_count[9].r.part1[12] 
	,\sa_count[9].r.part1[11] ,\sa_count[9].r.part1[10] 
	,\sa_count[9].r.part1[9] ,\sa_count[9].r.part1[8] 
	,\sa_count[9].r.part1[7] ,\sa_count[9].r.part1[6] 
	,\sa_count[9].r.part1[5] ,\sa_count[9].r.part1[4] 
	,\sa_count[9].r.part1[3] ,\sa_count[9].r.part1[2] 
	,\sa_count[9].r.part1[1] ,\sa_count[9].r.part1[0] 
	,\sa_count[9].r.part0[31] ,\sa_count[9].r.part0[30] 
	,\sa_count[9].r.part0[29] ,\sa_count[9].r.part0[28] 
	,\sa_count[9].r.part0[27] ,\sa_count[9].r.part0[26] 
	,\sa_count[9].r.part0[25] ,\sa_count[9].r.part0[24] 
	,\sa_count[9].r.part0[23] ,\sa_count[9].r.part0[22] 
	,\sa_count[9].r.part0[21] ,\sa_count[9].r.part0[20] 
	,\sa_count[9].r.part0[19] ,\sa_count[9].r.part0[18] 
	,\sa_count[9].r.part0[17] ,\sa_count[9].r.part0[16] 
	,\sa_count[9].r.part0[15] ,\sa_count[9].r.part0[14] 
	,\sa_count[9].r.part0[13] ,\sa_count[9].r.part0[12] 
	,\sa_count[9].r.part0[11] ,\sa_count[9].r.part0[10] 
	,\sa_count[9].r.part0[9] ,\sa_count[9].r.part0[8] 
	,\sa_count[9].r.part0[7] ,\sa_count[9].r.part0[6] 
	,\sa_count[9].r.part0[5] ,\sa_count[9].r.part0[4] 
	,\sa_count[9].r.part0[3] ,\sa_count[9].r.part0[2] 
	,\sa_count[9].r.part0[1] ,\sa_count[9].r.part0[0] 
	,\sa_count[8].r.part1[31] ,\sa_count[8].r.part1[30] 
	,\sa_count[8].r.part1[29] ,\sa_count[8].r.part1[28] 
	,\sa_count[8].r.part1[27] ,\sa_count[8].r.part1[26] 
	,\sa_count[8].r.part1[25] ,\sa_count[8].r.part1[24] 
	,\sa_count[8].r.part1[23] ,\sa_count[8].r.part1[22] 
	,\sa_count[8].r.part1[21] ,\sa_count[8].r.part1[20] 
	,\sa_count[8].r.part1[19] ,\sa_count[8].r.part1[18] 
	,\sa_count[8].r.part1[17] ,\sa_count[8].r.part1[16] 
	,\sa_count[8].r.part1[15] ,\sa_count[8].r.part1[14] 
	,\sa_count[8].r.part1[13] ,\sa_count[8].r.part1[12] 
	,\sa_count[8].r.part1[11] ,\sa_count[8].r.part1[10] 
	,\sa_count[8].r.part1[9] ,\sa_count[8].r.part1[8] 
	,\sa_count[8].r.part1[7] ,\sa_count[8].r.part1[6] 
	,\sa_count[8].r.part1[5] ,\sa_count[8].r.part1[4] 
	,\sa_count[8].r.part1[3] ,\sa_count[8].r.part1[2] 
	,\sa_count[8].r.part1[1] ,\sa_count[8].r.part1[0] 
	,\sa_count[8].r.part0[31] ,\sa_count[8].r.part0[30] 
	,\sa_count[8].r.part0[29] ,\sa_count[8].r.part0[28] 
	,\sa_count[8].r.part0[27] ,\sa_count[8].r.part0[26] 
	,\sa_count[8].r.part0[25] ,\sa_count[8].r.part0[24] 
	,\sa_count[8].r.part0[23] ,\sa_count[8].r.part0[22] 
	,\sa_count[8].r.part0[21] ,\sa_count[8].r.part0[20] 
	,\sa_count[8].r.part0[19] ,\sa_count[8].r.part0[18] 
	,\sa_count[8].r.part0[17] ,\sa_count[8].r.part0[16] 
	,\sa_count[8].r.part0[15] ,\sa_count[8].r.part0[14] 
	,\sa_count[8].r.part0[13] ,\sa_count[8].r.part0[12] 
	,\sa_count[8].r.part0[11] ,\sa_count[8].r.part0[10] 
	,\sa_count[8].r.part0[9] ,\sa_count[8].r.part0[8] 
	,\sa_count[8].r.part0[7] ,\sa_count[8].r.part0[6] 
	,\sa_count[8].r.part0[5] ,\sa_count[8].r.part0[4] 
	,\sa_count[8].r.part0[3] ,\sa_count[8].r.part0[2] 
	,\sa_count[8].r.part0[1] ,\sa_count[8].r.part0[0] 
	,\sa_count[7].r.part1[31] ,\sa_count[7].r.part1[30] 
	,\sa_count[7].r.part1[29] ,\sa_count[7].r.part1[28] 
	,\sa_count[7].r.part1[27] ,\sa_count[7].r.part1[26] 
	,\sa_count[7].r.part1[25] ,\sa_count[7].r.part1[24] 
	,\sa_count[7].r.part1[23] ,\sa_count[7].r.part1[22] 
	,\sa_count[7].r.part1[21] ,\sa_count[7].r.part1[20] 
	,\sa_count[7].r.part1[19] ,\sa_count[7].r.part1[18] 
	,\sa_count[7].r.part1[17] ,\sa_count[7].r.part1[16] 
	,\sa_count[7].r.part1[15] ,\sa_count[7].r.part1[14] 
	,\sa_count[7].r.part1[13] ,\sa_count[7].r.part1[12] 
	,\sa_count[7].r.part1[11] ,\sa_count[7].r.part1[10] 
	,\sa_count[7].r.part1[9] ,\sa_count[7].r.part1[8] 
	,\sa_count[7].r.part1[7] ,\sa_count[7].r.part1[6] 
	,\sa_count[7].r.part1[5] ,\sa_count[7].r.part1[4] 
	,\sa_count[7].r.part1[3] ,\sa_count[7].r.part1[2] 
	,\sa_count[7].r.part1[1] ,\sa_count[7].r.part1[0] 
	,\sa_count[7].r.part0[31] ,\sa_count[7].r.part0[30] 
	,\sa_count[7].r.part0[29] ,\sa_count[7].r.part0[28] 
	,\sa_count[7].r.part0[27] ,\sa_count[7].r.part0[26] 
	,\sa_count[7].r.part0[25] ,\sa_count[7].r.part0[24] 
	,\sa_count[7].r.part0[23] ,\sa_count[7].r.part0[22] 
	,\sa_count[7].r.part0[21] ,\sa_count[7].r.part0[20] 
	,\sa_count[7].r.part0[19] ,\sa_count[7].r.part0[18] 
	,\sa_count[7].r.part0[17] ,\sa_count[7].r.part0[16] 
	,\sa_count[7].r.part0[15] ,\sa_count[7].r.part0[14] 
	,\sa_count[7].r.part0[13] ,\sa_count[7].r.part0[12] 
	,\sa_count[7].r.part0[11] ,\sa_count[7].r.part0[10] 
	,\sa_count[7].r.part0[9] ,\sa_count[7].r.part0[8] 
	,\sa_count[7].r.part0[7] ,\sa_count[7].r.part0[6] 
	,\sa_count[7].r.part0[5] ,\sa_count[7].r.part0[4] 
	,\sa_count[7].r.part0[3] ,\sa_count[7].r.part0[2] 
	,\sa_count[7].r.part0[1] ,\sa_count[7].r.part0[0] 
	,\sa_count[6].r.part1[31] ,\sa_count[6].r.part1[30] 
	,\sa_count[6].r.part1[29] ,\sa_count[6].r.part1[28] 
	,\sa_count[6].r.part1[27] ,\sa_count[6].r.part1[26] 
	,\sa_count[6].r.part1[25] ,\sa_count[6].r.part1[24] 
	,\sa_count[6].r.part1[23] ,\sa_count[6].r.part1[22] 
	,\sa_count[6].r.part1[21] ,\sa_count[6].r.part1[20] 
	,\sa_count[6].r.part1[19] ,\sa_count[6].r.part1[18] 
	,\sa_count[6].r.part1[17] ,\sa_count[6].r.part1[16] 
	,\sa_count[6].r.part1[15] ,\sa_count[6].r.part1[14] 
	,\sa_count[6].r.part1[13] ,\sa_count[6].r.part1[12] 
	,\sa_count[6].r.part1[11] ,\sa_count[6].r.part1[10] 
	,\sa_count[6].r.part1[9] ,\sa_count[6].r.part1[8] 
	,\sa_count[6].r.part1[7] ,\sa_count[6].r.part1[6] 
	,\sa_count[6].r.part1[5] ,\sa_count[6].r.part1[4] 
	,\sa_count[6].r.part1[3] ,\sa_count[6].r.part1[2] 
	,\sa_count[6].r.part1[1] ,\sa_count[6].r.part1[0] 
	,\sa_count[6].r.part0[31] ,\sa_count[6].r.part0[30] 
	,\sa_count[6].r.part0[29] ,\sa_count[6].r.part0[28] 
	,\sa_count[6].r.part0[27] ,\sa_count[6].r.part0[26] 
	,\sa_count[6].r.part0[25] ,\sa_count[6].r.part0[24] 
	,\sa_count[6].r.part0[23] ,\sa_count[6].r.part0[22] 
	,\sa_count[6].r.part0[21] ,\sa_count[6].r.part0[20] 
	,\sa_count[6].r.part0[19] ,\sa_count[6].r.part0[18] 
	,\sa_count[6].r.part0[17] ,\sa_count[6].r.part0[16] 
	,\sa_count[6].r.part0[15] ,\sa_count[6].r.part0[14] 
	,\sa_count[6].r.part0[13] ,\sa_count[6].r.part0[12] 
	,\sa_count[6].r.part0[11] ,\sa_count[6].r.part0[10] 
	,\sa_count[6].r.part0[9] ,\sa_count[6].r.part0[8] 
	,\sa_count[6].r.part0[7] ,\sa_count[6].r.part0[6] 
	,\sa_count[6].r.part0[5] ,\sa_count[6].r.part0[4] 
	,\sa_count[6].r.part0[3] ,\sa_count[6].r.part0[2] 
	,\sa_count[6].r.part0[1] ,\sa_count[6].r.part0[0] 
	,\sa_count[5].r.part1[31] ,\sa_count[5].r.part1[30] 
	,\sa_count[5].r.part1[29] ,\sa_count[5].r.part1[28] 
	,\sa_count[5].r.part1[27] ,\sa_count[5].r.part1[26] 
	,\sa_count[5].r.part1[25] ,\sa_count[5].r.part1[24] 
	,\sa_count[5].r.part1[23] ,\sa_count[5].r.part1[22] 
	,\sa_count[5].r.part1[21] ,\sa_count[5].r.part1[20] 
	,\sa_count[5].r.part1[19] ,\sa_count[5].r.part1[18] 
	,\sa_count[5].r.part1[17] ,\sa_count[5].r.part1[16] 
	,\sa_count[5].r.part1[15] ,\sa_count[5].r.part1[14] 
	,\sa_count[5].r.part1[13] ,\sa_count[5].r.part1[12] 
	,\sa_count[5].r.part1[11] ,\sa_count[5].r.part1[10] 
	,\sa_count[5].r.part1[9] ,\sa_count[5].r.part1[8] 
	,\sa_count[5].r.part1[7] ,\sa_count[5].r.part1[6] 
	,\sa_count[5].r.part1[5] ,\sa_count[5].r.part1[4] 
	,\sa_count[5].r.part1[3] ,\sa_count[5].r.part1[2] 
	,\sa_count[5].r.part1[1] ,\sa_count[5].r.part1[0] 
	,\sa_count[5].r.part0[31] ,\sa_count[5].r.part0[30] 
	,\sa_count[5].r.part0[29] ,\sa_count[5].r.part0[28] 
	,\sa_count[5].r.part0[27] ,\sa_count[5].r.part0[26] 
	,\sa_count[5].r.part0[25] ,\sa_count[5].r.part0[24] 
	,\sa_count[5].r.part0[23] ,\sa_count[5].r.part0[22] 
	,\sa_count[5].r.part0[21] ,\sa_count[5].r.part0[20] 
	,\sa_count[5].r.part0[19] ,\sa_count[5].r.part0[18] 
	,\sa_count[5].r.part0[17] ,\sa_count[5].r.part0[16] 
	,\sa_count[5].r.part0[15] ,\sa_count[5].r.part0[14] 
	,\sa_count[5].r.part0[13] ,\sa_count[5].r.part0[12] 
	,\sa_count[5].r.part0[11] ,\sa_count[5].r.part0[10] 
	,\sa_count[5].r.part0[9] ,\sa_count[5].r.part0[8] 
	,\sa_count[5].r.part0[7] ,\sa_count[5].r.part0[6] 
	,\sa_count[5].r.part0[5] ,\sa_count[5].r.part0[4] 
	,\sa_count[5].r.part0[3] ,\sa_count[5].r.part0[2] 
	,\sa_count[5].r.part0[1] ,\sa_count[5].r.part0[0] 
	,\sa_count[4].r.part1[31] ,\sa_count[4].r.part1[30] 
	,\sa_count[4].r.part1[29] ,\sa_count[4].r.part1[28] 
	,\sa_count[4].r.part1[27] ,\sa_count[4].r.part1[26] 
	,\sa_count[4].r.part1[25] ,\sa_count[4].r.part1[24] 
	,\sa_count[4].r.part1[23] ,\sa_count[4].r.part1[22] 
	,\sa_count[4].r.part1[21] ,\sa_count[4].r.part1[20] 
	,\sa_count[4].r.part1[19] ,\sa_count[4].r.part1[18] 
	,\sa_count[4].r.part1[17] ,\sa_count[4].r.part1[16] 
	,\sa_count[4].r.part1[15] ,\sa_count[4].r.part1[14] 
	,\sa_count[4].r.part1[13] ,\sa_count[4].r.part1[12] 
	,\sa_count[4].r.part1[11] ,\sa_count[4].r.part1[10] 
	,\sa_count[4].r.part1[9] ,\sa_count[4].r.part1[8] 
	,\sa_count[4].r.part1[7] ,\sa_count[4].r.part1[6] 
	,\sa_count[4].r.part1[5] ,\sa_count[4].r.part1[4] 
	,\sa_count[4].r.part1[3] ,\sa_count[4].r.part1[2] 
	,\sa_count[4].r.part1[1] ,\sa_count[4].r.part1[0] 
	,\sa_count[4].r.part0[31] ,\sa_count[4].r.part0[30] 
	,\sa_count[4].r.part0[29] ,\sa_count[4].r.part0[28] 
	,\sa_count[4].r.part0[27] ,\sa_count[4].r.part0[26] 
	,\sa_count[4].r.part0[25] ,\sa_count[4].r.part0[24] 
	,\sa_count[4].r.part0[23] ,\sa_count[4].r.part0[22] 
	,\sa_count[4].r.part0[21] ,\sa_count[4].r.part0[20] 
	,\sa_count[4].r.part0[19] ,\sa_count[4].r.part0[18] 
	,\sa_count[4].r.part0[17] ,\sa_count[4].r.part0[16] 
	,\sa_count[4].r.part0[15] ,\sa_count[4].r.part0[14] 
	,\sa_count[4].r.part0[13] ,\sa_count[4].r.part0[12] 
	,\sa_count[4].r.part0[11] ,\sa_count[4].r.part0[10] 
	,\sa_count[4].r.part0[9] ,\sa_count[4].r.part0[8] 
	,\sa_count[4].r.part0[7] ,\sa_count[4].r.part0[6] 
	,\sa_count[4].r.part0[5] ,\sa_count[4].r.part0[4] 
	,\sa_count[4].r.part0[3] ,\sa_count[4].r.part0[2] 
	,\sa_count[4].r.part0[1] ,\sa_count[4].r.part0[0] 
	,\sa_count[3].r.part1[31] ,\sa_count[3].r.part1[30] 
	,\sa_count[3].r.part1[29] ,\sa_count[3].r.part1[28] 
	,\sa_count[3].r.part1[27] ,\sa_count[3].r.part1[26] 
	,\sa_count[3].r.part1[25] ,\sa_count[3].r.part1[24] 
	,\sa_count[3].r.part1[23] ,\sa_count[3].r.part1[22] 
	,\sa_count[3].r.part1[21] ,\sa_count[3].r.part1[20] 
	,\sa_count[3].r.part1[19] ,\sa_count[3].r.part1[18] 
	,\sa_count[3].r.part1[17] ,\sa_count[3].r.part1[16] 
	,\sa_count[3].r.part1[15] ,\sa_count[3].r.part1[14] 
	,\sa_count[3].r.part1[13] ,\sa_count[3].r.part1[12] 
	,\sa_count[3].r.part1[11] ,\sa_count[3].r.part1[10] 
	,\sa_count[3].r.part1[9] ,\sa_count[3].r.part1[8] 
	,\sa_count[3].r.part1[7] ,\sa_count[3].r.part1[6] 
	,\sa_count[3].r.part1[5] ,\sa_count[3].r.part1[4] 
	,\sa_count[3].r.part1[3] ,\sa_count[3].r.part1[2] 
	,\sa_count[3].r.part1[1] ,\sa_count[3].r.part1[0] 
	,\sa_count[3].r.part0[31] ,\sa_count[3].r.part0[30] 
	,\sa_count[3].r.part0[29] ,\sa_count[3].r.part0[28] 
	,\sa_count[3].r.part0[27] ,\sa_count[3].r.part0[26] 
	,\sa_count[3].r.part0[25] ,\sa_count[3].r.part0[24] 
	,\sa_count[3].r.part0[23] ,\sa_count[3].r.part0[22] 
	,\sa_count[3].r.part0[21] ,\sa_count[3].r.part0[20] 
	,\sa_count[3].r.part0[19] ,\sa_count[3].r.part0[18] 
	,\sa_count[3].r.part0[17] ,\sa_count[3].r.part0[16] 
	,\sa_count[3].r.part0[15] ,\sa_count[3].r.part0[14] 
	,\sa_count[3].r.part0[13] ,\sa_count[3].r.part0[12] 
	,\sa_count[3].r.part0[11] ,\sa_count[3].r.part0[10] 
	,\sa_count[3].r.part0[9] ,\sa_count[3].r.part0[8] 
	,\sa_count[3].r.part0[7] ,\sa_count[3].r.part0[6] 
	,\sa_count[3].r.part0[5] ,\sa_count[3].r.part0[4] 
	,\sa_count[3].r.part0[3] ,\sa_count[3].r.part0[2] 
	,\sa_count[3].r.part0[1] ,\sa_count[3].r.part0[0] 
	,\sa_count[2].r.part1[31] ,\sa_count[2].r.part1[30] 
	,\sa_count[2].r.part1[29] ,\sa_count[2].r.part1[28] 
	,\sa_count[2].r.part1[27] ,\sa_count[2].r.part1[26] 
	,\sa_count[2].r.part1[25] ,\sa_count[2].r.part1[24] 
	,\sa_count[2].r.part1[23] ,\sa_count[2].r.part1[22] 
	,\sa_count[2].r.part1[21] ,\sa_count[2].r.part1[20] 
	,\sa_count[2].r.part1[19] ,\sa_count[2].r.part1[18] 
	,\sa_count[2].r.part1[17] ,\sa_count[2].r.part1[16] 
	,\sa_count[2].r.part1[15] ,\sa_count[2].r.part1[14] 
	,\sa_count[2].r.part1[13] ,\sa_count[2].r.part1[12] 
	,\sa_count[2].r.part1[11] ,\sa_count[2].r.part1[10] 
	,\sa_count[2].r.part1[9] ,\sa_count[2].r.part1[8] 
	,\sa_count[2].r.part1[7] ,\sa_count[2].r.part1[6] 
	,\sa_count[2].r.part1[5] ,\sa_count[2].r.part1[4] 
	,\sa_count[2].r.part1[3] ,\sa_count[2].r.part1[2] 
	,\sa_count[2].r.part1[1] ,\sa_count[2].r.part1[0] 
	,\sa_count[2].r.part0[31] ,\sa_count[2].r.part0[30] 
	,\sa_count[2].r.part0[29] ,\sa_count[2].r.part0[28] 
	,\sa_count[2].r.part0[27] ,\sa_count[2].r.part0[26] 
	,\sa_count[2].r.part0[25] ,\sa_count[2].r.part0[24] 
	,\sa_count[2].r.part0[23] ,\sa_count[2].r.part0[22] 
	,\sa_count[2].r.part0[21] ,\sa_count[2].r.part0[20] 
	,\sa_count[2].r.part0[19] ,\sa_count[2].r.part0[18] 
	,\sa_count[2].r.part0[17] ,\sa_count[2].r.part0[16] 
	,\sa_count[2].r.part0[15] ,\sa_count[2].r.part0[14] 
	,\sa_count[2].r.part0[13] ,\sa_count[2].r.part0[12] 
	,\sa_count[2].r.part0[11] ,\sa_count[2].r.part0[10] 
	,\sa_count[2].r.part0[9] ,\sa_count[2].r.part0[8] 
	,\sa_count[2].r.part0[7] ,\sa_count[2].r.part0[6] 
	,\sa_count[2].r.part0[5] ,\sa_count[2].r.part0[4] 
	,\sa_count[2].r.part0[3] ,\sa_count[2].r.part0[2] 
	,\sa_count[2].r.part0[1] ,\sa_count[2].r.part0[0] 
	,\sa_count[1].r.part1[31] ,\sa_count[1].r.part1[30] 
	,\sa_count[1].r.part1[29] ,\sa_count[1].r.part1[28] 
	,\sa_count[1].r.part1[27] ,\sa_count[1].r.part1[26] 
	,\sa_count[1].r.part1[25] ,\sa_count[1].r.part1[24] 
	,\sa_count[1].r.part1[23] ,\sa_count[1].r.part1[22] 
	,\sa_count[1].r.part1[21] ,\sa_count[1].r.part1[20] 
	,\sa_count[1].r.part1[19] ,\sa_count[1].r.part1[18] 
	,\sa_count[1].r.part1[17] ,\sa_count[1].r.part1[16] 
	,\sa_count[1].r.part1[15] ,\sa_count[1].r.part1[14] 
	,\sa_count[1].r.part1[13] ,\sa_count[1].r.part1[12] 
	,\sa_count[1].r.part1[11] ,\sa_count[1].r.part1[10] 
	,\sa_count[1].r.part1[9] ,\sa_count[1].r.part1[8] 
	,\sa_count[1].r.part1[7] ,\sa_count[1].r.part1[6] 
	,\sa_count[1].r.part1[5] ,\sa_count[1].r.part1[4] 
	,\sa_count[1].r.part1[3] ,\sa_count[1].r.part1[2] 
	,\sa_count[1].r.part1[1] ,\sa_count[1].r.part1[0] 
	,\sa_count[1].r.part0[31] ,\sa_count[1].r.part0[30] 
	,\sa_count[1].r.part0[29] ,\sa_count[1].r.part0[28] 
	,\sa_count[1].r.part0[27] ,\sa_count[1].r.part0[26] 
	,\sa_count[1].r.part0[25] ,\sa_count[1].r.part0[24] 
	,\sa_count[1].r.part0[23] ,\sa_count[1].r.part0[22] 
	,\sa_count[1].r.part0[21] ,\sa_count[1].r.part0[20] 
	,\sa_count[1].r.part0[19] ,\sa_count[1].r.part0[18] 
	,\sa_count[1].r.part0[17] ,\sa_count[1].r.part0[16] 
	,\sa_count[1].r.part0[15] ,\sa_count[1].r.part0[14] 
	,\sa_count[1].r.part0[13] ,\sa_count[1].r.part0[12] 
	,\sa_count[1].r.part0[11] ,\sa_count[1].r.part0[10] 
	,\sa_count[1].r.part0[9] ,\sa_count[1].r.part0[8] 
	,\sa_count[1].r.part0[7] ,\sa_count[1].r.part0[6] 
	,\sa_count[1].r.part0[5] ,\sa_count[1].r.part0[4] 
	,\sa_count[1].r.part0[3] ,\sa_count[1].r.part0[2] 
	,\sa_count[1].r.part0[1] ,\sa_count[1].r.part0[0] 
	,\sa_count[0].r.part1[31] ,\sa_count[0].r.part1[30] 
	,\sa_count[0].r.part1[29] ,\sa_count[0].r.part1[28] 
	,\sa_count[0].r.part1[27] ,\sa_count[0].r.part1[26] 
	,\sa_count[0].r.part1[25] ,\sa_count[0].r.part1[24] 
	,\sa_count[0].r.part1[23] ,\sa_count[0].r.part1[22] 
	,\sa_count[0].r.part1[21] ,\sa_count[0].r.part1[20] 
	,\sa_count[0].r.part1[19] ,\sa_count[0].r.part1[18] 
	,\sa_count[0].r.part1[17] ,\sa_count[0].r.part1[16] 
	,\sa_count[0].r.part1[15] ,\sa_count[0].r.part1[14] 
	,\sa_count[0].r.part1[13] ,\sa_count[0].r.part1[12] 
	,\sa_count[0].r.part1[11] ,\sa_count[0].r.part1[10] 
	,\sa_count[0].r.part1[9] ,\sa_count[0].r.part1[8] 
	,\sa_count[0].r.part1[7] ,\sa_count[0].r.part1[6] 
	,\sa_count[0].r.part1[5] ,\sa_count[0].r.part1[4] 
	,\sa_count[0].r.part1[3] ,\sa_count[0].r.part1[2] 
	,\sa_count[0].r.part1[1] ,\sa_count[0].r.part1[0] 
	,\sa_count[0].r.part0[31] ,\sa_count[0].r.part0[30] 
	,\sa_count[0].r.part0[29] ,\sa_count[0].r.part0[28] 
	,\sa_count[0].r.part0[27] ,\sa_count[0].r.part0[26] 
	,\sa_count[0].r.part0[25] ,\sa_count[0].r.part0[24] 
	,\sa_count[0].r.part0[23] ,\sa_count[0].r.part0[22] 
	,\sa_count[0].r.part0[21] ,\sa_count[0].r.part0[20] 
	,\sa_count[0].r.part0[19] ,\sa_count[0].r.part0[18] 
	,\sa_count[0].r.part0[17] ,\sa_count[0].r.part0[16] 
	,\sa_count[0].r.part0[15] ,\sa_count[0].r.part0[14] 
	,\sa_count[0].r.part0[13] ,\sa_count[0].r.part0[12] 
	,\sa_count[0].r.part0[11] ,\sa_count[0].r.part0[10] 
	,\sa_count[0].r.part0[9] ,\sa_count[0].r.part0[8] 
	,\sa_count[0].r.part0[7] ,\sa_count[0].r.part0[6] 
	,\sa_count[0].r.part0[5] ,\sa_count[0].r.part0[4] 
	,\sa_count[0].r.part0[3] ,\sa_count[0].r.part0[2] 
	,\sa_count[0].r.part0[1] ,\sa_count[0].r.part0[0] ;
output kme_idle;
output [31:0] \idle_components.r.part0 ;
wire [19:0] \idle_components.f.num_key_tlvs_in_flight ;
wire \idle_components.f.cddip0_key_tlv_rsm_idle ;
wire \idle_components.f.cddip1_key_tlv_rsm_idle ;
wire \idle_components.f.cddip2_key_tlv_rsm_idle ;
wire \idle_components.f.cddip3_key_tlv_rsm_idle ;
wire \idle_components.f.cceip0_key_tlv_rsm_idle ;
wire \idle_components.f.cceip1_key_tlv_rsm_idle ;
wire \idle_components.f.cceip2_key_tlv_rsm_idle ;
wire \idle_components.f.cceip3_key_tlv_rsm_idle ;
wire \idle_components.f.no_key_tlv_in_flight ;
wire \idle_components.f.tlv_parser_idle ;
wire \idle_components.f.drng_idle ;
wire \idle_components.f.kme_slv_empty ;
wire [31:0] idle_components;
input clk;
input rst_n;
input disable_debug_cmd;
input cceip_encrypt_gcm_tag_fail_int;
input cceip_validate_gcm_tag_fail_int;
input cddip_decrypt_gcm_tag_fail_int;
input [3:0] cceip_ob_full;
input [3:0] cddip_ob_full;
input [8:0] \tready_override.r.part0 ;
wire \tready_override.f.txc_tready_override ;
wire \tready_override.f.engine_7_tready_override ;
wire \tready_override.f.engine_6_tready_override ;
wire \tready_override.f.engine_5_tready_override ;
wire \tready_override.f.engine_4_tready_override ;
wire \tready_override.f.engine_3_tready_override ;
wire \tready_override.f.engine_2_tready_override ;
wire \tready_override.f.engine_1_tready_override ;
wire \tready_override.f.engine_0_tready_override ;
wire [8:0] tready_override;
input \core_kme_ib_out.tready ;
wire [0:0] core_kme_ib_out;
input [31:0] \sa_global_ctrl.r.part0 ;
wire [29:0] \sa_global_ctrl.f.spare ;
wire \sa_global_ctrl.f.sa_snap ;
wire \sa_global_ctrl.f.sa_clear_live ;
wire [31:0] sa_global_ctrl;
input \sa_ctrl[31].r.part0[31] ,\sa_ctrl[31].r.part0[30] 
	,\sa_ctrl[31].r.part0[29] ,\sa_ctrl[31].r.part0[28] 
	,\sa_ctrl[31].r.part0[27] ,\sa_ctrl[31].r.part0[26] 
	,\sa_ctrl[31].r.part0[25] ,\sa_ctrl[31].r.part0[24] 
	,\sa_ctrl[31].r.part0[23] ,\sa_ctrl[31].r.part0[22] 
	,\sa_ctrl[31].r.part0[21] ,\sa_ctrl[31].r.part0[20] 
	,\sa_ctrl[31].r.part0[19] ,\sa_ctrl[31].r.part0[18] 
	,\sa_ctrl[31].r.part0[17] ,\sa_ctrl[31].r.part0[16] 
	,\sa_ctrl[31].r.part0[15] ,\sa_ctrl[31].r.part0[14] 
	,\sa_ctrl[31].r.part0[13] ,\sa_ctrl[31].r.part0[12] 
	,\sa_ctrl[31].r.part0[11] ,\sa_ctrl[31].r.part0[10] 
	,\sa_ctrl[31].r.part0[9] ,\sa_ctrl[31].r.part0[8] 
	,\sa_ctrl[31].r.part0[7] ,\sa_ctrl[31].r.part0[6] 
	,\sa_ctrl[31].r.part0[5] ,\sa_ctrl[31].r.part0[4] 
	,\sa_ctrl[31].r.part0[3] ,\sa_ctrl[31].r.part0[2] 
	,\sa_ctrl[31].r.part0[1] ,\sa_ctrl[31].r.part0[0] 
	,\sa_ctrl[30].r.part0[31] ,\sa_ctrl[30].r.part0[30] 
	,\sa_ctrl[30].r.part0[29] ,\sa_ctrl[30].r.part0[28] 
	,\sa_ctrl[30].r.part0[27] ,\sa_ctrl[30].r.part0[26] 
	,\sa_ctrl[30].r.part0[25] ,\sa_ctrl[30].r.part0[24] 
	,\sa_ctrl[30].r.part0[23] ,\sa_ctrl[30].r.part0[22] 
	,\sa_ctrl[30].r.part0[21] ,\sa_ctrl[30].r.part0[20] 
	,\sa_ctrl[30].r.part0[19] ,\sa_ctrl[30].r.part0[18] 
	,\sa_ctrl[30].r.part0[17] ,\sa_ctrl[30].r.part0[16] 
	,\sa_ctrl[30].r.part0[15] ,\sa_ctrl[30].r.part0[14] 
	,\sa_ctrl[30].r.part0[13] ,\sa_ctrl[30].r.part0[12] 
	,\sa_ctrl[30].r.part0[11] ,\sa_ctrl[30].r.part0[10] 
	,\sa_ctrl[30].r.part0[9] ,\sa_ctrl[30].r.part0[8] 
	,\sa_ctrl[30].r.part0[7] ,\sa_ctrl[30].r.part0[6] 
	,\sa_ctrl[30].r.part0[5] ,\sa_ctrl[30].r.part0[4] 
	,\sa_ctrl[30].r.part0[3] ,\sa_ctrl[30].r.part0[2] 
	,\sa_ctrl[30].r.part0[1] ,\sa_ctrl[30].r.part0[0] 
	,\sa_ctrl[29].r.part0[31] ,\sa_ctrl[29].r.part0[30] 
	,\sa_ctrl[29].r.part0[29] ,\sa_ctrl[29].r.part0[28] 
	,\sa_ctrl[29].r.part0[27] ,\sa_ctrl[29].r.part0[26] 
	,\sa_ctrl[29].r.part0[25] ,\sa_ctrl[29].r.part0[24] 
	,\sa_ctrl[29].r.part0[23] ,\sa_ctrl[29].r.part0[22] 
	,\sa_ctrl[29].r.part0[21] ,\sa_ctrl[29].r.part0[20] 
	,\sa_ctrl[29].r.part0[19] ,\sa_ctrl[29].r.part0[18] 
	,\sa_ctrl[29].r.part0[17] ,\sa_ctrl[29].r.part0[16] 
	,\sa_ctrl[29].r.part0[15] ,\sa_ctrl[29].r.part0[14] 
	,\sa_ctrl[29].r.part0[13] ,\sa_ctrl[29].r.part0[12] 
	,\sa_ctrl[29].r.part0[11] ,\sa_ctrl[29].r.part0[10] 
	,\sa_ctrl[29].r.part0[9] ,\sa_ctrl[29].r.part0[8] 
	,\sa_ctrl[29].r.part0[7] ,\sa_ctrl[29].r.part0[6] 
	,\sa_ctrl[29].r.part0[5] ,\sa_ctrl[29].r.part0[4] 
	,\sa_ctrl[29].r.part0[3] ,\sa_ctrl[29].r.part0[2] 
	,\sa_ctrl[29].r.part0[1] ,\sa_ctrl[29].r.part0[0] 
	,\sa_ctrl[28].r.part0[31] ,\sa_ctrl[28].r.part0[30] 
	,\sa_ctrl[28].r.part0[29] ,\sa_ctrl[28].r.part0[28] 
	,\sa_ctrl[28].r.part0[27] ,\sa_ctrl[28].r.part0[26] 
	,\sa_ctrl[28].r.part0[25] ,\sa_ctrl[28].r.part0[24] 
	,\sa_ctrl[28].r.part0[23] ,\sa_ctrl[28].r.part0[22] 
	,\sa_ctrl[28].r.part0[21] ,\sa_ctrl[28].r.part0[20] 
	,\sa_ctrl[28].r.part0[19] ,\sa_ctrl[28].r.part0[18] 
	,\sa_ctrl[28].r.part0[17] ,\sa_ctrl[28].r.part0[16] 
	,\sa_ctrl[28].r.part0[15] ,\sa_ctrl[28].r.part0[14] 
	,\sa_ctrl[28].r.part0[13] ,\sa_ctrl[28].r.part0[12] 
	,\sa_ctrl[28].r.part0[11] ,\sa_ctrl[28].r.part0[10] 
	,\sa_ctrl[28].r.part0[9] ,\sa_ctrl[28].r.part0[8] 
	,\sa_ctrl[28].r.part0[7] ,\sa_ctrl[28].r.part0[6] 
	,\sa_ctrl[28].r.part0[5] ,\sa_ctrl[28].r.part0[4] 
	,\sa_ctrl[28].r.part0[3] ,\sa_ctrl[28].r.part0[2] 
	,\sa_ctrl[28].r.part0[1] ,\sa_ctrl[28].r.part0[0] 
	,\sa_ctrl[27].r.part0[31] ,\sa_ctrl[27].r.part0[30] 
	,\sa_ctrl[27].r.part0[29] ,\sa_ctrl[27].r.part0[28] 
	,\sa_ctrl[27].r.part0[27] ,\sa_ctrl[27].r.part0[26] 
	,\sa_ctrl[27].r.part0[25] ,\sa_ctrl[27].r.part0[24] 
	,\sa_ctrl[27].r.part0[23] ,\sa_ctrl[27].r.part0[22] 
	,\sa_ctrl[27].r.part0[21] ,\sa_ctrl[27].r.part0[20] 
	,\sa_ctrl[27].r.part0[19] ,\sa_ctrl[27].r.part0[18] 
	,\sa_ctrl[27].r.part0[17] ,\sa_ctrl[27].r.part0[16] 
	,\sa_ctrl[27].r.part0[15] ,\sa_ctrl[27].r.part0[14] 
	,\sa_ctrl[27].r.part0[13] ,\sa_ctrl[27].r.part0[12] 
	,\sa_ctrl[27].r.part0[11] ,\sa_ctrl[27].r.part0[10] 
	,\sa_ctrl[27].r.part0[9] ,\sa_ctrl[27].r.part0[8] 
	,\sa_ctrl[27].r.part0[7] ,\sa_ctrl[27].r.part0[6] 
	,\sa_ctrl[27].r.part0[5] ,\sa_ctrl[27].r.part0[4] 
	,\sa_ctrl[27].r.part0[3] ,\sa_ctrl[27].r.part0[2] 
	,\sa_ctrl[27].r.part0[1] ,\sa_ctrl[27].r.part0[0] 
	,\sa_ctrl[26].r.part0[31] ,\sa_ctrl[26].r.part0[30] 
	,\sa_ctrl[26].r.part0[29] ,\sa_ctrl[26].r.part0[28] 
	,\sa_ctrl[26].r.part0[27] ,\sa_ctrl[26].r.part0[26] 
	,\sa_ctrl[26].r.part0[25] ,\sa_ctrl[26].r.part0[24] 
	,\sa_ctrl[26].r.part0[23] ,\sa_ctrl[26].r.part0[22] 
	,\sa_ctrl[26].r.part0[21] ,\sa_ctrl[26].r.part0[20] 
	,\sa_ctrl[26].r.part0[19] ,\sa_ctrl[26].r.part0[18] 
	,\sa_ctrl[26].r.part0[17] ,\sa_ctrl[26].r.part0[16] 
	,\sa_ctrl[26].r.part0[15] ,\sa_ctrl[26].r.part0[14] 
	,\sa_ctrl[26].r.part0[13] ,\sa_ctrl[26].r.part0[12] 
	,\sa_ctrl[26].r.part0[11] ,\sa_ctrl[26].r.part0[10] 
	,\sa_ctrl[26].r.part0[9] ,\sa_ctrl[26].r.part0[8] 
	,\sa_ctrl[26].r.part0[7] ,\sa_ctrl[26].r.part0[6] 
	,\sa_ctrl[26].r.part0[5] ,\sa_ctrl[26].r.part0[4] 
	,\sa_ctrl[26].r.part0[3] ,\sa_ctrl[26].r.part0[2] 
	,\sa_ctrl[26].r.part0[1] ,\sa_ctrl[26].r.part0[0] 
	,\sa_ctrl[25].r.part0[31] ,\sa_ctrl[25].r.part0[30] 
	,\sa_ctrl[25].r.part0[29] ,\sa_ctrl[25].r.part0[28] 
	,\sa_ctrl[25].r.part0[27] ,\sa_ctrl[25].r.part0[26] 
	,\sa_ctrl[25].r.part0[25] ,\sa_ctrl[25].r.part0[24] 
	,\sa_ctrl[25].r.part0[23] ,\sa_ctrl[25].r.part0[22] 
	,\sa_ctrl[25].r.part0[21] ,\sa_ctrl[25].r.part0[20] 
	,\sa_ctrl[25].r.part0[19] ,\sa_ctrl[25].r.part0[18] 
	,\sa_ctrl[25].r.part0[17] ,\sa_ctrl[25].r.part0[16] 
	,\sa_ctrl[25].r.part0[15] ,\sa_ctrl[25].r.part0[14] 
	,\sa_ctrl[25].r.part0[13] ,\sa_ctrl[25].r.part0[12] 
	,\sa_ctrl[25].r.part0[11] ,\sa_ctrl[25].r.part0[10] 
	,\sa_ctrl[25].r.part0[9] ,\sa_ctrl[25].r.part0[8] 
	,\sa_ctrl[25].r.part0[7] ,\sa_ctrl[25].r.part0[6] 
	,\sa_ctrl[25].r.part0[5] ,\sa_ctrl[25].r.part0[4] 
	,\sa_ctrl[25].r.part0[3] ,\sa_ctrl[25].r.part0[2] 
	,\sa_ctrl[25].r.part0[1] ,\sa_ctrl[25].r.part0[0] 
	,\sa_ctrl[24].r.part0[31] ,\sa_ctrl[24].r.part0[30] 
	,\sa_ctrl[24].r.part0[29] ,\sa_ctrl[24].r.part0[28] 
	,\sa_ctrl[24].r.part0[27] ,\sa_ctrl[24].r.part0[26] 
	,\sa_ctrl[24].r.part0[25] ,\sa_ctrl[24].r.part0[24] 
	,\sa_ctrl[24].r.part0[23] ,\sa_ctrl[24].r.part0[22] 
	,\sa_ctrl[24].r.part0[21] ,\sa_ctrl[24].r.part0[20] 
	,\sa_ctrl[24].r.part0[19] ,\sa_ctrl[24].r.part0[18] 
	,\sa_ctrl[24].r.part0[17] ,\sa_ctrl[24].r.part0[16] 
	,\sa_ctrl[24].r.part0[15] ,\sa_ctrl[24].r.part0[14] 
	,\sa_ctrl[24].r.part0[13] ,\sa_ctrl[24].r.part0[12] 
	,\sa_ctrl[24].r.part0[11] ,\sa_ctrl[24].r.part0[10] 
	,\sa_ctrl[24].r.part0[9] ,\sa_ctrl[24].r.part0[8] 
	,\sa_ctrl[24].r.part0[7] ,\sa_ctrl[24].r.part0[6] 
	,\sa_ctrl[24].r.part0[5] ,\sa_ctrl[24].r.part0[4] 
	,\sa_ctrl[24].r.part0[3] ,\sa_ctrl[24].r.part0[2] 
	,\sa_ctrl[24].r.part0[1] ,\sa_ctrl[24].r.part0[0] 
	,\sa_ctrl[23].r.part0[31] ,\sa_ctrl[23].r.part0[30] 
	,\sa_ctrl[23].r.part0[29] ,\sa_ctrl[23].r.part0[28] 
	,\sa_ctrl[23].r.part0[27] ,\sa_ctrl[23].r.part0[26] 
	,\sa_ctrl[23].r.part0[25] ,\sa_ctrl[23].r.part0[24] 
	,\sa_ctrl[23].r.part0[23] ,\sa_ctrl[23].r.part0[22] 
	,\sa_ctrl[23].r.part0[21] ,\sa_ctrl[23].r.part0[20] 
	,\sa_ctrl[23].r.part0[19] ,\sa_ctrl[23].r.part0[18] 
	,\sa_ctrl[23].r.part0[17] ,\sa_ctrl[23].r.part0[16] 
	,\sa_ctrl[23].r.part0[15] ,\sa_ctrl[23].r.part0[14] 
	,\sa_ctrl[23].r.part0[13] ,\sa_ctrl[23].r.part0[12] 
	,\sa_ctrl[23].r.part0[11] ,\sa_ctrl[23].r.part0[10] 
	,\sa_ctrl[23].r.part0[9] ,\sa_ctrl[23].r.part0[8] 
	,\sa_ctrl[23].r.part0[7] ,\sa_ctrl[23].r.part0[6] 
	,\sa_ctrl[23].r.part0[5] ,\sa_ctrl[23].r.part0[4] 
	,\sa_ctrl[23].r.part0[3] ,\sa_ctrl[23].r.part0[2] 
	,\sa_ctrl[23].r.part0[1] ,\sa_ctrl[23].r.part0[0] 
	,\sa_ctrl[22].r.part0[31] ,\sa_ctrl[22].r.part0[30] 
	,\sa_ctrl[22].r.part0[29] ,\sa_ctrl[22].r.part0[28] 
	,\sa_ctrl[22].r.part0[27] ,\sa_ctrl[22].r.part0[26] 
	,\sa_ctrl[22].r.part0[25] ,\sa_ctrl[22].r.part0[24] 
	,\sa_ctrl[22].r.part0[23] ,\sa_ctrl[22].r.part0[22] 
	,\sa_ctrl[22].r.part0[21] ,\sa_ctrl[22].r.part0[20] 
	,\sa_ctrl[22].r.part0[19] ,\sa_ctrl[22].r.part0[18] 
	,\sa_ctrl[22].r.part0[17] ,\sa_ctrl[22].r.part0[16] 
	,\sa_ctrl[22].r.part0[15] ,\sa_ctrl[22].r.part0[14] 
	,\sa_ctrl[22].r.part0[13] ,\sa_ctrl[22].r.part0[12] 
	,\sa_ctrl[22].r.part0[11] ,\sa_ctrl[22].r.part0[10] 
	,\sa_ctrl[22].r.part0[9] ,\sa_ctrl[22].r.part0[8] 
	,\sa_ctrl[22].r.part0[7] ,\sa_ctrl[22].r.part0[6] 
	,\sa_ctrl[22].r.part0[5] ,\sa_ctrl[22].r.part0[4] 
	,\sa_ctrl[22].r.part0[3] ,\sa_ctrl[22].r.part0[2] 
	,\sa_ctrl[22].r.part0[1] ,\sa_ctrl[22].r.part0[0] 
	,\sa_ctrl[21].r.part0[31] ,\sa_ctrl[21].r.part0[30] 
	,\sa_ctrl[21].r.part0[29] ,\sa_ctrl[21].r.part0[28] 
	,\sa_ctrl[21].r.part0[27] ,\sa_ctrl[21].r.part0[26] 
	,\sa_ctrl[21].r.part0[25] ,\sa_ctrl[21].r.part0[24] 
	,\sa_ctrl[21].r.part0[23] ,\sa_ctrl[21].r.part0[22] 
	,\sa_ctrl[21].r.part0[21] ,\sa_ctrl[21].r.part0[20] 
	,\sa_ctrl[21].r.part0[19] ,\sa_ctrl[21].r.part0[18] 
	,\sa_ctrl[21].r.part0[17] ,\sa_ctrl[21].r.part0[16] 
	,\sa_ctrl[21].r.part0[15] ,\sa_ctrl[21].r.part0[14] 
	,\sa_ctrl[21].r.part0[13] ,\sa_ctrl[21].r.part0[12] 
	,\sa_ctrl[21].r.part0[11] ,\sa_ctrl[21].r.part0[10] 
	,\sa_ctrl[21].r.part0[9] ,\sa_ctrl[21].r.part0[8] 
	,\sa_ctrl[21].r.part0[7] ,\sa_ctrl[21].r.part0[6] 
	,\sa_ctrl[21].r.part0[5] ,\sa_ctrl[21].r.part0[4] 
	,\sa_ctrl[21].r.part0[3] ,\sa_ctrl[21].r.part0[2] 
	,\sa_ctrl[21].r.part0[1] ,\sa_ctrl[21].r.part0[0] 
	,\sa_ctrl[20].r.part0[31] ,\sa_ctrl[20].r.part0[30] 
	,\sa_ctrl[20].r.part0[29] ,\sa_ctrl[20].r.part0[28] 
	,\sa_ctrl[20].r.part0[27] ,\sa_ctrl[20].r.part0[26] 
	,\sa_ctrl[20].r.part0[25] ,\sa_ctrl[20].r.part0[24] 
	,\sa_ctrl[20].r.part0[23] ,\sa_ctrl[20].r.part0[22] 
	,\sa_ctrl[20].r.part0[21] ,\sa_ctrl[20].r.part0[20] 
	,\sa_ctrl[20].r.part0[19] ,\sa_ctrl[20].r.part0[18] 
	,\sa_ctrl[20].r.part0[17] ,\sa_ctrl[20].r.part0[16] 
	,\sa_ctrl[20].r.part0[15] ,\sa_ctrl[20].r.part0[14] 
	,\sa_ctrl[20].r.part0[13] ,\sa_ctrl[20].r.part0[12] 
	,\sa_ctrl[20].r.part0[11] ,\sa_ctrl[20].r.part0[10] 
	,\sa_ctrl[20].r.part0[9] ,\sa_ctrl[20].r.part0[8] 
	,\sa_ctrl[20].r.part0[7] ,\sa_ctrl[20].r.part0[6] 
	,\sa_ctrl[20].r.part0[5] ,\sa_ctrl[20].r.part0[4] 
	,\sa_ctrl[20].r.part0[3] ,\sa_ctrl[20].r.part0[2] 
	,\sa_ctrl[20].r.part0[1] ,\sa_ctrl[20].r.part0[0] 
	,\sa_ctrl[19].r.part0[31] ,\sa_ctrl[19].r.part0[30] 
	,\sa_ctrl[19].r.part0[29] ,\sa_ctrl[19].r.part0[28] 
	,\sa_ctrl[19].r.part0[27] ,\sa_ctrl[19].r.part0[26] 
	,\sa_ctrl[19].r.part0[25] ,\sa_ctrl[19].r.part0[24] 
	,\sa_ctrl[19].r.part0[23] ,\sa_ctrl[19].r.part0[22] 
	,\sa_ctrl[19].r.part0[21] ,\sa_ctrl[19].r.part0[20] 
	,\sa_ctrl[19].r.part0[19] ,\sa_ctrl[19].r.part0[18] 
	,\sa_ctrl[19].r.part0[17] ,\sa_ctrl[19].r.part0[16] 
	,\sa_ctrl[19].r.part0[15] ,\sa_ctrl[19].r.part0[14] 
	,\sa_ctrl[19].r.part0[13] ,\sa_ctrl[19].r.part0[12] 
	,\sa_ctrl[19].r.part0[11] ,\sa_ctrl[19].r.part0[10] 
	,\sa_ctrl[19].r.part0[9] ,\sa_ctrl[19].r.part0[8] 
	,\sa_ctrl[19].r.part0[7] ,\sa_ctrl[19].r.part0[6] 
	,\sa_ctrl[19].r.part0[5] ,\sa_ctrl[19].r.part0[4] 
	,\sa_ctrl[19].r.part0[3] ,\sa_ctrl[19].r.part0[2] 
	,\sa_ctrl[19].r.part0[1] ,\sa_ctrl[19].r.part0[0] 
	,\sa_ctrl[18].r.part0[31] ,\sa_ctrl[18].r.part0[30] 
	,\sa_ctrl[18].r.part0[29] ,\sa_ctrl[18].r.part0[28] 
	,\sa_ctrl[18].r.part0[27] ,\sa_ctrl[18].r.part0[26] 
	,\sa_ctrl[18].r.part0[25] ,\sa_ctrl[18].r.part0[24] 
	,\sa_ctrl[18].r.part0[23] ,\sa_ctrl[18].r.part0[22] 
	,\sa_ctrl[18].r.part0[21] ,\sa_ctrl[18].r.part0[20] 
	,\sa_ctrl[18].r.part0[19] ,\sa_ctrl[18].r.part0[18] 
	,\sa_ctrl[18].r.part0[17] ,\sa_ctrl[18].r.part0[16] 
	,\sa_ctrl[18].r.part0[15] ,\sa_ctrl[18].r.part0[14] 
	,\sa_ctrl[18].r.part0[13] ,\sa_ctrl[18].r.part0[12] 
	,\sa_ctrl[18].r.part0[11] ,\sa_ctrl[18].r.part0[10] 
	,\sa_ctrl[18].r.part0[9] ,\sa_ctrl[18].r.part0[8] 
	,\sa_ctrl[18].r.part0[7] ,\sa_ctrl[18].r.part0[6] 
	,\sa_ctrl[18].r.part0[5] ,\sa_ctrl[18].r.part0[4] 
	,\sa_ctrl[18].r.part0[3] ,\sa_ctrl[18].r.part0[2] 
	,\sa_ctrl[18].r.part0[1] ,\sa_ctrl[18].r.part0[0] 
	,\sa_ctrl[17].r.part0[31] ,\sa_ctrl[17].r.part0[30] 
	,\sa_ctrl[17].r.part0[29] ,\sa_ctrl[17].r.part0[28] 
	,\sa_ctrl[17].r.part0[27] ,\sa_ctrl[17].r.part0[26] 
	,\sa_ctrl[17].r.part0[25] ,\sa_ctrl[17].r.part0[24] 
	,\sa_ctrl[17].r.part0[23] ,\sa_ctrl[17].r.part0[22] 
	,\sa_ctrl[17].r.part0[21] ,\sa_ctrl[17].r.part0[20] 
	,\sa_ctrl[17].r.part0[19] ,\sa_ctrl[17].r.part0[18] 
	,\sa_ctrl[17].r.part0[17] ,\sa_ctrl[17].r.part0[16] 
	,\sa_ctrl[17].r.part0[15] ,\sa_ctrl[17].r.part0[14] 
	,\sa_ctrl[17].r.part0[13] ,\sa_ctrl[17].r.part0[12] 
	,\sa_ctrl[17].r.part0[11] ,\sa_ctrl[17].r.part0[10] 
	,\sa_ctrl[17].r.part0[9] ,\sa_ctrl[17].r.part0[8] 
	,\sa_ctrl[17].r.part0[7] ,\sa_ctrl[17].r.part0[6] 
	,\sa_ctrl[17].r.part0[5] ,\sa_ctrl[17].r.part0[4] 
	,\sa_ctrl[17].r.part0[3] ,\sa_ctrl[17].r.part0[2] 
	,\sa_ctrl[17].r.part0[1] ,\sa_ctrl[17].r.part0[0] 
	,\sa_ctrl[16].r.part0[31] ,\sa_ctrl[16].r.part0[30] 
	,\sa_ctrl[16].r.part0[29] ,\sa_ctrl[16].r.part0[28] 
	,\sa_ctrl[16].r.part0[27] ,\sa_ctrl[16].r.part0[26] 
	,\sa_ctrl[16].r.part0[25] ,\sa_ctrl[16].r.part0[24] 
	,\sa_ctrl[16].r.part0[23] ,\sa_ctrl[16].r.part0[22] 
	,\sa_ctrl[16].r.part0[21] ,\sa_ctrl[16].r.part0[20] 
	,\sa_ctrl[16].r.part0[19] ,\sa_ctrl[16].r.part0[18] 
	,\sa_ctrl[16].r.part0[17] ,\sa_ctrl[16].r.part0[16] 
	,\sa_ctrl[16].r.part0[15] ,\sa_ctrl[16].r.part0[14] 
	,\sa_ctrl[16].r.part0[13] ,\sa_ctrl[16].r.part0[12] 
	,\sa_ctrl[16].r.part0[11] ,\sa_ctrl[16].r.part0[10] 
	,\sa_ctrl[16].r.part0[9] ,\sa_ctrl[16].r.part0[8] 
	,\sa_ctrl[16].r.part0[7] ,\sa_ctrl[16].r.part0[6] 
	,\sa_ctrl[16].r.part0[5] ,\sa_ctrl[16].r.part0[4] 
	,\sa_ctrl[16].r.part0[3] ,\sa_ctrl[16].r.part0[2] 
	,\sa_ctrl[16].r.part0[1] ,\sa_ctrl[16].r.part0[0] 
	,\sa_ctrl[15].r.part0[31] ,\sa_ctrl[15].r.part0[30] 
	,\sa_ctrl[15].r.part0[29] ,\sa_ctrl[15].r.part0[28] 
	,\sa_ctrl[15].r.part0[27] ,\sa_ctrl[15].r.part0[26] 
	,\sa_ctrl[15].r.part0[25] ,\sa_ctrl[15].r.part0[24] 
	,\sa_ctrl[15].r.part0[23] ,\sa_ctrl[15].r.part0[22] 
	,\sa_ctrl[15].r.part0[21] ,\sa_ctrl[15].r.part0[20] 
	,\sa_ctrl[15].r.part0[19] ,\sa_ctrl[15].r.part0[18] 
	,\sa_ctrl[15].r.part0[17] ,\sa_ctrl[15].r.part0[16] 
	,\sa_ctrl[15].r.part0[15] ,\sa_ctrl[15].r.part0[14] 
	,\sa_ctrl[15].r.part0[13] ,\sa_ctrl[15].r.part0[12] 
	,\sa_ctrl[15].r.part0[11] ,\sa_ctrl[15].r.part0[10] 
	,\sa_ctrl[15].r.part0[9] ,\sa_ctrl[15].r.part0[8] 
	,\sa_ctrl[15].r.part0[7] ,\sa_ctrl[15].r.part0[6] 
	,\sa_ctrl[15].r.part0[5] ,\sa_ctrl[15].r.part0[4] 
	,\sa_ctrl[15].r.part0[3] ,\sa_ctrl[15].r.part0[2] 
	,\sa_ctrl[15].r.part0[1] ,\sa_ctrl[15].r.part0[0] 
	,\sa_ctrl[14].r.part0[31] ,\sa_ctrl[14].r.part0[30] 
	,\sa_ctrl[14].r.part0[29] ,\sa_ctrl[14].r.part0[28] 
	,\sa_ctrl[14].r.part0[27] ,\sa_ctrl[14].r.part0[26] 
	,\sa_ctrl[14].r.part0[25] ,\sa_ctrl[14].r.part0[24] 
	,\sa_ctrl[14].r.part0[23] ,\sa_ctrl[14].r.part0[22] 
	,\sa_ctrl[14].r.part0[21] ,\sa_ctrl[14].r.part0[20] 
	,\sa_ctrl[14].r.part0[19] ,\sa_ctrl[14].r.part0[18] 
	,\sa_ctrl[14].r.part0[17] ,\sa_ctrl[14].r.part0[16] 
	,\sa_ctrl[14].r.part0[15] ,\sa_ctrl[14].r.part0[14] 
	,\sa_ctrl[14].r.part0[13] ,\sa_ctrl[14].r.part0[12] 
	,\sa_ctrl[14].r.part0[11] ,\sa_ctrl[14].r.part0[10] 
	,\sa_ctrl[14].r.part0[9] ,\sa_ctrl[14].r.part0[8] 
	,\sa_ctrl[14].r.part0[7] ,\sa_ctrl[14].r.part0[6] 
	,\sa_ctrl[14].r.part0[5] ,\sa_ctrl[14].r.part0[4] 
	,\sa_ctrl[14].r.part0[3] ,\sa_ctrl[14].r.part0[2] 
	,\sa_ctrl[14].r.part0[1] ,\sa_ctrl[14].r.part0[0] 
	,\sa_ctrl[13].r.part0[31] ,\sa_ctrl[13].r.part0[30] 
	,\sa_ctrl[13].r.part0[29] ,\sa_ctrl[13].r.part0[28] 
	,\sa_ctrl[13].r.part0[27] ,\sa_ctrl[13].r.part0[26] 
	,\sa_ctrl[13].r.part0[25] ,\sa_ctrl[13].r.part0[24] 
	,\sa_ctrl[13].r.part0[23] ,\sa_ctrl[13].r.part0[22] 
	,\sa_ctrl[13].r.part0[21] ,\sa_ctrl[13].r.part0[20] 
	,\sa_ctrl[13].r.part0[19] ,\sa_ctrl[13].r.part0[18] 
	,\sa_ctrl[13].r.part0[17] ,\sa_ctrl[13].r.part0[16] 
	,\sa_ctrl[13].r.part0[15] ,\sa_ctrl[13].r.part0[14] 
	,\sa_ctrl[13].r.part0[13] ,\sa_ctrl[13].r.part0[12] 
	,\sa_ctrl[13].r.part0[11] ,\sa_ctrl[13].r.part0[10] 
	,\sa_ctrl[13].r.part0[9] ,\sa_ctrl[13].r.part0[8] 
	,\sa_ctrl[13].r.part0[7] ,\sa_ctrl[13].r.part0[6] 
	,\sa_ctrl[13].r.part0[5] ,\sa_ctrl[13].r.part0[4] 
	,\sa_ctrl[13].r.part0[3] ,\sa_ctrl[13].r.part0[2] 
	,\sa_ctrl[13].r.part0[1] ,\sa_ctrl[13].r.part0[0] 
	,\sa_ctrl[12].r.part0[31] ,\sa_ctrl[12].r.part0[30] 
	,\sa_ctrl[12].r.part0[29] ,\sa_ctrl[12].r.part0[28] 
	,\sa_ctrl[12].r.part0[27] ,\sa_ctrl[12].r.part0[26] 
	,\sa_ctrl[12].r.part0[25] ,\sa_ctrl[12].r.part0[24] 
	,\sa_ctrl[12].r.part0[23] ,\sa_ctrl[12].r.part0[22] 
	,\sa_ctrl[12].r.part0[21] ,\sa_ctrl[12].r.part0[20] 
	,\sa_ctrl[12].r.part0[19] ,\sa_ctrl[12].r.part0[18] 
	,\sa_ctrl[12].r.part0[17] ,\sa_ctrl[12].r.part0[16] 
	,\sa_ctrl[12].r.part0[15] ,\sa_ctrl[12].r.part0[14] 
	,\sa_ctrl[12].r.part0[13] ,\sa_ctrl[12].r.part0[12] 
	,\sa_ctrl[12].r.part0[11] ,\sa_ctrl[12].r.part0[10] 
	,\sa_ctrl[12].r.part0[9] ,\sa_ctrl[12].r.part0[8] 
	,\sa_ctrl[12].r.part0[7] ,\sa_ctrl[12].r.part0[6] 
	,\sa_ctrl[12].r.part0[5] ,\sa_ctrl[12].r.part0[4] 
	,\sa_ctrl[12].r.part0[3] ,\sa_ctrl[12].r.part0[2] 
	,\sa_ctrl[12].r.part0[1] ,\sa_ctrl[12].r.part0[0] 
	,\sa_ctrl[11].r.part0[31] ,\sa_ctrl[11].r.part0[30] 
	,\sa_ctrl[11].r.part0[29] ,\sa_ctrl[11].r.part0[28] 
	,\sa_ctrl[11].r.part0[27] ,\sa_ctrl[11].r.part0[26] 
	,\sa_ctrl[11].r.part0[25] ,\sa_ctrl[11].r.part0[24] 
	,\sa_ctrl[11].r.part0[23] ,\sa_ctrl[11].r.part0[22] 
	,\sa_ctrl[11].r.part0[21] ,\sa_ctrl[11].r.part0[20] 
	,\sa_ctrl[11].r.part0[19] ,\sa_ctrl[11].r.part0[18] 
	,\sa_ctrl[11].r.part0[17] ,\sa_ctrl[11].r.part0[16] 
	,\sa_ctrl[11].r.part0[15] ,\sa_ctrl[11].r.part0[14] 
	,\sa_ctrl[11].r.part0[13] ,\sa_ctrl[11].r.part0[12] 
	,\sa_ctrl[11].r.part0[11] ,\sa_ctrl[11].r.part0[10] 
	,\sa_ctrl[11].r.part0[9] ,\sa_ctrl[11].r.part0[8] 
	,\sa_ctrl[11].r.part0[7] ,\sa_ctrl[11].r.part0[6] 
	,\sa_ctrl[11].r.part0[5] ,\sa_ctrl[11].r.part0[4] 
	,\sa_ctrl[11].r.part0[3] ,\sa_ctrl[11].r.part0[2] 
	,\sa_ctrl[11].r.part0[1] ,\sa_ctrl[11].r.part0[0] 
	,\sa_ctrl[10].r.part0[31] ,\sa_ctrl[10].r.part0[30] 
	,\sa_ctrl[10].r.part0[29] ,\sa_ctrl[10].r.part0[28] 
	,\sa_ctrl[10].r.part0[27] ,\sa_ctrl[10].r.part0[26] 
	,\sa_ctrl[10].r.part0[25] ,\sa_ctrl[10].r.part0[24] 
	,\sa_ctrl[10].r.part0[23] ,\sa_ctrl[10].r.part0[22] 
	,\sa_ctrl[10].r.part0[21] ,\sa_ctrl[10].r.part0[20] 
	,\sa_ctrl[10].r.part0[19] ,\sa_ctrl[10].r.part0[18] 
	,\sa_ctrl[10].r.part0[17] ,\sa_ctrl[10].r.part0[16] 
	,\sa_ctrl[10].r.part0[15] ,\sa_ctrl[10].r.part0[14] 
	,\sa_ctrl[10].r.part0[13] ,\sa_ctrl[10].r.part0[12] 
	,\sa_ctrl[10].r.part0[11] ,\sa_ctrl[10].r.part0[10] 
	,\sa_ctrl[10].r.part0[9] ,\sa_ctrl[10].r.part0[8] 
	,\sa_ctrl[10].r.part0[7] ,\sa_ctrl[10].r.part0[6] 
	,\sa_ctrl[10].r.part0[5] ,\sa_ctrl[10].r.part0[4] 
	,\sa_ctrl[10].r.part0[3] ,\sa_ctrl[10].r.part0[2] 
	,\sa_ctrl[10].r.part0[1] ,\sa_ctrl[10].r.part0[0] 
	,\sa_ctrl[9].r.part0[31] ,\sa_ctrl[9].r.part0[30] 
	,\sa_ctrl[9].r.part0[29] ,\sa_ctrl[9].r.part0[28] 
	,\sa_ctrl[9].r.part0[27] ,\sa_ctrl[9].r.part0[26] 
	,\sa_ctrl[9].r.part0[25] ,\sa_ctrl[9].r.part0[24] 
	,\sa_ctrl[9].r.part0[23] ,\sa_ctrl[9].r.part0[22] 
	,\sa_ctrl[9].r.part0[21] ,\sa_ctrl[9].r.part0[20] 
	,\sa_ctrl[9].r.part0[19] ,\sa_ctrl[9].r.part0[18] 
	,\sa_ctrl[9].r.part0[17] ,\sa_ctrl[9].r.part0[16] 
	,\sa_ctrl[9].r.part0[15] ,\sa_ctrl[9].r.part0[14] 
	,\sa_ctrl[9].r.part0[13] ,\sa_ctrl[9].r.part0[12] 
	,\sa_ctrl[9].r.part0[11] ,\sa_ctrl[9].r.part0[10] 
	,\sa_ctrl[9].r.part0[9] ,\sa_ctrl[9].r.part0[8] 
	,\sa_ctrl[9].r.part0[7] ,\sa_ctrl[9].r.part0[6] 
	,\sa_ctrl[9].r.part0[5] ,\sa_ctrl[9].r.part0[4] 
	,\sa_ctrl[9].r.part0[3] ,\sa_ctrl[9].r.part0[2] 
	,\sa_ctrl[9].r.part0[1] ,\sa_ctrl[9].r.part0[0] 
	,\sa_ctrl[8].r.part0[31] ,\sa_ctrl[8].r.part0[30] 
	,\sa_ctrl[8].r.part0[29] ,\sa_ctrl[8].r.part0[28] 
	,\sa_ctrl[8].r.part0[27] ,\sa_ctrl[8].r.part0[26] 
	,\sa_ctrl[8].r.part0[25] ,\sa_ctrl[8].r.part0[24] 
	,\sa_ctrl[8].r.part0[23] ,\sa_ctrl[8].r.part0[22] 
	,\sa_ctrl[8].r.part0[21] ,\sa_ctrl[8].r.part0[20] 
	,\sa_ctrl[8].r.part0[19] ,\sa_ctrl[8].r.part0[18] 
	,\sa_ctrl[8].r.part0[17] ,\sa_ctrl[8].r.part0[16] 
	,\sa_ctrl[8].r.part0[15] ,\sa_ctrl[8].r.part0[14] 
	,\sa_ctrl[8].r.part0[13] ,\sa_ctrl[8].r.part0[12] 
	,\sa_ctrl[8].r.part0[11] ,\sa_ctrl[8].r.part0[10] 
	,\sa_ctrl[8].r.part0[9] ,\sa_ctrl[8].r.part0[8] 
	,\sa_ctrl[8].r.part0[7] ,\sa_ctrl[8].r.part0[6] 
	,\sa_ctrl[8].r.part0[5] ,\sa_ctrl[8].r.part0[4] 
	,\sa_ctrl[8].r.part0[3] ,\sa_ctrl[8].r.part0[2] 
	,\sa_ctrl[8].r.part0[1] ,\sa_ctrl[8].r.part0[0] 
	,\sa_ctrl[7].r.part0[31] ,\sa_ctrl[7].r.part0[30] 
	,\sa_ctrl[7].r.part0[29] ,\sa_ctrl[7].r.part0[28] 
	,\sa_ctrl[7].r.part0[27] ,\sa_ctrl[7].r.part0[26] 
	,\sa_ctrl[7].r.part0[25] ,\sa_ctrl[7].r.part0[24] 
	,\sa_ctrl[7].r.part0[23] ,\sa_ctrl[7].r.part0[22] 
	,\sa_ctrl[7].r.part0[21] ,\sa_ctrl[7].r.part0[20] 
	,\sa_ctrl[7].r.part0[19] ,\sa_ctrl[7].r.part0[18] 
	,\sa_ctrl[7].r.part0[17] ,\sa_ctrl[7].r.part0[16] 
	,\sa_ctrl[7].r.part0[15] ,\sa_ctrl[7].r.part0[14] 
	,\sa_ctrl[7].r.part0[13] ,\sa_ctrl[7].r.part0[12] 
	,\sa_ctrl[7].r.part0[11] ,\sa_ctrl[7].r.part0[10] 
	,\sa_ctrl[7].r.part0[9] ,\sa_ctrl[7].r.part0[8] 
	,\sa_ctrl[7].r.part0[7] ,\sa_ctrl[7].r.part0[6] 
	,\sa_ctrl[7].r.part0[5] ,\sa_ctrl[7].r.part0[4] 
	,\sa_ctrl[7].r.part0[3] ,\sa_ctrl[7].r.part0[2] 
	,\sa_ctrl[7].r.part0[1] ,\sa_ctrl[7].r.part0[0] 
	,\sa_ctrl[6].r.part0[31] ,\sa_ctrl[6].r.part0[30] 
	,\sa_ctrl[6].r.part0[29] ,\sa_ctrl[6].r.part0[28] 
	,\sa_ctrl[6].r.part0[27] ,\sa_ctrl[6].r.part0[26] 
	,\sa_ctrl[6].r.part0[25] ,\sa_ctrl[6].r.part0[24] 
	,\sa_ctrl[6].r.part0[23] ,\sa_ctrl[6].r.part0[22] 
	,\sa_ctrl[6].r.part0[21] ,\sa_ctrl[6].r.part0[20] 
	,\sa_ctrl[6].r.part0[19] ,\sa_ctrl[6].r.part0[18] 
	,\sa_ctrl[6].r.part0[17] ,\sa_ctrl[6].r.part0[16] 
	,\sa_ctrl[6].r.part0[15] ,\sa_ctrl[6].r.part0[14] 
	,\sa_ctrl[6].r.part0[13] ,\sa_ctrl[6].r.part0[12] 
	,\sa_ctrl[6].r.part0[11] ,\sa_ctrl[6].r.part0[10] 
	,\sa_ctrl[6].r.part0[9] ,\sa_ctrl[6].r.part0[8] 
	,\sa_ctrl[6].r.part0[7] ,\sa_ctrl[6].r.part0[6] 
	,\sa_ctrl[6].r.part0[5] ,\sa_ctrl[6].r.part0[4] 
	,\sa_ctrl[6].r.part0[3] ,\sa_ctrl[6].r.part0[2] 
	,\sa_ctrl[6].r.part0[1] ,\sa_ctrl[6].r.part0[0] 
	,\sa_ctrl[5].r.part0[31] ,\sa_ctrl[5].r.part0[30] 
	,\sa_ctrl[5].r.part0[29] ,\sa_ctrl[5].r.part0[28] 
	,\sa_ctrl[5].r.part0[27] ,\sa_ctrl[5].r.part0[26] 
	,\sa_ctrl[5].r.part0[25] ,\sa_ctrl[5].r.part0[24] 
	,\sa_ctrl[5].r.part0[23] ,\sa_ctrl[5].r.part0[22] 
	,\sa_ctrl[5].r.part0[21] ,\sa_ctrl[5].r.part0[20] 
	,\sa_ctrl[5].r.part0[19] ,\sa_ctrl[5].r.part0[18] 
	,\sa_ctrl[5].r.part0[17] ,\sa_ctrl[5].r.part0[16] 
	,\sa_ctrl[5].r.part0[15] ,\sa_ctrl[5].r.part0[14] 
	,\sa_ctrl[5].r.part0[13] ,\sa_ctrl[5].r.part0[12] 
	,\sa_ctrl[5].r.part0[11] ,\sa_ctrl[5].r.part0[10] 
	,\sa_ctrl[5].r.part0[9] ,\sa_ctrl[5].r.part0[8] 
	,\sa_ctrl[5].r.part0[7] ,\sa_ctrl[5].r.part0[6] 
	,\sa_ctrl[5].r.part0[5] ,\sa_ctrl[5].r.part0[4] 
	,\sa_ctrl[5].r.part0[3] ,\sa_ctrl[5].r.part0[2] 
	,\sa_ctrl[5].r.part0[1] ,\sa_ctrl[5].r.part0[0] 
	,\sa_ctrl[4].r.part0[31] ,\sa_ctrl[4].r.part0[30] 
	,\sa_ctrl[4].r.part0[29] ,\sa_ctrl[4].r.part0[28] 
	,\sa_ctrl[4].r.part0[27] ,\sa_ctrl[4].r.part0[26] 
	,\sa_ctrl[4].r.part0[25] ,\sa_ctrl[4].r.part0[24] 
	,\sa_ctrl[4].r.part0[23] ,\sa_ctrl[4].r.part0[22] 
	,\sa_ctrl[4].r.part0[21] ,\sa_ctrl[4].r.part0[20] 
	,\sa_ctrl[4].r.part0[19] ,\sa_ctrl[4].r.part0[18] 
	,\sa_ctrl[4].r.part0[17] ,\sa_ctrl[4].r.part0[16] 
	,\sa_ctrl[4].r.part0[15] ,\sa_ctrl[4].r.part0[14] 
	,\sa_ctrl[4].r.part0[13] ,\sa_ctrl[4].r.part0[12] 
	,\sa_ctrl[4].r.part0[11] ,\sa_ctrl[4].r.part0[10] 
	,\sa_ctrl[4].r.part0[9] ,\sa_ctrl[4].r.part0[8] 
	,\sa_ctrl[4].r.part0[7] ,\sa_ctrl[4].r.part0[6] 
	,\sa_ctrl[4].r.part0[5] ,\sa_ctrl[4].r.part0[4] 
	,\sa_ctrl[4].r.part0[3] ,\sa_ctrl[4].r.part0[2] 
	,\sa_ctrl[4].r.part0[1] ,\sa_ctrl[4].r.part0[0] 
	,\sa_ctrl[3].r.part0[31] ,\sa_ctrl[3].r.part0[30] 
	,\sa_ctrl[3].r.part0[29] ,\sa_ctrl[3].r.part0[28] 
	,\sa_ctrl[3].r.part0[27] ,\sa_ctrl[3].r.part0[26] 
	,\sa_ctrl[3].r.part0[25] ,\sa_ctrl[3].r.part0[24] 
	,\sa_ctrl[3].r.part0[23] ,\sa_ctrl[3].r.part0[22] 
	,\sa_ctrl[3].r.part0[21] ,\sa_ctrl[3].r.part0[20] 
	,\sa_ctrl[3].r.part0[19] ,\sa_ctrl[3].r.part0[18] 
	,\sa_ctrl[3].r.part0[17] ,\sa_ctrl[3].r.part0[16] 
	,\sa_ctrl[3].r.part0[15] ,\sa_ctrl[3].r.part0[14] 
	,\sa_ctrl[3].r.part0[13] ,\sa_ctrl[3].r.part0[12] 
	,\sa_ctrl[3].r.part0[11] ,\sa_ctrl[3].r.part0[10] 
	,\sa_ctrl[3].r.part0[9] ,\sa_ctrl[3].r.part0[8] 
	,\sa_ctrl[3].r.part0[7] ,\sa_ctrl[3].r.part0[6] 
	,\sa_ctrl[3].r.part0[5] ,\sa_ctrl[3].r.part0[4] 
	,\sa_ctrl[3].r.part0[3] ,\sa_ctrl[3].r.part0[2] 
	,\sa_ctrl[3].r.part0[1] ,\sa_ctrl[3].r.part0[0] 
	,\sa_ctrl[2].r.part0[31] ,\sa_ctrl[2].r.part0[30] 
	,\sa_ctrl[2].r.part0[29] ,\sa_ctrl[2].r.part0[28] 
	,\sa_ctrl[2].r.part0[27] ,\sa_ctrl[2].r.part0[26] 
	,\sa_ctrl[2].r.part0[25] ,\sa_ctrl[2].r.part0[24] 
	,\sa_ctrl[2].r.part0[23] ,\sa_ctrl[2].r.part0[22] 
	,\sa_ctrl[2].r.part0[21] ,\sa_ctrl[2].r.part0[20] 
	,\sa_ctrl[2].r.part0[19] ,\sa_ctrl[2].r.part0[18] 
	,\sa_ctrl[2].r.part0[17] ,\sa_ctrl[2].r.part0[16] 
	,\sa_ctrl[2].r.part0[15] ,\sa_ctrl[2].r.part0[14] 
	,\sa_ctrl[2].r.part0[13] ,\sa_ctrl[2].r.part0[12] 
	,\sa_ctrl[2].r.part0[11] ,\sa_ctrl[2].r.part0[10] 
	,\sa_ctrl[2].r.part0[9] ,\sa_ctrl[2].r.part0[8] 
	,\sa_ctrl[2].r.part0[7] ,\sa_ctrl[2].r.part0[6] 
	,\sa_ctrl[2].r.part0[5] ,\sa_ctrl[2].r.part0[4] 
	,\sa_ctrl[2].r.part0[3] ,\sa_ctrl[2].r.part0[2] 
	,\sa_ctrl[2].r.part0[1] ,\sa_ctrl[2].r.part0[0] 
	,\sa_ctrl[1].r.part0[31] ,\sa_ctrl[1].r.part0[30] 
	,\sa_ctrl[1].r.part0[29] ,\sa_ctrl[1].r.part0[28] 
	,\sa_ctrl[1].r.part0[27] ,\sa_ctrl[1].r.part0[26] 
	,\sa_ctrl[1].r.part0[25] ,\sa_ctrl[1].r.part0[24] 
	,\sa_ctrl[1].r.part0[23] ,\sa_ctrl[1].r.part0[22] 
	,\sa_ctrl[1].r.part0[21] ,\sa_ctrl[1].r.part0[20] 
	,\sa_ctrl[1].r.part0[19] ,\sa_ctrl[1].r.part0[18] 
	,\sa_ctrl[1].r.part0[17] ,\sa_ctrl[1].r.part0[16] 
	,\sa_ctrl[1].r.part0[15] ,\sa_ctrl[1].r.part0[14] 
	,\sa_ctrl[1].r.part0[13] ,\sa_ctrl[1].r.part0[12] 
	,\sa_ctrl[1].r.part0[11] ,\sa_ctrl[1].r.part0[10] 
	,\sa_ctrl[1].r.part0[9] ,\sa_ctrl[1].r.part0[8] 
	,\sa_ctrl[1].r.part0[7] ,\sa_ctrl[1].r.part0[6] 
	,\sa_ctrl[1].r.part0[5] ,\sa_ctrl[1].r.part0[4] 
	,\sa_ctrl[1].r.part0[3] ,\sa_ctrl[1].r.part0[2] 
	,\sa_ctrl[1].r.part0[1] ,\sa_ctrl[1].r.part0[0] 
	,\sa_ctrl[0].r.part0[31] ,\sa_ctrl[0].r.part0[30] 
	,\sa_ctrl[0].r.part0[29] ,\sa_ctrl[0].r.part0[28] 
	,\sa_ctrl[0].r.part0[27] ,\sa_ctrl[0].r.part0[26] 
	,\sa_ctrl[0].r.part0[25] ,\sa_ctrl[0].r.part0[24] 
	,\sa_ctrl[0].r.part0[23] ,\sa_ctrl[0].r.part0[22] 
	,\sa_ctrl[0].r.part0[21] ,\sa_ctrl[0].r.part0[20] 
	,\sa_ctrl[0].r.part0[19] ,\sa_ctrl[0].r.part0[18] 
	,\sa_ctrl[0].r.part0[17] ,\sa_ctrl[0].r.part0[16] 
	,\sa_ctrl[0].r.part0[15] ,\sa_ctrl[0].r.part0[14] 
	,\sa_ctrl[0].r.part0[13] ,\sa_ctrl[0].r.part0[12] 
	,\sa_ctrl[0].r.part0[11] ,\sa_ctrl[0].r.part0[10] 
	,\sa_ctrl[0].r.part0[9] ,\sa_ctrl[0].r.part0[8] 
	,\sa_ctrl[0].r.part0[7] ,\sa_ctrl[0].r.part0[6] 
	,\sa_ctrl[0].r.part0[5] ,\sa_ctrl[0].r.part0[4] 
	,\sa_ctrl[0].r.part0[3] ,\sa_ctrl[0].r.part0[2] 
	,\sa_ctrl[0].r.part0[1] ,\sa_ctrl[0].r.part0[0] ;
input stat_drbg_reseed;
input stat_req_with_expired_seed;
input stat_aux_key_type_0;
input stat_aux_key_type_1;
input stat_aux_key_type_2;
input stat_aux_key_type_3;
input stat_aux_key_type_4;
input stat_aux_key_type_5;
input stat_aux_key_type_6;
input stat_aux_key_type_7;
input stat_aux_key_type_8;
input stat_aux_key_type_9;
input stat_aux_key_type_10;
input stat_aux_key_type_11;
input stat_aux_key_type_12;
input stat_aux_key_type_13;
input stat_cceip0_stall_on_valid_key;
input stat_cceip1_stall_on_valid_key;
input stat_cceip2_stall_on_valid_key;
input stat_cceip3_stall_on_valid_key;
input stat_cddip0_stall_on_valid_key;
input stat_cddip1_stall_on_valid_key;
input stat_cddip2_stall_on_valid_key;
input stat_cddip3_stall_on_valid_key;
input stat_aux_cmd_with_vf_pf_fail;
input kme_slv_empty;
input drng_idle;
input tlv_parser_idle;
input tlv_parser_int_tlv_start_pulse;
input [3:0] cceip_key_tlv_rsm_end_pulse;
input [3:0] cddip_key_tlv_rsm_end_pulse;
input [3:0] cceip_key_tlv_rsm_idle;
input [3:0] cddip_key_tlv_rsm_idle;
wire _zy_simnet_disable_debug_cmd_q_0_w$;
wire _zy_simnet_set_txc_bp_int_1_w$;
wire _zy_simnet_kme_ib_out_2_w$;
wire _zy_simnet_kme_idle_3_w$;
wire [0:31] _zy_simnet_idle_components_4_w$;
wire [31:0] k;
wire [31:0] num_key_tlv_in_flight;
wire sa_snap;
wire sa_clear;
wire regs_sa_snap_r;
wire regs_sa_clear_live_r;
wire [0:9] \num_0_._zy_simnet_tvar_7 ;
wire \num_0_._zy_simnet_sa_clear_8_w$ ;
wire \num_0_._zy_simnet_sa_snap_9_w$ ;
wire [0:49] \num_0_._zy_simnet_tvar_6 ;
wire [0:49] \num_0_._zy_simnet_tvar_5 ;
wire [0:9] \num_1_._zy_simnet_tvar_12 ;
wire \num_1_._zy_simnet_sa_clear_13_w$ ;
wire \num_1_._zy_simnet_sa_snap_14_w$ ;
wire [0:49] \num_1_._zy_simnet_tvar_11 ;
wire [0:49] \num_1_._zy_simnet_tvar_10 ;
wire [0:9] \num_2_._zy_simnet_tvar_17 ;
wire \num_2_._zy_simnet_sa_clear_18_w$ ;
wire \num_2_._zy_simnet_sa_snap_19_w$ ;
wire [0:49] \num_2_._zy_simnet_tvar_16 ;
wire [0:49] \num_2_._zy_simnet_tvar_15 ;
wire [0:9] \num_3_._zy_simnet_tvar_22 ;
wire \num_3_._zy_simnet_sa_clear_23_w$ ;
wire \num_3_._zy_simnet_sa_snap_24_w$ ;
wire [0:49] \num_3_._zy_simnet_tvar_21 ;
wire [0:49] \num_3_._zy_simnet_tvar_20 ;
wire [0:9] \num_4_._zy_simnet_tvar_27 ;
wire \num_4_._zy_simnet_sa_clear_28_w$ ;
wire \num_4_._zy_simnet_sa_snap_29_w$ ;
wire [0:49] \num_4_._zy_simnet_tvar_26 ;
wire [0:49] \num_4_._zy_simnet_tvar_25 ;
wire [0:9] \num_5_._zy_simnet_tvar_32 ;
wire \num_5_._zy_simnet_sa_clear_33_w$ ;
wire \num_5_._zy_simnet_sa_snap_34_w$ ;
wire [0:49] \num_5_._zy_simnet_tvar_31 ;
wire [0:49] \num_5_._zy_simnet_tvar_30 ;
wire [0:9] \num_6_._zy_simnet_tvar_37 ;
wire \num_6_._zy_simnet_sa_clear_38_w$ ;
wire \num_6_._zy_simnet_sa_snap_39_w$ ;
wire [0:49] \num_6_._zy_simnet_tvar_36 ;
wire [0:49] \num_6_._zy_simnet_tvar_35 ;
wire [0:9] \num_7_._zy_simnet_tvar_42 ;
wire \num_7_._zy_simnet_sa_clear_43_w$ ;
wire \num_7_._zy_simnet_sa_snap_44_w$ ;
wire [0:49] \num_7_._zy_simnet_tvar_41 ;
wire [0:49] \num_7_._zy_simnet_tvar_40 ;
wire [0:9] \num_8_._zy_simnet_tvar_47 ;
wire \num_8_._zy_simnet_sa_clear_48_w$ ;
wire \num_8_._zy_simnet_sa_snap_49_w$ ;
wire [0:49] \num_8_._zy_simnet_tvar_46 ;
wire [0:49] \num_8_._zy_simnet_tvar_45 ;
wire [0:9] \num_9_._zy_simnet_tvar_52 ;
wire \num_9_._zy_simnet_sa_clear_53_w$ ;
wire \num_9_._zy_simnet_sa_snap_54_w$ ;
wire [0:49] \num_9_._zy_simnet_tvar_51 ;
wire [0:49] \num_9_._zy_simnet_tvar_50 ;
wire [0:9] \num_10_._zy_simnet_tvar_57 ;
wire \num_10_._zy_simnet_sa_clear_58_w$ ;
wire \num_10_._zy_simnet_sa_snap_59_w$ ;
wire [0:49] \num_10_._zy_simnet_tvar_56 ;
wire [0:49] \num_10_._zy_simnet_tvar_55 ;
wire [0:9] \num_11_._zy_simnet_tvar_62 ;
wire \num_11_._zy_simnet_sa_clear_63_w$ ;
wire \num_11_._zy_simnet_sa_snap_64_w$ ;
wire [0:49] \num_11_._zy_simnet_tvar_61 ;
wire [0:49] \num_11_._zy_simnet_tvar_60 ;
wire [0:9] \num_12_._zy_simnet_tvar_67 ;
wire \num_12_._zy_simnet_sa_clear_68_w$ ;
wire \num_12_._zy_simnet_sa_snap_69_w$ ;
wire [0:49] \num_12_._zy_simnet_tvar_66 ;
wire [0:49] \num_12_._zy_simnet_tvar_65 ;
wire [0:9] \num_13_._zy_simnet_tvar_72 ;
wire \num_13_._zy_simnet_sa_clear_73_w$ ;
wire \num_13_._zy_simnet_sa_snap_74_w$ ;
wire [0:49] \num_13_._zy_simnet_tvar_71 ;
wire [0:49] \num_13_._zy_simnet_tvar_70 ;
wire [0:9] \num_14_._zy_simnet_tvar_77 ;
wire \num_14_._zy_simnet_sa_clear_78_w$ ;
wire \num_14_._zy_simnet_sa_snap_79_w$ ;
wire [0:49] \num_14_._zy_simnet_tvar_76 ;
wire [0:49] \num_14_._zy_simnet_tvar_75 ;
wire [0:9] \num_15_._zy_simnet_tvar_82 ;
wire \num_15_._zy_simnet_sa_clear_83_w$ ;
wire \num_15_._zy_simnet_sa_snap_84_w$ ;
wire [0:49] \num_15_._zy_simnet_tvar_81 ;
wire [0:49] \num_15_._zy_simnet_tvar_80 ;
wire [0:9] \num_16_._zy_simnet_tvar_87 ;
wire \num_16_._zy_simnet_sa_clear_88_w$ ;
wire \num_16_._zy_simnet_sa_snap_89_w$ ;
wire [0:49] \num_16_._zy_simnet_tvar_86 ;
wire [0:49] \num_16_._zy_simnet_tvar_85 ;
wire [0:9] \num_17_._zy_simnet_tvar_92 ;
wire \num_17_._zy_simnet_sa_clear_93_w$ ;
wire \num_17_._zy_simnet_sa_snap_94_w$ ;
wire [0:49] \num_17_._zy_simnet_tvar_91 ;
wire [0:49] \num_17_._zy_simnet_tvar_90 ;
wire [0:9] \num_18_._zy_simnet_tvar_97 ;
wire \num_18_._zy_simnet_sa_clear_98_w$ ;
wire \num_18_._zy_simnet_sa_snap_99_w$ ;
wire [0:49] \num_18_._zy_simnet_tvar_96 ;
wire [0:49] \num_18_._zy_simnet_tvar_95 ;
wire [0:9] \num_19_._zy_simnet_tvar_102 ;
wire \num_19_._zy_simnet_sa_clear_103_w$ ;
wire \num_19_._zy_simnet_sa_snap_104_w$ ;
wire [0:49] \num_19_._zy_simnet_tvar_101 ;
wire [0:49] \num_19_._zy_simnet_tvar_100 ;
wire [0:9] \num_20_._zy_simnet_tvar_107 ;
wire \num_20_._zy_simnet_sa_clear_108_w$ ;
wire \num_20_._zy_simnet_sa_snap_109_w$ ;
wire [0:49] \num_20_._zy_simnet_tvar_106 ;
wire [0:49] \num_20_._zy_simnet_tvar_105 ;
wire [0:9] \num_21_._zy_simnet_tvar_112 ;
wire \num_21_._zy_simnet_sa_clear_113_w$ ;
wire \num_21_._zy_simnet_sa_snap_114_w$ ;
wire [0:49] \num_21_._zy_simnet_tvar_111 ;
wire [0:49] \num_21_._zy_simnet_tvar_110 ;
wire [0:9] \num_22_._zy_simnet_tvar_117 ;
wire \num_22_._zy_simnet_sa_clear_118_w$ ;
wire \num_22_._zy_simnet_sa_snap_119_w$ ;
wire [0:49] \num_22_._zy_simnet_tvar_116 ;
wire [0:49] \num_22_._zy_simnet_tvar_115 ;
wire [0:9] \num_23_._zy_simnet_tvar_122 ;
wire \num_23_._zy_simnet_sa_clear_123_w$ ;
wire \num_23_._zy_simnet_sa_snap_124_w$ ;
wire [0:49] \num_23_._zy_simnet_tvar_121 ;
wire [0:49] \num_23_._zy_simnet_tvar_120 ;
wire [0:9] \num_24_._zy_simnet_tvar_127 ;
wire \num_24_._zy_simnet_sa_clear_128_w$ ;
wire \num_24_._zy_simnet_sa_snap_129_w$ ;
wire [0:49] \num_24_._zy_simnet_tvar_126 ;
wire [0:49] \num_24_._zy_simnet_tvar_125 ;
wire [0:9] \num_25_._zy_simnet_tvar_132 ;
wire \num_25_._zy_simnet_sa_clear_133_w$ ;
wire \num_25_._zy_simnet_sa_snap_134_w$ ;
wire [0:49] \num_25_._zy_simnet_tvar_131 ;
wire [0:49] \num_25_._zy_simnet_tvar_130 ;
wire [0:9] \num_26_._zy_simnet_tvar_137 ;
wire \num_26_._zy_simnet_sa_clear_138_w$ ;
wire \num_26_._zy_simnet_sa_snap_139_w$ ;
wire [0:49] \num_26_._zy_simnet_tvar_136 ;
wire [0:49] \num_26_._zy_simnet_tvar_135 ;
wire [0:9] \num_27_._zy_simnet_tvar_142 ;
wire \num_27_._zy_simnet_sa_clear_143_w$ ;
wire \num_27_._zy_simnet_sa_snap_144_w$ ;
wire [0:49] \num_27_._zy_simnet_tvar_141 ;
wire [0:49] \num_27_._zy_simnet_tvar_140 ;
wire [0:9] \num_28_._zy_simnet_tvar_147 ;
wire \num_28_._zy_simnet_sa_clear_148_w$ ;
wire \num_28_._zy_simnet_sa_snap_149_w$ ;
wire [0:49] \num_28_._zy_simnet_tvar_146 ;
wire [0:49] \num_28_._zy_simnet_tvar_145 ;
wire [0:9] \num_29_._zy_simnet_tvar_152 ;
wire \num_29_._zy_simnet_sa_clear_153_w$ ;
wire \num_29_._zy_simnet_sa_snap_154_w$ ;
wire [0:49] \num_29_._zy_simnet_tvar_151 ;
wire [0:49] \num_29_._zy_simnet_tvar_150 ;
wire [0:9] \num_30_._zy_simnet_tvar_157 ;
wire \num_30_._zy_simnet_sa_clear_158_w$ ;
wire \num_30_._zy_simnet_sa_snap_159_w$ ;
wire [0:49] \num_30_._zy_simnet_tvar_156 ;
wire [0:49] \num_30_._zy_simnet_tvar_155 ;
wire [0:9] \num_31_._zy_simnet_tvar_162 ;
wire \num_31_._zy_simnet_sa_clear_163_w$ ;
wire \num_31_._zy_simnet_sa_snap_164_w$ ;
wire [0:49] \num_31_._zy_simnet_tvar_161 ;
wire [0:49] \num_31_._zy_simnet_tvar_160 ;
supply0 n1;
supply0 n81;
supply0 n82;
supply0 n83;
supply0 n84;
supply0 n85;
supply0 n86;
supply0 n87;
supply0 n88;
supply0 n89;
supply0 n90;
supply0 n91;
supply0 n92;
supply0 n93;
supply0 n94;
supply0 n95;
supply0 n96;
supply0 n97;
supply0 n98;
supply0 n99;
supply0 n100;
supply0 n101;
supply0 n102;
supply0 n103;
supply0 n104;
supply0 n105;
supply0 n106;
supply0 n107;
supply0 n108;
supply0 n109;
supply0 n110;
supply0 n111;
supply0 n112;
supply0 n113;
supply0 n114;
supply0 n115;
supply0 n116;
supply0 n117;
supply0 n118;
supply0 n119;
supply0 n120;
supply0 n121;
supply0 n122;
supply0 n123;
supply0 n124;
supply0 n125;
supply0 n126;
supply0 n127;
supply0 n128;
supply0 n129;
supply0 n130;
supply0 n131;
supply0 n132;
supply0 n133;
supply0 n134;
supply0 n135;
supply0 n136;
supply0 n137;
supply0 n138;
supply0 n139;
supply0 n140;
supply0 n141;
supply0 n142;
supply0 n143;
supply0 n144;
supply0 n145;
supply0 n146;
supply0 n147;
supply0 n148;
supply0 n149;
supply0 n150;
supply0 n151;
supply0 n152;
supply0 n153;
supply0 n154;
supply0 n155;
supply0 n156;
supply0 n157;
supply0 n158;
supply0 n159;
supply0 n160;
supply0 n161;
supply0 n162;
supply0 n163;
supply0 n164;
supply0 n165;
supply0 n166;
supply0 n167;
supply0 n168;
supply0 n169;
supply0 n170;
supply0 n171;
supply0 n172;
supply0 n173;
supply0 n174;
supply0 n175;
supply0 n176;
supply0 n177;
supply0 n178;
supply0 n179;
supply0 n180;
supply0 n181;
supply0 n182;
supply0 n183;
supply0 n184;
supply0 n185;
supply0 n186;
supply0 n187;
supply0 n188;
supply0 n189;
supply0 n190;
supply0 n191;
supply0 n192;
supply0 n193;
supply0 n194;
supply0 n195;
supply0 n196;
supply0 n197;
supply0 n198;
supply0 n199;
supply0 n200;
supply0 n201;
supply0 n202;
supply0 n203;
supply0 n204;
supply0 n205;
supply0 n206;
supply0 n207;
supply0 n208;
supply0 n209;
supply0 n210;
supply0 n211;
supply0 n212;
supply0 n213;
supply0 n214;
supply0 n215;
supply0 n216;
supply0 n217;
supply0 n218;
supply0 n219;
supply0 n220;
supply0 n221;
supply0 n222;
supply0 n223;
supply0 n224;
supply0 n225;
supply0 n226;
supply0 n227;
supply0 n228;
supply0 n229;
supply0 n230;
supply0 n231;
supply0 n232;
supply0 n233;
supply0 n234;
supply0 n235;
supply0 n236;
supply0 n237;
supply0 n238;
supply0 n239;
supply0 n240;
tran (kme_ib_out[0], \kme_ib_out.tready );
tran (\sa_snapshot[0][0] , \sa_snapshot[0].r.part0[0] );
tran (\sa_snapshot[0][0] , \sa_snapshot[0].f.lower[0] );
tran (\sa_snapshot[0][1] , \sa_snapshot[0].r.part0[1] );
tran (\sa_snapshot[0][1] , \sa_snapshot[0].f.lower[1] );
tran (\sa_snapshot[0][2] , \sa_snapshot[0].r.part0[2] );
tran (\sa_snapshot[0][2] , \sa_snapshot[0].f.lower[2] );
tran (\sa_snapshot[0][3] , \sa_snapshot[0].r.part0[3] );
tran (\sa_snapshot[0][3] , \sa_snapshot[0].f.lower[3] );
tran (\sa_snapshot[0][4] , \sa_snapshot[0].r.part0[4] );
tran (\sa_snapshot[0][4] , \sa_snapshot[0].f.lower[4] );
tran (\sa_snapshot[0][5] , \sa_snapshot[0].r.part0[5] );
tran (\sa_snapshot[0][5] , \sa_snapshot[0].f.lower[5] );
tran (\sa_snapshot[0][6] , \sa_snapshot[0].r.part0[6] );
tran (\sa_snapshot[0][6] , \sa_snapshot[0].f.lower[6] );
tran (\sa_snapshot[0][7] , \sa_snapshot[0].r.part0[7] );
tran (\sa_snapshot[0][7] , \sa_snapshot[0].f.lower[7] );
tran (\sa_snapshot[0][8] , \sa_snapshot[0].r.part0[8] );
tran (\sa_snapshot[0][8] , \sa_snapshot[0].f.lower[8] );
tran (\sa_snapshot[0][9] , \sa_snapshot[0].r.part0[9] );
tran (\sa_snapshot[0][9] , \sa_snapshot[0].f.lower[9] );
tran (\sa_snapshot[0][10] , \sa_snapshot[0].r.part0[10] );
tran (\sa_snapshot[0][10] , \sa_snapshot[0].f.lower[10] );
tran (\sa_snapshot[0][11] , \sa_snapshot[0].r.part0[11] );
tran (\sa_snapshot[0][11] , \sa_snapshot[0].f.lower[11] );
tran (\sa_snapshot[0][12] , \sa_snapshot[0].r.part0[12] );
tran (\sa_snapshot[0][12] , \sa_snapshot[0].f.lower[12] );
tran (\sa_snapshot[0][13] , \sa_snapshot[0].r.part0[13] );
tran (\sa_snapshot[0][13] , \sa_snapshot[0].f.lower[13] );
tran (\sa_snapshot[0][14] , \sa_snapshot[0].r.part0[14] );
tran (\sa_snapshot[0][14] , \sa_snapshot[0].f.lower[14] );
tran (\sa_snapshot[0][15] , \sa_snapshot[0].r.part0[15] );
tran (\sa_snapshot[0][15] , \sa_snapshot[0].f.lower[15] );
tran (\sa_snapshot[0][16] , \sa_snapshot[0].r.part0[16] );
tran (\sa_snapshot[0][16] , \sa_snapshot[0].f.lower[16] );
tran (\sa_snapshot[0][17] , \sa_snapshot[0].r.part0[17] );
tran (\sa_snapshot[0][17] , \sa_snapshot[0].f.lower[17] );
tran (\sa_snapshot[0][18] , \sa_snapshot[0].r.part0[18] );
tran (\sa_snapshot[0][18] , \sa_snapshot[0].f.lower[18] );
tran (\sa_snapshot[0][19] , \sa_snapshot[0].r.part0[19] );
tran (\sa_snapshot[0][19] , \sa_snapshot[0].f.lower[19] );
tran (\sa_snapshot[0][20] , \sa_snapshot[0].r.part0[20] );
tran (\sa_snapshot[0][20] , \sa_snapshot[0].f.lower[20] );
tran (\sa_snapshot[0][21] , \sa_snapshot[0].r.part0[21] );
tran (\sa_snapshot[0][21] , \sa_snapshot[0].f.lower[21] );
tran (\sa_snapshot[0][22] , \sa_snapshot[0].r.part0[22] );
tran (\sa_snapshot[0][22] , \sa_snapshot[0].f.lower[22] );
tran (\sa_snapshot[0][23] , \sa_snapshot[0].r.part0[23] );
tran (\sa_snapshot[0][23] , \sa_snapshot[0].f.lower[23] );
tran (\sa_snapshot[0][24] , \sa_snapshot[0].r.part0[24] );
tran (\sa_snapshot[0][24] , \sa_snapshot[0].f.lower[24] );
tran (\sa_snapshot[0][25] , \sa_snapshot[0].r.part0[25] );
tran (\sa_snapshot[0][25] , \sa_snapshot[0].f.lower[25] );
tran (\sa_snapshot[0][26] , \sa_snapshot[0].r.part0[26] );
tran (\sa_snapshot[0][26] , \sa_snapshot[0].f.lower[26] );
tran (\sa_snapshot[0][27] , \sa_snapshot[0].r.part0[27] );
tran (\sa_snapshot[0][27] , \sa_snapshot[0].f.lower[27] );
tran (\sa_snapshot[0][28] , \sa_snapshot[0].r.part0[28] );
tran (\sa_snapshot[0][28] , \sa_snapshot[0].f.lower[28] );
tran (\sa_snapshot[0][29] , \sa_snapshot[0].r.part0[29] );
tran (\sa_snapshot[0][29] , \sa_snapshot[0].f.lower[29] );
tran (\sa_snapshot[0][30] , \sa_snapshot[0].r.part0[30] );
tran (\sa_snapshot[0][30] , \sa_snapshot[0].f.lower[30] );
tran (\sa_snapshot[0][31] , \sa_snapshot[0].r.part0[31] );
tran (\sa_snapshot[0][31] , \sa_snapshot[0].f.lower[31] );
tran (\sa_snapshot[0][32] , \sa_snapshot[0].r.part1[0] );
tran (\sa_snapshot[0][32] , \sa_snapshot[0].f.upper[0] );
tran (\sa_snapshot[0][33] , \sa_snapshot[0].r.part1[1] );
tran (\sa_snapshot[0][33] , \sa_snapshot[0].f.upper[1] );
tran (\sa_snapshot[0][34] , \sa_snapshot[0].r.part1[2] );
tran (\sa_snapshot[0][34] , \sa_snapshot[0].f.upper[2] );
tran (\sa_snapshot[0][35] , \sa_snapshot[0].r.part1[3] );
tran (\sa_snapshot[0][35] , \sa_snapshot[0].f.upper[3] );
tran (\sa_snapshot[0][36] , \sa_snapshot[0].r.part1[4] );
tran (\sa_snapshot[0][36] , \sa_snapshot[0].f.upper[4] );
tran (\sa_snapshot[0][37] , \sa_snapshot[0].r.part1[5] );
tran (\sa_snapshot[0][37] , \sa_snapshot[0].f.upper[5] );
tran (\sa_snapshot[0][38] , \sa_snapshot[0].r.part1[6] );
tran (\sa_snapshot[0][38] , \sa_snapshot[0].f.upper[6] );
tran (\sa_snapshot[0][39] , \sa_snapshot[0].r.part1[7] );
tran (\sa_snapshot[0][39] , \sa_snapshot[0].f.upper[7] );
tran (\sa_snapshot[0][40] , \sa_snapshot[0].r.part1[8] );
tran (\sa_snapshot[0][40] , \sa_snapshot[0].f.upper[8] );
tran (\sa_snapshot[0][41] , \sa_snapshot[0].r.part1[9] );
tran (\sa_snapshot[0][41] , \sa_snapshot[0].f.upper[9] );
tran (\sa_snapshot[0][42] , \sa_snapshot[0].r.part1[10] );
tran (\sa_snapshot[0][42] , \sa_snapshot[0].f.upper[10] );
tran (\sa_snapshot[0][43] , \sa_snapshot[0].r.part1[11] );
tran (\sa_snapshot[0][43] , \sa_snapshot[0].f.upper[11] );
tran (\sa_snapshot[0][44] , \sa_snapshot[0].r.part1[12] );
tran (\sa_snapshot[0][44] , \sa_snapshot[0].f.upper[12] );
tran (\sa_snapshot[0][45] , \sa_snapshot[0].r.part1[13] );
tran (\sa_snapshot[0][45] , \sa_snapshot[0].f.upper[13] );
tran (\sa_snapshot[0][46] , \sa_snapshot[0].r.part1[14] );
tran (\sa_snapshot[0][46] , \sa_snapshot[0].f.upper[14] );
tran (\sa_snapshot[0][47] , \sa_snapshot[0].r.part1[15] );
tran (\sa_snapshot[0][47] , \sa_snapshot[0].f.upper[15] );
tran (\sa_snapshot[0][48] , \sa_snapshot[0].r.part1[16] );
tran (\sa_snapshot[0][48] , \sa_snapshot[0].f.upper[16] );
tran (\sa_snapshot[0][49] , \sa_snapshot[0].r.part1[17] );
tran (\sa_snapshot[0][49] , \sa_snapshot[0].f.upper[17] );
tran (\sa_snapshot[0][50] , \sa_snapshot[0].r.part1[18] );
tran (\sa_snapshot[0][50] , \sa_snapshot[0].f.unused[0] );
tran (\sa_snapshot[0][51] , \sa_snapshot[0].r.part1[19] );
tran (\sa_snapshot[0][51] , \sa_snapshot[0].f.unused[1] );
tran (\sa_snapshot[0][52] , \sa_snapshot[0].r.part1[20] );
tran (\sa_snapshot[0][52] , \sa_snapshot[0].f.unused[2] );
tran (\sa_snapshot[0][53] , \sa_snapshot[0].r.part1[21] );
tran (\sa_snapshot[0][53] , \sa_snapshot[0].f.unused[3] );
tran (\sa_snapshot[0][54] , \sa_snapshot[0].r.part1[22] );
tran (\sa_snapshot[0][54] , \sa_snapshot[0].f.unused[4] );
tran (\sa_snapshot[0][55] , \sa_snapshot[0].r.part1[23] );
tran (\sa_snapshot[0][55] , \sa_snapshot[0].f.unused[5] );
tran (\sa_snapshot[0][56] , \sa_snapshot[0].r.part1[24] );
tran (\sa_snapshot[0][56] , \sa_snapshot[0].f.unused[6] );
tran (\sa_snapshot[0][57] , \sa_snapshot[0].r.part1[25] );
tran (\sa_snapshot[0][57] , \sa_snapshot[0].f.unused[7] );
tran (\sa_snapshot[0][58] , \sa_snapshot[0].r.part1[26] );
tran (\sa_snapshot[0][58] , \sa_snapshot[0].f.unused[8] );
tran (\sa_snapshot[0][59] , \sa_snapshot[0].r.part1[27] );
tran (\sa_snapshot[0][59] , \sa_snapshot[0].f.unused[9] );
tran (\sa_snapshot[0][60] , \sa_snapshot[0].r.part1[28] );
tran (\sa_snapshot[0][60] , \sa_snapshot[0].f.unused[10] );
tran (\sa_snapshot[0][61] , \sa_snapshot[0].r.part1[29] );
tran (\sa_snapshot[0][61] , \sa_snapshot[0].f.unused[11] );
tran (\sa_snapshot[0][62] , \sa_snapshot[0].r.part1[30] );
tran (\sa_snapshot[0][62] , \sa_snapshot[0].f.unused[12] );
tran (\sa_snapshot[0][63] , \sa_snapshot[0].r.part1[31] );
tran (\sa_snapshot[0][63] , \sa_snapshot[0].f.unused[13] );
tran (\sa_snapshot[1][0] , \sa_snapshot[1].r.part0[0] );
tran (\sa_snapshot[1][0] , \sa_snapshot[1].f.lower[0] );
tran (\sa_snapshot[1][1] , \sa_snapshot[1].r.part0[1] );
tran (\sa_snapshot[1][1] , \sa_snapshot[1].f.lower[1] );
tran (\sa_snapshot[1][2] , \sa_snapshot[1].r.part0[2] );
tran (\sa_snapshot[1][2] , \sa_snapshot[1].f.lower[2] );
tran (\sa_snapshot[1][3] , \sa_snapshot[1].r.part0[3] );
tran (\sa_snapshot[1][3] , \sa_snapshot[1].f.lower[3] );
tran (\sa_snapshot[1][4] , \sa_snapshot[1].r.part0[4] );
tran (\sa_snapshot[1][4] , \sa_snapshot[1].f.lower[4] );
tran (\sa_snapshot[1][5] , \sa_snapshot[1].r.part0[5] );
tran (\sa_snapshot[1][5] , \sa_snapshot[1].f.lower[5] );
tran (\sa_snapshot[1][6] , \sa_snapshot[1].r.part0[6] );
tran (\sa_snapshot[1][6] , \sa_snapshot[1].f.lower[6] );
tran (\sa_snapshot[1][7] , \sa_snapshot[1].r.part0[7] );
tran (\sa_snapshot[1][7] , \sa_snapshot[1].f.lower[7] );
tran (\sa_snapshot[1][8] , \sa_snapshot[1].r.part0[8] );
tran (\sa_snapshot[1][8] , \sa_snapshot[1].f.lower[8] );
tran (\sa_snapshot[1][9] , \sa_snapshot[1].r.part0[9] );
tran (\sa_snapshot[1][9] , \sa_snapshot[1].f.lower[9] );
tran (\sa_snapshot[1][10] , \sa_snapshot[1].r.part0[10] );
tran (\sa_snapshot[1][10] , \sa_snapshot[1].f.lower[10] );
tran (\sa_snapshot[1][11] , \sa_snapshot[1].r.part0[11] );
tran (\sa_snapshot[1][11] , \sa_snapshot[1].f.lower[11] );
tran (\sa_snapshot[1][12] , \sa_snapshot[1].r.part0[12] );
tran (\sa_snapshot[1][12] , \sa_snapshot[1].f.lower[12] );
tran (\sa_snapshot[1][13] , \sa_snapshot[1].r.part0[13] );
tran (\sa_snapshot[1][13] , \sa_snapshot[1].f.lower[13] );
tran (\sa_snapshot[1][14] , \sa_snapshot[1].r.part0[14] );
tran (\sa_snapshot[1][14] , \sa_snapshot[1].f.lower[14] );
tran (\sa_snapshot[1][15] , \sa_snapshot[1].r.part0[15] );
tran (\sa_snapshot[1][15] , \sa_snapshot[1].f.lower[15] );
tran (\sa_snapshot[1][16] , \sa_snapshot[1].r.part0[16] );
tran (\sa_snapshot[1][16] , \sa_snapshot[1].f.lower[16] );
tran (\sa_snapshot[1][17] , \sa_snapshot[1].r.part0[17] );
tran (\sa_snapshot[1][17] , \sa_snapshot[1].f.lower[17] );
tran (\sa_snapshot[1][18] , \sa_snapshot[1].r.part0[18] );
tran (\sa_snapshot[1][18] , \sa_snapshot[1].f.lower[18] );
tran (\sa_snapshot[1][19] , \sa_snapshot[1].r.part0[19] );
tran (\sa_snapshot[1][19] , \sa_snapshot[1].f.lower[19] );
tran (\sa_snapshot[1][20] , \sa_snapshot[1].r.part0[20] );
tran (\sa_snapshot[1][20] , \sa_snapshot[1].f.lower[20] );
tran (\sa_snapshot[1][21] , \sa_snapshot[1].r.part0[21] );
tran (\sa_snapshot[1][21] , \sa_snapshot[1].f.lower[21] );
tran (\sa_snapshot[1][22] , \sa_snapshot[1].r.part0[22] );
tran (\sa_snapshot[1][22] , \sa_snapshot[1].f.lower[22] );
tran (\sa_snapshot[1][23] , \sa_snapshot[1].r.part0[23] );
tran (\sa_snapshot[1][23] , \sa_snapshot[1].f.lower[23] );
tran (\sa_snapshot[1][24] , \sa_snapshot[1].r.part0[24] );
tran (\sa_snapshot[1][24] , \sa_snapshot[1].f.lower[24] );
tran (\sa_snapshot[1][25] , \sa_snapshot[1].r.part0[25] );
tran (\sa_snapshot[1][25] , \sa_snapshot[1].f.lower[25] );
tran (\sa_snapshot[1][26] , \sa_snapshot[1].r.part0[26] );
tran (\sa_snapshot[1][26] , \sa_snapshot[1].f.lower[26] );
tran (\sa_snapshot[1][27] , \sa_snapshot[1].r.part0[27] );
tran (\sa_snapshot[1][27] , \sa_snapshot[1].f.lower[27] );
tran (\sa_snapshot[1][28] , \sa_snapshot[1].r.part0[28] );
tran (\sa_snapshot[1][28] , \sa_snapshot[1].f.lower[28] );
tran (\sa_snapshot[1][29] , \sa_snapshot[1].r.part0[29] );
tran (\sa_snapshot[1][29] , \sa_snapshot[1].f.lower[29] );
tran (\sa_snapshot[1][30] , \sa_snapshot[1].r.part0[30] );
tran (\sa_snapshot[1][30] , \sa_snapshot[1].f.lower[30] );
tran (\sa_snapshot[1][31] , \sa_snapshot[1].r.part0[31] );
tran (\sa_snapshot[1][31] , \sa_snapshot[1].f.lower[31] );
tran (\sa_snapshot[1][32] , \sa_snapshot[1].r.part1[0] );
tran (\sa_snapshot[1][32] , \sa_snapshot[1].f.upper[0] );
tran (\sa_snapshot[1][33] , \sa_snapshot[1].r.part1[1] );
tran (\sa_snapshot[1][33] , \sa_snapshot[1].f.upper[1] );
tran (\sa_snapshot[1][34] , \sa_snapshot[1].r.part1[2] );
tran (\sa_snapshot[1][34] , \sa_snapshot[1].f.upper[2] );
tran (\sa_snapshot[1][35] , \sa_snapshot[1].r.part1[3] );
tran (\sa_snapshot[1][35] , \sa_snapshot[1].f.upper[3] );
tran (\sa_snapshot[1][36] , \sa_snapshot[1].r.part1[4] );
tran (\sa_snapshot[1][36] , \sa_snapshot[1].f.upper[4] );
tran (\sa_snapshot[1][37] , \sa_snapshot[1].r.part1[5] );
tran (\sa_snapshot[1][37] , \sa_snapshot[1].f.upper[5] );
tran (\sa_snapshot[1][38] , \sa_snapshot[1].r.part1[6] );
tran (\sa_snapshot[1][38] , \sa_snapshot[1].f.upper[6] );
tran (\sa_snapshot[1][39] , \sa_snapshot[1].r.part1[7] );
tran (\sa_snapshot[1][39] , \sa_snapshot[1].f.upper[7] );
tran (\sa_snapshot[1][40] , \sa_snapshot[1].r.part1[8] );
tran (\sa_snapshot[1][40] , \sa_snapshot[1].f.upper[8] );
tran (\sa_snapshot[1][41] , \sa_snapshot[1].r.part1[9] );
tran (\sa_snapshot[1][41] , \sa_snapshot[1].f.upper[9] );
tran (\sa_snapshot[1][42] , \sa_snapshot[1].r.part1[10] );
tran (\sa_snapshot[1][42] , \sa_snapshot[1].f.upper[10] );
tran (\sa_snapshot[1][43] , \sa_snapshot[1].r.part1[11] );
tran (\sa_snapshot[1][43] , \sa_snapshot[1].f.upper[11] );
tran (\sa_snapshot[1][44] , \sa_snapshot[1].r.part1[12] );
tran (\sa_snapshot[1][44] , \sa_snapshot[1].f.upper[12] );
tran (\sa_snapshot[1][45] , \sa_snapshot[1].r.part1[13] );
tran (\sa_snapshot[1][45] , \sa_snapshot[1].f.upper[13] );
tran (\sa_snapshot[1][46] , \sa_snapshot[1].r.part1[14] );
tran (\sa_snapshot[1][46] , \sa_snapshot[1].f.upper[14] );
tran (\sa_snapshot[1][47] , \sa_snapshot[1].r.part1[15] );
tran (\sa_snapshot[1][47] , \sa_snapshot[1].f.upper[15] );
tran (\sa_snapshot[1][48] , \sa_snapshot[1].r.part1[16] );
tran (\sa_snapshot[1][48] , \sa_snapshot[1].f.upper[16] );
tran (\sa_snapshot[1][49] , \sa_snapshot[1].r.part1[17] );
tran (\sa_snapshot[1][49] , \sa_snapshot[1].f.upper[17] );
tran (\sa_snapshot[1][50] , \sa_snapshot[1].r.part1[18] );
tran (\sa_snapshot[1][50] , \sa_snapshot[1].f.unused[0] );
tran (\sa_snapshot[1][51] , \sa_snapshot[1].r.part1[19] );
tran (\sa_snapshot[1][51] , \sa_snapshot[1].f.unused[1] );
tran (\sa_snapshot[1][52] , \sa_snapshot[1].r.part1[20] );
tran (\sa_snapshot[1][52] , \sa_snapshot[1].f.unused[2] );
tran (\sa_snapshot[1][53] , \sa_snapshot[1].r.part1[21] );
tran (\sa_snapshot[1][53] , \sa_snapshot[1].f.unused[3] );
tran (\sa_snapshot[1][54] , \sa_snapshot[1].r.part1[22] );
tran (\sa_snapshot[1][54] , \sa_snapshot[1].f.unused[4] );
tran (\sa_snapshot[1][55] , \sa_snapshot[1].r.part1[23] );
tran (\sa_snapshot[1][55] , \sa_snapshot[1].f.unused[5] );
tran (\sa_snapshot[1][56] , \sa_snapshot[1].r.part1[24] );
tran (\sa_snapshot[1][56] , \sa_snapshot[1].f.unused[6] );
tran (\sa_snapshot[1][57] , \sa_snapshot[1].r.part1[25] );
tran (\sa_snapshot[1][57] , \sa_snapshot[1].f.unused[7] );
tran (\sa_snapshot[1][58] , \sa_snapshot[1].r.part1[26] );
tran (\sa_snapshot[1][58] , \sa_snapshot[1].f.unused[8] );
tran (\sa_snapshot[1][59] , \sa_snapshot[1].r.part1[27] );
tran (\sa_snapshot[1][59] , \sa_snapshot[1].f.unused[9] );
tran (\sa_snapshot[1][60] , \sa_snapshot[1].r.part1[28] );
tran (\sa_snapshot[1][60] , \sa_snapshot[1].f.unused[10] );
tran (\sa_snapshot[1][61] , \sa_snapshot[1].r.part1[29] );
tran (\sa_snapshot[1][61] , \sa_snapshot[1].f.unused[11] );
tran (\sa_snapshot[1][62] , \sa_snapshot[1].r.part1[30] );
tran (\sa_snapshot[1][62] , \sa_snapshot[1].f.unused[12] );
tran (\sa_snapshot[1][63] , \sa_snapshot[1].r.part1[31] );
tran (\sa_snapshot[1][63] , \sa_snapshot[1].f.unused[13] );
tran (\sa_snapshot[2][0] , \sa_snapshot[2].r.part0[0] );
tran (\sa_snapshot[2][0] , \sa_snapshot[2].f.lower[0] );
tran (\sa_snapshot[2][1] , \sa_snapshot[2].r.part0[1] );
tran (\sa_snapshot[2][1] , \sa_snapshot[2].f.lower[1] );
tran (\sa_snapshot[2][2] , \sa_snapshot[2].r.part0[2] );
tran (\sa_snapshot[2][2] , \sa_snapshot[2].f.lower[2] );
tran (\sa_snapshot[2][3] , \sa_snapshot[2].r.part0[3] );
tran (\sa_snapshot[2][3] , \sa_snapshot[2].f.lower[3] );
tran (\sa_snapshot[2][4] , \sa_snapshot[2].r.part0[4] );
tran (\sa_snapshot[2][4] , \sa_snapshot[2].f.lower[4] );
tran (\sa_snapshot[2][5] , \sa_snapshot[2].r.part0[5] );
tran (\sa_snapshot[2][5] , \sa_snapshot[2].f.lower[5] );
tran (\sa_snapshot[2][6] , \sa_snapshot[2].r.part0[6] );
tran (\sa_snapshot[2][6] , \sa_snapshot[2].f.lower[6] );
tran (\sa_snapshot[2][7] , \sa_snapshot[2].r.part0[7] );
tran (\sa_snapshot[2][7] , \sa_snapshot[2].f.lower[7] );
tran (\sa_snapshot[2][8] , \sa_snapshot[2].r.part0[8] );
tran (\sa_snapshot[2][8] , \sa_snapshot[2].f.lower[8] );
tran (\sa_snapshot[2][9] , \sa_snapshot[2].r.part0[9] );
tran (\sa_snapshot[2][9] , \sa_snapshot[2].f.lower[9] );
tran (\sa_snapshot[2][10] , \sa_snapshot[2].r.part0[10] );
tran (\sa_snapshot[2][10] , \sa_snapshot[2].f.lower[10] );
tran (\sa_snapshot[2][11] , \sa_snapshot[2].r.part0[11] );
tran (\sa_snapshot[2][11] , \sa_snapshot[2].f.lower[11] );
tran (\sa_snapshot[2][12] , \sa_snapshot[2].r.part0[12] );
tran (\sa_snapshot[2][12] , \sa_snapshot[2].f.lower[12] );
tran (\sa_snapshot[2][13] , \sa_snapshot[2].r.part0[13] );
tran (\sa_snapshot[2][13] , \sa_snapshot[2].f.lower[13] );
tran (\sa_snapshot[2][14] , \sa_snapshot[2].r.part0[14] );
tran (\sa_snapshot[2][14] , \sa_snapshot[2].f.lower[14] );
tran (\sa_snapshot[2][15] , \sa_snapshot[2].r.part0[15] );
tran (\sa_snapshot[2][15] , \sa_snapshot[2].f.lower[15] );
tran (\sa_snapshot[2][16] , \sa_snapshot[2].r.part0[16] );
tran (\sa_snapshot[2][16] , \sa_snapshot[2].f.lower[16] );
tran (\sa_snapshot[2][17] , \sa_snapshot[2].r.part0[17] );
tran (\sa_snapshot[2][17] , \sa_snapshot[2].f.lower[17] );
tran (\sa_snapshot[2][18] , \sa_snapshot[2].r.part0[18] );
tran (\sa_snapshot[2][18] , \sa_snapshot[2].f.lower[18] );
tran (\sa_snapshot[2][19] , \sa_snapshot[2].r.part0[19] );
tran (\sa_snapshot[2][19] , \sa_snapshot[2].f.lower[19] );
tran (\sa_snapshot[2][20] , \sa_snapshot[2].r.part0[20] );
tran (\sa_snapshot[2][20] , \sa_snapshot[2].f.lower[20] );
tran (\sa_snapshot[2][21] , \sa_snapshot[2].r.part0[21] );
tran (\sa_snapshot[2][21] , \sa_snapshot[2].f.lower[21] );
tran (\sa_snapshot[2][22] , \sa_snapshot[2].r.part0[22] );
tran (\sa_snapshot[2][22] , \sa_snapshot[2].f.lower[22] );
tran (\sa_snapshot[2][23] , \sa_snapshot[2].r.part0[23] );
tran (\sa_snapshot[2][23] , \sa_snapshot[2].f.lower[23] );
tran (\sa_snapshot[2][24] , \sa_snapshot[2].r.part0[24] );
tran (\sa_snapshot[2][24] , \sa_snapshot[2].f.lower[24] );
tran (\sa_snapshot[2][25] , \sa_snapshot[2].r.part0[25] );
tran (\sa_snapshot[2][25] , \sa_snapshot[2].f.lower[25] );
tran (\sa_snapshot[2][26] , \sa_snapshot[2].r.part0[26] );
tran (\sa_snapshot[2][26] , \sa_snapshot[2].f.lower[26] );
tran (\sa_snapshot[2][27] , \sa_snapshot[2].r.part0[27] );
tran (\sa_snapshot[2][27] , \sa_snapshot[2].f.lower[27] );
tran (\sa_snapshot[2][28] , \sa_snapshot[2].r.part0[28] );
tran (\sa_snapshot[2][28] , \sa_snapshot[2].f.lower[28] );
tran (\sa_snapshot[2][29] , \sa_snapshot[2].r.part0[29] );
tran (\sa_snapshot[2][29] , \sa_snapshot[2].f.lower[29] );
tran (\sa_snapshot[2][30] , \sa_snapshot[2].r.part0[30] );
tran (\sa_snapshot[2][30] , \sa_snapshot[2].f.lower[30] );
tran (\sa_snapshot[2][31] , \sa_snapshot[2].r.part0[31] );
tran (\sa_snapshot[2][31] , \sa_snapshot[2].f.lower[31] );
tran (\sa_snapshot[2][32] , \sa_snapshot[2].r.part1[0] );
tran (\sa_snapshot[2][32] , \sa_snapshot[2].f.upper[0] );
tran (\sa_snapshot[2][33] , \sa_snapshot[2].r.part1[1] );
tran (\sa_snapshot[2][33] , \sa_snapshot[2].f.upper[1] );
tran (\sa_snapshot[2][34] , \sa_snapshot[2].r.part1[2] );
tran (\sa_snapshot[2][34] , \sa_snapshot[2].f.upper[2] );
tran (\sa_snapshot[2][35] , \sa_snapshot[2].r.part1[3] );
tran (\sa_snapshot[2][35] , \sa_snapshot[2].f.upper[3] );
tran (\sa_snapshot[2][36] , \sa_snapshot[2].r.part1[4] );
tran (\sa_snapshot[2][36] , \sa_snapshot[2].f.upper[4] );
tran (\sa_snapshot[2][37] , \sa_snapshot[2].r.part1[5] );
tran (\sa_snapshot[2][37] , \sa_snapshot[2].f.upper[5] );
tran (\sa_snapshot[2][38] , \sa_snapshot[2].r.part1[6] );
tran (\sa_snapshot[2][38] , \sa_snapshot[2].f.upper[6] );
tran (\sa_snapshot[2][39] , \sa_snapshot[2].r.part1[7] );
tran (\sa_snapshot[2][39] , \sa_snapshot[2].f.upper[7] );
tran (\sa_snapshot[2][40] , \sa_snapshot[2].r.part1[8] );
tran (\sa_snapshot[2][40] , \sa_snapshot[2].f.upper[8] );
tran (\sa_snapshot[2][41] , \sa_snapshot[2].r.part1[9] );
tran (\sa_snapshot[2][41] , \sa_snapshot[2].f.upper[9] );
tran (\sa_snapshot[2][42] , \sa_snapshot[2].r.part1[10] );
tran (\sa_snapshot[2][42] , \sa_snapshot[2].f.upper[10] );
tran (\sa_snapshot[2][43] , \sa_snapshot[2].r.part1[11] );
tran (\sa_snapshot[2][43] , \sa_snapshot[2].f.upper[11] );
tran (\sa_snapshot[2][44] , \sa_snapshot[2].r.part1[12] );
tran (\sa_snapshot[2][44] , \sa_snapshot[2].f.upper[12] );
tran (\sa_snapshot[2][45] , \sa_snapshot[2].r.part1[13] );
tran (\sa_snapshot[2][45] , \sa_snapshot[2].f.upper[13] );
tran (\sa_snapshot[2][46] , \sa_snapshot[2].r.part1[14] );
tran (\sa_snapshot[2][46] , \sa_snapshot[2].f.upper[14] );
tran (\sa_snapshot[2][47] , \sa_snapshot[2].r.part1[15] );
tran (\sa_snapshot[2][47] , \sa_snapshot[2].f.upper[15] );
tran (\sa_snapshot[2][48] , \sa_snapshot[2].r.part1[16] );
tran (\sa_snapshot[2][48] , \sa_snapshot[2].f.upper[16] );
tran (\sa_snapshot[2][49] , \sa_snapshot[2].r.part1[17] );
tran (\sa_snapshot[2][49] , \sa_snapshot[2].f.upper[17] );
tran (\sa_snapshot[2][50] , \sa_snapshot[2].r.part1[18] );
tran (\sa_snapshot[2][50] , \sa_snapshot[2].f.unused[0] );
tran (\sa_snapshot[2][51] , \sa_snapshot[2].r.part1[19] );
tran (\sa_snapshot[2][51] , \sa_snapshot[2].f.unused[1] );
tran (\sa_snapshot[2][52] , \sa_snapshot[2].r.part1[20] );
tran (\sa_snapshot[2][52] , \sa_snapshot[2].f.unused[2] );
tran (\sa_snapshot[2][53] , \sa_snapshot[2].r.part1[21] );
tran (\sa_snapshot[2][53] , \sa_snapshot[2].f.unused[3] );
tran (\sa_snapshot[2][54] , \sa_snapshot[2].r.part1[22] );
tran (\sa_snapshot[2][54] , \sa_snapshot[2].f.unused[4] );
tran (\sa_snapshot[2][55] , \sa_snapshot[2].r.part1[23] );
tran (\sa_snapshot[2][55] , \sa_snapshot[2].f.unused[5] );
tran (\sa_snapshot[2][56] , \sa_snapshot[2].r.part1[24] );
tran (\sa_snapshot[2][56] , \sa_snapshot[2].f.unused[6] );
tran (\sa_snapshot[2][57] , \sa_snapshot[2].r.part1[25] );
tran (\sa_snapshot[2][57] , \sa_snapshot[2].f.unused[7] );
tran (\sa_snapshot[2][58] , \sa_snapshot[2].r.part1[26] );
tran (\sa_snapshot[2][58] , \sa_snapshot[2].f.unused[8] );
tran (\sa_snapshot[2][59] , \sa_snapshot[2].r.part1[27] );
tran (\sa_snapshot[2][59] , \sa_snapshot[2].f.unused[9] );
tran (\sa_snapshot[2][60] , \sa_snapshot[2].r.part1[28] );
tran (\sa_snapshot[2][60] , \sa_snapshot[2].f.unused[10] );
tran (\sa_snapshot[2][61] , \sa_snapshot[2].r.part1[29] );
tran (\sa_snapshot[2][61] , \sa_snapshot[2].f.unused[11] );
tran (\sa_snapshot[2][62] , \sa_snapshot[2].r.part1[30] );
tran (\sa_snapshot[2][62] , \sa_snapshot[2].f.unused[12] );
tran (\sa_snapshot[2][63] , \sa_snapshot[2].r.part1[31] );
tran (\sa_snapshot[2][63] , \sa_snapshot[2].f.unused[13] );
tran (\sa_snapshot[3][0] , \sa_snapshot[3].r.part0[0] );
tran (\sa_snapshot[3][0] , \sa_snapshot[3].f.lower[0] );
tran (\sa_snapshot[3][1] , \sa_snapshot[3].r.part0[1] );
tran (\sa_snapshot[3][1] , \sa_snapshot[3].f.lower[1] );
tran (\sa_snapshot[3][2] , \sa_snapshot[3].r.part0[2] );
tran (\sa_snapshot[3][2] , \sa_snapshot[3].f.lower[2] );
tran (\sa_snapshot[3][3] , \sa_snapshot[3].r.part0[3] );
tran (\sa_snapshot[3][3] , \sa_snapshot[3].f.lower[3] );
tran (\sa_snapshot[3][4] , \sa_snapshot[3].r.part0[4] );
tran (\sa_snapshot[3][4] , \sa_snapshot[3].f.lower[4] );
tran (\sa_snapshot[3][5] , \sa_snapshot[3].r.part0[5] );
tran (\sa_snapshot[3][5] , \sa_snapshot[3].f.lower[5] );
tran (\sa_snapshot[3][6] , \sa_snapshot[3].r.part0[6] );
tran (\sa_snapshot[3][6] , \sa_snapshot[3].f.lower[6] );
tran (\sa_snapshot[3][7] , \sa_snapshot[3].r.part0[7] );
tran (\sa_snapshot[3][7] , \sa_snapshot[3].f.lower[7] );
tran (\sa_snapshot[3][8] , \sa_snapshot[3].r.part0[8] );
tran (\sa_snapshot[3][8] , \sa_snapshot[3].f.lower[8] );
tran (\sa_snapshot[3][9] , \sa_snapshot[3].r.part0[9] );
tran (\sa_snapshot[3][9] , \sa_snapshot[3].f.lower[9] );
tran (\sa_snapshot[3][10] , \sa_snapshot[3].r.part0[10] );
tran (\sa_snapshot[3][10] , \sa_snapshot[3].f.lower[10] );
tran (\sa_snapshot[3][11] , \sa_snapshot[3].r.part0[11] );
tran (\sa_snapshot[3][11] , \sa_snapshot[3].f.lower[11] );
tran (\sa_snapshot[3][12] , \sa_snapshot[3].r.part0[12] );
tran (\sa_snapshot[3][12] , \sa_snapshot[3].f.lower[12] );
tran (\sa_snapshot[3][13] , \sa_snapshot[3].r.part0[13] );
tran (\sa_snapshot[3][13] , \sa_snapshot[3].f.lower[13] );
tran (\sa_snapshot[3][14] , \sa_snapshot[3].r.part0[14] );
tran (\sa_snapshot[3][14] , \sa_snapshot[3].f.lower[14] );
tran (\sa_snapshot[3][15] , \sa_snapshot[3].r.part0[15] );
tran (\sa_snapshot[3][15] , \sa_snapshot[3].f.lower[15] );
tran (\sa_snapshot[3][16] , \sa_snapshot[3].r.part0[16] );
tran (\sa_snapshot[3][16] , \sa_snapshot[3].f.lower[16] );
tran (\sa_snapshot[3][17] , \sa_snapshot[3].r.part0[17] );
tran (\sa_snapshot[3][17] , \sa_snapshot[3].f.lower[17] );
tran (\sa_snapshot[3][18] , \sa_snapshot[3].r.part0[18] );
tran (\sa_snapshot[3][18] , \sa_snapshot[3].f.lower[18] );
tran (\sa_snapshot[3][19] , \sa_snapshot[3].r.part0[19] );
tran (\sa_snapshot[3][19] , \sa_snapshot[3].f.lower[19] );
tran (\sa_snapshot[3][20] , \sa_snapshot[3].r.part0[20] );
tran (\sa_snapshot[3][20] , \sa_snapshot[3].f.lower[20] );
tran (\sa_snapshot[3][21] , \sa_snapshot[3].r.part0[21] );
tran (\sa_snapshot[3][21] , \sa_snapshot[3].f.lower[21] );
tran (\sa_snapshot[3][22] , \sa_snapshot[3].r.part0[22] );
tran (\sa_snapshot[3][22] , \sa_snapshot[3].f.lower[22] );
tran (\sa_snapshot[3][23] , \sa_snapshot[3].r.part0[23] );
tran (\sa_snapshot[3][23] , \sa_snapshot[3].f.lower[23] );
tran (\sa_snapshot[3][24] , \sa_snapshot[3].r.part0[24] );
tran (\sa_snapshot[3][24] , \sa_snapshot[3].f.lower[24] );
tran (\sa_snapshot[3][25] , \sa_snapshot[3].r.part0[25] );
tran (\sa_snapshot[3][25] , \sa_snapshot[3].f.lower[25] );
tran (\sa_snapshot[3][26] , \sa_snapshot[3].r.part0[26] );
tran (\sa_snapshot[3][26] , \sa_snapshot[3].f.lower[26] );
tran (\sa_snapshot[3][27] , \sa_snapshot[3].r.part0[27] );
tran (\sa_snapshot[3][27] , \sa_snapshot[3].f.lower[27] );
tran (\sa_snapshot[3][28] , \sa_snapshot[3].r.part0[28] );
tran (\sa_snapshot[3][28] , \sa_snapshot[3].f.lower[28] );
tran (\sa_snapshot[3][29] , \sa_snapshot[3].r.part0[29] );
tran (\sa_snapshot[3][29] , \sa_snapshot[3].f.lower[29] );
tran (\sa_snapshot[3][30] , \sa_snapshot[3].r.part0[30] );
tran (\sa_snapshot[3][30] , \sa_snapshot[3].f.lower[30] );
tran (\sa_snapshot[3][31] , \sa_snapshot[3].r.part0[31] );
tran (\sa_snapshot[3][31] , \sa_snapshot[3].f.lower[31] );
tran (\sa_snapshot[3][32] , \sa_snapshot[3].r.part1[0] );
tran (\sa_snapshot[3][32] , \sa_snapshot[3].f.upper[0] );
tran (\sa_snapshot[3][33] , \sa_snapshot[3].r.part1[1] );
tran (\sa_snapshot[3][33] , \sa_snapshot[3].f.upper[1] );
tran (\sa_snapshot[3][34] , \sa_snapshot[3].r.part1[2] );
tran (\sa_snapshot[3][34] , \sa_snapshot[3].f.upper[2] );
tran (\sa_snapshot[3][35] , \sa_snapshot[3].r.part1[3] );
tran (\sa_snapshot[3][35] , \sa_snapshot[3].f.upper[3] );
tran (\sa_snapshot[3][36] , \sa_snapshot[3].r.part1[4] );
tran (\sa_snapshot[3][36] , \sa_snapshot[3].f.upper[4] );
tran (\sa_snapshot[3][37] , \sa_snapshot[3].r.part1[5] );
tran (\sa_snapshot[3][37] , \sa_snapshot[3].f.upper[5] );
tran (\sa_snapshot[3][38] , \sa_snapshot[3].r.part1[6] );
tran (\sa_snapshot[3][38] , \sa_snapshot[3].f.upper[6] );
tran (\sa_snapshot[3][39] , \sa_snapshot[3].r.part1[7] );
tran (\sa_snapshot[3][39] , \sa_snapshot[3].f.upper[7] );
tran (\sa_snapshot[3][40] , \sa_snapshot[3].r.part1[8] );
tran (\sa_snapshot[3][40] , \sa_snapshot[3].f.upper[8] );
tran (\sa_snapshot[3][41] , \sa_snapshot[3].r.part1[9] );
tran (\sa_snapshot[3][41] , \sa_snapshot[3].f.upper[9] );
tran (\sa_snapshot[3][42] , \sa_snapshot[3].r.part1[10] );
tran (\sa_snapshot[3][42] , \sa_snapshot[3].f.upper[10] );
tran (\sa_snapshot[3][43] , \sa_snapshot[3].r.part1[11] );
tran (\sa_snapshot[3][43] , \sa_snapshot[3].f.upper[11] );
tran (\sa_snapshot[3][44] , \sa_snapshot[3].r.part1[12] );
tran (\sa_snapshot[3][44] , \sa_snapshot[3].f.upper[12] );
tran (\sa_snapshot[3][45] , \sa_snapshot[3].r.part1[13] );
tran (\sa_snapshot[3][45] , \sa_snapshot[3].f.upper[13] );
tran (\sa_snapshot[3][46] , \sa_snapshot[3].r.part1[14] );
tran (\sa_snapshot[3][46] , \sa_snapshot[3].f.upper[14] );
tran (\sa_snapshot[3][47] , \sa_snapshot[3].r.part1[15] );
tran (\sa_snapshot[3][47] , \sa_snapshot[3].f.upper[15] );
tran (\sa_snapshot[3][48] , \sa_snapshot[3].r.part1[16] );
tran (\sa_snapshot[3][48] , \sa_snapshot[3].f.upper[16] );
tran (\sa_snapshot[3][49] , \sa_snapshot[3].r.part1[17] );
tran (\sa_snapshot[3][49] , \sa_snapshot[3].f.upper[17] );
tran (\sa_snapshot[3][50] , \sa_snapshot[3].r.part1[18] );
tran (\sa_snapshot[3][50] , \sa_snapshot[3].f.unused[0] );
tran (\sa_snapshot[3][51] , \sa_snapshot[3].r.part1[19] );
tran (\sa_snapshot[3][51] , \sa_snapshot[3].f.unused[1] );
tran (\sa_snapshot[3][52] , \sa_snapshot[3].r.part1[20] );
tran (\sa_snapshot[3][52] , \sa_snapshot[3].f.unused[2] );
tran (\sa_snapshot[3][53] , \sa_snapshot[3].r.part1[21] );
tran (\sa_snapshot[3][53] , \sa_snapshot[3].f.unused[3] );
tran (\sa_snapshot[3][54] , \sa_snapshot[3].r.part1[22] );
tran (\sa_snapshot[3][54] , \sa_snapshot[3].f.unused[4] );
tran (\sa_snapshot[3][55] , \sa_snapshot[3].r.part1[23] );
tran (\sa_snapshot[3][55] , \sa_snapshot[3].f.unused[5] );
tran (\sa_snapshot[3][56] , \sa_snapshot[3].r.part1[24] );
tran (\sa_snapshot[3][56] , \sa_snapshot[3].f.unused[6] );
tran (\sa_snapshot[3][57] , \sa_snapshot[3].r.part1[25] );
tran (\sa_snapshot[3][57] , \sa_snapshot[3].f.unused[7] );
tran (\sa_snapshot[3][58] , \sa_snapshot[3].r.part1[26] );
tran (\sa_snapshot[3][58] , \sa_snapshot[3].f.unused[8] );
tran (\sa_snapshot[3][59] , \sa_snapshot[3].r.part1[27] );
tran (\sa_snapshot[3][59] , \sa_snapshot[3].f.unused[9] );
tran (\sa_snapshot[3][60] , \sa_snapshot[3].r.part1[28] );
tran (\sa_snapshot[3][60] , \sa_snapshot[3].f.unused[10] );
tran (\sa_snapshot[3][61] , \sa_snapshot[3].r.part1[29] );
tran (\sa_snapshot[3][61] , \sa_snapshot[3].f.unused[11] );
tran (\sa_snapshot[3][62] , \sa_snapshot[3].r.part1[30] );
tran (\sa_snapshot[3][62] , \sa_snapshot[3].f.unused[12] );
tran (\sa_snapshot[3][63] , \sa_snapshot[3].r.part1[31] );
tran (\sa_snapshot[3][63] , \sa_snapshot[3].f.unused[13] );
tran (\sa_snapshot[4][0] , \sa_snapshot[4].r.part0[0] );
tran (\sa_snapshot[4][0] , \sa_snapshot[4].f.lower[0] );
tran (\sa_snapshot[4][1] , \sa_snapshot[4].r.part0[1] );
tran (\sa_snapshot[4][1] , \sa_snapshot[4].f.lower[1] );
tran (\sa_snapshot[4][2] , \sa_snapshot[4].r.part0[2] );
tran (\sa_snapshot[4][2] , \sa_snapshot[4].f.lower[2] );
tran (\sa_snapshot[4][3] , \sa_snapshot[4].r.part0[3] );
tran (\sa_snapshot[4][3] , \sa_snapshot[4].f.lower[3] );
tran (\sa_snapshot[4][4] , \sa_snapshot[4].r.part0[4] );
tran (\sa_snapshot[4][4] , \sa_snapshot[4].f.lower[4] );
tran (\sa_snapshot[4][5] , \sa_snapshot[4].r.part0[5] );
tran (\sa_snapshot[4][5] , \sa_snapshot[4].f.lower[5] );
tran (\sa_snapshot[4][6] , \sa_snapshot[4].r.part0[6] );
tran (\sa_snapshot[4][6] , \sa_snapshot[4].f.lower[6] );
tran (\sa_snapshot[4][7] , \sa_snapshot[4].r.part0[7] );
tran (\sa_snapshot[4][7] , \sa_snapshot[4].f.lower[7] );
tran (\sa_snapshot[4][8] , \sa_snapshot[4].r.part0[8] );
tran (\sa_snapshot[4][8] , \sa_snapshot[4].f.lower[8] );
tran (\sa_snapshot[4][9] , \sa_snapshot[4].r.part0[9] );
tran (\sa_snapshot[4][9] , \sa_snapshot[4].f.lower[9] );
tran (\sa_snapshot[4][10] , \sa_snapshot[4].r.part0[10] );
tran (\sa_snapshot[4][10] , \sa_snapshot[4].f.lower[10] );
tran (\sa_snapshot[4][11] , \sa_snapshot[4].r.part0[11] );
tran (\sa_snapshot[4][11] , \sa_snapshot[4].f.lower[11] );
tran (\sa_snapshot[4][12] , \sa_snapshot[4].r.part0[12] );
tran (\sa_snapshot[4][12] , \sa_snapshot[4].f.lower[12] );
tran (\sa_snapshot[4][13] , \sa_snapshot[4].r.part0[13] );
tran (\sa_snapshot[4][13] , \sa_snapshot[4].f.lower[13] );
tran (\sa_snapshot[4][14] , \sa_snapshot[4].r.part0[14] );
tran (\sa_snapshot[4][14] , \sa_snapshot[4].f.lower[14] );
tran (\sa_snapshot[4][15] , \sa_snapshot[4].r.part0[15] );
tran (\sa_snapshot[4][15] , \sa_snapshot[4].f.lower[15] );
tran (\sa_snapshot[4][16] , \sa_snapshot[4].r.part0[16] );
tran (\sa_snapshot[4][16] , \sa_snapshot[4].f.lower[16] );
tran (\sa_snapshot[4][17] , \sa_snapshot[4].r.part0[17] );
tran (\sa_snapshot[4][17] , \sa_snapshot[4].f.lower[17] );
tran (\sa_snapshot[4][18] , \sa_snapshot[4].r.part0[18] );
tran (\sa_snapshot[4][18] , \sa_snapshot[4].f.lower[18] );
tran (\sa_snapshot[4][19] , \sa_snapshot[4].r.part0[19] );
tran (\sa_snapshot[4][19] , \sa_snapshot[4].f.lower[19] );
tran (\sa_snapshot[4][20] , \sa_snapshot[4].r.part0[20] );
tran (\sa_snapshot[4][20] , \sa_snapshot[4].f.lower[20] );
tran (\sa_snapshot[4][21] , \sa_snapshot[4].r.part0[21] );
tran (\sa_snapshot[4][21] , \sa_snapshot[4].f.lower[21] );
tran (\sa_snapshot[4][22] , \sa_snapshot[4].r.part0[22] );
tran (\sa_snapshot[4][22] , \sa_snapshot[4].f.lower[22] );
tran (\sa_snapshot[4][23] , \sa_snapshot[4].r.part0[23] );
tran (\sa_snapshot[4][23] , \sa_snapshot[4].f.lower[23] );
tran (\sa_snapshot[4][24] , \sa_snapshot[4].r.part0[24] );
tran (\sa_snapshot[4][24] , \sa_snapshot[4].f.lower[24] );
tran (\sa_snapshot[4][25] , \sa_snapshot[4].r.part0[25] );
tran (\sa_snapshot[4][25] , \sa_snapshot[4].f.lower[25] );
tran (\sa_snapshot[4][26] , \sa_snapshot[4].r.part0[26] );
tran (\sa_snapshot[4][26] , \sa_snapshot[4].f.lower[26] );
tran (\sa_snapshot[4][27] , \sa_snapshot[4].r.part0[27] );
tran (\sa_snapshot[4][27] , \sa_snapshot[4].f.lower[27] );
tran (\sa_snapshot[4][28] , \sa_snapshot[4].r.part0[28] );
tran (\sa_snapshot[4][28] , \sa_snapshot[4].f.lower[28] );
tran (\sa_snapshot[4][29] , \sa_snapshot[4].r.part0[29] );
tran (\sa_snapshot[4][29] , \sa_snapshot[4].f.lower[29] );
tran (\sa_snapshot[4][30] , \sa_snapshot[4].r.part0[30] );
tran (\sa_snapshot[4][30] , \sa_snapshot[4].f.lower[30] );
tran (\sa_snapshot[4][31] , \sa_snapshot[4].r.part0[31] );
tran (\sa_snapshot[4][31] , \sa_snapshot[4].f.lower[31] );
tran (\sa_snapshot[4][32] , \sa_snapshot[4].r.part1[0] );
tran (\sa_snapshot[4][32] , \sa_snapshot[4].f.upper[0] );
tran (\sa_snapshot[4][33] , \sa_snapshot[4].r.part1[1] );
tran (\sa_snapshot[4][33] , \sa_snapshot[4].f.upper[1] );
tran (\sa_snapshot[4][34] , \sa_snapshot[4].r.part1[2] );
tran (\sa_snapshot[4][34] , \sa_snapshot[4].f.upper[2] );
tran (\sa_snapshot[4][35] , \sa_snapshot[4].r.part1[3] );
tran (\sa_snapshot[4][35] , \sa_snapshot[4].f.upper[3] );
tran (\sa_snapshot[4][36] , \sa_snapshot[4].r.part1[4] );
tran (\sa_snapshot[4][36] , \sa_snapshot[4].f.upper[4] );
tran (\sa_snapshot[4][37] , \sa_snapshot[4].r.part1[5] );
tran (\sa_snapshot[4][37] , \sa_snapshot[4].f.upper[5] );
tran (\sa_snapshot[4][38] , \sa_snapshot[4].r.part1[6] );
tran (\sa_snapshot[4][38] , \sa_snapshot[4].f.upper[6] );
tran (\sa_snapshot[4][39] , \sa_snapshot[4].r.part1[7] );
tran (\sa_snapshot[4][39] , \sa_snapshot[4].f.upper[7] );
tran (\sa_snapshot[4][40] , \sa_snapshot[4].r.part1[8] );
tran (\sa_snapshot[4][40] , \sa_snapshot[4].f.upper[8] );
tran (\sa_snapshot[4][41] , \sa_snapshot[4].r.part1[9] );
tran (\sa_snapshot[4][41] , \sa_snapshot[4].f.upper[9] );
tran (\sa_snapshot[4][42] , \sa_snapshot[4].r.part1[10] );
tran (\sa_snapshot[4][42] , \sa_snapshot[4].f.upper[10] );
tran (\sa_snapshot[4][43] , \sa_snapshot[4].r.part1[11] );
tran (\sa_snapshot[4][43] , \sa_snapshot[4].f.upper[11] );
tran (\sa_snapshot[4][44] , \sa_snapshot[4].r.part1[12] );
tran (\sa_snapshot[4][44] , \sa_snapshot[4].f.upper[12] );
tran (\sa_snapshot[4][45] , \sa_snapshot[4].r.part1[13] );
tran (\sa_snapshot[4][45] , \sa_snapshot[4].f.upper[13] );
tran (\sa_snapshot[4][46] , \sa_snapshot[4].r.part1[14] );
tran (\sa_snapshot[4][46] , \sa_snapshot[4].f.upper[14] );
tran (\sa_snapshot[4][47] , \sa_snapshot[4].r.part1[15] );
tran (\sa_snapshot[4][47] , \sa_snapshot[4].f.upper[15] );
tran (\sa_snapshot[4][48] , \sa_snapshot[4].r.part1[16] );
tran (\sa_snapshot[4][48] , \sa_snapshot[4].f.upper[16] );
tran (\sa_snapshot[4][49] , \sa_snapshot[4].r.part1[17] );
tran (\sa_snapshot[4][49] , \sa_snapshot[4].f.upper[17] );
tran (\sa_snapshot[4][50] , \sa_snapshot[4].r.part1[18] );
tran (\sa_snapshot[4][50] , \sa_snapshot[4].f.unused[0] );
tran (\sa_snapshot[4][51] , \sa_snapshot[4].r.part1[19] );
tran (\sa_snapshot[4][51] , \sa_snapshot[4].f.unused[1] );
tran (\sa_snapshot[4][52] , \sa_snapshot[4].r.part1[20] );
tran (\sa_snapshot[4][52] , \sa_snapshot[4].f.unused[2] );
tran (\sa_snapshot[4][53] , \sa_snapshot[4].r.part1[21] );
tran (\sa_snapshot[4][53] , \sa_snapshot[4].f.unused[3] );
tran (\sa_snapshot[4][54] , \sa_snapshot[4].r.part1[22] );
tran (\sa_snapshot[4][54] , \sa_snapshot[4].f.unused[4] );
tran (\sa_snapshot[4][55] , \sa_snapshot[4].r.part1[23] );
tran (\sa_snapshot[4][55] , \sa_snapshot[4].f.unused[5] );
tran (\sa_snapshot[4][56] , \sa_snapshot[4].r.part1[24] );
tran (\sa_snapshot[4][56] , \sa_snapshot[4].f.unused[6] );
tran (\sa_snapshot[4][57] , \sa_snapshot[4].r.part1[25] );
tran (\sa_snapshot[4][57] , \sa_snapshot[4].f.unused[7] );
tran (\sa_snapshot[4][58] , \sa_snapshot[4].r.part1[26] );
tran (\sa_snapshot[4][58] , \sa_snapshot[4].f.unused[8] );
tran (\sa_snapshot[4][59] , \sa_snapshot[4].r.part1[27] );
tran (\sa_snapshot[4][59] , \sa_snapshot[4].f.unused[9] );
tran (\sa_snapshot[4][60] , \sa_snapshot[4].r.part1[28] );
tran (\sa_snapshot[4][60] , \sa_snapshot[4].f.unused[10] );
tran (\sa_snapshot[4][61] , \sa_snapshot[4].r.part1[29] );
tran (\sa_snapshot[4][61] , \sa_snapshot[4].f.unused[11] );
tran (\sa_snapshot[4][62] , \sa_snapshot[4].r.part1[30] );
tran (\sa_snapshot[4][62] , \sa_snapshot[4].f.unused[12] );
tran (\sa_snapshot[4][63] , \sa_snapshot[4].r.part1[31] );
tran (\sa_snapshot[4][63] , \sa_snapshot[4].f.unused[13] );
tran (\sa_snapshot[5][0] , \sa_snapshot[5].r.part0[0] );
tran (\sa_snapshot[5][0] , \sa_snapshot[5].f.lower[0] );
tran (\sa_snapshot[5][1] , \sa_snapshot[5].r.part0[1] );
tran (\sa_snapshot[5][1] , \sa_snapshot[5].f.lower[1] );
tran (\sa_snapshot[5][2] , \sa_snapshot[5].r.part0[2] );
tran (\sa_snapshot[5][2] , \sa_snapshot[5].f.lower[2] );
tran (\sa_snapshot[5][3] , \sa_snapshot[5].r.part0[3] );
tran (\sa_snapshot[5][3] , \sa_snapshot[5].f.lower[3] );
tran (\sa_snapshot[5][4] , \sa_snapshot[5].r.part0[4] );
tran (\sa_snapshot[5][4] , \sa_snapshot[5].f.lower[4] );
tran (\sa_snapshot[5][5] , \sa_snapshot[5].r.part0[5] );
tran (\sa_snapshot[5][5] , \sa_snapshot[5].f.lower[5] );
tran (\sa_snapshot[5][6] , \sa_snapshot[5].r.part0[6] );
tran (\sa_snapshot[5][6] , \sa_snapshot[5].f.lower[6] );
tran (\sa_snapshot[5][7] , \sa_snapshot[5].r.part0[7] );
tran (\sa_snapshot[5][7] , \sa_snapshot[5].f.lower[7] );
tran (\sa_snapshot[5][8] , \sa_snapshot[5].r.part0[8] );
tran (\sa_snapshot[5][8] , \sa_snapshot[5].f.lower[8] );
tran (\sa_snapshot[5][9] , \sa_snapshot[5].r.part0[9] );
tran (\sa_snapshot[5][9] , \sa_snapshot[5].f.lower[9] );
tran (\sa_snapshot[5][10] , \sa_snapshot[5].r.part0[10] );
tran (\sa_snapshot[5][10] , \sa_snapshot[5].f.lower[10] );
tran (\sa_snapshot[5][11] , \sa_snapshot[5].r.part0[11] );
tran (\sa_snapshot[5][11] , \sa_snapshot[5].f.lower[11] );
tran (\sa_snapshot[5][12] , \sa_snapshot[5].r.part0[12] );
tran (\sa_snapshot[5][12] , \sa_snapshot[5].f.lower[12] );
tran (\sa_snapshot[5][13] , \sa_snapshot[5].r.part0[13] );
tran (\sa_snapshot[5][13] , \sa_snapshot[5].f.lower[13] );
tran (\sa_snapshot[5][14] , \sa_snapshot[5].r.part0[14] );
tran (\sa_snapshot[5][14] , \sa_snapshot[5].f.lower[14] );
tran (\sa_snapshot[5][15] , \sa_snapshot[5].r.part0[15] );
tran (\sa_snapshot[5][15] , \sa_snapshot[5].f.lower[15] );
tran (\sa_snapshot[5][16] , \sa_snapshot[5].r.part0[16] );
tran (\sa_snapshot[5][16] , \sa_snapshot[5].f.lower[16] );
tran (\sa_snapshot[5][17] , \sa_snapshot[5].r.part0[17] );
tran (\sa_snapshot[5][17] , \sa_snapshot[5].f.lower[17] );
tran (\sa_snapshot[5][18] , \sa_snapshot[5].r.part0[18] );
tran (\sa_snapshot[5][18] , \sa_snapshot[5].f.lower[18] );
tran (\sa_snapshot[5][19] , \sa_snapshot[5].r.part0[19] );
tran (\sa_snapshot[5][19] , \sa_snapshot[5].f.lower[19] );
tran (\sa_snapshot[5][20] , \sa_snapshot[5].r.part0[20] );
tran (\sa_snapshot[5][20] , \sa_snapshot[5].f.lower[20] );
tran (\sa_snapshot[5][21] , \sa_snapshot[5].r.part0[21] );
tran (\sa_snapshot[5][21] , \sa_snapshot[5].f.lower[21] );
tran (\sa_snapshot[5][22] , \sa_snapshot[5].r.part0[22] );
tran (\sa_snapshot[5][22] , \sa_snapshot[5].f.lower[22] );
tran (\sa_snapshot[5][23] , \sa_snapshot[5].r.part0[23] );
tran (\sa_snapshot[5][23] , \sa_snapshot[5].f.lower[23] );
tran (\sa_snapshot[5][24] , \sa_snapshot[5].r.part0[24] );
tran (\sa_snapshot[5][24] , \sa_snapshot[5].f.lower[24] );
tran (\sa_snapshot[5][25] , \sa_snapshot[5].r.part0[25] );
tran (\sa_snapshot[5][25] , \sa_snapshot[5].f.lower[25] );
tran (\sa_snapshot[5][26] , \sa_snapshot[5].r.part0[26] );
tran (\sa_snapshot[5][26] , \sa_snapshot[5].f.lower[26] );
tran (\sa_snapshot[5][27] , \sa_snapshot[5].r.part0[27] );
tran (\sa_snapshot[5][27] , \sa_snapshot[5].f.lower[27] );
tran (\sa_snapshot[5][28] , \sa_snapshot[5].r.part0[28] );
tran (\sa_snapshot[5][28] , \sa_snapshot[5].f.lower[28] );
tran (\sa_snapshot[5][29] , \sa_snapshot[5].r.part0[29] );
tran (\sa_snapshot[5][29] , \sa_snapshot[5].f.lower[29] );
tran (\sa_snapshot[5][30] , \sa_snapshot[5].r.part0[30] );
tran (\sa_snapshot[5][30] , \sa_snapshot[5].f.lower[30] );
tran (\sa_snapshot[5][31] , \sa_snapshot[5].r.part0[31] );
tran (\sa_snapshot[5][31] , \sa_snapshot[5].f.lower[31] );
tran (\sa_snapshot[5][32] , \sa_snapshot[5].r.part1[0] );
tran (\sa_snapshot[5][32] , \sa_snapshot[5].f.upper[0] );
tran (\sa_snapshot[5][33] , \sa_snapshot[5].r.part1[1] );
tran (\sa_snapshot[5][33] , \sa_snapshot[5].f.upper[1] );
tran (\sa_snapshot[5][34] , \sa_snapshot[5].r.part1[2] );
tran (\sa_snapshot[5][34] , \sa_snapshot[5].f.upper[2] );
tran (\sa_snapshot[5][35] , \sa_snapshot[5].r.part1[3] );
tran (\sa_snapshot[5][35] , \sa_snapshot[5].f.upper[3] );
tran (\sa_snapshot[5][36] , \sa_snapshot[5].r.part1[4] );
tran (\sa_snapshot[5][36] , \sa_snapshot[5].f.upper[4] );
tran (\sa_snapshot[5][37] , \sa_snapshot[5].r.part1[5] );
tran (\sa_snapshot[5][37] , \sa_snapshot[5].f.upper[5] );
tran (\sa_snapshot[5][38] , \sa_snapshot[5].r.part1[6] );
tran (\sa_snapshot[5][38] , \sa_snapshot[5].f.upper[6] );
tran (\sa_snapshot[5][39] , \sa_snapshot[5].r.part1[7] );
tran (\sa_snapshot[5][39] , \sa_snapshot[5].f.upper[7] );
tran (\sa_snapshot[5][40] , \sa_snapshot[5].r.part1[8] );
tran (\sa_snapshot[5][40] , \sa_snapshot[5].f.upper[8] );
tran (\sa_snapshot[5][41] , \sa_snapshot[5].r.part1[9] );
tran (\sa_snapshot[5][41] , \sa_snapshot[5].f.upper[9] );
tran (\sa_snapshot[5][42] , \sa_snapshot[5].r.part1[10] );
tran (\sa_snapshot[5][42] , \sa_snapshot[5].f.upper[10] );
tran (\sa_snapshot[5][43] , \sa_snapshot[5].r.part1[11] );
tran (\sa_snapshot[5][43] , \sa_snapshot[5].f.upper[11] );
tran (\sa_snapshot[5][44] , \sa_snapshot[5].r.part1[12] );
tran (\sa_snapshot[5][44] , \sa_snapshot[5].f.upper[12] );
tran (\sa_snapshot[5][45] , \sa_snapshot[5].r.part1[13] );
tran (\sa_snapshot[5][45] , \sa_snapshot[5].f.upper[13] );
tran (\sa_snapshot[5][46] , \sa_snapshot[5].r.part1[14] );
tran (\sa_snapshot[5][46] , \sa_snapshot[5].f.upper[14] );
tran (\sa_snapshot[5][47] , \sa_snapshot[5].r.part1[15] );
tran (\sa_snapshot[5][47] , \sa_snapshot[5].f.upper[15] );
tran (\sa_snapshot[5][48] , \sa_snapshot[5].r.part1[16] );
tran (\sa_snapshot[5][48] , \sa_snapshot[5].f.upper[16] );
tran (\sa_snapshot[5][49] , \sa_snapshot[5].r.part1[17] );
tran (\sa_snapshot[5][49] , \sa_snapshot[5].f.upper[17] );
tran (\sa_snapshot[5][50] , \sa_snapshot[5].r.part1[18] );
tran (\sa_snapshot[5][50] , \sa_snapshot[5].f.unused[0] );
tran (\sa_snapshot[5][51] , \sa_snapshot[5].r.part1[19] );
tran (\sa_snapshot[5][51] , \sa_snapshot[5].f.unused[1] );
tran (\sa_snapshot[5][52] , \sa_snapshot[5].r.part1[20] );
tran (\sa_snapshot[5][52] , \sa_snapshot[5].f.unused[2] );
tran (\sa_snapshot[5][53] , \sa_snapshot[5].r.part1[21] );
tran (\sa_snapshot[5][53] , \sa_snapshot[5].f.unused[3] );
tran (\sa_snapshot[5][54] , \sa_snapshot[5].r.part1[22] );
tran (\sa_snapshot[5][54] , \sa_snapshot[5].f.unused[4] );
tran (\sa_snapshot[5][55] , \sa_snapshot[5].r.part1[23] );
tran (\sa_snapshot[5][55] , \sa_snapshot[5].f.unused[5] );
tran (\sa_snapshot[5][56] , \sa_snapshot[5].r.part1[24] );
tran (\sa_snapshot[5][56] , \sa_snapshot[5].f.unused[6] );
tran (\sa_snapshot[5][57] , \sa_snapshot[5].r.part1[25] );
tran (\sa_snapshot[5][57] , \sa_snapshot[5].f.unused[7] );
tran (\sa_snapshot[5][58] , \sa_snapshot[5].r.part1[26] );
tran (\sa_snapshot[5][58] , \sa_snapshot[5].f.unused[8] );
tran (\sa_snapshot[5][59] , \sa_snapshot[5].r.part1[27] );
tran (\sa_snapshot[5][59] , \sa_snapshot[5].f.unused[9] );
tran (\sa_snapshot[5][60] , \sa_snapshot[5].r.part1[28] );
tran (\sa_snapshot[5][60] , \sa_snapshot[5].f.unused[10] );
tran (\sa_snapshot[5][61] , \sa_snapshot[5].r.part1[29] );
tran (\sa_snapshot[5][61] , \sa_snapshot[5].f.unused[11] );
tran (\sa_snapshot[5][62] , \sa_snapshot[5].r.part1[30] );
tran (\sa_snapshot[5][62] , \sa_snapshot[5].f.unused[12] );
tran (\sa_snapshot[5][63] , \sa_snapshot[5].r.part1[31] );
tran (\sa_snapshot[5][63] , \sa_snapshot[5].f.unused[13] );
tran (\sa_snapshot[6][0] , \sa_snapshot[6].r.part0[0] );
tran (\sa_snapshot[6][0] , \sa_snapshot[6].f.lower[0] );
tran (\sa_snapshot[6][1] , \sa_snapshot[6].r.part0[1] );
tran (\sa_snapshot[6][1] , \sa_snapshot[6].f.lower[1] );
tran (\sa_snapshot[6][2] , \sa_snapshot[6].r.part0[2] );
tran (\sa_snapshot[6][2] , \sa_snapshot[6].f.lower[2] );
tran (\sa_snapshot[6][3] , \sa_snapshot[6].r.part0[3] );
tran (\sa_snapshot[6][3] , \sa_snapshot[6].f.lower[3] );
tran (\sa_snapshot[6][4] , \sa_snapshot[6].r.part0[4] );
tran (\sa_snapshot[6][4] , \sa_snapshot[6].f.lower[4] );
tran (\sa_snapshot[6][5] , \sa_snapshot[6].r.part0[5] );
tran (\sa_snapshot[6][5] , \sa_snapshot[6].f.lower[5] );
tran (\sa_snapshot[6][6] , \sa_snapshot[6].r.part0[6] );
tran (\sa_snapshot[6][6] , \sa_snapshot[6].f.lower[6] );
tran (\sa_snapshot[6][7] , \sa_snapshot[6].r.part0[7] );
tran (\sa_snapshot[6][7] , \sa_snapshot[6].f.lower[7] );
tran (\sa_snapshot[6][8] , \sa_snapshot[6].r.part0[8] );
tran (\sa_snapshot[6][8] , \sa_snapshot[6].f.lower[8] );
tran (\sa_snapshot[6][9] , \sa_snapshot[6].r.part0[9] );
tran (\sa_snapshot[6][9] , \sa_snapshot[6].f.lower[9] );
tran (\sa_snapshot[6][10] , \sa_snapshot[6].r.part0[10] );
tran (\sa_snapshot[6][10] , \sa_snapshot[6].f.lower[10] );
tran (\sa_snapshot[6][11] , \sa_snapshot[6].r.part0[11] );
tran (\sa_snapshot[6][11] , \sa_snapshot[6].f.lower[11] );
tran (\sa_snapshot[6][12] , \sa_snapshot[6].r.part0[12] );
tran (\sa_snapshot[6][12] , \sa_snapshot[6].f.lower[12] );
tran (\sa_snapshot[6][13] , \sa_snapshot[6].r.part0[13] );
tran (\sa_snapshot[6][13] , \sa_snapshot[6].f.lower[13] );
tran (\sa_snapshot[6][14] , \sa_snapshot[6].r.part0[14] );
tran (\sa_snapshot[6][14] , \sa_snapshot[6].f.lower[14] );
tran (\sa_snapshot[6][15] , \sa_snapshot[6].r.part0[15] );
tran (\sa_snapshot[6][15] , \sa_snapshot[6].f.lower[15] );
tran (\sa_snapshot[6][16] , \sa_snapshot[6].r.part0[16] );
tran (\sa_snapshot[6][16] , \sa_snapshot[6].f.lower[16] );
tran (\sa_snapshot[6][17] , \sa_snapshot[6].r.part0[17] );
tran (\sa_snapshot[6][17] , \sa_snapshot[6].f.lower[17] );
tran (\sa_snapshot[6][18] , \sa_snapshot[6].r.part0[18] );
tran (\sa_snapshot[6][18] , \sa_snapshot[6].f.lower[18] );
tran (\sa_snapshot[6][19] , \sa_snapshot[6].r.part0[19] );
tran (\sa_snapshot[6][19] , \sa_snapshot[6].f.lower[19] );
tran (\sa_snapshot[6][20] , \sa_snapshot[6].r.part0[20] );
tran (\sa_snapshot[6][20] , \sa_snapshot[6].f.lower[20] );
tran (\sa_snapshot[6][21] , \sa_snapshot[6].r.part0[21] );
tran (\sa_snapshot[6][21] , \sa_snapshot[6].f.lower[21] );
tran (\sa_snapshot[6][22] , \sa_snapshot[6].r.part0[22] );
tran (\sa_snapshot[6][22] , \sa_snapshot[6].f.lower[22] );
tran (\sa_snapshot[6][23] , \sa_snapshot[6].r.part0[23] );
tran (\sa_snapshot[6][23] , \sa_snapshot[6].f.lower[23] );
tran (\sa_snapshot[6][24] , \sa_snapshot[6].r.part0[24] );
tran (\sa_snapshot[6][24] , \sa_snapshot[6].f.lower[24] );
tran (\sa_snapshot[6][25] , \sa_snapshot[6].r.part0[25] );
tran (\sa_snapshot[6][25] , \sa_snapshot[6].f.lower[25] );
tran (\sa_snapshot[6][26] , \sa_snapshot[6].r.part0[26] );
tran (\sa_snapshot[6][26] , \sa_snapshot[6].f.lower[26] );
tran (\sa_snapshot[6][27] , \sa_snapshot[6].r.part0[27] );
tran (\sa_snapshot[6][27] , \sa_snapshot[6].f.lower[27] );
tran (\sa_snapshot[6][28] , \sa_snapshot[6].r.part0[28] );
tran (\sa_snapshot[6][28] , \sa_snapshot[6].f.lower[28] );
tran (\sa_snapshot[6][29] , \sa_snapshot[6].r.part0[29] );
tran (\sa_snapshot[6][29] , \sa_snapshot[6].f.lower[29] );
tran (\sa_snapshot[6][30] , \sa_snapshot[6].r.part0[30] );
tran (\sa_snapshot[6][30] , \sa_snapshot[6].f.lower[30] );
tran (\sa_snapshot[6][31] , \sa_snapshot[6].r.part0[31] );
tran (\sa_snapshot[6][31] , \sa_snapshot[6].f.lower[31] );
tran (\sa_snapshot[6][32] , \sa_snapshot[6].r.part1[0] );
tran (\sa_snapshot[6][32] , \sa_snapshot[6].f.upper[0] );
tran (\sa_snapshot[6][33] , \sa_snapshot[6].r.part1[1] );
tran (\sa_snapshot[6][33] , \sa_snapshot[6].f.upper[1] );
tran (\sa_snapshot[6][34] , \sa_snapshot[6].r.part1[2] );
tran (\sa_snapshot[6][34] , \sa_snapshot[6].f.upper[2] );
tran (\sa_snapshot[6][35] , \sa_snapshot[6].r.part1[3] );
tran (\sa_snapshot[6][35] , \sa_snapshot[6].f.upper[3] );
tran (\sa_snapshot[6][36] , \sa_snapshot[6].r.part1[4] );
tran (\sa_snapshot[6][36] , \sa_snapshot[6].f.upper[4] );
tran (\sa_snapshot[6][37] , \sa_snapshot[6].r.part1[5] );
tran (\sa_snapshot[6][37] , \sa_snapshot[6].f.upper[5] );
tran (\sa_snapshot[6][38] , \sa_snapshot[6].r.part1[6] );
tran (\sa_snapshot[6][38] , \sa_snapshot[6].f.upper[6] );
tran (\sa_snapshot[6][39] , \sa_snapshot[6].r.part1[7] );
tran (\sa_snapshot[6][39] , \sa_snapshot[6].f.upper[7] );
tran (\sa_snapshot[6][40] , \sa_snapshot[6].r.part1[8] );
tran (\sa_snapshot[6][40] , \sa_snapshot[6].f.upper[8] );
tran (\sa_snapshot[6][41] , \sa_snapshot[6].r.part1[9] );
tran (\sa_snapshot[6][41] , \sa_snapshot[6].f.upper[9] );
tran (\sa_snapshot[6][42] , \sa_snapshot[6].r.part1[10] );
tran (\sa_snapshot[6][42] , \sa_snapshot[6].f.upper[10] );
tran (\sa_snapshot[6][43] , \sa_snapshot[6].r.part1[11] );
tran (\sa_snapshot[6][43] , \sa_snapshot[6].f.upper[11] );
tran (\sa_snapshot[6][44] , \sa_snapshot[6].r.part1[12] );
tran (\sa_snapshot[6][44] , \sa_snapshot[6].f.upper[12] );
tran (\sa_snapshot[6][45] , \sa_snapshot[6].r.part1[13] );
tran (\sa_snapshot[6][45] , \sa_snapshot[6].f.upper[13] );
tran (\sa_snapshot[6][46] , \sa_snapshot[6].r.part1[14] );
tran (\sa_snapshot[6][46] , \sa_snapshot[6].f.upper[14] );
tran (\sa_snapshot[6][47] , \sa_snapshot[6].r.part1[15] );
tran (\sa_snapshot[6][47] , \sa_snapshot[6].f.upper[15] );
tran (\sa_snapshot[6][48] , \sa_snapshot[6].r.part1[16] );
tran (\sa_snapshot[6][48] , \sa_snapshot[6].f.upper[16] );
tran (\sa_snapshot[6][49] , \sa_snapshot[6].r.part1[17] );
tran (\sa_snapshot[6][49] , \sa_snapshot[6].f.upper[17] );
tran (\sa_snapshot[6][50] , \sa_snapshot[6].r.part1[18] );
tran (\sa_snapshot[6][50] , \sa_snapshot[6].f.unused[0] );
tran (\sa_snapshot[6][51] , \sa_snapshot[6].r.part1[19] );
tran (\sa_snapshot[6][51] , \sa_snapshot[6].f.unused[1] );
tran (\sa_snapshot[6][52] , \sa_snapshot[6].r.part1[20] );
tran (\sa_snapshot[6][52] , \sa_snapshot[6].f.unused[2] );
tran (\sa_snapshot[6][53] , \sa_snapshot[6].r.part1[21] );
tran (\sa_snapshot[6][53] , \sa_snapshot[6].f.unused[3] );
tran (\sa_snapshot[6][54] , \sa_snapshot[6].r.part1[22] );
tran (\sa_snapshot[6][54] , \sa_snapshot[6].f.unused[4] );
tran (\sa_snapshot[6][55] , \sa_snapshot[6].r.part1[23] );
tran (\sa_snapshot[6][55] , \sa_snapshot[6].f.unused[5] );
tran (\sa_snapshot[6][56] , \sa_snapshot[6].r.part1[24] );
tran (\sa_snapshot[6][56] , \sa_snapshot[6].f.unused[6] );
tran (\sa_snapshot[6][57] , \sa_snapshot[6].r.part1[25] );
tran (\sa_snapshot[6][57] , \sa_snapshot[6].f.unused[7] );
tran (\sa_snapshot[6][58] , \sa_snapshot[6].r.part1[26] );
tran (\sa_snapshot[6][58] , \sa_snapshot[6].f.unused[8] );
tran (\sa_snapshot[6][59] , \sa_snapshot[6].r.part1[27] );
tran (\sa_snapshot[6][59] , \sa_snapshot[6].f.unused[9] );
tran (\sa_snapshot[6][60] , \sa_snapshot[6].r.part1[28] );
tran (\sa_snapshot[6][60] , \sa_snapshot[6].f.unused[10] );
tran (\sa_snapshot[6][61] , \sa_snapshot[6].r.part1[29] );
tran (\sa_snapshot[6][61] , \sa_snapshot[6].f.unused[11] );
tran (\sa_snapshot[6][62] , \sa_snapshot[6].r.part1[30] );
tran (\sa_snapshot[6][62] , \sa_snapshot[6].f.unused[12] );
tran (\sa_snapshot[6][63] , \sa_snapshot[6].r.part1[31] );
tran (\sa_snapshot[6][63] , \sa_snapshot[6].f.unused[13] );
tran (\sa_snapshot[7][0] , \sa_snapshot[7].r.part0[0] );
tran (\sa_snapshot[7][0] , \sa_snapshot[7].f.lower[0] );
tran (\sa_snapshot[7][1] , \sa_snapshot[7].r.part0[1] );
tran (\sa_snapshot[7][1] , \sa_snapshot[7].f.lower[1] );
tran (\sa_snapshot[7][2] , \sa_snapshot[7].r.part0[2] );
tran (\sa_snapshot[7][2] , \sa_snapshot[7].f.lower[2] );
tran (\sa_snapshot[7][3] , \sa_snapshot[7].r.part0[3] );
tran (\sa_snapshot[7][3] , \sa_snapshot[7].f.lower[3] );
tran (\sa_snapshot[7][4] , \sa_snapshot[7].r.part0[4] );
tran (\sa_snapshot[7][4] , \sa_snapshot[7].f.lower[4] );
tran (\sa_snapshot[7][5] , \sa_snapshot[7].r.part0[5] );
tran (\sa_snapshot[7][5] , \sa_snapshot[7].f.lower[5] );
tran (\sa_snapshot[7][6] , \sa_snapshot[7].r.part0[6] );
tran (\sa_snapshot[7][6] , \sa_snapshot[7].f.lower[6] );
tran (\sa_snapshot[7][7] , \sa_snapshot[7].r.part0[7] );
tran (\sa_snapshot[7][7] , \sa_snapshot[7].f.lower[7] );
tran (\sa_snapshot[7][8] , \sa_snapshot[7].r.part0[8] );
tran (\sa_snapshot[7][8] , \sa_snapshot[7].f.lower[8] );
tran (\sa_snapshot[7][9] , \sa_snapshot[7].r.part0[9] );
tran (\sa_snapshot[7][9] , \sa_snapshot[7].f.lower[9] );
tran (\sa_snapshot[7][10] , \sa_snapshot[7].r.part0[10] );
tran (\sa_snapshot[7][10] , \sa_snapshot[7].f.lower[10] );
tran (\sa_snapshot[7][11] , \sa_snapshot[7].r.part0[11] );
tran (\sa_snapshot[7][11] , \sa_snapshot[7].f.lower[11] );
tran (\sa_snapshot[7][12] , \sa_snapshot[7].r.part0[12] );
tran (\sa_snapshot[7][12] , \sa_snapshot[7].f.lower[12] );
tran (\sa_snapshot[7][13] , \sa_snapshot[7].r.part0[13] );
tran (\sa_snapshot[7][13] , \sa_snapshot[7].f.lower[13] );
tran (\sa_snapshot[7][14] , \sa_snapshot[7].r.part0[14] );
tran (\sa_snapshot[7][14] , \sa_snapshot[7].f.lower[14] );
tran (\sa_snapshot[7][15] , \sa_snapshot[7].r.part0[15] );
tran (\sa_snapshot[7][15] , \sa_snapshot[7].f.lower[15] );
tran (\sa_snapshot[7][16] , \sa_snapshot[7].r.part0[16] );
tran (\sa_snapshot[7][16] , \sa_snapshot[7].f.lower[16] );
tran (\sa_snapshot[7][17] , \sa_snapshot[7].r.part0[17] );
tran (\sa_snapshot[7][17] , \sa_snapshot[7].f.lower[17] );
tran (\sa_snapshot[7][18] , \sa_snapshot[7].r.part0[18] );
tran (\sa_snapshot[7][18] , \sa_snapshot[7].f.lower[18] );
tran (\sa_snapshot[7][19] , \sa_snapshot[7].r.part0[19] );
tran (\sa_snapshot[7][19] , \sa_snapshot[7].f.lower[19] );
tran (\sa_snapshot[7][20] , \sa_snapshot[7].r.part0[20] );
tran (\sa_snapshot[7][20] , \sa_snapshot[7].f.lower[20] );
tran (\sa_snapshot[7][21] , \sa_snapshot[7].r.part0[21] );
tran (\sa_snapshot[7][21] , \sa_snapshot[7].f.lower[21] );
tran (\sa_snapshot[7][22] , \sa_snapshot[7].r.part0[22] );
tran (\sa_snapshot[7][22] , \sa_snapshot[7].f.lower[22] );
tran (\sa_snapshot[7][23] , \sa_snapshot[7].r.part0[23] );
tran (\sa_snapshot[7][23] , \sa_snapshot[7].f.lower[23] );
tran (\sa_snapshot[7][24] , \sa_snapshot[7].r.part0[24] );
tran (\sa_snapshot[7][24] , \sa_snapshot[7].f.lower[24] );
tran (\sa_snapshot[7][25] , \sa_snapshot[7].r.part0[25] );
tran (\sa_snapshot[7][25] , \sa_snapshot[7].f.lower[25] );
tran (\sa_snapshot[7][26] , \sa_snapshot[7].r.part0[26] );
tran (\sa_snapshot[7][26] , \sa_snapshot[7].f.lower[26] );
tran (\sa_snapshot[7][27] , \sa_snapshot[7].r.part0[27] );
tran (\sa_snapshot[7][27] , \sa_snapshot[7].f.lower[27] );
tran (\sa_snapshot[7][28] , \sa_snapshot[7].r.part0[28] );
tran (\sa_snapshot[7][28] , \sa_snapshot[7].f.lower[28] );
tran (\sa_snapshot[7][29] , \sa_snapshot[7].r.part0[29] );
tran (\sa_snapshot[7][29] , \sa_snapshot[7].f.lower[29] );
tran (\sa_snapshot[7][30] , \sa_snapshot[7].r.part0[30] );
tran (\sa_snapshot[7][30] , \sa_snapshot[7].f.lower[30] );
tran (\sa_snapshot[7][31] , \sa_snapshot[7].r.part0[31] );
tran (\sa_snapshot[7][31] , \sa_snapshot[7].f.lower[31] );
tran (\sa_snapshot[7][32] , \sa_snapshot[7].r.part1[0] );
tran (\sa_snapshot[7][32] , \sa_snapshot[7].f.upper[0] );
tran (\sa_snapshot[7][33] , \sa_snapshot[7].r.part1[1] );
tran (\sa_snapshot[7][33] , \sa_snapshot[7].f.upper[1] );
tran (\sa_snapshot[7][34] , \sa_snapshot[7].r.part1[2] );
tran (\sa_snapshot[7][34] , \sa_snapshot[7].f.upper[2] );
tran (\sa_snapshot[7][35] , \sa_snapshot[7].r.part1[3] );
tran (\sa_snapshot[7][35] , \sa_snapshot[7].f.upper[3] );
tran (\sa_snapshot[7][36] , \sa_snapshot[7].r.part1[4] );
tran (\sa_snapshot[7][36] , \sa_snapshot[7].f.upper[4] );
tran (\sa_snapshot[7][37] , \sa_snapshot[7].r.part1[5] );
tran (\sa_snapshot[7][37] , \sa_snapshot[7].f.upper[5] );
tran (\sa_snapshot[7][38] , \sa_snapshot[7].r.part1[6] );
tran (\sa_snapshot[7][38] , \sa_snapshot[7].f.upper[6] );
tran (\sa_snapshot[7][39] , \sa_snapshot[7].r.part1[7] );
tran (\sa_snapshot[7][39] , \sa_snapshot[7].f.upper[7] );
tran (\sa_snapshot[7][40] , \sa_snapshot[7].r.part1[8] );
tran (\sa_snapshot[7][40] , \sa_snapshot[7].f.upper[8] );
tran (\sa_snapshot[7][41] , \sa_snapshot[7].r.part1[9] );
tran (\sa_snapshot[7][41] , \sa_snapshot[7].f.upper[9] );
tran (\sa_snapshot[7][42] , \sa_snapshot[7].r.part1[10] );
tran (\sa_snapshot[7][42] , \sa_snapshot[7].f.upper[10] );
tran (\sa_snapshot[7][43] , \sa_snapshot[7].r.part1[11] );
tran (\sa_snapshot[7][43] , \sa_snapshot[7].f.upper[11] );
tran (\sa_snapshot[7][44] , \sa_snapshot[7].r.part1[12] );
tran (\sa_snapshot[7][44] , \sa_snapshot[7].f.upper[12] );
tran (\sa_snapshot[7][45] , \sa_snapshot[7].r.part1[13] );
tran (\sa_snapshot[7][45] , \sa_snapshot[7].f.upper[13] );
tran (\sa_snapshot[7][46] , \sa_snapshot[7].r.part1[14] );
tran (\sa_snapshot[7][46] , \sa_snapshot[7].f.upper[14] );
tran (\sa_snapshot[7][47] , \sa_snapshot[7].r.part1[15] );
tran (\sa_snapshot[7][47] , \sa_snapshot[7].f.upper[15] );
tran (\sa_snapshot[7][48] , \sa_snapshot[7].r.part1[16] );
tran (\sa_snapshot[7][48] , \sa_snapshot[7].f.upper[16] );
tran (\sa_snapshot[7][49] , \sa_snapshot[7].r.part1[17] );
tran (\sa_snapshot[7][49] , \sa_snapshot[7].f.upper[17] );
tran (\sa_snapshot[7][50] , \sa_snapshot[7].r.part1[18] );
tran (\sa_snapshot[7][50] , \sa_snapshot[7].f.unused[0] );
tran (\sa_snapshot[7][51] , \sa_snapshot[7].r.part1[19] );
tran (\sa_snapshot[7][51] , \sa_snapshot[7].f.unused[1] );
tran (\sa_snapshot[7][52] , \sa_snapshot[7].r.part1[20] );
tran (\sa_snapshot[7][52] , \sa_snapshot[7].f.unused[2] );
tran (\sa_snapshot[7][53] , \sa_snapshot[7].r.part1[21] );
tran (\sa_snapshot[7][53] , \sa_snapshot[7].f.unused[3] );
tran (\sa_snapshot[7][54] , \sa_snapshot[7].r.part1[22] );
tran (\sa_snapshot[7][54] , \sa_snapshot[7].f.unused[4] );
tran (\sa_snapshot[7][55] , \sa_snapshot[7].r.part1[23] );
tran (\sa_snapshot[7][55] , \sa_snapshot[7].f.unused[5] );
tran (\sa_snapshot[7][56] , \sa_snapshot[7].r.part1[24] );
tran (\sa_snapshot[7][56] , \sa_snapshot[7].f.unused[6] );
tran (\sa_snapshot[7][57] , \sa_snapshot[7].r.part1[25] );
tran (\sa_snapshot[7][57] , \sa_snapshot[7].f.unused[7] );
tran (\sa_snapshot[7][58] , \sa_snapshot[7].r.part1[26] );
tran (\sa_snapshot[7][58] , \sa_snapshot[7].f.unused[8] );
tran (\sa_snapshot[7][59] , \sa_snapshot[7].r.part1[27] );
tran (\sa_snapshot[7][59] , \sa_snapshot[7].f.unused[9] );
tran (\sa_snapshot[7][60] , \sa_snapshot[7].r.part1[28] );
tran (\sa_snapshot[7][60] , \sa_snapshot[7].f.unused[10] );
tran (\sa_snapshot[7][61] , \sa_snapshot[7].r.part1[29] );
tran (\sa_snapshot[7][61] , \sa_snapshot[7].f.unused[11] );
tran (\sa_snapshot[7][62] , \sa_snapshot[7].r.part1[30] );
tran (\sa_snapshot[7][62] , \sa_snapshot[7].f.unused[12] );
tran (\sa_snapshot[7][63] , \sa_snapshot[7].r.part1[31] );
tran (\sa_snapshot[7][63] , \sa_snapshot[7].f.unused[13] );
tran (\sa_snapshot[8][0] , \sa_snapshot[8].r.part0[0] );
tran (\sa_snapshot[8][0] , \sa_snapshot[8].f.lower[0] );
tran (\sa_snapshot[8][1] , \sa_snapshot[8].r.part0[1] );
tran (\sa_snapshot[8][1] , \sa_snapshot[8].f.lower[1] );
tran (\sa_snapshot[8][2] , \sa_snapshot[8].r.part0[2] );
tran (\sa_snapshot[8][2] , \sa_snapshot[8].f.lower[2] );
tran (\sa_snapshot[8][3] , \sa_snapshot[8].r.part0[3] );
tran (\sa_snapshot[8][3] , \sa_snapshot[8].f.lower[3] );
tran (\sa_snapshot[8][4] , \sa_snapshot[8].r.part0[4] );
tran (\sa_snapshot[8][4] , \sa_snapshot[8].f.lower[4] );
tran (\sa_snapshot[8][5] , \sa_snapshot[8].r.part0[5] );
tran (\sa_snapshot[8][5] , \sa_snapshot[8].f.lower[5] );
tran (\sa_snapshot[8][6] , \sa_snapshot[8].r.part0[6] );
tran (\sa_snapshot[8][6] , \sa_snapshot[8].f.lower[6] );
tran (\sa_snapshot[8][7] , \sa_snapshot[8].r.part0[7] );
tran (\sa_snapshot[8][7] , \sa_snapshot[8].f.lower[7] );
tran (\sa_snapshot[8][8] , \sa_snapshot[8].r.part0[8] );
tran (\sa_snapshot[8][8] , \sa_snapshot[8].f.lower[8] );
tran (\sa_snapshot[8][9] , \sa_snapshot[8].r.part0[9] );
tran (\sa_snapshot[8][9] , \sa_snapshot[8].f.lower[9] );
tran (\sa_snapshot[8][10] , \sa_snapshot[8].r.part0[10] );
tran (\sa_snapshot[8][10] , \sa_snapshot[8].f.lower[10] );
tran (\sa_snapshot[8][11] , \sa_snapshot[8].r.part0[11] );
tran (\sa_snapshot[8][11] , \sa_snapshot[8].f.lower[11] );
tran (\sa_snapshot[8][12] , \sa_snapshot[8].r.part0[12] );
tran (\sa_snapshot[8][12] , \sa_snapshot[8].f.lower[12] );
tran (\sa_snapshot[8][13] , \sa_snapshot[8].r.part0[13] );
tran (\sa_snapshot[8][13] , \sa_snapshot[8].f.lower[13] );
tran (\sa_snapshot[8][14] , \sa_snapshot[8].r.part0[14] );
tran (\sa_snapshot[8][14] , \sa_snapshot[8].f.lower[14] );
tran (\sa_snapshot[8][15] , \sa_snapshot[8].r.part0[15] );
tran (\sa_snapshot[8][15] , \sa_snapshot[8].f.lower[15] );
tran (\sa_snapshot[8][16] , \sa_snapshot[8].r.part0[16] );
tran (\sa_snapshot[8][16] , \sa_snapshot[8].f.lower[16] );
tran (\sa_snapshot[8][17] , \sa_snapshot[8].r.part0[17] );
tran (\sa_snapshot[8][17] , \sa_snapshot[8].f.lower[17] );
tran (\sa_snapshot[8][18] , \sa_snapshot[8].r.part0[18] );
tran (\sa_snapshot[8][18] , \sa_snapshot[8].f.lower[18] );
tran (\sa_snapshot[8][19] , \sa_snapshot[8].r.part0[19] );
tran (\sa_snapshot[8][19] , \sa_snapshot[8].f.lower[19] );
tran (\sa_snapshot[8][20] , \sa_snapshot[8].r.part0[20] );
tran (\sa_snapshot[8][20] , \sa_snapshot[8].f.lower[20] );
tran (\sa_snapshot[8][21] , \sa_snapshot[8].r.part0[21] );
tran (\sa_snapshot[8][21] , \sa_snapshot[8].f.lower[21] );
tran (\sa_snapshot[8][22] , \sa_snapshot[8].r.part0[22] );
tran (\sa_snapshot[8][22] , \sa_snapshot[8].f.lower[22] );
tran (\sa_snapshot[8][23] , \sa_snapshot[8].r.part0[23] );
tran (\sa_snapshot[8][23] , \sa_snapshot[8].f.lower[23] );
tran (\sa_snapshot[8][24] , \sa_snapshot[8].r.part0[24] );
tran (\sa_snapshot[8][24] , \sa_snapshot[8].f.lower[24] );
tran (\sa_snapshot[8][25] , \sa_snapshot[8].r.part0[25] );
tran (\sa_snapshot[8][25] , \sa_snapshot[8].f.lower[25] );
tran (\sa_snapshot[8][26] , \sa_snapshot[8].r.part0[26] );
tran (\sa_snapshot[8][26] , \sa_snapshot[8].f.lower[26] );
tran (\sa_snapshot[8][27] , \sa_snapshot[8].r.part0[27] );
tran (\sa_snapshot[8][27] , \sa_snapshot[8].f.lower[27] );
tran (\sa_snapshot[8][28] , \sa_snapshot[8].r.part0[28] );
tran (\sa_snapshot[8][28] , \sa_snapshot[8].f.lower[28] );
tran (\sa_snapshot[8][29] , \sa_snapshot[8].r.part0[29] );
tran (\sa_snapshot[8][29] , \sa_snapshot[8].f.lower[29] );
tran (\sa_snapshot[8][30] , \sa_snapshot[8].r.part0[30] );
tran (\sa_snapshot[8][30] , \sa_snapshot[8].f.lower[30] );
tran (\sa_snapshot[8][31] , \sa_snapshot[8].r.part0[31] );
tran (\sa_snapshot[8][31] , \sa_snapshot[8].f.lower[31] );
tran (\sa_snapshot[8][32] , \sa_snapshot[8].r.part1[0] );
tran (\sa_snapshot[8][32] , \sa_snapshot[8].f.upper[0] );
tran (\sa_snapshot[8][33] , \sa_snapshot[8].r.part1[1] );
tran (\sa_snapshot[8][33] , \sa_snapshot[8].f.upper[1] );
tran (\sa_snapshot[8][34] , \sa_snapshot[8].r.part1[2] );
tran (\sa_snapshot[8][34] , \sa_snapshot[8].f.upper[2] );
tran (\sa_snapshot[8][35] , \sa_snapshot[8].r.part1[3] );
tran (\sa_snapshot[8][35] , \sa_snapshot[8].f.upper[3] );
tran (\sa_snapshot[8][36] , \sa_snapshot[8].r.part1[4] );
tran (\sa_snapshot[8][36] , \sa_snapshot[8].f.upper[4] );
tran (\sa_snapshot[8][37] , \sa_snapshot[8].r.part1[5] );
tran (\sa_snapshot[8][37] , \sa_snapshot[8].f.upper[5] );
tran (\sa_snapshot[8][38] , \sa_snapshot[8].r.part1[6] );
tran (\sa_snapshot[8][38] , \sa_snapshot[8].f.upper[6] );
tran (\sa_snapshot[8][39] , \sa_snapshot[8].r.part1[7] );
tran (\sa_snapshot[8][39] , \sa_snapshot[8].f.upper[7] );
tran (\sa_snapshot[8][40] , \sa_snapshot[8].r.part1[8] );
tran (\sa_snapshot[8][40] , \sa_snapshot[8].f.upper[8] );
tran (\sa_snapshot[8][41] , \sa_snapshot[8].r.part1[9] );
tran (\sa_snapshot[8][41] , \sa_snapshot[8].f.upper[9] );
tran (\sa_snapshot[8][42] , \sa_snapshot[8].r.part1[10] );
tran (\sa_snapshot[8][42] , \sa_snapshot[8].f.upper[10] );
tran (\sa_snapshot[8][43] , \sa_snapshot[8].r.part1[11] );
tran (\sa_snapshot[8][43] , \sa_snapshot[8].f.upper[11] );
tran (\sa_snapshot[8][44] , \sa_snapshot[8].r.part1[12] );
tran (\sa_snapshot[8][44] , \sa_snapshot[8].f.upper[12] );
tran (\sa_snapshot[8][45] , \sa_snapshot[8].r.part1[13] );
tran (\sa_snapshot[8][45] , \sa_snapshot[8].f.upper[13] );
tran (\sa_snapshot[8][46] , \sa_snapshot[8].r.part1[14] );
tran (\sa_snapshot[8][46] , \sa_snapshot[8].f.upper[14] );
tran (\sa_snapshot[8][47] , \sa_snapshot[8].r.part1[15] );
tran (\sa_snapshot[8][47] , \sa_snapshot[8].f.upper[15] );
tran (\sa_snapshot[8][48] , \sa_snapshot[8].r.part1[16] );
tran (\sa_snapshot[8][48] , \sa_snapshot[8].f.upper[16] );
tran (\sa_snapshot[8][49] , \sa_snapshot[8].r.part1[17] );
tran (\sa_snapshot[8][49] , \sa_snapshot[8].f.upper[17] );
tran (\sa_snapshot[8][50] , \sa_snapshot[8].r.part1[18] );
tran (\sa_snapshot[8][50] , \sa_snapshot[8].f.unused[0] );
tran (\sa_snapshot[8][51] , \sa_snapshot[8].r.part1[19] );
tran (\sa_snapshot[8][51] , \sa_snapshot[8].f.unused[1] );
tran (\sa_snapshot[8][52] , \sa_snapshot[8].r.part1[20] );
tran (\sa_snapshot[8][52] , \sa_snapshot[8].f.unused[2] );
tran (\sa_snapshot[8][53] , \sa_snapshot[8].r.part1[21] );
tran (\sa_snapshot[8][53] , \sa_snapshot[8].f.unused[3] );
tran (\sa_snapshot[8][54] , \sa_snapshot[8].r.part1[22] );
tran (\sa_snapshot[8][54] , \sa_snapshot[8].f.unused[4] );
tran (\sa_snapshot[8][55] , \sa_snapshot[8].r.part1[23] );
tran (\sa_snapshot[8][55] , \sa_snapshot[8].f.unused[5] );
tran (\sa_snapshot[8][56] , \sa_snapshot[8].r.part1[24] );
tran (\sa_snapshot[8][56] , \sa_snapshot[8].f.unused[6] );
tran (\sa_snapshot[8][57] , \sa_snapshot[8].r.part1[25] );
tran (\sa_snapshot[8][57] , \sa_snapshot[8].f.unused[7] );
tran (\sa_snapshot[8][58] , \sa_snapshot[8].r.part1[26] );
tran (\sa_snapshot[8][58] , \sa_snapshot[8].f.unused[8] );
tran (\sa_snapshot[8][59] , \sa_snapshot[8].r.part1[27] );
tran (\sa_snapshot[8][59] , \sa_snapshot[8].f.unused[9] );
tran (\sa_snapshot[8][60] , \sa_snapshot[8].r.part1[28] );
tran (\sa_snapshot[8][60] , \sa_snapshot[8].f.unused[10] );
tran (\sa_snapshot[8][61] , \sa_snapshot[8].r.part1[29] );
tran (\sa_snapshot[8][61] , \sa_snapshot[8].f.unused[11] );
tran (\sa_snapshot[8][62] , \sa_snapshot[8].r.part1[30] );
tran (\sa_snapshot[8][62] , \sa_snapshot[8].f.unused[12] );
tran (\sa_snapshot[8][63] , \sa_snapshot[8].r.part1[31] );
tran (\sa_snapshot[8][63] , \sa_snapshot[8].f.unused[13] );
tran (\sa_snapshot[9][0] , \sa_snapshot[9].r.part0[0] );
tran (\sa_snapshot[9][0] , \sa_snapshot[9].f.lower[0] );
tran (\sa_snapshot[9][1] , \sa_snapshot[9].r.part0[1] );
tran (\sa_snapshot[9][1] , \sa_snapshot[9].f.lower[1] );
tran (\sa_snapshot[9][2] , \sa_snapshot[9].r.part0[2] );
tran (\sa_snapshot[9][2] , \sa_snapshot[9].f.lower[2] );
tran (\sa_snapshot[9][3] , \sa_snapshot[9].r.part0[3] );
tran (\sa_snapshot[9][3] , \sa_snapshot[9].f.lower[3] );
tran (\sa_snapshot[9][4] , \sa_snapshot[9].r.part0[4] );
tran (\sa_snapshot[9][4] , \sa_snapshot[9].f.lower[4] );
tran (\sa_snapshot[9][5] , \sa_snapshot[9].r.part0[5] );
tran (\sa_snapshot[9][5] , \sa_snapshot[9].f.lower[5] );
tran (\sa_snapshot[9][6] , \sa_snapshot[9].r.part0[6] );
tran (\sa_snapshot[9][6] , \sa_snapshot[9].f.lower[6] );
tran (\sa_snapshot[9][7] , \sa_snapshot[9].r.part0[7] );
tran (\sa_snapshot[9][7] , \sa_snapshot[9].f.lower[7] );
tran (\sa_snapshot[9][8] , \sa_snapshot[9].r.part0[8] );
tran (\sa_snapshot[9][8] , \sa_snapshot[9].f.lower[8] );
tran (\sa_snapshot[9][9] , \sa_snapshot[9].r.part0[9] );
tran (\sa_snapshot[9][9] , \sa_snapshot[9].f.lower[9] );
tran (\sa_snapshot[9][10] , \sa_snapshot[9].r.part0[10] );
tran (\sa_snapshot[9][10] , \sa_snapshot[9].f.lower[10] );
tran (\sa_snapshot[9][11] , \sa_snapshot[9].r.part0[11] );
tran (\sa_snapshot[9][11] , \sa_snapshot[9].f.lower[11] );
tran (\sa_snapshot[9][12] , \sa_snapshot[9].r.part0[12] );
tran (\sa_snapshot[9][12] , \sa_snapshot[9].f.lower[12] );
tran (\sa_snapshot[9][13] , \sa_snapshot[9].r.part0[13] );
tran (\sa_snapshot[9][13] , \sa_snapshot[9].f.lower[13] );
tran (\sa_snapshot[9][14] , \sa_snapshot[9].r.part0[14] );
tran (\sa_snapshot[9][14] , \sa_snapshot[9].f.lower[14] );
tran (\sa_snapshot[9][15] , \sa_snapshot[9].r.part0[15] );
tran (\sa_snapshot[9][15] , \sa_snapshot[9].f.lower[15] );
tran (\sa_snapshot[9][16] , \sa_snapshot[9].r.part0[16] );
tran (\sa_snapshot[9][16] , \sa_snapshot[9].f.lower[16] );
tran (\sa_snapshot[9][17] , \sa_snapshot[9].r.part0[17] );
tran (\sa_snapshot[9][17] , \sa_snapshot[9].f.lower[17] );
tran (\sa_snapshot[9][18] , \sa_snapshot[9].r.part0[18] );
tran (\sa_snapshot[9][18] , \sa_snapshot[9].f.lower[18] );
tran (\sa_snapshot[9][19] , \sa_snapshot[9].r.part0[19] );
tran (\sa_snapshot[9][19] , \sa_snapshot[9].f.lower[19] );
tran (\sa_snapshot[9][20] , \sa_snapshot[9].r.part0[20] );
tran (\sa_snapshot[9][20] , \sa_snapshot[9].f.lower[20] );
tran (\sa_snapshot[9][21] , \sa_snapshot[9].r.part0[21] );
tran (\sa_snapshot[9][21] , \sa_snapshot[9].f.lower[21] );
tran (\sa_snapshot[9][22] , \sa_snapshot[9].r.part0[22] );
tran (\sa_snapshot[9][22] , \sa_snapshot[9].f.lower[22] );
tran (\sa_snapshot[9][23] , \sa_snapshot[9].r.part0[23] );
tran (\sa_snapshot[9][23] , \sa_snapshot[9].f.lower[23] );
tran (\sa_snapshot[9][24] , \sa_snapshot[9].r.part0[24] );
tran (\sa_snapshot[9][24] , \sa_snapshot[9].f.lower[24] );
tran (\sa_snapshot[9][25] , \sa_snapshot[9].r.part0[25] );
tran (\sa_snapshot[9][25] , \sa_snapshot[9].f.lower[25] );
tran (\sa_snapshot[9][26] , \sa_snapshot[9].r.part0[26] );
tran (\sa_snapshot[9][26] , \sa_snapshot[9].f.lower[26] );
tran (\sa_snapshot[9][27] , \sa_snapshot[9].r.part0[27] );
tran (\sa_snapshot[9][27] , \sa_snapshot[9].f.lower[27] );
tran (\sa_snapshot[9][28] , \sa_snapshot[9].r.part0[28] );
tran (\sa_snapshot[9][28] , \sa_snapshot[9].f.lower[28] );
tran (\sa_snapshot[9][29] , \sa_snapshot[9].r.part0[29] );
tran (\sa_snapshot[9][29] , \sa_snapshot[9].f.lower[29] );
tran (\sa_snapshot[9][30] , \sa_snapshot[9].r.part0[30] );
tran (\sa_snapshot[9][30] , \sa_snapshot[9].f.lower[30] );
tran (\sa_snapshot[9][31] , \sa_snapshot[9].r.part0[31] );
tran (\sa_snapshot[9][31] , \sa_snapshot[9].f.lower[31] );
tran (\sa_snapshot[9][32] , \sa_snapshot[9].r.part1[0] );
tran (\sa_snapshot[9][32] , \sa_snapshot[9].f.upper[0] );
tran (\sa_snapshot[9][33] , \sa_snapshot[9].r.part1[1] );
tran (\sa_snapshot[9][33] , \sa_snapshot[9].f.upper[1] );
tran (\sa_snapshot[9][34] , \sa_snapshot[9].r.part1[2] );
tran (\sa_snapshot[9][34] , \sa_snapshot[9].f.upper[2] );
tran (\sa_snapshot[9][35] , \sa_snapshot[9].r.part1[3] );
tran (\sa_snapshot[9][35] , \sa_snapshot[9].f.upper[3] );
tran (\sa_snapshot[9][36] , \sa_snapshot[9].r.part1[4] );
tran (\sa_snapshot[9][36] , \sa_snapshot[9].f.upper[4] );
tran (\sa_snapshot[9][37] , \sa_snapshot[9].r.part1[5] );
tran (\sa_snapshot[9][37] , \sa_snapshot[9].f.upper[5] );
tran (\sa_snapshot[9][38] , \sa_snapshot[9].r.part1[6] );
tran (\sa_snapshot[9][38] , \sa_snapshot[9].f.upper[6] );
tran (\sa_snapshot[9][39] , \sa_snapshot[9].r.part1[7] );
tran (\sa_snapshot[9][39] , \sa_snapshot[9].f.upper[7] );
tran (\sa_snapshot[9][40] , \sa_snapshot[9].r.part1[8] );
tran (\sa_snapshot[9][40] , \sa_snapshot[9].f.upper[8] );
tran (\sa_snapshot[9][41] , \sa_snapshot[9].r.part1[9] );
tran (\sa_snapshot[9][41] , \sa_snapshot[9].f.upper[9] );
tran (\sa_snapshot[9][42] , \sa_snapshot[9].r.part1[10] );
tran (\sa_snapshot[9][42] , \sa_snapshot[9].f.upper[10] );
tran (\sa_snapshot[9][43] , \sa_snapshot[9].r.part1[11] );
tran (\sa_snapshot[9][43] , \sa_snapshot[9].f.upper[11] );
tran (\sa_snapshot[9][44] , \sa_snapshot[9].r.part1[12] );
tran (\sa_snapshot[9][44] , \sa_snapshot[9].f.upper[12] );
tran (\sa_snapshot[9][45] , \sa_snapshot[9].r.part1[13] );
tran (\sa_snapshot[9][45] , \sa_snapshot[9].f.upper[13] );
tran (\sa_snapshot[9][46] , \sa_snapshot[9].r.part1[14] );
tran (\sa_snapshot[9][46] , \sa_snapshot[9].f.upper[14] );
tran (\sa_snapshot[9][47] , \sa_snapshot[9].r.part1[15] );
tran (\sa_snapshot[9][47] , \sa_snapshot[9].f.upper[15] );
tran (\sa_snapshot[9][48] , \sa_snapshot[9].r.part1[16] );
tran (\sa_snapshot[9][48] , \sa_snapshot[9].f.upper[16] );
tran (\sa_snapshot[9][49] , \sa_snapshot[9].r.part1[17] );
tran (\sa_snapshot[9][49] , \sa_snapshot[9].f.upper[17] );
tran (\sa_snapshot[9][50] , \sa_snapshot[9].r.part1[18] );
tran (\sa_snapshot[9][50] , \sa_snapshot[9].f.unused[0] );
tran (\sa_snapshot[9][51] , \sa_snapshot[9].r.part1[19] );
tran (\sa_snapshot[9][51] , \sa_snapshot[9].f.unused[1] );
tran (\sa_snapshot[9][52] , \sa_snapshot[9].r.part1[20] );
tran (\sa_snapshot[9][52] , \sa_snapshot[9].f.unused[2] );
tran (\sa_snapshot[9][53] , \sa_snapshot[9].r.part1[21] );
tran (\sa_snapshot[9][53] , \sa_snapshot[9].f.unused[3] );
tran (\sa_snapshot[9][54] , \sa_snapshot[9].r.part1[22] );
tran (\sa_snapshot[9][54] , \sa_snapshot[9].f.unused[4] );
tran (\sa_snapshot[9][55] , \sa_snapshot[9].r.part1[23] );
tran (\sa_snapshot[9][55] , \sa_snapshot[9].f.unused[5] );
tran (\sa_snapshot[9][56] , \sa_snapshot[9].r.part1[24] );
tran (\sa_snapshot[9][56] , \sa_snapshot[9].f.unused[6] );
tran (\sa_snapshot[9][57] , \sa_snapshot[9].r.part1[25] );
tran (\sa_snapshot[9][57] , \sa_snapshot[9].f.unused[7] );
tran (\sa_snapshot[9][58] , \sa_snapshot[9].r.part1[26] );
tran (\sa_snapshot[9][58] , \sa_snapshot[9].f.unused[8] );
tran (\sa_snapshot[9][59] , \sa_snapshot[9].r.part1[27] );
tran (\sa_snapshot[9][59] , \sa_snapshot[9].f.unused[9] );
tran (\sa_snapshot[9][60] , \sa_snapshot[9].r.part1[28] );
tran (\sa_snapshot[9][60] , \sa_snapshot[9].f.unused[10] );
tran (\sa_snapshot[9][61] , \sa_snapshot[9].r.part1[29] );
tran (\sa_snapshot[9][61] , \sa_snapshot[9].f.unused[11] );
tran (\sa_snapshot[9][62] , \sa_snapshot[9].r.part1[30] );
tran (\sa_snapshot[9][62] , \sa_snapshot[9].f.unused[12] );
tran (\sa_snapshot[9][63] , \sa_snapshot[9].r.part1[31] );
tran (\sa_snapshot[9][63] , \sa_snapshot[9].f.unused[13] );
tran (\sa_snapshot[10][0] , \sa_snapshot[10].r.part0[0] );
tran (\sa_snapshot[10][0] , \sa_snapshot[10].f.lower[0] );
tran (\sa_snapshot[10][1] , \sa_snapshot[10].r.part0[1] );
tran (\sa_snapshot[10][1] , \sa_snapshot[10].f.lower[1] );
tran (\sa_snapshot[10][2] , \sa_snapshot[10].r.part0[2] );
tran (\sa_snapshot[10][2] , \sa_snapshot[10].f.lower[2] );
tran (\sa_snapshot[10][3] , \sa_snapshot[10].r.part0[3] );
tran (\sa_snapshot[10][3] , \sa_snapshot[10].f.lower[3] );
tran (\sa_snapshot[10][4] , \sa_snapshot[10].r.part0[4] );
tran (\sa_snapshot[10][4] , \sa_snapshot[10].f.lower[4] );
tran (\sa_snapshot[10][5] , \sa_snapshot[10].r.part0[5] );
tran (\sa_snapshot[10][5] , \sa_snapshot[10].f.lower[5] );
tran (\sa_snapshot[10][6] , \sa_snapshot[10].r.part0[6] );
tran (\sa_snapshot[10][6] , \sa_snapshot[10].f.lower[6] );
tran (\sa_snapshot[10][7] , \sa_snapshot[10].r.part0[7] );
tran (\sa_snapshot[10][7] , \sa_snapshot[10].f.lower[7] );
tran (\sa_snapshot[10][8] , \sa_snapshot[10].r.part0[8] );
tran (\sa_snapshot[10][8] , \sa_snapshot[10].f.lower[8] );
tran (\sa_snapshot[10][9] , \sa_snapshot[10].r.part0[9] );
tran (\sa_snapshot[10][9] , \sa_snapshot[10].f.lower[9] );
tran (\sa_snapshot[10][10] , \sa_snapshot[10].r.part0[10] );
tran (\sa_snapshot[10][10] , \sa_snapshot[10].f.lower[10] );
tran (\sa_snapshot[10][11] , \sa_snapshot[10].r.part0[11] );
tran (\sa_snapshot[10][11] , \sa_snapshot[10].f.lower[11] );
tran (\sa_snapshot[10][12] , \sa_snapshot[10].r.part0[12] );
tran (\sa_snapshot[10][12] , \sa_snapshot[10].f.lower[12] );
tran (\sa_snapshot[10][13] , \sa_snapshot[10].r.part0[13] );
tran (\sa_snapshot[10][13] , \sa_snapshot[10].f.lower[13] );
tran (\sa_snapshot[10][14] , \sa_snapshot[10].r.part0[14] );
tran (\sa_snapshot[10][14] , \sa_snapshot[10].f.lower[14] );
tran (\sa_snapshot[10][15] , \sa_snapshot[10].r.part0[15] );
tran (\sa_snapshot[10][15] , \sa_snapshot[10].f.lower[15] );
tran (\sa_snapshot[10][16] , \sa_snapshot[10].r.part0[16] );
tran (\sa_snapshot[10][16] , \sa_snapshot[10].f.lower[16] );
tran (\sa_snapshot[10][17] , \sa_snapshot[10].r.part0[17] );
tran (\sa_snapshot[10][17] , \sa_snapshot[10].f.lower[17] );
tran (\sa_snapshot[10][18] , \sa_snapshot[10].r.part0[18] );
tran (\sa_snapshot[10][18] , \sa_snapshot[10].f.lower[18] );
tran (\sa_snapshot[10][19] , \sa_snapshot[10].r.part0[19] );
tran (\sa_snapshot[10][19] , \sa_snapshot[10].f.lower[19] );
tran (\sa_snapshot[10][20] , \sa_snapshot[10].r.part0[20] );
tran (\sa_snapshot[10][20] , \sa_snapshot[10].f.lower[20] );
tran (\sa_snapshot[10][21] , \sa_snapshot[10].r.part0[21] );
tran (\sa_snapshot[10][21] , \sa_snapshot[10].f.lower[21] );
tran (\sa_snapshot[10][22] , \sa_snapshot[10].r.part0[22] );
tran (\sa_snapshot[10][22] , \sa_snapshot[10].f.lower[22] );
tran (\sa_snapshot[10][23] , \sa_snapshot[10].r.part0[23] );
tran (\sa_snapshot[10][23] , \sa_snapshot[10].f.lower[23] );
tran (\sa_snapshot[10][24] , \sa_snapshot[10].r.part0[24] );
tran (\sa_snapshot[10][24] , \sa_snapshot[10].f.lower[24] );
tran (\sa_snapshot[10][25] , \sa_snapshot[10].r.part0[25] );
tran (\sa_snapshot[10][25] , \sa_snapshot[10].f.lower[25] );
tran (\sa_snapshot[10][26] , \sa_snapshot[10].r.part0[26] );
tran (\sa_snapshot[10][26] , \sa_snapshot[10].f.lower[26] );
tran (\sa_snapshot[10][27] , \sa_snapshot[10].r.part0[27] );
tran (\sa_snapshot[10][27] , \sa_snapshot[10].f.lower[27] );
tran (\sa_snapshot[10][28] , \sa_snapshot[10].r.part0[28] );
tran (\sa_snapshot[10][28] , \sa_snapshot[10].f.lower[28] );
tran (\sa_snapshot[10][29] , \sa_snapshot[10].r.part0[29] );
tran (\sa_snapshot[10][29] , \sa_snapshot[10].f.lower[29] );
tran (\sa_snapshot[10][30] , \sa_snapshot[10].r.part0[30] );
tran (\sa_snapshot[10][30] , \sa_snapshot[10].f.lower[30] );
tran (\sa_snapshot[10][31] , \sa_snapshot[10].r.part0[31] );
tran (\sa_snapshot[10][31] , \sa_snapshot[10].f.lower[31] );
tran (\sa_snapshot[10][32] , \sa_snapshot[10].r.part1[0] );
tran (\sa_snapshot[10][32] , \sa_snapshot[10].f.upper[0] );
tran (\sa_snapshot[10][33] , \sa_snapshot[10].r.part1[1] );
tran (\sa_snapshot[10][33] , \sa_snapshot[10].f.upper[1] );
tran (\sa_snapshot[10][34] , \sa_snapshot[10].r.part1[2] );
tran (\sa_snapshot[10][34] , \sa_snapshot[10].f.upper[2] );
tran (\sa_snapshot[10][35] , \sa_snapshot[10].r.part1[3] );
tran (\sa_snapshot[10][35] , \sa_snapshot[10].f.upper[3] );
tran (\sa_snapshot[10][36] , \sa_snapshot[10].r.part1[4] );
tran (\sa_snapshot[10][36] , \sa_snapshot[10].f.upper[4] );
tran (\sa_snapshot[10][37] , \sa_snapshot[10].r.part1[5] );
tran (\sa_snapshot[10][37] , \sa_snapshot[10].f.upper[5] );
tran (\sa_snapshot[10][38] , \sa_snapshot[10].r.part1[6] );
tran (\sa_snapshot[10][38] , \sa_snapshot[10].f.upper[6] );
tran (\sa_snapshot[10][39] , \sa_snapshot[10].r.part1[7] );
tran (\sa_snapshot[10][39] , \sa_snapshot[10].f.upper[7] );
tran (\sa_snapshot[10][40] , \sa_snapshot[10].r.part1[8] );
tran (\sa_snapshot[10][40] , \sa_snapshot[10].f.upper[8] );
tran (\sa_snapshot[10][41] , \sa_snapshot[10].r.part1[9] );
tran (\sa_snapshot[10][41] , \sa_snapshot[10].f.upper[9] );
tran (\sa_snapshot[10][42] , \sa_snapshot[10].r.part1[10] );
tran (\sa_snapshot[10][42] , \sa_snapshot[10].f.upper[10] );
tran (\sa_snapshot[10][43] , \sa_snapshot[10].r.part1[11] );
tran (\sa_snapshot[10][43] , \sa_snapshot[10].f.upper[11] );
tran (\sa_snapshot[10][44] , \sa_snapshot[10].r.part1[12] );
tran (\sa_snapshot[10][44] , \sa_snapshot[10].f.upper[12] );
tran (\sa_snapshot[10][45] , \sa_snapshot[10].r.part1[13] );
tran (\sa_snapshot[10][45] , \sa_snapshot[10].f.upper[13] );
tran (\sa_snapshot[10][46] , \sa_snapshot[10].r.part1[14] );
tran (\sa_snapshot[10][46] , \sa_snapshot[10].f.upper[14] );
tran (\sa_snapshot[10][47] , \sa_snapshot[10].r.part1[15] );
tran (\sa_snapshot[10][47] , \sa_snapshot[10].f.upper[15] );
tran (\sa_snapshot[10][48] , \sa_snapshot[10].r.part1[16] );
tran (\sa_snapshot[10][48] , \sa_snapshot[10].f.upper[16] );
tran (\sa_snapshot[10][49] , \sa_snapshot[10].r.part1[17] );
tran (\sa_snapshot[10][49] , \sa_snapshot[10].f.upper[17] );
tran (\sa_snapshot[10][50] , \sa_snapshot[10].r.part1[18] );
tran (\sa_snapshot[10][50] , \sa_snapshot[10].f.unused[0] );
tran (\sa_snapshot[10][51] , \sa_snapshot[10].r.part1[19] );
tran (\sa_snapshot[10][51] , \sa_snapshot[10].f.unused[1] );
tran (\sa_snapshot[10][52] , \sa_snapshot[10].r.part1[20] );
tran (\sa_snapshot[10][52] , \sa_snapshot[10].f.unused[2] );
tran (\sa_snapshot[10][53] , \sa_snapshot[10].r.part1[21] );
tran (\sa_snapshot[10][53] , \sa_snapshot[10].f.unused[3] );
tran (\sa_snapshot[10][54] , \sa_snapshot[10].r.part1[22] );
tran (\sa_snapshot[10][54] , \sa_snapshot[10].f.unused[4] );
tran (\sa_snapshot[10][55] , \sa_snapshot[10].r.part1[23] );
tran (\sa_snapshot[10][55] , \sa_snapshot[10].f.unused[5] );
tran (\sa_snapshot[10][56] , \sa_snapshot[10].r.part1[24] );
tran (\sa_snapshot[10][56] , \sa_snapshot[10].f.unused[6] );
tran (\sa_snapshot[10][57] , \sa_snapshot[10].r.part1[25] );
tran (\sa_snapshot[10][57] , \sa_snapshot[10].f.unused[7] );
tran (\sa_snapshot[10][58] , \sa_snapshot[10].r.part1[26] );
tran (\sa_snapshot[10][58] , \sa_snapshot[10].f.unused[8] );
tran (\sa_snapshot[10][59] , \sa_snapshot[10].r.part1[27] );
tran (\sa_snapshot[10][59] , \sa_snapshot[10].f.unused[9] );
tran (\sa_snapshot[10][60] , \sa_snapshot[10].r.part1[28] );
tran (\sa_snapshot[10][60] , \sa_snapshot[10].f.unused[10] );
tran (\sa_snapshot[10][61] , \sa_snapshot[10].r.part1[29] );
tran (\sa_snapshot[10][61] , \sa_snapshot[10].f.unused[11] );
tran (\sa_snapshot[10][62] , \sa_snapshot[10].r.part1[30] );
tran (\sa_snapshot[10][62] , \sa_snapshot[10].f.unused[12] );
tran (\sa_snapshot[10][63] , \sa_snapshot[10].r.part1[31] );
tran (\sa_snapshot[10][63] , \sa_snapshot[10].f.unused[13] );
tran (\sa_snapshot[11][0] , \sa_snapshot[11].r.part0[0] );
tran (\sa_snapshot[11][0] , \sa_snapshot[11].f.lower[0] );
tran (\sa_snapshot[11][1] , \sa_snapshot[11].r.part0[1] );
tran (\sa_snapshot[11][1] , \sa_snapshot[11].f.lower[1] );
tran (\sa_snapshot[11][2] , \sa_snapshot[11].r.part0[2] );
tran (\sa_snapshot[11][2] , \sa_snapshot[11].f.lower[2] );
tran (\sa_snapshot[11][3] , \sa_snapshot[11].r.part0[3] );
tran (\sa_snapshot[11][3] , \sa_snapshot[11].f.lower[3] );
tran (\sa_snapshot[11][4] , \sa_snapshot[11].r.part0[4] );
tran (\sa_snapshot[11][4] , \sa_snapshot[11].f.lower[4] );
tran (\sa_snapshot[11][5] , \sa_snapshot[11].r.part0[5] );
tran (\sa_snapshot[11][5] , \sa_snapshot[11].f.lower[5] );
tran (\sa_snapshot[11][6] , \sa_snapshot[11].r.part0[6] );
tran (\sa_snapshot[11][6] , \sa_snapshot[11].f.lower[6] );
tran (\sa_snapshot[11][7] , \sa_snapshot[11].r.part0[7] );
tran (\sa_snapshot[11][7] , \sa_snapshot[11].f.lower[7] );
tran (\sa_snapshot[11][8] , \sa_snapshot[11].r.part0[8] );
tran (\sa_snapshot[11][8] , \sa_snapshot[11].f.lower[8] );
tran (\sa_snapshot[11][9] , \sa_snapshot[11].r.part0[9] );
tran (\sa_snapshot[11][9] , \sa_snapshot[11].f.lower[9] );
tran (\sa_snapshot[11][10] , \sa_snapshot[11].r.part0[10] );
tran (\sa_snapshot[11][10] , \sa_snapshot[11].f.lower[10] );
tran (\sa_snapshot[11][11] , \sa_snapshot[11].r.part0[11] );
tran (\sa_snapshot[11][11] , \sa_snapshot[11].f.lower[11] );
tran (\sa_snapshot[11][12] , \sa_snapshot[11].r.part0[12] );
tran (\sa_snapshot[11][12] , \sa_snapshot[11].f.lower[12] );
tran (\sa_snapshot[11][13] , \sa_snapshot[11].r.part0[13] );
tran (\sa_snapshot[11][13] , \sa_snapshot[11].f.lower[13] );
tran (\sa_snapshot[11][14] , \sa_snapshot[11].r.part0[14] );
tran (\sa_snapshot[11][14] , \sa_snapshot[11].f.lower[14] );
tran (\sa_snapshot[11][15] , \sa_snapshot[11].r.part0[15] );
tran (\sa_snapshot[11][15] , \sa_snapshot[11].f.lower[15] );
tran (\sa_snapshot[11][16] , \sa_snapshot[11].r.part0[16] );
tran (\sa_snapshot[11][16] , \sa_snapshot[11].f.lower[16] );
tran (\sa_snapshot[11][17] , \sa_snapshot[11].r.part0[17] );
tran (\sa_snapshot[11][17] , \sa_snapshot[11].f.lower[17] );
tran (\sa_snapshot[11][18] , \sa_snapshot[11].r.part0[18] );
tran (\sa_snapshot[11][18] , \sa_snapshot[11].f.lower[18] );
tran (\sa_snapshot[11][19] , \sa_snapshot[11].r.part0[19] );
tran (\sa_snapshot[11][19] , \sa_snapshot[11].f.lower[19] );
tran (\sa_snapshot[11][20] , \sa_snapshot[11].r.part0[20] );
tran (\sa_snapshot[11][20] , \sa_snapshot[11].f.lower[20] );
tran (\sa_snapshot[11][21] , \sa_snapshot[11].r.part0[21] );
tran (\sa_snapshot[11][21] , \sa_snapshot[11].f.lower[21] );
tran (\sa_snapshot[11][22] , \sa_snapshot[11].r.part0[22] );
tran (\sa_snapshot[11][22] , \sa_snapshot[11].f.lower[22] );
tran (\sa_snapshot[11][23] , \sa_snapshot[11].r.part0[23] );
tran (\sa_snapshot[11][23] , \sa_snapshot[11].f.lower[23] );
tran (\sa_snapshot[11][24] , \sa_snapshot[11].r.part0[24] );
tran (\sa_snapshot[11][24] , \sa_snapshot[11].f.lower[24] );
tran (\sa_snapshot[11][25] , \sa_snapshot[11].r.part0[25] );
tran (\sa_snapshot[11][25] , \sa_snapshot[11].f.lower[25] );
tran (\sa_snapshot[11][26] , \sa_snapshot[11].r.part0[26] );
tran (\sa_snapshot[11][26] , \sa_snapshot[11].f.lower[26] );
tran (\sa_snapshot[11][27] , \sa_snapshot[11].r.part0[27] );
tran (\sa_snapshot[11][27] , \sa_snapshot[11].f.lower[27] );
tran (\sa_snapshot[11][28] , \sa_snapshot[11].r.part0[28] );
tran (\sa_snapshot[11][28] , \sa_snapshot[11].f.lower[28] );
tran (\sa_snapshot[11][29] , \sa_snapshot[11].r.part0[29] );
tran (\sa_snapshot[11][29] , \sa_snapshot[11].f.lower[29] );
tran (\sa_snapshot[11][30] , \sa_snapshot[11].r.part0[30] );
tran (\sa_snapshot[11][30] , \sa_snapshot[11].f.lower[30] );
tran (\sa_snapshot[11][31] , \sa_snapshot[11].r.part0[31] );
tran (\sa_snapshot[11][31] , \sa_snapshot[11].f.lower[31] );
tran (\sa_snapshot[11][32] , \sa_snapshot[11].r.part1[0] );
tran (\sa_snapshot[11][32] , \sa_snapshot[11].f.upper[0] );
tran (\sa_snapshot[11][33] , \sa_snapshot[11].r.part1[1] );
tran (\sa_snapshot[11][33] , \sa_snapshot[11].f.upper[1] );
tran (\sa_snapshot[11][34] , \sa_snapshot[11].r.part1[2] );
tran (\sa_snapshot[11][34] , \sa_snapshot[11].f.upper[2] );
tran (\sa_snapshot[11][35] , \sa_snapshot[11].r.part1[3] );
tran (\sa_snapshot[11][35] , \sa_snapshot[11].f.upper[3] );
tran (\sa_snapshot[11][36] , \sa_snapshot[11].r.part1[4] );
tran (\sa_snapshot[11][36] , \sa_snapshot[11].f.upper[4] );
tran (\sa_snapshot[11][37] , \sa_snapshot[11].r.part1[5] );
tran (\sa_snapshot[11][37] , \sa_snapshot[11].f.upper[5] );
tran (\sa_snapshot[11][38] , \sa_snapshot[11].r.part1[6] );
tran (\sa_snapshot[11][38] , \sa_snapshot[11].f.upper[6] );
tran (\sa_snapshot[11][39] , \sa_snapshot[11].r.part1[7] );
tran (\sa_snapshot[11][39] , \sa_snapshot[11].f.upper[7] );
tran (\sa_snapshot[11][40] , \sa_snapshot[11].r.part1[8] );
tran (\sa_snapshot[11][40] , \sa_snapshot[11].f.upper[8] );
tran (\sa_snapshot[11][41] , \sa_snapshot[11].r.part1[9] );
tran (\sa_snapshot[11][41] , \sa_snapshot[11].f.upper[9] );
tran (\sa_snapshot[11][42] , \sa_snapshot[11].r.part1[10] );
tran (\sa_snapshot[11][42] , \sa_snapshot[11].f.upper[10] );
tran (\sa_snapshot[11][43] , \sa_snapshot[11].r.part1[11] );
tran (\sa_snapshot[11][43] , \sa_snapshot[11].f.upper[11] );
tran (\sa_snapshot[11][44] , \sa_snapshot[11].r.part1[12] );
tran (\sa_snapshot[11][44] , \sa_snapshot[11].f.upper[12] );
tran (\sa_snapshot[11][45] , \sa_snapshot[11].r.part1[13] );
tran (\sa_snapshot[11][45] , \sa_snapshot[11].f.upper[13] );
tran (\sa_snapshot[11][46] , \sa_snapshot[11].r.part1[14] );
tran (\sa_snapshot[11][46] , \sa_snapshot[11].f.upper[14] );
tran (\sa_snapshot[11][47] , \sa_snapshot[11].r.part1[15] );
tran (\sa_snapshot[11][47] , \sa_snapshot[11].f.upper[15] );
tran (\sa_snapshot[11][48] , \sa_snapshot[11].r.part1[16] );
tran (\sa_snapshot[11][48] , \sa_snapshot[11].f.upper[16] );
tran (\sa_snapshot[11][49] , \sa_snapshot[11].r.part1[17] );
tran (\sa_snapshot[11][49] , \sa_snapshot[11].f.upper[17] );
tran (\sa_snapshot[11][50] , \sa_snapshot[11].r.part1[18] );
tran (\sa_snapshot[11][50] , \sa_snapshot[11].f.unused[0] );
tran (\sa_snapshot[11][51] , \sa_snapshot[11].r.part1[19] );
tran (\sa_snapshot[11][51] , \sa_snapshot[11].f.unused[1] );
tran (\sa_snapshot[11][52] , \sa_snapshot[11].r.part1[20] );
tran (\sa_snapshot[11][52] , \sa_snapshot[11].f.unused[2] );
tran (\sa_snapshot[11][53] , \sa_snapshot[11].r.part1[21] );
tran (\sa_snapshot[11][53] , \sa_snapshot[11].f.unused[3] );
tran (\sa_snapshot[11][54] , \sa_snapshot[11].r.part1[22] );
tran (\sa_snapshot[11][54] , \sa_snapshot[11].f.unused[4] );
tran (\sa_snapshot[11][55] , \sa_snapshot[11].r.part1[23] );
tran (\sa_snapshot[11][55] , \sa_snapshot[11].f.unused[5] );
tran (\sa_snapshot[11][56] , \sa_snapshot[11].r.part1[24] );
tran (\sa_snapshot[11][56] , \sa_snapshot[11].f.unused[6] );
tran (\sa_snapshot[11][57] , \sa_snapshot[11].r.part1[25] );
tran (\sa_snapshot[11][57] , \sa_snapshot[11].f.unused[7] );
tran (\sa_snapshot[11][58] , \sa_snapshot[11].r.part1[26] );
tran (\sa_snapshot[11][58] , \sa_snapshot[11].f.unused[8] );
tran (\sa_snapshot[11][59] , \sa_snapshot[11].r.part1[27] );
tran (\sa_snapshot[11][59] , \sa_snapshot[11].f.unused[9] );
tran (\sa_snapshot[11][60] , \sa_snapshot[11].r.part1[28] );
tran (\sa_snapshot[11][60] , \sa_snapshot[11].f.unused[10] );
tran (\sa_snapshot[11][61] , \sa_snapshot[11].r.part1[29] );
tran (\sa_snapshot[11][61] , \sa_snapshot[11].f.unused[11] );
tran (\sa_snapshot[11][62] , \sa_snapshot[11].r.part1[30] );
tran (\sa_snapshot[11][62] , \sa_snapshot[11].f.unused[12] );
tran (\sa_snapshot[11][63] , \sa_snapshot[11].r.part1[31] );
tran (\sa_snapshot[11][63] , \sa_snapshot[11].f.unused[13] );
tran (\sa_snapshot[12][0] , \sa_snapshot[12].r.part0[0] );
tran (\sa_snapshot[12][0] , \sa_snapshot[12].f.lower[0] );
tran (\sa_snapshot[12][1] , \sa_snapshot[12].r.part0[1] );
tran (\sa_snapshot[12][1] , \sa_snapshot[12].f.lower[1] );
tran (\sa_snapshot[12][2] , \sa_snapshot[12].r.part0[2] );
tran (\sa_snapshot[12][2] , \sa_snapshot[12].f.lower[2] );
tran (\sa_snapshot[12][3] , \sa_snapshot[12].r.part0[3] );
tran (\sa_snapshot[12][3] , \sa_snapshot[12].f.lower[3] );
tran (\sa_snapshot[12][4] , \sa_snapshot[12].r.part0[4] );
tran (\sa_snapshot[12][4] , \sa_snapshot[12].f.lower[4] );
tran (\sa_snapshot[12][5] , \sa_snapshot[12].r.part0[5] );
tran (\sa_snapshot[12][5] , \sa_snapshot[12].f.lower[5] );
tran (\sa_snapshot[12][6] , \sa_snapshot[12].r.part0[6] );
tran (\sa_snapshot[12][6] , \sa_snapshot[12].f.lower[6] );
tran (\sa_snapshot[12][7] , \sa_snapshot[12].r.part0[7] );
tran (\sa_snapshot[12][7] , \sa_snapshot[12].f.lower[7] );
tran (\sa_snapshot[12][8] , \sa_snapshot[12].r.part0[8] );
tran (\sa_snapshot[12][8] , \sa_snapshot[12].f.lower[8] );
tran (\sa_snapshot[12][9] , \sa_snapshot[12].r.part0[9] );
tran (\sa_snapshot[12][9] , \sa_snapshot[12].f.lower[9] );
tran (\sa_snapshot[12][10] , \sa_snapshot[12].r.part0[10] );
tran (\sa_snapshot[12][10] , \sa_snapshot[12].f.lower[10] );
tran (\sa_snapshot[12][11] , \sa_snapshot[12].r.part0[11] );
tran (\sa_snapshot[12][11] , \sa_snapshot[12].f.lower[11] );
tran (\sa_snapshot[12][12] , \sa_snapshot[12].r.part0[12] );
tran (\sa_snapshot[12][12] , \sa_snapshot[12].f.lower[12] );
tran (\sa_snapshot[12][13] , \sa_snapshot[12].r.part0[13] );
tran (\sa_snapshot[12][13] , \sa_snapshot[12].f.lower[13] );
tran (\sa_snapshot[12][14] , \sa_snapshot[12].r.part0[14] );
tran (\sa_snapshot[12][14] , \sa_snapshot[12].f.lower[14] );
tran (\sa_snapshot[12][15] , \sa_snapshot[12].r.part0[15] );
tran (\sa_snapshot[12][15] , \sa_snapshot[12].f.lower[15] );
tran (\sa_snapshot[12][16] , \sa_snapshot[12].r.part0[16] );
tran (\sa_snapshot[12][16] , \sa_snapshot[12].f.lower[16] );
tran (\sa_snapshot[12][17] , \sa_snapshot[12].r.part0[17] );
tran (\sa_snapshot[12][17] , \sa_snapshot[12].f.lower[17] );
tran (\sa_snapshot[12][18] , \sa_snapshot[12].r.part0[18] );
tran (\sa_snapshot[12][18] , \sa_snapshot[12].f.lower[18] );
tran (\sa_snapshot[12][19] , \sa_snapshot[12].r.part0[19] );
tran (\sa_snapshot[12][19] , \sa_snapshot[12].f.lower[19] );
tran (\sa_snapshot[12][20] , \sa_snapshot[12].r.part0[20] );
tran (\sa_snapshot[12][20] , \sa_snapshot[12].f.lower[20] );
tran (\sa_snapshot[12][21] , \sa_snapshot[12].r.part0[21] );
tran (\sa_snapshot[12][21] , \sa_snapshot[12].f.lower[21] );
tran (\sa_snapshot[12][22] , \sa_snapshot[12].r.part0[22] );
tran (\sa_snapshot[12][22] , \sa_snapshot[12].f.lower[22] );
tran (\sa_snapshot[12][23] , \sa_snapshot[12].r.part0[23] );
tran (\sa_snapshot[12][23] , \sa_snapshot[12].f.lower[23] );
tran (\sa_snapshot[12][24] , \sa_snapshot[12].r.part0[24] );
tran (\sa_snapshot[12][24] , \sa_snapshot[12].f.lower[24] );
tran (\sa_snapshot[12][25] , \sa_snapshot[12].r.part0[25] );
tran (\sa_snapshot[12][25] , \sa_snapshot[12].f.lower[25] );
tran (\sa_snapshot[12][26] , \sa_snapshot[12].r.part0[26] );
tran (\sa_snapshot[12][26] , \sa_snapshot[12].f.lower[26] );
tran (\sa_snapshot[12][27] , \sa_snapshot[12].r.part0[27] );
tran (\sa_snapshot[12][27] , \sa_snapshot[12].f.lower[27] );
tran (\sa_snapshot[12][28] , \sa_snapshot[12].r.part0[28] );
tran (\sa_snapshot[12][28] , \sa_snapshot[12].f.lower[28] );
tran (\sa_snapshot[12][29] , \sa_snapshot[12].r.part0[29] );
tran (\sa_snapshot[12][29] , \sa_snapshot[12].f.lower[29] );
tran (\sa_snapshot[12][30] , \sa_snapshot[12].r.part0[30] );
tran (\sa_snapshot[12][30] , \sa_snapshot[12].f.lower[30] );
tran (\sa_snapshot[12][31] , \sa_snapshot[12].r.part0[31] );
tran (\sa_snapshot[12][31] , \sa_snapshot[12].f.lower[31] );
tran (\sa_snapshot[12][32] , \sa_snapshot[12].r.part1[0] );
tran (\sa_snapshot[12][32] , \sa_snapshot[12].f.upper[0] );
tran (\sa_snapshot[12][33] , \sa_snapshot[12].r.part1[1] );
tran (\sa_snapshot[12][33] , \sa_snapshot[12].f.upper[1] );
tran (\sa_snapshot[12][34] , \sa_snapshot[12].r.part1[2] );
tran (\sa_snapshot[12][34] , \sa_snapshot[12].f.upper[2] );
tran (\sa_snapshot[12][35] , \sa_snapshot[12].r.part1[3] );
tran (\sa_snapshot[12][35] , \sa_snapshot[12].f.upper[3] );
tran (\sa_snapshot[12][36] , \sa_snapshot[12].r.part1[4] );
tran (\sa_snapshot[12][36] , \sa_snapshot[12].f.upper[4] );
tran (\sa_snapshot[12][37] , \sa_snapshot[12].r.part1[5] );
tran (\sa_snapshot[12][37] , \sa_snapshot[12].f.upper[5] );
tran (\sa_snapshot[12][38] , \sa_snapshot[12].r.part1[6] );
tran (\sa_snapshot[12][38] , \sa_snapshot[12].f.upper[6] );
tran (\sa_snapshot[12][39] , \sa_snapshot[12].r.part1[7] );
tran (\sa_snapshot[12][39] , \sa_snapshot[12].f.upper[7] );
tran (\sa_snapshot[12][40] , \sa_snapshot[12].r.part1[8] );
tran (\sa_snapshot[12][40] , \sa_snapshot[12].f.upper[8] );
tran (\sa_snapshot[12][41] , \sa_snapshot[12].r.part1[9] );
tran (\sa_snapshot[12][41] , \sa_snapshot[12].f.upper[9] );
tran (\sa_snapshot[12][42] , \sa_snapshot[12].r.part1[10] );
tran (\sa_snapshot[12][42] , \sa_snapshot[12].f.upper[10] );
tran (\sa_snapshot[12][43] , \sa_snapshot[12].r.part1[11] );
tran (\sa_snapshot[12][43] , \sa_snapshot[12].f.upper[11] );
tran (\sa_snapshot[12][44] , \sa_snapshot[12].r.part1[12] );
tran (\sa_snapshot[12][44] , \sa_snapshot[12].f.upper[12] );
tran (\sa_snapshot[12][45] , \sa_snapshot[12].r.part1[13] );
tran (\sa_snapshot[12][45] , \sa_snapshot[12].f.upper[13] );
tran (\sa_snapshot[12][46] , \sa_snapshot[12].r.part1[14] );
tran (\sa_snapshot[12][46] , \sa_snapshot[12].f.upper[14] );
tran (\sa_snapshot[12][47] , \sa_snapshot[12].r.part1[15] );
tran (\sa_snapshot[12][47] , \sa_snapshot[12].f.upper[15] );
tran (\sa_snapshot[12][48] , \sa_snapshot[12].r.part1[16] );
tran (\sa_snapshot[12][48] , \sa_snapshot[12].f.upper[16] );
tran (\sa_snapshot[12][49] , \sa_snapshot[12].r.part1[17] );
tran (\sa_snapshot[12][49] , \sa_snapshot[12].f.upper[17] );
tran (\sa_snapshot[12][50] , \sa_snapshot[12].r.part1[18] );
tran (\sa_snapshot[12][50] , \sa_snapshot[12].f.unused[0] );
tran (\sa_snapshot[12][51] , \sa_snapshot[12].r.part1[19] );
tran (\sa_snapshot[12][51] , \sa_snapshot[12].f.unused[1] );
tran (\sa_snapshot[12][52] , \sa_snapshot[12].r.part1[20] );
tran (\sa_snapshot[12][52] , \sa_snapshot[12].f.unused[2] );
tran (\sa_snapshot[12][53] , \sa_snapshot[12].r.part1[21] );
tran (\sa_snapshot[12][53] , \sa_snapshot[12].f.unused[3] );
tran (\sa_snapshot[12][54] , \sa_snapshot[12].r.part1[22] );
tran (\sa_snapshot[12][54] , \sa_snapshot[12].f.unused[4] );
tran (\sa_snapshot[12][55] , \sa_snapshot[12].r.part1[23] );
tran (\sa_snapshot[12][55] , \sa_snapshot[12].f.unused[5] );
tran (\sa_snapshot[12][56] , \sa_snapshot[12].r.part1[24] );
tran (\sa_snapshot[12][56] , \sa_snapshot[12].f.unused[6] );
tran (\sa_snapshot[12][57] , \sa_snapshot[12].r.part1[25] );
tran (\sa_snapshot[12][57] , \sa_snapshot[12].f.unused[7] );
tran (\sa_snapshot[12][58] , \sa_snapshot[12].r.part1[26] );
tran (\sa_snapshot[12][58] , \sa_snapshot[12].f.unused[8] );
tran (\sa_snapshot[12][59] , \sa_snapshot[12].r.part1[27] );
tran (\sa_snapshot[12][59] , \sa_snapshot[12].f.unused[9] );
tran (\sa_snapshot[12][60] , \sa_snapshot[12].r.part1[28] );
tran (\sa_snapshot[12][60] , \sa_snapshot[12].f.unused[10] );
tran (\sa_snapshot[12][61] , \sa_snapshot[12].r.part1[29] );
tran (\sa_snapshot[12][61] , \sa_snapshot[12].f.unused[11] );
tran (\sa_snapshot[12][62] , \sa_snapshot[12].r.part1[30] );
tran (\sa_snapshot[12][62] , \sa_snapshot[12].f.unused[12] );
tran (\sa_snapshot[12][63] , \sa_snapshot[12].r.part1[31] );
tran (\sa_snapshot[12][63] , \sa_snapshot[12].f.unused[13] );
tran (\sa_snapshot[13][0] , \sa_snapshot[13].r.part0[0] );
tran (\sa_snapshot[13][0] , \sa_snapshot[13].f.lower[0] );
tran (\sa_snapshot[13][1] , \sa_snapshot[13].r.part0[1] );
tran (\sa_snapshot[13][1] , \sa_snapshot[13].f.lower[1] );
tran (\sa_snapshot[13][2] , \sa_snapshot[13].r.part0[2] );
tran (\sa_snapshot[13][2] , \sa_snapshot[13].f.lower[2] );
tran (\sa_snapshot[13][3] , \sa_snapshot[13].r.part0[3] );
tran (\sa_snapshot[13][3] , \sa_snapshot[13].f.lower[3] );
tran (\sa_snapshot[13][4] , \sa_snapshot[13].r.part0[4] );
tran (\sa_snapshot[13][4] , \sa_snapshot[13].f.lower[4] );
tran (\sa_snapshot[13][5] , \sa_snapshot[13].r.part0[5] );
tran (\sa_snapshot[13][5] , \sa_snapshot[13].f.lower[5] );
tran (\sa_snapshot[13][6] , \sa_snapshot[13].r.part0[6] );
tran (\sa_snapshot[13][6] , \sa_snapshot[13].f.lower[6] );
tran (\sa_snapshot[13][7] , \sa_snapshot[13].r.part0[7] );
tran (\sa_snapshot[13][7] , \sa_snapshot[13].f.lower[7] );
tran (\sa_snapshot[13][8] , \sa_snapshot[13].r.part0[8] );
tran (\sa_snapshot[13][8] , \sa_snapshot[13].f.lower[8] );
tran (\sa_snapshot[13][9] , \sa_snapshot[13].r.part0[9] );
tran (\sa_snapshot[13][9] , \sa_snapshot[13].f.lower[9] );
tran (\sa_snapshot[13][10] , \sa_snapshot[13].r.part0[10] );
tran (\sa_snapshot[13][10] , \sa_snapshot[13].f.lower[10] );
tran (\sa_snapshot[13][11] , \sa_snapshot[13].r.part0[11] );
tran (\sa_snapshot[13][11] , \sa_snapshot[13].f.lower[11] );
tran (\sa_snapshot[13][12] , \sa_snapshot[13].r.part0[12] );
tran (\sa_snapshot[13][12] , \sa_snapshot[13].f.lower[12] );
tran (\sa_snapshot[13][13] , \sa_snapshot[13].r.part0[13] );
tran (\sa_snapshot[13][13] , \sa_snapshot[13].f.lower[13] );
tran (\sa_snapshot[13][14] , \sa_snapshot[13].r.part0[14] );
tran (\sa_snapshot[13][14] , \sa_snapshot[13].f.lower[14] );
tran (\sa_snapshot[13][15] , \sa_snapshot[13].r.part0[15] );
tran (\sa_snapshot[13][15] , \sa_snapshot[13].f.lower[15] );
tran (\sa_snapshot[13][16] , \sa_snapshot[13].r.part0[16] );
tran (\sa_snapshot[13][16] , \sa_snapshot[13].f.lower[16] );
tran (\sa_snapshot[13][17] , \sa_snapshot[13].r.part0[17] );
tran (\sa_snapshot[13][17] , \sa_snapshot[13].f.lower[17] );
tran (\sa_snapshot[13][18] , \sa_snapshot[13].r.part0[18] );
tran (\sa_snapshot[13][18] , \sa_snapshot[13].f.lower[18] );
tran (\sa_snapshot[13][19] , \sa_snapshot[13].r.part0[19] );
tran (\sa_snapshot[13][19] , \sa_snapshot[13].f.lower[19] );
tran (\sa_snapshot[13][20] , \sa_snapshot[13].r.part0[20] );
tran (\sa_snapshot[13][20] , \sa_snapshot[13].f.lower[20] );
tran (\sa_snapshot[13][21] , \sa_snapshot[13].r.part0[21] );
tran (\sa_snapshot[13][21] , \sa_snapshot[13].f.lower[21] );
tran (\sa_snapshot[13][22] , \sa_snapshot[13].r.part0[22] );
tran (\sa_snapshot[13][22] , \sa_snapshot[13].f.lower[22] );
tran (\sa_snapshot[13][23] , \sa_snapshot[13].r.part0[23] );
tran (\sa_snapshot[13][23] , \sa_snapshot[13].f.lower[23] );
tran (\sa_snapshot[13][24] , \sa_snapshot[13].r.part0[24] );
tran (\sa_snapshot[13][24] , \sa_snapshot[13].f.lower[24] );
tran (\sa_snapshot[13][25] , \sa_snapshot[13].r.part0[25] );
tran (\sa_snapshot[13][25] , \sa_snapshot[13].f.lower[25] );
tran (\sa_snapshot[13][26] , \sa_snapshot[13].r.part0[26] );
tran (\sa_snapshot[13][26] , \sa_snapshot[13].f.lower[26] );
tran (\sa_snapshot[13][27] , \sa_snapshot[13].r.part0[27] );
tran (\sa_snapshot[13][27] , \sa_snapshot[13].f.lower[27] );
tran (\sa_snapshot[13][28] , \sa_snapshot[13].r.part0[28] );
tran (\sa_snapshot[13][28] , \sa_snapshot[13].f.lower[28] );
tran (\sa_snapshot[13][29] , \sa_snapshot[13].r.part0[29] );
tran (\sa_snapshot[13][29] , \sa_snapshot[13].f.lower[29] );
tran (\sa_snapshot[13][30] , \sa_snapshot[13].r.part0[30] );
tran (\sa_snapshot[13][30] , \sa_snapshot[13].f.lower[30] );
tran (\sa_snapshot[13][31] , \sa_snapshot[13].r.part0[31] );
tran (\sa_snapshot[13][31] , \sa_snapshot[13].f.lower[31] );
tran (\sa_snapshot[13][32] , \sa_snapshot[13].r.part1[0] );
tran (\sa_snapshot[13][32] , \sa_snapshot[13].f.upper[0] );
tran (\sa_snapshot[13][33] , \sa_snapshot[13].r.part1[1] );
tran (\sa_snapshot[13][33] , \sa_snapshot[13].f.upper[1] );
tran (\sa_snapshot[13][34] , \sa_snapshot[13].r.part1[2] );
tran (\sa_snapshot[13][34] , \sa_snapshot[13].f.upper[2] );
tran (\sa_snapshot[13][35] , \sa_snapshot[13].r.part1[3] );
tran (\sa_snapshot[13][35] , \sa_snapshot[13].f.upper[3] );
tran (\sa_snapshot[13][36] , \sa_snapshot[13].r.part1[4] );
tran (\sa_snapshot[13][36] , \sa_snapshot[13].f.upper[4] );
tran (\sa_snapshot[13][37] , \sa_snapshot[13].r.part1[5] );
tran (\sa_snapshot[13][37] , \sa_snapshot[13].f.upper[5] );
tran (\sa_snapshot[13][38] , \sa_snapshot[13].r.part1[6] );
tran (\sa_snapshot[13][38] , \sa_snapshot[13].f.upper[6] );
tran (\sa_snapshot[13][39] , \sa_snapshot[13].r.part1[7] );
tran (\sa_snapshot[13][39] , \sa_snapshot[13].f.upper[7] );
tran (\sa_snapshot[13][40] , \sa_snapshot[13].r.part1[8] );
tran (\sa_snapshot[13][40] , \sa_snapshot[13].f.upper[8] );
tran (\sa_snapshot[13][41] , \sa_snapshot[13].r.part1[9] );
tran (\sa_snapshot[13][41] , \sa_snapshot[13].f.upper[9] );
tran (\sa_snapshot[13][42] , \sa_snapshot[13].r.part1[10] );
tran (\sa_snapshot[13][42] , \sa_snapshot[13].f.upper[10] );
tran (\sa_snapshot[13][43] , \sa_snapshot[13].r.part1[11] );
tran (\sa_snapshot[13][43] , \sa_snapshot[13].f.upper[11] );
tran (\sa_snapshot[13][44] , \sa_snapshot[13].r.part1[12] );
tran (\sa_snapshot[13][44] , \sa_snapshot[13].f.upper[12] );
tran (\sa_snapshot[13][45] , \sa_snapshot[13].r.part1[13] );
tran (\sa_snapshot[13][45] , \sa_snapshot[13].f.upper[13] );
tran (\sa_snapshot[13][46] , \sa_snapshot[13].r.part1[14] );
tran (\sa_snapshot[13][46] , \sa_snapshot[13].f.upper[14] );
tran (\sa_snapshot[13][47] , \sa_snapshot[13].r.part1[15] );
tran (\sa_snapshot[13][47] , \sa_snapshot[13].f.upper[15] );
tran (\sa_snapshot[13][48] , \sa_snapshot[13].r.part1[16] );
tran (\sa_snapshot[13][48] , \sa_snapshot[13].f.upper[16] );
tran (\sa_snapshot[13][49] , \sa_snapshot[13].r.part1[17] );
tran (\sa_snapshot[13][49] , \sa_snapshot[13].f.upper[17] );
tran (\sa_snapshot[13][50] , \sa_snapshot[13].r.part1[18] );
tran (\sa_snapshot[13][50] , \sa_snapshot[13].f.unused[0] );
tran (\sa_snapshot[13][51] , \sa_snapshot[13].r.part1[19] );
tran (\sa_snapshot[13][51] , \sa_snapshot[13].f.unused[1] );
tran (\sa_snapshot[13][52] , \sa_snapshot[13].r.part1[20] );
tran (\sa_snapshot[13][52] , \sa_snapshot[13].f.unused[2] );
tran (\sa_snapshot[13][53] , \sa_snapshot[13].r.part1[21] );
tran (\sa_snapshot[13][53] , \sa_snapshot[13].f.unused[3] );
tran (\sa_snapshot[13][54] , \sa_snapshot[13].r.part1[22] );
tran (\sa_snapshot[13][54] , \sa_snapshot[13].f.unused[4] );
tran (\sa_snapshot[13][55] , \sa_snapshot[13].r.part1[23] );
tran (\sa_snapshot[13][55] , \sa_snapshot[13].f.unused[5] );
tran (\sa_snapshot[13][56] , \sa_snapshot[13].r.part1[24] );
tran (\sa_snapshot[13][56] , \sa_snapshot[13].f.unused[6] );
tran (\sa_snapshot[13][57] , \sa_snapshot[13].r.part1[25] );
tran (\sa_snapshot[13][57] , \sa_snapshot[13].f.unused[7] );
tran (\sa_snapshot[13][58] , \sa_snapshot[13].r.part1[26] );
tran (\sa_snapshot[13][58] , \sa_snapshot[13].f.unused[8] );
tran (\sa_snapshot[13][59] , \sa_snapshot[13].r.part1[27] );
tran (\sa_snapshot[13][59] , \sa_snapshot[13].f.unused[9] );
tran (\sa_snapshot[13][60] , \sa_snapshot[13].r.part1[28] );
tran (\sa_snapshot[13][60] , \sa_snapshot[13].f.unused[10] );
tran (\sa_snapshot[13][61] , \sa_snapshot[13].r.part1[29] );
tran (\sa_snapshot[13][61] , \sa_snapshot[13].f.unused[11] );
tran (\sa_snapshot[13][62] , \sa_snapshot[13].r.part1[30] );
tran (\sa_snapshot[13][62] , \sa_snapshot[13].f.unused[12] );
tran (\sa_snapshot[13][63] , \sa_snapshot[13].r.part1[31] );
tran (\sa_snapshot[13][63] , \sa_snapshot[13].f.unused[13] );
tran (\sa_snapshot[14][0] , \sa_snapshot[14].r.part0[0] );
tran (\sa_snapshot[14][0] , \sa_snapshot[14].f.lower[0] );
tran (\sa_snapshot[14][1] , \sa_snapshot[14].r.part0[1] );
tran (\sa_snapshot[14][1] , \sa_snapshot[14].f.lower[1] );
tran (\sa_snapshot[14][2] , \sa_snapshot[14].r.part0[2] );
tran (\sa_snapshot[14][2] , \sa_snapshot[14].f.lower[2] );
tran (\sa_snapshot[14][3] , \sa_snapshot[14].r.part0[3] );
tran (\sa_snapshot[14][3] , \sa_snapshot[14].f.lower[3] );
tran (\sa_snapshot[14][4] , \sa_snapshot[14].r.part0[4] );
tran (\sa_snapshot[14][4] , \sa_snapshot[14].f.lower[4] );
tran (\sa_snapshot[14][5] , \sa_snapshot[14].r.part0[5] );
tran (\sa_snapshot[14][5] , \sa_snapshot[14].f.lower[5] );
tran (\sa_snapshot[14][6] , \sa_snapshot[14].r.part0[6] );
tran (\sa_snapshot[14][6] , \sa_snapshot[14].f.lower[6] );
tran (\sa_snapshot[14][7] , \sa_snapshot[14].r.part0[7] );
tran (\sa_snapshot[14][7] , \sa_snapshot[14].f.lower[7] );
tran (\sa_snapshot[14][8] , \sa_snapshot[14].r.part0[8] );
tran (\sa_snapshot[14][8] , \sa_snapshot[14].f.lower[8] );
tran (\sa_snapshot[14][9] , \sa_snapshot[14].r.part0[9] );
tran (\sa_snapshot[14][9] , \sa_snapshot[14].f.lower[9] );
tran (\sa_snapshot[14][10] , \sa_snapshot[14].r.part0[10] );
tran (\sa_snapshot[14][10] , \sa_snapshot[14].f.lower[10] );
tran (\sa_snapshot[14][11] , \sa_snapshot[14].r.part0[11] );
tran (\sa_snapshot[14][11] , \sa_snapshot[14].f.lower[11] );
tran (\sa_snapshot[14][12] , \sa_snapshot[14].r.part0[12] );
tran (\sa_snapshot[14][12] , \sa_snapshot[14].f.lower[12] );
tran (\sa_snapshot[14][13] , \sa_snapshot[14].r.part0[13] );
tran (\sa_snapshot[14][13] , \sa_snapshot[14].f.lower[13] );
tran (\sa_snapshot[14][14] , \sa_snapshot[14].r.part0[14] );
tran (\sa_snapshot[14][14] , \sa_snapshot[14].f.lower[14] );
tran (\sa_snapshot[14][15] , \sa_snapshot[14].r.part0[15] );
tran (\sa_snapshot[14][15] , \sa_snapshot[14].f.lower[15] );
tran (\sa_snapshot[14][16] , \sa_snapshot[14].r.part0[16] );
tran (\sa_snapshot[14][16] , \sa_snapshot[14].f.lower[16] );
tran (\sa_snapshot[14][17] , \sa_snapshot[14].r.part0[17] );
tran (\sa_snapshot[14][17] , \sa_snapshot[14].f.lower[17] );
tran (\sa_snapshot[14][18] , \sa_snapshot[14].r.part0[18] );
tran (\sa_snapshot[14][18] , \sa_snapshot[14].f.lower[18] );
tran (\sa_snapshot[14][19] , \sa_snapshot[14].r.part0[19] );
tran (\sa_snapshot[14][19] , \sa_snapshot[14].f.lower[19] );
tran (\sa_snapshot[14][20] , \sa_snapshot[14].r.part0[20] );
tran (\sa_snapshot[14][20] , \sa_snapshot[14].f.lower[20] );
tran (\sa_snapshot[14][21] , \sa_snapshot[14].r.part0[21] );
tran (\sa_snapshot[14][21] , \sa_snapshot[14].f.lower[21] );
tran (\sa_snapshot[14][22] , \sa_snapshot[14].r.part0[22] );
tran (\sa_snapshot[14][22] , \sa_snapshot[14].f.lower[22] );
tran (\sa_snapshot[14][23] , \sa_snapshot[14].r.part0[23] );
tran (\sa_snapshot[14][23] , \sa_snapshot[14].f.lower[23] );
tran (\sa_snapshot[14][24] , \sa_snapshot[14].r.part0[24] );
tran (\sa_snapshot[14][24] , \sa_snapshot[14].f.lower[24] );
tran (\sa_snapshot[14][25] , \sa_snapshot[14].r.part0[25] );
tran (\sa_snapshot[14][25] , \sa_snapshot[14].f.lower[25] );
tran (\sa_snapshot[14][26] , \sa_snapshot[14].r.part0[26] );
tran (\sa_snapshot[14][26] , \sa_snapshot[14].f.lower[26] );
tran (\sa_snapshot[14][27] , \sa_snapshot[14].r.part0[27] );
tran (\sa_snapshot[14][27] , \sa_snapshot[14].f.lower[27] );
tran (\sa_snapshot[14][28] , \sa_snapshot[14].r.part0[28] );
tran (\sa_snapshot[14][28] , \sa_snapshot[14].f.lower[28] );
tran (\sa_snapshot[14][29] , \sa_snapshot[14].r.part0[29] );
tran (\sa_snapshot[14][29] , \sa_snapshot[14].f.lower[29] );
tran (\sa_snapshot[14][30] , \sa_snapshot[14].r.part0[30] );
tran (\sa_snapshot[14][30] , \sa_snapshot[14].f.lower[30] );
tran (\sa_snapshot[14][31] , \sa_snapshot[14].r.part0[31] );
tran (\sa_snapshot[14][31] , \sa_snapshot[14].f.lower[31] );
tran (\sa_snapshot[14][32] , \sa_snapshot[14].r.part1[0] );
tran (\sa_snapshot[14][32] , \sa_snapshot[14].f.upper[0] );
tran (\sa_snapshot[14][33] , \sa_snapshot[14].r.part1[1] );
tran (\sa_snapshot[14][33] , \sa_snapshot[14].f.upper[1] );
tran (\sa_snapshot[14][34] , \sa_snapshot[14].r.part1[2] );
tran (\sa_snapshot[14][34] , \sa_snapshot[14].f.upper[2] );
tran (\sa_snapshot[14][35] , \sa_snapshot[14].r.part1[3] );
tran (\sa_snapshot[14][35] , \sa_snapshot[14].f.upper[3] );
tran (\sa_snapshot[14][36] , \sa_snapshot[14].r.part1[4] );
tran (\sa_snapshot[14][36] , \sa_snapshot[14].f.upper[4] );
tran (\sa_snapshot[14][37] , \sa_snapshot[14].r.part1[5] );
tran (\sa_snapshot[14][37] , \sa_snapshot[14].f.upper[5] );
tran (\sa_snapshot[14][38] , \sa_snapshot[14].r.part1[6] );
tran (\sa_snapshot[14][38] , \sa_snapshot[14].f.upper[6] );
tran (\sa_snapshot[14][39] , \sa_snapshot[14].r.part1[7] );
tran (\sa_snapshot[14][39] , \sa_snapshot[14].f.upper[7] );
tran (\sa_snapshot[14][40] , \sa_snapshot[14].r.part1[8] );
tran (\sa_snapshot[14][40] , \sa_snapshot[14].f.upper[8] );
tran (\sa_snapshot[14][41] , \sa_snapshot[14].r.part1[9] );
tran (\sa_snapshot[14][41] , \sa_snapshot[14].f.upper[9] );
tran (\sa_snapshot[14][42] , \sa_snapshot[14].r.part1[10] );
tran (\sa_snapshot[14][42] , \sa_snapshot[14].f.upper[10] );
tran (\sa_snapshot[14][43] , \sa_snapshot[14].r.part1[11] );
tran (\sa_snapshot[14][43] , \sa_snapshot[14].f.upper[11] );
tran (\sa_snapshot[14][44] , \sa_snapshot[14].r.part1[12] );
tran (\sa_snapshot[14][44] , \sa_snapshot[14].f.upper[12] );
tran (\sa_snapshot[14][45] , \sa_snapshot[14].r.part1[13] );
tran (\sa_snapshot[14][45] , \sa_snapshot[14].f.upper[13] );
tran (\sa_snapshot[14][46] , \sa_snapshot[14].r.part1[14] );
tran (\sa_snapshot[14][46] , \sa_snapshot[14].f.upper[14] );
tran (\sa_snapshot[14][47] , \sa_snapshot[14].r.part1[15] );
tran (\sa_snapshot[14][47] , \sa_snapshot[14].f.upper[15] );
tran (\sa_snapshot[14][48] , \sa_snapshot[14].r.part1[16] );
tran (\sa_snapshot[14][48] , \sa_snapshot[14].f.upper[16] );
tran (\sa_snapshot[14][49] , \sa_snapshot[14].r.part1[17] );
tran (\sa_snapshot[14][49] , \sa_snapshot[14].f.upper[17] );
tran (\sa_snapshot[14][50] , \sa_snapshot[14].r.part1[18] );
tran (\sa_snapshot[14][50] , \sa_snapshot[14].f.unused[0] );
tran (\sa_snapshot[14][51] , \sa_snapshot[14].r.part1[19] );
tran (\sa_snapshot[14][51] , \sa_snapshot[14].f.unused[1] );
tran (\sa_snapshot[14][52] , \sa_snapshot[14].r.part1[20] );
tran (\sa_snapshot[14][52] , \sa_snapshot[14].f.unused[2] );
tran (\sa_snapshot[14][53] , \sa_snapshot[14].r.part1[21] );
tran (\sa_snapshot[14][53] , \sa_snapshot[14].f.unused[3] );
tran (\sa_snapshot[14][54] , \sa_snapshot[14].r.part1[22] );
tran (\sa_snapshot[14][54] , \sa_snapshot[14].f.unused[4] );
tran (\sa_snapshot[14][55] , \sa_snapshot[14].r.part1[23] );
tran (\sa_snapshot[14][55] , \sa_snapshot[14].f.unused[5] );
tran (\sa_snapshot[14][56] , \sa_snapshot[14].r.part1[24] );
tran (\sa_snapshot[14][56] , \sa_snapshot[14].f.unused[6] );
tran (\sa_snapshot[14][57] , \sa_snapshot[14].r.part1[25] );
tran (\sa_snapshot[14][57] , \sa_snapshot[14].f.unused[7] );
tran (\sa_snapshot[14][58] , \sa_snapshot[14].r.part1[26] );
tran (\sa_snapshot[14][58] , \sa_snapshot[14].f.unused[8] );
tran (\sa_snapshot[14][59] , \sa_snapshot[14].r.part1[27] );
tran (\sa_snapshot[14][59] , \sa_snapshot[14].f.unused[9] );
tran (\sa_snapshot[14][60] , \sa_snapshot[14].r.part1[28] );
tran (\sa_snapshot[14][60] , \sa_snapshot[14].f.unused[10] );
tran (\sa_snapshot[14][61] , \sa_snapshot[14].r.part1[29] );
tran (\sa_snapshot[14][61] , \sa_snapshot[14].f.unused[11] );
tran (\sa_snapshot[14][62] , \sa_snapshot[14].r.part1[30] );
tran (\sa_snapshot[14][62] , \sa_snapshot[14].f.unused[12] );
tran (\sa_snapshot[14][63] , \sa_snapshot[14].r.part1[31] );
tran (\sa_snapshot[14][63] , \sa_snapshot[14].f.unused[13] );
tran (\sa_snapshot[15][0] , \sa_snapshot[15].r.part0[0] );
tran (\sa_snapshot[15][0] , \sa_snapshot[15].f.lower[0] );
tran (\sa_snapshot[15][1] , \sa_snapshot[15].r.part0[1] );
tran (\sa_snapshot[15][1] , \sa_snapshot[15].f.lower[1] );
tran (\sa_snapshot[15][2] , \sa_snapshot[15].r.part0[2] );
tran (\sa_snapshot[15][2] , \sa_snapshot[15].f.lower[2] );
tran (\sa_snapshot[15][3] , \sa_snapshot[15].r.part0[3] );
tran (\sa_snapshot[15][3] , \sa_snapshot[15].f.lower[3] );
tran (\sa_snapshot[15][4] , \sa_snapshot[15].r.part0[4] );
tran (\sa_snapshot[15][4] , \sa_snapshot[15].f.lower[4] );
tran (\sa_snapshot[15][5] , \sa_snapshot[15].r.part0[5] );
tran (\sa_snapshot[15][5] , \sa_snapshot[15].f.lower[5] );
tran (\sa_snapshot[15][6] , \sa_snapshot[15].r.part0[6] );
tran (\sa_snapshot[15][6] , \sa_snapshot[15].f.lower[6] );
tran (\sa_snapshot[15][7] , \sa_snapshot[15].r.part0[7] );
tran (\sa_snapshot[15][7] , \sa_snapshot[15].f.lower[7] );
tran (\sa_snapshot[15][8] , \sa_snapshot[15].r.part0[8] );
tran (\sa_snapshot[15][8] , \sa_snapshot[15].f.lower[8] );
tran (\sa_snapshot[15][9] , \sa_snapshot[15].r.part0[9] );
tran (\sa_snapshot[15][9] , \sa_snapshot[15].f.lower[9] );
tran (\sa_snapshot[15][10] , \sa_snapshot[15].r.part0[10] );
tran (\sa_snapshot[15][10] , \sa_snapshot[15].f.lower[10] );
tran (\sa_snapshot[15][11] , \sa_snapshot[15].r.part0[11] );
tran (\sa_snapshot[15][11] , \sa_snapshot[15].f.lower[11] );
tran (\sa_snapshot[15][12] , \sa_snapshot[15].r.part0[12] );
tran (\sa_snapshot[15][12] , \sa_snapshot[15].f.lower[12] );
tran (\sa_snapshot[15][13] , \sa_snapshot[15].r.part0[13] );
tran (\sa_snapshot[15][13] , \sa_snapshot[15].f.lower[13] );
tran (\sa_snapshot[15][14] , \sa_snapshot[15].r.part0[14] );
tran (\sa_snapshot[15][14] , \sa_snapshot[15].f.lower[14] );
tran (\sa_snapshot[15][15] , \sa_snapshot[15].r.part0[15] );
tran (\sa_snapshot[15][15] , \sa_snapshot[15].f.lower[15] );
tran (\sa_snapshot[15][16] , \sa_snapshot[15].r.part0[16] );
tran (\sa_snapshot[15][16] , \sa_snapshot[15].f.lower[16] );
tran (\sa_snapshot[15][17] , \sa_snapshot[15].r.part0[17] );
tran (\sa_snapshot[15][17] , \sa_snapshot[15].f.lower[17] );
tran (\sa_snapshot[15][18] , \sa_snapshot[15].r.part0[18] );
tran (\sa_snapshot[15][18] , \sa_snapshot[15].f.lower[18] );
tran (\sa_snapshot[15][19] , \sa_snapshot[15].r.part0[19] );
tran (\sa_snapshot[15][19] , \sa_snapshot[15].f.lower[19] );
tran (\sa_snapshot[15][20] , \sa_snapshot[15].r.part0[20] );
tran (\sa_snapshot[15][20] , \sa_snapshot[15].f.lower[20] );
tran (\sa_snapshot[15][21] , \sa_snapshot[15].r.part0[21] );
tran (\sa_snapshot[15][21] , \sa_snapshot[15].f.lower[21] );
tran (\sa_snapshot[15][22] , \sa_snapshot[15].r.part0[22] );
tran (\sa_snapshot[15][22] , \sa_snapshot[15].f.lower[22] );
tran (\sa_snapshot[15][23] , \sa_snapshot[15].r.part0[23] );
tran (\sa_snapshot[15][23] , \sa_snapshot[15].f.lower[23] );
tran (\sa_snapshot[15][24] , \sa_snapshot[15].r.part0[24] );
tran (\sa_snapshot[15][24] , \sa_snapshot[15].f.lower[24] );
tran (\sa_snapshot[15][25] , \sa_snapshot[15].r.part0[25] );
tran (\sa_snapshot[15][25] , \sa_snapshot[15].f.lower[25] );
tran (\sa_snapshot[15][26] , \sa_snapshot[15].r.part0[26] );
tran (\sa_snapshot[15][26] , \sa_snapshot[15].f.lower[26] );
tran (\sa_snapshot[15][27] , \sa_snapshot[15].r.part0[27] );
tran (\sa_snapshot[15][27] , \sa_snapshot[15].f.lower[27] );
tran (\sa_snapshot[15][28] , \sa_snapshot[15].r.part0[28] );
tran (\sa_snapshot[15][28] , \sa_snapshot[15].f.lower[28] );
tran (\sa_snapshot[15][29] , \sa_snapshot[15].r.part0[29] );
tran (\sa_snapshot[15][29] , \sa_snapshot[15].f.lower[29] );
tran (\sa_snapshot[15][30] , \sa_snapshot[15].r.part0[30] );
tran (\sa_snapshot[15][30] , \sa_snapshot[15].f.lower[30] );
tran (\sa_snapshot[15][31] , \sa_snapshot[15].r.part0[31] );
tran (\sa_snapshot[15][31] , \sa_snapshot[15].f.lower[31] );
tran (\sa_snapshot[15][32] , \sa_snapshot[15].r.part1[0] );
tran (\sa_snapshot[15][32] , \sa_snapshot[15].f.upper[0] );
tran (\sa_snapshot[15][33] , \sa_snapshot[15].r.part1[1] );
tran (\sa_snapshot[15][33] , \sa_snapshot[15].f.upper[1] );
tran (\sa_snapshot[15][34] , \sa_snapshot[15].r.part1[2] );
tran (\sa_snapshot[15][34] , \sa_snapshot[15].f.upper[2] );
tran (\sa_snapshot[15][35] , \sa_snapshot[15].r.part1[3] );
tran (\sa_snapshot[15][35] , \sa_snapshot[15].f.upper[3] );
tran (\sa_snapshot[15][36] , \sa_snapshot[15].r.part1[4] );
tran (\sa_snapshot[15][36] , \sa_snapshot[15].f.upper[4] );
tran (\sa_snapshot[15][37] , \sa_snapshot[15].r.part1[5] );
tran (\sa_snapshot[15][37] , \sa_snapshot[15].f.upper[5] );
tran (\sa_snapshot[15][38] , \sa_snapshot[15].r.part1[6] );
tran (\sa_snapshot[15][38] , \sa_snapshot[15].f.upper[6] );
tran (\sa_snapshot[15][39] , \sa_snapshot[15].r.part1[7] );
tran (\sa_snapshot[15][39] , \sa_snapshot[15].f.upper[7] );
tran (\sa_snapshot[15][40] , \sa_snapshot[15].r.part1[8] );
tran (\sa_snapshot[15][40] , \sa_snapshot[15].f.upper[8] );
tran (\sa_snapshot[15][41] , \sa_snapshot[15].r.part1[9] );
tran (\sa_snapshot[15][41] , \sa_snapshot[15].f.upper[9] );
tran (\sa_snapshot[15][42] , \sa_snapshot[15].r.part1[10] );
tran (\sa_snapshot[15][42] , \sa_snapshot[15].f.upper[10] );
tran (\sa_snapshot[15][43] , \sa_snapshot[15].r.part1[11] );
tran (\sa_snapshot[15][43] , \sa_snapshot[15].f.upper[11] );
tran (\sa_snapshot[15][44] , \sa_snapshot[15].r.part1[12] );
tran (\sa_snapshot[15][44] , \sa_snapshot[15].f.upper[12] );
tran (\sa_snapshot[15][45] , \sa_snapshot[15].r.part1[13] );
tran (\sa_snapshot[15][45] , \sa_snapshot[15].f.upper[13] );
tran (\sa_snapshot[15][46] , \sa_snapshot[15].r.part1[14] );
tran (\sa_snapshot[15][46] , \sa_snapshot[15].f.upper[14] );
tran (\sa_snapshot[15][47] , \sa_snapshot[15].r.part1[15] );
tran (\sa_snapshot[15][47] , \sa_snapshot[15].f.upper[15] );
tran (\sa_snapshot[15][48] , \sa_snapshot[15].r.part1[16] );
tran (\sa_snapshot[15][48] , \sa_snapshot[15].f.upper[16] );
tran (\sa_snapshot[15][49] , \sa_snapshot[15].r.part1[17] );
tran (\sa_snapshot[15][49] , \sa_snapshot[15].f.upper[17] );
tran (\sa_snapshot[15][50] , \sa_snapshot[15].r.part1[18] );
tran (\sa_snapshot[15][50] , \sa_snapshot[15].f.unused[0] );
tran (\sa_snapshot[15][51] , \sa_snapshot[15].r.part1[19] );
tran (\sa_snapshot[15][51] , \sa_snapshot[15].f.unused[1] );
tran (\sa_snapshot[15][52] , \sa_snapshot[15].r.part1[20] );
tran (\sa_snapshot[15][52] , \sa_snapshot[15].f.unused[2] );
tran (\sa_snapshot[15][53] , \sa_snapshot[15].r.part1[21] );
tran (\sa_snapshot[15][53] , \sa_snapshot[15].f.unused[3] );
tran (\sa_snapshot[15][54] , \sa_snapshot[15].r.part1[22] );
tran (\sa_snapshot[15][54] , \sa_snapshot[15].f.unused[4] );
tran (\sa_snapshot[15][55] , \sa_snapshot[15].r.part1[23] );
tran (\sa_snapshot[15][55] , \sa_snapshot[15].f.unused[5] );
tran (\sa_snapshot[15][56] , \sa_snapshot[15].r.part1[24] );
tran (\sa_snapshot[15][56] , \sa_snapshot[15].f.unused[6] );
tran (\sa_snapshot[15][57] , \sa_snapshot[15].r.part1[25] );
tran (\sa_snapshot[15][57] , \sa_snapshot[15].f.unused[7] );
tran (\sa_snapshot[15][58] , \sa_snapshot[15].r.part1[26] );
tran (\sa_snapshot[15][58] , \sa_snapshot[15].f.unused[8] );
tran (\sa_snapshot[15][59] , \sa_snapshot[15].r.part1[27] );
tran (\sa_snapshot[15][59] , \sa_snapshot[15].f.unused[9] );
tran (\sa_snapshot[15][60] , \sa_snapshot[15].r.part1[28] );
tran (\sa_snapshot[15][60] , \sa_snapshot[15].f.unused[10] );
tran (\sa_snapshot[15][61] , \sa_snapshot[15].r.part1[29] );
tran (\sa_snapshot[15][61] , \sa_snapshot[15].f.unused[11] );
tran (\sa_snapshot[15][62] , \sa_snapshot[15].r.part1[30] );
tran (\sa_snapshot[15][62] , \sa_snapshot[15].f.unused[12] );
tran (\sa_snapshot[15][63] , \sa_snapshot[15].r.part1[31] );
tran (\sa_snapshot[15][63] , \sa_snapshot[15].f.unused[13] );
tran (\sa_snapshot[16][0] , \sa_snapshot[16].r.part0[0] );
tran (\sa_snapshot[16][0] , \sa_snapshot[16].f.lower[0] );
tran (\sa_snapshot[16][1] , \sa_snapshot[16].r.part0[1] );
tran (\sa_snapshot[16][1] , \sa_snapshot[16].f.lower[1] );
tran (\sa_snapshot[16][2] , \sa_snapshot[16].r.part0[2] );
tran (\sa_snapshot[16][2] , \sa_snapshot[16].f.lower[2] );
tran (\sa_snapshot[16][3] , \sa_snapshot[16].r.part0[3] );
tran (\sa_snapshot[16][3] , \sa_snapshot[16].f.lower[3] );
tran (\sa_snapshot[16][4] , \sa_snapshot[16].r.part0[4] );
tran (\sa_snapshot[16][4] , \sa_snapshot[16].f.lower[4] );
tran (\sa_snapshot[16][5] , \sa_snapshot[16].r.part0[5] );
tran (\sa_snapshot[16][5] , \sa_snapshot[16].f.lower[5] );
tran (\sa_snapshot[16][6] , \sa_snapshot[16].r.part0[6] );
tran (\sa_snapshot[16][6] , \sa_snapshot[16].f.lower[6] );
tran (\sa_snapshot[16][7] , \sa_snapshot[16].r.part0[7] );
tran (\sa_snapshot[16][7] , \sa_snapshot[16].f.lower[7] );
tran (\sa_snapshot[16][8] , \sa_snapshot[16].r.part0[8] );
tran (\sa_snapshot[16][8] , \sa_snapshot[16].f.lower[8] );
tran (\sa_snapshot[16][9] , \sa_snapshot[16].r.part0[9] );
tran (\sa_snapshot[16][9] , \sa_snapshot[16].f.lower[9] );
tran (\sa_snapshot[16][10] , \sa_snapshot[16].r.part0[10] );
tran (\sa_snapshot[16][10] , \sa_snapshot[16].f.lower[10] );
tran (\sa_snapshot[16][11] , \sa_snapshot[16].r.part0[11] );
tran (\sa_snapshot[16][11] , \sa_snapshot[16].f.lower[11] );
tran (\sa_snapshot[16][12] , \sa_snapshot[16].r.part0[12] );
tran (\sa_snapshot[16][12] , \sa_snapshot[16].f.lower[12] );
tran (\sa_snapshot[16][13] , \sa_snapshot[16].r.part0[13] );
tran (\sa_snapshot[16][13] , \sa_snapshot[16].f.lower[13] );
tran (\sa_snapshot[16][14] , \sa_snapshot[16].r.part0[14] );
tran (\sa_snapshot[16][14] , \sa_snapshot[16].f.lower[14] );
tran (\sa_snapshot[16][15] , \sa_snapshot[16].r.part0[15] );
tran (\sa_snapshot[16][15] , \sa_snapshot[16].f.lower[15] );
tran (\sa_snapshot[16][16] , \sa_snapshot[16].r.part0[16] );
tran (\sa_snapshot[16][16] , \sa_snapshot[16].f.lower[16] );
tran (\sa_snapshot[16][17] , \sa_snapshot[16].r.part0[17] );
tran (\sa_snapshot[16][17] , \sa_snapshot[16].f.lower[17] );
tran (\sa_snapshot[16][18] , \sa_snapshot[16].r.part0[18] );
tran (\sa_snapshot[16][18] , \sa_snapshot[16].f.lower[18] );
tran (\sa_snapshot[16][19] , \sa_snapshot[16].r.part0[19] );
tran (\sa_snapshot[16][19] , \sa_snapshot[16].f.lower[19] );
tran (\sa_snapshot[16][20] , \sa_snapshot[16].r.part0[20] );
tran (\sa_snapshot[16][20] , \sa_snapshot[16].f.lower[20] );
tran (\sa_snapshot[16][21] , \sa_snapshot[16].r.part0[21] );
tran (\sa_snapshot[16][21] , \sa_snapshot[16].f.lower[21] );
tran (\sa_snapshot[16][22] , \sa_snapshot[16].r.part0[22] );
tran (\sa_snapshot[16][22] , \sa_snapshot[16].f.lower[22] );
tran (\sa_snapshot[16][23] , \sa_snapshot[16].r.part0[23] );
tran (\sa_snapshot[16][23] , \sa_snapshot[16].f.lower[23] );
tran (\sa_snapshot[16][24] , \sa_snapshot[16].r.part0[24] );
tran (\sa_snapshot[16][24] , \sa_snapshot[16].f.lower[24] );
tran (\sa_snapshot[16][25] , \sa_snapshot[16].r.part0[25] );
tran (\sa_snapshot[16][25] , \sa_snapshot[16].f.lower[25] );
tran (\sa_snapshot[16][26] , \sa_snapshot[16].r.part0[26] );
tran (\sa_snapshot[16][26] , \sa_snapshot[16].f.lower[26] );
tran (\sa_snapshot[16][27] , \sa_snapshot[16].r.part0[27] );
tran (\sa_snapshot[16][27] , \sa_snapshot[16].f.lower[27] );
tran (\sa_snapshot[16][28] , \sa_snapshot[16].r.part0[28] );
tran (\sa_snapshot[16][28] , \sa_snapshot[16].f.lower[28] );
tran (\sa_snapshot[16][29] , \sa_snapshot[16].r.part0[29] );
tran (\sa_snapshot[16][29] , \sa_snapshot[16].f.lower[29] );
tran (\sa_snapshot[16][30] , \sa_snapshot[16].r.part0[30] );
tran (\sa_snapshot[16][30] , \sa_snapshot[16].f.lower[30] );
tran (\sa_snapshot[16][31] , \sa_snapshot[16].r.part0[31] );
tran (\sa_snapshot[16][31] , \sa_snapshot[16].f.lower[31] );
tran (\sa_snapshot[16][32] , \sa_snapshot[16].r.part1[0] );
tran (\sa_snapshot[16][32] , \sa_snapshot[16].f.upper[0] );
tran (\sa_snapshot[16][33] , \sa_snapshot[16].r.part1[1] );
tran (\sa_snapshot[16][33] , \sa_snapshot[16].f.upper[1] );
tran (\sa_snapshot[16][34] , \sa_snapshot[16].r.part1[2] );
tran (\sa_snapshot[16][34] , \sa_snapshot[16].f.upper[2] );
tran (\sa_snapshot[16][35] , \sa_snapshot[16].r.part1[3] );
tran (\sa_snapshot[16][35] , \sa_snapshot[16].f.upper[3] );
tran (\sa_snapshot[16][36] , \sa_snapshot[16].r.part1[4] );
tran (\sa_snapshot[16][36] , \sa_snapshot[16].f.upper[4] );
tran (\sa_snapshot[16][37] , \sa_snapshot[16].r.part1[5] );
tran (\sa_snapshot[16][37] , \sa_snapshot[16].f.upper[5] );
tran (\sa_snapshot[16][38] , \sa_snapshot[16].r.part1[6] );
tran (\sa_snapshot[16][38] , \sa_snapshot[16].f.upper[6] );
tran (\sa_snapshot[16][39] , \sa_snapshot[16].r.part1[7] );
tran (\sa_snapshot[16][39] , \sa_snapshot[16].f.upper[7] );
tran (\sa_snapshot[16][40] , \sa_snapshot[16].r.part1[8] );
tran (\sa_snapshot[16][40] , \sa_snapshot[16].f.upper[8] );
tran (\sa_snapshot[16][41] , \sa_snapshot[16].r.part1[9] );
tran (\sa_snapshot[16][41] , \sa_snapshot[16].f.upper[9] );
tran (\sa_snapshot[16][42] , \sa_snapshot[16].r.part1[10] );
tran (\sa_snapshot[16][42] , \sa_snapshot[16].f.upper[10] );
tran (\sa_snapshot[16][43] , \sa_snapshot[16].r.part1[11] );
tran (\sa_snapshot[16][43] , \sa_snapshot[16].f.upper[11] );
tran (\sa_snapshot[16][44] , \sa_snapshot[16].r.part1[12] );
tran (\sa_snapshot[16][44] , \sa_snapshot[16].f.upper[12] );
tran (\sa_snapshot[16][45] , \sa_snapshot[16].r.part1[13] );
tran (\sa_snapshot[16][45] , \sa_snapshot[16].f.upper[13] );
tran (\sa_snapshot[16][46] , \sa_snapshot[16].r.part1[14] );
tran (\sa_snapshot[16][46] , \sa_snapshot[16].f.upper[14] );
tran (\sa_snapshot[16][47] , \sa_snapshot[16].r.part1[15] );
tran (\sa_snapshot[16][47] , \sa_snapshot[16].f.upper[15] );
tran (\sa_snapshot[16][48] , \sa_snapshot[16].r.part1[16] );
tran (\sa_snapshot[16][48] , \sa_snapshot[16].f.upper[16] );
tran (\sa_snapshot[16][49] , \sa_snapshot[16].r.part1[17] );
tran (\sa_snapshot[16][49] , \sa_snapshot[16].f.upper[17] );
tran (\sa_snapshot[16][50] , \sa_snapshot[16].r.part1[18] );
tran (\sa_snapshot[16][50] , \sa_snapshot[16].f.unused[0] );
tran (\sa_snapshot[16][51] , \sa_snapshot[16].r.part1[19] );
tran (\sa_snapshot[16][51] , \sa_snapshot[16].f.unused[1] );
tran (\sa_snapshot[16][52] , \sa_snapshot[16].r.part1[20] );
tran (\sa_snapshot[16][52] , \sa_snapshot[16].f.unused[2] );
tran (\sa_snapshot[16][53] , \sa_snapshot[16].r.part1[21] );
tran (\sa_snapshot[16][53] , \sa_snapshot[16].f.unused[3] );
tran (\sa_snapshot[16][54] , \sa_snapshot[16].r.part1[22] );
tran (\sa_snapshot[16][54] , \sa_snapshot[16].f.unused[4] );
tran (\sa_snapshot[16][55] , \sa_snapshot[16].r.part1[23] );
tran (\sa_snapshot[16][55] , \sa_snapshot[16].f.unused[5] );
tran (\sa_snapshot[16][56] , \sa_snapshot[16].r.part1[24] );
tran (\sa_snapshot[16][56] , \sa_snapshot[16].f.unused[6] );
tran (\sa_snapshot[16][57] , \sa_snapshot[16].r.part1[25] );
tran (\sa_snapshot[16][57] , \sa_snapshot[16].f.unused[7] );
tran (\sa_snapshot[16][58] , \sa_snapshot[16].r.part1[26] );
tran (\sa_snapshot[16][58] , \sa_snapshot[16].f.unused[8] );
tran (\sa_snapshot[16][59] , \sa_snapshot[16].r.part1[27] );
tran (\sa_snapshot[16][59] , \sa_snapshot[16].f.unused[9] );
tran (\sa_snapshot[16][60] , \sa_snapshot[16].r.part1[28] );
tran (\sa_snapshot[16][60] , \sa_snapshot[16].f.unused[10] );
tran (\sa_snapshot[16][61] , \sa_snapshot[16].r.part1[29] );
tran (\sa_snapshot[16][61] , \sa_snapshot[16].f.unused[11] );
tran (\sa_snapshot[16][62] , \sa_snapshot[16].r.part1[30] );
tran (\sa_snapshot[16][62] , \sa_snapshot[16].f.unused[12] );
tran (\sa_snapshot[16][63] , \sa_snapshot[16].r.part1[31] );
tran (\sa_snapshot[16][63] , \sa_snapshot[16].f.unused[13] );
tran (\sa_snapshot[17][0] , \sa_snapshot[17].r.part0[0] );
tran (\sa_snapshot[17][0] , \sa_snapshot[17].f.lower[0] );
tran (\sa_snapshot[17][1] , \sa_snapshot[17].r.part0[1] );
tran (\sa_snapshot[17][1] , \sa_snapshot[17].f.lower[1] );
tran (\sa_snapshot[17][2] , \sa_snapshot[17].r.part0[2] );
tran (\sa_snapshot[17][2] , \sa_snapshot[17].f.lower[2] );
tran (\sa_snapshot[17][3] , \sa_snapshot[17].r.part0[3] );
tran (\sa_snapshot[17][3] , \sa_snapshot[17].f.lower[3] );
tran (\sa_snapshot[17][4] , \sa_snapshot[17].r.part0[4] );
tran (\sa_snapshot[17][4] , \sa_snapshot[17].f.lower[4] );
tran (\sa_snapshot[17][5] , \sa_snapshot[17].r.part0[5] );
tran (\sa_snapshot[17][5] , \sa_snapshot[17].f.lower[5] );
tran (\sa_snapshot[17][6] , \sa_snapshot[17].r.part0[6] );
tran (\sa_snapshot[17][6] , \sa_snapshot[17].f.lower[6] );
tran (\sa_snapshot[17][7] , \sa_snapshot[17].r.part0[7] );
tran (\sa_snapshot[17][7] , \sa_snapshot[17].f.lower[7] );
tran (\sa_snapshot[17][8] , \sa_snapshot[17].r.part0[8] );
tran (\sa_snapshot[17][8] , \sa_snapshot[17].f.lower[8] );
tran (\sa_snapshot[17][9] , \sa_snapshot[17].r.part0[9] );
tran (\sa_snapshot[17][9] , \sa_snapshot[17].f.lower[9] );
tran (\sa_snapshot[17][10] , \sa_snapshot[17].r.part0[10] );
tran (\sa_snapshot[17][10] , \sa_snapshot[17].f.lower[10] );
tran (\sa_snapshot[17][11] , \sa_snapshot[17].r.part0[11] );
tran (\sa_snapshot[17][11] , \sa_snapshot[17].f.lower[11] );
tran (\sa_snapshot[17][12] , \sa_snapshot[17].r.part0[12] );
tran (\sa_snapshot[17][12] , \sa_snapshot[17].f.lower[12] );
tran (\sa_snapshot[17][13] , \sa_snapshot[17].r.part0[13] );
tran (\sa_snapshot[17][13] , \sa_snapshot[17].f.lower[13] );
tran (\sa_snapshot[17][14] , \sa_snapshot[17].r.part0[14] );
tran (\sa_snapshot[17][14] , \sa_snapshot[17].f.lower[14] );
tran (\sa_snapshot[17][15] , \sa_snapshot[17].r.part0[15] );
tran (\sa_snapshot[17][15] , \sa_snapshot[17].f.lower[15] );
tran (\sa_snapshot[17][16] , \sa_snapshot[17].r.part0[16] );
tran (\sa_snapshot[17][16] , \sa_snapshot[17].f.lower[16] );
tran (\sa_snapshot[17][17] , \sa_snapshot[17].r.part0[17] );
tran (\sa_snapshot[17][17] , \sa_snapshot[17].f.lower[17] );
tran (\sa_snapshot[17][18] , \sa_snapshot[17].r.part0[18] );
tran (\sa_snapshot[17][18] , \sa_snapshot[17].f.lower[18] );
tran (\sa_snapshot[17][19] , \sa_snapshot[17].r.part0[19] );
tran (\sa_snapshot[17][19] , \sa_snapshot[17].f.lower[19] );
tran (\sa_snapshot[17][20] , \sa_snapshot[17].r.part0[20] );
tran (\sa_snapshot[17][20] , \sa_snapshot[17].f.lower[20] );
tran (\sa_snapshot[17][21] , \sa_snapshot[17].r.part0[21] );
tran (\sa_snapshot[17][21] , \sa_snapshot[17].f.lower[21] );
tran (\sa_snapshot[17][22] , \sa_snapshot[17].r.part0[22] );
tran (\sa_snapshot[17][22] , \sa_snapshot[17].f.lower[22] );
tran (\sa_snapshot[17][23] , \sa_snapshot[17].r.part0[23] );
tran (\sa_snapshot[17][23] , \sa_snapshot[17].f.lower[23] );
tran (\sa_snapshot[17][24] , \sa_snapshot[17].r.part0[24] );
tran (\sa_snapshot[17][24] , \sa_snapshot[17].f.lower[24] );
tran (\sa_snapshot[17][25] , \sa_snapshot[17].r.part0[25] );
tran (\sa_snapshot[17][25] , \sa_snapshot[17].f.lower[25] );
tran (\sa_snapshot[17][26] , \sa_snapshot[17].r.part0[26] );
tran (\sa_snapshot[17][26] , \sa_snapshot[17].f.lower[26] );
tran (\sa_snapshot[17][27] , \sa_snapshot[17].r.part0[27] );
tran (\sa_snapshot[17][27] , \sa_snapshot[17].f.lower[27] );
tran (\sa_snapshot[17][28] , \sa_snapshot[17].r.part0[28] );
tran (\sa_snapshot[17][28] , \sa_snapshot[17].f.lower[28] );
tran (\sa_snapshot[17][29] , \sa_snapshot[17].r.part0[29] );
tran (\sa_snapshot[17][29] , \sa_snapshot[17].f.lower[29] );
tran (\sa_snapshot[17][30] , \sa_snapshot[17].r.part0[30] );
tran (\sa_snapshot[17][30] , \sa_snapshot[17].f.lower[30] );
tran (\sa_snapshot[17][31] , \sa_snapshot[17].r.part0[31] );
tran (\sa_snapshot[17][31] , \sa_snapshot[17].f.lower[31] );
tran (\sa_snapshot[17][32] , \sa_snapshot[17].r.part1[0] );
tran (\sa_snapshot[17][32] , \sa_snapshot[17].f.upper[0] );
tran (\sa_snapshot[17][33] , \sa_snapshot[17].r.part1[1] );
tran (\sa_snapshot[17][33] , \sa_snapshot[17].f.upper[1] );
tran (\sa_snapshot[17][34] , \sa_snapshot[17].r.part1[2] );
tran (\sa_snapshot[17][34] , \sa_snapshot[17].f.upper[2] );
tran (\sa_snapshot[17][35] , \sa_snapshot[17].r.part1[3] );
tran (\sa_snapshot[17][35] , \sa_snapshot[17].f.upper[3] );
tran (\sa_snapshot[17][36] , \sa_snapshot[17].r.part1[4] );
tran (\sa_snapshot[17][36] , \sa_snapshot[17].f.upper[4] );
tran (\sa_snapshot[17][37] , \sa_snapshot[17].r.part1[5] );
tran (\sa_snapshot[17][37] , \sa_snapshot[17].f.upper[5] );
tran (\sa_snapshot[17][38] , \sa_snapshot[17].r.part1[6] );
tran (\sa_snapshot[17][38] , \sa_snapshot[17].f.upper[6] );
tran (\sa_snapshot[17][39] , \sa_snapshot[17].r.part1[7] );
tran (\sa_snapshot[17][39] , \sa_snapshot[17].f.upper[7] );
tran (\sa_snapshot[17][40] , \sa_snapshot[17].r.part1[8] );
tran (\sa_snapshot[17][40] , \sa_snapshot[17].f.upper[8] );
tran (\sa_snapshot[17][41] , \sa_snapshot[17].r.part1[9] );
tran (\sa_snapshot[17][41] , \sa_snapshot[17].f.upper[9] );
tran (\sa_snapshot[17][42] , \sa_snapshot[17].r.part1[10] );
tran (\sa_snapshot[17][42] , \sa_snapshot[17].f.upper[10] );
tran (\sa_snapshot[17][43] , \sa_snapshot[17].r.part1[11] );
tran (\sa_snapshot[17][43] , \sa_snapshot[17].f.upper[11] );
tran (\sa_snapshot[17][44] , \sa_snapshot[17].r.part1[12] );
tran (\sa_snapshot[17][44] , \sa_snapshot[17].f.upper[12] );
tran (\sa_snapshot[17][45] , \sa_snapshot[17].r.part1[13] );
tran (\sa_snapshot[17][45] , \sa_snapshot[17].f.upper[13] );
tran (\sa_snapshot[17][46] , \sa_snapshot[17].r.part1[14] );
tran (\sa_snapshot[17][46] , \sa_snapshot[17].f.upper[14] );
tran (\sa_snapshot[17][47] , \sa_snapshot[17].r.part1[15] );
tran (\sa_snapshot[17][47] , \sa_snapshot[17].f.upper[15] );
tran (\sa_snapshot[17][48] , \sa_snapshot[17].r.part1[16] );
tran (\sa_snapshot[17][48] , \sa_snapshot[17].f.upper[16] );
tran (\sa_snapshot[17][49] , \sa_snapshot[17].r.part1[17] );
tran (\sa_snapshot[17][49] , \sa_snapshot[17].f.upper[17] );
tran (\sa_snapshot[17][50] , \sa_snapshot[17].r.part1[18] );
tran (\sa_snapshot[17][50] , \sa_snapshot[17].f.unused[0] );
tran (\sa_snapshot[17][51] , \sa_snapshot[17].r.part1[19] );
tran (\sa_snapshot[17][51] , \sa_snapshot[17].f.unused[1] );
tran (\sa_snapshot[17][52] , \sa_snapshot[17].r.part1[20] );
tran (\sa_snapshot[17][52] , \sa_snapshot[17].f.unused[2] );
tran (\sa_snapshot[17][53] , \sa_snapshot[17].r.part1[21] );
tran (\sa_snapshot[17][53] , \sa_snapshot[17].f.unused[3] );
tran (\sa_snapshot[17][54] , \sa_snapshot[17].r.part1[22] );
tran (\sa_snapshot[17][54] , \sa_snapshot[17].f.unused[4] );
tran (\sa_snapshot[17][55] , \sa_snapshot[17].r.part1[23] );
tran (\sa_snapshot[17][55] , \sa_snapshot[17].f.unused[5] );
tran (\sa_snapshot[17][56] , \sa_snapshot[17].r.part1[24] );
tran (\sa_snapshot[17][56] , \sa_snapshot[17].f.unused[6] );
tran (\sa_snapshot[17][57] , \sa_snapshot[17].r.part1[25] );
tran (\sa_snapshot[17][57] , \sa_snapshot[17].f.unused[7] );
tran (\sa_snapshot[17][58] , \sa_snapshot[17].r.part1[26] );
tran (\sa_snapshot[17][58] , \sa_snapshot[17].f.unused[8] );
tran (\sa_snapshot[17][59] , \sa_snapshot[17].r.part1[27] );
tran (\sa_snapshot[17][59] , \sa_snapshot[17].f.unused[9] );
tran (\sa_snapshot[17][60] , \sa_snapshot[17].r.part1[28] );
tran (\sa_snapshot[17][60] , \sa_snapshot[17].f.unused[10] );
tran (\sa_snapshot[17][61] , \sa_snapshot[17].r.part1[29] );
tran (\sa_snapshot[17][61] , \sa_snapshot[17].f.unused[11] );
tran (\sa_snapshot[17][62] , \sa_snapshot[17].r.part1[30] );
tran (\sa_snapshot[17][62] , \sa_snapshot[17].f.unused[12] );
tran (\sa_snapshot[17][63] , \sa_snapshot[17].r.part1[31] );
tran (\sa_snapshot[17][63] , \sa_snapshot[17].f.unused[13] );
tran (\sa_snapshot[18][0] , \sa_snapshot[18].r.part0[0] );
tran (\sa_snapshot[18][0] , \sa_snapshot[18].f.lower[0] );
tran (\sa_snapshot[18][1] , \sa_snapshot[18].r.part0[1] );
tran (\sa_snapshot[18][1] , \sa_snapshot[18].f.lower[1] );
tran (\sa_snapshot[18][2] , \sa_snapshot[18].r.part0[2] );
tran (\sa_snapshot[18][2] , \sa_snapshot[18].f.lower[2] );
tran (\sa_snapshot[18][3] , \sa_snapshot[18].r.part0[3] );
tran (\sa_snapshot[18][3] , \sa_snapshot[18].f.lower[3] );
tran (\sa_snapshot[18][4] , \sa_snapshot[18].r.part0[4] );
tran (\sa_snapshot[18][4] , \sa_snapshot[18].f.lower[4] );
tran (\sa_snapshot[18][5] , \sa_snapshot[18].r.part0[5] );
tran (\sa_snapshot[18][5] , \sa_snapshot[18].f.lower[5] );
tran (\sa_snapshot[18][6] , \sa_snapshot[18].r.part0[6] );
tran (\sa_snapshot[18][6] , \sa_snapshot[18].f.lower[6] );
tran (\sa_snapshot[18][7] , \sa_snapshot[18].r.part0[7] );
tran (\sa_snapshot[18][7] , \sa_snapshot[18].f.lower[7] );
tran (\sa_snapshot[18][8] , \sa_snapshot[18].r.part0[8] );
tran (\sa_snapshot[18][8] , \sa_snapshot[18].f.lower[8] );
tran (\sa_snapshot[18][9] , \sa_snapshot[18].r.part0[9] );
tran (\sa_snapshot[18][9] , \sa_snapshot[18].f.lower[9] );
tran (\sa_snapshot[18][10] , \sa_snapshot[18].r.part0[10] );
tran (\sa_snapshot[18][10] , \sa_snapshot[18].f.lower[10] );
tran (\sa_snapshot[18][11] , \sa_snapshot[18].r.part0[11] );
tran (\sa_snapshot[18][11] , \sa_snapshot[18].f.lower[11] );
tran (\sa_snapshot[18][12] , \sa_snapshot[18].r.part0[12] );
tran (\sa_snapshot[18][12] , \sa_snapshot[18].f.lower[12] );
tran (\sa_snapshot[18][13] , \sa_snapshot[18].r.part0[13] );
tran (\sa_snapshot[18][13] , \sa_snapshot[18].f.lower[13] );
tran (\sa_snapshot[18][14] , \sa_snapshot[18].r.part0[14] );
tran (\sa_snapshot[18][14] , \sa_snapshot[18].f.lower[14] );
tran (\sa_snapshot[18][15] , \sa_snapshot[18].r.part0[15] );
tran (\sa_snapshot[18][15] , \sa_snapshot[18].f.lower[15] );
tran (\sa_snapshot[18][16] , \sa_snapshot[18].r.part0[16] );
tran (\sa_snapshot[18][16] , \sa_snapshot[18].f.lower[16] );
tran (\sa_snapshot[18][17] , \sa_snapshot[18].r.part0[17] );
tran (\sa_snapshot[18][17] , \sa_snapshot[18].f.lower[17] );
tran (\sa_snapshot[18][18] , \sa_snapshot[18].r.part0[18] );
tran (\sa_snapshot[18][18] , \sa_snapshot[18].f.lower[18] );
tran (\sa_snapshot[18][19] , \sa_snapshot[18].r.part0[19] );
tran (\sa_snapshot[18][19] , \sa_snapshot[18].f.lower[19] );
tran (\sa_snapshot[18][20] , \sa_snapshot[18].r.part0[20] );
tran (\sa_snapshot[18][20] , \sa_snapshot[18].f.lower[20] );
tran (\sa_snapshot[18][21] , \sa_snapshot[18].r.part0[21] );
tran (\sa_snapshot[18][21] , \sa_snapshot[18].f.lower[21] );
tran (\sa_snapshot[18][22] , \sa_snapshot[18].r.part0[22] );
tran (\sa_snapshot[18][22] , \sa_snapshot[18].f.lower[22] );
tran (\sa_snapshot[18][23] , \sa_snapshot[18].r.part0[23] );
tran (\sa_snapshot[18][23] , \sa_snapshot[18].f.lower[23] );
tran (\sa_snapshot[18][24] , \sa_snapshot[18].r.part0[24] );
tran (\sa_snapshot[18][24] , \sa_snapshot[18].f.lower[24] );
tran (\sa_snapshot[18][25] , \sa_snapshot[18].r.part0[25] );
tran (\sa_snapshot[18][25] , \sa_snapshot[18].f.lower[25] );
tran (\sa_snapshot[18][26] , \sa_snapshot[18].r.part0[26] );
tran (\sa_snapshot[18][26] , \sa_snapshot[18].f.lower[26] );
tran (\sa_snapshot[18][27] , \sa_snapshot[18].r.part0[27] );
tran (\sa_snapshot[18][27] , \sa_snapshot[18].f.lower[27] );
tran (\sa_snapshot[18][28] , \sa_snapshot[18].r.part0[28] );
tran (\sa_snapshot[18][28] , \sa_snapshot[18].f.lower[28] );
tran (\sa_snapshot[18][29] , \sa_snapshot[18].r.part0[29] );
tran (\sa_snapshot[18][29] , \sa_snapshot[18].f.lower[29] );
tran (\sa_snapshot[18][30] , \sa_snapshot[18].r.part0[30] );
tran (\sa_snapshot[18][30] , \sa_snapshot[18].f.lower[30] );
tran (\sa_snapshot[18][31] , \sa_snapshot[18].r.part0[31] );
tran (\sa_snapshot[18][31] , \sa_snapshot[18].f.lower[31] );
tran (\sa_snapshot[18][32] , \sa_snapshot[18].r.part1[0] );
tran (\sa_snapshot[18][32] , \sa_snapshot[18].f.upper[0] );
tran (\sa_snapshot[18][33] , \sa_snapshot[18].r.part1[1] );
tran (\sa_snapshot[18][33] , \sa_snapshot[18].f.upper[1] );
tran (\sa_snapshot[18][34] , \sa_snapshot[18].r.part1[2] );
tran (\sa_snapshot[18][34] , \sa_snapshot[18].f.upper[2] );
tran (\sa_snapshot[18][35] , \sa_snapshot[18].r.part1[3] );
tran (\sa_snapshot[18][35] , \sa_snapshot[18].f.upper[3] );
tran (\sa_snapshot[18][36] , \sa_snapshot[18].r.part1[4] );
tran (\sa_snapshot[18][36] , \sa_snapshot[18].f.upper[4] );
tran (\sa_snapshot[18][37] , \sa_snapshot[18].r.part1[5] );
tran (\sa_snapshot[18][37] , \sa_snapshot[18].f.upper[5] );
tran (\sa_snapshot[18][38] , \sa_snapshot[18].r.part1[6] );
tran (\sa_snapshot[18][38] , \sa_snapshot[18].f.upper[6] );
tran (\sa_snapshot[18][39] , \sa_snapshot[18].r.part1[7] );
tran (\sa_snapshot[18][39] , \sa_snapshot[18].f.upper[7] );
tran (\sa_snapshot[18][40] , \sa_snapshot[18].r.part1[8] );
tran (\sa_snapshot[18][40] , \sa_snapshot[18].f.upper[8] );
tran (\sa_snapshot[18][41] , \sa_snapshot[18].r.part1[9] );
tran (\sa_snapshot[18][41] , \sa_snapshot[18].f.upper[9] );
tran (\sa_snapshot[18][42] , \sa_snapshot[18].r.part1[10] );
tran (\sa_snapshot[18][42] , \sa_snapshot[18].f.upper[10] );
tran (\sa_snapshot[18][43] , \sa_snapshot[18].r.part1[11] );
tran (\sa_snapshot[18][43] , \sa_snapshot[18].f.upper[11] );
tran (\sa_snapshot[18][44] , \sa_snapshot[18].r.part1[12] );
tran (\sa_snapshot[18][44] , \sa_snapshot[18].f.upper[12] );
tran (\sa_snapshot[18][45] , \sa_snapshot[18].r.part1[13] );
tran (\sa_snapshot[18][45] , \sa_snapshot[18].f.upper[13] );
tran (\sa_snapshot[18][46] , \sa_snapshot[18].r.part1[14] );
tran (\sa_snapshot[18][46] , \sa_snapshot[18].f.upper[14] );
tran (\sa_snapshot[18][47] , \sa_snapshot[18].r.part1[15] );
tran (\sa_snapshot[18][47] , \sa_snapshot[18].f.upper[15] );
tran (\sa_snapshot[18][48] , \sa_snapshot[18].r.part1[16] );
tran (\sa_snapshot[18][48] , \sa_snapshot[18].f.upper[16] );
tran (\sa_snapshot[18][49] , \sa_snapshot[18].r.part1[17] );
tran (\sa_snapshot[18][49] , \sa_snapshot[18].f.upper[17] );
tran (\sa_snapshot[18][50] , \sa_snapshot[18].r.part1[18] );
tran (\sa_snapshot[18][50] , \sa_snapshot[18].f.unused[0] );
tran (\sa_snapshot[18][51] , \sa_snapshot[18].r.part1[19] );
tran (\sa_snapshot[18][51] , \sa_snapshot[18].f.unused[1] );
tran (\sa_snapshot[18][52] , \sa_snapshot[18].r.part1[20] );
tran (\sa_snapshot[18][52] , \sa_snapshot[18].f.unused[2] );
tran (\sa_snapshot[18][53] , \sa_snapshot[18].r.part1[21] );
tran (\sa_snapshot[18][53] , \sa_snapshot[18].f.unused[3] );
tran (\sa_snapshot[18][54] , \sa_snapshot[18].r.part1[22] );
tran (\sa_snapshot[18][54] , \sa_snapshot[18].f.unused[4] );
tran (\sa_snapshot[18][55] , \sa_snapshot[18].r.part1[23] );
tran (\sa_snapshot[18][55] , \sa_snapshot[18].f.unused[5] );
tran (\sa_snapshot[18][56] , \sa_snapshot[18].r.part1[24] );
tran (\sa_snapshot[18][56] , \sa_snapshot[18].f.unused[6] );
tran (\sa_snapshot[18][57] , \sa_snapshot[18].r.part1[25] );
tran (\sa_snapshot[18][57] , \sa_snapshot[18].f.unused[7] );
tran (\sa_snapshot[18][58] , \sa_snapshot[18].r.part1[26] );
tran (\sa_snapshot[18][58] , \sa_snapshot[18].f.unused[8] );
tran (\sa_snapshot[18][59] , \sa_snapshot[18].r.part1[27] );
tran (\sa_snapshot[18][59] , \sa_snapshot[18].f.unused[9] );
tran (\sa_snapshot[18][60] , \sa_snapshot[18].r.part1[28] );
tran (\sa_snapshot[18][60] , \sa_snapshot[18].f.unused[10] );
tran (\sa_snapshot[18][61] , \sa_snapshot[18].r.part1[29] );
tran (\sa_snapshot[18][61] , \sa_snapshot[18].f.unused[11] );
tran (\sa_snapshot[18][62] , \sa_snapshot[18].r.part1[30] );
tran (\sa_snapshot[18][62] , \sa_snapshot[18].f.unused[12] );
tran (\sa_snapshot[18][63] , \sa_snapshot[18].r.part1[31] );
tran (\sa_snapshot[18][63] , \sa_snapshot[18].f.unused[13] );
tran (\sa_snapshot[19][0] , \sa_snapshot[19].r.part0[0] );
tran (\sa_snapshot[19][0] , \sa_snapshot[19].f.lower[0] );
tran (\sa_snapshot[19][1] , \sa_snapshot[19].r.part0[1] );
tran (\sa_snapshot[19][1] , \sa_snapshot[19].f.lower[1] );
tran (\sa_snapshot[19][2] , \sa_snapshot[19].r.part0[2] );
tran (\sa_snapshot[19][2] , \sa_snapshot[19].f.lower[2] );
tran (\sa_snapshot[19][3] , \sa_snapshot[19].r.part0[3] );
tran (\sa_snapshot[19][3] , \sa_snapshot[19].f.lower[3] );
tran (\sa_snapshot[19][4] , \sa_snapshot[19].r.part0[4] );
tran (\sa_snapshot[19][4] , \sa_snapshot[19].f.lower[4] );
tran (\sa_snapshot[19][5] , \sa_snapshot[19].r.part0[5] );
tran (\sa_snapshot[19][5] , \sa_snapshot[19].f.lower[5] );
tran (\sa_snapshot[19][6] , \sa_snapshot[19].r.part0[6] );
tran (\sa_snapshot[19][6] , \sa_snapshot[19].f.lower[6] );
tran (\sa_snapshot[19][7] , \sa_snapshot[19].r.part0[7] );
tran (\sa_snapshot[19][7] , \sa_snapshot[19].f.lower[7] );
tran (\sa_snapshot[19][8] , \sa_snapshot[19].r.part0[8] );
tran (\sa_snapshot[19][8] , \sa_snapshot[19].f.lower[8] );
tran (\sa_snapshot[19][9] , \sa_snapshot[19].r.part0[9] );
tran (\sa_snapshot[19][9] , \sa_snapshot[19].f.lower[9] );
tran (\sa_snapshot[19][10] , \sa_snapshot[19].r.part0[10] );
tran (\sa_snapshot[19][10] , \sa_snapshot[19].f.lower[10] );
tran (\sa_snapshot[19][11] , \sa_snapshot[19].r.part0[11] );
tran (\sa_snapshot[19][11] , \sa_snapshot[19].f.lower[11] );
tran (\sa_snapshot[19][12] , \sa_snapshot[19].r.part0[12] );
tran (\sa_snapshot[19][12] , \sa_snapshot[19].f.lower[12] );
tran (\sa_snapshot[19][13] , \sa_snapshot[19].r.part0[13] );
tran (\sa_snapshot[19][13] , \sa_snapshot[19].f.lower[13] );
tran (\sa_snapshot[19][14] , \sa_snapshot[19].r.part0[14] );
tran (\sa_snapshot[19][14] , \sa_snapshot[19].f.lower[14] );
tran (\sa_snapshot[19][15] , \sa_snapshot[19].r.part0[15] );
tran (\sa_snapshot[19][15] , \sa_snapshot[19].f.lower[15] );
tran (\sa_snapshot[19][16] , \sa_snapshot[19].r.part0[16] );
tran (\sa_snapshot[19][16] , \sa_snapshot[19].f.lower[16] );
tran (\sa_snapshot[19][17] , \sa_snapshot[19].r.part0[17] );
tran (\sa_snapshot[19][17] , \sa_snapshot[19].f.lower[17] );
tran (\sa_snapshot[19][18] , \sa_snapshot[19].r.part0[18] );
tran (\sa_snapshot[19][18] , \sa_snapshot[19].f.lower[18] );
tran (\sa_snapshot[19][19] , \sa_snapshot[19].r.part0[19] );
tran (\sa_snapshot[19][19] , \sa_snapshot[19].f.lower[19] );
tran (\sa_snapshot[19][20] , \sa_snapshot[19].r.part0[20] );
tran (\sa_snapshot[19][20] , \sa_snapshot[19].f.lower[20] );
tran (\sa_snapshot[19][21] , \sa_snapshot[19].r.part0[21] );
tran (\sa_snapshot[19][21] , \sa_snapshot[19].f.lower[21] );
tran (\sa_snapshot[19][22] , \sa_snapshot[19].r.part0[22] );
tran (\sa_snapshot[19][22] , \sa_snapshot[19].f.lower[22] );
tran (\sa_snapshot[19][23] , \sa_snapshot[19].r.part0[23] );
tran (\sa_snapshot[19][23] , \sa_snapshot[19].f.lower[23] );
tran (\sa_snapshot[19][24] , \sa_snapshot[19].r.part0[24] );
tran (\sa_snapshot[19][24] , \sa_snapshot[19].f.lower[24] );
tran (\sa_snapshot[19][25] , \sa_snapshot[19].r.part0[25] );
tran (\sa_snapshot[19][25] , \sa_snapshot[19].f.lower[25] );
tran (\sa_snapshot[19][26] , \sa_snapshot[19].r.part0[26] );
tran (\sa_snapshot[19][26] , \sa_snapshot[19].f.lower[26] );
tran (\sa_snapshot[19][27] , \sa_snapshot[19].r.part0[27] );
tran (\sa_snapshot[19][27] , \sa_snapshot[19].f.lower[27] );
tran (\sa_snapshot[19][28] , \sa_snapshot[19].r.part0[28] );
tran (\sa_snapshot[19][28] , \sa_snapshot[19].f.lower[28] );
tran (\sa_snapshot[19][29] , \sa_snapshot[19].r.part0[29] );
tran (\sa_snapshot[19][29] , \sa_snapshot[19].f.lower[29] );
tran (\sa_snapshot[19][30] , \sa_snapshot[19].r.part0[30] );
tran (\sa_snapshot[19][30] , \sa_snapshot[19].f.lower[30] );
tran (\sa_snapshot[19][31] , \sa_snapshot[19].r.part0[31] );
tran (\sa_snapshot[19][31] , \sa_snapshot[19].f.lower[31] );
tran (\sa_snapshot[19][32] , \sa_snapshot[19].r.part1[0] );
tran (\sa_snapshot[19][32] , \sa_snapshot[19].f.upper[0] );
tran (\sa_snapshot[19][33] , \sa_snapshot[19].r.part1[1] );
tran (\sa_snapshot[19][33] , \sa_snapshot[19].f.upper[1] );
tran (\sa_snapshot[19][34] , \sa_snapshot[19].r.part1[2] );
tran (\sa_snapshot[19][34] , \sa_snapshot[19].f.upper[2] );
tran (\sa_snapshot[19][35] , \sa_snapshot[19].r.part1[3] );
tran (\sa_snapshot[19][35] , \sa_snapshot[19].f.upper[3] );
tran (\sa_snapshot[19][36] , \sa_snapshot[19].r.part1[4] );
tran (\sa_snapshot[19][36] , \sa_snapshot[19].f.upper[4] );
tran (\sa_snapshot[19][37] , \sa_snapshot[19].r.part1[5] );
tran (\sa_snapshot[19][37] , \sa_snapshot[19].f.upper[5] );
tran (\sa_snapshot[19][38] , \sa_snapshot[19].r.part1[6] );
tran (\sa_snapshot[19][38] , \sa_snapshot[19].f.upper[6] );
tran (\sa_snapshot[19][39] , \sa_snapshot[19].r.part1[7] );
tran (\sa_snapshot[19][39] , \sa_snapshot[19].f.upper[7] );
tran (\sa_snapshot[19][40] , \sa_snapshot[19].r.part1[8] );
tran (\sa_snapshot[19][40] , \sa_snapshot[19].f.upper[8] );
tran (\sa_snapshot[19][41] , \sa_snapshot[19].r.part1[9] );
tran (\sa_snapshot[19][41] , \sa_snapshot[19].f.upper[9] );
tran (\sa_snapshot[19][42] , \sa_snapshot[19].r.part1[10] );
tran (\sa_snapshot[19][42] , \sa_snapshot[19].f.upper[10] );
tran (\sa_snapshot[19][43] , \sa_snapshot[19].r.part1[11] );
tran (\sa_snapshot[19][43] , \sa_snapshot[19].f.upper[11] );
tran (\sa_snapshot[19][44] , \sa_snapshot[19].r.part1[12] );
tran (\sa_snapshot[19][44] , \sa_snapshot[19].f.upper[12] );
tran (\sa_snapshot[19][45] , \sa_snapshot[19].r.part1[13] );
tran (\sa_snapshot[19][45] , \sa_snapshot[19].f.upper[13] );
tran (\sa_snapshot[19][46] , \sa_snapshot[19].r.part1[14] );
tran (\sa_snapshot[19][46] , \sa_snapshot[19].f.upper[14] );
tran (\sa_snapshot[19][47] , \sa_snapshot[19].r.part1[15] );
tran (\sa_snapshot[19][47] , \sa_snapshot[19].f.upper[15] );
tran (\sa_snapshot[19][48] , \sa_snapshot[19].r.part1[16] );
tran (\sa_snapshot[19][48] , \sa_snapshot[19].f.upper[16] );
tran (\sa_snapshot[19][49] , \sa_snapshot[19].r.part1[17] );
tran (\sa_snapshot[19][49] , \sa_snapshot[19].f.upper[17] );
tran (\sa_snapshot[19][50] , \sa_snapshot[19].r.part1[18] );
tran (\sa_snapshot[19][50] , \sa_snapshot[19].f.unused[0] );
tran (\sa_snapshot[19][51] , \sa_snapshot[19].r.part1[19] );
tran (\sa_snapshot[19][51] , \sa_snapshot[19].f.unused[1] );
tran (\sa_snapshot[19][52] , \sa_snapshot[19].r.part1[20] );
tran (\sa_snapshot[19][52] , \sa_snapshot[19].f.unused[2] );
tran (\sa_snapshot[19][53] , \sa_snapshot[19].r.part1[21] );
tran (\sa_snapshot[19][53] , \sa_snapshot[19].f.unused[3] );
tran (\sa_snapshot[19][54] , \sa_snapshot[19].r.part1[22] );
tran (\sa_snapshot[19][54] , \sa_snapshot[19].f.unused[4] );
tran (\sa_snapshot[19][55] , \sa_snapshot[19].r.part1[23] );
tran (\sa_snapshot[19][55] , \sa_snapshot[19].f.unused[5] );
tran (\sa_snapshot[19][56] , \sa_snapshot[19].r.part1[24] );
tran (\sa_snapshot[19][56] , \sa_snapshot[19].f.unused[6] );
tran (\sa_snapshot[19][57] , \sa_snapshot[19].r.part1[25] );
tran (\sa_snapshot[19][57] , \sa_snapshot[19].f.unused[7] );
tran (\sa_snapshot[19][58] , \sa_snapshot[19].r.part1[26] );
tran (\sa_snapshot[19][58] , \sa_snapshot[19].f.unused[8] );
tran (\sa_snapshot[19][59] , \sa_snapshot[19].r.part1[27] );
tran (\sa_snapshot[19][59] , \sa_snapshot[19].f.unused[9] );
tran (\sa_snapshot[19][60] , \sa_snapshot[19].r.part1[28] );
tran (\sa_snapshot[19][60] , \sa_snapshot[19].f.unused[10] );
tran (\sa_snapshot[19][61] , \sa_snapshot[19].r.part1[29] );
tran (\sa_snapshot[19][61] , \sa_snapshot[19].f.unused[11] );
tran (\sa_snapshot[19][62] , \sa_snapshot[19].r.part1[30] );
tran (\sa_snapshot[19][62] , \sa_snapshot[19].f.unused[12] );
tran (\sa_snapshot[19][63] , \sa_snapshot[19].r.part1[31] );
tran (\sa_snapshot[19][63] , \sa_snapshot[19].f.unused[13] );
tran (\sa_snapshot[20][0] , \sa_snapshot[20].r.part0[0] );
tran (\sa_snapshot[20][0] , \sa_snapshot[20].f.lower[0] );
tran (\sa_snapshot[20][1] , \sa_snapshot[20].r.part0[1] );
tran (\sa_snapshot[20][1] , \sa_snapshot[20].f.lower[1] );
tran (\sa_snapshot[20][2] , \sa_snapshot[20].r.part0[2] );
tran (\sa_snapshot[20][2] , \sa_snapshot[20].f.lower[2] );
tran (\sa_snapshot[20][3] , \sa_snapshot[20].r.part0[3] );
tran (\sa_snapshot[20][3] , \sa_snapshot[20].f.lower[3] );
tran (\sa_snapshot[20][4] , \sa_snapshot[20].r.part0[4] );
tran (\sa_snapshot[20][4] , \sa_snapshot[20].f.lower[4] );
tran (\sa_snapshot[20][5] , \sa_snapshot[20].r.part0[5] );
tran (\sa_snapshot[20][5] , \sa_snapshot[20].f.lower[5] );
tran (\sa_snapshot[20][6] , \sa_snapshot[20].r.part0[6] );
tran (\sa_snapshot[20][6] , \sa_snapshot[20].f.lower[6] );
tran (\sa_snapshot[20][7] , \sa_snapshot[20].r.part0[7] );
tran (\sa_snapshot[20][7] , \sa_snapshot[20].f.lower[7] );
tran (\sa_snapshot[20][8] , \sa_snapshot[20].r.part0[8] );
tran (\sa_snapshot[20][8] , \sa_snapshot[20].f.lower[8] );
tran (\sa_snapshot[20][9] , \sa_snapshot[20].r.part0[9] );
tran (\sa_snapshot[20][9] , \sa_snapshot[20].f.lower[9] );
tran (\sa_snapshot[20][10] , \sa_snapshot[20].r.part0[10] );
tran (\sa_snapshot[20][10] , \sa_snapshot[20].f.lower[10] );
tran (\sa_snapshot[20][11] , \sa_snapshot[20].r.part0[11] );
tran (\sa_snapshot[20][11] , \sa_snapshot[20].f.lower[11] );
tran (\sa_snapshot[20][12] , \sa_snapshot[20].r.part0[12] );
tran (\sa_snapshot[20][12] , \sa_snapshot[20].f.lower[12] );
tran (\sa_snapshot[20][13] , \sa_snapshot[20].r.part0[13] );
tran (\sa_snapshot[20][13] , \sa_snapshot[20].f.lower[13] );
tran (\sa_snapshot[20][14] , \sa_snapshot[20].r.part0[14] );
tran (\sa_snapshot[20][14] , \sa_snapshot[20].f.lower[14] );
tran (\sa_snapshot[20][15] , \sa_snapshot[20].r.part0[15] );
tran (\sa_snapshot[20][15] , \sa_snapshot[20].f.lower[15] );
tran (\sa_snapshot[20][16] , \sa_snapshot[20].r.part0[16] );
tran (\sa_snapshot[20][16] , \sa_snapshot[20].f.lower[16] );
tran (\sa_snapshot[20][17] , \sa_snapshot[20].r.part0[17] );
tran (\sa_snapshot[20][17] , \sa_snapshot[20].f.lower[17] );
tran (\sa_snapshot[20][18] , \sa_snapshot[20].r.part0[18] );
tran (\sa_snapshot[20][18] , \sa_snapshot[20].f.lower[18] );
tran (\sa_snapshot[20][19] , \sa_snapshot[20].r.part0[19] );
tran (\sa_snapshot[20][19] , \sa_snapshot[20].f.lower[19] );
tran (\sa_snapshot[20][20] , \sa_snapshot[20].r.part0[20] );
tran (\sa_snapshot[20][20] , \sa_snapshot[20].f.lower[20] );
tran (\sa_snapshot[20][21] , \sa_snapshot[20].r.part0[21] );
tran (\sa_snapshot[20][21] , \sa_snapshot[20].f.lower[21] );
tran (\sa_snapshot[20][22] , \sa_snapshot[20].r.part0[22] );
tran (\sa_snapshot[20][22] , \sa_snapshot[20].f.lower[22] );
tran (\sa_snapshot[20][23] , \sa_snapshot[20].r.part0[23] );
tran (\sa_snapshot[20][23] , \sa_snapshot[20].f.lower[23] );
tran (\sa_snapshot[20][24] , \sa_snapshot[20].r.part0[24] );
tran (\sa_snapshot[20][24] , \sa_snapshot[20].f.lower[24] );
tran (\sa_snapshot[20][25] , \sa_snapshot[20].r.part0[25] );
tran (\sa_snapshot[20][25] , \sa_snapshot[20].f.lower[25] );
tran (\sa_snapshot[20][26] , \sa_snapshot[20].r.part0[26] );
tran (\sa_snapshot[20][26] , \sa_snapshot[20].f.lower[26] );
tran (\sa_snapshot[20][27] , \sa_snapshot[20].r.part0[27] );
tran (\sa_snapshot[20][27] , \sa_snapshot[20].f.lower[27] );
tran (\sa_snapshot[20][28] , \sa_snapshot[20].r.part0[28] );
tran (\sa_snapshot[20][28] , \sa_snapshot[20].f.lower[28] );
tran (\sa_snapshot[20][29] , \sa_snapshot[20].r.part0[29] );
tran (\sa_snapshot[20][29] , \sa_snapshot[20].f.lower[29] );
tran (\sa_snapshot[20][30] , \sa_snapshot[20].r.part0[30] );
tran (\sa_snapshot[20][30] , \sa_snapshot[20].f.lower[30] );
tran (\sa_snapshot[20][31] , \sa_snapshot[20].r.part0[31] );
tran (\sa_snapshot[20][31] , \sa_snapshot[20].f.lower[31] );
tran (\sa_snapshot[20][32] , \sa_snapshot[20].r.part1[0] );
tran (\sa_snapshot[20][32] , \sa_snapshot[20].f.upper[0] );
tran (\sa_snapshot[20][33] , \sa_snapshot[20].r.part1[1] );
tran (\sa_snapshot[20][33] , \sa_snapshot[20].f.upper[1] );
tran (\sa_snapshot[20][34] , \sa_snapshot[20].r.part1[2] );
tran (\sa_snapshot[20][34] , \sa_snapshot[20].f.upper[2] );
tran (\sa_snapshot[20][35] , \sa_snapshot[20].r.part1[3] );
tran (\sa_snapshot[20][35] , \sa_snapshot[20].f.upper[3] );
tran (\sa_snapshot[20][36] , \sa_snapshot[20].r.part1[4] );
tran (\sa_snapshot[20][36] , \sa_snapshot[20].f.upper[4] );
tran (\sa_snapshot[20][37] , \sa_snapshot[20].r.part1[5] );
tran (\sa_snapshot[20][37] , \sa_snapshot[20].f.upper[5] );
tran (\sa_snapshot[20][38] , \sa_snapshot[20].r.part1[6] );
tran (\sa_snapshot[20][38] , \sa_snapshot[20].f.upper[6] );
tran (\sa_snapshot[20][39] , \sa_snapshot[20].r.part1[7] );
tran (\sa_snapshot[20][39] , \sa_snapshot[20].f.upper[7] );
tran (\sa_snapshot[20][40] , \sa_snapshot[20].r.part1[8] );
tran (\sa_snapshot[20][40] , \sa_snapshot[20].f.upper[8] );
tran (\sa_snapshot[20][41] , \sa_snapshot[20].r.part1[9] );
tran (\sa_snapshot[20][41] , \sa_snapshot[20].f.upper[9] );
tran (\sa_snapshot[20][42] , \sa_snapshot[20].r.part1[10] );
tran (\sa_snapshot[20][42] , \sa_snapshot[20].f.upper[10] );
tran (\sa_snapshot[20][43] , \sa_snapshot[20].r.part1[11] );
tran (\sa_snapshot[20][43] , \sa_snapshot[20].f.upper[11] );
tran (\sa_snapshot[20][44] , \sa_snapshot[20].r.part1[12] );
tran (\sa_snapshot[20][44] , \sa_snapshot[20].f.upper[12] );
tran (\sa_snapshot[20][45] , \sa_snapshot[20].r.part1[13] );
tran (\sa_snapshot[20][45] , \sa_snapshot[20].f.upper[13] );
tran (\sa_snapshot[20][46] , \sa_snapshot[20].r.part1[14] );
tran (\sa_snapshot[20][46] , \sa_snapshot[20].f.upper[14] );
tran (\sa_snapshot[20][47] , \sa_snapshot[20].r.part1[15] );
tran (\sa_snapshot[20][47] , \sa_snapshot[20].f.upper[15] );
tran (\sa_snapshot[20][48] , \sa_snapshot[20].r.part1[16] );
tran (\sa_snapshot[20][48] , \sa_snapshot[20].f.upper[16] );
tran (\sa_snapshot[20][49] , \sa_snapshot[20].r.part1[17] );
tran (\sa_snapshot[20][49] , \sa_snapshot[20].f.upper[17] );
tran (\sa_snapshot[20][50] , \sa_snapshot[20].r.part1[18] );
tran (\sa_snapshot[20][50] , \sa_snapshot[20].f.unused[0] );
tran (\sa_snapshot[20][51] , \sa_snapshot[20].r.part1[19] );
tran (\sa_snapshot[20][51] , \sa_snapshot[20].f.unused[1] );
tran (\sa_snapshot[20][52] , \sa_snapshot[20].r.part1[20] );
tran (\sa_snapshot[20][52] , \sa_snapshot[20].f.unused[2] );
tran (\sa_snapshot[20][53] , \sa_snapshot[20].r.part1[21] );
tran (\sa_snapshot[20][53] , \sa_snapshot[20].f.unused[3] );
tran (\sa_snapshot[20][54] , \sa_snapshot[20].r.part1[22] );
tran (\sa_snapshot[20][54] , \sa_snapshot[20].f.unused[4] );
tran (\sa_snapshot[20][55] , \sa_snapshot[20].r.part1[23] );
tran (\sa_snapshot[20][55] , \sa_snapshot[20].f.unused[5] );
tran (\sa_snapshot[20][56] , \sa_snapshot[20].r.part1[24] );
tran (\sa_snapshot[20][56] , \sa_snapshot[20].f.unused[6] );
tran (\sa_snapshot[20][57] , \sa_snapshot[20].r.part1[25] );
tran (\sa_snapshot[20][57] , \sa_snapshot[20].f.unused[7] );
tran (\sa_snapshot[20][58] , \sa_snapshot[20].r.part1[26] );
tran (\sa_snapshot[20][58] , \sa_snapshot[20].f.unused[8] );
tran (\sa_snapshot[20][59] , \sa_snapshot[20].r.part1[27] );
tran (\sa_snapshot[20][59] , \sa_snapshot[20].f.unused[9] );
tran (\sa_snapshot[20][60] , \sa_snapshot[20].r.part1[28] );
tran (\sa_snapshot[20][60] , \sa_snapshot[20].f.unused[10] );
tran (\sa_snapshot[20][61] , \sa_snapshot[20].r.part1[29] );
tran (\sa_snapshot[20][61] , \sa_snapshot[20].f.unused[11] );
tran (\sa_snapshot[20][62] , \sa_snapshot[20].r.part1[30] );
tran (\sa_snapshot[20][62] , \sa_snapshot[20].f.unused[12] );
tran (\sa_snapshot[20][63] , \sa_snapshot[20].r.part1[31] );
tran (\sa_snapshot[20][63] , \sa_snapshot[20].f.unused[13] );
tran (\sa_snapshot[21][0] , \sa_snapshot[21].r.part0[0] );
tran (\sa_snapshot[21][0] , \sa_snapshot[21].f.lower[0] );
tran (\sa_snapshot[21][1] , \sa_snapshot[21].r.part0[1] );
tran (\sa_snapshot[21][1] , \sa_snapshot[21].f.lower[1] );
tran (\sa_snapshot[21][2] , \sa_snapshot[21].r.part0[2] );
tran (\sa_snapshot[21][2] , \sa_snapshot[21].f.lower[2] );
tran (\sa_snapshot[21][3] , \sa_snapshot[21].r.part0[3] );
tran (\sa_snapshot[21][3] , \sa_snapshot[21].f.lower[3] );
tran (\sa_snapshot[21][4] , \sa_snapshot[21].r.part0[4] );
tran (\sa_snapshot[21][4] , \sa_snapshot[21].f.lower[4] );
tran (\sa_snapshot[21][5] , \sa_snapshot[21].r.part0[5] );
tran (\sa_snapshot[21][5] , \sa_snapshot[21].f.lower[5] );
tran (\sa_snapshot[21][6] , \sa_snapshot[21].r.part0[6] );
tran (\sa_snapshot[21][6] , \sa_snapshot[21].f.lower[6] );
tran (\sa_snapshot[21][7] , \sa_snapshot[21].r.part0[7] );
tran (\sa_snapshot[21][7] , \sa_snapshot[21].f.lower[7] );
tran (\sa_snapshot[21][8] , \sa_snapshot[21].r.part0[8] );
tran (\sa_snapshot[21][8] , \sa_snapshot[21].f.lower[8] );
tran (\sa_snapshot[21][9] , \sa_snapshot[21].r.part0[9] );
tran (\sa_snapshot[21][9] , \sa_snapshot[21].f.lower[9] );
tran (\sa_snapshot[21][10] , \sa_snapshot[21].r.part0[10] );
tran (\sa_snapshot[21][10] , \sa_snapshot[21].f.lower[10] );
tran (\sa_snapshot[21][11] , \sa_snapshot[21].r.part0[11] );
tran (\sa_snapshot[21][11] , \sa_snapshot[21].f.lower[11] );
tran (\sa_snapshot[21][12] , \sa_snapshot[21].r.part0[12] );
tran (\sa_snapshot[21][12] , \sa_snapshot[21].f.lower[12] );
tran (\sa_snapshot[21][13] , \sa_snapshot[21].r.part0[13] );
tran (\sa_snapshot[21][13] , \sa_snapshot[21].f.lower[13] );
tran (\sa_snapshot[21][14] , \sa_snapshot[21].r.part0[14] );
tran (\sa_snapshot[21][14] , \sa_snapshot[21].f.lower[14] );
tran (\sa_snapshot[21][15] , \sa_snapshot[21].r.part0[15] );
tran (\sa_snapshot[21][15] , \sa_snapshot[21].f.lower[15] );
tran (\sa_snapshot[21][16] , \sa_snapshot[21].r.part0[16] );
tran (\sa_snapshot[21][16] , \sa_snapshot[21].f.lower[16] );
tran (\sa_snapshot[21][17] , \sa_snapshot[21].r.part0[17] );
tran (\sa_snapshot[21][17] , \sa_snapshot[21].f.lower[17] );
tran (\sa_snapshot[21][18] , \sa_snapshot[21].r.part0[18] );
tran (\sa_snapshot[21][18] , \sa_snapshot[21].f.lower[18] );
tran (\sa_snapshot[21][19] , \sa_snapshot[21].r.part0[19] );
tran (\sa_snapshot[21][19] , \sa_snapshot[21].f.lower[19] );
tran (\sa_snapshot[21][20] , \sa_snapshot[21].r.part0[20] );
tran (\sa_snapshot[21][20] , \sa_snapshot[21].f.lower[20] );
tran (\sa_snapshot[21][21] , \sa_snapshot[21].r.part0[21] );
tran (\sa_snapshot[21][21] , \sa_snapshot[21].f.lower[21] );
tran (\sa_snapshot[21][22] , \sa_snapshot[21].r.part0[22] );
tran (\sa_snapshot[21][22] , \sa_snapshot[21].f.lower[22] );
tran (\sa_snapshot[21][23] , \sa_snapshot[21].r.part0[23] );
tran (\sa_snapshot[21][23] , \sa_snapshot[21].f.lower[23] );
tran (\sa_snapshot[21][24] , \sa_snapshot[21].r.part0[24] );
tran (\sa_snapshot[21][24] , \sa_snapshot[21].f.lower[24] );
tran (\sa_snapshot[21][25] , \sa_snapshot[21].r.part0[25] );
tran (\sa_snapshot[21][25] , \sa_snapshot[21].f.lower[25] );
tran (\sa_snapshot[21][26] , \sa_snapshot[21].r.part0[26] );
tran (\sa_snapshot[21][26] , \sa_snapshot[21].f.lower[26] );
tran (\sa_snapshot[21][27] , \sa_snapshot[21].r.part0[27] );
tran (\sa_snapshot[21][27] , \sa_snapshot[21].f.lower[27] );
tran (\sa_snapshot[21][28] , \sa_snapshot[21].r.part0[28] );
tran (\sa_snapshot[21][28] , \sa_snapshot[21].f.lower[28] );
tran (\sa_snapshot[21][29] , \sa_snapshot[21].r.part0[29] );
tran (\sa_snapshot[21][29] , \sa_snapshot[21].f.lower[29] );
tran (\sa_snapshot[21][30] , \sa_snapshot[21].r.part0[30] );
tran (\sa_snapshot[21][30] , \sa_snapshot[21].f.lower[30] );
tran (\sa_snapshot[21][31] , \sa_snapshot[21].r.part0[31] );
tran (\sa_snapshot[21][31] , \sa_snapshot[21].f.lower[31] );
tran (\sa_snapshot[21][32] , \sa_snapshot[21].r.part1[0] );
tran (\sa_snapshot[21][32] , \sa_snapshot[21].f.upper[0] );
tran (\sa_snapshot[21][33] , \sa_snapshot[21].r.part1[1] );
tran (\sa_snapshot[21][33] , \sa_snapshot[21].f.upper[1] );
tran (\sa_snapshot[21][34] , \sa_snapshot[21].r.part1[2] );
tran (\sa_snapshot[21][34] , \sa_snapshot[21].f.upper[2] );
tran (\sa_snapshot[21][35] , \sa_snapshot[21].r.part1[3] );
tran (\sa_snapshot[21][35] , \sa_snapshot[21].f.upper[3] );
tran (\sa_snapshot[21][36] , \sa_snapshot[21].r.part1[4] );
tran (\sa_snapshot[21][36] , \sa_snapshot[21].f.upper[4] );
tran (\sa_snapshot[21][37] , \sa_snapshot[21].r.part1[5] );
tran (\sa_snapshot[21][37] , \sa_snapshot[21].f.upper[5] );
tran (\sa_snapshot[21][38] , \sa_snapshot[21].r.part1[6] );
tran (\sa_snapshot[21][38] , \sa_snapshot[21].f.upper[6] );
tran (\sa_snapshot[21][39] , \sa_snapshot[21].r.part1[7] );
tran (\sa_snapshot[21][39] , \sa_snapshot[21].f.upper[7] );
tran (\sa_snapshot[21][40] , \sa_snapshot[21].r.part1[8] );
tran (\sa_snapshot[21][40] , \sa_snapshot[21].f.upper[8] );
tran (\sa_snapshot[21][41] , \sa_snapshot[21].r.part1[9] );
tran (\sa_snapshot[21][41] , \sa_snapshot[21].f.upper[9] );
tran (\sa_snapshot[21][42] , \sa_snapshot[21].r.part1[10] );
tran (\sa_snapshot[21][42] , \sa_snapshot[21].f.upper[10] );
tran (\sa_snapshot[21][43] , \sa_snapshot[21].r.part1[11] );
tran (\sa_snapshot[21][43] , \sa_snapshot[21].f.upper[11] );
tran (\sa_snapshot[21][44] , \sa_snapshot[21].r.part1[12] );
tran (\sa_snapshot[21][44] , \sa_snapshot[21].f.upper[12] );
tran (\sa_snapshot[21][45] , \sa_snapshot[21].r.part1[13] );
tran (\sa_snapshot[21][45] , \sa_snapshot[21].f.upper[13] );
tran (\sa_snapshot[21][46] , \sa_snapshot[21].r.part1[14] );
tran (\sa_snapshot[21][46] , \sa_snapshot[21].f.upper[14] );
tran (\sa_snapshot[21][47] , \sa_snapshot[21].r.part1[15] );
tran (\sa_snapshot[21][47] , \sa_snapshot[21].f.upper[15] );
tran (\sa_snapshot[21][48] , \sa_snapshot[21].r.part1[16] );
tran (\sa_snapshot[21][48] , \sa_snapshot[21].f.upper[16] );
tran (\sa_snapshot[21][49] , \sa_snapshot[21].r.part1[17] );
tran (\sa_snapshot[21][49] , \sa_snapshot[21].f.upper[17] );
tran (\sa_snapshot[21][50] , \sa_snapshot[21].r.part1[18] );
tran (\sa_snapshot[21][50] , \sa_snapshot[21].f.unused[0] );
tran (\sa_snapshot[21][51] , \sa_snapshot[21].r.part1[19] );
tran (\sa_snapshot[21][51] , \sa_snapshot[21].f.unused[1] );
tran (\sa_snapshot[21][52] , \sa_snapshot[21].r.part1[20] );
tran (\sa_snapshot[21][52] , \sa_snapshot[21].f.unused[2] );
tran (\sa_snapshot[21][53] , \sa_snapshot[21].r.part1[21] );
tran (\sa_snapshot[21][53] , \sa_snapshot[21].f.unused[3] );
tran (\sa_snapshot[21][54] , \sa_snapshot[21].r.part1[22] );
tran (\sa_snapshot[21][54] , \sa_snapshot[21].f.unused[4] );
tran (\sa_snapshot[21][55] , \sa_snapshot[21].r.part1[23] );
tran (\sa_snapshot[21][55] , \sa_snapshot[21].f.unused[5] );
tran (\sa_snapshot[21][56] , \sa_snapshot[21].r.part1[24] );
tran (\sa_snapshot[21][56] , \sa_snapshot[21].f.unused[6] );
tran (\sa_snapshot[21][57] , \sa_snapshot[21].r.part1[25] );
tran (\sa_snapshot[21][57] , \sa_snapshot[21].f.unused[7] );
tran (\sa_snapshot[21][58] , \sa_snapshot[21].r.part1[26] );
tran (\sa_snapshot[21][58] , \sa_snapshot[21].f.unused[8] );
tran (\sa_snapshot[21][59] , \sa_snapshot[21].r.part1[27] );
tran (\sa_snapshot[21][59] , \sa_snapshot[21].f.unused[9] );
tran (\sa_snapshot[21][60] , \sa_snapshot[21].r.part1[28] );
tran (\sa_snapshot[21][60] , \sa_snapshot[21].f.unused[10] );
tran (\sa_snapshot[21][61] , \sa_snapshot[21].r.part1[29] );
tran (\sa_snapshot[21][61] , \sa_snapshot[21].f.unused[11] );
tran (\sa_snapshot[21][62] , \sa_snapshot[21].r.part1[30] );
tran (\sa_snapshot[21][62] , \sa_snapshot[21].f.unused[12] );
tran (\sa_snapshot[21][63] , \sa_snapshot[21].r.part1[31] );
tran (\sa_snapshot[21][63] , \sa_snapshot[21].f.unused[13] );
tran (\sa_snapshot[22][0] , \sa_snapshot[22].r.part0[0] );
tran (\sa_snapshot[22][0] , \sa_snapshot[22].f.lower[0] );
tran (\sa_snapshot[22][1] , \sa_snapshot[22].r.part0[1] );
tran (\sa_snapshot[22][1] , \sa_snapshot[22].f.lower[1] );
tran (\sa_snapshot[22][2] , \sa_snapshot[22].r.part0[2] );
tran (\sa_snapshot[22][2] , \sa_snapshot[22].f.lower[2] );
tran (\sa_snapshot[22][3] , \sa_snapshot[22].r.part0[3] );
tran (\sa_snapshot[22][3] , \sa_snapshot[22].f.lower[3] );
tran (\sa_snapshot[22][4] , \sa_snapshot[22].r.part0[4] );
tran (\sa_snapshot[22][4] , \sa_snapshot[22].f.lower[4] );
tran (\sa_snapshot[22][5] , \sa_snapshot[22].r.part0[5] );
tran (\sa_snapshot[22][5] , \sa_snapshot[22].f.lower[5] );
tran (\sa_snapshot[22][6] , \sa_snapshot[22].r.part0[6] );
tran (\sa_snapshot[22][6] , \sa_snapshot[22].f.lower[6] );
tran (\sa_snapshot[22][7] , \sa_snapshot[22].r.part0[7] );
tran (\sa_snapshot[22][7] , \sa_snapshot[22].f.lower[7] );
tran (\sa_snapshot[22][8] , \sa_snapshot[22].r.part0[8] );
tran (\sa_snapshot[22][8] , \sa_snapshot[22].f.lower[8] );
tran (\sa_snapshot[22][9] , \sa_snapshot[22].r.part0[9] );
tran (\sa_snapshot[22][9] , \sa_snapshot[22].f.lower[9] );
tran (\sa_snapshot[22][10] , \sa_snapshot[22].r.part0[10] );
tran (\sa_snapshot[22][10] , \sa_snapshot[22].f.lower[10] );
tran (\sa_snapshot[22][11] , \sa_snapshot[22].r.part0[11] );
tran (\sa_snapshot[22][11] , \sa_snapshot[22].f.lower[11] );
tran (\sa_snapshot[22][12] , \sa_snapshot[22].r.part0[12] );
tran (\sa_snapshot[22][12] , \sa_snapshot[22].f.lower[12] );
tran (\sa_snapshot[22][13] , \sa_snapshot[22].r.part0[13] );
tran (\sa_snapshot[22][13] , \sa_snapshot[22].f.lower[13] );
tran (\sa_snapshot[22][14] , \sa_snapshot[22].r.part0[14] );
tran (\sa_snapshot[22][14] , \sa_snapshot[22].f.lower[14] );
tran (\sa_snapshot[22][15] , \sa_snapshot[22].r.part0[15] );
tran (\sa_snapshot[22][15] , \sa_snapshot[22].f.lower[15] );
tran (\sa_snapshot[22][16] , \sa_snapshot[22].r.part0[16] );
tran (\sa_snapshot[22][16] , \sa_snapshot[22].f.lower[16] );
tran (\sa_snapshot[22][17] , \sa_snapshot[22].r.part0[17] );
tran (\sa_snapshot[22][17] , \sa_snapshot[22].f.lower[17] );
tran (\sa_snapshot[22][18] , \sa_snapshot[22].r.part0[18] );
tran (\sa_snapshot[22][18] , \sa_snapshot[22].f.lower[18] );
tran (\sa_snapshot[22][19] , \sa_snapshot[22].r.part0[19] );
tran (\sa_snapshot[22][19] , \sa_snapshot[22].f.lower[19] );
tran (\sa_snapshot[22][20] , \sa_snapshot[22].r.part0[20] );
tran (\sa_snapshot[22][20] , \sa_snapshot[22].f.lower[20] );
tran (\sa_snapshot[22][21] , \sa_snapshot[22].r.part0[21] );
tran (\sa_snapshot[22][21] , \sa_snapshot[22].f.lower[21] );
tran (\sa_snapshot[22][22] , \sa_snapshot[22].r.part0[22] );
tran (\sa_snapshot[22][22] , \sa_snapshot[22].f.lower[22] );
tran (\sa_snapshot[22][23] , \sa_snapshot[22].r.part0[23] );
tran (\sa_snapshot[22][23] , \sa_snapshot[22].f.lower[23] );
tran (\sa_snapshot[22][24] , \sa_snapshot[22].r.part0[24] );
tran (\sa_snapshot[22][24] , \sa_snapshot[22].f.lower[24] );
tran (\sa_snapshot[22][25] , \sa_snapshot[22].r.part0[25] );
tran (\sa_snapshot[22][25] , \sa_snapshot[22].f.lower[25] );
tran (\sa_snapshot[22][26] , \sa_snapshot[22].r.part0[26] );
tran (\sa_snapshot[22][26] , \sa_snapshot[22].f.lower[26] );
tran (\sa_snapshot[22][27] , \sa_snapshot[22].r.part0[27] );
tran (\sa_snapshot[22][27] , \sa_snapshot[22].f.lower[27] );
tran (\sa_snapshot[22][28] , \sa_snapshot[22].r.part0[28] );
tran (\sa_snapshot[22][28] , \sa_snapshot[22].f.lower[28] );
tran (\sa_snapshot[22][29] , \sa_snapshot[22].r.part0[29] );
tran (\sa_snapshot[22][29] , \sa_snapshot[22].f.lower[29] );
tran (\sa_snapshot[22][30] , \sa_snapshot[22].r.part0[30] );
tran (\sa_snapshot[22][30] , \sa_snapshot[22].f.lower[30] );
tran (\sa_snapshot[22][31] , \sa_snapshot[22].r.part0[31] );
tran (\sa_snapshot[22][31] , \sa_snapshot[22].f.lower[31] );
tran (\sa_snapshot[22][32] , \sa_snapshot[22].r.part1[0] );
tran (\sa_snapshot[22][32] , \sa_snapshot[22].f.upper[0] );
tran (\sa_snapshot[22][33] , \sa_snapshot[22].r.part1[1] );
tran (\sa_snapshot[22][33] , \sa_snapshot[22].f.upper[1] );
tran (\sa_snapshot[22][34] , \sa_snapshot[22].r.part1[2] );
tran (\sa_snapshot[22][34] , \sa_snapshot[22].f.upper[2] );
tran (\sa_snapshot[22][35] , \sa_snapshot[22].r.part1[3] );
tran (\sa_snapshot[22][35] , \sa_snapshot[22].f.upper[3] );
tran (\sa_snapshot[22][36] , \sa_snapshot[22].r.part1[4] );
tran (\sa_snapshot[22][36] , \sa_snapshot[22].f.upper[4] );
tran (\sa_snapshot[22][37] , \sa_snapshot[22].r.part1[5] );
tran (\sa_snapshot[22][37] , \sa_snapshot[22].f.upper[5] );
tran (\sa_snapshot[22][38] , \sa_snapshot[22].r.part1[6] );
tran (\sa_snapshot[22][38] , \sa_snapshot[22].f.upper[6] );
tran (\sa_snapshot[22][39] , \sa_snapshot[22].r.part1[7] );
tran (\sa_snapshot[22][39] , \sa_snapshot[22].f.upper[7] );
tran (\sa_snapshot[22][40] , \sa_snapshot[22].r.part1[8] );
tran (\sa_snapshot[22][40] , \sa_snapshot[22].f.upper[8] );
tran (\sa_snapshot[22][41] , \sa_snapshot[22].r.part1[9] );
tran (\sa_snapshot[22][41] , \sa_snapshot[22].f.upper[9] );
tran (\sa_snapshot[22][42] , \sa_snapshot[22].r.part1[10] );
tran (\sa_snapshot[22][42] , \sa_snapshot[22].f.upper[10] );
tran (\sa_snapshot[22][43] , \sa_snapshot[22].r.part1[11] );
tran (\sa_snapshot[22][43] , \sa_snapshot[22].f.upper[11] );
tran (\sa_snapshot[22][44] , \sa_snapshot[22].r.part1[12] );
tran (\sa_snapshot[22][44] , \sa_snapshot[22].f.upper[12] );
tran (\sa_snapshot[22][45] , \sa_snapshot[22].r.part1[13] );
tran (\sa_snapshot[22][45] , \sa_snapshot[22].f.upper[13] );
tran (\sa_snapshot[22][46] , \sa_snapshot[22].r.part1[14] );
tran (\sa_snapshot[22][46] , \sa_snapshot[22].f.upper[14] );
tran (\sa_snapshot[22][47] , \sa_snapshot[22].r.part1[15] );
tran (\sa_snapshot[22][47] , \sa_snapshot[22].f.upper[15] );
tran (\sa_snapshot[22][48] , \sa_snapshot[22].r.part1[16] );
tran (\sa_snapshot[22][48] , \sa_snapshot[22].f.upper[16] );
tran (\sa_snapshot[22][49] , \sa_snapshot[22].r.part1[17] );
tran (\sa_snapshot[22][49] , \sa_snapshot[22].f.upper[17] );
tran (\sa_snapshot[22][50] , \sa_snapshot[22].r.part1[18] );
tran (\sa_snapshot[22][50] , \sa_snapshot[22].f.unused[0] );
tran (\sa_snapshot[22][51] , \sa_snapshot[22].r.part1[19] );
tran (\sa_snapshot[22][51] , \sa_snapshot[22].f.unused[1] );
tran (\sa_snapshot[22][52] , \sa_snapshot[22].r.part1[20] );
tran (\sa_snapshot[22][52] , \sa_snapshot[22].f.unused[2] );
tran (\sa_snapshot[22][53] , \sa_snapshot[22].r.part1[21] );
tran (\sa_snapshot[22][53] , \sa_snapshot[22].f.unused[3] );
tran (\sa_snapshot[22][54] , \sa_snapshot[22].r.part1[22] );
tran (\sa_snapshot[22][54] , \sa_snapshot[22].f.unused[4] );
tran (\sa_snapshot[22][55] , \sa_snapshot[22].r.part1[23] );
tran (\sa_snapshot[22][55] , \sa_snapshot[22].f.unused[5] );
tran (\sa_snapshot[22][56] , \sa_snapshot[22].r.part1[24] );
tran (\sa_snapshot[22][56] , \sa_snapshot[22].f.unused[6] );
tran (\sa_snapshot[22][57] , \sa_snapshot[22].r.part1[25] );
tran (\sa_snapshot[22][57] , \sa_snapshot[22].f.unused[7] );
tran (\sa_snapshot[22][58] , \sa_snapshot[22].r.part1[26] );
tran (\sa_snapshot[22][58] , \sa_snapshot[22].f.unused[8] );
tran (\sa_snapshot[22][59] , \sa_snapshot[22].r.part1[27] );
tran (\sa_snapshot[22][59] , \sa_snapshot[22].f.unused[9] );
tran (\sa_snapshot[22][60] , \sa_snapshot[22].r.part1[28] );
tran (\sa_snapshot[22][60] , \sa_snapshot[22].f.unused[10] );
tran (\sa_snapshot[22][61] , \sa_snapshot[22].r.part1[29] );
tran (\sa_snapshot[22][61] , \sa_snapshot[22].f.unused[11] );
tran (\sa_snapshot[22][62] , \sa_snapshot[22].r.part1[30] );
tran (\sa_snapshot[22][62] , \sa_snapshot[22].f.unused[12] );
tran (\sa_snapshot[22][63] , \sa_snapshot[22].r.part1[31] );
tran (\sa_snapshot[22][63] , \sa_snapshot[22].f.unused[13] );
tran (\sa_snapshot[23][0] , \sa_snapshot[23].r.part0[0] );
tran (\sa_snapshot[23][0] , \sa_snapshot[23].f.lower[0] );
tran (\sa_snapshot[23][1] , \sa_snapshot[23].r.part0[1] );
tran (\sa_snapshot[23][1] , \sa_snapshot[23].f.lower[1] );
tran (\sa_snapshot[23][2] , \sa_snapshot[23].r.part0[2] );
tran (\sa_snapshot[23][2] , \sa_snapshot[23].f.lower[2] );
tran (\sa_snapshot[23][3] , \sa_snapshot[23].r.part0[3] );
tran (\sa_snapshot[23][3] , \sa_snapshot[23].f.lower[3] );
tran (\sa_snapshot[23][4] , \sa_snapshot[23].r.part0[4] );
tran (\sa_snapshot[23][4] , \sa_snapshot[23].f.lower[4] );
tran (\sa_snapshot[23][5] , \sa_snapshot[23].r.part0[5] );
tran (\sa_snapshot[23][5] , \sa_snapshot[23].f.lower[5] );
tran (\sa_snapshot[23][6] , \sa_snapshot[23].r.part0[6] );
tran (\sa_snapshot[23][6] , \sa_snapshot[23].f.lower[6] );
tran (\sa_snapshot[23][7] , \sa_snapshot[23].r.part0[7] );
tran (\sa_snapshot[23][7] , \sa_snapshot[23].f.lower[7] );
tran (\sa_snapshot[23][8] , \sa_snapshot[23].r.part0[8] );
tran (\sa_snapshot[23][8] , \sa_snapshot[23].f.lower[8] );
tran (\sa_snapshot[23][9] , \sa_snapshot[23].r.part0[9] );
tran (\sa_snapshot[23][9] , \sa_snapshot[23].f.lower[9] );
tran (\sa_snapshot[23][10] , \sa_snapshot[23].r.part0[10] );
tran (\sa_snapshot[23][10] , \sa_snapshot[23].f.lower[10] );
tran (\sa_snapshot[23][11] , \sa_snapshot[23].r.part0[11] );
tran (\sa_snapshot[23][11] , \sa_snapshot[23].f.lower[11] );
tran (\sa_snapshot[23][12] , \sa_snapshot[23].r.part0[12] );
tran (\sa_snapshot[23][12] , \sa_snapshot[23].f.lower[12] );
tran (\sa_snapshot[23][13] , \sa_snapshot[23].r.part0[13] );
tran (\sa_snapshot[23][13] , \sa_snapshot[23].f.lower[13] );
tran (\sa_snapshot[23][14] , \sa_snapshot[23].r.part0[14] );
tran (\sa_snapshot[23][14] , \sa_snapshot[23].f.lower[14] );
tran (\sa_snapshot[23][15] , \sa_snapshot[23].r.part0[15] );
tran (\sa_snapshot[23][15] , \sa_snapshot[23].f.lower[15] );
tran (\sa_snapshot[23][16] , \sa_snapshot[23].r.part0[16] );
tran (\sa_snapshot[23][16] , \sa_snapshot[23].f.lower[16] );
tran (\sa_snapshot[23][17] , \sa_snapshot[23].r.part0[17] );
tran (\sa_snapshot[23][17] , \sa_snapshot[23].f.lower[17] );
tran (\sa_snapshot[23][18] , \sa_snapshot[23].r.part0[18] );
tran (\sa_snapshot[23][18] , \sa_snapshot[23].f.lower[18] );
tran (\sa_snapshot[23][19] , \sa_snapshot[23].r.part0[19] );
tran (\sa_snapshot[23][19] , \sa_snapshot[23].f.lower[19] );
tran (\sa_snapshot[23][20] , \sa_snapshot[23].r.part0[20] );
tran (\sa_snapshot[23][20] , \sa_snapshot[23].f.lower[20] );
tran (\sa_snapshot[23][21] , \sa_snapshot[23].r.part0[21] );
tran (\sa_snapshot[23][21] , \sa_snapshot[23].f.lower[21] );
tran (\sa_snapshot[23][22] , \sa_snapshot[23].r.part0[22] );
tran (\sa_snapshot[23][22] , \sa_snapshot[23].f.lower[22] );
tran (\sa_snapshot[23][23] , \sa_snapshot[23].r.part0[23] );
tran (\sa_snapshot[23][23] , \sa_snapshot[23].f.lower[23] );
tran (\sa_snapshot[23][24] , \sa_snapshot[23].r.part0[24] );
tran (\sa_snapshot[23][24] , \sa_snapshot[23].f.lower[24] );
tran (\sa_snapshot[23][25] , \sa_snapshot[23].r.part0[25] );
tran (\sa_snapshot[23][25] , \sa_snapshot[23].f.lower[25] );
tran (\sa_snapshot[23][26] , \sa_snapshot[23].r.part0[26] );
tran (\sa_snapshot[23][26] , \sa_snapshot[23].f.lower[26] );
tran (\sa_snapshot[23][27] , \sa_snapshot[23].r.part0[27] );
tran (\sa_snapshot[23][27] , \sa_snapshot[23].f.lower[27] );
tran (\sa_snapshot[23][28] , \sa_snapshot[23].r.part0[28] );
tran (\sa_snapshot[23][28] , \sa_snapshot[23].f.lower[28] );
tran (\sa_snapshot[23][29] , \sa_snapshot[23].r.part0[29] );
tran (\sa_snapshot[23][29] , \sa_snapshot[23].f.lower[29] );
tran (\sa_snapshot[23][30] , \sa_snapshot[23].r.part0[30] );
tran (\sa_snapshot[23][30] , \sa_snapshot[23].f.lower[30] );
tran (\sa_snapshot[23][31] , \sa_snapshot[23].r.part0[31] );
tran (\sa_snapshot[23][31] , \sa_snapshot[23].f.lower[31] );
tran (\sa_snapshot[23][32] , \sa_snapshot[23].r.part1[0] );
tran (\sa_snapshot[23][32] , \sa_snapshot[23].f.upper[0] );
tran (\sa_snapshot[23][33] , \sa_snapshot[23].r.part1[1] );
tran (\sa_snapshot[23][33] , \sa_snapshot[23].f.upper[1] );
tran (\sa_snapshot[23][34] , \sa_snapshot[23].r.part1[2] );
tran (\sa_snapshot[23][34] , \sa_snapshot[23].f.upper[2] );
tran (\sa_snapshot[23][35] , \sa_snapshot[23].r.part1[3] );
tran (\sa_snapshot[23][35] , \sa_snapshot[23].f.upper[3] );
tran (\sa_snapshot[23][36] , \sa_snapshot[23].r.part1[4] );
tran (\sa_snapshot[23][36] , \sa_snapshot[23].f.upper[4] );
tran (\sa_snapshot[23][37] , \sa_snapshot[23].r.part1[5] );
tran (\sa_snapshot[23][37] , \sa_snapshot[23].f.upper[5] );
tran (\sa_snapshot[23][38] , \sa_snapshot[23].r.part1[6] );
tran (\sa_snapshot[23][38] , \sa_snapshot[23].f.upper[6] );
tran (\sa_snapshot[23][39] , \sa_snapshot[23].r.part1[7] );
tran (\sa_snapshot[23][39] , \sa_snapshot[23].f.upper[7] );
tran (\sa_snapshot[23][40] , \sa_snapshot[23].r.part1[8] );
tran (\sa_snapshot[23][40] , \sa_snapshot[23].f.upper[8] );
tran (\sa_snapshot[23][41] , \sa_snapshot[23].r.part1[9] );
tran (\sa_snapshot[23][41] , \sa_snapshot[23].f.upper[9] );
tran (\sa_snapshot[23][42] , \sa_snapshot[23].r.part1[10] );
tran (\sa_snapshot[23][42] , \sa_snapshot[23].f.upper[10] );
tran (\sa_snapshot[23][43] , \sa_snapshot[23].r.part1[11] );
tran (\sa_snapshot[23][43] , \sa_snapshot[23].f.upper[11] );
tran (\sa_snapshot[23][44] , \sa_snapshot[23].r.part1[12] );
tran (\sa_snapshot[23][44] , \sa_snapshot[23].f.upper[12] );
tran (\sa_snapshot[23][45] , \sa_snapshot[23].r.part1[13] );
tran (\sa_snapshot[23][45] , \sa_snapshot[23].f.upper[13] );
tran (\sa_snapshot[23][46] , \sa_snapshot[23].r.part1[14] );
tran (\sa_snapshot[23][46] , \sa_snapshot[23].f.upper[14] );
tran (\sa_snapshot[23][47] , \sa_snapshot[23].r.part1[15] );
tran (\sa_snapshot[23][47] , \sa_snapshot[23].f.upper[15] );
tran (\sa_snapshot[23][48] , \sa_snapshot[23].r.part1[16] );
tran (\sa_snapshot[23][48] , \sa_snapshot[23].f.upper[16] );
tran (\sa_snapshot[23][49] , \sa_snapshot[23].r.part1[17] );
tran (\sa_snapshot[23][49] , \sa_snapshot[23].f.upper[17] );
tran (\sa_snapshot[23][50] , \sa_snapshot[23].r.part1[18] );
tran (\sa_snapshot[23][50] , \sa_snapshot[23].f.unused[0] );
tran (\sa_snapshot[23][51] , \sa_snapshot[23].r.part1[19] );
tran (\sa_snapshot[23][51] , \sa_snapshot[23].f.unused[1] );
tran (\sa_snapshot[23][52] , \sa_snapshot[23].r.part1[20] );
tran (\sa_snapshot[23][52] , \sa_snapshot[23].f.unused[2] );
tran (\sa_snapshot[23][53] , \sa_snapshot[23].r.part1[21] );
tran (\sa_snapshot[23][53] , \sa_snapshot[23].f.unused[3] );
tran (\sa_snapshot[23][54] , \sa_snapshot[23].r.part1[22] );
tran (\sa_snapshot[23][54] , \sa_snapshot[23].f.unused[4] );
tran (\sa_snapshot[23][55] , \sa_snapshot[23].r.part1[23] );
tran (\sa_snapshot[23][55] , \sa_snapshot[23].f.unused[5] );
tran (\sa_snapshot[23][56] , \sa_snapshot[23].r.part1[24] );
tran (\sa_snapshot[23][56] , \sa_snapshot[23].f.unused[6] );
tran (\sa_snapshot[23][57] , \sa_snapshot[23].r.part1[25] );
tran (\sa_snapshot[23][57] , \sa_snapshot[23].f.unused[7] );
tran (\sa_snapshot[23][58] , \sa_snapshot[23].r.part1[26] );
tran (\sa_snapshot[23][58] , \sa_snapshot[23].f.unused[8] );
tran (\sa_snapshot[23][59] , \sa_snapshot[23].r.part1[27] );
tran (\sa_snapshot[23][59] , \sa_snapshot[23].f.unused[9] );
tran (\sa_snapshot[23][60] , \sa_snapshot[23].r.part1[28] );
tran (\sa_snapshot[23][60] , \sa_snapshot[23].f.unused[10] );
tran (\sa_snapshot[23][61] , \sa_snapshot[23].r.part1[29] );
tran (\sa_snapshot[23][61] , \sa_snapshot[23].f.unused[11] );
tran (\sa_snapshot[23][62] , \sa_snapshot[23].r.part1[30] );
tran (\sa_snapshot[23][62] , \sa_snapshot[23].f.unused[12] );
tran (\sa_snapshot[23][63] , \sa_snapshot[23].r.part1[31] );
tran (\sa_snapshot[23][63] , \sa_snapshot[23].f.unused[13] );
tran (\sa_snapshot[24][0] , \sa_snapshot[24].r.part0[0] );
tran (\sa_snapshot[24][0] , \sa_snapshot[24].f.lower[0] );
tran (\sa_snapshot[24][1] , \sa_snapshot[24].r.part0[1] );
tran (\sa_snapshot[24][1] , \sa_snapshot[24].f.lower[1] );
tran (\sa_snapshot[24][2] , \sa_snapshot[24].r.part0[2] );
tran (\sa_snapshot[24][2] , \sa_snapshot[24].f.lower[2] );
tran (\sa_snapshot[24][3] , \sa_snapshot[24].r.part0[3] );
tran (\sa_snapshot[24][3] , \sa_snapshot[24].f.lower[3] );
tran (\sa_snapshot[24][4] , \sa_snapshot[24].r.part0[4] );
tran (\sa_snapshot[24][4] , \sa_snapshot[24].f.lower[4] );
tran (\sa_snapshot[24][5] , \sa_snapshot[24].r.part0[5] );
tran (\sa_snapshot[24][5] , \sa_snapshot[24].f.lower[5] );
tran (\sa_snapshot[24][6] , \sa_snapshot[24].r.part0[6] );
tran (\sa_snapshot[24][6] , \sa_snapshot[24].f.lower[6] );
tran (\sa_snapshot[24][7] , \sa_snapshot[24].r.part0[7] );
tran (\sa_snapshot[24][7] , \sa_snapshot[24].f.lower[7] );
tran (\sa_snapshot[24][8] , \sa_snapshot[24].r.part0[8] );
tran (\sa_snapshot[24][8] , \sa_snapshot[24].f.lower[8] );
tran (\sa_snapshot[24][9] , \sa_snapshot[24].r.part0[9] );
tran (\sa_snapshot[24][9] , \sa_snapshot[24].f.lower[9] );
tran (\sa_snapshot[24][10] , \sa_snapshot[24].r.part0[10] );
tran (\sa_snapshot[24][10] , \sa_snapshot[24].f.lower[10] );
tran (\sa_snapshot[24][11] , \sa_snapshot[24].r.part0[11] );
tran (\sa_snapshot[24][11] , \sa_snapshot[24].f.lower[11] );
tran (\sa_snapshot[24][12] , \sa_snapshot[24].r.part0[12] );
tran (\sa_snapshot[24][12] , \sa_snapshot[24].f.lower[12] );
tran (\sa_snapshot[24][13] , \sa_snapshot[24].r.part0[13] );
tran (\sa_snapshot[24][13] , \sa_snapshot[24].f.lower[13] );
tran (\sa_snapshot[24][14] , \sa_snapshot[24].r.part0[14] );
tran (\sa_snapshot[24][14] , \sa_snapshot[24].f.lower[14] );
tran (\sa_snapshot[24][15] , \sa_snapshot[24].r.part0[15] );
tran (\sa_snapshot[24][15] , \sa_snapshot[24].f.lower[15] );
tran (\sa_snapshot[24][16] , \sa_snapshot[24].r.part0[16] );
tran (\sa_snapshot[24][16] , \sa_snapshot[24].f.lower[16] );
tran (\sa_snapshot[24][17] , \sa_snapshot[24].r.part0[17] );
tran (\sa_snapshot[24][17] , \sa_snapshot[24].f.lower[17] );
tran (\sa_snapshot[24][18] , \sa_snapshot[24].r.part0[18] );
tran (\sa_snapshot[24][18] , \sa_snapshot[24].f.lower[18] );
tran (\sa_snapshot[24][19] , \sa_snapshot[24].r.part0[19] );
tran (\sa_snapshot[24][19] , \sa_snapshot[24].f.lower[19] );
tran (\sa_snapshot[24][20] , \sa_snapshot[24].r.part0[20] );
tran (\sa_snapshot[24][20] , \sa_snapshot[24].f.lower[20] );
tran (\sa_snapshot[24][21] , \sa_snapshot[24].r.part0[21] );
tran (\sa_snapshot[24][21] , \sa_snapshot[24].f.lower[21] );
tran (\sa_snapshot[24][22] , \sa_snapshot[24].r.part0[22] );
tran (\sa_snapshot[24][22] , \sa_snapshot[24].f.lower[22] );
tran (\sa_snapshot[24][23] , \sa_snapshot[24].r.part0[23] );
tran (\sa_snapshot[24][23] , \sa_snapshot[24].f.lower[23] );
tran (\sa_snapshot[24][24] , \sa_snapshot[24].r.part0[24] );
tran (\sa_snapshot[24][24] , \sa_snapshot[24].f.lower[24] );
tran (\sa_snapshot[24][25] , \sa_snapshot[24].r.part0[25] );
tran (\sa_snapshot[24][25] , \sa_snapshot[24].f.lower[25] );
tran (\sa_snapshot[24][26] , \sa_snapshot[24].r.part0[26] );
tran (\sa_snapshot[24][26] , \sa_snapshot[24].f.lower[26] );
tran (\sa_snapshot[24][27] , \sa_snapshot[24].r.part0[27] );
tran (\sa_snapshot[24][27] , \sa_snapshot[24].f.lower[27] );
tran (\sa_snapshot[24][28] , \sa_snapshot[24].r.part0[28] );
tran (\sa_snapshot[24][28] , \sa_snapshot[24].f.lower[28] );
tran (\sa_snapshot[24][29] , \sa_snapshot[24].r.part0[29] );
tran (\sa_snapshot[24][29] , \sa_snapshot[24].f.lower[29] );
tran (\sa_snapshot[24][30] , \sa_snapshot[24].r.part0[30] );
tran (\sa_snapshot[24][30] , \sa_snapshot[24].f.lower[30] );
tran (\sa_snapshot[24][31] , \sa_snapshot[24].r.part0[31] );
tran (\sa_snapshot[24][31] , \sa_snapshot[24].f.lower[31] );
tran (\sa_snapshot[24][32] , \sa_snapshot[24].r.part1[0] );
tran (\sa_snapshot[24][32] , \sa_snapshot[24].f.upper[0] );
tran (\sa_snapshot[24][33] , \sa_snapshot[24].r.part1[1] );
tran (\sa_snapshot[24][33] , \sa_snapshot[24].f.upper[1] );
tran (\sa_snapshot[24][34] , \sa_snapshot[24].r.part1[2] );
tran (\sa_snapshot[24][34] , \sa_snapshot[24].f.upper[2] );
tran (\sa_snapshot[24][35] , \sa_snapshot[24].r.part1[3] );
tran (\sa_snapshot[24][35] , \sa_snapshot[24].f.upper[3] );
tran (\sa_snapshot[24][36] , \sa_snapshot[24].r.part1[4] );
tran (\sa_snapshot[24][36] , \sa_snapshot[24].f.upper[4] );
tran (\sa_snapshot[24][37] , \sa_snapshot[24].r.part1[5] );
tran (\sa_snapshot[24][37] , \sa_snapshot[24].f.upper[5] );
tran (\sa_snapshot[24][38] , \sa_snapshot[24].r.part1[6] );
tran (\sa_snapshot[24][38] , \sa_snapshot[24].f.upper[6] );
tran (\sa_snapshot[24][39] , \sa_snapshot[24].r.part1[7] );
tran (\sa_snapshot[24][39] , \sa_snapshot[24].f.upper[7] );
tran (\sa_snapshot[24][40] , \sa_snapshot[24].r.part1[8] );
tran (\sa_snapshot[24][40] , \sa_snapshot[24].f.upper[8] );
tran (\sa_snapshot[24][41] , \sa_snapshot[24].r.part1[9] );
tran (\sa_snapshot[24][41] , \sa_snapshot[24].f.upper[9] );
tran (\sa_snapshot[24][42] , \sa_snapshot[24].r.part1[10] );
tran (\sa_snapshot[24][42] , \sa_snapshot[24].f.upper[10] );
tran (\sa_snapshot[24][43] , \sa_snapshot[24].r.part1[11] );
tran (\sa_snapshot[24][43] , \sa_snapshot[24].f.upper[11] );
tran (\sa_snapshot[24][44] , \sa_snapshot[24].r.part1[12] );
tran (\sa_snapshot[24][44] , \sa_snapshot[24].f.upper[12] );
tran (\sa_snapshot[24][45] , \sa_snapshot[24].r.part1[13] );
tran (\sa_snapshot[24][45] , \sa_snapshot[24].f.upper[13] );
tran (\sa_snapshot[24][46] , \sa_snapshot[24].r.part1[14] );
tran (\sa_snapshot[24][46] , \sa_snapshot[24].f.upper[14] );
tran (\sa_snapshot[24][47] , \sa_snapshot[24].r.part1[15] );
tran (\sa_snapshot[24][47] , \sa_snapshot[24].f.upper[15] );
tran (\sa_snapshot[24][48] , \sa_snapshot[24].r.part1[16] );
tran (\sa_snapshot[24][48] , \sa_snapshot[24].f.upper[16] );
tran (\sa_snapshot[24][49] , \sa_snapshot[24].r.part1[17] );
tran (\sa_snapshot[24][49] , \sa_snapshot[24].f.upper[17] );
tran (\sa_snapshot[24][50] , \sa_snapshot[24].r.part1[18] );
tran (\sa_snapshot[24][50] , \sa_snapshot[24].f.unused[0] );
tran (\sa_snapshot[24][51] , \sa_snapshot[24].r.part1[19] );
tran (\sa_snapshot[24][51] , \sa_snapshot[24].f.unused[1] );
tran (\sa_snapshot[24][52] , \sa_snapshot[24].r.part1[20] );
tran (\sa_snapshot[24][52] , \sa_snapshot[24].f.unused[2] );
tran (\sa_snapshot[24][53] , \sa_snapshot[24].r.part1[21] );
tran (\sa_snapshot[24][53] , \sa_snapshot[24].f.unused[3] );
tran (\sa_snapshot[24][54] , \sa_snapshot[24].r.part1[22] );
tran (\sa_snapshot[24][54] , \sa_snapshot[24].f.unused[4] );
tran (\sa_snapshot[24][55] , \sa_snapshot[24].r.part1[23] );
tran (\sa_snapshot[24][55] , \sa_snapshot[24].f.unused[5] );
tran (\sa_snapshot[24][56] , \sa_snapshot[24].r.part1[24] );
tran (\sa_snapshot[24][56] , \sa_snapshot[24].f.unused[6] );
tran (\sa_snapshot[24][57] , \sa_snapshot[24].r.part1[25] );
tran (\sa_snapshot[24][57] , \sa_snapshot[24].f.unused[7] );
tran (\sa_snapshot[24][58] , \sa_snapshot[24].r.part1[26] );
tran (\sa_snapshot[24][58] , \sa_snapshot[24].f.unused[8] );
tran (\sa_snapshot[24][59] , \sa_snapshot[24].r.part1[27] );
tran (\sa_snapshot[24][59] , \sa_snapshot[24].f.unused[9] );
tran (\sa_snapshot[24][60] , \sa_snapshot[24].r.part1[28] );
tran (\sa_snapshot[24][60] , \sa_snapshot[24].f.unused[10] );
tran (\sa_snapshot[24][61] , \sa_snapshot[24].r.part1[29] );
tran (\sa_snapshot[24][61] , \sa_snapshot[24].f.unused[11] );
tran (\sa_snapshot[24][62] , \sa_snapshot[24].r.part1[30] );
tran (\sa_snapshot[24][62] , \sa_snapshot[24].f.unused[12] );
tran (\sa_snapshot[24][63] , \sa_snapshot[24].r.part1[31] );
tran (\sa_snapshot[24][63] , \sa_snapshot[24].f.unused[13] );
tran (\sa_snapshot[25][0] , \sa_snapshot[25].r.part0[0] );
tran (\sa_snapshot[25][0] , \sa_snapshot[25].f.lower[0] );
tran (\sa_snapshot[25][1] , \sa_snapshot[25].r.part0[1] );
tran (\sa_snapshot[25][1] , \sa_snapshot[25].f.lower[1] );
tran (\sa_snapshot[25][2] , \sa_snapshot[25].r.part0[2] );
tran (\sa_snapshot[25][2] , \sa_snapshot[25].f.lower[2] );
tran (\sa_snapshot[25][3] , \sa_snapshot[25].r.part0[3] );
tran (\sa_snapshot[25][3] , \sa_snapshot[25].f.lower[3] );
tran (\sa_snapshot[25][4] , \sa_snapshot[25].r.part0[4] );
tran (\sa_snapshot[25][4] , \sa_snapshot[25].f.lower[4] );
tran (\sa_snapshot[25][5] , \sa_snapshot[25].r.part0[5] );
tran (\sa_snapshot[25][5] , \sa_snapshot[25].f.lower[5] );
tran (\sa_snapshot[25][6] , \sa_snapshot[25].r.part0[6] );
tran (\sa_snapshot[25][6] , \sa_snapshot[25].f.lower[6] );
tran (\sa_snapshot[25][7] , \sa_snapshot[25].r.part0[7] );
tran (\sa_snapshot[25][7] , \sa_snapshot[25].f.lower[7] );
tran (\sa_snapshot[25][8] , \sa_snapshot[25].r.part0[8] );
tran (\sa_snapshot[25][8] , \sa_snapshot[25].f.lower[8] );
tran (\sa_snapshot[25][9] , \sa_snapshot[25].r.part0[9] );
tran (\sa_snapshot[25][9] , \sa_snapshot[25].f.lower[9] );
tran (\sa_snapshot[25][10] , \sa_snapshot[25].r.part0[10] );
tran (\sa_snapshot[25][10] , \sa_snapshot[25].f.lower[10] );
tran (\sa_snapshot[25][11] , \sa_snapshot[25].r.part0[11] );
tran (\sa_snapshot[25][11] , \sa_snapshot[25].f.lower[11] );
tran (\sa_snapshot[25][12] , \sa_snapshot[25].r.part0[12] );
tran (\sa_snapshot[25][12] , \sa_snapshot[25].f.lower[12] );
tran (\sa_snapshot[25][13] , \sa_snapshot[25].r.part0[13] );
tran (\sa_snapshot[25][13] , \sa_snapshot[25].f.lower[13] );
tran (\sa_snapshot[25][14] , \sa_snapshot[25].r.part0[14] );
tran (\sa_snapshot[25][14] , \sa_snapshot[25].f.lower[14] );
tran (\sa_snapshot[25][15] , \sa_snapshot[25].r.part0[15] );
tran (\sa_snapshot[25][15] , \sa_snapshot[25].f.lower[15] );
tran (\sa_snapshot[25][16] , \sa_snapshot[25].r.part0[16] );
tran (\sa_snapshot[25][16] , \sa_snapshot[25].f.lower[16] );
tran (\sa_snapshot[25][17] , \sa_snapshot[25].r.part0[17] );
tran (\sa_snapshot[25][17] , \sa_snapshot[25].f.lower[17] );
tran (\sa_snapshot[25][18] , \sa_snapshot[25].r.part0[18] );
tran (\sa_snapshot[25][18] , \sa_snapshot[25].f.lower[18] );
tran (\sa_snapshot[25][19] , \sa_snapshot[25].r.part0[19] );
tran (\sa_snapshot[25][19] , \sa_snapshot[25].f.lower[19] );
tran (\sa_snapshot[25][20] , \sa_snapshot[25].r.part0[20] );
tran (\sa_snapshot[25][20] , \sa_snapshot[25].f.lower[20] );
tran (\sa_snapshot[25][21] , \sa_snapshot[25].r.part0[21] );
tran (\sa_snapshot[25][21] , \sa_snapshot[25].f.lower[21] );
tran (\sa_snapshot[25][22] , \sa_snapshot[25].r.part0[22] );
tran (\sa_snapshot[25][22] , \sa_snapshot[25].f.lower[22] );
tran (\sa_snapshot[25][23] , \sa_snapshot[25].r.part0[23] );
tran (\sa_snapshot[25][23] , \sa_snapshot[25].f.lower[23] );
tran (\sa_snapshot[25][24] , \sa_snapshot[25].r.part0[24] );
tran (\sa_snapshot[25][24] , \sa_snapshot[25].f.lower[24] );
tran (\sa_snapshot[25][25] , \sa_snapshot[25].r.part0[25] );
tran (\sa_snapshot[25][25] , \sa_snapshot[25].f.lower[25] );
tran (\sa_snapshot[25][26] , \sa_snapshot[25].r.part0[26] );
tran (\sa_snapshot[25][26] , \sa_snapshot[25].f.lower[26] );
tran (\sa_snapshot[25][27] , \sa_snapshot[25].r.part0[27] );
tran (\sa_snapshot[25][27] , \sa_snapshot[25].f.lower[27] );
tran (\sa_snapshot[25][28] , \sa_snapshot[25].r.part0[28] );
tran (\sa_snapshot[25][28] , \sa_snapshot[25].f.lower[28] );
tran (\sa_snapshot[25][29] , \sa_snapshot[25].r.part0[29] );
tran (\sa_snapshot[25][29] , \sa_snapshot[25].f.lower[29] );
tran (\sa_snapshot[25][30] , \sa_snapshot[25].r.part0[30] );
tran (\sa_snapshot[25][30] , \sa_snapshot[25].f.lower[30] );
tran (\sa_snapshot[25][31] , \sa_snapshot[25].r.part0[31] );
tran (\sa_snapshot[25][31] , \sa_snapshot[25].f.lower[31] );
tran (\sa_snapshot[25][32] , \sa_snapshot[25].r.part1[0] );
tran (\sa_snapshot[25][32] , \sa_snapshot[25].f.upper[0] );
tran (\sa_snapshot[25][33] , \sa_snapshot[25].r.part1[1] );
tran (\sa_snapshot[25][33] , \sa_snapshot[25].f.upper[1] );
tran (\sa_snapshot[25][34] , \sa_snapshot[25].r.part1[2] );
tran (\sa_snapshot[25][34] , \sa_snapshot[25].f.upper[2] );
tran (\sa_snapshot[25][35] , \sa_snapshot[25].r.part1[3] );
tran (\sa_snapshot[25][35] , \sa_snapshot[25].f.upper[3] );
tran (\sa_snapshot[25][36] , \sa_snapshot[25].r.part1[4] );
tran (\sa_snapshot[25][36] , \sa_snapshot[25].f.upper[4] );
tran (\sa_snapshot[25][37] , \sa_snapshot[25].r.part1[5] );
tran (\sa_snapshot[25][37] , \sa_snapshot[25].f.upper[5] );
tran (\sa_snapshot[25][38] , \sa_snapshot[25].r.part1[6] );
tran (\sa_snapshot[25][38] , \sa_snapshot[25].f.upper[6] );
tran (\sa_snapshot[25][39] , \sa_snapshot[25].r.part1[7] );
tran (\sa_snapshot[25][39] , \sa_snapshot[25].f.upper[7] );
tran (\sa_snapshot[25][40] , \sa_snapshot[25].r.part1[8] );
tran (\sa_snapshot[25][40] , \sa_snapshot[25].f.upper[8] );
tran (\sa_snapshot[25][41] , \sa_snapshot[25].r.part1[9] );
tran (\sa_snapshot[25][41] , \sa_snapshot[25].f.upper[9] );
tran (\sa_snapshot[25][42] , \sa_snapshot[25].r.part1[10] );
tran (\sa_snapshot[25][42] , \sa_snapshot[25].f.upper[10] );
tran (\sa_snapshot[25][43] , \sa_snapshot[25].r.part1[11] );
tran (\sa_snapshot[25][43] , \sa_snapshot[25].f.upper[11] );
tran (\sa_snapshot[25][44] , \sa_snapshot[25].r.part1[12] );
tran (\sa_snapshot[25][44] , \sa_snapshot[25].f.upper[12] );
tran (\sa_snapshot[25][45] , \sa_snapshot[25].r.part1[13] );
tran (\sa_snapshot[25][45] , \sa_snapshot[25].f.upper[13] );
tran (\sa_snapshot[25][46] , \sa_snapshot[25].r.part1[14] );
tran (\sa_snapshot[25][46] , \sa_snapshot[25].f.upper[14] );
tran (\sa_snapshot[25][47] , \sa_snapshot[25].r.part1[15] );
tran (\sa_snapshot[25][47] , \sa_snapshot[25].f.upper[15] );
tran (\sa_snapshot[25][48] , \sa_snapshot[25].r.part1[16] );
tran (\sa_snapshot[25][48] , \sa_snapshot[25].f.upper[16] );
tran (\sa_snapshot[25][49] , \sa_snapshot[25].r.part1[17] );
tran (\sa_snapshot[25][49] , \sa_snapshot[25].f.upper[17] );
tran (\sa_snapshot[25][50] , \sa_snapshot[25].r.part1[18] );
tran (\sa_snapshot[25][50] , \sa_snapshot[25].f.unused[0] );
tran (\sa_snapshot[25][51] , \sa_snapshot[25].r.part1[19] );
tran (\sa_snapshot[25][51] , \sa_snapshot[25].f.unused[1] );
tran (\sa_snapshot[25][52] , \sa_snapshot[25].r.part1[20] );
tran (\sa_snapshot[25][52] , \sa_snapshot[25].f.unused[2] );
tran (\sa_snapshot[25][53] , \sa_snapshot[25].r.part1[21] );
tran (\sa_snapshot[25][53] , \sa_snapshot[25].f.unused[3] );
tran (\sa_snapshot[25][54] , \sa_snapshot[25].r.part1[22] );
tran (\sa_snapshot[25][54] , \sa_snapshot[25].f.unused[4] );
tran (\sa_snapshot[25][55] , \sa_snapshot[25].r.part1[23] );
tran (\sa_snapshot[25][55] , \sa_snapshot[25].f.unused[5] );
tran (\sa_snapshot[25][56] , \sa_snapshot[25].r.part1[24] );
tran (\sa_snapshot[25][56] , \sa_snapshot[25].f.unused[6] );
tran (\sa_snapshot[25][57] , \sa_snapshot[25].r.part1[25] );
tran (\sa_snapshot[25][57] , \sa_snapshot[25].f.unused[7] );
tran (\sa_snapshot[25][58] , \sa_snapshot[25].r.part1[26] );
tran (\sa_snapshot[25][58] , \sa_snapshot[25].f.unused[8] );
tran (\sa_snapshot[25][59] , \sa_snapshot[25].r.part1[27] );
tran (\sa_snapshot[25][59] , \sa_snapshot[25].f.unused[9] );
tran (\sa_snapshot[25][60] , \sa_snapshot[25].r.part1[28] );
tran (\sa_snapshot[25][60] , \sa_snapshot[25].f.unused[10] );
tran (\sa_snapshot[25][61] , \sa_snapshot[25].r.part1[29] );
tran (\sa_snapshot[25][61] , \sa_snapshot[25].f.unused[11] );
tran (\sa_snapshot[25][62] , \sa_snapshot[25].r.part1[30] );
tran (\sa_snapshot[25][62] , \sa_snapshot[25].f.unused[12] );
tran (\sa_snapshot[25][63] , \sa_snapshot[25].r.part1[31] );
tran (\sa_snapshot[25][63] , \sa_snapshot[25].f.unused[13] );
tran (\sa_snapshot[26][0] , \sa_snapshot[26].r.part0[0] );
tran (\sa_snapshot[26][0] , \sa_snapshot[26].f.lower[0] );
tran (\sa_snapshot[26][1] , \sa_snapshot[26].r.part0[1] );
tran (\sa_snapshot[26][1] , \sa_snapshot[26].f.lower[1] );
tran (\sa_snapshot[26][2] , \sa_snapshot[26].r.part0[2] );
tran (\sa_snapshot[26][2] , \sa_snapshot[26].f.lower[2] );
tran (\sa_snapshot[26][3] , \sa_snapshot[26].r.part0[3] );
tran (\sa_snapshot[26][3] , \sa_snapshot[26].f.lower[3] );
tran (\sa_snapshot[26][4] , \sa_snapshot[26].r.part0[4] );
tran (\sa_snapshot[26][4] , \sa_snapshot[26].f.lower[4] );
tran (\sa_snapshot[26][5] , \sa_snapshot[26].r.part0[5] );
tran (\sa_snapshot[26][5] , \sa_snapshot[26].f.lower[5] );
tran (\sa_snapshot[26][6] , \sa_snapshot[26].r.part0[6] );
tran (\sa_snapshot[26][6] , \sa_snapshot[26].f.lower[6] );
tran (\sa_snapshot[26][7] , \sa_snapshot[26].r.part0[7] );
tran (\sa_snapshot[26][7] , \sa_snapshot[26].f.lower[7] );
tran (\sa_snapshot[26][8] , \sa_snapshot[26].r.part0[8] );
tran (\sa_snapshot[26][8] , \sa_snapshot[26].f.lower[8] );
tran (\sa_snapshot[26][9] , \sa_snapshot[26].r.part0[9] );
tran (\sa_snapshot[26][9] , \sa_snapshot[26].f.lower[9] );
tran (\sa_snapshot[26][10] , \sa_snapshot[26].r.part0[10] );
tran (\sa_snapshot[26][10] , \sa_snapshot[26].f.lower[10] );
tran (\sa_snapshot[26][11] , \sa_snapshot[26].r.part0[11] );
tran (\sa_snapshot[26][11] , \sa_snapshot[26].f.lower[11] );
tran (\sa_snapshot[26][12] , \sa_snapshot[26].r.part0[12] );
tran (\sa_snapshot[26][12] , \sa_snapshot[26].f.lower[12] );
tran (\sa_snapshot[26][13] , \sa_snapshot[26].r.part0[13] );
tran (\sa_snapshot[26][13] , \sa_snapshot[26].f.lower[13] );
tran (\sa_snapshot[26][14] , \sa_snapshot[26].r.part0[14] );
tran (\sa_snapshot[26][14] , \sa_snapshot[26].f.lower[14] );
tran (\sa_snapshot[26][15] , \sa_snapshot[26].r.part0[15] );
tran (\sa_snapshot[26][15] , \sa_snapshot[26].f.lower[15] );
tran (\sa_snapshot[26][16] , \sa_snapshot[26].r.part0[16] );
tran (\sa_snapshot[26][16] , \sa_snapshot[26].f.lower[16] );
tran (\sa_snapshot[26][17] , \sa_snapshot[26].r.part0[17] );
tran (\sa_snapshot[26][17] , \sa_snapshot[26].f.lower[17] );
tran (\sa_snapshot[26][18] , \sa_snapshot[26].r.part0[18] );
tran (\sa_snapshot[26][18] , \sa_snapshot[26].f.lower[18] );
tran (\sa_snapshot[26][19] , \sa_snapshot[26].r.part0[19] );
tran (\sa_snapshot[26][19] , \sa_snapshot[26].f.lower[19] );
tran (\sa_snapshot[26][20] , \sa_snapshot[26].r.part0[20] );
tran (\sa_snapshot[26][20] , \sa_snapshot[26].f.lower[20] );
tran (\sa_snapshot[26][21] , \sa_snapshot[26].r.part0[21] );
tran (\sa_snapshot[26][21] , \sa_snapshot[26].f.lower[21] );
tran (\sa_snapshot[26][22] , \sa_snapshot[26].r.part0[22] );
tran (\sa_snapshot[26][22] , \sa_snapshot[26].f.lower[22] );
tran (\sa_snapshot[26][23] , \sa_snapshot[26].r.part0[23] );
tran (\sa_snapshot[26][23] , \sa_snapshot[26].f.lower[23] );
tran (\sa_snapshot[26][24] , \sa_snapshot[26].r.part0[24] );
tran (\sa_snapshot[26][24] , \sa_snapshot[26].f.lower[24] );
tran (\sa_snapshot[26][25] , \sa_snapshot[26].r.part0[25] );
tran (\sa_snapshot[26][25] , \sa_snapshot[26].f.lower[25] );
tran (\sa_snapshot[26][26] , \sa_snapshot[26].r.part0[26] );
tran (\sa_snapshot[26][26] , \sa_snapshot[26].f.lower[26] );
tran (\sa_snapshot[26][27] , \sa_snapshot[26].r.part0[27] );
tran (\sa_snapshot[26][27] , \sa_snapshot[26].f.lower[27] );
tran (\sa_snapshot[26][28] , \sa_snapshot[26].r.part0[28] );
tran (\sa_snapshot[26][28] , \sa_snapshot[26].f.lower[28] );
tran (\sa_snapshot[26][29] , \sa_snapshot[26].r.part0[29] );
tran (\sa_snapshot[26][29] , \sa_snapshot[26].f.lower[29] );
tran (\sa_snapshot[26][30] , \sa_snapshot[26].r.part0[30] );
tran (\sa_snapshot[26][30] , \sa_snapshot[26].f.lower[30] );
tran (\sa_snapshot[26][31] , \sa_snapshot[26].r.part0[31] );
tran (\sa_snapshot[26][31] , \sa_snapshot[26].f.lower[31] );
tran (\sa_snapshot[26][32] , \sa_snapshot[26].r.part1[0] );
tran (\sa_snapshot[26][32] , \sa_snapshot[26].f.upper[0] );
tran (\sa_snapshot[26][33] , \sa_snapshot[26].r.part1[1] );
tran (\sa_snapshot[26][33] , \sa_snapshot[26].f.upper[1] );
tran (\sa_snapshot[26][34] , \sa_snapshot[26].r.part1[2] );
tran (\sa_snapshot[26][34] , \sa_snapshot[26].f.upper[2] );
tran (\sa_snapshot[26][35] , \sa_snapshot[26].r.part1[3] );
tran (\sa_snapshot[26][35] , \sa_snapshot[26].f.upper[3] );
tran (\sa_snapshot[26][36] , \sa_snapshot[26].r.part1[4] );
tran (\sa_snapshot[26][36] , \sa_snapshot[26].f.upper[4] );
tran (\sa_snapshot[26][37] , \sa_snapshot[26].r.part1[5] );
tran (\sa_snapshot[26][37] , \sa_snapshot[26].f.upper[5] );
tran (\sa_snapshot[26][38] , \sa_snapshot[26].r.part1[6] );
tran (\sa_snapshot[26][38] , \sa_snapshot[26].f.upper[6] );
tran (\sa_snapshot[26][39] , \sa_snapshot[26].r.part1[7] );
tran (\sa_snapshot[26][39] , \sa_snapshot[26].f.upper[7] );
tran (\sa_snapshot[26][40] , \sa_snapshot[26].r.part1[8] );
tran (\sa_snapshot[26][40] , \sa_snapshot[26].f.upper[8] );
tran (\sa_snapshot[26][41] , \sa_snapshot[26].r.part1[9] );
tran (\sa_snapshot[26][41] , \sa_snapshot[26].f.upper[9] );
tran (\sa_snapshot[26][42] , \sa_snapshot[26].r.part1[10] );
tran (\sa_snapshot[26][42] , \sa_snapshot[26].f.upper[10] );
tran (\sa_snapshot[26][43] , \sa_snapshot[26].r.part1[11] );
tran (\sa_snapshot[26][43] , \sa_snapshot[26].f.upper[11] );
tran (\sa_snapshot[26][44] , \sa_snapshot[26].r.part1[12] );
tran (\sa_snapshot[26][44] , \sa_snapshot[26].f.upper[12] );
tran (\sa_snapshot[26][45] , \sa_snapshot[26].r.part1[13] );
tran (\sa_snapshot[26][45] , \sa_snapshot[26].f.upper[13] );
tran (\sa_snapshot[26][46] , \sa_snapshot[26].r.part1[14] );
tran (\sa_snapshot[26][46] , \sa_snapshot[26].f.upper[14] );
tran (\sa_snapshot[26][47] , \sa_snapshot[26].r.part1[15] );
tran (\sa_snapshot[26][47] , \sa_snapshot[26].f.upper[15] );
tran (\sa_snapshot[26][48] , \sa_snapshot[26].r.part1[16] );
tran (\sa_snapshot[26][48] , \sa_snapshot[26].f.upper[16] );
tran (\sa_snapshot[26][49] , \sa_snapshot[26].r.part1[17] );
tran (\sa_snapshot[26][49] , \sa_snapshot[26].f.upper[17] );
tran (\sa_snapshot[26][50] , \sa_snapshot[26].r.part1[18] );
tran (\sa_snapshot[26][50] , \sa_snapshot[26].f.unused[0] );
tran (\sa_snapshot[26][51] , \sa_snapshot[26].r.part1[19] );
tran (\sa_snapshot[26][51] , \sa_snapshot[26].f.unused[1] );
tran (\sa_snapshot[26][52] , \sa_snapshot[26].r.part1[20] );
tran (\sa_snapshot[26][52] , \sa_snapshot[26].f.unused[2] );
tran (\sa_snapshot[26][53] , \sa_snapshot[26].r.part1[21] );
tran (\sa_snapshot[26][53] , \sa_snapshot[26].f.unused[3] );
tran (\sa_snapshot[26][54] , \sa_snapshot[26].r.part1[22] );
tran (\sa_snapshot[26][54] , \sa_snapshot[26].f.unused[4] );
tran (\sa_snapshot[26][55] , \sa_snapshot[26].r.part1[23] );
tran (\sa_snapshot[26][55] , \sa_snapshot[26].f.unused[5] );
tran (\sa_snapshot[26][56] , \sa_snapshot[26].r.part1[24] );
tran (\sa_snapshot[26][56] , \sa_snapshot[26].f.unused[6] );
tran (\sa_snapshot[26][57] , \sa_snapshot[26].r.part1[25] );
tran (\sa_snapshot[26][57] , \sa_snapshot[26].f.unused[7] );
tran (\sa_snapshot[26][58] , \sa_snapshot[26].r.part1[26] );
tran (\sa_snapshot[26][58] , \sa_snapshot[26].f.unused[8] );
tran (\sa_snapshot[26][59] , \sa_snapshot[26].r.part1[27] );
tran (\sa_snapshot[26][59] , \sa_snapshot[26].f.unused[9] );
tran (\sa_snapshot[26][60] , \sa_snapshot[26].r.part1[28] );
tran (\sa_snapshot[26][60] , \sa_snapshot[26].f.unused[10] );
tran (\sa_snapshot[26][61] , \sa_snapshot[26].r.part1[29] );
tran (\sa_snapshot[26][61] , \sa_snapshot[26].f.unused[11] );
tran (\sa_snapshot[26][62] , \sa_snapshot[26].r.part1[30] );
tran (\sa_snapshot[26][62] , \sa_snapshot[26].f.unused[12] );
tran (\sa_snapshot[26][63] , \sa_snapshot[26].r.part1[31] );
tran (\sa_snapshot[26][63] , \sa_snapshot[26].f.unused[13] );
tran (\sa_snapshot[27][0] , \sa_snapshot[27].r.part0[0] );
tran (\sa_snapshot[27][0] , \sa_snapshot[27].f.lower[0] );
tran (\sa_snapshot[27][1] , \sa_snapshot[27].r.part0[1] );
tran (\sa_snapshot[27][1] , \sa_snapshot[27].f.lower[1] );
tran (\sa_snapshot[27][2] , \sa_snapshot[27].r.part0[2] );
tran (\sa_snapshot[27][2] , \sa_snapshot[27].f.lower[2] );
tran (\sa_snapshot[27][3] , \sa_snapshot[27].r.part0[3] );
tran (\sa_snapshot[27][3] , \sa_snapshot[27].f.lower[3] );
tran (\sa_snapshot[27][4] , \sa_snapshot[27].r.part0[4] );
tran (\sa_snapshot[27][4] , \sa_snapshot[27].f.lower[4] );
tran (\sa_snapshot[27][5] , \sa_snapshot[27].r.part0[5] );
tran (\sa_snapshot[27][5] , \sa_snapshot[27].f.lower[5] );
tran (\sa_snapshot[27][6] , \sa_snapshot[27].r.part0[6] );
tran (\sa_snapshot[27][6] , \sa_snapshot[27].f.lower[6] );
tran (\sa_snapshot[27][7] , \sa_snapshot[27].r.part0[7] );
tran (\sa_snapshot[27][7] , \sa_snapshot[27].f.lower[7] );
tran (\sa_snapshot[27][8] , \sa_snapshot[27].r.part0[8] );
tran (\sa_snapshot[27][8] , \sa_snapshot[27].f.lower[8] );
tran (\sa_snapshot[27][9] , \sa_snapshot[27].r.part0[9] );
tran (\sa_snapshot[27][9] , \sa_snapshot[27].f.lower[9] );
tran (\sa_snapshot[27][10] , \sa_snapshot[27].r.part0[10] );
tran (\sa_snapshot[27][10] , \sa_snapshot[27].f.lower[10] );
tran (\sa_snapshot[27][11] , \sa_snapshot[27].r.part0[11] );
tran (\sa_snapshot[27][11] , \sa_snapshot[27].f.lower[11] );
tran (\sa_snapshot[27][12] , \sa_snapshot[27].r.part0[12] );
tran (\sa_snapshot[27][12] , \sa_snapshot[27].f.lower[12] );
tran (\sa_snapshot[27][13] , \sa_snapshot[27].r.part0[13] );
tran (\sa_snapshot[27][13] , \sa_snapshot[27].f.lower[13] );
tran (\sa_snapshot[27][14] , \sa_snapshot[27].r.part0[14] );
tran (\sa_snapshot[27][14] , \sa_snapshot[27].f.lower[14] );
tran (\sa_snapshot[27][15] , \sa_snapshot[27].r.part0[15] );
tran (\sa_snapshot[27][15] , \sa_snapshot[27].f.lower[15] );
tran (\sa_snapshot[27][16] , \sa_snapshot[27].r.part0[16] );
tran (\sa_snapshot[27][16] , \sa_snapshot[27].f.lower[16] );
tran (\sa_snapshot[27][17] , \sa_snapshot[27].r.part0[17] );
tran (\sa_snapshot[27][17] , \sa_snapshot[27].f.lower[17] );
tran (\sa_snapshot[27][18] , \sa_snapshot[27].r.part0[18] );
tran (\sa_snapshot[27][18] , \sa_snapshot[27].f.lower[18] );
tran (\sa_snapshot[27][19] , \sa_snapshot[27].r.part0[19] );
tran (\sa_snapshot[27][19] , \sa_snapshot[27].f.lower[19] );
tran (\sa_snapshot[27][20] , \sa_snapshot[27].r.part0[20] );
tran (\sa_snapshot[27][20] , \sa_snapshot[27].f.lower[20] );
tran (\sa_snapshot[27][21] , \sa_snapshot[27].r.part0[21] );
tran (\sa_snapshot[27][21] , \sa_snapshot[27].f.lower[21] );
tran (\sa_snapshot[27][22] , \sa_snapshot[27].r.part0[22] );
tran (\sa_snapshot[27][22] , \sa_snapshot[27].f.lower[22] );
tran (\sa_snapshot[27][23] , \sa_snapshot[27].r.part0[23] );
tran (\sa_snapshot[27][23] , \sa_snapshot[27].f.lower[23] );
tran (\sa_snapshot[27][24] , \sa_snapshot[27].r.part0[24] );
tran (\sa_snapshot[27][24] , \sa_snapshot[27].f.lower[24] );
tran (\sa_snapshot[27][25] , \sa_snapshot[27].r.part0[25] );
tran (\sa_snapshot[27][25] , \sa_snapshot[27].f.lower[25] );
tran (\sa_snapshot[27][26] , \sa_snapshot[27].r.part0[26] );
tran (\sa_snapshot[27][26] , \sa_snapshot[27].f.lower[26] );
tran (\sa_snapshot[27][27] , \sa_snapshot[27].r.part0[27] );
tran (\sa_snapshot[27][27] , \sa_snapshot[27].f.lower[27] );
tran (\sa_snapshot[27][28] , \sa_snapshot[27].r.part0[28] );
tran (\sa_snapshot[27][28] , \sa_snapshot[27].f.lower[28] );
tran (\sa_snapshot[27][29] , \sa_snapshot[27].r.part0[29] );
tran (\sa_snapshot[27][29] , \sa_snapshot[27].f.lower[29] );
tran (\sa_snapshot[27][30] , \sa_snapshot[27].r.part0[30] );
tran (\sa_snapshot[27][30] , \sa_snapshot[27].f.lower[30] );
tran (\sa_snapshot[27][31] , \sa_snapshot[27].r.part0[31] );
tran (\sa_snapshot[27][31] , \sa_snapshot[27].f.lower[31] );
tran (\sa_snapshot[27][32] , \sa_snapshot[27].r.part1[0] );
tran (\sa_snapshot[27][32] , \sa_snapshot[27].f.upper[0] );
tran (\sa_snapshot[27][33] , \sa_snapshot[27].r.part1[1] );
tran (\sa_snapshot[27][33] , \sa_snapshot[27].f.upper[1] );
tran (\sa_snapshot[27][34] , \sa_snapshot[27].r.part1[2] );
tran (\sa_snapshot[27][34] , \sa_snapshot[27].f.upper[2] );
tran (\sa_snapshot[27][35] , \sa_snapshot[27].r.part1[3] );
tran (\sa_snapshot[27][35] , \sa_snapshot[27].f.upper[3] );
tran (\sa_snapshot[27][36] , \sa_snapshot[27].r.part1[4] );
tran (\sa_snapshot[27][36] , \sa_snapshot[27].f.upper[4] );
tran (\sa_snapshot[27][37] , \sa_snapshot[27].r.part1[5] );
tran (\sa_snapshot[27][37] , \sa_snapshot[27].f.upper[5] );
tran (\sa_snapshot[27][38] , \sa_snapshot[27].r.part1[6] );
tran (\sa_snapshot[27][38] , \sa_snapshot[27].f.upper[6] );
tran (\sa_snapshot[27][39] , \sa_snapshot[27].r.part1[7] );
tran (\sa_snapshot[27][39] , \sa_snapshot[27].f.upper[7] );
tran (\sa_snapshot[27][40] , \sa_snapshot[27].r.part1[8] );
tran (\sa_snapshot[27][40] , \sa_snapshot[27].f.upper[8] );
tran (\sa_snapshot[27][41] , \sa_snapshot[27].r.part1[9] );
tran (\sa_snapshot[27][41] , \sa_snapshot[27].f.upper[9] );
tran (\sa_snapshot[27][42] , \sa_snapshot[27].r.part1[10] );
tran (\sa_snapshot[27][42] , \sa_snapshot[27].f.upper[10] );
tran (\sa_snapshot[27][43] , \sa_snapshot[27].r.part1[11] );
tran (\sa_snapshot[27][43] , \sa_snapshot[27].f.upper[11] );
tran (\sa_snapshot[27][44] , \sa_snapshot[27].r.part1[12] );
tran (\sa_snapshot[27][44] , \sa_snapshot[27].f.upper[12] );
tran (\sa_snapshot[27][45] , \sa_snapshot[27].r.part1[13] );
tran (\sa_snapshot[27][45] , \sa_snapshot[27].f.upper[13] );
tran (\sa_snapshot[27][46] , \sa_snapshot[27].r.part1[14] );
tran (\sa_snapshot[27][46] , \sa_snapshot[27].f.upper[14] );
tran (\sa_snapshot[27][47] , \sa_snapshot[27].r.part1[15] );
tran (\sa_snapshot[27][47] , \sa_snapshot[27].f.upper[15] );
tran (\sa_snapshot[27][48] , \sa_snapshot[27].r.part1[16] );
tran (\sa_snapshot[27][48] , \sa_snapshot[27].f.upper[16] );
tran (\sa_snapshot[27][49] , \sa_snapshot[27].r.part1[17] );
tran (\sa_snapshot[27][49] , \sa_snapshot[27].f.upper[17] );
tran (\sa_snapshot[27][50] , \sa_snapshot[27].r.part1[18] );
tran (\sa_snapshot[27][50] , \sa_snapshot[27].f.unused[0] );
tran (\sa_snapshot[27][51] , \sa_snapshot[27].r.part1[19] );
tran (\sa_snapshot[27][51] , \sa_snapshot[27].f.unused[1] );
tran (\sa_snapshot[27][52] , \sa_snapshot[27].r.part1[20] );
tran (\sa_snapshot[27][52] , \sa_snapshot[27].f.unused[2] );
tran (\sa_snapshot[27][53] , \sa_snapshot[27].r.part1[21] );
tran (\sa_snapshot[27][53] , \sa_snapshot[27].f.unused[3] );
tran (\sa_snapshot[27][54] , \sa_snapshot[27].r.part1[22] );
tran (\sa_snapshot[27][54] , \sa_snapshot[27].f.unused[4] );
tran (\sa_snapshot[27][55] , \sa_snapshot[27].r.part1[23] );
tran (\sa_snapshot[27][55] , \sa_snapshot[27].f.unused[5] );
tran (\sa_snapshot[27][56] , \sa_snapshot[27].r.part1[24] );
tran (\sa_snapshot[27][56] , \sa_snapshot[27].f.unused[6] );
tran (\sa_snapshot[27][57] , \sa_snapshot[27].r.part1[25] );
tran (\sa_snapshot[27][57] , \sa_snapshot[27].f.unused[7] );
tran (\sa_snapshot[27][58] , \sa_snapshot[27].r.part1[26] );
tran (\sa_snapshot[27][58] , \sa_snapshot[27].f.unused[8] );
tran (\sa_snapshot[27][59] , \sa_snapshot[27].r.part1[27] );
tran (\sa_snapshot[27][59] , \sa_snapshot[27].f.unused[9] );
tran (\sa_snapshot[27][60] , \sa_snapshot[27].r.part1[28] );
tran (\sa_snapshot[27][60] , \sa_snapshot[27].f.unused[10] );
tran (\sa_snapshot[27][61] , \sa_snapshot[27].r.part1[29] );
tran (\sa_snapshot[27][61] , \sa_snapshot[27].f.unused[11] );
tran (\sa_snapshot[27][62] , \sa_snapshot[27].r.part1[30] );
tran (\sa_snapshot[27][62] , \sa_snapshot[27].f.unused[12] );
tran (\sa_snapshot[27][63] , \sa_snapshot[27].r.part1[31] );
tran (\sa_snapshot[27][63] , \sa_snapshot[27].f.unused[13] );
tran (\sa_snapshot[28][0] , \sa_snapshot[28].r.part0[0] );
tran (\sa_snapshot[28][0] , \sa_snapshot[28].f.lower[0] );
tran (\sa_snapshot[28][1] , \sa_snapshot[28].r.part0[1] );
tran (\sa_snapshot[28][1] , \sa_snapshot[28].f.lower[1] );
tran (\sa_snapshot[28][2] , \sa_snapshot[28].r.part0[2] );
tran (\sa_snapshot[28][2] , \sa_snapshot[28].f.lower[2] );
tran (\sa_snapshot[28][3] , \sa_snapshot[28].r.part0[3] );
tran (\sa_snapshot[28][3] , \sa_snapshot[28].f.lower[3] );
tran (\sa_snapshot[28][4] , \sa_snapshot[28].r.part0[4] );
tran (\sa_snapshot[28][4] , \sa_snapshot[28].f.lower[4] );
tran (\sa_snapshot[28][5] , \sa_snapshot[28].r.part0[5] );
tran (\sa_snapshot[28][5] , \sa_snapshot[28].f.lower[5] );
tran (\sa_snapshot[28][6] , \sa_snapshot[28].r.part0[6] );
tran (\sa_snapshot[28][6] , \sa_snapshot[28].f.lower[6] );
tran (\sa_snapshot[28][7] , \sa_snapshot[28].r.part0[7] );
tran (\sa_snapshot[28][7] , \sa_snapshot[28].f.lower[7] );
tran (\sa_snapshot[28][8] , \sa_snapshot[28].r.part0[8] );
tran (\sa_snapshot[28][8] , \sa_snapshot[28].f.lower[8] );
tran (\sa_snapshot[28][9] , \sa_snapshot[28].r.part0[9] );
tran (\sa_snapshot[28][9] , \sa_snapshot[28].f.lower[9] );
tran (\sa_snapshot[28][10] , \sa_snapshot[28].r.part0[10] );
tran (\sa_snapshot[28][10] , \sa_snapshot[28].f.lower[10] );
tran (\sa_snapshot[28][11] , \sa_snapshot[28].r.part0[11] );
tran (\sa_snapshot[28][11] , \sa_snapshot[28].f.lower[11] );
tran (\sa_snapshot[28][12] , \sa_snapshot[28].r.part0[12] );
tran (\sa_snapshot[28][12] , \sa_snapshot[28].f.lower[12] );
tran (\sa_snapshot[28][13] , \sa_snapshot[28].r.part0[13] );
tran (\sa_snapshot[28][13] , \sa_snapshot[28].f.lower[13] );
tran (\sa_snapshot[28][14] , \sa_snapshot[28].r.part0[14] );
tran (\sa_snapshot[28][14] , \sa_snapshot[28].f.lower[14] );
tran (\sa_snapshot[28][15] , \sa_snapshot[28].r.part0[15] );
tran (\sa_snapshot[28][15] , \sa_snapshot[28].f.lower[15] );
tran (\sa_snapshot[28][16] , \sa_snapshot[28].r.part0[16] );
tran (\sa_snapshot[28][16] , \sa_snapshot[28].f.lower[16] );
tran (\sa_snapshot[28][17] , \sa_snapshot[28].r.part0[17] );
tran (\sa_snapshot[28][17] , \sa_snapshot[28].f.lower[17] );
tran (\sa_snapshot[28][18] , \sa_snapshot[28].r.part0[18] );
tran (\sa_snapshot[28][18] , \sa_snapshot[28].f.lower[18] );
tran (\sa_snapshot[28][19] , \sa_snapshot[28].r.part0[19] );
tran (\sa_snapshot[28][19] , \sa_snapshot[28].f.lower[19] );
tran (\sa_snapshot[28][20] , \sa_snapshot[28].r.part0[20] );
tran (\sa_snapshot[28][20] , \sa_snapshot[28].f.lower[20] );
tran (\sa_snapshot[28][21] , \sa_snapshot[28].r.part0[21] );
tran (\sa_snapshot[28][21] , \sa_snapshot[28].f.lower[21] );
tran (\sa_snapshot[28][22] , \sa_snapshot[28].r.part0[22] );
tran (\sa_snapshot[28][22] , \sa_snapshot[28].f.lower[22] );
tran (\sa_snapshot[28][23] , \sa_snapshot[28].r.part0[23] );
tran (\sa_snapshot[28][23] , \sa_snapshot[28].f.lower[23] );
tran (\sa_snapshot[28][24] , \sa_snapshot[28].r.part0[24] );
tran (\sa_snapshot[28][24] , \sa_snapshot[28].f.lower[24] );
tran (\sa_snapshot[28][25] , \sa_snapshot[28].r.part0[25] );
tran (\sa_snapshot[28][25] , \sa_snapshot[28].f.lower[25] );
tran (\sa_snapshot[28][26] , \sa_snapshot[28].r.part0[26] );
tran (\sa_snapshot[28][26] , \sa_snapshot[28].f.lower[26] );
tran (\sa_snapshot[28][27] , \sa_snapshot[28].r.part0[27] );
tran (\sa_snapshot[28][27] , \sa_snapshot[28].f.lower[27] );
tran (\sa_snapshot[28][28] , \sa_snapshot[28].r.part0[28] );
tran (\sa_snapshot[28][28] , \sa_snapshot[28].f.lower[28] );
tran (\sa_snapshot[28][29] , \sa_snapshot[28].r.part0[29] );
tran (\sa_snapshot[28][29] , \sa_snapshot[28].f.lower[29] );
tran (\sa_snapshot[28][30] , \sa_snapshot[28].r.part0[30] );
tran (\sa_snapshot[28][30] , \sa_snapshot[28].f.lower[30] );
tran (\sa_snapshot[28][31] , \sa_snapshot[28].r.part0[31] );
tran (\sa_snapshot[28][31] , \sa_snapshot[28].f.lower[31] );
tran (\sa_snapshot[28][32] , \sa_snapshot[28].r.part1[0] );
tran (\sa_snapshot[28][32] , \sa_snapshot[28].f.upper[0] );
tran (\sa_snapshot[28][33] , \sa_snapshot[28].r.part1[1] );
tran (\sa_snapshot[28][33] , \sa_snapshot[28].f.upper[1] );
tran (\sa_snapshot[28][34] , \sa_snapshot[28].r.part1[2] );
tran (\sa_snapshot[28][34] , \sa_snapshot[28].f.upper[2] );
tran (\sa_snapshot[28][35] , \sa_snapshot[28].r.part1[3] );
tran (\sa_snapshot[28][35] , \sa_snapshot[28].f.upper[3] );
tran (\sa_snapshot[28][36] , \sa_snapshot[28].r.part1[4] );
tran (\sa_snapshot[28][36] , \sa_snapshot[28].f.upper[4] );
tran (\sa_snapshot[28][37] , \sa_snapshot[28].r.part1[5] );
tran (\sa_snapshot[28][37] , \sa_snapshot[28].f.upper[5] );
tran (\sa_snapshot[28][38] , \sa_snapshot[28].r.part1[6] );
tran (\sa_snapshot[28][38] , \sa_snapshot[28].f.upper[6] );
tran (\sa_snapshot[28][39] , \sa_snapshot[28].r.part1[7] );
tran (\sa_snapshot[28][39] , \sa_snapshot[28].f.upper[7] );
tran (\sa_snapshot[28][40] , \sa_snapshot[28].r.part1[8] );
tran (\sa_snapshot[28][40] , \sa_snapshot[28].f.upper[8] );
tran (\sa_snapshot[28][41] , \sa_snapshot[28].r.part1[9] );
tran (\sa_snapshot[28][41] , \sa_snapshot[28].f.upper[9] );
tran (\sa_snapshot[28][42] , \sa_snapshot[28].r.part1[10] );
tran (\sa_snapshot[28][42] , \sa_snapshot[28].f.upper[10] );
tran (\sa_snapshot[28][43] , \sa_snapshot[28].r.part1[11] );
tran (\sa_snapshot[28][43] , \sa_snapshot[28].f.upper[11] );
tran (\sa_snapshot[28][44] , \sa_snapshot[28].r.part1[12] );
tran (\sa_snapshot[28][44] , \sa_snapshot[28].f.upper[12] );
tran (\sa_snapshot[28][45] , \sa_snapshot[28].r.part1[13] );
tran (\sa_snapshot[28][45] , \sa_snapshot[28].f.upper[13] );
tran (\sa_snapshot[28][46] , \sa_snapshot[28].r.part1[14] );
tran (\sa_snapshot[28][46] , \sa_snapshot[28].f.upper[14] );
tran (\sa_snapshot[28][47] , \sa_snapshot[28].r.part1[15] );
tran (\sa_snapshot[28][47] , \sa_snapshot[28].f.upper[15] );
tran (\sa_snapshot[28][48] , \sa_snapshot[28].r.part1[16] );
tran (\sa_snapshot[28][48] , \sa_snapshot[28].f.upper[16] );
tran (\sa_snapshot[28][49] , \sa_snapshot[28].r.part1[17] );
tran (\sa_snapshot[28][49] , \sa_snapshot[28].f.upper[17] );
tran (\sa_snapshot[28][50] , \sa_snapshot[28].r.part1[18] );
tran (\sa_snapshot[28][50] , \sa_snapshot[28].f.unused[0] );
tran (\sa_snapshot[28][51] , \sa_snapshot[28].r.part1[19] );
tran (\sa_snapshot[28][51] , \sa_snapshot[28].f.unused[1] );
tran (\sa_snapshot[28][52] , \sa_snapshot[28].r.part1[20] );
tran (\sa_snapshot[28][52] , \sa_snapshot[28].f.unused[2] );
tran (\sa_snapshot[28][53] , \sa_snapshot[28].r.part1[21] );
tran (\sa_snapshot[28][53] , \sa_snapshot[28].f.unused[3] );
tran (\sa_snapshot[28][54] , \sa_snapshot[28].r.part1[22] );
tran (\sa_snapshot[28][54] , \sa_snapshot[28].f.unused[4] );
tran (\sa_snapshot[28][55] , \sa_snapshot[28].r.part1[23] );
tran (\sa_snapshot[28][55] , \sa_snapshot[28].f.unused[5] );
tran (\sa_snapshot[28][56] , \sa_snapshot[28].r.part1[24] );
tran (\sa_snapshot[28][56] , \sa_snapshot[28].f.unused[6] );
tran (\sa_snapshot[28][57] , \sa_snapshot[28].r.part1[25] );
tran (\sa_snapshot[28][57] , \sa_snapshot[28].f.unused[7] );
tran (\sa_snapshot[28][58] , \sa_snapshot[28].r.part1[26] );
tran (\sa_snapshot[28][58] , \sa_snapshot[28].f.unused[8] );
tran (\sa_snapshot[28][59] , \sa_snapshot[28].r.part1[27] );
tran (\sa_snapshot[28][59] , \sa_snapshot[28].f.unused[9] );
tran (\sa_snapshot[28][60] , \sa_snapshot[28].r.part1[28] );
tran (\sa_snapshot[28][60] , \sa_snapshot[28].f.unused[10] );
tran (\sa_snapshot[28][61] , \sa_snapshot[28].r.part1[29] );
tran (\sa_snapshot[28][61] , \sa_snapshot[28].f.unused[11] );
tran (\sa_snapshot[28][62] , \sa_snapshot[28].r.part1[30] );
tran (\sa_snapshot[28][62] , \sa_snapshot[28].f.unused[12] );
tran (\sa_snapshot[28][63] , \sa_snapshot[28].r.part1[31] );
tran (\sa_snapshot[28][63] , \sa_snapshot[28].f.unused[13] );
tran (\sa_snapshot[29][0] , \sa_snapshot[29].r.part0[0] );
tran (\sa_snapshot[29][0] , \sa_snapshot[29].f.lower[0] );
tran (\sa_snapshot[29][1] , \sa_snapshot[29].r.part0[1] );
tran (\sa_snapshot[29][1] , \sa_snapshot[29].f.lower[1] );
tran (\sa_snapshot[29][2] , \sa_snapshot[29].r.part0[2] );
tran (\sa_snapshot[29][2] , \sa_snapshot[29].f.lower[2] );
tran (\sa_snapshot[29][3] , \sa_snapshot[29].r.part0[3] );
tran (\sa_snapshot[29][3] , \sa_snapshot[29].f.lower[3] );
tran (\sa_snapshot[29][4] , \sa_snapshot[29].r.part0[4] );
tran (\sa_snapshot[29][4] , \sa_snapshot[29].f.lower[4] );
tran (\sa_snapshot[29][5] , \sa_snapshot[29].r.part0[5] );
tran (\sa_snapshot[29][5] , \sa_snapshot[29].f.lower[5] );
tran (\sa_snapshot[29][6] , \sa_snapshot[29].r.part0[6] );
tran (\sa_snapshot[29][6] , \sa_snapshot[29].f.lower[6] );
tran (\sa_snapshot[29][7] , \sa_snapshot[29].r.part0[7] );
tran (\sa_snapshot[29][7] , \sa_snapshot[29].f.lower[7] );
tran (\sa_snapshot[29][8] , \sa_snapshot[29].r.part0[8] );
tran (\sa_snapshot[29][8] , \sa_snapshot[29].f.lower[8] );
tran (\sa_snapshot[29][9] , \sa_snapshot[29].r.part0[9] );
tran (\sa_snapshot[29][9] , \sa_snapshot[29].f.lower[9] );
tran (\sa_snapshot[29][10] , \sa_snapshot[29].r.part0[10] );
tran (\sa_snapshot[29][10] , \sa_snapshot[29].f.lower[10] );
tran (\sa_snapshot[29][11] , \sa_snapshot[29].r.part0[11] );
tran (\sa_snapshot[29][11] , \sa_snapshot[29].f.lower[11] );
tran (\sa_snapshot[29][12] , \sa_snapshot[29].r.part0[12] );
tran (\sa_snapshot[29][12] , \sa_snapshot[29].f.lower[12] );
tran (\sa_snapshot[29][13] , \sa_snapshot[29].r.part0[13] );
tran (\sa_snapshot[29][13] , \sa_snapshot[29].f.lower[13] );
tran (\sa_snapshot[29][14] , \sa_snapshot[29].r.part0[14] );
tran (\sa_snapshot[29][14] , \sa_snapshot[29].f.lower[14] );
tran (\sa_snapshot[29][15] , \sa_snapshot[29].r.part0[15] );
tran (\sa_snapshot[29][15] , \sa_snapshot[29].f.lower[15] );
tran (\sa_snapshot[29][16] , \sa_snapshot[29].r.part0[16] );
tran (\sa_snapshot[29][16] , \sa_snapshot[29].f.lower[16] );
tran (\sa_snapshot[29][17] , \sa_snapshot[29].r.part0[17] );
tran (\sa_snapshot[29][17] , \sa_snapshot[29].f.lower[17] );
tran (\sa_snapshot[29][18] , \sa_snapshot[29].r.part0[18] );
tran (\sa_snapshot[29][18] , \sa_snapshot[29].f.lower[18] );
tran (\sa_snapshot[29][19] , \sa_snapshot[29].r.part0[19] );
tran (\sa_snapshot[29][19] , \sa_snapshot[29].f.lower[19] );
tran (\sa_snapshot[29][20] , \sa_snapshot[29].r.part0[20] );
tran (\sa_snapshot[29][20] , \sa_snapshot[29].f.lower[20] );
tran (\sa_snapshot[29][21] , \sa_snapshot[29].r.part0[21] );
tran (\sa_snapshot[29][21] , \sa_snapshot[29].f.lower[21] );
tran (\sa_snapshot[29][22] , \sa_snapshot[29].r.part0[22] );
tran (\sa_snapshot[29][22] , \sa_snapshot[29].f.lower[22] );
tran (\sa_snapshot[29][23] , \sa_snapshot[29].r.part0[23] );
tran (\sa_snapshot[29][23] , \sa_snapshot[29].f.lower[23] );
tran (\sa_snapshot[29][24] , \sa_snapshot[29].r.part0[24] );
tran (\sa_snapshot[29][24] , \sa_snapshot[29].f.lower[24] );
tran (\sa_snapshot[29][25] , \sa_snapshot[29].r.part0[25] );
tran (\sa_snapshot[29][25] , \sa_snapshot[29].f.lower[25] );
tran (\sa_snapshot[29][26] , \sa_snapshot[29].r.part0[26] );
tran (\sa_snapshot[29][26] , \sa_snapshot[29].f.lower[26] );
tran (\sa_snapshot[29][27] , \sa_snapshot[29].r.part0[27] );
tran (\sa_snapshot[29][27] , \sa_snapshot[29].f.lower[27] );
tran (\sa_snapshot[29][28] , \sa_snapshot[29].r.part0[28] );
tran (\sa_snapshot[29][28] , \sa_snapshot[29].f.lower[28] );
tran (\sa_snapshot[29][29] , \sa_snapshot[29].r.part0[29] );
tran (\sa_snapshot[29][29] , \sa_snapshot[29].f.lower[29] );
tran (\sa_snapshot[29][30] , \sa_snapshot[29].r.part0[30] );
tran (\sa_snapshot[29][30] , \sa_snapshot[29].f.lower[30] );
tran (\sa_snapshot[29][31] , \sa_snapshot[29].r.part0[31] );
tran (\sa_snapshot[29][31] , \sa_snapshot[29].f.lower[31] );
tran (\sa_snapshot[29][32] , \sa_snapshot[29].r.part1[0] );
tran (\sa_snapshot[29][32] , \sa_snapshot[29].f.upper[0] );
tran (\sa_snapshot[29][33] , \sa_snapshot[29].r.part1[1] );
tran (\sa_snapshot[29][33] , \sa_snapshot[29].f.upper[1] );
tran (\sa_snapshot[29][34] , \sa_snapshot[29].r.part1[2] );
tran (\sa_snapshot[29][34] , \sa_snapshot[29].f.upper[2] );
tran (\sa_snapshot[29][35] , \sa_snapshot[29].r.part1[3] );
tran (\sa_snapshot[29][35] , \sa_snapshot[29].f.upper[3] );
tran (\sa_snapshot[29][36] , \sa_snapshot[29].r.part1[4] );
tran (\sa_snapshot[29][36] , \sa_snapshot[29].f.upper[4] );
tran (\sa_snapshot[29][37] , \sa_snapshot[29].r.part1[5] );
tran (\sa_snapshot[29][37] , \sa_snapshot[29].f.upper[5] );
tran (\sa_snapshot[29][38] , \sa_snapshot[29].r.part1[6] );
tran (\sa_snapshot[29][38] , \sa_snapshot[29].f.upper[6] );
tran (\sa_snapshot[29][39] , \sa_snapshot[29].r.part1[7] );
tran (\sa_snapshot[29][39] , \sa_snapshot[29].f.upper[7] );
tran (\sa_snapshot[29][40] , \sa_snapshot[29].r.part1[8] );
tran (\sa_snapshot[29][40] , \sa_snapshot[29].f.upper[8] );
tran (\sa_snapshot[29][41] , \sa_snapshot[29].r.part1[9] );
tran (\sa_snapshot[29][41] , \sa_snapshot[29].f.upper[9] );
tran (\sa_snapshot[29][42] , \sa_snapshot[29].r.part1[10] );
tran (\sa_snapshot[29][42] , \sa_snapshot[29].f.upper[10] );
tran (\sa_snapshot[29][43] , \sa_snapshot[29].r.part1[11] );
tran (\sa_snapshot[29][43] , \sa_snapshot[29].f.upper[11] );
tran (\sa_snapshot[29][44] , \sa_snapshot[29].r.part1[12] );
tran (\sa_snapshot[29][44] , \sa_snapshot[29].f.upper[12] );
tran (\sa_snapshot[29][45] , \sa_snapshot[29].r.part1[13] );
tran (\sa_snapshot[29][45] , \sa_snapshot[29].f.upper[13] );
tran (\sa_snapshot[29][46] , \sa_snapshot[29].r.part1[14] );
tran (\sa_snapshot[29][46] , \sa_snapshot[29].f.upper[14] );
tran (\sa_snapshot[29][47] , \sa_snapshot[29].r.part1[15] );
tran (\sa_snapshot[29][47] , \sa_snapshot[29].f.upper[15] );
tran (\sa_snapshot[29][48] , \sa_snapshot[29].r.part1[16] );
tran (\sa_snapshot[29][48] , \sa_snapshot[29].f.upper[16] );
tran (\sa_snapshot[29][49] , \sa_snapshot[29].r.part1[17] );
tran (\sa_snapshot[29][49] , \sa_snapshot[29].f.upper[17] );
tran (\sa_snapshot[29][50] , \sa_snapshot[29].r.part1[18] );
tran (\sa_snapshot[29][50] , \sa_snapshot[29].f.unused[0] );
tran (\sa_snapshot[29][51] , \sa_snapshot[29].r.part1[19] );
tran (\sa_snapshot[29][51] , \sa_snapshot[29].f.unused[1] );
tran (\sa_snapshot[29][52] , \sa_snapshot[29].r.part1[20] );
tran (\sa_snapshot[29][52] , \sa_snapshot[29].f.unused[2] );
tran (\sa_snapshot[29][53] , \sa_snapshot[29].r.part1[21] );
tran (\sa_snapshot[29][53] , \sa_snapshot[29].f.unused[3] );
tran (\sa_snapshot[29][54] , \sa_snapshot[29].r.part1[22] );
tran (\sa_snapshot[29][54] , \sa_snapshot[29].f.unused[4] );
tran (\sa_snapshot[29][55] , \sa_snapshot[29].r.part1[23] );
tran (\sa_snapshot[29][55] , \sa_snapshot[29].f.unused[5] );
tran (\sa_snapshot[29][56] , \sa_snapshot[29].r.part1[24] );
tran (\sa_snapshot[29][56] , \sa_snapshot[29].f.unused[6] );
tran (\sa_snapshot[29][57] , \sa_snapshot[29].r.part1[25] );
tran (\sa_snapshot[29][57] , \sa_snapshot[29].f.unused[7] );
tran (\sa_snapshot[29][58] , \sa_snapshot[29].r.part1[26] );
tran (\sa_snapshot[29][58] , \sa_snapshot[29].f.unused[8] );
tran (\sa_snapshot[29][59] , \sa_snapshot[29].r.part1[27] );
tran (\sa_snapshot[29][59] , \sa_snapshot[29].f.unused[9] );
tran (\sa_snapshot[29][60] , \sa_snapshot[29].r.part1[28] );
tran (\sa_snapshot[29][60] , \sa_snapshot[29].f.unused[10] );
tran (\sa_snapshot[29][61] , \sa_snapshot[29].r.part1[29] );
tran (\sa_snapshot[29][61] , \sa_snapshot[29].f.unused[11] );
tran (\sa_snapshot[29][62] , \sa_snapshot[29].r.part1[30] );
tran (\sa_snapshot[29][62] , \sa_snapshot[29].f.unused[12] );
tran (\sa_snapshot[29][63] , \sa_snapshot[29].r.part1[31] );
tran (\sa_snapshot[29][63] , \sa_snapshot[29].f.unused[13] );
tran (\sa_snapshot[30][0] , \sa_snapshot[30].r.part0[0] );
tran (\sa_snapshot[30][0] , \sa_snapshot[30].f.lower[0] );
tran (\sa_snapshot[30][1] , \sa_snapshot[30].r.part0[1] );
tran (\sa_snapshot[30][1] , \sa_snapshot[30].f.lower[1] );
tran (\sa_snapshot[30][2] , \sa_snapshot[30].r.part0[2] );
tran (\sa_snapshot[30][2] , \sa_snapshot[30].f.lower[2] );
tran (\sa_snapshot[30][3] , \sa_snapshot[30].r.part0[3] );
tran (\sa_snapshot[30][3] , \sa_snapshot[30].f.lower[3] );
tran (\sa_snapshot[30][4] , \sa_snapshot[30].r.part0[4] );
tran (\sa_snapshot[30][4] , \sa_snapshot[30].f.lower[4] );
tran (\sa_snapshot[30][5] , \sa_snapshot[30].r.part0[5] );
tran (\sa_snapshot[30][5] , \sa_snapshot[30].f.lower[5] );
tran (\sa_snapshot[30][6] , \sa_snapshot[30].r.part0[6] );
tran (\sa_snapshot[30][6] , \sa_snapshot[30].f.lower[6] );
tran (\sa_snapshot[30][7] , \sa_snapshot[30].r.part0[7] );
tran (\sa_snapshot[30][7] , \sa_snapshot[30].f.lower[7] );
tran (\sa_snapshot[30][8] , \sa_snapshot[30].r.part0[8] );
tran (\sa_snapshot[30][8] , \sa_snapshot[30].f.lower[8] );
tran (\sa_snapshot[30][9] , \sa_snapshot[30].r.part0[9] );
tran (\sa_snapshot[30][9] , \sa_snapshot[30].f.lower[9] );
tran (\sa_snapshot[30][10] , \sa_snapshot[30].r.part0[10] );
tran (\sa_snapshot[30][10] , \sa_snapshot[30].f.lower[10] );
tran (\sa_snapshot[30][11] , \sa_snapshot[30].r.part0[11] );
tran (\sa_snapshot[30][11] , \sa_snapshot[30].f.lower[11] );
tran (\sa_snapshot[30][12] , \sa_snapshot[30].r.part0[12] );
tran (\sa_snapshot[30][12] , \sa_snapshot[30].f.lower[12] );
tran (\sa_snapshot[30][13] , \sa_snapshot[30].r.part0[13] );
tran (\sa_snapshot[30][13] , \sa_snapshot[30].f.lower[13] );
tran (\sa_snapshot[30][14] , \sa_snapshot[30].r.part0[14] );
tran (\sa_snapshot[30][14] , \sa_snapshot[30].f.lower[14] );
tran (\sa_snapshot[30][15] , \sa_snapshot[30].r.part0[15] );
tran (\sa_snapshot[30][15] , \sa_snapshot[30].f.lower[15] );
tran (\sa_snapshot[30][16] , \sa_snapshot[30].r.part0[16] );
tran (\sa_snapshot[30][16] , \sa_snapshot[30].f.lower[16] );
tran (\sa_snapshot[30][17] , \sa_snapshot[30].r.part0[17] );
tran (\sa_snapshot[30][17] , \sa_snapshot[30].f.lower[17] );
tran (\sa_snapshot[30][18] , \sa_snapshot[30].r.part0[18] );
tran (\sa_snapshot[30][18] , \sa_snapshot[30].f.lower[18] );
tran (\sa_snapshot[30][19] , \sa_snapshot[30].r.part0[19] );
tran (\sa_snapshot[30][19] , \sa_snapshot[30].f.lower[19] );
tran (\sa_snapshot[30][20] , \sa_snapshot[30].r.part0[20] );
tran (\sa_snapshot[30][20] , \sa_snapshot[30].f.lower[20] );
tran (\sa_snapshot[30][21] , \sa_snapshot[30].r.part0[21] );
tran (\sa_snapshot[30][21] , \sa_snapshot[30].f.lower[21] );
tran (\sa_snapshot[30][22] , \sa_snapshot[30].r.part0[22] );
tran (\sa_snapshot[30][22] , \sa_snapshot[30].f.lower[22] );
tran (\sa_snapshot[30][23] , \sa_snapshot[30].r.part0[23] );
tran (\sa_snapshot[30][23] , \sa_snapshot[30].f.lower[23] );
tran (\sa_snapshot[30][24] , \sa_snapshot[30].r.part0[24] );
tran (\sa_snapshot[30][24] , \sa_snapshot[30].f.lower[24] );
tran (\sa_snapshot[30][25] , \sa_snapshot[30].r.part0[25] );
tran (\sa_snapshot[30][25] , \sa_snapshot[30].f.lower[25] );
tran (\sa_snapshot[30][26] , \sa_snapshot[30].r.part0[26] );
tran (\sa_snapshot[30][26] , \sa_snapshot[30].f.lower[26] );
tran (\sa_snapshot[30][27] , \sa_snapshot[30].r.part0[27] );
tran (\sa_snapshot[30][27] , \sa_snapshot[30].f.lower[27] );
tran (\sa_snapshot[30][28] , \sa_snapshot[30].r.part0[28] );
tran (\sa_snapshot[30][28] , \sa_snapshot[30].f.lower[28] );
tran (\sa_snapshot[30][29] , \sa_snapshot[30].r.part0[29] );
tran (\sa_snapshot[30][29] , \sa_snapshot[30].f.lower[29] );
tran (\sa_snapshot[30][30] , \sa_snapshot[30].r.part0[30] );
tran (\sa_snapshot[30][30] , \sa_snapshot[30].f.lower[30] );
tran (\sa_snapshot[30][31] , \sa_snapshot[30].r.part0[31] );
tran (\sa_snapshot[30][31] , \sa_snapshot[30].f.lower[31] );
tran (\sa_snapshot[30][32] , \sa_snapshot[30].r.part1[0] );
tran (\sa_snapshot[30][32] , \sa_snapshot[30].f.upper[0] );
tran (\sa_snapshot[30][33] , \sa_snapshot[30].r.part1[1] );
tran (\sa_snapshot[30][33] , \sa_snapshot[30].f.upper[1] );
tran (\sa_snapshot[30][34] , \sa_snapshot[30].r.part1[2] );
tran (\sa_snapshot[30][34] , \sa_snapshot[30].f.upper[2] );
tran (\sa_snapshot[30][35] , \sa_snapshot[30].r.part1[3] );
tran (\sa_snapshot[30][35] , \sa_snapshot[30].f.upper[3] );
tran (\sa_snapshot[30][36] , \sa_snapshot[30].r.part1[4] );
tran (\sa_snapshot[30][36] , \sa_snapshot[30].f.upper[4] );
tran (\sa_snapshot[30][37] , \sa_snapshot[30].r.part1[5] );
tran (\sa_snapshot[30][37] , \sa_snapshot[30].f.upper[5] );
tran (\sa_snapshot[30][38] , \sa_snapshot[30].r.part1[6] );
tran (\sa_snapshot[30][38] , \sa_snapshot[30].f.upper[6] );
tran (\sa_snapshot[30][39] , \sa_snapshot[30].r.part1[7] );
tran (\sa_snapshot[30][39] , \sa_snapshot[30].f.upper[7] );
tran (\sa_snapshot[30][40] , \sa_snapshot[30].r.part1[8] );
tran (\sa_snapshot[30][40] , \sa_snapshot[30].f.upper[8] );
tran (\sa_snapshot[30][41] , \sa_snapshot[30].r.part1[9] );
tran (\sa_snapshot[30][41] , \sa_snapshot[30].f.upper[9] );
tran (\sa_snapshot[30][42] , \sa_snapshot[30].r.part1[10] );
tran (\sa_snapshot[30][42] , \sa_snapshot[30].f.upper[10] );
tran (\sa_snapshot[30][43] , \sa_snapshot[30].r.part1[11] );
tran (\sa_snapshot[30][43] , \sa_snapshot[30].f.upper[11] );
tran (\sa_snapshot[30][44] , \sa_snapshot[30].r.part1[12] );
tran (\sa_snapshot[30][44] , \sa_snapshot[30].f.upper[12] );
tran (\sa_snapshot[30][45] , \sa_snapshot[30].r.part1[13] );
tran (\sa_snapshot[30][45] , \sa_snapshot[30].f.upper[13] );
tran (\sa_snapshot[30][46] , \sa_snapshot[30].r.part1[14] );
tran (\sa_snapshot[30][46] , \sa_snapshot[30].f.upper[14] );
tran (\sa_snapshot[30][47] , \sa_snapshot[30].r.part1[15] );
tran (\sa_snapshot[30][47] , \sa_snapshot[30].f.upper[15] );
tran (\sa_snapshot[30][48] , \sa_snapshot[30].r.part1[16] );
tran (\sa_snapshot[30][48] , \sa_snapshot[30].f.upper[16] );
tran (\sa_snapshot[30][49] , \sa_snapshot[30].r.part1[17] );
tran (\sa_snapshot[30][49] , \sa_snapshot[30].f.upper[17] );
tran (\sa_snapshot[30][50] , \sa_snapshot[30].r.part1[18] );
tran (\sa_snapshot[30][50] , \sa_snapshot[30].f.unused[0] );
tran (\sa_snapshot[30][51] , \sa_snapshot[30].r.part1[19] );
tran (\sa_snapshot[30][51] , \sa_snapshot[30].f.unused[1] );
tran (\sa_snapshot[30][52] , \sa_snapshot[30].r.part1[20] );
tran (\sa_snapshot[30][52] , \sa_snapshot[30].f.unused[2] );
tran (\sa_snapshot[30][53] , \sa_snapshot[30].r.part1[21] );
tran (\sa_snapshot[30][53] , \sa_snapshot[30].f.unused[3] );
tran (\sa_snapshot[30][54] , \sa_snapshot[30].r.part1[22] );
tran (\sa_snapshot[30][54] , \sa_snapshot[30].f.unused[4] );
tran (\sa_snapshot[30][55] , \sa_snapshot[30].r.part1[23] );
tran (\sa_snapshot[30][55] , \sa_snapshot[30].f.unused[5] );
tran (\sa_snapshot[30][56] , \sa_snapshot[30].r.part1[24] );
tran (\sa_snapshot[30][56] , \sa_snapshot[30].f.unused[6] );
tran (\sa_snapshot[30][57] , \sa_snapshot[30].r.part1[25] );
tran (\sa_snapshot[30][57] , \sa_snapshot[30].f.unused[7] );
tran (\sa_snapshot[30][58] , \sa_snapshot[30].r.part1[26] );
tran (\sa_snapshot[30][58] , \sa_snapshot[30].f.unused[8] );
tran (\sa_snapshot[30][59] , \sa_snapshot[30].r.part1[27] );
tran (\sa_snapshot[30][59] , \sa_snapshot[30].f.unused[9] );
tran (\sa_snapshot[30][60] , \sa_snapshot[30].r.part1[28] );
tran (\sa_snapshot[30][60] , \sa_snapshot[30].f.unused[10] );
tran (\sa_snapshot[30][61] , \sa_snapshot[30].r.part1[29] );
tran (\sa_snapshot[30][61] , \sa_snapshot[30].f.unused[11] );
tran (\sa_snapshot[30][62] , \sa_snapshot[30].r.part1[30] );
tran (\sa_snapshot[30][62] , \sa_snapshot[30].f.unused[12] );
tran (\sa_snapshot[30][63] , \sa_snapshot[30].r.part1[31] );
tran (\sa_snapshot[30][63] , \sa_snapshot[30].f.unused[13] );
tran (\sa_snapshot[31][0] , \sa_snapshot[31].r.part0[0] );
tran (\sa_snapshot[31][0] , \sa_snapshot[31].f.lower[0] );
tran (\sa_snapshot[31][1] , \sa_snapshot[31].r.part0[1] );
tran (\sa_snapshot[31][1] , \sa_snapshot[31].f.lower[1] );
tran (\sa_snapshot[31][2] , \sa_snapshot[31].r.part0[2] );
tran (\sa_snapshot[31][2] , \sa_snapshot[31].f.lower[2] );
tran (\sa_snapshot[31][3] , \sa_snapshot[31].r.part0[3] );
tran (\sa_snapshot[31][3] , \sa_snapshot[31].f.lower[3] );
tran (\sa_snapshot[31][4] , \sa_snapshot[31].r.part0[4] );
tran (\sa_snapshot[31][4] , \sa_snapshot[31].f.lower[4] );
tran (\sa_snapshot[31][5] , \sa_snapshot[31].r.part0[5] );
tran (\sa_snapshot[31][5] , \sa_snapshot[31].f.lower[5] );
tran (\sa_snapshot[31][6] , \sa_snapshot[31].r.part0[6] );
tran (\sa_snapshot[31][6] , \sa_snapshot[31].f.lower[6] );
tran (\sa_snapshot[31][7] , \sa_snapshot[31].r.part0[7] );
tran (\sa_snapshot[31][7] , \sa_snapshot[31].f.lower[7] );
tran (\sa_snapshot[31][8] , \sa_snapshot[31].r.part0[8] );
tran (\sa_snapshot[31][8] , \sa_snapshot[31].f.lower[8] );
tran (\sa_snapshot[31][9] , \sa_snapshot[31].r.part0[9] );
tran (\sa_snapshot[31][9] , \sa_snapshot[31].f.lower[9] );
tran (\sa_snapshot[31][10] , \sa_snapshot[31].r.part0[10] );
tran (\sa_snapshot[31][10] , \sa_snapshot[31].f.lower[10] );
tran (\sa_snapshot[31][11] , \sa_snapshot[31].r.part0[11] );
tran (\sa_snapshot[31][11] , \sa_snapshot[31].f.lower[11] );
tran (\sa_snapshot[31][12] , \sa_snapshot[31].r.part0[12] );
tran (\sa_snapshot[31][12] , \sa_snapshot[31].f.lower[12] );
tran (\sa_snapshot[31][13] , \sa_snapshot[31].r.part0[13] );
tran (\sa_snapshot[31][13] , \sa_snapshot[31].f.lower[13] );
tran (\sa_snapshot[31][14] , \sa_snapshot[31].r.part0[14] );
tran (\sa_snapshot[31][14] , \sa_snapshot[31].f.lower[14] );
tran (\sa_snapshot[31][15] , \sa_snapshot[31].r.part0[15] );
tran (\sa_snapshot[31][15] , \sa_snapshot[31].f.lower[15] );
tran (\sa_snapshot[31][16] , \sa_snapshot[31].r.part0[16] );
tran (\sa_snapshot[31][16] , \sa_snapshot[31].f.lower[16] );
tran (\sa_snapshot[31][17] , \sa_snapshot[31].r.part0[17] );
tran (\sa_snapshot[31][17] , \sa_snapshot[31].f.lower[17] );
tran (\sa_snapshot[31][18] , \sa_snapshot[31].r.part0[18] );
tran (\sa_snapshot[31][18] , \sa_snapshot[31].f.lower[18] );
tran (\sa_snapshot[31][19] , \sa_snapshot[31].r.part0[19] );
tran (\sa_snapshot[31][19] , \sa_snapshot[31].f.lower[19] );
tran (\sa_snapshot[31][20] , \sa_snapshot[31].r.part0[20] );
tran (\sa_snapshot[31][20] , \sa_snapshot[31].f.lower[20] );
tran (\sa_snapshot[31][21] , \sa_snapshot[31].r.part0[21] );
tran (\sa_snapshot[31][21] , \sa_snapshot[31].f.lower[21] );
tran (\sa_snapshot[31][22] , \sa_snapshot[31].r.part0[22] );
tran (\sa_snapshot[31][22] , \sa_snapshot[31].f.lower[22] );
tran (\sa_snapshot[31][23] , \sa_snapshot[31].r.part0[23] );
tran (\sa_snapshot[31][23] , \sa_snapshot[31].f.lower[23] );
tran (\sa_snapshot[31][24] , \sa_snapshot[31].r.part0[24] );
tran (\sa_snapshot[31][24] , \sa_snapshot[31].f.lower[24] );
tran (\sa_snapshot[31][25] , \sa_snapshot[31].r.part0[25] );
tran (\sa_snapshot[31][25] , \sa_snapshot[31].f.lower[25] );
tran (\sa_snapshot[31][26] , \sa_snapshot[31].r.part0[26] );
tran (\sa_snapshot[31][26] , \sa_snapshot[31].f.lower[26] );
tran (\sa_snapshot[31][27] , \sa_snapshot[31].r.part0[27] );
tran (\sa_snapshot[31][27] , \sa_snapshot[31].f.lower[27] );
tran (\sa_snapshot[31][28] , \sa_snapshot[31].r.part0[28] );
tran (\sa_snapshot[31][28] , \sa_snapshot[31].f.lower[28] );
tran (\sa_snapshot[31][29] , \sa_snapshot[31].r.part0[29] );
tran (\sa_snapshot[31][29] , \sa_snapshot[31].f.lower[29] );
tran (\sa_snapshot[31][30] , \sa_snapshot[31].r.part0[30] );
tran (\sa_snapshot[31][30] , \sa_snapshot[31].f.lower[30] );
tran (\sa_snapshot[31][31] , \sa_snapshot[31].r.part0[31] );
tran (\sa_snapshot[31][31] , \sa_snapshot[31].f.lower[31] );
tran (\sa_snapshot[31][32] , \sa_snapshot[31].r.part1[0] );
tran (\sa_snapshot[31][32] , \sa_snapshot[31].f.upper[0] );
tran (\sa_snapshot[31][33] , \sa_snapshot[31].r.part1[1] );
tran (\sa_snapshot[31][33] , \sa_snapshot[31].f.upper[1] );
tran (\sa_snapshot[31][34] , \sa_snapshot[31].r.part1[2] );
tran (\sa_snapshot[31][34] , \sa_snapshot[31].f.upper[2] );
tran (\sa_snapshot[31][35] , \sa_snapshot[31].r.part1[3] );
tran (\sa_snapshot[31][35] , \sa_snapshot[31].f.upper[3] );
tran (\sa_snapshot[31][36] , \sa_snapshot[31].r.part1[4] );
tran (\sa_snapshot[31][36] , \sa_snapshot[31].f.upper[4] );
tran (\sa_snapshot[31][37] , \sa_snapshot[31].r.part1[5] );
tran (\sa_snapshot[31][37] , \sa_snapshot[31].f.upper[5] );
tran (\sa_snapshot[31][38] , \sa_snapshot[31].r.part1[6] );
tran (\sa_snapshot[31][38] , \sa_snapshot[31].f.upper[6] );
tran (\sa_snapshot[31][39] , \sa_snapshot[31].r.part1[7] );
tran (\sa_snapshot[31][39] , \sa_snapshot[31].f.upper[7] );
tran (\sa_snapshot[31][40] , \sa_snapshot[31].r.part1[8] );
tran (\sa_snapshot[31][40] , \sa_snapshot[31].f.upper[8] );
tran (\sa_snapshot[31][41] , \sa_snapshot[31].r.part1[9] );
tran (\sa_snapshot[31][41] , \sa_snapshot[31].f.upper[9] );
tran (\sa_snapshot[31][42] , \sa_snapshot[31].r.part1[10] );
tran (\sa_snapshot[31][42] , \sa_snapshot[31].f.upper[10] );
tran (\sa_snapshot[31][43] , \sa_snapshot[31].r.part1[11] );
tran (\sa_snapshot[31][43] , \sa_snapshot[31].f.upper[11] );
tran (\sa_snapshot[31][44] , \sa_snapshot[31].r.part1[12] );
tran (\sa_snapshot[31][44] , \sa_snapshot[31].f.upper[12] );
tran (\sa_snapshot[31][45] , \sa_snapshot[31].r.part1[13] );
tran (\sa_snapshot[31][45] , \sa_snapshot[31].f.upper[13] );
tran (\sa_snapshot[31][46] , \sa_snapshot[31].r.part1[14] );
tran (\sa_snapshot[31][46] , \sa_snapshot[31].f.upper[14] );
tran (\sa_snapshot[31][47] , \sa_snapshot[31].r.part1[15] );
tran (\sa_snapshot[31][47] , \sa_snapshot[31].f.upper[15] );
tran (\sa_snapshot[31][48] , \sa_snapshot[31].r.part1[16] );
tran (\sa_snapshot[31][48] , \sa_snapshot[31].f.upper[16] );
tran (\sa_snapshot[31][49] , \sa_snapshot[31].r.part1[17] );
tran (\sa_snapshot[31][49] , \sa_snapshot[31].f.upper[17] );
tran (\sa_snapshot[31][50] , \sa_snapshot[31].r.part1[18] );
tran (\sa_snapshot[31][50] , \sa_snapshot[31].f.unused[0] );
tran (\sa_snapshot[31][51] , \sa_snapshot[31].r.part1[19] );
tran (\sa_snapshot[31][51] , \sa_snapshot[31].f.unused[1] );
tran (\sa_snapshot[31][52] , \sa_snapshot[31].r.part1[20] );
tran (\sa_snapshot[31][52] , \sa_snapshot[31].f.unused[2] );
tran (\sa_snapshot[31][53] , \sa_snapshot[31].r.part1[21] );
tran (\sa_snapshot[31][53] , \sa_snapshot[31].f.unused[3] );
tran (\sa_snapshot[31][54] , \sa_snapshot[31].r.part1[22] );
tran (\sa_snapshot[31][54] , \sa_snapshot[31].f.unused[4] );
tran (\sa_snapshot[31][55] , \sa_snapshot[31].r.part1[23] );
tran (\sa_snapshot[31][55] , \sa_snapshot[31].f.unused[5] );
tran (\sa_snapshot[31][56] , \sa_snapshot[31].r.part1[24] );
tran (\sa_snapshot[31][56] , \sa_snapshot[31].f.unused[6] );
tran (\sa_snapshot[31][57] , \sa_snapshot[31].r.part1[25] );
tran (\sa_snapshot[31][57] , \sa_snapshot[31].f.unused[7] );
tran (\sa_snapshot[31][58] , \sa_snapshot[31].r.part1[26] );
tran (\sa_snapshot[31][58] , \sa_snapshot[31].f.unused[8] );
tran (\sa_snapshot[31][59] , \sa_snapshot[31].r.part1[27] );
tran (\sa_snapshot[31][59] , \sa_snapshot[31].f.unused[9] );
tran (\sa_snapshot[31][60] , \sa_snapshot[31].r.part1[28] );
tran (\sa_snapshot[31][60] , \sa_snapshot[31].f.unused[10] );
tran (\sa_snapshot[31][61] , \sa_snapshot[31].r.part1[29] );
tran (\sa_snapshot[31][61] , \sa_snapshot[31].f.unused[11] );
tran (\sa_snapshot[31][62] , \sa_snapshot[31].r.part1[30] );
tran (\sa_snapshot[31][62] , \sa_snapshot[31].f.unused[12] );
tran (\sa_snapshot[31][63] , \sa_snapshot[31].r.part1[31] );
tran (\sa_snapshot[31][63] , \sa_snapshot[31].f.unused[13] );
tran (\sa_count[0][0] , \sa_count[0].r.part0[0] );
tran (\sa_count[0][0] , \sa_count[0].f.lower[0] );
tran (\sa_count[0][1] , \sa_count[0].r.part0[1] );
tran (\sa_count[0][1] , \sa_count[0].f.lower[1] );
tran (\sa_count[0][2] , \sa_count[0].r.part0[2] );
tran (\sa_count[0][2] , \sa_count[0].f.lower[2] );
tran (\sa_count[0][3] , \sa_count[0].r.part0[3] );
tran (\sa_count[0][3] , \sa_count[0].f.lower[3] );
tran (\sa_count[0][4] , \sa_count[0].r.part0[4] );
tran (\sa_count[0][4] , \sa_count[0].f.lower[4] );
tran (\sa_count[0][5] , \sa_count[0].r.part0[5] );
tran (\sa_count[0][5] , \sa_count[0].f.lower[5] );
tran (\sa_count[0][6] , \sa_count[0].r.part0[6] );
tran (\sa_count[0][6] , \sa_count[0].f.lower[6] );
tran (\sa_count[0][7] , \sa_count[0].r.part0[7] );
tran (\sa_count[0][7] , \sa_count[0].f.lower[7] );
tran (\sa_count[0][8] , \sa_count[0].r.part0[8] );
tran (\sa_count[0][8] , \sa_count[0].f.lower[8] );
tran (\sa_count[0][9] , \sa_count[0].r.part0[9] );
tran (\sa_count[0][9] , \sa_count[0].f.lower[9] );
tran (\sa_count[0][10] , \sa_count[0].r.part0[10] );
tran (\sa_count[0][10] , \sa_count[0].f.lower[10] );
tran (\sa_count[0][11] , \sa_count[0].r.part0[11] );
tran (\sa_count[0][11] , \sa_count[0].f.lower[11] );
tran (\sa_count[0][12] , \sa_count[0].r.part0[12] );
tran (\sa_count[0][12] , \sa_count[0].f.lower[12] );
tran (\sa_count[0][13] , \sa_count[0].r.part0[13] );
tran (\sa_count[0][13] , \sa_count[0].f.lower[13] );
tran (\sa_count[0][14] , \sa_count[0].r.part0[14] );
tran (\sa_count[0][14] , \sa_count[0].f.lower[14] );
tran (\sa_count[0][15] , \sa_count[0].r.part0[15] );
tran (\sa_count[0][15] , \sa_count[0].f.lower[15] );
tran (\sa_count[0][16] , \sa_count[0].r.part0[16] );
tran (\sa_count[0][16] , \sa_count[0].f.lower[16] );
tran (\sa_count[0][17] , \sa_count[0].r.part0[17] );
tran (\sa_count[0][17] , \sa_count[0].f.lower[17] );
tran (\sa_count[0][18] , \sa_count[0].r.part0[18] );
tran (\sa_count[0][18] , \sa_count[0].f.lower[18] );
tran (\sa_count[0][19] , \sa_count[0].r.part0[19] );
tran (\sa_count[0][19] , \sa_count[0].f.lower[19] );
tran (\sa_count[0][20] , \sa_count[0].r.part0[20] );
tran (\sa_count[0][20] , \sa_count[0].f.lower[20] );
tran (\sa_count[0][21] , \sa_count[0].r.part0[21] );
tran (\sa_count[0][21] , \sa_count[0].f.lower[21] );
tran (\sa_count[0][22] , \sa_count[0].r.part0[22] );
tran (\sa_count[0][22] , \sa_count[0].f.lower[22] );
tran (\sa_count[0][23] , \sa_count[0].r.part0[23] );
tran (\sa_count[0][23] , \sa_count[0].f.lower[23] );
tran (\sa_count[0][24] , \sa_count[0].r.part0[24] );
tran (\sa_count[0][24] , \sa_count[0].f.lower[24] );
tran (\sa_count[0][25] , \sa_count[0].r.part0[25] );
tran (\sa_count[0][25] , \sa_count[0].f.lower[25] );
tran (\sa_count[0][26] , \sa_count[0].r.part0[26] );
tran (\sa_count[0][26] , \sa_count[0].f.lower[26] );
tran (\sa_count[0][27] , \sa_count[0].r.part0[27] );
tran (\sa_count[0][27] , \sa_count[0].f.lower[27] );
tran (\sa_count[0][28] , \sa_count[0].r.part0[28] );
tran (\sa_count[0][28] , \sa_count[0].f.lower[28] );
tran (\sa_count[0][29] , \sa_count[0].r.part0[29] );
tran (\sa_count[0][29] , \sa_count[0].f.lower[29] );
tran (\sa_count[0][30] , \sa_count[0].r.part0[30] );
tran (\sa_count[0][30] , \sa_count[0].f.lower[30] );
tran (\sa_count[0][31] , \sa_count[0].r.part0[31] );
tran (\sa_count[0][31] , \sa_count[0].f.lower[31] );
tran (\sa_count[0][32] , \sa_count[0].r.part1[0] );
tran (\sa_count[0][32] , \sa_count[0].f.upper[0] );
tran (\sa_count[0][33] , \sa_count[0].r.part1[1] );
tran (\sa_count[0][33] , \sa_count[0].f.upper[1] );
tran (\sa_count[0][34] , \sa_count[0].r.part1[2] );
tran (\sa_count[0][34] , \sa_count[0].f.upper[2] );
tran (\sa_count[0][35] , \sa_count[0].r.part1[3] );
tran (\sa_count[0][35] , \sa_count[0].f.upper[3] );
tran (\sa_count[0][36] , \sa_count[0].r.part1[4] );
tran (\sa_count[0][36] , \sa_count[0].f.upper[4] );
tran (\sa_count[0][37] , \sa_count[0].r.part1[5] );
tran (\sa_count[0][37] , \sa_count[0].f.upper[5] );
tran (\sa_count[0][38] , \sa_count[0].r.part1[6] );
tran (\sa_count[0][38] , \sa_count[0].f.upper[6] );
tran (\sa_count[0][39] , \sa_count[0].r.part1[7] );
tran (\sa_count[0][39] , \sa_count[0].f.upper[7] );
tran (\sa_count[0][40] , \sa_count[0].r.part1[8] );
tran (\sa_count[0][40] , \sa_count[0].f.upper[8] );
tran (\sa_count[0][41] , \sa_count[0].r.part1[9] );
tran (\sa_count[0][41] , \sa_count[0].f.upper[9] );
tran (\sa_count[0][42] , \sa_count[0].r.part1[10] );
tran (\sa_count[0][42] , \sa_count[0].f.upper[10] );
tran (\sa_count[0][43] , \sa_count[0].r.part1[11] );
tran (\sa_count[0][43] , \sa_count[0].f.upper[11] );
tran (\sa_count[0][44] , \sa_count[0].r.part1[12] );
tran (\sa_count[0][44] , \sa_count[0].f.upper[12] );
tran (\sa_count[0][45] , \sa_count[0].r.part1[13] );
tran (\sa_count[0][45] , \sa_count[0].f.upper[13] );
tran (\sa_count[0][46] , \sa_count[0].r.part1[14] );
tran (\sa_count[0][46] , \sa_count[0].f.upper[14] );
tran (\sa_count[0][47] , \sa_count[0].r.part1[15] );
tran (\sa_count[0][47] , \sa_count[0].f.upper[15] );
tran (\sa_count[0][48] , \sa_count[0].r.part1[16] );
tran (\sa_count[0][48] , \sa_count[0].f.upper[16] );
tran (\sa_count[0][49] , \sa_count[0].r.part1[17] );
tran (\sa_count[0][49] , \sa_count[0].f.upper[17] );
tran (\sa_count[0][50] , \sa_count[0].r.part1[18] );
tran (\sa_count[0][50] , \sa_count[0].f.unused[0] );
tran (\sa_count[0][51] , \sa_count[0].r.part1[19] );
tran (\sa_count[0][51] , \sa_count[0].f.unused[1] );
tran (\sa_count[0][52] , \sa_count[0].r.part1[20] );
tran (\sa_count[0][52] , \sa_count[0].f.unused[2] );
tran (\sa_count[0][53] , \sa_count[0].r.part1[21] );
tran (\sa_count[0][53] , \sa_count[0].f.unused[3] );
tran (\sa_count[0][54] , \sa_count[0].r.part1[22] );
tran (\sa_count[0][54] , \sa_count[0].f.unused[4] );
tran (\sa_count[0][55] , \sa_count[0].r.part1[23] );
tran (\sa_count[0][55] , \sa_count[0].f.unused[5] );
tran (\sa_count[0][56] , \sa_count[0].r.part1[24] );
tran (\sa_count[0][56] , \sa_count[0].f.unused[6] );
tran (\sa_count[0][57] , \sa_count[0].r.part1[25] );
tran (\sa_count[0][57] , \sa_count[0].f.unused[7] );
tran (\sa_count[0][58] , \sa_count[0].r.part1[26] );
tran (\sa_count[0][58] , \sa_count[0].f.unused[8] );
tran (\sa_count[0][59] , \sa_count[0].r.part1[27] );
tran (\sa_count[0][59] , \sa_count[0].f.unused[9] );
tran (\sa_count[0][60] , \sa_count[0].r.part1[28] );
tran (\sa_count[0][60] , \sa_count[0].f.unused[10] );
tran (\sa_count[0][61] , \sa_count[0].r.part1[29] );
tran (\sa_count[0][61] , \sa_count[0].f.unused[11] );
tran (\sa_count[0][62] , \sa_count[0].r.part1[30] );
tran (\sa_count[0][62] , \sa_count[0].f.unused[12] );
tran (\sa_count[0][63] , \sa_count[0].r.part1[31] );
tran (\sa_count[0][63] , \sa_count[0].f.unused[13] );
tran (\sa_count[1][0] , \sa_count[1].r.part0[0] );
tran (\sa_count[1][0] , \sa_count[1].f.lower[0] );
tran (\sa_count[1][1] , \sa_count[1].r.part0[1] );
tran (\sa_count[1][1] , \sa_count[1].f.lower[1] );
tran (\sa_count[1][2] , \sa_count[1].r.part0[2] );
tran (\sa_count[1][2] , \sa_count[1].f.lower[2] );
tran (\sa_count[1][3] , \sa_count[1].r.part0[3] );
tran (\sa_count[1][3] , \sa_count[1].f.lower[3] );
tran (\sa_count[1][4] , \sa_count[1].r.part0[4] );
tran (\sa_count[1][4] , \sa_count[1].f.lower[4] );
tran (\sa_count[1][5] , \sa_count[1].r.part0[5] );
tran (\sa_count[1][5] , \sa_count[1].f.lower[5] );
tran (\sa_count[1][6] , \sa_count[1].r.part0[6] );
tran (\sa_count[1][6] , \sa_count[1].f.lower[6] );
tran (\sa_count[1][7] , \sa_count[1].r.part0[7] );
tran (\sa_count[1][7] , \sa_count[1].f.lower[7] );
tran (\sa_count[1][8] , \sa_count[1].r.part0[8] );
tran (\sa_count[1][8] , \sa_count[1].f.lower[8] );
tran (\sa_count[1][9] , \sa_count[1].r.part0[9] );
tran (\sa_count[1][9] , \sa_count[1].f.lower[9] );
tran (\sa_count[1][10] , \sa_count[1].r.part0[10] );
tran (\sa_count[1][10] , \sa_count[1].f.lower[10] );
tran (\sa_count[1][11] , \sa_count[1].r.part0[11] );
tran (\sa_count[1][11] , \sa_count[1].f.lower[11] );
tran (\sa_count[1][12] , \sa_count[1].r.part0[12] );
tran (\sa_count[1][12] , \sa_count[1].f.lower[12] );
tran (\sa_count[1][13] , \sa_count[1].r.part0[13] );
tran (\sa_count[1][13] , \sa_count[1].f.lower[13] );
tran (\sa_count[1][14] , \sa_count[1].r.part0[14] );
tran (\sa_count[1][14] , \sa_count[1].f.lower[14] );
tran (\sa_count[1][15] , \sa_count[1].r.part0[15] );
tran (\sa_count[1][15] , \sa_count[1].f.lower[15] );
tran (\sa_count[1][16] , \sa_count[1].r.part0[16] );
tran (\sa_count[1][16] , \sa_count[1].f.lower[16] );
tran (\sa_count[1][17] , \sa_count[1].r.part0[17] );
tran (\sa_count[1][17] , \sa_count[1].f.lower[17] );
tran (\sa_count[1][18] , \sa_count[1].r.part0[18] );
tran (\sa_count[1][18] , \sa_count[1].f.lower[18] );
tran (\sa_count[1][19] , \sa_count[1].r.part0[19] );
tran (\sa_count[1][19] , \sa_count[1].f.lower[19] );
tran (\sa_count[1][20] , \sa_count[1].r.part0[20] );
tran (\sa_count[1][20] , \sa_count[1].f.lower[20] );
tran (\sa_count[1][21] , \sa_count[1].r.part0[21] );
tran (\sa_count[1][21] , \sa_count[1].f.lower[21] );
tran (\sa_count[1][22] , \sa_count[1].r.part0[22] );
tran (\sa_count[1][22] , \sa_count[1].f.lower[22] );
tran (\sa_count[1][23] , \sa_count[1].r.part0[23] );
tran (\sa_count[1][23] , \sa_count[1].f.lower[23] );
tran (\sa_count[1][24] , \sa_count[1].r.part0[24] );
tran (\sa_count[1][24] , \sa_count[1].f.lower[24] );
tran (\sa_count[1][25] , \sa_count[1].r.part0[25] );
tran (\sa_count[1][25] , \sa_count[1].f.lower[25] );
tran (\sa_count[1][26] , \sa_count[1].r.part0[26] );
tran (\sa_count[1][26] , \sa_count[1].f.lower[26] );
tran (\sa_count[1][27] , \sa_count[1].r.part0[27] );
tran (\sa_count[1][27] , \sa_count[1].f.lower[27] );
tran (\sa_count[1][28] , \sa_count[1].r.part0[28] );
tran (\sa_count[1][28] , \sa_count[1].f.lower[28] );
tran (\sa_count[1][29] , \sa_count[1].r.part0[29] );
tran (\sa_count[1][29] , \sa_count[1].f.lower[29] );
tran (\sa_count[1][30] , \sa_count[1].r.part0[30] );
tran (\sa_count[1][30] , \sa_count[1].f.lower[30] );
tran (\sa_count[1][31] , \sa_count[1].r.part0[31] );
tran (\sa_count[1][31] , \sa_count[1].f.lower[31] );
tran (\sa_count[1][32] , \sa_count[1].r.part1[0] );
tran (\sa_count[1][32] , \sa_count[1].f.upper[0] );
tran (\sa_count[1][33] , \sa_count[1].r.part1[1] );
tran (\sa_count[1][33] , \sa_count[1].f.upper[1] );
tran (\sa_count[1][34] , \sa_count[1].r.part1[2] );
tran (\sa_count[1][34] , \sa_count[1].f.upper[2] );
tran (\sa_count[1][35] , \sa_count[1].r.part1[3] );
tran (\sa_count[1][35] , \sa_count[1].f.upper[3] );
tran (\sa_count[1][36] , \sa_count[1].r.part1[4] );
tran (\sa_count[1][36] , \sa_count[1].f.upper[4] );
tran (\sa_count[1][37] , \sa_count[1].r.part1[5] );
tran (\sa_count[1][37] , \sa_count[1].f.upper[5] );
tran (\sa_count[1][38] , \sa_count[1].r.part1[6] );
tran (\sa_count[1][38] , \sa_count[1].f.upper[6] );
tran (\sa_count[1][39] , \sa_count[1].r.part1[7] );
tran (\sa_count[1][39] , \sa_count[1].f.upper[7] );
tran (\sa_count[1][40] , \sa_count[1].r.part1[8] );
tran (\sa_count[1][40] , \sa_count[1].f.upper[8] );
tran (\sa_count[1][41] , \sa_count[1].r.part1[9] );
tran (\sa_count[1][41] , \sa_count[1].f.upper[9] );
tran (\sa_count[1][42] , \sa_count[1].r.part1[10] );
tran (\sa_count[1][42] , \sa_count[1].f.upper[10] );
tran (\sa_count[1][43] , \sa_count[1].r.part1[11] );
tran (\sa_count[1][43] , \sa_count[1].f.upper[11] );
tran (\sa_count[1][44] , \sa_count[1].r.part1[12] );
tran (\sa_count[1][44] , \sa_count[1].f.upper[12] );
tran (\sa_count[1][45] , \sa_count[1].r.part1[13] );
tran (\sa_count[1][45] , \sa_count[1].f.upper[13] );
tran (\sa_count[1][46] , \sa_count[1].r.part1[14] );
tran (\sa_count[1][46] , \sa_count[1].f.upper[14] );
tran (\sa_count[1][47] , \sa_count[1].r.part1[15] );
tran (\sa_count[1][47] , \sa_count[1].f.upper[15] );
tran (\sa_count[1][48] , \sa_count[1].r.part1[16] );
tran (\sa_count[1][48] , \sa_count[1].f.upper[16] );
tran (\sa_count[1][49] , \sa_count[1].r.part1[17] );
tran (\sa_count[1][49] , \sa_count[1].f.upper[17] );
tran (\sa_count[1][50] , \sa_count[1].r.part1[18] );
tran (\sa_count[1][50] , \sa_count[1].f.unused[0] );
tran (\sa_count[1][51] , \sa_count[1].r.part1[19] );
tran (\sa_count[1][51] , \sa_count[1].f.unused[1] );
tran (\sa_count[1][52] , \sa_count[1].r.part1[20] );
tran (\sa_count[1][52] , \sa_count[1].f.unused[2] );
tran (\sa_count[1][53] , \sa_count[1].r.part1[21] );
tran (\sa_count[1][53] , \sa_count[1].f.unused[3] );
tran (\sa_count[1][54] , \sa_count[1].r.part1[22] );
tran (\sa_count[1][54] , \sa_count[1].f.unused[4] );
tran (\sa_count[1][55] , \sa_count[1].r.part1[23] );
tran (\sa_count[1][55] , \sa_count[1].f.unused[5] );
tran (\sa_count[1][56] , \sa_count[1].r.part1[24] );
tran (\sa_count[1][56] , \sa_count[1].f.unused[6] );
tran (\sa_count[1][57] , \sa_count[1].r.part1[25] );
tran (\sa_count[1][57] , \sa_count[1].f.unused[7] );
tran (\sa_count[1][58] , \sa_count[1].r.part1[26] );
tran (\sa_count[1][58] , \sa_count[1].f.unused[8] );
tran (\sa_count[1][59] , \sa_count[1].r.part1[27] );
tran (\sa_count[1][59] , \sa_count[1].f.unused[9] );
tran (\sa_count[1][60] , \sa_count[1].r.part1[28] );
tran (\sa_count[1][60] , \sa_count[1].f.unused[10] );
tran (\sa_count[1][61] , \sa_count[1].r.part1[29] );
tran (\sa_count[1][61] , \sa_count[1].f.unused[11] );
tran (\sa_count[1][62] , \sa_count[1].r.part1[30] );
tran (\sa_count[1][62] , \sa_count[1].f.unused[12] );
tran (\sa_count[1][63] , \sa_count[1].r.part1[31] );
tran (\sa_count[1][63] , \sa_count[1].f.unused[13] );
tran (\sa_count[2][0] , \sa_count[2].r.part0[0] );
tran (\sa_count[2][0] , \sa_count[2].f.lower[0] );
tran (\sa_count[2][1] , \sa_count[2].r.part0[1] );
tran (\sa_count[2][1] , \sa_count[2].f.lower[1] );
tran (\sa_count[2][2] , \sa_count[2].r.part0[2] );
tran (\sa_count[2][2] , \sa_count[2].f.lower[2] );
tran (\sa_count[2][3] , \sa_count[2].r.part0[3] );
tran (\sa_count[2][3] , \sa_count[2].f.lower[3] );
tran (\sa_count[2][4] , \sa_count[2].r.part0[4] );
tran (\sa_count[2][4] , \sa_count[2].f.lower[4] );
tran (\sa_count[2][5] , \sa_count[2].r.part0[5] );
tran (\sa_count[2][5] , \sa_count[2].f.lower[5] );
tran (\sa_count[2][6] , \sa_count[2].r.part0[6] );
tran (\sa_count[2][6] , \sa_count[2].f.lower[6] );
tran (\sa_count[2][7] , \sa_count[2].r.part0[7] );
tran (\sa_count[2][7] , \sa_count[2].f.lower[7] );
tran (\sa_count[2][8] , \sa_count[2].r.part0[8] );
tran (\sa_count[2][8] , \sa_count[2].f.lower[8] );
tran (\sa_count[2][9] , \sa_count[2].r.part0[9] );
tran (\sa_count[2][9] , \sa_count[2].f.lower[9] );
tran (\sa_count[2][10] , \sa_count[2].r.part0[10] );
tran (\sa_count[2][10] , \sa_count[2].f.lower[10] );
tran (\sa_count[2][11] , \sa_count[2].r.part0[11] );
tran (\sa_count[2][11] , \sa_count[2].f.lower[11] );
tran (\sa_count[2][12] , \sa_count[2].r.part0[12] );
tran (\sa_count[2][12] , \sa_count[2].f.lower[12] );
tran (\sa_count[2][13] , \sa_count[2].r.part0[13] );
tran (\sa_count[2][13] , \sa_count[2].f.lower[13] );
tran (\sa_count[2][14] , \sa_count[2].r.part0[14] );
tran (\sa_count[2][14] , \sa_count[2].f.lower[14] );
tran (\sa_count[2][15] , \sa_count[2].r.part0[15] );
tran (\sa_count[2][15] , \sa_count[2].f.lower[15] );
tran (\sa_count[2][16] , \sa_count[2].r.part0[16] );
tran (\sa_count[2][16] , \sa_count[2].f.lower[16] );
tran (\sa_count[2][17] , \sa_count[2].r.part0[17] );
tran (\sa_count[2][17] , \sa_count[2].f.lower[17] );
tran (\sa_count[2][18] , \sa_count[2].r.part0[18] );
tran (\sa_count[2][18] , \sa_count[2].f.lower[18] );
tran (\sa_count[2][19] , \sa_count[2].r.part0[19] );
tran (\sa_count[2][19] , \sa_count[2].f.lower[19] );
tran (\sa_count[2][20] , \sa_count[2].r.part0[20] );
tran (\sa_count[2][20] , \sa_count[2].f.lower[20] );
tran (\sa_count[2][21] , \sa_count[2].r.part0[21] );
tran (\sa_count[2][21] , \sa_count[2].f.lower[21] );
tran (\sa_count[2][22] , \sa_count[2].r.part0[22] );
tran (\sa_count[2][22] , \sa_count[2].f.lower[22] );
tran (\sa_count[2][23] , \sa_count[2].r.part0[23] );
tran (\sa_count[2][23] , \sa_count[2].f.lower[23] );
tran (\sa_count[2][24] , \sa_count[2].r.part0[24] );
tran (\sa_count[2][24] , \sa_count[2].f.lower[24] );
tran (\sa_count[2][25] , \sa_count[2].r.part0[25] );
tran (\sa_count[2][25] , \sa_count[2].f.lower[25] );
tran (\sa_count[2][26] , \sa_count[2].r.part0[26] );
tran (\sa_count[2][26] , \sa_count[2].f.lower[26] );
tran (\sa_count[2][27] , \sa_count[2].r.part0[27] );
tran (\sa_count[2][27] , \sa_count[2].f.lower[27] );
tran (\sa_count[2][28] , \sa_count[2].r.part0[28] );
tran (\sa_count[2][28] , \sa_count[2].f.lower[28] );
tran (\sa_count[2][29] , \sa_count[2].r.part0[29] );
tran (\sa_count[2][29] , \sa_count[2].f.lower[29] );
tran (\sa_count[2][30] , \sa_count[2].r.part0[30] );
tran (\sa_count[2][30] , \sa_count[2].f.lower[30] );
tran (\sa_count[2][31] , \sa_count[2].r.part0[31] );
tran (\sa_count[2][31] , \sa_count[2].f.lower[31] );
tran (\sa_count[2][32] , \sa_count[2].r.part1[0] );
tran (\sa_count[2][32] , \sa_count[2].f.upper[0] );
tran (\sa_count[2][33] , \sa_count[2].r.part1[1] );
tran (\sa_count[2][33] , \sa_count[2].f.upper[1] );
tran (\sa_count[2][34] , \sa_count[2].r.part1[2] );
tran (\sa_count[2][34] , \sa_count[2].f.upper[2] );
tran (\sa_count[2][35] , \sa_count[2].r.part1[3] );
tran (\sa_count[2][35] , \sa_count[2].f.upper[3] );
tran (\sa_count[2][36] , \sa_count[2].r.part1[4] );
tran (\sa_count[2][36] , \sa_count[2].f.upper[4] );
tran (\sa_count[2][37] , \sa_count[2].r.part1[5] );
tran (\sa_count[2][37] , \sa_count[2].f.upper[5] );
tran (\sa_count[2][38] , \sa_count[2].r.part1[6] );
tran (\sa_count[2][38] , \sa_count[2].f.upper[6] );
tran (\sa_count[2][39] , \sa_count[2].r.part1[7] );
tran (\sa_count[2][39] , \sa_count[2].f.upper[7] );
tran (\sa_count[2][40] , \sa_count[2].r.part1[8] );
tran (\sa_count[2][40] , \sa_count[2].f.upper[8] );
tran (\sa_count[2][41] , \sa_count[2].r.part1[9] );
tran (\sa_count[2][41] , \sa_count[2].f.upper[9] );
tran (\sa_count[2][42] , \sa_count[2].r.part1[10] );
tran (\sa_count[2][42] , \sa_count[2].f.upper[10] );
tran (\sa_count[2][43] , \sa_count[2].r.part1[11] );
tran (\sa_count[2][43] , \sa_count[2].f.upper[11] );
tran (\sa_count[2][44] , \sa_count[2].r.part1[12] );
tran (\sa_count[2][44] , \sa_count[2].f.upper[12] );
tran (\sa_count[2][45] , \sa_count[2].r.part1[13] );
tran (\sa_count[2][45] , \sa_count[2].f.upper[13] );
tran (\sa_count[2][46] , \sa_count[2].r.part1[14] );
tran (\sa_count[2][46] , \sa_count[2].f.upper[14] );
tran (\sa_count[2][47] , \sa_count[2].r.part1[15] );
tran (\sa_count[2][47] , \sa_count[2].f.upper[15] );
tran (\sa_count[2][48] , \sa_count[2].r.part1[16] );
tran (\sa_count[2][48] , \sa_count[2].f.upper[16] );
tran (\sa_count[2][49] , \sa_count[2].r.part1[17] );
tran (\sa_count[2][49] , \sa_count[2].f.upper[17] );
tran (\sa_count[2][50] , \sa_count[2].r.part1[18] );
tran (\sa_count[2][50] , \sa_count[2].f.unused[0] );
tran (\sa_count[2][51] , \sa_count[2].r.part1[19] );
tran (\sa_count[2][51] , \sa_count[2].f.unused[1] );
tran (\sa_count[2][52] , \sa_count[2].r.part1[20] );
tran (\sa_count[2][52] , \sa_count[2].f.unused[2] );
tran (\sa_count[2][53] , \sa_count[2].r.part1[21] );
tran (\sa_count[2][53] , \sa_count[2].f.unused[3] );
tran (\sa_count[2][54] , \sa_count[2].r.part1[22] );
tran (\sa_count[2][54] , \sa_count[2].f.unused[4] );
tran (\sa_count[2][55] , \sa_count[2].r.part1[23] );
tran (\sa_count[2][55] , \sa_count[2].f.unused[5] );
tran (\sa_count[2][56] , \sa_count[2].r.part1[24] );
tran (\sa_count[2][56] , \sa_count[2].f.unused[6] );
tran (\sa_count[2][57] , \sa_count[2].r.part1[25] );
tran (\sa_count[2][57] , \sa_count[2].f.unused[7] );
tran (\sa_count[2][58] , \sa_count[2].r.part1[26] );
tran (\sa_count[2][58] , \sa_count[2].f.unused[8] );
tran (\sa_count[2][59] , \sa_count[2].r.part1[27] );
tran (\sa_count[2][59] , \sa_count[2].f.unused[9] );
tran (\sa_count[2][60] , \sa_count[2].r.part1[28] );
tran (\sa_count[2][60] , \sa_count[2].f.unused[10] );
tran (\sa_count[2][61] , \sa_count[2].r.part1[29] );
tran (\sa_count[2][61] , \sa_count[2].f.unused[11] );
tran (\sa_count[2][62] , \sa_count[2].r.part1[30] );
tran (\sa_count[2][62] , \sa_count[2].f.unused[12] );
tran (\sa_count[2][63] , \sa_count[2].r.part1[31] );
tran (\sa_count[2][63] , \sa_count[2].f.unused[13] );
tran (\sa_count[3][0] , \sa_count[3].r.part0[0] );
tran (\sa_count[3][0] , \sa_count[3].f.lower[0] );
tran (\sa_count[3][1] , \sa_count[3].r.part0[1] );
tran (\sa_count[3][1] , \sa_count[3].f.lower[1] );
tran (\sa_count[3][2] , \sa_count[3].r.part0[2] );
tran (\sa_count[3][2] , \sa_count[3].f.lower[2] );
tran (\sa_count[3][3] , \sa_count[3].r.part0[3] );
tran (\sa_count[3][3] , \sa_count[3].f.lower[3] );
tran (\sa_count[3][4] , \sa_count[3].r.part0[4] );
tran (\sa_count[3][4] , \sa_count[3].f.lower[4] );
tran (\sa_count[3][5] , \sa_count[3].r.part0[5] );
tran (\sa_count[3][5] , \sa_count[3].f.lower[5] );
tran (\sa_count[3][6] , \sa_count[3].r.part0[6] );
tran (\sa_count[3][6] , \sa_count[3].f.lower[6] );
tran (\sa_count[3][7] , \sa_count[3].r.part0[7] );
tran (\sa_count[3][7] , \sa_count[3].f.lower[7] );
tran (\sa_count[3][8] , \sa_count[3].r.part0[8] );
tran (\sa_count[3][8] , \sa_count[3].f.lower[8] );
tran (\sa_count[3][9] , \sa_count[3].r.part0[9] );
tran (\sa_count[3][9] , \sa_count[3].f.lower[9] );
tran (\sa_count[3][10] , \sa_count[3].r.part0[10] );
tran (\sa_count[3][10] , \sa_count[3].f.lower[10] );
tran (\sa_count[3][11] , \sa_count[3].r.part0[11] );
tran (\sa_count[3][11] , \sa_count[3].f.lower[11] );
tran (\sa_count[3][12] , \sa_count[3].r.part0[12] );
tran (\sa_count[3][12] , \sa_count[3].f.lower[12] );
tran (\sa_count[3][13] , \sa_count[3].r.part0[13] );
tran (\sa_count[3][13] , \sa_count[3].f.lower[13] );
tran (\sa_count[3][14] , \sa_count[3].r.part0[14] );
tran (\sa_count[3][14] , \sa_count[3].f.lower[14] );
tran (\sa_count[3][15] , \sa_count[3].r.part0[15] );
tran (\sa_count[3][15] , \sa_count[3].f.lower[15] );
tran (\sa_count[3][16] , \sa_count[3].r.part0[16] );
tran (\sa_count[3][16] , \sa_count[3].f.lower[16] );
tran (\sa_count[3][17] , \sa_count[3].r.part0[17] );
tran (\sa_count[3][17] , \sa_count[3].f.lower[17] );
tran (\sa_count[3][18] , \sa_count[3].r.part0[18] );
tran (\sa_count[3][18] , \sa_count[3].f.lower[18] );
tran (\sa_count[3][19] , \sa_count[3].r.part0[19] );
tran (\sa_count[3][19] , \sa_count[3].f.lower[19] );
tran (\sa_count[3][20] , \sa_count[3].r.part0[20] );
tran (\sa_count[3][20] , \sa_count[3].f.lower[20] );
tran (\sa_count[3][21] , \sa_count[3].r.part0[21] );
tran (\sa_count[3][21] , \sa_count[3].f.lower[21] );
tran (\sa_count[3][22] , \sa_count[3].r.part0[22] );
tran (\sa_count[3][22] , \sa_count[3].f.lower[22] );
tran (\sa_count[3][23] , \sa_count[3].r.part0[23] );
tran (\sa_count[3][23] , \sa_count[3].f.lower[23] );
tran (\sa_count[3][24] , \sa_count[3].r.part0[24] );
tran (\sa_count[3][24] , \sa_count[3].f.lower[24] );
tran (\sa_count[3][25] , \sa_count[3].r.part0[25] );
tran (\sa_count[3][25] , \sa_count[3].f.lower[25] );
tran (\sa_count[3][26] , \sa_count[3].r.part0[26] );
tran (\sa_count[3][26] , \sa_count[3].f.lower[26] );
tran (\sa_count[3][27] , \sa_count[3].r.part0[27] );
tran (\sa_count[3][27] , \sa_count[3].f.lower[27] );
tran (\sa_count[3][28] , \sa_count[3].r.part0[28] );
tran (\sa_count[3][28] , \sa_count[3].f.lower[28] );
tran (\sa_count[3][29] , \sa_count[3].r.part0[29] );
tran (\sa_count[3][29] , \sa_count[3].f.lower[29] );
tran (\sa_count[3][30] , \sa_count[3].r.part0[30] );
tran (\sa_count[3][30] , \sa_count[3].f.lower[30] );
tran (\sa_count[3][31] , \sa_count[3].r.part0[31] );
tran (\sa_count[3][31] , \sa_count[3].f.lower[31] );
tran (\sa_count[3][32] , \sa_count[3].r.part1[0] );
tran (\sa_count[3][32] , \sa_count[3].f.upper[0] );
tran (\sa_count[3][33] , \sa_count[3].r.part1[1] );
tran (\sa_count[3][33] , \sa_count[3].f.upper[1] );
tran (\sa_count[3][34] , \sa_count[3].r.part1[2] );
tran (\sa_count[3][34] , \sa_count[3].f.upper[2] );
tran (\sa_count[3][35] , \sa_count[3].r.part1[3] );
tran (\sa_count[3][35] , \sa_count[3].f.upper[3] );
tran (\sa_count[3][36] , \sa_count[3].r.part1[4] );
tran (\sa_count[3][36] , \sa_count[3].f.upper[4] );
tran (\sa_count[3][37] , \sa_count[3].r.part1[5] );
tran (\sa_count[3][37] , \sa_count[3].f.upper[5] );
tran (\sa_count[3][38] , \sa_count[3].r.part1[6] );
tran (\sa_count[3][38] , \sa_count[3].f.upper[6] );
tran (\sa_count[3][39] , \sa_count[3].r.part1[7] );
tran (\sa_count[3][39] , \sa_count[3].f.upper[7] );
tran (\sa_count[3][40] , \sa_count[3].r.part1[8] );
tran (\sa_count[3][40] , \sa_count[3].f.upper[8] );
tran (\sa_count[3][41] , \sa_count[3].r.part1[9] );
tran (\sa_count[3][41] , \sa_count[3].f.upper[9] );
tran (\sa_count[3][42] , \sa_count[3].r.part1[10] );
tran (\sa_count[3][42] , \sa_count[3].f.upper[10] );
tran (\sa_count[3][43] , \sa_count[3].r.part1[11] );
tran (\sa_count[3][43] , \sa_count[3].f.upper[11] );
tran (\sa_count[3][44] , \sa_count[3].r.part1[12] );
tran (\sa_count[3][44] , \sa_count[3].f.upper[12] );
tran (\sa_count[3][45] , \sa_count[3].r.part1[13] );
tran (\sa_count[3][45] , \sa_count[3].f.upper[13] );
tran (\sa_count[3][46] , \sa_count[3].r.part1[14] );
tran (\sa_count[3][46] , \sa_count[3].f.upper[14] );
tran (\sa_count[3][47] , \sa_count[3].r.part1[15] );
tran (\sa_count[3][47] , \sa_count[3].f.upper[15] );
tran (\sa_count[3][48] , \sa_count[3].r.part1[16] );
tran (\sa_count[3][48] , \sa_count[3].f.upper[16] );
tran (\sa_count[3][49] , \sa_count[3].r.part1[17] );
tran (\sa_count[3][49] , \sa_count[3].f.upper[17] );
tran (\sa_count[3][50] , \sa_count[3].r.part1[18] );
tran (\sa_count[3][50] , \sa_count[3].f.unused[0] );
tran (\sa_count[3][51] , \sa_count[3].r.part1[19] );
tran (\sa_count[3][51] , \sa_count[3].f.unused[1] );
tran (\sa_count[3][52] , \sa_count[3].r.part1[20] );
tran (\sa_count[3][52] , \sa_count[3].f.unused[2] );
tran (\sa_count[3][53] , \sa_count[3].r.part1[21] );
tran (\sa_count[3][53] , \sa_count[3].f.unused[3] );
tran (\sa_count[3][54] , \sa_count[3].r.part1[22] );
tran (\sa_count[3][54] , \sa_count[3].f.unused[4] );
tran (\sa_count[3][55] , \sa_count[3].r.part1[23] );
tran (\sa_count[3][55] , \sa_count[3].f.unused[5] );
tran (\sa_count[3][56] , \sa_count[3].r.part1[24] );
tran (\sa_count[3][56] , \sa_count[3].f.unused[6] );
tran (\sa_count[3][57] , \sa_count[3].r.part1[25] );
tran (\sa_count[3][57] , \sa_count[3].f.unused[7] );
tran (\sa_count[3][58] , \sa_count[3].r.part1[26] );
tran (\sa_count[3][58] , \sa_count[3].f.unused[8] );
tran (\sa_count[3][59] , \sa_count[3].r.part1[27] );
tran (\sa_count[3][59] , \sa_count[3].f.unused[9] );
tran (\sa_count[3][60] , \sa_count[3].r.part1[28] );
tran (\sa_count[3][60] , \sa_count[3].f.unused[10] );
tran (\sa_count[3][61] , \sa_count[3].r.part1[29] );
tran (\sa_count[3][61] , \sa_count[3].f.unused[11] );
tran (\sa_count[3][62] , \sa_count[3].r.part1[30] );
tran (\sa_count[3][62] , \sa_count[3].f.unused[12] );
tran (\sa_count[3][63] , \sa_count[3].r.part1[31] );
tran (\sa_count[3][63] , \sa_count[3].f.unused[13] );
tran (\sa_count[4][0] , \sa_count[4].r.part0[0] );
tran (\sa_count[4][0] , \sa_count[4].f.lower[0] );
tran (\sa_count[4][1] , \sa_count[4].r.part0[1] );
tran (\sa_count[4][1] , \sa_count[4].f.lower[1] );
tran (\sa_count[4][2] , \sa_count[4].r.part0[2] );
tran (\sa_count[4][2] , \sa_count[4].f.lower[2] );
tran (\sa_count[4][3] , \sa_count[4].r.part0[3] );
tran (\sa_count[4][3] , \sa_count[4].f.lower[3] );
tran (\sa_count[4][4] , \sa_count[4].r.part0[4] );
tran (\sa_count[4][4] , \sa_count[4].f.lower[4] );
tran (\sa_count[4][5] , \sa_count[4].r.part0[5] );
tran (\sa_count[4][5] , \sa_count[4].f.lower[5] );
tran (\sa_count[4][6] , \sa_count[4].r.part0[6] );
tran (\sa_count[4][6] , \sa_count[4].f.lower[6] );
tran (\sa_count[4][7] , \sa_count[4].r.part0[7] );
tran (\sa_count[4][7] , \sa_count[4].f.lower[7] );
tran (\sa_count[4][8] , \sa_count[4].r.part0[8] );
tran (\sa_count[4][8] , \sa_count[4].f.lower[8] );
tran (\sa_count[4][9] , \sa_count[4].r.part0[9] );
tran (\sa_count[4][9] , \sa_count[4].f.lower[9] );
tran (\sa_count[4][10] , \sa_count[4].r.part0[10] );
tran (\sa_count[4][10] , \sa_count[4].f.lower[10] );
tran (\sa_count[4][11] , \sa_count[4].r.part0[11] );
tran (\sa_count[4][11] , \sa_count[4].f.lower[11] );
tran (\sa_count[4][12] , \sa_count[4].r.part0[12] );
tran (\sa_count[4][12] , \sa_count[4].f.lower[12] );
tran (\sa_count[4][13] , \sa_count[4].r.part0[13] );
tran (\sa_count[4][13] , \sa_count[4].f.lower[13] );
tran (\sa_count[4][14] , \sa_count[4].r.part0[14] );
tran (\sa_count[4][14] , \sa_count[4].f.lower[14] );
tran (\sa_count[4][15] , \sa_count[4].r.part0[15] );
tran (\sa_count[4][15] , \sa_count[4].f.lower[15] );
tran (\sa_count[4][16] , \sa_count[4].r.part0[16] );
tran (\sa_count[4][16] , \sa_count[4].f.lower[16] );
tran (\sa_count[4][17] , \sa_count[4].r.part0[17] );
tran (\sa_count[4][17] , \sa_count[4].f.lower[17] );
tran (\sa_count[4][18] , \sa_count[4].r.part0[18] );
tran (\sa_count[4][18] , \sa_count[4].f.lower[18] );
tran (\sa_count[4][19] , \sa_count[4].r.part0[19] );
tran (\sa_count[4][19] , \sa_count[4].f.lower[19] );
tran (\sa_count[4][20] , \sa_count[4].r.part0[20] );
tran (\sa_count[4][20] , \sa_count[4].f.lower[20] );
tran (\sa_count[4][21] , \sa_count[4].r.part0[21] );
tran (\sa_count[4][21] , \sa_count[4].f.lower[21] );
tran (\sa_count[4][22] , \sa_count[4].r.part0[22] );
tran (\sa_count[4][22] , \sa_count[4].f.lower[22] );
tran (\sa_count[4][23] , \sa_count[4].r.part0[23] );
tran (\sa_count[4][23] , \sa_count[4].f.lower[23] );
tran (\sa_count[4][24] , \sa_count[4].r.part0[24] );
tran (\sa_count[4][24] , \sa_count[4].f.lower[24] );
tran (\sa_count[4][25] , \sa_count[4].r.part0[25] );
tran (\sa_count[4][25] , \sa_count[4].f.lower[25] );
tran (\sa_count[4][26] , \sa_count[4].r.part0[26] );
tran (\sa_count[4][26] , \sa_count[4].f.lower[26] );
tran (\sa_count[4][27] , \sa_count[4].r.part0[27] );
tran (\sa_count[4][27] , \sa_count[4].f.lower[27] );
tran (\sa_count[4][28] , \sa_count[4].r.part0[28] );
tran (\sa_count[4][28] , \sa_count[4].f.lower[28] );
tran (\sa_count[4][29] , \sa_count[4].r.part0[29] );
tran (\sa_count[4][29] , \sa_count[4].f.lower[29] );
tran (\sa_count[4][30] , \sa_count[4].r.part0[30] );
tran (\sa_count[4][30] , \sa_count[4].f.lower[30] );
tran (\sa_count[4][31] , \sa_count[4].r.part0[31] );
tran (\sa_count[4][31] , \sa_count[4].f.lower[31] );
tran (\sa_count[4][32] , \sa_count[4].r.part1[0] );
tran (\sa_count[4][32] , \sa_count[4].f.upper[0] );
tran (\sa_count[4][33] , \sa_count[4].r.part1[1] );
tran (\sa_count[4][33] , \sa_count[4].f.upper[1] );
tran (\sa_count[4][34] , \sa_count[4].r.part1[2] );
tran (\sa_count[4][34] , \sa_count[4].f.upper[2] );
tran (\sa_count[4][35] , \sa_count[4].r.part1[3] );
tran (\sa_count[4][35] , \sa_count[4].f.upper[3] );
tran (\sa_count[4][36] , \sa_count[4].r.part1[4] );
tran (\sa_count[4][36] , \sa_count[4].f.upper[4] );
tran (\sa_count[4][37] , \sa_count[4].r.part1[5] );
tran (\sa_count[4][37] , \sa_count[4].f.upper[5] );
tran (\sa_count[4][38] , \sa_count[4].r.part1[6] );
tran (\sa_count[4][38] , \sa_count[4].f.upper[6] );
tran (\sa_count[4][39] , \sa_count[4].r.part1[7] );
tran (\sa_count[4][39] , \sa_count[4].f.upper[7] );
tran (\sa_count[4][40] , \sa_count[4].r.part1[8] );
tran (\sa_count[4][40] , \sa_count[4].f.upper[8] );
tran (\sa_count[4][41] , \sa_count[4].r.part1[9] );
tran (\sa_count[4][41] , \sa_count[4].f.upper[9] );
tran (\sa_count[4][42] , \sa_count[4].r.part1[10] );
tran (\sa_count[4][42] , \sa_count[4].f.upper[10] );
tran (\sa_count[4][43] , \sa_count[4].r.part1[11] );
tran (\sa_count[4][43] , \sa_count[4].f.upper[11] );
tran (\sa_count[4][44] , \sa_count[4].r.part1[12] );
tran (\sa_count[4][44] , \sa_count[4].f.upper[12] );
tran (\sa_count[4][45] , \sa_count[4].r.part1[13] );
tran (\sa_count[4][45] , \sa_count[4].f.upper[13] );
tran (\sa_count[4][46] , \sa_count[4].r.part1[14] );
tran (\sa_count[4][46] , \sa_count[4].f.upper[14] );
tran (\sa_count[4][47] , \sa_count[4].r.part1[15] );
tran (\sa_count[4][47] , \sa_count[4].f.upper[15] );
tran (\sa_count[4][48] , \sa_count[4].r.part1[16] );
tran (\sa_count[4][48] , \sa_count[4].f.upper[16] );
tran (\sa_count[4][49] , \sa_count[4].r.part1[17] );
tran (\sa_count[4][49] , \sa_count[4].f.upper[17] );
tran (\sa_count[4][50] , \sa_count[4].r.part1[18] );
tran (\sa_count[4][50] , \sa_count[4].f.unused[0] );
tran (\sa_count[4][51] , \sa_count[4].r.part1[19] );
tran (\sa_count[4][51] , \sa_count[4].f.unused[1] );
tran (\sa_count[4][52] , \sa_count[4].r.part1[20] );
tran (\sa_count[4][52] , \sa_count[4].f.unused[2] );
tran (\sa_count[4][53] , \sa_count[4].r.part1[21] );
tran (\sa_count[4][53] , \sa_count[4].f.unused[3] );
tran (\sa_count[4][54] , \sa_count[4].r.part1[22] );
tran (\sa_count[4][54] , \sa_count[4].f.unused[4] );
tran (\sa_count[4][55] , \sa_count[4].r.part1[23] );
tran (\sa_count[4][55] , \sa_count[4].f.unused[5] );
tran (\sa_count[4][56] , \sa_count[4].r.part1[24] );
tran (\sa_count[4][56] , \sa_count[4].f.unused[6] );
tran (\sa_count[4][57] , \sa_count[4].r.part1[25] );
tran (\sa_count[4][57] , \sa_count[4].f.unused[7] );
tran (\sa_count[4][58] , \sa_count[4].r.part1[26] );
tran (\sa_count[4][58] , \sa_count[4].f.unused[8] );
tran (\sa_count[4][59] , \sa_count[4].r.part1[27] );
tran (\sa_count[4][59] , \sa_count[4].f.unused[9] );
tran (\sa_count[4][60] , \sa_count[4].r.part1[28] );
tran (\sa_count[4][60] , \sa_count[4].f.unused[10] );
tran (\sa_count[4][61] , \sa_count[4].r.part1[29] );
tran (\sa_count[4][61] , \sa_count[4].f.unused[11] );
tran (\sa_count[4][62] , \sa_count[4].r.part1[30] );
tran (\sa_count[4][62] , \sa_count[4].f.unused[12] );
tran (\sa_count[4][63] , \sa_count[4].r.part1[31] );
tran (\sa_count[4][63] , \sa_count[4].f.unused[13] );
tran (\sa_count[5][0] , \sa_count[5].r.part0[0] );
tran (\sa_count[5][0] , \sa_count[5].f.lower[0] );
tran (\sa_count[5][1] , \sa_count[5].r.part0[1] );
tran (\sa_count[5][1] , \sa_count[5].f.lower[1] );
tran (\sa_count[5][2] , \sa_count[5].r.part0[2] );
tran (\sa_count[5][2] , \sa_count[5].f.lower[2] );
tran (\sa_count[5][3] , \sa_count[5].r.part0[3] );
tran (\sa_count[5][3] , \sa_count[5].f.lower[3] );
tran (\sa_count[5][4] , \sa_count[5].r.part0[4] );
tran (\sa_count[5][4] , \sa_count[5].f.lower[4] );
tran (\sa_count[5][5] , \sa_count[5].r.part0[5] );
tran (\sa_count[5][5] , \sa_count[5].f.lower[5] );
tran (\sa_count[5][6] , \sa_count[5].r.part0[6] );
tran (\sa_count[5][6] , \sa_count[5].f.lower[6] );
tran (\sa_count[5][7] , \sa_count[5].r.part0[7] );
tran (\sa_count[5][7] , \sa_count[5].f.lower[7] );
tran (\sa_count[5][8] , \sa_count[5].r.part0[8] );
tran (\sa_count[5][8] , \sa_count[5].f.lower[8] );
tran (\sa_count[5][9] , \sa_count[5].r.part0[9] );
tran (\sa_count[5][9] , \sa_count[5].f.lower[9] );
tran (\sa_count[5][10] , \sa_count[5].r.part0[10] );
tran (\sa_count[5][10] , \sa_count[5].f.lower[10] );
tran (\sa_count[5][11] , \sa_count[5].r.part0[11] );
tran (\sa_count[5][11] , \sa_count[5].f.lower[11] );
tran (\sa_count[5][12] , \sa_count[5].r.part0[12] );
tran (\sa_count[5][12] , \sa_count[5].f.lower[12] );
tran (\sa_count[5][13] , \sa_count[5].r.part0[13] );
tran (\sa_count[5][13] , \sa_count[5].f.lower[13] );
tran (\sa_count[5][14] , \sa_count[5].r.part0[14] );
tran (\sa_count[5][14] , \sa_count[5].f.lower[14] );
tran (\sa_count[5][15] , \sa_count[5].r.part0[15] );
tran (\sa_count[5][15] , \sa_count[5].f.lower[15] );
tran (\sa_count[5][16] , \sa_count[5].r.part0[16] );
tran (\sa_count[5][16] , \sa_count[5].f.lower[16] );
tran (\sa_count[5][17] , \sa_count[5].r.part0[17] );
tran (\sa_count[5][17] , \sa_count[5].f.lower[17] );
tran (\sa_count[5][18] , \sa_count[5].r.part0[18] );
tran (\sa_count[5][18] , \sa_count[5].f.lower[18] );
tran (\sa_count[5][19] , \sa_count[5].r.part0[19] );
tran (\sa_count[5][19] , \sa_count[5].f.lower[19] );
tran (\sa_count[5][20] , \sa_count[5].r.part0[20] );
tran (\sa_count[5][20] , \sa_count[5].f.lower[20] );
tran (\sa_count[5][21] , \sa_count[5].r.part0[21] );
tran (\sa_count[5][21] , \sa_count[5].f.lower[21] );
tran (\sa_count[5][22] , \sa_count[5].r.part0[22] );
tran (\sa_count[5][22] , \sa_count[5].f.lower[22] );
tran (\sa_count[5][23] , \sa_count[5].r.part0[23] );
tran (\sa_count[5][23] , \sa_count[5].f.lower[23] );
tran (\sa_count[5][24] , \sa_count[5].r.part0[24] );
tran (\sa_count[5][24] , \sa_count[5].f.lower[24] );
tran (\sa_count[5][25] , \sa_count[5].r.part0[25] );
tran (\sa_count[5][25] , \sa_count[5].f.lower[25] );
tran (\sa_count[5][26] , \sa_count[5].r.part0[26] );
tran (\sa_count[5][26] , \sa_count[5].f.lower[26] );
tran (\sa_count[5][27] , \sa_count[5].r.part0[27] );
tran (\sa_count[5][27] , \sa_count[5].f.lower[27] );
tran (\sa_count[5][28] , \sa_count[5].r.part0[28] );
tran (\sa_count[5][28] , \sa_count[5].f.lower[28] );
tran (\sa_count[5][29] , \sa_count[5].r.part0[29] );
tran (\sa_count[5][29] , \sa_count[5].f.lower[29] );
tran (\sa_count[5][30] , \sa_count[5].r.part0[30] );
tran (\sa_count[5][30] , \sa_count[5].f.lower[30] );
tran (\sa_count[5][31] , \sa_count[5].r.part0[31] );
tran (\sa_count[5][31] , \sa_count[5].f.lower[31] );
tran (\sa_count[5][32] , \sa_count[5].r.part1[0] );
tran (\sa_count[5][32] , \sa_count[5].f.upper[0] );
tran (\sa_count[5][33] , \sa_count[5].r.part1[1] );
tran (\sa_count[5][33] , \sa_count[5].f.upper[1] );
tran (\sa_count[5][34] , \sa_count[5].r.part1[2] );
tran (\sa_count[5][34] , \sa_count[5].f.upper[2] );
tran (\sa_count[5][35] , \sa_count[5].r.part1[3] );
tran (\sa_count[5][35] , \sa_count[5].f.upper[3] );
tran (\sa_count[5][36] , \sa_count[5].r.part1[4] );
tran (\sa_count[5][36] , \sa_count[5].f.upper[4] );
tran (\sa_count[5][37] , \sa_count[5].r.part1[5] );
tran (\sa_count[5][37] , \sa_count[5].f.upper[5] );
tran (\sa_count[5][38] , \sa_count[5].r.part1[6] );
tran (\sa_count[5][38] , \sa_count[5].f.upper[6] );
tran (\sa_count[5][39] , \sa_count[5].r.part1[7] );
tran (\sa_count[5][39] , \sa_count[5].f.upper[7] );
tran (\sa_count[5][40] , \sa_count[5].r.part1[8] );
tran (\sa_count[5][40] , \sa_count[5].f.upper[8] );
tran (\sa_count[5][41] , \sa_count[5].r.part1[9] );
tran (\sa_count[5][41] , \sa_count[5].f.upper[9] );
tran (\sa_count[5][42] , \sa_count[5].r.part1[10] );
tran (\sa_count[5][42] , \sa_count[5].f.upper[10] );
tran (\sa_count[5][43] , \sa_count[5].r.part1[11] );
tran (\sa_count[5][43] , \sa_count[5].f.upper[11] );
tran (\sa_count[5][44] , \sa_count[5].r.part1[12] );
tran (\sa_count[5][44] , \sa_count[5].f.upper[12] );
tran (\sa_count[5][45] , \sa_count[5].r.part1[13] );
tran (\sa_count[5][45] , \sa_count[5].f.upper[13] );
tran (\sa_count[5][46] , \sa_count[5].r.part1[14] );
tran (\sa_count[5][46] , \sa_count[5].f.upper[14] );
tran (\sa_count[5][47] , \sa_count[5].r.part1[15] );
tran (\sa_count[5][47] , \sa_count[5].f.upper[15] );
tran (\sa_count[5][48] , \sa_count[5].r.part1[16] );
tran (\sa_count[5][48] , \sa_count[5].f.upper[16] );
tran (\sa_count[5][49] , \sa_count[5].r.part1[17] );
tran (\sa_count[5][49] , \sa_count[5].f.upper[17] );
tran (\sa_count[5][50] , \sa_count[5].r.part1[18] );
tran (\sa_count[5][50] , \sa_count[5].f.unused[0] );
tran (\sa_count[5][51] , \sa_count[5].r.part1[19] );
tran (\sa_count[5][51] , \sa_count[5].f.unused[1] );
tran (\sa_count[5][52] , \sa_count[5].r.part1[20] );
tran (\sa_count[5][52] , \sa_count[5].f.unused[2] );
tran (\sa_count[5][53] , \sa_count[5].r.part1[21] );
tran (\sa_count[5][53] , \sa_count[5].f.unused[3] );
tran (\sa_count[5][54] , \sa_count[5].r.part1[22] );
tran (\sa_count[5][54] , \sa_count[5].f.unused[4] );
tran (\sa_count[5][55] , \sa_count[5].r.part1[23] );
tran (\sa_count[5][55] , \sa_count[5].f.unused[5] );
tran (\sa_count[5][56] , \sa_count[5].r.part1[24] );
tran (\sa_count[5][56] , \sa_count[5].f.unused[6] );
tran (\sa_count[5][57] , \sa_count[5].r.part1[25] );
tran (\sa_count[5][57] , \sa_count[5].f.unused[7] );
tran (\sa_count[5][58] , \sa_count[5].r.part1[26] );
tran (\sa_count[5][58] , \sa_count[5].f.unused[8] );
tran (\sa_count[5][59] , \sa_count[5].r.part1[27] );
tran (\sa_count[5][59] , \sa_count[5].f.unused[9] );
tran (\sa_count[5][60] , \sa_count[5].r.part1[28] );
tran (\sa_count[5][60] , \sa_count[5].f.unused[10] );
tran (\sa_count[5][61] , \sa_count[5].r.part1[29] );
tran (\sa_count[5][61] , \sa_count[5].f.unused[11] );
tran (\sa_count[5][62] , \sa_count[5].r.part1[30] );
tran (\sa_count[5][62] , \sa_count[5].f.unused[12] );
tran (\sa_count[5][63] , \sa_count[5].r.part1[31] );
tran (\sa_count[5][63] , \sa_count[5].f.unused[13] );
tran (\sa_count[6][0] , \sa_count[6].r.part0[0] );
tran (\sa_count[6][0] , \sa_count[6].f.lower[0] );
tran (\sa_count[6][1] , \sa_count[6].r.part0[1] );
tran (\sa_count[6][1] , \sa_count[6].f.lower[1] );
tran (\sa_count[6][2] , \sa_count[6].r.part0[2] );
tran (\sa_count[6][2] , \sa_count[6].f.lower[2] );
tran (\sa_count[6][3] , \sa_count[6].r.part0[3] );
tran (\sa_count[6][3] , \sa_count[6].f.lower[3] );
tran (\sa_count[6][4] , \sa_count[6].r.part0[4] );
tran (\sa_count[6][4] , \sa_count[6].f.lower[4] );
tran (\sa_count[6][5] , \sa_count[6].r.part0[5] );
tran (\sa_count[6][5] , \sa_count[6].f.lower[5] );
tran (\sa_count[6][6] , \sa_count[6].r.part0[6] );
tran (\sa_count[6][6] , \sa_count[6].f.lower[6] );
tran (\sa_count[6][7] , \sa_count[6].r.part0[7] );
tran (\sa_count[6][7] , \sa_count[6].f.lower[7] );
tran (\sa_count[6][8] , \sa_count[6].r.part0[8] );
tran (\sa_count[6][8] , \sa_count[6].f.lower[8] );
tran (\sa_count[6][9] , \sa_count[6].r.part0[9] );
tran (\sa_count[6][9] , \sa_count[6].f.lower[9] );
tran (\sa_count[6][10] , \sa_count[6].r.part0[10] );
tran (\sa_count[6][10] , \sa_count[6].f.lower[10] );
tran (\sa_count[6][11] , \sa_count[6].r.part0[11] );
tran (\sa_count[6][11] , \sa_count[6].f.lower[11] );
tran (\sa_count[6][12] , \sa_count[6].r.part0[12] );
tran (\sa_count[6][12] , \sa_count[6].f.lower[12] );
tran (\sa_count[6][13] , \sa_count[6].r.part0[13] );
tran (\sa_count[6][13] , \sa_count[6].f.lower[13] );
tran (\sa_count[6][14] , \sa_count[6].r.part0[14] );
tran (\sa_count[6][14] , \sa_count[6].f.lower[14] );
tran (\sa_count[6][15] , \sa_count[6].r.part0[15] );
tran (\sa_count[6][15] , \sa_count[6].f.lower[15] );
tran (\sa_count[6][16] , \sa_count[6].r.part0[16] );
tran (\sa_count[6][16] , \sa_count[6].f.lower[16] );
tran (\sa_count[6][17] , \sa_count[6].r.part0[17] );
tran (\sa_count[6][17] , \sa_count[6].f.lower[17] );
tran (\sa_count[6][18] , \sa_count[6].r.part0[18] );
tran (\sa_count[6][18] , \sa_count[6].f.lower[18] );
tran (\sa_count[6][19] , \sa_count[6].r.part0[19] );
tran (\sa_count[6][19] , \sa_count[6].f.lower[19] );
tran (\sa_count[6][20] , \sa_count[6].r.part0[20] );
tran (\sa_count[6][20] , \sa_count[6].f.lower[20] );
tran (\sa_count[6][21] , \sa_count[6].r.part0[21] );
tran (\sa_count[6][21] , \sa_count[6].f.lower[21] );
tran (\sa_count[6][22] , \sa_count[6].r.part0[22] );
tran (\sa_count[6][22] , \sa_count[6].f.lower[22] );
tran (\sa_count[6][23] , \sa_count[6].r.part0[23] );
tran (\sa_count[6][23] , \sa_count[6].f.lower[23] );
tran (\sa_count[6][24] , \sa_count[6].r.part0[24] );
tran (\sa_count[6][24] , \sa_count[6].f.lower[24] );
tran (\sa_count[6][25] , \sa_count[6].r.part0[25] );
tran (\sa_count[6][25] , \sa_count[6].f.lower[25] );
tran (\sa_count[6][26] , \sa_count[6].r.part0[26] );
tran (\sa_count[6][26] , \sa_count[6].f.lower[26] );
tran (\sa_count[6][27] , \sa_count[6].r.part0[27] );
tran (\sa_count[6][27] , \sa_count[6].f.lower[27] );
tran (\sa_count[6][28] , \sa_count[6].r.part0[28] );
tran (\sa_count[6][28] , \sa_count[6].f.lower[28] );
tran (\sa_count[6][29] , \sa_count[6].r.part0[29] );
tran (\sa_count[6][29] , \sa_count[6].f.lower[29] );
tran (\sa_count[6][30] , \sa_count[6].r.part0[30] );
tran (\sa_count[6][30] , \sa_count[6].f.lower[30] );
tran (\sa_count[6][31] , \sa_count[6].r.part0[31] );
tran (\sa_count[6][31] , \sa_count[6].f.lower[31] );
tran (\sa_count[6][32] , \sa_count[6].r.part1[0] );
tran (\sa_count[6][32] , \sa_count[6].f.upper[0] );
tran (\sa_count[6][33] , \sa_count[6].r.part1[1] );
tran (\sa_count[6][33] , \sa_count[6].f.upper[1] );
tran (\sa_count[6][34] , \sa_count[6].r.part1[2] );
tran (\sa_count[6][34] , \sa_count[6].f.upper[2] );
tran (\sa_count[6][35] , \sa_count[6].r.part1[3] );
tran (\sa_count[6][35] , \sa_count[6].f.upper[3] );
tran (\sa_count[6][36] , \sa_count[6].r.part1[4] );
tran (\sa_count[6][36] , \sa_count[6].f.upper[4] );
tran (\sa_count[6][37] , \sa_count[6].r.part1[5] );
tran (\sa_count[6][37] , \sa_count[6].f.upper[5] );
tran (\sa_count[6][38] , \sa_count[6].r.part1[6] );
tran (\sa_count[6][38] , \sa_count[6].f.upper[6] );
tran (\sa_count[6][39] , \sa_count[6].r.part1[7] );
tran (\sa_count[6][39] , \sa_count[6].f.upper[7] );
tran (\sa_count[6][40] , \sa_count[6].r.part1[8] );
tran (\sa_count[6][40] , \sa_count[6].f.upper[8] );
tran (\sa_count[6][41] , \sa_count[6].r.part1[9] );
tran (\sa_count[6][41] , \sa_count[6].f.upper[9] );
tran (\sa_count[6][42] , \sa_count[6].r.part1[10] );
tran (\sa_count[6][42] , \sa_count[6].f.upper[10] );
tran (\sa_count[6][43] , \sa_count[6].r.part1[11] );
tran (\sa_count[6][43] , \sa_count[6].f.upper[11] );
tran (\sa_count[6][44] , \sa_count[6].r.part1[12] );
tran (\sa_count[6][44] , \sa_count[6].f.upper[12] );
tran (\sa_count[6][45] , \sa_count[6].r.part1[13] );
tran (\sa_count[6][45] , \sa_count[6].f.upper[13] );
tran (\sa_count[6][46] , \sa_count[6].r.part1[14] );
tran (\sa_count[6][46] , \sa_count[6].f.upper[14] );
tran (\sa_count[6][47] , \sa_count[6].r.part1[15] );
tran (\sa_count[6][47] , \sa_count[6].f.upper[15] );
tran (\sa_count[6][48] , \sa_count[6].r.part1[16] );
tran (\sa_count[6][48] , \sa_count[6].f.upper[16] );
tran (\sa_count[6][49] , \sa_count[6].r.part1[17] );
tran (\sa_count[6][49] , \sa_count[6].f.upper[17] );
tran (\sa_count[6][50] , \sa_count[6].r.part1[18] );
tran (\sa_count[6][50] , \sa_count[6].f.unused[0] );
tran (\sa_count[6][51] , \sa_count[6].r.part1[19] );
tran (\sa_count[6][51] , \sa_count[6].f.unused[1] );
tran (\sa_count[6][52] , \sa_count[6].r.part1[20] );
tran (\sa_count[6][52] , \sa_count[6].f.unused[2] );
tran (\sa_count[6][53] , \sa_count[6].r.part1[21] );
tran (\sa_count[6][53] , \sa_count[6].f.unused[3] );
tran (\sa_count[6][54] , \sa_count[6].r.part1[22] );
tran (\sa_count[6][54] , \sa_count[6].f.unused[4] );
tran (\sa_count[6][55] , \sa_count[6].r.part1[23] );
tran (\sa_count[6][55] , \sa_count[6].f.unused[5] );
tran (\sa_count[6][56] , \sa_count[6].r.part1[24] );
tran (\sa_count[6][56] , \sa_count[6].f.unused[6] );
tran (\sa_count[6][57] , \sa_count[6].r.part1[25] );
tran (\sa_count[6][57] , \sa_count[6].f.unused[7] );
tran (\sa_count[6][58] , \sa_count[6].r.part1[26] );
tran (\sa_count[6][58] , \sa_count[6].f.unused[8] );
tran (\sa_count[6][59] , \sa_count[6].r.part1[27] );
tran (\sa_count[6][59] , \sa_count[6].f.unused[9] );
tran (\sa_count[6][60] , \sa_count[6].r.part1[28] );
tran (\sa_count[6][60] , \sa_count[6].f.unused[10] );
tran (\sa_count[6][61] , \sa_count[6].r.part1[29] );
tran (\sa_count[6][61] , \sa_count[6].f.unused[11] );
tran (\sa_count[6][62] , \sa_count[6].r.part1[30] );
tran (\sa_count[6][62] , \sa_count[6].f.unused[12] );
tran (\sa_count[6][63] , \sa_count[6].r.part1[31] );
tran (\sa_count[6][63] , \sa_count[6].f.unused[13] );
tran (\sa_count[7][0] , \sa_count[7].r.part0[0] );
tran (\sa_count[7][0] , \sa_count[7].f.lower[0] );
tran (\sa_count[7][1] , \sa_count[7].r.part0[1] );
tran (\sa_count[7][1] , \sa_count[7].f.lower[1] );
tran (\sa_count[7][2] , \sa_count[7].r.part0[2] );
tran (\sa_count[7][2] , \sa_count[7].f.lower[2] );
tran (\sa_count[7][3] , \sa_count[7].r.part0[3] );
tran (\sa_count[7][3] , \sa_count[7].f.lower[3] );
tran (\sa_count[7][4] , \sa_count[7].r.part0[4] );
tran (\sa_count[7][4] , \sa_count[7].f.lower[4] );
tran (\sa_count[7][5] , \sa_count[7].r.part0[5] );
tran (\sa_count[7][5] , \sa_count[7].f.lower[5] );
tran (\sa_count[7][6] , \sa_count[7].r.part0[6] );
tran (\sa_count[7][6] , \sa_count[7].f.lower[6] );
tran (\sa_count[7][7] , \sa_count[7].r.part0[7] );
tran (\sa_count[7][7] , \sa_count[7].f.lower[7] );
tran (\sa_count[7][8] , \sa_count[7].r.part0[8] );
tran (\sa_count[7][8] , \sa_count[7].f.lower[8] );
tran (\sa_count[7][9] , \sa_count[7].r.part0[9] );
tran (\sa_count[7][9] , \sa_count[7].f.lower[9] );
tran (\sa_count[7][10] , \sa_count[7].r.part0[10] );
tran (\sa_count[7][10] , \sa_count[7].f.lower[10] );
tran (\sa_count[7][11] , \sa_count[7].r.part0[11] );
tran (\sa_count[7][11] , \sa_count[7].f.lower[11] );
tran (\sa_count[7][12] , \sa_count[7].r.part0[12] );
tran (\sa_count[7][12] , \sa_count[7].f.lower[12] );
tran (\sa_count[7][13] , \sa_count[7].r.part0[13] );
tran (\sa_count[7][13] , \sa_count[7].f.lower[13] );
tran (\sa_count[7][14] , \sa_count[7].r.part0[14] );
tran (\sa_count[7][14] , \sa_count[7].f.lower[14] );
tran (\sa_count[7][15] , \sa_count[7].r.part0[15] );
tran (\sa_count[7][15] , \sa_count[7].f.lower[15] );
tran (\sa_count[7][16] , \sa_count[7].r.part0[16] );
tran (\sa_count[7][16] , \sa_count[7].f.lower[16] );
tran (\sa_count[7][17] , \sa_count[7].r.part0[17] );
tran (\sa_count[7][17] , \sa_count[7].f.lower[17] );
tran (\sa_count[7][18] , \sa_count[7].r.part0[18] );
tran (\sa_count[7][18] , \sa_count[7].f.lower[18] );
tran (\sa_count[7][19] , \sa_count[7].r.part0[19] );
tran (\sa_count[7][19] , \sa_count[7].f.lower[19] );
tran (\sa_count[7][20] , \sa_count[7].r.part0[20] );
tran (\sa_count[7][20] , \sa_count[7].f.lower[20] );
tran (\sa_count[7][21] , \sa_count[7].r.part0[21] );
tran (\sa_count[7][21] , \sa_count[7].f.lower[21] );
tran (\sa_count[7][22] , \sa_count[7].r.part0[22] );
tran (\sa_count[7][22] , \sa_count[7].f.lower[22] );
tran (\sa_count[7][23] , \sa_count[7].r.part0[23] );
tran (\sa_count[7][23] , \sa_count[7].f.lower[23] );
tran (\sa_count[7][24] , \sa_count[7].r.part0[24] );
tran (\sa_count[7][24] , \sa_count[7].f.lower[24] );
tran (\sa_count[7][25] , \sa_count[7].r.part0[25] );
tran (\sa_count[7][25] , \sa_count[7].f.lower[25] );
tran (\sa_count[7][26] , \sa_count[7].r.part0[26] );
tran (\sa_count[7][26] , \sa_count[7].f.lower[26] );
tran (\sa_count[7][27] , \sa_count[7].r.part0[27] );
tran (\sa_count[7][27] , \sa_count[7].f.lower[27] );
tran (\sa_count[7][28] , \sa_count[7].r.part0[28] );
tran (\sa_count[7][28] , \sa_count[7].f.lower[28] );
tran (\sa_count[7][29] , \sa_count[7].r.part0[29] );
tran (\sa_count[7][29] , \sa_count[7].f.lower[29] );
tran (\sa_count[7][30] , \sa_count[7].r.part0[30] );
tran (\sa_count[7][30] , \sa_count[7].f.lower[30] );
tran (\sa_count[7][31] , \sa_count[7].r.part0[31] );
tran (\sa_count[7][31] , \sa_count[7].f.lower[31] );
tran (\sa_count[7][32] , \sa_count[7].r.part1[0] );
tran (\sa_count[7][32] , \sa_count[7].f.upper[0] );
tran (\sa_count[7][33] , \sa_count[7].r.part1[1] );
tran (\sa_count[7][33] , \sa_count[7].f.upper[1] );
tran (\sa_count[7][34] , \sa_count[7].r.part1[2] );
tran (\sa_count[7][34] , \sa_count[7].f.upper[2] );
tran (\sa_count[7][35] , \sa_count[7].r.part1[3] );
tran (\sa_count[7][35] , \sa_count[7].f.upper[3] );
tran (\sa_count[7][36] , \sa_count[7].r.part1[4] );
tran (\sa_count[7][36] , \sa_count[7].f.upper[4] );
tran (\sa_count[7][37] , \sa_count[7].r.part1[5] );
tran (\sa_count[7][37] , \sa_count[7].f.upper[5] );
tran (\sa_count[7][38] , \sa_count[7].r.part1[6] );
tran (\sa_count[7][38] , \sa_count[7].f.upper[6] );
tran (\sa_count[7][39] , \sa_count[7].r.part1[7] );
tran (\sa_count[7][39] , \sa_count[7].f.upper[7] );
tran (\sa_count[7][40] , \sa_count[7].r.part1[8] );
tran (\sa_count[7][40] , \sa_count[7].f.upper[8] );
tran (\sa_count[7][41] , \sa_count[7].r.part1[9] );
tran (\sa_count[7][41] , \sa_count[7].f.upper[9] );
tran (\sa_count[7][42] , \sa_count[7].r.part1[10] );
tran (\sa_count[7][42] , \sa_count[7].f.upper[10] );
tran (\sa_count[7][43] , \sa_count[7].r.part1[11] );
tran (\sa_count[7][43] , \sa_count[7].f.upper[11] );
tran (\sa_count[7][44] , \sa_count[7].r.part1[12] );
tran (\sa_count[7][44] , \sa_count[7].f.upper[12] );
tran (\sa_count[7][45] , \sa_count[7].r.part1[13] );
tran (\sa_count[7][45] , \sa_count[7].f.upper[13] );
tran (\sa_count[7][46] , \sa_count[7].r.part1[14] );
tran (\sa_count[7][46] , \sa_count[7].f.upper[14] );
tran (\sa_count[7][47] , \sa_count[7].r.part1[15] );
tran (\sa_count[7][47] , \sa_count[7].f.upper[15] );
tran (\sa_count[7][48] , \sa_count[7].r.part1[16] );
tran (\sa_count[7][48] , \sa_count[7].f.upper[16] );
tran (\sa_count[7][49] , \sa_count[7].r.part1[17] );
tran (\sa_count[7][49] , \sa_count[7].f.upper[17] );
tran (\sa_count[7][50] , \sa_count[7].r.part1[18] );
tran (\sa_count[7][50] , \sa_count[7].f.unused[0] );
tran (\sa_count[7][51] , \sa_count[7].r.part1[19] );
tran (\sa_count[7][51] , \sa_count[7].f.unused[1] );
tran (\sa_count[7][52] , \sa_count[7].r.part1[20] );
tran (\sa_count[7][52] , \sa_count[7].f.unused[2] );
tran (\sa_count[7][53] , \sa_count[7].r.part1[21] );
tran (\sa_count[7][53] , \sa_count[7].f.unused[3] );
tran (\sa_count[7][54] , \sa_count[7].r.part1[22] );
tran (\sa_count[7][54] , \sa_count[7].f.unused[4] );
tran (\sa_count[7][55] , \sa_count[7].r.part1[23] );
tran (\sa_count[7][55] , \sa_count[7].f.unused[5] );
tran (\sa_count[7][56] , \sa_count[7].r.part1[24] );
tran (\sa_count[7][56] , \sa_count[7].f.unused[6] );
tran (\sa_count[7][57] , \sa_count[7].r.part1[25] );
tran (\sa_count[7][57] , \sa_count[7].f.unused[7] );
tran (\sa_count[7][58] , \sa_count[7].r.part1[26] );
tran (\sa_count[7][58] , \sa_count[7].f.unused[8] );
tran (\sa_count[7][59] , \sa_count[7].r.part1[27] );
tran (\sa_count[7][59] , \sa_count[7].f.unused[9] );
tran (\sa_count[7][60] , \sa_count[7].r.part1[28] );
tran (\sa_count[7][60] , \sa_count[7].f.unused[10] );
tran (\sa_count[7][61] , \sa_count[7].r.part1[29] );
tran (\sa_count[7][61] , \sa_count[7].f.unused[11] );
tran (\sa_count[7][62] , \sa_count[7].r.part1[30] );
tran (\sa_count[7][62] , \sa_count[7].f.unused[12] );
tran (\sa_count[7][63] , \sa_count[7].r.part1[31] );
tran (\sa_count[7][63] , \sa_count[7].f.unused[13] );
tran (\sa_count[8][0] , \sa_count[8].r.part0[0] );
tran (\sa_count[8][0] , \sa_count[8].f.lower[0] );
tran (\sa_count[8][1] , \sa_count[8].r.part0[1] );
tran (\sa_count[8][1] , \sa_count[8].f.lower[1] );
tran (\sa_count[8][2] , \sa_count[8].r.part0[2] );
tran (\sa_count[8][2] , \sa_count[8].f.lower[2] );
tran (\sa_count[8][3] , \sa_count[8].r.part0[3] );
tran (\sa_count[8][3] , \sa_count[8].f.lower[3] );
tran (\sa_count[8][4] , \sa_count[8].r.part0[4] );
tran (\sa_count[8][4] , \sa_count[8].f.lower[4] );
tran (\sa_count[8][5] , \sa_count[8].r.part0[5] );
tran (\sa_count[8][5] , \sa_count[8].f.lower[5] );
tran (\sa_count[8][6] , \sa_count[8].r.part0[6] );
tran (\sa_count[8][6] , \sa_count[8].f.lower[6] );
tran (\sa_count[8][7] , \sa_count[8].r.part0[7] );
tran (\sa_count[8][7] , \sa_count[8].f.lower[7] );
tran (\sa_count[8][8] , \sa_count[8].r.part0[8] );
tran (\sa_count[8][8] , \sa_count[8].f.lower[8] );
tran (\sa_count[8][9] , \sa_count[8].r.part0[9] );
tran (\sa_count[8][9] , \sa_count[8].f.lower[9] );
tran (\sa_count[8][10] , \sa_count[8].r.part0[10] );
tran (\sa_count[8][10] , \sa_count[8].f.lower[10] );
tran (\sa_count[8][11] , \sa_count[8].r.part0[11] );
tran (\sa_count[8][11] , \sa_count[8].f.lower[11] );
tran (\sa_count[8][12] , \sa_count[8].r.part0[12] );
tran (\sa_count[8][12] , \sa_count[8].f.lower[12] );
tran (\sa_count[8][13] , \sa_count[8].r.part0[13] );
tran (\sa_count[8][13] , \sa_count[8].f.lower[13] );
tran (\sa_count[8][14] , \sa_count[8].r.part0[14] );
tran (\sa_count[8][14] , \sa_count[8].f.lower[14] );
tran (\sa_count[8][15] , \sa_count[8].r.part0[15] );
tran (\sa_count[8][15] , \sa_count[8].f.lower[15] );
tran (\sa_count[8][16] , \sa_count[8].r.part0[16] );
tran (\sa_count[8][16] , \sa_count[8].f.lower[16] );
tran (\sa_count[8][17] , \sa_count[8].r.part0[17] );
tran (\sa_count[8][17] , \sa_count[8].f.lower[17] );
tran (\sa_count[8][18] , \sa_count[8].r.part0[18] );
tran (\sa_count[8][18] , \sa_count[8].f.lower[18] );
tran (\sa_count[8][19] , \sa_count[8].r.part0[19] );
tran (\sa_count[8][19] , \sa_count[8].f.lower[19] );
tran (\sa_count[8][20] , \sa_count[8].r.part0[20] );
tran (\sa_count[8][20] , \sa_count[8].f.lower[20] );
tran (\sa_count[8][21] , \sa_count[8].r.part0[21] );
tran (\sa_count[8][21] , \sa_count[8].f.lower[21] );
tran (\sa_count[8][22] , \sa_count[8].r.part0[22] );
tran (\sa_count[8][22] , \sa_count[8].f.lower[22] );
tran (\sa_count[8][23] , \sa_count[8].r.part0[23] );
tran (\sa_count[8][23] , \sa_count[8].f.lower[23] );
tran (\sa_count[8][24] , \sa_count[8].r.part0[24] );
tran (\sa_count[8][24] , \sa_count[8].f.lower[24] );
tran (\sa_count[8][25] , \sa_count[8].r.part0[25] );
tran (\sa_count[8][25] , \sa_count[8].f.lower[25] );
tran (\sa_count[8][26] , \sa_count[8].r.part0[26] );
tran (\sa_count[8][26] , \sa_count[8].f.lower[26] );
tran (\sa_count[8][27] , \sa_count[8].r.part0[27] );
tran (\sa_count[8][27] , \sa_count[8].f.lower[27] );
tran (\sa_count[8][28] , \sa_count[8].r.part0[28] );
tran (\sa_count[8][28] , \sa_count[8].f.lower[28] );
tran (\sa_count[8][29] , \sa_count[8].r.part0[29] );
tran (\sa_count[8][29] , \sa_count[8].f.lower[29] );
tran (\sa_count[8][30] , \sa_count[8].r.part0[30] );
tran (\sa_count[8][30] , \sa_count[8].f.lower[30] );
tran (\sa_count[8][31] , \sa_count[8].r.part0[31] );
tran (\sa_count[8][31] , \sa_count[8].f.lower[31] );
tran (\sa_count[8][32] , \sa_count[8].r.part1[0] );
tran (\sa_count[8][32] , \sa_count[8].f.upper[0] );
tran (\sa_count[8][33] , \sa_count[8].r.part1[1] );
tran (\sa_count[8][33] , \sa_count[8].f.upper[1] );
tran (\sa_count[8][34] , \sa_count[8].r.part1[2] );
tran (\sa_count[8][34] , \sa_count[8].f.upper[2] );
tran (\sa_count[8][35] , \sa_count[8].r.part1[3] );
tran (\sa_count[8][35] , \sa_count[8].f.upper[3] );
tran (\sa_count[8][36] , \sa_count[8].r.part1[4] );
tran (\sa_count[8][36] , \sa_count[8].f.upper[4] );
tran (\sa_count[8][37] , \sa_count[8].r.part1[5] );
tran (\sa_count[8][37] , \sa_count[8].f.upper[5] );
tran (\sa_count[8][38] , \sa_count[8].r.part1[6] );
tran (\sa_count[8][38] , \sa_count[8].f.upper[6] );
tran (\sa_count[8][39] , \sa_count[8].r.part1[7] );
tran (\sa_count[8][39] , \sa_count[8].f.upper[7] );
tran (\sa_count[8][40] , \sa_count[8].r.part1[8] );
tran (\sa_count[8][40] , \sa_count[8].f.upper[8] );
tran (\sa_count[8][41] , \sa_count[8].r.part1[9] );
tran (\sa_count[8][41] , \sa_count[8].f.upper[9] );
tran (\sa_count[8][42] , \sa_count[8].r.part1[10] );
tran (\sa_count[8][42] , \sa_count[8].f.upper[10] );
tran (\sa_count[8][43] , \sa_count[8].r.part1[11] );
tran (\sa_count[8][43] , \sa_count[8].f.upper[11] );
tran (\sa_count[8][44] , \sa_count[8].r.part1[12] );
tran (\sa_count[8][44] , \sa_count[8].f.upper[12] );
tran (\sa_count[8][45] , \sa_count[8].r.part1[13] );
tran (\sa_count[8][45] , \sa_count[8].f.upper[13] );
tran (\sa_count[8][46] , \sa_count[8].r.part1[14] );
tran (\sa_count[8][46] , \sa_count[8].f.upper[14] );
tran (\sa_count[8][47] , \sa_count[8].r.part1[15] );
tran (\sa_count[8][47] , \sa_count[8].f.upper[15] );
tran (\sa_count[8][48] , \sa_count[8].r.part1[16] );
tran (\sa_count[8][48] , \sa_count[8].f.upper[16] );
tran (\sa_count[8][49] , \sa_count[8].r.part1[17] );
tran (\sa_count[8][49] , \sa_count[8].f.upper[17] );
tran (\sa_count[8][50] , \sa_count[8].r.part1[18] );
tran (\sa_count[8][50] , \sa_count[8].f.unused[0] );
tran (\sa_count[8][51] , \sa_count[8].r.part1[19] );
tran (\sa_count[8][51] , \sa_count[8].f.unused[1] );
tran (\sa_count[8][52] , \sa_count[8].r.part1[20] );
tran (\sa_count[8][52] , \sa_count[8].f.unused[2] );
tran (\sa_count[8][53] , \sa_count[8].r.part1[21] );
tran (\sa_count[8][53] , \sa_count[8].f.unused[3] );
tran (\sa_count[8][54] , \sa_count[8].r.part1[22] );
tran (\sa_count[8][54] , \sa_count[8].f.unused[4] );
tran (\sa_count[8][55] , \sa_count[8].r.part1[23] );
tran (\sa_count[8][55] , \sa_count[8].f.unused[5] );
tran (\sa_count[8][56] , \sa_count[8].r.part1[24] );
tran (\sa_count[8][56] , \sa_count[8].f.unused[6] );
tran (\sa_count[8][57] , \sa_count[8].r.part1[25] );
tran (\sa_count[8][57] , \sa_count[8].f.unused[7] );
tran (\sa_count[8][58] , \sa_count[8].r.part1[26] );
tran (\sa_count[8][58] , \sa_count[8].f.unused[8] );
tran (\sa_count[8][59] , \sa_count[8].r.part1[27] );
tran (\sa_count[8][59] , \sa_count[8].f.unused[9] );
tran (\sa_count[8][60] , \sa_count[8].r.part1[28] );
tran (\sa_count[8][60] , \sa_count[8].f.unused[10] );
tran (\sa_count[8][61] , \sa_count[8].r.part1[29] );
tran (\sa_count[8][61] , \sa_count[8].f.unused[11] );
tran (\sa_count[8][62] , \sa_count[8].r.part1[30] );
tran (\sa_count[8][62] , \sa_count[8].f.unused[12] );
tran (\sa_count[8][63] , \sa_count[8].r.part1[31] );
tran (\sa_count[8][63] , \sa_count[8].f.unused[13] );
tran (\sa_count[9][0] , \sa_count[9].r.part0[0] );
tran (\sa_count[9][0] , \sa_count[9].f.lower[0] );
tran (\sa_count[9][1] , \sa_count[9].r.part0[1] );
tran (\sa_count[9][1] , \sa_count[9].f.lower[1] );
tran (\sa_count[9][2] , \sa_count[9].r.part0[2] );
tran (\sa_count[9][2] , \sa_count[9].f.lower[2] );
tran (\sa_count[9][3] , \sa_count[9].r.part0[3] );
tran (\sa_count[9][3] , \sa_count[9].f.lower[3] );
tran (\sa_count[9][4] , \sa_count[9].r.part0[4] );
tran (\sa_count[9][4] , \sa_count[9].f.lower[4] );
tran (\sa_count[9][5] , \sa_count[9].r.part0[5] );
tran (\sa_count[9][5] , \sa_count[9].f.lower[5] );
tran (\sa_count[9][6] , \sa_count[9].r.part0[6] );
tran (\sa_count[9][6] , \sa_count[9].f.lower[6] );
tran (\sa_count[9][7] , \sa_count[9].r.part0[7] );
tran (\sa_count[9][7] , \sa_count[9].f.lower[7] );
tran (\sa_count[9][8] , \sa_count[9].r.part0[8] );
tran (\sa_count[9][8] , \sa_count[9].f.lower[8] );
tran (\sa_count[9][9] , \sa_count[9].r.part0[9] );
tran (\sa_count[9][9] , \sa_count[9].f.lower[9] );
tran (\sa_count[9][10] , \sa_count[9].r.part0[10] );
tran (\sa_count[9][10] , \sa_count[9].f.lower[10] );
tran (\sa_count[9][11] , \sa_count[9].r.part0[11] );
tran (\sa_count[9][11] , \sa_count[9].f.lower[11] );
tran (\sa_count[9][12] , \sa_count[9].r.part0[12] );
tran (\sa_count[9][12] , \sa_count[9].f.lower[12] );
tran (\sa_count[9][13] , \sa_count[9].r.part0[13] );
tran (\sa_count[9][13] , \sa_count[9].f.lower[13] );
tran (\sa_count[9][14] , \sa_count[9].r.part0[14] );
tran (\sa_count[9][14] , \sa_count[9].f.lower[14] );
tran (\sa_count[9][15] , \sa_count[9].r.part0[15] );
tran (\sa_count[9][15] , \sa_count[9].f.lower[15] );
tran (\sa_count[9][16] , \sa_count[9].r.part0[16] );
tran (\sa_count[9][16] , \sa_count[9].f.lower[16] );
tran (\sa_count[9][17] , \sa_count[9].r.part0[17] );
tran (\sa_count[9][17] , \sa_count[9].f.lower[17] );
tran (\sa_count[9][18] , \sa_count[9].r.part0[18] );
tran (\sa_count[9][18] , \sa_count[9].f.lower[18] );
tran (\sa_count[9][19] , \sa_count[9].r.part0[19] );
tran (\sa_count[9][19] , \sa_count[9].f.lower[19] );
tran (\sa_count[9][20] , \sa_count[9].r.part0[20] );
tran (\sa_count[9][20] , \sa_count[9].f.lower[20] );
tran (\sa_count[9][21] , \sa_count[9].r.part0[21] );
tran (\sa_count[9][21] , \sa_count[9].f.lower[21] );
tran (\sa_count[9][22] , \sa_count[9].r.part0[22] );
tran (\sa_count[9][22] , \sa_count[9].f.lower[22] );
tran (\sa_count[9][23] , \sa_count[9].r.part0[23] );
tran (\sa_count[9][23] , \sa_count[9].f.lower[23] );
tran (\sa_count[9][24] , \sa_count[9].r.part0[24] );
tran (\sa_count[9][24] , \sa_count[9].f.lower[24] );
tran (\sa_count[9][25] , \sa_count[9].r.part0[25] );
tran (\sa_count[9][25] , \sa_count[9].f.lower[25] );
tran (\sa_count[9][26] , \sa_count[9].r.part0[26] );
tran (\sa_count[9][26] , \sa_count[9].f.lower[26] );
tran (\sa_count[9][27] , \sa_count[9].r.part0[27] );
tran (\sa_count[9][27] , \sa_count[9].f.lower[27] );
tran (\sa_count[9][28] , \sa_count[9].r.part0[28] );
tran (\sa_count[9][28] , \sa_count[9].f.lower[28] );
tran (\sa_count[9][29] , \sa_count[9].r.part0[29] );
tran (\sa_count[9][29] , \sa_count[9].f.lower[29] );
tran (\sa_count[9][30] , \sa_count[9].r.part0[30] );
tran (\sa_count[9][30] , \sa_count[9].f.lower[30] );
tran (\sa_count[9][31] , \sa_count[9].r.part0[31] );
tran (\sa_count[9][31] , \sa_count[9].f.lower[31] );
tran (\sa_count[9][32] , \sa_count[9].r.part1[0] );
tran (\sa_count[9][32] , \sa_count[9].f.upper[0] );
tran (\sa_count[9][33] , \sa_count[9].r.part1[1] );
tran (\sa_count[9][33] , \sa_count[9].f.upper[1] );
tran (\sa_count[9][34] , \sa_count[9].r.part1[2] );
tran (\sa_count[9][34] , \sa_count[9].f.upper[2] );
tran (\sa_count[9][35] , \sa_count[9].r.part1[3] );
tran (\sa_count[9][35] , \sa_count[9].f.upper[3] );
tran (\sa_count[9][36] , \sa_count[9].r.part1[4] );
tran (\sa_count[9][36] , \sa_count[9].f.upper[4] );
tran (\sa_count[9][37] , \sa_count[9].r.part1[5] );
tran (\sa_count[9][37] , \sa_count[9].f.upper[5] );
tran (\sa_count[9][38] , \sa_count[9].r.part1[6] );
tran (\sa_count[9][38] , \sa_count[9].f.upper[6] );
tran (\sa_count[9][39] , \sa_count[9].r.part1[7] );
tran (\sa_count[9][39] , \sa_count[9].f.upper[7] );
tran (\sa_count[9][40] , \sa_count[9].r.part1[8] );
tran (\sa_count[9][40] , \sa_count[9].f.upper[8] );
tran (\sa_count[9][41] , \sa_count[9].r.part1[9] );
tran (\sa_count[9][41] , \sa_count[9].f.upper[9] );
tran (\sa_count[9][42] , \sa_count[9].r.part1[10] );
tran (\sa_count[9][42] , \sa_count[9].f.upper[10] );
tran (\sa_count[9][43] , \sa_count[9].r.part1[11] );
tran (\sa_count[9][43] , \sa_count[9].f.upper[11] );
tran (\sa_count[9][44] , \sa_count[9].r.part1[12] );
tran (\sa_count[9][44] , \sa_count[9].f.upper[12] );
tran (\sa_count[9][45] , \sa_count[9].r.part1[13] );
tran (\sa_count[9][45] , \sa_count[9].f.upper[13] );
tran (\sa_count[9][46] , \sa_count[9].r.part1[14] );
tran (\sa_count[9][46] , \sa_count[9].f.upper[14] );
tran (\sa_count[9][47] , \sa_count[9].r.part1[15] );
tran (\sa_count[9][47] , \sa_count[9].f.upper[15] );
tran (\sa_count[9][48] , \sa_count[9].r.part1[16] );
tran (\sa_count[9][48] , \sa_count[9].f.upper[16] );
tran (\sa_count[9][49] , \sa_count[9].r.part1[17] );
tran (\sa_count[9][49] , \sa_count[9].f.upper[17] );
tran (\sa_count[9][50] , \sa_count[9].r.part1[18] );
tran (\sa_count[9][50] , \sa_count[9].f.unused[0] );
tran (\sa_count[9][51] , \sa_count[9].r.part1[19] );
tran (\sa_count[9][51] , \sa_count[9].f.unused[1] );
tran (\sa_count[9][52] , \sa_count[9].r.part1[20] );
tran (\sa_count[9][52] , \sa_count[9].f.unused[2] );
tran (\sa_count[9][53] , \sa_count[9].r.part1[21] );
tran (\sa_count[9][53] , \sa_count[9].f.unused[3] );
tran (\sa_count[9][54] , \sa_count[9].r.part1[22] );
tran (\sa_count[9][54] , \sa_count[9].f.unused[4] );
tran (\sa_count[9][55] , \sa_count[9].r.part1[23] );
tran (\sa_count[9][55] , \sa_count[9].f.unused[5] );
tran (\sa_count[9][56] , \sa_count[9].r.part1[24] );
tran (\sa_count[9][56] , \sa_count[9].f.unused[6] );
tran (\sa_count[9][57] , \sa_count[9].r.part1[25] );
tran (\sa_count[9][57] , \sa_count[9].f.unused[7] );
tran (\sa_count[9][58] , \sa_count[9].r.part1[26] );
tran (\sa_count[9][58] , \sa_count[9].f.unused[8] );
tran (\sa_count[9][59] , \sa_count[9].r.part1[27] );
tran (\sa_count[9][59] , \sa_count[9].f.unused[9] );
tran (\sa_count[9][60] , \sa_count[9].r.part1[28] );
tran (\sa_count[9][60] , \sa_count[9].f.unused[10] );
tran (\sa_count[9][61] , \sa_count[9].r.part1[29] );
tran (\sa_count[9][61] , \sa_count[9].f.unused[11] );
tran (\sa_count[9][62] , \sa_count[9].r.part1[30] );
tran (\sa_count[9][62] , \sa_count[9].f.unused[12] );
tran (\sa_count[9][63] , \sa_count[9].r.part1[31] );
tran (\sa_count[9][63] , \sa_count[9].f.unused[13] );
tran (\sa_count[10][0] , \sa_count[10].r.part0[0] );
tran (\sa_count[10][0] , \sa_count[10].f.lower[0] );
tran (\sa_count[10][1] , \sa_count[10].r.part0[1] );
tran (\sa_count[10][1] , \sa_count[10].f.lower[1] );
tran (\sa_count[10][2] , \sa_count[10].r.part0[2] );
tran (\sa_count[10][2] , \sa_count[10].f.lower[2] );
tran (\sa_count[10][3] , \sa_count[10].r.part0[3] );
tran (\sa_count[10][3] , \sa_count[10].f.lower[3] );
tran (\sa_count[10][4] , \sa_count[10].r.part0[4] );
tran (\sa_count[10][4] , \sa_count[10].f.lower[4] );
tran (\sa_count[10][5] , \sa_count[10].r.part0[5] );
tran (\sa_count[10][5] , \sa_count[10].f.lower[5] );
tran (\sa_count[10][6] , \sa_count[10].r.part0[6] );
tran (\sa_count[10][6] , \sa_count[10].f.lower[6] );
tran (\sa_count[10][7] , \sa_count[10].r.part0[7] );
tran (\sa_count[10][7] , \sa_count[10].f.lower[7] );
tran (\sa_count[10][8] , \sa_count[10].r.part0[8] );
tran (\sa_count[10][8] , \sa_count[10].f.lower[8] );
tran (\sa_count[10][9] , \sa_count[10].r.part0[9] );
tran (\sa_count[10][9] , \sa_count[10].f.lower[9] );
tran (\sa_count[10][10] , \sa_count[10].r.part0[10] );
tran (\sa_count[10][10] , \sa_count[10].f.lower[10] );
tran (\sa_count[10][11] , \sa_count[10].r.part0[11] );
tran (\sa_count[10][11] , \sa_count[10].f.lower[11] );
tran (\sa_count[10][12] , \sa_count[10].r.part0[12] );
tran (\sa_count[10][12] , \sa_count[10].f.lower[12] );
tran (\sa_count[10][13] , \sa_count[10].r.part0[13] );
tran (\sa_count[10][13] , \sa_count[10].f.lower[13] );
tran (\sa_count[10][14] , \sa_count[10].r.part0[14] );
tran (\sa_count[10][14] , \sa_count[10].f.lower[14] );
tran (\sa_count[10][15] , \sa_count[10].r.part0[15] );
tran (\sa_count[10][15] , \sa_count[10].f.lower[15] );
tran (\sa_count[10][16] , \sa_count[10].r.part0[16] );
tran (\sa_count[10][16] , \sa_count[10].f.lower[16] );
tran (\sa_count[10][17] , \sa_count[10].r.part0[17] );
tran (\sa_count[10][17] , \sa_count[10].f.lower[17] );
tran (\sa_count[10][18] , \sa_count[10].r.part0[18] );
tran (\sa_count[10][18] , \sa_count[10].f.lower[18] );
tran (\sa_count[10][19] , \sa_count[10].r.part0[19] );
tran (\sa_count[10][19] , \sa_count[10].f.lower[19] );
tran (\sa_count[10][20] , \sa_count[10].r.part0[20] );
tran (\sa_count[10][20] , \sa_count[10].f.lower[20] );
tran (\sa_count[10][21] , \sa_count[10].r.part0[21] );
tran (\sa_count[10][21] , \sa_count[10].f.lower[21] );
tran (\sa_count[10][22] , \sa_count[10].r.part0[22] );
tran (\sa_count[10][22] , \sa_count[10].f.lower[22] );
tran (\sa_count[10][23] , \sa_count[10].r.part0[23] );
tran (\sa_count[10][23] , \sa_count[10].f.lower[23] );
tran (\sa_count[10][24] , \sa_count[10].r.part0[24] );
tran (\sa_count[10][24] , \sa_count[10].f.lower[24] );
tran (\sa_count[10][25] , \sa_count[10].r.part0[25] );
tran (\sa_count[10][25] , \sa_count[10].f.lower[25] );
tran (\sa_count[10][26] , \sa_count[10].r.part0[26] );
tran (\sa_count[10][26] , \sa_count[10].f.lower[26] );
tran (\sa_count[10][27] , \sa_count[10].r.part0[27] );
tran (\sa_count[10][27] , \sa_count[10].f.lower[27] );
tran (\sa_count[10][28] , \sa_count[10].r.part0[28] );
tran (\sa_count[10][28] , \sa_count[10].f.lower[28] );
tran (\sa_count[10][29] , \sa_count[10].r.part0[29] );
tran (\sa_count[10][29] , \sa_count[10].f.lower[29] );
tran (\sa_count[10][30] , \sa_count[10].r.part0[30] );
tran (\sa_count[10][30] , \sa_count[10].f.lower[30] );
tran (\sa_count[10][31] , \sa_count[10].r.part0[31] );
tran (\sa_count[10][31] , \sa_count[10].f.lower[31] );
tran (\sa_count[10][32] , \sa_count[10].r.part1[0] );
tran (\sa_count[10][32] , \sa_count[10].f.upper[0] );
tran (\sa_count[10][33] , \sa_count[10].r.part1[1] );
tran (\sa_count[10][33] , \sa_count[10].f.upper[1] );
tran (\sa_count[10][34] , \sa_count[10].r.part1[2] );
tran (\sa_count[10][34] , \sa_count[10].f.upper[2] );
tran (\sa_count[10][35] , \sa_count[10].r.part1[3] );
tran (\sa_count[10][35] , \sa_count[10].f.upper[3] );
tran (\sa_count[10][36] , \sa_count[10].r.part1[4] );
tran (\sa_count[10][36] , \sa_count[10].f.upper[4] );
tran (\sa_count[10][37] , \sa_count[10].r.part1[5] );
tran (\sa_count[10][37] , \sa_count[10].f.upper[5] );
tran (\sa_count[10][38] , \sa_count[10].r.part1[6] );
tran (\sa_count[10][38] , \sa_count[10].f.upper[6] );
tran (\sa_count[10][39] , \sa_count[10].r.part1[7] );
tran (\sa_count[10][39] , \sa_count[10].f.upper[7] );
tran (\sa_count[10][40] , \sa_count[10].r.part1[8] );
tran (\sa_count[10][40] , \sa_count[10].f.upper[8] );
tran (\sa_count[10][41] , \sa_count[10].r.part1[9] );
tran (\sa_count[10][41] , \sa_count[10].f.upper[9] );
tran (\sa_count[10][42] , \sa_count[10].r.part1[10] );
tran (\sa_count[10][42] , \sa_count[10].f.upper[10] );
tran (\sa_count[10][43] , \sa_count[10].r.part1[11] );
tran (\sa_count[10][43] , \sa_count[10].f.upper[11] );
tran (\sa_count[10][44] , \sa_count[10].r.part1[12] );
tran (\sa_count[10][44] , \sa_count[10].f.upper[12] );
tran (\sa_count[10][45] , \sa_count[10].r.part1[13] );
tran (\sa_count[10][45] , \sa_count[10].f.upper[13] );
tran (\sa_count[10][46] , \sa_count[10].r.part1[14] );
tran (\sa_count[10][46] , \sa_count[10].f.upper[14] );
tran (\sa_count[10][47] , \sa_count[10].r.part1[15] );
tran (\sa_count[10][47] , \sa_count[10].f.upper[15] );
tran (\sa_count[10][48] , \sa_count[10].r.part1[16] );
tran (\sa_count[10][48] , \sa_count[10].f.upper[16] );
tran (\sa_count[10][49] , \sa_count[10].r.part1[17] );
tran (\sa_count[10][49] , \sa_count[10].f.upper[17] );
tran (\sa_count[10][50] , \sa_count[10].r.part1[18] );
tran (\sa_count[10][50] , \sa_count[10].f.unused[0] );
tran (\sa_count[10][51] , \sa_count[10].r.part1[19] );
tran (\sa_count[10][51] , \sa_count[10].f.unused[1] );
tran (\sa_count[10][52] , \sa_count[10].r.part1[20] );
tran (\sa_count[10][52] , \sa_count[10].f.unused[2] );
tran (\sa_count[10][53] , \sa_count[10].r.part1[21] );
tran (\sa_count[10][53] , \sa_count[10].f.unused[3] );
tran (\sa_count[10][54] , \sa_count[10].r.part1[22] );
tran (\sa_count[10][54] , \sa_count[10].f.unused[4] );
tran (\sa_count[10][55] , \sa_count[10].r.part1[23] );
tran (\sa_count[10][55] , \sa_count[10].f.unused[5] );
tran (\sa_count[10][56] , \sa_count[10].r.part1[24] );
tran (\sa_count[10][56] , \sa_count[10].f.unused[6] );
tran (\sa_count[10][57] , \sa_count[10].r.part1[25] );
tran (\sa_count[10][57] , \sa_count[10].f.unused[7] );
tran (\sa_count[10][58] , \sa_count[10].r.part1[26] );
tran (\sa_count[10][58] , \sa_count[10].f.unused[8] );
tran (\sa_count[10][59] , \sa_count[10].r.part1[27] );
tran (\sa_count[10][59] , \sa_count[10].f.unused[9] );
tran (\sa_count[10][60] , \sa_count[10].r.part1[28] );
tran (\sa_count[10][60] , \sa_count[10].f.unused[10] );
tran (\sa_count[10][61] , \sa_count[10].r.part1[29] );
tran (\sa_count[10][61] , \sa_count[10].f.unused[11] );
tran (\sa_count[10][62] , \sa_count[10].r.part1[30] );
tran (\sa_count[10][62] , \sa_count[10].f.unused[12] );
tran (\sa_count[10][63] , \sa_count[10].r.part1[31] );
tran (\sa_count[10][63] , \sa_count[10].f.unused[13] );
tran (\sa_count[11][0] , \sa_count[11].r.part0[0] );
tran (\sa_count[11][0] , \sa_count[11].f.lower[0] );
tran (\sa_count[11][1] , \sa_count[11].r.part0[1] );
tran (\sa_count[11][1] , \sa_count[11].f.lower[1] );
tran (\sa_count[11][2] , \sa_count[11].r.part0[2] );
tran (\sa_count[11][2] , \sa_count[11].f.lower[2] );
tran (\sa_count[11][3] , \sa_count[11].r.part0[3] );
tran (\sa_count[11][3] , \sa_count[11].f.lower[3] );
tran (\sa_count[11][4] , \sa_count[11].r.part0[4] );
tran (\sa_count[11][4] , \sa_count[11].f.lower[4] );
tran (\sa_count[11][5] , \sa_count[11].r.part0[5] );
tran (\sa_count[11][5] , \sa_count[11].f.lower[5] );
tran (\sa_count[11][6] , \sa_count[11].r.part0[6] );
tran (\sa_count[11][6] , \sa_count[11].f.lower[6] );
tran (\sa_count[11][7] , \sa_count[11].r.part0[7] );
tran (\sa_count[11][7] , \sa_count[11].f.lower[7] );
tran (\sa_count[11][8] , \sa_count[11].r.part0[8] );
tran (\sa_count[11][8] , \sa_count[11].f.lower[8] );
tran (\sa_count[11][9] , \sa_count[11].r.part0[9] );
tran (\sa_count[11][9] , \sa_count[11].f.lower[9] );
tran (\sa_count[11][10] , \sa_count[11].r.part0[10] );
tran (\sa_count[11][10] , \sa_count[11].f.lower[10] );
tran (\sa_count[11][11] , \sa_count[11].r.part0[11] );
tran (\sa_count[11][11] , \sa_count[11].f.lower[11] );
tran (\sa_count[11][12] , \sa_count[11].r.part0[12] );
tran (\sa_count[11][12] , \sa_count[11].f.lower[12] );
tran (\sa_count[11][13] , \sa_count[11].r.part0[13] );
tran (\sa_count[11][13] , \sa_count[11].f.lower[13] );
tran (\sa_count[11][14] , \sa_count[11].r.part0[14] );
tran (\sa_count[11][14] , \sa_count[11].f.lower[14] );
tran (\sa_count[11][15] , \sa_count[11].r.part0[15] );
tran (\sa_count[11][15] , \sa_count[11].f.lower[15] );
tran (\sa_count[11][16] , \sa_count[11].r.part0[16] );
tran (\sa_count[11][16] , \sa_count[11].f.lower[16] );
tran (\sa_count[11][17] , \sa_count[11].r.part0[17] );
tran (\sa_count[11][17] , \sa_count[11].f.lower[17] );
tran (\sa_count[11][18] , \sa_count[11].r.part0[18] );
tran (\sa_count[11][18] , \sa_count[11].f.lower[18] );
tran (\sa_count[11][19] , \sa_count[11].r.part0[19] );
tran (\sa_count[11][19] , \sa_count[11].f.lower[19] );
tran (\sa_count[11][20] , \sa_count[11].r.part0[20] );
tran (\sa_count[11][20] , \sa_count[11].f.lower[20] );
tran (\sa_count[11][21] , \sa_count[11].r.part0[21] );
tran (\sa_count[11][21] , \sa_count[11].f.lower[21] );
tran (\sa_count[11][22] , \sa_count[11].r.part0[22] );
tran (\sa_count[11][22] , \sa_count[11].f.lower[22] );
tran (\sa_count[11][23] , \sa_count[11].r.part0[23] );
tran (\sa_count[11][23] , \sa_count[11].f.lower[23] );
tran (\sa_count[11][24] , \sa_count[11].r.part0[24] );
tran (\sa_count[11][24] , \sa_count[11].f.lower[24] );
tran (\sa_count[11][25] , \sa_count[11].r.part0[25] );
tran (\sa_count[11][25] , \sa_count[11].f.lower[25] );
tran (\sa_count[11][26] , \sa_count[11].r.part0[26] );
tran (\sa_count[11][26] , \sa_count[11].f.lower[26] );
tran (\sa_count[11][27] , \sa_count[11].r.part0[27] );
tran (\sa_count[11][27] , \sa_count[11].f.lower[27] );
tran (\sa_count[11][28] , \sa_count[11].r.part0[28] );
tran (\sa_count[11][28] , \sa_count[11].f.lower[28] );
tran (\sa_count[11][29] , \sa_count[11].r.part0[29] );
tran (\sa_count[11][29] , \sa_count[11].f.lower[29] );
tran (\sa_count[11][30] , \sa_count[11].r.part0[30] );
tran (\sa_count[11][30] , \sa_count[11].f.lower[30] );
tran (\sa_count[11][31] , \sa_count[11].r.part0[31] );
tran (\sa_count[11][31] , \sa_count[11].f.lower[31] );
tran (\sa_count[11][32] , \sa_count[11].r.part1[0] );
tran (\sa_count[11][32] , \sa_count[11].f.upper[0] );
tran (\sa_count[11][33] , \sa_count[11].r.part1[1] );
tran (\sa_count[11][33] , \sa_count[11].f.upper[1] );
tran (\sa_count[11][34] , \sa_count[11].r.part1[2] );
tran (\sa_count[11][34] , \sa_count[11].f.upper[2] );
tran (\sa_count[11][35] , \sa_count[11].r.part1[3] );
tran (\sa_count[11][35] , \sa_count[11].f.upper[3] );
tran (\sa_count[11][36] , \sa_count[11].r.part1[4] );
tran (\sa_count[11][36] , \sa_count[11].f.upper[4] );
tran (\sa_count[11][37] , \sa_count[11].r.part1[5] );
tran (\sa_count[11][37] , \sa_count[11].f.upper[5] );
tran (\sa_count[11][38] , \sa_count[11].r.part1[6] );
tran (\sa_count[11][38] , \sa_count[11].f.upper[6] );
tran (\sa_count[11][39] , \sa_count[11].r.part1[7] );
tran (\sa_count[11][39] , \sa_count[11].f.upper[7] );
tran (\sa_count[11][40] , \sa_count[11].r.part1[8] );
tran (\sa_count[11][40] , \sa_count[11].f.upper[8] );
tran (\sa_count[11][41] , \sa_count[11].r.part1[9] );
tran (\sa_count[11][41] , \sa_count[11].f.upper[9] );
tran (\sa_count[11][42] , \sa_count[11].r.part1[10] );
tran (\sa_count[11][42] , \sa_count[11].f.upper[10] );
tran (\sa_count[11][43] , \sa_count[11].r.part1[11] );
tran (\sa_count[11][43] , \sa_count[11].f.upper[11] );
tran (\sa_count[11][44] , \sa_count[11].r.part1[12] );
tran (\sa_count[11][44] , \sa_count[11].f.upper[12] );
tran (\sa_count[11][45] , \sa_count[11].r.part1[13] );
tran (\sa_count[11][45] , \sa_count[11].f.upper[13] );
tran (\sa_count[11][46] , \sa_count[11].r.part1[14] );
tran (\sa_count[11][46] , \sa_count[11].f.upper[14] );
tran (\sa_count[11][47] , \sa_count[11].r.part1[15] );
tran (\sa_count[11][47] , \sa_count[11].f.upper[15] );
tran (\sa_count[11][48] , \sa_count[11].r.part1[16] );
tran (\sa_count[11][48] , \sa_count[11].f.upper[16] );
tran (\sa_count[11][49] , \sa_count[11].r.part1[17] );
tran (\sa_count[11][49] , \sa_count[11].f.upper[17] );
tran (\sa_count[11][50] , \sa_count[11].r.part1[18] );
tran (\sa_count[11][50] , \sa_count[11].f.unused[0] );
tran (\sa_count[11][51] , \sa_count[11].r.part1[19] );
tran (\sa_count[11][51] , \sa_count[11].f.unused[1] );
tran (\sa_count[11][52] , \sa_count[11].r.part1[20] );
tran (\sa_count[11][52] , \sa_count[11].f.unused[2] );
tran (\sa_count[11][53] , \sa_count[11].r.part1[21] );
tran (\sa_count[11][53] , \sa_count[11].f.unused[3] );
tran (\sa_count[11][54] , \sa_count[11].r.part1[22] );
tran (\sa_count[11][54] , \sa_count[11].f.unused[4] );
tran (\sa_count[11][55] , \sa_count[11].r.part1[23] );
tran (\sa_count[11][55] , \sa_count[11].f.unused[5] );
tran (\sa_count[11][56] , \sa_count[11].r.part1[24] );
tran (\sa_count[11][56] , \sa_count[11].f.unused[6] );
tran (\sa_count[11][57] , \sa_count[11].r.part1[25] );
tran (\sa_count[11][57] , \sa_count[11].f.unused[7] );
tran (\sa_count[11][58] , \sa_count[11].r.part1[26] );
tran (\sa_count[11][58] , \sa_count[11].f.unused[8] );
tran (\sa_count[11][59] , \sa_count[11].r.part1[27] );
tran (\sa_count[11][59] , \sa_count[11].f.unused[9] );
tran (\sa_count[11][60] , \sa_count[11].r.part1[28] );
tran (\sa_count[11][60] , \sa_count[11].f.unused[10] );
tran (\sa_count[11][61] , \sa_count[11].r.part1[29] );
tran (\sa_count[11][61] , \sa_count[11].f.unused[11] );
tran (\sa_count[11][62] , \sa_count[11].r.part1[30] );
tran (\sa_count[11][62] , \sa_count[11].f.unused[12] );
tran (\sa_count[11][63] , \sa_count[11].r.part1[31] );
tran (\sa_count[11][63] , \sa_count[11].f.unused[13] );
tran (\sa_count[12][0] , \sa_count[12].r.part0[0] );
tran (\sa_count[12][0] , \sa_count[12].f.lower[0] );
tran (\sa_count[12][1] , \sa_count[12].r.part0[1] );
tran (\sa_count[12][1] , \sa_count[12].f.lower[1] );
tran (\sa_count[12][2] , \sa_count[12].r.part0[2] );
tran (\sa_count[12][2] , \sa_count[12].f.lower[2] );
tran (\sa_count[12][3] , \sa_count[12].r.part0[3] );
tran (\sa_count[12][3] , \sa_count[12].f.lower[3] );
tran (\sa_count[12][4] , \sa_count[12].r.part0[4] );
tran (\sa_count[12][4] , \sa_count[12].f.lower[4] );
tran (\sa_count[12][5] , \sa_count[12].r.part0[5] );
tran (\sa_count[12][5] , \sa_count[12].f.lower[5] );
tran (\sa_count[12][6] , \sa_count[12].r.part0[6] );
tran (\sa_count[12][6] , \sa_count[12].f.lower[6] );
tran (\sa_count[12][7] , \sa_count[12].r.part0[7] );
tran (\sa_count[12][7] , \sa_count[12].f.lower[7] );
tran (\sa_count[12][8] , \sa_count[12].r.part0[8] );
tran (\sa_count[12][8] , \sa_count[12].f.lower[8] );
tran (\sa_count[12][9] , \sa_count[12].r.part0[9] );
tran (\sa_count[12][9] , \sa_count[12].f.lower[9] );
tran (\sa_count[12][10] , \sa_count[12].r.part0[10] );
tran (\sa_count[12][10] , \sa_count[12].f.lower[10] );
tran (\sa_count[12][11] , \sa_count[12].r.part0[11] );
tran (\sa_count[12][11] , \sa_count[12].f.lower[11] );
tran (\sa_count[12][12] , \sa_count[12].r.part0[12] );
tran (\sa_count[12][12] , \sa_count[12].f.lower[12] );
tran (\sa_count[12][13] , \sa_count[12].r.part0[13] );
tran (\sa_count[12][13] , \sa_count[12].f.lower[13] );
tran (\sa_count[12][14] , \sa_count[12].r.part0[14] );
tran (\sa_count[12][14] , \sa_count[12].f.lower[14] );
tran (\sa_count[12][15] , \sa_count[12].r.part0[15] );
tran (\sa_count[12][15] , \sa_count[12].f.lower[15] );
tran (\sa_count[12][16] , \sa_count[12].r.part0[16] );
tran (\sa_count[12][16] , \sa_count[12].f.lower[16] );
tran (\sa_count[12][17] , \sa_count[12].r.part0[17] );
tran (\sa_count[12][17] , \sa_count[12].f.lower[17] );
tran (\sa_count[12][18] , \sa_count[12].r.part0[18] );
tran (\sa_count[12][18] , \sa_count[12].f.lower[18] );
tran (\sa_count[12][19] , \sa_count[12].r.part0[19] );
tran (\sa_count[12][19] , \sa_count[12].f.lower[19] );
tran (\sa_count[12][20] , \sa_count[12].r.part0[20] );
tran (\sa_count[12][20] , \sa_count[12].f.lower[20] );
tran (\sa_count[12][21] , \sa_count[12].r.part0[21] );
tran (\sa_count[12][21] , \sa_count[12].f.lower[21] );
tran (\sa_count[12][22] , \sa_count[12].r.part0[22] );
tran (\sa_count[12][22] , \sa_count[12].f.lower[22] );
tran (\sa_count[12][23] , \sa_count[12].r.part0[23] );
tran (\sa_count[12][23] , \sa_count[12].f.lower[23] );
tran (\sa_count[12][24] , \sa_count[12].r.part0[24] );
tran (\sa_count[12][24] , \sa_count[12].f.lower[24] );
tran (\sa_count[12][25] , \sa_count[12].r.part0[25] );
tran (\sa_count[12][25] , \sa_count[12].f.lower[25] );
tran (\sa_count[12][26] , \sa_count[12].r.part0[26] );
tran (\sa_count[12][26] , \sa_count[12].f.lower[26] );
tran (\sa_count[12][27] , \sa_count[12].r.part0[27] );
tran (\sa_count[12][27] , \sa_count[12].f.lower[27] );
tran (\sa_count[12][28] , \sa_count[12].r.part0[28] );
tran (\sa_count[12][28] , \sa_count[12].f.lower[28] );
tran (\sa_count[12][29] , \sa_count[12].r.part0[29] );
tran (\sa_count[12][29] , \sa_count[12].f.lower[29] );
tran (\sa_count[12][30] , \sa_count[12].r.part0[30] );
tran (\sa_count[12][30] , \sa_count[12].f.lower[30] );
tran (\sa_count[12][31] , \sa_count[12].r.part0[31] );
tran (\sa_count[12][31] , \sa_count[12].f.lower[31] );
tran (\sa_count[12][32] , \sa_count[12].r.part1[0] );
tran (\sa_count[12][32] , \sa_count[12].f.upper[0] );
tran (\sa_count[12][33] , \sa_count[12].r.part1[1] );
tran (\sa_count[12][33] , \sa_count[12].f.upper[1] );
tran (\sa_count[12][34] , \sa_count[12].r.part1[2] );
tran (\sa_count[12][34] , \sa_count[12].f.upper[2] );
tran (\sa_count[12][35] , \sa_count[12].r.part1[3] );
tran (\sa_count[12][35] , \sa_count[12].f.upper[3] );
tran (\sa_count[12][36] , \sa_count[12].r.part1[4] );
tran (\sa_count[12][36] , \sa_count[12].f.upper[4] );
tran (\sa_count[12][37] , \sa_count[12].r.part1[5] );
tran (\sa_count[12][37] , \sa_count[12].f.upper[5] );
tran (\sa_count[12][38] , \sa_count[12].r.part1[6] );
tran (\sa_count[12][38] , \sa_count[12].f.upper[6] );
tran (\sa_count[12][39] , \sa_count[12].r.part1[7] );
tran (\sa_count[12][39] , \sa_count[12].f.upper[7] );
tran (\sa_count[12][40] , \sa_count[12].r.part1[8] );
tran (\sa_count[12][40] , \sa_count[12].f.upper[8] );
tran (\sa_count[12][41] , \sa_count[12].r.part1[9] );
tran (\sa_count[12][41] , \sa_count[12].f.upper[9] );
tran (\sa_count[12][42] , \sa_count[12].r.part1[10] );
tran (\sa_count[12][42] , \sa_count[12].f.upper[10] );
tran (\sa_count[12][43] , \sa_count[12].r.part1[11] );
tran (\sa_count[12][43] , \sa_count[12].f.upper[11] );
tran (\sa_count[12][44] , \sa_count[12].r.part1[12] );
tran (\sa_count[12][44] , \sa_count[12].f.upper[12] );
tran (\sa_count[12][45] , \sa_count[12].r.part1[13] );
tran (\sa_count[12][45] , \sa_count[12].f.upper[13] );
tran (\sa_count[12][46] , \sa_count[12].r.part1[14] );
tran (\sa_count[12][46] , \sa_count[12].f.upper[14] );
tran (\sa_count[12][47] , \sa_count[12].r.part1[15] );
tran (\sa_count[12][47] , \sa_count[12].f.upper[15] );
tran (\sa_count[12][48] , \sa_count[12].r.part1[16] );
tran (\sa_count[12][48] , \sa_count[12].f.upper[16] );
tran (\sa_count[12][49] , \sa_count[12].r.part1[17] );
tran (\sa_count[12][49] , \sa_count[12].f.upper[17] );
tran (\sa_count[12][50] , \sa_count[12].r.part1[18] );
tran (\sa_count[12][50] , \sa_count[12].f.unused[0] );
tran (\sa_count[12][51] , \sa_count[12].r.part1[19] );
tran (\sa_count[12][51] , \sa_count[12].f.unused[1] );
tran (\sa_count[12][52] , \sa_count[12].r.part1[20] );
tran (\sa_count[12][52] , \sa_count[12].f.unused[2] );
tran (\sa_count[12][53] , \sa_count[12].r.part1[21] );
tran (\sa_count[12][53] , \sa_count[12].f.unused[3] );
tran (\sa_count[12][54] , \sa_count[12].r.part1[22] );
tran (\sa_count[12][54] , \sa_count[12].f.unused[4] );
tran (\sa_count[12][55] , \sa_count[12].r.part1[23] );
tran (\sa_count[12][55] , \sa_count[12].f.unused[5] );
tran (\sa_count[12][56] , \sa_count[12].r.part1[24] );
tran (\sa_count[12][56] , \sa_count[12].f.unused[6] );
tran (\sa_count[12][57] , \sa_count[12].r.part1[25] );
tran (\sa_count[12][57] , \sa_count[12].f.unused[7] );
tran (\sa_count[12][58] , \sa_count[12].r.part1[26] );
tran (\sa_count[12][58] , \sa_count[12].f.unused[8] );
tran (\sa_count[12][59] , \sa_count[12].r.part1[27] );
tran (\sa_count[12][59] , \sa_count[12].f.unused[9] );
tran (\sa_count[12][60] , \sa_count[12].r.part1[28] );
tran (\sa_count[12][60] , \sa_count[12].f.unused[10] );
tran (\sa_count[12][61] , \sa_count[12].r.part1[29] );
tran (\sa_count[12][61] , \sa_count[12].f.unused[11] );
tran (\sa_count[12][62] , \sa_count[12].r.part1[30] );
tran (\sa_count[12][62] , \sa_count[12].f.unused[12] );
tran (\sa_count[12][63] , \sa_count[12].r.part1[31] );
tran (\sa_count[12][63] , \sa_count[12].f.unused[13] );
tran (\sa_count[13][0] , \sa_count[13].r.part0[0] );
tran (\sa_count[13][0] , \sa_count[13].f.lower[0] );
tran (\sa_count[13][1] , \sa_count[13].r.part0[1] );
tran (\sa_count[13][1] , \sa_count[13].f.lower[1] );
tran (\sa_count[13][2] , \sa_count[13].r.part0[2] );
tran (\sa_count[13][2] , \sa_count[13].f.lower[2] );
tran (\sa_count[13][3] , \sa_count[13].r.part0[3] );
tran (\sa_count[13][3] , \sa_count[13].f.lower[3] );
tran (\sa_count[13][4] , \sa_count[13].r.part0[4] );
tran (\sa_count[13][4] , \sa_count[13].f.lower[4] );
tran (\sa_count[13][5] , \sa_count[13].r.part0[5] );
tran (\sa_count[13][5] , \sa_count[13].f.lower[5] );
tran (\sa_count[13][6] , \sa_count[13].r.part0[6] );
tran (\sa_count[13][6] , \sa_count[13].f.lower[6] );
tran (\sa_count[13][7] , \sa_count[13].r.part0[7] );
tran (\sa_count[13][7] , \sa_count[13].f.lower[7] );
tran (\sa_count[13][8] , \sa_count[13].r.part0[8] );
tran (\sa_count[13][8] , \sa_count[13].f.lower[8] );
tran (\sa_count[13][9] , \sa_count[13].r.part0[9] );
tran (\sa_count[13][9] , \sa_count[13].f.lower[9] );
tran (\sa_count[13][10] , \sa_count[13].r.part0[10] );
tran (\sa_count[13][10] , \sa_count[13].f.lower[10] );
tran (\sa_count[13][11] , \sa_count[13].r.part0[11] );
tran (\sa_count[13][11] , \sa_count[13].f.lower[11] );
tran (\sa_count[13][12] , \sa_count[13].r.part0[12] );
tran (\sa_count[13][12] , \sa_count[13].f.lower[12] );
tran (\sa_count[13][13] , \sa_count[13].r.part0[13] );
tran (\sa_count[13][13] , \sa_count[13].f.lower[13] );
tran (\sa_count[13][14] , \sa_count[13].r.part0[14] );
tran (\sa_count[13][14] , \sa_count[13].f.lower[14] );
tran (\sa_count[13][15] , \sa_count[13].r.part0[15] );
tran (\sa_count[13][15] , \sa_count[13].f.lower[15] );
tran (\sa_count[13][16] , \sa_count[13].r.part0[16] );
tran (\sa_count[13][16] , \sa_count[13].f.lower[16] );
tran (\sa_count[13][17] , \sa_count[13].r.part0[17] );
tran (\sa_count[13][17] , \sa_count[13].f.lower[17] );
tran (\sa_count[13][18] , \sa_count[13].r.part0[18] );
tran (\sa_count[13][18] , \sa_count[13].f.lower[18] );
tran (\sa_count[13][19] , \sa_count[13].r.part0[19] );
tran (\sa_count[13][19] , \sa_count[13].f.lower[19] );
tran (\sa_count[13][20] , \sa_count[13].r.part0[20] );
tran (\sa_count[13][20] , \sa_count[13].f.lower[20] );
tran (\sa_count[13][21] , \sa_count[13].r.part0[21] );
tran (\sa_count[13][21] , \sa_count[13].f.lower[21] );
tran (\sa_count[13][22] , \sa_count[13].r.part0[22] );
tran (\sa_count[13][22] , \sa_count[13].f.lower[22] );
tran (\sa_count[13][23] , \sa_count[13].r.part0[23] );
tran (\sa_count[13][23] , \sa_count[13].f.lower[23] );
tran (\sa_count[13][24] , \sa_count[13].r.part0[24] );
tran (\sa_count[13][24] , \sa_count[13].f.lower[24] );
tran (\sa_count[13][25] , \sa_count[13].r.part0[25] );
tran (\sa_count[13][25] , \sa_count[13].f.lower[25] );
tran (\sa_count[13][26] , \sa_count[13].r.part0[26] );
tran (\sa_count[13][26] , \sa_count[13].f.lower[26] );
tran (\sa_count[13][27] , \sa_count[13].r.part0[27] );
tran (\sa_count[13][27] , \sa_count[13].f.lower[27] );
tran (\sa_count[13][28] , \sa_count[13].r.part0[28] );
tran (\sa_count[13][28] , \sa_count[13].f.lower[28] );
tran (\sa_count[13][29] , \sa_count[13].r.part0[29] );
tran (\sa_count[13][29] , \sa_count[13].f.lower[29] );
tran (\sa_count[13][30] , \sa_count[13].r.part0[30] );
tran (\sa_count[13][30] , \sa_count[13].f.lower[30] );
tran (\sa_count[13][31] , \sa_count[13].r.part0[31] );
tran (\sa_count[13][31] , \sa_count[13].f.lower[31] );
tran (\sa_count[13][32] , \sa_count[13].r.part1[0] );
tran (\sa_count[13][32] , \sa_count[13].f.upper[0] );
tran (\sa_count[13][33] , \sa_count[13].r.part1[1] );
tran (\sa_count[13][33] , \sa_count[13].f.upper[1] );
tran (\sa_count[13][34] , \sa_count[13].r.part1[2] );
tran (\sa_count[13][34] , \sa_count[13].f.upper[2] );
tran (\sa_count[13][35] , \sa_count[13].r.part1[3] );
tran (\sa_count[13][35] , \sa_count[13].f.upper[3] );
tran (\sa_count[13][36] , \sa_count[13].r.part1[4] );
tran (\sa_count[13][36] , \sa_count[13].f.upper[4] );
tran (\sa_count[13][37] , \sa_count[13].r.part1[5] );
tran (\sa_count[13][37] , \sa_count[13].f.upper[5] );
tran (\sa_count[13][38] , \sa_count[13].r.part1[6] );
tran (\sa_count[13][38] , \sa_count[13].f.upper[6] );
tran (\sa_count[13][39] , \sa_count[13].r.part1[7] );
tran (\sa_count[13][39] , \sa_count[13].f.upper[7] );
tran (\sa_count[13][40] , \sa_count[13].r.part1[8] );
tran (\sa_count[13][40] , \sa_count[13].f.upper[8] );
tran (\sa_count[13][41] , \sa_count[13].r.part1[9] );
tran (\sa_count[13][41] , \sa_count[13].f.upper[9] );
tran (\sa_count[13][42] , \sa_count[13].r.part1[10] );
tran (\sa_count[13][42] , \sa_count[13].f.upper[10] );
tran (\sa_count[13][43] , \sa_count[13].r.part1[11] );
tran (\sa_count[13][43] , \sa_count[13].f.upper[11] );
tran (\sa_count[13][44] , \sa_count[13].r.part1[12] );
tran (\sa_count[13][44] , \sa_count[13].f.upper[12] );
tran (\sa_count[13][45] , \sa_count[13].r.part1[13] );
tran (\sa_count[13][45] , \sa_count[13].f.upper[13] );
tran (\sa_count[13][46] , \sa_count[13].r.part1[14] );
tran (\sa_count[13][46] , \sa_count[13].f.upper[14] );
tran (\sa_count[13][47] , \sa_count[13].r.part1[15] );
tran (\sa_count[13][47] , \sa_count[13].f.upper[15] );
tran (\sa_count[13][48] , \sa_count[13].r.part1[16] );
tran (\sa_count[13][48] , \sa_count[13].f.upper[16] );
tran (\sa_count[13][49] , \sa_count[13].r.part1[17] );
tran (\sa_count[13][49] , \sa_count[13].f.upper[17] );
tran (\sa_count[13][50] , \sa_count[13].r.part1[18] );
tran (\sa_count[13][50] , \sa_count[13].f.unused[0] );
tran (\sa_count[13][51] , \sa_count[13].r.part1[19] );
tran (\sa_count[13][51] , \sa_count[13].f.unused[1] );
tran (\sa_count[13][52] , \sa_count[13].r.part1[20] );
tran (\sa_count[13][52] , \sa_count[13].f.unused[2] );
tran (\sa_count[13][53] , \sa_count[13].r.part1[21] );
tran (\sa_count[13][53] , \sa_count[13].f.unused[3] );
tran (\sa_count[13][54] , \sa_count[13].r.part1[22] );
tran (\sa_count[13][54] , \sa_count[13].f.unused[4] );
tran (\sa_count[13][55] , \sa_count[13].r.part1[23] );
tran (\sa_count[13][55] , \sa_count[13].f.unused[5] );
tran (\sa_count[13][56] , \sa_count[13].r.part1[24] );
tran (\sa_count[13][56] , \sa_count[13].f.unused[6] );
tran (\sa_count[13][57] , \sa_count[13].r.part1[25] );
tran (\sa_count[13][57] , \sa_count[13].f.unused[7] );
tran (\sa_count[13][58] , \sa_count[13].r.part1[26] );
tran (\sa_count[13][58] , \sa_count[13].f.unused[8] );
tran (\sa_count[13][59] , \sa_count[13].r.part1[27] );
tran (\sa_count[13][59] , \sa_count[13].f.unused[9] );
tran (\sa_count[13][60] , \sa_count[13].r.part1[28] );
tran (\sa_count[13][60] , \sa_count[13].f.unused[10] );
tran (\sa_count[13][61] , \sa_count[13].r.part1[29] );
tran (\sa_count[13][61] , \sa_count[13].f.unused[11] );
tran (\sa_count[13][62] , \sa_count[13].r.part1[30] );
tran (\sa_count[13][62] , \sa_count[13].f.unused[12] );
tran (\sa_count[13][63] , \sa_count[13].r.part1[31] );
tran (\sa_count[13][63] , \sa_count[13].f.unused[13] );
tran (\sa_count[14][0] , \sa_count[14].r.part0[0] );
tran (\sa_count[14][0] , \sa_count[14].f.lower[0] );
tran (\sa_count[14][1] , \sa_count[14].r.part0[1] );
tran (\sa_count[14][1] , \sa_count[14].f.lower[1] );
tran (\sa_count[14][2] , \sa_count[14].r.part0[2] );
tran (\sa_count[14][2] , \sa_count[14].f.lower[2] );
tran (\sa_count[14][3] , \sa_count[14].r.part0[3] );
tran (\sa_count[14][3] , \sa_count[14].f.lower[3] );
tran (\sa_count[14][4] , \sa_count[14].r.part0[4] );
tran (\sa_count[14][4] , \sa_count[14].f.lower[4] );
tran (\sa_count[14][5] , \sa_count[14].r.part0[5] );
tran (\sa_count[14][5] , \sa_count[14].f.lower[5] );
tran (\sa_count[14][6] , \sa_count[14].r.part0[6] );
tran (\sa_count[14][6] , \sa_count[14].f.lower[6] );
tran (\sa_count[14][7] , \sa_count[14].r.part0[7] );
tran (\sa_count[14][7] , \sa_count[14].f.lower[7] );
tran (\sa_count[14][8] , \sa_count[14].r.part0[8] );
tran (\sa_count[14][8] , \sa_count[14].f.lower[8] );
tran (\sa_count[14][9] , \sa_count[14].r.part0[9] );
tran (\sa_count[14][9] , \sa_count[14].f.lower[9] );
tran (\sa_count[14][10] , \sa_count[14].r.part0[10] );
tran (\sa_count[14][10] , \sa_count[14].f.lower[10] );
tran (\sa_count[14][11] , \sa_count[14].r.part0[11] );
tran (\sa_count[14][11] , \sa_count[14].f.lower[11] );
tran (\sa_count[14][12] , \sa_count[14].r.part0[12] );
tran (\sa_count[14][12] , \sa_count[14].f.lower[12] );
tran (\sa_count[14][13] , \sa_count[14].r.part0[13] );
tran (\sa_count[14][13] , \sa_count[14].f.lower[13] );
tran (\sa_count[14][14] , \sa_count[14].r.part0[14] );
tran (\sa_count[14][14] , \sa_count[14].f.lower[14] );
tran (\sa_count[14][15] , \sa_count[14].r.part0[15] );
tran (\sa_count[14][15] , \sa_count[14].f.lower[15] );
tran (\sa_count[14][16] , \sa_count[14].r.part0[16] );
tran (\sa_count[14][16] , \sa_count[14].f.lower[16] );
tran (\sa_count[14][17] , \sa_count[14].r.part0[17] );
tran (\sa_count[14][17] , \sa_count[14].f.lower[17] );
tran (\sa_count[14][18] , \sa_count[14].r.part0[18] );
tran (\sa_count[14][18] , \sa_count[14].f.lower[18] );
tran (\sa_count[14][19] , \sa_count[14].r.part0[19] );
tran (\sa_count[14][19] , \sa_count[14].f.lower[19] );
tran (\sa_count[14][20] , \sa_count[14].r.part0[20] );
tran (\sa_count[14][20] , \sa_count[14].f.lower[20] );
tran (\sa_count[14][21] , \sa_count[14].r.part0[21] );
tran (\sa_count[14][21] , \sa_count[14].f.lower[21] );
tran (\sa_count[14][22] , \sa_count[14].r.part0[22] );
tran (\sa_count[14][22] , \sa_count[14].f.lower[22] );
tran (\sa_count[14][23] , \sa_count[14].r.part0[23] );
tran (\sa_count[14][23] , \sa_count[14].f.lower[23] );
tran (\sa_count[14][24] , \sa_count[14].r.part0[24] );
tran (\sa_count[14][24] , \sa_count[14].f.lower[24] );
tran (\sa_count[14][25] , \sa_count[14].r.part0[25] );
tran (\sa_count[14][25] , \sa_count[14].f.lower[25] );
tran (\sa_count[14][26] , \sa_count[14].r.part0[26] );
tran (\sa_count[14][26] , \sa_count[14].f.lower[26] );
tran (\sa_count[14][27] , \sa_count[14].r.part0[27] );
tran (\sa_count[14][27] , \sa_count[14].f.lower[27] );
tran (\sa_count[14][28] , \sa_count[14].r.part0[28] );
tran (\sa_count[14][28] , \sa_count[14].f.lower[28] );
tran (\sa_count[14][29] , \sa_count[14].r.part0[29] );
tran (\sa_count[14][29] , \sa_count[14].f.lower[29] );
tran (\sa_count[14][30] , \sa_count[14].r.part0[30] );
tran (\sa_count[14][30] , \sa_count[14].f.lower[30] );
tran (\sa_count[14][31] , \sa_count[14].r.part0[31] );
tran (\sa_count[14][31] , \sa_count[14].f.lower[31] );
tran (\sa_count[14][32] , \sa_count[14].r.part1[0] );
tran (\sa_count[14][32] , \sa_count[14].f.upper[0] );
tran (\sa_count[14][33] , \sa_count[14].r.part1[1] );
tran (\sa_count[14][33] , \sa_count[14].f.upper[1] );
tran (\sa_count[14][34] , \sa_count[14].r.part1[2] );
tran (\sa_count[14][34] , \sa_count[14].f.upper[2] );
tran (\sa_count[14][35] , \sa_count[14].r.part1[3] );
tran (\sa_count[14][35] , \sa_count[14].f.upper[3] );
tran (\sa_count[14][36] , \sa_count[14].r.part1[4] );
tran (\sa_count[14][36] , \sa_count[14].f.upper[4] );
tran (\sa_count[14][37] , \sa_count[14].r.part1[5] );
tran (\sa_count[14][37] , \sa_count[14].f.upper[5] );
tran (\sa_count[14][38] , \sa_count[14].r.part1[6] );
tran (\sa_count[14][38] , \sa_count[14].f.upper[6] );
tran (\sa_count[14][39] , \sa_count[14].r.part1[7] );
tran (\sa_count[14][39] , \sa_count[14].f.upper[7] );
tran (\sa_count[14][40] , \sa_count[14].r.part1[8] );
tran (\sa_count[14][40] , \sa_count[14].f.upper[8] );
tran (\sa_count[14][41] , \sa_count[14].r.part1[9] );
tran (\sa_count[14][41] , \sa_count[14].f.upper[9] );
tran (\sa_count[14][42] , \sa_count[14].r.part1[10] );
tran (\sa_count[14][42] , \sa_count[14].f.upper[10] );
tran (\sa_count[14][43] , \sa_count[14].r.part1[11] );
tran (\sa_count[14][43] , \sa_count[14].f.upper[11] );
tran (\sa_count[14][44] , \sa_count[14].r.part1[12] );
tran (\sa_count[14][44] , \sa_count[14].f.upper[12] );
tran (\sa_count[14][45] , \sa_count[14].r.part1[13] );
tran (\sa_count[14][45] , \sa_count[14].f.upper[13] );
tran (\sa_count[14][46] , \sa_count[14].r.part1[14] );
tran (\sa_count[14][46] , \sa_count[14].f.upper[14] );
tran (\sa_count[14][47] , \sa_count[14].r.part1[15] );
tran (\sa_count[14][47] , \sa_count[14].f.upper[15] );
tran (\sa_count[14][48] , \sa_count[14].r.part1[16] );
tran (\sa_count[14][48] , \sa_count[14].f.upper[16] );
tran (\sa_count[14][49] , \sa_count[14].r.part1[17] );
tran (\sa_count[14][49] , \sa_count[14].f.upper[17] );
tran (\sa_count[14][50] , \sa_count[14].r.part1[18] );
tran (\sa_count[14][50] , \sa_count[14].f.unused[0] );
tran (\sa_count[14][51] , \sa_count[14].r.part1[19] );
tran (\sa_count[14][51] , \sa_count[14].f.unused[1] );
tran (\sa_count[14][52] , \sa_count[14].r.part1[20] );
tran (\sa_count[14][52] , \sa_count[14].f.unused[2] );
tran (\sa_count[14][53] , \sa_count[14].r.part1[21] );
tran (\sa_count[14][53] , \sa_count[14].f.unused[3] );
tran (\sa_count[14][54] , \sa_count[14].r.part1[22] );
tran (\sa_count[14][54] , \sa_count[14].f.unused[4] );
tran (\sa_count[14][55] , \sa_count[14].r.part1[23] );
tran (\sa_count[14][55] , \sa_count[14].f.unused[5] );
tran (\sa_count[14][56] , \sa_count[14].r.part1[24] );
tran (\sa_count[14][56] , \sa_count[14].f.unused[6] );
tran (\sa_count[14][57] , \sa_count[14].r.part1[25] );
tran (\sa_count[14][57] , \sa_count[14].f.unused[7] );
tran (\sa_count[14][58] , \sa_count[14].r.part1[26] );
tran (\sa_count[14][58] , \sa_count[14].f.unused[8] );
tran (\sa_count[14][59] , \sa_count[14].r.part1[27] );
tran (\sa_count[14][59] , \sa_count[14].f.unused[9] );
tran (\sa_count[14][60] , \sa_count[14].r.part1[28] );
tran (\sa_count[14][60] , \sa_count[14].f.unused[10] );
tran (\sa_count[14][61] , \sa_count[14].r.part1[29] );
tran (\sa_count[14][61] , \sa_count[14].f.unused[11] );
tran (\sa_count[14][62] , \sa_count[14].r.part1[30] );
tran (\sa_count[14][62] , \sa_count[14].f.unused[12] );
tran (\sa_count[14][63] , \sa_count[14].r.part1[31] );
tran (\sa_count[14][63] , \sa_count[14].f.unused[13] );
tran (\sa_count[15][0] , \sa_count[15].r.part0[0] );
tran (\sa_count[15][0] , \sa_count[15].f.lower[0] );
tran (\sa_count[15][1] , \sa_count[15].r.part0[1] );
tran (\sa_count[15][1] , \sa_count[15].f.lower[1] );
tran (\sa_count[15][2] , \sa_count[15].r.part0[2] );
tran (\sa_count[15][2] , \sa_count[15].f.lower[2] );
tran (\sa_count[15][3] , \sa_count[15].r.part0[3] );
tran (\sa_count[15][3] , \sa_count[15].f.lower[3] );
tran (\sa_count[15][4] , \sa_count[15].r.part0[4] );
tran (\sa_count[15][4] , \sa_count[15].f.lower[4] );
tran (\sa_count[15][5] , \sa_count[15].r.part0[5] );
tran (\sa_count[15][5] , \sa_count[15].f.lower[5] );
tran (\sa_count[15][6] , \sa_count[15].r.part0[6] );
tran (\sa_count[15][6] , \sa_count[15].f.lower[6] );
tran (\sa_count[15][7] , \sa_count[15].r.part0[7] );
tran (\sa_count[15][7] , \sa_count[15].f.lower[7] );
tran (\sa_count[15][8] , \sa_count[15].r.part0[8] );
tran (\sa_count[15][8] , \sa_count[15].f.lower[8] );
tran (\sa_count[15][9] , \sa_count[15].r.part0[9] );
tran (\sa_count[15][9] , \sa_count[15].f.lower[9] );
tran (\sa_count[15][10] , \sa_count[15].r.part0[10] );
tran (\sa_count[15][10] , \sa_count[15].f.lower[10] );
tran (\sa_count[15][11] , \sa_count[15].r.part0[11] );
tran (\sa_count[15][11] , \sa_count[15].f.lower[11] );
tran (\sa_count[15][12] , \sa_count[15].r.part0[12] );
tran (\sa_count[15][12] , \sa_count[15].f.lower[12] );
tran (\sa_count[15][13] , \sa_count[15].r.part0[13] );
tran (\sa_count[15][13] , \sa_count[15].f.lower[13] );
tran (\sa_count[15][14] , \sa_count[15].r.part0[14] );
tran (\sa_count[15][14] , \sa_count[15].f.lower[14] );
tran (\sa_count[15][15] , \sa_count[15].r.part0[15] );
tran (\sa_count[15][15] , \sa_count[15].f.lower[15] );
tran (\sa_count[15][16] , \sa_count[15].r.part0[16] );
tran (\sa_count[15][16] , \sa_count[15].f.lower[16] );
tran (\sa_count[15][17] , \sa_count[15].r.part0[17] );
tran (\sa_count[15][17] , \sa_count[15].f.lower[17] );
tran (\sa_count[15][18] , \sa_count[15].r.part0[18] );
tran (\sa_count[15][18] , \sa_count[15].f.lower[18] );
tran (\sa_count[15][19] , \sa_count[15].r.part0[19] );
tran (\sa_count[15][19] , \sa_count[15].f.lower[19] );
tran (\sa_count[15][20] , \sa_count[15].r.part0[20] );
tran (\sa_count[15][20] , \sa_count[15].f.lower[20] );
tran (\sa_count[15][21] , \sa_count[15].r.part0[21] );
tran (\sa_count[15][21] , \sa_count[15].f.lower[21] );
tran (\sa_count[15][22] , \sa_count[15].r.part0[22] );
tran (\sa_count[15][22] , \sa_count[15].f.lower[22] );
tran (\sa_count[15][23] , \sa_count[15].r.part0[23] );
tran (\sa_count[15][23] , \sa_count[15].f.lower[23] );
tran (\sa_count[15][24] , \sa_count[15].r.part0[24] );
tran (\sa_count[15][24] , \sa_count[15].f.lower[24] );
tran (\sa_count[15][25] , \sa_count[15].r.part0[25] );
tran (\sa_count[15][25] , \sa_count[15].f.lower[25] );
tran (\sa_count[15][26] , \sa_count[15].r.part0[26] );
tran (\sa_count[15][26] , \sa_count[15].f.lower[26] );
tran (\sa_count[15][27] , \sa_count[15].r.part0[27] );
tran (\sa_count[15][27] , \sa_count[15].f.lower[27] );
tran (\sa_count[15][28] , \sa_count[15].r.part0[28] );
tran (\sa_count[15][28] , \sa_count[15].f.lower[28] );
tran (\sa_count[15][29] , \sa_count[15].r.part0[29] );
tran (\sa_count[15][29] , \sa_count[15].f.lower[29] );
tran (\sa_count[15][30] , \sa_count[15].r.part0[30] );
tran (\sa_count[15][30] , \sa_count[15].f.lower[30] );
tran (\sa_count[15][31] , \sa_count[15].r.part0[31] );
tran (\sa_count[15][31] , \sa_count[15].f.lower[31] );
tran (\sa_count[15][32] , \sa_count[15].r.part1[0] );
tran (\sa_count[15][32] , \sa_count[15].f.upper[0] );
tran (\sa_count[15][33] , \sa_count[15].r.part1[1] );
tran (\sa_count[15][33] , \sa_count[15].f.upper[1] );
tran (\sa_count[15][34] , \sa_count[15].r.part1[2] );
tran (\sa_count[15][34] , \sa_count[15].f.upper[2] );
tran (\sa_count[15][35] , \sa_count[15].r.part1[3] );
tran (\sa_count[15][35] , \sa_count[15].f.upper[3] );
tran (\sa_count[15][36] , \sa_count[15].r.part1[4] );
tran (\sa_count[15][36] , \sa_count[15].f.upper[4] );
tran (\sa_count[15][37] , \sa_count[15].r.part1[5] );
tran (\sa_count[15][37] , \sa_count[15].f.upper[5] );
tran (\sa_count[15][38] , \sa_count[15].r.part1[6] );
tran (\sa_count[15][38] , \sa_count[15].f.upper[6] );
tran (\sa_count[15][39] , \sa_count[15].r.part1[7] );
tran (\sa_count[15][39] , \sa_count[15].f.upper[7] );
tran (\sa_count[15][40] , \sa_count[15].r.part1[8] );
tran (\sa_count[15][40] , \sa_count[15].f.upper[8] );
tran (\sa_count[15][41] , \sa_count[15].r.part1[9] );
tran (\sa_count[15][41] , \sa_count[15].f.upper[9] );
tran (\sa_count[15][42] , \sa_count[15].r.part1[10] );
tran (\sa_count[15][42] , \sa_count[15].f.upper[10] );
tran (\sa_count[15][43] , \sa_count[15].r.part1[11] );
tran (\sa_count[15][43] , \sa_count[15].f.upper[11] );
tran (\sa_count[15][44] , \sa_count[15].r.part1[12] );
tran (\sa_count[15][44] , \sa_count[15].f.upper[12] );
tran (\sa_count[15][45] , \sa_count[15].r.part1[13] );
tran (\sa_count[15][45] , \sa_count[15].f.upper[13] );
tran (\sa_count[15][46] , \sa_count[15].r.part1[14] );
tran (\sa_count[15][46] , \sa_count[15].f.upper[14] );
tran (\sa_count[15][47] , \sa_count[15].r.part1[15] );
tran (\sa_count[15][47] , \sa_count[15].f.upper[15] );
tran (\sa_count[15][48] , \sa_count[15].r.part1[16] );
tran (\sa_count[15][48] , \sa_count[15].f.upper[16] );
tran (\sa_count[15][49] , \sa_count[15].r.part1[17] );
tran (\sa_count[15][49] , \sa_count[15].f.upper[17] );
tran (\sa_count[15][50] , \sa_count[15].r.part1[18] );
tran (\sa_count[15][50] , \sa_count[15].f.unused[0] );
tran (\sa_count[15][51] , \sa_count[15].r.part1[19] );
tran (\sa_count[15][51] , \sa_count[15].f.unused[1] );
tran (\sa_count[15][52] , \sa_count[15].r.part1[20] );
tran (\sa_count[15][52] , \sa_count[15].f.unused[2] );
tran (\sa_count[15][53] , \sa_count[15].r.part1[21] );
tran (\sa_count[15][53] , \sa_count[15].f.unused[3] );
tran (\sa_count[15][54] , \sa_count[15].r.part1[22] );
tran (\sa_count[15][54] , \sa_count[15].f.unused[4] );
tran (\sa_count[15][55] , \sa_count[15].r.part1[23] );
tran (\sa_count[15][55] , \sa_count[15].f.unused[5] );
tran (\sa_count[15][56] , \sa_count[15].r.part1[24] );
tran (\sa_count[15][56] , \sa_count[15].f.unused[6] );
tran (\sa_count[15][57] , \sa_count[15].r.part1[25] );
tran (\sa_count[15][57] , \sa_count[15].f.unused[7] );
tran (\sa_count[15][58] , \sa_count[15].r.part1[26] );
tran (\sa_count[15][58] , \sa_count[15].f.unused[8] );
tran (\sa_count[15][59] , \sa_count[15].r.part1[27] );
tran (\sa_count[15][59] , \sa_count[15].f.unused[9] );
tran (\sa_count[15][60] , \sa_count[15].r.part1[28] );
tran (\sa_count[15][60] , \sa_count[15].f.unused[10] );
tran (\sa_count[15][61] , \sa_count[15].r.part1[29] );
tran (\sa_count[15][61] , \sa_count[15].f.unused[11] );
tran (\sa_count[15][62] , \sa_count[15].r.part1[30] );
tran (\sa_count[15][62] , \sa_count[15].f.unused[12] );
tran (\sa_count[15][63] , \sa_count[15].r.part1[31] );
tran (\sa_count[15][63] , \sa_count[15].f.unused[13] );
tran (\sa_count[16][0] , \sa_count[16].r.part0[0] );
tran (\sa_count[16][0] , \sa_count[16].f.lower[0] );
tran (\sa_count[16][1] , \sa_count[16].r.part0[1] );
tran (\sa_count[16][1] , \sa_count[16].f.lower[1] );
tran (\sa_count[16][2] , \sa_count[16].r.part0[2] );
tran (\sa_count[16][2] , \sa_count[16].f.lower[2] );
tran (\sa_count[16][3] , \sa_count[16].r.part0[3] );
tran (\sa_count[16][3] , \sa_count[16].f.lower[3] );
tran (\sa_count[16][4] , \sa_count[16].r.part0[4] );
tran (\sa_count[16][4] , \sa_count[16].f.lower[4] );
tran (\sa_count[16][5] , \sa_count[16].r.part0[5] );
tran (\sa_count[16][5] , \sa_count[16].f.lower[5] );
tran (\sa_count[16][6] , \sa_count[16].r.part0[6] );
tran (\sa_count[16][6] , \sa_count[16].f.lower[6] );
tran (\sa_count[16][7] , \sa_count[16].r.part0[7] );
tran (\sa_count[16][7] , \sa_count[16].f.lower[7] );
tran (\sa_count[16][8] , \sa_count[16].r.part0[8] );
tran (\sa_count[16][8] , \sa_count[16].f.lower[8] );
tran (\sa_count[16][9] , \sa_count[16].r.part0[9] );
tran (\sa_count[16][9] , \sa_count[16].f.lower[9] );
tran (\sa_count[16][10] , \sa_count[16].r.part0[10] );
tran (\sa_count[16][10] , \sa_count[16].f.lower[10] );
tran (\sa_count[16][11] , \sa_count[16].r.part0[11] );
tran (\sa_count[16][11] , \sa_count[16].f.lower[11] );
tran (\sa_count[16][12] , \sa_count[16].r.part0[12] );
tran (\sa_count[16][12] , \sa_count[16].f.lower[12] );
tran (\sa_count[16][13] , \sa_count[16].r.part0[13] );
tran (\sa_count[16][13] , \sa_count[16].f.lower[13] );
tran (\sa_count[16][14] , \sa_count[16].r.part0[14] );
tran (\sa_count[16][14] , \sa_count[16].f.lower[14] );
tran (\sa_count[16][15] , \sa_count[16].r.part0[15] );
tran (\sa_count[16][15] , \sa_count[16].f.lower[15] );
tran (\sa_count[16][16] , \sa_count[16].r.part0[16] );
tran (\sa_count[16][16] , \sa_count[16].f.lower[16] );
tran (\sa_count[16][17] , \sa_count[16].r.part0[17] );
tran (\sa_count[16][17] , \sa_count[16].f.lower[17] );
tran (\sa_count[16][18] , \sa_count[16].r.part0[18] );
tran (\sa_count[16][18] , \sa_count[16].f.lower[18] );
tran (\sa_count[16][19] , \sa_count[16].r.part0[19] );
tran (\sa_count[16][19] , \sa_count[16].f.lower[19] );
tran (\sa_count[16][20] , \sa_count[16].r.part0[20] );
tran (\sa_count[16][20] , \sa_count[16].f.lower[20] );
tran (\sa_count[16][21] , \sa_count[16].r.part0[21] );
tran (\sa_count[16][21] , \sa_count[16].f.lower[21] );
tran (\sa_count[16][22] , \sa_count[16].r.part0[22] );
tran (\sa_count[16][22] , \sa_count[16].f.lower[22] );
tran (\sa_count[16][23] , \sa_count[16].r.part0[23] );
tran (\sa_count[16][23] , \sa_count[16].f.lower[23] );
tran (\sa_count[16][24] , \sa_count[16].r.part0[24] );
tran (\sa_count[16][24] , \sa_count[16].f.lower[24] );
tran (\sa_count[16][25] , \sa_count[16].r.part0[25] );
tran (\sa_count[16][25] , \sa_count[16].f.lower[25] );
tran (\sa_count[16][26] , \sa_count[16].r.part0[26] );
tran (\sa_count[16][26] , \sa_count[16].f.lower[26] );
tran (\sa_count[16][27] , \sa_count[16].r.part0[27] );
tran (\sa_count[16][27] , \sa_count[16].f.lower[27] );
tran (\sa_count[16][28] , \sa_count[16].r.part0[28] );
tran (\sa_count[16][28] , \sa_count[16].f.lower[28] );
tran (\sa_count[16][29] , \sa_count[16].r.part0[29] );
tran (\sa_count[16][29] , \sa_count[16].f.lower[29] );
tran (\sa_count[16][30] , \sa_count[16].r.part0[30] );
tran (\sa_count[16][30] , \sa_count[16].f.lower[30] );
tran (\sa_count[16][31] , \sa_count[16].r.part0[31] );
tran (\sa_count[16][31] , \sa_count[16].f.lower[31] );
tran (\sa_count[16][32] , \sa_count[16].r.part1[0] );
tran (\sa_count[16][32] , \sa_count[16].f.upper[0] );
tran (\sa_count[16][33] , \sa_count[16].r.part1[1] );
tran (\sa_count[16][33] , \sa_count[16].f.upper[1] );
tran (\sa_count[16][34] , \sa_count[16].r.part1[2] );
tran (\sa_count[16][34] , \sa_count[16].f.upper[2] );
tran (\sa_count[16][35] , \sa_count[16].r.part1[3] );
tran (\sa_count[16][35] , \sa_count[16].f.upper[3] );
tran (\sa_count[16][36] , \sa_count[16].r.part1[4] );
tran (\sa_count[16][36] , \sa_count[16].f.upper[4] );
tran (\sa_count[16][37] , \sa_count[16].r.part1[5] );
tran (\sa_count[16][37] , \sa_count[16].f.upper[5] );
tran (\sa_count[16][38] , \sa_count[16].r.part1[6] );
tran (\sa_count[16][38] , \sa_count[16].f.upper[6] );
tran (\sa_count[16][39] , \sa_count[16].r.part1[7] );
tran (\sa_count[16][39] , \sa_count[16].f.upper[7] );
tran (\sa_count[16][40] , \sa_count[16].r.part1[8] );
tran (\sa_count[16][40] , \sa_count[16].f.upper[8] );
tran (\sa_count[16][41] , \sa_count[16].r.part1[9] );
tran (\sa_count[16][41] , \sa_count[16].f.upper[9] );
tran (\sa_count[16][42] , \sa_count[16].r.part1[10] );
tran (\sa_count[16][42] , \sa_count[16].f.upper[10] );
tran (\sa_count[16][43] , \sa_count[16].r.part1[11] );
tran (\sa_count[16][43] , \sa_count[16].f.upper[11] );
tran (\sa_count[16][44] , \sa_count[16].r.part1[12] );
tran (\sa_count[16][44] , \sa_count[16].f.upper[12] );
tran (\sa_count[16][45] , \sa_count[16].r.part1[13] );
tran (\sa_count[16][45] , \sa_count[16].f.upper[13] );
tran (\sa_count[16][46] , \sa_count[16].r.part1[14] );
tran (\sa_count[16][46] , \sa_count[16].f.upper[14] );
tran (\sa_count[16][47] , \sa_count[16].r.part1[15] );
tran (\sa_count[16][47] , \sa_count[16].f.upper[15] );
tran (\sa_count[16][48] , \sa_count[16].r.part1[16] );
tran (\sa_count[16][48] , \sa_count[16].f.upper[16] );
tran (\sa_count[16][49] , \sa_count[16].r.part1[17] );
tran (\sa_count[16][49] , \sa_count[16].f.upper[17] );
tran (\sa_count[16][50] , \sa_count[16].r.part1[18] );
tran (\sa_count[16][50] , \sa_count[16].f.unused[0] );
tran (\sa_count[16][51] , \sa_count[16].r.part1[19] );
tran (\sa_count[16][51] , \sa_count[16].f.unused[1] );
tran (\sa_count[16][52] , \sa_count[16].r.part1[20] );
tran (\sa_count[16][52] , \sa_count[16].f.unused[2] );
tran (\sa_count[16][53] , \sa_count[16].r.part1[21] );
tran (\sa_count[16][53] , \sa_count[16].f.unused[3] );
tran (\sa_count[16][54] , \sa_count[16].r.part1[22] );
tran (\sa_count[16][54] , \sa_count[16].f.unused[4] );
tran (\sa_count[16][55] , \sa_count[16].r.part1[23] );
tran (\sa_count[16][55] , \sa_count[16].f.unused[5] );
tran (\sa_count[16][56] , \sa_count[16].r.part1[24] );
tran (\sa_count[16][56] , \sa_count[16].f.unused[6] );
tran (\sa_count[16][57] , \sa_count[16].r.part1[25] );
tran (\sa_count[16][57] , \sa_count[16].f.unused[7] );
tran (\sa_count[16][58] , \sa_count[16].r.part1[26] );
tran (\sa_count[16][58] , \sa_count[16].f.unused[8] );
tran (\sa_count[16][59] , \sa_count[16].r.part1[27] );
tran (\sa_count[16][59] , \sa_count[16].f.unused[9] );
tran (\sa_count[16][60] , \sa_count[16].r.part1[28] );
tran (\sa_count[16][60] , \sa_count[16].f.unused[10] );
tran (\sa_count[16][61] , \sa_count[16].r.part1[29] );
tran (\sa_count[16][61] , \sa_count[16].f.unused[11] );
tran (\sa_count[16][62] , \sa_count[16].r.part1[30] );
tran (\sa_count[16][62] , \sa_count[16].f.unused[12] );
tran (\sa_count[16][63] , \sa_count[16].r.part1[31] );
tran (\sa_count[16][63] , \sa_count[16].f.unused[13] );
tran (\sa_count[17][0] , \sa_count[17].r.part0[0] );
tran (\sa_count[17][0] , \sa_count[17].f.lower[0] );
tran (\sa_count[17][1] , \sa_count[17].r.part0[1] );
tran (\sa_count[17][1] , \sa_count[17].f.lower[1] );
tran (\sa_count[17][2] , \sa_count[17].r.part0[2] );
tran (\sa_count[17][2] , \sa_count[17].f.lower[2] );
tran (\sa_count[17][3] , \sa_count[17].r.part0[3] );
tran (\sa_count[17][3] , \sa_count[17].f.lower[3] );
tran (\sa_count[17][4] , \sa_count[17].r.part0[4] );
tran (\sa_count[17][4] , \sa_count[17].f.lower[4] );
tran (\sa_count[17][5] , \sa_count[17].r.part0[5] );
tran (\sa_count[17][5] , \sa_count[17].f.lower[5] );
tran (\sa_count[17][6] , \sa_count[17].r.part0[6] );
tran (\sa_count[17][6] , \sa_count[17].f.lower[6] );
tran (\sa_count[17][7] , \sa_count[17].r.part0[7] );
tran (\sa_count[17][7] , \sa_count[17].f.lower[7] );
tran (\sa_count[17][8] , \sa_count[17].r.part0[8] );
tran (\sa_count[17][8] , \sa_count[17].f.lower[8] );
tran (\sa_count[17][9] , \sa_count[17].r.part0[9] );
tran (\sa_count[17][9] , \sa_count[17].f.lower[9] );
tran (\sa_count[17][10] , \sa_count[17].r.part0[10] );
tran (\sa_count[17][10] , \sa_count[17].f.lower[10] );
tran (\sa_count[17][11] , \sa_count[17].r.part0[11] );
tran (\sa_count[17][11] , \sa_count[17].f.lower[11] );
tran (\sa_count[17][12] , \sa_count[17].r.part0[12] );
tran (\sa_count[17][12] , \sa_count[17].f.lower[12] );
tran (\sa_count[17][13] , \sa_count[17].r.part0[13] );
tran (\sa_count[17][13] , \sa_count[17].f.lower[13] );
tran (\sa_count[17][14] , \sa_count[17].r.part0[14] );
tran (\sa_count[17][14] , \sa_count[17].f.lower[14] );
tran (\sa_count[17][15] , \sa_count[17].r.part0[15] );
tran (\sa_count[17][15] , \sa_count[17].f.lower[15] );
tran (\sa_count[17][16] , \sa_count[17].r.part0[16] );
tran (\sa_count[17][16] , \sa_count[17].f.lower[16] );
tran (\sa_count[17][17] , \sa_count[17].r.part0[17] );
tran (\sa_count[17][17] , \sa_count[17].f.lower[17] );
tran (\sa_count[17][18] , \sa_count[17].r.part0[18] );
tran (\sa_count[17][18] , \sa_count[17].f.lower[18] );
tran (\sa_count[17][19] , \sa_count[17].r.part0[19] );
tran (\sa_count[17][19] , \sa_count[17].f.lower[19] );
tran (\sa_count[17][20] , \sa_count[17].r.part0[20] );
tran (\sa_count[17][20] , \sa_count[17].f.lower[20] );
tran (\sa_count[17][21] , \sa_count[17].r.part0[21] );
tran (\sa_count[17][21] , \sa_count[17].f.lower[21] );
tran (\sa_count[17][22] , \sa_count[17].r.part0[22] );
tran (\sa_count[17][22] , \sa_count[17].f.lower[22] );
tran (\sa_count[17][23] , \sa_count[17].r.part0[23] );
tran (\sa_count[17][23] , \sa_count[17].f.lower[23] );
tran (\sa_count[17][24] , \sa_count[17].r.part0[24] );
tran (\sa_count[17][24] , \sa_count[17].f.lower[24] );
tran (\sa_count[17][25] , \sa_count[17].r.part0[25] );
tran (\sa_count[17][25] , \sa_count[17].f.lower[25] );
tran (\sa_count[17][26] , \sa_count[17].r.part0[26] );
tran (\sa_count[17][26] , \sa_count[17].f.lower[26] );
tran (\sa_count[17][27] , \sa_count[17].r.part0[27] );
tran (\sa_count[17][27] , \sa_count[17].f.lower[27] );
tran (\sa_count[17][28] , \sa_count[17].r.part0[28] );
tran (\sa_count[17][28] , \sa_count[17].f.lower[28] );
tran (\sa_count[17][29] , \sa_count[17].r.part0[29] );
tran (\sa_count[17][29] , \sa_count[17].f.lower[29] );
tran (\sa_count[17][30] , \sa_count[17].r.part0[30] );
tran (\sa_count[17][30] , \sa_count[17].f.lower[30] );
tran (\sa_count[17][31] , \sa_count[17].r.part0[31] );
tran (\sa_count[17][31] , \sa_count[17].f.lower[31] );
tran (\sa_count[17][32] , \sa_count[17].r.part1[0] );
tran (\sa_count[17][32] , \sa_count[17].f.upper[0] );
tran (\sa_count[17][33] , \sa_count[17].r.part1[1] );
tran (\sa_count[17][33] , \sa_count[17].f.upper[1] );
tran (\sa_count[17][34] , \sa_count[17].r.part1[2] );
tran (\sa_count[17][34] , \sa_count[17].f.upper[2] );
tran (\sa_count[17][35] , \sa_count[17].r.part1[3] );
tran (\sa_count[17][35] , \sa_count[17].f.upper[3] );
tran (\sa_count[17][36] , \sa_count[17].r.part1[4] );
tran (\sa_count[17][36] , \sa_count[17].f.upper[4] );
tran (\sa_count[17][37] , \sa_count[17].r.part1[5] );
tran (\sa_count[17][37] , \sa_count[17].f.upper[5] );
tran (\sa_count[17][38] , \sa_count[17].r.part1[6] );
tran (\sa_count[17][38] , \sa_count[17].f.upper[6] );
tran (\sa_count[17][39] , \sa_count[17].r.part1[7] );
tran (\sa_count[17][39] , \sa_count[17].f.upper[7] );
tran (\sa_count[17][40] , \sa_count[17].r.part1[8] );
tran (\sa_count[17][40] , \sa_count[17].f.upper[8] );
tran (\sa_count[17][41] , \sa_count[17].r.part1[9] );
tran (\sa_count[17][41] , \sa_count[17].f.upper[9] );
tran (\sa_count[17][42] , \sa_count[17].r.part1[10] );
tran (\sa_count[17][42] , \sa_count[17].f.upper[10] );
tran (\sa_count[17][43] , \sa_count[17].r.part1[11] );
tran (\sa_count[17][43] , \sa_count[17].f.upper[11] );
tran (\sa_count[17][44] , \sa_count[17].r.part1[12] );
tran (\sa_count[17][44] , \sa_count[17].f.upper[12] );
tran (\sa_count[17][45] , \sa_count[17].r.part1[13] );
tran (\sa_count[17][45] , \sa_count[17].f.upper[13] );
tran (\sa_count[17][46] , \sa_count[17].r.part1[14] );
tran (\sa_count[17][46] , \sa_count[17].f.upper[14] );
tran (\sa_count[17][47] , \sa_count[17].r.part1[15] );
tran (\sa_count[17][47] , \sa_count[17].f.upper[15] );
tran (\sa_count[17][48] , \sa_count[17].r.part1[16] );
tran (\sa_count[17][48] , \sa_count[17].f.upper[16] );
tran (\sa_count[17][49] , \sa_count[17].r.part1[17] );
tran (\sa_count[17][49] , \sa_count[17].f.upper[17] );
tran (\sa_count[17][50] , \sa_count[17].r.part1[18] );
tran (\sa_count[17][50] , \sa_count[17].f.unused[0] );
tran (\sa_count[17][51] , \sa_count[17].r.part1[19] );
tran (\sa_count[17][51] , \sa_count[17].f.unused[1] );
tran (\sa_count[17][52] , \sa_count[17].r.part1[20] );
tran (\sa_count[17][52] , \sa_count[17].f.unused[2] );
tran (\sa_count[17][53] , \sa_count[17].r.part1[21] );
tran (\sa_count[17][53] , \sa_count[17].f.unused[3] );
tran (\sa_count[17][54] , \sa_count[17].r.part1[22] );
tran (\sa_count[17][54] , \sa_count[17].f.unused[4] );
tran (\sa_count[17][55] , \sa_count[17].r.part1[23] );
tran (\sa_count[17][55] , \sa_count[17].f.unused[5] );
tran (\sa_count[17][56] , \sa_count[17].r.part1[24] );
tran (\sa_count[17][56] , \sa_count[17].f.unused[6] );
tran (\sa_count[17][57] , \sa_count[17].r.part1[25] );
tran (\sa_count[17][57] , \sa_count[17].f.unused[7] );
tran (\sa_count[17][58] , \sa_count[17].r.part1[26] );
tran (\sa_count[17][58] , \sa_count[17].f.unused[8] );
tran (\sa_count[17][59] , \sa_count[17].r.part1[27] );
tran (\sa_count[17][59] , \sa_count[17].f.unused[9] );
tran (\sa_count[17][60] , \sa_count[17].r.part1[28] );
tran (\sa_count[17][60] , \sa_count[17].f.unused[10] );
tran (\sa_count[17][61] , \sa_count[17].r.part1[29] );
tran (\sa_count[17][61] , \sa_count[17].f.unused[11] );
tran (\sa_count[17][62] , \sa_count[17].r.part1[30] );
tran (\sa_count[17][62] , \sa_count[17].f.unused[12] );
tran (\sa_count[17][63] , \sa_count[17].r.part1[31] );
tran (\sa_count[17][63] , \sa_count[17].f.unused[13] );
tran (\sa_count[18][0] , \sa_count[18].r.part0[0] );
tran (\sa_count[18][0] , \sa_count[18].f.lower[0] );
tran (\sa_count[18][1] , \sa_count[18].r.part0[1] );
tran (\sa_count[18][1] , \sa_count[18].f.lower[1] );
tran (\sa_count[18][2] , \sa_count[18].r.part0[2] );
tran (\sa_count[18][2] , \sa_count[18].f.lower[2] );
tran (\sa_count[18][3] , \sa_count[18].r.part0[3] );
tran (\sa_count[18][3] , \sa_count[18].f.lower[3] );
tran (\sa_count[18][4] , \sa_count[18].r.part0[4] );
tran (\sa_count[18][4] , \sa_count[18].f.lower[4] );
tran (\sa_count[18][5] , \sa_count[18].r.part0[5] );
tran (\sa_count[18][5] , \sa_count[18].f.lower[5] );
tran (\sa_count[18][6] , \sa_count[18].r.part0[6] );
tran (\sa_count[18][6] , \sa_count[18].f.lower[6] );
tran (\sa_count[18][7] , \sa_count[18].r.part0[7] );
tran (\sa_count[18][7] , \sa_count[18].f.lower[7] );
tran (\sa_count[18][8] , \sa_count[18].r.part0[8] );
tran (\sa_count[18][8] , \sa_count[18].f.lower[8] );
tran (\sa_count[18][9] , \sa_count[18].r.part0[9] );
tran (\sa_count[18][9] , \sa_count[18].f.lower[9] );
tran (\sa_count[18][10] , \sa_count[18].r.part0[10] );
tran (\sa_count[18][10] , \sa_count[18].f.lower[10] );
tran (\sa_count[18][11] , \sa_count[18].r.part0[11] );
tran (\sa_count[18][11] , \sa_count[18].f.lower[11] );
tran (\sa_count[18][12] , \sa_count[18].r.part0[12] );
tran (\sa_count[18][12] , \sa_count[18].f.lower[12] );
tran (\sa_count[18][13] , \sa_count[18].r.part0[13] );
tran (\sa_count[18][13] , \sa_count[18].f.lower[13] );
tran (\sa_count[18][14] , \sa_count[18].r.part0[14] );
tran (\sa_count[18][14] , \sa_count[18].f.lower[14] );
tran (\sa_count[18][15] , \sa_count[18].r.part0[15] );
tran (\sa_count[18][15] , \sa_count[18].f.lower[15] );
tran (\sa_count[18][16] , \sa_count[18].r.part0[16] );
tran (\sa_count[18][16] , \sa_count[18].f.lower[16] );
tran (\sa_count[18][17] , \sa_count[18].r.part0[17] );
tran (\sa_count[18][17] , \sa_count[18].f.lower[17] );
tran (\sa_count[18][18] , \sa_count[18].r.part0[18] );
tran (\sa_count[18][18] , \sa_count[18].f.lower[18] );
tran (\sa_count[18][19] , \sa_count[18].r.part0[19] );
tran (\sa_count[18][19] , \sa_count[18].f.lower[19] );
tran (\sa_count[18][20] , \sa_count[18].r.part0[20] );
tran (\sa_count[18][20] , \sa_count[18].f.lower[20] );
tran (\sa_count[18][21] , \sa_count[18].r.part0[21] );
tran (\sa_count[18][21] , \sa_count[18].f.lower[21] );
tran (\sa_count[18][22] , \sa_count[18].r.part0[22] );
tran (\sa_count[18][22] , \sa_count[18].f.lower[22] );
tran (\sa_count[18][23] , \sa_count[18].r.part0[23] );
tran (\sa_count[18][23] , \sa_count[18].f.lower[23] );
tran (\sa_count[18][24] , \sa_count[18].r.part0[24] );
tran (\sa_count[18][24] , \sa_count[18].f.lower[24] );
tran (\sa_count[18][25] , \sa_count[18].r.part0[25] );
tran (\sa_count[18][25] , \sa_count[18].f.lower[25] );
tran (\sa_count[18][26] , \sa_count[18].r.part0[26] );
tran (\sa_count[18][26] , \sa_count[18].f.lower[26] );
tran (\sa_count[18][27] , \sa_count[18].r.part0[27] );
tran (\sa_count[18][27] , \sa_count[18].f.lower[27] );
tran (\sa_count[18][28] , \sa_count[18].r.part0[28] );
tran (\sa_count[18][28] , \sa_count[18].f.lower[28] );
tran (\sa_count[18][29] , \sa_count[18].r.part0[29] );
tran (\sa_count[18][29] , \sa_count[18].f.lower[29] );
tran (\sa_count[18][30] , \sa_count[18].r.part0[30] );
tran (\sa_count[18][30] , \sa_count[18].f.lower[30] );
tran (\sa_count[18][31] , \sa_count[18].r.part0[31] );
tran (\sa_count[18][31] , \sa_count[18].f.lower[31] );
tran (\sa_count[18][32] , \sa_count[18].r.part1[0] );
tran (\sa_count[18][32] , \sa_count[18].f.upper[0] );
tran (\sa_count[18][33] , \sa_count[18].r.part1[1] );
tran (\sa_count[18][33] , \sa_count[18].f.upper[1] );
tran (\sa_count[18][34] , \sa_count[18].r.part1[2] );
tran (\sa_count[18][34] , \sa_count[18].f.upper[2] );
tran (\sa_count[18][35] , \sa_count[18].r.part1[3] );
tran (\sa_count[18][35] , \sa_count[18].f.upper[3] );
tran (\sa_count[18][36] , \sa_count[18].r.part1[4] );
tran (\sa_count[18][36] , \sa_count[18].f.upper[4] );
tran (\sa_count[18][37] , \sa_count[18].r.part1[5] );
tran (\sa_count[18][37] , \sa_count[18].f.upper[5] );
tran (\sa_count[18][38] , \sa_count[18].r.part1[6] );
tran (\sa_count[18][38] , \sa_count[18].f.upper[6] );
tran (\sa_count[18][39] , \sa_count[18].r.part1[7] );
tran (\sa_count[18][39] , \sa_count[18].f.upper[7] );
tran (\sa_count[18][40] , \sa_count[18].r.part1[8] );
tran (\sa_count[18][40] , \sa_count[18].f.upper[8] );
tran (\sa_count[18][41] , \sa_count[18].r.part1[9] );
tran (\sa_count[18][41] , \sa_count[18].f.upper[9] );
tran (\sa_count[18][42] , \sa_count[18].r.part1[10] );
tran (\sa_count[18][42] , \sa_count[18].f.upper[10] );
tran (\sa_count[18][43] , \sa_count[18].r.part1[11] );
tran (\sa_count[18][43] , \sa_count[18].f.upper[11] );
tran (\sa_count[18][44] , \sa_count[18].r.part1[12] );
tran (\sa_count[18][44] , \sa_count[18].f.upper[12] );
tran (\sa_count[18][45] , \sa_count[18].r.part1[13] );
tran (\sa_count[18][45] , \sa_count[18].f.upper[13] );
tran (\sa_count[18][46] , \sa_count[18].r.part1[14] );
tran (\sa_count[18][46] , \sa_count[18].f.upper[14] );
tran (\sa_count[18][47] , \sa_count[18].r.part1[15] );
tran (\sa_count[18][47] , \sa_count[18].f.upper[15] );
tran (\sa_count[18][48] , \sa_count[18].r.part1[16] );
tran (\sa_count[18][48] , \sa_count[18].f.upper[16] );
tran (\sa_count[18][49] , \sa_count[18].r.part1[17] );
tran (\sa_count[18][49] , \sa_count[18].f.upper[17] );
tran (\sa_count[18][50] , \sa_count[18].r.part1[18] );
tran (\sa_count[18][50] , \sa_count[18].f.unused[0] );
tran (\sa_count[18][51] , \sa_count[18].r.part1[19] );
tran (\sa_count[18][51] , \sa_count[18].f.unused[1] );
tran (\sa_count[18][52] , \sa_count[18].r.part1[20] );
tran (\sa_count[18][52] , \sa_count[18].f.unused[2] );
tran (\sa_count[18][53] , \sa_count[18].r.part1[21] );
tran (\sa_count[18][53] , \sa_count[18].f.unused[3] );
tran (\sa_count[18][54] , \sa_count[18].r.part1[22] );
tran (\sa_count[18][54] , \sa_count[18].f.unused[4] );
tran (\sa_count[18][55] , \sa_count[18].r.part1[23] );
tran (\sa_count[18][55] , \sa_count[18].f.unused[5] );
tran (\sa_count[18][56] , \sa_count[18].r.part1[24] );
tran (\sa_count[18][56] , \sa_count[18].f.unused[6] );
tran (\sa_count[18][57] , \sa_count[18].r.part1[25] );
tran (\sa_count[18][57] , \sa_count[18].f.unused[7] );
tran (\sa_count[18][58] , \sa_count[18].r.part1[26] );
tran (\sa_count[18][58] , \sa_count[18].f.unused[8] );
tran (\sa_count[18][59] , \sa_count[18].r.part1[27] );
tran (\sa_count[18][59] , \sa_count[18].f.unused[9] );
tran (\sa_count[18][60] , \sa_count[18].r.part1[28] );
tran (\sa_count[18][60] , \sa_count[18].f.unused[10] );
tran (\sa_count[18][61] , \sa_count[18].r.part1[29] );
tran (\sa_count[18][61] , \sa_count[18].f.unused[11] );
tran (\sa_count[18][62] , \sa_count[18].r.part1[30] );
tran (\sa_count[18][62] , \sa_count[18].f.unused[12] );
tran (\sa_count[18][63] , \sa_count[18].r.part1[31] );
tran (\sa_count[18][63] , \sa_count[18].f.unused[13] );
tran (\sa_count[19][0] , \sa_count[19].r.part0[0] );
tran (\sa_count[19][0] , \sa_count[19].f.lower[0] );
tran (\sa_count[19][1] , \sa_count[19].r.part0[1] );
tran (\sa_count[19][1] , \sa_count[19].f.lower[1] );
tran (\sa_count[19][2] , \sa_count[19].r.part0[2] );
tran (\sa_count[19][2] , \sa_count[19].f.lower[2] );
tran (\sa_count[19][3] , \sa_count[19].r.part0[3] );
tran (\sa_count[19][3] , \sa_count[19].f.lower[3] );
tran (\sa_count[19][4] , \sa_count[19].r.part0[4] );
tran (\sa_count[19][4] , \sa_count[19].f.lower[4] );
tran (\sa_count[19][5] , \sa_count[19].r.part0[5] );
tran (\sa_count[19][5] , \sa_count[19].f.lower[5] );
tran (\sa_count[19][6] , \sa_count[19].r.part0[6] );
tran (\sa_count[19][6] , \sa_count[19].f.lower[6] );
tran (\sa_count[19][7] , \sa_count[19].r.part0[7] );
tran (\sa_count[19][7] , \sa_count[19].f.lower[7] );
tran (\sa_count[19][8] , \sa_count[19].r.part0[8] );
tran (\sa_count[19][8] , \sa_count[19].f.lower[8] );
tran (\sa_count[19][9] , \sa_count[19].r.part0[9] );
tran (\sa_count[19][9] , \sa_count[19].f.lower[9] );
tran (\sa_count[19][10] , \sa_count[19].r.part0[10] );
tran (\sa_count[19][10] , \sa_count[19].f.lower[10] );
tran (\sa_count[19][11] , \sa_count[19].r.part0[11] );
tran (\sa_count[19][11] , \sa_count[19].f.lower[11] );
tran (\sa_count[19][12] , \sa_count[19].r.part0[12] );
tran (\sa_count[19][12] , \sa_count[19].f.lower[12] );
tran (\sa_count[19][13] , \sa_count[19].r.part0[13] );
tran (\sa_count[19][13] , \sa_count[19].f.lower[13] );
tran (\sa_count[19][14] , \sa_count[19].r.part0[14] );
tran (\sa_count[19][14] , \sa_count[19].f.lower[14] );
tran (\sa_count[19][15] , \sa_count[19].r.part0[15] );
tran (\sa_count[19][15] , \sa_count[19].f.lower[15] );
tran (\sa_count[19][16] , \sa_count[19].r.part0[16] );
tran (\sa_count[19][16] , \sa_count[19].f.lower[16] );
tran (\sa_count[19][17] , \sa_count[19].r.part0[17] );
tran (\sa_count[19][17] , \sa_count[19].f.lower[17] );
tran (\sa_count[19][18] , \sa_count[19].r.part0[18] );
tran (\sa_count[19][18] , \sa_count[19].f.lower[18] );
tran (\sa_count[19][19] , \sa_count[19].r.part0[19] );
tran (\sa_count[19][19] , \sa_count[19].f.lower[19] );
tran (\sa_count[19][20] , \sa_count[19].r.part0[20] );
tran (\sa_count[19][20] , \sa_count[19].f.lower[20] );
tran (\sa_count[19][21] , \sa_count[19].r.part0[21] );
tran (\sa_count[19][21] , \sa_count[19].f.lower[21] );
tran (\sa_count[19][22] , \sa_count[19].r.part0[22] );
tran (\sa_count[19][22] , \sa_count[19].f.lower[22] );
tran (\sa_count[19][23] , \sa_count[19].r.part0[23] );
tran (\sa_count[19][23] , \sa_count[19].f.lower[23] );
tran (\sa_count[19][24] , \sa_count[19].r.part0[24] );
tran (\sa_count[19][24] , \sa_count[19].f.lower[24] );
tran (\sa_count[19][25] , \sa_count[19].r.part0[25] );
tran (\sa_count[19][25] , \sa_count[19].f.lower[25] );
tran (\sa_count[19][26] , \sa_count[19].r.part0[26] );
tran (\sa_count[19][26] , \sa_count[19].f.lower[26] );
tran (\sa_count[19][27] , \sa_count[19].r.part0[27] );
tran (\sa_count[19][27] , \sa_count[19].f.lower[27] );
tran (\sa_count[19][28] , \sa_count[19].r.part0[28] );
tran (\sa_count[19][28] , \sa_count[19].f.lower[28] );
tran (\sa_count[19][29] , \sa_count[19].r.part0[29] );
tran (\sa_count[19][29] , \sa_count[19].f.lower[29] );
tran (\sa_count[19][30] , \sa_count[19].r.part0[30] );
tran (\sa_count[19][30] , \sa_count[19].f.lower[30] );
tran (\sa_count[19][31] , \sa_count[19].r.part0[31] );
tran (\sa_count[19][31] , \sa_count[19].f.lower[31] );
tran (\sa_count[19][32] , \sa_count[19].r.part1[0] );
tran (\sa_count[19][32] , \sa_count[19].f.upper[0] );
tran (\sa_count[19][33] , \sa_count[19].r.part1[1] );
tran (\sa_count[19][33] , \sa_count[19].f.upper[1] );
tran (\sa_count[19][34] , \sa_count[19].r.part1[2] );
tran (\sa_count[19][34] , \sa_count[19].f.upper[2] );
tran (\sa_count[19][35] , \sa_count[19].r.part1[3] );
tran (\sa_count[19][35] , \sa_count[19].f.upper[3] );
tran (\sa_count[19][36] , \sa_count[19].r.part1[4] );
tran (\sa_count[19][36] , \sa_count[19].f.upper[4] );
tran (\sa_count[19][37] , \sa_count[19].r.part1[5] );
tran (\sa_count[19][37] , \sa_count[19].f.upper[5] );
tran (\sa_count[19][38] , \sa_count[19].r.part1[6] );
tran (\sa_count[19][38] , \sa_count[19].f.upper[6] );
tran (\sa_count[19][39] , \sa_count[19].r.part1[7] );
tran (\sa_count[19][39] , \sa_count[19].f.upper[7] );
tran (\sa_count[19][40] , \sa_count[19].r.part1[8] );
tran (\sa_count[19][40] , \sa_count[19].f.upper[8] );
tran (\sa_count[19][41] , \sa_count[19].r.part1[9] );
tran (\sa_count[19][41] , \sa_count[19].f.upper[9] );
tran (\sa_count[19][42] , \sa_count[19].r.part1[10] );
tran (\sa_count[19][42] , \sa_count[19].f.upper[10] );
tran (\sa_count[19][43] , \sa_count[19].r.part1[11] );
tran (\sa_count[19][43] , \sa_count[19].f.upper[11] );
tran (\sa_count[19][44] , \sa_count[19].r.part1[12] );
tran (\sa_count[19][44] , \sa_count[19].f.upper[12] );
tran (\sa_count[19][45] , \sa_count[19].r.part1[13] );
tran (\sa_count[19][45] , \sa_count[19].f.upper[13] );
tran (\sa_count[19][46] , \sa_count[19].r.part1[14] );
tran (\sa_count[19][46] , \sa_count[19].f.upper[14] );
tran (\sa_count[19][47] , \sa_count[19].r.part1[15] );
tran (\sa_count[19][47] , \sa_count[19].f.upper[15] );
tran (\sa_count[19][48] , \sa_count[19].r.part1[16] );
tran (\sa_count[19][48] , \sa_count[19].f.upper[16] );
tran (\sa_count[19][49] , \sa_count[19].r.part1[17] );
tran (\sa_count[19][49] , \sa_count[19].f.upper[17] );
tran (\sa_count[19][50] , \sa_count[19].r.part1[18] );
tran (\sa_count[19][50] , \sa_count[19].f.unused[0] );
tran (\sa_count[19][51] , \sa_count[19].r.part1[19] );
tran (\sa_count[19][51] , \sa_count[19].f.unused[1] );
tran (\sa_count[19][52] , \sa_count[19].r.part1[20] );
tran (\sa_count[19][52] , \sa_count[19].f.unused[2] );
tran (\sa_count[19][53] , \sa_count[19].r.part1[21] );
tran (\sa_count[19][53] , \sa_count[19].f.unused[3] );
tran (\sa_count[19][54] , \sa_count[19].r.part1[22] );
tran (\sa_count[19][54] , \sa_count[19].f.unused[4] );
tran (\sa_count[19][55] , \sa_count[19].r.part1[23] );
tran (\sa_count[19][55] , \sa_count[19].f.unused[5] );
tran (\sa_count[19][56] , \sa_count[19].r.part1[24] );
tran (\sa_count[19][56] , \sa_count[19].f.unused[6] );
tran (\sa_count[19][57] , \sa_count[19].r.part1[25] );
tran (\sa_count[19][57] , \sa_count[19].f.unused[7] );
tran (\sa_count[19][58] , \sa_count[19].r.part1[26] );
tran (\sa_count[19][58] , \sa_count[19].f.unused[8] );
tran (\sa_count[19][59] , \sa_count[19].r.part1[27] );
tran (\sa_count[19][59] , \sa_count[19].f.unused[9] );
tran (\sa_count[19][60] , \sa_count[19].r.part1[28] );
tran (\sa_count[19][60] , \sa_count[19].f.unused[10] );
tran (\sa_count[19][61] , \sa_count[19].r.part1[29] );
tran (\sa_count[19][61] , \sa_count[19].f.unused[11] );
tran (\sa_count[19][62] , \sa_count[19].r.part1[30] );
tran (\sa_count[19][62] , \sa_count[19].f.unused[12] );
tran (\sa_count[19][63] , \sa_count[19].r.part1[31] );
tran (\sa_count[19][63] , \sa_count[19].f.unused[13] );
tran (\sa_count[20][0] , \sa_count[20].r.part0[0] );
tran (\sa_count[20][0] , \sa_count[20].f.lower[0] );
tran (\sa_count[20][1] , \sa_count[20].r.part0[1] );
tran (\sa_count[20][1] , \sa_count[20].f.lower[1] );
tran (\sa_count[20][2] , \sa_count[20].r.part0[2] );
tran (\sa_count[20][2] , \sa_count[20].f.lower[2] );
tran (\sa_count[20][3] , \sa_count[20].r.part0[3] );
tran (\sa_count[20][3] , \sa_count[20].f.lower[3] );
tran (\sa_count[20][4] , \sa_count[20].r.part0[4] );
tran (\sa_count[20][4] , \sa_count[20].f.lower[4] );
tran (\sa_count[20][5] , \sa_count[20].r.part0[5] );
tran (\sa_count[20][5] , \sa_count[20].f.lower[5] );
tran (\sa_count[20][6] , \sa_count[20].r.part0[6] );
tran (\sa_count[20][6] , \sa_count[20].f.lower[6] );
tran (\sa_count[20][7] , \sa_count[20].r.part0[7] );
tran (\sa_count[20][7] , \sa_count[20].f.lower[7] );
tran (\sa_count[20][8] , \sa_count[20].r.part0[8] );
tran (\sa_count[20][8] , \sa_count[20].f.lower[8] );
tran (\sa_count[20][9] , \sa_count[20].r.part0[9] );
tran (\sa_count[20][9] , \sa_count[20].f.lower[9] );
tran (\sa_count[20][10] , \sa_count[20].r.part0[10] );
tran (\sa_count[20][10] , \sa_count[20].f.lower[10] );
tran (\sa_count[20][11] , \sa_count[20].r.part0[11] );
tran (\sa_count[20][11] , \sa_count[20].f.lower[11] );
tran (\sa_count[20][12] , \sa_count[20].r.part0[12] );
tran (\sa_count[20][12] , \sa_count[20].f.lower[12] );
tran (\sa_count[20][13] , \sa_count[20].r.part0[13] );
tran (\sa_count[20][13] , \sa_count[20].f.lower[13] );
tran (\sa_count[20][14] , \sa_count[20].r.part0[14] );
tran (\sa_count[20][14] , \sa_count[20].f.lower[14] );
tran (\sa_count[20][15] , \sa_count[20].r.part0[15] );
tran (\sa_count[20][15] , \sa_count[20].f.lower[15] );
tran (\sa_count[20][16] , \sa_count[20].r.part0[16] );
tran (\sa_count[20][16] , \sa_count[20].f.lower[16] );
tran (\sa_count[20][17] , \sa_count[20].r.part0[17] );
tran (\sa_count[20][17] , \sa_count[20].f.lower[17] );
tran (\sa_count[20][18] , \sa_count[20].r.part0[18] );
tran (\sa_count[20][18] , \sa_count[20].f.lower[18] );
tran (\sa_count[20][19] , \sa_count[20].r.part0[19] );
tran (\sa_count[20][19] , \sa_count[20].f.lower[19] );
tran (\sa_count[20][20] , \sa_count[20].r.part0[20] );
tran (\sa_count[20][20] , \sa_count[20].f.lower[20] );
tran (\sa_count[20][21] , \sa_count[20].r.part0[21] );
tran (\sa_count[20][21] , \sa_count[20].f.lower[21] );
tran (\sa_count[20][22] , \sa_count[20].r.part0[22] );
tran (\sa_count[20][22] , \sa_count[20].f.lower[22] );
tran (\sa_count[20][23] , \sa_count[20].r.part0[23] );
tran (\sa_count[20][23] , \sa_count[20].f.lower[23] );
tran (\sa_count[20][24] , \sa_count[20].r.part0[24] );
tran (\sa_count[20][24] , \sa_count[20].f.lower[24] );
tran (\sa_count[20][25] , \sa_count[20].r.part0[25] );
tran (\sa_count[20][25] , \sa_count[20].f.lower[25] );
tran (\sa_count[20][26] , \sa_count[20].r.part0[26] );
tran (\sa_count[20][26] , \sa_count[20].f.lower[26] );
tran (\sa_count[20][27] , \sa_count[20].r.part0[27] );
tran (\sa_count[20][27] , \sa_count[20].f.lower[27] );
tran (\sa_count[20][28] , \sa_count[20].r.part0[28] );
tran (\sa_count[20][28] , \sa_count[20].f.lower[28] );
tran (\sa_count[20][29] , \sa_count[20].r.part0[29] );
tran (\sa_count[20][29] , \sa_count[20].f.lower[29] );
tran (\sa_count[20][30] , \sa_count[20].r.part0[30] );
tran (\sa_count[20][30] , \sa_count[20].f.lower[30] );
tran (\sa_count[20][31] , \sa_count[20].r.part0[31] );
tran (\sa_count[20][31] , \sa_count[20].f.lower[31] );
tran (\sa_count[20][32] , \sa_count[20].r.part1[0] );
tran (\sa_count[20][32] , \sa_count[20].f.upper[0] );
tran (\sa_count[20][33] , \sa_count[20].r.part1[1] );
tran (\sa_count[20][33] , \sa_count[20].f.upper[1] );
tran (\sa_count[20][34] , \sa_count[20].r.part1[2] );
tran (\sa_count[20][34] , \sa_count[20].f.upper[2] );
tran (\sa_count[20][35] , \sa_count[20].r.part1[3] );
tran (\sa_count[20][35] , \sa_count[20].f.upper[3] );
tran (\sa_count[20][36] , \sa_count[20].r.part1[4] );
tran (\sa_count[20][36] , \sa_count[20].f.upper[4] );
tran (\sa_count[20][37] , \sa_count[20].r.part1[5] );
tran (\sa_count[20][37] , \sa_count[20].f.upper[5] );
tran (\sa_count[20][38] , \sa_count[20].r.part1[6] );
tran (\sa_count[20][38] , \sa_count[20].f.upper[6] );
tran (\sa_count[20][39] , \sa_count[20].r.part1[7] );
tran (\sa_count[20][39] , \sa_count[20].f.upper[7] );
tran (\sa_count[20][40] , \sa_count[20].r.part1[8] );
tran (\sa_count[20][40] , \sa_count[20].f.upper[8] );
tran (\sa_count[20][41] , \sa_count[20].r.part1[9] );
tran (\sa_count[20][41] , \sa_count[20].f.upper[9] );
tran (\sa_count[20][42] , \sa_count[20].r.part1[10] );
tran (\sa_count[20][42] , \sa_count[20].f.upper[10] );
tran (\sa_count[20][43] , \sa_count[20].r.part1[11] );
tran (\sa_count[20][43] , \sa_count[20].f.upper[11] );
tran (\sa_count[20][44] , \sa_count[20].r.part1[12] );
tran (\sa_count[20][44] , \sa_count[20].f.upper[12] );
tran (\sa_count[20][45] , \sa_count[20].r.part1[13] );
tran (\sa_count[20][45] , \sa_count[20].f.upper[13] );
tran (\sa_count[20][46] , \sa_count[20].r.part1[14] );
tran (\sa_count[20][46] , \sa_count[20].f.upper[14] );
tran (\sa_count[20][47] , \sa_count[20].r.part1[15] );
tran (\sa_count[20][47] , \sa_count[20].f.upper[15] );
tran (\sa_count[20][48] , \sa_count[20].r.part1[16] );
tran (\sa_count[20][48] , \sa_count[20].f.upper[16] );
tran (\sa_count[20][49] , \sa_count[20].r.part1[17] );
tran (\sa_count[20][49] , \sa_count[20].f.upper[17] );
tran (\sa_count[20][50] , \sa_count[20].r.part1[18] );
tran (\sa_count[20][50] , \sa_count[20].f.unused[0] );
tran (\sa_count[20][51] , \sa_count[20].r.part1[19] );
tran (\sa_count[20][51] , \sa_count[20].f.unused[1] );
tran (\sa_count[20][52] , \sa_count[20].r.part1[20] );
tran (\sa_count[20][52] , \sa_count[20].f.unused[2] );
tran (\sa_count[20][53] , \sa_count[20].r.part1[21] );
tran (\sa_count[20][53] , \sa_count[20].f.unused[3] );
tran (\sa_count[20][54] , \sa_count[20].r.part1[22] );
tran (\sa_count[20][54] , \sa_count[20].f.unused[4] );
tran (\sa_count[20][55] , \sa_count[20].r.part1[23] );
tran (\sa_count[20][55] , \sa_count[20].f.unused[5] );
tran (\sa_count[20][56] , \sa_count[20].r.part1[24] );
tran (\sa_count[20][56] , \sa_count[20].f.unused[6] );
tran (\sa_count[20][57] , \sa_count[20].r.part1[25] );
tran (\sa_count[20][57] , \sa_count[20].f.unused[7] );
tran (\sa_count[20][58] , \sa_count[20].r.part1[26] );
tran (\sa_count[20][58] , \sa_count[20].f.unused[8] );
tran (\sa_count[20][59] , \sa_count[20].r.part1[27] );
tran (\sa_count[20][59] , \sa_count[20].f.unused[9] );
tran (\sa_count[20][60] , \sa_count[20].r.part1[28] );
tran (\sa_count[20][60] , \sa_count[20].f.unused[10] );
tran (\sa_count[20][61] , \sa_count[20].r.part1[29] );
tran (\sa_count[20][61] , \sa_count[20].f.unused[11] );
tran (\sa_count[20][62] , \sa_count[20].r.part1[30] );
tran (\sa_count[20][62] , \sa_count[20].f.unused[12] );
tran (\sa_count[20][63] , \sa_count[20].r.part1[31] );
tran (\sa_count[20][63] , \sa_count[20].f.unused[13] );
tran (\sa_count[21][0] , \sa_count[21].r.part0[0] );
tran (\sa_count[21][0] , \sa_count[21].f.lower[0] );
tran (\sa_count[21][1] , \sa_count[21].r.part0[1] );
tran (\sa_count[21][1] , \sa_count[21].f.lower[1] );
tran (\sa_count[21][2] , \sa_count[21].r.part0[2] );
tran (\sa_count[21][2] , \sa_count[21].f.lower[2] );
tran (\sa_count[21][3] , \sa_count[21].r.part0[3] );
tran (\sa_count[21][3] , \sa_count[21].f.lower[3] );
tran (\sa_count[21][4] , \sa_count[21].r.part0[4] );
tran (\sa_count[21][4] , \sa_count[21].f.lower[4] );
tran (\sa_count[21][5] , \sa_count[21].r.part0[5] );
tran (\sa_count[21][5] , \sa_count[21].f.lower[5] );
tran (\sa_count[21][6] , \sa_count[21].r.part0[6] );
tran (\sa_count[21][6] , \sa_count[21].f.lower[6] );
tran (\sa_count[21][7] , \sa_count[21].r.part0[7] );
tran (\sa_count[21][7] , \sa_count[21].f.lower[7] );
tran (\sa_count[21][8] , \sa_count[21].r.part0[8] );
tran (\sa_count[21][8] , \sa_count[21].f.lower[8] );
tran (\sa_count[21][9] , \sa_count[21].r.part0[9] );
tran (\sa_count[21][9] , \sa_count[21].f.lower[9] );
tran (\sa_count[21][10] , \sa_count[21].r.part0[10] );
tran (\sa_count[21][10] , \sa_count[21].f.lower[10] );
tran (\sa_count[21][11] , \sa_count[21].r.part0[11] );
tran (\sa_count[21][11] , \sa_count[21].f.lower[11] );
tran (\sa_count[21][12] , \sa_count[21].r.part0[12] );
tran (\sa_count[21][12] , \sa_count[21].f.lower[12] );
tran (\sa_count[21][13] , \sa_count[21].r.part0[13] );
tran (\sa_count[21][13] , \sa_count[21].f.lower[13] );
tran (\sa_count[21][14] , \sa_count[21].r.part0[14] );
tran (\sa_count[21][14] , \sa_count[21].f.lower[14] );
tran (\sa_count[21][15] , \sa_count[21].r.part0[15] );
tran (\sa_count[21][15] , \sa_count[21].f.lower[15] );
tran (\sa_count[21][16] , \sa_count[21].r.part0[16] );
tran (\sa_count[21][16] , \sa_count[21].f.lower[16] );
tran (\sa_count[21][17] , \sa_count[21].r.part0[17] );
tran (\sa_count[21][17] , \sa_count[21].f.lower[17] );
tran (\sa_count[21][18] , \sa_count[21].r.part0[18] );
tran (\sa_count[21][18] , \sa_count[21].f.lower[18] );
tran (\sa_count[21][19] , \sa_count[21].r.part0[19] );
tran (\sa_count[21][19] , \sa_count[21].f.lower[19] );
tran (\sa_count[21][20] , \sa_count[21].r.part0[20] );
tran (\sa_count[21][20] , \sa_count[21].f.lower[20] );
tran (\sa_count[21][21] , \sa_count[21].r.part0[21] );
tran (\sa_count[21][21] , \sa_count[21].f.lower[21] );
tran (\sa_count[21][22] , \sa_count[21].r.part0[22] );
tran (\sa_count[21][22] , \sa_count[21].f.lower[22] );
tran (\sa_count[21][23] , \sa_count[21].r.part0[23] );
tran (\sa_count[21][23] , \sa_count[21].f.lower[23] );
tran (\sa_count[21][24] , \sa_count[21].r.part0[24] );
tran (\sa_count[21][24] , \sa_count[21].f.lower[24] );
tran (\sa_count[21][25] , \sa_count[21].r.part0[25] );
tran (\sa_count[21][25] , \sa_count[21].f.lower[25] );
tran (\sa_count[21][26] , \sa_count[21].r.part0[26] );
tran (\sa_count[21][26] , \sa_count[21].f.lower[26] );
tran (\sa_count[21][27] , \sa_count[21].r.part0[27] );
tran (\sa_count[21][27] , \sa_count[21].f.lower[27] );
tran (\sa_count[21][28] , \sa_count[21].r.part0[28] );
tran (\sa_count[21][28] , \sa_count[21].f.lower[28] );
tran (\sa_count[21][29] , \sa_count[21].r.part0[29] );
tran (\sa_count[21][29] , \sa_count[21].f.lower[29] );
tran (\sa_count[21][30] , \sa_count[21].r.part0[30] );
tran (\sa_count[21][30] , \sa_count[21].f.lower[30] );
tran (\sa_count[21][31] , \sa_count[21].r.part0[31] );
tran (\sa_count[21][31] , \sa_count[21].f.lower[31] );
tran (\sa_count[21][32] , \sa_count[21].r.part1[0] );
tran (\sa_count[21][32] , \sa_count[21].f.upper[0] );
tran (\sa_count[21][33] , \sa_count[21].r.part1[1] );
tran (\sa_count[21][33] , \sa_count[21].f.upper[1] );
tran (\sa_count[21][34] , \sa_count[21].r.part1[2] );
tran (\sa_count[21][34] , \sa_count[21].f.upper[2] );
tran (\sa_count[21][35] , \sa_count[21].r.part1[3] );
tran (\sa_count[21][35] , \sa_count[21].f.upper[3] );
tran (\sa_count[21][36] , \sa_count[21].r.part1[4] );
tran (\sa_count[21][36] , \sa_count[21].f.upper[4] );
tran (\sa_count[21][37] , \sa_count[21].r.part1[5] );
tran (\sa_count[21][37] , \sa_count[21].f.upper[5] );
tran (\sa_count[21][38] , \sa_count[21].r.part1[6] );
tran (\sa_count[21][38] , \sa_count[21].f.upper[6] );
tran (\sa_count[21][39] , \sa_count[21].r.part1[7] );
tran (\sa_count[21][39] , \sa_count[21].f.upper[7] );
tran (\sa_count[21][40] , \sa_count[21].r.part1[8] );
tran (\sa_count[21][40] , \sa_count[21].f.upper[8] );
tran (\sa_count[21][41] , \sa_count[21].r.part1[9] );
tran (\sa_count[21][41] , \sa_count[21].f.upper[9] );
tran (\sa_count[21][42] , \sa_count[21].r.part1[10] );
tran (\sa_count[21][42] , \sa_count[21].f.upper[10] );
tran (\sa_count[21][43] , \sa_count[21].r.part1[11] );
tran (\sa_count[21][43] , \sa_count[21].f.upper[11] );
tran (\sa_count[21][44] , \sa_count[21].r.part1[12] );
tran (\sa_count[21][44] , \sa_count[21].f.upper[12] );
tran (\sa_count[21][45] , \sa_count[21].r.part1[13] );
tran (\sa_count[21][45] , \sa_count[21].f.upper[13] );
tran (\sa_count[21][46] , \sa_count[21].r.part1[14] );
tran (\sa_count[21][46] , \sa_count[21].f.upper[14] );
tran (\sa_count[21][47] , \sa_count[21].r.part1[15] );
tran (\sa_count[21][47] , \sa_count[21].f.upper[15] );
tran (\sa_count[21][48] , \sa_count[21].r.part1[16] );
tran (\sa_count[21][48] , \sa_count[21].f.upper[16] );
tran (\sa_count[21][49] , \sa_count[21].r.part1[17] );
tran (\sa_count[21][49] , \sa_count[21].f.upper[17] );
tran (\sa_count[21][50] , \sa_count[21].r.part1[18] );
tran (\sa_count[21][50] , \sa_count[21].f.unused[0] );
tran (\sa_count[21][51] , \sa_count[21].r.part1[19] );
tran (\sa_count[21][51] , \sa_count[21].f.unused[1] );
tran (\sa_count[21][52] , \sa_count[21].r.part1[20] );
tran (\sa_count[21][52] , \sa_count[21].f.unused[2] );
tran (\sa_count[21][53] , \sa_count[21].r.part1[21] );
tran (\sa_count[21][53] , \sa_count[21].f.unused[3] );
tran (\sa_count[21][54] , \sa_count[21].r.part1[22] );
tran (\sa_count[21][54] , \sa_count[21].f.unused[4] );
tran (\sa_count[21][55] , \sa_count[21].r.part1[23] );
tran (\sa_count[21][55] , \sa_count[21].f.unused[5] );
tran (\sa_count[21][56] , \sa_count[21].r.part1[24] );
tran (\sa_count[21][56] , \sa_count[21].f.unused[6] );
tran (\sa_count[21][57] , \sa_count[21].r.part1[25] );
tran (\sa_count[21][57] , \sa_count[21].f.unused[7] );
tran (\sa_count[21][58] , \sa_count[21].r.part1[26] );
tran (\sa_count[21][58] , \sa_count[21].f.unused[8] );
tran (\sa_count[21][59] , \sa_count[21].r.part1[27] );
tran (\sa_count[21][59] , \sa_count[21].f.unused[9] );
tran (\sa_count[21][60] , \sa_count[21].r.part1[28] );
tran (\sa_count[21][60] , \sa_count[21].f.unused[10] );
tran (\sa_count[21][61] , \sa_count[21].r.part1[29] );
tran (\sa_count[21][61] , \sa_count[21].f.unused[11] );
tran (\sa_count[21][62] , \sa_count[21].r.part1[30] );
tran (\sa_count[21][62] , \sa_count[21].f.unused[12] );
tran (\sa_count[21][63] , \sa_count[21].r.part1[31] );
tran (\sa_count[21][63] , \sa_count[21].f.unused[13] );
tran (\sa_count[22][0] , \sa_count[22].r.part0[0] );
tran (\sa_count[22][0] , \sa_count[22].f.lower[0] );
tran (\sa_count[22][1] , \sa_count[22].r.part0[1] );
tran (\sa_count[22][1] , \sa_count[22].f.lower[1] );
tran (\sa_count[22][2] , \sa_count[22].r.part0[2] );
tran (\sa_count[22][2] , \sa_count[22].f.lower[2] );
tran (\sa_count[22][3] , \sa_count[22].r.part0[3] );
tran (\sa_count[22][3] , \sa_count[22].f.lower[3] );
tran (\sa_count[22][4] , \sa_count[22].r.part0[4] );
tran (\sa_count[22][4] , \sa_count[22].f.lower[4] );
tran (\sa_count[22][5] , \sa_count[22].r.part0[5] );
tran (\sa_count[22][5] , \sa_count[22].f.lower[5] );
tran (\sa_count[22][6] , \sa_count[22].r.part0[6] );
tran (\sa_count[22][6] , \sa_count[22].f.lower[6] );
tran (\sa_count[22][7] , \sa_count[22].r.part0[7] );
tran (\sa_count[22][7] , \sa_count[22].f.lower[7] );
tran (\sa_count[22][8] , \sa_count[22].r.part0[8] );
tran (\sa_count[22][8] , \sa_count[22].f.lower[8] );
tran (\sa_count[22][9] , \sa_count[22].r.part0[9] );
tran (\sa_count[22][9] , \sa_count[22].f.lower[9] );
tran (\sa_count[22][10] , \sa_count[22].r.part0[10] );
tran (\sa_count[22][10] , \sa_count[22].f.lower[10] );
tran (\sa_count[22][11] , \sa_count[22].r.part0[11] );
tran (\sa_count[22][11] , \sa_count[22].f.lower[11] );
tran (\sa_count[22][12] , \sa_count[22].r.part0[12] );
tran (\sa_count[22][12] , \sa_count[22].f.lower[12] );
tran (\sa_count[22][13] , \sa_count[22].r.part0[13] );
tran (\sa_count[22][13] , \sa_count[22].f.lower[13] );
tran (\sa_count[22][14] , \sa_count[22].r.part0[14] );
tran (\sa_count[22][14] , \sa_count[22].f.lower[14] );
tran (\sa_count[22][15] , \sa_count[22].r.part0[15] );
tran (\sa_count[22][15] , \sa_count[22].f.lower[15] );
tran (\sa_count[22][16] , \sa_count[22].r.part0[16] );
tran (\sa_count[22][16] , \sa_count[22].f.lower[16] );
tran (\sa_count[22][17] , \sa_count[22].r.part0[17] );
tran (\sa_count[22][17] , \sa_count[22].f.lower[17] );
tran (\sa_count[22][18] , \sa_count[22].r.part0[18] );
tran (\sa_count[22][18] , \sa_count[22].f.lower[18] );
tran (\sa_count[22][19] , \sa_count[22].r.part0[19] );
tran (\sa_count[22][19] , \sa_count[22].f.lower[19] );
tran (\sa_count[22][20] , \sa_count[22].r.part0[20] );
tran (\sa_count[22][20] , \sa_count[22].f.lower[20] );
tran (\sa_count[22][21] , \sa_count[22].r.part0[21] );
tran (\sa_count[22][21] , \sa_count[22].f.lower[21] );
tran (\sa_count[22][22] , \sa_count[22].r.part0[22] );
tran (\sa_count[22][22] , \sa_count[22].f.lower[22] );
tran (\sa_count[22][23] , \sa_count[22].r.part0[23] );
tran (\sa_count[22][23] , \sa_count[22].f.lower[23] );
tran (\sa_count[22][24] , \sa_count[22].r.part0[24] );
tran (\sa_count[22][24] , \sa_count[22].f.lower[24] );
tran (\sa_count[22][25] , \sa_count[22].r.part0[25] );
tran (\sa_count[22][25] , \sa_count[22].f.lower[25] );
tran (\sa_count[22][26] , \sa_count[22].r.part0[26] );
tran (\sa_count[22][26] , \sa_count[22].f.lower[26] );
tran (\sa_count[22][27] , \sa_count[22].r.part0[27] );
tran (\sa_count[22][27] , \sa_count[22].f.lower[27] );
tran (\sa_count[22][28] , \sa_count[22].r.part0[28] );
tran (\sa_count[22][28] , \sa_count[22].f.lower[28] );
tran (\sa_count[22][29] , \sa_count[22].r.part0[29] );
tran (\sa_count[22][29] , \sa_count[22].f.lower[29] );
tran (\sa_count[22][30] , \sa_count[22].r.part0[30] );
tran (\sa_count[22][30] , \sa_count[22].f.lower[30] );
tran (\sa_count[22][31] , \sa_count[22].r.part0[31] );
tran (\sa_count[22][31] , \sa_count[22].f.lower[31] );
tran (\sa_count[22][32] , \sa_count[22].r.part1[0] );
tran (\sa_count[22][32] , \sa_count[22].f.upper[0] );
tran (\sa_count[22][33] , \sa_count[22].r.part1[1] );
tran (\sa_count[22][33] , \sa_count[22].f.upper[1] );
tran (\sa_count[22][34] , \sa_count[22].r.part1[2] );
tran (\sa_count[22][34] , \sa_count[22].f.upper[2] );
tran (\sa_count[22][35] , \sa_count[22].r.part1[3] );
tran (\sa_count[22][35] , \sa_count[22].f.upper[3] );
tran (\sa_count[22][36] , \sa_count[22].r.part1[4] );
tran (\sa_count[22][36] , \sa_count[22].f.upper[4] );
tran (\sa_count[22][37] , \sa_count[22].r.part1[5] );
tran (\sa_count[22][37] , \sa_count[22].f.upper[5] );
tran (\sa_count[22][38] , \sa_count[22].r.part1[6] );
tran (\sa_count[22][38] , \sa_count[22].f.upper[6] );
tran (\sa_count[22][39] , \sa_count[22].r.part1[7] );
tran (\sa_count[22][39] , \sa_count[22].f.upper[7] );
tran (\sa_count[22][40] , \sa_count[22].r.part1[8] );
tran (\sa_count[22][40] , \sa_count[22].f.upper[8] );
tran (\sa_count[22][41] , \sa_count[22].r.part1[9] );
tran (\sa_count[22][41] , \sa_count[22].f.upper[9] );
tran (\sa_count[22][42] , \sa_count[22].r.part1[10] );
tran (\sa_count[22][42] , \sa_count[22].f.upper[10] );
tran (\sa_count[22][43] , \sa_count[22].r.part1[11] );
tran (\sa_count[22][43] , \sa_count[22].f.upper[11] );
tran (\sa_count[22][44] , \sa_count[22].r.part1[12] );
tran (\sa_count[22][44] , \sa_count[22].f.upper[12] );
tran (\sa_count[22][45] , \sa_count[22].r.part1[13] );
tran (\sa_count[22][45] , \sa_count[22].f.upper[13] );
tran (\sa_count[22][46] , \sa_count[22].r.part1[14] );
tran (\sa_count[22][46] , \sa_count[22].f.upper[14] );
tran (\sa_count[22][47] , \sa_count[22].r.part1[15] );
tran (\sa_count[22][47] , \sa_count[22].f.upper[15] );
tran (\sa_count[22][48] , \sa_count[22].r.part1[16] );
tran (\sa_count[22][48] , \sa_count[22].f.upper[16] );
tran (\sa_count[22][49] , \sa_count[22].r.part1[17] );
tran (\sa_count[22][49] , \sa_count[22].f.upper[17] );
tran (\sa_count[22][50] , \sa_count[22].r.part1[18] );
tran (\sa_count[22][50] , \sa_count[22].f.unused[0] );
tran (\sa_count[22][51] , \sa_count[22].r.part1[19] );
tran (\sa_count[22][51] , \sa_count[22].f.unused[1] );
tran (\sa_count[22][52] , \sa_count[22].r.part1[20] );
tran (\sa_count[22][52] , \sa_count[22].f.unused[2] );
tran (\sa_count[22][53] , \sa_count[22].r.part1[21] );
tran (\sa_count[22][53] , \sa_count[22].f.unused[3] );
tran (\sa_count[22][54] , \sa_count[22].r.part1[22] );
tran (\sa_count[22][54] , \sa_count[22].f.unused[4] );
tran (\sa_count[22][55] , \sa_count[22].r.part1[23] );
tran (\sa_count[22][55] , \sa_count[22].f.unused[5] );
tran (\sa_count[22][56] , \sa_count[22].r.part1[24] );
tran (\sa_count[22][56] , \sa_count[22].f.unused[6] );
tran (\sa_count[22][57] , \sa_count[22].r.part1[25] );
tran (\sa_count[22][57] , \sa_count[22].f.unused[7] );
tran (\sa_count[22][58] , \sa_count[22].r.part1[26] );
tran (\sa_count[22][58] , \sa_count[22].f.unused[8] );
tran (\sa_count[22][59] , \sa_count[22].r.part1[27] );
tran (\sa_count[22][59] , \sa_count[22].f.unused[9] );
tran (\sa_count[22][60] , \sa_count[22].r.part1[28] );
tran (\sa_count[22][60] , \sa_count[22].f.unused[10] );
tran (\sa_count[22][61] , \sa_count[22].r.part1[29] );
tran (\sa_count[22][61] , \sa_count[22].f.unused[11] );
tran (\sa_count[22][62] , \sa_count[22].r.part1[30] );
tran (\sa_count[22][62] , \sa_count[22].f.unused[12] );
tran (\sa_count[22][63] , \sa_count[22].r.part1[31] );
tran (\sa_count[22][63] , \sa_count[22].f.unused[13] );
tran (\sa_count[23][0] , \sa_count[23].r.part0[0] );
tran (\sa_count[23][0] , \sa_count[23].f.lower[0] );
tran (\sa_count[23][1] , \sa_count[23].r.part0[1] );
tran (\sa_count[23][1] , \sa_count[23].f.lower[1] );
tran (\sa_count[23][2] , \sa_count[23].r.part0[2] );
tran (\sa_count[23][2] , \sa_count[23].f.lower[2] );
tran (\sa_count[23][3] , \sa_count[23].r.part0[3] );
tran (\sa_count[23][3] , \sa_count[23].f.lower[3] );
tran (\sa_count[23][4] , \sa_count[23].r.part0[4] );
tran (\sa_count[23][4] , \sa_count[23].f.lower[4] );
tran (\sa_count[23][5] , \sa_count[23].r.part0[5] );
tran (\sa_count[23][5] , \sa_count[23].f.lower[5] );
tran (\sa_count[23][6] , \sa_count[23].r.part0[6] );
tran (\sa_count[23][6] , \sa_count[23].f.lower[6] );
tran (\sa_count[23][7] , \sa_count[23].r.part0[7] );
tran (\sa_count[23][7] , \sa_count[23].f.lower[7] );
tran (\sa_count[23][8] , \sa_count[23].r.part0[8] );
tran (\sa_count[23][8] , \sa_count[23].f.lower[8] );
tran (\sa_count[23][9] , \sa_count[23].r.part0[9] );
tran (\sa_count[23][9] , \sa_count[23].f.lower[9] );
tran (\sa_count[23][10] , \sa_count[23].r.part0[10] );
tran (\sa_count[23][10] , \sa_count[23].f.lower[10] );
tran (\sa_count[23][11] , \sa_count[23].r.part0[11] );
tran (\sa_count[23][11] , \sa_count[23].f.lower[11] );
tran (\sa_count[23][12] , \sa_count[23].r.part0[12] );
tran (\sa_count[23][12] , \sa_count[23].f.lower[12] );
tran (\sa_count[23][13] , \sa_count[23].r.part0[13] );
tran (\sa_count[23][13] , \sa_count[23].f.lower[13] );
tran (\sa_count[23][14] , \sa_count[23].r.part0[14] );
tran (\sa_count[23][14] , \sa_count[23].f.lower[14] );
tran (\sa_count[23][15] , \sa_count[23].r.part0[15] );
tran (\sa_count[23][15] , \sa_count[23].f.lower[15] );
tran (\sa_count[23][16] , \sa_count[23].r.part0[16] );
tran (\sa_count[23][16] , \sa_count[23].f.lower[16] );
tran (\sa_count[23][17] , \sa_count[23].r.part0[17] );
tran (\sa_count[23][17] , \sa_count[23].f.lower[17] );
tran (\sa_count[23][18] , \sa_count[23].r.part0[18] );
tran (\sa_count[23][18] , \sa_count[23].f.lower[18] );
tran (\sa_count[23][19] , \sa_count[23].r.part0[19] );
tran (\sa_count[23][19] , \sa_count[23].f.lower[19] );
tran (\sa_count[23][20] , \sa_count[23].r.part0[20] );
tran (\sa_count[23][20] , \sa_count[23].f.lower[20] );
tran (\sa_count[23][21] , \sa_count[23].r.part0[21] );
tran (\sa_count[23][21] , \sa_count[23].f.lower[21] );
tran (\sa_count[23][22] , \sa_count[23].r.part0[22] );
tran (\sa_count[23][22] , \sa_count[23].f.lower[22] );
tran (\sa_count[23][23] , \sa_count[23].r.part0[23] );
tran (\sa_count[23][23] , \sa_count[23].f.lower[23] );
tran (\sa_count[23][24] , \sa_count[23].r.part0[24] );
tran (\sa_count[23][24] , \sa_count[23].f.lower[24] );
tran (\sa_count[23][25] , \sa_count[23].r.part0[25] );
tran (\sa_count[23][25] , \sa_count[23].f.lower[25] );
tran (\sa_count[23][26] , \sa_count[23].r.part0[26] );
tran (\sa_count[23][26] , \sa_count[23].f.lower[26] );
tran (\sa_count[23][27] , \sa_count[23].r.part0[27] );
tran (\sa_count[23][27] , \sa_count[23].f.lower[27] );
tran (\sa_count[23][28] , \sa_count[23].r.part0[28] );
tran (\sa_count[23][28] , \sa_count[23].f.lower[28] );
tran (\sa_count[23][29] , \sa_count[23].r.part0[29] );
tran (\sa_count[23][29] , \sa_count[23].f.lower[29] );
tran (\sa_count[23][30] , \sa_count[23].r.part0[30] );
tran (\sa_count[23][30] , \sa_count[23].f.lower[30] );
tran (\sa_count[23][31] , \sa_count[23].r.part0[31] );
tran (\sa_count[23][31] , \sa_count[23].f.lower[31] );
tran (\sa_count[23][32] , \sa_count[23].r.part1[0] );
tran (\sa_count[23][32] , \sa_count[23].f.upper[0] );
tran (\sa_count[23][33] , \sa_count[23].r.part1[1] );
tran (\sa_count[23][33] , \sa_count[23].f.upper[1] );
tran (\sa_count[23][34] , \sa_count[23].r.part1[2] );
tran (\sa_count[23][34] , \sa_count[23].f.upper[2] );
tran (\sa_count[23][35] , \sa_count[23].r.part1[3] );
tran (\sa_count[23][35] , \sa_count[23].f.upper[3] );
tran (\sa_count[23][36] , \sa_count[23].r.part1[4] );
tran (\sa_count[23][36] , \sa_count[23].f.upper[4] );
tran (\sa_count[23][37] , \sa_count[23].r.part1[5] );
tran (\sa_count[23][37] , \sa_count[23].f.upper[5] );
tran (\sa_count[23][38] , \sa_count[23].r.part1[6] );
tran (\sa_count[23][38] , \sa_count[23].f.upper[6] );
tran (\sa_count[23][39] , \sa_count[23].r.part1[7] );
tran (\sa_count[23][39] , \sa_count[23].f.upper[7] );
tran (\sa_count[23][40] , \sa_count[23].r.part1[8] );
tran (\sa_count[23][40] , \sa_count[23].f.upper[8] );
tran (\sa_count[23][41] , \sa_count[23].r.part1[9] );
tran (\sa_count[23][41] , \sa_count[23].f.upper[9] );
tran (\sa_count[23][42] , \sa_count[23].r.part1[10] );
tran (\sa_count[23][42] , \sa_count[23].f.upper[10] );
tran (\sa_count[23][43] , \sa_count[23].r.part1[11] );
tran (\sa_count[23][43] , \sa_count[23].f.upper[11] );
tran (\sa_count[23][44] , \sa_count[23].r.part1[12] );
tran (\sa_count[23][44] , \sa_count[23].f.upper[12] );
tran (\sa_count[23][45] , \sa_count[23].r.part1[13] );
tran (\sa_count[23][45] , \sa_count[23].f.upper[13] );
tran (\sa_count[23][46] , \sa_count[23].r.part1[14] );
tran (\sa_count[23][46] , \sa_count[23].f.upper[14] );
tran (\sa_count[23][47] , \sa_count[23].r.part1[15] );
tran (\sa_count[23][47] , \sa_count[23].f.upper[15] );
tran (\sa_count[23][48] , \sa_count[23].r.part1[16] );
tran (\sa_count[23][48] , \sa_count[23].f.upper[16] );
tran (\sa_count[23][49] , \sa_count[23].r.part1[17] );
tran (\sa_count[23][49] , \sa_count[23].f.upper[17] );
tran (\sa_count[23][50] , \sa_count[23].r.part1[18] );
tran (\sa_count[23][50] , \sa_count[23].f.unused[0] );
tran (\sa_count[23][51] , \sa_count[23].r.part1[19] );
tran (\sa_count[23][51] , \sa_count[23].f.unused[1] );
tran (\sa_count[23][52] , \sa_count[23].r.part1[20] );
tran (\sa_count[23][52] , \sa_count[23].f.unused[2] );
tran (\sa_count[23][53] , \sa_count[23].r.part1[21] );
tran (\sa_count[23][53] , \sa_count[23].f.unused[3] );
tran (\sa_count[23][54] , \sa_count[23].r.part1[22] );
tran (\sa_count[23][54] , \sa_count[23].f.unused[4] );
tran (\sa_count[23][55] , \sa_count[23].r.part1[23] );
tran (\sa_count[23][55] , \sa_count[23].f.unused[5] );
tran (\sa_count[23][56] , \sa_count[23].r.part1[24] );
tran (\sa_count[23][56] , \sa_count[23].f.unused[6] );
tran (\sa_count[23][57] , \sa_count[23].r.part1[25] );
tran (\sa_count[23][57] , \sa_count[23].f.unused[7] );
tran (\sa_count[23][58] , \sa_count[23].r.part1[26] );
tran (\sa_count[23][58] , \sa_count[23].f.unused[8] );
tran (\sa_count[23][59] , \sa_count[23].r.part1[27] );
tran (\sa_count[23][59] , \sa_count[23].f.unused[9] );
tran (\sa_count[23][60] , \sa_count[23].r.part1[28] );
tran (\sa_count[23][60] , \sa_count[23].f.unused[10] );
tran (\sa_count[23][61] , \sa_count[23].r.part1[29] );
tran (\sa_count[23][61] , \sa_count[23].f.unused[11] );
tran (\sa_count[23][62] , \sa_count[23].r.part1[30] );
tran (\sa_count[23][62] , \sa_count[23].f.unused[12] );
tran (\sa_count[23][63] , \sa_count[23].r.part1[31] );
tran (\sa_count[23][63] , \sa_count[23].f.unused[13] );
tran (\sa_count[24][0] , \sa_count[24].r.part0[0] );
tran (\sa_count[24][0] , \sa_count[24].f.lower[0] );
tran (\sa_count[24][1] , \sa_count[24].r.part0[1] );
tran (\sa_count[24][1] , \sa_count[24].f.lower[1] );
tran (\sa_count[24][2] , \sa_count[24].r.part0[2] );
tran (\sa_count[24][2] , \sa_count[24].f.lower[2] );
tran (\sa_count[24][3] , \sa_count[24].r.part0[3] );
tran (\sa_count[24][3] , \sa_count[24].f.lower[3] );
tran (\sa_count[24][4] , \sa_count[24].r.part0[4] );
tran (\sa_count[24][4] , \sa_count[24].f.lower[4] );
tran (\sa_count[24][5] , \sa_count[24].r.part0[5] );
tran (\sa_count[24][5] , \sa_count[24].f.lower[5] );
tran (\sa_count[24][6] , \sa_count[24].r.part0[6] );
tran (\sa_count[24][6] , \sa_count[24].f.lower[6] );
tran (\sa_count[24][7] , \sa_count[24].r.part0[7] );
tran (\sa_count[24][7] , \sa_count[24].f.lower[7] );
tran (\sa_count[24][8] , \sa_count[24].r.part0[8] );
tran (\sa_count[24][8] , \sa_count[24].f.lower[8] );
tran (\sa_count[24][9] , \sa_count[24].r.part0[9] );
tran (\sa_count[24][9] , \sa_count[24].f.lower[9] );
tran (\sa_count[24][10] , \sa_count[24].r.part0[10] );
tran (\sa_count[24][10] , \sa_count[24].f.lower[10] );
tran (\sa_count[24][11] , \sa_count[24].r.part0[11] );
tran (\sa_count[24][11] , \sa_count[24].f.lower[11] );
tran (\sa_count[24][12] , \sa_count[24].r.part0[12] );
tran (\sa_count[24][12] , \sa_count[24].f.lower[12] );
tran (\sa_count[24][13] , \sa_count[24].r.part0[13] );
tran (\sa_count[24][13] , \sa_count[24].f.lower[13] );
tran (\sa_count[24][14] , \sa_count[24].r.part0[14] );
tran (\sa_count[24][14] , \sa_count[24].f.lower[14] );
tran (\sa_count[24][15] , \sa_count[24].r.part0[15] );
tran (\sa_count[24][15] , \sa_count[24].f.lower[15] );
tran (\sa_count[24][16] , \sa_count[24].r.part0[16] );
tran (\sa_count[24][16] , \sa_count[24].f.lower[16] );
tran (\sa_count[24][17] , \sa_count[24].r.part0[17] );
tran (\sa_count[24][17] , \sa_count[24].f.lower[17] );
tran (\sa_count[24][18] , \sa_count[24].r.part0[18] );
tran (\sa_count[24][18] , \sa_count[24].f.lower[18] );
tran (\sa_count[24][19] , \sa_count[24].r.part0[19] );
tran (\sa_count[24][19] , \sa_count[24].f.lower[19] );
tran (\sa_count[24][20] , \sa_count[24].r.part0[20] );
tran (\sa_count[24][20] , \sa_count[24].f.lower[20] );
tran (\sa_count[24][21] , \sa_count[24].r.part0[21] );
tran (\sa_count[24][21] , \sa_count[24].f.lower[21] );
tran (\sa_count[24][22] , \sa_count[24].r.part0[22] );
tran (\sa_count[24][22] , \sa_count[24].f.lower[22] );
tran (\sa_count[24][23] , \sa_count[24].r.part0[23] );
tran (\sa_count[24][23] , \sa_count[24].f.lower[23] );
tran (\sa_count[24][24] , \sa_count[24].r.part0[24] );
tran (\sa_count[24][24] , \sa_count[24].f.lower[24] );
tran (\sa_count[24][25] , \sa_count[24].r.part0[25] );
tran (\sa_count[24][25] , \sa_count[24].f.lower[25] );
tran (\sa_count[24][26] , \sa_count[24].r.part0[26] );
tran (\sa_count[24][26] , \sa_count[24].f.lower[26] );
tran (\sa_count[24][27] , \sa_count[24].r.part0[27] );
tran (\sa_count[24][27] , \sa_count[24].f.lower[27] );
tran (\sa_count[24][28] , \sa_count[24].r.part0[28] );
tran (\sa_count[24][28] , \sa_count[24].f.lower[28] );
tran (\sa_count[24][29] , \sa_count[24].r.part0[29] );
tran (\sa_count[24][29] , \sa_count[24].f.lower[29] );
tran (\sa_count[24][30] , \sa_count[24].r.part0[30] );
tran (\sa_count[24][30] , \sa_count[24].f.lower[30] );
tran (\sa_count[24][31] , \sa_count[24].r.part0[31] );
tran (\sa_count[24][31] , \sa_count[24].f.lower[31] );
tran (\sa_count[24][32] , \sa_count[24].r.part1[0] );
tran (\sa_count[24][32] , \sa_count[24].f.upper[0] );
tran (\sa_count[24][33] , \sa_count[24].r.part1[1] );
tran (\sa_count[24][33] , \sa_count[24].f.upper[1] );
tran (\sa_count[24][34] , \sa_count[24].r.part1[2] );
tran (\sa_count[24][34] , \sa_count[24].f.upper[2] );
tran (\sa_count[24][35] , \sa_count[24].r.part1[3] );
tran (\sa_count[24][35] , \sa_count[24].f.upper[3] );
tran (\sa_count[24][36] , \sa_count[24].r.part1[4] );
tran (\sa_count[24][36] , \sa_count[24].f.upper[4] );
tran (\sa_count[24][37] , \sa_count[24].r.part1[5] );
tran (\sa_count[24][37] , \sa_count[24].f.upper[5] );
tran (\sa_count[24][38] , \sa_count[24].r.part1[6] );
tran (\sa_count[24][38] , \sa_count[24].f.upper[6] );
tran (\sa_count[24][39] , \sa_count[24].r.part1[7] );
tran (\sa_count[24][39] , \sa_count[24].f.upper[7] );
tran (\sa_count[24][40] , \sa_count[24].r.part1[8] );
tran (\sa_count[24][40] , \sa_count[24].f.upper[8] );
tran (\sa_count[24][41] , \sa_count[24].r.part1[9] );
tran (\sa_count[24][41] , \sa_count[24].f.upper[9] );
tran (\sa_count[24][42] , \sa_count[24].r.part1[10] );
tran (\sa_count[24][42] , \sa_count[24].f.upper[10] );
tran (\sa_count[24][43] , \sa_count[24].r.part1[11] );
tran (\sa_count[24][43] , \sa_count[24].f.upper[11] );
tran (\sa_count[24][44] , \sa_count[24].r.part1[12] );
tran (\sa_count[24][44] , \sa_count[24].f.upper[12] );
tran (\sa_count[24][45] , \sa_count[24].r.part1[13] );
tran (\sa_count[24][45] , \sa_count[24].f.upper[13] );
tran (\sa_count[24][46] , \sa_count[24].r.part1[14] );
tran (\sa_count[24][46] , \sa_count[24].f.upper[14] );
tran (\sa_count[24][47] , \sa_count[24].r.part1[15] );
tran (\sa_count[24][47] , \sa_count[24].f.upper[15] );
tran (\sa_count[24][48] , \sa_count[24].r.part1[16] );
tran (\sa_count[24][48] , \sa_count[24].f.upper[16] );
tran (\sa_count[24][49] , \sa_count[24].r.part1[17] );
tran (\sa_count[24][49] , \sa_count[24].f.upper[17] );
tran (\sa_count[24][50] , \sa_count[24].r.part1[18] );
tran (\sa_count[24][50] , \sa_count[24].f.unused[0] );
tran (\sa_count[24][51] , \sa_count[24].r.part1[19] );
tran (\sa_count[24][51] , \sa_count[24].f.unused[1] );
tran (\sa_count[24][52] , \sa_count[24].r.part1[20] );
tran (\sa_count[24][52] , \sa_count[24].f.unused[2] );
tran (\sa_count[24][53] , \sa_count[24].r.part1[21] );
tran (\sa_count[24][53] , \sa_count[24].f.unused[3] );
tran (\sa_count[24][54] , \sa_count[24].r.part1[22] );
tran (\sa_count[24][54] , \sa_count[24].f.unused[4] );
tran (\sa_count[24][55] , \sa_count[24].r.part1[23] );
tran (\sa_count[24][55] , \sa_count[24].f.unused[5] );
tran (\sa_count[24][56] , \sa_count[24].r.part1[24] );
tran (\sa_count[24][56] , \sa_count[24].f.unused[6] );
tran (\sa_count[24][57] , \sa_count[24].r.part1[25] );
tran (\sa_count[24][57] , \sa_count[24].f.unused[7] );
tran (\sa_count[24][58] , \sa_count[24].r.part1[26] );
tran (\sa_count[24][58] , \sa_count[24].f.unused[8] );
tran (\sa_count[24][59] , \sa_count[24].r.part1[27] );
tran (\sa_count[24][59] , \sa_count[24].f.unused[9] );
tran (\sa_count[24][60] , \sa_count[24].r.part1[28] );
tran (\sa_count[24][60] , \sa_count[24].f.unused[10] );
tran (\sa_count[24][61] , \sa_count[24].r.part1[29] );
tran (\sa_count[24][61] , \sa_count[24].f.unused[11] );
tran (\sa_count[24][62] , \sa_count[24].r.part1[30] );
tran (\sa_count[24][62] , \sa_count[24].f.unused[12] );
tran (\sa_count[24][63] , \sa_count[24].r.part1[31] );
tran (\sa_count[24][63] , \sa_count[24].f.unused[13] );
tran (\sa_count[25][0] , \sa_count[25].r.part0[0] );
tran (\sa_count[25][0] , \sa_count[25].f.lower[0] );
tran (\sa_count[25][1] , \sa_count[25].r.part0[1] );
tran (\sa_count[25][1] , \sa_count[25].f.lower[1] );
tran (\sa_count[25][2] , \sa_count[25].r.part0[2] );
tran (\sa_count[25][2] , \sa_count[25].f.lower[2] );
tran (\sa_count[25][3] , \sa_count[25].r.part0[3] );
tran (\sa_count[25][3] , \sa_count[25].f.lower[3] );
tran (\sa_count[25][4] , \sa_count[25].r.part0[4] );
tran (\sa_count[25][4] , \sa_count[25].f.lower[4] );
tran (\sa_count[25][5] , \sa_count[25].r.part0[5] );
tran (\sa_count[25][5] , \sa_count[25].f.lower[5] );
tran (\sa_count[25][6] , \sa_count[25].r.part0[6] );
tran (\sa_count[25][6] , \sa_count[25].f.lower[6] );
tran (\sa_count[25][7] , \sa_count[25].r.part0[7] );
tran (\sa_count[25][7] , \sa_count[25].f.lower[7] );
tran (\sa_count[25][8] , \sa_count[25].r.part0[8] );
tran (\sa_count[25][8] , \sa_count[25].f.lower[8] );
tran (\sa_count[25][9] , \sa_count[25].r.part0[9] );
tran (\sa_count[25][9] , \sa_count[25].f.lower[9] );
tran (\sa_count[25][10] , \sa_count[25].r.part0[10] );
tran (\sa_count[25][10] , \sa_count[25].f.lower[10] );
tran (\sa_count[25][11] , \sa_count[25].r.part0[11] );
tran (\sa_count[25][11] , \sa_count[25].f.lower[11] );
tran (\sa_count[25][12] , \sa_count[25].r.part0[12] );
tran (\sa_count[25][12] , \sa_count[25].f.lower[12] );
tran (\sa_count[25][13] , \sa_count[25].r.part0[13] );
tran (\sa_count[25][13] , \sa_count[25].f.lower[13] );
tran (\sa_count[25][14] , \sa_count[25].r.part0[14] );
tran (\sa_count[25][14] , \sa_count[25].f.lower[14] );
tran (\sa_count[25][15] , \sa_count[25].r.part0[15] );
tran (\sa_count[25][15] , \sa_count[25].f.lower[15] );
tran (\sa_count[25][16] , \sa_count[25].r.part0[16] );
tran (\sa_count[25][16] , \sa_count[25].f.lower[16] );
tran (\sa_count[25][17] , \sa_count[25].r.part0[17] );
tran (\sa_count[25][17] , \sa_count[25].f.lower[17] );
tran (\sa_count[25][18] , \sa_count[25].r.part0[18] );
tran (\sa_count[25][18] , \sa_count[25].f.lower[18] );
tran (\sa_count[25][19] , \sa_count[25].r.part0[19] );
tran (\sa_count[25][19] , \sa_count[25].f.lower[19] );
tran (\sa_count[25][20] , \sa_count[25].r.part0[20] );
tran (\sa_count[25][20] , \sa_count[25].f.lower[20] );
tran (\sa_count[25][21] , \sa_count[25].r.part0[21] );
tran (\sa_count[25][21] , \sa_count[25].f.lower[21] );
tran (\sa_count[25][22] , \sa_count[25].r.part0[22] );
tran (\sa_count[25][22] , \sa_count[25].f.lower[22] );
tran (\sa_count[25][23] , \sa_count[25].r.part0[23] );
tran (\sa_count[25][23] , \sa_count[25].f.lower[23] );
tran (\sa_count[25][24] , \sa_count[25].r.part0[24] );
tran (\sa_count[25][24] , \sa_count[25].f.lower[24] );
tran (\sa_count[25][25] , \sa_count[25].r.part0[25] );
tran (\sa_count[25][25] , \sa_count[25].f.lower[25] );
tran (\sa_count[25][26] , \sa_count[25].r.part0[26] );
tran (\sa_count[25][26] , \sa_count[25].f.lower[26] );
tran (\sa_count[25][27] , \sa_count[25].r.part0[27] );
tran (\sa_count[25][27] , \sa_count[25].f.lower[27] );
tran (\sa_count[25][28] , \sa_count[25].r.part0[28] );
tran (\sa_count[25][28] , \sa_count[25].f.lower[28] );
tran (\sa_count[25][29] , \sa_count[25].r.part0[29] );
tran (\sa_count[25][29] , \sa_count[25].f.lower[29] );
tran (\sa_count[25][30] , \sa_count[25].r.part0[30] );
tran (\sa_count[25][30] , \sa_count[25].f.lower[30] );
tran (\sa_count[25][31] , \sa_count[25].r.part0[31] );
tran (\sa_count[25][31] , \sa_count[25].f.lower[31] );
tran (\sa_count[25][32] , \sa_count[25].r.part1[0] );
tran (\sa_count[25][32] , \sa_count[25].f.upper[0] );
tran (\sa_count[25][33] , \sa_count[25].r.part1[1] );
tran (\sa_count[25][33] , \sa_count[25].f.upper[1] );
tran (\sa_count[25][34] , \sa_count[25].r.part1[2] );
tran (\sa_count[25][34] , \sa_count[25].f.upper[2] );
tran (\sa_count[25][35] , \sa_count[25].r.part1[3] );
tran (\sa_count[25][35] , \sa_count[25].f.upper[3] );
tran (\sa_count[25][36] , \sa_count[25].r.part1[4] );
tran (\sa_count[25][36] , \sa_count[25].f.upper[4] );
tran (\sa_count[25][37] , \sa_count[25].r.part1[5] );
tran (\sa_count[25][37] , \sa_count[25].f.upper[5] );
tran (\sa_count[25][38] , \sa_count[25].r.part1[6] );
tran (\sa_count[25][38] , \sa_count[25].f.upper[6] );
tran (\sa_count[25][39] , \sa_count[25].r.part1[7] );
tran (\sa_count[25][39] , \sa_count[25].f.upper[7] );
tran (\sa_count[25][40] , \sa_count[25].r.part1[8] );
tran (\sa_count[25][40] , \sa_count[25].f.upper[8] );
tran (\sa_count[25][41] , \sa_count[25].r.part1[9] );
tran (\sa_count[25][41] , \sa_count[25].f.upper[9] );
tran (\sa_count[25][42] , \sa_count[25].r.part1[10] );
tran (\sa_count[25][42] , \sa_count[25].f.upper[10] );
tran (\sa_count[25][43] , \sa_count[25].r.part1[11] );
tran (\sa_count[25][43] , \sa_count[25].f.upper[11] );
tran (\sa_count[25][44] , \sa_count[25].r.part1[12] );
tran (\sa_count[25][44] , \sa_count[25].f.upper[12] );
tran (\sa_count[25][45] , \sa_count[25].r.part1[13] );
tran (\sa_count[25][45] , \sa_count[25].f.upper[13] );
tran (\sa_count[25][46] , \sa_count[25].r.part1[14] );
tran (\sa_count[25][46] , \sa_count[25].f.upper[14] );
tran (\sa_count[25][47] , \sa_count[25].r.part1[15] );
tran (\sa_count[25][47] , \sa_count[25].f.upper[15] );
tran (\sa_count[25][48] , \sa_count[25].r.part1[16] );
tran (\sa_count[25][48] , \sa_count[25].f.upper[16] );
tran (\sa_count[25][49] , \sa_count[25].r.part1[17] );
tran (\sa_count[25][49] , \sa_count[25].f.upper[17] );
tran (\sa_count[25][50] , \sa_count[25].r.part1[18] );
tran (\sa_count[25][50] , \sa_count[25].f.unused[0] );
tran (\sa_count[25][51] , \sa_count[25].r.part1[19] );
tran (\sa_count[25][51] , \sa_count[25].f.unused[1] );
tran (\sa_count[25][52] , \sa_count[25].r.part1[20] );
tran (\sa_count[25][52] , \sa_count[25].f.unused[2] );
tran (\sa_count[25][53] , \sa_count[25].r.part1[21] );
tran (\sa_count[25][53] , \sa_count[25].f.unused[3] );
tran (\sa_count[25][54] , \sa_count[25].r.part1[22] );
tran (\sa_count[25][54] , \sa_count[25].f.unused[4] );
tran (\sa_count[25][55] , \sa_count[25].r.part1[23] );
tran (\sa_count[25][55] , \sa_count[25].f.unused[5] );
tran (\sa_count[25][56] , \sa_count[25].r.part1[24] );
tran (\sa_count[25][56] , \sa_count[25].f.unused[6] );
tran (\sa_count[25][57] , \sa_count[25].r.part1[25] );
tran (\sa_count[25][57] , \sa_count[25].f.unused[7] );
tran (\sa_count[25][58] , \sa_count[25].r.part1[26] );
tran (\sa_count[25][58] , \sa_count[25].f.unused[8] );
tran (\sa_count[25][59] , \sa_count[25].r.part1[27] );
tran (\sa_count[25][59] , \sa_count[25].f.unused[9] );
tran (\sa_count[25][60] , \sa_count[25].r.part1[28] );
tran (\sa_count[25][60] , \sa_count[25].f.unused[10] );
tran (\sa_count[25][61] , \sa_count[25].r.part1[29] );
tran (\sa_count[25][61] , \sa_count[25].f.unused[11] );
tran (\sa_count[25][62] , \sa_count[25].r.part1[30] );
tran (\sa_count[25][62] , \sa_count[25].f.unused[12] );
tran (\sa_count[25][63] , \sa_count[25].r.part1[31] );
tran (\sa_count[25][63] , \sa_count[25].f.unused[13] );
tran (\sa_count[26][0] , \sa_count[26].r.part0[0] );
tran (\sa_count[26][0] , \sa_count[26].f.lower[0] );
tran (\sa_count[26][1] , \sa_count[26].r.part0[1] );
tran (\sa_count[26][1] , \sa_count[26].f.lower[1] );
tran (\sa_count[26][2] , \sa_count[26].r.part0[2] );
tran (\sa_count[26][2] , \sa_count[26].f.lower[2] );
tran (\sa_count[26][3] , \sa_count[26].r.part0[3] );
tran (\sa_count[26][3] , \sa_count[26].f.lower[3] );
tran (\sa_count[26][4] , \sa_count[26].r.part0[4] );
tran (\sa_count[26][4] , \sa_count[26].f.lower[4] );
tran (\sa_count[26][5] , \sa_count[26].r.part0[5] );
tran (\sa_count[26][5] , \sa_count[26].f.lower[5] );
tran (\sa_count[26][6] , \sa_count[26].r.part0[6] );
tran (\sa_count[26][6] , \sa_count[26].f.lower[6] );
tran (\sa_count[26][7] , \sa_count[26].r.part0[7] );
tran (\sa_count[26][7] , \sa_count[26].f.lower[7] );
tran (\sa_count[26][8] , \sa_count[26].r.part0[8] );
tran (\sa_count[26][8] , \sa_count[26].f.lower[8] );
tran (\sa_count[26][9] , \sa_count[26].r.part0[9] );
tran (\sa_count[26][9] , \sa_count[26].f.lower[9] );
tran (\sa_count[26][10] , \sa_count[26].r.part0[10] );
tran (\sa_count[26][10] , \sa_count[26].f.lower[10] );
tran (\sa_count[26][11] , \sa_count[26].r.part0[11] );
tran (\sa_count[26][11] , \sa_count[26].f.lower[11] );
tran (\sa_count[26][12] , \sa_count[26].r.part0[12] );
tran (\sa_count[26][12] , \sa_count[26].f.lower[12] );
tran (\sa_count[26][13] , \sa_count[26].r.part0[13] );
tran (\sa_count[26][13] , \sa_count[26].f.lower[13] );
tran (\sa_count[26][14] , \sa_count[26].r.part0[14] );
tran (\sa_count[26][14] , \sa_count[26].f.lower[14] );
tran (\sa_count[26][15] , \sa_count[26].r.part0[15] );
tran (\sa_count[26][15] , \sa_count[26].f.lower[15] );
tran (\sa_count[26][16] , \sa_count[26].r.part0[16] );
tran (\sa_count[26][16] , \sa_count[26].f.lower[16] );
tran (\sa_count[26][17] , \sa_count[26].r.part0[17] );
tran (\sa_count[26][17] , \sa_count[26].f.lower[17] );
tran (\sa_count[26][18] , \sa_count[26].r.part0[18] );
tran (\sa_count[26][18] , \sa_count[26].f.lower[18] );
tran (\sa_count[26][19] , \sa_count[26].r.part0[19] );
tran (\sa_count[26][19] , \sa_count[26].f.lower[19] );
tran (\sa_count[26][20] , \sa_count[26].r.part0[20] );
tran (\sa_count[26][20] , \sa_count[26].f.lower[20] );
tran (\sa_count[26][21] , \sa_count[26].r.part0[21] );
tran (\sa_count[26][21] , \sa_count[26].f.lower[21] );
tran (\sa_count[26][22] , \sa_count[26].r.part0[22] );
tran (\sa_count[26][22] , \sa_count[26].f.lower[22] );
tran (\sa_count[26][23] , \sa_count[26].r.part0[23] );
tran (\sa_count[26][23] , \sa_count[26].f.lower[23] );
tran (\sa_count[26][24] , \sa_count[26].r.part0[24] );
tran (\sa_count[26][24] , \sa_count[26].f.lower[24] );
tran (\sa_count[26][25] , \sa_count[26].r.part0[25] );
tran (\sa_count[26][25] , \sa_count[26].f.lower[25] );
tran (\sa_count[26][26] , \sa_count[26].r.part0[26] );
tran (\sa_count[26][26] , \sa_count[26].f.lower[26] );
tran (\sa_count[26][27] , \sa_count[26].r.part0[27] );
tran (\sa_count[26][27] , \sa_count[26].f.lower[27] );
tran (\sa_count[26][28] , \sa_count[26].r.part0[28] );
tran (\sa_count[26][28] , \sa_count[26].f.lower[28] );
tran (\sa_count[26][29] , \sa_count[26].r.part0[29] );
tran (\sa_count[26][29] , \sa_count[26].f.lower[29] );
tran (\sa_count[26][30] , \sa_count[26].r.part0[30] );
tran (\sa_count[26][30] , \sa_count[26].f.lower[30] );
tran (\sa_count[26][31] , \sa_count[26].r.part0[31] );
tran (\sa_count[26][31] , \sa_count[26].f.lower[31] );
tran (\sa_count[26][32] , \sa_count[26].r.part1[0] );
tran (\sa_count[26][32] , \sa_count[26].f.upper[0] );
tran (\sa_count[26][33] , \sa_count[26].r.part1[1] );
tran (\sa_count[26][33] , \sa_count[26].f.upper[1] );
tran (\sa_count[26][34] , \sa_count[26].r.part1[2] );
tran (\sa_count[26][34] , \sa_count[26].f.upper[2] );
tran (\sa_count[26][35] , \sa_count[26].r.part1[3] );
tran (\sa_count[26][35] , \sa_count[26].f.upper[3] );
tran (\sa_count[26][36] , \sa_count[26].r.part1[4] );
tran (\sa_count[26][36] , \sa_count[26].f.upper[4] );
tran (\sa_count[26][37] , \sa_count[26].r.part1[5] );
tran (\sa_count[26][37] , \sa_count[26].f.upper[5] );
tran (\sa_count[26][38] , \sa_count[26].r.part1[6] );
tran (\sa_count[26][38] , \sa_count[26].f.upper[6] );
tran (\sa_count[26][39] , \sa_count[26].r.part1[7] );
tran (\sa_count[26][39] , \sa_count[26].f.upper[7] );
tran (\sa_count[26][40] , \sa_count[26].r.part1[8] );
tran (\sa_count[26][40] , \sa_count[26].f.upper[8] );
tran (\sa_count[26][41] , \sa_count[26].r.part1[9] );
tran (\sa_count[26][41] , \sa_count[26].f.upper[9] );
tran (\sa_count[26][42] , \sa_count[26].r.part1[10] );
tran (\sa_count[26][42] , \sa_count[26].f.upper[10] );
tran (\sa_count[26][43] , \sa_count[26].r.part1[11] );
tran (\sa_count[26][43] , \sa_count[26].f.upper[11] );
tran (\sa_count[26][44] , \sa_count[26].r.part1[12] );
tran (\sa_count[26][44] , \sa_count[26].f.upper[12] );
tran (\sa_count[26][45] , \sa_count[26].r.part1[13] );
tran (\sa_count[26][45] , \sa_count[26].f.upper[13] );
tran (\sa_count[26][46] , \sa_count[26].r.part1[14] );
tran (\sa_count[26][46] , \sa_count[26].f.upper[14] );
tran (\sa_count[26][47] , \sa_count[26].r.part1[15] );
tran (\sa_count[26][47] , \sa_count[26].f.upper[15] );
tran (\sa_count[26][48] , \sa_count[26].r.part1[16] );
tran (\sa_count[26][48] , \sa_count[26].f.upper[16] );
tran (\sa_count[26][49] , \sa_count[26].r.part1[17] );
tran (\sa_count[26][49] , \sa_count[26].f.upper[17] );
tran (\sa_count[26][50] , \sa_count[26].r.part1[18] );
tran (\sa_count[26][50] , \sa_count[26].f.unused[0] );
tran (\sa_count[26][51] , \sa_count[26].r.part1[19] );
tran (\sa_count[26][51] , \sa_count[26].f.unused[1] );
tran (\sa_count[26][52] , \sa_count[26].r.part1[20] );
tran (\sa_count[26][52] , \sa_count[26].f.unused[2] );
tran (\sa_count[26][53] , \sa_count[26].r.part1[21] );
tran (\sa_count[26][53] , \sa_count[26].f.unused[3] );
tran (\sa_count[26][54] , \sa_count[26].r.part1[22] );
tran (\sa_count[26][54] , \sa_count[26].f.unused[4] );
tran (\sa_count[26][55] , \sa_count[26].r.part1[23] );
tran (\sa_count[26][55] , \sa_count[26].f.unused[5] );
tran (\sa_count[26][56] , \sa_count[26].r.part1[24] );
tran (\sa_count[26][56] , \sa_count[26].f.unused[6] );
tran (\sa_count[26][57] , \sa_count[26].r.part1[25] );
tran (\sa_count[26][57] , \sa_count[26].f.unused[7] );
tran (\sa_count[26][58] , \sa_count[26].r.part1[26] );
tran (\sa_count[26][58] , \sa_count[26].f.unused[8] );
tran (\sa_count[26][59] , \sa_count[26].r.part1[27] );
tran (\sa_count[26][59] , \sa_count[26].f.unused[9] );
tran (\sa_count[26][60] , \sa_count[26].r.part1[28] );
tran (\sa_count[26][60] , \sa_count[26].f.unused[10] );
tran (\sa_count[26][61] , \sa_count[26].r.part1[29] );
tran (\sa_count[26][61] , \sa_count[26].f.unused[11] );
tran (\sa_count[26][62] , \sa_count[26].r.part1[30] );
tran (\sa_count[26][62] , \sa_count[26].f.unused[12] );
tran (\sa_count[26][63] , \sa_count[26].r.part1[31] );
tran (\sa_count[26][63] , \sa_count[26].f.unused[13] );
tran (\sa_count[27][0] , \sa_count[27].r.part0[0] );
tran (\sa_count[27][0] , \sa_count[27].f.lower[0] );
tran (\sa_count[27][1] , \sa_count[27].r.part0[1] );
tran (\sa_count[27][1] , \sa_count[27].f.lower[1] );
tran (\sa_count[27][2] , \sa_count[27].r.part0[2] );
tran (\sa_count[27][2] , \sa_count[27].f.lower[2] );
tran (\sa_count[27][3] , \sa_count[27].r.part0[3] );
tran (\sa_count[27][3] , \sa_count[27].f.lower[3] );
tran (\sa_count[27][4] , \sa_count[27].r.part0[4] );
tran (\sa_count[27][4] , \sa_count[27].f.lower[4] );
tran (\sa_count[27][5] , \sa_count[27].r.part0[5] );
tran (\sa_count[27][5] , \sa_count[27].f.lower[5] );
tran (\sa_count[27][6] , \sa_count[27].r.part0[6] );
tran (\sa_count[27][6] , \sa_count[27].f.lower[6] );
tran (\sa_count[27][7] , \sa_count[27].r.part0[7] );
tran (\sa_count[27][7] , \sa_count[27].f.lower[7] );
tran (\sa_count[27][8] , \sa_count[27].r.part0[8] );
tran (\sa_count[27][8] , \sa_count[27].f.lower[8] );
tran (\sa_count[27][9] , \sa_count[27].r.part0[9] );
tran (\sa_count[27][9] , \sa_count[27].f.lower[9] );
tran (\sa_count[27][10] , \sa_count[27].r.part0[10] );
tran (\sa_count[27][10] , \sa_count[27].f.lower[10] );
tran (\sa_count[27][11] , \sa_count[27].r.part0[11] );
tran (\sa_count[27][11] , \sa_count[27].f.lower[11] );
tran (\sa_count[27][12] , \sa_count[27].r.part0[12] );
tran (\sa_count[27][12] , \sa_count[27].f.lower[12] );
tran (\sa_count[27][13] , \sa_count[27].r.part0[13] );
tran (\sa_count[27][13] , \sa_count[27].f.lower[13] );
tran (\sa_count[27][14] , \sa_count[27].r.part0[14] );
tran (\sa_count[27][14] , \sa_count[27].f.lower[14] );
tran (\sa_count[27][15] , \sa_count[27].r.part0[15] );
tran (\sa_count[27][15] , \sa_count[27].f.lower[15] );
tran (\sa_count[27][16] , \sa_count[27].r.part0[16] );
tran (\sa_count[27][16] , \sa_count[27].f.lower[16] );
tran (\sa_count[27][17] , \sa_count[27].r.part0[17] );
tran (\sa_count[27][17] , \sa_count[27].f.lower[17] );
tran (\sa_count[27][18] , \sa_count[27].r.part0[18] );
tran (\sa_count[27][18] , \sa_count[27].f.lower[18] );
tran (\sa_count[27][19] , \sa_count[27].r.part0[19] );
tran (\sa_count[27][19] , \sa_count[27].f.lower[19] );
tran (\sa_count[27][20] , \sa_count[27].r.part0[20] );
tran (\sa_count[27][20] , \sa_count[27].f.lower[20] );
tran (\sa_count[27][21] , \sa_count[27].r.part0[21] );
tran (\sa_count[27][21] , \sa_count[27].f.lower[21] );
tran (\sa_count[27][22] , \sa_count[27].r.part0[22] );
tran (\sa_count[27][22] , \sa_count[27].f.lower[22] );
tran (\sa_count[27][23] , \sa_count[27].r.part0[23] );
tran (\sa_count[27][23] , \sa_count[27].f.lower[23] );
tran (\sa_count[27][24] , \sa_count[27].r.part0[24] );
tran (\sa_count[27][24] , \sa_count[27].f.lower[24] );
tran (\sa_count[27][25] , \sa_count[27].r.part0[25] );
tran (\sa_count[27][25] , \sa_count[27].f.lower[25] );
tran (\sa_count[27][26] , \sa_count[27].r.part0[26] );
tran (\sa_count[27][26] , \sa_count[27].f.lower[26] );
tran (\sa_count[27][27] , \sa_count[27].r.part0[27] );
tran (\sa_count[27][27] , \sa_count[27].f.lower[27] );
tran (\sa_count[27][28] , \sa_count[27].r.part0[28] );
tran (\sa_count[27][28] , \sa_count[27].f.lower[28] );
tran (\sa_count[27][29] , \sa_count[27].r.part0[29] );
tran (\sa_count[27][29] , \sa_count[27].f.lower[29] );
tran (\sa_count[27][30] , \sa_count[27].r.part0[30] );
tran (\sa_count[27][30] , \sa_count[27].f.lower[30] );
tran (\sa_count[27][31] , \sa_count[27].r.part0[31] );
tran (\sa_count[27][31] , \sa_count[27].f.lower[31] );
tran (\sa_count[27][32] , \sa_count[27].r.part1[0] );
tran (\sa_count[27][32] , \sa_count[27].f.upper[0] );
tran (\sa_count[27][33] , \sa_count[27].r.part1[1] );
tran (\sa_count[27][33] , \sa_count[27].f.upper[1] );
tran (\sa_count[27][34] , \sa_count[27].r.part1[2] );
tran (\sa_count[27][34] , \sa_count[27].f.upper[2] );
tran (\sa_count[27][35] , \sa_count[27].r.part1[3] );
tran (\sa_count[27][35] , \sa_count[27].f.upper[3] );
tran (\sa_count[27][36] , \sa_count[27].r.part1[4] );
tran (\sa_count[27][36] , \sa_count[27].f.upper[4] );
tran (\sa_count[27][37] , \sa_count[27].r.part1[5] );
tran (\sa_count[27][37] , \sa_count[27].f.upper[5] );
tran (\sa_count[27][38] , \sa_count[27].r.part1[6] );
tran (\sa_count[27][38] , \sa_count[27].f.upper[6] );
tran (\sa_count[27][39] , \sa_count[27].r.part1[7] );
tran (\sa_count[27][39] , \sa_count[27].f.upper[7] );
tran (\sa_count[27][40] , \sa_count[27].r.part1[8] );
tran (\sa_count[27][40] , \sa_count[27].f.upper[8] );
tran (\sa_count[27][41] , \sa_count[27].r.part1[9] );
tran (\sa_count[27][41] , \sa_count[27].f.upper[9] );
tran (\sa_count[27][42] , \sa_count[27].r.part1[10] );
tran (\sa_count[27][42] , \sa_count[27].f.upper[10] );
tran (\sa_count[27][43] , \sa_count[27].r.part1[11] );
tran (\sa_count[27][43] , \sa_count[27].f.upper[11] );
tran (\sa_count[27][44] , \sa_count[27].r.part1[12] );
tran (\sa_count[27][44] , \sa_count[27].f.upper[12] );
tran (\sa_count[27][45] , \sa_count[27].r.part1[13] );
tran (\sa_count[27][45] , \sa_count[27].f.upper[13] );
tran (\sa_count[27][46] , \sa_count[27].r.part1[14] );
tran (\sa_count[27][46] , \sa_count[27].f.upper[14] );
tran (\sa_count[27][47] , \sa_count[27].r.part1[15] );
tran (\sa_count[27][47] , \sa_count[27].f.upper[15] );
tran (\sa_count[27][48] , \sa_count[27].r.part1[16] );
tran (\sa_count[27][48] , \sa_count[27].f.upper[16] );
tran (\sa_count[27][49] , \sa_count[27].r.part1[17] );
tran (\sa_count[27][49] , \sa_count[27].f.upper[17] );
tran (\sa_count[27][50] , \sa_count[27].r.part1[18] );
tran (\sa_count[27][50] , \sa_count[27].f.unused[0] );
tran (\sa_count[27][51] , \sa_count[27].r.part1[19] );
tran (\sa_count[27][51] , \sa_count[27].f.unused[1] );
tran (\sa_count[27][52] , \sa_count[27].r.part1[20] );
tran (\sa_count[27][52] , \sa_count[27].f.unused[2] );
tran (\sa_count[27][53] , \sa_count[27].r.part1[21] );
tran (\sa_count[27][53] , \sa_count[27].f.unused[3] );
tran (\sa_count[27][54] , \sa_count[27].r.part1[22] );
tran (\sa_count[27][54] , \sa_count[27].f.unused[4] );
tran (\sa_count[27][55] , \sa_count[27].r.part1[23] );
tran (\sa_count[27][55] , \sa_count[27].f.unused[5] );
tran (\sa_count[27][56] , \sa_count[27].r.part1[24] );
tran (\sa_count[27][56] , \sa_count[27].f.unused[6] );
tran (\sa_count[27][57] , \sa_count[27].r.part1[25] );
tran (\sa_count[27][57] , \sa_count[27].f.unused[7] );
tran (\sa_count[27][58] , \sa_count[27].r.part1[26] );
tran (\sa_count[27][58] , \sa_count[27].f.unused[8] );
tran (\sa_count[27][59] , \sa_count[27].r.part1[27] );
tran (\sa_count[27][59] , \sa_count[27].f.unused[9] );
tran (\sa_count[27][60] , \sa_count[27].r.part1[28] );
tran (\sa_count[27][60] , \sa_count[27].f.unused[10] );
tran (\sa_count[27][61] , \sa_count[27].r.part1[29] );
tran (\sa_count[27][61] , \sa_count[27].f.unused[11] );
tran (\sa_count[27][62] , \sa_count[27].r.part1[30] );
tran (\sa_count[27][62] , \sa_count[27].f.unused[12] );
tran (\sa_count[27][63] , \sa_count[27].r.part1[31] );
tran (\sa_count[27][63] , \sa_count[27].f.unused[13] );
tran (\sa_count[28][0] , \sa_count[28].r.part0[0] );
tran (\sa_count[28][0] , \sa_count[28].f.lower[0] );
tran (\sa_count[28][1] , \sa_count[28].r.part0[1] );
tran (\sa_count[28][1] , \sa_count[28].f.lower[1] );
tran (\sa_count[28][2] , \sa_count[28].r.part0[2] );
tran (\sa_count[28][2] , \sa_count[28].f.lower[2] );
tran (\sa_count[28][3] , \sa_count[28].r.part0[3] );
tran (\sa_count[28][3] , \sa_count[28].f.lower[3] );
tran (\sa_count[28][4] , \sa_count[28].r.part0[4] );
tran (\sa_count[28][4] , \sa_count[28].f.lower[4] );
tran (\sa_count[28][5] , \sa_count[28].r.part0[5] );
tran (\sa_count[28][5] , \sa_count[28].f.lower[5] );
tran (\sa_count[28][6] , \sa_count[28].r.part0[6] );
tran (\sa_count[28][6] , \sa_count[28].f.lower[6] );
tran (\sa_count[28][7] , \sa_count[28].r.part0[7] );
tran (\sa_count[28][7] , \sa_count[28].f.lower[7] );
tran (\sa_count[28][8] , \sa_count[28].r.part0[8] );
tran (\sa_count[28][8] , \sa_count[28].f.lower[8] );
tran (\sa_count[28][9] , \sa_count[28].r.part0[9] );
tran (\sa_count[28][9] , \sa_count[28].f.lower[9] );
tran (\sa_count[28][10] , \sa_count[28].r.part0[10] );
tran (\sa_count[28][10] , \sa_count[28].f.lower[10] );
tran (\sa_count[28][11] , \sa_count[28].r.part0[11] );
tran (\sa_count[28][11] , \sa_count[28].f.lower[11] );
tran (\sa_count[28][12] , \sa_count[28].r.part0[12] );
tran (\sa_count[28][12] , \sa_count[28].f.lower[12] );
tran (\sa_count[28][13] , \sa_count[28].r.part0[13] );
tran (\sa_count[28][13] , \sa_count[28].f.lower[13] );
tran (\sa_count[28][14] , \sa_count[28].r.part0[14] );
tran (\sa_count[28][14] , \sa_count[28].f.lower[14] );
tran (\sa_count[28][15] , \sa_count[28].r.part0[15] );
tran (\sa_count[28][15] , \sa_count[28].f.lower[15] );
tran (\sa_count[28][16] , \sa_count[28].r.part0[16] );
tran (\sa_count[28][16] , \sa_count[28].f.lower[16] );
tran (\sa_count[28][17] , \sa_count[28].r.part0[17] );
tran (\sa_count[28][17] , \sa_count[28].f.lower[17] );
tran (\sa_count[28][18] , \sa_count[28].r.part0[18] );
tran (\sa_count[28][18] , \sa_count[28].f.lower[18] );
tran (\sa_count[28][19] , \sa_count[28].r.part0[19] );
tran (\sa_count[28][19] , \sa_count[28].f.lower[19] );
tran (\sa_count[28][20] , \sa_count[28].r.part0[20] );
tran (\sa_count[28][20] , \sa_count[28].f.lower[20] );
tran (\sa_count[28][21] , \sa_count[28].r.part0[21] );
tran (\sa_count[28][21] , \sa_count[28].f.lower[21] );
tran (\sa_count[28][22] , \sa_count[28].r.part0[22] );
tran (\sa_count[28][22] , \sa_count[28].f.lower[22] );
tran (\sa_count[28][23] , \sa_count[28].r.part0[23] );
tran (\sa_count[28][23] , \sa_count[28].f.lower[23] );
tran (\sa_count[28][24] , \sa_count[28].r.part0[24] );
tran (\sa_count[28][24] , \sa_count[28].f.lower[24] );
tran (\sa_count[28][25] , \sa_count[28].r.part0[25] );
tran (\sa_count[28][25] , \sa_count[28].f.lower[25] );
tran (\sa_count[28][26] , \sa_count[28].r.part0[26] );
tran (\sa_count[28][26] , \sa_count[28].f.lower[26] );
tran (\sa_count[28][27] , \sa_count[28].r.part0[27] );
tran (\sa_count[28][27] , \sa_count[28].f.lower[27] );
tran (\sa_count[28][28] , \sa_count[28].r.part0[28] );
tran (\sa_count[28][28] , \sa_count[28].f.lower[28] );
tran (\sa_count[28][29] , \sa_count[28].r.part0[29] );
tran (\sa_count[28][29] , \sa_count[28].f.lower[29] );
tran (\sa_count[28][30] , \sa_count[28].r.part0[30] );
tran (\sa_count[28][30] , \sa_count[28].f.lower[30] );
tran (\sa_count[28][31] , \sa_count[28].r.part0[31] );
tran (\sa_count[28][31] , \sa_count[28].f.lower[31] );
tran (\sa_count[28][32] , \sa_count[28].r.part1[0] );
tran (\sa_count[28][32] , \sa_count[28].f.upper[0] );
tran (\sa_count[28][33] , \sa_count[28].r.part1[1] );
tran (\sa_count[28][33] , \sa_count[28].f.upper[1] );
tran (\sa_count[28][34] , \sa_count[28].r.part1[2] );
tran (\sa_count[28][34] , \sa_count[28].f.upper[2] );
tran (\sa_count[28][35] , \sa_count[28].r.part1[3] );
tran (\sa_count[28][35] , \sa_count[28].f.upper[3] );
tran (\sa_count[28][36] , \sa_count[28].r.part1[4] );
tran (\sa_count[28][36] , \sa_count[28].f.upper[4] );
tran (\sa_count[28][37] , \sa_count[28].r.part1[5] );
tran (\sa_count[28][37] , \sa_count[28].f.upper[5] );
tran (\sa_count[28][38] , \sa_count[28].r.part1[6] );
tran (\sa_count[28][38] , \sa_count[28].f.upper[6] );
tran (\sa_count[28][39] , \sa_count[28].r.part1[7] );
tran (\sa_count[28][39] , \sa_count[28].f.upper[7] );
tran (\sa_count[28][40] , \sa_count[28].r.part1[8] );
tran (\sa_count[28][40] , \sa_count[28].f.upper[8] );
tran (\sa_count[28][41] , \sa_count[28].r.part1[9] );
tran (\sa_count[28][41] , \sa_count[28].f.upper[9] );
tran (\sa_count[28][42] , \sa_count[28].r.part1[10] );
tran (\sa_count[28][42] , \sa_count[28].f.upper[10] );
tran (\sa_count[28][43] , \sa_count[28].r.part1[11] );
tran (\sa_count[28][43] , \sa_count[28].f.upper[11] );
tran (\sa_count[28][44] , \sa_count[28].r.part1[12] );
tran (\sa_count[28][44] , \sa_count[28].f.upper[12] );
tran (\sa_count[28][45] , \sa_count[28].r.part1[13] );
tran (\sa_count[28][45] , \sa_count[28].f.upper[13] );
tran (\sa_count[28][46] , \sa_count[28].r.part1[14] );
tran (\sa_count[28][46] , \sa_count[28].f.upper[14] );
tran (\sa_count[28][47] , \sa_count[28].r.part1[15] );
tran (\sa_count[28][47] , \sa_count[28].f.upper[15] );
tran (\sa_count[28][48] , \sa_count[28].r.part1[16] );
tran (\sa_count[28][48] , \sa_count[28].f.upper[16] );
tran (\sa_count[28][49] , \sa_count[28].r.part1[17] );
tran (\sa_count[28][49] , \sa_count[28].f.upper[17] );
tran (\sa_count[28][50] , \sa_count[28].r.part1[18] );
tran (\sa_count[28][50] , \sa_count[28].f.unused[0] );
tran (\sa_count[28][51] , \sa_count[28].r.part1[19] );
tran (\sa_count[28][51] , \sa_count[28].f.unused[1] );
tran (\sa_count[28][52] , \sa_count[28].r.part1[20] );
tran (\sa_count[28][52] , \sa_count[28].f.unused[2] );
tran (\sa_count[28][53] , \sa_count[28].r.part1[21] );
tran (\sa_count[28][53] , \sa_count[28].f.unused[3] );
tran (\sa_count[28][54] , \sa_count[28].r.part1[22] );
tran (\sa_count[28][54] , \sa_count[28].f.unused[4] );
tran (\sa_count[28][55] , \sa_count[28].r.part1[23] );
tran (\sa_count[28][55] , \sa_count[28].f.unused[5] );
tran (\sa_count[28][56] , \sa_count[28].r.part1[24] );
tran (\sa_count[28][56] , \sa_count[28].f.unused[6] );
tran (\sa_count[28][57] , \sa_count[28].r.part1[25] );
tran (\sa_count[28][57] , \sa_count[28].f.unused[7] );
tran (\sa_count[28][58] , \sa_count[28].r.part1[26] );
tran (\sa_count[28][58] , \sa_count[28].f.unused[8] );
tran (\sa_count[28][59] , \sa_count[28].r.part1[27] );
tran (\sa_count[28][59] , \sa_count[28].f.unused[9] );
tran (\sa_count[28][60] , \sa_count[28].r.part1[28] );
tran (\sa_count[28][60] , \sa_count[28].f.unused[10] );
tran (\sa_count[28][61] , \sa_count[28].r.part1[29] );
tran (\sa_count[28][61] , \sa_count[28].f.unused[11] );
tran (\sa_count[28][62] , \sa_count[28].r.part1[30] );
tran (\sa_count[28][62] , \sa_count[28].f.unused[12] );
tran (\sa_count[28][63] , \sa_count[28].r.part1[31] );
tran (\sa_count[28][63] , \sa_count[28].f.unused[13] );
tran (\sa_count[29][0] , \sa_count[29].r.part0[0] );
tran (\sa_count[29][0] , \sa_count[29].f.lower[0] );
tran (\sa_count[29][1] , \sa_count[29].r.part0[1] );
tran (\sa_count[29][1] , \sa_count[29].f.lower[1] );
tran (\sa_count[29][2] , \sa_count[29].r.part0[2] );
tran (\sa_count[29][2] , \sa_count[29].f.lower[2] );
tran (\sa_count[29][3] , \sa_count[29].r.part0[3] );
tran (\sa_count[29][3] , \sa_count[29].f.lower[3] );
tran (\sa_count[29][4] , \sa_count[29].r.part0[4] );
tran (\sa_count[29][4] , \sa_count[29].f.lower[4] );
tran (\sa_count[29][5] , \sa_count[29].r.part0[5] );
tran (\sa_count[29][5] , \sa_count[29].f.lower[5] );
tran (\sa_count[29][6] , \sa_count[29].r.part0[6] );
tran (\sa_count[29][6] , \sa_count[29].f.lower[6] );
tran (\sa_count[29][7] , \sa_count[29].r.part0[7] );
tran (\sa_count[29][7] , \sa_count[29].f.lower[7] );
tran (\sa_count[29][8] , \sa_count[29].r.part0[8] );
tran (\sa_count[29][8] , \sa_count[29].f.lower[8] );
tran (\sa_count[29][9] , \sa_count[29].r.part0[9] );
tran (\sa_count[29][9] , \sa_count[29].f.lower[9] );
tran (\sa_count[29][10] , \sa_count[29].r.part0[10] );
tran (\sa_count[29][10] , \sa_count[29].f.lower[10] );
tran (\sa_count[29][11] , \sa_count[29].r.part0[11] );
tran (\sa_count[29][11] , \sa_count[29].f.lower[11] );
tran (\sa_count[29][12] , \sa_count[29].r.part0[12] );
tran (\sa_count[29][12] , \sa_count[29].f.lower[12] );
tran (\sa_count[29][13] , \sa_count[29].r.part0[13] );
tran (\sa_count[29][13] , \sa_count[29].f.lower[13] );
tran (\sa_count[29][14] , \sa_count[29].r.part0[14] );
tran (\sa_count[29][14] , \sa_count[29].f.lower[14] );
tran (\sa_count[29][15] , \sa_count[29].r.part0[15] );
tran (\sa_count[29][15] , \sa_count[29].f.lower[15] );
tran (\sa_count[29][16] , \sa_count[29].r.part0[16] );
tran (\sa_count[29][16] , \sa_count[29].f.lower[16] );
tran (\sa_count[29][17] , \sa_count[29].r.part0[17] );
tran (\sa_count[29][17] , \sa_count[29].f.lower[17] );
tran (\sa_count[29][18] , \sa_count[29].r.part0[18] );
tran (\sa_count[29][18] , \sa_count[29].f.lower[18] );
tran (\sa_count[29][19] , \sa_count[29].r.part0[19] );
tran (\sa_count[29][19] , \sa_count[29].f.lower[19] );
tran (\sa_count[29][20] , \sa_count[29].r.part0[20] );
tran (\sa_count[29][20] , \sa_count[29].f.lower[20] );
tran (\sa_count[29][21] , \sa_count[29].r.part0[21] );
tran (\sa_count[29][21] , \sa_count[29].f.lower[21] );
tran (\sa_count[29][22] , \sa_count[29].r.part0[22] );
tran (\sa_count[29][22] , \sa_count[29].f.lower[22] );
tran (\sa_count[29][23] , \sa_count[29].r.part0[23] );
tran (\sa_count[29][23] , \sa_count[29].f.lower[23] );
tran (\sa_count[29][24] , \sa_count[29].r.part0[24] );
tran (\sa_count[29][24] , \sa_count[29].f.lower[24] );
tran (\sa_count[29][25] , \sa_count[29].r.part0[25] );
tran (\sa_count[29][25] , \sa_count[29].f.lower[25] );
tran (\sa_count[29][26] , \sa_count[29].r.part0[26] );
tran (\sa_count[29][26] , \sa_count[29].f.lower[26] );
tran (\sa_count[29][27] , \sa_count[29].r.part0[27] );
tran (\sa_count[29][27] , \sa_count[29].f.lower[27] );
tran (\sa_count[29][28] , \sa_count[29].r.part0[28] );
tran (\sa_count[29][28] , \sa_count[29].f.lower[28] );
tran (\sa_count[29][29] , \sa_count[29].r.part0[29] );
tran (\sa_count[29][29] , \sa_count[29].f.lower[29] );
tran (\sa_count[29][30] , \sa_count[29].r.part0[30] );
tran (\sa_count[29][30] , \sa_count[29].f.lower[30] );
tran (\sa_count[29][31] , \sa_count[29].r.part0[31] );
tran (\sa_count[29][31] , \sa_count[29].f.lower[31] );
tran (\sa_count[29][32] , \sa_count[29].r.part1[0] );
tran (\sa_count[29][32] , \sa_count[29].f.upper[0] );
tran (\sa_count[29][33] , \sa_count[29].r.part1[1] );
tran (\sa_count[29][33] , \sa_count[29].f.upper[1] );
tran (\sa_count[29][34] , \sa_count[29].r.part1[2] );
tran (\sa_count[29][34] , \sa_count[29].f.upper[2] );
tran (\sa_count[29][35] , \sa_count[29].r.part1[3] );
tran (\sa_count[29][35] , \sa_count[29].f.upper[3] );
tran (\sa_count[29][36] , \sa_count[29].r.part1[4] );
tran (\sa_count[29][36] , \sa_count[29].f.upper[4] );
tran (\sa_count[29][37] , \sa_count[29].r.part1[5] );
tran (\sa_count[29][37] , \sa_count[29].f.upper[5] );
tran (\sa_count[29][38] , \sa_count[29].r.part1[6] );
tran (\sa_count[29][38] , \sa_count[29].f.upper[6] );
tran (\sa_count[29][39] , \sa_count[29].r.part1[7] );
tran (\sa_count[29][39] , \sa_count[29].f.upper[7] );
tran (\sa_count[29][40] , \sa_count[29].r.part1[8] );
tran (\sa_count[29][40] , \sa_count[29].f.upper[8] );
tran (\sa_count[29][41] , \sa_count[29].r.part1[9] );
tran (\sa_count[29][41] , \sa_count[29].f.upper[9] );
tran (\sa_count[29][42] , \sa_count[29].r.part1[10] );
tran (\sa_count[29][42] , \sa_count[29].f.upper[10] );
tran (\sa_count[29][43] , \sa_count[29].r.part1[11] );
tran (\sa_count[29][43] , \sa_count[29].f.upper[11] );
tran (\sa_count[29][44] , \sa_count[29].r.part1[12] );
tran (\sa_count[29][44] , \sa_count[29].f.upper[12] );
tran (\sa_count[29][45] , \sa_count[29].r.part1[13] );
tran (\sa_count[29][45] , \sa_count[29].f.upper[13] );
tran (\sa_count[29][46] , \sa_count[29].r.part1[14] );
tran (\sa_count[29][46] , \sa_count[29].f.upper[14] );
tran (\sa_count[29][47] , \sa_count[29].r.part1[15] );
tran (\sa_count[29][47] , \sa_count[29].f.upper[15] );
tran (\sa_count[29][48] , \sa_count[29].r.part1[16] );
tran (\sa_count[29][48] , \sa_count[29].f.upper[16] );
tran (\sa_count[29][49] , \sa_count[29].r.part1[17] );
tran (\sa_count[29][49] , \sa_count[29].f.upper[17] );
tran (\sa_count[29][50] , \sa_count[29].r.part1[18] );
tran (\sa_count[29][50] , \sa_count[29].f.unused[0] );
tran (\sa_count[29][51] , \sa_count[29].r.part1[19] );
tran (\sa_count[29][51] , \sa_count[29].f.unused[1] );
tran (\sa_count[29][52] , \sa_count[29].r.part1[20] );
tran (\sa_count[29][52] , \sa_count[29].f.unused[2] );
tran (\sa_count[29][53] , \sa_count[29].r.part1[21] );
tran (\sa_count[29][53] , \sa_count[29].f.unused[3] );
tran (\sa_count[29][54] , \sa_count[29].r.part1[22] );
tran (\sa_count[29][54] , \sa_count[29].f.unused[4] );
tran (\sa_count[29][55] , \sa_count[29].r.part1[23] );
tran (\sa_count[29][55] , \sa_count[29].f.unused[5] );
tran (\sa_count[29][56] , \sa_count[29].r.part1[24] );
tran (\sa_count[29][56] , \sa_count[29].f.unused[6] );
tran (\sa_count[29][57] , \sa_count[29].r.part1[25] );
tran (\sa_count[29][57] , \sa_count[29].f.unused[7] );
tran (\sa_count[29][58] , \sa_count[29].r.part1[26] );
tran (\sa_count[29][58] , \sa_count[29].f.unused[8] );
tran (\sa_count[29][59] , \sa_count[29].r.part1[27] );
tran (\sa_count[29][59] , \sa_count[29].f.unused[9] );
tran (\sa_count[29][60] , \sa_count[29].r.part1[28] );
tran (\sa_count[29][60] , \sa_count[29].f.unused[10] );
tran (\sa_count[29][61] , \sa_count[29].r.part1[29] );
tran (\sa_count[29][61] , \sa_count[29].f.unused[11] );
tran (\sa_count[29][62] , \sa_count[29].r.part1[30] );
tran (\sa_count[29][62] , \sa_count[29].f.unused[12] );
tran (\sa_count[29][63] , \sa_count[29].r.part1[31] );
tran (\sa_count[29][63] , \sa_count[29].f.unused[13] );
tran (\sa_count[30][0] , \sa_count[30].r.part0[0] );
tran (\sa_count[30][0] , \sa_count[30].f.lower[0] );
tran (\sa_count[30][1] , \sa_count[30].r.part0[1] );
tran (\sa_count[30][1] , \sa_count[30].f.lower[1] );
tran (\sa_count[30][2] , \sa_count[30].r.part0[2] );
tran (\sa_count[30][2] , \sa_count[30].f.lower[2] );
tran (\sa_count[30][3] , \sa_count[30].r.part0[3] );
tran (\sa_count[30][3] , \sa_count[30].f.lower[3] );
tran (\sa_count[30][4] , \sa_count[30].r.part0[4] );
tran (\sa_count[30][4] , \sa_count[30].f.lower[4] );
tran (\sa_count[30][5] , \sa_count[30].r.part0[5] );
tran (\sa_count[30][5] , \sa_count[30].f.lower[5] );
tran (\sa_count[30][6] , \sa_count[30].r.part0[6] );
tran (\sa_count[30][6] , \sa_count[30].f.lower[6] );
tran (\sa_count[30][7] , \sa_count[30].r.part0[7] );
tran (\sa_count[30][7] , \sa_count[30].f.lower[7] );
tran (\sa_count[30][8] , \sa_count[30].r.part0[8] );
tran (\sa_count[30][8] , \sa_count[30].f.lower[8] );
tran (\sa_count[30][9] , \sa_count[30].r.part0[9] );
tran (\sa_count[30][9] , \sa_count[30].f.lower[9] );
tran (\sa_count[30][10] , \sa_count[30].r.part0[10] );
tran (\sa_count[30][10] , \sa_count[30].f.lower[10] );
tran (\sa_count[30][11] , \sa_count[30].r.part0[11] );
tran (\sa_count[30][11] , \sa_count[30].f.lower[11] );
tran (\sa_count[30][12] , \sa_count[30].r.part0[12] );
tran (\sa_count[30][12] , \sa_count[30].f.lower[12] );
tran (\sa_count[30][13] , \sa_count[30].r.part0[13] );
tran (\sa_count[30][13] , \sa_count[30].f.lower[13] );
tran (\sa_count[30][14] , \sa_count[30].r.part0[14] );
tran (\sa_count[30][14] , \sa_count[30].f.lower[14] );
tran (\sa_count[30][15] , \sa_count[30].r.part0[15] );
tran (\sa_count[30][15] , \sa_count[30].f.lower[15] );
tran (\sa_count[30][16] , \sa_count[30].r.part0[16] );
tran (\sa_count[30][16] , \sa_count[30].f.lower[16] );
tran (\sa_count[30][17] , \sa_count[30].r.part0[17] );
tran (\sa_count[30][17] , \sa_count[30].f.lower[17] );
tran (\sa_count[30][18] , \sa_count[30].r.part0[18] );
tran (\sa_count[30][18] , \sa_count[30].f.lower[18] );
tran (\sa_count[30][19] , \sa_count[30].r.part0[19] );
tran (\sa_count[30][19] , \sa_count[30].f.lower[19] );
tran (\sa_count[30][20] , \sa_count[30].r.part0[20] );
tran (\sa_count[30][20] , \sa_count[30].f.lower[20] );
tran (\sa_count[30][21] , \sa_count[30].r.part0[21] );
tran (\sa_count[30][21] , \sa_count[30].f.lower[21] );
tran (\sa_count[30][22] , \sa_count[30].r.part0[22] );
tran (\sa_count[30][22] , \sa_count[30].f.lower[22] );
tran (\sa_count[30][23] , \sa_count[30].r.part0[23] );
tran (\sa_count[30][23] , \sa_count[30].f.lower[23] );
tran (\sa_count[30][24] , \sa_count[30].r.part0[24] );
tran (\sa_count[30][24] , \sa_count[30].f.lower[24] );
tran (\sa_count[30][25] , \sa_count[30].r.part0[25] );
tran (\sa_count[30][25] , \sa_count[30].f.lower[25] );
tran (\sa_count[30][26] , \sa_count[30].r.part0[26] );
tran (\sa_count[30][26] , \sa_count[30].f.lower[26] );
tran (\sa_count[30][27] , \sa_count[30].r.part0[27] );
tran (\sa_count[30][27] , \sa_count[30].f.lower[27] );
tran (\sa_count[30][28] , \sa_count[30].r.part0[28] );
tran (\sa_count[30][28] , \sa_count[30].f.lower[28] );
tran (\sa_count[30][29] , \sa_count[30].r.part0[29] );
tran (\sa_count[30][29] , \sa_count[30].f.lower[29] );
tran (\sa_count[30][30] , \sa_count[30].r.part0[30] );
tran (\sa_count[30][30] , \sa_count[30].f.lower[30] );
tran (\sa_count[30][31] , \sa_count[30].r.part0[31] );
tran (\sa_count[30][31] , \sa_count[30].f.lower[31] );
tran (\sa_count[30][32] , \sa_count[30].r.part1[0] );
tran (\sa_count[30][32] , \sa_count[30].f.upper[0] );
tran (\sa_count[30][33] , \sa_count[30].r.part1[1] );
tran (\sa_count[30][33] , \sa_count[30].f.upper[1] );
tran (\sa_count[30][34] , \sa_count[30].r.part1[2] );
tran (\sa_count[30][34] , \sa_count[30].f.upper[2] );
tran (\sa_count[30][35] , \sa_count[30].r.part1[3] );
tran (\sa_count[30][35] , \sa_count[30].f.upper[3] );
tran (\sa_count[30][36] , \sa_count[30].r.part1[4] );
tran (\sa_count[30][36] , \sa_count[30].f.upper[4] );
tran (\sa_count[30][37] , \sa_count[30].r.part1[5] );
tran (\sa_count[30][37] , \sa_count[30].f.upper[5] );
tran (\sa_count[30][38] , \sa_count[30].r.part1[6] );
tran (\sa_count[30][38] , \sa_count[30].f.upper[6] );
tran (\sa_count[30][39] , \sa_count[30].r.part1[7] );
tran (\sa_count[30][39] , \sa_count[30].f.upper[7] );
tran (\sa_count[30][40] , \sa_count[30].r.part1[8] );
tran (\sa_count[30][40] , \sa_count[30].f.upper[8] );
tran (\sa_count[30][41] , \sa_count[30].r.part1[9] );
tran (\sa_count[30][41] , \sa_count[30].f.upper[9] );
tran (\sa_count[30][42] , \sa_count[30].r.part1[10] );
tran (\sa_count[30][42] , \sa_count[30].f.upper[10] );
tran (\sa_count[30][43] , \sa_count[30].r.part1[11] );
tran (\sa_count[30][43] , \sa_count[30].f.upper[11] );
tran (\sa_count[30][44] , \sa_count[30].r.part1[12] );
tran (\sa_count[30][44] , \sa_count[30].f.upper[12] );
tran (\sa_count[30][45] , \sa_count[30].r.part1[13] );
tran (\sa_count[30][45] , \sa_count[30].f.upper[13] );
tran (\sa_count[30][46] , \sa_count[30].r.part1[14] );
tran (\sa_count[30][46] , \sa_count[30].f.upper[14] );
tran (\sa_count[30][47] , \sa_count[30].r.part1[15] );
tran (\sa_count[30][47] , \sa_count[30].f.upper[15] );
tran (\sa_count[30][48] , \sa_count[30].r.part1[16] );
tran (\sa_count[30][48] , \sa_count[30].f.upper[16] );
tran (\sa_count[30][49] , \sa_count[30].r.part1[17] );
tran (\sa_count[30][49] , \sa_count[30].f.upper[17] );
tran (\sa_count[30][50] , \sa_count[30].r.part1[18] );
tran (\sa_count[30][50] , \sa_count[30].f.unused[0] );
tran (\sa_count[30][51] , \sa_count[30].r.part1[19] );
tran (\sa_count[30][51] , \sa_count[30].f.unused[1] );
tran (\sa_count[30][52] , \sa_count[30].r.part1[20] );
tran (\sa_count[30][52] , \sa_count[30].f.unused[2] );
tran (\sa_count[30][53] , \sa_count[30].r.part1[21] );
tran (\sa_count[30][53] , \sa_count[30].f.unused[3] );
tran (\sa_count[30][54] , \sa_count[30].r.part1[22] );
tran (\sa_count[30][54] , \sa_count[30].f.unused[4] );
tran (\sa_count[30][55] , \sa_count[30].r.part1[23] );
tran (\sa_count[30][55] , \sa_count[30].f.unused[5] );
tran (\sa_count[30][56] , \sa_count[30].r.part1[24] );
tran (\sa_count[30][56] , \sa_count[30].f.unused[6] );
tran (\sa_count[30][57] , \sa_count[30].r.part1[25] );
tran (\sa_count[30][57] , \sa_count[30].f.unused[7] );
tran (\sa_count[30][58] , \sa_count[30].r.part1[26] );
tran (\sa_count[30][58] , \sa_count[30].f.unused[8] );
tran (\sa_count[30][59] , \sa_count[30].r.part1[27] );
tran (\sa_count[30][59] , \sa_count[30].f.unused[9] );
tran (\sa_count[30][60] , \sa_count[30].r.part1[28] );
tran (\sa_count[30][60] , \sa_count[30].f.unused[10] );
tran (\sa_count[30][61] , \sa_count[30].r.part1[29] );
tran (\sa_count[30][61] , \sa_count[30].f.unused[11] );
tran (\sa_count[30][62] , \sa_count[30].r.part1[30] );
tran (\sa_count[30][62] , \sa_count[30].f.unused[12] );
tran (\sa_count[30][63] , \sa_count[30].r.part1[31] );
tran (\sa_count[30][63] , \sa_count[30].f.unused[13] );
tran (\sa_count[31][0] , \sa_count[31].r.part0[0] );
tran (\sa_count[31][0] , \sa_count[31].f.lower[0] );
tran (\sa_count[31][1] , \sa_count[31].r.part0[1] );
tran (\sa_count[31][1] , \sa_count[31].f.lower[1] );
tran (\sa_count[31][2] , \sa_count[31].r.part0[2] );
tran (\sa_count[31][2] , \sa_count[31].f.lower[2] );
tran (\sa_count[31][3] , \sa_count[31].r.part0[3] );
tran (\sa_count[31][3] , \sa_count[31].f.lower[3] );
tran (\sa_count[31][4] , \sa_count[31].r.part0[4] );
tran (\sa_count[31][4] , \sa_count[31].f.lower[4] );
tran (\sa_count[31][5] , \sa_count[31].r.part0[5] );
tran (\sa_count[31][5] , \sa_count[31].f.lower[5] );
tran (\sa_count[31][6] , \sa_count[31].r.part0[6] );
tran (\sa_count[31][6] , \sa_count[31].f.lower[6] );
tran (\sa_count[31][7] , \sa_count[31].r.part0[7] );
tran (\sa_count[31][7] , \sa_count[31].f.lower[7] );
tran (\sa_count[31][8] , \sa_count[31].r.part0[8] );
tran (\sa_count[31][8] , \sa_count[31].f.lower[8] );
tran (\sa_count[31][9] , \sa_count[31].r.part0[9] );
tran (\sa_count[31][9] , \sa_count[31].f.lower[9] );
tran (\sa_count[31][10] , \sa_count[31].r.part0[10] );
tran (\sa_count[31][10] , \sa_count[31].f.lower[10] );
tran (\sa_count[31][11] , \sa_count[31].r.part0[11] );
tran (\sa_count[31][11] , \sa_count[31].f.lower[11] );
tran (\sa_count[31][12] , \sa_count[31].r.part0[12] );
tran (\sa_count[31][12] , \sa_count[31].f.lower[12] );
tran (\sa_count[31][13] , \sa_count[31].r.part0[13] );
tran (\sa_count[31][13] , \sa_count[31].f.lower[13] );
tran (\sa_count[31][14] , \sa_count[31].r.part0[14] );
tran (\sa_count[31][14] , \sa_count[31].f.lower[14] );
tran (\sa_count[31][15] , \sa_count[31].r.part0[15] );
tran (\sa_count[31][15] , \sa_count[31].f.lower[15] );
tran (\sa_count[31][16] , \sa_count[31].r.part0[16] );
tran (\sa_count[31][16] , \sa_count[31].f.lower[16] );
tran (\sa_count[31][17] , \sa_count[31].r.part0[17] );
tran (\sa_count[31][17] , \sa_count[31].f.lower[17] );
tran (\sa_count[31][18] , \sa_count[31].r.part0[18] );
tran (\sa_count[31][18] , \sa_count[31].f.lower[18] );
tran (\sa_count[31][19] , \sa_count[31].r.part0[19] );
tran (\sa_count[31][19] , \sa_count[31].f.lower[19] );
tran (\sa_count[31][20] , \sa_count[31].r.part0[20] );
tran (\sa_count[31][20] , \sa_count[31].f.lower[20] );
tran (\sa_count[31][21] , \sa_count[31].r.part0[21] );
tran (\sa_count[31][21] , \sa_count[31].f.lower[21] );
tran (\sa_count[31][22] , \sa_count[31].r.part0[22] );
tran (\sa_count[31][22] , \sa_count[31].f.lower[22] );
tran (\sa_count[31][23] , \sa_count[31].r.part0[23] );
tran (\sa_count[31][23] , \sa_count[31].f.lower[23] );
tran (\sa_count[31][24] , \sa_count[31].r.part0[24] );
tran (\sa_count[31][24] , \sa_count[31].f.lower[24] );
tran (\sa_count[31][25] , \sa_count[31].r.part0[25] );
tran (\sa_count[31][25] , \sa_count[31].f.lower[25] );
tran (\sa_count[31][26] , \sa_count[31].r.part0[26] );
tran (\sa_count[31][26] , \sa_count[31].f.lower[26] );
tran (\sa_count[31][27] , \sa_count[31].r.part0[27] );
tran (\sa_count[31][27] , \sa_count[31].f.lower[27] );
tran (\sa_count[31][28] , \sa_count[31].r.part0[28] );
tran (\sa_count[31][28] , \sa_count[31].f.lower[28] );
tran (\sa_count[31][29] , \sa_count[31].r.part0[29] );
tran (\sa_count[31][29] , \sa_count[31].f.lower[29] );
tran (\sa_count[31][30] , \sa_count[31].r.part0[30] );
tran (\sa_count[31][30] , \sa_count[31].f.lower[30] );
tran (\sa_count[31][31] , \sa_count[31].r.part0[31] );
tran (\sa_count[31][31] , \sa_count[31].f.lower[31] );
tran (\sa_count[31][32] , \sa_count[31].r.part1[0] );
tran (\sa_count[31][32] , \sa_count[31].f.upper[0] );
tran (\sa_count[31][33] , \sa_count[31].r.part1[1] );
tran (\sa_count[31][33] , \sa_count[31].f.upper[1] );
tran (\sa_count[31][34] , \sa_count[31].r.part1[2] );
tran (\sa_count[31][34] , \sa_count[31].f.upper[2] );
tran (\sa_count[31][35] , \sa_count[31].r.part1[3] );
tran (\sa_count[31][35] , \sa_count[31].f.upper[3] );
tran (\sa_count[31][36] , \sa_count[31].r.part1[4] );
tran (\sa_count[31][36] , \sa_count[31].f.upper[4] );
tran (\sa_count[31][37] , \sa_count[31].r.part1[5] );
tran (\sa_count[31][37] , \sa_count[31].f.upper[5] );
tran (\sa_count[31][38] , \sa_count[31].r.part1[6] );
tran (\sa_count[31][38] , \sa_count[31].f.upper[6] );
tran (\sa_count[31][39] , \sa_count[31].r.part1[7] );
tran (\sa_count[31][39] , \sa_count[31].f.upper[7] );
tran (\sa_count[31][40] , \sa_count[31].r.part1[8] );
tran (\sa_count[31][40] , \sa_count[31].f.upper[8] );
tran (\sa_count[31][41] , \sa_count[31].r.part1[9] );
tran (\sa_count[31][41] , \sa_count[31].f.upper[9] );
tran (\sa_count[31][42] , \sa_count[31].r.part1[10] );
tran (\sa_count[31][42] , \sa_count[31].f.upper[10] );
tran (\sa_count[31][43] , \sa_count[31].r.part1[11] );
tran (\sa_count[31][43] , \sa_count[31].f.upper[11] );
tran (\sa_count[31][44] , \sa_count[31].r.part1[12] );
tran (\sa_count[31][44] , \sa_count[31].f.upper[12] );
tran (\sa_count[31][45] , \sa_count[31].r.part1[13] );
tran (\sa_count[31][45] , \sa_count[31].f.upper[13] );
tran (\sa_count[31][46] , \sa_count[31].r.part1[14] );
tran (\sa_count[31][46] , \sa_count[31].f.upper[14] );
tran (\sa_count[31][47] , \sa_count[31].r.part1[15] );
tran (\sa_count[31][47] , \sa_count[31].f.upper[15] );
tran (\sa_count[31][48] , \sa_count[31].r.part1[16] );
tran (\sa_count[31][48] , \sa_count[31].f.upper[16] );
tran (\sa_count[31][49] , \sa_count[31].r.part1[17] );
tran (\sa_count[31][49] , \sa_count[31].f.upper[17] );
tran (\sa_count[31][50] , \sa_count[31].r.part1[18] );
tran (\sa_count[31][50] , \sa_count[31].f.unused[0] );
tran (\sa_count[31][51] , \sa_count[31].r.part1[19] );
tran (\sa_count[31][51] , \sa_count[31].f.unused[1] );
tran (\sa_count[31][52] , \sa_count[31].r.part1[20] );
tran (\sa_count[31][52] , \sa_count[31].f.unused[2] );
tran (\sa_count[31][53] , \sa_count[31].r.part1[21] );
tran (\sa_count[31][53] , \sa_count[31].f.unused[3] );
tran (\sa_count[31][54] , \sa_count[31].r.part1[22] );
tran (\sa_count[31][54] , \sa_count[31].f.unused[4] );
tran (\sa_count[31][55] , \sa_count[31].r.part1[23] );
tran (\sa_count[31][55] , \sa_count[31].f.unused[5] );
tran (\sa_count[31][56] , \sa_count[31].r.part1[24] );
tran (\sa_count[31][56] , \sa_count[31].f.unused[6] );
tran (\sa_count[31][57] , \sa_count[31].r.part1[25] );
tran (\sa_count[31][57] , \sa_count[31].f.unused[7] );
tran (\sa_count[31][58] , \sa_count[31].r.part1[26] );
tran (\sa_count[31][58] , \sa_count[31].f.unused[8] );
tran (\sa_count[31][59] , \sa_count[31].r.part1[27] );
tran (\sa_count[31][59] , \sa_count[31].f.unused[9] );
tran (\sa_count[31][60] , \sa_count[31].r.part1[28] );
tran (\sa_count[31][60] , \sa_count[31].f.unused[10] );
tran (\sa_count[31][61] , \sa_count[31].r.part1[29] );
tran (\sa_count[31][61] , \sa_count[31].f.unused[11] );
tran (\sa_count[31][62] , \sa_count[31].r.part1[30] );
tran (\sa_count[31][62] , \sa_count[31].f.unused[12] );
tran (\sa_count[31][63] , \sa_count[31].r.part1[31] );
tran (\sa_count[31][63] , \sa_count[31].f.unused[13] );
tran (idle_components[31], \idle_components.r.part0 [31]);
tran (idle_components[31], \idle_components.f.num_key_tlvs_in_flight [19]);
tran (idle_components[30], \idle_components.r.part0 [30]);
tran (idle_components[30], \idle_components.f.num_key_tlvs_in_flight [18]);
tran (idle_components[29], \idle_components.r.part0 [29]);
tran (idle_components[29], \idle_components.f.num_key_tlvs_in_flight [17]);
tran (idle_components[28], \idle_components.r.part0 [28]);
tran (idle_components[28], \idle_components.f.num_key_tlvs_in_flight [16]);
tran (idle_components[27], \idle_components.r.part0 [27]);
tran (idle_components[27], \idle_components.f.num_key_tlvs_in_flight [15]);
tran (idle_components[26], \idle_components.r.part0 [26]);
tran (idle_components[26], \idle_components.f.num_key_tlvs_in_flight [14]);
tran (idle_components[25], \idle_components.r.part0 [25]);
tran (idle_components[25], \idle_components.f.num_key_tlvs_in_flight [13]);
tran (idle_components[24], \idle_components.r.part0 [24]);
tran (idle_components[24], \idle_components.f.num_key_tlvs_in_flight [12]);
tran (idle_components[23], \idle_components.r.part0 [23]);
tran (idle_components[23], \idle_components.f.num_key_tlvs_in_flight [11]);
tran (idle_components[22], \idle_components.r.part0 [22]);
tran (idle_components[22], \idle_components.f.num_key_tlvs_in_flight [10]);
tran (idle_components[21], \idle_components.r.part0 [21]);
tran (idle_components[21], \idle_components.f.num_key_tlvs_in_flight [9]);
tran (idle_components[20], \idle_components.r.part0 [20]);
tran (idle_components[20], \idle_components.f.num_key_tlvs_in_flight [8]);
tran (idle_components[19], \idle_components.r.part0 [19]);
tran (idle_components[19], \idle_components.f.num_key_tlvs_in_flight [7]);
tran (idle_components[18], \idle_components.r.part0 [18]);
tran (idle_components[18], \idle_components.f.num_key_tlvs_in_flight [6]);
tran (idle_components[17], \idle_components.r.part0 [17]);
tran (idle_components[17], \idle_components.f.num_key_tlvs_in_flight [5]);
tran (idle_components[16], \idle_components.r.part0 [16]);
tran (idle_components[16], \idle_components.f.num_key_tlvs_in_flight [4]);
tran (idle_components[15], \idle_components.r.part0 [15]);
tran (idle_components[15], \idle_components.f.num_key_tlvs_in_flight [3]);
tran (idle_components[14], \idle_components.r.part0 [14]);
tran (idle_components[14], \idle_components.f.num_key_tlvs_in_flight [2]);
tran (idle_components[13], \idle_components.r.part0 [13]);
tran (idle_components[13], \idle_components.f.num_key_tlvs_in_flight [1]);
tran (idle_components[12], \idle_components.r.part0 [12]);
tran (idle_components[12], \idle_components.f.num_key_tlvs_in_flight [0]);
tran (idle_components[11], \idle_components.r.part0 [11]);
tran (idle_components[11], \idle_components.f.cddip0_key_tlv_rsm_idle );
tran (idle_components[10], \idle_components.r.part0 [10]);
tran (idle_components[10], \idle_components.f.cddip1_key_tlv_rsm_idle );
tran (idle_components[9], \idle_components.r.part0 [9]);
tran (idle_components[9], \idle_components.f.cddip2_key_tlv_rsm_idle );
tran (idle_components[8], \idle_components.r.part0 [8]);
tran (idle_components[8], \idle_components.f.cddip3_key_tlv_rsm_idle );
tran (idle_components[7], \idle_components.r.part0 [7]);
tran (idle_components[7], \idle_components.f.cceip0_key_tlv_rsm_idle );
tran (idle_components[6], \idle_components.r.part0 [6]);
tran (idle_components[6], \idle_components.f.cceip1_key_tlv_rsm_idle );
tran (idle_components[5], \idle_components.r.part0 [5]);
tran (idle_components[5], \idle_components.f.cceip2_key_tlv_rsm_idle );
tran (idle_components[4], \idle_components.r.part0 [4]);
tran (idle_components[4], \idle_components.f.cceip3_key_tlv_rsm_idle );
tran (idle_components[3], \idle_components.r.part0 [3]);
tran (idle_components[3], \idle_components.f.no_key_tlv_in_flight );
tran (idle_components[2], \idle_components.r.part0 [2]);
tran (idle_components[2], \idle_components.f.tlv_parser_idle );
tran (idle_components[1], \idle_components.r.part0 [1]);
tran (idle_components[1], \idle_components.f.drng_idle );
tran (idle_components[0], \idle_components.r.part0 [0]);
tran (idle_components[0], \idle_components.f.kme_slv_empty );
tran (tready_override[8], \tready_override.r.part0 [8]);
tran (tready_override[8], \tready_override.f.txc_tready_override );
tran (tready_override[7], \tready_override.r.part0 [7]);
tran (tready_override[7], \tready_override.f.engine_7_tready_override );
tran (tready_override[6], \tready_override.r.part0 [6]);
tran (tready_override[6], \tready_override.f.engine_6_tready_override );
tran (tready_override[5], \tready_override.r.part0 [5]);
tran (tready_override[5], \tready_override.f.engine_5_tready_override );
tran (tready_override[4], \tready_override.r.part0 [4]);
tran (tready_override[4], \tready_override.f.engine_4_tready_override );
tran (tready_override[3], \tready_override.r.part0 [3]);
tran (tready_override[3], \tready_override.f.engine_3_tready_override );
tran (tready_override[2], \tready_override.r.part0 [2]);
tran (tready_override[2], \tready_override.f.engine_2_tready_override );
tran (tready_override[1], \tready_override.r.part0 [1]);
tran (tready_override[1], \tready_override.f.engine_1_tready_override );
tran (tready_override[0], \tready_override.r.part0 [0]);
tran (tready_override[0], \tready_override.f.engine_0_tready_override );
tran (core_kme_ib_out[0], \core_kme_ib_out.tready );
tran (sa_global_ctrl[31], \sa_global_ctrl.r.part0 [31]);
tran (sa_global_ctrl[31], \sa_global_ctrl.f.spare [29]);
tran (sa_global_ctrl[30], \sa_global_ctrl.r.part0 [30]);
tran (sa_global_ctrl[30], \sa_global_ctrl.f.spare [28]);
tran (sa_global_ctrl[29], \sa_global_ctrl.r.part0 [29]);
tran (sa_global_ctrl[29], \sa_global_ctrl.f.spare [27]);
tran (sa_global_ctrl[28], \sa_global_ctrl.r.part0 [28]);
tran (sa_global_ctrl[28], \sa_global_ctrl.f.spare [26]);
tran (sa_global_ctrl[27], \sa_global_ctrl.r.part0 [27]);
tran (sa_global_ctrl[27], \sa_global_ctrl.f.spare [25]);
tran (sa_global_ctrl[26], \sa_global_ctrl.r.part0 [26]);
tran (sa_global_ctrl[26], \sa_global_ctrl.f.spare [24]);
tran (sa_global_ctrl[25], \sa_global_ctrl.r.part0 [25]);
tran (sa_global_ctrl[25], \sa_global_ctrl.f.spare [23]);
tran (sa_global_ctrl[24], \sa_global_ctrl.r.part0 [24]);
tran (sa_global_ctrl[24], \sa_global_ctrl.f.spare [22]);
tran (sa_global_ctrl[23], \sa_global_ctrl.r.part0 [23]);
tran (sa_global_ctrl[23], \sa_global_ctrl.f.spare [21]);
tran (sa_global_ctrl[22], \sa_global_ctrl.r.part0 [22]);
tran (sa_global_ctrl[22], \sa_global_ctrl.f.spare [20]);
tran (sa_global_ctrl[21], \sa_global_ctrl.r.part0 [21]);
tran (sa_global_ctrl[21], \sa_global_ctrl.f.spare [19]);
tran (sa_global_ctrl[20], \sa_global_ctrl.r.part0 [20]);
tran (sa_global_ctrl[20], \sa_global_ctrl.f.spare [18]);
tran (sa_global_ctrl[19], \sa_global_ctrl.r.part0 [19]);
tran (sa_global_ctrl[19], \sa_global_ctrl.f.spare [17]);
tran (sa_global_ctrl[18], \sa_global_ctrl.r.part0 [18]);
tran (sa_global_ctrl[18], \sa_global_ctrl.f.spare [16]);
tran (sa_global_ctrl[17], \sa_global_ctrl.r.part0 [17]);
tran (sa_global_ctrl[17], \sa_global_ctrl.f.spare [15]);
tran (sa_global_ctrl[16], \sa_global_ctrl.r.part0 [16]);
tran (sa_global_ctrl[16], \sa_global_ctrl.f.spare [14]);
tran (sa_global_ctrl[15], \sa_global_ctrl.r.part0 [15]);
tran (sa_global_ctrl[15], \sa_global_ctrl.f.spare [13]);
tran (sa_global_ctrl[14], \sa_global_ctrl.r.part0 [14]);
tran (sa_global_ctrl[14], \sa_global_ctrl.f.spare [12]);
tran (sa_global_ctrl[13], \sa_global_ctrl.r.part0 [13]);
tran (sa_global_ctrl[13], \sa_global_ctrl.f.spare [11]);
tran (sa_global_ctrl[12], \sa_global_ctrl.r.part0 [12]);
tran (sa_global_ctrl[12], \sa_global_ctrl.f.spare [10]);
tran (sa_global_ctrl[11], \sa_global_ctrl.r.part0 [11]);
tran (sa_global_ctrl[11], \sa_global_ctrl.f.spare [9]);
tran (sa_global_ctrl[10], \sa_global_ctrl.r.part0 [10]);
tran (sa_global_ctrl[10], \sa_global_ctrl.f.spare [8]);
tran (sa_global_ctrl[9], \sa_global_ctrl.r.part0 [9]);
tran (sa_global_ctrl[9], \sa_global_ctrl.f.spare [7]);
tran (sa_global_ctrl[8], \sa_global_ctrl.r.part0 [8]);
tran (sa_global_ctrl[8], \sa_global_ctrl.f.spare [6]);
tran (sa_global_ctrl[7], \sa_global_ctrl.r.part0 [7]);
tran (sa_global_ctrl[7], \sa_global_ctrl.f.spare [5]);
tran (sa_global_ctrl[6], \sa_global_ctrl.r.part0 [6]);
tran (sa_global_ctrl[6], \sa_global_ctrl.f.spare [4]);
tran (sa_global_ctrl[5], \sa_global_ctrl.r.part0 [5]);
tran (sa_global_ctrl[5], \sa_global_ctrl.f.spare [3]);
tran (sa_global_ctrl[4], \sa_global_ctrl.r.part0 [4]);
tran (sa_global_ctrl[4], \sa_global_ctrl.f.spare [2]);
tran (sa_global_ctrl[3], \sa_global_ctrl.r.part0 [3]);
tran (sa_global_ctrl[3], \sa_global_ctrl.f.spare [1]);
tran (sa_global_ctrl[2], \sa_global_ctrl.r.part0 [2]);
tran (sa_global_ctrl[2], \sa_global_ctrl.f.spare [0]);
tran (sa_global_ctrl[1], \sa_global_ctrl.r.part0 [1]);
tran (sa_global_ctrl[1], \sa_global_ctrl.f.sa_snap );
tran (sa_global_ctrl[0], \sa_global_ctrl.r.part0 [0]);
tran (sa_global_ctrl[0], \sa_global_ctrl.f.sa_clear_live );
tran (\sa_ctrl[0][0] , \sa_ctrl[0].r.part0[0] );
tran (\sa_ctrl[0][0] , \sa_ctrl[0].f.sa_event_sel[0] );
tran (\sa_ctrl[0][1] , \sa_ctrl[0].r.part0[1] );
tran (\sa_ctrl[0][1] , \sa_ctrl[0].f.sa_event_sel[1] );
tran (\sa_ctrl[0][2] , \sa_ctrl[0].r.part0[2] );
tran (\sa_ctrl[0][2] , \sa_ctrl[0].f.sa_event_sel[2] );
tran (\sa_ctrl[0][3] , \sa_ctrl[0].r.part0[3] );
tran (\sa_ctrl[0][3] , \sa_ctrl[0].f.sa_event_sel[3] );
tran (\sa_ctrl[0][4] , \sa_ctrl[0].r.part0[4] );
tran (\sa_ctrl[0][4] , \sa_ctrl[0].f.sa_event_sel[4] );
tran (\sa_ctrl[0][5] , \sa_ctrl[0].r.part0[5] );
tran (\sa_ctrl[0][5] , \sa_ctrl[0].f.spare[0] );
tran (\sa_ctrl[0][6] , \sa_ctrl[0].r.part0[6] );
tran (\sa_ctrl[0][6] , \sa_ctrl[0].f.spare[1] );
tran (\sa_ctrl[0][7] , \sa_ctrl[0].r.part0[7] );
tran (\sa_ctrl[0][7] , \sa_ctrl[0].f.spare[2] );
tran (\sa_ctrl[0][8] , \sa_ctrl[0].r.part0[8] );
tran (\sa_ctrl[0][8] , \sa_ctrl[0].f.spare[3] );
tran (\sa_ctrl[0][9] , \sa_ctrl[0].r.part0[9] );
tran (\sa_ctrl[0][9] , \sa_ctrl[0].f.spare[4] );
tran (\sa_ctrl[0][10] , \sa_ctrl[0].r.part0[10] );
tran (\sa_ctrl[0][10] , \sa_ctrl[0].f.spare[5] );
tran (\sa_ctrl[0][11] , \sa_ctrl[0].r.part0[11] );
tran (\sa_ctrl[0][11] , \sa_ctrl[0].f.spare[6] );
tran (\sa_ctrl[0][12] , \sa_ctrl[0].r.part0[12] );
tran (\sa_ctrl[0][12] , \sa_ctrl[0].f.spare[7] );
tran (\sa_ctrl[0][13] , \sa_ctrl[0].r.part0[13] );
tran (\sa_ctrl[0][13] , \sa_ctrl[0].f.spare[8] );
tran (\sa_ctrl[0][14] , \sa_ctrl[0].r.part0[14] );
tran (\sa_ctrl[0][14] , \sa_ctrl[0].f.spare[9] );
tran (\sa_ctrl[0][15] , \sa_ctrl[0].r.part0[15] );
tran (\sa_ctrl[0][15] , \sa_ctrl[0].f.spare[10] );
tran (\sa_ctrl[0][16] , \sa_ctrl[0].r.part0[16] );
tran (\sa_ctrl[0][16] , \sa_ctrl[0].f.spare[11] );
tran (\sa_ctrl[0][17] , \sa_ctrl[0].r.part0[17] );
tran (\sa_ctrl[0][17] , \sa_ctrl[0].f.spare[12] );
tran (\sa_ctrl[0][18] , \sa_ctrl[0].r.part0[18] );
tran (\sa_ctrl[0][18] , \sa_ctrl[0].f.spare[13] );
tran (\sa_ctrl[0][19] , \sa_ctrl[0].r.part0[19] );
tran (\sa_ctrl[0][19] , \sa_ctrl[0].f.spare[14] );
tran (\sa_ctrl[0][20] , \sa_ctrl[0].r.part0[20] );
tran (\sa_ctrl[0][20] , \sa_ctrl[0].f.spare[15] );
tran (\sa_ctrl[0][21] , \sa_ctrl[0].r.part0[21] );
tran (\sa_ctrl[0][21] , \sa_ctrl[0].f.spare[16] );
tran (\sa_ctrl[0][22] , \sa_ctrl[0].r.part0[22] );
tran (\sa_ctrl[0][22] , \sa_ctrl[0].f.spare[17] );
tran (\sa_ctrl[0][23] , \sa_ctrl[0].r.part0[23] );
tran (\sa_ctrl[0][23] , \sa_ctrl[0].f.spare[18] );
tran (\sa_ctrl[0][24] , \sa_ctrl[0].r.part0[24] );
tran (\sa_ctrl[0][24] , \sa_ctrl[0].f.spare[19] );
tran (\sa_ctrl[0][25] , \sa_ctrl[0].r.part0[25] );
tran (\sa_ctrl[0][25] , \sa_ctrl[0].f.spare[20] );
tran (\sa_ctrl[0][26] , \sa_ctrl[0].r.part0[26] );
tran (\sa_ctrl[0][26] , \sa_ctrl[0].f.spare[21] );
tran (\sa_ctrl[0][27] , \sa_ctrl[0].r.part0[27] );
tran (\sa_ctrl[0][27] , \sa_ctrl[0].f.spare[22] );
tran (\sa_ctrl[0][28] , \sa_ctrl[0].r.part0[28] );
tran (\sa_ctrl[0][28] , \sa_ctrl[0].f.spare[23] );
tran (\sa_ctrl[0][29] , \sa_ctrl[0].r.part0[29] );
tran (\sa_ctrl[0][29] , \sa_ctrl[0].f.spare[24] );
tran (\sa_ctrl[0][30] , \sa_ctrl[0].r.part0[30] );
tran (\sa_ctrl[0][30] , \sa_ctrl[0].f.spare[25] );
tran (\sa_ctrl[0][31] , \sa_ctrl[0].r.part0[31] );
tran (\sa_ctrl[0][31] , \sa_ctrl[0].f.spare[26] );
tran (\sa_ctrl[1][0] , \sa_ctrl[1].r.part0[0] );
tran (\sa_ctrl[1][0] , \sa_ctrl[1].f.sa_event_sel[0] );
tran (\sa_ctrl[1][1] , \sa_ctrl[1].r.part0[1] );
tran (\sa_ctrl[1][1] , \sa_ctrl[1].f.sa_event_sel[1] );
tran (\sa_ctrl[1][2] , \sa_ctrl[1].r.part0[2] );
tran (\sa_ctrl[1][2] , \sa_ctrl[1].f.sa_event_sel[2] );
tran (\sa_ctrl[1][3] , \sa_ctrl[1].r.part0[3] );
tran (\sa_ctrl[1][3] , \sa_ctrl[1].f.sa_event_sel[3] );
tran (\sa_ctrl[1][4] , \sa_ctrl[1].r.part0[4] );
tran (\sa_ctrl[1][4] , \sa_ctrl[1].f.sa_event_sel[4] );
tran (\sa_ctrl[1][5] , \sa_ctrl[1].r.part0[5] );
tran (\sa_ctrl[1][5] , \sa_ctrl[1].f.spare[0] );
tran (\sa_ctrl[1][6] , \sa_ctrl[1].r.part0[6] );
tran (\sa_ctrl[1][6] , \sa_ctrl[1].f.spare[1] );
tran (\sa_ctrl[1][7] , \sa_ctrl[1].r.part0[7] );
tran (\sa_ctrl[1][7] , \sa_ctrl[1].f.spare[2] );
tran (\sa_ctrl[1][8] , \sa_ctrl[1].r.part0[8] );
tran (\sa_ctrl[1][8] , \sa_ctrl[1].f.spare[3] );
tran (\sa_ctrl[1][9] , \sa_ctrl[1].r.part0[9] );
tran (\sa_ctrl[1][9] , \sa_ctrl[1].f.spare[4] );
tran (\sa_ctrl[1][10] , \sa_ctrl[1].r.part0[10] );
tran (\sa_ctrl[1][10] , \sa_ctrl[1].f.spare[5] );
tran (\sa_ctrl[1][11] , \sa_ctrl[1].r.part0[11] );
tran (\sa_ctrl[1][11] , \sa_ctrl[1].f.spare[6] );
tran (\sa_ctrl[1][12] , \sa_ctrl[1].r.part0[12] );
tran (\sa_ctrl[1][12] , \sa_ctrl[1].f.spare[7] );
tran (\sa_ctrl[1][13] , \sa_ctrl[1].r.part0[13] );
tran (\sa_ctrl[1][13] , \sa_ctrl[1].f.spare[8] );
tran (\sa_ctrl[1][14] , \sa_ctrl[1].r.part0[14] );
tran (\sa_ctrl[1][14] , \sa_ctrl[1].f.spare[9] );
tran (\sa_ctrl[1][15] , \sa_ctrl[1].r.part0[15] );
tran (\sa_ctrl[1][15] , \sa_ctrl[1].f.spare[10] );
tran (\sa_ctrl[1][16] , \sa_ctrl[1].r.part0[16] );
tran (\sa_ctrl[1][16] , \sa_ctrl[1].f.spare[11] );
tran (\sa_ctrl[1][17] , \sa_ctrl[1].r.part0[17] );
tran (\sa_ctrl[1][17] , \sa_ctrl[1].f.spare[12] );
tran (\sa_ctrl[1][18] , \sa_ctrl[1].r.part0[18] );
tran (\sa_ctrl[1][18] , \sa_ctrl[1].f.spare[13] );
tran (\sa_ctrl[1][19] , \sa_ctrl[1].r.part0[19] );
tran (\sa_ctrl[1][19] , \sa_ctrl[1].f.spare[14] );
tran (\sa_ctrl[1][20] , \sa_ctrl[1].r.part0[20] );
tran (\sa_ctrl[1][20] , \sa_ctrl[1].f.spare[15] );
tran (\sa_ctrl[1][21] , \sa_ctrl[1].r.part0[21] );
tran (\sa_ctrl[1][21] , \sa_ctrl[1].f.spare[16] );
tran (\sa_ctrl[1][22] , \sa_ctrl[1].r.part0[22] );
tran (\sa_ctrl[1][22] , \sa_ctrl[1].f.spare[17] );
tran (\sa_ctrl[1][23] , \sa_ctrl[1].r.part0[23] );
tran (\sa_ctrl[1][23] , \sa_ctrl[1].f.spare[18] );
tran (\sa_ctrl[1][24] , \sa_ctrl[1].r.part0[24] );
tran (\sa_ctrl[1][24] , \sa_ctrl[1].f.spare[19] );
tran (\sa_ctrl[1][25] , \sa_ctrl[1].r.part0[25] );
tran (\sa_ctrl[1][25] , \sa_ctrl[1].f.spare[20] );
tran (\sa_ctrl[1][26] , \sa_ctrl[1].r.part0[26] );
tran (\sa_ctrl[1][26] , \sa_ctrl[1].f.spare[21] );
tran (\sa_ctrl[1][27] , \sa_ctrl[1].r.part0[27] );
tran (\sa_ctrl[1][27] , \sa_ctrl[1].f.spare[22] );
tran (\sa_ctrl[1][28] , \sa_ctrl[1].r.part0[28] );
tran (\sa_ctrl[1][28] , \sa_ctrl[1].f.spare[23] );
tran (\sa_ctrl[1][29] , \sa_ctrl[1].r.part0[29] );
tran (\sa_ctrl[1][29] , \sa_ctrl[1].f.spare[24] );
tran (\sa_ctrl[1][30] , \sa_ctrl[1].r.part0[30] );
tran (\sa_ctrl[1][30] , \sa_ctrl[1].f.spare[25] );
tran (\sa_ctrl[1][31] , \sa_ctrl[1].r.part0[31] );
tran (\sa_ctrl[1][31] , \sa_ctrl[1].f.spare[26] );
tran (\sa_ctrl[2][0] , \sa_ctrl[2].r.part0[0] );
tran (\sa_ctrl[2][0] , \sa_ctrl[2].f.sa_event_sel[0] );
tran (\sa_ctrl[2][1] , \sa_ctrl[2].r.part0[1] );
tran (\sa_ctrl[2][1] , \sa_ctrl[2].f.sa_event_sel[1] );
tran (\sa_ctrl[2][2] , \sa_ctrl[2].r.part0[2] );
tran (\sa_ctrl[2][2] , \sa_ctrl[2].f.sa_event_sel[2] );
tran (\sa_ctrl[2][3] , \sa_ctrl[2].r.part0[3] );
tran (\sa_ctrl[2][3] , \sa_ctrl[2].f.sa_event_sel[3] );
tran (\sa_ctrl[2][4] , \sa_ctrl[2].r.part0[4] );
tran (\sa_ctrl[2][4] , \sa_ctrl[2].f.sa_event_sel[4] );
tran (\sa_ctrl[2][5] , \sa_ctrl[2].r.part0[5] );
tran (\sa_ctrl[2][5] , \sa_ctrl[2].f.spare[0] );
tran (\sa_ctrl[2][6] , \sa_ctrl[2].r.part0[6] );
tran (\sa_ctrl[2][6] , \sa_ctrl[2].f.spare[1] );
tran (\sa_ctrl[2][7] , \sa_ctrl[2].r.part0[7] );
tran (\sa_ctrl[2][7] , \sa_ctrl[2].f.spare[2] );
tran (\sa_ctrl[2][8] , \sa_ctrl[2].r.part0[8] );
tran (\sa_ctrl[2][8] , \sa_ctrl[2].f.spare[3] );
tran (\sa_ctrl[2][9] , \sa_ctrl[2].r.part0[9] );
tran (\sa_ctrl[2][9] , \sa_ctrl[2].f.spare[4] );
tran (\sa_ctrl[2][10] , \sa_ctrl[2].r.part0[10] );
tran (\sa_ctrl[2][10] , \sa_ctrl[2].f.spare[5] );
tran (\sa_ctrl[2][11] , \sa_ctrl[2].r.part0[11] );
tran (\sa_ctrl[2][11] , \sa_ctrl[2].f.spare[6] );
tran (\sa_ctrl[2][12] , \sa_ctrl[2].r.part0[12] );
tran (\sa_ctrl[2][12] , \sa_ctrl[2].f.spare[7] );
tran (\sa_ctrl[2][13] , \sa_ctrl[2].r.part0[13] );
tran (\sa_ctrl[2][13] , \sa_ctrl[2].f.spare[8] );
tran (\sa_ctrl[2][14] , \sa_ctrl[2].r.part0[14] );
tran (\sa_ctrl[2][14] , \sa_ctrl[2].f.spare[9] );
tran (\sa_ctrl[2][15] , \sa_ctrl[2].r.part0[15] );
tran (\sa_ctrl[2][15] , \sa_ctrl[2].f.spare[10] );
tran (\sa_ctrl[2][16] , \sa_ctrl[2].r.part0[16] );
tran (\sa_ctrl[2][16] , \sa_ctrl[2].f.spare[11] );
tran (\sa_ctrl[2][17] , \sa_ctrl[2].r.part0[17] );
tran (\sa_ctrl[2][17] , \sa_ctrl[2].f.spare[12] );
tran (\sa_ctrl[2][18] , \sa_ctrl[2].r.part0[18] );
tran (\sa_ctrl[2][18] , \sa_ctrl[2].f.spare[13] );
tran (\sa_ctrl[2][19] , \sa_ctrl[2].r.part0[19] );
tran (\sa_ctrl[2][19] , \sa_ctrl[2].f.spare[14] );
tran (\sa_ctrl[2][20] , \sa_ctrl[2].r.part0[20] );
tran (\sa_ctrl[2][20] , \sa_ctrl[2].f.spare[15] );
tran (\sa_ctrl[2][21] , \sa_ctrl[2].r.part0[21] );
tran (\sa_ctrl[2][21] , \sa_ctrl[2].f.spare[16] );
tran (\sa_ctrl[2][22] , \sa_ctrl[2].r.part0[22] );
tran (\sa_ctrl[2][22] , \sa_ctrl[2].f.spare[17] );
tran (\sa_ctrl[2][23] , \sa_ctrl[2].r.part0[23] );
tran (\sa_ctrl[2][23] , \sa_ctrl[2].f.spare[18] );
tran (\sa_ctrl[2][24] , \sa_ctrl[2].r.part0[24] );
tran (\sa_ctrl[2][24] , \sa_ctrl[2].f.spare[19] );
tran (\sa_ctrl[2][25] , \sa_ctrl[2].r.part0[25] );
tran (\sa_ctrl[2][25] , \sa_ctrl[2].f.spare[20] );
tran (\sa_ctrl[2][26] , \sa_ctrl[2].r.part0[26] );
tran (\sa_ctrl[2][26] , \sa_ctrl[2].f.spare[21] );
tran (\sa_ctrl[2][27] , \sa_ctrl[2].r.part0[27] );
tran (\sa_ctrl[2][27] , \sa_ctrl[2].f.spare[22] );
tran (\sa_ctrl[2][28] , \sa_ctrl[2].r.part0[28] );
tran (\sa_ctrl[2][28] , \sa_ctrl[2].f.spare[23] );
tran (\sa_ctrl[2][29] , \sa_ctrl[2].r.part0[29] );
tran (\sa_ctrl[2][29] , \sa_ctrl[2].f.spare[24] );
tran (\sa_ctrl[2][30] , \sa_ctrl[2].r.part0[30] );
tran (\sa_ctrl[2][30] , \sa_ctrl[2].f.spare[25] );
tran (\sa_ctrl[2][31] , \sa_ctrl[2].r.part0[31] );
tran (\sa_ctrl[2][31] , \sa_ctrl[2].f.spare[26] );
tran (\sa_ctrl[3][0] , \sa_ctrl[3].r.part0[0] );
tran (\sa_ctrl[3][0] , \sa_ctrl[3].f.sa_event_sel[0] );
tran (\sa_ctrl[3][1] , \sa_ctrl[3].r.part0[1] );
tran (\sa_ctrl[3][1] , \sa_ctrl[3].f.sa_event_sel[1] );
tran (\sa_ctrl[3][2] , \sa_ctrl[3].r.part0[2] );
tran (\sa_ctrl[3][2] , \sa_ctrl[3].f.sa_event_sel[2] );
tran (\sa_ctrl[3][3] , \sa_ctrl[3].r.part0[3] );
tran (\sa_ctrl[3][3] , \sa_ctrl[3].f.sa_event_sel[3] );
tran (\sa_ctrl[3][4] , \sa_ctrl[3].r.part0[4] );
tran (\sa_ctrl[3][4] , \sa_ctrl[3].f.sa_event_sel[4] );
tran (\sa_ctrl[3][5] , \sa_ctrl[3].r.part0[5] );
tran (\sa_ctrl[3][5] , \sa_ctrl[3].f.spare[0] );
tran (\sa_ctrl[3][6] , \sa_ctrl[3].r.part0[6] );
tran (\sa_ctrl[3][6] , \sa_ctrl[3].f.spare[1] );
tran (\sa_ctrl[3][7] , \sa_ctrl[3].r.part0[7] );
tran (\sa_ctrl[3][7] , \sa_ctrl[3].f.spare[2] );
tran (\sa_ctrl[3][8] , \sa_ctrl[3].r.part0[8] );
tran (\sa_ctrl[3][8] , \sa_ctrl[3].f.spare[3] );
tran (\sa_ctrl[3][9] , \sa_ctrl[3].r.part0[9] );
tran (\sa_ctrl[3][9] , \sa_ctrl[3].f.spare[4] );
tran (\sa_ctrl[3][10] , \sa_ctrl[3].r.part0[10] );
tran (\sa_ctrl[3][10] , \sa_ctrl[3].f.spare[5] );
tran (\sa_ctrl[3][11] , \sa_ctrl[3].r.part0[11] );
tran (\sa_ctrl[3][11] , \sa_ctrl[3].f.spare[6] );
tran (\sa_ctrl[3][12] , \sa_ctrl[3].r.part0[12] );
tran (\sa_ctrl[3][12] , \sa_ctrl[3].f.spare[7] );
tran (\sa_ctrl[3][13] , \sa_ctrl[3].r.part0[13] );
tran (\sa_ctrl[3][13] , \sa_ctrl[3].f.spare[8] );
tran (\sa_ctrl[3][14] , \sa_ctrl[3].r.part0[14] );
tran (\sa_ctrl[3][14] , \sa_ctrl[3].f.spare[9] );
tran (\sa_ctrl[3][15] , \sa_ctrl[3].r.part0[15] );
tran (\sa_ctrl[3][15] , \sa_ctrl[3].f.spare[10] );
tran (\sa_ctrl[3][16] , \sa_ctrl[3].r.part0[16] );
tran (\sa_ctrl[3][16] , \sa_ctrl[3].f.spare[11] );
tran (\sa_ctrl[3][17] , \sa_ctrl[3].r.part0[17] );
tran (\sa_ctrl[3][17] , \sa_ctrl[3].f.spare[12] );
tran (\sa_ctrl[3][18] , \sa_ctrl[3].r.part0[18] );
tran (\sa_ctrl[3][18] , \sa_ctrl[3].f.spare[13] );
tran (\sa_ctrl[3][19] , \sa_ctrl[3].r.part0[19] );
tran (\sa_ctrl[3][19] , \sa_ctrl[3].f.spare[14] );
tran (\sa_ctrl[3][20] , \sa_ctrl[3].r.part0[20] );
tran (\sa_ctrl[3][20] , \sa_ctrl[3].f.spare[15] );
tran (\sa_ctrl[3][21] , \sa_ctrl[3].r.part0[21] );
tran (\sa_ctrl[3][21] , \sa_ctrl[3].f.spare[16] );
tran (\sa_ctrl[3][22] , \sa_ctrl[3].r.part0[22] );
tran (\sa_ctrl[3][22] , \sa_ctrl[3].f.spare[17] );
tran (\sa_ctrl[3][23] , \sa_ctrl[3].r.part0[23] );
tran (\sa_ctrl[3][23] , \sa_ctrl[3].f.spare[18] );
tran (\sa_ctrl[3][24] , \sa_ctrl[3].r.part0[24] );
tran (\sa_ctrl[3][24] , \sa_ctrl[3].f.spare[19] );
tran (\sa_ctrl[3][25] , \sa_ctrl[3].r.part0[25] );
tran (\sa_ctrl[3][25] , \sa_ctrl[3].f.spare[20] );
tran (\sa_ctrl[3][26] , \sa_ctrl[3].r.part0[26] );
tran (\sa_ctrl[3][26] , \sa_ctrl[3].f.spare[21] );
tran (\sa_ctrl[3][27] , \sa_ctrl[3].r.part0[27] );
tran (\sa_ctrl[3][27] , \sa_ctrl[3].f.spare[22] );
tran (\sa_ctrl[3][28] , \sa_ctrl[3].r.part0[28] );
tran (\sa_ctrl[3][28] , \sa_ctrl[3].f.spare[23] );
tran (\sa_ctrl[3][29] , \sa_ctrl[3].r.part0[29] );
tran (\sa_ctrl[3][29] , \sa_ctrl[3].f.spare[24] );
tran (\sa_ctrl[3][30] , \sa_ctrl[3].r.part0[30] );
tran (\sa_ctrl[3][30] , \sa_ctrl[3].f.spare[25] );
tran (\sa_ctrl[3][31] , \sa_ctrl[3].r.part0[31] );
tran (\sa_ctrl[3][31] , \sa_ctrl[3].f.spare[26] );
tran (\sa_ctrl[4][0] , \sa_ctrl[4].r.part0[0] );
tran (\sa_ctrl[4][0] , \sa_ctrl[4].f.sa_event_sel[0] );
tran (\sa_ctrl[4][1] , \sa_ctrl[4].r.part0[1] );
tran (\sa_ctrl[4][1] , \sa_ctrl[4].f.sa_event_sel[1] );
tran (\sa_ctrl[4][2] , \sa_ctrl[4].r.part0[2] );
tran (\sa_ctrl[4][2] , \sa_ctrl[4].f.sa_event_sel[2] );
tran (\sa_ctrl[4][3] , \sa_ctrl[4].r.part0[3] );
tran (\sa_ctrl[4][3] , \sa_ctrl[4].f.sa_event_sel[3] );
tran (\sa_ctrl[4][4] , \sa_ctrl[4].r.part0[4] );
tran (\sa_ctrl[4][4] , \sa_ctrl[4].f.sa_event_sel[4] );
tran (\sa_ctrl[4][5] , \sa_ctrl[4].r.part0[5] );
tran (\sa_ctrl[4][5] , \sa_ctrl[4].f.spare[0] );
tran (\sa_ctrl[4][6] , \sa_ctrl[4].r.part0[6] );
tran (\sa_ctrl[4][6] , \sa_ctrl[4].f.spare[1] );
tran (\sa_ctrl[4][7] , \sa_ctrl[4].r.part0[7] );
tran (\sa_ctrl[4][7] , \sa_ctrl[4].f.spare[2] );
tran (\sa_ctrl[4][8] , \sa_ctrl[4].r.part0[8] );
tran (\sa_ctrl[4][8] , \sa_ctrl[4].f.spare[3] );
tran (\sa_ctrl[4][9] , \sa_ctrl[4].r.part0[9] );
tran (\sa_ctrl[4][9] , \sa_ctrl[4].f.spare[4] );
tran (\sa_ctrl[4][10] , \sa_ctrl[4].r.part0[10] );
tran (\sa_ctrl[4][10] , \sa_ctrl[4].f.spare[5] );
tran (\sa_ctrl[4][11] , \sa_ctrl[4].r.part0[11] );
tran (\sa_ctrl[4][11] , \sa_ctrl[4].f.spare[6] );
tran (\sa_ctrl[4][12] , \sa_ctrl[4].r.part0[12] );
tran (\sa_ctrl[4][12] , \sa_ctrl[4].f.spare[7] );
tran (\sa_ctrl[4][13] , \sa_ctrl[4].r.part0[13] );
tran (\sa_ctrl[4][13] , \sa_ctrl[4].f.spare[8] );
tran (\sa_ctrl[4][14] , \sa_ctrl[4].r.part0[14] );
tran (\sa_ctrl[4][14] , \sa_ctrl[4].f.spare[9] );
tran (\sa_ctrl[4][15] , \sa_ctrl[4].r.part0[15] );
tran (\sa_ctrl[4][15] , \sa_ctrl[4].f.spare[10] );
tran (\sa_ctrl[4][16] , \sa_ctrl[4].r.part0[16] );
tran (\sa_ctrl[4][16] , \sa_ctrl[4].f.spare[11] );
tran (\sa_ctrl[4][17] , \sa_ctrl[4].r.part0[17] );
tran (\sa_ctrl[4][17] , \sa_ctrl[4].f.spare[12] );
tran (\sa_ctrl[4][18] , \sa_ctrl[4].r.part0[18] );
tran (\sa_ctrl[4][18] , \sa_ctrl[4].f.spare[13] );
tran (\sa_ctrl[4][19] , \sa_ctrl[4].r.part0[19] );
tran (\sa_ctrl[4][19] , \sa_ctrl[4].f.spare[14] );
tran (\sa_ctrl[4][20] , \sa_ctrl[4].r.part0[20] );
tran (\sa_ctrl[4][20] , \sa_ctrl[4].f.spare[15] );
tran (\sa_ctrl[4][21] , \sa_ctrl[4].r.part0[21] );
tran (\sa_ctrl[4][21] , \sa_ctrl[4].f.spare[16] );
tran (\sa_ctrl[4][22] , \sa_ctrl[4].r.part0[22] );
tran (\sa_ctrl[4][22] , \sa_ctrl[4].f.spare[17] );
tran (\sa_ctrl[4][23] , \sa_ctrl[4].r.part0[23] );
tran (\sa_ctrl[4][23] , \sa_ctrl[4].f.spare[18] );
tran (\sa_ctrl[4][24] , \sa_ctrl[4].r.part0[24] );
tran (\sa_ctrl[4][24] , \sa_ctrl[4].f.spare[19] );
tran (\sa_ctrl[4][25] , \sa_ctrl[4].r.part0[25] );
tran (\sa_ctrl[4][25] , \sa_ctrl[4].f.spare[20] );
tran (\sa_ctrl[4][26] , \sa_ctrl[4].r.part0[26] );
tran (\sa_ctrl[4][26] , \sa_ctrl[4].f.spare[21] );
tran (\sa_ctrl[4][27] , \sa_ctrl[4].r.part0[27] );
tran (\sa_ctrl[4][27] , \sa_ctrl[4].f.spare[22] );
tran (\sa_ctrl[4][28] , \sa_ctrl[4].r.part0[28] );
tran (\sa_ctrl[4][28] , \sa_ctrl[4].f.spare[23] );
tran (\sa_ctrl[4][29] , \sa_ctrl[4].r.part0[29] );
tran (\sa_ctrl[4][29] , \sa_ctrl[4].f.spare[24] );
tran (\sa_ctrl[4][30] , \sa_ctrl[4].r.part0[30] );
tran (\sa_ctrl[4][30] , \sa_ctrl[4].f.spare[25] );
tran (\sa_ctrl[4][31] , \sa_ctrl[4].r.part0[31] );
tran (\sa_ctrl[4][31] , \sa_ctrl[4].f.spare[26] );
tran (\sa_ctrl[5][0] , \sa_ctrl[5].r.part0[0] );
tran (\sa_ctrl[5][0] , \sa_ctrl[5].f.sa_event_sel[0] );
tran (\sa_ctrl[5][1] , \sa_ctrl[5].r.part0[1] );
tran (\sa_ctrl[5][1] , \sa_ctrl[5].f.sa_event_sel[1] );
tran (\sa_ctrl[5][2] , \sa_ctrl[5].r.part0[2] );
tran (\sa_ctrl[5][2] , \sa_ctrl[5].f.sa_event_sel[2] );
tran (\sa_ctrl[5][3] , \sa_ctrl[5].r.part0[3] );
tran (\sa_ctrl[5][3] , \sa_ctrl[5].f.sa_event_sel[3] );
tran (\sa_ctrl[5][4] , \sa_ctrl[5].r.part0[4] );
tran (\sa_ctrl[5][4] , \sa_ctrl[5].f.sa_event_sel[4] );
tran (\sa_ctrl[5][5] , \sa_ctrl[5].r.part0[5] );
tran (\sa_ctrl[5][5] , \sa_ctrl[5].f.spare[0] );
tran (\sa_ctrl[5][6] , \sa_ctrl[5].r.part0[6] );
tran (\sa_ctrl[5][6] , \sa_ctrl[5].f.spare[1] );
tran (\sa_ctrl[5][7] , \sa_ctrl[5].r.part0[7] );
tran (\sa_ctrl[5][7] , \sa_ctrl[5].f.spare[2] );
tran (\sa_ctrl[5][8] , \sa_ctrl[5].r.part0[8] );
tran (\sa_ctrl[5][8] , \sa_ctrl[5].f.spare[3] );
tran (\sa_ctrl[5][9] , \sa_ctrl[5].r.part0[9] );
tran (\sa_ctrl[5][9] , \sa_ctrl[5].f.spare[4] );
tran (\sa_ctrl[5][10] , \sa_ctrl[5].r.part0[10] );
tran (\sa_ctrl[5][10] , \sa_ctrl[5].f.spare[5] );
tran (\sa_ctrl[5][11] , \sa_ctrl[5].r.part0[11] );
tran (\sa_ctrl[5][11] , \sa_ctrl[5].f.spare[6] );
tran (\sa_ctrl[5][12] , \sa_ctrl[5].r.part0[12] );
tran (\sa_ctrl[5][12] , \sa_ctrl[5].f.spare[7] );
tran (\sa_ctrl[5][13] , \sa_ctrl[5].r.part0[13] );
tran (\sa_ctrl[5][13] , \sa_ctrl[5].f.spare[8] );
tran (\sa_ctrl[5][14] , \sa_ctrl[5].r.part0[14] );
tran (\sa_ctrl[5][14] , \sa_ctrl[5].f.spare[9] );
tran (\sa_ctrl[5][15] , \sa_ctrl[5].r.part0[15] );
tran (\sa_ctrl[5][15] , \sa_ctrl[5].f.spare[10] );
tran (\sa_ctrl[5][16] , \sa_ctrl[5].r.part0[16] );
tran (\sa_ctrl[5][16] , \sa_ctrl[5].f.spare[11] );
tran (\sa_ctrl[5][17] , \sa_ctrl[5].r.part0[17] );
tran (\sa_ctrl[5][17] , \sa_ctrl[5].f.spare[12] );
tran (\sa_ctrl[5][18] , \sa_ctrl[5].r.part0[18] );
tran (\sa_ctrl[5][18] , \sa_ctrl[5].f.spare[13] );
tran (\sa_ctrl[5][19] , \sa_ctrl[5].r.part0[19] );
tran (\sa_ctrl[5][19] , \sa_ctrl[5].f.spare[14] );
tran (\sa_ctrl[5][20] , \sa_ctrl[5].r.part0[20] );
tran (\sa_ctrl[5][20] , \sa_ctrl[5].f.spare[15] );
tran (\sa_ctrl[5][21] , \sa_ctrl[5].r.part0[21] );
tran (\sa_ctrl[5][21] , \sa_ctrl[5].f.spare[16] );
tran (\sa_ctrl[5][22] , \sa_ctrl[5].r.part0[22] );
tran (\sa_ctrl[5][22] , \sa_ctrl[5].f.spare[17] );
tran (\sa_ctrl[5][23] , \sa_ctrl[5].r.part0[23] );
tran (\sa_ctrl[5][23] , \sa_ctrl[5].f.spare[18] );
tran (\sa_ctrl[5][24] , \sa_ctrl[5].r.part0[24] );
tran (\sa_ctrl[5][24] , \sa_ctrl[5].f.spare[19] );
tran (\sa_ctrl[5][25] , \sa_ctrl[5].r.part0[25] );
tran (\sa_ctrl[5][25] , \sa_ctrl[5].f.spare[20] );
tran (\sa_ctrl[5][26] , \sa_ctrl[5].r.part0[26] );
tran (\sa_ctrl[5][26] , \sa_ctrl[5].f.spare[21] );
tran (\sa_ctrl[5][27] , \sa_ctrl[5].r.part0[27] );
tran (\sa_ctrl[5][27] , \sa_ctrl[5].f.spare[22] );
tran (\sa_ctrl[5][28] , \sa_ctrl[5].r.part0[28] );
tran (\sa_ctrl[5][28] , \sa_ctrl[5].f.spare[23] );
tran (\sa_ctrl[5][29] , \sa_ctrl[5].r.part0[29] );
tran (\sa_ctrl[5][29] , \sa_ctrl[5].f.spare[24] );
tran (\sa_ctrl[5][30] , \sa_ctrl[5].r.part0[30] );
tran (\sa_ctrl[5][30] , \sa_ctrl[5].f.spare[25] );
tran (\sa_ctrl[5][31] , \sa_ctrl[5].r.part0[31] );
tran (\sa_ctrl[5][31] , \sa_ctrl[5].f.spare[26] );
tran (\sa_ctrl[6][0] , \sa_ctrl[6].r.part0[0] );
tran (\sa_ctrl[6][0] , \sa_ctrl[6].f.sa_event_sel[0] );
tran (\sa_ctrl[6][1] , \sa_ctrl[6].r.part0[1] );
tran (\sa_ctrl[6][1] , \sa_ctrl[6].f.sa_event_sel[1] );
tran (\sa_ctrl[6][2] , \sa_ctrl[6].r.part0[2] );
tran (\sa_ctrl[6][2] , \sa_ctrl[6].f.sa_event_sel[2] );
tran (\sa_ctrl[6][3] , \sa_ctrl[6].r.part0[3] );
tran (\sa_ctrl[6][3] , \sa_ctrl[6].f.sa_event_sel[3] );
tran (\sa_ctrl[6][4] , \sa_ctrl[6].r.part0[4] );
tran (\sa_ctrl[6][4] , \sa_ctrl[6].f.sa_event_sel[4] );
tran (\sa_ctrl[6][5] , \sa_ctrl[6].r.part0[5] );
tran (\sa_ctrl[6][5] , \sa_ctrl[6].f.spare[0] );
tran (\sa_ctrl[6][6] , \sa_ctrl[6].r.part0[6] );
tran (\sa_ctrl[6][6] , \sa_ctrl[6].f.spare[1] );
tran (\sa_ctrl[6][7] , \sa_ctrl[6].r.part0[7] );
tran (\sa_ctrl[6][7] , \sa_ctrl[6].f.spare[2] );
tran (\sa_ctrl[6][8] , \sa_ctrl[6].r.part0[8] );
tran (\sa_ctrl[6][8] , \sa_ctrl[6].f.spare[3] );
tran (\sa_ctrl[6][9] , \sa_ctrl[6].r.part0[9] );
tran (\sa_ctrl[6][9] , \sa_ctrl[6].f.spare[4] );
tran (\sa_ctrl[6][10] , \sa_ctrl[6].r.part0[10] );
tran (\sa_ctrl[6][10] , \sa_ctrl[6].f.spare[5] );
tran (\sa_ctrl[6][11] , \sa_ctrl[6].r.part0[11] );
tran (\sa_ctrl[6][11] , \sa_ctrl[6].f.spare[6] );
tran (\sa_ctrl[6][12] , \sa_ctrl[6].r.part0[12] );
tran (\sa_ctrl[6][12] , \sa_ctrl[6].f.spare[7] );
tran (\sa_ctrl[6][13] , \sa_ctrl[6].r.part0[13] );
tran (\sa_ctrl[6][13] , \sa_ctrl[6].f.spare[8] );
tran (\sa_ctrl[6][14] , \sa_ctrl[6].r.part0[14] );
tran (\sa_ctrl[6][14] , \sa_ctrl[6].f.spare[9] );
tran (\sa_ctrl[6][15] , \sa_ctrl[6].r.part0[15] );
tran (\sa_ctrl[6][15] , \sa_ctrl[6].f.spare[10] );
tran (\sa_ctrl[6][16] , \sa_ctrl[6].r.part0[16] );
tran (\sa_ctrl[6][16] , \sa_ctrl[6].f.spare[11] );
tran (\sa_ctrl[6][17] , \sa_ctrl[6].r.part0[17] );
tran (\sa_ctrl[6][17] , \sa_ctrl[6].f.spare[12] );
tran (\sa_ctrl[6][18] , \sa_ctrl[6].r.part0[18] );
tran (\sa_ctrl[6][18] , \sa_ctrl[6].f.spare[13] );
tran (\sa_ctrl[6][19] , \sa_ctrl[6].r.part0[19] );
tran (\sa_ctrl[6][19] , \sa_ctrl[6].f.spare[14] );
tran (\sa_ctrl[6][20] , \sa_ctrl[6].r.part0[20] );
tran (\sa_ctrl[6][20] , \sa_ctrl[6].f.spare[15] );
tran (\sa_ctrl[6][21] , \sa_ctrl[6].r.part0[21] );
tran (\sa_ctrl[6][21] , \sa_ctrl[6].f.spare[16] );
tran (\sa_ctrl[6][22] , \sa_ctrl[6].r.part0[22] );
tran (\sa_ctrl[6][22] , \sa_ctrl[6].f.spare[17] );
tran (\sa_ctrl[6][23] , \sa_ctrl[6].r.part0[23] );
tran (\sa_ctrl[6][23] , \sa_ctrl[6].f.spare[18] );
tran (\sa_ctrl[6][24] , \sa_ctrl[6].r.part0[24] );
tran (\sa_ctrl[6][24] , \sa_ctrl[6].f.spare[19] );
tran (\sa_ctrl[6][25] , \sa_ctrl[6].r.part0[25] );
tran (\sa_ctrl[6][25] , \sa_ctrl[6].f.spare[20] );
tran (\sa_ctrl[6][26] , \sa_ctrl[6].r.part0[26] );
tran (\sa_ctrl[6][26] , \sa_ctrl[6].f.spare[21] );
tran (\sa_ctrl[6][27] , \sa_ctrl[6].r.part0[27] );
tran (\sa_ctrl[6][27] , \sa_ctrl[6].f.spare[22] );
tran (\sa_ctrl[6][28] , \sa_ctrl[6].r.part0[28] );
tran (\sa_ctrl[6][28] , \sa_ctrl[6].f.spare[23] );
tran (\sa_ctrl[6][29] , \sa_ctrl[6].r.part0[29] );
tran (\sa_ctrl[6][29] , \sa_ctrl[6].f.spare[24] );
tran (\sa_ctrl[6][30] , \sa_ctrl[6].r.part0[30] );
tran (\sa_ctrl[6][30] , \sa_ctrl[6].f.spare[25] );
tran (\sa_ctrl[6][31] , \sa_ctrl[6].r.part0[31] );
tran (\sa_ctrl[6][31] , \sa_ctrl[6].f.spare[26] );
tran (\sa_ctrl[7][0] , \sa_ctrl[7].r.part0[0] );
tran (\sa_ctrl[7][0] , \sa_ctrl[7].f.sa_event_sel[0] );
tran (\sa_ctrl[7][1] , \sa_ctrl[7].r.part0[1] );
tran (\sa_ctrl[7][1] , \sa_ctrl[7].f.sa_event_sel[1] );
tran (\sa_ctrl[7][2] , \sa_ctrl[7].r.part0[2] );
tran (\sa_ctrl[7][2] , \sa_ctrl[7].f.sa_event_sel[2] );
tran (\sa_ctrl[7][3] , \sa_ctrl[7].r.part0[3] );
tran (\sa_ctrl[7][3] , \sa_ctrl[7].f.sa_event_sel[3] );
tran (\sa_ctrl[7][4] , \sa_ctrl[7].r.part0[4] );
tran (\sa_ctrl[7][4] , \sa_ctrl[7].f.sa_event_sel[4] );
tran (\sa_ctrl[7][5] , \sa_ctrl[7].r.part0[5] );
tran (\sa_ctrl[7][5] , \sa_ctrl[7].f.spare[0] );
tran (\sa_ctrl[7][6] , \sa_ctrl[7].r.part0[6] );
tran (\sa_ctrl[7][6] , \sa_ctrl[7].f.spare[1] );
tran (\sa_ctrl[7][7] , \sa_ctrl[7].r.part0[7] );
tran (\sa_ctrl[7][7] , \sa_ctrl[7].f.spare[2] );
tran (\sa_ctrl[7][8] , \sa_ctrl[7].r.part0[8] );
tran (\sa_ctrl[7][8] , \sa_ctrl[7].f.spare[3] );
tran (\sa_ctrl[7][9] , \sa_ctrl[7].r.part0[9] );
tran (\sa_ctrl[7][9] , \sa_ctrl[7].f.spare[4] );
tran (\sa_ctrl[7][10] , \sa_ctrl[7].r.part0[10] );
tran (\sa_ctrl[7][10] , \sa_ctrl[7].f.spare[5] );
tran (\sa_ctrl[7][11] , \sa_ctrl[7].r.part0[11] );
tran (\sa_ctrl[7][11] , \sa_ctrl[7].f.spare[6] );
tran (\sa_ctrl[7][12] , \sa_ctrl[7].r.part0[12] );
tran (\sa_ctrl[7][12] , \sa_ctrl[7].f.spare[7] );
tran (\sa_ctrl[7][13] , \sa_ctrl[7].r.part0[13] );
tran (\sa_ctrl[7][13] , \sa_ctrl[7].f.spare[8] );
tran (\sa_ctrl[7][14] , \sa_ctrl[7].r.part0[14] );
tran (\sa_ctrl[7][14] , \sa_ctrl[7].f.spare[9] );
tran (\sa_ctrl[7][15] , \sa_ctrl[7].r.part0[15] );
tran (\sa_ctrl[7][15] , \sa_ctrl[7].f.spare[10] );
tran (\sa_ctrl[7][16] , \sa_ctrl[7].r.part0[16] );
tran (\sa_ctrl[7][16] , \sa_ctrl[7].f.spare[11] );
tran (\sa_ctrl[7][17] , \sa_ctrl[7].r.part0[17] );
tran (\sa_ctrl[7][17] , \sa_ctrl[7].f.spare[12] );
tran (\sa_ctrl[7][18] , \sa_ctrl[7].r.part0[18] );
tran (\sa_ctrl[7][18] , \sa_ctrl[7].f.spare[13] );
tran (\sa_ctrl[7][19] , \sa_ctrl[7].r.part0[19] );
tran (\sa_ctrl[7][19] , \sa_ctrl[7].f.spare[14] );
tran (\sa_ctrl[7][20] , \sa_ctrl[7].r.part0[20] );
tran (\sa_ctrl[7][20] , \sa_ctrl[7].f.spare[15] );
tran (\sa_ctrl[7][21] , \sa_ctrl[7].r.part0[21] );
tran (\sa_ctrl[7][21] , \sa_ctrl[7].f.spare[16] );
tran (\sa_ctrl[7][22] , \sa_ctrl[7].r.part0[22] );
tran (\sa_ctrl[7][22] , \sa_ctrl[7].f.spare[17] );
tran (\sa_ctrl[7][23] , \sa_ctrl[7].r.part0[23] );
tran (\sa_ctrl[7][23] , \sa_ctrl[7].f.spare[18] );
tran (\sa_ctrl[7][24] , \sa_ctrl[7].r.part0[24] );
tran (\sa_ctrl[7][24] , \sa_ctrl[7].f.spare[19] );
tran (\sa_ctrl[7][25] , \sa_ctrl[7].r.part0[25] );
tran (\sa_ctrl[7][25] , \sa_ctrl[7].f.spare[20] );
tran (\sa_ctrl[7][26] , \sa_ctrl[7].r.part0[26] );
tran (\sa_ctrl[7][26] , \sa_ctrl[7].f.spare[21] );
tran (\sa_ctrl[7][27] , \sa_ctrl[7].r.part0[27] );
tran (\sa_ctrl[7][27] , \sa_ctrl[7].f.spare[22] );
tran (\sa_ctrl[7][28] , \sa_ctrl[7].r.part0[28] );
tran (\sa_ctrl[7][28] , \sa_ctrl[7].f.spare[23] );
tran (\sa_ctrl[7][29] , \sa_ctrl[7].r.part0[29] );
tran (\sa_ctrl[7][29] , \sa_ctrl[7].f.spare[24] );
tran (\sa_ctrl[7][30] , \sa_ctrl[7].r.part0[30] );
tran (\sa_ctrl[7][30] , \sa_ctrl[7].f.spare[25] );
tran (\sa_ctrl[7][31] , \sa_ctrl[7].r.part0[31] );
tran (\sa_ctrl[7][31] , \sa_ctrl[7].f.spare[26] );
tran (\sa_ctrl[8][0] , \sa_ctrl[8].r.part0[0] );
tran (\sa_ctrl[8][0] , \sa_ctrl[8].f.sa_event_sel[0] );
tran (\sa_ctrl[8][1] , \sa_ctrl[8].r.part0[1] );
tran (\sa_ctrl[8][1] , \sa_ctrl[8].f.sa_event_sel[1] );
tran (\sa_ctrl[8][2] , \sa_ctrl[8].r.part0[2] );
tran (\sa_ctrl[8][2] , \sa_ctrl[8].f.sa_event_sel[2] );
tran (\sa_ctrl[8][3] , \sa_ctrl[8].r.part0[3] );
tran (\sa_ctrl[8][3] , \sa_ctrl[8].f.sa_event_sel[3] );
tran (\sa_ctrl[8][4] , \sa_ctrl[8].r.part0[4] );
tran (\sa_ctrl[8][4] , \sa_ctrl[8].f.sa_event_sel[4] );
tran (\sa_ctrl[8][5] , \sa_ctrl[8].r.part0[5] );
tran (\sa_ctrl[8][5] , \sa_ctrl[8].f.spare[0] );
tran (\sa_ctrl[8][6] , \sa_ctrl[8].r.part0[6] );
tran (\sa_ctrl[8][6] , \sa_ctrl[8].f.spare[1] );
tran (\sa_ctrl[8][7] , \sa_ctrl[8].r.part0[7] );
tran (\sa_ctrl[8][7] , \sa_ctrl[8].f.spare[2] );
tran (\sa_ctrl[8][8] , \sa_ctrl[8].r.part0[8] );
tran (\sa_ctrl[8][8] , \sa_ctrl[8].f.spare[3] );
tran (\sa_ctrl[8][9] , \sa_ctrl[8].r.part0[9] );
tran (\sa_ctrl[8][9] , \sa_ctrl[8].f.spare[4] );
tran (\sa_ctrl[8][10] , \sa_ctrl[8].r.part0[10] );
tran (\sa_ctrl[8][10] , \sa_ctrl[8].f.spare[5] );
tran (\sa_ctrl[8][11] , \sa_ctrl[8].r.part0[11] );
tran (\sa_ctrl[8][11] , \sa_ctrl[8].f.spare[6] );
tran (\sa_ctrl[8][12] , \sa_ctrl[8].r.part0[12] );
tran (\sa_ctrl[8][12] , \sa_ctrl[8].f.spare[7] );
tran (\sa_ctrl[8][13] , \sa_ctrl[8].r.part0[13] );
tran (\sa_ctrl[8][13] , \sa_ctrl[8].f.spare[8] );
tran (\sa_ctrl[8][14] , \sa_ctrl[8].r.part0[14] );
tran (\sa_ctrl[8][14] , \sa_ctrl[8].f.spare[9] );
tran (\sa_ctrl[8][15] , \sa_ctrl[8].r.part0[15] );
tran (\sa_ctrl[8][15] , \sa_ctrl[8].f.spare[10] );
tran (\sa_ctrl[8][16] , \sa_ctrl[8].r.part0[16] );
tran (\sa_ctrl[8][16] , \sa_ctrl[8].f.spare[11] );
tran (\sa_ctrl[8][17] , \sa_ctrl[8].r.part0[17] );
tran (\sa_ctrl[8][17] , \sa_ctrl[8].f.spare[12] );
tran (\sa_ctrl[8][18] , \sa_ctrl[8].r.part0[18] );
tran (\sa_ctrl[8][18] , \sa_ctrl[8].f.spare[13] );
tran (\sa_ctrl[8][19] , \sa_ctrl[8].r.part0[19] );
tran (\sa_ctrl[8][19] , \sa_ctrl[8].f.spare[14] );
tran (\sa_ctrl[8][20] , \sa_ctrl[8].r.part0[20] );
tran (\sa_ctrl[8][20] , \sa_ctrl[8].f.spare[15] );
tran (\sa_ctrl[8][21] , \sa_ctrl[8].r.part0[21] );
tran (\sa_ctrl[8][21] , \sa_ctrl[8].f.spare[16] );
tran (\sa_ctrl[8][22] , \sa_ctrl[8].r.part0[22] );
tran (\sa_ctrl[8][22] , \sa_ctrl[8].f.spare[17] );
tran (\sa_ctrl[8][23] , \sa_ctrl[8].r.part0[23] );
tran (\sa_ctrl[8][23] , \sa_ctrl[8].f.spare[18] );
tran (\sa_ctrl[8][24] , \sa_ctrl[8].r.part0[24] );
tran (\sa_ctrl[8][24] , \sa_ctrl[8].f.spare[19] );
tran (\sa_ctrl[8][25] , \sa_ctrl[8].r.part0[25] );
tran (\sa_ctrl[8][25] , \sa_ctrl[8].f.spare[20] );
tran (\sa_ctrl[8][26] , \sa_ctrl[8].r.part0[26] );
tran (\sa_ctrl[8][26] , \sa_ctrl[8].f.spare[21] );
tran (\sa_ctrl[8][27] , \sa_ctrl[8].r.part0[27] );
tran (\sa_ctrl[8][27] , \sa_ctrl[8].f.spare[22] );
tran (\sa_ctrl[8][28] , \sa_ctrl[8].r.part0[28] );
tran (\sa_ctrl[8][28] , \sa_ctrl[8].f.spare[23] );
tran (\sa_ctrl[8][29] , \sa_ctrl[8].r.part0[29] );
tran (\sa_ctrl[8][29] , \sa_ctrl[8].f.spare[24] );
tran (\sa_ctrl[8][30] , \sa_ctrl[8].r.part0[30] );
tran (\sa_ctrl[8][30] , \sa_ctrl[8].f.spare[25] );
tran (\sa_ctrl[8][31] , \sa_ctrl[8].r.part0[31] );
tran (\sa_ctrl[8][31] , \sa_ctrl[8].f.spare[26] );
tran (\sa_ctrl[9][0] , \sa_ctrl[9].r.part0[0] );
tran (\sa_ctrl[9][0] , \sa_ctrl[9].f.sa_event_sel[0] );
tran (\sa_ctrl[9][1] , \sa_ctrl[9].r.part0[1] );
tran (\sa_ctrl[9][1] , \sa_ctrl[9].f.sa_event_sel[1] );
tran (\sa_ctrl[9][2] , \sa_ctrl[9].r.part0[2] );
tran (\sa_ctrl[9][2] , \sa_ctrl[9].f.sa_event_sel[2] );
tran (\sa_ctrl[9][3] , \sa_ctrl[9].r.part0[3] );
tran (\sa_ctrl[9][3] , \sa_ctrl[9].f.sa_event_sel[3] );
tran (\sa_ctrl[9][4] , \sa_ctrl[9].r.part0[4] );
tran (\sa_ctrl[9][4] , \sa_ctrl[9].f.sa_event_sel[4] );
tran (\sa_ctrl[9][5] , \sa_ctrl[9].r.part0[5] );
tran (\sa_ctrl[9][5] , \sa_ctrl[9].f.spare[0] );
tran (\sa_ctrl[9][6] , \sa_ctrl[9].r.part0[6] );
tran (\sa_ctrl[9][6] , \sa_ctrl[9].f.spare[1] );
tran (\sa_ctrl[9][7] , \sa_ctrl[9].r.part0[7] );
tran (\sa_ctrl[9][7] , \sa_ctrl[9].f.spare[2] );
tran (\sa_ctrl[9][8] , \sa_ctrl[9].r.part0[8] );
tran (\sa_ctrl[9][8] , \sa_ctrl[9].f.spare[3] );
tran (\sa_ctrl[9][9] , \sa_ctrl[9].r.part0[9] );
tran (\sa_ctrl[9][9] , \sa_ctrl[9].f.spare[4] );
tran (\sa_ctrl[9][10] , \sa_ctrl[9].r.part0[10] );
tran (\sa_ctrl[9][10] , \sa_ctrl[9].f.spare[5] );
tran (\sa_ctrl[9][11] , \sa_ctrl[9].r.part0[11] );
tran (\sa_ctrl[9][11] , \sa_ctrl[9].f.spare[6] );
tran (\sa_ctrl[9][12] , \sa_ctrl[9].r.part0[12] );
tran (\sa_ctrl[9][12] , \sa_ctrl[9].f.spare[7] );
tran (\sa_ctrl[9][13] , \sa_ctrl[9].r.part0[13] );
tran (\sa_ctrl[9][13] , \sa_ctrl[9].f.spare[8] );
tran (\sa_ctrl[9][14] , \sa_ctrl[9].r.part0[14] );
tran (\sa_ctrl[9][14] , \sa_ctrl[9].f.spare[9] );
tran (\sa_ctrl[9][15] , \sa_ctrl[9].r.part0[15] );
tran (\sa_ctrl[9][15] , \sa_ctrl[9].f.spare[10] );
tran (\sa_ctrl[9][16] , \sa_ctrl[9].r.part0[16] );
tran (\sa_ctrl[9][16] , \sa_ctrl[9].f.spare[11] );
tran (\sa_ctrl[9][17] , \sa_ctrl[9].r.part0[17] );
tran (\sa_ctrl[9][17] , \sa_ctrl[9].f.spare[12] );
tran (\sa_ctrl[9][18] , \sa_ctrl[9].r.part0[18] );
tran (\sa_ctrl[9][18] , \sa_ctrl[9].f.spare[13] );
tran (\sa_ctrl[9][19] , \sa_ctrl[9].r.part0[19] );
tran (\sa_ctrl[9][19] , \sa_ctrl[9].f.spare[14] );
tran (\sa_ctrl[9][20] , \sa_ctrl[9].r.part0[20] );
tran (\sa_ctrl[9][20] , \sa_ctrl[9].f.spare[15] );
tran (\sa_ctrl[9][21] , \sa_ctrl[9].r.part0[21] );
tran (\sa_ctrl[9][21] , \sa_ctrl[9].f.spare[16] );
tran (\sa_ctrl[9][22] , \sa_ctrl[9].r.part0[22] );
tran (\sa_ctrl[9][22] , \sa_ctrl[9].f.spare[17] );
tran (\sa_ctrl[9][23] , \sa_ctrl[9].r.part0[23] );
tran (\sa_ctrl[9][23] , \sa_ctrl[9].f.spare[18] );
tran (\sa_ctrl[9][24] , \sa_ctrl[9].r.part0[24] );
tran (\sa_ctrl[9][24] , \sa_ctrl[9].f.spare[19] );
tran (\sa_ctrl[9][25] , \sa_ctrl[9].r.part0[25] );
tran (\sa_ctrl[9][25] , \sa_ctrl[9].f.spare[20] );
tran (\sa_ctrl[9][26] , \sa_ctrl[9].r.part0[26] );
tran (\sa_ctrl[9][26] , \sa_ctrl[9].f.spare[21] );
tran (\sa_ctrl[9][27] , \sa_ctrl[9].r.part0[27] );
tran (\sa_ctrl[9][27] , \sa_ctrl[9].f.spare[22] );
tran (\sa_ctrl[9][28] , \sa_ctrl[9].r.part0[28] );
tran (\sa_ctrl[9][28] , \sa_ctrl[9].f.spare[23] );
tran (\sa_ctrl[9][29] , \sa_ctrl[9].r.part0[29] );
tran (\sa_ctrl[9][29] , \sa_ctrl[9].f.spare[24] );
tran (\sa_ctrl[9][30] , \sa_ctrl[9].r.part0[30] );
tran (\sa_ctrl[9][30] , \sa_ctrl[9].f.spare[25] );
tran (\sa_ctrl[9][31] , \sa_ctrl[9].r.part0[31] );
tran (\sa_ctrl[9][31] , \sa_ctrl[9].f.spare[26] );
tran (\sa_ctrl[10][0] , \sa_ctrl[10].r.part0[0] );
tran (\sa_ctrl[10][0] , \sa_ctrl[10].f.sa_event_sel[0] );
tran (\sa_ctrl[10][1] , \sa_ctrl[10].r.part0[1] );
tran (\sa_ctrl[10][1] , \sa_ctrl[10].f.sa_event_sel[1] );
tran (\sa_ctrl[10][2] , \sa_ctrl[10].r.part0[2] );
tran (\sa_ctrl[10][2] , \sa_ctrl[10].f.sa_event_sel[2] );
tran (\sa_ctrl[10][3] , \sa_ctrl[10].r.part0[3] );
tran (\sa_ctrl[10][3] , \sa_ctrl[10].f.sa_event_sel[3] );
tran (\sa_ctrl[10][4] , \sa_ctrl[10].r.part0[4] );
tran (\sa_ctrl[10][4] , \sa_ctrl[10].f.sa_event_sel[4] );
tran (\sa_ctrl[10][5] , \sa_ctrl[10].r.part0[5] );
tran (\sa_ctrl[10][5] , \sa_ctrl[10].f.spare[0] );
tran (\sa_ctrl[10][6] , \sa_ctrl[10].r.part0[6] );
tran (\sa_ctrl[10][6] , \sa_ctrl[10].f.spare[1] );
tran (\sa_ctrl[10][7] , \sa_ctrl[10].r.part0[7] );
tran (\sa_ctrl[10][7] , \sa_ctrl[10].f.spare[2] );
tran (\sa_ctrl[10][8] , \sa_ctrl[10].r.part0[8] );
tran (\sa_ctrl[10][8] , \sa_ctrl[10].f.spare[3] );
tran (\sa_ctrl[10][9] , \sa_ctrl[10].r.part0[9] );
tran (\sa_ctrl[10][9] , \sa_ctrl[10].f.spare[4] );
tran (\sa_ctrl[10][10] , \sa_ctrl[10].r.part0[10] );
tran (\sa_ctrl[10][10] , \sa_ctrl[10].f.spare[5] );
tran (\sa_ctrl[10][11] , \sa_ctrl[10].r.part0[11] );
tran (\sa_ctrl[10][11] , \sa_ctrl[10].f.spare[6] );
tran (\sa_ctrl[10][12] , \sa_ctrl[10].r.part0[12] );
tran (\sa_ctrl[10][12] , \sa_ctrl[10].f.spare[7] );
tran (\sa_ctrl[10][13] , \sa_ctrl[10].r.part0[13] );
tran (\sa_ctrl[10][13] , \sa_ctrl[10].f.spare[8] );
tran (\sa_ctrl[10][14] , \sa_ctrl[10].r.part0[14] );
tran (\sa_ctrl[10][14] , \sa_ctrl[10].f.spare[9] );
tran (\sa_ctrl[10][15] , \sa_ctrl[10].r.part0[15] );
tran (\sa_ctrl[10][15] , \sa_ctrl[10].f.spare[10] );
tran (\sa_ctrl[10][16] , \sa_ctrl[10].r.part0[16] );
tran (\sa_ctrl[10][16] , \sa_ctrl[10].f.spare[11] );
tran (\sa_ctrl[10][17] , \sa_ctrl[10].r.part0[17] );
tran (\sa_ctrl[10][17] , \sa_ctrl[10].f.spare[12] );
tran (\sa_ctrl[10][18] , \sa_ctrl[10].r.part0[18] );
tran (\sa_ctrl[10][18] , \sa_ctrl[10].f.spare[13] );
tran (\sa_ctrl[10][19] , \sa_ctrl[10].r.part0[19] );
tran (\sa_ctrl[10][19] , \sa_ctrl[10].f.spare[14] );
tran (\sa_ctrl[10][20] , \sa_ctrl[10].r.part0[20] );
tran (\sa_ctrl[10][20] , \sa_ctrl[10].f.spare[15] );
tran (\sa_ctrl[10][21] , \sa_ctrl[10].r.part0[21] );
tran (\sa_ctrl[10][21] , \sa_ctrl[10].f.spare[16] );
tran (\sa_ctrl[10][22] , \sa_ctrl[10].r.part0[22] );
tran (\sa_ctrl[10][22] , \sa_ctrl[10].f.spare[17] );
tran (\sa_ctrl[10][23] , \sa_ctrl[10].r.part0[23] );
tran (\sa_ctrl[10][23] , \sa_ctrl[10].f.spare[18] );
tran (\sa_ctrl[10][24] , \sa_ctrl[10].r.part0[24] );
tran (\sa_ctrl[10][24] , \sa_ctrl[10].f.spare[19] );
tran (\sa_ctrl[10][25] , \sa_ctrl[10].r.part0[25] );
tran (\sa_ctrl[10][25] , \sa_ctrl[10].f.spare[20] );
tran (\sa_ctrl[10][26] , \sa_ctrl[10].r.part0[26] );
tran (\sa_ctrl[10][26] , \sa_ctrl[10].f.spare[21] );
tran (\sa_ctrl[10][27] , \sa_ctrl[10].r.part0[27] );
tran (\sa_ctrl[10][27] , \sa_ctrl[10].f.spare[22] );
tran (\sa_ctrl[10][28] , \sa_ctrl[10].r.part0[28] );
tran (\sa_ctrl[10][28] , \sa_ctrl[10].f.spare[23] );
tran (\sa_ctrl[10][29] , \sa_ctrl[10].r.part0[29] );
tran (\sa_ctrl[10][29] , \sa_ctrl[10].f.spare[24] );
tran (\sa_ctrl[10][30] , \sa_ctrl[10].r.part0[30] );
tran (\sa_ctrl[10][30] , \sa_ctrl[10].f.spare[25] );
tran (\sa_ctrl[10][31] , \sa_ctrl[10].r.part0[31] );
tran (\sa_ctrl[10][31] , \sa_ctrl[10].f.spare[26] );
tran (\sa_ctrl[11][0] , \sa_ctrl[11].r.part0[0] );
tran (\sa_ctrl[11][0] , \sa_ctrl[11].f.sa_event_sel[0] );
tran (\sa_ctrl[11][1] , \sa_ctrl[11].r.part0[1] );
tran (\sa_ctrl[11][1] , \sa_ctrl[11].f.sa_event_sel[1] );
tran (\sa_ctrl[11][2] , \sa_ctrl[11].r.part0[2] );
tran (\sa_ctrl[11][2] , \sa_ctrl[11].f.sa_event_sel[2] );
tran (\sa_ctrl[11][3] , \sa_ctrl[11].r.part0[3] );
tran (\sa_ctrl[11][3] , \sa_ctrl[11].f.sa_event_sel[3] );
tran (\sa_ctrl[11][4] , \sa_ctrl[11].r.part0[4] );
tran (\sa_ctrl[11][4] , \sa_ctrl[11].f.sa_event_sel[4] );
tran (\sa_ctrl[11][5] , \sa_ctrl[11].r.part0[5] );
tran (\sa_ctrl[11][5] , \sa_ctrl[11].f.spare[0] );
tran (\sa_ctrl[11][6] , \sa_ctrl[11].r.part0[6] );
tran (\sa_ctrl[11][6] , \sa_ctrl[11].f.spare[1] );
tran (\sa_ctrl[11][7] , \sa_ctrl[11].r.part0[7] );
tran (\sa_ctrl[11][7] , \sa_ctrl[11].f.spare[2] );
tran (\sa_ctrl[11][8] , \sa_ctrl[11].r.part0[8] );
tran (\sa_ctrl[11][8] , \sa_ctrl[11].f.spare[3] );
tran (\sa_ctrl[11][9] , \sa_ctrl[11].r.part0[9] );
tran (\sa_ctrl[11][9] , \sa_ctrl[11].f.spare[4] );
tran (\sa_ctrl[11][10] , \sa_ctrl[11].r.part0[10] );
tran (\sa_ctrl[11][10] , \sa_ctrl[11].f.spare[5] );
tran (\sa_ctrl[11][11] , \sa_ctrl[11].r.part0[11] );
tran (\sa_ctrl[11][11] , \sa_ctrl[11].f.spare[6] );
tran (\sa_ctrl[11][12] , \sa_ctrl[11].r.part0[12] );
tran (\sa_ctrl[11][12] , \sa_ctrl[11].f.spare[7] );
tran (\sa_ctrl[11][13] , \sa_ctrl[11].r.part0[13] );
tran (\sa_ctrl[11][13] , \sa_ctrl[11].f.spare[8] );
tran (\sa_ctrl[11][14] , \sa_ctrl[11].r.part0[14] );
tran (\sa_ctrl[11][14] , \sa_ctrl[11].f.spare[9] );
tran (\sa_ctrl[11][15] , \sa_ctrl[11].r.part0[15] );
tran (\sa_ctrl[11][15] , \sa_ctrl[11].f.spare[10] );
tran (\sa_ctrl[11][16] , \sa_ctrl[11].r.part0[16] );
tran (\sa_ctrl[11][16] , \sa_ctrl[11].f.spare[11] );
tran (\sa_ctrl[11][17] , \sa_ctrl[11].r.part0[17] );
tran (\sa_ctrl[11][17] , \sa_ctrl[11].f.spare[12] );
tran (\sa_ctrl[11][18] , \sa_ctrl[11].r.part0[18] );
tran (\sa_ctrl[11][18] , \sa_ctrl[11].f.spare[13] );
tran (\sa_ctrl[11][19] , \sa_ctrl[11].r.part0[19] );
tran (\sa_ctrl[11][19] , \sa_ctrl[11].f.spare[14] );
tran (\sa_ctrl[11][20] , \sa_ctrl[11].r.part0[20] );
tran (\sa_ctrl[11][20] , \sa_ctrl[11].f.spare[15] );
tran (\sa_ctrl[11][21] , \sa_ctrl[11].r.part0[21] );
tran (\sa_ctrl[11][21] , \sa_ctrl[11].f.spare[16] );
tran (\sa_ctrl[11][22] , \sa_ctrl[11].r.part0[22] );
tran (\sa_ctrl[11][22] , \sa_ctrl[11].f.spare[17] );
tran (\sa_ctrl[11][23] , \sa_ctrl[11].r.part0[23] );
tran (\sa_ctrl[11][23] , \sa_ctrl[11].f.spare[18] );
tran (\sa_ctrl[11][24] , \sa_ctrl[11].r.part0[24] );
tran (\sa_ctrl[11][24] , \sa_ctrl[11].f.spare[19] );
tran (\sa_ctrl[11][25] , \sa_ctrl[11].r.part0[25] );
tran (\sa_ctrl[11][25] , \sa_ctrl[11].f.spare[20] );
tran (\sa_ctrl[11][26] , \sa_ctrl[11].r.part0[26] );
tran (\sa_ctrl[11][26] , \sa_ctrl[11].f.spare[21] );
tran (\sa_ctrl[11][27] , \sa_ctrl[11].r.part0[27] );
tran (\sa_ctrl[11][27] , \sa_ctrl[11].f.spare[22] );
tran (\sa_ctrl[11][28] , \sa_ctrl[11].r.part0[28] );
tran (\sa_ctrl[11][28] , \sa_ctrl[11].f.spare[23] );
tran (\sa_ctrl[11][29] , \sa_ctrl[11].r.part0[29] );
tran (\sa_ctrl[11][29] , \sa_ctrl[11].f.spare[24] );
tran (\sa_ctrl[11][30] , \sa_ctrl[11].r.part0[30] );
tran (\sa_ctrl[11][30] , \sa_ctrl[11].f.spare[25] );
tran (\sa_ctrl[11][31] , \sa_ctrl[11].r.part0[31] );
tran (\sa_ctrl[11][31] , \sa_ctrl[11].f.spare[26] );
tran (\sa_ctrl[12][0] , \sa_ctrl[12].r.part0[0] );
tran (\sa_ctrl[12][0] , \sa_ctrl[12].f.sa_event_sel[0] );
tran (\sa_ctrl[12][1] , \sa_ctrl[12].r.part0[1] );
tran (\sa_ctrl[12][1] , \sa_ctrl[12].f.sa_event_sel[1] );
tran (\sa_ctrl[12][2] , \sa_ctrl[12].r.part0[2] );
tran (\sa_ctrl[12][2] , \sa_ctrl[12].f.sa_event_sel[2] );
tran (\sa_ctrl[12][3] , \sa_ctrl[12].r.part0[3] );
tran (\sa_ctrl[12][3] , \sa_ctrl[12].f.sa_event_sel[3] );
tran (\sa_ctrl[12][4] , \sa_ctrl[12].r.part0[4] );
tran (\sa_ctrl[12][4] , \sa_ctrl[12].f.sa_event_sel[4] );
tran (\sa_ctrl[12][5] , \sa_ctrl[12].r.part0[5] );
tran (\sa_ctrl[12][5] , \sa_ctrl[12].f.spare[0] );
tran (\sa_ctrl[12][6] , \sa_ctrl[12].r.part0[6] );
tran (\sa_ctrl[12][6] , \sa_ctrl[12].f.spare[1] );
tran (\sa_ctrl[12][7] , \sa_ctrl[12].r.part0[7] );
tran (\sa_ctrl[12][7] , \sa_ctrl[12].f.spare[2] );
tran (\sa_ctrl[12][8] , \sa_ctrl[12].r.part0[8] );
tran (\sa_ctrl[12][8] , \sa_ctrl[12].f.spare[3] );
tran (\sa_ctrl[12][9] , \sa_ctrl[12].r.part0[9] );
tran (\sa_ctrl[12][9] , \sa_ctrl[12].f.spare[4] );
tran (\sa_ctrl[12][10] , \sa_ctrl[12].r.part0[10] );
tran (\sa_ctrl[12][10] , \sa_ctrl[12].f.spare[5] );
tran (\sa_ctrl[12][11] , \sa_ctrl[12].r.part0[11] );
tran (\sa_ctrl[12][11] , \sa_ctrl[12].f.spare[6] );
tran (\sa_ctrl[12][12] , \sa_ctrl[12].r.part0[12] );
tran (\sa_ctrl[12][12] , \sa_ctrl[12].f.spare[7] );
tran (\sa_ctrl[12][13] , \sa_ctrl[12].r.part0[13] );
tran (\sa_ctrl[12][13] , \sa_ctrl[12].f.spare[8] );
tran (\sa_ctrl[12][14] , \sa_ctrl[12].r.part0[14] );
tran (\sa_ctrl[12][14] , \sa_ctrl[12].f.spare[9] );
tran (\sa_ctrl[12][15] , \sa_ctrl[12].r.part0[15] );
tran (\sa_ctrl[12][15] , \sa_ctrl[12].f.spare[10] );
tran (\sa_ctrl[12][16] , \sa_ctrl[12].r.part0[16] );
tran (\sa_ctrl[12][16] , \sa_ctrl[12].f.spare[11] );
tran (\sa_ctrl[12][17] , \sa_ctrl[12].r.part0[17] );
tran (\sa_ctrl[12][17] , \sa_ctrl[12].f.spare[12] );
tran (\sa_ctrl[12][18] , \sa_ctrl[12].r.part0[18] );
tran (\sa_ctrl[12][18] , \sa_ctrl[12].f.spare[13] );
tran (\sa_ctrl[12][19] , \sa_ctrl[12].r.part0[19] );
tran (\sa_ctrl[12][19] , \sa_ctrl[12].f.spare[14] );
tran (\sa_ctrl[12][20] , \sa_ctrl[12].r.part0[20] );
tran (\sa_ctrl[12][20] , \sa_ctrl[12].f.spare[15] );
tran (\sa_ctrl[12][21] , \sa_ctrl[12].r.part0[21] );
tran (\sa_ctrl[12][21] , \sa_ctrl[12].f.spare[16] );
tran (\sa_ctrl[12][22] , \sa_ctrl[12].r.part0[22] );
tran (\sa_ctrl[12][22] , \sa_ctrl[12].f.spare[17] );
tran (\sa_ctrl[12][23] , \sa_ctrl[12].r.part0[23] );
tran (\sa_ctrl[12][23] , \sa_ctrl[12].f.spare[18] );
tran (\sa_ctrl[12][24] , \sa_ctrl[12].r.part0[24] );
tran (\sa_ctrl[12][24] , \sa_ctrl[12].f.spare[19] );
tran (\sa_ctrl[12][25] , \sa_ctrl[12].r.part0[25] );
tran (\sa_ctrl[12][25] , \sa_ctrl[12].f.spare[20] );
tran (\sa_ctrl[12][26] , \sa_ctrl[12].r.part0[26] );
tran (\sa_ctrl[12][26] , \sa_ctrl[12].f.spare[21] );
tran (\sa_ctrl[12][27] , \sa_ctrl[12].r.part0[27] );
tran (\sa_ctrl[12][27] , \sa_ctrl[12].f.spare[22] );
tran (\sa_ctrl[12][28] , \sa_ctrl[12].r.part0[28] );
tran (\sa_ctrl[12][28] , \sa_ctrl[12].f.spare[23] );
tran (\sa_ctrl[12][29] , \sa_ctrl[12].r.part0[29] );
tran (\sa_ctrl[12][29] , \sa_ctrl[12].f.spare[24] );
tran (\sa_ctrl[12][30] , \sa_ctrl[12].r.part0[30] );
tran (\sa_ctrl[12][30] , \sa_ctrl[12].f.spare[25] );
tran (\sa_ctrl[12][31] , \sa_ctrl[12].r.part0[31] );
tran (\sa_ctrl[12][31] , \sa_ctrl[12].f.spare[26] );
tran (\sa_ctrl[13][0] , \sa_ctrl[13].r.part0[0] );
tran (\sa_ctrl[13][0] , \sa_ctrl[13].f.sa_event_sel[0] );
tran (\sa_ctrl[13][1] , \sa_ctrl[13].r.part0[1] );
tran (\sa_ctrl[13][1] , \sa_ctrl[13].f.sa_event_sel[1] );
tran (\sa_ctrl[13][2] , \sa_ctrl[13].r.part0[2] );
tran (\sa_ctrl[13][2] , \sa_ctrl[13].f.sa_event_sel[2] );
tran (\sa_ctrl[13][3] , \sa_ctrl[13].r.part0[3] );
tran (\sa_ctrl[13][3] , \sa_ctrl[13].f.sa_event_sel[3] );
tran (\sa_ctrl[13][4] , \sa_ctrl[13].r.part0[4] );
tran (\sa_ctrl[13][4] , \sa_ctrl[13].f.sa_event_sel[4] );
tran (\sa_ctrl[13][5] , \sa_ctrl[13].r.part0[5] );
tran (\sa_ctrl[13][5] , \sa_ctrl[13].f.spare[0] );
tran (\sa_ctrl[13][6] , \sa_ctrl[13].r.part0[6] );
tran (\sa_ctrl[13][6] , \sa_ctrl[13].f.spare[1] );
tran (\sa_ctrl[13][7] , \sa_ctrl[13].r.part0[7] );
tran (\sa_ctrl[13][7] , \sa_ctrl[13].f.spare[2] );
tran (\sa_ctrl[13][8] , \sa_ctrl[13].r.part0[8] );
tran (\sa_ctrl[13][8] , \sa_ctrl[13].f.spare[3] );
tran (\sa_ctrl[13][9] , \sa_ctrl[13].r.part0[9] );
tran (\sa_ctrl[13][9] , \sa_ctrl[13].f.spare[4] );
tran (\sa_ctrl[13][10] , \sa_ctrl[13].r.part0[10] );
tran (\sa_ctrl[13][10] , \sa_ctrl[13].f.spare[5] );
tran (\sa_ctrl[13][11] , \sa_ctrl[13].r.part0[11] );
tran (\sa_ctrl[13][11] , \sa_ctrl[13].f.spare[6] );
tran (\sa_ctrl[13][12] , \sa_ctrl[13].r.part0[12] );
tran (\sa_ctrl[13][12] , \sa_ctrl[13].f.spare[7] );
tran (\sa_ctrl[13][13] , \sa_ctrl[13].r.part0[13] );
tran (\sa_ctrl[13][13] , \sa_ctrl[13].f.spare[8] );
tran (\sa_ctrl[13][14] , \sa_ctrl[13].r.part0[14] );
tran (\sa_ctrl[13][14] , \sa_ctrl[13].f.spare[9] );
tran (\sa_ctrl[13][15] , \sa_ctrl[13].r.part0[15] );
tran (\sa_ctrl[13][15] , \sa_ctrl[13].f.spare[10] );
tran (\sa_ctrl[13][16] , \sa_ctrl[13].r.part0[16] );
tran (\sa_ctrl[13][16] , \sa_ctrl[13].f.spare[11] );
tran (\sa_ctrl[13][17] , \sa_ctrl[13].r.part0[17] );
tran (\sa_ctrl[13][17] , \sa_ctrl[13].f.spare[12] );
tran (\sa_ctrl[13][18] , \sa_ctrl[13].r.part0[18] );
tran (\sa_ctrl[13][18] , \sa_ctrl[13].f.spare[13] );
tran (\sa_ctrl[13][19] , \sa_ctrl[13].r.part0[19] );
tran (\sa_ctrl[13][19] , \sa_ctrl[13].f.spare[14] );
tran (\sa_ctrl[13][20] , \sa_ctrl[13].r.part0[20] );
tran (\sa_ctrl[13][20] , \sa_ctrl[13].f.spare[15] );
tran (\sa_ctrl[13][21] , \sa_ctrl[13].r.part0[21] );
tran (\sa_ctrl[13][21] , \sa_ctrl[13].f.spare[16] );
tran (\sa_ctrl[13][22] , \sa_ctrl[13].r.part0[22] );
tran (\sa_ctrl[13][22] , \sa_ctrl[13].f.spare[17] );
tran (\sa_ctrl[13][23] , \sa_ctrl[13].r.part0[23] );
tran (\sa_ctrl[13][23] , \sa_ctrl[13].f.spare[18] );
tran (\sa_ctrl[13][24] , \sa_ctrl[13].r.part0[24] );
tran (\sa_ctrl[13][24] , \sa_ctrl[13].f.spare[19] );
tran (\sa_ctrl[13][25] , \sa_ctrl[13].r.part0[25] );
tran (\sa_ctrl[13][25] , \sa_ctrl[13].f.spare[20] );
tran (\sa_ctrl[13][26] , \sa_ctrl[13].r.part0[26] );
tran (\sa_ctrl[13][26] , \sa_ctrl[13].f.spare[21] );
tran (\sa_ctrl[13][27] , \sa_ctrl[13].r.part0[27] );
tran (\sa_ctrl[13][27] , \sa_ctrl[13].f.spare[22] );
tran (\sa_ctrl[13][28] , \sa_ctrl[13].r.part0[28] );
tran (\sa_ctrl[13][28] , \sa_ctrl[13].f.spare[23] );
tran (\sa_ctrl[13][29] , \sa_ctrl[13].r.part0[29] );
tran (\sa_ctrl[13][29] , \sa_ctrl[13].f.spare[24] );
tran (\sa_ctrl[13][30] , \sa_ctrl[13].r.part0[30] );
tran (\sa_ctrl[13][30] , \sa_ctrl[13].f.spare[25] );
tran (\sa_ctrl[13][31] , \sa_ctrl[13].r.part0[31] );
tran (\sa_ctrl[13][31] , \sa_ctrl[13].f.spare[26] );
tran (\sa_ctrl[14][0] , \sa_ctrl[14].r.part0[0] );
tran (\sa_ctrl[14][0] , \sa_ctrl[14].f.sa_event_sel[0] );
tran (\sa_ctrl[14][1] , \sa_ctrl[14].r.part0[1] );
tran (\sa_ctrl[14][1] , \sa_ctrl[14].f.sa_event_sel[1] );
tran (\sa_ctrl[14][2] , \sa_ctrl[14].r.part0[2] );
tran (\sa_ctrl[14][2] , \sa_ctrl[14].f.sa_event_sel[2] );
tran (\sa_ctrl[14][3] , \sa_ctrl[14].r.part0[3] );
tran (\sa_ctrl[14][3] , \sa_ctrl[14].f.sa_event_sel[3] );
tran (\sa_ctrl[14][4] , \sa_ctrl[14].r.part0[4] );
tran (\sa_ctrl[14][4] , \sa_ctrl[14].f.sa_event_sel[4] );
tran (\sa_ctrl[14][5] , \sa_ctrl[14].r.part0[5] );
tran (\sa_ctrl[14][5] , \sa_ctrl[14].f.spare[0] );
tran (\sa_ctrl[14][6] , \sa_ctrl[14].r.part0[6] );
tran (\sa_ctrl[14][6] , \sa_ctrl[14].f.spare[1] );
tran (\sa_ctrl[14][7] , \sa_ctrl[14].r.part0[7] );
tran (\sa_ctrl[14][7] , \sa_ctrl[14].f.spare[2] );
tran (\sa_ctrl[14][8] , \sa_ctrl[14].r.part0[8] );
tran (\sa_ctrl[14][8] , \sa_ctrl[14].f.spare[3] );
tran (\sa_ctrl[14][9] , \sa_ctrl[14].r.part0[9] );
tran (\sa_ctrl[14][9] , \sa_ctrl[14].f.spare[4] );
tran (\sa_ctrl[14][10] , \sa_ctrl[14].r.part0[10] );
tran (\sa_ctrl[14][10] , \sa_ctrl[14].f.spare[5] );
tran (\sa_ctrl[14][11] , \sa_ctrl[14].r.part0[11] );
tran (\sa_ctrl[14][11] , \sa_ctrl[14].f.spare[6] );
tran (\sa_ctrl[14][12] , \sa_ctrl[14].r.part0[12] );
tran (\sa_ctrl[14][12] , \sa_ctrl[14].f.spare[7] );
tran (\sa_ctrl[14][13] , \sa_ctrl[14].r.part0[13] );
tran (\sa_ctrl[14][13] , \sa_ctrl[14].f.spare[8] );
tran (\sa_ctrl[14][14] , \sa_ctrl[14].r.part0[14] );
tran (\sa_ctrl[14][14] , \sa_ctrl[14].f.spare[9] );
tran (\sa_ctrl[14][15] , \sa_ctrl[14].r.part0[15] );
tran (\sa_ctrl[14][15] , \sa_ctrl[14].f.spare[10] );
tran (\sa_ctrl[14][16] , \sa_ctrl[14].r.part0[16] );
tran (\sa_ctrl[14][16] , \sa_ctrl[14].f.spare[11] );
tran (\sa_ctrl[14][17] , \sa_ctrl[14].r.part0[17] );
tran (\sa_ctrl[14][17] , \sa_ctrl[14].f.spare[12] );
tran (\sa_ctrl[14][18] , \sa_ctrl[14].r.part0[18] );
tran (\sa_ctrl[14][18] , \sa_ctrl[14].f.spare[13] );
tran (\sa_ctrl[14][19] , \sa_ctrl[14].r.part0[19] );
tran (\sa_ctrl[14][19] , \sa_ctrl[14].f.spare[14] );
tran (\sa_ctrl[14][20] , \sa_ctrl[14].r.part0[20] );
tran (\sa_ctrl[14][20] , \sa_ctrl[14].f.spare[15] );
tran (\sa_ctrl[14][21] , \sa_ctrl[14].r.part0[21] );
tran (\sa_ctrl[14][21] , \sa_ctrl[14].f.spare[16] );
tran (\sa_ctrl[14][22] , \sa_ctrl[14].r.part0[22] );
tran (\sa_ctrl[14][22] , \sa_ctrl[14].f.spare[17] );
tran (\sa_ctrl[14][23] , \sa_ctrl[14].r.part0[23] );
tran (\sa_ctrl[14][23] , \sa_ctrl[14].f.spare[18] );
tran (\sa_ctrl[14][24] , \sa_ctrl[14].r.part0[24] );
tran (\sa_ctrl[14][24] , \sa_ctrl[14].f.spare[19] );
tran (\sa_ctrl[14][25] , \sa_ctrl[14].r.part0[25] );
tran (\sa_ctrl[14][25] , \sa_ctrl[14].f.spare[20] );
tran (\sa_ctrl[14][26] , \sa_ctrl[14].r.part0[26] );
tran (\sa_ctrl[14][26] , \sa_ctrl[14].f.spare[21] );
tran (\sa_ctrl[14][27] , \sa_ctrl[14].r.part0[27] );
tran (\sa_ctrl[14][27] , \sa_ctrl[14].f.spare[22] );
tran (\sa_ctrl[14][28] , \sa_ctrl[14].r.part0[28] );
tran (\sa_ctrl[14][28] , \sa_ctrl[14].f.spare[23] );
tran (\sa_ctrl[14][29] , \sa_ctrl[14].r.part0[29] );
tran (\sa_ctrl[14][29] , \sa_ctrl[14].f.spare[24] );
tran (\sa_ctrl[14][30] , \sa_ctrl[14].r.part0[30] );
tran (\sa_ctrl[14][30] , \sa_ctrl[14].f.spare[25] );
tran (\sa_ctrl[14][31] , \sa_ctrl[14].r.part0[31] );
tran (\sa_ctrl[14][31] , \sa_ctrl[14].f.spare[26] );
tran (\sa_ctrl[15][0] , \sa_ctrl[15].r.part0[0] );
tran (\sa_ctrl[15][0] , \sa_ctrl[15].f.sa_event_sel[0] );
tran (\sa_ctrl[15][1] , \sa_ctrl[15].r.part0[1] );
tran (\sa_ctrl[15][1] , \sa_ctrl[15].f.sa_event_sel[1] );
tran (\sa_ctrl[15][2] , \sa_ctrl[15].r.part0[2] );
tran (\sa_ctrl[15][2] , \sa_ctrl[15].f.sa_event_sel[2] );
tran (\sa_ctrl[15][3] , \sa_ctrl[15].r.part0[3] );
tran (\sa_ctrl[15][3] , \sa_ctrl[15].f.sa_event_sel[3] );
tran (\sa_ctrl[15][4] , \sa_ctrl[15].r.part0[4] );
tran (\sa_ctrl[15][4] , \sa_ctrl[15].f.sa_event_sel[4] );
tran (\sa_ctrl[15][5] , \sa_ctrl[15].r.part0[5] );
tran (\sa_ctrl[15][5] , \sa_ctrl[15].f.spare[0] );
tran (\sa_ctrl[15][6] , \sa_ctrl[15].r.part0[6] );
tran (\sa_ctrl[15][6] , \sa_ctrl[15].f.spare[1] );
tran (\sa_ctrl[15][7] , \sa_ctrl[15].r.part0[7] );
tran (\sa_ctrl[15][7] , \sa_ctrl[15].f.spare[2] );
tran (\sa_ctrl[15][8] , \sa_ctrl[15].r.part0[8] );
tran (\sa_ctrl[15][8] , \sa_ctrl[15].f.spare[3] );
tran (\sa_ctrl[15][9] , \sa_ctrl[15].r.part0[9] );
tran (\sa_ctrl[15][9] , \sa_ctrl[15].f.spare[4] );
tran (\sa_ctrl[15][10] , \sa_ctrl[15].r.part0[10] );
tran (\sa_ctrl[15][10] , \sa_ctrl[15].f.spare[5] );
tran (\sa_ctrl[15][11] , \sa_ctrl[15].r.part0[11] );
tran (\sa_ctrl[15][11] , \sa_ctrl[15].f.spare[6] );
tran (\sa_ctrl[15][12] , \sa_ctrl[15].r.part0[12] );
tran (\sa_ctrl[15][12] , \sa_ctrl[15].f.spare[7] );
tran (\sa_ctrl[15][13] , \sa_ctrl[15].r.part0[13] );
tran (\sa_ctrl[15][13] , \sa_ctrl[15].f.spare[8] );
tran (\sa_ctrl[15][14] , \sa_ctrl[15].r.part0[14] );
tran (\sa_ctrl[15][14] , \sa_ctrl[15].f.spare[9] );
tran (\sa_ctrl[15][15] , \sa_ctrl[15].r.part0[15] );
tran (\sa_ctrl[15][15] , \sa_ctrl[15].f.spare[10] );
tran (\sa_ctrl[15][16] , \sa_ctrl[15].r.part0[16] );
tran (\sa_ctrl[15][16] , \sa_ctrl[15].f.spare[11] );
tran (\sa_ctrl[15][17] , \sa_ctrl[15].r.part0[17] );
tran (\sa_ctrl[15][17] , \sa_ctrl[15].f.spare[12] );
tran (\sa_ctrl[15][18] , \sa_ctrl[15].r.part0[18] );
tran (\sa_ctrl[15][18] , \sa_ctrl[15].f.spare[13] );
tran (\sa_ctrl[15][19] , \sa_ctrl[15].r.part0[19] );
tran (\sa_ctrl[15][19] , \sa_ctrl[15].f.spare[14] );
tran (\sa_ctrl[15][20] , \sa_ctrl[15].r.part0[20] );
tran (\sa_ctrl[15][20] , \sa_ctrl[15].f.spare[15] );
tran (\sa_ctrl[15][21] , \sa_ctrl[15].r.part0[21] );
tran (\sa_ctrl[15][21] , \sa_ctrl[15].f.spare[16] );
tran (\sa_ctrl[15][22] , \sa_ctrl[15].r.part0[22] );
tran (\sa_ctrl[15][22] , \sa_ctrl[15].f.spare[17] );
tran (\sa_ctrl[15][23] , \sa_ctrl[15].r.part0[23] );
tran (\sa_ctrl[15][23] , \sa_ctrl[15].f.spare[18] );
tran (\sa_ctrl[15][24] , \sa_ctrl[15].r.part0[24] );
tran (\sa_ctrl[15][24] , \sa_ctrl[15].f.spare[19] );
tran (\sa_ctrl[15][25] , \sa_ctrl[15].r.part0[25] );
tran (\sa_ctrl[15][25] , \sa_ctrl[15].f.spare[20] );
tran (\sa_ctrl[15][26] , \sa_ctrl[15].r.part0[26] );
tran (\sa_ctrl[15][26] , \sa_ctrl[15].f.spare[21] );
tran (\sa_ctrl[15][27] , \sa_ctrl[15].r.part0[27] );
tran (\sa_ctrl[15][27] , \sa_ctrl[15].f.spare[22] );
tran (\sa_ctrl[15][28] , \sa_ctrl[15].r.part0[28] );
tran (\sa_ctrl[15][28] , \sa_ctrl[15].f.spare[23] );
tran (\sa_ctrl[15][29] , \sa_ctrl[15].r.part0[29] );
tran (\sa_ctrl[15][29] , \sa_ctrl[15].f.spare[24] );
tran (\sa_ctrl[15][30] , \sa_ctrl[15].r.part0[30] );
tran (\sa_ctrl[15][30] , \sa_ctrl[15].f.spare[25] );
tran (\sa_ctrl[15][31] , \sa_ctrl[15].r.part0[31] );
tran (\sa_ctrl[15][31] , \sa_ctrl[15].f.spare[26] );
tran (\sa_ctrl[16][0] , \sa_ctrl[16].r.part0[0] );
tran (\sa_ctrl[16][0] , \sa_ctrl[16].f.sa_event_sel[0] );
tran (\sa_ctrl[16][1] , \sa_ctrl[16].r.part0[1] );
tran (\sa_ctrl[16][1] , \sa_ctrl[16].f.sa_event_sel[1] );
tran (\sa_ctrl[16][2] , \sa_ctrl[16].r.part0[2] );
tran (\sa_ctrl[16][2] , \sa_ctrl[16].f.sa_event_sel[2] );
tran (\sa_ctrl[16][3] , \sa_ctrl[16].r.part0[3] );
tran (\sa_ctrl[16][3] , \sa_ctrl[16].f.sa_event_sel[3] );
tran (\sa_ctrl[16][4] , \sa_ctrl[16].r.part0[4] );
tran (\sa_ctrl[16][4] , \sa_ctrl[16].f.sa_event_sel[4] );
tran (\sa_ctrl[16][5] , \sa_ctrl[16].r.part0[5] );
tran (\sa_ctrl[16][5] , \sa_ctrl[16].f.spare[0] );
tran (\sa_ctrl[16][6] , \sa_ctrl[16].r.part0[6] );
tran (\sa_ctrl[16][6] , \sa_ctrl[16].f.spare[1] );
tran (\sa_ctrl[16][7] , \sa_ctrl[16].r.part0[7] );
tran (\sa_ctrl[16][7] , \sa_ctrl[16].f.spare[2] );
tran (\sa_ctrl[16][8] , \sa_ctrl[16].r.part0[8] );
tran (\sa_ctrl[16][8] , \sa_ctrl[16].f.spare[3] );
tran (\sa_ctrl[16][9] , \sa_ctrl[16].r.part0[9] );
tran (\sa_ctrl[16][9] , \sa_ctrl[16].f.spare[4] );
tran (\sa_ctrl[16][10] , \sa_ctrl[16].r.part0[10] );
tran (\sa_ctrl[16][10] , \sa_ctrl[16].f.spare[5] );
tran (\sa_ctrl[16][11] , \sa_ctrl[16].r.part0[11] );
tran (\sa_ctrl[16][11] , \sa_ctrl[16].f.spare[6] );
tran (\sa_ctrl[16][12] , \sa_ctrl[16].r.part0[12] );
tran (\sa_ctrl[16][12] , \sa_ctrl[16].f.spare[7] );
tran (\sa_ctrl[16][13] , \sa_ctrl[16].r.part0[13] );
tran (\sa_ctrl[16][13] , \sa_ctrl[16].f.spare[8] );
tran (\sa_ctrl[16][14] , \sa_ctrl[16].r.part0[14] );
tran (\sa_ctrl[16][14] , \sa_ctrl[16].f.spare[9] );
tran (\sa_ctrl[16][15] , \sa_ctrl[16].r.part0[15] );
tran (\sa_ctrl[16][15] , \sa_ctrl[16].f.spare[10] );
tran (\sa_ctrl[16][16] , \sa_ctrl[16].r.part0[16] );
tran (\sa_ctrl[16][16] , \sa_ctrl[16].f.spare[11] );
tran (\sa_ctrl[16][17] , \sa_ctrl[16].r.part0[17] );
tran (\sa_ctrl[16][17] , \sa_ctrl[16].f.spare[12] );
tran (\sa_ctrl[16][18] , \sa_ctrl[16].r.part0[18] );
tran (\sa_ctrl[16][18] , \sa_ctrl[16].f.spare[13] );
tran (\sa_ctrl[16][19] , \sa_ctrl[16].r.part0[19] );
tran (\sa_ctrl[16][19] , \sa_ctrl[16].f.spare[14] );
tran (\sa_ctrl[16][20] , \sa_ctrl[16].r.part0[20] );
tran (\sa_ctrl[16][20] , \sa_ctrl[16].f.spare[15] );
tran (\sa_ctrl[16][21] , \sa_ctrl[16].r.part0[21] );
tran (\sa_ctrl[16][21] , \sa_ctrl[16].f.spare[16] );
tran (\sa_ctrl[16][22] , \sa_ctrl[16].r.part0[22] );
tran (\sa_ctrl[16][22] , \sa_ctrl[16].f.spare[17] );
tran (\sa_ctrl[16][23] , \sa_ctrl[16].r.part0[23] );
tran (\sa_ctrl[16][23] , \sa_ctrl[16].f.spare[18] );
tran (\sa_ctrl[16][24] , \sa_ctrl[16].r.part0[24] );
tran (\sa_ctrl[16][24] , \sa_ctrl[16].f.spare[19] );
tran (\sa_ctrl[16][25] , \sa_ctrl[16].r.part0[25] );
tran (\sa_ctrl[16][25] , \sa_ctrl[16].f.spare[20] );
tran (\sa_ctrl[16][26] , \sa_ctrl[16].r.part0[26] );
tran (\sa_ctrl[16][26] , \sa_ctrl[16].f.spare[21] );
tran (\sa_ctrl[16][27] , \sa_ctrl[16].r.part0[27] );
tran (\sa_ctrl[16][27] , \sa_ctrl[16].f.spare[22] );
tran (\sa_ctrl[16][28] , \sa_ctrl[16].r.part0[28] );
tran (\sa_ctrl[16][28] , \sa_ctrl[16].f.spare[23] );
tran (\sa_ctrl[16][29] , \sa_ctrl[16].r.part0[29] );
tran (\sa_ctrl[16][29] , \sa_ctrl[16].f.spare[24] );
tran (\sa_ctrl[16][30] , \sa_ctrl[16].r.part0[30] );
tran (\sa_ctrl[16][30] , \sa_ctrl[16].f.spare[25] );
tran (\sa_ctrl[16][31] , \sa_ctrl[16].r.part0[31] );
tran (\sa_ctrl[16][31] , \sa_ctrl[16].f.spare[26] );
tran (\sa_ctrl[17][0] , \sa_ctrl[17].r.part0[0] );
tran (\sa_ctrl[17][0] , \sa_ctrl[17].f.sa_event_sel[0] );
tran (\sa_ctrl[17][1] , \sa_ctrl[17].r.part0[1] );
tran (\sa_ctrl[17][1] , \sa_ctrl[17].f.sa_event_sel[1] );
tran (\sa_ctrl[17][2] , \sa_ctrl[17].r.part0[2] );
tran (\sa_ctrl[17][2] , \sa_ctrl[17].f.sa_event_sel[2] );
tran (\sa_ctrl[17][3] , \sa_ctrl[17].r.part0[3] );
tran (\sa_ctrl[17][3] , \sa_ctrl[17].f.sa_event_sel[3] );
tran (\sa_ctrl[17][4] , \sa_ctrl[17].r.part0[4] );
tran (\sa_ctrl[17][4] , \sa_ctrl[17].f.sa_event_sel[4] );
tran (\sa_ctrl[17][5] , \sa_ctrl[17].r.part0[5] );
tran (\sa_ctrl[17][5] , \sa_ctrl[17].f.spare[0] );
tran (\sa_ctrl[17][6] , \sa_ctrl[17].r.part0[6] );
tran (\sa_ctrl[17][6] , \sa_ctrl[17].f.spare[1] );
tran (\sa_ctrl[17][7] , \sa_ctrl[17].r.part0[7] );
tran (\sa_ctrl[17][7] , \sa_ctrl[17].f.spare[2] );
tran (\sa_ctrl[17][8] , \sa_ctrl[17].r.part0[8] );
tran (\sa_ctrl[17][8] , \sa_ctrl[17].f.spare[3] );
tran (\sa_ctrl[17][9] , \sa_ctrl[17].r.part0[9] );
tran (\sa_ctrl[17][9] , \sa_ctrl[17].f.spare[4] );
tran (\sa_ctrl[17][10] , \sa_ctrl[17].r.part0[10] );
tran (\sa_ctrl[17][10] , \sa_ctrl[17].f.spare[5] );
tran (\sa_ctrl[17][11] , \sa_ctrl[17].r.part0[11] );
tran (\sa_ctrl[17][11] , \sa_ctrl[17].f.spare[6] );
tran (\sa_ctrl[17][12] , \sa_ctrl[17].r.part0[12] );
tran (\sa_ctrl[17][12] , \sa_ctrl[17].f.spare[7] );
tran (\sa_ctrl[17][13] , \sa_ctrl[17].r.part0[13] );
tran (\sa_ctrl[17][13] , \sa_ctrl[17].f.spare[8] );
tran (\sa_ctrl[17][14] , \sa_ctrl[17].r.part0[14] );
tran (\sa_ctrl[17][14] , \sa_ctrl[17].f.spare[9] );
tran (\sa_ctrl[17][15] , \sa_ctrl[17].r.part0[15] );
tran (\sa_ctrl[17][15] , \sa_ctrl[17].f.spare[10] );
tran (\sa_ctrl[17][16] , \sa_ctrl[17].r.part0[16] );
tran (\sa_ctrl[17][16] , \sa_ctrl[17].f.spare[11] );
tran (\sa_ctrl[17][17] , \sa_ctrl[17].r.part0[17] );
tran (\sa_ctrl[17][17] , \sa_ctrl[17].f.spare[12] );
tran (\sa_ctrl[17][18] , \sa_ctrl[17].r.part0[18] );
tran (\sa_ctrl[17][18] , \sa_ctrl[17].f.spare[13] );
tran (\sa_ctrl[17][19] , \sa_ctrl[17].r.part0[19] );
tran (\sa_ctrl[17][19] , \sa_ctrl[17].f.spare[14] );
tran (\sa_ctrl[17][20] , \sa_ctrl[17].r.part0[20] );
tran (\sa_ctrl[17][20] , \sa_ctrl[17].f.spare[15] );
tran (\sa_ctrl[17][21] , \sa_ctrl[17].r.part0[21] );
tran (\sa_ctrl[17][21] , \sa_ctrl[17].f.spare[16] );
tran (\sa_ctrl[17][22] , \sa_ctrl[17].r.part0[22] );
tran (\sa_ctrl[17][22] , \sa_ctrl[17].f.spare[17] );
tran (\sa_ctrl[17][23] , \sa_ctrl[17].r.part0[23] );
tran (\sa_ctrl[17][23] , \sa_ctrl[17].f.spare[18] );
tran (\sa_ctrl[17][24] , \sa_ctrl[17].r.part0[24] );
tran (\sa_ctrl[17][24] , \sa_ctrl[17].f.spare[19] );
tran (\sa_ctrl[17][25] , \sa_ctrl[17].r.part0[25] );
tran (\sa_ctrl[17][25] , \sa_ctrl[17].f.spare[20] );
tran (\sa_ctrl[17][26] , \sa_ctrl[17].r.part0[26] );
tran (\sa_ctrl[17][26] , \sa_ctrl[17].f.spare[21] );
tran (\sa_ctrl[17][27] , \sa_ctrl[17].r.part0[27] );
tran (\sa_ctrl[17][27] , \sa_ctrl[17].f.spare[22] );
tran (\sa_ctrl[17][28] , \sa_ctrl[17].r.part0[28] );
tran (\sa_ctrl[17][28] , \sa_ctrl[17].f.spare[23] );
tran (\sa_ctrl[17][29] , \sa_ctrl[17].r.part0[29] );
tran (\sa_ctrl[17][29] , \sa_ctrl[17].f.spare[24] );
tran (\sa_ctrl[17][30] , \sa_ctrl[17].r.part0[30] );
tran (\sa_ctrl[17][30] , \sa_ctrl[17].f.spare[25] );
tran (\sa_ctrl[17][31] , \sa_ctrl[17].r.part0[31] );
tran (\sa_ctrl[17][31] , \sa_ctrl[17].f.spare[26] );
tran (\sa_ctrl[18][0] , \sa_ctrl[18].r.part0[0] );
tran (\sa_ctrl[18][0] , \sa_ctrl[18].f.sa_event_sel[0] );
tran (\sa_ctrl[18][1] , \sa_ctrl[18].r.part0[1] );
tran (\sa_ctrl[18][1] , \sa_ctrl[18].f.sa_event_sel[1] );
tran (\sa_ctrl[18][2] , \sa_ctrl[18].r.part0[2] );
tran (\sa_ctrl[18][2] , \sa_ctrl[18].f.sa_event_sel[2] );
tran (\sa_ctrl[18][3] , \sa_ctrl[18].r.part0[3] );
tran (\sa_ctrl[18][3] , \sa_ctrl[18].f.sa_event_sel[3] );
tran (\sa_ctrl[18][4] , \sa_ctrl[18].r.part0[4] );
tran (\sa_ctrl[18][4] , \sa_ctrl[18].f.sa_event_sel[4] );
tran (\sa_ctrl[18][5] , \sa_ctrl[18].r.part0[5] );
tran (\sa_ctrl[18][5] , \sa_ctrl[18].f.spare[0] );
tran (\sa_ctrl[18][6] , \sa_ctrl[18].r.part0[6] );
tran (\sa_ctrl[18][6] , \sa_ctrl[18].f.spare[1] );
tran (\sa_ctrl[18][7] , \sa_ctrl[18].r.part0[7] );
tran (\sa_ctrl[18][7] , \sa_ctrl[18].f.spare[2] );
tran (\sa_ctrl[18][8] , \sa_ctrl[18].r.part0[8] );
tran (\sa_ctrl[18][8] , \sa_ctrl[18].f.spare[3] );
tran (\sa_ctrl[18][9] , \sa_ctrl[18].r.part0[9] );
tran (\sa_ctrl[18][9] , \sa_ctrl[18].f.spare[4] );
tran (\sa_ctrl[18][10] , \sa_ctrl[18].r.part0[10] );
tran (\sa_ctrl[18][10] , \sa_ctrl[18].f.spare[5] );
tran (\sa_ctrl[18][11] , \sa_ctrl[18].r.part0[11] );
tran (\sa_ctrl[18][11] , \sa_ctrl[18].f.spare[6] );
tran (\sa_ctrl[18][12] , \sa_ctrl[18].r.part0[12] );
tran (\sa_ctrl[18][12] , \sa_ctrl[18].f.spare[7] );
tran (\sa_ctrl[18][13] , \sa_ctrl[18].r.part0[13] );
tran (\sa_ctrl[18][13] , \sa_ctrl[18].f.spare[8] );
tran (\sa_ctrl[18][14] , \sa_ctrl[18].r.part0[14] );
tran (\sa_ctrl[18][14] , \sa_ctrl[18].f.spare[9] );
tran (\sa_ctrl[18][15] , \sa_ctrl[18].r.part0[15] );
tran (\sa_ctrl[18][15] , \sa_ctrl[18].f.spare[10] );
tran (\sa_ctrl[18][16] , \sa_ctrl[18].r.part0[16] );
tran (\sa_ctrl[18][16] , \sa_ctrl[18].f.spare[11] );
tran (\sa_ctrl[18][17] , \sa_ctrl[18].r.part0[17] );
tran (\sa_ctrl[18][17] , \sa_ctrl[18].f.spare[12] );
tran (\sa_ctrl[18][18] , \sa_ctrl[18].r.part0[18] );
tran (\sa_ctrl[18][18] , \sa_ctrl[18].f.spare[13] );
tran (\sa_ctrl[18][19] , \sa_ctrl[18].r.part0[19] );
tran (\sa_ctrl[18][19] , \sa_ctrl[18].f.spare[14] );
tran (\sa_ctrl[18][20] , \sa_ctrl[18].r.part0[20] );
tran (\sa_ctrl[18][20] , \sa_ctrl[18].f.spare[15] );
tran (\sa_ctrl[18][21] , \sa_ctrl[18].r.part0[21] );
tran (\sa_ctrl[18][21] , \sa_ctrl[18].f.spare[16] );
tran (\sa_ctrl[18][22] , \sa_ctrl[18].r.part0[22] );
tran (\sa_ctrl[18][22] , \sa_ctrl[18].f.spare[17] );
tran (\sa_ctrl[18][23] , \sa_ctrl[18].r.part0[23] );
tran (\sa_ctrl[18][23] , \sa_ctrl[18].f.spare[18] );
tran (\sa_ctrl[18][24] , \sa_ctrl[18].r.part0[24] );
tran (\sa_ctrl[18][24] , \sa_ctrl[18].f.spare[19] );
tran (\sa_ctrl[18][25] , \sa_ctrl[18].r.part0[25] );
tran (\sa_ctrl[18][25] , \sa_ctrl[18].f.spare[20] );
tran (\sa_ctrl[18][26] , \sa_ctrl[18].r.part0[26] );
tran (\sa_ctrl[18][26] , \sa_ctrl[18].f.spare[21] );
tran (\sa_ctrl[18][27] , \sa_ctrl[18].r.part0[27] );
tran (\sa_ctrl[18][27] , \sa_ctrl[18].f.spare[22] );
tran (\sa_ctrl[18][28] , \sa_ctrl[18].r.part0[28] );
tran (\sa_ctrl[18][28] , \sa_ctrl[18].f.spare[23] );
tran (\sa_ctrl[18][29] , \sa_ctrl[18].r.part0[29] );
tran (\sa_ctrl[18][29] , \sa_ctrl[18].f.spare[24] );
tran (\sa_ctrl[18][30] , \sa_ctrl[18].r.part0[30] );
tran (\sa_ctrl[18][30] , \sa_ctrl[18].f.spare[25] );
tran (\sa_ctrl[18][31] , \sa_ctrl[18].r.part0[31] );
tran (\sa_ctrl[18][31] , \sa_ctrl[18].f.spare[26] );
tran (\sa_ctrl[19][0] , \sa_ctrl[19].r.part0[0] );
tran (\sa_ctrl[19][0] , \sa_ctrl[19].f.sa_event_sel[0] );
tran (\sa_ctrl[19][1] , \sa_ctrl[19].r.part0[1] );
tran (\sa_ctrl[19][1] , \sa_ctrl[19].f.sa_event_sel[1] );
tran (\sa_ctrl[19][2] , \sa_ctrl[19].r.part0[2] );
tran (\sa_ctrl[19][2] , \sa_ctrl[19].f.sa_event_sel[2] );
tran (\sa_ctrl[19][3] , \sa_ctrl[19].r.part0[3] );
tran (\sa_ctrl[19][3] , \sa_ctrl[19].f.sa_event_sel[3] );
tran (\sa_ctrl[19][4] , \sa_ctrl[19].r.part0[4] );
tran (\sa_ctrl[19][4] , \sa_ctrl[19].f.sa_event_sel[4] );
tran (\sa_ctrl[19][5] , \sa_ctrl[19].r.part0[5] );
tran (\sa_ctrl[19][5] , \sa_ctrl[19].f.spare[0] );
tran (\sa_ctrl[19][6] , \sa_ctrl[19].r.part0[6] );
tran (\sa_ctrl[19][6] , \sa_ctrl[19].f.spare[1] );
tran (\sa_ctrl[19][7] , \sa_ctrl[19].r.part0[7] );
tran (\sa_ctrl[19][7] , \sa_ctrl[19].f.spare[2] );
tran (\sa_ctrl[19][8] , \sa_ctrl[19].r.part0[8] );
tran (\sa_ctrl[19][8] , \sa_ctrl[19].f.spare[3] );
tran (\sa_ctrl[19][9] , \sa_ctrl[19].r.part0[9] );
tran (\sa_ctrl[19][9] , \sa_ctrl[19].f.spare[4] );
tran (\sa_ctrl[19][10] , \sa_ctrl[19].r.part0[10] );
tran (\sa_ctrl[19][10] , \sa_ctrl[19].f.spare[5] );
tran (\sa_ctrl[19][11] , \sa_ctrl[19].r.part0[11] );
tran (\sa_ctrl[19][11] , \sa_ctrl[19].f.spare[6] );
tran (\sa_ctrl[19][12] , \sa_ctrl[19].r.part0[12] );
tran (\sa_ctrl[19][12] , \sa_ctrl[19].f.spare[7] );
tran (\sa_ctrl[19][13] , \sa_ctrl[19].r.part0[13] );
tran (\sa_ctrl[19][13] , \sa_ctrl[19].f.spare[8] );
tran (\sa_ctrl[19][14] , \sa_ctrl[19].r.part0[14] );
tran (\sa_ctrl[19][14] , \sa_ctrl[19].f.spare[9] );
tran (\sa_ctrl[19][15] , \sa_ctrl[19].r.part0[15] );
tran (\sa_ctrl[19][15] , \sa_ctrl[19].f.spare[10] );
tran (\sa_ctrl[19][16] , \sa_ctrl[19].r.part0[16] );
tran (\sa_ctrl[19][16] , \sa_ctrl[19].f.spare[11] );
tran (\sa_ctrl[19][17] , \sa_ctrl[19].r.part0[17] );
tran (\sa_ctrl[19][17] , \sa_ctrl[19].f.spare[12] );
tran (\sa_ctrl[19][18] , \sa_ctrl[19].r.part0[18] );
tran (\sa_ctrl[19][18] , \sa_ctrl[19].f.spare[13] );
tran (\sa_ctrl[19][19] , \sa_ctrl[19].r.part0[19] );
tran (\sa_ctrl[19][19] , \sa_ctrl[19].f.spare[14] );
tran (\sa_ctrl[19][20] , \sa_ctrl[19].r.part0[20] );
tran (\sa_ctrl[19][20] , \sa_ctrl[19].f.spare[15] );
tran (\sa_ctrl[19][21] , \sa_ctrl[19].r.part0[21] );
tran (\sa_ctrl[19][21] , \sa_ctrl[19].f.spare[16] );
tran (\sa_ctrl[19][22] , \sa_ctrl[19].r.part0[22] );
tran (\sa_ctrl[19][22] , \sa_ctrl[19].f.spare[17] );
tran (\sa_ctrl[19][23] , \sa_ctrl[19].r.part0[23] );
tran (\sa_ctrl[19][23] , \sa_ctrl[19].f.spare[18] );
tran (\sa_ctrl[19][24] , \sa_ctrl[19].r.part0[24] );
tran (\sa_ctrl[19][24] , \sa_ctrl[19].f.spare[19] );
tran (\sa_ctrl[19][25] , \sa_ctrl[19].r.part0[25] );
tran (\sa_ctrl[19][25] , \sa_ctrl[19].f.spare[20] );
tran (\sa_ctrl[19][26] , \sa_ctrl[19].r.part0[26] );
tran (\sa_ctrl[19][26] , \sa_ctrl[19].f.spare[21] );
tran (\sa_ctrl[19][27] , \sa_ctrl[19].r.part0[27] );
tran (\sa_ctrl[19][27] , \sa_ctrl[19].f.spare[22] );
tran (\sa_ctrl[19][28] , \sa_ctrl[19].r.part0[28] );
tran (\sa_ctrl[19][28] , \sa_ctrl[19].f.spare[23] );
tran (\sa_ctrl[19][29] , \sa_ctrl[19].r.part0[29] );
tran (\sa_ctrl[19][29] , \sa_ctrl[19].f.spare[24] );
tran (\sa_ctrl[19][30] , \sa_ctrl[19].r.part0[30] );
tran (\sa_ctrl[19][30] , \sa_ctrl[19].f.spare[25] );
tran (\sa_ctrl[19][31] , \sa_ctrl[19].r.part0[31] );
tran (\sa_ctrl[19][31] , \sa_ctrl[19].f.spare[26] );
tran (\sa_ctrl[20][0] , \sa_ctrl[20].r.part0[0] );
tran (\sa_ctrl[20][0] , \sa_ctrl[20].f.sa_event_sel[0] );
tran (\sa_ctrl[20][1] , \sa_ctrl[20].r.part0[1] );
tran (\sa_ctrl[20][1] , \sa_ctrl[20].f.sa_event_sel[1] );
tran (\sa_ctrl[20][2] , \sa_ctrl[20].r.part0[2] );
tran (\sa_ctrl[20][2] , \sa_ctrl[20].f.sa_event_sel[2] );
tran (\sa_ctrl[20][3] , \sa_ctrl[20].r.part0[3] );
tran (\sa_ctrl[20][3] , \sa_ctrl[20].f.sa_event_sel[3] );
tran (\sa_ctrl[20][4] , \sa_ctrl[20].r.part0[4] );
tran (\sa_ctrl[20][4] , \sa_ctrl[20].f.sa_event_sel[4] );
tran (\sa_ctrl[20][5] , \sa_ctrl[20].r.part0[5] );
tran (\sa_ctrl[20][5] , \sa_ctrl[20].f.spare[0] );
tran (\sa_ctrl[20][6] , \sa_ctrl[20].r.part0[6] );
tran (\sa_ctrl[20][6] , \sa_ctrl[20].f.spare[1] );
tran (\sa_ctrl[20][7] , \sa_ctrl[20].r.part0[7] );
tran (\sa_ctrl[20][7] , \sa_ctrl[20].f.spare[2] );
tran (\sa_ctrl[20][8] , \sa_ctrl[20].r.part0[8] );
tran (\sa_ctrl[20][8] , \sa_ctrl[20].f.spare[3] );
tran (\sa_ctrl[20][9] , \sa_ctrl[20].r.part0[9] );
tran (\sa_ctrl[20][9] , \sa_ctrl[20].f.spare[4] );
tran (\sa_ctrl[20][10] , \sa_ctrl[20].r.part0[10] );
tran (\sa_ctrl[20][10] , \sa_ctrl[20].f.spare[5] );
tran (\sa_ctrl[20][11] , \sa_ctrl[20].r.part0[11] );
tran (\sa_ctrl[20][11] , \sa_ctrl[20].f.spare[6] );
tran (\sa_ctrl[20][12] , \sa_ctrl[20].r.part0[12] );
tran (\sa_ctrl[20][12] , \sa_ctrl[20].f.spare[7] );
tran (\sa_ctrl[20][13] , \sa_ctrl[20].r.part0[13] );
tran (\sa_ctrl[20][13] , \sa_ctrl[20].f.spare[8] );
tran (\sa_ctrl[20][14] , \sa_ctrl[20].r.part0[14] );
tran (\sa_ctrl[20][14] , \sa_ctrl[20].f.spare[9] );
tran (\sa_ctrl[20][15] , \sa_ctrl[20].r.part0[15] );
tran (\sa_ctrl[20][15] , \sa_ctrl[20].f.spare[10] );
tran (\sa_ctrl[20][16] , \sa_ctrl[20].r.part0[16] );
tran (\sa_ctrl[20][16] , \sa_ctrl[20].f.spare[11] );
tran (\sa_ctrl[20][17] , \sa_ctrl[20].r.part0[17] );
tran (\sa_ctrl[20][17] , \sa_ctrl[20].f.spare[12] );
tran (\sa_ctrl[20][18] , \sa_ctrl[20].r.part0[18] );
tran (\sa_ctrl[20][18] , \sa_ctrl[20].f.spare[13] );
tran (\sa_ctrl[20][19] , \sa_ctrl[20].r.part0[19] );
tran (\sa_ctrl[20][19] , \sa_ctrl[20].f.spare[14] );
tran (\sa_ctrl[20][20] , \sa_ctrl[20].r.part0[20] );
tran (\sa_ctrl[20][20] , \sa_ctrl[20].f.spare[15] );
tran (\sa_ctrl[20][21] , \sa_ctrl[20].r.part0[21] );
tran (\sa_ctrl[20][21] , \sa_ctrl[20].f.spare[16] );
tran (\sa_ctrl[20][22] , \sa_ctrl[20].r.part0[22] );
tran (\sa_ctrl[20][22] , \sa_ctrl[20].f.spare[17] );
tran (\sa_ctrl[20][23] , \sa_ctrl[20].r.part0[23] );
tran (\sa_ctrl[20][23] , \sa_ctrl[20].f.spare[18] );
tran (\sa_ctrl[20][24] , \sa_ctrl[20].r.part0[24] );
tran (\sa_ctrl[20][24] , \sa_ctrl[20].f.spare[19] );
tran (\sa_ctrl[20][25] , \sa_ctrl[20].r.part0[25] );
tran (\sa_ctrl[20][25] , \sa_ctrl[20].f.spare[20] );
tran (\sa_ctrl[20][26] , \sa_ctrl[20].r.part0[26] );
tran (\sa_ctrl[20][26] , \sa_ctrl[20].f.spare[21] );
tran (\sa_ctrl[20][27] , \sa_ctrl[20].r.part0[27] );
tran (\sa_ctrl[20][27] , \sa_ctrl[20].f.spare[22] );
tran (\sa_ctrl[20][28] , \sa_ctrl[20].r.part0[28] );
tran (\sa_ctrl[20][28] , \sa_ctrl[20].f.spare[23] );
tran (\sa_ctrl[20][29] , \sa_ctrl[20].r.part0[29] );
tran (\sa_ctrl[20][29] , \sa_ctrl[20].f.spare[24] );
tran (\sa_ctrl[20][30] , \sa_ctrl[20].r.part0[30] );
tran (\sa_ctrl[20][30] , \sa_ctrl[20].f.spare[25] );
tran (\sa_ctrl[20][31] , \sa_ctrl[20].r.part0[31] );
tran (\sa_ctrl[20][31] , \sa_ctrl[20].f.spare[26] );
tran (\sa_ctrl[21][0] , \sa_ctrl[21].r.part0[0] );
tran (\sa_ctrl[21][0] , \sa_ctrl[21].f.sa_event_sel[0] );
tran (\sa_ctrl[21][1] , \sa_ctrl[21].r.part0[1] );
tran (\sa_ctrl[21][1] , \sa_ctrl[21].f.sa_event_sel[1] );
tran (\sa_ctrl[21][2] , \sa_ctrl[21].r.part0[2] );
tran (\sa_ctrl[21][2] , \sa_ctrl[21].f.sa_event_sel[2] );
tran (\sa_ctrl[21][3] , \sa_ctrl[21].r.part0[3] );
tran (\sa_ctrl[21][3] , \sa_ctrl[21].f.sa_event_sel[3] );
tran (\sa_ctrl[21][4] , \sa_ctrl[21].r.part0[4] );
tran (\sa_ctrl[21][4] , \sa_ctrl[21].f.sa_event_sel[4] );
tran (\sa_ctrl[21][5] , \sa_ctrl[21].r.part0[5] );
tran (\sa_ctrl[21][5] , \sa_ctrl[21].f.spare[0] );
tran (\sa_ctrl[21][6] , \sa_ctrl[21].r.part0[6] );
tran (\sa_ctrl[21][6] , \sa_ctrl[21].f.spare[1] );
tran (\sa_ctrl[21][7] , \sa_ctrl[21].r.part0[7] );
tran (\sa_ctrl[21][7] , \sa_ctrl[21].f.spare[2] );
tran (\sa_ctrl[21][8] , \sa_ctrl[21].r.part0[8] );
tran (\sa_ctrl[21][8] , \sa_ctrl[21].f.spare[3] );
tran (\sa_ctrl[21][9] , \sa_ctrl[21].r.part0[9] );
tran (\sa_ctrl[21][9] , \sa_ctrl[21].f.spare[4] );
tran (\sa_ctrl[21][10] , \sa_ctrl[21].r.part0[10] );
tran (\sa_ctrl[21][10] , \sa_ctrl[21].f.spare[5] );
tran (\sa_ctrl[21][11] , \sa_ctrl[21].r.part0[11] );
tran (\sa_ctrl[21][11] , \sa_ctrl[21].f.spare[6] );
tran (\sa_ctrl[21][12] , \sa_ctrl[21].r.part0[12] );
tran (\sa_ctrl[21][12] , \sa_ctrl[21].f.spare[7] );
tran (\sa_ctrl[21][13] , \sa_ctrl[21].r.part0[13] );
tran (\sa_ctrl[21][13] , \sa_ctrl[21].f.spare[8] );
tran (\sa_ctrl[21][14] , \sa_ctrl[21].r.part0[14] );
tran (\sa_ctrl[21][14] , \sa_ctrl[21].f.spare[9] );
tran (\sa_ctrl[21][15] , \sa_ctrl[21].r.part0[15] );
tran (\sa_ctrl[21][15] , \sa_ctrl[21].f.spare[10] );
tran (\sa_ctrl[21][16] , \sa_ctrl[21].r.part0[16] );
tran (\sa_ctrl[21][16] , \sa_ctrl[21].f.spare[11] );
tran (\sa_ctrl[21][17] , \sa_ctrl[21].r.part0[17] );
tran (\sa_ctrl[21][17] , \sa_ctrl[21].f.spare[12] );
tran (\sa_ctrl[21][18] , \sa_ctrl[21].r.part0[18] );
tran (\sa_ctrl[21][18] , \sa_ctrl[21].f.spare[13] );
tran (\sa_ctrl[21][19] , \sa_ctrl[21].r.part0[19] );
tran (\sa_ctrl[21][19] , \sa_ctrl[21].f.spare[14] );
tran (\sa_ctrl[21][20] , \sa_ctrl[21].r.part0[20] );
tran (\sa_ctrl[21][20] , \sa_ctrl[21].f.spare[15] );
tran (\sa_ctrl[21][21] , \sa_ctrl[21].r.part0[21] );
tran (\sa_ctrl[21][21] , \sa_ctrl[21].f.spare[16] );
tran (\sa_ctrl[21][22] , \sa_ctrl[21].r.part0[22] );
tran (\sa_ctrl[21][22] , \sa_ctrl[21].f.spare[17] );
tran (\sa_ctrl[21][23] , \sa_ctrl[21].r.part0[23] );
tran (\sa_ctrl[21][23] , \sa_ctrl[21].f.spare[18] );
tran (\sa_ctrl[21][24] , \sa_ctrl[21].r.part0[24] );
tran (\sa_ctrl[21][24] , \sa_ctrl[21].f.spare[19] );
tran (\sa_ctrl[21][25] , \sa_ctrl[21].r.part0[25] );
tran (\sa_ctrl[21][25] , \sa_ctrl[21].f.spare[20] );
tran (\sa_ctrl[21][26] , \sa_ctrl[21].r.part0[26] );
tran (\sa_ctrl[21][26] , \sa_ctrl[21].f.spare[21] );
tran (\sa_ctrl[21][27] , \sa_ctrl[21].r.part0[27] );
tran (\sa_ctrl[21][27] , \sa_ctrl[21].f.spare[22] );
tran (\sa_ctrl[21][28] , \sa_ctrl[21].r.part0[28] );
tran (\sa_ctrl[21][28] , \sa_ctrl[21].f.spare[23] );
tran (\sa_ctrl[21][29] , \sa_ctrl[21].r.part0[29] );
tran (\sa_ctrl[21][29] , \sa_ctrl[21].f.spare[24] );
tran (\sa_ctrl[21][30] , \sa_ctrl[21].r.part0[30] );
tran (\sa_ctrl[21][30] , \sa_ctrl[21].f.spare[25] );
tran (\sa_ctrl[21][31] , \sa_ctrl[21].r.part0[31] );
tran (\sa_ctrl[21][31] , \sa_ctrl[21].f.spare[26] );
tran (\sa_ctrl[22][0] , \sa_ctrl[22].r.part0[0] );
tran (\sa_ctrl[22][0] , \sa_ctrl[22].f.sa_event_sel[0] );
tran (\sa_ctrl[22][1] , \sa_ctrl[22].r.part0[1] );
tran (\sa_ctrl[22][1] , \sa_ctrl[22].f.sa_event_sel[1] );
tran (\sa_ctrl[22][2] , \sa_ctrl[22].r.part0[2] );
tran (\sa_ctrl[22][2] , \sa_ctrl[22].f.sa_event_sel[2] );
tran (\sa_ctrl[22][3] , \sa_ctrl[22].r.part0[3] );
tran (\sa_ctrl[22][3] , \sa_ctrl[22].f.sa_event_sel[3] );
tran (\sa_ctrl[22][4] , \sa_ctrl[22].r.part0[4] );
tran (\sa_ctrl[22][4] , \sa_ctrl[22].f.sa_event_sel[4] );
tran (\sa_ctrl[22][5] , \sa_ctrl[22].r.part0[5] );
tran (\sa_ctrl[22][5] , \sa_ctrl[22].f.spare[0] );
tran (\sa_ctrl[22][6] , \sa_ctrl[22].r.part0[6] );
tran (\sa_ctrl[22][6] , \sa_ctrl[22].f.spare[1] );
tran (\sa_ctrl[22][7] , \sa_ctrl[22].r.part0[7] );
tran (\sa_ctrl[22][7] , \sa_ctrl[22].f.spare[2] );
tran (\sa_ctrl[22][8] , \sa_ctrl[22].r.part0[8] );
tran (\sa_ctrl[22][8] , \sa_ctrl[22].f.spare[3] );
tran (\sa_ctrl[22][9] , \sa_ctrl[22].r.part0[9] );
tran (\sa_ctrl[22][9] , \sa_ctrl[22].f.spare[4] );
tran (\sa_ctrl[22][10] , \sa_ctrl[22].r.part0[10] );
tran (\sa_ctrl[22][10] , \sa_ctrl[22].f.spare[5] );
tran (\sa_ctrl[22][11] , \sa_ctrl[22].r.part0[11] );
tran (\sa_ctrl[22][11] , \sa_ctrl[22].f.spare[6] );
tran (\sa_ctrl[22][12] , \sa_ctrl[22].r.part0[12] );
tran (\sa_ctrl[22][12] , \sa_ctrl[22].f.spare[7] );
tran (\sa_ctrl[22][13] , \sa_ctrl[22].r.part0[13] );
tran (\sa_ctrl[22][13] , \sa_ctrl[22].f.spare[8] );
tran (\sa_ctrl[22][14] , \sa_ctrl[22].r.part0[14] );
tran (\sa_ctrl[22][14] , \sa_ctrl[22].f.spare[9] );
tran (\sa_ctrl[22][15] , \sa_ctrl[22].r.part0[15] );
tran (\sa_ctrl[22][15] , \sa_ctrl[22].f.spare[10] );
tran (\sa_ctrl[22][16] , \sa_ctrl[22].r.part0[16] );
tran (\sa_ctrl[22][16] , \sa_ctrl[22].f.spare[11] );
tran (\sa_ctrl[22][17] , \sa_ctrl[22].r.part0[17] );
tran (\sa_ctrl[22][17] , \sa_ctrl[22].f.spare[12] );
tran (\sa_ctrl[22][18] , \sa_ctrl[22].r.part0[18] );
tran (\sa_ctrl[22][18] , \sa_ctrl[22].f.spare[13] );
tran (\sa_ctrl[22][19] , \sa_ctrl[22].r.part0[19] );
tran (\sa_ctrl[22][19] , \sa_ctrl[22].f.spare[14] );
tran (\sa_ctrl[22][20] , \sa_ctrl[22].r.part0[20] );
tran (\sa_ctrl[22][20] , \sa_ctrl[22].f.spare[15] );
tran (\sa_ctrl[22][21] , \sa_ctrl[22].r.part0[21] );
tran (\sa_ctrl[22][21] , \sa_ctrl[22].f.spare[16] );
tran (\sa_ctrl[22][22] , \sa_ctrl[22].r.part0[22] );
tran (\sa_ctrl[22][22] , \sa_ctrl[22].f.spare[17] );
tran (\sa_ctrl[22][23] , \sa_ctrl[22].r.part0[23] );
tran (\sa_ctrl[22][23] , \sa_ctrl[22].f.spare[18] );
tran (\sa_ctrl[22][24] , \sa_ctrl[22].r.part0[24] );
tran (\sa_ctrl[22][24] , \sa_ctrl[22].f.spare[19] );
tran (\sa_ctrl[22][25] , \sa_ctrl[22].r.part0[25] );
tran (\sa_ctrl[22][25] , \sa_ctrl[22].f.spare[20] );
tran (\sa_ctrl[22][26] , \sa_ctrl[22].r.part0[26] );
tran (\sa_ctrl[22][26] , \sa_ctrl[22].f.spare[21] );
tran (\sa_ctrl[22][27] , \sa_ctrl[22].r.part0[27] );
tran (\sa_ctrl[22][27] , \sa_ctrl[22].f.spare[22] );
tran (\sa_ctrl[22][28] , \sa_ctrl[22].r.part0[28] );
tran (\sa_ctrl[22][28] , \sa_ctrl[22].f.spare[23] );
tran (\sa_ctrl[22][29] , \sa_ctrl[22].r.part0[29] );
tran (\sa_ctrl[22][29] , \sa_ctrl[22].f.spare[24] );
tran (\sa_ctrl[22][30] , \sa_ctrl[22].r.part0[30] );
tran (\sa_ctrl[22][30] , \sa_ctrl[22].f.spare[25] );
tran (\sa_ctrl[22][31] , \sa_ctrl[22].r.part0[31] );
tran (\sa_ctrl[22][31] , \sa_ctrl[22].f.spare[26] );
tran (\sa_ctrl[23][0] , \sa_ctrl[23].r.part0[0] );
tran (\sa_ctrl[23][0] , \sa_ctrl[23].f.sa_event_sel[0] );
tran (\sa_ctrl[23][1] , \sa_ctrl[23].r.part0[1] );
tran (\sa_ctrl[23][1] , \sa_ctrl[23].f.sa_event_sel[1] );
tran (\sa_ctrl[23][2] , \sa_ctrl[23].r.part0[2] );
tran (\sa_ctrl[23][2] , \sa_ctrl[23].f.sa_event_sel[2] );
tran (\sa_ctrl[23][3] , \sa_ctrl[23].r.part0[3] );
tran (\sa_ctrl[23][3] , \sa_ctrl[23].f.sa_event_sel[3] );
tran (\sa_ctrl[23][4] , \sa_ctrl[23].r.part0[4] );
tran (\sa_ctrl[23][4] , \sa_ctrl[23].f.sa_event_sel[4] );
tran (\sa_ctrl[23][5] , \sa_ctrl[23].r.part0[5] );
tran (\sa_ctrl[23][5] , \sa_ctrl[23].f.spare[0] );
tran (\sa_ctrl[23][6] , \sa_ctrl[23].r.part0[6] );
tran (\sa_ctrl[23][6] , \sa_ctrl[23].f.spare[1] );
tran (\sa_ctrl[23][7] , \sa_ctrl[23].r.part0[7] );
tran (\sa_ctrl[23][7] , \sa_ctrl[23].f.spare[2] );
tran (\sa_ctrl[23][8] , \sa_ctrl[23].r.part0[8] );
tran (\sa_ctrl[23][8] , \sa_ctrl[23].f.spare[3] );
tran (\sa_ctrl[23][9] , \sa_ctrl[23].r.part0[9] );
tran (\sa_ctrl[23][9] , \sa_ctrl[23].f.spare[4] );
tran (\sa_ctrl[23][10] , \sa_ctrl[23].r.part0[10] );
tran (\sa_ctrl[23][10] , \sa_ctrl[23].f.spare[5] );
tran (\sa_ctrl[23][11] , \sa_ctrl[23].r.part0[11] );
tran (\sa_ctrl[23][11] , \sa_ctrl[23].f.spare[6] );
tran (\sa_ctrl[23][12] , \sa_ctrl[23].r.part0[12] );
tran (\sa_ctrl[23][12] , \sa_ctrl[23].f.spare[7] );
tran (\sa_ctrl[23][13] , \sa_ctrl[23].r.part0[13] );
tran (\sa_ctrl[23][13] , \sa_ctrl[23].f.spare[8] );
tran (\sa_ctrl[23][14] , \sa_ctrl[23].r.part0[14] );
tran (\sa_ctrl[23][14] , \sa_ctrl[23].f.spare[9] );
tran (\sa_ctrl[23][15] , \sa_ctrl[23].r.part0[15] );
tran (\sa_ctrl[23][15] , \sa_ctrl[23].f.spare[10] );
tran (\sa_ctrl[23][16] , \sa_ctrl[23].r.part0[16] );
tran (\sa_ctrl[23][16] , \sa_ctrl[23].f.spare[11] );
tran (\sa_ctrl[23][17] , \sa_ctrl[23].r.part0[17] );
tran (\sa_ctrl[23][17] , \sa_ctrl[23].f.spare[12] );
tran (\sa_ctrl[23][18] , \sa_ctrl[23].r.part0[18] );
tran (\sa_ctrl[23][18] , \sa_ctrl[23].f.spare[13] );
tran (\sa_ctrl[23][19] , \sa_ctrl[23].r.part0[19] );
tran (\sa_ctrl[23][19] , \sa_ctrl[23].f.spare[14] );
tran (\sa_ctrl[23][20] , \sa_ctrl[23].r.part0[20] );
tran (\sa_ctrl[23][20] , \sa_ctrl[23].f.spare[15] );
tran (\sa_ctrl[23][21] , \sa_ctrl[23].r.part0[21] );
tran (\sa_ctrl[23][21] , \sa_ctrl[23].f.spare[16] );
tran (\sa_ctrl[23][22] , \sa_ctrl[23].r.part0[22] );
tran (\sa_ctrl[23][22] , \sa_ctrl[23].f.spare[17] );
tran (\sa_ctrl[23][23] , \sa_ctrl[23].r.part0[23] );
tran (\sa_ctrl[23][23] , \sa_ctrl[23].f.spare[18] );
tran (\sa_ctrl[23][24] , \sa_ctrl[23].r.part0[24] );
tran (\sa_ctrl[23][24] , \sa_ctrl[23].f.spare[19] );
tran (\sa_ctrl[23][25] , \sa_ctrl[23].r.part0[25] );
tran (\sa_ctrl[23][25] , \sa_ctrl[23].f.spare[20] );
tran (\sa_ctrl[23][26] , \sa_ctrl[23].r.part0[26] );
tran (\sa_ctrl[23][26] , \sa_ctrl[23].f.spare[21] );
tran (\sa_ctrl[23][27] , \sa_ctrl[23].r.part0[27] );
tran (\sa_ctrl[23][27] , \sa_ctrl[23].f.spare[22] );
tran (\sa_ctrl[23][28] , \sa_ctrl[23].r.part0[28] );
tran (\sa_ctrl[23][28] , \sa_ctrl[23].f.spare[23] );
tran (\sa_ctrl[23][29] , \sa_ctrl[23].r.part0[29] );
tran (\sa_ctrl[23][29] , \sa_ctrl[23].f.spare[24] );
tran (\sa_ctrl[23][30] , \sa_ctrl[23].r.part0[30] );
tran (\sa_ctrl[23][30] , \sa_ctrl[23].f.spare[25] );
tran (\sa_ctrl[23][31] , \sa_ctrl[23].r.part0[31] );
tran (\sa_ctrl[23][31] , \sa_ctrl[23].f.spare[26] );
tran (\sa_ctrl[24][0] , \sa_ctrl[24].r.part0[0] );
tran (\sa_ctrl[24][0] , \sa_ctrl[24].f.sa_event_sel[0] );
tran (\sa_ctrl[24][1] , \sa_ctrl[24].r.part0[1] );
tran (\sa_ctrl[24][1] , \sa_ctrl[24].f.sa_event_sel[1] );
tran (\sa_ctrl[24][2] , \sa_ctrl[24].r.part0[2] );
tran (\sa_ctrl[24][2] , \sa_ctrl[24].f.sa_event_sel[2] );
tran (\sa_ctrl[24][3] , \sa_ctrl[24].r.part0[3] );
tran (\sa_ctrl[24][3] , \sa_ctrl[24].f.sa_event_sel[3] );
tran (\sa_ctrl[24][4] , \sa_ctrl[24].r.part0[4] );
tran (\sa_ctrl[24][4] , \sa_ctrl[24].f.sa_event_sel[4] );
tran (\sa_ctrl[24][5] , \sa_ctrl[24].r.part0[5] );
tran (\sa_ctrl[24][5] , \sa_ctrl[24].f.spare[0] );
tran (\sa_ctrl[24][6] , \sa_ctrl[24].r.part0[6] );
tran (\sa_ctrl[24][6] , \sa_ctrl[24].f.spare[1] );
tran (\sa_ctrl[24][7] , \sa_ctrl[24].r.part0[7] );
tran (\sa_ctrl[24][7] , \sa_ctrl[24].f.spare[2] );
tran (\sa_ctrl[24][8] , \sa_ctrl[24].r.part0[8] );
tran (\sa_ctrl[24][8] , \sa_ctrl[24].f.spare[3] );
tran (\sa_ctrl[24][9] , \sa_ctrl[24].r.part0[9] );
tran (\sa_ctrl[24][9] , \sa_ctrl[24].f.spare[4] );
tran (\sa_ctrl[24][10] , \sa_ctrl[24].r.part0[10] );
tran (\sa_ctrl[24][10] , \sa_ctrl[24].f.spare[5] );
tran (\sa_ctrl[24][11] , \sa_ctrl[24].r.part0[11] );
tran (\sa_ctrl[24][11] , \sa_ctrl[24].f.spare[6] );
tran (\sa_ctrl[24][12] , \sa_ctrl[24].r.part0[12] );
tran (\sa_ctrl[24][12] , \sa_ctrl[24].f.spare[7] );
tran (\sa_ctrl[24][13] , \sa_ctrl[24].r.part0[13] );
tran (\sa_ctrl[24][13] , \sa_ctrl[24].f.spare[8] );
tran (\sa_ctrl[24][14] , \sa_ctrl[24].r.part0[14] );
tran (\sa_ctrl[24][14] , \sa_ctrl[24].f.spare[9] );
tran (\sa_ctrl[24][15] , \sa_ctrl[24].r.part0[15] );
tran (\sa_ctrl[24][15] , \sa_ctrl[24].f.spare[10] );
tran (\sa_ctrl[24][16] , \sa_ctrl[24].r.part0[16] );
tran (\sa_ctrl[24][16] , \sa_ctrl[24].f.spare[11] );
tran (\sa_ctrl[24][17] , \sa_ctrl[24].r.part0[17] );
tran (\sa_ctrl[24][17] , \sa_ctrl[24].f.spare[12] );
tran (\sa_ctrl[24][18] , \sa_ctrl[24].r.part0[18] );
tran (\sa_ctrl[24][18] , \sa_ctrl[24].f.spare[13] );
tran (\sa_ctrl[24][19] , \sa_ctrl[24].r.part0[19] );
tran (\sa_ctrl[24][19] , \sa_ctrl[24].f.spare[14] );
tran (\sa_ctrl[24][20] , \sa_ctrl[24].r.part0[20] );
tran (\sa_ctrl[24][20] , \sa_ctrl[24].f.spare[15] );
tran (\sa_ctrl[24][21] , \sa_ctrl[24].r.part0[21] );
tran (\sa_ctrl[24][21] , \sa_ctrl[24].f.spare[16] );
tran (\sa_ctrl[24][22] , \sa_ctrl[24].r.part0[22] );
tran (\sa_ctrl[24][22] , \sa_ctrl[24].f.spare[17] );
tran (\sa_ctrl[24][23] , \sa_ctrl[24].r.part0[23] );
tran (\sa_ctrl[24][23] , \sa_ctrl[24].f.spare[18] );
tran (\sa_ctrl[24][24] , \sa_ctrl[24].r.part0[24] );
tran (\sa_ctrl[24][24] , \sa_ctrl[24].f.spare[19] );
tran (\sa_ctrl[24][25] , \sa_ctrl[24].r.part0[25] );
tran (\sa_ctrl[24][25] , \sa_ctrl[24].f.spare[20] );
tran (\sa_ctrl[24][26] , \sa_ctrl[24].r.part0[26] );
tran (\sa_ctrl[24][26] , \sa_ctrl[24].f.spare[21] );
tran (\sa_ctrl[24][27] , \sa_ctrl[24].r.part0[27] );
tran (\sa_ctrl[24][27] , \sa_ctrl[24].f.spare[22] );
tran (\sa_ctrl[24][28] , \sa_ctrl[24].r.part0[28] );
tran (\sa_ctrl[24][28] , \sa_ctrl[24].f.spare[23] );
tran (\sa_ctrl[24][29] , \sa_ctrl[24].r.part0[29] );
tran (\sa_ctrl[24][29] , \sa_ctrl[24].f.spare[24] );
tran (\sa_ctrl[24][30] , \sa_ctrl[24].r.part0[30] );
tran (\sa_ctrl[24][30] , \sa_ctrl[24].f.spare[25] );
tran (\sa_ctrl[24][31] , \sa_ctrl[24].r.part0[31] );
tran (\sa_ctrl[24][31] , \sa_ctrl[24].f.spare[26] );
tran (\sa_ctrl[25][0] , \sa_ctrl[25].r.part0[0] );
tran (\sa_ctrl[25][0] , \sa_ctrl[25].f.sa_event_sel[0] );
tran (\sa_ctrl[25][1] , \sa_ctrl[25].r.part0[1] );
tran (\sa_ctrl[25][1] , \sa_ctrl[25].f.sa_event_sel[1] );
tran (\sa_ctrl[25][2] , \sa_ctrl[25].r.part0[2] );
tran (\sa_ctrl[25][2] , \sa_ctrl[25].f.sa_event_sel[2] );
tran (\sa_ctrl[25][3] , \sa_ctrl[25].r.part0[3] );
tran (\sa_ctrl[25][3] , \sa_ctrl[25].f.sa_event_sel[3] );
tran (\sa_ctrl[25][4] , \sa_ctrl[25].r.part0[4] );
tran (\sa_ctrl[25][4] , \sa_ctrl[25].f.sa_event_sel[4] );
tran (\sa_ctrl[25][5] , \sa_ctrl[25].r.part0[5] );
tran (\sa_ctrl[25][5] , \sa_ctrl[25].f.spare[0] );
tran (\sa_ctrl[25][6] , \sa_ctrl[25].r.part0[6] );
tran (\sa_ctrl[25][6] , \sa_ctrl[25].f.spare[1] );
tran (\sa_ctrl[25][7] , \sa_ctrl[25].r.part0[7] );
tran (\sa_ctrl[25][7] , \sa_ctrl[25].f.spare[2] );
tran (\sa_ctrl[25][8] , \sa_ctrl[25].r.part0[8] );
tran (\sa_ctrl[25][8] , \sa_ctrl[25].f.spare[3] );
tran (\sa_ctrl[25][9] , \sa_ctrl[25].r.part0[9] );
tran (\sa_ctrl[25][9] , \sa_ctrl[25].f.spare[4] );
tran (\sa_ctrl[25][10] , \sa_ctrl[25].r.part0[10] );
tran (\sa_ctrl[25][10] , \sa_ctrl[25].f.spare[5] );
tran (\sa_ctrl[25][11] , \sa_ctrl[25].r.part0[11] );
tran (\sa_ctrl[25][11] , \sa_ctrl[25].f.spare[6] );
tran (\sa_ctrl[25][12] , \sa_ctrl[25].r.part0[12] );
tran (\sa_ctrl[25][12] , \sa_ctrl[25].f.spare[7] );
tran (\sa_ctrl[25][13] , \sa_ctrl[25].r.part0[13] );
tran (\sa_ctrl[25][13] , \sa_ctrl[25].f.spare[8] );
tran (\sa_ctrl[25][14] , \sa_ctrl[25].r.part0[14] );
tran (\sa_ctrl[25][14] , \sa_ctrl[25].f.spare[9] );
tran (\sa_ctrl[25][15] , \sa_ctrl[25].r.part0[15] );
tran (\sa_ctrl[25][15] , \sa_ctrl[25].f.spare[10] );
tran (\sa_ctrl[25][16] , \sa_ctrl[25].r.part0[16] );
tran (\sa_ctrl[25][16] , \sa_ctrl[25].f.spare[11] );
tran (\sa_ctrl[25][17] , \sa_ctrl[25].r.part0[17] );
tran (\sa_ctrl[25][17] , \sa_ctrl[25].f.spare[12] );
tran (\sa_ctrl[25][18] , \sa_ctrl[25].r.part0[18] );
tran (\sa_ctrl[25][18] , \sa_ctrl[25].f.spare[13] );
tran (\sa_ctrl[25][19] , \sa_ctrl[25].r.part0[19] );
tran (\sa_ctrl[25][19] , \sa_ctrl[25].f.spare[14] );
tran (\sa_ctrl[25][20] , \sa_ctrl[25].r.part0[20] );
tran (\sa_ctrl[25][20] , \sa_ctrl[25].f.spare[15] );
tran (\sa_ctrl[25][21] , \sa_ctrl[25].r.part0[21] );
tran (\sa_ctrl[25][21] , \sa_ctrl[25].f.spare[16] );
tran (\sa_ctrl[25][22] , \sa_ctrl[25].r.part0[22] );
tran (\sa_ctrl[25][22] , \sa_ctrl[25].f.spare[17] );
tran (\sa_ctrl[25][23] , \sa_ctrl[25].r.part0[23] );
tran (\sa_ctrl[25][23] , \sa_ctrl[25].f.spare[18] );
tran (\sa_ctrl[25][24] , \sa_ctrl[25].r.part0[24] );
tran (\sa_ctrl[25][24] , \sa_ctrl[25].f.spare[19] );
tran (\sa_ctrl[25][25] , \sa_ctrl[25].r.part0[25] );
tran (\sa_ctrl[25][25] , \sa_ctrl[25].f.spare[20] );
tran (\sa_ctrl[25][26] , \sa_ctrl[25].r.part0[26] );
tran (\sa_ctrl[25][26] , \sa_ctrl[25].f.spare[21] );
tran (\sa_ctrl[25][27] , \sa_ctrl[25].r.part0[27] );
tran (\sa_ctrl[25][27] , \sa_ctrl[25].f.spare[22] );
tran (\sa_ctrl[25][28] , \sa_ctrl[25].r.part0[28] );
tran (\sa_ctrl[25][28] , \sa_ctrl[25].f.spare[23] );
tran (\sa_ctrl[25][29] , \sa_ctrl[25].r.part0[29] );
tran (\sa_ctrl[25][29] , \sa_ctrl[25].f.spare[24] );
tran (\sa_ctrl[25][30] , \sa_ctrl[25].r.part0[30] );
tran (\sa_ctrl[25][30] , \sa_ctrl[25].f.spare[25] );
tran (\sa_ctrl[25][31] , \sa_ctrl[25].r.part0[31] );
tran (\sa_ctrl[25][31] , \sa_ctrl[25].f.spare[26] );
tran (\sa_ctrl[26][0] , \sa_ctrl[26].r.part0[0] );
tran (\sa_ctrl[26][0] , \sa_ctrl[26].f.sa_event_sel[0] );
tran (\sa_ctrl[26][1] , \sa_ctrl[26].r.part0[1] );
tran (\sa_ctrl[26][1] , \sa_ctrl[26].f.sa_event_sel[1] );
tran (\sa_ctrl[26][2] , \sa_ctrl[26].r.part0[2] );
tran (\sa_ctrl[26][2] , \sa_ctrl[26].f.sa_event_sel[2] );
tran (\sa_ctrl[26][3] , \sa_ctrl[26].r.part0[3] );
tran (\sa_ctrl[26][3] , \sa_ctrl[26].f.sa_event_sel[3] );
tran (\sa_ctrl[26][4] , \sa_ctrl[26].r.part0[4] );
tran (\sa_ctrl[26][4] , \sa_ctrl[26].f.sa_event_sel[4] );
tran (\sa_ctrl[26][5] , \sa_ctrl[26].r.part0[5] );
tran (\sa_ctrl[26][5] , \sa_ctrl[26].f.spare[0] );
tran (\sa_ctrl[26][6] , \sa_ctrl[26].r.part0[6] );
tran (\sa_ctrl[26][6] , \sa_ctrl[26].f.spare[1] );
tran (\sa_ctrl[26][7] , \sa_ctrl[26].r.part0[7] );
tran (\sa_ctrl[26][7] , \sa_ctrl[26].f.spare[2] );
tran (\sa_ctrl[26][8] , \sa_ctrl[26].r.part0[8] );
tran (\sa_ctrl[26][8] , \sa_ctrl[26].f.spare[3] );
tran (\sa_ctrl[26][9] , \sa_ctrl[26].r.part0[9] );
tran (\sa_ctrl[26][9] , \sa_ctrl[26].f.spare[4] );
tran (\sa_ctrl[26][10] , \sa_ctrl[26].r.part0[10] );
tran (\sa_ctrl[26][10] , \sa_ctrl[26].f.spare[5] );
tran (\sa_ctrl[26][11] , \sa_ctrl[26].r.part0[11] );
tran (\sa_ctrl[26][11] , \sa_ctrl[26].f.spare[6] );
tran (\sa_ctrl[26][12] , \sa_ctrl[26].r.part0[12] );
tran (\sa_ctrl[26][12] , \sa_ctrl[26].f.spare[7] );
tran (\sa_ctrl[26][13] , \sa_ctrl[26].r.part0[13] );
tran (\sa_ctrl[26][13] , \sa_ctrl[26].f.spare[8] );
tran (\sa_ctrl[26][14] , \sa_ctrl[26].r.part0[14] );
tran (\sa_ctrl[26][14] , \sa_ctrl[26].f.spare[9] );
tran (\sa_ctrl[26][15] , \sa_ctrl[26].r.part0[15] );
tran (\sa_ctrl[26][15] , \sa_ctrl[26].f.spare[10] );
tran (\sa_ctrl[26][16] , \sa_ctrl[26].r.part0[16] );
tran (\sa_ctrl[26][16] , \sa_ctrl[26].f.spare[11] );
tran (\sa_ctrl[26][17] , \sa_ctrl[26].r.part0[17] );
tran (\sa_ctrl[26][17] , \sa_ctrl[26].f.spare[12] );
tran (\sa_ctrl[26][18] , \sa_ctrl[26].r.part0[18] );
tran (\sa_ctrl[26][18] , \sa_ctrl[26].f.spare[13] );
tran (\sa_ctrl[26][19] , \sa_ctrl[26].r.part0[19] );
tran (\sa_ctrl[26][19] , \sa_ctrl[26].f.spare[14] );
tran (\sa_ctrl[26][20] , \sa_ctrl[26].r.part0[20] );
tran (\sa_ctrl[26][20] , \sa_ctrl[26].f.spare[15] );
tran (\sa_ctrl[26][21] , \sa_ctrl[26].r.part0[21] );
tran (\sa_ctrl[26][21] , \sa_ctrl[26].f.spare[16] );
tran (\sa_ctrl[26][22] , \sa_ctrl[26].r.part0[22] );
tran (\sa_ctrl[26][22] , \sa_ctrl[26].f.spare[17] );
tran (\sa_ctrl[26][23] , \sa_ctrl[26].r.part0[23] );
tran (\sa_ctrl[26][23] , \sa_ctrl[26].f.spare[18] );
tran (\sa_ctrl[26][24] , \sa_ctrl[26].r.part0[24] );
tran (\sa_ctrl[26][24] , \sa_ctrl[26].f.spare[19] );
tran (\sa_ctrl[26][25] , \sa_ctrl[26].r.part0[25] );
tran (\sa_ctrl[26][25] , \sa_ctrl[26].f.spare[20] );
tran (\sa_ctrl[26][26] , \sa_ctrl[26].r.part0[26] );
tran (\sa_ctrl[26][26] , \sa_ctrl[26].f.spare[21] );
tran (\sa_ctrl[26][27] , \sa_ctrl[26].r.part0[27] );
tran (\sa_ctrl[26][27] , \sa_ctrl[26].f.spare[22] );
tran (\sa_ctrl[26][28] , \sa_ctrl[26].r.part0[28] );
tran (\sa_ctrl[26][28] , \sa_ctrl[26].f.spare[23] );
tran (\sa_ctrl[26][29] , \sa_ctrl[26].r.part0[29] );
tran (\sa_ctrl[26][29] , \sa_ctrl[26].f.spare[24] );
tran (\sa_ctrl[26][30] , \sa_ctrl[26].r.part0[30] );
tran (\sa_ctrl[26][30] , \sa_ctrl[26].f.spare[25] );
tran (\sa_ctrl[26][31] , \sa_ctrl[26].r.part0[31] );
tran (\sa_ctrl[26][31] , \sa_ctrl[26].f.spare[26] );
tran (\sa_ctrl[27][0] , \sa_ctrl[27].r.part0[0] );
tran (\sa_ctrl[27][0] , \sa_ctrl[27].f.sa_event_sel[0] );
tran (\sa_ctrl[27][1] , \sa_ctrl[27].r.part0[1] );
tran (\sa_ctrl[27][1] , \sa_ctrl[27].f.sa_event_sel[1] );
tran (\sa_ctrl[27][2] , \sa_ctrl[27].r.part0[2] );
tran (\sa_ctrl[27][2] , \sa_ctrl[27].f.sa_event_sel[2] );
tran (\sa_ctrl[27][3] , \sa_ctrl[27].r.part0[3] );
tran (\sa_ctrl[27][3] , \sa_ctrl[27].f.sa_event_sel[3] );
tran (\sa_ctrl[27][4] , \sa_ctrl[27].r.part0[4] );
tran (\sa_ctrl[27][4] , \sa_ctrl[27].f.sa_event_sel[4] );
tran (\sa_ctrl[27][5] , \sa_ctrl[27].r.part0[5] );
tran (\sa_ctrl[27][5] , \sa_ctrl[27].f.spare[0] );
tran (\sa_ctrl[27][6] , \sa_ctrl[27].r.part0[6] );
tran (\sa_ctrl[27][6] , \sa_ctrl[27].f.spare[1] );
tran (\sa_ctrl[27][7] , \sa_ctrl[27].r.part0[7] );
tran (\sa_ctrl[27][7] , \sa_ctrl[27].f.spare[2] );
tran (\sa_ctrl[27][8] , \sa_ctrl[27].r.part0[8] );
tran (\sa_ctrl[27][8] , \sa_ctrl[27].f.spare[3] );
tran (\sa_ctrl[27][9] , \sa_ctrl[27].r.part0[9] );
tran (\sa_ctrl[27][9] , \sa_ctrl[27].f.spare[4] );
tran (\sa_ctrl[27][10] , \sa_ctrl[27].r.part0[10] );
tran (\sa_ctrl[27][10] , \sa_ctrl[27].f.spare[5] );
tran (\sa_ctrl[27][11] , \sa_ctrl[27].r.part0[11] );
tran (\sa_ctrl[27][11] , \sa_ctrl[27].f.spare[6] );
tran (\sa_ctrl[27][12] , \sa_ctrl[27].r.part0[12] );
tran (\sa_ctrl[27][12] , \sa_ctrl[27].f.spare[7] );
tran (\sa_ctrl[27][13] , \sa_ctrl[27].r.part0[13] );
tran (\sa_ctrl[27][13] , \sa_ctrl[27].f.spare[8] );
tran (\sa_ctrl[27][14] , \sa_ctrl[27].r.part0[14] );
tran (\sa_ctrl[27][14] , \sa_ctrl[27].f.spare[9] );
tran (\sa_ctrl[27][15] , \sa_ctrl[27].r.part0[15] );
tran (\sa_ctrl[27][15] , \sa_ctrl[27].f.spare[10] );
tran (\sa_ctrl[27][16] , \sa_ctrl[27].r.part0[16] );
tran (\sa_ctrl[27][16] , \sa_ctrl[27].f.spare[11] );
tran (\sa_ctrl[27][17] , \sa_ctrl[27].r.part0[17] );
tran (\sa_ctrl[27][17] , \sa_ctrl[27].f.spare[12] );
tran (\sa_ctrl[27][18] , \sa_ctrl[27].r.part0[18] );
tran (\sa_ctrl[27][18] , \sa_ctrl[27].f.spare[13] );
tran (\sa_ctrl[27][19] , \sa_ctrl[27].r.part0[19] );
tran (\sa_ctrl[27][19] , \sa_ctrl[27].f.spare[14] );
tran (\sa_ctrl[27][20] , \sa_ctrl[27].r.part0[20] );
tran (\sa_ctrl[27][20] , \sa_ctrl[27].f.spare[15] );
tran (\sa_ctrl[27][21] , \sa_ctrl[27].r.part0[21] );
tran (\sa_ctrl[27][21] , \sa_ctrl[27].f.spare[16] );
tran (\sa_ctrl[27][22] , \sa_ctrl[27].r.part0[22] );
tran (\sa_ctrl[27][22] , \sa_ctrl[27].f.spare[17] );
tran (\sa_ctrl[27][23] , \sa_ctrl[27].r.part0[23] );
tran (\sa_ctrl[27][23] , \sa_ctrl[27].f.spare[18] );
tran (\sa_ctrl[27][24] , \sa_ctrl[27].r.part0[24] );
tran (\sa_ctrl[27][24] , \sa_ctrl[27].f.spare[19] );
tran (\sa_ctrl[27][25] , \sa_ctrl[27].r.part0[25] );
tran (\sa_ctrl[27][25] , \sa_ctrl[27].f.spare[20] );
tran (\sa_ctrl[27][26] , \sa_ctrl[27].r.part0[26] );
tran (\sa_ctrl[27][26] , \sa_ctrl[27].f.spare[21] );
tran (\sa_ctrl[27][27] , \sa_ctrl[27].r.part0[27] );
tran (\sa_ctrl[27][27] , \sa_ctrl[27].f.spare[22] );
tran (\sa_ctrl[27][28] , \sa_ctrl[27].r.part0[28] );
tran (\sa_ctrl[27][28] , \sa_ctrl[27].f.spare[23] );
tran (\sa_ctrl[27][29] , \sa_ctrl[27].r.part0[29] );
tran (\sa_ctrl[27][29] , \sa_ctrl[27].f.spare[24] );
tran (\sa_ctrl[27][30] , \sa_ctrl[27].r.part0[30] );
tran (\sa_ctrl[27][30] , \sa_ctrl[27].f.spare[25] );
tran (\sa_ctrl[27][31] , \sa_ctrl[27].r.part0[31] );
tran (\sa_ctrl[27][31] , \sa_ctrl[27].f.spare[26] );
tran (\sa_ctrl[28][0] , \sa_ctrl[28].r.part0[0] );
tran (\sa_ctrl[28][0] , \sa_ctrl[28].f.sa_event_sel[0] );
tran (\sa_ctrl[28][1] , \sa_ctrl[28].r.part0[1] );
tran (\sa_ctrl[28][1] , \sa_ctrl[28].f.sa_event_sel[1] );
tran (\sa_ctrl[28][2] , \sa_ctrl[28].r.part0[2] );
tran (\sa_ctrl[28][2] , \sa_ctrl[28].f.sa_event_sel[2] );
tran (\sa_ctrl[28][3] , \sa_ctrl[28].r.part0[3] );
tran (\sa_ctrl[28][3] , \sa_ctrl[28].f.sa_event_sel[3] );
tran (\sa_ctrl[28][4] , \sa_ctrl[28].r.part0[4] );
tran (\sa_ctrl[28][4] , \sa_ctrl[28].f.sa_event_sel[4] );
tran (\sa_ctrl[28][5] , \sa_ctrl[28].r.part0[5] );
tran (\sa_ctrl[28][5] , \sa_ctrl[28].f.spare[0] );
tran (\sa_ctrl[28][6] , \sa_ctrl[28].r.part0[6] );
tran (\sa_ctrl[28][6] , \sa_ctrl[28].f.spare[1] );
tran (\sa_ctrl[28][7] , \sa_ctrl[28].r.part0[7] );
tran (\sa_ctrl[28][7] , \sa_ctrl[28].f.spare[2] );
tran (\sa_ctrl[28][8] , \sa_ctrl[28].r.part0[8] );
tran (\sa_ctrl[28][8] , \sa_ctrl[28].f.spare[3] );
tran (\sa_ctrl[28][9] , \sa_ctrl[28].r.part0[9] );
tran (\sa_ctrl[28][9] , \sa_ctrl[28].f.spare[4] );
tran (\sa_ctrl[28][10] , \sa_ctrl[28].r.part0[10] );
tran (\sa_ctrl[28][10] , \sa_ctrl[28].f.spare[5] );
tran (\sa_ctrl[28][11] , \sa_ctrl[28].r.part0[11] );
tran (\sa_ctrl[28][11] , \sa_ctrl[28].f.spare[6] );
tran (\sa_ctrl[28][12] , \sa_ctrl[28].r.part0[12] );
tran (\sa_ctrl[28][12] , \sa_ctrl[28].f.spare[7] );
tran (\sa_ctrl[28][13] , \sa_ctrl[28].r.part0[13] );
tran (\sa_ctrl[28][13] , \sa_ctrl[28].f.spare[8] );
tran (\sa_ctrl[28][14] , \sa_ctrl[28].r.part0[14] );
tran (\sa_ctrl[28][14] , \sa_ctrl[28].f.spare[9] );
tran (\sa_ctrl[28][15] , \sa_ctrl[28].r.part0[15] );
tran (\sa_ctrl[28][15] , \sa_ctrl[28].f.spare[10] );
tran (\sa_ctrl[28][16] , \sa_ctrl[28].r.part0[16] );
tran (\sa_ctrl[28][16] , \sa_ctrl[28].f.spare[11] );
tran (\sa_ctrl[28][17] , \sa_ctrl[28].r.part0[17] );
tran (\sa_ctrl[28][17] , \sa_ctrl[28].f.spare[12] );
tran (\sa_ctrl[28][18] , \sa_ctrl[28].r.part0[18] );
tran (\sa_ctrl[28][18] , \sa_ctrl[28].f.spare[13] );
tran (\sa_ctrl[28][19] , \sa_ctrl[28].r.part0[19] );
tran (\sa_ctrl[28][19] , \sa_ctrl[28].f.spare[14] );
tran (\sa_ctrl[28][20] , \sa_ctrl[28].r.part0[20] );
tran (\sa_ctrl[28][20] , \sa_ctrl[28].f.spare[15] );
tran (\sa_ctrl[28][21] , \sa_ctrl[28].r.part0[21] );
tran (\sa_ctrl[28][21] , \sa_ctrl[28].f.spare[16] );
tran (\sa_ctrl[28][22] , \sa_ctrl[28].r.part0[22] );
tran (\sa_ctrl[28][22] , \sa_ctrl[28].f.spare[17] );
tran (\sa_ctrl[28][23] , \sa_ctrl[28].r.part0[23] );
tran (\sa_ctrl[28][23] , \sa_ctrl[28].f.spare[18] );
tran (\sa_ctrl[28][24] , \sa_ctrl[28].r.part0[24] );
tran (\sa_ctrl[28][24] , \sa_ctrl[28].f.spare[19] );
tran (\sa_ctrl[28][25] , \sa_ctrl[28].r.part0[25] );
tran (\sa_ctrl[28][25] , \sa_ctrl[28].f.spare[20] );
tran (\sa_ctrl[28][26] , \sa_ctrl[28].r.part0[26] );
tran (\sa_ctrl[28][26] , \sa_ctrl[28].f.spare[21] );
tran (\sa_ctrl[28][27] , \sa_ctrl[28].r.part0[27] );
tran (\sa_ctrl[28][27] , \sa_ctrl[28].f.spare[22] );
tran (\sa_ctrl[28][28] , \sa_ctrl[28].r.part0[28] );
tran (\sa_ctrl[28][28] , \sa_ctrl[28].f.spare[23] );
tran (\sa_ctrl[28][29] , \sa_ctrl[28].r.part0[29] );
tran (\sa_ctrl[28][29] , \sa_ctrl[28].f.spare[24] );
tran (\sa_ctrl[28][30] , \sa_ctrl[28].r.part0[30] );
tran (\sa_ctrl[28][30] , \sa_ctrl[28].f.spare[25] );
tran (\sa_ctrl[28][31] , \sa_ctrl[28].r.part0[31] );
tran (\sa_ctrl[28][31] , \sa_ctrl[28].f.spare[26] );
tran (\sa_ctrl[29][0] , \sa_ctrl[29].r.part0[0] );
tran (\sa_ctrl[29][0] , \sa_ctrl[29].f.sa_event_sel[0] );
tran (\sa_ctrl[29][1] , \sa_ctrl[29].r.part0[1] );
tran (\sa_ctrl[29][1] , \sa_ctrl[29].f.sa_event_sel[1] );
tran (\sa_ctrl[29][2] , \sa_ctrl[29].r.part0[2] );
tran (\sa_ctrl[29][2] , \sa_ctrl[29].f.sa_event_sel[2] );
tran (\sa_ctrl[29][3] , \sa_ctrl[29].r.part0[3] );
tran (\sa_ctrl[29][3] , \sa_ctrl[29].f.sa_event_sel[3] );
tran (\sa_ctrl[29][4] , \sa_ctrl[29].r.part0[4] );
tran (\sa_ctrl[29][4] , \sa_ctrl[29].f.sa_event_sel[4] );
tran (\sa_ctrl[29][5] , \sa_ctrl[29].r.part0[5] );
tran (\sa_ctrl[29][5] , \sa_ctrl[29].f.spare[0] );
tran (\sa_ctrl[29][6] , \sa_ctrl[29].r.part0[6] );
tran (\sa_ctrl[29][6] , \sa_ctrl[29].f.spare[1] );
tran (\sa_ctrl[29][7] , \sa_ctrl[29].r.part0[7] );
tran (\sa_ctrl[29][7] , \sa_ctrl[29].f.spare[2] );
tran (\sa_ctrl[29][8] , \sa_ctrl[29].r.part0[8] );
tran (\sa_ctrl[29][8] , \sa_ctrl[29].f.spare[3] );
tran (\sa_ctrl[29][9] , \sa_ctrl[29].r.part0[9] );
tran (\sa_ctrl[29][9] , \sa_ctrl[29].f.spare[4] );
tran (\sa_ctrl[29][10] , \sa_ctrl[29].r.part0[10] );
tran (\sa_ctrl[29][10] , \sa_ctrl[29].f.spare[5] );
tran (\sa_ctrl[29][11] , \sa_ctrl[29].r.part0[11] );
tran (\sa_ctrl[29][11] , \sa_ctrl[29].f.spare[6] );
tran (\sa_ctrl[29][12] , \sa_ctrl[29].r.part0[12] );
tran (\sa_ctrl[29][12] , \sa_ctrl[29].f.spare[7] );
tran (\sa_ctrl[29][13] , \sa_ctrl[29].r.part0[13] );
tran (\sa_ctrl[29][13] , \sa_ctrl[29].f.spare[8] );
tran (\sa_ctrl[29][14] , \sa_ctrl[29].r.part0[14] );
tran (\sa_ctrl[29][14] , \sa_ctrl[29].f.spare[9] );
tran (\sa_ctrl[29][15] , \sa_ctrl[29].r.part0[15] );
tran (\sa_ctrl[29][15] , \sa_ctrl[29].f.spare[10] );
tran (\sa_ctrl[29][16] , \sa_ctrl[29].r.part0[16] );
tran (\sa_ctrl[29][16] , \sa_ctrl[29].f.spare[11] );
tran (\sa_ctrl[29][17] , \sa_ctrl[29].r.part0[17] );
tran (\sa_ctrl[29][17] , \sa_ctrl[29].f.spare[12] );
tran (\sa_ctrl[29][18] , \sa_ctrl[29].r.part0[18] );
tran (\sa_ctrl[29][18] , \sa_ctrl[29].f.spare[13] );
tran (\sa_ctrl[29][19] , \sa_ctrl[29].r.part0[19] );
tran (\sa_ctrl[29][19] , \sa_ctrl[29].f.spare[14] );
tran (\sa_ctrl[29][20] , \sa_ctrl[29].r.part0[20] );
tran (\sa_ctrl[29][20] , \sa_ctrl[29].f.spare[15] );
tran (\sa_ctrl[29][21] , \sa_ctrl[29].r.part0[21] );
tran (\sa_ctrl[29][21] , \sa_ctrl[29].f.spare[16] );
tran (\sa_ctrl[29][22] , \sa_ctrl[29].r.part0[22] );
tran (\sa_ctrl[29][22] , \sa_ctrl[29].f.spare[17] );
tran (\sa_ctrl[29][23] , \sa_ctrl[29].r.part0[23] );
tran (\sa_ctrl[29][23] , \sa_ctrl[29].f.spare[18] );
tran (\sa_ctrl[29][24] , \sa_ctrl[29].r.part0[24] );
tran (\sa_ctrl[29][24] , \sa_ctrl[29].f.spare[19] );
tran (\sa_ctrl[29][25] , \sa_ctrl[29].r.part0[25] );
tran (\sa_ctrl[29][25] , \sa_ctrl[29].f.spare[20] );
tran (\sa_ctrl[29][26] , \sa_ctrl[29].r.part0[26] );
tran (\sa_ctrl[29][26] , \sa_ctrl[29].f.spare[21] );
tran (\sa_ctrl[29][27] , \sa_ctrl[29].r.part0[27] );
tran (\sa_ctrl[29][27] , \sa_ctrl[29].f.spare[22] );
tran (\sa_ctrl[29][28] , \sa_ctrl[29].r.part0[28] );
tran (\sa_ctrl[29][28] , \sa_ctrl[29].f.spare[23] );
tran (\sa_ctrl[29][29] , \sa_ctrl[29].r.part0[29] );
tran (\sa_ctrl[29][29] , \sa_ctrl[29].f.spare[24] );
tran (\sa_ctrl[29][30] , \sa_ctrl[29].r.part0[30] );
tran (\sa_ctrl[29][30] , \sa_ctrl[29].f.spare[25] );
tran (\sa_ctrl[29][31] , \sa_ctrl[29].r.part0[31] );
tran (\sa_ctrl[29][31] , \sa_ctrl[29].f.spare[26] );
tran (\sa_ctrl[30][0] , \sa_ctrl[30].r.part0[0] );
tran (\sa_ctrl[30][0] , \sa_ctrl[30].f.sa_event_sel[0] );
tran (\sa_ctrl[30][1] , \sa_ctrl[30].r.part0[1] );
tran (\sa_ctrl[30][1] , \sa_ctrl[30].f.sa_event_sel[1] );
tran (\sa_ctrl[30][2] , \sa_ctrl[30].r.part0[2] );
tran (\sa_ctrl[30][2] , \sa_ctrl[30].f.sa_event_sel[2] );
tran (\sa_ctrl[30][3] , \sa_ctrl[30].r.part0[3] );
tran (\sa_ctrl[30][3] , \sa_ctrl[30].f.sa_event_sel[3] );
tran (\sa_ctrl[30][4] , \sa_ctrl[30].r.part0[4] );
tran (\sa_ctrl[30][4] , \sa_ctrl[30].f.sa_event_sel[4] );
tran (\sa_ctrl[30][5] , \sa_ctrl[30].r.part0[5] );
tran (\sa_ctrl[30][5] , \sa_ctrl[30].f.spare[0] );
tran (\sa_ctrl[30][6] , \sa_ctrl[30].r.part0[6] );
tran (\sa_ctrl[30][6] , \sa_ctrl[30].f.spare[1] );
tran (\sa_ctrl[30][7] , \sa_ctrl[30].r.part0[7] );
tran (\sa_ctrl[30][7] , \sa_ctrl[30].f.spare[2] );
tran (\sa_ctrl[30][8] , \sa_ctrl[30].r.part0[8] );
tran (\sa_ctrl[30][8] , \sa_ctrl[30].f.spare[3] );
tran (\sa_ctrl[30][9] , \sa_ctrl[30].r.part0[9] );
tran (\sa_ctrl[30][9] , \sa_ctrl[30].f.spare[4] );
tran (\sa_ctrl[30][10] , \sa_ctrl[30].r.part0[10] );
tran (\sa_ctrl[30][10] , \sa_ctrl[30].f.spare[5] );
tran (\sa_ctrl[30][11] , \sa_ctrl[30].r.part0[11] );
tran (\sa_ctrl[30][11] , \sa_ctrl[30].f.spare[6] );
tran (\sa_ctrl[30][12] , \sa_ctrl[30].r.part0[12] );
tran (\sa_ctrl[30][12] , \sa_ctrl[30].f.spare[7] );
tran (\sa_ctrl[30][13] , \sa_ctrl[30].r.part0[13] );
tran (\sa_ctrl[30][13] , \sa_ctrl[30].f.spare[8] );
tran (\sa_ctrl[30][14] , \sa_ctrl[30].r.part0[14] );
tran (\sa_ctrl[30][14] , \sa_ctrl[30].f.spare[9] );
tran (\sa_ctrl[30][15] , \sa_ctrl[30].r.part0[15] );
tran (\sa_ctrl[30][15] , \sa_ctrl[30].f.spare[10] );
tran (\sa_ctrl[30][16] , \sa_ctrl[30].r.part0[16] );
tran (\sa_ctrl[30][16] , \sa_ctrl[30].f.spare[11] );
tran (\sa_ctrl[30][17] , \sa_ctrl[30].r.part0[17] );
tran (\sa_ctrl[30][17] , \sa_ctrl[30].f.spare[12] );
tran (\sa_ctrl[30][18] , \sa_ctrl[30].r.part0[18] );
tran (\sa_ctrl[30][18] , \sa_ctrl[30].f.spare[13] );
tran (\sa_ctrl[30][19] , \sa_ctrl[30].r.part0[19] );
tran (\sa_ctrl[30][19] , \sa_ctrl[30].f.spare[14] );
tran (\sa_ctrl[30][20] , \sa_ctrl[30].r.part0[20] );
tran (\sa_ctrl[30][20] , \sa_ctrl[30].f.spare[15] );
tran (\sa_ctrl[30][21] , \sa_ctrl[30].r.part0[21] );
tran (\sa_ctrl[30][21] , \sa_ctrl[30].f.spare[16] );
tran (\sa_ctrl[30][22] , \sa_ctrl[30].r.part0[22] );
tran (\sa_ctrl[30][22] , \sa_ctrl[30].f.spare[17] );
tran (\sa_ctrl[30][23] , \sa_ctrl[30].r.part0[23] );
tran (\sa_ctrl[30][23] , \sa_ctrl[30].f.spare[18] );
tran (\sa_ctrl[30][24] , \sa_ctrl[30].r.part0[24] );
tran (\sa_ctrl[30][24] , \sa_ctrl[30].f.spare[19] );
tran (\sa_ctrl[30][25] , \sa_ctrl[30].r.part0[25] );
tran (\sa_ctrl[30][25] , \sa_ctrl[30].f.spare[20] );
tran (\sa_ctrl[30][26] , \sa_ctrl[30].r.part0[26] );
tran (\sa_ctrl[30][26] , \sa_ctrl[30].f.spare[21] );
tran (\sa_ctrl[30][27] , \sa_ctrl[30].r.part0[27] );
tran (\sa_ctrl[30][27] , \sa_ctrl[30].f.spare[22] );
tran (\sa_ctrl[30][28] , \sa_ctrl[30].r.part0[28] );
tran (\sa_ctrl[30][28] , \sa_ctrl[30].f.spare[23] );
tran (\sa_ctrl[30][29] , \sa_ctrl[30].r.part0[29] );
tran (\sa_ctrl[30][29] , \sa_ctrl[30].f.spare[24] );
tran (\sa_ctrl[30][30] , \sa_ctrl[30].r.part0[30] );
tran (\sa_ctrl[30][30] , \sa_ctrl[30].f.spare[25] );
tran (\sa_ctrl[30][31] , \sa_ctrl[30].r.part0[31] );
tran (\sa_ctrl[30][31] , \sa_ctrl[30].f.spare[26] );
tran (\sa_ctrl[31][0] , \sa_ctrl[31].r.part0[0] );
tran (\sa_ctrl[31][0] , \sa_ctrl[31].f.sa_event_sel[0] );
tran (\sa_ctrl[31][1] , \sa_ctrl[31].r.part0[1] );
tran (\sa_ctrl[31][1] , \sa_ctrl[31].f.sa_event_sel[1] );
tran (\sa_ctrl[31][2] , \sa_ctrl[31].r.part0[2] );
tran (\sa_ctrl[31][2] , \sa_ctrl[31].f.sa_event_sel[2] );
tran (\sa_ctrl[31][3] , \sa_ctrl[31].r.part0[3] );
tran (\sa_ctrl[31][3] , \sa_ctrl[31].f.sa_event_sel[3] );
tran (\sa_ctrl[31][4] , \sa_ctrl[31].r.part0[4] );
tran (\sa_ctrl[31][4] , \sa_ctrl[31].f.sa_event_sel[4] );
tran (\sa_ctrl[31][5] , \sa_ctrl[31].r.part0[5] );
tran (\sa_ctrl[31][5] , \sa_ctrl[31].f.spare[0] );
tran (\sa_ctrl[31][6] , \sa_ctrl[31].r.part0[6] );
tran (\sa_ctrl[31][6] , \sa_ctrl[31].f.spare[1] );
tran (\sa_ctrl[31][7] , \sa_ctrl[31].r.part0[7] );
tran (\sa_ctrl[31][7] , \sa_ctrl[31].f.spare[2] );
tran (\sa_ctrl[31][8] , \sa_ctrl[31].r.part0[8] );
tran (\sa_ctrl[31][8] , \sa_ctrl[31].f.spare[3] );
tran (\sa_ctrl[31][9] , \sa_ctrl[31].r.part0[9] );
tran (\sa_ctrl[31][9] , \sa_ctrl[31].f.spare[4] );
tran (\sa_ctrl[31][10] , \sa_ctrl[31].r.part0[10] );
tran (\sa_ctrl[31][10] , \sa_ctrl[31].f.spare[5] );
tran (\sa_ctrl[31][11] , \sa_ctrl[31].r.part0[11] );
tran (\sa_ctrl[31][11] , \sa_ctrl[31].f.spare[6] );
tran (\sa_ctrl[31][12] , \sa_ctrl[31].r.part0[12] );
tran (\sa_ctrl[31][12] , \sa_ctrl[31].f.spare[7] );
tran (\sa_ctrl[31][13] , \sa_ctrl[31].r.part0[13] );
tran (\sa_ctrl[31][13] , \sa_ctrl[31].f.spare[8] );
tran (\sa_ctrl[31][14] , \sa_ctrl[31].r.part0[14] );
tran (\sa_ctrl[31][14] , \sa_ctrl[31].f.spare[9] );
tran (\sa_ctrl[31][15] , \sa_ctrl[31].r.part0[15] );
tran (\sa_ctrl[31][15] , \sa_ctrl[31].f.spare[10] );
tran (\sa_ctrl[31][16] , \sa_ctrl[31].r.part0[16] );
tran (\sa_ctrl[31][16] , \sa_ctrl[31].f.spare[11] );
tran (\sa_ctrl[31][17] , \sa_ctrl[31].r.part0[17] );
tran (\sa_ctrl[31][17] , \sa_ctrl[31].f.spare[12] );
tran (\sa_ctrl[31][18] , \sa_ctrl[31].r.part0[18] );
tran (\sa_ctrl[31][18] , \sa_ctrl[31].f.spare[13] );
tran (\sa_ctrl[31][19] , \sa_ctrl[31].r.part0[19] );
tran (\sa_ctrl[31][19] , \sa_ctrl[31].f.spare[14] );
tran (\sa_ctrl[31][20] , \sa_ctrl[31].r.part0[20] );
tran (\sa_ctrl[31][20] , \sa_ctrl[31].f.spare[15] );
tran (\sa_ctrl[31][21] , \sa_ctrl[31].r.part0[21] );
tran (\sa_ctrl[31][21] , \sa_ctrl[31].f.spare[16] );
tran (\sa_ctrl[31][22] , \sa_ctrl[31].r.part0[22] );
tran (\sa_ctrl[31][22] , \sa_ctrl[31].f.spare[17] );
tran (\sa_ctrl[31][23] , \sa_ctrl[31].r.part0[23] );
tran (\sa_ctrl[31][23] , \sa_ctrl[31].f.spare[18] );
tran (\sa_ctrl[31][24] , \sa_ctrl[31].r.part0[24] );
tran (\sa_ctrl[31][24] , \sa_ctrl[31].f.spare[19] );
tran (\sa_ctrl[31][25] , \sa_ctrl[31].r.part0[25] );
tran (\sa_ctrl[31][25] , \sa_ctrl[31].f.spare[20] );
tran (\sa_ctrl[31][26] , \sa_ctrl[31].r.part0[26] );
tran (\sa_ctrl[31][26] , \sa_ctrl[31].f.spare[21] );
tran (\sa_ctrl[31][27] , \sa_ctrl[31].r.part0[27] );
tran (\sa_ctrl[31][27] , \sa_ctrl[31].f.spare[22] );
tran (\sa_ctrl[31][28] , \sa_ctrl[31].r.part0[28] );
tran (\sa_ctrl[31][28] , \sa_ctrl[31].f.spare[23] );
tran (\sa_ctrl[31][29] , \sa_ctrl[31].r.part0[29] );
tran (\sa_ctrl[31][29] , \sa_ctrl[31].f.spare[24] );
tran (\sa_ctrl[31][30] , \sa_ctrl[31].r.part0[30] );
tran (\sa_ctrl[31][30] , \sa_ctrl[31].f.spare[25] );
tran (\sa_ctrl[31][31] , \sa_ctrl[31].r.part0[31] );
tran (\sa_ctrl[31][31] , \sa_ctrl[31].f.spare[26] );
Q_BUF U0 ( .A(n1), .Z(\sa_snapshot[31][63] ));
Q_BUF U1 ( .A(n1), .Z(\sa_snapshot[31][62] ));
Q_BUF U2 ( .A(n1), .Z(\sa_snapshot[31][61] ));
Q_BUF U3 ( .A(n1), .Z(\sa_snapshot[31][60] ));
Q_BUF U4 ( .A(n1), .Z(\sa_snapshot[31][59] ));
Q_BUF U5 ( .A(n1), .Z(\sa_snapshot[31][58] ));
Q_BUF U6 ( .A(n1), .Z(\sa_snapshot[31][57] ));
Q_BUF U7 ( .A(n1), .Z(\sa_snapshot[31][56] ));
Q_BUF U8 ( .A(n1), .Z(\sa_snapshot[31][55] ));
Q_BUF U9 ( .A(n1), .Z(\sa_snapshot[31][54] ));
Q_BUF U10 ( .A(n1), .Z(\sa_snapshot[31][53] ));
Q_BUF U11 ( .A(n1), .Z(\sa_snapshot[31][52] ));
Q_BUF U12 ( .A(n1), .Z(\sa_snapshot[31][51] ));
Q_BUF U13 ( .A(n1), .Z(\sa_snapshot[31][50] ));
Q_BUF U14 ( .A(n1), .Z(\sa_snapshot[30][63] ));
Q_BUF U15 ( .A(n1), .Z(\sa_snapshot[30][62] ));
Q_BUF U16 ( .A(n1), .Z(\sa_snapshot[30][61] ));
Q_BUF U17 ( .A(n1), .Z(\sa_snapshot[30][60] ));
Q_BUF U18 ( .A(n1), .Z(\sa_snapshot[30][59] ));
Q_BUF U19 ( .A(n1), .Z(\sa_snapshot[30][58] ));
Q_BUF U20 ( .A(n1), .Z(\sa_snapshot[30][57] ));
Q_BUF U21 ( .A(n1), .Z(\sa_snapshot[30][56] ));
Q_BUF U22 ( .A(n1), .Z(\sa_snapshot[30][55] ));
Q_BUF U23 ( .A(n1), .Z(\sa_snapshot[30][54] ));
Q_BUF U24 ( .A(n1), .Z(\sa_snapshot[30][53] ));
Q_BUF U25 ( .A(n1), .Z(\sa_snapshot[30][52] ));
Q_BUF U26 ( .A(n1), .Z(\sa_snapshot[30][51] ));
Q_BUF U27 ( .A(n1), .Z(\sa_snapshot[30][50] ));
Q_BUF U28 ( .A(n1), .Z(\sa_snapshot[29][63] ));
Q_BUF U29 ( .A(n1), .Z(\sa_snapshot[29][62] ));
Q_BUF U30 ( .A(n1), .Z(\sa_snapshot[29][61] ));
Q_BUF U31 ( .A(n1), .Z(\sa_snapshot[29][60] ));
Q_BUF U32 ( .A(n1), .Z(\sa_snapshot[29][59] ));
Q_BUF U33 ( .A(n1), .Z(\sa_snapshot[29][58] ));
Q_BUF U34 ( .A(n1), .Z(\sa_snapshot[29][57] ));
Q_BUF U35 ( .A(n1), .Z(\sa_snapshot[29][56] ));
Q_BUF U36 ( .A(n1), .Z(\sa_snapshot[29][55] ));
Q_BUF U37 ( .A(n1), .Z(\sa_snapshot[29][54] ));
Q_BUF U38 ( .A(n1), .Z(\sa_snapshot[29][53] ));
Q_BUF U39 ( .A(n1), .Z(\sa_snapshot[29][52] ));
Q_BUF U40 ( .A(n1), .Z(\sa_snapshot[29][51] ));
Q_BUF U41 ( .A(n1), .Z(\sa_snapshot[29][50] ));
Q_BUF U42 ( .A(n1), .Z(\sa_snapshot[28][63] ));
Q_BUF U43 ( .A(n1), .Z(\sa_snapshot[28][62] ));
Q_BUF U44 ( .A(n1), .Z(\sa_snapshot[28][61] ));
Q_BUF U45 ( .A(n1), .Z(\sa_snapshot[28][60] ));
Q_BUF U46 ( .A(n1), .Z(\sa_snapshot[28][59] ));
Q_BUF U47 ( .A(n1), .Z(\sa_snapshot[28][58] ));
Q_BUF U48 ( .A(n1), .Z(\sa_snapshot[28][57] ));
Q_BUF U49 ( .A(n1), .Z(\sa_snapshot[28][56] ));
Q_BUF U50 ( .A(n1), .Z(\sa_snapshot[28][55] ));
Q_BUF U51 ( .A(n1), .Z(\sa_snapshot[28][54] ));
Q_BUF U52 ( .A(n1), .Z(\sa_snapshot[28][53] ));
Q_BUF U53 ( .A(n1), .Z(\sa_snapshot[28][52] ));
Q_BUF U54 ( .A(n1), .Z(\sa_snapshot[28][51] ));
Q_BUF U55 ( .A(n1), .Z(\sa_snapshot[28][50] ));
Q_BUF U56 ( .A(n1), .Z(\sa_snapshot[27][63] ));
Q_BUF U57 ( .A(n1), .Z(\sa_snapshot[27][62] ));
Q_BUF U58 ( .A(n1), .Z(\sa_snapshot[27][61] ));
Q_BUF U59 ( .A(n1), .Z(\sa_snapshot[27][60] ));
Q_BUF U60 ( .A(n1), .Z(\sa_snapshot[27][59] ));
Q_BUF U61 ( .A(n1), .Z(\sa_snapshot[27][58] ));
Q_BUF U62 ( .A(n1), .Z(\sa_snapshot[27][57] ));
Q_BUF U63 ( .A(n1), .Z(\sa_snapshot[27][56] ));
Q_BUF U64 ( .A(n1), .Z(\sa_snapshot[27][55] ));
Q_BUF U65 ( .A(n1), .Z(\sa_snapshot[27][54] ));
Q_BUF U66 ( .A(n1), .Z(\sa_snapshot[27][53] ));
Q_BUF U67 ( .A(n1), .Z(\sa_snapshot[27][52] ));
Q_BUF U68 ( .A(n1), .Z(\sa_snapshot[27][51] ));
Q_BUF U69 ( .A(n1), .Z(\sa_snapshot[27][50] ));
Q_BUF U70 ( .A(n1), .Z(\sa_snapshot[26][63] ));
Q_BUF U71 ( .A(n1), .Z(\sa_snapshot[26][62] ));
Q_BUF U72 ( .A(n1), .Z(\sa_snapshot[26][61] ));
Q_BUF U73 ( .A(n1), .Z(\sa_snapshot[26][60] ));
Q_BUF U74 ( .A(n1), .Z(\sa_snapshot[26][59] ));
Q_BUF U75 ( .A(n1), .Z(\sa_snapshot[26][58] ));
Q_BUF U76 ( .A(n1), .Z(\sa_snapshot[26][57] ));
Q_BUF U77 ( .A(n1), .Z(\sa_snapshot[26][56] ));
Q_BUF U78 ( .A(n1), .Z(\sa_snapshot[26][55] ));
Q_BUF U79 ( .A(n1), .Z(\sa_snapshot[26][54] ));
Q_BUF U80 ( .A(n1), .Z(\sa_snapshot[26][53] ));
Q_BUF U81 ( .A(n1), .Z(\sa_snapshot[26][52] ));
Q_BUF U82 ( .A(n1), .Z(\sa_snapshot[26][51] ));
Q_BUF U83 ( .A(n1), .Z(\sa_snapshot[26][50] ));
Q_BUF U84 ( .A(n1), .Z(\sa_snapshot[25][63] ));
Q_BUF U85 ( .A(n1), .Z(\sa_snapshot[25][62] ));
Q_BUF U86 ( .A(n1), .Z(\sa_snapshot[25][61] ));
Q_BUF U87 ( .A(n1), .Z(\sa_snapshot[25][60] ));
Q_BUF U88 ( .A(n1), .Z(\sa_snapshot[25][59] ));
Q_BUF U89 ( .A(n1), .Z(\sa_snapshot[25][58] ));
Q_BUF U90 ( .A(n1), .Z(\sa_snapshot[25][57] ));
Q_BUF U91 ( .A(n1), .Z(\sa_snapshot[25][56] ));
Q_BUF U92 ( .A(n1), .Z(\sa_snapshot[25][55] ));
Q_BUF U93 ( .A(n1), .Z(\sa_snapshot[25][54] ));
Q_BUF U94 ( .A(n1), .Z(\sa_snapshot[25][53] ));
Q_BUF U95 ( .A(n1), .Z(\sa_snapshot[25][52] ));
Q_BUF U96 ( .A(n1), .Z(\sa_snapshot[25][51] ));
Q_BUF U97 ( .A(n1), .Z(\sa_snapshot[25][50] ));
Q_BUF U98 ( .A(n1), .Z(\sa_snapshot[24][63] ));
Q_BUF U99 ( .A(n1), .Z(\sa_snapshot[24][62] ));
Q_BUF U100 ( .A(n1), .Z(\sa_snapshot[24][61] ));
Q_BUF U101 ( .A(n1), .Z(\sa_snapshot[24][60] ));
Q_BUF U102 ( .A(n1), .Z(\sa_snapshot[24][59] ));
Q_BUF U103 ( .A(n1), .Z(\sa_snapshot[24][58] ));
Q_BUF U104 ( .A(n1), .Z(\sa_snapshot[24][57] ));
Q_BUF U105 ( .A(n1), .Z(\sa_snapshot[24][56] ));
Q_BUF U106 ( .A(n1), .Z(\sa_snapshot[24][55] ));
Q_BUF U107 ( .A(n1), .Z(\sa_snapshot[24][54] ));
Q_BUF U108 ( .A(n1), .Z(\sa_snapshot[24][53] ));
Q_BUF U109 ( .A(n1), .Z(\sa_snapshot[24][52] ));
Q_BUF U110 ( .A(n1), .Z(\sa_snapshot[24][51] ));
Q_BUF U111 ( .A(n1), .Z(\sa_snapshot[24][50] ));
Q_BUF U112 ( .A(n1), .Z(\sa_snapshot[23][63] ));
Q_BUF U113 ( .A(n1), .Z(\sa_snapshot[23][62] ));
Q_BUF U114 ( .A(n1), .Z(\sa_snapshot[23][61] ));
Q_BUF U115 ( .A(n1), .Z(\sa_snapshot[23][60] ));
Q_BUF U116 ( .A(n1), .Z(\sa_snapshot[23][59] ));
Q_BUF U117 ( .A(n1), .Z(\sa_snapshot[23][58] ));
Q_BUF U118 ( .A(n1), .Z(\sa_snapshot[23][57] ));
Q_BUF U119 ( .A(n1), .Z(\sa_snapshot[23][56] ));
Q_BUF U120 ( .A(n1), .Z(\sa_snapshot[23][55] ));
Q_BUF U121 ( .A(n1), .Z(\sa_snapshot[23][54] ));
Q_BUF U122 ( .A(n1), .Z(\sa_snapshot[23][53] ));
Q_BUF U123 ( .A(n1), .Z(\sa_snapshot[23][52] ));
Q_BUF U124 ( .A(n1), .Z(\sa_snapshot[23][51] ));
Q_BUF U125 ( .A(n1), .Z(\sa_snapshot[23][50] ));
Q_BUF U126 ( .A(n1), .Z(\sa_snapshot[22][63] ));
Q_BUF U127 ( .A(n1), .Z(\sa_snapshot[22][62] ));
Q_BUF U128 ( .A(n1), .Z(\sa_snapshot[22][61] ));
Q_BUF U129 ( .A(n1), .Z(\sa_snapshot[22][60] ));
Q_BUF U130 ( .A(n1), .Z(\sa_snapshot[22][59] ));
Q_BUF U131 ( .A(n1), .Z(\sa_snapshot[22][58] ));
Q_BUF U132 ( .A(n1), .Z(\sa_snapshot[22][57] ));
Q_BUF U133 ( .A(n1), .Z(\sa_snapshot[22][56] ));
Q_BUF U134 ( .A(n1), .Z(\sa_snapshot[22][55] ));
Q_BUF U135 ( .A(n1), .Z(\sa_snapshot[22][54] ));
Q_BUF U136 ( .A(n1), .Z(\sa_snapshot[22][53] ));
Q_BUF U137 ( .A(n1), .Z(\sa_snapshot[22][52] ));
Q_BUF U138 ( .A(n1), .Z(\sa_snapshot[22][51] ));
Q_BUF U139 ( .A(n1), .Z(\sa_snapshot[22][50] ));
Q_BUF U140 ( .A(n1), .Z(\sa_snapshot[21][63] ));
Q_BUF U141 ( .A(n1), .Z(\sa_snapshot[21][62] ));
Q_BUF U142 ( .A(n1), .Z(\sa_snapshot[21][61] ));
Q_BUF U143 ( .A(n1), .Z(\sa_snapshot[21][60] ));
Q_BUF U144 ( .A(n1), .Z(\sa_snapshot[21][59] ));
Q_BUF U145 ( .A(n1), .Z(\sa_snapshot[21][58] ));
Q_BUF U146 ( .A(n1), .Z(\sa_snapshot[21][57] ));
Q_BUF U147 ( .A(n1), .Z(\sa_snapshot[21][56] ));
Q_BUF U148 ( .A(n1), .Z(\sa_snapshot[21][55] ));
Q_BUF U149 ( .A(n1), .Z(\sa_snapshot[21][54] ));
Q_BUF U150 ( .A(n1), .Z(\sa_snapshot[21][53] ));
Q_BUF U151 ( .A(n1), .Z(\sa_snapshot[21][52] ));
Q_BUF U152 ( .A(n1), .Z(\sa_snapshot[21][51] ));
Q_BUF U153 ( .A(n1), .Z(\sa_snapshot[21][50] ));
Q_BUF U154 ( .A(n1), .Z(\sa_snapshot[20][63] ));
Q_BUF U155 ( .A(n1), .Z(\sa_snapshot[20][62] ));
Q_BUF U156 ( .A(n1), .Z(\sa_snapshot[20][61] ));
Q_BUF U157 ( .A(n1), .Z(\sa_snapshot[20][60] ));
Q_BUF U158 ( .A(n1), .Z(\sa_snapshot[20][59] ));
Q_BUF U159 ( .A(n1), .Z(\sa_snapshot[20][58] ));
Q_BUF U160 ( .A(n1), .Z(\sa_snapshot[20][57] ));
Q_BUF U161 ( .A(n1), .Z(\sa_snapshot[20][56] ));
Q_BUF U162 ( .A(n1), .Z(\sa_snapshot[20][55] ));
Q_BUF U163 ( .A(n1), .Z(\sa_snapshot[20][54] ));
Q_BUF U164 ( .A(n1), .Z(\sa_snapshot[20][53] ));
Q_BUF U165 ( .A(n1), .Z(\sa_snapshot[20][52] ));
Q_BUF U166 ( .A(n1), .Z(\sa_snapshot[20][51] ));
Q_BUF U167 ( .A(n1), .Z(\sa_snapshot[20][50] ));
Q_BUF U168 ( .A(n1), .Z(\sa_snapshot[19][63] ));
Q_BUF U169 ( .A(n1), .Z(\sa_snapshot[19][62] ));
Q_BUF U170 ( .A(n1), .Z(\sa_snapshot[19][61] ));
Q_BUF U171 ( .A(n1), .Z(\sa_snapshot[19][60] ));
Q_BUF U172 ( .A(n1), .Z(\sa_snapshot[19][59] ));
Q_BUF U173 ( .A(n1), .Z(\sa_snapshot[19][58] ));
Q_BUF U174 ( .A(n1), .Z(\sa_snapshot[19][57] ));
Q_BUF U175 ( .A(n1), .Z(\sa_snapshot[19][56] ));
Q_BUF U176 ( .A(n1), .Z(\sa_snapshot[19][55] ));
Q_BUF U177 ( .A(n1), .Z(\sa_snapshot[19][54] ));
Q_BUF U178 ( .A(n1), .Z(\sa_snapshot[19][53] ));
Q_BUF U179 ( .A(n1), .Z(\sa_snapshot[19][52] ));
Q_BUF U180 ( .A(n1), .Z(\sa_snapshot[19][51] ));
Q_BUF U181 ( .A(n1), .Z(\sa_snapshot[19][50] ));
Q_BUF U182 ( .A(n1), .Z(\sa_snapshot[18][63] ));
Q_BUF U183 ( .A(n1), .Z(\sa_snapshot[18][62] ));
Q_BUF U184 ( .A(n1), .Z(\sa_snapshot[18][61] ));
Q_BUF U185 ( .A(n1), .Z(\sa_snapshot[18][60] ));
Q_BUF U186 ( .A(n1), .Z(\sa_snapshot[18][59] ));
Q_BUF U187 ( .A(n1), .Z(\sa_snapshot[18][58] ));
Q_BUF U188 ( .A(n1), .Z(\sa_snapshot[18][57] ));
Q_BUF U189 ( .A(n1), .Z(\sa_snapshot[18][56] ));
Q_BUF U190 ( .A(n1), .Z(\sa_snapshot[18][55] ));
Q_BUF U191 ( .A(n1), .Z(\sa_snapshot[18][54] ));
Q_BUF U192 ( .A(n1), .Z(\sa_snapshot[18][53] ));
Q_BUF U193 ( .A(n1), .Z(\sa_snapshot[18][52] ));
Q_BUF U194 ( .A(n1), .Z(\sa_snapshot[18][51] ));
Q_BUF U195 ( .A(n1), .Z(\sa_snapshot[18][50] ));
Q_BUF U196 ( .A(n1), .Z(\sa_snapshot[17][63] ));
Q_BUF U197 ( .A(n1), .Z(\sa_snapshot[17][62] ));
Q_BUF U198 ( .A(n1), .Z(\sa_snapshot[17][61] ));
Q_BUF U199 ( .A(n1), .Z(\sa_snapshot[17][60] ));
Q_BUF U200 ( .A(n1), .Z(\sa_snapshot[17][59] ));
Q_BUF U201 ( .A(n1), .Z(\sa_snapshot[17][58] ));
Q_BUF U202 ( .A(n1), .Z(\sa_snapshot[17][57] ));
Q_BUF U203 ( .A(n1), .Z(\sa_snapshot[17][56] ));
Q_BUF U204 ( .A(n1), .Z(\sa_snapshot[17][55] ));
Q_BUF U205 ( .A(n1), .Z(\sa_snapshot[17][54] ));
Q_BUF U206 ( .A(n1), .Z(\sa_snapshot[17][53] ));
Q_BUF U207 ( .A(n1), .Z(\sa_snapshot[17][52] ));
Q_BUF U208 ( .A(n1), .Z(\sa_snapshot[17][51] ));
Q_BUF U209 ( .A(n1), .Z(\sa_snapshot[17][50] ));
Q_BUF U210 ( .A(n1), .Z(\sa_snapshot[16][63] ));
Q_BUF U211 ( .A(n1), .Z(\sa_snapshot[16][62] ));
Q_BUF U212 ( .A(n1), .Z(\sa_snapshot[16][61] ));
Q_BUF U213 ( .A(n1), .Z(\sa_snapshot[16][60] ));
Q_BUF U214 ( .A(n1), .Z(\sa_snapshot[16][59] ));
Q_BUF U215 ( .A(n1), .Z(\sa_snapshot[16][58] ));
Q_BUF U216 ( .A(n1), .Z(\sa_snapshot[16][57] ));
Q_BUF U217 ( .A(n1), .Z(\sa_snapshot[16][56] ));
Q_BUF U218 ( .A(n1), .Z(\sa_snapshot[16][55] ));
Q_BUF U219 ( .A(n1), .Z(\sa_snapshot[16][54] ));
Q_BUF U220 ( .A(n1), .Z(\sa_snapshot[16][53] ));
Q_BUF U221 ( .A(n1), .Z(\sa_snapshot[16][52] ));
Q_BUF U222 ( .A(n1), .Z(\sa_snapshot[16][51] ));
Q_BUF U223 ( .A(n1), .Z(\sa_snapshot[16][50] ));
Q_BUF U224 ( .A(n1), .Z(\sa_snapshot[15][63] ));
Q_BUF U225 ( .A(n1), .Z(\sa_snapshot[15][62] ));
Q_BUF U226 ( .A(n1), .Z(\sa_snapshot[15][61] ));
Q_BUF U227 ( .A(n1), .Z(\sa_snapshot[15][60] ));
Q_BUF U228 ( .A(n1), .Z(\sa_snapshot[15][59] ));
Q_BUF U229 ( .A(n1), .Z(\sa_snapshot[15][58] ));
Q_BUF U230 ( .A(n1), .Z(\sa_snapshot[15][57] ));
Q_BUF U231 ( .A(n1), .Z(\sa_snapshot[15][56] ));
Q_BUF U232 ( .A(n1), .Z(\sa_snapshot[15][55] ));
Q_BUF U233 ( .A(n1), .Z(\sa_snapshot[15][54] ));
Q_BUF U234 ( .A(n1), .Z(\sa_snapshot[15][53] ));
Q_BUF U235 ( .A(n1), .Z(\sa_snapshot[15][52] ));
Q_BUF U236 ( .A(n1), .Z(\sa_snapshot[15][51] ));
Q_BUF U237 ( .A(n1), .Z(\sa_snapshot[15][50] ));
Q_BUF U238 ( .A(n1), .Z(\sa_snapshot[14][63] ));
Q_BUF U239 ( .A(n1), .Z(\sa_snapshot[14][62] ));
Q_BUF U240 ( .A(n1), .Z(\sa_snapshot[14][61] ));
Q_BUF U241 ( .A(n1), .Z(\sa_snapshot[14][60] ));
Q_BUF U242 ( .A(n1), .Z(\sa_snapshot[14][59] ));
Q_BUF U243 ( .A(n1), .Z(\sa_snapshot[14][58] ));
Q_BUF U244 ( .A(n1), .Z(\sa_snapshot[14][57] ));
Q_BUF U245 ( .A(n1), .Z(\sa_snapshot[14][56] ));
Q_BUF U246 ( .A(n1), .Z(\sa_snapshot[14][55] ));
Q_BUF U247 ( .A(n1), .Z(\sa_snapshot[14][54] ));
Q_BUF U248 ( .A(n1), .Z(\sa_snapshot[14][53] ));
Q_BUF U249 ( .A(n1), .Z(\sa_snapshot[14][52] ));
Q_BUF U250 ( .A(n1), .Z(\sa_snapshot[14][51] ));
Q_BUF U251 ( .A(n1), .Z(\sa_snapshot[14][50] ));
Q_BUF U252 ( .A(n1), .Z(\sa_snapshot[13][63] ));
Q_BUF U253 ( .A(n1), .Z(\sa_snapshot[13][62] ));
Q_BUF U254 ( .A(n1), .Z(\sa_snapshot[13][61] ));
Q_BUF U255 ( .A(n1), .Z(\sa_snapshot[13][60] ));
Q_BUF U256 ( .A(n1), .Z(\sa_snapshot[13][59] ));
Q_BUF U257 ( .A(n1), .Z(\sa_snapshot[13][58] ));
Q_BUF U258 ( .A(n1), .Z(\sa_snapshot[13][57] ));
Q_BUF U259 ( .A(n1), .Z(\sa_snapshot[13][56] ));
Q_BUF U260 ( .A(n1), .Z(\sa_snapshot[13][55] ));
Q_BUF U261 ( .A(n1), .Z(\sa_snapshot[13][54] ));
Q_BUF U262 ( .A(n1), .Z(\sa_snapshot[13][53] ));
Q_BUF U263 ( .A(n1), .Z(\sa_snapshot[13][52] ));
Q_BUF U264 ( .A(n1), .Z(\sa_snapshot[13][51] ));
Q_BUF U265 ( .A(n1), .Z(\sa_snapshot[13][50] ));
Q_BUF U266 ( .A(n1), .Z(\sa_snapshot[12][63] ));
Q_BUF U267 ( .A(n1), .Z(\sa_snapshot[12][62] ));
Q_BUF U268 ( .A(n1), .Z(\sa_snapshot[12][61] ));
Q_BUF U269 ( .A(n1), .Z(\sa_snapshot[12][60] ));
Q_BUF U270 ( .A(n1), .Z(\sa_snapshot[12][59] ));
Q_BUF U271 ( .A(n1), .Z(\sa_snapshot[12][58] ));
Q_BUF U272 ( .A(n1), .Z(\sa_snapshot[12][57] ));
Q_BUF U273 ( .A(n1), .Z(\sa_snapshot[12][56] ));
Q_BUF U274 ( .A(n1), .Z(\sa_snapshot[12][55] ));
Q_BUF U275 ( .A(n1), .Z(\sa_snapshot[12][54] ));
Q_BUF U276 ( .A(n1), .Z(\sa_snapshot[12][53] ));
Q_BUF U277 ( .A(n1), .Z(\sa_snapshot[12][52] ));
Q_BUF U278 ( .A(n1), .Z(\sa_snapshot[12][51] ));
Q_BUF U279 ( .A(n1), .Z(\sa_snapshot[12][50] ));
Q_BUF U280 ( .A(n1), .Z(\sa_snapshot[11][63] ));
Q_BUF U281 ( .A(n1), .Z(\sa_snapshot[11][62] ));
Q_BUF U282 ( .A(n1), .Z(\sa_snapshot[11][61] ));
Q_BUF U283 ( .A(n1), .Z(\sa_snapshot[11][60] ));
Q_BUF U284 ( .A(n1), .Z(\sa_snapshot[11][59] ));
Q_BUF U285 ( .A(n1), .Z(\sa_snapshot[11][58] ));
Q_BUF U286 ( .A(n1), .Z(\sa_snapshot[11][57] ));
Q_BUF U287 ( .A(n1), .Z(\sa_snapshot[11][56] ));
Q_BUF U288 ( .A(n1), .Z(\sa_snapshot[11][55] ));
Q_BUF U289 ( .A(n1), .Z(\sa_snapshot[11][54] ));
Q_BUF U290 ( .A(n1), .Z(\sa_snapshot[11][53] ));
Q_BUF U291 ( .A(n1), .Z(\sa_snapshot[11][52] ));
Q_BUF U292 ( .A(n1), .Z(\sa_snapshot[11][51] ));
Q_BUF U293 ( .A(n1), .Z(\sa_snapshot[11][50] ));
Q_BUF U294 ( .A(n1), .Z(\sa_snapshot[10][63] ));
Q_BUF U295 ( .A(n1), .Z(\sa_snapshot[10][62] ));
Q_BUF U296 ( .A(n1), .Z(\sa_snapshot[10][61] ));
Q_BUF U297 ( .A(n1), .Z(\sa_snapshot[10][60] ));
Q_BUF U298 ( .A(n1), .Z(\sa_snapshot[10][59] ));
Q_BUF U299 ( .A(n1), .Z(\sa_snapshot[10][58] ));
Q_BUF U300 ( .A(n1), .Z(\sa_snapshot[10][57] ));
Q_BUF U301 ( .A(n1), .Z(\sa_snapshot[10][56] ));
Q_BUF U302 ( .A(n1), .Z(\sa_snapshot[10][55] ));
Q_BUF U303 ( .A(n1), .Z(\sa_snapshot[10][54] ));
Q_BUF U304 ( .A(n1), .Z(\sa_snapshot[10][53] ));
Q_BUF U305 ( .A(n1), .Z(\sa_snapshot[10][52] ));
Q_BUF U306 ( .A(n1), .Z(\sa_snapshot[10][51] ));
Q_BUF U307 ( .A(n1), .Z(\sa_snapshot[10][50] ));
Q_BUF U308 ( .A(n1), .Z(\sa_snapshot[9][63] ));
Q_BUF U309 ( .A(n1), .Z(\sa_snapshot[9][62] ));
Q_BUF U310 ( .A(n1), .Z(\sa_snapshot[9][61] ));
Q_BUF U311 ( .A(n1), .Z(\sa_snapshot[9][60] ));
Q_BUF U312 ( .A(n1), .Z(\sa_snapshot[9][59] ));
Q_BUF U313 ( .A(n1), .Z(\sa_snapshot[9][58] ));
Q_BUF U314 ( .A(n1), .Z(\sa_snapshot[9][57] ));
Q_BUF U315 ( .A(n1), .Z(\sa_snapshot[9][56] ));
Q_BUF U316 ( .A(n1), .Z(\sa_snapshot[9][55] ));
Q_BUF U317 ( .A(n1), .Z(\sa_snapshot[9][54] ));
Q_BUF U318 ( .A(n1), .Z(\sa_snapshot[9][53] ));
Q_BUF U319 ( .A(n1), .Z(\sa_snapshot[9][52] ));
Q_BUF U320 ( .A(n1), .Z(\sa_snapshot[9][51] ));
Q_BUF U321 ( .A(n1), .Z(\sa_snapshot[9][50] ));
Q_BUF U322 ( .A(n1), .Z(\sa_snapshot[8][63] ));
Q_BUF U323 ( .A(n1), .Z(\sa_snapshot[8][62] ));
Q_BUF U324 ( .A(n1), .Z(\sa_snapshot[8][61] ));
Q_BUF U325 ( .A(n1), .Z(\sa_snapshot[8][60] ));
Q_BUF U326 ( .A(n1), .Z(\sa_snapshot[8][59] ));
Q_BUF U327 ( .A(n1), .Z(\sa_snapshot[8][58] ));
Q_BUF U328 ( .A(n1), .Z(\sa_snapshot[8][57] ));
Q_BUF U329 ( .A(n1), .Z(\sa_snapshot[8][56] ));
Q_BUF U330 ( .A(n1), .Z(\sa_snapshot[8][55] ));
Q_BUF U331 ( .A(n1), .Z(\sa_snapshot[8][54] ));
Q_BUF U332 ( .A(n1), .Z(\sa_snapshot[8][53] ));
Q_BUF U333 ( .A(n1), .Z(\sa_snapshot[8][52] ));
Q_BUF U334 ( .A(n1), .Z(\sa_snapshot[8][51] ));
Q_BUF U335 ( .A(n1), .Z(\sa_snapshot[8][50] ));
Q_BUF U336 ( .A(n1), .Z(\sa_snapshot[7][63] ));
Q_BUF U337 ( .A(n1), .Z(\sa_snapshot[7][62] ));
Q_BUF U338 ( .A(n1), .Z(\sa_snapshot[7][61] ));
Q_BUF U339 ( .A(n1), .Z(\sa_snapshot[7][60] ));
Q_BUF U340 ( .A(n1), .Z(\sa_snapshot[7][59] ));
Q_BUF U341 ( .A(n1), .Z(\sa_snapshot[7][58] ));
Q_BUF U342 ( .A(n1), .Z(\sa_snapshot[7][57] ));
Q_BUF U343 ( .A(n1), .Z(\sa_snapshot[7][56] ));
Q_BUF U344 ( .A(n1), .Z(\sa_snapshot[7][55] ));
Q_BUF U345 ( .A(n1), .Z(\sa_snapshot[7][54] ));
Q_BUF U346 ( .A(n1), .Z(\sa_snapshot[7][53] ));
Q_BUF U347 ( .A(n1), .Z(\sa_snapshot[7][52] ));
Q_BUF U348 ( .A(n1), .Z(\sa_snapshot[7][51] ));
Q_BUF U349 ( .A(n1), .Z(\sa_snapshot[7][50] ));
Q_BUF U350 ( .A(n1), .Z(\sa_snapshot[6][63] ));
Q_BUF U351 ( .A(n1), .Z(\sa_snapshot[6][62] ));
Q_BUF U352 ( .A(n1), .Z(\sa_snapshot[6][61] ));
Q_BUF U353 ( .A(n1), .Z(\sa_snapshot[6][60] ));
Q_BUF U354 ( .A(n1), .Z(\sa_snapshot[6][59] ));
Q_BUF U355 ( .A(n1), .Z(\sa_snapshot[6][58] ));
Q_BUF U356 ( .A(n1), .Z(\sa_snapshot[6][57] ));
Q_BUF U357 ( .A(n1), .Z(\sa_snapshot[6][56] ));
Q_BUF U358 ( .A(n1), .Z(\sa_snapshot[6][55] ));
Q_BUF U359 ( .A(n1), .Z(\sa_snapshot[6][54] ));
Q_BUF U360 ( .A(n1), .Z(\sa_snapshot[6][53] ));
Q_BUF U361 ( .A(n1), .Z(\sa_snapshot[6][52] ));
Q_BUF U362 ( .A(n1), .Z(\sa_snapshot[6][51] ));
Q_BUF U363 ( .A(n1), .Z(\sa_snapshot[6][50] ));
Q_BUF U364 ( .A(n1), .Z(\sa_snapshot[5][63] ));
Q_BUF U365 ( .A(n1), .Z(\sa_snapshot[5][62] ));
Q_BUF U366 ( .A(n1), .Z(\sa_snapshot[5][61] ));
Q_BUF U367 ( .A(n1), .Z(\sa_snapshot[5][60] ));
Q_BUF U368 ( .A(n1), .Z(\sa_snapshot[5][59] ));
Q_BUF U369 ( .A(n1), .Z(\sa_snapshot[5][58] ));
Q_BUF U370 ( .A(n1), .Z(\sa_snapshot[5][57] ));
Q_BUF U371 ( .A(n1), .Z(\sa_snapshot[5][56] ));
Q_BUF U372 ( .A(n1), .Z(\sa_snapshot[5][55] ));
Q_BUF U373 ( .A(n1), .Z(\sa_snapshot[5][54] ));
Q_BUF U374 ( .A(n1), .Z(\sa_snapshot[5][53] ));
Q_BUF U375 ( .A(n1), .Z(\sa_snapshot[5][52] ));
Q_BUF U376 ( .A(n1), .Z(\sa_snapshot[5][51] ));
Q_BUF U377 ( .A(n1), .Z(\sa_snapshot[5][50] ));
Q_BUF U378 ( .A(n1), .Z(\sa_snapshot[4][63] ));
Q_BUF U379 ( .A(n1), .Z(\sa_snapshot[4][62] ));
Q_BUF U380 ( .A(n1), .Z(\sa_snapshot[4][61] ));
Q_BUF U381 ( .A(n1), .Z(\sa_snapshot[4][60] ));
Q_BUF U382 ( .A(n1), .Z(\sa_snapshot[4][59] ));
Q_BUF U383 ( .A(n1), .Z(\sa_snapshot[4][58] ));
Q_BUF U384 ( .A(n1), .Z(\sa_snapshot[4][57] ));
Q_BUF U385 ( .A(n1), .Z(\sa_snapshot[4][56] ));
Q_BUF U386 ( .A(n1), .Z(\sa_snapshot[4][55] ));
Q_BUF U387 ( .A(n1), .Z(\sa_snapshot[4][54] ));
Q_BUF U388 ( .A(n1), .Z(\sa_snapshot[4][53] ));
Q_BUF U389 ( .A(n1), .Z(\sa_snapshot[4][52] ));
Q_BUF U390 ( .A(n1), .Z(\sa_snapshot[4][51] ));
Q_BUF U391 ( .A(n1), .Z(\sa_snapshot[4][50] ));
Q_BUF U392 ( .A(n1), .Z(\sa_snapshot[3][63] ));
Q_BUF U393 ( .A(n1), .Z(\sa_snapshot[3][62] ));
Q_BUF U394 ( .A(n1), .Z(\sa_snapshot[3][61] ));
Q_BUF U395 ( .A(n1), .Z(\sa_snapshot[3][60] ));
Q_BUF U396 ( .A(n1), .Z(\sa_snapshot[3][59] ));
Q_BUF U397 ( .A(n1), .Z(\sa_snapshot[3][58] ));
Q_BUF U398 ( .A(n1), .Z(\sa_snapshot[3][57] ));
Q_BUF U399 ( .A(n1), .Z(\sa_snapshot[3][56] ));
Q_BUF U400 ( .A(n1), .Z(\sa_snapshot[3][55] ));
Q_BUF U401 ( .A(n1), .Z(\sa_snapshot[3][54] ));
Q_BUF U402 ( .A(n1), .Z(\sa_snapshot[3][53] ));
Q_BUF U403 ( .A(n1), .Z(\sa_snapshot[3][52] ));
Q_BUF U404 ( .A(n1), .Z(\sa_snapshot[3][51] ));
Q_BUF U405 ( .A(n1), .Z(\sa_snapshot[3][50] ));
Q_BUF U406 ( .A(n1), .Z(\sa_snapshot[2][63] ));
Q_BUF U407 ( .A(n1), .Z(\sa_snapshot[2][62] ));
Q_BUF U408 ( .A(n1), .Z(\sa_snapshot[2][61] ));
Q_BUF U409 ( .A(n1), .Z(\sa_snapshot[2][60] ));
Q_BUF U410 ( .A(n1), .Z(\sa_snapshot[2][59] ));
Q_BUF U411 ( .A(n1), .Z(\sa_snapshot[2][58] ));
Q_BUF U412 ( .A(n1), .Z(\sa_snapshot[2][57] ));
Q_BUF U413 ( .A(n1), .Z(\sa_snapshot[2][56] ));
Q_BUF U414 ( .A(n1), .Z(\sa_snapshot[2][55] ));
Q_BUF U415 ( .A(n1), .Z(\sa_snapshot[2][54] ));
Q_BUF U416 ( .A(n1), .Z(\sa_snapshot[2][53] ));
Q_BUF U417 ( .A(n1), .Z(\sa_snapshot[2][52] ));
Q_BUF U418 ( .A(n1), .Z(\sa_snapshot[2][51] ));
Q_BUF U419 ( .A(n1), .Z(\sa_snapshot[2][50] ));
Q_BUF U420 ( .A(n1), .Z(\sa_snapshot[1][63] ));
Q_BUF U421 ( .A(n1), .Z(\sa_snapshot[1][62] ));
Q_BUF U422 ( .A(n1), .Z(\sa_snapshot[1][61] ));
Q_BUF U423 ( .A(n1), .Z(\sa_snapshot[1][60] ));
Q_BUF U424 ( .A(n1), .Z(\sa_snapshot[1][59] ));
Q_BUF U425 ( .A(n1), .Z(\sa_snapshot[1][58] ));
Q_BUF U426 ( .A(n1), .Z(\sa_snapshot[1][57] ));
Q_BUF U427 ( .A(n1), .Z(\sa_snapshot[1][56] ));
Q_BUF U428 ( .A(n1), .Z(\sa_snapshot[1][55] ));
Q_BUF U429 ( .A(n1), .Z(\sa_snapshot[1][54] ));
Q_BUF U430 ( .A(n1), .Z(\sa_snapshot[1][53] ));
Q_BUF U431 ( .A(n1), .Z(\sa_snapshot[1][52] ));
Q_BUF U432 ( .A(n1), .Z(\sa_snapshot[1][51] ));
Q_BUF U433 ( .A(n1), .Z(\sa_snapshot[1][50] ));
Q_BUF U434 ( .A(n1), .Z(\sa_snapshot[0][63] ));
Q_BUF U435 ( .A(n1), .Z(\sa_snapshot[0][62] ));
Q_BUF U436 ( .A(n1), .Z(\sa_snapshot[0][61] ));
Q_BUF U437 ( .A(n1), .Z(\sa_snapshot[0][60] ));
Q_BUF U438 ( .A(n1), .Z(\sa_snapshot[0][59] ));
Q_BUF U439 ( .A(n1), .Z(\sa_snapshot[0][58] ));
Q_BUF U440 ( .A(n1), .Z(\sa_snapshot[0][57] ));
Q_BUF U441 ( .A(n1), .Z(\sa_snapshot[0][56] ));
Q_BUF U442 ( .A(n1), .Z(\sa_snapshot[0][55] ));
Q_BUF U443 ( .A(n1), .Z(\sa_snapshot[0][54] ));
Q_BUF U444 ( .A(n1), .Z(\sa_snapshot[0][53] ));
Q_BUF U445 ( .A(n1), .Z(\sa_snapshot[0][52] ));
Q_BUF U446 ( .A(n1), .Z(\sa_snapshot[0][51] ));
Q_BUF U447 ( .A(n1), .Z(\sa_snapshot[0][50] ));
Q_BUF U448 ( .A(n1), .Z(\sa_count[31][63] ));
Q_BUF U449 ( .A(n1), .Z(\sa_count[31][62] ));
Q_BUF U450 ( .A(n1), .Z(\sa_count[31][61] ));
Q_BUF U451 ( .A(n1), .Z(\sa_count[31][60] ));
Q_BUF U452 ( .A(n1), .Z(\sa_count[31][59] ));
Q_BUF U453 ( .A(n1), .Z(\sa_count[31][58] ));
Q_BUF U454 ( .A(n1), .Z(\sa_count[31][57] ));
Q_BUF U455 ( .A(n1), .Z(\sa_count[31][56] ));
Q_BUF U456 ( .A(n1), .Z(\sa_count[31][55] ));
Q_BUF U457 ( .A(n1), .Z(\sa_count[31][54] ));
Q_BUF U458 ( .A(n1), .Z(\sa_count[31][53] ));
Q_BUF U459 ( .A(n1), .Z(\sa_count[31][52] ));
Q_BUF U460 ( .A(n1), .Z(\sa_count[31][51] ));
Q_BUF U461 ( .A(n1), .Z(\sa_count[31][50] ));
Q_BUF U462 ( .A(n1), .Z(\sa_count[30][63] ));
Q_BUF U463 ( .A(n1), .Z(\sa_count[30][62] ));
Q_BUF U464 ( .A(n1), .Z(\sa_count[30][61] ));
Q_BUF U465 ( .A(n1), .Z(\sa_count[30][60] ));
Q_BUF U466 ( .A(n1), .Z(\sa_count[30][59] ));
Q_BUF U467 ( .A(n1), .Z(\sa_count[30][58] ));
Q_BUF U468 ( .A(n1), .Z(\sa_count[30][57] ));
Q_BUF U469 ( .A(n1), .Z(\sa_count[30][56] ));
Q_BUF U470 ( .A(n1), .Z(\sa_count[30][55] ));
Q_BUF U471 ( .A(n1), .Z(\sa_count[30][54] ));
Q_BUF U472 ( .A(n1), .Z(\sa_count[30][53] ));
Q_BUF U473 ( .A(n1), .Z(\sa_count[30][52] ));
Q_BUF U474 ( .A(n1), .Z(\sa_count[30][51] ));
Q_BUF U475 ( .A(n1), .Z(\sa_count[30][50] ));
Q_BUF U476 ( .A(n1), .Z(\sa_count[29][63] ));
Q_BUF U477 ( .A(n1), .Z(\sa_count[29][62] ));
Q_BUF U478 ( .A(n1), .Z(\sa_count[29][61] ));
Q_BUF U479 ( .A(n1), .Z(\sa_count[29][60] ));
Q_BUF U480 ( .A(n1), .Z(\sa_count[29][59] ));
Q_BUF U481 ( .A(n1), .Z(\sa_count[29][58] ));
Q_BUF U482 ( .A(n1), .Z(\sa_count[29][57] ));
Q_BUF U483 ( .A(n1), .Z(\sa_count[29][56] ));
Q_BUF U484 ( .A(n1), .Z(\sa_count[29][55] ));
Q_BUF U485 ( .A(n1), .Z(\sa_count[29][54] ));
Q_BUF U486 ( .A(n1), .Z(\sa_count[29][53] ));
Q_BUF U487 ( .A(n1), .Z(\sa_count[29][52] ));
Q_BUF U488 ( .A(n1), .Z(\sa_count[29][51] ));
Q_BUF U489 ( .A(n1), .Z(\sa_count[29][50] ));
Q_BUF U490 ( .A(n1), .Z(\sa_count[28][63] ));
Q_BUF U491 ( .A(n1), .Z(\sa_count[28][62] ));
Q_BUF U492 ( .A(n1), .Z(\sa_count[28][61] ));
Q_BUF U493 ( .A(n1), .Z(\sa_count[28][60] ));
Q_BUF U494 ( .A(n1), .Z(\sa_count[28][59] ));
Q_BUF U495 ( .A(n1), .Z(\sa_count[28][58] ));
Q_BUF U496 ( .A(n1), .Z(\sa_count[28][57] ));
Q_BUF U497 ( .A(n1), .Z(\sa_count[28][56] ));
Q_BUF U498 ( .A(n1), .Z(\sa_count[28][55] ));
Q_BUF U499 ( .A(n1), .Z(\sa_count[28][54] ));
Q_BUF U500 ( .A(n1), .Z(\sa_count[28][53] ));
Q_BUF U501 ( .A(n1), .Z(\sa_count[28][52] ));
Q_BUF U502 ( .A(n1), .Z(\sa_count[28][51] ));
Q_BUF U503 ( .A(n1), .Z(\sa_count[28][50] ));
Q_BUF U504 ( .A(n1), .Z(\sa_count[27][63] ));
Q_BUF U505 ( .A(n1), .Z(\sa_count[27][62] ));
Q_BUF U506 ( .A(n1), .Z(\sa_count[27][61] ));
Q_BUF U507 ( .A(n1), .Z(\sa_count[27][60] ));
Q_BUF U508 ( .A(n1), .Z(\sa_count[27][59] ));
Q_BUF U509 ( .A(n1), .Z(\sa_count[27][58] ));
Q_BUF U510 ( .A(n1), .Z(\sa_count[27][57] ));
Q_BUF U511 ( .A(n1), .Z(\sa_count[27][56] ));
Q_BUF U512 ( .A(n1), .Z(\sa_count[27][55] ));
Q_BUF U513 ( .A(n1), .Z(\sa_count[27][54] ));
Q_BUF U514 ( .A(n1), .Z(\sa_count[27][53] ));
Q_BUF U515 ( .A(n1), .Z(\sa_count[27][52] ));
Q_BUF U516 ( .A(n1), .Z(\sa_count[27][51] ));
Q_BUF U517 ( .A(n1), .Z(\sa_count[27][50] ));
Q_BUF U518 ( .A(n1), .Z(\sa_count[26][63] ));
Q_BUF U519 ( .A(n1), .Z(\sa_count[26][62] ));
Q_BUF U520 ( .A(n1), .Z(\sa_count[26][61] ));
Q_BUF U521 ( .A(n1), .Z(\sa_count[26][60] ));
Q_BUF U522 ( .A(n1), .Z(\sa_count[26][59] ));
Q_BUF U523 ( .A(n1), .Z(\sa_count[26][58] ));
Q_BUF U524 ( .A(n1), .Z(\sa_count[26][57] ));
Q_BUF U525 ( .A(n1), .Z(\sa_count[26][56] ));
Q_BUF U526 ( .A(n1), .Z(\sa_count[26][55] ));
Q_BUF U527 ( .A(n1), .Z(\sa_count[26][54] ));
Q_BUF U528 ( .A(n1), .Z(\sa_count[26][53] ));
Q_BUF U529 ( .A(n1), .Z(\sa_count[26][52] ));
Q_BUF U530 ( .A(n1), .Z(\sa_count[26][51] ));
Q_BUF U531 ( .A(n1), .Z(\sa_count[26][50] ));
Q_BUF U532 ( .A(n1), .Z(\sa_count[25][63] ));
Q_BUF U533 ( .A(n1), .Z(\sa_count[25][62] ));
Q_BUF U534 ( .A(n1), .Z(\sa_count[25][61] ));
Q_BUF U535 ( .A(n1), .Z(\sa_count[25][60] ));
Q_BUF U536 ( .A(n1), .Z(\sa_count[25][59] ));
Q_BUF U537 ( .A(n1), .Z(\sa_count[25][58] ));
Q_BUF U538 ( .A(n1), .Z(\sa_count[25][57] ));
Q_BUF U539 ( .A(n1), .Z(\sa_count[25][56] ));
Q_BUF U540 ( .A(n1), .Z(\sa_count[25][55] ));
Q_BUF U541 ( .A(n1), .Z(\sa_count[25][54] ));
Q_BUF U542 ( .A(n1), .Z(\sa_count[25][53] ));
Q_BUF U543 ( .A(n1), .Z(\sa_count[25][52] ));
Q_BUF U544 ( .A(n1), .Z(\sa_count[25][51] ));
Q_BUF U545 ( .A(n1), .Z(\sa_count[25][50] ));
Q_BUF U546 ( .A(n1), .Z(\sa_count[24][63] ));
Q_BUF U547 ( .A(n1), .Z(\sa_count[24][62] ));
Q_BUF U548 ( .A(n1), .Z(\sa_count[24][61] ));
Q_BUF U549 ( .A(n1), .Z(\sa_count[24][60] ));
Q_BUF U550 ( .A(n1), .Z(\sa_count[24][59] ));
Q_BUF U551 ( .A(n1), .Z(\sa_count[24][58] ));
Q_BUF U552 ( .A(n1), .Z(\sa_count[24][57] ));
Q_BUF U553 ( .A(n1), .Z(\sa_count[24][56] ));
Q_BUF U554 ( .A(n1), .Z(\sa_count[24][55] ));
Q_BUF U555 ( .A(n1), .Z(\sa_count[24][54] ));
Q_BUF U556 ( .A(n1), .Z(\sa_count[24][53] ));
Q_BUF U557 ( .A(n1), .Z(\sa_count[24][52] ));
Q_BUF U558 ( .A(n1), .Z(\sa_count[24][51] ));
Q_BUF U559 ( .A(n1), .Z(\sa_count[24][50] ));
Q_BUF U560 ( .A(n1), .Z(\sa_count[23][63] ));
Q_BUF U561 ( .A(n1), .Z(\sa_count[23][62] ));
Q_BUF U562 ( .A(n1), .Z(\sa_count[23][61] ));
Q_BUF U563 ( .A(n1), .Z(\sa_count[23][60] ));
Q_BUF U564 ( .A(n1), .Z(\sa_count[23][59] ));
Q_BUF U565 ( .A(n1), .Z(\sa_count[23][58] ));
Q_BUF U566 ( .A(n1), .Z(\sa_count[23][57] ));
Q_BUF U567 ( .A(n1), .Z(\sa_count[23][56] ));
Q_BUF U568 ( .A(n1), .Z(\sa_count[23][55] ));
Q_BUF U569 ( .A(n1), .Z(\sa_count[23][54] ));
Q_BUF U570 ( .A(n1), .Z(\sa_count[23][53] ));
Q_BUF U571 ( .A(n1), .Z(\sa_count[23][52] ));
Q_BUF U572 ( .A(n1), .Z(\sa_count[23][51] ));
Q_BUF U573 ( .A(n1), .Z(\sa_count[23][50] ));
Q_BUF U574 ( .A(n1), .Z(\sa_count[22][63] ));
Q_BUF U575 ( .A(n1), .Z(\sa_count[22][62] ));
Q_BUF U576 ( .A(n1), .Z(\sa_count[22][61] ));
Q_BUF U577 ( .A(n1), .Z(\sa_count[22][60] ));
Q_BUF U578 ( .A(n1), .Z(\sa_count[22][59] ));
Q_BUF U579 ( .A(n1), .Z(\sa_count[22][58] ));
Q_BUF U580 ( .A(n1), .Z(\sa_count[22][57] ));
Q_BUF U581 ( .A(n1), .Z(\sa_count[22][56] ));
Q_BUF U582 ( .A(n1), .Z(\sa_count[22][55] ));
Q_BUF U583 ( .A(n1), .Z(\sa_count[22][54] ));
Q_BUF U584 ( .A(n1), .Z(\sa_count[22][53] ));
Q_BUF U585 ( .A(n1), .Z(\sa_count[22][52] ));
Q_BUF U586 ( .A(n1), .Z(\sa_count[22][51] ));
Q_BUF U587 ( .A(n1), .Z(\sa_count[22][50] ));
Q_BUF U588 ( .A(n1), .Z(\sa_count[21][63] ));
Q_BUF U589 ( .A(n1), .Z(\sa_count[21][62] ));
Q_BUF U590 ( .A(n1), .Z(\sa_count[21][61] ));
Q_BUF U591 ( .A(n1), .Z(\sa_count[21][60] ));
Q_BUF U592 ( .A(n1), .Z(\sa_count[21][59] ));
Q_BUF U593 ( .A(n1), .Z(\sa_count[21][58] ));
Q_BUF U594 ( .A(n1), .Z(\sa_count[21][57] ));
Q_BUF U595 ( .A(n1), .Z(\sa_count[21][56] ));
Q_BUF U596 ( .A(n1), .Z(\sa_count[21][55] ));
Q_BUF U597 ( .A(n1), .Z(\sa_count[21][54] ));
Q_BUF U598 ( .A(n1), .Z(\sa_count[21][53] ));
Q_BUF U599 ( .A(n1), .Z(\sa_count[21][52] ));
Q_BUF U600 ( .A(n1), .Z(\sa_count[21][51] ));
Q_BUF U601 ( .A(n1), .Z(\sa_count[21][50] ));
Q_BUF U602 ( .A(n1), .Z(\sa_count[20][63] ));
Q_BUF U603 ( .A(n1), .Z(\sa_count[20][62] ));
Q_BUF U604 ( .A(n1), .Z(\sa_count[20][61] ));
Q_BUF U605 ( .A(n1), .Z(\sa_count[20][60] ));
Q_BUF U606 ( .A(n1), .Z(\sa_count[20][59] ));
Q_BUF U607 ( .A(n1), .Z(\sa_count[20][58] ));
Q_BUF U608 ( .A(n1), .Z(\sa_count[20][57] ));
Q_BUF U609 ( .A(n1), .Z(\sa_count[20][56] ));
Q_BUF U610 ( .A(n1), .Z(\sa_count[20][55] ));
Q_BUF U611 ( .A(n1), .Z(\sa_count[20][54] ));
Q_BUF U612 ( .A(n1), .Z(\sa_count[20][53] ));
Q_BUF U613 ( .A(n1), .Z(\sa_count[20][52] ));
Q_BUF U614 ( .A(n1), .Z(\sa_count[20][51] ));
Q_BUF U615 ( .A(n1), .Z(\sa_count[20][50] ));
Q_BUF U616 ( .A(n1), .Z(\sa_count[19][63] ));
Q_BUF U617 ( .A(n1), .Z(\sa_count[19][62] ));
Q_BUF U618 ( .A(n1), .Z(\sa_count[19][61] ));
Q_BUF U619 ( .A(n1), .Z(\sa_count[19][60] ));
Q_BUF U620 ( .A(n1), .Z(\sa_count[19][59] ));
Q_BUF U621 ( .A(n1), .Z(\sa_count[19][58] ));
Q_BUF U622 ( .A(n1), .Z(\sa_count[19][57] ));
Q_BUF U623 ( .A(n1), .Z(\sa_count[19][56] ));
Q_BUF U624 ( .A(n1), .Z(\sa_count[19][55] ));
Q_BUF U625 ( .A(n1), .Z(\sa_count[19][54] ));
Q_BUF U626 ( .A(n1), .Z(\sa_count[19][53] ));
Q_BUF U627 ( .A(n1), .Z(\sa_count[19][52] ));
Q_BUF U628 ( .A(n1), .Z(\sa_count[19][51] ));
Q_BUF U629 ( .A(n1), .Z(\sa_count[19][50] ));
Q_BUF U630 ( .A(n1), .Z(\sa_count[18][63] ));
Q_BUF U631 ( .A(n1), .Z(\sa_count[18][62] ));
Q_BUF U632 ( .A(n1), .Z(\sa_count[18][61] ));
Q_BUF U633 ( .A(n1), .Z(\sa_count[18][60] ));
Q_BUF U634 ( .A(n1), .Z(\sa_count[18][59] ));
Q_BUF U635 ( .A(n1), .Z(\sa_count[18][58] ));
Q_BUF U636 ( .A(n1), .Z(\sa_count[18][57] ));
Q_BUF U637 ( .A(n1), .Z(\sa_count[18][56] ));
Q_BUF U638 ( .A(n1), .Z(\sa_count[18][55] ));
Q_BUF U639 ( .A(n1), .Z(\sa_count[18][54] ));
Q_BUF U640 ( .A(n1), .Z(\sa_count[18][53] ));
Q_BUF U641 ( .A(n1), .Z(\sa_count[18][52] ));
Q_BUF U642 ( .A(n1), .Z(\sa_count[18][51] ));
Q_BUF U643 ( .A(n1), .Z(\sa_count[18][50] ));
Q_BUF U644 ( .A(n1), .Z(\sa_count[17][63] ));
Q_BUF U645 ( .A(n1), .Z(\sa_count[17][62] ));
Q_BUF U646 ( .A(n1), .Z(\sa_count[17][61] ));
Q_BUF U647 ( .A(n1), .Z(\sa_count[17][60] ));
Q_BUF U648 ( .A(n1), .Z(\sa_count[17][59] ));
Q_BUF U649 ( .A(n1), .Z(\sa_count[17][58] ));
Q_BUF U650 ( .A(n1), .Z(\sa_count[17][57] ));
Q_BUF U651 ( .A(n1), .Z(\sa_count[17][56] ));
Q_BUF U652 ( .A(n1), .Z(\sa_count[17][55] ));
Q_BUF U653 ( .A(n1), .Z(\sa_count[17][54] ));
Q_BUF U654 ( .A(n1), .Z(\sa_count[17][53] ));
Q_BUF U655 ( .A(n1), .Z(\sa_count[17][52] ));
Q_BUF U656 ( .A(n1), .Z(\sa_count[17][51] ));
Q_BUF U657 ( .A(n1), .Z(\sa_count[17][50] ));
Q_BUF U658 ( .A(n1), .Z(\sa_count[16][63] ));
Q_BUF U659 ( .A(n1), .Z(\sa_count[16][62] ));
Q_BUF U660 ( .A(n1), .Z(\sa_count[16][61] ));
Q_BUF U661 ( .A(n1), .Z(\sa_count[16][60] ));
Q_BUF U662 ( .A(n1), .Z(\sa_count[16][59] ));
Q_BUF U663 ( .A(n1), .Z(\sa_count[16][58] ));
Q_BUF U664 ( .A(n1), .Z(\sa_count[16][57] ));
Q_BUF U665 ( .A(n1), .Z(\sa_count[16][56] ));
Q_BUF U666 ( .A(n1), .Z(\sa_count[16][55] ));
Q_BUF U667 ( .A(n1), .Z(\sa_count[16][54] ));
Q_BUF U668 ( .A(n1), .Z(\sa_count[16][53] ));
Q_BUF U669 ( .A(n1), .Z(\sa_count[16][52] ));
Q_BUF U670 ( .A(n1), .Z(\sa_count[16][51] ));
Q_BUF U671 ( .A(n1), .Z(\sa_count[16][50] ));
Q_BUF U672 ( .A(n1), .Z(\sa_count[15][63] ));
Q_BUF U673 ( .A(n1), .Z(\sa_count[15][62] ));
Q_BUF U674 ( .A(n1), .Z(\sa_count[15][61] ));
Q_BUF U675 ( .A(n1), .Z(\sa_count[15][60] ));
Q_BUF U676 ( .A(n1), .Z(\sa_count[15][59] ));
Q_BUF U677 ( .A(n1), .Z(\sa_count[15][58] ));
Q_BUF U678 ( .A(n1), .Z(\sa_count[15][57] ));
Q_BUF U679 ( .A(n1), .Z(\sa_count[15][56] ));
Q_BUF U680 ( .A(n1), .Z(\sa_count[15][55] ));
Q_BUF U681 ( .A(n1), .Z(\sa_count[15][54] ));
Q_BUF U682 ( .A(n1), .Z(\sa_count[15][53] ));
Q_BUF U683 ( .A(n1), .Z(\sa_count[15][52] ));
Q_BUF U684 ( .A(n1), .Z(\sa_count[15][51] ));
Q_BUF U685 ( .A(n1), .Z(\sa_count[15][50] ));
Q_BUF U686 ( .A(n1), .Z(\sa_count[14][63] ));
Q_BUF U687 ( .A(n1), .Z(\sa_count[14][62] ));
Q_BUF U688 ( .A(n1), .Z(\sa_count[14][61] ));
Q_BUF U689 ( .A(n1), .Z(\sa_count[14][60] ));
Q_BUF U690 ( .A(n1), .Z(\sa_count[14][59] ));
Q_BUF U691 ( .A(n1), .Z(\sa_count[14][58] ));
Q_BUF U692 ( .A(n1), .Z(\sa_count[14][57] ));
Q_BUF U693 ( .A(n1), .Z(\sa_count[14][56] ));
Q_BUF U694 ( .A(n1), .Z(\sa_count[14][55] ));
Q_BUF U695 ( .A(n1), .Z(\sa_count[14][54] ));
Q_BUF U696 ( .A(n1), .Z(\sa_count[14][53] ));
Q_BUF U697 ( .A(n1), .Z(\sa_count[14][52] ));
Q_BUF U698 ( .A(n1), .Z(\sa_count[14][51] ));
Q_BUF U699 ( .A(n1), .Z(\sa_count[14][50] ));
Q_BUF U700 ( .A(n1), .Z(\sa_count[13][63] ));
Q_BUF U701 ( .A(n1), .Z(\sa_count[13][62] ));
Q_BUF U702 ( .A(n1), .Z(\sa_count[13][61] ));
Q_BUF U703 ( .A(n1), .Z(\sa_count[13][60] ));
Q_BUF U704 ( .A(n1), .Z(\sa_count[13][59] ));
Q_BUF U705 ( .A(n1), .Z(\sa_count[13][58] ));
Q_BUF U706 ( .A(n1), .Z(\sa_count[13][57] ));
Q_BUF U707 ( .A(n1), .Z(\sa_count[13][56] ));
Q_BUF U708 ( .A(n1), .Z(\sa_count[13][55] ));
Q_BUF U709 ( .A(n1), .Z(\sa_count[13][54] ));
Q_BUF U710 ( .A(n1), .Z(\sa_count[13][53] ));
Q_BUF U711 ( .A(n1), .Z(\sa_count[13][52] ));
Q_BUF U712 ( .A(n1), .Z(\sa_count[13][51] ));
Q_BUF U713 ( .A(n1), .Z(\sa_count[13][50] ));
Q_BUF U714 ( .A(n1), .Z(\sa_count[12][63] ));
Q_BUF U715 ( .A(n1), .Z(\sa_count[12][62] ));
Q_BUF U716 ( .A(n1), .Z(\sa_count[12][61] ));
Q_BUF U717 ( .A(n1), .Z(\sa_count[12][60] ));
Q_BUF U718 ( .A(n1), .Z(\sa_count[12][59] ));
Q_BUF U719 ( .A(n1), .Z(\sa_count[12][58] ));
Q_BUF U720 ( .A(n1), .Z(\sa_count[12][57] ));
Q_BUF U721 ( .A(n1), .Z(\sa_count[12][56] ));
Q_BUF U722 ( .A(n1), .Z(\sa_count[12][55] ));
Q_BUF U723 ( .A(n1), .Z(\sa_count[12][54] ));
Q_BUF U724 ( .A(n1), .Z(\sa_count[12][53] ));
Q_BUF U725 ( .A(n1), .Z(\sa_count[12][52] ));
Q_BUF U726 ( .A(n1), .Z(\sa_count[12][51] ));
Q_BUF U727 ( .A(n1), .Z(\sa_count[12][50] ));
Q_BUF U728 ( .A(n1), .Z(\sa_count[11][63] ));
Q_BUF U729 ( .A(n1), .Z(\sa_count[11][62] ));
Q_BUF U730 ( .A(n1), .Z(\sa_count[11][61] ));
Q_BUF U731 ( .A(n1), .Z(\sa_count[11][60] ));
Q_BUF U732 ( .A(n1), .Z(\sa_count[11][59] ));
Q_BUF U733 ( .A(n1), .Z(\sa_count[11][58] ));
Q_BUF U734 ( .A(n1), .Z(\sa_count[11][57] ));
Q_BUF U735 ( .A(n1), .Z(\sa_count[11][56] ));
Q_BUF U736 ( .A(n1), .Z(\sa_count[11][55] ));
Q_BUF U737 ( .A(n1), .Z(\sa_count[11][54] ));
Q_BUF U738 ( .A(n1), .Z(\sa_count[11][53] ));
Q_BUF U739 ( .A(n1), .Z(\sa_count[11][52] ));
Q_BUF U740 ( .A(n1), .Z(\sa_count[11][51] ));
Q_BUF U741 ( .A(n1), .Z(\sa_count[11][50] ));
Q_BUF U742 ( .A(n1), .Z(\sa_count[10][63] ));
Q_BUF U743 ( .A(n1), .Z(\sa_count[10][62] ));
Q_BUF U744 ( .A(n1), .Z(\sa_count[10][61] ));
Q_BUF U745 ( .A(n1), .Z(\sa_count[10][60] ));
Q_BUF U746 ( .A(n1), .Z(\sa_count[10][59] ));
Q_BUF U747 ( .A(n1), .Z(\sa_count[10][58] ));
Q_BUF U748 ( .A(n1), .Z(\sa_count[10][57] ));
Q_BUF U749 ( .A(n1), .Z(\sa_count[10][56] ));
Q_BUF U750 ( .A(n1), .Z(\sa_count[10][55] ));
Q_BUF U751 ( .A(n1), .Z(\sa_count[10][54] ));
Q_BUF U752 ( .A(n1), .Z(\sa_count[10][53] ));
Q_BUF U753 ( .A(n1), .Z(\sa_count[10][52] ));
Q_BUF U754 ( .A(n1), .Z(\sa_count[10][51] ));
Q_BUF U755 ( .A(n1), .Z(\sa_count[10][50] ));
Q_BUF U756 ( .A(n1), .Z(\sa_count[9][63] ));
Q_BUF U757 ( .A(n1), .Z(\sa_count[9][62] ));
Q_BUF U758 ( .A(n1), .Z(\sa_count[9][61] ));
Q_BUF U759 ( .A(n1), .Z(\sa_count[9][60] ));
Q_BUF U760 ( .A(n1), .Z(\sa_count[9][59] ));
Q_BUF U761 ( .A(n1), .Z(\sa_count[9][58] ));
Q_BUF U762 ( .A(n1), .Z(\sa_count[9][57] ));
Q_BUF U763 ( .A(n1), .Z(\sa_count[9][56] ));
Q_BUF U764 ( .A(n1), .Z(\sa_count[9][55] ));
Q_BUF U765 ( .A(n1), .Z(\sa_count[9][54] ));
Q_BUF U766 ( .A(n1), .Z(\sa_count[9][53] ));
Q_BUF U767 ( .A(n1), .Z(\sa_count[9][52] ));
Q_BUF U768 ( .A(n1), .Z(\sa_count[9][51] ));
Q_BUF U769 ( .A(n1), .Z(\sa_count[9][50] ));
Q_BUF U770 ( .A(n1), .Z(\sa_count[8][63] ));
Q_BUF U771 ( .A(n1), .Z(\sa_count[8][62] ));
Q_BUF U772 ( .A(n1), .Z(\sa_count[8][61] ));
Q_BUF U773 ( .A(n1), .Z(\sa_count[8][60] ));
Q_BUF U774 ( .A(n1), .Z(\sa_count[8][59] ));
Q_BUF U775 ( .A(n1), .Z(\sa_count[8][58] ));
Q_BUF U776 ( .A(n1), .Z(\sa_count[8][57] ));
Q_BUF U777 ( .A(n1), .Z(\sa_count[8][56] ));
Q_BUF U778 ( .A(n1), .Z(\sa_count[8][55] ));
Q_BUF U779 ( .A(n1), .Z(\sa_count[8][54] ));
Q_BUF U780 ( .A(n1), .Z(\sa_count[8][53] ));
Q_BUF U781 ( .A(n1), .Z(\sa_count[8][52] ));
Q_BUF U782 ( .A(n1), .Z(\sa_count[8][51] ));
Q_BUF U783 ( .A(n1), .Z(\sa_count[8][50] ));
Q_BUF U784 ( .A(n1), .Z(\sa_count[7][63] ));
Q_BUF U785 ( .A(n1), .Z(\sa_count[7][62] ));
Q_BUF U786 ( .A(n1), .Z(\sa_count[7][61] ));
Q_BUF U787 ( .A(n1), .Z(\sa_count[7][60] ));
Q_BUF U788 ( .A(n1), .Z(\sa_count[7][59] ));
Q_BUF U789 ( .A(n1), .Z(\sa_count[7][58] ));
Q_BUF U790 ( .A(n1), .Z(\sa_count[7][57] ));
Q_BUF U791 ( .A(n1), .Z(\sa_count[7][56] ));
Q_BUF U792 ( .A(n1), .Z(\sa_count[7][55] ));
Q_BUF U793 ( .A(n1), .Z(\sa_count[7][54] ));
Q_BUF U794 ( .A(n1), .Z(\sa_count[7][53] ));
Q_BUF U795 ( .A(n1), .Z(\sa_count[7][52] ));
Q_BUF U796 ( .A(n1), .Z(\sa_count[7][51] ));
Q_BUF U797 ( .A(n1), .Z(\sa_count[7][50] ));
Q_BUF U798 ( .A(n1), .Z(\sa_count[6][63] ));
Q_BUF U799 ( .A(n1), .Z(\sa_count[6][62] ));
Q_BUF U800 ( .A(n1), .Z(\sa_count[6][61] ));
Q_BUF U801 ( .A(n1), .Z(\sa_count[6][60] ));
Q_BUF U802 ( .A(n1), .Z(\sa_count[6][59] ));
Q_BUF U803 ( .A(n1), .Z(\sa_count[6][58] ));
Q_BUF U804 ( .A(n1), .Z(\sa_count[6][57] ));
Q_BUF U805 ( .A(n1), .Z(\sa_count[6][56] ));
Q_BUF U806 ( .A(n1), .Z(\sa_count[6][55] ));
Q_BUF U807 ( .A(n1), .Z(\sa_count[6][54] ));
Q_BUF U808 ( .A(n1), .Z(\sa_count[6][53] ));
Q_BUF U809 ( .A(n1), .Z(\sa_count[6][52] ));
Q_BUF U810 ( .A(n1), .Z(\sa_count[6][51] ));
Q_BUF U811 ( .A(n1), .Z(\sa_count[6][50] ));
Q_BUF U812 ( .A(n1), .Z(\sa_count[5][63] ));
Q_BUF U813 ( .A(n1), .Z(\sa_count[5][62] ));
Q_BUF U814 ( .A(n1), .Z(\sa_count[5][61] ));
Q_BUF U815 ( .A(n1), .Z(\sa_count[5][60] ));
Q_BUF U816 ( .A(n1), .Z(\sa_count[5][59] ));
Q_BUF U817 ( .A(n1), .Z(\sa_count[5][58] ));
Q_BUF U818 ( .A(n1), .Z(\sa_count[5][57] ));
Q_BUF U819 ( .A(n1), .Z(\sa_count[5][56] ));
Q_BUF U820 ( .A(n1), .Z(\sa_count[5][55] ));
Q_BUF U821 ( .A(n1), .Z(\sa_count[5][54] ));
Q_BUF U822 ( .A(n1), .Z(\sa_count[5][53] ));
Q_BUF U823 ( .A(n1), .Z(\sa_count[5][52] ));
Q_BUF U824 ( .A(n1), .Z(\sa_count[5][51] ));
Q_BUF U825 ( .A(n1), .Z(\sa_count[5][50] ));
Q_BUF U826 ( .A(n1), .Z(\sa_count[4][63] ));
Q_BUF U827 ( .A(n1), .Z(\sa_count[4][62] ));
Q_BUF U828 ( .A(n1), .Z(\sa_count[4][61] ));
Q_BUF U829 ( .A(n1), .Z(\sa_count[4][60] ));
Q_BUF U830 ( .A(n1), .Z(\sa_count[4][59] ));
Q_BUF U831 ( .A(n1), .Z(\sa_count[4][58] ));
Q_BUF U832 ( .A(n1), .Z(\sa_count[4][57] ));
Q_BUF U833 ( .A(n1), .Z(\sa_count[4][56] ));
Q_BUF U834 ( .A(n1), .Z(\sa_count[4][55] ));
Q_BUF U835 ( .A(n1), .Z(\sa_count[4][54] ));
Q_BUF U836 ( .A(n1), .Z(\sa_count[4][53] ));
Q_BUF U837 ( .A(n1), .Z(\sa_count[4][52] ));
Q_BUF U838 ( .A(n1), .Z(\sa_count[4][51] ));
Q_BUF U839 ( .A(n1), .Z(\sa_count[4][50] ));
Q_BUF U840 ( .A(n1), .Z(\sa_count[3][63] ));
Q_BUF U841 ( .A(n1), .Z(\sa_count[3][62] ));
Q_BUF U842 ( .A(n1), .Z(\sa_count[3][61] ));
Q_BUF U843 ( .A(n1), .Z(\sa_count[3][60] ));
Q_BUF U844 ( .A(n1), .Z(\sa_count[3][59] ));
Q_BUF U845 ( .A(n1), .Z(\sa_count[3][58] ));
Q_BUF U846 ( .A(n1), .Z(\sa_count[3][57] ));
Q_BUF U847 ( .A(n1), .Z(\sa_count[3][56] ));
Q_BUF U848 ( .A(n1), .Z(\sa_count[3][55] ));
Q_BUF U849 ( .A(n1), .Z(\sa_count[3][54] ));
Q_BUF U850 ( .A(n1), .Z(\sa_count[3][53] ));
Q_BUF U851 ( .A(n1), .Z(\sa_count[3][52] ));
Q_BUF U852 ( .A(n1), .Z(\sa_count[3][51] ));
Q_BUF U853 ( .A(n1), .Z(\sa_count[3][50] ));
Q_BUF U854 ( .A(n1), .Z(\sa_count[2][63] ));
Q_BUF U855 ( .A(n1), .Z(\sa_count[2][62] ));
Q_BUF U856 ( .A(n1), .Z(\sa_count[2][61] ));
Q_BUF U857 ( .A(n1), .Z(\sa_count[2][60] ));
Q_BUF U858 ( .A(n1), .Z(\sa_count[2][59] ));
Q_BUF U859 ( .A(n1), .Z(\sa_count[2][58] ));
Q_BUF U860 ( .A(n1), .Z(\sa_count[2][57] ));
Q_BUF U861 ( .A(n1), .Z(\sa_count[2][56] ));
Q_BUF U862 ( .A(n1), .Z(\sa_count[2][55] ));
Q_BUF U863 ( .A(n1), .Z(\sa_count[2][54] ));
Q_BUF U864 ( .A(n1), .Z(\sa_count[2][53] ));
Q_BUF U865 ( .A(n1), .Z(\sa_count[2][52] ));
Q_BUF U866 ( .A(n1), .Z(\sa_count[2][51] ));
Q_BUF U867 ( .A(n1), .Z(\sa_count[2][50] ));
Q_BUF U868 ( .A(n1), .Z(\sa_count[1][63] ));
Q_BUF U869 ( .A(n1), .Z(\sa_count[1][62] ));
Q_BUF U870 ( .A(n1), .Z(\sa_count[1][61] ));
Q_BUF U871 ( .A(n1), .Z(\sa_count[1][60] ));
Q_BUF U872 ( .A(n1), .Z(\sa_count[1][59] ));
Q_BUF U873 ( .A(n1), .Z(\sa_count[1][58] ));
Q_BUF U874 ( .A(n1), .Z(\sa_count[1][57] ));
Q_BUF U875 ( .A(n1), .Z(\sa_count[1][56] ));
Q_BUF U876 ( .A(n1), .Z(\sa_count[1][55] ));
Q_BUF U877 ( .A(n1), .Z(\sa_count[1][54] ));
Q_BUF U878 ( .A(n1), .Z(\sa_count[1][53] ));
Q_BUF U879 ( .A(n1), .Z(\sa_count[1][52] ));
Q_BUF U880 ( .A(n1), .Z(\sa_count[1][51] ));
Q_BUF U881 ( .A(n1), .Z(\sa_count[1][50] ));
Q_BUF U882 ( .A(n1), .Z(\sa_count[0][63] ));
Q_BUF U883 ( .A(n1), .Z(\sa_count[0][62] ));
Q_BUF U884 ( .A(n1), .Z(\sa_count[0][61] ));
Q_BUF U885 ( .A(n1), .Z(\sa_count[0][60] ));
Q_BUF U886 ( .A(n1), .Z(\sa_count[0][59] ));
Q_BUF U887 ( .A(n1), .Z(\sa_count[0][58] ));
Q_BUF U888 ( .A(n1), .Z(\sa_count[0][57] ));
Q_BUF U889 ( .A(n1), .Z(\sa_count[0][56] ));
Q_BUF U890 ( .A(n1), .Z(\sa_count[0][55] ));
Q_BUF U891 ( .A(n1), .Z(\sa_count[0][54] ));
Q_BUF U892 ( .A(n1), .Z(\sa_count[0][53] ));
Q_BUF U893 ( .A(n1), .Z(\sa_count[0][52] ));
Q_BUF U894 ( .A(n1), .Z(\sa_count[0][51] ));
Q_BUF U895 ( .A(n1), .Z(\sa_count[0][50] ));
Q_BUF U896 ( .A(n1), .Z(\sa_events[0][63] ));
Q_BUF U897 ( .A(n1), .Z(\sa_events[0][62] ));
Q_BUF U898 ( .A(n1), .Z(\sa_events[0][61] ));
Q_BUF U899 ( .A(n1), .Z(\sa_events[0][60] ));
Q_BUF U900 ( .A(n1), .Z(\sa_events[0][59] ));
Q_BUF U901 ( .A(n1), .Z(\sa_events[0][58] ));
Q_BUF U902 ( .A(n1), .Z(\sa_events[0][57] ));
Q_BUF U903 ( .A(n1), .Z(\sa_events[0][56] ));
Q_BUF U904 ( .A(n1), .Z(\sa_events[0][55] ));
Q_BUF U905 ( .A(n1), .Z(\sa_events[0][54] ));
Q_BUF U906 ( .A(n1), .Z(\sa_events[0][53] ));
Q_BUF U907 ( .A(n1), .Z(\sa_events[0][52] ));
Q_BUF U908 ( .A(n1), .Z(\sa_events[0][51] ));
Q_BUF U909 ( .A(n1), .Z(\sa_events[0][50] ));
Q_BUF U910 ( .A(n1), .Z(\sa_events[0][49] ));
Q_BUF U911 ( .A(n1), .Z(\sa_events[0][48] ));
Q_BUF U912 ( .A(n1), .Z(\sa_events[0][47] ));
Q_BUF U913 ( .A(n1), .Z(\sa_events[0][46] ));
Q_BUF U914 ( .A(n1), .Z(\sa_events[0][45] ));
Q_BUF U915 ( .A(n1), .Z(\sa_events[0][44] ));
Q_BUF U916 ( .A(n1), .Z(\sa_events[0][43] ));
Q_BUF U917 ( .A(n1), .Z(\sa_events[0][42] ));
Q_BUF U918 ( .A(n1), .Z(\sa_events[0][41] ));
Q_BUF U919 ( .A(n1), .Z(\sa_events[0][40] ));
Q_BUF U920 ( .A(n1), .Z(\sa_events[0][39] ));
Q_BUF U921 ( .A(n1), .Z(\sa_events[0][38] ));
Q_BUF U922 ( .A(n1), .Z(\sa_events[0][37] ));
Q_BUF U923 ( .A(n1), .Z(\sa_events[0][36] ));
Q_BUF U924 ( .A(n1), .Z(\sa_events[0][35] ));
Q_BUF U925 ( .A(n1), .Z(\sa_events[0][34] ));
Q_BUF U926 ( .A(n1), .Z(\sa_events[0][33] ));
Q_BUF U927 ( .A(n1), .Z(\sa_events[0][32] ));
Q_BUF U928 ( .A(n1), .Z(\sa_events[0][31] ));
Q_BUF U929 ( .A(n1), .Z(\sa_events[0][30] ));
Q_BUF U930 ( .A(n1), .Z(\sa_events[0][29] ));
Q_BUF U931 ( .A(n1), .Z(\sa_events[0][28] ));
Q_BUF U932 ( .A(n1), .Z(\sa_events[0][27] ));
Q_BUF U933 ( .A(n1), .Z(\sa_events[0][26] ));
Q_BUF U934 ( .A(n1), .Z(\sa_events[0][25] ));
Q_BUF U935 ( .A(n1), .Z(\sa_events[1][63] ));
Q_BUF U936 ( .A(n1), .Z(\sa_events[1][62] ));
Q_BUF U937 ( .A(n1), .Z(\sa_events[1][61] ));
Q_BUF U938 ( .A(n1), .Z(\sa_events[1][60] ));
Q_BUF U939 ( .A(n1), .Z(\sa_events[1][59] ));
Q_BUF U940 ( .A(n1), .Z(\sa_events[1][58] ));
Q_BUF U941 ( .A(n1), .Z(\sa_events[1][57] ));
Q_BUF U942 ( .A(n1), .Z(\sa_events[1][56] ));
Q_BUF U943 ( .A(n1), .Z(\sa_events[1][55] ));
Q_BUF U944 ( .A(n1), .Z(\sa_events[1][54] ));
Q_BUF U945 ( .A(n1), .Z(\sa_events[1][53] ));
Q_BUF U946 ( .A(n1), .Z(\sa_events[1][52] ));
Q_BUF U947 ( .A(n1), .Z(\sa_events[1][51] ));
Q_BUF U948 ( .A(n1), .Z(\sa_events[1][50] ));
Q_BUF U949 ( .A(n1), .Z(\sa_events[1][49] ));
Q_BUF U950 ( .A(n1), .Z(\sa_events[1][48] ));
Q_BUF U951 ( .A(n1), .Z(\sa_events[1][47] ));
Q_BUF U952 ( .A(n1), .Z(\sa_events[1][46] ));
Q_BUF U953 ( .A(n1), .Z(\sa_events[1][45] ));
Q_BUF U954 ( .A(n1), .Z(\sa_events[1][44] ));
Q_BUF U955 ( .A(n1), .Z(\sa_events[1][43] ));
Q_BUF U956 ( .A(n1), .Z(\sa_events[1][42] ));
Q_BUF U957 ( .A(n1), .Z(\sa_events[1][41] ));
Q_BUF U958 ( .A(n1), .Z(\sa_events[1][40] ));
Q_BUF U959 ( .A(n1), .Z(\sa_events[1][39] ));
Q_BUF U960 ( .A(n1), .Z(\sa_events[1][38] ));
Q_BUF U961 ( .A(n1), .Z(\sa_events[1][37] ));
Q_BUF U962 ( .A(n1), .Z(\sa_events[1][36] ));
Q_BUF U963 ( .A(n1), .Z(\sa_events[1][35] ));
Q_BUF U964 ( .A(n1), .Z(\sa_events[1][34] ));
Q_BUF U965 ( .A(n1), .Z(\sa_events[1][33] ));
Q_BUF U966 ( .A(n1), .Z(\sa_events[1][32] ));
Q_BUF U967 ( .A(n1), .Z(\sa_events[1][31] ));
Q_BUF U968 ( .A(n1), .Z(\sa_events[1][30] ));
Q_BUF U969 ( .A(n1), .Z(\sa_events[1][29] ));
Q_BUF U970 ( .A(n1), .Z(\sa_events[1][28] ));
Q_BUF U971 ( .A(n1), .Z(\sa_events[1][27] ));
Q_BUF U972 ( .A(n1), .Z(\sa_events[1][26] ));
Q_BUF U973 ( .A(n1), .Z(\sa_events[1][25] ));
Q_BUF U974 ( .A(n1), .Z(\sa_events[1][24] ));
Q_BUF U975 ( .A(n1), .Z(\sa_events[1][23] ));
Q_BUF U976 ( .A(n1), .Z(\sa_events[1][22] ));
Q_BUF U977 ( .A(n1), .Z(\sa_events[1][21] ));
Q_BUF U978 ( .A(n1), .Z(\sa_events[1][20] ));
Q_BUF U979 ( .A(n1), .Z(\sa_events[1][19] ));
Q_BUF U980 ( .A(n1), .Z(\sa_events[1][18] ));
Q_BUF U981 ( .A(n1), .Z(\sa_events[1][17] ));
Q_BUF U982 ( .A(n1), .Z(\sa_events[1][16] ));
Q_BUF U983 ( .A(n1), .Z(\sa_events[1][15] ));
Q_BUF U984 ( .A(n1), .Z(\sa_events[1][14] ));
Q_BUF U985 ( .A(n1), .Z(\sa_events[1][13] ));
Q_BUF U986 ( .A(n1), .Z(\sa_events[1][12] ));
Q_BUF U987 ( .A(n1), .Z(\sa_events[1][11] ));
Q_BUF U988 ( .A(n1), .Z(\sa_events[1][10] ));
Q_BUF U989 ( .A(n1), .Z(\sa_events[1][9] ));
Q_BUF U990 ( .A(n1), .Z(\sa_events[1][8] ));
Q_BUF U991 ( .A(n1), .Z(\sa_events[1][7] ));
Q_BUF U992 ( .A(n1), .Z(\sa_events[1][6] ));
Q_BUF U993 ( .A(n1), .Z(\sa_events[1][5] ));
Q_BUF U994 ( .A(n1), .Z(\sa_events[1][4] ));
Q_BUF U995 ( .A(n1), .Z(\sa_events[1][3] ));
Q_BUF U996 ( .A(n1), .Z(\sa_events[1][2] ));
Q_BUF U997 ( .A(n1), .Z(\sa_events[1][1] ));
Q_BUF U998 ( .A(n1), .Z(\sa_events[1][0] ));
Q_BUF U999 ( .A(n1), .Z(\sa_events[2][63] ));
Q_BUF U1000 ( .A(n1), .Z(\sa_events[2][62] ));
Q_BUF U1001 ( .A(n1), .Z(\sa_events[2][61] ));
Q_BUF U1002 ( .A(n1), .Z(\sa_events[2][60] ));
Q_BUF U1003 ( .A(n1), .Z(\sa_events[2][59] ));
Q_BUF U1004 ( .A(n1), .Z(\sa_events[2][58] ));
Q_BUF U1005 ( .A(n1), .Z(\sa_events[2][57] ));
Q_BUF U1006 ( .A(n1), .Z(\sa_events[2][56] ));
Q_BUF U1007 ( .A(n1), .Z(\sa_events[2][55] ));
Q_BUF U1008 ( .A(n1), .Z(\sa_events[2][54] ));
Q_BUF U1009 ( .A(n1), .Z(\sa_events[2][53] ));
Q_BUF U1010 ( .A(n1), .Z(\sa_events[2][52] ));
Q_BUF U1011 ( .A(n1), .Z(\sa_events[2][51] ));
Q_BUF U1012 ( .A(n1), .Z(\sa_events[2][50] ));
Q_BUF U1013 ( .A(n1), .Z(\sa_events[2][49] ));
Q_BUF U1014 ( .A(n1), .Z(\sa_events[2][48] ));
Q_BUF U1015 ( .A(n1), .Z(\sa_events[2][47] ));
Q_BUF U1016 ( .A(n1), .Z(\sa_events[2][46] ));
Q_BUF U1017 ( .A(n1), .Z(\sa_events[2][45] ));
Q_BUF U1018 ( .A(n1), .Z(\sa_events[2][44] ));
Q_BUF U1019 ( .A(n1), .Z(\sa_events[2][43] ));
Q_BUF U1020 ( .A(n1), .Z(\sa_events[2][42] ));
Q_BUF U1021 ( .A(n1), .Z(\sa_events[2][41] ));
Q_BUF U1022 ( .A(n1), .Z(\sa_events[2][40] ));
Q_BUF U1023 ( .A(n1), .Z(\sa_events[2][39] ));
Q_BUF U1024 ( .A(n1), .Z(\sa_events[2][38] ));
Q_BUF U1025 ( .A(n1), .Z(\sa_events[2][37] ));
Q_BUF U1026 ( .A(n1), .Z(\sa_events[2][36] ));
Q_BUF U1027 ( .A(n1), .Z(\sa_events[2][35] ));
Q_BUF U1028 ( .A(n1), .Z(\sa_events[2][34] ));
Q_BUF U1029 ( .A(n1), .Z(\sa_events[2][33] ));
Q_BUF U1030 ( .A(n1), .Z(\sa_events[2][32] ));
Q_BUF U1031 ( .A(n1), .Z(\sa_events[2][31] ));
Q_BUF U1032 ( .A(n1), .Z(\sa_events[2][30] ));
Q_BUF U1033 ( .A(n1), .Z(\sa_events[2][29] ));
Q_BUF U1034 ( .A(n1), .Z(\sa_events[2][28] ));
Q_BUF U1035 ( .A(n1), .Z(\sa_events[2][27] ));
Q_BUF U1036 ( .A(n1), .Z(\sa_events[2][26] ));
Q_BUF U1037 ( .A(n1), .Z(\sa_events[2][25] ));
Q_BUF U1038 ( .A(n1), .Z(\sa_events[2][24] ));
Q_BUF U1039 ( .A(n1), .Z(\sa_events[2][23] ));
Q_BUF U1040 ( .A(n1), .Z(\sa_events[2][22] ));
Q_BUF U1041 ( .A(n1), .Z(\sa_events[2][21] ));
Q_BUF U1042 ( .A(n1), .Z(\sa_events[2][20] ));
Q_BUF U1043 ( .A(n1), .Z(\sa_events[2][19] ));
Q_BUF U1044 ( .A(n1), .Z(\sa_events[2][18] ));
Q_BUF U1045 ( .A(n1), .Z(\sa_events[2][17] ));
Q_BUF U1046 ( .A(n1), .Z(\sa_events[2][16] ));
Q_BUF U1047 ( .A(n1), .Z(\sa_events[2][15] ));
Q_BUF U1048 ( .A(n1), .Z(\sa_events[2][14] ));
Q_BUF U1049 ( .A(n1), .Z(\sa_events[2][13] ));
Q_BUF U1050 ( .A(n1), .Z(\sa_events[2][12] ));
Q_BUF U1051 ( .A(n1), .Z(\sa_events[2][11] ));
Q_BUF U1052 ( .A(n1), .Z(\sa_events[2][10] ));
Q_BUF U1053 ( .A(n1), .Z(\sa_events[2][9] ));
Q_BUF U1054 ( .A(n1), .Z(\sa_events[2][8] ));
Q_BUF U1055 ( .A(n1), .Z(\sa_events[2][7] ));
Q_BUF U1056 ( .A(n1), .Z(\sa_events[2][6] ));
Q_BUF U1057 ( .A(n1), .Z(\sa_events[2][5] ));
Q_BUF U1058 ( .A(n1), .Z(\sa_events[2][4] ));
Q_BUF U1059 ( .A(n1), .Z(\sa_events[2][3] ));
Q_BUF U1060 ( .A(n1), .Z(\sa_events[2][2] ));
Q_BUF U1061 ( .A(n1), .Z(\sa_events[2][1] ));
Q_BUF U1062 ( .A(n1), .Z(\sa_events[2][0] ));
Q_BUF U1063 ( .A(n1), .Z(\sa_events[3][63] ));
Q_BUF U1064 ( .A(n1), .Z(\sa_events[3][62] ));
Q_BUF U1065 ( .A(n1), .Z(\sa_events[3][61] ));
Q_BUF U1066 ( .A(n1), .Z(\sa_events[3][60] ));
Q_BUF U1067 ( .A(n1), .Z(\sa_events[3][59] ));
Q_BUF U1068 ( .A(n1), .Z(\sa_events[3][58] ));
Q_BUF U1069 ( .A(n1), .Z(\sa_events[3][57] ));
Q_BUF U1070 ( .A(n1), .Z(\sa_events[3][56] ));
Q_BUF U1071 ( .A(n1), .Z(\sa_events[3][55] ));
Q_BUF U1072 ( .A(n1), .Z(\sa_events[3][54] ));
Q_BUF U1073 ( .A(n1), .Z(\sa_events[3][53] ));
Q_BUF U1074 ( .A(n1), .Z(\sa_events[3][52] ));
Q_BUF U1075 ( .A(n1), .Z(\sa_events[3][51] ));
Q_BUF U1076 ( .A(n1), .Z(\sa_events[3][50] ));
Q_BUF U1077 ( .A(n1), .Z(\sa_events[3][49] ));
Q_BUF U1078 ( .A(n1), .Z(\sa_events[3][48] ));
Q_BUF U1079 ( .A(n1), .Z(\sa_events[3][47] ));
Q_BUF U1080 ( .A(n1), .Z(\sa_events[3][46] ));
Q_BUF U1081 ( .A(n1), .Z(\sa_events[3][45] ));
Q_BUF U1082 ( .A(n1), .Z(\sa_events[3][44] ));
Q_BUF U1083 ( .A(n1), .Z(\sa_events[3][43] ));
Q_BUF U1084 ( .A(n1), .Z(\sa_events[3][42] ));
Q_BUF U1085 ( .A(n1), .Z(\sa_events[3][41] ));
Q_BUF U1086 ( .A(n1), .Z(\sa_events[3][40] ));
Q_BUF U1087 ( .A(n1), .Z(\sa_events[3][39] ));
Q_BUF U1088 ( .A(n1), .Z(\sa_events[3][38] ));
Q_BUF U1089 ( .A(n1), .Z(\sa_events[3][37] ));
Q_BUF U1090 ( .A(n1), .Z(\sa_events[3][36] ));
Q_BUF U1091 ( .A(n1), .Z(\sa_events[3][35] ));
Q_BUF U1092 ( .A(n1), .Z(\sa_events[3][34] ));
Q_BUF U1093 ( .A(n1), .Z(\sa_events[3][33] ));
Q_BUF U1094 ( .A(n1), .Z(\sa_events[3][32] ));
Q_BUF U1095 ( .A(n1), .Z(\sa_events[3][31] ));
Q_BUF U1096 ( .A(n1), .Z(\sa_events[3][30] ));
Q_BUF U1097 ( .A(n1), .Z(\sa_events[3][29] ));
Q_BUF U1098 ( .A(n1), .Z(\sa_events[3][28] ));
Q_BUF U1099 ( .A(n1), .Z(\sa_events[3][27] ));
Q_BUF U1100 ( .A(n1), .Z(\sa_events[3][26] ));
Q_BUF U1101 ( .A(n1), .Z(\sa_events[3][25] ));
Q_BUF U1102 ( .A(n1), .Z(\sa_events[3][24] ));
Q_BUF U1103 ( .A(n1), .Z(\sa_events[3][23] ));
Q_BUF U1104 ( .A(n1), .Z(\sa_events[3][22] ));
Q_BUF U1105 ( .A(n1), .Z(\sa_events[3][21] ));
Q_BUF U1106 ( .A(n1), .Z(\sa_events[3][20] ));
Q_BUF U1107 ( .A(n1), .Z(\sa_events[3][19] ));
Q_BUF U1108 ( .A(n1), .Z(\sa_events[3][18] ));
Q_BUF U1109 ( .A(n1), .Z(\sa_events[3][17] ));
Q_BUF U1110 ( .A(n1), .Z(\sa_events[3][16] ));
Q_BUF U1111 ( .A(n1), .Z(\sa_events[3][15] ));
Q_BUF U1112 ( .A(n1), .Z(\sa_events[3][14] ));
Q_BUF U1113 ( .A(n1), .Z(\sa_events[3][13] ));
Q_BUF U1114 ( .A(n1), .Z(\sa_events[3][12] ));
Q_BUF U1115 ( .A(n1), .Z(\sa_events[3][11] ));
Q_BUF U1116 ( .A(n1), .Z(\sa_events[3][10] ));
Q_BUF U1117 ( .A(n1), .Z(\sa_events[3][9] ));
Q_BUF U1118 ( .A(n1), .Z(\sa_events[3][8] ));
Q_BUF U1119 ( .A(n1), .Z(\sa_events[3][7] ));
Q_BUF U1120 ( .A(n1), .Z(\sa_events[3][6] ));
Q_BUF U1121 ( .A(n1), .Z(\sa_events[3][5] ));
Q_BUF U1122 ( .A(n1), .Z(\sa_events[3][4] ));
Q_BUF U1123 ( .A(n1), .Z(\sa_events[3][3] ));
Q_BUF U1124 ( .A(n1), .Z(\sa_events[3][2] ));
Q_BUF U1125 ( .A(n1), .Z(\sa_events[3][1] ));
Q_BUF U1126 ( .A(n1), .Z(\sa_events[3][0] ));
Q_BUF U1127 ( .A(n1), .Z(\sa_events[4][63] ));
Q_BUF U1128 ( .A(n1), .Z(\sa_events[4][62] ));
Q_BUF U1129 ( .A(n1), .Z(\sa_events[4][61] ));
Q_BUF U1130 ( .A(n1), .Z(\sa_events[4][60] ));
Q_BUF U1131 ( .A(n1), .Z(\sa_events[4][59] ));
Q_BUF U1132 ( .A(n1), .Z(\sa_events[4][58] ));
Q_BUF U1133 ( .A(n1), .Z(\sa_events[4][57] ));
Q_BUF U1134 ( .A(n1), .Z(\sa_events[4][56] ));
Q_BUF U1135 ( .A(n1), .Z(\sa_events[4][55] ));
Q_BUF U1136 ( .A(n1), .Z(\sa_events[4][54] ));
Q_BUF U1137 ( .A(n1), .Z(\sa_events[4][53] ));
Q_BUF U1138 ( .A(n1), .Z(\sa_events[4][52] ));
Q_BUF U1139 ( .A(n1), .Z(\sa_events[4][51] ));
Q_BUF U1140 ( .A(n1), .Z(\sa_events[4][50] ));
Q_BUF U1141 ( .A(n1), .Z(\sa_events[4][49] ));
Q_BUF U1142 ( .A(n1), .Z(\sa_events[4][48] ));
Q_BUF U1143 ( .A(n1), .Z(\sa_events[4][47] ));
Q_BUF U1144 ( .A(n1), .Z(\sa_events[4][46] ));
Q_BUF U1145 ( .A(n1), .Z(\sa_events[4][45] ));
Q_BUF U1146 ( .A(n1), .Z(\sa_events[4][44] ));
Q_BUF U1147 ( .A(n1), .Z(\sa_events[4][43] ));
Q_BUF U1148 ( .A(n1), .Z(\sa_events[4][42] ));
Q_BUF U1149 ( .A(n1), .Z(\sa_events[4][41] ));
Q_BUF U1150 ( .A(n1), .Z(\sa_events[4][40] ));
Q_BUF U1151 ( .A(n1), .Z(\sa_events[4][39] ));
Q_BUF U1152 ( .A(n1), .Z(\sa_events[4][38] ));
Q_BUF U1153 ( .A(n1), .Z(\sa_events[4][37] ));
Q_BUF U1154 ( .A(n1), .Z(\sa_events[4][36] ));
Q_BUF U1155 ( .A(n1), .Z(\sa_events[4][35] ));
Q_BUF U1156 ( .A(n1), .Z(\sa_events[4][34] ));
Q_BUF U1157 ( .A(n1), .Z(\sa_events[4][33] ));
Q_BUF U1158 ( .A(n1), .Z(\sa_events[4][32] ));
Q_BUF U1159 ( .A(n1), .Z(\sa_events[4][31] ));
Q_BUF U1160 ( .A(n1), .Z(\sa_events[4][30] ));
Q_BUF U1161 ( .A(n1), .Z(\sa_events[4][29] ));
Q_BUF U1162 ( .A(n1), .Z(\sa_events[4][28] ));
Q_BUF U1163 ( .A(n1), .Z(\sa_events[4][27] ));
Q_BUF U1164 ( .A(n1), .Z(\sa_events[4][26] ));
Q_BUF U1165 ( .A(n1), .Z(\sa_events[4][25] ));
Q_BUF U1166 ( .A(n1), .Z(\sa_events[4][24] ));
Q_BUF U1167 ( .A(n1), .Z(\sa_events[4][23] ));
Q_BUF U1168 ( .A(n1), .Z(\sa_events[4][22] ));
Q_BUF U1169 ( .A(n1), .Z(\sa_events[4][21] ));
Q_BUF U1170 ( .A(n1), .Z(\sa_events[4][20] ));
Q_BUF U1171 ( .A(n1), .Z(\sa_events[4][19] ));
Q_BUF U1172 ( .A(n1), .Z(\sa_events[4][18] ));
Q_BUF U1173 ( .A(n1), .Z(\sa_events[4][17] ));
Q_BUF U1174 ( .A(n1), .Z(\sa_events[4][16] ));
Q_BUF U1175 ( .A(n1), .Z(\sa_events[4][15] ));
Q_BUF U1176 ( .A(n1), .Z(\sa_events[4][14] ));
Q_BUF U1177 ( .A(n1), .Z(\sa_events[4][13] ));
Q_BUF U1178 ( .A(n1), .Z(\sa_events[4][12] ));
Q_BUF U1179 ( .A(n1), .Z(\sa_events[4][11] ));
Q_BUF U1180 ( .A(n1), .Z(\sa_events[4][10] ));
Q_BUF U1181 ( .A(n1), .Z(\sa_events[4][9] ));
Q_BUF U1182 ( .A(n1), .Z(\sa_events[4][8] ));
Q_BUF U1183 ( .A(n1), .Z(\sa_events[4][7] ));
Q_BUF U1184 ( .A(n1), .Z(\sa_events[4][6] ));
Q_BUF U1185 ( .A(n1), .Z(\sa_events[4][5] ));
Q_BUF U1186 ( .A(n1), .Z(\sa_events[4][4] ));
Q_BUF U1187 ( .A(n1), .Z(\sa_events[4][3] ));
Q_BUF U1188 ( .A(n1), .Z(\sa_events[4][2] ));
Q_BUF U1189 ( .A(n1), .Z(\sa_events[4][1] ));
Q_BUF U1190 ( .A(n1), .Z(\sa_events[4][0] ));
Q_BUF U1191 ( .A(n1), .Z(\sa_events[5][63] ));
Q_BUF U1192 ( .A(n1), .Z(\sa_events[5][62] ));
Q_BUF U1193 ( .A(n1), .Z(\sa_events[5][61] ));
Q_BUF U1194 ( .A(n1), .Z(\sa_events[5][60] ));
Q_BUF U1195 ( .A(n1), .Z(\sa_events[5][59] ));
Q_BUF U1196 ( .A(n1), .Z(\sa_events[5][58] ));
Q_BUF U1197 ( .A(n1), .Z(\sa_events[5][57] ));
Q_BUF U1198 ( .A(n1), .Z(\sa_events[5][56] ));
Q_BUF U1199 ( .A(n1), .Z(\sa_events[5][55] ));
Q_BUF U1200 ( .A(n1), .Z(\sa_events[5][54] ));
Q_BUF U1201 ( .A(n1), .Z(\sa_events[5][53] ));
Q_BUF U1202 ( .A(n1), .Z(\sa_events[5][52] ));
Q_BUF U1203 ( .A(n1), .Z(\sa_events[5][51] ));
Q_BUF U1204 ( .A(n1), .Z(\sa_events[5][50] ));
Q_BUF U1205 ( .A(n1), .Z(\sa_events[5][49] ));
Q_BUF U1206 ( .A(n1), .Z(\sa_events[5][48] ));
Q_BUF U1207 ( .A(n1), .Z(\sa_events[5][47] ));
Q_BUF U1208 ( .A(n1), .Z(\sa_events[5][46] ));
Q_BUF U1209 ( .A(n1), .Z(\sa_events[5][45] ));
Q_BUF U1210 ( .A(n1), .Z(\sa_events[5][44] ));
Q_BUF U1211 ( .A(n1), .Z(\sa_events[5][43] ));
Q_BUF U1212 ( .A(n1), .Z(\sa_events[5][42] ));
Q_BUF U1213 ( .A(n1), .Z(\sa_events[5][41] ));
Q_BUF U1214 ( .A(n1), .Z(\sa_events[5][40] ));
Q_BUF U1215 ( .A(n1), .Z(\sa_events[5][39] ));
Q_BUF U1216 ( .A(n1), .Z(\sa_events[5][38] ));
Q_BUF U1217 ( .A(n1), .Z(\sa_events[5][37] ));
Q_BUF U1218 ( .A(n1), .Z(\sa_events[5][36] ));
Q_BUF U1219 ( .A(n1), .Z(\sa_events[5][35] ));
Q_BUF U1220 ( .A(n1), .Z(\sa_events[5][34] ));
Q_BUF U1221 ( .A(n1), .Z(\sa_events[5][33] ));
Q_BUF U1222 ( .A(n1), .Z(\sa_events[5][32] ));
Q_BUF U1223 ( .A(n1), .Z(\sa_events[5][31] ));
Q_BUF U1224 ( .A(n1), .Z(\sa_events[5][30] ));
Q_BUF U1225 ( .A(n1), .Z(\sa_events[5][29] ));
Q_BUF U1226 ( .A(n1), .Z(\sa_events[5][28] ));
Q_BUF U1227 ( .A(n1), .Z(\sa_events[5][27] ));
Q_BUF U1228 ( .A(n1), .Z(\sa_events[5][26] ));
Q_BUF U1229 ( .A(n1), .Z(\sa_events[5][25] ));
Q_BUF U1230 ( .A(n1), .Z(\sa_events[5][24] ));
Q_BUF U1231 ( .A(n1), .Z(\sa_events[5][23] ));
Q_BUF U1232 ( .A(n1), .Z(\sa_events[5][22] ));
Q_BUF U1233 ( .A(n1), .Z(\sa_events[5][21] ));
Q_BUF U1234 ( .A(n1), .Z(\sa_events[5][20] ));
Q_BUF U1235 ( .A(n1), .Z(\sa_events[5][19] ));
Q_BUF U1236 ( .A(n1), .Z(\sa_events[5][18] ));
Q_BUF U1237 ( .A(n1), .Z(\sa_events[5][17] ));
Q_BUF U1238 ( .A(n1), .Z(\sa_events[5][16] ));
Q_BUF U1239 ( .A(n1), .Z(\sa_events[5][15] ));
Q_BUF U1240 ( .A(n1), .Z(\sa_events[5][14] ));
Q_BUF U1241 ( .A(n1), .Z(\sa_events[5][13] ));
Q_BUF U1242 ( .A(n1), .Z(\sa_events[5][12] ));
Q_BUF U1243 ( .A(n1), .Z(\sa_events[5][11] ));
Q_BUF U1244 ( .A(n1), .Z(\sa_events[5][10] ));
Q_BUF U1245 ( .A(n1), .Z(\sa_events[5][9] ));
Q_BUF U1246 ( .A(n1), .Z(\sa_events[5][8] ));
Q_BUF U1247 ( .A(n1), .Z(\sa_events[5][7] ));
Q_BUF U1248 ( .A(n1), .Z(\sa_events[5][6] ));
Q_BUF U1249 ( .A(n1), .Z(\sa_events[5][5] ));
Q_BUF U1250 ( .A(n1), .Z(\sa_events[5][4] ));
Q_BUF U1251 ( .A(n1), .Z(\sa_events[5][3] ));
Q_BUF U1252 ( .A(n1), .Z(\sa_events[5][2] ));
Q_BUF U1253 ( .A(n1), .Z(\sa_events[5][1] ));
Q_BUF U1254 ( .A(n1), .Z(\sa_events[5][0] ));
Q_BUF U1255 ( .A(n1), .Z(\sa_events[6][63] ));
Q_BUF U1256 ( .A(n1), .Z(\sa_events[6][62] ));
Q_BUF U1257 ( .A(n1), .Z(\sa_events[6][61] ));
Q_BUF U1258 ( .A(n1), .Z(\sa_events[6][60] ));
Q_BUF U1259 ( .A(n1), .Z(\sa_events[6][59] ));
Q_BUF U1260 ( .A(n1), .Z(\sa_events[6][58] ));
Q_BUF U1261 ( .A(n1), .Z(\sa_events[6][57] ));
Q_BUF U1262 ( .A(n1), .Z(\sa_events[6][56] ));
Q_BUF U1263 ( .A(n1), .Z(\sa_events[6][55] ));
Q_BUF U1264 ( .A(n1), .Z(\sa_events[6][54] ));
Q_BUF U1265 ( .A(n1), .Z(\sa_events[6][53] ));
Q_BUF U1266 ( .A(n1), .Z(\sa_events[6][52] ));
Q_BUF U1267 ( .A(n1), .Z(\sa_events[6][51] ));
Q_BUF U1268 ( .A(n1), .Z(\sa_events[6][50] ));
Q_BUF U1269 ( .A(n1), .Z(\sa_events[6][49] ));
Q_BUF U1270 ( .A(n1), .Z(\sa_events[6][48] ));
Q_BUF U1271 ( .A(n1), .Z(\sa_events[6][47] ));
Q_BUF U1272 ( .A(n1), .Z(\sa_events[6][46] ));
Q_BUF U1273 ( .A(n1), .Z(\sa_events[6][45] ));
Q_BUF U1274 ( .A(n1), .Z(\sa_events[6][44] ));
Q_BUF U1275 ( .A(n1), .Z(\sa_events[6][43] ));
Q_BUF U1276 ( .A(n1), .Z(\sa_events[6][42] ));
Q_BUF U1277 ( .A(n1), .Z(\sa_events[6][41] ));
Q_BUF U1278 ( .A(n1), .Z(\sa_events[6][40] ));
Q_BUF U1279 ( .A(n1), .Z(\sa_events[6][39] ));
Q_BUF U1280 ( .A(n1), .Z(\sa_events[6][38] ));
Q_BUF U1281 ( .A(n1), .Z(\sa_events[6][37] ));
Q_BUF U1282 ( .A(n1), .Z(\sa_events[6][36] ));
Q_BUF U1283 ( .A(n1), .Z(\sa_events[6][35] ));
Q_BUF U1284 ( .A(n1), .Z(\sa_events[6][34] ));
Q_BUF U1285 ( .A(n1), .Z(\sa_events[6][33] ));
Q_BUF U1286 ( .A(n1), .Z(\sa_events[6][32] ));
Q_BUF U1287 ( .A(n1), .Z(\sa_events[6][31] ));
Q_BUF U1288 ( .A(n1), .Z(\sa_events[6][30] ));
Q_BUF U1289 ( .A(n1), .Z(\sa_events[6][29] ));
Q_BUF U1290 ( .A(n1), .Z(\sa_events[6][28] ));
Q_BUF U1291 ( .A(n1), .Z(\sa_events[6][27] ));
Q_BUF U1292 ( .A(n1), .Z(\sa_events[6][26] ));
Q_BUF U1293 ( .A(n1), .Z(\sa_events[6][25] ));
Q_BUF U1294 ( .A(n1), .Z(\sa_events[6][24] ));
Q_BUF U1295 ( .A(n1), .Z(\sa_events[6][23] ));
Q_BUF U1296 ( .A(n1), .Z(\sa_events[6][22] ));
Q_BUF U1297 ( .A(n1), .Z(\sa_events[6][21] ));
Q_BUF U1298 ( .A(n1), .Z(\sa_events[6][20] ));
Q_BUF U1299 ( .A(n1), .Z(\sa_events[6][19] ));
Q_BUF U1300 ( .A(n1), .Z(\sa_events[6][18] ));
Q_BUF U1301 ( .A(n1), .Z(\sa_events[6][17] ));
Q_BUF U1302 ( .A(n1), .Z(\sa_events[6][16] ));
Q_BUF U1303 ( .A(n1), .Z(\sa_events[6][15] ));
Q_BUF U1304 ( .A(n1), .Z(\sa_events[6][14] ));
Q_BUF U1305 ( .A(n1), .Z(\sa_events[6][13] ));
Q_BUF U1306 ( .A(n1), .Z(\sa_events[6][12] ));
Q_BUF U1307 ( .A(n1), .Z(\sa_events[6][11] ));
Q_BUF U1308 ( .A(n1), .Z(\sa_events[6][10] ));
Q_BUF U1309 ( .A(n1), .Z(\sa_events[6][9] ));
Q_BUF U1310 ( .A(n1), .Z(\sa_events[6][8] ));
Q_BUF U1311 ( .A(n1), .Z(\sa_events[6][7] ));
Q_BUF U1312 ( .A(n1), .Z(\sa_events[6][6] ));
Q_BUF U1313 ( .A(n1), .Z(\sa_events[6][5] ));
Q_BUF U1314 ( .A(n1), .Z(\sa_events[6][4] ));
Q_BUF U1315 ( .A(n1), .Z(\sa_events[6][3] ));
Q_BUF U1316 ( .A(n1), .Z(\sa_events[6][2] ));
Q_BUF U1317 ( .A(n1), .Z(\sa_events[6][1] ));
Q_BUF U1318 ( .A(n1), .Z(\sa_events[6][0] ));
Q_BUF U1319 ( .A(n1), .Z(\sa_events[7][63] ));
Q_BUF U1320 ( .A(n1), .Z(\sa_events[7][62] ));
Q_BUF U1321 ( .A(n1), .Z(\sa_events[7][61] ));
Q_BUF U1322 ( .A(n1), .Z(\sa_events[7][60] ));
Q_BUF U1323 ( .A(n1), .Z(\sa_events[7][59] ));
Q_BUF U1324 ( .A(n1), .Z(\sa_events[7][58] ));
Q_BUF U1325 ( .A(n1), .Z(\sa_events[7][57] ));
Q_BUF U1326 ( .A(n1), .Z(\sa_events[7][56] ));
Q_BUF U1327 ( .A(n1), .Z(\sa_events[7][55] ));
Q_BUF U1328 ( .A(n1), .Z(\sa_events[7][54] ));
Q_BUF U1329 ( .A(n1), .Z(\sa_events[7][53] ));
Q_BUF U1330 ( .A(n1), .Z(\sa_events[7][52] ));
Q_BUF U1331 ( .A(n1), .Z(\sa_events[7][51] ));
Q_BUF U1332 ( .A(n1), .Z(\sa_events[7][50] ));
Q_BUF U1333 ( .A(n1), .Z(\sa_events[7][49] ));
Q_BUF U1334 ( .A(n1), .Z(\sa_events[7][48] ));
Q_BUF U1335 ( .A(n1), .Z(\sa_events[7][47] ));
Q_BUF U1336 ( .A(n1), .Z(\sa_events[7][46] ));
Q_BUF U1337 ( .A(n1), .Z(\sa_events[7][45] ));
Q_BUF U1338 ( .A(n1), .Z(\sa_events[7][44] ));
Q_BUF U1339 ( .A(n1), .Z(\sa_events[7][43] ));
Q_BUF U1340 ( .A(n1), .Z(\sa_events[7][42] ));
Q_BUF U1341 ( .A(n1), .Z(\sa_events[7][41] ));
Q_BUF U1342 ( .A(n1), .Z(\sa_events[7][40] ));
Q_BUF U1343 ( .A(n1), .Z(\sa_events[7][39] ));
Q_BUF U1344 ( .A(n1), .Z(\sa_events[7][38] ));
Q_BUF U1345 ( .A(n1), .Z(\sa_events[7][37] ));
Q_BUF U1346 ( .A(n1), .Z(\sa_events[7][36] ));
Q_BUF U1347 ( .A(n1), .Z(\sa_events[7][35] ));
Q_BUF U1348 ( .A(n1), .Z(\sa_events[7][34] ));
Q_BUF U1349 ( .A(n1), .Z(\sa_events[7][33] ));
Q_BUF U1350 ( .A(n1), .Z(\sa_events[7][32] ));
Q_BUF U1351 ( .A(n1), .Z(\sa_events[7][31] ));
Q_BUF U1352 ( .A(n1), .Z(\sa_events[7][30] ));
Q_BUF U1353 ( .A(n1), .Z(\sa_events[7][29] ));
Q_BUF U1354 ( .A(n1), .Z(\sa_events[7][28] ));
Q_BUF U1355 ( .A(n1), .Z(\sa_events[7][27] ));
Q_BUF U1356 ( .A(n1), .Z(\sa_events[7][26] ));
Q_BUF U1357 ( .A(n1), .Z(\sa_events[7][25] ));
Q_BUF U1358 ( .A(n1), .Z(\sa_events[7][24] ));
Q_BUF U1359 ( .A(n1), .Z(\sa_events[7][23] ));
Q_BUF U1360 ( .A(n1), .Z(\sa_events[7][22] ));
Q_BUF U1361 ( .A(n1), .Z(\sa_events[7][21] ));
Q_BUF U1362 ( .A(n1), .Z(\sa_events[7][20] ));
Q_BUF U1363 ( .A(n1), .Z(\sa_events[7][19] ));
Q_BUF U1364 ( .A(n1), .Z(\sa_events[7][18] ));
Q_BUF U1365 ( .A(n1), .Z(\sa_events[7][17] ));
Q_BUF U1366 ( .A(n1), .Z(\sa_events[7][16] ));
Q_BUF U1367 ( .A(n1), .Z(\sa_events[7][15] ));
Q_BUF U1368 ( .A(n1), .Z(\sa_events[7][14] ));
Q_BUF U1369 ( .A(n1), .Z(\sa_events[7][13] ));
Q_BUF U1370 ( .A(n1), .Z(\sa_events[7][12] ));
Q_BUF U1371 ( .A(n1), .Z(\sa_events[7][11] ));
Q_BUF U1372 ( .A(n1), .Z(\sa_events[7][10] ));
Q_BUF U1373 ( .A(n1), .Z(\sa_events[7][9] ));
Q_BUF U1374 ( .A(n1), .Z(\sa_events[7][8] ));
Q_BUF U1375 ( .A(n1), .Z(\sa_events[7][7] ));
Q_BUF U1376 ( .A(n1), .Z(\sa_events[7][6] ));
Q_BUF U1377 ( .A(n1), .Z(\sa_events[7][5] ));
Q_BUF U1378 ( .A(n1), .Z(\sa_events[7][4] ));
Q_BUF U1379 ( .A(n1), .Z(\sa_events[7][3] ));
Q_BUF U1380 ( .A(n1), .Z(\sa_events[7][2] ));
Q_BUF U1381 ( .A(n1), .Z(\sa_events[7][1] ));
Q_BUF U1382 ( .A(n1), .Z(\sa_events[7][0] ));
Q_BUF U1383 ( .A(n1), .Z(\sa_events[8][63] ));
Q_BUF U1384 ( .A(n1), .Z(\sa_events[8][62] ));
Q_BUF U1385 ( .A(n1), .Z(\sa_events[8][61] ));
Q_BUF U1386 ( .A(n1), .Z(\sa_events[8][60] ));
Q_BUF U1387 ( .A(n1), .Z(\sa_events[8][59] ));
Q_BUF U1388 ( .A(n1), .Z(\sa_events[8][58] ));
Q_BUF U1389 ( .A(n1), .Z(\sa_events[8][57] ));
Q_BUF U1390 ( .A(n1), .Z(\sa_events[8][56] ));
Q_BUF U1391 ( .A(n1), .Z(\sa_events[8][55] ));
Q_BUF U1392 ( .A(n1), .Z(\sa_events[8][54] ));
Q_BUF U1393 ( .A(n1), .Z(\sa_events[8][53] ));
Q_BUF U1394 ( .A(n1), .Z(\sa_events[8][52] ));
Q_BUF U1395 ( .A(n1), .Z(\sa_events[8][51] ));
Q_BUF U1396 ( .A(n1), .Z(\sa_events[8][50] ));
Q_BUF U1397 ( .A(n1), .Z(\sa_events[8][49] ));
Q_BUF U1398 ( .A(n1), .Z(\sa_events[8][48] ));
Q_BUF U1399 ( .A(n1), .Z(\sa_events[8][47] ));
Q_BUF U1400 ( .A(n1), .Z(\sa_events[8][46] ));
Q_BUF U1401 ( .A(n1), .Z(\sa_events[8][45] ));
Q_BUF U1402 ( .A(n1), .Z(\sa_events[8][44] ));
Q_BUF U1403 ( .A(n1), .Z(\sa_events[8][43] ));
Q_BUF U1404 ( .A(n1), .Z(\sa_events[8][42] ));
Q_BUF U1405 ( .A(n1), .Z(\sa_events[8][41] ));
Q_BUF U1406 ( .A(n1), .Z(\sa_events[8][40] ));
Q_BUF U1407 ( .A(n1), .Z(\sa_events[8][39] ));
Q_BUF U1408 ( .A(n1), .Z(\sa_events[8][38] ));
Q_BUF U1409 ( .A(n1), .Z(\sa_events[8][37] ));
Q_BUF U1410 ( .A(n1), .Z(\sa_events[8][36] ));
Q_BUF U1411 ( .A(n1), .Z(\sa_events[8][35] ));
Q_BUF U1412 ( .A(n1), .Z(\sa_events[8][34] ));
Q_BUF U1413 ( .A(n1), .Z(\sa_events[8][33] ));
Q_BUF U1414 ( .A(n1), .Z(\sa_events[8][32] ));
Q_BUF U1415 ( .A(n1), .Z(\sa_events[8][31] ));
Q_BUF U1416 ( .A(n1), .Z(\sa_events[8][30] ));
Q_BUF U1417 ( .A(n1), .Z(\sa_events[8][29] ));
Q_BUF U1418 ( .A(n1), .Z(\sa_events[8][28] ));
Q_BUF U1419 ( .A(n1), .Z(\sa_events[8][27] ));
Q_BUF U1420 ( .A(n1), .Z(\sa_events[8][26] ));
Q_BUF U1421 ( .A(n1), .Z(\sa_events[8][25] ));
Q_BUF U1422 ( .A(n1), .Z(\sa_events[8][24] ));
Q_BUF U1423 ( .A(n1), .Z(\sa_events[8][23] ));
Q_BUF U1424 ( .A(n1), .Z(\sa_events[8][22] ));
Q_BUF U1425 ( .A(n1), .Z(\sa_events[8][21] ));
Q_BUF U1426 ( .A(n1), .Z(\sa_events[8][20] ));
Q_BUF U1427 ( .A(n1), .Z(\sa_events[8][19] ));
Q_BUF U1428 ( .A(n1), .Z(\sa_events[8][18] ));
Q_BUF U1429 ( .A(n1), .Z(\sa_events[8][17] ));
Q_BUF U1430 ( .A(n1), .Z(\sa_events[8][16] ));
Q_BUF U1431 ( .A(n1), .Z(\sa_events[8][15] ));
Q_BUF U1432 ( .A(n1), .Z(\sa_events[8][14] ));
Q_BUF U1433 ( .A(n1), .Z(\sa_events[8][13] ));
Q_BUF U1434 ( .A(n1), .Z(\sa_events[8][12] ));
Q_BUF U1435 ( .A(n1), .Z(\sa_events[8][11] ));
Q_BUF U1436 ( .A(n1), .Z(\sa_events[8][10] ));
Q_BUF U1437 ( .A(n1), .Z(\sa_events[8][9] ));
Q_BUF U1438 ( .A(n1), .Z(\sa_events[8][8] ));
Q_BUF U1439 ( .A(n1), .Z(\sa_events[8][7] ));
Q_BUF U1440 ( .A(n1), .Z(\sa_events[8][6] ));
Q_BUF U1441 ( .A(n1), .Z(\sa_events[8][5] ));
Q_BUF U1442 ( .A(n1), .Z(\sa_events[8][4] ));
Q_BUF U1443 ( .A(n1), .Z(\sa_events[8][3] ));
Q_BUF U1444 ( .A(n1), .Z(\sa_events[8][2] ));
Q_BUF U1445 ( .A(n1), .Z(\sa_events[8][1] ));
Q_BUF U1446 ( .A(n1), .Z(\sa_events[8][0] ));
Q_BUF U1447 ( .A(n1), .Z(\sa_events[9][63] ));
Q_BUF U1448 ( .A(n1), .Z(\sa_events[9][62] ));
Q_BUF U1449 ( .A(n1), .Z(\sa_events[9][61] ));
Q_BUF U1450 ( .A(n1), .Z(\sa_events[9][60] ));
Q_BUF U1451 ( .A(n1), .Z(\sa_events[9][59] ));
Q_BUF U1452 ( .A(n1), .Z(\sa_events[9][58] ));
Q_BUF U1453 ( .A(n1), .Z(\sa_events[9][57] ));
Q_BUF U1454 ( .A(n1), .Z(\sa_events[9][56] ));
Q_BUF U1455 ( .A(n1), .Z(\sa_events[9][55] ));
Q_BUF U1456 ( .A(n1), .Z(\sa_events[9][54] ));
Q_BUF U1457 ( .A(n1), .Z(\sa_events[9][53] ));
Q_BUF U1458 ( .A(n1), .Z(\sa_events[9][52] ));
Q_BUF U1459 ( .A(n1), .Z(\sa_events[9][51] ));
Q_BUF U1460 ( .A(n1), .Z(\sa_events[9][50] ));
Q_BUF U1461 ( .A(n1), .Z(\sa_events[9][49] ));
Q_BUF U1462 ( .A(n1), .Z(\sa_events[9][48] ));
Q_BUF U1463 ( .A(n1), .Z(\sa_events[9][47] ));
Q_BUF U1464 ( .A(n1), .Z(\sa_events[9][46] ));
Q_BUF U1465 ( .A(n1), .Z(\sa_events[9][45] ));
Q_BUF U1466 ( .A(n1), .Z(\sa_events[9][44] ));
Q_BUF U1467 ( .A(n1), .Z(\sa_events[9][43] ));
Q_BUF U1468 ( .A(n1), .Z(\sa_events[9][42] ));
Q_BUF U1469 ( .A(n1), .Z(\sa_events[9][41] ));
Q_BUF U1470 ( .A(n1), .Z(\sa_events[9][40] ));
Q_BUF U1471 ( .A(n1), .Z(\sa_events[9][39] ));
Q_BUF U1472 ( .A(n1), .Z(\sa_events[9][38] ));
Q_BUF U1473 ( .A(n1), .Z(\sa_events[9][37] ));
Q_BUF U1474 ( .A(n1), .Z(\sa_events[9][36] ));
Q_BUF U1475 ( .A(n1), .Z(\sa_events[9][35] ));
Q_BUF U1476 ( .A(n1), .Z(\sa_events[9][34] ));
Q_BUF U1477 ( .A(n1), .Z(\sa_events[9][33] ));
Q_BUF U1478 ( .A(n1), .Z(\sa_events[9][32] ));
Q_BUF U1479 ( .A(n1), .Z(\sa_events[9][31] ));
Q_BUF U1480 ( .A(n1), .Z(\sa_events[9][30] ));
Q_BUF U1481 ( .A(n1), .Z(\sa_events[9][29] ));
Q_BUF U1482 ( .A(n1), .Z(\sa_events[9][28] ));
Q_BUF U1483 ( .A(n1), .Z(\sa_events[9][27] ));
Q_BUF U1484 ( .A(n1), .Z(\sa_events[9][26] ));
Q_BUF U1485 ( .A(n1), .Z(\sa_events[9][25] ));
Q_BUF U1486 ( .A(n1), .Z(\sa_events[9][24] ));
Q_BUF U1487 ( .A(n1), .Z(\sa_events[9][23] ));
Q_BUF U1488 ( .A(n1), .Z(\sa_events[9][22] ));
Q_BUF U1489 ( .A(n1), .Z(\sa_events[9][21] ));
Q_BUF U1490 ( .A(n1), .Z(\sa_events[9][20] ));
Q_BUF U1491 ( .A(n1), .Z(\sa_events[9][19] ));
Q_BUF U1492 ( .A(n1), .Z(\sa_events[9][18] ));
Q_BUF U1493 ( .A(n1), .Z(\sa_events[9][17] ));
Q_BUF U1494 ( .A(n1), .Z(\sa_events[9][16] ));
Q_BUF U1495 ( .A(n1), .Z(\sa_events[9][15] ));
Q_BUF U1496 ( .A(n1), .Z(\sa_events[9][14] ));
Q_BUF U1497 ( .A(n1), .Z(\sa_events[9][13] ));
Q_BUF U1498 ( .A(n1), .Z(\sa_events[9][12] ));
Q_BUF U1499 ( .A(n1), .Z(\sa_events[9][11] ));
Q_BUF U1500 ( .A(n1), .Z(\sa_events[9][10] ));
Q_BUF U1501 ( .A(n1), .Z(\sa_events[9][9] ));
Q_BUF U1502 ( .A(n1), .Z(\sa_events[9][8] ));
Q_BUF U1503 ( .A(n1), .Z(\sa_events[9][7] ));
Q_BUF U1504 ( .A(n1), .Z(\sa_events[9][6] ));
Q_BUF U1505 ( .A(n1), .Z(\sa_events[9][5] ));
Q_BUF U1506 ( .A(n1), .Z(\sa_events[9][4] ));
Q_BUF U1507 ( .A(n1), .Z(\sa_events[9][3] ));
Q_BUF U1508 ( .A(n1), .Z(\sa_events[9][2] ));
Q_BUF U1509 ( .A(n1), .Z(\sa_events[9][1] ));
Q_BUF U1510 ( .A(n1), .Z(\sa_events[9][0] ));
Q_BUF U1511 ( .A(n1), .Z(\sa_events[10][63] ));
Q_BUF U1512 ( .A(n1), .Z(\sa_events[10][62] ));
Q_BUF U1513 ( .A(n1), .Z(\sa_events[10][61] ));
Q_BUF U1514 ( .A(n1), .Z(\sa_events[10][60] ));
Q_BUF U1515 ( .A(n1), .Z(\sa_events[10][59] ));
Q_BUF U1516 ( .A(n1), .Z(\sa_events[10][58] ));
Q_BUF U1517 ( .A(n1), .Z(\sa_events[10][57] ));
Q_BUF U1518 ( .A(n1), .Z(\sa_events[10][56] ));
Q_BUF U1519 ( .A(n1), .Z(\sa_events[10][55] ));
Q_BUF U1520 ( .A(n1), .Z(\sa_events[10][54] ));
Q_BUF U1521 ( .A(n1), .Z(\sa_events[10][53] ));
Q_BUF U1522 ( .A(n1), .Z(\sa_events[10][52] ));
Q_BUF U1523 ( .A(n1), .Z(\sa_events[10][51] ));
Q_BUF U1524 ( .A(n1), .Z(\sa_events[10][50] ));
Q_BUF U1525 ( .A(n1), .Z(\sa_events[10][49] ));
Q_BUF U1526 ( .A(n1), .Z(\sa_events[10][48] ));
Q_BUF U1527 ( .A(n1), .Z(\sa_events[10][47] ));
Q_BUF U1528 ( .A(n1), .Z(\sa_events[10][46] ));
Q_BUF U1529 ( .A(n1), .Z(\sa_events[10][45] ));
Q_BUF U1530 ( .A(n1), .Z(\sa_events[10][44] ));
Q_BUF U1531 ( .A(n1), .Z(\sa_events[10][43] ));
Q_BUF U1532 ( .A(n1), .Z(\sa_events[10][42] ));
Q_BUF U1533 ( .A(n1), .Z(\sa_events[10][41] ));
Q_BUF U1534 ( .A(n1), .Z(\sa_events[10][40] ));
Q_BUF U1535 ( .A(n1), .Z(\sa_events[10][39] ));
Q_BUF U1536 ( .A(n1), .Z(\sa_events[10][38] ));
Q_BUF U1537 ( .A(n1), .Z(\sa_events[10][37] ));
Q_BUF U1538 ( .A(n1), .Z(\sa_events[10][36] ));
Q_BUF U1539 ( .A(n1), .Z(\sa_events[10][35] ));
Q_BUF U1540 ( .A(n1), .Z(\sa_events[10][34] ));
Q_BUF U1541 ( .A(n1), .Z(\sa_events[10][33] ));
Q_BUF U1542 ( .A(n1), .Z(\sa_events[10][32] ));
Q_BUF U1543 ( .A(n1), .Z(\sa_events[10][31] ));
Q_BUF U1544 ( .A(n1), .Z(\sa_events[10][30] ));
Q_BUF U1545 ( .A(n1), .Z(\sa_events[10][29] ));
Q_BUF U1546 ( .A(n1), .Z(\sa_events[10][28] ));
Q_BUF U1547 ( .A(n1), .Z(\sa_events[10][27] ));
Q_BUF U1548 ( .A(n1), .Z(\sa_events[10][26] ));
Q_BUF U1549 ( .A(n1), .Z(\sa_events[10][25] ));
Q_BUF U1550 ( .A(n1), .Z(\sa_events[10][24] ));
Q_BUF U1551 ( .A(n1), .Z(\sa_events[10][23] ));
Q_BUF U1552 ( .A(n1), .Z(\sa_events[10][22] ));
Q_BUF U1553 ( .A(n1), .Z(\sa_events[10][21] ));
Q_BUF U1554 ( .A(n1), .Z(\sa_events[10][20] ));
Q_BUF U1555 ( .A(n1), .Z(\sa_events[10][19] ));
Q_BUF U1556 ( .A(n1), .Z(\sa_events[10][18] ));
Q_BUF U1557 ( .A(n1), .Z(\sa_events[10][17] ));
Q_BUF U1558 ( .A(n1), .Z(\sa_events[10][16] ));
Q_BUF U1559 ( .A(n1), .Z(\sa_events[10][15] ));
Q_BUF U1560 ( .A(n1), .Z(\sa_events[10][14] ));
Q_BUF U1561 ( .A(n1), .Z(\sa_events[10][13] ));
Q_BUF U1562 ( .A(n1), .Z(\sa_events[10][12] ));
Q_BUF U1563 ( .A(n1), .Z(\sa_events[10][11] ));
Q_BUF U1564 ( .A(n1), .Z(\sa_events[10][10] ));
Q_BUF U1565 ( .A(n1), .Z(\sa_events[10][9] ));
Q_BUF U1566 ( .A(n1), .Z(\sa_events[10][8] ));
Q_BUF U1567 ( .A(n1), .Z(\sa_events[10][7] ));
Q_BUF U1568 ( .A(n1), .Z(\sa_events[10][6] ));
Q_BUF U1569 ( .A(n1), .Z(\sa_events[10][5] ));
Q_BUF U1570 ( .A(n1), .Z(\sa_events[10][4] ));
Q_BUF U1571 ( .A(n1), .Z(\sa_events[10][3] ));
Q_BUF U1572 ( .A(n1), .Z(\sa_events[10][2] ));
Q_BUF U1573 ( .A(n1), .Z(\sa_events[10][1] ));
Q_BUF U1574 ( .A(n1), .Z(\sa_events[10][0] ));
Q_BUF U1575 ( .A(n1), .Z(\sa_events[11][63] ));
Q_BUF U1576 ( .A(n1), .Z(\sa_events[11][62] ));
Q_BUF U1577 ( .A(n1), .Z(\sa_events[11][61] ));
Q_BUF U1578 ( .A(n1), .Z(\sa_events[11][60] ));
Q_BUF U1579 ( .A(n1), .Z(\sa_events[11][59] ));
Q_BUF U1580 ( .A(n1), .Z(\sa_events[11][58] ));
Q_BUF U1581 ( .A(n1), .Z(\sa_events[11][57] ));
Q_BUF U1582 ( .A(n1), .Z(\sa_events[11][56] ));
Q_BUF U1583 ( .A(n1), .Z(\sa_events[11][55] ));
Q_BUF U1584 ( .A(n1), .Z(\sa_events[11][54] ));
Q_BUF U1585 ( .A(n1), .Z(\sa_events[11][53] ));
Q_BUF U1586 ( .A(n1), .Z(\sa_events[11][52] ));
Q_BUF U1587 ( .A(n1), .Z(\sa_events[11][51] ));
Q_BUF U1588 ( .A(n1), .Z(\sa_events[11][50] ));
Q_BUF U1589 ( .A(n1), .Z(\sa_events[11][49] ));
Q_BUF U1590 ( .A(n1), .Z(\sa_events[11][48] ));
Q_BUF U1591 ( .A(n1), .Z(\sa_events[11][47] ));
Q_BUF U1592 ( .A(n1), .Z(\sa_events[11][46] ));
Q_BUF U1593 ( .A(n1), .Z(\sa_events[11][45] ));
Q_BUF U1594 ( .A(n1), .Z(\sa_events[11][44] ));
Q_BUF U1595 ( .A(n1), .Z(\sa_events[11][43] ));
Q_BUF U1596 ( .A(n1), .Z(\sa_events[11][42] ));
Q_BUF U1597 ( .A(n1), .Z(\sa_events[11][41] ));
Q_BUF U1598 ( .A(n1), .Z(\sa_events[11][40] ));
Q_BUF U1599 ( .A(n1), .Z(\sa_events[11][39] ));
Q_BUF U1600 ( .A(n1), .Z(\sa_events[11][38] ));
Q_BUF U1601 ( .A(n1), .Z(\sa_events[11][37] ));
Q_BUF U1602 ( .A(n1), .Z(\sa_events[11][36] ));
Q_BUF U1603 ( .A(n1), .Z(\sa_events[11][35] ));
Q_BUF U1604 ( .A(n1), .Z(\sa_events[11][34] ));
Q_BUF U1605 ( .A(n1), .Z(\sa_events[11][33] ));
Q_BUF U1606 ( .A(n1), .Z(\sa_events[11][32] ));
Q_BUF U1607 ( .A(n1), .Z(\sa_events[11][31] ));
Q_BUF U1608 ( .A(n1), .Z(\sa_events[11][30] ));
Q_BUF U1609 ( .A(n1), .Z(\sa_events[11][29] ));
Q_BUF U1610 ( .A(n1), .Z(\sa_events[11][28] ));
Q_BUF U1611 ( .A(n1), .Z(\sa_events[11][27] ));
Q_BUF U1612 ( .A(n1), .Z(\sa_events[11][26] ));
Q_BUF U1613 ( .A(n1), .Z(\sa_events[11][25] ));
Q_BUF U1614 ( .A(n1), .Z(\sa_events[11][24] ));
Q_BUF U1615 ( .A(n1), .Z(\sa_events[11][23] ));
Q_BUF U1616 ( .A(n1), .Z(\sa_events[11][22] ));
Q_BUF U1617 ( .A(n1), .Z(\sa_events[11][21] ));
Q_BUF U1618 ( .A(n1), .Z(\sa_events[11][20] ));
Q_BUF U1619 ( .A(n1), .Z(\sa_events[11][19] ));
Q_BUF U1620 ( .A(n1), .Z(\sa_events[11][18] ));
Q_BUF U1621 ( .A(n1), .Z(\sa_events[11][17] ));
Q_BUF U1622 ( .A(n1), .Z(\sa_events[11][16] ));
Q_BUF U1623 ( .A(n1), .Z(\sa_events[11][15] ));
Q_BUF U1624 ( .A(n1), .Z(\sa_events[11][14] ));
Q_BUF U1625 ( .A(n1), .Z(\sa_events[11][13] ));
Q_BUF U1626 ( .A(n1), .Z(\sa_events[11][12] ));
Q_BUF U1627 ( .A(n1), .Z(\sa_events[11][11] ));
Q_BUF U1628 ( .A(n1), .Z(\sa_events[11][10] ));
Q_BUF U1629 ( .A(n1), .Z(\sa_events[11][9] ));
Q_BUF U1630 ( .A(n1), .Z(\sa_events[11][8] ));
Q_BUF U1631 ( .A(n1), .Z(\sa_events[11][7] ));
Q_BUF U1632 ( .A(n1), .Z(\sa_events[11][6] ));
Q_BUF U1633 ( .A(n1), .Z(\sa_events[11][5] ));
Q_BUF U1634 ( .A(n1), .Z(\sa_events[11][4] ));
Q_BUF U1635 ( .A(n1), .Z(\sa_events[11][3] ));
Q_BUF U1636 ( .A(n1), .Z(\sa_events[11][2] ));
Q_BUF U1637 ( .A(n1), .Z(\sa_events[11][1] ));
Q_BUF U1638 ( .A(n1), .Z(\sa_events[11][0] ));
Q_BUF U1639 ( .A(n1), .Z(\sa_events[12][63] ));
Q_BUF U1640 ( .A(n1), .Z(\sa_events[12][62] ));
Q_BUF U1641 ( .A(n1), .Z(\sa_events[12][61] ));
Q_BUF U1642 ( .A(n1), .Z(\sa_events[12][60] ));
Q_BUF U1643 ( .A(n1), .Z(\sa_events[12][59] ));
Q_BUF U1644 ( .A(n1), .Z(\sa_events[12][58] ));
Q_BUF U1645 ( .A(n1), .Z(\sa_events[12][57] ));
Q_BUF U1646 ( .A(n1), .Z(\sa_events[12][56] ));
Q_BUF U1647 ( .A(n1), .Z(\sa_events[12][55] ));
Q_BUF U1648 ( .A(n1), .Z(\sa_events[12][54] ));
Q_BUF U1649 ( .A(n1), .Z(\sa_events[12][53] ));
Q_BUF U1650 ( .A(n1), .Z(\sa_events[12][52] ));
Q_BUF U1651 ( .A(n1), .Z(\sa_events[12][51] ));
Q_BUF U1652 ( .A(n1), .Z(\sa_events[12][50] ));
Q_BUF U1653 ( .A(n1), .Z(\sa_events[12][49] ));
Q_BUF U1654 ( .A(n1), .Z(\sa_events[12][48] ));
Q_BUF U1655 ( .A(n1), .Z(\sa_events[12][47] ));
Q_BUF U1656 ( .A(n1), .Z(\sa_events[12][46] ));
Q_BUF U1657 ( .A(n1), .Z(\sa_events[12][45] ));
Q_BUF U1658 ( .A(n1), .Z(\sa_events[12][44] ));
Q_BUF U1659 ( .A(n1), .Z(\sa_events[12][43] ));
Q_BUF U1660 ( .A(n1), .Z(\sa_events[12][42] ));
Q_BUF U1661 ( .A(n1), .Z(\sa_events[12][41] ));
Q_BUF U1662 ( .A(n1), .Z(\sa_events[12][40] ));
Q_BUF U1663 ( .A(n1), .Z(\sa_events[12][39] ));
Q_BUF U1664 ( .A(n1), .Z(\sa_events[12][38] ));
Q_BUF U1665 ( .A(n1), .Z(\sa_events[12][37] ));
Q_BUF U1666 ( .A(n1), .Z(\sa_events[12][36] ));
Q_BUF U1667 ( .A(n1), .Z(\sa_events[12][35] ));
Q_BUF U1668 ( .A(n1), .Z(\sa_events[12][34] ));
Q_BUF U1669 ( .A(n1), .Z(\sa_events[12][33] ));
Q_BUF U1670 ( .A(n1), .Z(\sa_events[12][32] ));
Q_BUF U1671 ( .A(n1), .Z(\sa_events[12][31] ));
Q_BUF U1672 ( .A(n1), .Z(\sa_events[12][30] ));
Q_BUF U1673 ( .A(n1), .Z(\sa_events[12][29] ));
Q_BUF U1674 ( .A(n1), .Z(\sa_events[12][28] ));
Q_BUF U1675 ( .A(n1), .Z(\sa_events[12][27] ));
Q_BUF U1676 ( .A(n1), .Z(\sa_events[12][26] ));
Q_BUF U1677 ( .A(n1), .Z(\sa_events[12][25] ));
Q_BUF U1678 ( .A(n1), .Z(\sa_events[12][24] ));
Q_BUF U1679 ( .A(n1), .Z(\sa_events[12][23] ));
Q_BUF U1680 ( .A(n1), .Z(\sa_events[12][22] ));
Q_BUF U1681 ( .A(n1), .Z(\sa_events[12][21] ));
Q_BUF U1682 ( .A(n1), .Z(\sa_events[12][20] ));
Q_BUF U1683 ( .A(n1), .Z(\sa_events[12][19] ));
Q_BUF U1684 ( .A(n1), .Z(\sa_events[12][18] ));
Q_BUF U1685 ( .A(n1), .Z(\sa_events[12][17] ));
Q_BUF U1686 ( .A(n1), .Z(\sa_events[12][16] ));
Q_BUF U1687 ( .A(n1), .Z(\sa_events[12][15] ));
Q_BUF U1688 ( .A(n1), .Z(\sa_events[12][14] ));
Q_BUF U1689 ( .A(n1), .Z(\sa_events[12][13] ));
Q_BUF U1690 ( .A(n1), .Z(\sa_events[12][12] ));
Q_BUF U1691 ( .A(n1), .Z(\sa_events[12][11] ));
Q_BUF U1692 ( .A(n1), .Z(\sa_events[12][10] ));
Q_BUF U1693 ( .A(n1), .Z(\sa_events[12][9] ));
Q_BUF U1694 ( .A(n1), .Z(\sa_events[12][8] ));
Q_BUF U1695 ( .A(n1), .Z(\sa_events[12][7] ));
Q_BUF U1696 ( .A(n1), .Z(\sa_events[12][6] ));
Q_BUF U1697 ( .A(n1), .Z(\sa_events[12][5] ));
Q_BUF U1698 ( .A(n1), .Z(\sa_events[12][4] ));
Q_BUF U1699 ( .A(n1), .Z(\sa_events[12][3] ));
Q_BUF U1700 ( .A(n1), .Z(\sa_events[12][2] ));
Q_BUF U1701 ( .A(n1), .Z(\sa_events[12][1] ));
Q_BUF U1702 ( .A(n1), .Z(\sa_events[12][0] ));
Q_BUF U1703 ( .A(n1), .Z(\sa_events[13][63] ));
Q_BUF U1704 ( .A(n1), .Z(\sa_events[13][62] ));
Q_BUF U1705 ( .A(n1), .Z(\sa_events[13][61] ));
Q_BUF U1706 ( .A(n1), .Z(\sa_events[13][60] ));
Q_BUF U1707 ( .A(n1), .Z(\sa_events[13][59] ));
Q_BUF U1708 ( .A(n1), .Z(\sa_events[13][58] ));
Q_BUF U1709 ( .A(n1), .Z(\sa_events[13][57] ));
Q_BUF U1710 ( .A(n1), .Z(\sa_events[13][56] ));
Q_BUF U1711 ( .A(n1), .Z(\sa_events[13][55] ));
Q_BUF U1712 ( .A(n1), .Z(\sa_events[13][54] ));
Q_BUF U1713 ( .A(n1), .Z(\sa_events[13][53] ));
Q_BUF U1714 ( .A(n1), .Z(\sa_events[13][52] ));
Q_BUF U1715 ( .A(n1), .Z(\sa_events[13][51] ));
Q_BUF U1716 ( .A(n1), .Z(\sa_events[13][50] ));
Q_BUF U1717 ( .A(n1), .Z(\sa_events[13][49] ));
Q_BUF U1718 ( .A(n1), .Z(\sa_events[13][48] ));
Q_BUF U1719 ( .A(n1), .Z(\sa_events[13][47] ));
Q_BUF U1720 ( .A(n1), .Z(\sa_events[13][46] ));
Q_BUF U1721 ( .A(n1), .Z(\sa_events[13][45] ));
Q_BUF U1722 ( .A(n1), .Z(\sa_events[13][44] ));
Q_BUF U1723 ( .A(n1), .Z(\sa_events[13][43] ));
Q_BUF U1724 ( .A(n1), .Z(\sa_events[13][42] ));
Q_BUF U1725 ( .A(n1), .Z(\sa_events[13][41] ));
Q_BUF U1726 ( .A(n1), .Z(\sa_events[13][40] ));
Q_BUF U1727 ( .A(n1), .Z(\sa_events[13][39] ));
Q_BUF U1728 ( .A(n1), .Z(\sa_events[13][38] ));
Q_BUF U1729 ( .A(n1), .Z(\sa_events[13][37] ));
Q_BUF U1730 ( .A(n1), .Z(\sa_events[13][36] ));
Q_BUF U1731 ( .A(n1), .Z(\sa_events[13][35] ));
Q_BUF U1732 ( .A(n1), .Z(\sa_events[13][34] ));
Q_BUF U1733 ( .A(n1), .Z(\sa_events[13][33] ));
Q_BUF U1734 ( .A(n1), .Z(\sa_events[13][32] ));
Q_BUF U1735 ( .A(n1), .Z(\sa_events[13][31] ));
Q_BUF U1736 ( .A(n1), .Z(\sa_events[13][30] ));
Q_BUF U1737 ( .A(n1), .Z(\sa_events[13][29] ));
Q_BUF U1738 ( .A(n1), .Z(\sa_events[13][28] ));
Q_BUF U1739 ( .A(n1), .Z(\sa_events[13][27] ));
Q_BUF U1740 ( .A(n1), .Z(\sa_events[13][26] ));
Q_BUF U1741 ( .A(n1), .Z(\sa_events[13][25] ));
Q_BUF U1742 ( .A(n1), .Z(\sa_events[13][24] ));
Q_BUF U1743 ( .A(n1), .Z(\sa_events[13][23] ));
Q_BUF U1744 ( .A(n1), .Z(\sa_events[13][22] ));
Q_BUF U1745 ( .A(n1), .Z(\sa_events[13][21] ));
Q_BUF U1746 ( .A(n1), .Z(\sa_events[13][20] ));
Q_BUF U1747 ( .A(n1), .Z(\sa_events[13][19] ));
Q_BUF U1748 ( .A(n1), .Z(\sa_events[13][18] ));
Q_BUF U1749 ( .A(n1), .Z(\sa_events[13][17] ));
Q_BUF U1750 ( .A(n1), .Z(\sa_events[13][16] ));
Q_BUF U1751 ( .A(n1), .Z(\sa_events[13][15] ));
Q_BUF U1752 ( .A(n1), .Z(\sa_events[13][14] ));
Q_BUF U1753 ( .A(n1), .Z(\sa_events[13][13] ));
Q_BUF U1754 ( .A(n1), .Z(\sa_events[13][12] ));
Q_BUF U1755 ( .A(n1), .Z(\sa_events[13][11] ));
Q_BUF U1756 ( .A(n1), .Z(\sa_events[13][10] ));
Q_BUF U1757 ( .A(n1), .Z(\sa_events[13][9] ));
Q_BUF U1758 ( .A(n1), .Z(\sa_events[13][8] ));
Q_BUF U1759 ( .A(n1), .Z(\sa_events[13][7] ));
Q_BUF U1760 ( .A(n1), .Z(\sa_events[13][6] ));
Q_BUF U1761 ( .A(n1), .Z(\sa_events[13][5] ));
Q_BUF U1762 ( .A(n1), .Z(\sa_events[13][4] ));
Q_BUF U1763 ( .A(n1), .Z(\sa_events[13][3] ));
Q_BUF U1764 ( .A(n1), .Z(\sa_events[13][2] ));
Q_BUF U1765 ( .A(n1), .Z(\sa_events[13][1] ));
Q_BUF U1766 ( .A(n1), .Z(\sa_events[13][0] ));
Q_BUF U1767 ( .A(n1), .Z(\sa_events[14][63] ));
Q_BUF U1768 ( .A(n1), .Z(\sa_events[14][62] ));
Q_BUF U1769 ( .A(n1), .Z(\sa_events[14][61] ));
Q_BUF U1770 ( .A(n1), .Z(\sa_events[14][60] ));
Q_BUF U1771 ( .A(n1), .Z(\sa_events[14][59] ));
Q_BUF U1772 ( .A(n1), .Z(\sa_events[14][58] ));
Q_BUF U1773 ( .A(n1), .Z(\sa_events[14][57] ));
Q_BUF U1774 ( .A(n1), .Z(\sa_events[14][56] ));
Q_BUF U1775 ( .A(n1), .Z(\sa_events[14][55] ));
Q_BUF U1776 ( .A(n1), .Z(\sa_events[14][54] ));
Q_BUF U1777 ( .A(n1), .Z(\sa_events[14][53] ));
Q_BUF U1778 ( .A(n1), .Z(\sa_events[14][52] ));
Q_BUF U1779 ( .A(n1), .Z(\sa_events[14][51] ));
Q_BUF U1780 ( .A(n1), .Z(\sa_events[14][50] ));
Q_BUF U1781 ( .A(n1), .Z(\sa_events[14][49] ));
Q_BUF U1782 ( .A(n1), .Z(\sa_events[14][48] ));
Q_BUF U1783 ( .A(n1), .Z(\sa_events[14][47] ));
Q_BUF U1784 ( .A(n1), .Z(\sa_events[14][46] ));
Q_BUF U1785 ( .A(n1), .Z(\sa_events[14][45] ));
Q_BUF U1786 ( .A(n1), .Z(\sa_events[14][44] ));
Q_BUF U1787 ( .A(n1), .Z(\sa_events[14][43] ));
Q_BUF U1788 ( .A(n1), .Z(\sa_events[14][42] ));
Q_BUF U1789 ( .A(n1), .Z(\sa_events[14][41] ));
Q_BUF U1790 ( .A(n1), .Z(\sa_events[14][40] ));
Q_BUF U1791 ( .A(n1), .Z(\sa_events[14][39] ));
Q_BUF U1792 ( .A(n1), .Z(\sa_events[14][38] ));
Q_BUF U1793 ( .A(n1), .Z(\sa_events[14][37] ));
Q_BUF U1794 ( .A(n1), .Z(\sa_events[14][36] ));
Q_BUF U1795 ( .A(n1), .Z(\sa_events[14][35] ));
Q_BUF U1796 ( .A(n1), .Z(\sa_events[14][34] ));
Q_BUF U1797 ( .A(n1), .Z(\sa_events[14][33] ));
Q_BUF U1798 ( .A(n1), .Z(\sa_events[14][32] ));
Q_BUF U1799 ( .A(n1), .Z(\sa_events[14][31] ));
Q_BUF U1800 ( .A(n1), .Z(\sa_events[14][30] ));
Q_BUF U1801 ( .A(n1), .Z(\sa_events[14][29] ));
Q_BUF U1802 ( .A(n1), .Z(\sa_events[14][28] ));
Q_BUF U1803 ( .A(n1), .Z(\sa_events[14][27] ));
Q_BUF U1804 ( .A(n1), .Z(\sa_events[14][26] ));
Q_BUF U1805 ( .A(n1), .Z(\sa_events[14][25] ));
Q_BUF U1806 ( .A(n1), .Z(\sa_events[14][24] ));
Q_BUF U1807 ( .A(n1), .Z(\sa_events[14][23] ));
Q_BUF U1808 ( .A(n1), .Z(\sa_events[14][22] ));
Q_BUF U1809 ( .A(n1), .Z(\sa_events[14][21] ));
Q_BUF U1810 ( .A(n1), .Z(\sa_events[14][20] ));
Q_BUF U1811 ( .A(n1), .Z(\sa_events[14][19] ));
Q_BUF U1812 ( .A(n1), .Z(\sa_events[14][18] ));
Q_BUF U1813 ( .A(n1), .Z(\sa_events[14][17] ));
Q_BUF U1814 ( .A(n1), .Z(\sa_events[14][16] ));
Q_BUF U1815 ( .A(n1), .Z(\sa_events[14][15] ));
Q_BUF U1816 ( .A(n1), .Z(\sa_events[14][14] ));
Q_BUF U1817 ( .A(n1), .Z(\sa_events[14][13] ));
Q_BUF U1818 ( .A(n1), .Z(\sa_events[14][12] ));
Q_BUF U1819 ( .A(n1), .Z(\sa_events[14][11] ));
Q_BUF U1820 ( .A(n1), .Z(\sa_events[14][10] ));
Q_BUF U1821 ( .A(n1), .Z(\sa_events[14][9] ));
Q_BUF U1822 ( .A(n1), .Z(\sa_events[14][8] ));
Q_BUF U1823 ( .A(n1), .Z(\sa_events[14][7] ));
Q_BUF U1824 ( .A(n1), .Z(\sa_events[14][6] ));
Q_BUF U1825 ( .A(n1), .Z(\sa_events[14][5] ));
Q_BUF U1826 ( .A(n1), .Z(\sa_events[14][4] ));
Q_BUF U1827 ( .A(n1), .Z(\sa_events[14][3] ));
Q_BUF U1828 ( .A(n1), .Z(\sa_events[14][2] ));
Q_BUF U1829 ( .A(n1), .Z(\sa_events[14][1] ));
Q_BUF U1830 ( .A(n1), .Z(\sa_events[14][0] ));
Q_BUF U1831 ( .A(n1), .Z(\sa_events[15][63] ));
Q_BUF U1832 ( .A(n1), .Z(\sa_events[15][62] ));
Q_BUF U1833 ( .A(n1), .Z(\sa_events[15][61] ));
Q_BUF U1834 ( .A(n1), .Z(\sa_events[15][60] ));
Q_BUF U1835 ( .A(n1), .Z(\sa_events[15][59] ));
Q_BUF U1836 ( .A(n1), .Z(\sa_events[15][58] ));
Q_BUF U1837 ( .A(n1), .Z(\sa_events[15][57] ));
Q_BUF U1838 ( .A(n1), .Z(\sa_events[15][56] ));
Q_BUF U1839 ( .A(n1), .Z(\sa_events[15][55] ));
Q_BUF U1840 ( .A(n1), .Z(\sa_events[15][54] ));
Q_BUF U1841 ( .A(n1), .Z(\sa_events[15][53] ));
Q_BUF U1842 ( .A(n1), .Z(\sa_events[15][52] ));
Q_BUF U1843 ( .A(n1), .Z(\sa_events[15][51] ));
Q_BUF U1844 ( .A(n1), .Z(\sa_events[15][50] ));
Q_BUF U1845 ( .A(n1), .Z(\sa_events[15][49] ));
Q_BUF U1846 ( .A(n1), .Z(\sa_events[15][48] ));
Q_BUF U1847 ( .A(n1), .Z(\sa_events[15][47] ));
Q_BUF U1848 ( .A(n1), .Z(\sa_events[15][46] ));
Q_BUF U1849 ( .A(n1), .Z(\sa_events[15][45] ));
Q_BUF U1850 ( .A(n1), .Z(\sa_events[15][44] ));
Q_BUF U1851 ( .A(n1), .Z(\sa_events[15][43] ));
Q_BUF U1852 ( .A(n1), .Z(\sa_events[15][42] ));
Q_BUF U1853 ( .A(n1), .Z(\sa_events[15][41] ));
Q_BUF U1854 ( .A(n1), .Z(\sa_events[15][40] ));
Q_BUF U1855 ( .A(n1), .Z(\sa_events[15][39] ));
Q_BUF U1856 ( .A(n1), .Z(\sa_events[15][38] ));
Q_BUF U1857 ( .A(n1), .Z(\sa_events[15][37] ));
Q_BUF U1858 ( .A(n1), .Z(\sa_events[15][36] ));
Q_BUF U1859 ( .A(n1), .Z(\sa_events[15][35] ));
Q_BUF U1860 ( .A(n1), .Z(\sa_events[15][34] ));
Q_BUF U1861 ( .A(n1), .Z(\sa_events[15][33] ));
Q_BUF U1862 ( .A(n1), .Z(\sa_events[15][32] ));
Q_BUF U1863 ( .A(n1), .Z(\sa_events[15][31] ));
Q_BUF U1864 ( .A(n1), .Z(\sa_events[15][30] ));
Q_BUF U1865 ( .A(n1), .Z(\sa_events[15][29] ));
Q_BUF U1866 ( .A(n1), .Z(\sa_events[15][28] ));
Q_BUF U1867 ( .A(n1), .Z(\sa_events[15][27] ));
Q_BUF U1868 ( .A(n1), .Z(\sa_events[15][26] ));
Q_BUF U1869 ( .A(n1), .Z(\sa_events[15][25] ));
Q_BUF U1870 ( .A(n1), .Z(\sa_events[15][24] ));
Q_BUF U1871 ( .A(n1), .Z(\sa_events[15][23] ));
Q_BUF U1872 ( .A(n1), .Z(\sa_events[15][22] ));
Q_BUF U1873 ( .A(n1), .Z(\sa_events[15][21] ));
Q_BUF U1874 ( .A(n1), .Z(\sa_events[15][20] ));
Q_BUF U1875 ( .A(n1), .Z(\sa_events[15][19] ));
Q_BUF U1876 ( .A(n1), .Z(\sa_events[15][18] ));
Q_BUF U1877 ( .A(n1), .Z(\sa_events[15][17] ));
Q_BUF U1878 ( .A(n1), .Z(\sa_events[15][16] ));
Q_BUF U1879 ( .A(n1), .Z(\sa_events[15][15] ));
Q_BUF U1880 ( .A(n1), .Z(\sa_events[15][14] ));
Q_BUF U1881 ( .A(n1), .Z(\sa_events[15][13] ));
Q_BUF U1882 ( .A(n1), .Z(\sa_events[15][12] ));
Q_BUF U1883 ( .A(n1), .Z(\sa_events[15][11] ));
Q_BUF U1884 ( .A(n1), .Z(\sa_events[15][10] ));
Q_BUF U1885 ( .A(n1), .Z(\sa_events[15][9] ));
Q_BUF U1886 ( .A(n1), .Z(\sa_events[15][8] ));
Q_BUF U1887 ( .A(n1), .Z(\sa_events[15][7] ));
Q_BUF U1888 ( .A(n1), .Z(\sa_events[15][6] ));
Q_BUF U1889 ( .A(n1), .Z(\sa_events[15][5] ));
Q_BUF U1890 ( .A(n1), .Z(\sa_events[15][4] ));
Q_BUF U1891 ( .A(n1), .Z(\sa_events[15][3] ));
Q_BUF U1892 ( .A(n1), .Z(\sa_events[15][2] ));
Q_BUF U1893 ( .A(n1), .Z(\sa_events[15][1] ));
Q_BUF U1894 ( .A(n1), .Z(\sa_events[15][0] ));
Q_ASSIGN U1895 ( .B(stat_aux_cmd_with_vf_pf_fail), .A(\sa_events[0][24] ));
Q_ASSIGN U1896 ( .B(stat_cddip3_stall_on_valid_key), .A(\sa_events[0][23] ));
Q_ASSIGN U1897 ( .B(stat_cddip2_stall_on_valid_key), .A(\sa_events[0][22] ));
Q_ASSIGN U1898 ( .B(stat_cddip1_stall_on_valid_key), .A(\sa_events[0][21] ));
Q_ASSIGN U1899 ( .B(stat_cddip0_stall_on_valid_key), .A(\sa_events[0][20] ));
Q_ASSIGN U1900 ( .B(stat_cceip3_stall_on_valid_key), .A(\sa_events[0][19] ));
Q_ASSIGN U1901 ( .B(stat_cceip2_stall_on_valid_key), .A(\sa_events[0][18] ));
Q_ASSIGN U1902 ( .B(stat_cceip1_stall_on_valid_key), .A(\sa_events[0][17] ));
Q_ASSIGN U1903 ( .B(stat_cceip0_stall_on_valid_key), .A(\sa_events[0][16] ));
Q_ASSIGN U1904 ( .B(stat_aux_key_type_13), .A(\sa_events[0][15] ));
Q_ASSIGN U1905 ( .B(stat_aux_key_type_12), .A(\sa_events[0][14] ));
Q_ASSIGN U1906 ( .B(stat_aux_key_type_11), .A(\sa_events[0][13] ));
Q_ASSIGN U1907 ( .B(stat_aux_key_type_10), .A(\sa_events[0][12] ));
Q_ASSIGN U1908 ( .B(stat_aux_key_type_9), .A(\sa_events[0][11] ));
Q_ASSIGN U1909 ( .B(stat_aux_key_type_8), .A(\sa_events[0][10] ));
Q_ASSIGN U1910 ( .B(stat_aux_key_type_7), .A(\sa_events[0][9] ));
Q_ASSIGN U1911 ( .B(stat_aux_key_type_6), .A(\sa_events[0][8] ));
Q_ASSIGN U1912 ( .B(stat_aux_key_type_5), .A(\sa_events[0][7] ));
Q_ASSIGN U1913 ( .B(stat_aux_key_type_4), .A(\sa_events[0][6] ));
Q_ASSIGN U1914 ( .B(stat_aux_key_type_3), .A(\sa_events[0][5] ));
Q_ASSIGN U1915 ( .B(stat_aux_key_type_2), .A(\sa_events[0][4] ));
Q_ASSIGN U1916 ( .B(stat_aux_key_type_1), .A(\sa_events[0][3] ));
Q_ASSIGN U1917 ( .B(stat_aux_key_type_0), .A(\sa_events[0][2] ));
Q_ASSIGN U1918 ( .B(stat_req_with_expired_seed), .A(\sa_events[0][1] ));
Q_ASSIGN U1919 ( .B(stat_drbg_reseed), .A(\sa_events[0][0] ));
ixc_assign _zz_strnp_169 ( idle_components[4], cceip_key_tlv_rsm_idle[3]);
ixc_assign _zz_strnp_168 ( idle_components[5], cceip_key_tlv_rsm_idle[2]);
ixc_assign _zz_strnp_167 ( idle_components[6], cceip_key_tlv_rsm_idle[1]);
ixc_assign _zz_strnp_166 ( idle_components[7], cceip_key_tlv_rsm_idle[0]);
ixc_assign _zz_strnp_165 ( idle_components[8], cddip_key_tlv_rsm_idle[3]);
ixc_assign _zz_strnp_164 ( idle_components[9], cddip_key_tlv_rsm_idle[2]);
ixc_assign _zz_strnp_163 ( idle_components[10], cddip_key_tlv_rsm_idle[1]);
ixc_assign _zz_strnp_162 ( idle_components[11], cddip_key_tlv_rsm_idle[0]);
ixc_assign_32 _zz_strnp_177 ( _zy_simnet_idle_components_4_w$[0:31], 
	idle_components[31:0]);
ixc_assign _zz_strnp_176 ( _zy_simnet_kme_idle_3_w$, kme_idle);
ixc_assign _zz_strnp_175 ( _zy_simnet_kme_ib_out_2_w$, kme_ib_out[0]);
ixc_assign _zz_strnp_174 ( _zy_simnet_set_txc_bp_int_1_w$, set_txc_bp_int);
ixc_assign _zz_strnp_173 ( _zy_simnet_disable_debug_cmd_q_0_w$, 
	disable_debug_cmd_q);
ixc_assign _zz_strnp_172 ( idle_components[0], kme_slv_empty);
ixc_assign _zz_strnp_171 ( idle_components[1], drng_idle);
ixc_assign _zz_strnp_170 ( idle_components[2], tlv_parser_idle);
Q_NR02 U1936 ( .A0(n15), .A1(n16), .Z(idle_components[3]));
Q_OR03 U1937 ( .A0(n12), .A1(n13), .A2(n14), .Z(n16));
Q_OR03 U1938 ( .A0(n9), .A1(n10), .A2(n11), .Z(n15));
Q_OR03 U1939 ( .A0(n6), .A1(n7), .A2(n8), .Z(n14));
Q_OR03 U1940 ( .A0(n3), .A1(n4), .A2(n5), .Z(n13));
Q_OR03 U1941 ( .A0(num_key_tlv_in_flight[1]), .A1(num_key_tlv_in_flight[0]), .A2(n2), .Z(n12));
Q_OR03 U1942 ( .A0(num_key_tlv_in_flight[4]), .A1(num_key_tlv_in_flight[3]), .A2(num_key_tlv_in_flight[2]), .Z(n11));
Q_OR03 U1943 ( .A0(num_key_tlv_in_flight[7]), .A1(num_key_tlv_in_flight[6]), .A2(num_key_tlv_in_flight[5]), .Z(n10));
Q_OR03 U1944 ( .A0(num_key_tlv_in_flight[10]), .A1(num_key_tlv_in_flight[9]), .A2(num_key_tlv_in_flight[8]), .Z(n9));
Q_OR03 U1945 ( .A0(num_key_tlv_in_flight[13]), .A1(num_key_tlv_in_flight[12]), .A2(num_key_tlv_in_flight[11]), .Z(n8));
Q_OR03 U1946 ( .A0(num_key_tlv_in_flight[16]), .A1(num_key_tlv_in_flight[15]), .A2(num_key_tlv_in_flight[14]), .Z(n7));
Q_OR03 U1947 ( .A0(num_key_tlv_in_flight[19]), .A1(num_key_tlv_in_flight[18]), .A2(num_key_tlv_in_flight[17]), .Z(n6));
Q_OR03 U1948 ( .A0(num_key_tlv_in_flight[22]), .A1(num_key_tlv_in_flight[21]), .A2(num_key_tlv_in_flight[20]), .Z(n5));
Q_OR03 U1949 ( .A0(num_key_tlv_in_flight[25]), .A1(num_key_tlv_in_flight[24]), .A2(num_key_tlv_in_flight[23]), .Z(n4));
Q_OR03 U1950 ( .A0(num_key_tlv_in_flight[28]), .A1(num_key_tlv_in_flight[27]), .A2(num_key_tlv_in_flight[26]), .Z(n3));
Q_OR03 U1951 ( .A0(num_key_tlv_in_flight[31]), .A1(num_key_tlv_in_flight[30]), .A2(num_key_tlv_in_flight[29]), .Z(n2));
ixc_assign_20 _zz_strnp_161 ( idle_components[31:12], 
	num_key_tlv_in_flight[19:0]);
ixc_assign_8 _zz_strnp_160 ( set_rsm_is_backpressuring[7:0], { 
	cddip_ob_full[3], cddip_ob_full[2], cddip_ob_full[1], 
	cddip_ob_full[0], cceip_ob_full[3], cceip_ob_full[2], 
	cceip_ob_full[1], cceip_ob_full[0]});
Q_OR03 U1954 ( .A0(cceip_encrypt_gcm_tag_fail_int), .A1(cceip_validate_gcm_tag_fail_int), .A2(cddip_decrypt_gcm_tag_fail_int), .Z(set_gcm_tag_fail_int));
Q_AN02 U1955 ( .A0(n17), .A1(core_kme_ib_out[0]), .Z(kme_ib_out[0]));
Q_INV U1956 ( .A(tready_override[8]), .Z(n17));
Q_FDP1 disable_debug_cmd_q_REG  ( .CK(clk), .R(rst_n), .D(disable_debug_cmd), .Q(disable_debug_cmd_q), .QN( ));
Q_FDP1 set_txc_bp_int_REG  ( .CK(clk), .R(rst_n), .D(n18), .Q(set_txc_bp_int), .QN( ));
Q_INV U1959 ( .A(kme_ib_out[0]), .Z(n18));
Q_FDP1 sa_clear_REG  ( .CK(clk), .R(rst_n), .D(n19), .Q(sa_clear), .QN( ));
Q_AN02 U1961 ( .A0(sa_global_ctrl[0]), .A1(n20), .Z(n19));
Q_FDP1 sa_snap_REG  ( .CK(clk), .R(rst_n), .D(n21), .Q(sa_snap), .QN( ));
Q_AN02 U1963 ( .A0(sa_global_ctrl[1]), .A1(n22), .Z(n21));
Q_FDP1 regs_sa_clear_live_r_REG  ( .CK(clk), .R(rst_n), .D(sa_global_ctrl[0]), .Q(regs_sa_clear_live_r), .QN(n20));
Q_FDP1 regs_sa_snap_r_REG  ( .CK(clk), .R(rst_n), .D(sa_global_ctrl[1]), .Q(regs_sa_snap_r), .QN(n22));
Q_OR03 U1966 ( .A0(cceip_key_tlv_rsm_end_pulse[3]), .A1(cceip_key_tlv_rsm_end_pulse[2]), .A2(cceip_key_tlv_rsm_end_pulse[1]), .Z(n23));
Q_OR03 U1967 ( .A0(cceip_key_tlv_rsm_end_pulse[0]), .A1(n23), .A2(n25), .Z(n73));
Q_OR03 U1968 ( .A0(cddip_key_tlv_rsm_end_pulse[3]), .A1(cddip_key_tlv_rsm_end_pulse[2]), .A2(cddip_key_tlv_rsm_end_pulse[1]), .Z(n24));
Q_OR02 U1969 ( .A0(cddip_key_tlv_rsm_end_pulse[0]), .A1(n24), .Z(n25));
Q_XOR3 U1970 ( .A0(num_key_tlv_in_flight[31]), .A1(n73), .A2(n70), .Z(n71));
Q_AD02 U1971 ( .CI(num_key_tlv_in_flight[0]), .A0(num_key_tlv_in_flight[1]), .A1(num_key_tlv_in_flight[2]), .B0(n73), .B1(n73), .S0(n26), .S1(n27), .CO(n28));
Q_AD02 U1972 ( .CI(n28), .A0(num_key_tlv_in_flight[3]), .A1(num_key_tlv_in_flight[4]), .B0(n73), .B1(n73), .S0(n29), .S1(n30), .CO(n31));
Q_AD02 U1973 ( .CI(n31), .A0(num_key_tlv_in_flight[5]), .A1(num_key_tlv_in_flight[6]), .B0(n73), .B1(n73), .S0(n32), .S1(n33), .CO(n34));
Q_AD02 U1974 ( .CI(n34), .A0(num_key_tlv_in_flight[7]), .A1(num_key_tlv_in_flight[8]), .B0(n73), .B1(n73), .S0(n35), .S1(n36), .CO(n37));
Q_AD02 U1975 ( .CI(n37), .A0(num_key_tlv_in_flight[9]), .A1(num_key_tlv_in_flight[10]), .B0(n73), .B1(n73), .S0(n38), .S1(n39), .CO(n40));
Q_AD02 U1976 ( .CI(n40), .A0(num_key_tlv_in_flight[11]), .A1(num_key_tlv_in_flight[12]), .B0(n73), .B1(n73), .S0(n41), .S1(n42), .CO(n43));
Q_AD02 U1977 ( .CI(n43), .A0(num_key_tlv_in_flight[13]), .A1(num_key_tlv_in_flight[14]), .B0(n73), .B1(n73), .S0(n44), .S1(n45), .CO(n46));
Q_AD02 U1978 ( .CI(n46), .A0(num_key_tlv_in_flight[15]), .A1(num_key_tlv_in_flight[16]), .B0(n73), .B1(n73), .S0(n47), .S1(n48), .CO(n49));
Q_AD02 U1979 ( .CI(n49), .A0(num_key_tlv_in_flight[17]), .A1(num_key_tlv_in_flight[18]), .B0(n73), .B1(n73), .S0(n50), .S1(n51), .CO(n52));
Q_AD02 U1980 ( .CI(n52), .A0(num_key_tlv_in_flight[19]), .A1(num_key_tlv_in_flight[20]), .B0(n73), .B1(n73), .S0(n53), .S1(n54), .CO(n55));
Q_AD02 U1981 ( .CI(n55), .A0(num_key_tlv_in_flight[21]), .A1(num_key_tlv_in_flight[22]), .B0(n73), .B1(n73), .S0(n56), .S1(n57), .CO(n58));
Q_AD02 U1982 ( .CI(n58), .A0(num_key_tlv_in_flight[23]), .A1(num_key_tlv_in_flight[24]), .B0(n73), .B1(n73), .S0(n59), .S1(n60), .CO(n61));
Q_AD02 U1983 ( .CI(n61), .A0(num_key_tlv_in_flight[25]), .A1(num_key_tlv_in_flight[26]), .B0(n73), .B1(n73), .S0(n62), .S1(n63), .CO(n64));
Q_AD02 U1984 ( .CI(n64), .A0(num_key_tlv_in_flight[27]), .A1(num_key_tlv_in_flight[28]), .B0(n73), .B1(n73), .S0(n65), .S1(n66), .CO(n67));
Q_AD02 U1985 ( .CI(n67), .A0(num_key_tlv_in_flight[29]), .A1(num_key_tlv_in_flight[30]), .B0(n73), .B1(n73), .S0(n68), .S1(n69), .CO(n70));
Q_XOR2 U1986 ( .A0(tlv_parser_int_tlv_start_pulse), .A1(n73), .Z(n72));
Q_FDP1 kme_idle_REG  ( .CK(clk), .R(rst_n), .D(n74), .Q(kme_idle), .QN( ));
Q_AN02 U1988 ( .A0(n75), .A1(idle_components[3]), .Z(n74));
Q_AN03 U1989 ( .A0(n76), .A1(n77), .A2(n79), .Z(n75));
Q_AN03 U1990 ( .A0(tlv_parser_idle), .A1(drng_idle), .A2(kme_slv_empty), .Z(n76));
Q_AN02 U1991 ( .A0(cddip_key_tlv_rsm_idle[0]), .A1(n78), .Z(n77));
Q_AN03 U1992 ( .A0(cddip_key_tlv_rsm_idle[3]), .A1(cddip_key_tlv_rsm_idle[2]), .A2(cddip_key_tlv_rsm_idle[1]), .Z(n78));
Q_AN02 U1993 ( .A0(cceip_key_tlv_rsm_idle[0]), .A1(n80), .Z(n79));
Q_AN03 U1994 ( .A0(cceip_key_tlv_rsm_idle[3]), .A1(cceip_key_tlv_rsm_idle[2]), .A2(cceip_key_tlv_rsm_idle[1]), .Z(n80));
ixc_assign_10 \num_0_._zz_strnp_2 ( \num_0_._zy_simnet_tvar_7 [0:9], { n85, 
	n84, n83, n82, n81, \sa_ctrl[0][4] , \sa_ctrl[0][3] , 
	\sa_ctrl[0][2] , \sa_ctrl[0][1] , \sa_ctrl[0][0] });
cr_sa_counter \num_0_.sa_counter_i ( .sa_count( 
	\num_0_._zy_simnet_tvar_5 [0:49]), .sa_snapshot( 
	\num_0_._zy_simnet_tvar_6 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_0_._zy_simnet_tvar_7 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_0_._zy_simnet_sa_clear_8_w$ ), 
	.sa_snap( \num_0_._zy_simnet_sa_snap_9_w$ ));
ixc_assign \num_0_._zz_strnp_4 ( \num_0_._zy_simnet_sa_snap_9_w$ , sa_snap);
ixc_assign \num_0_._zz_strnp_3 ( \num_0_._zy_simnet_sa_clear_8_w$ , sa_clear);
ixc_assign_50 \num_0_._zz_strnp_1 ( { \sa_snapshot[0][49] , 
	\sa_snapshot[0][48] , \sa_snapshot[0][47] , \sa_snapshot[0][46] , 
	\sa_snapshot[0][45] , \sa_snapshot[0][44] , \sa_snapshot[0][43] , 
	\sa_snapshot[0][42] , \sa_snapshot[0][41] , \sa_snapshot[0][40] , 
	\sa_snapshot[0][39] , \sa_snapshot[0][38] , \sa_snapshot[0][37] , 
	\sa_snapshot[0][36] , \sa_snapshot[0][35] , \sa_snapshot[0][34] , 
	\sa_snapshot[0][33] , \sa_snapshot[0][32] , \sa_snapshot[0][31] , 
	\sa_snapshot[0][30] , \sa_snapshot[0][29] , \sa_snapshot[0][28] , 
	\sa_snapshot[0][27] , \sa_snapshot[0][26] , \sa_snapshot[0][25] , 
	\sa_snapshot[0][24] , \sa_snapshot[0][23] , \sa_snapshot[0][22] , 
	\sa_snapshot[0][21] , \sa_snapshot[0][20] , \sa_snapshot[0][19] , 
	\sa_snapshot[0][18] , \sa_snapshot[0][17] , \sa_snapshot[0][16] , 
	\sa_snapshot[0][15] , \sa_snapshot[0][14] , \sa_snapshot[0][13] , 
	\sa_snapshot[0][12] , \sa_snapshot[0][11] , \sa_snapshot[0][10] , 
	\sa_snapshot[0][9] , \sa_snapshot[0][8] , \sa_snapshot[0][7] , 
	\sa_snapshot[0][6] , \sa_snapshot[0][5] , \sa_snapshot[0][4] , 
	\sa_snapshot[0][3] , \sa_snapshot[0][2] , \sa_snapshot[0][1] , 
	\sa_snapshot[0][0] }, \num_0_._zy_simnet_tvar_6 [0:49]);
ixc_assign_50 \num_0_._zz_strnp_0 ( { \sa_count[0][49] , \sa_count[0][48] , 
	\sa_count[0][47] , \sa_count[0][46] , \sa_count[0][45] , 
	\sa_count[0][44] , \sa_count[0][43] , \sa_count[0][42] , 
	\sa_count[0][41] , \sa_count[0][40] , \sa_count[0][39] , 
	\sa_count[0][38] , \sa_count[0][37] , \sa_count[0][36] , 
	\sa_count[0][35] , \sa_count[0][34] , \sa_count[0][33] , 
	\sa_count[0][32] , \sa_count[0][31] , \sa_count[0][30] , 
	\sa_count[0][29] , \sa_count[0][28] , \sa_count[0][27] , 
	\sa_count[0][26] , \sa_count[0][25] , \sa_count[0][24] , 
	\sa_count[0][23] , \sa_count[0][22] , \sa_count[0][21] , 
	\sa_count[0][20] , \sa_count[0][19] , \sa_count[0][18] , 
	\sa_count[0][17] , \sa_count[0][16] , \sa_count[0][15] , 
	\sa_count[0][14] , \sa_count[0][13] , \sa_count[0][12] , 
	\sa_count[0][11] , \sa_count[0][10] , \sa_count[0][9] , 
	\sa_count[0][8] , \sa_count[0][7] , \sa_count[0][6] , 
	\sa_count[0][5] , \sa_count[0][4] , \sa_count[0][3] , 
	\sa_count[0][2] , \sa_count[0][1] , \sa_count[0][0] }, 
	\num_0_._zy_simnet_tvar_5 [0:49]);
ixc_assign_10 \num_1_._zz_strnp_7 ( \num_1_._zy_simnet_tvar_12 [0:9], { n90, 
	n89, n88, n87, n86, \sa_ctrl[1][4] , \sa_ctrl[1][3] , 
	\sa_ctrl[1][2] , \sa_ctrl[1][1] , \sa_ctrl[1][0] });
cr_sa_counter \num_1_.sa_counter_i ( .sa_count( 
	\num_1_._zy_simnet_tvar_10 [0:49]), .sa_snapshot( 
	\num_1_._zy_simnet_tvar_11 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_1_._zy_simnet_tvar_12 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_1_._zy_simnet_sa_clear_13_w$ ), 
	.sa_snap( \num_1_._zy_simnet_sa_snap_14_w$ ));
ixc_assign \num_1_._zz_strnp_9 ( \num_1_._zy_simnet_sa_snap_14_w$ , sa_snap);
ixc_assign \num_1_._zz_strnp_8 ( \num_1_._zy_simnet_sa_clear_13_w$ , sa_clear);
ixc_assign_50 \num_1_._zz_strnp_6 ( { \sa_snapshot[1][49] , 
	\sa_snapshot[1][48] , \sa_snapshot[1][47] , \sa_snapshot[1][46] , 
	\sa_snapshot[1][45] , \sa_snapshot[1][44] , \sa_snapshot[1][43] , 
	\sa_snapshot[1][42] , \sa_snapshot[1][41] , \sa_snapshot[1][40] , 
	\sa_snapshot[1][39] , \sa_snapshot[1][38] , \sa_snapshot[1][37] , 
	\sa_snapshot[1][36] , \sa_snapshot[1][35] , \sa_snapshot[1][34] , 
	\sa_snapshot[1][33] , \sa_snapshot[1][32] , \sa_snapshot[1][31] , 
	\sa_snapshot[1][30] , \sa_snapshot[1][29] , \sa_snapshot[1][28] , 
	\sa_snapshot[1][27] , \sa_snapshot[1][26] , \sa_snapshot[1][25] , 
	\sa_snapshot[1][24] , \sa_snapshot[1][23] , \sa_snapshot[1][22] , 
	\sa_snapshot[1][21] , \sa_snapshot[1][20] , \sa_snapshot[1][19] , 
	\sa_snapshot[1][18] , \sa_snapshot[1][17] , \sa_snapshot[1][16] , 
	\sa_snapshot[1][15] , \sa_snapshot[1][14] , \sa_snapshot[1][13] , 
	\sa_snapshot[1][12] , \sa_snapshot[1][11] , \sa_snapshot[1][10] , 
	\sa_snapshot[1][9] , \sa_snapshot[1][8] , \sa_snapshot[1][7] , 
	\sa_snapshot[1][6] , \sa_snapshot[1][5] , \sa_snapshot[1][4] , 
	\sa_snapshot[1][3] , \sa_snapshot[1][2] , \sa_snapshot[1][1] , 
	\sa_snapshot[1][0] }, \num_1_._zy_simnet_tvar_11 [0:49]);
ixc_assign_50 \num_1_._zz_strnp_5 ( { \sa_count[1][49] , \sa_count[1][48] , 
	\sa_count[1][47] , \sa_count[1][46] , \sa_count[1][45] , 
	\sa_count[1][44] , \sa_count[1][43] , \sa_count[1][42] , 
	\sa_count[1][41] , \sa_count[1][40] , \sa_count[1][39] , 
	\sa_count[1][38] , \sa_count[1][37] , \sa_count[1][36] , 
	\sa_count[1][35] , \sa_count[1][34] , \sa_count[1][33] , 
	\sa_count[1][32] , \sa_count[1][31] , \sa_count[1][30] , 
	\sa_count[1][29] , \sa_count[1][28] , \sa_count[1][27] , 
	\sa_count[1][26] , \sa_count[1][25] , \sa_count[1][24] , 
	\sa_count[1][23] , \sa_count[1][22] , \sa_count[1][21] , 
	\sa_count[1][20] , \sa_count[1][19] , \sa_count[1][18] , 
	\sa_count[1][17] , \sa_count[1][16] , \sa_count[1][15] , 
	\sa_count[1][14] , \sa_count[1][13] , \sa_count[1][12] , 
	\sa_count[1][11] , \sa_count[1][10] , \sa_count[1][9] , 
	\sa_count[1][8] , \sa_count[1][7] , \sa_count[1][6] , 
	\sa_count[1][5] , \sa_count[1][4] , \sa_count[1][3] , 
	\sa_count[1][2] , \sa_count[1][1] , \sa_count[1][0] }, 
	\num_1_._zy_simnet_tvar_10 [0:49]);
ixc_assign_10 \num_2_._zz_strnp_12 ( \num_2_._zy_simnet_tvar_17 [0:9], { n95, 
	n94, n93, n92, n91, \sa_ctrl[2][4] , \sa_ctrl[2][3] , 
	\sa_ctrl[2][2] , \sa_ctrl[2][1] , \sa_ctrl[2][0] });
cr_sa_counter \num_2_.sa_counter_i ( .sa_count( 
	\num_2_._zy_simnet_tvar_15 [0:49]), .sa_snapshot( 
	\num_2_._zy_simnet_tvar_16 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_2_._zy_simnet_tvar_17 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_2_._zy_simnet_sa_clear_18_w$ ), 
	.sa_snap( \num_2_._zy_simnet_sa_snap_19_w$ ));
ixc_assign \num_2_._zz_strnp_14 ( \num_2_._zy_simnet_sa_snap_19_w$ , sa_snap);
ixc_assign \num_2_._zz_strnp_13 ( \num_2_._zy_simnet_sa_clear_18_w$ , 
	sa_clear);
ixc_assign_50 \num_2_._zz_strnp_11 ( { \sa_snapshot[2][49] , 
	\sa_snapshot[2][48] , \sa_snapshot[2][47] , \sa_snapshot[2][46] , 
	\sa_snapshot[2][45] , \sa_snapshot[2][44] , \sa_snapshot[2][43] , 
	\sa_snapshot[2][42] , \sa_snapshot[2][41] , \sa_snapshot[2][40] , 
	\sa_snapshot[2][39] , \sa_snapshot[2][38] , \sa_snapshot[2][37] , 
	\sa_snapshot[2][36] , \sa_snapshot[2][35] , \sa_snapshot[2][34] , 
	\sa_snapshot[2][33] , \sa_snapshot[2][32] , \sa_snapshot[2][31] , 
	\sa_snapshot[2][30] , \sa_snapshot[2][29] , \sa_snapshot[2][28] , 
	\sa_snapshot[2][27] , \sa_snapshot[2][26] , \sa_snapshot[2][25] , 
	\sa_snapshot[2][24] , \sa_snapshot[2][23] , \sa_snapshot[2][22] , 
	\sa_snapshot[2][21] , \sa_snapshot[2][20] , \sa_snapshot[2][19] , 
	\sa_snapshot[2][18] , \sa_snapshot[2][17] , \sa_snapshot[2][16] , 
	\sa_snapshot[2][15] , \sa_snapshot[2][14] , \sa_snapshot[2][13] , 
	\sa_snapshot[2][12] , \sa_snapshot[2][11] , \sa_snapshot[2][10] , 
	\sa_snapshot[2][9] , \sa_snapshot[2][8] , \sa_snapshot[2][7] , 
	\sa_snapshot[2][6] , \sa_snapshot[2][5] , \sa_snapshot[2][4] , 
	\sa_snapshot[2][3] , \sa_snapshot[2][2] , \sa_snapshot[2][1] , 
	\sa_snapshot[2][0] }, \num_2_._zy_simnet_tvar_16 [0:49]);
ixc_assign_50 \num_2_._zz_strnp_10 ( { \sa_count[2][49] , \sa_count[2][48] , 
	\sa_count[2][47] , \sa_count[2][46] , \sa_count[2][45] , 
	\sa_count[2][44] , \sa_count[2][43] , \sa_count[2][42] , 
	\sa_count[2][41] , \sa_count[2][40] , \sa_count[2][39] , 
	\sa_count[2][38] , \sa_count[2][37] , \sa_count[2][36] , 
	\sa_count[2][35] , \sa_count[2][34] , \sa_count[2][33] , 
	\sa_count[2][32] , \sa_count[2][31] , \sa_count[2][30] , 
	\sa_count[2][29] , \sa_count[2][28] , \sa_count[2][27] , 
	\sa_count[2][26] , \sa_count[2][25] , \sa_count[2][24] , 
	\sa_count[2][23] , \sa_count[2][22] , \sa_count[2][21] , 
	\sa_count[2][20] , \sa_count[2][19] , \sa_count[2][18] , 
	\sa_count[2][17] , \sa_count[2][16] , \sa_count[2][15] , 
	\sa_count[2][14] , \sa_count[2][13] , \sa_count[2][12] , 
	\sa_count[2][11] , \sa_count[2][10] , \sa_count[2][9] , 
	\sa_count[2][8] , \sa_count[2][7] , \sa_count[2][6] , 
	\sa_count[2][5] , \sa_count[2][4] , \sa_count[2][3] , 
	\sa_count[2][2] , \sa_count[2][1] , \sa_count[2][0] }, 
	\num_2_._zy_simnet_tvar_15 [0:49]);
ixc_assign_10 \num_3_._zz_strnp_17 ( \num_3_._zy_simnet_tvar_22 [0:9], { n100, 
	n99, n98, n97, n96, \sa_ctrl[3][4] , \sa_ctrl[3][3] , 
	\sa_ctrl[3][2] , \sa_ctrl[3][1] , \sa_ctrl[3][0] });
cr_sa_counter \num_3_.sa_counter_i ( .sa_count( 
	\num_3_._zy_simnet_tvar_20 [0:49]), .sa_snapshot( 
	\num_3_._zy_simnet_tvar_21 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_3_._zy_simnet_tvar_22 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_3_._zy_simnet_sa_clear_23_w$ ), 
	.sa_snap( \num_3_._zy_simnet_sa_snap_24_w$ ));
ixc_assign \num_3_._zz_strnp_19 ( \num_3_._zy_simnet_sa_snap_24_w$ , sa_snap);
ixc_assign \num_3_._zz_strnp_18 ( \num_3_._zy_simnet_sa_clear_23_w$ , 
	sa_clear);
ixc_assign_50 \num_3_._zz_strnp_16 ( { \sa_snapshot[3][49] , 
	\sa_snapshot[3][48] , \sa_snapshot[3][47] , \sa_snapshot[3][46] , 
	\sa_snapshot[3][45] , \sa_snapshot[3][44] , \sa_snapshot[3][43] , 
	\sa_snapshot[3][42] , \sa_snapshot[3][41] , \sa_snapshot[3][40] , 
	\sa_snapshot[3][39] , \sa_snapshot[3][38] , \sa_snapshot[3][37] , 
	\sa_snapshot[3][36] , \sa_snapshot[3][35] , \sa_snapshot[3][34] , 
	\sa_snapshot[3][33] , \sa_snapshot[3][32] , \sa_snapshot[3][31] , 
	\sa_snapshot[3][30] , \sa_snapshot[3][29] , \sa_snapshot[3][28] , 
	\sa_snapshot[3][27] , \sa_snapshot[3][26] , \sa_snapshot[3][25] , 
	\sa_snapshot[3][24] , \sa_snapshot[3][23] , \sa_snapshot[3][22] , 
	\sa_snapshot[3][21] , \sa_snapshot[3][20] , \sa_snapshot[3][19] , 
	\sa_snapshot[3][18] , \sa_snapshot[3][17] , \sa_snapshot[3][16] , 
	\sa_snapshot[3][15] , \sa_snapshot[3][14] , \sa_snapshot[3][13] , 
	\sa_snapshot[3][12] , \sa_snapshot[3][11] , \sa_snapshot[3][10] , 
	\sa_snapshot[3][9] , \sa_snapshot[3][8] , \sa_snapshot[3][7] , 
	\sa_snapshot[3][6] , \sa_snapshot[3][5] , \sa_snapshot[3][4] , 
	\sa_snapshot[3][3] , \sa_snapshot[3][2] , \sa_snapshot[3][1] , 
	\sa_snapshot[3][0] }, \num_3_._zy_simnet_tvar_21 [0:49]);
ixc_assign_50 \num_3_._zz_strnp_15 ( { \sa_count[3][49] , \sa_count[3][48] , 
	\sa_count[3][47] , \sa_count[3][46] , \sa_count[3][45] , 
	\sa_count[3][44] , \sa_count[3][43] , \sa_count[3][42] , 
	\sa_count[3][41] , \sa_count[3][40] , \sa_count[3][39] , 
	\sa_count[3][38] , \sa_count[3][37] , \sa_count[3][36] , 
	\sa_count[3][35] , \sa_count[3][34] , \sa_count[3][33] , 
	\sa_count[3][32] , \sa_count[3][31] , \sa_count[3][30] , 
	\sa_count[3][29] , \sa_count[3][28] , \sa_count[3][27] , 
	\sa_count[3][26] , \sa_count[3][25] , \sa_count[3][24] , 
	\sa_count[3][23] , \sa_count[3][22] , \sa_count[3][21] , 
	\sa_count[3][20] , \sa_count[3][19] , \sa_count[3][18] , 
	\sa_count[3][17] , \sa_count[3][16] , \sa_count[3][15] , 
	\sa_count[3][14] , \sa_count[3][13] , \sa_count[3][12] , 
	\sa_count[3][11] , \sa_count[3][10] , \sa_count[3][9] , 
	\sa_count[3][8] , \sa_count[3][7] , \sa_count[3][6] , 
	\sa_count[3][5] , \sa_count[3][4] , \sa_count[3][3] , 
	\sa_count[3][2] , \sa_count[3][1] , \sa_count[3][0] }, 
	\num_3_._zy_simnet_tvar_20 [0:49]);
ixc_assign_10 \num_4_._zz_strnp_22 ( \num_4_._zy_simnet_tvar_27 [0:9], { n105, 
	n104, n103, n102, n101, \sa_ctrl[4][4] , \sa_ctrl[4][3] , 
	\sa_ctrl[4][2] , \sa_ctrl[4][1] , \sa_ctrl[4][0] });
cr_sa_counter \num_4_.sa_counter_i ( .sa_count( 
	\num_4_._zy_simnet_tvar_25 [0:49]), .sa_snapshot( 
	\num_4_._zy_simnet_tvar_26 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_4_._zy_simnet_tvar_27 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_4_._zy_simnet_sa_clear_28_w$ ), 
	.sa_snap( \num_4_._zy_simnet_sa_snap_29_w$ ));
ixc_assign \num_4_._zz_strnp_24 ( \num_4_._zy_simnet_sa_snap_29_w$ , sa_snap);
ixc_assign \num_4_._zz_strnp_23 ( \num_4_._zy_simnet_sa_clear_28_w$ , 
	sa_clear);
ixc_assign_50 \num_4_._zz_strnp_21 ( { \sa_snapshot[4][49] , 
	\sa_snapshot[4][48] , \sa_snapshot[4][47] , \sa_snapshot[4][46] , 
	\sa_snapshot[4][45] , \sa_snapshot[4][44] , \sa_snapshot[4][43] , 
	\sa_snapshot[4][42] , \sa_snapshot[4][41] , \sa_snapshot[4][40] , 
	\sa_snapshot[4][39] , \sa_snapshot[4][38] , \sa_snapshot[4][37] , 
	\sa_snapshot[4][36] , \sa_snapshot[4][35] , \sa_snapshot[4][34] , 
	\sa_snapshot[4][33] , \sa_snapshot[4][32] , \sa_snapshot[4][31] , 
	\sa_snapshot[4][30] , \sa_snapshot[4][29] , \sa_snapshot[4][28] , 
	\sa_snapshot[4][27] , \sa_snapshot[4][26] , \sa_snapshot[4][25] , 
	\sa_snapshot[4][24] , \sa_snapshot[4][23] , \sa_snapshot[4][22] , 
	\sa_snapshot[4][21] , \sa_snapshot[4][20] , \sa_snapshot[4][19] , 
	\sa_snapshot[4][18] , \sa_snapshot[4][17] , \sa_snapshot[4][16] , 
	\sa_snapshot[4][15] , \sa_snapshot[4][14] , \sa_snapshot[4][13] , 
	\sa_snapshot[4][12] , \sa_snapshot[4][11] , \sa_snapshot[4][10] , 
	\sa_snapshot[4][9] , \sa_snapshot[4][8] , \sa_snapshot[4][7] , 
	\sa_snapshot[4][6] , \sa_snapshot[4][5] , \sa_snapshot[4][4] , 
	\sa_snapshot[4][3] , \sa_snapshot[4][2] , \sa_snapshot[4][1] , 
	\sa_snapshot[4][0] }, \num_4_._zy_simnet_tvar_26 [0:49]);
ixc_assign_50 \num_4_._zz_strnp_20 ( { \sa_count[4][49] , \sa_count[4][48] , 
	\sa_count[4][47] , \sa_count[4][46] , \sa_count[4][45] , 
	\sa_count[4][44] , \sa_count[4][43] , \sa_count[4][42] , 
	\sa_count[4][41] , \sa_count[4][40] , \sa_count[4][39] , 
	\sa_count[4][38] , \sa_count[4][37] , \sa_count[4][36] , 
	\sa_count[4][35] , \sa_count[4][34] , \sa_count[4][33] , 
	\sa_count[4][32] , \sa_count[4][31] , \sa_count[4][30] , 
	\sa_count[4][29] , \sa_count[4][28] , \sa_count[4][27] , 
	\sa_count[4][26] , \sa_count[4][25] , \sa_count[4][24] , 
	\sa_count[4][23] , \sa_count[4][22] , \sa_count[4][21] , 
	\sa_count[4][20] , \sa_count[4][19] , \sa_count[4][18] , 
	\sa_count[4][17] , \sa_count[4][16] , \sa_count[4][15] , 
	\sa_count[4][14] , \sa_count[4][13] , \sa_count[4][12] , 
	\sa_count[4][11] , \sa_count[4][10] , \sa_count[4][9] , 
	\sa_count[4][8] , \sa_count[4][7] , \sa_count[4][6] , 
	\sa_count[4][5] , \sa_count[4][4] , \sa_count[4][3] , 
	\sa_count[4][2] , \sa_count[4][1] , \sa_count[4][0] }, 
	\num_4_._zy_simnet_tvar_25 [0:49]);
ixc_assign_10 \num_5_._zz_strnp_27 ( \num_5_._zy_simnet_tvar_32 [0:9], { n110, 
	n109, n108, n107, n106, \sa_ctrl[5][4] , \sa_ctrl[5][3] , 
	\sa_ctrl[5][2] , \sa_ctrl[5][1] , \sa_ctrl[5][0] });
cr_sa_counter \num_5_.sa_counter_i ( .sa_count( 
	\num_5_._zy_simnet_tvar_30 [0:49]), .sa_snapshot( 
	\num_5_._zy_simnet_tvar_31 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_5_._zy_simnet_tvar_32 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_5_._zy_simnet_sa_clear_33_w$ ), 
	.sa_snap( \num_5_._zy_simnet_sa_snap_34_w$ ));
ixc_assign \num_5_._zz_strnp_29 ( \num_5_._zy_simnet_sa_snap_34_w$ , sa_snap);
ixc_assign \num_5_._zz_strnp_28 ( \num_5_._zy_simnet_sa_clear_33_w$ , 
	sa_clear);
ixc_assign_50 \num_5_._zz_strnp_26 ( { \sa_snapshot[5][49] , 
	\sa_snapshot[5][48] , \sa_snapshot[5][47] , \sa_snapshot[5][46] , 
	\sa_snapshot[5][45] , \sa_snapshot[5][44] , \sa_snapshot[5][43] , 
	\sa_snapshot[5][42] , \sa_snapshot[5][41] , \sa_snapshot[5][40] , 
	\sa_snapshot[5][39] , \sa_snapshot[5][38] , \sa_snapshot[5][37] , 
	\sa_snapshot[5][36] , \sa_snapshot[5][35] , \sa_snapshot[5][34] , 
	\sa_snapshot[5][33] , \sa_snapshot[5][32] , \sa_snapshot[5][31] , 
	\sa_snapshot[5][30] , \sa_snapshot[5][29] , \sa_snapshot[5][28] , 
	\sa_snapshot[5][27] , \sa_snapshot[5][26] , \sa_snapshot[5][25] , 
	\sa_snapshot[5][24] , \sa_snapshot[5][23] , \sa_snapshot[5][22] , 
	\sa_snapshot[5][21] , \sa_snapshot[5][20] , \sa_snapshot[5][19] , 
	\sa_snapshot[5][18] , \sa_snapshot[5][17] , \sa_snapshot[5][16] , 
	\sa_snapshot[5][15] , \sa_snapshot[5][14] , \sa_snapshot[5][13] , 
	\sa_snapshot[5][12] , \sa_snapshot[5][11] , \sa_snapshot[5][10] , 
	\sa_snapshot[5][9] , \sa_snapshot[5][8] , \sa_snapshot[5][7] , 
	\sa_snapshot[5][6] , \sa_snapshot[5][5] , \sa_snapshot[5][4] , 
	\sa_snapshot[5][3] , \sa_snapshot[5][2] , \sa_snapshot[5][1] , 
	\sa_snapshot[5][0] }, \num_5_._zy_simnet_tvar_31 [0:49]);
ixc_assign_50 \num_5_._zz_strnp_25 ( { \sa_count[5][49] , \sa_count[5][48] , 
	\sa_count[5][47] , \sa_count[5][46] , \sa_count[5][45] , 
	\sa_count[5][44] , \sa_count[5][43] , \sa_count[5][42] , 
	\sa_count[5][41] , \sa_count[5][40] , \sa_count[5][39] , 
	\sa_count[5][38] , \sa_count[5][37] , \sa_count[5][36] , 
	\sa_count[5][35] , \sa_count[5][34] , \sa_count[5][33] , 
	\sa_count[5][32] , \sa_count[5][31] , \sa_count[5][30] , 
	\sa_count[5][29] , \sa_count[5][28] , \sa_count[5][27] , 
	\sa_count[5][26] , \sa_count[5][25] , \sa_count[5][24] , 
	\sa_count[5][23] , \sa_count[5][22] , \sa_count[5][21] , 
	\sa_count[5][20] , \sa_count[5][19] , \sa_count[5][18] , 
	\sa_count[5][17] , \sa_count[5][16] , \sa_count[5][15] , 
	\sa_count[5][14] , \sa_count[5][13] , \sa_count[5][12] , 
	\sa_count[5][11] , \sa_count[5][10] , \sa_count[5][9] , 
	\sa_count[5][8] , \sa_count[5][7] , \sa_count[5][6] , 
	\sa_count[5][5] , \sa_count[5][4] , \sa_count[5][3] , 
	\sa_count[5][2] , \sa_count[5][1] , \sa_count[5][0] }, 
	\num_5_._zy_simnet_tvar_30 [0:49]);
ixc_assign_10 \num_6_._zz_strnp_32 ( \num_6_._zy_simnet_tvar_37 [0:9], { n115, 
	n114, n113, n112, n111, \sa_ctrl[6][4] , \sa_ctrl[6][3] , 
	\sa_ctrl[6][2] , \sa_ctrl[6][1] , \sa_ctrl[6][0] });
cr_sa_counter \num_6_.sa_counter_i ( .sa_count( 
	\num_6_._zy_simnet_tvar_35 [0:49]), .sa_snapshot( 
	\num_6_._zy_simnet_tvar_36 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_6_._zy_simnet_tvar_37 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_6_._zy_simnet_sa_clear_38_w$ ), 
	.sa_snap( \num_6_._zy_simnet_sa_snap_39_w$ ));
ixc_assign \num_6_._zz_strnp_34 ( \num_6_._zy_simnet_sa_snap_39_w$ , sa_snap);
ixc_assign \num_6_._zz_strnp_33 ( \num_6_._zy_simnet_sa_clear_38_w$ , 
	sa_clear);
ixc_assign_50 \num_6_._zz_strnp_31 ( { \sa_snapshot[6][49] , 
	\sa_snapshot[6][48] , \sa_snapshot[6][47] , \sa_snapshot[6][46] , 
	\sa_snapshot[6][45] , \sa_snapshot[6][44] , \sa_snapshot[6][43] , 
	\sa_snapshot[6][42] , \sa_snapshot[6][41] , \sa_snapshot[6][40] , 
	\sa_snapshot[6][39] , \sa_snapshot[6][38] , \sa_snapshot[6][37] , 
	\sa_snapshot[6][36] , \sa_snapshot[6][35] , \sa_snapshot[6][34] , 
	\sa_snapshot[6][33] , \sa_snapshot[6][32] , \sa_snapshot[6][31] , 
	\sa_snapshot[6][30] , \sa_snapshot[6][29] , \sa_snapshot[6][28] , 
	\sa_snapshot[6][27] , \sa_snapshot[6][26] , \sa_snapshot[6][25] , 
	\sa_snapshot[6][24] , \sa_snapshot[6][23] , \sa_snapshot[6][22] , 
	\sa_snapshot[6][21] , \sa_snapshot[6][20] , \sa_snapshot[6][19] , 
	\sa_snapshot[6][18] , \sa_snapshot[6][17] , \sa_snapshot[6][16] , 
	\sa_snapshot[6][15] , \sa_snapshot[6][14] , \sa_snapshot[6][13] , 
	\sa_snapshot[6][12] , \sa_snapshot[6][11] , \sa_snapshot[6][10] , 
	\sa_snapshot[6][9] , \sa_snapshot[6][8] , \sa_snapshot[6][7] , 
	\sa_snapshot[6][6] , \sa_snapshot[6][5] , \sa_snapshot[6][4] , 
	\sa_snapshot[6][3] , \sa_snapshot[6][2] , \sa_snapshot[6][1] , 
	\sa_snapshot[6][0] }, \num_6_._zy_simnet_tvar_36 [0:49]);
ixc_assign_50 \num_6_._zz_strnp_30 ( { \sa_count[6][49] , \sa_count[6][48] , 
	\sa_count[6][47] , \sa_count[6][46] , \sa_count[6][45] , 
	\sa_count[6][44] , \sa_count[6][43] , \sa_count[6][42] , 
	\sa_count[6][41] , \sa_count[6][40] , \sa_count[6][39] , 
	\sa_count[6][38] , \sa_count[6][37] , \sa_count[6][36] , 
	\sa_count[6][35] , \sa_count[6][34] , \sa_count[6][33] , 
	\sa_count[6][32] , \sa_count[6][31] , \sa_count[6][30] , 
	\sa_count[6][29] , \sa_count[6][28] , \sa_count[6][27] , 
	\sa_count[6][26] , \sa_count[6][25] , \sa_count[6][24] , 
	\sa_count[6][23] , \sa_count[6][22] , \sa_count[6][21] , 
	\sa_count[6][20] , \sa_count[6][19] , \sa_count[6][18] , 
	\sa_count[6][17] , \sa_count[6][16] , \sa_count[6][15] , 
	\sa_count[6][14] , \sa_count[6][13] , \sa_count[6][12] , 
	\sa_count[6][11] , \sa_count[6][10] , \sa_count[6][9] , 
	\sa_count[6][8] , \sa_count[6][7] , \sa_count[6][6] , 
	\sa_count[6][5] , \sa_count[6][4] , \sa_count[6][3] , 
	\sa_count[6][2] , \sa_count[6][1] , \sa_count[6][0] }, 
	\num_6_._zy_simnet_tvar_35 [0:49]);
ixc_assign_10 \num_7_._zz_strnp_37 ( \num_7_._zy_simnet_tvar_42 [0:9], { n120, 
	n119, n118, n117, n116, \sa_ctrl[7][4] , \sa_ctrl[7][3] , 
	\sa_ctrl[7][2] , \sa_ctrl[7][1] , \sa_ctrl[7][0] });
cr_sa_counter \num_7_.sa_counter_i ( .sa_count( 
	\num_7_._zy_simnet_tvar_40 [0:49]), .sa_snapshot( 
	\num_7_._zy_simnet_tvar_41 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_7_._zy_simnet_tvar_42 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_7_._zy_simnet_sa_clear_43_w$ ), 
	.sa_snap( \num_7_._zy_simnet_sa_snap_44_w$ ));
ixc_assign \num_7_._zz_strnp_39 ( \num_7_._zy_simnet_sa_snap_44_w$ , sa_snap);
ixc_assign \num_7_._zz_strnp_38 ( \num_7_._zy_simnet_sa_clear_43_w$ , 
	sa_clear);
ixc_assign_50 \num_7_._zz_strnp_36 ( { \sa_snapshot[7][49] , 
	\sa_snapshot[7][48] , \sa_snapshot[7][47] , \sa_snapshot[7][46] , 
	\sa_snapshot[7][45] , \sa_snapshot[7][44] , \sa_snapshot[7][43] , 
	\sa_snapshot[7][42] , \sa_snapshot[7][41] , \sa_snapshot[7][40] , 
	\sa_snapshot[7][39] , \sa_snapshot[7][38] , \sa_snapshot[7][37] , 
	\sa_snapshot[7][36] , \sa_snapshot[7][35] , \sa_snapshot[7][34] , 
	\sa_snapshot[7][33] , \sa_snapshot[7][32] , \sa_snapshot[7][31] , 
	\sa_snapshot[7][30] , \sa_snapshot[7][29] , \sa_snapshot[7][28] , 
	\sa_snapshot[7][27] , \sa_snapshot[7][26] , \sa_snapshot[7][25] , 
	\sa_snapshot[7][24] , \sa_snapshot[7][23] , \sa_snapshot[7][22] , 
	\sa_snapshot[7][21] , \sa_snapshot[7][20] , \sa_snapshot[7][19] , 
	\sa_snapshot[7][18] , \sa_snapshot[7][17] , \sa_snapshot[7][16] , 
	\sa_snapshot[7][15] , \sa_snapshot[7][14] , \sa_snapshot[7][13] , 
	\sa_snapshot[7][12] , \sa_snapshot[7][11] , \sa_snapshot[7][10] , 
	\sa_snapshot[7][9] , \sa_snapshot[7][8] , \sa_snapshot[7][7] , 
	\sa_snapshot[7][6] , \sa_snapshot[7][5] , \sa_snapshot[7][4] , 
	\sa_snapshot[7][3] , \sa_snapshot[7][2] , \sa_snapshot[7][1] , 
	\sa_snapshot[7][0] }, \num_7_._zy_simnet_tvar_41 [0:49]);
ixc_assign_50 \num_7_._zz_strnp_35 ( { \sa_count[7][49] , \sa_count[7][48] , 
	\sa_count[7][47] , \sa_count[7][46] , \sa_count[7][45] , 
	\sa_count[7][44] , \sa_count[7][43] , \sa_count[7][42] , 
	\sa_count[7][41] , \sa_count[7][40] , \sa_count[7][39] , 
	\sa_count[7][38] , \sa_count[7][37] , \sa_count[7][36] , 
	\sa_count[7][35] , \sa_count[7][34] , \sa_count[7][33] , 
	\sa_count[7][32] , \sa_count[7][31] , \sa_count[7][30] , 
	\sa_count[7][29] , \sa_count[7][28] , \sa_count[7][27] , 
	\sa_count[7][26] , \sa_count[7][25] , \sa_count[7][24] , 
	\sa_count[7][23] , \sa_count[7][22] , \sa_count[7][21] , 
	\sa_count[7][20] , \sa_count[7][19] , \sa_count[7][18] , 
	\sa_count[7][17] , \sa_count[7][16] , \sa_count[7][15] , 
	\sa_count[7][14] , \sa_count[7][13] , \sa_count[7][12] , 
	\sa_count[7][11] , \sa_count[7][10] , \sa_count[7][9] , 
	\sa_count[7][8] , \sa_count[7][7] , \sa_count[7][6] , 
	\sa_count[7][5] , \sa_count[7][4] , \sa_count[7][3] , 
	\sa_count[7][2] , \sa_count[7][1] , \sa_count[7][0] }, 
	\num_7_._zy_simnet_tvar_40 [0:49]);
ixc_assign_10 \num_8_._zz_strnp_42 ( \num_8_._zy_simnet_tvar_47 [0:9], { n125, 
	n124, n123, n122, n121, \sa_ctrl[8][4] , \sa_ctrl[8][3] , 
	\sa_ctrl[8][2] , \sa_ctrl[8][1] , \sa_ctrl[8][0] });
cr_sa_counter \num_8_.sa_counter_i ( .sa_count( 
	\num_8_._zy_simnet_tvar_45 [0:49]), .sa_snapshot( 
	\num_8_._zy_simnet_tvar_46 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_8_._zy_simnet_tvar_47 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_8_._zy_simnet_sa_clear_48_w$ ), 
	.sa_snap( \num_8_._zy_simnet_sa_snap_49_w$ ));
ixc_assign \num_8_._zz_strnp_44 ( \num_8_._zy_simnet_sa_snap_49_w$ , sa_snap);
ixc_assign \num_8_._zz_strnp_43 ( \num_8_._zy_simnet_sa_clear_48_w$ , 
	sa_clear);
ixc_assign_50 \num_8_._zz_strnp_41 ( { \sa_snapshot[8][49] , 
	\sa_snapshot[8][48] , \sa_snapshot[8][47] , \sa_snapshot[8][46] , 
	\sa_snapshot[8][45] , \sa_snapshot[8][44] , \sa_snapshot[8][43] , 
	\sa_snapshot[8][42] , \sa_snapshot[8][41] , \sa_snapshot[8][40] , 
	\sa_snapshot[8][39] , \sa_snapshot[8][38] , \sa_snapshot[8][37] , 
	\sa_snapshot[8][36] , \sa_snapshot[8][35] , \sa_snapshot[8][34] , 
	\sa_snapshot[8][33] , \sa_snapshot[8][32] , \sa_snapshot[8][31] , 
	\sa_snapshot[8][30] , \sa_snapshot[8][29] , \sa_snapshot[8][28] , 
	\sa_snapshot[8][27] , \sa_snapshot[8][26] , \sa_snapshot[8][25] , 
	\sa_snapshot[8][24] , \sa_snapshot[8][23] , \sa_snapshot[8][22] , 
	\sa_snapshot[8][21] , \sa_snapshot[8][20] , \sa_snapshot[8][19] , 
	\sa_snapshot[8][18] , \sa_snapshot[8][17] , \sa_snapshot[8][16] , 
	\sa_snapshot[8][15] , \sa_snapshot[8][14] , \sa_snapshot[8][13] , 
	\sa_snapshot[8][12] , \sa_snapshot[8][11] , \sa_snapshot[8][10] , 
	\sa_snapshot[8][9] , \sa_snapshot[8][8] , \sa_snapshot[8][7] , 
	\sa_snapshot[8][6] , \sa_snapshot[8][5] , \sa_snapshot[8][4] , 
	\sa_snapshot[8][3] , \sa_snapshot[8][2] , \sa_snapshot[8][1] , 
	\sa_snapshot[8][0] }, \num_8_._zy_simnet_tvar_46 [0:49]);
ixc_assign_50 \num_8_._zz_strnp_40 ( { \sa_count[8][49] , \sa_count[8][48] , 
	\sa_count[8][47] , \sa_count[8][46] , \sa_count[8][45] , 
	\sa_count[8][44] , \sa_count[8][43] , \sa_count[8][42] , 
	\sa_count[8][41] , \sa_count[8][40] , \sa_count[8][39] , 
	\sa_count[8][38] , \sa_count[8][37] , \sa_count[8][36] , 
	\sa_count[8][35] , \sa_count[8][34] , \sa_count[8][33] , 
	\sa_count[8][32] , \sa_count[8][31] , \sa_count[8][30] , 
	\sa_count[8][29] , \sa_count[8][28] , \sa_count[8][27] , 
	\sa_count[8][26] , \sa_count[8][25] , \sa_count[8][24] , 
	\sa_count[8][23] , \sa_count[8][22] , \sa_count[8][21] , 
	\sa_count[8][20] , \sa_count[8][19] , \sa_count[8][18] , 
	\sa_count[8][17] , \sa_count[8][16] , \sa_count[8][15] , 
	\sa_count[8][14] , \sa_count[8][13] , \sa_count[8][12] , 
	\sa_count[8][11] , \sa_count[8][10] , \sa_count[8][9] , 
	\sa_count[8][8] , \sa_count[8][7] , \sa_count[8][6] , 
	\sa_count[8][5] , \sa_count[8][4] , \sa_count[8][3] , 
	\sa_count[8][2] , \sa_count[8][1] , \sa_count[8][0] }, 
	\num_8_._zy_simnet_tvar_45 [0:49]);
ixc_assign_10 \num_9_._zz_strnp_47 ( \num_9_._zy_simnet_tvar_52 [0:9], { n130, 
	n129, n128, n127, n126, \sa_ctrl[9][4] , \sa_ctrl[9][3] , 
	\sa_ctrl[9][2] , \sa_ctrl[9][1] , \sa_ctrl[9][0] });
cr_sa_counter \num_9_.sa_counter_i ( .sa_count( 
	\num_9_._zy_simnet_tvar_50 [0:49]), .sa_snapshot( 
	\num_9_._zy_simnet_tvar_51 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_9_._zy_simnet_tvar_52 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_9_._zy_simnet_sa_clear_53_w$ ), 
	.sa_snap( \num_9_._zy_simnet_sa_snap_54_w$ ));
ixc_assign \num_9_._zz_strnp_49 ( \num_9_._zy_simnet_sa_snap_54_w$ , sa_snap);
ixc_assign \num_9_._zz_strnp_48 ( \num_9_._zy_simnet_sa_clear_53_w$ , 
	sa_clear);
ixc_assign_50 \num_9_._zz_strnp_46 ( { \sa_snapshot[9][49] , 
	\sa_snapshot[9][48] , \sa_snapshot[9][47] , \sa_snapshot[9][46] , 
	\sa_snapshot[9][45] , \sa_snapshot[9][44] , \sa_snapshot[9][43] , 
	\sa_snapshot[9][42] , \sa_snapshot[9][41] , \sa_snapshot[9][40] , 
	\sa_snapshot[9][39] , \sa_snapshot[9][38] , \sa_snapshot[9][37] , 
	\sa_snapshot[9][36] , \sa_snapshot[9][35] , \sa_snapshot[9][34] , 
	\sa_snapshot[9][33] , \sa_snapshot[9][32] , \sa_snapshot[9][31] , 
	\sa_snapshot[9][30] , \sa_snapshot[9][29] , \sa_snapshot[9][28] , 
	\sa_snapshot[9][27] , \sa_snapshot[9][26] , \sa_snapshot[9][25] , 
	\sa_snapshot[9][24] , \sa_snapshot[9][23] , \sa_snapshot[9][22] , 
	\sa_snapshot[9][21] , \sa_snapshot[9][20] , \sa_snapshot[9][19] , 
	\sa_snapshot[9][18] , \sa_snapshot[9][17] , \sa_snapshot[9][16] , 
	\sa_snapshot[9][15] , \sa_snapshot[9][14] , \sa_snapshot[9][13] , 
	\sa_snapshot[9][12] , \sa_snapshot[9][11] , \sa_snapshot[9][10] , 
	\sa_snapshot[9][9] , \sa_snapshot[9][8] , \sa_snapshot[9][7] , 
	\sa_snapshot[9][6] , \sa_snapshot[9][5] , \sa_snapshot[9][4] , 
	\sa_snapshot[9][3] , \sa_snapshot[9][2] , \sa_snapshot[9][1] , 
	\sa_snapshot[9][0] }, \num_9_._zy_simnet_tvar_51 [0:49]);
ixc_assign_50 \num_9_._zz_strnp_45 ( { \sa_count[9][49] , \sa_count[9][48] , 
	\sa_count[9][47] , \sa_count[9][46] , \sa_count[9][45] , 
	\sa_count[9][44] , \sa_count[9][43] , \sa_count[9][42] , 
	\sa_count[9][41] , \sa_count[9][40] , \sa_count[9][39] , 
	\sa_count[9][38] , \sa_count[9][37] , \sa_count[9][36] , 
	\sa_count[9][35] , \sa_count[9][34] , \sa_count[9][33] , 
	\sa_count[9][32] , \sa_count[9][31] , \sa_count[9][30] , 
	\sa_count[9][29] , \sa_count[9][28] , \sa_count[9][27] , 
	\sa_count[9][26] , \sa_count[9][25] , \sa_count[9][24] , 
	\sa_count[9][23] , \sa_count[9][22] , \sa_count[9][21] , 
	\sa_count[9][20] , \sa_count[9][19] , \sa_count[9][18] , 
	\sa_count[9][17] , \sa_count[9][16] , \sa_count[9][15] , 
	\sa_count[9][14] , \sa_count[9][13] , \sa_count[9][12] , 
	\sa_count[9][11] , \sa_count[9][10] , \sa_count[9][9] , 
	\sa_count[9][8] , \sa_count[9][7] , \sa_count[9][6] , 
	\sa_count[9][5] , \sa_count[9][4] , \sa_count[9][3] , 
	\sa_count[9][2] , \sa_count[9][1] , \sa_count[9][0] }, 
	\num_9_._zy_simnet_tvar_50 [0:49]);
ixc_assign_10 \num_10_._zz_strnp_52 ( \num_10_._zy_simnet_tvar_57 [0:9], { 
	n135, n134, n133, n132, n131, \sa_ctrl[10][4] , \sa_ctrl[10][3] , 
	\sa_ctrl[10][2] , \sa_ctrl[10][1] , \sa_ctrl[10][0] });
cr_sa_counter \num_10_.sa_counter_i ( .sa_count( 
	\num_10_._zy_simnet_tvar_55 [0:49]), .sa_snapshot( 
	\num_10_._zy_simnet_tvar_56 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_10_._zy_simnet_tvar_57 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_10_._zy_simnet_sa_clear_58_w$ ), 
	.sa_snap( \num_10_._zy_simnet_sa_snap_59_w$ ));
ixc_assign \num_10_._zz_strnp_54 ( \num_10_._zy_simnet_sa_snap_59_w$ , 
	sa_snap);
ixc_assign \num_10_._zz_strnp_53 ( \num_10_._zy_simnet_sa_clear_58_w$ , 
	sa_clear);
ixc_assign_50 \num_10_._zz_strnp_51 ( { \sa_snapshot[10][49] , 
	\sa_snapshot[10][48] , \sa_snapshot[10][47] , \sa_snapshot[10][46] , 
	\sa_snapshot[10][45] , \sa_snapshot[10][44] , \sa_snapshot[10][43] , 
	\sa_snapshot[10][42] , \sa_snapshot[10][41] , \sa_snapshot[10][40] , 
	\sa_snapshot[10][39] , \sa_snapshot[10][38] , \sa_snapshot[10][37] , 
	\sa_snapshot[10][36] , \sa_snapshot[10][35] , \sa_snapshot[10][34] , 
	\sa_snapshot[10][33] , \sa_snapshot[10][32] , \sa_snapshot[10][31] , 
	\sa_snapshot[10][30] , \sa_snapshot[10][29] , \sa_snapshot[10][28] , 
	\sa_snapshot[10][27] , \sa_snapshot[10][26] , \sa_snapshot[10][25] , 
	\sa_snapshot[10][24] , \sa_snapshot[10][23] , \sa_snapshot[10][22] , 
	\sa_snapshot[10][21] , \sa_snapshot[10][20] , \sa_snapshot[10][19] , 
	\sa_snapshot[10][18] , \sa_snapshot[10][17] , \sa_snapshot[10][16] , 
	\sa_snapshot[10][15] , \sa_snapshot[10][14] , \sa_snapshot[10][13] , 
	\sa_snapshot[10][12] , \sa_snapshot[10][11] , \sa_snapshot[10][10] , 
	\sa_snapshot[10][9] , \sa_snapshot[10][8] , \sa_snapshot[10][7] , 
	\sa_snapshot[10][6] , \sa_snapshot[10][5] , \sa_snapshot[10][4] , 
	\sa_snapshot[10][3] , \sa_snapshot[10][2] , \sa_snapshot[10][1] , 
	\sa_snapshot[10][0] }, \num_10_._zy_simnet_tvar_56 [0:49]);
ixc_assign_50 \num_10_._zz_strnp_50 ( { \sa_count[10][49] , 
	\sa_count[10][48] , \sa_count[10][47] , \sa_count[10][46] , 
	\sa_count[10][45] , \sa_count[10][44] , \sa_count[10][43] , 
	\sa_count[10][42] , \sa_count[10][41] , \sa_count[10][40] , 
	\sa_count[10][39] , \sa_count[10][38] , \sa_count[10][37] , 
	\sa_count[10][36] , \sa_count[10][35] , \sa_count[10][34] , 
	\sa_count[10][33] , \sa_count[10][32] , \sa_count[10][31] , 
	\sa_count[10][30] , \sa_count[10][29] , \sa_count[10][28] , 
	\sa_count[10][27] , \sa_count[10][26] , \sa_count[10][25] , 
	\sa_count[10][24] , \sa_count[10][23] , \sa_count[10][22] , 
	\sa_count[10][21] , \sa_count[10][20] , \sa_count[10][19] , 
	\sa_count[10][18] , \sa_count[10][17] , \sa_count[10][16] , 
	\sa_count[10][15] , \sa_count[10][14] , \sa_count[10][13] , 
	\sa_count[10][12] , \sa_count[10][11] , \sa_count[10][10] , 
	\sa_count[10][9] , \sa_count[10][8] , \sa_count[10][7] , 
	\sa_count[10][6] , \sa_count[10][5] , \sa_count[10][4] , 
	\sa_count[10][3] , \sa_count[10][2] , \sa_count[10][1] , 
	\sa_count[10][0] }, \num_10_._zy_simnet_tvar_55 [0:49]);
ixc_assign_10 \num_11_._zz_strnp_57 ( \num_11_._zy_simnet_tvar_62 [0:9], { 
	n140, n139, n138, n137, n136, \sa_ctrl[11][4] , \sa_ctrl[11][3] , 
	\sa_ctrl[11][2] , \sa_ctrl[11][1] , \sa_ctrl[11][0] });
cr_sa_counter \num_11_.sa_counter_i ( .sa_count( 
	\num_11_._zy_simnet_tvar_60 [0:49]), .sa_snapshot( 
	\num_11_._zy_simnet_tvar_61 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_11_._zy_simnet_tvar_62 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_11_._zy_simnet_sa_clear_63_w$ ), 
	.sa_snap( \num_11_._zy_simnet_sa_snap_64_w$ ));
ixc_assign \num_11_._zz_strnp_59 ( \num_11_._zy_simnet_sa_snap_64_w$ , 
	sa_snap);
ixc_assign \num_11_._zz_strnp_58 ( \num_11_._zy_simnet_sa_clear_63_w$ , 
	sa_clear);
ixc_assign_50 \num_11_._zz_strnp_56 ( { \sa_snapshot[11][49] , 
	\sa_snapshot[11][48] , \sa_snapshot[11][47] , \sa_snapshot[11][46] , 
	\sa_snapshot[11][45] , \sa_snapshot[11][44] , \sa_snapshot[11][43] , 
	\sa_snapshot[11][42] , \sa_snapshot[11][41] , \sa_snapshot[11][40] , 
	\sa_snapshot[11][39] , \sa_snapshot[11][38] , \sa_snapshot[11][37] , 
	\sa_snapshot[11][36] , \sa_snapshot[11][35] , \sa_snapshot[11][34] , 
	\sa_snapshot[11][33] , \sa_snapshot[11][32] , \sa_snapshot[11][31] , 
	\sa_snapshot[11][30] , \sa_snapshot[11][29] , \sa_snapshot[11][28] , 
	\sa_snapshot[11][27] , \sa_snapshot[11][26] , \sa_snapshot[11][25] , 
	\sa_snapshot[11][24] , \sa_snapshot[11][23] , \sa_snapshot[11][22] , 
	\sa_snapshot[11][21] , \sa_snapshot[11][20] , \sa_snapshot[11][19] , 
	\sa_snapshot[11][18] , \sa_snapshot[11][17] , \sa_snapshot[11][16] , 
	\sa_snapshot[11][15] , \sa_snapshot[11][14] , \sa_snapshot[11][13] , 
	\sa_snapshot[11][12] , \sa_snapshot[11][11] , \sa_snapshot[11][10] , 
	\sa_snapshot[11][9] , \sa_snapshot[11][8] , \sa_snapshot[11][7] , 
	\sa_snapshot[11][6] , \sa_snapshot[11][5] , \sa_snapshot[11][4] , 
	\sa_snapshot[11][3] , \sa_snapshot[11][2] , \sa_snapshot[11][1] , 
	\sa_snapshot[11][0] }, \num_11_._zy_simnet_tvar_61 [0:49]);
ixc_assign_50 \num_11_._zz_strnp_55 ( { \sa_count[11][49] , 
	\sa_count[11][48] , \sa_count[11][47] , \sa_count[11][46] , 
	\sa_count[11][45] , \sa_count[11][44] , \sa_count[11][43] , 
	\sa_count[11][42] , \sa_count[11][41] , \sa_count[11][40] , 
	\sa_count[11][39] , \sa_count[11][38] , \sa_count[11][37] , 
	\sa_count[11][36] , \sa_count[11][35] , \sa_count[11][34] , 
	\sa_count[11][33] , \sa_count[11][32] , \sa_count[11][31] , 
	\sa_count[11][30] , \sa_count[11][29] , \sa_count[11][28] , 
	\sa_count[11][27] , \sa_count[11][26] , \sa_count[11][25] , 
	\sa_count[11][24] , \sa_count[11][23] , \sa_count[11][22] , 
	\sa_count[11][21] , \sa_count[11][20] , \sa_count[11][19] , 
	\sa_count[11][18] , \sa_count[11][17] , \sa_count[11][16] , 
	\sa_count[11][15] , \sa_count[11][14] , \sa_count[11][13] , 
	\sa_count[11][12] , \sa_count[11][11] , \sa_count[11][10] , 
	\sa_count[11][9] , \sa_count[11][8] , \sa_count[11][7] , 
	\sa_count[11][6] , \sa_count[11][5] , \sa_count[11][4] , 
	\sa_count[11][3] , \sa_count[11][2] , \sa_count[11][1] , 
	\sa_count[11][0] }, \num_11_._zy_simnet_tvar_60 [0:49]);
ixc_assign_10 \num_12_._zz_strnp_62 ( \num_12_._zy_simnet_tvar_67 [0:9], { 
	n145, n144, n143, n142, n141, \sa_ctrl[12][4] , \sa_ctrl[12][3] , 
	\sa_ctrl[12][2] , \sa_ctrl[12][1] , \sa_ctrl[12][0] });
cr_sa_counter \num_12_.sa_counter_i ( .sa_count( 
	\num_12_._zy_simnet_tvar_65 [0:49]), .sa_snapshot( 
	\num_12_._zy_simnet_tvar_66 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_12_._zy_simnet_tvar_67 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_12_._zy_simnet_sa_clear_68_w$ ), 
	.sa_snap( \num_12_._zy_simnet_sa_snap_69_w$ ));
ixc_assign \num_12_._zz_strnp_64 ( \num_12_._zy_simnet_sa_snap_69_w$ , 
	sa_snap);
ixc_assign \num_12_._zz_strnp_63 ( \num_12_._zy_simnet_sa_clear_68_w$ , 
	sa_clear);
ixc_assign_50 \num_12_._zz_strnp_61 ( { \sa_snapshot[12][49] , 
	\sa_snapshot[12][48] , \sa_snapshot[12][47] , \sa_snapshot[12][46] , 
	\sa_snapshot[12][45] , \sa_snapshot[12][44] , \sa_snapshot[12][43] , 
	\sa_snapshot[12][42] , \sa_snapshot[12][41] , \sa_snapshot[12][40] , 
	\sa_snapshot[12][39] , \sa_snapshot[12][38] , \sa_snapshot[12][37] , 
	\sa_snapshot[12][36] , \sa_snapshot[12][35] , \sa_snapshot[12][34] , 
	\sa_snapshot[12][33] , \sa_snapshot[12][32] , \sa_snapshot[12][31] , 
	\sa_snapshot[12][30] , \sa_snapshot[12][29] , \sa_snapshot[12][28] , 
	\sa_snapshot[12][27] , \sa_snapshot[12][26] , \sa_snapshot[12][25] , 
	\sa_snapshot[12][24] , \sa_snapshot[12][23] , \sa_snapshot[12][22] , 
	\sa_snapshot[12][21] , \sa_snapshot[12][20] , \sa_snapshot[12][19] , 
	\sa_snapshot[12][18] , \sa_snapshot[12][17] , \sa_snapshot[12][16] , 
	\sa_snapshot[12][15] , \sa_snapshot[12][14] , \sa_snapshot[12][13] , 
	\sa_snapshot[12][12] , \sa_snapshot[12][11] , \sa_snapshot[12][10] , 
	\sa_snapshot[12][9] , \sa_snapshot[12][8] , \sa_snapshot[12][7] , 
	\sa_snapshot[12][6] , \sa_snapshot[12][5] , \sa_snapshot[12][4] , 
	\sa_snapshot[12][3] , \sa_snapshot[12][2] , \sa_snapshot[12][1] , 
	\sa_snapshot[12][0] }, \num_12_._zy_simnet_tvar_66 [0:49]);
ixc_assign_50 \num_12_._zz_strnp_60 ( { \sa_count[12][49] , 
	\sa_count[12][48] , \sa_count[12][47] , \sa_count[12][46] , 
	\sa_count[12][45] , \sa_count[12][44] , \sa_count[12][43] , 
	\sa_count[12][42] , \sa_count[12][41] , \sa_count[12][40] , 
	\sa_count[12][39] , \sa_count[12][38] , \sa_count[12][37] , 
	\sa_count[12][36] , \sa_count[12][35] , \sa_count[12][34] , 
	\sa_count[12][33] , \sa_count[12][32] , \sa_count[12][31] , 
	\sa_count[12][30] , \sa_count[12][29] , \sa_count[12][28] , 
	\sa_count[12][27] , \sa_count[12][26] , \sa_count[12][25] , 
	\sa_count[12][24] , \sa_count[12][23] , \sa_count[12][22] , 
	\sa_count[12][21] , \sa_count[12][20] , \sa_count[12][19] , 
	\sa_count[12][18] , \sa_count[12][17] , \sa_count[12][16] , 
	\sa_count[12][15] , \sa_count[12][14] , \sa_count[12][13] , 
	\sa_count[12][12] , \sa_count[12][11] , \sa_count[12][10] , 
	\sa_count[12][9] , \sa_count[12][8] , \sa_count[12][7] , 
	\sa_count[12][6] , \sa_count[12][5] , \sa_count[12][4] , 
	\sa_count[12][3] , \sa_count[12][2] , \sa_count[12][1] , 
	\sa_count[12][0] }, \num_12_._zy_simnet_tvar_65 [0:49]);
ixc_assign_10 \num_13_._zz_strnp_67 ( \num_13_._zy_simnet_tvar_72 [0:9], { 
	n150, n149, n148, n147, n146, \sa_ctrl[13][4] , \sa_ctrl[13][3] , 
	\sa_ctrl[13][2] , \sa_ctrl[13][1] , \sa_ctrl[13][0] });
cr_sa_counter \num_13_.sa_counter_i ( .sa_count( 
	\num_13_._zy_simnet_tvar_70 [0:49]), .sa_snapshot( 
	\num_13_._zy_simnet_tvar_71 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_13_._zy_simnet_tvar_72 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_13_._zy_simnet_sa_clear_73_w$ ), 
	.sa_snap( \num_13_._zy_simnet_sa_snap_74_w$ ));
ixc_assign \num_13_._zz_strnp_69 ( \num_13_._zy_simnet_sa_snap_74_w$ , 
	sa_snap);
ixc_assign \num_13_._zz_strnp_68 ( \num_13_._zy_simnet_sa_clear_73_w$ , 
	sa_clear);
ixc_assign_50 \num_13_._zz_strnp_66 ( { \sa_snapshot[13][49] , 
	\sa_snapshot[13][48] , \sa_snapshot[13][47] , \sa_snapshot[13][46] , 
	\sa_snapshot[13][45] , \sa_snapshot[13][44] , \sa_snapshot[13][43] , 
	\sa_snapshot[13][42] , \sa_snapshot[13][41] , \sa_snapshot[13][40] , 
	\sa_snapshot[13][39] , \sa_snapshot[13][38] , \sa_snapshot[13][37] , 
	\sa_snapshot[13][36] , \sa_snapshot[13][35] , \sa_snapshot[13][34] , 
	\sa_snapshot[13][33] , \sa_snapshot[13][32] , \sa_snapshot[13][31] , 
	\sa_snapshot[13][30] , \sa_snapshot[13][29] , \sa_snapshot[13][28] , 
	\sa_snapshot[13][27] , \sa_snapshot[13][26] , \sa_snapshot[13][25] , 
	\sa_snapshot[13][24] , \sa_snapshot[13][23] , \sa_snapshot[13][22] , 
	\sa_snapshot[13][21] , \sa_snapshot[13][20] , \sa_snapshot[13][19] , 
	\sa_snapshot[13][18] , \sa_snapshot[13][17] , \sa_snapshot[13][16] , 
	\sa_snapshot[13][15] , \sa_snapshot[13][14] , \sa_snapshot[13][13] , 
	\sa_snapshot[13][12] , \sa_snapshot[13][11] , \sa_snapshot[13][10] , 
	\sa_snapshot[13][9] , \sa_snapshot[13][8] , \sa_snapshot[13][7] , 
	\sa_snapshot[13][6] , \sa_snapshot[13][5] , \sa_snapshot[13][4] , 
	\sa_snapshot[13][3] , \sa_snapshot[13][2] , \sa_snapshot[13][1] , 
	\sa_snapshot[13][0] }, \num_13_._zy_simnet_tvar_71 [0:49]);
ixc_assign_50 \num_13_._zz_strnp_65 ( { \sa_count[13][49] , 
	\sa_count[13][48] , \sa_count[13][47] , \sa_count[13][46] , 
	\sa_count[13][45] , \sa_count[13][44] , \sa_count[13][43] , 
	\sa_count[13][42] , \sa_count[13][41] , \sa_count[13][40] , 
	\sa_count[13][39] , \sa_count[13][38] , \sa_count[13][37] , 
	\sa_count[13][36] , \sa_count[13][35] , \sa_count[13][34] , 
	\sa_count[13][33] , \sa_count[13][32] , \sa_count[13][31] , 
	\sa_count[13][30] , \sa_count[13][29] , \sa_count[13][28] , 
	\sa_count[13][27] , \sa_count[13][26] , \sa_count[13][25] , 
	\sa_count[13][24] , \sa_count[13][23] , \sa_count[13][22] , 
	\sa_count[13][21] , \sa_count[13][20] , \sa_count[13][19] , 
	\sa_count[13][18] , \sa_count[13][17] , \sa_count[13][16] , 
	\sa_count[13][15] , \sa_count[13][14] , \sa_count[13][13] , 
	\sa_count[13][12] , \sa_count[13][11] , \sa_count[13][10] , 
	\sa_count[13][9] , \sa_count[13][8] , \sa_count[13][7] , 
	\sa_count[13][6] , \sa_count[13][5] , \sa_count[13][4] , 
	\sa_count[13][3] , \sa_count[13][2] , \sa_count[13][1] , 
	\sa_count[13][0] }, \num_13_._zy_simnet_tvar_70 [0:49]);
ixc_assign_10 \num_14_._zz_strnp_72 ( \num_14_._zy_simnet_tvar_77 [0:9], { 
	n155, n154, n153, n152, n151, \sa_ctrl[14][4] , \sa_ctrl[14][3] , 
	\sa_ctrl[14][2] , \sa_ctrl[14][1] , \sa_ctrl[14][0] });
cr_sa_counter \num_14_.sa_counter_i ( .sa_count( 
	\num_14_._zy_simnet_tvar_75 [0:49]), .sa_snapshot( 
	\num_14_._zy_simnet_tvar_76 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_14_._zy_simnet_tvar_77 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_14_._zy_simnet_sa_clear_78_w$ ), 
	.sa_snap( \num_14_._zy_simnet_sa_snap_79_w$ ));
ixc_assign \num_14_._zz_strnp_74 ( \num_14_._zy_simnet_sa_snap_79_w$ , 
	sa_snap);
ixc_assign \num_14_._zz_strnp_73 ( \num_14_._zy_simnet_sa_clear_78_w$ , 
	sa_clear);
ixc_assign_50 \num_14_._zz_strnp_71 ( { \sa_snapshot[14][49] , 
	\sa_snapshot[14][48] , \sa_snapshot[14][47] , \sa_snapshot[14][46] , 
	\sa_snapshot[14][45] , \sa_snapshot[14][44] , \sa_snapshot[14][43] , 
	\sa_snapshot[14][42] , \sa_snapshot[14][41] , \sa_snapshot[14][40] , 
	\sa_snapshot[14][39] , \sa_snapshot[14][38] , \sa_snapshot[14][37] , 
	\sa_snapshot[14][36] , \sa_snapshot[14][35] , \sa_snapshot[14][34] , 
	\sa_snapshot[14][33] , \sa_snapshot[14][32] , \sa_snapshot[14][31] , 
	\sa_snapshot[14][30] , \sa_snapshot[14][29] , \sa_snapshot[14][28] , 
	\sa_snapshot[14][27] , \sa_snapshot[14][26] , \sa_snapshot[14][25] , 
	\sa_snapshot[14][24] , \sa_snapshot[14][23] , \sa_snapshot[14][22] , 
	\sa_snapshot[14][21] , \sa_snapshot[14][20] , \sa_snapshot[14][19] , 
	\sa_snapshot[14][18] , \sa_snapshot[14][17] , \sa_snapshot[14][16] , 
	\sa_snapshot[14][15] , \sa_snapshot[14][14] , \sa_snapshot[14][13] , 
	\sa_snapshot[14][12] , \sa_snapshot[14][11] , \sa_snapshot[14][10] , 
	\sa_snapshot[14][9] , \sa_snapshot[14][8] , \sa_snapshot[14][7] , 
	\sa_snapshot[14][6] , \sa_snapshot[14][5] , \sa_snapshot[14][4] , 
	\sa_snapshot[14][3] , \sa_snapshot[14][2] , \sa_snapshot[14][1] , 
	\sa_snapshot[14][0] }, \num_14_._zy_simnet_tvar_76 [0:49]);
ixc_assign_50 \num_14_._zz_strnp_70 ( { \sa_count[14][49] , 
	\sa_count[14][48] , \sa_count[14][47] , \sa_count[14][46] , 
	\sa_count[14][45] , \sa_count[14][44] , \sa_count[14][43] , 
	\sa_count[14][42] , \sa_count[14][41] , \sa_count[14][40] , 
	\sa_count[14][39] , \sa_count[14][38] , \sa_count[14][37] , 
	\sa_count[14][36] , \sa_count[14][35] , \sa_count[14][34] , 
	\sa_count[14][33] , \sa_count[14][32] , \sa_count[14][31] , 
	\sa_count[14][30] , \sa_count[14][29] , \sa_count[14][28] , 
	\sa_count[14][27] , \sa_count[14][26] , \sa_count[14][25] , 
	\sa_count[14][24] , \sa_count[14][23] , \sa_count[14][22] , 
	\sa_count[14][21] , \sa_count[14][20] , \sa_count[14][19] , 
	\sa_count[14][18] , \sa_count[14][17] , \sa_count[14][16] , 
	\sa_count[14][15] , \sa_count[14][14] , \sa_count[14][13] , 
	\sa_count[14][12] , \sa_count[14][11] , \sa_count[14][10] , 
	\sa_count[14][9] , \sa_count[14][8] , \sa_count[14][7] , 
	\sa_count[14][6] , \sa_count[14][5] , \sa_count[14][4] , 
	\sa_count[14][3] , \sa_count[14][2] , \sa_count[14][1] , 
	\sa_count[14][0] }, \num_14_._zy_simnet_tvar_75 [0:49]);
ixc_assign_10 \num_15_._zz_strnp_77 ( \num_15_._zy_simnet_tvar_82 [0:9], { 
	n160, n159, n158, n157, n156, \sa_ctrl[15][4] , \sa_ctrl[15][3] , 
	\sa_ctrl[15][2] , \sa_ctrl[15][1] , \sa_ctrl[15][0] });
cr_sa_counter \num_15_.sa_counter_i ( .sa_count( 
	\num_15_._zy_simnet_tvar_80 [0:49]), .sa_snapshot( 
	\num_15_._zy_simnet_tvar_81 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_15_._zy_simnet_tvar_82 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_15_._zy_simnet_sa_clear_83_w$ ), 
	.sa_snap( \num_15_._zy_simnet_sa_snap_84_w$ ));
ixc_assign \num_15_._zz_strnp_79 ( \num_15_._zy_simnet_sa_snap_84_w$ , 
	sa_snap);
ixc_assign \num_15_._zz_strnp_78 ( \num_15_._zy_simnet_sa_clear_83_w$ , 
	sa_clear);
ixc_assign_50 \num_15_._zz_strnp_76 ( { \sa_snapshot[15][49] , 
	\sa_snapshot[15][48] , \sa_snapshot[15][47] , \sa_snapshot[15][46] , 
	\sa_snapshot[15][45] , \sa_snapshot[15][44] , \sa_snapshot[15][43] , 
	\sa_snapshot[15][42] , \sa_snapshot[15][41] , \sa_snapshot[15][40] , 
	\sa_snapshot[15][39] , \sa_snapshot[15][38] , \sa_snapshot[15][37] , 
	\sa_snapshot[15][36] , \sa_snapshot[15][35] , \sa_snapshot[15][34] , 
	\sa_snapshot[15][33] , \sa_snapshot[15][32] , \sa_snapshot[15][31] , 
	\sa_snapshot[15][30] , \sa_snapshot[15][29] , \sa_snapshot[15][28] , 
	\sa_snapshot[15][27] , \sa_snapshot[15][26] , \sa_snapshot[15][25] , 
	\sa_snapshot[15][24] , \sa_snapshot[15][23] , \sa_snapshot[15][22] , 
	\sa_snapshot[15][21] , \sa_snapshot[15][20] , \sa_snapshot[15][19] , 
	\sa_snapshot[15][18] , \sa_snapshot[15][17] , \sa_snapshot[15][16] , 
	\sa_snapshot[15][15] , \sa_snapshot[15][14] , \sa_snapshot[15][13] , 
	\sa_snapshot[15][12] , \sa_snapshot[15][11] , \sa_snapshot[15][10] , 
	\sa_snapshot[15][9] , \sa_snapshot[15][8] , \sa_snapshot[15][7] , 
	\sa_snapshot[15][6] , \sa_snapshot[15][5] , \sa_snapshot[15][4] , 
	\sa_snapshot[15][3] , \sa_snapshot[15][2] , \sa_snapshot[15][1] , 
	\sa_snapshot[15][0] }, \num_15_._zy_simnet_tvar_81 [0:49]);
ixc_assign_50 \num_15_._zz_strnp_75 ( { \sa_count[15][49] , 
	\sa_count[15][48] , \sa_count[15][47] , \sa_count[15][46] , 
	\sa_count[15][45] , \sa_count[15][44] , \sa_count[15][43] , 
	\sa_count[15][42] , \sa_count[15][41] , \sa_count[15][40] , 
	\sa_count[15][39] , \sa_count[15][38] , \sa_count[15][37] , 
	\sa_count[15][36] , \sa_count[15][35] , \sa_count[15][34] , 
	\sa_count[15][33] , \sa_count[15][32] , \sa_count[15][31] , 
	\sa_count[15][30] , \sa_count[15][29] , \sa_count[15][28] , 
	\sa_count[15][27] , \sa_count[15][26] , \sa_count[15][25] , 
	\sa_count[15][24] , \sa_count[15][23] , \sa_count[15][22] , 
	\sa_count[15][21] , \sa_count[15][20] , \sa_count[15][19] , 
	\sa_count[15][18] , \sa_count[15][17] , \sa_count[15][16] , 
	\sa_count[15][15] , \sa_count[15][14] , \sa_count[15][13] , 
	\sa_count[15][12] , \sa_count[15][11] , \sa_count[15][10] , 
	\sa_count[15][9] , \sa_count[15][8] , \sa_count[15][7] , 
	\sa_count[15][6] , \sa_count[15][5] , \sa_count[15][4] , 
	\sa_count[15][3] , \sa_count[15][2] , \sa_count[15][1] , 
	\sa_count[15][0] }, \num_15_._zy_simnet_tvar_80 [0:49]);
ixc_assign_10 \num_16_._zz_strnp_82 ( \num_16_._zy_simnet_tvar_87 [0:9], { 
	n165, n164, n163, n162, n161, \sa_ctrl[16][4] , \sa_ctrl[16][3] , 
	\sa_ctrl[16][2] , \sa_ctrl[16][1] , \sa_ctrl[16][0] });
cr_sa_counter \num_16_.sa_counter_i ( .sa_count( 
	\num_16_._zy_simnet_tvar_85 [0:49]), .sa_snapshot( 
	\num_16_._zy_simnet_tvar_86 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_16_._zy_simnet_tvar_87 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_16_._zy_simnet_sa_clear_88_w$ ), 
	.sa_snap( \num_16_._zy_simnet_sa_snap_89_w$ ));
ixc_assign \num_16_._zz_strnp_84 ( \num_16_._zy_simnet_sa_snap_89_w$ , 
	sa_snap);
ixc_assign \num_16_._zz_strnp_83 ( \num_16_._zy_simnet_sa_clear_88_w$ , 
	sa_clear);
ixc_assign_50 \num_16_._zz_strnp_81 ( { \sa_snapshot[16][49] , 
	\sa_snapshot[16][48] , \sa_snapshot[16][47] , \sa_snapshot[16][46] , 
	\sa_snapshot[16][45] , \sa_snapshot[16][44] , \sa_snapshot[16][43] , 
	\sa_snapshot[16][42] , \sa_snapshot[16][41] , \sa_snapshot[16][40] , 
	\sa_snapshot[16][39] , \sa_snapshot[16][38] , \sa_snapshot[16][37] , 
	\sa_snapshot[16][36] , \sa_snapshot[16][35] , \sa_snapshot[16][34] , 
	\sa_snapshot[16][33] , \sa_snapshot[16][32] , \sa_snapshot[16][31] , 
	\sa_snapshot[16][30] , \sa_snapshot[16][29] , \sa_snapshot[16][28] , 
	\sa_snapshot[16][27] , \sa_snapshot[16][26] , \sa_snapshot[16][25] , 
	\sa_snapshot[16][24] , \sa_snapshot[16][23] , \sa_snapshot[16][22] , 
	\sa_snapshot[16][21] , \sa_snapshot[16][20] , \sa_snapshot[16][19] , 
	\sa_snapshot[16][18] , \sa_snapshot[16][17] , \sa_snapshot[16][16] , 
	\sa_snapshot[16][15] , \sa_snapshot[16][14] , \sa_snapshot[16][13] , 
	\sa_snapshot[16][12] , \sa_snapshot[16][11] , \sa_snapshot[16][10] , 
	\sa_snapshot[16][9] , \sa_snapshot[16][8] , \sa_snapshot[16][7] , 
	\sa_snapshot[16][6] , \sa_snapshot[16][5] , \sa_snapshot[16][4] , 
	\sa_snapshot[16][3] , \sa_snapshot[16][2] , \sa_snapshot[16][1] , 
	\sa_snapshot[16][0] }, \num_16_._zy_simnet_tvar_86 [0:49]);
ixc_assign_50 \num_16_._zz_strnp_80 ( { \sa_count[16][49] , 
	\sa_count[16][48] , \sa_count[16][47] , \sa_count[16][46] , 
	\sa_count[16][45] , \sa_count[16][44] , \sa_count[16][43] , 
	\sa_count[16][42] , \sa_count[16][41] , \sa_count[16][40] , 
	\sa_count[16][39] , \sa_count[16][38] , \sa_count[16][37] , 
	\sa_count[16][36] , \sa_count[16][35] , \sa_count[16][34] , 
	\sa_count[16][33] , \sa_count[16][32] , \sa_count[16][31] , 
	\sa_count[16][30] , \sa_count[16][29] , \sa_count[16][28] , 
	\sa_count[16][27] , \sa_count[16][26] , \sa_count[16][25] , 
	\sa_count[16][24] , \sa_count[16][23] , \sa_count[16][22] , 
	\sa_count[16][21] , \sa_count[16][20] , \sa_count[16][19] , 
	\sa_count[16][18] , \sa_count[16][17] , \sa_count[16][16] , 
	\sa_count[16][15] , \sa_count[16][14] , \sa_count[16][13] , 
	\sa_count[16][12] , \sa_count[16][11] , \sa_count[16][10] , 
	\sa_count[16][9] , \sa_count[16][8] , \sa_count[16][7] , 
	\sa_count[16][6] , \sa_count[16][5] , \sa_count[16][4] , 
	\sa_count[16][3] , \sa_count[16][2] , \sa_count[16][1] , 
	\sa_count[16][0] }, \num_16_._zy_simnet_tvar_85 [0:49]);
ixc_assign_10 \num_17_._zz_strnp_87 ( \num_17_._zy_simnet_tvar_92 [0:9], { 
	n170, n169, n168, n167, n166, \sa_ctrl[17][4] , \sa_ctrl[17][3] , 
	\sa_ctrl[17][2] , \sa_ctrl[17][1] , \sa_ctrl[17][0] });
cr_sa_counter \num_17_.sa_counter_i ( .sa_count( 
	\num_17_._zy_simnet_tvar_90 [0:49]), .sa_snapshot( 
	\num_17_._zy_simnet_tvar_91 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_17_._zy_simnet_tvar_92 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_17_._zy_simnet_sa_clear_93_w$ ), 
	.sa_snap( \num_17_._zy_simnet_sa_snap_94_w$ ));
ixc_assign \num_17_._zz_strnp_89 ( \num_17_._zy_simnet_sa_snap_94_w$ , 
	sa_snap);
ixc_assign \num_17_._zz_strnp_88 ( \num_17_._zy_simnet_sa_clear_93_w$ , 
	sa_clear);
ixc_assign_50 \num_17_._zz_strnp_86 ( { \sa_snapshot[17][49] , 
	\sa_snapshot[17][48] , \sa_snapshot[17][47] , \sa_snapshot[17][46] , 
	\sa_snapshot[17][45] , \sa_snapshot[17][44] , \sa_snapshot[17][43] , 
	\sa_snapshot[17][42] , \sa_snapshot[17][41] , \sa_snapshot[17][40] , 
	\sa_snapshot[17][39] , \sa_snapshot[17][38] , \sa_snapshot[17][37] , 
	\sa_snapshot[17][36] , \sa_snapshot[17][35] , \sa_snapshot[17][34] , 
	\sa_snapshot[17][33] , \sa_snapshot[17][32] , \sa_snapshot[17][31] , 
	\sa_snapshot[17][30] , \sa_snapshot[17][29] , \sa_snapshot[17][28] , 
	\sa_snapshot[17][27] , \sa_snapshot[17][26] , \sa_snapshot[17][25] , 
	\sa_snapshot[17][24] , \sa_snapshot[17][23] , \sa_snapshot[17][22] , 
	\sa_snapshot[17][21] , \sa_snapshot[17][20] , \sa_snapshot[17][19] , 
	\sa_snapshot[17][18] , \sa_snapshot[17][17] , \sa_snapshot[17][16] , 
	\sa_snapshot[17][15] , \sa_snapshot[17][14] , \sa_snapshot[17][13] , 
	\sa_snapshot[17][12] , \sa_snapshot[17][11] , \sa_snapshot[17][10] , 
	\sa_snapshot[17][9] , \sa_snapshot[17][8] , \sa_snapshot[17][7] , 
	\sa_snapshot[17][6] , \sa_snapshot[17][5] , \sa_snapshot[17][4] , 
	\sa_snapshot[17][3] , \sa_snapshot[17][2] , \sa_snapshot[17][1] , 
	\sa_snapshot[17][0] }, \num_17_._zy_simnet_tvar_91 [0:49]);
ixc_assign_50 \num_17_._zz_strnp_85 ( { \sa_count[17][49] , 
	\sa_count[17][48] , \sa_count[17][47] , \sa_count[17][46] , 
	\sa_count[17][45] , \sa_count[17][44] , \sa_count[17][43] , 
	\sa_count[17][42] , \sa_count[17][41] , \sa_count[17][40] , 
	\sa_count[17][39] , \sa_count[17][38] , \sa_count[17][37] , 
	\sa_count[17][36] , \sa_count[17][35] , \sa_count[17][34] , 
	\sa_count[17][33] , \sa_count[17][32] , \sa_count[17][31] , 
	\sa_count[17][30] , \sa_count[17][29] , \sa_count[17][28] , 
	\sa_count[17][27] , \sa_count[17][26] , \sa_count[17][25] , 
	\sa_count[17][24] , \sa_count[17][23] , \sa_count[17][22] , 
	\sa_count[17][21] , \sa_count[17][20] , \sa_count[17][19] , 
	\sa_count[17][18] , \sa_count[17][17] , \sa_count[17][16] , 
	\sa_count[17][15] , \sa_count[17][14] , \sa_count[17][13] , 
	\sa_count[17][12] , \sa_count[17][11] , \sa_count[17][10] , 
	\sa_count[17][9] , \sa_count[17][8] , \sa_count[17][7] , 
	\sa_count[17][6] , \sa_count[17][5] , \sa_count[17][4] , 
	\sa_count[17][3] , \sa_count[17][2] , \sa_count[17][1] , 
	\sa_count[17][0] }, \num_17_._zy_simnet_tvar_90 [0:49]);
ixc_assign_10 \num_18_._zz_strnp_92 ( \num_18_._zy_simnet_tvar_97 [0:9], { 
	n175, n174, n173, n172, n171, \sa_ctrl[18][4] , \sa_ctrl[18][3] , 
	\sa_ctrl[18][2] , \sa_ctrl[18][1] , \sa_ctrl[18][0] });
cr_sa_counter \num_18_.sa_counter_i ( .sa_count( 
	\num_18_._zy_simnet_tvar_95 [0:49]), .sa_snapshot( 
	\num_18_._zy_simnet_tvar_96 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_18_._zy_simnet_tvar_97 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( \num_18_._zy_simnet_sa_clear_98_w$ ), 
	.sa_snap( \num_18_._zy_simnet_sa_snap_99_w$ ));
ixc_assign \num_18_._zz_strnp_94 ( \num_18_._zy_simnet_sa_snap_99_w$ , 
	sa_snap);
ixc_assign \num_18_._zz_strnp_93 ( \num_18_._zy_simnet_sa_clear_98_w$ , 
	sa_clear);
ixc_assign_50 \num_18_._zz_strnp_91 ( { \sa_snapshot[18][49] , 
	\sa_snapshot[18][48] , \sa_snapshot[18][47] , \sa_snapshot[18][46] , 
	\sa_snapshot[18][45] , \sa_snapshot[18][44] , \sa_snapshot[18][43] , 
	\sa_snapshot[18][42] , \sa_snapshot[18][41] , \sa_snapshot[18][40] , 
	\sa_snapshot[18][39] , \sa_snapshot[18][38] , \sa_snapshot[18][37] , 
	\sa_snapshot[18][36] , \sa_snapshot[18][35] , \sa_snapshot[18][34] , 
	\sa_snapshot[18][33] , \sa_snapshot[18][32] , \sa_snapshot[18][31] , 
	\sa_snapshot[18][30] , \sa_snapshot[18][29] , \sa_snapshot[18][28] , 
	\sa_snapshot[18][27] , \sa_snapshot[18][26] , \sa_snapshot[18][25] , 
	\sa_snapshot[18][24] , \sa_snapshot[18][23] , \sa_snapshot[18][22] , 
	\sa_snapshot[18][21] , \sa_snapshot[18][20] , \sa_snapshot[18][19] , 
	\sa_snapshot[18][18] , \sa_snapshot[18][17] , \sa_snapshot[18][16] , 
	\sa_snapshot[18][15] , \sa_snapshot[18][14] , \sa_snapshot[18][13] , 
	\sa_snapshot[18][12] , \sa_snapshot[18][11] , \sa_snapshot[18][10] , 
	\sa_snapshot[18][9] , \sa_snapshot[18][8] , \sa_snapshot[18][7] , 
	\sa_snapshot[18][6] , \sa_snapshot[18][5] , \sa_snapshot[18][4] , 
	\sa_snapshot[18][3] , \sa_snapshot[18][2] , \sa_snapshot[18][1] , 
	\sa_snapshot[18][0] }, \num_18_._zy_simnet_tvar_96 [0:49]);
ixc_assign_50 \num_18_._zz_strnp_90 ( { \sa_count[18][49] , 
	\sa_count[18][48] , \sa_count[18][47] , \sa_count[18][46] , 
	\sa_count[18][45] , \sa_count[18][44] , \sa_count[18][43] , 
	\sa_count[18][42] , \sa_count[18][41] , \sa_count[18][40] , 
	\sa_count[18][39] , \sa_count[18][38] , \sa_count[18][37] , 
	\sa_count[18][36] , \sa_count[18][35] , \sa_count[18][34] , 
	\sa_count[18][33] , \sa_count[18][32] , \sa_count[18][31] , 
	\sa_count[18][30] , \sa_count[18][29] , \sa_count[18][28] , 
	\sa_count[18][27] , \sa_count[18][26] , \sa_count[18][25] , 
	\sa_count[18][24] , \sa_count[18][23] , \sa_count[18][22] , 
	\sa_count[18][21] , \sa_count[18][20] , \sa_count[18][19] , 
	\sa_count[18][18] , \sa_count[18][17] , \sa_count[18][16] , 
	\sa_count[18][15] , \sa_count[18][14] , \sa_count[18][13] , 
	\sa_count[18][12] , \sa_count[18][11] , \sa_count[18][10] , 
	\sa_count[18][9] , \sa_count[18][8] , \sa_count[18][7] , 
	\sa_count[18][6] , \sa_count[18][5] , \sa_count[18][4] , 
	\sa_count[18][3] , \sa_count[18][2] , \sa_count[18][1] , 
	\sa_count[18][0] }, \num_18_._zy_simnet_tvar_95 [0:49]);
ixc_assign_10 \num_19_._zz_strnp_97 ( \num_19_._zy_simnet_tvar_102 [0:9], { 
	n180, n179, n178, n177, n176, \sa_ctrl[19][4] , \sa_ctrl[19][3] , 
	\sa_ctrl[19][2] , \sa_ctrl[19][1] , \sa_ctrl[19][0] });
cr_sa_counter \num_19_.sa_counter_i ( .sa_count( 
	\num_19_._zy_simnet_tvar_100 [0:49]), .sa_snapshot( 
	\num_19_._zy_simnet_tvar_101 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_19_._zy_simnet_tvar_102 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_19_._zy_simnet_sa_clear_103_w$ ), .sa_snap( 
	\num_19_._zy_simnet_sa_snap_104_w$ ));
ixc_assign \num_19_._zz_strnp_99 ( \num_19_._zy_simnet_sa_snap_104_w$ , 
	sa_snap);
ixc_assign \num_19_._zz_strnp_98 ( \num_19_._zy_simnet_sa_clear_103_w$ , 
	sa_clear);
ixc_assign_50 \num_19_._zz_strnp_96 ( { \sa_snapshot[19][49] , 
	\sa_snapshot[19][48] , \sa_snapshot[19][47] , \sa_snapshot[19][46] , 
	\sa_snapshot[19][45] , \sa_snapshot[19][44] , \sa_snapshot[19][43] , 
	\sa_snapshot[19][42] , \sa_snapshot[19][41] , \sa_snapshot[19][40] , 
	\sa_snapshot[19][39] , \sa_snapshot[19][38] , \sa_snapshot[19][37] , 
	\sa_snapshot[19][36] , \sa_snapshot[19][35] , \sa_snapshot[19][34] , 
	\sa_snapshot[19][33] , \sa_snapshot[19][32] , \sa_snapshot[19][31] , 
	\sa_snapshot[19][30] , \sa_snapshot[19][29] , \sa_snapshot[19][28] , 
	\sa_snapshot[19][27] , \sa_snapshot[19][26] , \sa_snapshot[19][25] , 
	\sa_snapshot[19][24] , \sa_snapshot[19][23] , \sa_snapshot[19][22] , 
	\sa_snapshot[19][21] , \sa_snapshot[19][20] , \sa_snapshot[19][19] , 
	\sa_snapshot[19][18] , \sa_snapshot[19][17] , \sa_snapshot[19][16] , 
	\sa_snapshot[19][15] , \sa_snapshot[19][14] , \sa_snapshot[19][13] , 
	\sa_snapshot[19][12] , \sa_snapshot[19][11] , \sa_snapshot[19][10] , 
	\sa_snapshot[19][9] , \sa_snapshot[19][8] , \sa_snapshot[19][7] , 
	\sa_snapshot[19][6] , \sa_snapshot[19][5] , \sa_snapshot[19][4] , 
	\sa_snapshot[19][3] , \sa_snapshot[19][2] , \sa_snapshot[19][1] , 
	\sa_snapshot[19][0] }, \num_19_._zy_simnet_tvar_101 [0:49]);
ixc_assign_50 \num_19_._zz_strnp_95 ( { \sa_count[19][49] , 
	\sa_count[19][48] , \sa_count[19][47] , \sa_count[19][46] , 
	\sa_count[19][45] , \sa_count[19][44] , \sa_count[19][43] , 
	\sa_count[19][42] , \sa_count[19][41] , \sa_count[19][40] , 
	\sa_count[19][39] , \sa_count[19][38] , \sa_count[19][37] , 
	\sa_count[19][36] , \sa_count[19][35] , \sa_count[19][34] , 
	\sa_count[19][33] , \sa_count[19][32] , \sa_count[19][31] , 
	\sa_count[19][30] , \sa_count[19][29] , \sa_count[19][28] , 
	\sa_count[19][27] , \sa_count[19][26] , \sa_count[19][25] , 
	\sa_count[19][24] , \sa_count[19][23] , \sa_count[19][22] , 
	\sa_count[19][21] , \sa_count[19][20] , \sa_count[19][19] , 
	\sa_count[19][18] , \sa_count[19][17] , \sa_count[19][16] , 
	\sa_count[19][15] , \sa_count[19][14] , \sa_count[19][13] , 
	\sa_count[19][12] , \sa_count[19][11] , \sa_count[19][10] , 
	\sa_count[19][9] , \sa_count[19][8] , \sa_count[19][7] , 
	\sa_count[19][6] , \sa_count[19][5] , \sa_count[19][4] , 
	\sa_count[19][3] , \sa_count[19][2] , \sa_count[19][1] , 
	\sa_count[19][0] }, \num_19_._zy_simnet_tvar_100 [0:49]);
ixc_assign_10 \num_20_._zz_strnp_102 ( \num_20_._zy_simnet_tvar_107 [0:9], { 
	n185, n184, n183, n182, n181, \sa_ctrl[20][4] , \sa_ctrl[20][3] , 
	\sa_ctrl[20][2] , \sa_ctrl[20][1] , \sa_ctrl[20][0] });
cr_sa_counter \num_20_.sa_counter_i ( .sa_count( 
	\num_20_._zy_simnet_tvar_105 [0:49]), .sa_snapshot( 
	\num_20_._zy_simnet_tvar_106 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_20_._zy_simnet_tvar_107 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_20_._zy_simnet_sa_clear_108_w$ ), .sa_snap( 
	\num_20_._zy_simnet_sa_snap_109_w$ ));
ixc_assign \num_20_._zz_strnp_104 ( \num_20_._zy_simnet_sa_snap_109_w$ , 
	sa_snap);
ixc_assign \num_20_._zz_strnp_103 ( \num_20_._zy_simnet_sa_clear_108_w$ , 
	sa_clear);
ixc_assign_50 \num_20_._zz_strnp_101 ( { \sa_snapshot[20][49] , 
	\sa_snapshot[20][48] , \sa_snapshot[20][47] , \sa_snapshot[20][46] , 
	\sa_snapshot[20][45] , \sa_snapshot[20][44] , \sa_snapshot[20][43] , 
	\sa_snapshot[20][42] , \sa_snapshot[20][41] , \sa_snapshot[20][40] , 
	\sa_snapshot[20][39] , \sa_snapshot[20][38] , \sa_snapshot[20][37] , 
	\sa_snapshot[20][36] , \sa_snapshot[20][35] , \sa_snapshot[20][34] , 
	\sa_snapshot[20][33] , \sa_snapshot[20][32] , \sa_snapshot[20][31] , 
	\sa_snapshot[20][30] , \sa_snapshot[20][29] , \sa_snapshot[20][28] , 
	\sa_snapshot[20][27] , \sa_snapshot[20][26] , \sa_snapshot[20][25] , 
	\sa_snapshot[20][24] , \sa_snapshot[20][23] , \sa_snapshot[20][22] , 
	\sa_snapshot[20][21] , \sa_snapshot[20][20] , \sa_snapshot[20][19] , 
	\sa_snapshot[20][18] , \sa_snapshot[20][17] , \sa_snapshot[20][16] , 
	\sa_snapshot[20][15] , \sa_snapshot[20][14] , \sa_snapshot[20][13] , 
	\sa_snapshot[20][12] , \sa_snapshot[20][11] , \sa_snapshot[20][10] , 
	\sa_snapshot[20][9] , \sa_snapshot[20][8] , \sa_snapshot[20][7] , 
	\sa_snapshot[20][6] , \sa_snapshot[20][5] , \sa_snapshot[20][4] , 
	\sa_snapshot[20][3] , \sa_snapshot[20][2] , \sa_snapshot[20][1] , 
	\sa_snapshot[20][0] }, \num_20_._zy_simnet_tvar_106 [0:49]);
ixc_assign_50 \num_20_._zz_strnp_100 ( { \sa_count[20][49] , 
	\sa_count[20][48] , \sa_count[20][47] , \sa_count[20][46] , 
	\sa_count[20][45] , \sa_count[20][44] , \sa_count[20][43] , 
	\sa_count[20][42] , \sa_count[20][41] , \sa_count[20][40] , 
	\sa_count[20][39] , \sa_count[20][38] , \sa_count[20][37] , 
	\sa_count[20][36] , \sa_count[20][35] , \sa_count[20][34] , 
	\sa_count[20][33] , \sa_count[20][32] , \sa_count[20][31] , 
	\sa_count[20][30] , \sa_count[20][29] , \sa_count[20][28] , 
	\sa_count[20][27] , \sa_count[20][26] , \sa_count[20][25] , 
	\sa_count[20][24] , \sa_count[20][23] , \sa_count[20][22] , 
	\sa_count[20][21] , \sa_count[20][20] , \sa_count[20][19] , 
	\sa_count[20][18] , \sa_count[20][17] , \sa_count[20][16] , 
	\sa_count[20][15] , \sa_count[20][14] , \sa_count[20][13] , 
	\sa_count[20][12] , \sa_count[20][11] , \sa_count[20][10] , 
	\sa_count[20][9] , \sa_count[20][8] , \sa_count[20][7] , 
	\sa_count[20][6] , \sa_count[20][5] , \sa_count[20][4] , 
	\sa_count[20][3] , \sa_count[20][2] , \sa_count[20][1] , 
	\sa_count[20][0] }, \num_20_._zy_simnet_tvar_105 [0:49]);
ixc_assign_10 \num_21_._zz_strnp_107 ( \num_21_._zy_simnet_tvar_112 [0:9], { 
	n190, n189, n188, n187, n186, \sa_ctrl[21][4] , \sa_ctrl[21][3] , 
	\sa_ctrl[21][2] , \sa_ctrl[21][1] , \sa_ctrl[21][0] });
cr_sa_counter \num_21_.sa_counter_i ( .sa_count( 
	\num_21_._zy_simnet_tvar_110 [0:49]), .sa_snapshot( 
	\num_21_._zy_simnet_tvar_111 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_21_._zy_simnet_tvar_112 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_21_._zy_simnet_sa_clear_113_w$ ), .sa_snap( 
	\num_21_._zy_simnet_sa_snap_114_w$ ));
ixc_assign \num_21_._zz_strnp_109 ( \num_21_._zy_simnet_sa_snap_114_w$ , 
	sa_snap);
ixc_assign \num_21_._zz_strnp_108 ( \num_21_._zy_simnet_sa_clear_113_w$ , 
	sa_clear);
ixc_assign_50 \num_21_._zz_strnp_106 ( { \sa_snapshot[21][49] , 
	\sa_snapshot[21][48] , \sa_snapshot[21][47] , \sa_snapshot[21][46] , 
	\sa_snapshot[21][45] , \sa_snapshot[21][44] , \sa_snapshot[21][43] , 
	\sa_snapshot[21][42] , \sa_snapshot[21][41] , \sa_snapshot[21][40] , 
	\sa_snapshot[21][39] , \sa_snapshot[21][38] , \sa_snapshot[21][37] , 
	\sa_snapshot[21][36] , \sa_snapshot[21][35] , \sa_snapshot[21][34] , 
	\sa_snapshot[21][33] , \sa_snapshot[21][32] , \sa_snapshot[21][31] , 
	\sa_snapshot[21][30] , \sa_snapshot[21][29] , \sa_snapshot[21][28] , 
	\sa_snapshot[21][27] , \sa_snapshot[21][26] , \sa_snapshot[21][25] , 
	\sa_snapshot[21][24] , \sa_snapshot[21][23] , \sa_snapshot[21][22] , 
	\sa_snapshot[21][21] , \sa_snapshot[21][20] , \sa_snapshot[21][19] , 
	\sa_snapshot[21][18] , \sa_snapshot[21][17] , \sa_snapshot[21][16] , 
	\sa_snapshot[21][15] , \sa_snapshot[21][14] , \sa_snapshot[21][13] , 
	\sa_snapshot[21][12] , \sa_snapshot[21][11] , \sa_snapshot[21][10] , 
	\sa_snapshot[21][9] , \sa_snapshot[21][8] , \sa_snapshot[21][7] , 
	\sa_snapshot[21][6] , \sa_snapshot[21][5] , \sa_snapshot[21][4] , 
	\sa_snapshot[21][3] , \sa_snapshot[21][2] , \sa_snapshot[21][1] , 
	\sa_snapshot[21][0] }, \num_21_._zy_simnet_tvar_111 [0:49]);
ixc_assign_50 \num_21_._zz_strnp_105 ( { \sa_count[21][49] , 
	\sa_count[21][48] , \sa_count[21][47] , \sa_count[21][46] , 
	\sa_count[21][45] , \sa_count[21][44] , \sa_count[21][43] , 
	\sa_count[21][42] , \sa_count[21][41] , \sa_count[21][40] , 
	\sa_count[21][39] , \sa_count[21][38] , \sa_count[21][37] , 
	\sa_count[21][36] , \sa_count[21][35] , \sa_count[21][34] , 
	\sa_count[21][33] , \sa_count[21][32] , \sa_count[21][31] , 
	\sa_count[21][30] , \sa_count[21][29] , \sa_count[21][28] , 
	\sa_count[21][27] , \sa_count[21][26] , \sa_count[21][25] , 
	\sa_count[21][24] , \sa_count[21][23] , \sa_count[21][22] , 
	\sa_count[21][21] , \sa_count[21][20] , \sa_count[21][19] , 
	\sa_count[21][18] , \sa_count[21][17] , \sa_count[21][16] , 
	\sa_count[21][15] , \sa_count[21][14] , \sa_count[21][13] , 
	\sa_count[21][12] , \sa_count[21][11] , \sa_count[21][10] , 
	\sa_count[21][9] , \sa_count[21][8] , \sa_count[21][7] , 
	\sa_count[21][6] , \sa_count[21][5] , \sa_count[21][4] , 
	\sa_count[21][3] , \sa_count[21][2] , \sa_count[21][1] , 
	\sa_count[21][0] }, \num_21_._zy_simnet_tvar_110 [0:49]);
ixc_assign_10 \num_22_._zz_strnp_112 ( \num_22_._zy_simnet_tvar_117 [0:9], { 
	n195, n194, n193, n192, n191, \sa_ctrl[22][4] , \sa_ctrl[22][3] , 
	\sa_ctrl[22][2] , \sa_ctrl[22][1] , \sa_ctrl[22][0] });
cr_sa_counter \num_22_.sa_counter_i ( .sa_count( 
	\num_22_._zy_simnet_tvar_115 [0:49]), .sa_snapshot( 
	\num_22_._zy_simnet_tvar_116 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_22_._zy_simnet_tvar_117 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_22_._zy_simnet_sa_clear_118_w$ ), .sa_snap( 
	\num_22_._zy_simnet_sa_snap_119_w$ ));
ixc_assign \num_22_._zz_strnp_114 ( \num_22_._zy_simnet_sa_snap_119_w$ , 
	sa_snap);
ixc_assign \num_22_._zz_strnp_113 ( \num_22_._zy_simnet_sa_clear_118_w$ , 
	sa_clear);
ixc_assign_50 \num_22_._zz_strnp_111 ( { \sa_snapshot[22][49] , 
	\sa_snapshot[22][48] , \sa_snapshot[22][47] , \sa_snapshot[22][46] , 
	\sa_snapshot[22][45] , \sa_snapshot[22][44] , \sa_snapshot[22][43] , 
	\sa_snapshot[22][42] , \sa_snapshot[22][41] , \sa_snapshot[22][40] , 
	\sa_snapshot[22][39] , \sa_snapshot[22][38] , \sa_snapshot[22][37] , 
	\sa_snapshot[22][36] , \sa_snapshot[22][35] , \sa_snapshot[22][34] , 
	\sa_snapshot[22][33] , \sa_snapshot[22][32] , \sa_snapshot[22][31] , 
	\sa_snapshot[22][30] , \sa_snapshot[22][29] , \sa_snapshot[22][28] , 
	\sa_snapshot[22][27] , \sa_snapshot[22][26] , \sa_snapshot[22][25] , 
	\sa_snapshot[22][24] , \sa_snapshot[22][23] , \sa_snapshot[22][22] , 
	\sa_snapshot[22][21] , \sa_snapshot[22][20] , \sa_snapshot[22][19] , 
	\sa_snapshot[22][18] , \sa_snapshot[22][17] , \sa_snapshot[22][16] , 
	\sa_snapshot[22][15] , \sa_snapshot[22][14] , \sa_snapshot[22][13] , 
	\sa_snapshot[22][12] , \sa_snapshot[22][11] , \sa_snapshot[22][10] , 
	\sa_snapshot[22][9] , \sa_snapshot[22][8] , \sa_snapshot[22][7] , 
	\sa_snapshot[22][6] , \sa_snapshot[22][5] , \sa_snapshot[22][4] , 
	\sa_snapshot[22][3] , \sa_snapshot[22][2] , \sa_snapshot[22][1] , 
	\sa_snapshot[22][0] }, \num_22_._zy_simnet_tvar_116 [0:49]);
ixc_assign_50 \num_22_._zz_strnp_110 ( { \sa_count[22][49] , 
	\sa_count[22][48] , \sa_count[22][47] , \sa_count[22][46] , 
	\sa_count[22][45] , \sa_count[22][44] , \sa_count[22][43] , 
	\sa_count[22][42] , \sa_count[22][41] , \sa_count[22][40] , 
	\sa_count[22][39] , \sa_count[22][38] , \sa_count[22][37] , 
	\sa_count[22][36] , \sa_count[22][35] , \sa_count[22][34] , 
	\sa_count[22][33] , \sa_count[22][32] , \sa_count[22][31] , 
	\sa_count[22][30] , \sa_count[22][29] , \sa_count[22][28] , 
	\sa_count[22][27] , \sa_count[22][26] , \sa_count[22][25] , 
	\sa_count[22][24] , \sa_count[22][23] , \sa_count[22][22] , 
	\sa_count[22][21] , \sa_count[22][20] , \sa_count[22][19] , 
	\sa_count[22][18] , \sa_count[22][17] , \sa_count[22][16] , 
	\sa_count[22][15] , \sa_count[22][14] , \sa_count[22][13] , 
	\sa_count[22][12] , \sa_count[22][11] , \sa_count[22][10] , 
	\sa_count[22][9] , \sa_count[22][8] , \sa_count[22][7] , 
	\sa_count[22][6] , \sa_count[22][5] , \sa_count[22][4] , 
	\sa_count[22][3] , \sa_count[22][2] , \sa_count[22][1] , 
	\sa_count[22][0] }, \num_22_._zy_simnet_tvar_115 [0:49]);
ixc_assign_10 \num_23_._zz_strnp_117 ( \num_23_._zy_simnet_tvar_122 [0:9], { 
	n200, n199, n198, n197, n196, \sa_ctrl[23][4] , \sa_ctrl[23][3] , 
	\sa_ctrl[23][2] , \sa_ctrl[23][1] , \sa_ctrl[23][0] });
cr_sa_counter \num_23_.sa_counter_i ( .sa_count( 
	\num_23_._zy_simnet_tvar_120 [0:49]), .sa_snapshot( 
	\num_23_._zy_simnet_tvar_121 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_23_._zy_simnet_tvar_122 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_23_._zy_simnet_sa_clear_123_w$ ), .sa_snap( 
	\num_23_._zy_simnet_sa_snap_124_w$ ));
ixc_assign \num_23_._zz_strnp_119 ( \num_23_._zy_simnet_sa_snap_124_w$ , 
	sa_snap);
ixc_assign \num_23_._zz_strnp_118 ( \num_23_._zy_simnet_sa_clear_123_w$ , 
	sa_clear);
ixc_assign_50 \num_23_._zz_strnp_116 ( { \sa_snapshot[23][49] , 
	\sa_snapshot[23][48] , \sa_snapshot[23][47] , \sa_snapshot[23][46] , 
	\sa_snapshot[23][45] , \sa_snapshot[23][44] , \sa_snapshot[23][43] , 
	\sa_snapshot[23][42] , \sa_snapshot[23][41] , \sa_snapshot[23][40] , 
	\sa_snapshot[23][39] , \sa_snapshot[23][38] , \sa_snapshot[23][37] , 
	\sa_snapshot[23][36] , \sa_snapshot[23][35] , \sa_snapshot[23][34] , 
	\sa_snapshot[23][33] , \sa_snapshot[23][32] , \sa_snapshot[23][31] , 
	\sa_snapshot[23][30] , \sa_snapshot[23][29] , \sa_snapshot[23][28] , 
	\sa_snapshot[23][27] , \sa_snapshot[23][26] , \sa_snapshot[23][25] , 
	\sa_snapshot[23][24] , \sa_snapshot[23][23] , \sa_snapshot[23][22] , 
	\sa_snapshot[23][21] , \sa_snapshot[23][20] , \sa_snapshot[23][19] , 
	\sa_snapshot[23][18] , \sa_snapshot[23][17] , \sa_snapshot[23][16] , 
	\sa_snapshot[23][15] , \sa_snapshot[23][14] , \sa_snapshot[23][13] , 
	\sa_snapshot[23][12] , \sa_snapshot[23][11] , \sa_snapshot[23][10] , 
	\sa_snapshot[23][9] , \sa_snapshot[23][8] , \sa_snapshot[23][7] , 
	\sa_snapshot[23][6] , \sa_snapshot[23][5] , \sa_snapshot[23][4] , 
	\sa_snapshot[23][3] , \sa_snapshot[23][2] , \sa_snapshot[23][1] , 
	\sa_snapshot[23][0] }, \num_23_._zy_simnet_tvar_121 [0:49]);
ixc_assign_50 \num_23_._zz_strnp_115 ( { \sa_count[23][49] , 
	\sa_count[23][48] , \sa_count[23][47] , \sa_count[23][46] , 
	\sa_count[23][45] , \sa_count[23][44] , \sa_count[23][43] , 
	\sa_count[23][42] , \sa_count[23][41] , \sa_count[23][40] , 
	\sa_count[23][39] , \sa_count[23][38] , \sa_count[23][37] , 
	\sa_count[23][36] , \sa_count[23][35] , \sa_count[23][34] , 
	\sa_count[23][33] , \sa_count[23][32] , \sa_count[23][31] , 
	\sa_count[23][30] , \sa_count[23][29] , \sa_count[23][28] , 
	\sa_count[23][27] , \sa_count[23][26] , \sa_count[23][25] , 
	\sa_count[23][24] , \sa_count[23][23] , \sa_count[23][22] , 
	\sa_count[23][21] , \sa_count[23][20] , \sa_count[23][19] , 
	\sa_count[23][18] , \sa_count[23][17] , \sa_count[23][16] , 
	\sa_count[23][15] , \sa_count[23][14] , \sa_count[23][13] , 
	\sa_count[23][12] , \sa_count[23][11] , \sa_count[23][10] , 
	\sa_count[23][9] , \sa_count[23][8] , \sa_count[23][7] , 
	\sa_count[23][6] , \sa_count[23][5] , \sa_count[23][4] , 
	\sa_count[23][3] , \sa_count[23][2] , \sa_count[23][1] , 
	\sa_count[23][0] }, \num_23_._zy_simnet_tvar_120 [0:49]);
ixc_assign_10 \num_24_._zz_strnp_122 ( \num_24_._zy_simnet_tvar_127 [0:9], { 
	n205, n204, n203, n202, n201, \sa_ctrl[24][4] , \sa_ctrl[24][3] , 
	\sa_ctrl[24][2] , \sa_ctrl[24][1] , \sa_ctrl[24][0] });
cr_sa_counter \num_24_.sa_counter_i ( .sa_count( 
	\num_24_._zy_simnet_tvar_125 [0:49]), .sa_snapshot( 
	\num_24_._zy_simnet_tvar_126 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_24_._zy_simnet_tvar_127 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_24_._zy_simnet_sa_clear_128_w$ ), .sa_snap( 
	\num_24_._zy_simnet_sa_snap_129_w$ ));
ixc_assign \num_24_._zz_strnp_124 ( \num_24_._zy_simnet_sa_snap_129_w$ , 
	sa_snap);
ixc_assign \num_24_._zz_strnp_123 ( \num_24_._zy_simnet_sa_clear_128_w$ , 
	sa_clear);
ixc_assign_50 \num_24_._zz_strnp_121 ( { \sa_snapshot[24][49] , 
	\sa_snapshot[24][48] , \sa_snapshot[24][47] , \sa_snapshot[24][46] , 
	\sa_snapshot[24][45] , \sa_snapshot[24][44] , \sa_snapshot[24][43] , 
	\sa_snapshot[24][42] , \sa_snapshot[24][41] , \sa_snapshot[24][40] , 
	\sa_snapshot[24][39] , \sa_snapshot[24][38] , \sa_snapshot[24][37] , 
	\sa_snapshot[24][36] , \sa_snapshot[24][35] , \sa_snapshot[24][34] , 
	\sa_snapshot[24][33] , \sa_snapshot[24][32] , \sa_snapshot[24][31] , 
	\sa_snapshot[24][30] , \sa_snapshot[24][29] , \sa_snapshot[24][28] , 
	\sa_snapshot[24][27] , \sa_snapshot[24][26] , \sa_snapshot[24][25] , 
	\sa_snapshot[24][24] , \sa_snapshot[24][23] , \sa_snapshot[24][22] , 
	\sa_snapshot[24][21] , \sa_snapshot[24][20] , \sa_snapshot[24][19] , 
	\sa_snapshot[24][18] , \sa_snapshot[24][17] , \sa_snapshot[24][16] , 
	\sa_snapshot[24][15] , \sa_snapshot[24][14] , \sa_snapshot[24][13] , 
	\sa_snapshot[24][12] , \sa_snapshot[24][11] , \sa_snapshot[24][10] , 
	\sa_snapshot[24][9] , \sa_snapshot[24][8] , \sa_snapshot[24][7] , 
	\sa_snapshot[24][6] , \sa_snapshot[24][5] , \sa_snapshot[24][4] , 
	\sa_snapshot[24][3] , \sa_snapshot[24][2] , \sa_snapshot[24][1] , 
	\sa_snapshot[24][0] }, \num_24_._zy_simnet_tvar_126 [0:49]);
ixc_assign_50 \num_24_._zz_strnp_120 ( { \sa_count[24][49] , 
	\sa_count[24][48] , \sa_count[24][47] , \sa_count[24][46] , 
	\sa_count[24][45] , \sa_count[24][44] , \sa_count[24][43] , 
	\sa_count[24][42] , \sa_count[24][41] , \sa_count[24][40] , 
	\sa_count[24][39] , \sa_count[24][38] , \sa_count[24][37] , 
	\sa_count[24][36] , \sa_count[24][35] , \sa_count[24][34] , 
	\sa_count[24][33] , \sa_count[24][32] , \sa_count[24][31] , 
	\sa_count[24][30] , \sa_count[24][29] , \sa_count[24][28] , 
	\sa_count[24][27] , \sa_count[24][26] , \sa_count[24][25] , 
	\sa_count[24][24] , \sa_count[24][23] , \sa_count[24][22] , 
	\sa_count[24][21] , \sa_count[24][20] , \sa_count[24][19] , 
	\sa_count[24][18] , \sa_count[24][17] , \sa_count[24][16] , 
	\sa_count[24][15] , \sa_count[24][14] , \sa_count[24][13] , 
	\sa_count[24][12] , \sa_count[24][11] , \sa_count[24][10] , 
	\sa_count[24][9] , \sa_count[24][8] , \sa_count[24][7] , 
	\sa_count[24][6] , \sa_count[24][5] , \sa_count[24][4] , 
	\sa_count[24][3] , \sa_count[24][2] , \sa_count[24][1] , 
	\sa_count[24][0] }, \num_24_._zy_simnet_tvar_125 [0:49]);
ixc_assign_10 \num_25_._zz_strnp_127 ( \num_25_._zy_simnet_tvar_132 [0:9], { 
	n210, n209, n208, n207, n206, \sa_ctrl[25][4] , \sa_ctrl[25][3] , 
	\sa_ctrl[25][2] , \sa_ctrl[25][1] , \sa_ctrl[25][0] });
cr_sa_counter \num_25_.sa_counter_i ( .sa_count( 
	\num_25_._zy_simnet_tvar_130 [0:49]), .sa_snapshot( 
	\num_25_._zy_simnet_tvar_131 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_25_._zy_simnet_tvar_132 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_25_._zy_simnet_sa_clear_133_w$ ), .sa_snap( 
	\num_25_._zy_simnet_sa_snap_134_w$ ));
ixc_assign \num_25_._zz_strnp_129 ( \num_25_._zy_simnet_sa_snap_134_w$ , 
	sa_snap);
ixc_assign \num_25_._zz_strnp_128 ( \num_25_._zy_simnet_sa_clear_133_w$ , 
	sa_clear);
ixc_assign_50 \num_25_._zz_strnp_126 ( { \sa_snapshot[25][49] , 
	\sa_snapshot[25][48] , \sa_snapshot[25][47] , \sa_snapshot[25][46] , 
	\sa_snapshot[25][45] , \sa_snapshot[25][44] , \sa_snapshot[25][43] , 
	\sa_snapshot[25][42] , \sa_snapshot[25][41] , \sa_snapshot[25][40] , 
	\sa_snapshot[25][39] , \sa_snapshot[25][38] , \sa_snapshot[25][37] , 
	\sa_snapshot[25][36] , \sa_snapshot[25][35] , \sa_snapshot[25][34] , 
	\sa_snapshot[25][33] , \sa_snapshot[25][32] , \sa_snapshot[25][31] , 
	\sa_snapshot[25][30] , \sa_snapshot[25][29] , \sa_snapshot[25][28] , 
	\sa_snapshot[25][27] , \sa_snapshot[25][26] , \sa_snapshot[25][25] , 
	\sa_snapshot[25][24] , \sa_snapshot[25][23] , \sa_snapshot[25][22] , 
	\sa_snapshot[25][21] , \sa_snapshot[25][20] , \sa_snapshot[25][19] , 
	\sa_snapshot[25][18] , \sa_snapshot[25][17] , \sa_snapshot[25][16] , 
	\sa_snapshot[25][15] , \sa_snapshot[25][14] , \sa_snapshot[25][13] , 
	\sa_snapshot[25][12] , \sa_snapshot[25][11] , \sa_snapshot[25][10] , 
	\sa_snapshot[25][9] , \sa_snapshot[25][8] , \sa_snapshot[25][7] , 
	\sa_snapshot[25][6] , \sa_snapshot[25][5] , \sa_snapshot[25][4] , 
	\sa_snapshot[25][3] , \sa_snapshot[25][2] , \sa_snapshot[25][1] , 
	\sa_snapshot[25][0] }, \num_25_._zy_simnet_tvar_131 [0:49]);
ixc_assign_50 \num_25_._zz_strnp_125 ( { \sa_count[25][49] , 
	\sa_count[25][48] , \sa_count[25][47] , \sa_count[25][46] , 
	\sa_count[25][45] , \sa_count[25][44] , \sa_count[25][43] , 
	\sa_count[25][42] , \sa_count[25][41] , \sa_count[25][40] , 
	\sa_count[25][39] , \sa_count[25][38] , \sa_count[25][37] , 
	\sa_count[25][36] , \sa_count[25][35] , \sa_count[25][34] , 
	\sa_count[25][33] , \sa_count[25][32] , \sa_count[25][31] , 
	\sa_count[25][30] , \sa_count[25][29] , \sa_count[25][28] , 
	\sa_count[25][27] , \sa_count[25][26] , \sa_count[25][25] , 
	\sa_count[25][24] , \sa_count[25][23] , \sa_count[25][22] , 
	\sa_count[25][21] , \sa_count[25][20] , \sa_count[25][19] , 
	\sa_count[25][18] , \sa_count[25][17] , \sa_count[25][16] , 
	\sa_count[25][15] , \sa_count[25][14] , \sa_count[25][13] , 
	\sa_count[25][12] , \sa_count[25][11] , \sa_count[25][10] , 
	\sa_count[25][9] , \sa_count[25][8] , \sa_count[25][7] , 
	\sa_count[25][6] , \sa_count[25][5] , \sa_count[25][4] , 
	\sa_count[25][3] , \sa_count[25][2] , \sa_count[25][1] , 
	\sa_count[25][0] }, \num_25_._zy_simnet_tvar_130 [0:49]);
ixc_assign_10 \num_26_._zz_strnp_132 ( \num_26_._zy_simnet_tvar_137 [0:9], { 
	n215, n214, n213, n212, n211, \sa_ctrl[26][4] , \sa_ctrl[26][3] , 
	\sa_ctrl[26][2] , \sa_ctrl[26][1] , \sa_ctrl[26][0] });
cr_sa_counter \num_26_.sa_counter_i ( .sa_count( 
	\num_26_._zy_simnet_tvar_135 [0:49]), .sa_snapshot( 
	\num_26_._zy_simnet_tvar_136 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_26_._zy_simnet_tvar_137 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_26_._zy_simnet_sa_clear_138_w$ ), .sa_snap( 
	\num_26_._zy_simnet_sa_snap_139_w$ ));
ixc_assign \num_26_._zz_strnp_134 ( \num_26_._zy_simnet_sa_snap_139_w$ , 
	sa_snap);
ixc_assign \num_26_._zz_strnp_133 ( \num_26_._zy_simnet_sa_clear_138_w$ , 
	sa_clear);
ixc_assign_50 \num_26_._zz_strnp_131 ( { \sa_snapshot[26][49] , 
	\sa_snapshot[26][48] , \sa_snapshot[26][47] , \sa_snapshot[26][46] , 
	\sa_snapshot[26][45] , \sa_snapshot[26][44] , \sa_snapshot[26][43] , 
	\sa_snapshot[26][42] , \sa_snapshot[26][41] , \sa_snapshot[26][40] , 
	\sa_snapshot[26][39] , \sa_snapshot[26][38] , \sa_snapshot[26][37] , 
	\sa_snapshot[26][36] , \sa_snapshot[26][35] , \sa_snapshot[26][34] , 
	\sa_snapshot[26][33] , \sa_snapshot[26][32] , \sa_snapshot[26][31] , 
	\sa_snapshot[26][30] , \sa_snapshot[26][29] , \sa_snapshot[26][28] , 
	\sa_snapshot[26][27] , \sa_snapshot[26][26] , \sa_snapshot[26][25] , 
	\sa_snapshot[26][24] , \sa_snapshot[26][23] , \sa_snapshot[26][22] , 
	\sa_snapshot[26][21] , \sa_snapshot[26][20] , \sa_snapshot[26][19] , 
	\sa_snapshot[26][18] , \sa_snapshot[26][17] , \sa_snapshot[26][16] , 
	\sa_snapshot[26][15] , \sa_snapshot[26][14] , \sa_snapshot[26][13] , 
	\sa_snapshot[26][12] , \sa_snapshot[26][11] , \sa_snapshot[26][10] , 
	\sa_snapshot[26][9] , \sa_snapshot[26][8] , \sa_snapshot[26][7] , 
	\sa_snapshot[26][6] , \sa_snapshot[26][5] , \sa_snapshot[26][4] , 
	\sa_snapshot[26][3] , \sa_snapshot[26][2] , \sa_snapshot[26][1] , 
	\sa_snapshot[26][0] }, \num_26_._zy_simnet_tvar_136 [0:49]);
ixc_assign_50 \num_26_._zz_strnp_130 ( { \sa_count[26][49] , 
	\sa_count[26][48] , \sa_count[26][47] , \sa_count[26][46] , 
	\sa_count[26][45] , \sa_count[26][44] , \sa_count[26][43] , 
	\sa_count[26][42] , \sa_count[26][41] , \sa_count[26][40] , 
	\sa_count[26][39] , \sa_count[26][38] , \sa_count[26][37] , 
	\sa_count[26][36] , \sa_count[26][35] , \sa_count[26][34] , 
	\sa_count[26][33] , \sa_count[26][32] , \sa_count[26][31] , 
	\sa_count[26][30] , \sa_count[26][29] , \sa_count[26][28] , 
	\sa_count[26][27] , \sa_count[26][26] , \sa_count[26][25] , 
	\sa_count[26][24] , \sa_count[26][23] , \sa_count[26][22] , 
	\sa_count[26][21] , \sa_count[26][20] , \sa_count[26][19] , 
	\sa_count[26][18] , \sa_count[26][17] , \sa_count[26][16] , 
	\sa_count[26][15] , \sa_count[26][14] , \sa_count[26][13] , 
	\sa_count[26][12] , \sa_count[26][11] , \sa_count[26][10] , 
	\sa_count[26][9] , \sa_count[26][8] , \sa_count[26][7] , 
	\sa_count[26][6] , \sa_count[26][5] , \sa_count[26][4] , 
	\sa_count[26][3] , \sa_count[26][2] , \sa_count[26][1] , 
	\sa_count[26][0] }, \num_26_._zy_simnet_tvar_135 [0:49]);
ixc_assign_10 \num_27_._zz_strnp_137 ( \num_27_._zy_simnet_tvar_142 [0:9], { 
	n220, n219, n218, n217, n216, \sa_ctrl[27][4] , \sa_ctrl[27][3] , 
	\sa_ctrl[27][2] , \sa_ctrl[27][1] , \sa_ctrl[27][0] });
cr_sa_counter \num_27_.sa_counter_i ( .sa_count( 
	\num_27_._zy_simnet_tvar_140 [0:49]), .sa_snapshot( 
	\num_27_._zy_simnet_tvar_141 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_27_._zy_simnet_tvar_142 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_27_._zy_simnet_sa_clear_143_w$ ), .sa_snap( 
	\num_27_._zy_simnet_sa_snap_144_w$ ));
ixc_assign \num_27_._zz_strnp_139 ( \num_27_._zy_simnet_sa_snap_144_w$ , 
	sa_snap);
ixc_assign \num_27_._zz_strnp_138 ( \num_27_._zy_simnet_sa_clear_143_w$ , 
	sa_clear);
ixc_assign_50 \num_27_._zz_strnp_136 ( { \sa_snapshot[27][49] , 
	\sa_snapshot[27][48] , \sa_snapshot[27][47] , \sa_snapshot[27][46] , 
	\sa_snapshot[27][45] , \sa_snapshot[27][44] , \sa_snapshot[27][43] , 
	\sa_snapshot[27][42] , \sa_snapshot[27][41] , \sa_snapshot[27][40] , 
	\sa_snapshot[27][39] , \sa_snapshot[27][38] , \sa_snapshot[27][37] , 
	\sa_snapshot[27][36] , \sa_snapshot[27][35] , \sa_snapshot[27][34] , 
	\sa_snapshot[27][33] , \sa_snapshot[27][32] , \sa_snapshot[27][31] , 
	\sa_snapshot[27][30] , \sa_snapshot[27][29] , \sa_snapshot[27][28] , 
	\sa_snapshot[27][27] , \sa_snapshot[27][26] , \sa_snapshot[27][25] , 
	\sa_snapshot[27][24] , \sa_snapshot[27][23] , \sa_snapshot[27][22] , 
	\sa_snapshot[27][21] , \sa_snapshot[27][20] , \sa_snapshot[27][19] , 
	\sa_snapshot[27][18] , \sa_snapshot[27][17] , \sa_snapshot[27][16] , 
	\sa_snapshot[27][15] , \sa_snapshot[27][14] , \sa_snapshot[27][13] , 
	\sa_snapshot[27][12] , \sa_snapshot[27][11] , \sa_snapshot[27][10] , 
	\sa_snapshot[27][9] , \sa_snapshot[27][8] , \sa_snapshot[27][7] , 
	\sa_snapshot[27][6] , \sa_snapshot[27][5] , \sa_snapshot[27][4] , 
	\sa_snapshot[27][3] , \sa_snapshot[27][2] , \sa_snapshot[27][1] , 
	\sa_snapshot[27][0] }, \num_27_._zy_simnet_tvar_141 [0:49]);
ixc_assign_50 \num_27_._zz_strnp_135 ( { \sa_count[27][49] , 
	\sa_count[27][48] , \sa_count[27][47] , \sa_count[27][46] , 
	\sa_count[27][45] , \sa_count[27][44] , \sa_count[27][43] , 
	\sa_count[27][42] , \sa_count[27][41] , \sa_count[27][40] , 
	\sa_count[27][39] , \sa_count[27][38] , \sa_count[27][37] , 
	\sa_count[27][36] , \sa_count[27][35] , \sa_count[27][34] , 
	\sa_count[27][33] , \sa_count[27][32] , \sa_count[27][31] , 
	\sa_count[27][30] , \sa_count[27][29] , \sa_count[27][28] , 
	\sa_count[27][27] , \sa_count[27][26] , \sa_count[27][25] , 
	\sa_count[27][24] , \sa_count[27][23] , \sa_count[27][22] , 
	\sa_count[27][21] , \sa_count[27][20] , \sa_count[27][19] , 
	\sa_count[27][18] , \sa_count[27][17] , \sa_count[27][16] , 
	\sa_count[27][15] , \sa_count[27][14] , \sa_count[27][13] , 
	\sa_count[27][12] , \sa_count[27][11] , \sa_count[27][10] , 
	\sa_count[27][9] , \sa_count[27][8] , \sa_count[27][7] , 
	\sa_count[27][6] , \sa_count[27][5] , \sa_count[27][4] , 
	\sa_count[27][3] , \sa_count[27][2] , \sa_count[27][1] , 
	\sa_count[27][0] }, \num_27_._zy_simnet_tvar_140 [0:49]);
ixc_assign_10 \num_28_._zz_strnp_142 ( \num_28_._zy_simnet_tvar_147 [0:9], { 
	n225, n224, n223, n222, n221, \sa_ctrl[28][4] , \sa_ctrl[28][3] , 
	\sa_ctrl[28][2] , \sa_ctrl[28][1] , \sa_ctrl[28][0] });
cr_sa_counter \num_28_.sa_counter_i ( .sa_count( 
	\num_28_._zy_simnet_tvar_145 [0:49]), .sa_snapshot( 
	\num_28_._zy_simnet_tvar_146 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_28_._zy_simnet_tvar_147 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_28_._zy_simnet_sa_clear_148_w$ ), .sa_snap( 
	\num_28_._zy_simnet_sa_snap_149_w$ ));
ixc_assign \num_28_._zz_strnp_144 ( \num_28_._zy_simnet_sa_snap_149_w$ , 
	sa_snap);
ixc_assign \num_28_._zz_strnp_143 ( \num_28_._zy_simnet_sa_clear_148_w$ , 
	sa_clear);
ixc_assign_50 \num_28_._zz_strnp_141 ( { \sa_snapshot[28][49] , 
	\sa_snapshot[28][48] , \sa_snapshot[28][47] , \sa_snapshot[28][46] , 
	\sa_snapshot[28][45] , \sa_snapshot[28][44] , \sa_snapshot[28][43] , 
	\sa_snapshot[28][42] , \sa_snapshot[28][41] , \sa_snapshot[28][40] , 
	\sa_snapshot[28][39] , \sa_snapshot[28][38] , \sa_snapshot[28][37] , 
	\sa_snapshot[28][36] , \sa_snapshot[28][35] , \sa_snapshot[28][34] , 
	\sa_snapshot[28][33] , \sa_snapshot[28][32] , \sa_snapshot[28][31] , 
	\sa_snapshot[28][30] , \sa_snapshot[28][29] , \sa_snapshot[28][28] , 
	\sa_snapshot[28][27] , \sa_snapshot[28][26] , \sa_snapshot[28][25] , 
	\sa_snapshot[28][24] , \sa_snapshot[28][23] , \sa_snapshot[28][22] , 
	\sa_snapshot[28][21] , \sa_snapshot[28][20] , \sa_snapshot[28][19] , 
	\sa_snapshot[28][18] , \sa_snapshot[28][17] , \sa_snapshot[28][16] , 
	\sa_snapshot[28][15] , \sa_snapshot[28][14] , \sa_snapshot[28][13] , 
	\sa_snapshot[28][12] , \sa_snapshot[28][11] , \sa_snapshot[28][10] , 
	\sa_snapshot[28][9] , \sa_snapshot[28][8] , \sa_snapshot[28][7] , 
	\sa_snapshot[28][6] , \sa_snapshot[28][5] , \sa_snapshot[28][4] , 
	\sa_snapshot[28][3] , \sa_snapshot[28][2] , \sa_snapshot[28][1] , 
	\sa_snapshot[28][0] }, \num_28_._zy_simnet_tvar_146 [0:49]);
ixc_assign_50 \num_28_._zz_strnp_140 ( { \sa_count[28][49] , 
	\sa_count[28][48] , \sa_count[28][47] , \sa_count[28][46] , 
	\sa_count[28][45] , \sa_count[28][44] , \sa_count[28][43] , 
	\sa_count[28][42] , \sa_count[28][41] , \sa_count[28][40] , 
	\sa_count[28][39] , \sa_count[28][38] , \sa_count[28][37] , 
	\sa_count[28][36] , \sa_count[28][35] , \sa_count[28][34] , 
	\sa_count[28][33] , \sa_count[28][32] , \sa_count[28][31] , 
	\sa_count[28][30] , \sa_count[28][29] , \sa_count[28][28] , 
	\sa_count[28][27] , \sa_count[28][26] , \sa_count[28][25] , 
	\sa_count[28][24] , \sa_count[28][23] , \sa_count[28][22] , 
	\sa_count[28][21] , \sa_count[28][20] , \sa_count[28][19] , 
	\sa_count[28][18] , \sa_count[28][17] , \sa_count[28][16] , 
	\sa_count[28][15] , \sa_count[28][14] , \sa_count[28][13] , 
	\sa_count[28][12] , \sa_count[28][11] , \sa_count[28][10] , 
	\sa_count[28][9] , \sa_count[28][8] , \sa_count[28][7] , 
	\sa_count[28][6] , \sa_count[28][5] , \sa_count[28][4] , 
	\sa_count[28][3] , \sa_count[28][2] , \sa_count[28][1] , 
	\sa_count[28][0] }, \num_28_._zy_simnet_tvar_145 [0:49]);
ixc_assign_10 \num_29_._zz_strnp_147 ( \num_29_._zy_simnet_tvar_152 [0:9], { 
	n230, n229, n228, n227, n226, \sa_ctrl[29][4] , \sa_ctrl[29][3] , 
	\sa_ctrl[29][2] , \sa_ctrl[29][1] , \sa_ctrl[29][0] });
cr_sa_counter \num_29_.sa_counter_i ( .sa_count( 
	\num_29_._zy_simnet_tvar_150 [0:49]), .sa_snapshot( 
	\num_29_._zy_simnet_tvar_151 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_29_._zy_simnet_tvar_152 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_29_._zy_simnet_sa_clear_153_w$ ), .sa_snap( 
	\num_29_._zy_simnet_sa_snap_154_w$ ));
ixc_assign \num_29_._zz_strnp_149 ( \num_29_._zy_simnet_sa_snap_154_w$ , 
	sa_snap);
ixc_assign \num_29_._zz_strnp_148 ( \num_29_._zy_simnet_sa_clear_153_w$ , 
	sa_clear);
ixc_assign_50 \num_29_._zz_strnp_146 ( { \sa_snapshot[29][49] , 
	\sa_snapshot[29][48] , \sa_snapshot[29][47] , \sa_snapshot[29][46] , 
	\sa_snapshot[29][45] , \sa_snapshot[29][44] , \sa_snapshot[29][43] , 
	\sa_snapshot[29][42] , \sa_snapshot[29][41] , \sa_snapshot[29][40] , 
	\sa_snapshot[29][39] , \sa_snapshot[29][38] , \sa_snapshot[29][37] , 
	\sa_snapshot[29][36] , \sa_snapshot[29][35] , \sa_snapshot[29][34] , 
	\sa_snapshot[29][33] , \sa_snapshot[29][32] , \sa_snapshot[29][31] , 
	\sa_snapshot[29][30] , \sa_snapshot[29][29] , \sa_snapshot[29][28] , 
	\sa_snapshot[29][27] , \sa_snapshot[29][26] , \sa_snapshot[29][25] , 
	\sa_snapshot[29][24] , \sa_snapshot[29][23] , \sa_snapshot[29][22] , 
	\sa_snapshot[29][21] , \sa_snapshot[29][20] , \sa_snapshot[29][19] , 
	\sa_snapshot[29][18] , \sa_snapshot[29][17] , \sa_snapshot[29][16] , 
	\sa_snapshot[29][15] , \sa_snapshot[29][14] , \sa_snapshot[29][13] , 
	\sa_snapshot[29][12] , \sa_snapshot[29][11] , \sa_snapshot[29][10] , 
	\sa_snapshot[29][9] , \sa_snapshot[29][8] , \sa_snapshot[29][7] , 
	\sa_snapshot[29][6] , \sa_snapshot[29][5] , \sa_snapshot[29][4] , 
	\sa_snapshot[29][3] , \sa_snapshot[29][2] , \sa_snapshot[29][1] , 
	\sa_snapshot[29][0] }, \num_29_._zy_simnet_tvar_151 [0:49]);
ixc_assign_50 \num_29_._zz_strnp_145 ( { \sa_count[29][49] , 
	\sa_count[29][48] , \sa_count[29][47] , \sa_count[29][46] , 
	\sa_count[29][45] , \sa_count[29][44] , \sa_count[29][43] , 
	\sa_count[29][42] , \sa_count[29][41] , \sa_count[29][40] , 
	\sa_count[29][39] , \sa_count[29][38] , \sa_count[29][37] , 
	\sa_count[29][36] , \sa_count[29][35] , \sa_count[29][34] , 
	\sa_count[29][33] , \sa_count[29][32] , \sa_count[29][31] , 
	\sa_count[29][30] , \sa_count[29][29] , \sa_count[29][28] , 
	\sa_count[29][27] , \sa_count[29][26] , \sa_count[29][25] , 
	\sa_count[29][24] , \sa_count[29][23] , \sa_count[29][22] , 
	\sa_count[29][21] , \sa_count[29][20] , \sa_count[29][19] , 
	\sa_count[29][18] , \sa_count[29][17] , \sa_count[29][16] , 
	\sa_count[29][15] , \sa_count[29][14] , \sa_count[29][13] , 
	\sa_count[29][12] , \sa_count[29][11] , \sa_count[29][10] , 
	\sa_count[29][9] , \sa_count[29][8] , \sa_count[29][7] , 
	\sa_count[29][6] , \sa_count[29][5] , \sa_count[29][4] , 
	\sa_count[29][3] , \sa_count[29][2] , \sa_count[29][1] , 
	\sa_count[29][0] }, \num_29_._zy_simnet_tvar_150 [0:49]);
ixc_assign_10 \num_30_._zz_strnp_152 ( \num_30_._zy_simnet_tvar_157 [0:9], { 
	n235, n234, n233, n232, n231, \sa_ctrl[30][4] , \sa_ctrl[30][3] , 
	\sa_ctrl[30][2] , \sa_ctrl[30][1] , \sa_ctrl[30][0] });
cr_sa_counter \num_30_.sa_counter_i ( .sa_count( 
	\num_30_._zy_simnet_tvar_155 [0:49]), .sa_snapshot( 
	\num_30_._zy_simnet_tvar_156 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_30_._zy_simnet_tvar_157 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_30_._zy_simnet_sa_clear_158_w$ ), .sa_snap( 
	\num_30_._zy_simnet_sa_snap_159_w$ ));
ixc_assign \num_30_._zz_strnp_154 ( \num_30_._zy_simnet_sa_snap_159_w$ , 
	sa_snap);
ixc_assign \num_30_._zz_strnp_153 ( \num_30_._zy_simnet_sa_clear_158_w$ , 
	sa_clear);
ixc_assign_50 \num_30_._zz_strnp_151 ( { \sa_snapshot[30][49] , 
	\sa_snapshot[30][48] , \sa_snapshot[30][47] , \sa_snapshot[30][46] , 
	\sa_snapshot[30][45] , \sa_snapshot[30][44] , \sa_snapshot[30][43] , 
	\sa_snapshot[30][42] , \sa_snapshot[30][41] , \sa_snapshot[30][40] , 
	\sa_snapshot[30][39] , \sa_snapshot[30][38] , \sa_snapshot[30][37] , 
	\sa_snapshot[30][36] , \sa_snapshot[30][35] , \sa_snapshot[30][34] , 
	\sa_snapshot[30][33] , \sa_snapshot[30][32] , \sa_snapshot[30][31] , 
	\sa_snapshot[30][30] , \sa_snapshot[30][29] , \sa_snapshot[30][28] , 
	\sa_snapshot[30][27] , \sa_snapshot[30][26] , \sa_snapshot[30][25] , 
	\sa_snapshot[30][24] , \sa_snapshot[30][23] , \sa_snapshot[30][22] , 
	\sa_snapshot[30][21] , \sa_snapshot[30][20] , \sa_snapshot[30][19] , 
	\sa_snapshot[30][18] , \sa_snapshot[30][17] , \sa_snapshot[30][16] , 
	\sa_snapshot[30][15] , \sa_snapshot[30][14] , \sa_snapshot[30][13] , 
	\sa_snapshot[30][12] , \sa_snapshot[30][11] , \sa_snapshot[30][10] , 
	\sa_snapshot[30][9] , \sa_snapshot[30][8] , \sa_snapshot[30][7] , 
	\sa_snapshot[30][6] , \sa_snapshot[30][5] , \sa_snapshot[30][4] , 
	\sa_snapshot[30][3] , \sa_snapshot[30][2] , \sa_snapshot[30][1] , 
	\sa_snapshot[30][0] }, \num_30_._zy_simnet_tvar_156 [0:49]);
ixc_assign_50 \num_30_._zz_strnp_150 ( { \sa_count[30][49] , 
	\sa_count[30][48] , \sa_count[30][47] , \sa_count[30][46] , 
	\sa_count[30][45] , \sa_count[30][44] , \sa_count[30][43] , 
	\sa_count[30][42] , \sa_count[30][41] , \sa_count[30][40] , 
	\sa_count[30][39] , \sa_count[30][38] , \sa_count[30][37] , 
	\sa_count[30][36] , \sa_count[30][35] , \sa_count[30][34] , 
	\sa_count[30][33] , \sa_count[30][32] , \sa_count[30][31] , 
	\sa_count[30][30] , \sa_count[30][29] , \sa_count[30][28] , 
	\sa_count[30][27] , \sa_count[30][26] , \sa_count[30][25] , 
	\sa_count[30][24] , \sa_count[30][23] , \sa_count[30][22] , 
	\sa_count[30][21] , \sa_count[30][20] , \sa_count[30][19] , 
	\sa_count[30][18] , \sa_count[30][17] , \sa_count[30][16] , 
	\sa_count[30][15] , \sa_count[30][14] , \sa_count[30][13] , 
	\sa_count[30][12] , \sa_count[30][11] , \sa_count[30][10] , 
	\sa_count[30][9] , \sa_count[30][8] , \sa_count[30][7] , 
	\sa_count[30][6] , \sa_count[30][5] , \sa_count[30][4] , 
	\sa_count[30][3] , \sa_count[30][2] , \sa_count[30][1] , 
	\sa_count[30][0] }, \num_30_._zy_simnet_tvar_155 [0:49]);
ixc_assign_10 \num_31_._zz_strnp_157 ( \num_31_._zy_simnet_tvar_162 [0:9], { 
	n240, n239, n238, n237, n236, \sa_ctrl[31][4] , \sa_ctrl[31][3] , 
	\sa_ctrl[31][2] , \sa_ctrl[31][1] , \sa_ctrl[31][0] });
cr_sa_counter \num_31_.sa_counter_i ( .sa_count( 
	\num_31_._zy_simnet_tvar_160 [0:49]), .sa_snapshot( 
	\num_31_._zy_simnet_tvar_161 [0:49]), .clk( clk), .rst_n( rst_n), 
	.sa_event_sel( \num_31_._zy_simnet_tvar_162 [0:9]), .sa_events( { 
	\sa_events[15][63] , \sa_events[15][62] , \sa_events[15][61] , 
	\sa_events[15][60] , \sa_events[15][59] , \sa_events[15][58] , 
	\sa_events[15][57] , \sa_events[15][56] , \sa_events[15][55] , 
	\sa_events[15][54] , \sa_events[15][53] , \sa_events[15][52] , 
	\sa_events[15][51] , \sa_events[15][50] , \sa_events[15][49] , 
	\sa_events[15][48] , \sa_events[15][47] , \sa_events[15][46] , 
	\sa_events[15][45] , \sa_events[15][44] , \sa_events[15][43] , 
	\sa_events[15][42] , \sa_events[15][41] , \sa_events[15][40] , 
	\sa_events[15][39] , \sa_events[15][38] , \sa_events[15][37] , 
	\sa_events[15][36] , \sa_events[15][35] , \sa_events[15][34] , 
	\sa_events[15][33] , \sa_events[15][32] , \sa_events[15][31] , 
	\sa_events[15][30] , \sa_events[15][29] , \sa_events[15][28] , 
	\sa_events[15][27] , \sa_events[15][26] , \sa_events[15][25] , 
	\sa_events[15][24] , \sa_events[15][23] , \sa_events[15][22] , 
	\sa_events[15][21] , \sa_events[15][20] , \sa_events[15][19] , 
	\sa_events[15][18] , \sa_events[15][17] , \sa_events[15][16] , 
	\sa_events[15][15] , \sa_events[15][14] , \sa_events[15][13] , 
	\sa_events[15][12] , \sa_events[15][11] , \sa_events[15][10] , 
	\sa_events[15][9] , \sa_events[15][8] , \sa_events[15][7] , 
	\sa_events[15][6] , \sa_events[15][5] , \sa_events[15][4] , 
	\sa_events[15][3] , \sa_events[15][2] , \sa_events[15][1] , 
	\sa_events[15][0] , \sa_events[14][63] , \sa_events[14][62] , 
	\sa_events[14][61] , \sa_events[14][60] , \sa_events[14][59] , 
	\sa_events[14][58] , \sa_events[14][57] , \sa_events[14][56] , 
	\sa_events[14][55] , \sa_events[14][54] , \sa_events[14][53] , 
	\sa_events[14][52] , \sa_events[14][51] , \sa_events[14][50] , 
	\sa_events[14][49] , \sa_events[14][48] , \sa_events[14][47] , 
	\sa_events[14][46] , \sa_events[14][45] , \sa_events[14][44] , 
	\sa_events[14][43] , \sa_events[14][42] , \sa_events[14][41] , 
	\sa_events[14][40] , \sa_events[14][39] , \sa_events[14][38] , 
	\sa_events[14][37] , \sa_events[14][36] , \sa_events[14][35] , 
	\sa_events[14][34] , \sa_events[14][33] , \sa_events[14][32] , 
	\sa_events[14][31] , \sa_events[14][30] , \sa_events[14][29] , 
	\sa_events[14][28] , \sa_events[14][27] , \sa_events[14][26] , 
	\sa_events[14][25] , \sa_events[14][24] , \sa_events[14][23] , 
	\sa_events[14][22] , \sa_events[14][21] , \sa_events[14][20] , 
	\sa_events[14][19] , \sa_events[14][18] , \sa_events[14][17] , 
	\sa_events[14][16] , \sa_events[14][15] , \sa_events[14][14] , 
	\sa_events[14][13] , \sa_events[14][12] , \sa_events[14][11] , 
	\sa_events[14][10] , \sa_events[14][9] , \sa_events[14][8] , 
	\sa_events[14][7] , \sa_events[14][6] , \sa_events[14][5] , 
	\sa_events[14][4] , \sa_events[14][3] , \sa_events[14][2] , 
	\sa_events[14][1] , \sa_events[14][0] , \sa_events[13][63] , 
	\sa_events[13][62] , \sa_events[13][61] , \sa_events[13][60] , 
	\sa_events[13][59] , \sa_events[13][58] , \sa_events[13][57] , 
	\sa_events[13][56] , \sa_events[13][55] , \sa_events[13][54] , 
	\sa_events[13][53] , \sa_events[13][52] , \sa_events[13][51] , 
	\sa_events[13][50] , \sa_events[13][49] , \sa_events[13][48] , 
	\sa_events[13][47] , \sa_events[13][46] , \sa_events[13][45] , 
	\sa_events[13][44] , \sa_events[13][43] , \sa_events[13][42] , 
	\sa_events[13][41] , \sa_events[13][40] , \sa_events[13][39] , 
	\sa_events[13][38] , \sa_events[13][37] , \sa_events[13][36] , 
	\sa_events[13][35] , \sa_events[13][34] , \sa_events[13][33] , 
	\sa_events[13][32] , \sa_events[13][31] , \sa_events[13][30] , 
	\sa_events[13][29] , \sa_events[13][28] , \sa_events[13][27] , 
	\sa_events[13][26] , \sa_events[13][25] , \sa_events[13][24] , 
	\sa_events[13][23] , \sa_events[13][22] , \sa_events[13][21] , 
	\sa_events[13][20] , \sa_events[13][19] , \sa_events[13][18] , 
	\sa_events[13][17] , \sa_events[13][16] , \sa_events[13][15] , 
	\sa_events[13][14] , \sa_events[13][13] , \sa_events[13][12] , 
	\sa_events[13][11] , \sa_events[13][10] , \sa_events[13][9] , 
	\sa_events[13][8] , \sa_events[13][7] , \sa_events[13][6] , 
	\sa_events[13][5] , \sa_events[13][4] , \sa_events[13][3] , 
	\sa_events[13][2] , \sa_events[13][1] , \sa_events[13][0] , 
	\sa_events[12][63] , \sa_events[12][62] , \sa_events[12][61] , 
	\sa_events[12][60] , \sa_events[12][59] , \sa_events[12][58] , 
	\sa_events[12][57] , \sa_events[12][56] , \sa_events[12][55] , 
	\sa_events[12][54] , \sa_events[12][53] , \sa_events[12][52] , 
	\sa_events[12][51] , \sa_events[12][50] , \sa_events[12][49] , 
	\sa_events[12][48] , \sa_events[12][47] , \sa_events[12][46] , 
	\sa_events[12][45] , \sa_events[12][44] , \sa_events[12][43] , 
	\sa_events[12][42] , \sa_events[12][41] , \sa_events[12][40] , 
	\sa_events[12][39] , \sa_events[12][38] , \sa_events[12][37] , 
	\sa_events[12][36] , \sa_events[12][35] , \sa_events[12][34] , 
	\sa_events[12][33] , \sa_events[12][32] , \sa_events[12][31] , 
	\sa_events[12][30] , \sa_events[12][29] , \sa_events[12][28] , 
	\sa_events[12][27] , \sa_events[12][26] , \sa_events[12][25] , 
	\sa_events[12][24] , \sa_events[12][23] , \sa_events[12][22] , 
	\sa_events[12][21] , \sa_events[12][20] , \sa_events[12][19] , 
	\sa_events[12][18] , \sa_events[12][17] , \sa_events[12][16] , 
	\sa_events[12][15] , \sa_events[12][14] , \sa_events[12][13] , 
	\sa_events[12][12] , \sa_events[12][11] , \sa_events[12][10] , 
	\sa_events[12][9] , \sa_events[12][8] , \sa_events[12][7] , 
	\sa_events[12][6] , \sa_events[12][5] , \sa_events[12][4] , 
	\sa_events[12][3] , \sa_events[12][2] , \sa_events[12][1] , 
	\sa_events[12][0] , \sa_events[11][63] , \sa_events[11][62] , 
	\sa_events[11][61] , \sa_events[11][60] , \sa_events[11][59] , 
	\sa_events[11][58] , \sa_events[11][57] , \sa_events[11][56] , 
	\sa_events[11][55] , \sa_events[11][54] , \sa_events[11][53] , 
	\sa_events[11][52] , \sa_events[11][51] , \sa_events[11][50] , 
	\sa_events[11][49] , \sa_events[11][48] , \sa_events[11][47] , 
	\sa_events[11][46] , \sa_events[11][45] , \sa_events[11][44] , 
	\sa_events[11][43] , \sa_events[11][42] , \sa_events[11][41] , 
	\sa_events[11][40] , \sa_events[11][39] , \sa_events[11][38] , 
	\sa_events[11][37] , \sa_events[11][36] , \sa_events[11][35] , 
	\sa_events[11][34] , \sa_events[11][33] , \sa_events[11][32] , 
	\sa_events[11][31] , \sa_events[11][30] , \sa_events[11][29] , 
	\sa_events[11][28] , \sa_events[11][27] , \sa_events[11][26] , 
	\sa_events[11][25] , \sa_events[11][24] , \sa_events[11][23] , 
	\sa_events[11][22] , \sa_events[11][21] , \sa_events[11][20] , 
	\sa_events[11][19] , \sa_events[11][18] , \sa_events[11][17] , 
	\sa_events[11][16] , \sa_events[11][15] , \sa_events[11][14] , 
	\sa_events[11][13] , \sa_events[11][12] , \sa_events[11][11] , 
	\sa_events[11][10] , \sa_events[11][9] , \sa_events[11][8] , 
	\sa_events[11][7] , \sa_events[11][6] , \sa_events[11][5] , 
	\sa_events[11][4] , \sa_events[11][3] , \sa_events[11][2] , 
	\sa_events[11][1] , \sa_events[11][0] , \sa_events[10][63] , 
	\sa_events[10][62] , \sa_events[10][61] , \sa_events[10][60] , 
	\sa_events[10][59] , \sa_events[10][58] , \sa_events[10][57] , 
	\sa_events[10][56] , \sa_events[10][55] , \sa_events[10][54] , 
	\sa_events[10][53] , \sa_events[10][52] , \sa_events[10][51] , 
	\sa_events[10][50] , \sa_events[10][49] , \sa_events[10][48] , 
	\sa_events[10][47] , \sa_events[10][46] , \sa_events[10][45] , 
	\sa_events[10][44] , \sa_events[10][43] , \sa_events[10][42] , 
	\sa_events[10][41] , \sa_events[10][40] , \sa_events[10][39] , 
	\sa_events[10][38] , \sa_events[10][37] , \sa_events[10][36] , 
	\sa_events[10][35] , \sa_events[10][34] , \sa_events[10][33] , 
	\sa_events[10][32] , \sa_events[10][31] , \sa_events[10][30] , 
	\sa_events[10][29] , \sa_events[10][28] , \sa_events[10][27] , 
	\sa_events[10][26] , \sa_events[10][25] , \sa_events[10][24] , 
	\sa_events[10][23] , \sa_events[10][22] , \sa_events[10][21] , 
	\sa_events[10][20] , \sa_events[10][19] , \sa_events[10][18] , 
	\sa_events[10][17] , \sa_events[10][16] , \sa_events[10][15] , 
	\sa_events[10][14] , \sa_events[10][13] , \sa_events[10][12] , 
	\sa_events[10][11] , \sa_events[10][10] , \sa_events[10][9] , 
	\sa_events[10][8] , \sa_events[10][7] , \sa_events[10][6] , 
	\sa_events[10][5] , \sa_events[10][4] , \sa_events[10][3] , 
	\sa_events[10][2] , \sa_events[10][1] , \sa_events[10][0] , 
	\sa_events[9][63] , \sa_events[9][62] , \sa_events[9][61] , 
	\sa_events[9][60] , \sa_events[9][59] , \sa_events[9][58] , 
	\sa_events[9][57] , \sa_events[9][56] , \sa_events[9][55] , 
	\sa_events[9][54] , \sa_events[9][53] , \sa_events[9][52] , 
	\sa_events[9][51] , \sa_events[9][50] , \sa_events[9][49] , 
	\sa_events[9][48] , \sa_events[9][47] , \sa_events[9][46] , 
	\sa_events[9][45] , \sa_events[9][44] , \sa_events[9][43] , 
	\sa_events[9][42] , \sa_events[9][41] , \sa_events[9][40] , 
	\sa_events[9][39] , \sa_events[9][38] , \sa_events[9][37] , 
	\sa_events[9][36] , \sa_events[9][35] , \sa_events[9][34] , 
	\sa_events[9][33] , \sa_events[9][32] , \sa_events[9][31] , 
	\sa_events[9][30] , \sa_events[9][29] , \sa_events[9][28] , 
	\sa_events[9][27] , \sa_events[9][26] , \sa_events[9][25] , 
	\sa_events[9][24] , \sa_events[9][23] , \sa_events[9][22] , 
	\sa_events[9][21] , \sa_events[9][20] , \sa_events[9][19] , 
	\sa_events[9][18] , \sa_events[9][17] , \sa_events[9][16] , 
	\sa_events[9][15] , \sa_events[9][14] , \sa_events[9][13] , 
	\sa_events[9][12] , \sa_events[9][11] , \sa_events[9][10] , 
	\sa_events[9][9] , \sa_events[9][8] , \sa_events[9][7] , 
	\sa_events[9][6] , \sa_events[9][5] , \sa_events[9][4] , 
	\sa_events[9][3] , \sa_events[9][2] , \sa_events[9][1] , 
	\sa_events[9][0] , \sa_events[8][63] , \sa_events[8][62] , 
	\sa_events[8][61] , \sa_events[8][60] , \sa_events[8][59] , 
	\sa_events[8][58] , \sa_events[8][57] , \sa_events[8][56] , 
	\sa_events[8][55] , \sa_events[8][54] , \sa_events[8][53] , 
	\sa_events[8][52] , \sa_events[8][51] , \sa_events[8][50] , 
	\sa_events[8][49] , \sa_events[8][48] , \sa_events[8][47] , 
	\sa_events[8][46] , \sa_events[8][45] , \sa_events[8][44] , 
	\sa_events[8][43] , \sa_events[8][42] , \sa_events[8][41] , 
	\sa_events[8][40] , \sa_events[8][39] , \sa_events[8][38] , 
	\sa_events[8][37] , \sa_events[8][36] , \sa_events[8][35] , 
	\sa_events[8][34] , \sa_events[8][33] , \sa_events[8][32] , 
	\sa_events[8][31] , \sa_events[8][30] , \sa_events[8][29] , 
	\sa_events[8][28] , \sa_events[8][27] , \sa_events[8][26] , 
	\sa_events[8][25] , \sa_events[8][24] , \sa_events[8][23] , 
	\sa_events[8][22] , \sa_events[8][21] , \sa_events[8][20] , 
	\sa_events[8][19] , \sa_events[8][18] , \sa_events[8][17] , 
	\sa_events[8][16] , \sa_events[8][15] , \sa_events[8][14] , 
	\sa_events[8][13] , \sa_events[8][12] , \sa_events[8][11] , 
	\sa_events[8][10] , \sa_events[8][9] , \sa_events[8][8] , 
	\sa_events[8][7] , \sa_events[8][6] , \sa_events[8][5] , 
	\sa_events[8][4] , \sa_events[8][3] , \sa_events[8][2] , 
	\sa_events[8][1] , \sa_events[8][0] , \sa_events[7][63] , 
	\sa_events[7][62] , \sa_events[7][61] , \sa_events[7][60] , 
	\sa_events[7][59] , \sa_events[7][58] , \sa_events[7][57] , 
	\sa_events[7][56] , \sa_events[7][55] , \sa_events[7][54] , 
	\sa_events[7][53] , \sa_events[7][52] , \sa_events[7][51] , 
	\sa_events[7][50] , \sa_events[7][49] , \sa_events[7][48] , 
	\sa_events[7][47] , \sa_events[7][46] , \sa_events[7][45] , 
	\sa_events[7][44] , \sa_events[7][43] , \sa_events[7][42] , 
	\sa_events[7][41] , \sa_events[7][40] , \sa_events[7][39] , 
	\sa_events[7][38] , \sa_events[7][37] , \sa_events[7][36] , 
	\sa_events[7][35] , \sa_events[7][34] , \sa_events[7][33] , 
	\sa_events[7][32] , \sa_events[7][31] , \sa_events[7][30] , 
	\sa_events[7][29] , \sa_events[7][28] , \sa_events[7][27] , 
	\sa_events[7][26] , \sa_events[7][25] , \sa_events[7][24] , 
	\sa_events[7][23] , \sa_events[7][22] , \sa_events[7][21] , 
	\sa_events[7][20] , \sa_events[7][19] , \sa_events[7][18] , 
	\sa_events[7][17] , \sa_events[7][16] , \sa_events[7][15] , 
	\sa_events[7][14] , \sa_events[7][13] , \sa_events[7][12] , 
	\sa_events[7][11] , \sa_events[7][10] , \sa_events[7][9] , 
	\sa_events[7][8] , \sa_events[7][7] , \sa_events[7][6] , 
	\sa_events[7][5] , \sa_events[7][4] , \sa_events[7][3] , 
	\sa_events[7][2] , \sa_events[7][1] , \sa_events[7][0] , 
	\sa_events[6][63] , \sa_events[6][62] , \sa_events[6][61] , 
	\sa_events[6][60] , \sa_events[6][59] , \sa_events[6][58] , 
	\sa_events[6][57] , \sa_events[6][56] , \sa_events[6][55] , 
	\sa_events[6][54] , \sa_events[6][53] , \sa_events[6][52] , 
	\sa_events[6][51] , \sa_events[6][50] , \sa_events[6][49] , 
	\sa_events[6][48] , \sa_events[6][47] , \sa_events[6][46] , 
	\sa_events[6][45] , \sa_events[6][44] , \sa_events[6][43] , 
	\sa_events[6][42] , \sa_events[6][41] , \sa_events[6][40] , 
	\sa_events[6][39] , \sa_events[6][38] , \sa_events[6][37] , 
	\sa_events[6][36] , \sa_events[6][35] , \sa_events[6][34] , 
	\sa_events[6][33] , \sa_events[6][32] , \sa_events[6][31] , 
	\sa_events[6][30] , \sa_events[6][29] , \sa_events[6][28] , 
	\sa_events[6][27] , \sa_events[6][26] , \sa_events[6][25] , 
	\sa_events[6][24] , \sa_events[6][23] , \sa_events[6][22] , 
	\sa_events[6][21] , \sa_events[6][20] , \sa_events[6][19] , 
	\sa_events[6][18] , \sa_events[6][17] , \sa_events[6][16] , 
	\sa_events[6][15] , \sa_events[6][14] , \sa_events[6][13] , 
	\sa_events[6][12] , \sa_events[6][11] , \sa_events[6][10] , 
	\sa_events[6][9] , \sa_events[6][8] , \sa_events[6][7] , 
	\sa_events[6][6] , \sa_events[6][5] , \sa_events[6][4] , 
	\sa_events[6][3] , \sa_events[6][2] , \sa_events[6][1] , 
	\sa_events[6][0] , \sa_events[5][63] , \sa_events[5][62] , 
	\sa_events[5][61] , \sa_events[5][60] , \sa_events[5][59] , 
	\sa_events[5][58] , \sa_events[5][57] , \sa_events[5][56] , 
	\sa_events[5][55] , \sa_events[5][54] , \sa_events[5][53] , 
	\sa_events[5][52] , \sa_events[5][51] , \sa_events[5][50] , 
	\sa_events[5][49] , \sa_events[5][48] , \sa_events[5][47] , 
	\sa_events[5][46] , \sa_events[5][45] , \sa_events[5][44] , 
	\sa_events[5][43] , \sa_events[5][42] , \sa_events[5][41] , 
	\sa_events[5][40] , \sa_events[5][39] , \sa_events[5][38] , 
	\sa_events[5][37] , \sa_events[5][36] , \sa_events[5][35] , 
	\sa_events[5][34] , \sa_events[5][33] , \sa_events[5][32] , 
	\sa_events[5][31] , \sa_events[5][30] , \sa_events[5][29] , 
	\sa_events[5][28] , \sa_events[5][27] , \sa_events[5][26] , 
	\sa_events[5][25] , \sa_events[5][24] , \sa_events[5][23] , 
	\sa_events[5][22] , \sa_events[5][21] , \sa_events[5][20] , 
	\sa_events[5][19] , \sa_events[5][18] , \sa_events[5][17] , 
	\sa_events[5][16] , \sa_events[5][15] , \sa_events[5][14] , 
	\sa_events[5][13] , \sa_events[5][12] , \sa_events[5][11] , 
	\sa_events[5][10] , \sa_events[5][9] , \sa_events[5][8] , 
	\sa_events[5][7] , \sa_events[5][6] , \sa_events[5][5] , 
	\sa_events[5][4] , \sa_events[5][3] , \sa_events[5][2] , 
	\sa_events[5][1] , \sa_events[5][0] , \sa_events[4][63] , 
	\sa_events[4][62] , \sa_events[4][61] , \sa_events[4][60] , 
	\sa_events[4][59] , \sa_events[4][58] , \sa_events[4][57] , 
	\sa_events[4][56] , \sa_events[4][55] , \sa_events[4][54] , 
	\sa_events[4][53] , \sa_events[4][52] , \sa_events[4][51] , 
	\sa_events[4][50] , \sa_events[4][49] , \sa_events[4][48] , 
	\sa_events[4][47] , \sa_events[4][46] , \sa_events[4][45] , 
	\sa_events[4][44] , \sa_events[4][43] , \sa_events[4][42] , 
	\sa_events[4][41] , \sa_events[4][40] , \sa_events[4][39] , 
	\sa_events[4][38] , \sa_events[4][37] , \sa_events[4][36] , 
	\sa_events[4][35] , \sa_events[4][34] , \sa_events[4][33] , 
	\sa_events[4][32] , \sa_events[4][31] , \sa_events[4][30] , 
	\sa_events[4][29] , \sa_events[4][28] , \sa_events[4][27] , 
	\sa_events[4][26] , \sa_events[4][25] , \sa_events[4][24] , 
	\sa_events[4][23] , \sa_events[4][22] , \sa_events[4][21] , 
	\sa_events[4][20] , \sa_events[4][19] , \sa_events[4][18] , 
	\sa_events[4][17] , \sa_events[4][16] , \sa_events[4][15] , 
	\sa_events[4][14] , \sa_events[4][13] , \sa_events[4][12] , 
	\sa_events[4][11] , \sa_events[4][10] , \sa_events[4][9] , 
	\sa_events[4][8] , \sa_events[4][7] , \sa_events[4][6] , 
	\sa_events[4][5] , \sa_events[4][4] , \sa_events[4][3] , 
	\sa_events[4][2] , \sa_events[4][1] , \sa_events[4][0] , 
	\sa_events[3][63] , \sa_events[3][62] , \sa_events[3][61] , 
	\sa_events[3][60] , \sa_events[3][59] , \sa_events[3][58] , 
	\sa_events[3][57] , \sa_events[3][56] , \sa_events[3][55] , 
	\sa_events[3][54] , \sa_events[3][53] , \sa_events[3][52] , 
	\sa_events[3][51] , \sa_events[3][50] , \sa_events[3][49] , 
	\sa_events[3][48] , \sa_events[3][47] , \sa_events[3][46] , 
	\sa_events[3][45] , \sa_events[3][44] , \sa_events[3][43] , 
	\sa_events[3][42] , \sa_events[3][41] , \sa_events[3][40] , 
	\sa_events[3][39] , \sa_events[3][38] , \sa_events[3][37] , 
	\sa_events[3][36] , \sa_events[3][35] , \sa_events[3][34] , 
	\sa_events[3][33] , \sa_events[3][32] , \sa_events[3][31] , 
	\sa_events[3][30] , \sa_events[3][29] , \sa_events[3][28] , 
	\sa_events[3][27] , \sa_events[3][26] , \sa_events[3][25] , 
	\sa_events[3][24] , \sa_events[3][23] , \sa_events[3][22] , 
	\sa_events[3][21] , \sa_events[3][20] , \sa_events[3][19] , 
	\sa_events[3][18] , \sa_events[3][17] , \sa_events[3][16] , 
	\sa_events[3][15] , \sa_events[3][14] , \sa_events[3][13] , 
	\sa_events[3][12] , \sa_events[3][11] , \sa_events[3][10] , 
	\sa_events[3][9] , \sa_events[3][8] , \sa_events[3][7] , 
	\sa_events[3][6] , \sa_events[3][5] , \sa_events[3][4] , 
	\sa_events[3][3] , \sa_events[3][2] , \sa_events[3][1] , 
	\sa_events[3][0] , \sa_events[2][63] , \sa_events[2][62] , 
	\sa_events[2][61] , \sa_events[2][60] , \sa_events[2][59] , 
	\sa_events[2][58] , \sa_events[2][57] , \sa_events[2][56] , 
	\sa_events[2][55] , \sa_events[2][54] , \sa_events[2][53] , 
	\sa_events[2][52] , \sa_events[2][51] , \sa_events[2][50] , 
	\sa_events[2][49] , \sa_events[2][48] , \sa_events[2][47] , 
	\sa_events[2][46] , \sa_events[2][45] , \sa_events[2][44] , 
	\sa_events[2][43] , \sa_events[2][42] , \sa_events[2][41] , 
	\sa_events[2][40] , \sa_events[2][39] , \sa_events[2][38] , 
	\sa_events[2][37] , \sa_events[2][36] , \sa_events[2][35] , 
	\sa_events[2][34] , \sa_events[2][33] , \sa_events[2][32] , 
	\sa_events[2][31] , \sa_events[2][30] , \sa_events[2][29] , 
	\sa_events[2][28] , \sa_events[2][27] , \sa_events[2][26] , 
	\sa_events[2][25] , \sa_events[2][24] , \sa_events[2][23] , 
	\sa_events[2][22] , \sa_events[2][21] , \sa_events[2][20] , 
	\sa_events[2][19] , \sa_events[2][18] , \sa_events[2][17] , 
	\sa_events[2][16] , \sa_events[2][15] , \sa_events[2][14] , 
	\sa_events[2][13] , \sa_events[2][12] , \sa_events[2][11] , 
	\sa_events[2][10] , \sa_events[2][9] , \sa_events[2][8] , 
	\sa_events[2][7] , \sa_events[2][6] , \sa_events[2][5] , 
	\sa_events[2][4] , \sa_events[2][3] , \sa_events[2][2] , 
	\sa_events[2][1] , \sa_events[2][0] , \sa_events[1][63] , 
	\sa_events[1][62] , \sa_events[1][61] , \sa_events[1][60] , 
	\sa_events[1][59] , \sa_events[1][58] , \sa_events[1][57] , 
	\sa_events[1][56] , \sa_events[1][55] , \sa_events[1][54] , 
	\sa_events[1][53] , \sa_events[1][52] , \sa_events[1][51] , 
	\sa_events[1][50] , \sa_events[1][49] , \sa_events[1][48] , 
	\sa_events[1][47] , \sa_events[1][46] , \sa_events[1][45] , 
	\sa_events[1][44] , \sa_events[1][43] , \sa_events[1][42] , 
	\sa_events[1][41] , \sa_events[1][40] , \sa_events[1][39] , 
	\sa_events[1][38] , \sa_events[1][37] , \sa_events[1][36] , 
	\sa_events[1][35] , \sa_events[1][34] , \sa_events[1][33] , 
	\sa_events[1][32] , \sa_events[1][31] , \sa_events[1][30] , 
	\sa_events[1][29] , \sa_events[1][28] , \sa_events[1][27] , 
	\sa_events[1][26] , \sa_events[1][25] , \sa_events[1][24] , 
	\sa_events[1][23] , \sa_events[1][22] , \sa_events[1][21] , 
	\sa_events[1][20] , \sa_events[1][19] , \sa_events[1][18] , 
	\sa_events[1][17] , \sa_events[1][16] , \sa_events[1][15] , 
	\sa_events[1][14] , \sa_events[1][13] , \sa_events[1][12] , 
	\sa_events[1][11] , \sa_events[1][10] , \sa_events[1][9] , 
	\sa_events[1][8] , \sa_events[1][7] , \sa_events[1][6] , 
	\sa_events[1][5] , \sa_events[1][4] , \sa_events[1][3] , 
	\sa_events[1][2] , \sa_events[1][1] , \sa_events[1][0] , 
	\sa_events[0][63] , \sa_events[0][62] , \sa_events[0][61] , 
	\sa_events[0][60] , \sa_events[0][59] , \sa_events[0][58] , 
	\sa_events[0][57] , \sa_events[0][56] , \sa_events[0][55] , 
	\sa_events[0][54] , \sa_events[0][53] , \sa_events[0][52] , 
	\sa_events[0][51] , \sa_events[0][50] , \sa_events[0][49] , 
	\sa_events[0][48] , \sa_events[0][47] , \sa_events[0][46] , 
	\sa_events[0][45] , \sa_events[0][44] , \sa_events[0][43] , 
	\sa_events[0][42] , \sa_events[0][41] , \sa_events[0][40] , 
	\sa_events[0][39] , \sa_events[0][38] , \sa_events[0][37] , 
	\sa_events[0][36] , \sa_events[0][35] , \sa_events[0][34] , 
	\sa_events[0][33] , \sa_events[0][32] , \sa_events[0][31] , 
	\sa_events[0][30] , \sa_events[0][29] , \sa_events[0][28] , 
	\sa_events[0][27] , \sa_events[0][26] , \sa_events[0][25] , 
	\sa_events[0][24] , \sa_events[0][23] , \sa_events[0][22] , 
	\sa_events[0][21] , \sa_events[0][20] , \sa_events[0][19] , 
	\sa_events[0][18] , \sa_events[0][17] , \sa_events[0][16] , 
	\sa_events[0][15] , \sa_events[0][14] , \sa_events[0][13] , 
	\sa_events[0][12] , \sa_events[0][11] , \sa_events[0][10] , 
	\sa_events[0][9] , \sa_events[0][8] , \sa_events[0][7] , 
	\sa_events[0][6] , \sa_events[0][5] , \sa_events[0][4] , 
	\sa_events[0][3] , \sa_events[0][2] , \sa_events[0][1] , 
	\sa_events[0][0] }), .sa_clear( 
	\num_31_._zy_simnet_sa_clear_163_w$ ), .sa_snap( 
	\num_31_._zy_simnet_sa_snap_164_w$ ));
ixc_assign \num_31_._zz_strnp_159 ( \num_31_._zy_simnet_sa_snap_164_w$ , 
	sa_snap);
ixc_assign \num_31_._zz_strnp_158 ( \num_31_._zy_simnet_sa_clear_163_w$ , 
	sa_clear);
ixc_assign_50 \num_31_._zz_strnp_156 ( { \sa_snapshot[31][49] , 
	\sa_snapshot[31][48] , \sa_snapshot[31][47] , \sa_snapshot[31][46] , 
	\sa_snapshot[31][45] , \sa_snapshot[31][44] , \sa_snapshot[31][43] , 
	\sa_snapshot[31][42] , \sa_snapshot[31][41] , \sa_snapshot[31][40] , 
	\sa_snapshot[31][39] , \sa_snapshot[31][38] , \sa_snapshot[31][37] , 
	\sa_snapshot[31][36] , \sa_snapshot[31][35] , \sa_snapshot[31][34] , 
	\sa_snapshot[31][33] , \sa_snapshot[31][32] , \sa_snapshot[31][31] , 
	\sa_snapshot[31][30] , \sa_snapshot[31][29] , \sa_snapshot[31][28] , 
	\sa_snapshot[31][27] , \sa_snapshot[31][26] , \sa_snapshot[31][25] , 
	\sa_snapshot[31][24] , \sa_snapshot[31][23] , \sa_snapshot[31][22] , 
	\sa_snapshot[31][21] , \sa_snapshot[31][20] , \sa_snapshot[31][19] , 
	\sa_snapshot[31][18] , \sa_snapshot[31][17] , \sa_snapshot[31][16] , 
	\sa_snapshot[31][15] , \sa_snapshot[31][14] , \sa_snapshot[31][13] , 
	\sa_snapshot[31][12] , \sa_snapshot[31][11] , \sa_snapshot[31][10] , 
	\sa_snapshot[31][9] , \sa_snapshot[31][8] , \sa_snapshot[31][7] , 
	\sa_snapshot[31][6] , \sa_snapshot[31][5] , \sa_snapshot[31][4] , 
	\sa_snapshot[31][3] , \sa_snapshot[31][2] , \sa_snapshot[31][1] , 
	\sa_snapshot[31][0] }, \num_31_._zy_simnet_tvar_161 [0:49]);
ixc_assign_50 \num_31_._zz_strnp_155 ( { \sa_count[31][49] , 
	\sa_count[31][48] , \sa_count[31][47] , \sa_count[31][46] , 
	\sa_count[31][45] , \sa_count[31][44] , \sa_count[31][43] , 
	\sa_count[31][42] , \sa_count[31][41] , \sa_count[31][40] , 
	\sa_count[31][39] , \sa_count[31][38] , \sa_count[31][37] , 
	\sa_count[31][36] , \sa_count[31][35] , \sa_count[31][34] , 
	\sa_count[31][33] , \sa_count[31][32] , \sa_count[31][31] , 
	\sa_count[31][30] , \sa_count[31][29] , \sa_count[31][28] , 
	\sa_count[31][27] , \sa_count[31][26] , \sa_count[31][25] , 
	\sa_count[31][24] , \sa_count[31][23] , \sa_count[31][22] , 
	\sa_count[31][21] , \sa_count[31][20] , \sa_count[31][19] , 
	\sa_count[31][18] , \sa_count[31][17] , \sa_count[31][16] , 
	\sa_count[31][15] , \sa_count[31][14] , \sa_count[31][13] , 
	\sa_count[31][12] , \sa_count[31][11] , \sa_count[31][10] , 
	\sa_count[31][9] , \sa_count[31][8] , \sa_count[31][7] , 
	\sa_count[31][6] , \sa_count[31][5] , \sa_count[31][4] , 
	\sa_count[31][3] , \sa_count[31][2] , \sa_count[31][1] , 
	\sa_count[31][0] }, \num_31_._zy_simnet_tvar_160 [0:49]);
Q_INV U2187 ( .A(num_key_tlv_in_flight[0]), .Z(n241));
Q_FDP4EP \num_key_tlv_in_flight_REG[0] ( .CK(clk), .CE(n72), .R(n242), .D(n241), .Q(num_key_tlv_in_flight[0]));
Q_INV U2189 ( .A(rst_n), .Z(n242));
Q_FDP4EP \num_key_tlv_in_flight_REG[1] ( .CK(clk), .CE(n72), .R(n242), .D(n26), .Q(num_key_tlv_in_flight[1]));
Q_FDP4EP \num_key_tlv_in_flight_REG[2] ( .CK(clk), .CE(n72), .R(n242), .D(n27), .Q(num_key_tlv_in_flight[2]));
Q_FDP4EP \num_key_tlv_in_flight_REG[3] ( .CK(clk), .CE(n72), .R(n242), .D(n29), .Q(num_key_tlv_in_flight[3]));
Q_FDP4EP \num_key_tlv_in_flight_REG[4] ( .CK(clk), .CE(n72), .R(n242), .D(n30), .Q(num_key_tlv_in_flight[4]));
Q_FDP4EP \num_key_tlv_in_flight_REG[5] ( .CK(clk), .CE(n72), .R(n242), .D(n32), .Q(num_key_tlv_in_flight[5]));
Q_FDP4EP \num_key_tlv_in_flight_REG[6] ( .CK(clk), .CE(n72), .R(n242), .D(n33), .Q(num_key_tlv_in_flight[6]));
Q_FDP4EP \num_key_tlv_in_flight_REG[7] ( .CK(clk), .CE(n72), .R(n242), .D(n35), .Q(num_key_tlv_in_flight[7]));
Q_FDP4EP \num_key_tlv_in_flight_REG[8] ( .CK(clk), .CE(n72), .R(n242), .D(n36), .Q(num_key_tlv_in_flight[8]));
Q_FDP4EP \num_key_tlv_in_flight_REG[9] ( .CK(clk), .CE(n72), .R(n242), .D(n38), .Q(num_key_tlv_in_flight[9]));
Q_FDP4EP \num_key_tlv_in_flight_REG[10] ( .CK(clk), .CE(n72), .R(n242), .D(n39), .Q(num_key_tlv_in_flight[10]));
Q_FDP4EP \num_key_tlv_in_flight_REG[11] ( .CK(clk), .CE(n72), .R(n242), .D(n41), .Q(num_key_tlv_in_flight[11]));
Q_FDP4EP \num_key_tlv_in_flight_REG[12] ( .CK(clk), .CE(n72), .R(n242), .D(n42), .Q(num_key_tlv_in_flight[12]));
Q_FDP4EP \num_key_tlv_in_flight_REG[13] ( .CK(clk), .CE(n72), .R(n242), .D(n44), .Q(num_key_tlv_in_flight[13]));
Q_FDP4EP \num_key_tlv_in_flight_REG[14] ( .CK(clk), .CE(n72), .R(n242), .D(n45), .Q(num_key_tlv_in_flight[14]));
Q_FDP4EP \num_key_tlv_in_flight_REG[15] ( .CK(clk), .CE(n72), .R(n242), .D(n47), .Q(num_key_tlv_in_flight[15]));
Q_FDP4EP \num_key_tlv_in_flight_REG[16] ( .CK(clk), .CE(n72), .R(n242), .D(n48), .Q(num_key_tlv_in_flight[16]));
Q_FDP4EP \num_key_tlv_in_flight_REG[17] ( .CK(clk), .CE(n72), .R(n242), .D(n50), .Q(num_key_tlv_in_flight[17]));
Q_FDP4EP \num_key_tlv_in_flight_REG[18] ( .CK(clk), .CE(n72), .R(n242), .D(n51), .Q(num_key_tlv_in_flight[18]));
Q_FDP4EP \num_key_tlv_in_flight_REG[19] ( .CK(clk), .CE(n72), .R(n242), .D(n53), .Q(num_key_tlv_in_flight[19]));
Q_FDP4EP \num_key_tlv_in_flight_REG[20] ( .CK(clk), .CE(n72), .R(n242), .D(n54), .Q(num_key_tlv_in_flight[20]));
Q_FDP4EP \num_key_tlv_in_flight_REG[21] ( .CK(clk), .CE(n72), .R(n242), .D(n56), .Q(num_key_tlv_in_flight[21]));
Q_FDP4EP \num_key_tlv_in_flight_REG[22] ( .CK(clk), .CE(n72), .R(n242), .D(n57), .Q(num_key_tlv_in_flight[22]));
Q_FDP4EP \num_key_tlv_in_flight_REG[23] ( .CK(clk), .CE(n72), .R(n242), .D(n59), .Q(num_key_tlv_in_flight[23]));
Q_FDP4EP \num_key_tlv_in_flight_REG[24] ( .CK(clk), .CE(n72), .R(n242), .D(n60), .Q(num_key_tlv_in_flight[24]));
Q_FDP4EP \num_key_tlv_in_flight_REG[25] ( .CK(clk), .CE(n72), .R(n242), .D(n62), .Q(num_key_tlv_in_flight[25]));
Q_FDP4EP \num_key_tlv_in_flight_REG[26] ( .CK(clk), .CE(n72), .R(n242), .D(n63), .Q(num_key_tlv_in_flight[26]));
Q_FDP4EP \num_key_tlv_in_flight_REG[27] ( .CK(clk), .CE(n72), .R(n242), .D(n65), .Q(num_key_tlv_in_flight[27]));
Q_FDP4EP \num_key_tlv_in_flight_REG[28] ( .CK(clk), .CE(n72), .R(n242), .D(n66), .Q(num_key_tlv_in_flight[28]));
Q_FDP4EP \num_key_tlv_in_flight_REG[29] ( .CK(clk), .CE(n72), .R(n242), .D(n68), .Q(num_key_tlv_in_flight[29]));
Q_FDP4EP \num_key_tlv_in_flight_REG[30] ( .CK(clk), .CE(n72), .R(n242), .D(n69), .Q(num_key_tlv_in_flight[30]));
Q_FDP4EP \num_key_tlv_in_flight_REG[31] ( .CK(clk), .CE(n72), .R(n242), .D(n71), .Q(num_key_tlv_in_flight[31]));
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m1 "sa_snapshot 1 63 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m2 "sa_count 1 63 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_DECL_m3 "sa_events 1 63 0 15 0"
// pragma CVASTRPROP MODULE HDLICE HDL_MEMORY_NON_CMM "3"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\sa_snapshot%s.r.part1  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\sa_snapshot%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\sa_snapshot%s.f.unused  1 13 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\sa_snapshot%s.f.upper  1 17 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\sa_snapshot%s.f.lower  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\sa_count%s.r.part1  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\sa_count%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\sa_count%s.f.unused  1 13 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\sa_count%s.f.upper  1 17 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\sa_count%s.f.lower  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\idle_components.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\idle_components.f.num_key_tlvs_in_flight  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\tready_override.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\sa_global_ctrl.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\sa_global_ctrl.f.spare  (1,0) 1 29 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\sa_ctrl%s.r.part0  1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\sa_ctrl%s.f.spare  1 26 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\sa_ctrl%s.f.sa_event_sel  1 4 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "sa_ctrl 1 31 0 31 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "19"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "kme_ib_out 1 \kme_ib_out.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r1 "sa_snapshot%s 2 \sa_snapshot%s.r  { \sa_snapshot%s.r.part1  \sa_snapshot%s.r.part0  } \sa_snapshot%s.f  { \sa_snapshot%s.f.unused  \sa_snapshot%s.f.upper  \sa_snapshot%s.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r2 "sa_count%s 2 \sa_count%s.r  { \sa_count%s.r.part1  \sa_count%s.r.part0  } \sa_count%s.f  { \sa_count%s.f.unused  \sa_count%s.f.upper  \sa_count%s.f.lower  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r3 "idle_components 2 \idle_components.r  { \idle_components.r.part0  } \idle_components.f  { \idle_components.f.num_key_tlvs_in_flight  \idle_components.f.cddip0_key_tlv_rsm_idle  \idle_components.f.cddip1_key_tlv_rsm_idle  \idle_components.f.cddip2_key_tlv_rsm_idle  \idle_components.f.cddip3_key_tlv_rsm_idle  \idle_components.f.cceip0_key_tlv_rsm_idle  \idle_components.f.cceip1_key_tlv_rsm_idle  \idle_components.f.cceip2_key_tlv_rsm_idle  \idle_components.f.cceip3_key_tlv_rsm_idle  \idle_components.f.no_key_tlv_in_flight  \idle_components.f.tlv_parser_idle  \idle_components.f.drng_idle  \idle_components.f.kme_slv_empty  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r4 "tready_override 2 \tready_override.r  { \tready_override.r.part0  } \tready_override.f  { \tready_override.f.txc_tready_override  \tready_override.f.engine_7_tready_override  \tready_override.f.engine_6_tready_override  \tready_override.f.engine_5_tready_override  \tready_override.f.engine_4_tready_override  \tready_override.f.engine_3_tready_override  \tready_override.f.engine_2_tready_override  \tready_override.f.engine_1_tready_override  \tready_override.f.engine_0_tready_override  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "core_kme_ib_out 1 \core_kme_ib_out.tready "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r5 "sa_global_ctrl 2 \sa_global_ctrl.r  { \sa_global_ctrl.r.part0  } \sa_global_ctrl.f  { \sa_global_ctrl.f.spare  \sa_global_ctrl.f.sa_snap  \sa_global_ctrl.f.sa_clear_live  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r6 "sa_ctrl%s 2 \sa_ctrl%s.r  { \sa_ctrl%s.r.part0  } \sa_ctrl%s.f  { \sa_ctrl%s.f.spare  \sa_ctrl%s.f.sa_event_sel  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "2"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_NUM "6"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 num 0 31 "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[31]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[30]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[29]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[28]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[27]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[26]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[25]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[24]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[23]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[22]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[21]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[20]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[19]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[18]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[17]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[16]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[15]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[14]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[13]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[12]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[11]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[10]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[9]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[8]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[7]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[6]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[5]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[4]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[3]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[2]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[1]"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "num[0]"
endmodule
