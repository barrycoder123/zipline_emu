library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
use work.cr_kme_regfilePKG.all ;
entity kme_tb is
  attribute _2_state_: integer;
end kme_tb ;
