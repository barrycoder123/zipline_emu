
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_upsizer_x2_xcm72 ( upsizer_in_stall, upsizer_out_valid, 
	upsizer_out_eof, upsizer_out_data, clk, rst_n, in_upsizer_valid, 
	in_upsizer_eof, in_upsizer_data, out_upsizer_stall);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output upsizer_in_stall;
output upsizer_out_valid;
output upsizer_out_eof;
output [127:0] upsizer_out_data;
input clk;
input rst_n;
input in_upsizer_valid;
input in_upsizer_eof;
input [63:0] in_upsizer_data;
input out_upsizer_stall;
wire _zy_simnet_upsizer_in_stall_0_w$;
wire _zy_simnet_upsizer_out_valid_1_w$;
wire _zy_simnet_upsizer_out_eof_2_w$;
wire [0:127] _zy_simnet_upsizer_out_data_3_w$;
wire send_data;
wire [63:0] buffer;
Q_BUF U0 ( .A(out_upsizer_stall), .Z(upsizer_in_stall));
ixc_assign_128 _zz_strnp_3 ( _zy_simnet_upsizer_out_data_3_w$[0:127], 
	upsizer_out_data[127:0]);
ixc_assign _zz_strnp_2 ( _zy_simnet_upsizer_out_eof_2_w$, upsizer_out_eof);
ixc_assign _zz_strnp_1 ( _zy_simnet_upsizer_out_valid_1_w$, upsizer_out_valid);
ixc_assign _zz_strnp_0 ( _zy_simnet_upsizer_in_stall_0_w$, out_upsizer_stall);
Q_AN02 U5 ( .A0(n1), .A1(in_upsizer_valid), .Z(n2));
Q_AN02 U6 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[0]), .Z(upsizer_out_data[0]));
Q_AN02 U7 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[1]), .Z(upsizer_out_data[1]));
Q_AN02 U8 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[2]), .Z(upsizer_out_data[2]));
Q_AN02 U9 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[3]), .Z(upsizer_out_data[3]));
Q_AN02 U10 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[4]), .Z(upsizer_out_data[4]));
Q_AN02 U11 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[5]), .Z(upsizer_out_data[5]));
Q_AN02 U12 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[6]), .Z(upsizer_out_data[6]));
Q_AN02 U13 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[7]), .Z(upsizer_out_data[7]));
Q_AN02 U14 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[8]), .Z(upsizer_out_data[8]));
Q_AN02 U15 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[9]), .Z(upsizer_out_data[9]));
Q_AN02 U16 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[10]), .Z(upsizer_out_data[10]));
Q_AN02 U17 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[11]), .Z(upsizer_out_data[11]));
Q_AN02 U18 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[12]), .Z(upsizer_out_data[12]));
Q_AN02 U19 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[13]), .Z(upsizer_out_data[13]));
Q_AN02 U20 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[14]), .Z(upsizer_out_data[14]));
Q_AN02 U21 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[15]), .Z(upsizer_out_data[15]));
Q_AN02 U22 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[16]), .Z(upsizer_out_data[16]));
Q_AN02 U23 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[17]), .Z(upsizer_out_data[17]));
Q_AN02 U24 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[18]), .Z(upsizer_out_data[18]));
Q_AN02 U25 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[19]), .Z(upsizer_out_data[19]));
Q_AN02 U26 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[20]), .Z(upsizer_out_data[20]));
Q_AN02 U27 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[21]), .Z(upsizer_out_data[21]));
Q_AN02 U28 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[22]), .Z(upsizer_out_data[22]));
Q_AN02 U29 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[23]), .Z(upsizer_out_data[23]));
Q_AN02 U30 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[24]), .Z(upsizer_out_data[24]));
Q_AN02 U31 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[25]), .Z(upsizer_out_data[25]));
Q_AN02 U32 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[26]), .Z(upsizer_out_data[26]));
Q_AN02 U33 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[27]), .Z(upsizer_out_data[27]));
Q_AN02 U34 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[28]), .Z(upsizer_out_data[28]));
Q_AN02 U35 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[29]), .Z(upsizer_out_data[29]));
Q_AN02 U36 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[30]), .Z(upsizer_out_data[30]));
Q_AN02 U37 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[31]), .Z(upsizer_out_data[31]));
Q_AN02 U38 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[32]), .Z(upsizer_out_data[32]));
Q_AN02 U39 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[33]), .Z(upsizer_out_data[33]));
Q_AN02 U40 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[34]), .Z(upsizer_out_data[34]));
Q_AN02 U41 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[35]), .Z(upsizer_out_data[35]));
Q_AN02 U42 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[36]), .Z(upsizer_out_data[36]));
Q_AN02 U43 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[37]), .Z(upsizer_out_data[37]));
Q_AN02 U44 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[38]), .Z(upsizer_out_data[38]));
Q_AN02 U45 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[39]), .Z(upsizer_out_data[39]));
Q_AN02 U46 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[40]), .Z(upsizer_out_data[40]));
Q_AN02 U47 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[41]), .Z(upsizer_out_data[41]));
Q_AN02 U48 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[42]), .Z(upsizer_out_data[42]));
Q_AN02 U49 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[43]), .Z(upsizer_out_data[43]));
Q_AN02 U50 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[44]), .Z(upsizer_out_data[44]));
Q_AN02 U51 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[45]), .Z(upsizer_out_data[45]));
Q_AN02 U52 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[46]), .Z(upsizer_out_data[46]));
Q_AN02 U53 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[47]), .Z(upsizer_out_data[47]));
Q_AN02 U54 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[48]), .Z(upsizer_out_data[48]));
Q_AN02 U55 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[49]), .Z(upsizer_out_data[49]));
Q_AN02 U56 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[50]), .Z(upsizer_out_data[50]));
Q_AN02 U57 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[51]), .Z(upsizer_out_data[51]));
Q_AN02 U58 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[52]), .Z(upsizer_out_data[52]));
Q_AN02 U59 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[53]), .Z(upsizer_out_data[53]));
Q_AN02 U60 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[54]), .Z(upsizer_out_data[54]));
Q_AN02 U61 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[55]), .Z(upsizer_out_data[55]));
Q_AN02 U62 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[56]), .Z(upsizer_out_data[56]));
Q_AN02 U63 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[57]), .Z(upsizer_out_data[57]));
Q_AN02 U64 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[58]), .Z(upsizer_out_data[58]));
Q_AN02 U65 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[59]), .Z(upsizer_out_data[59]));
Q_AN02 U66 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[60]), .Z(upsizer_out_data[60]));
Q_AN02 U67 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[61]), .Z(upsizer_out_data[61]));
Q_AN02 U68 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[62]), .Z(upsizer_out_data[62]));
Q_AN02 U69 ( .A0(upsizer_out_valid), .A1(in_upsizer_data[63]), .Z(upsizer_out_data[63]));
Q_AN02 U70 ( .A0(upsizer_out_valid), .A1(buffer[0]), .Z(upsizer_out_data[64]));
Q_AN02 U71 ( .A0(upsizer_out_valid), .A1(buffer[1]), .Z(upsizer_out_data[65]));
Q_AN02 U72 ( .A0(upsizer_out_valid), .A1(buffer[2]), .Z(upsizer_out_data[66]));
Q_AN02 U73 ( .A0(upsizer_out_valid), .A1(buffer[3]), .Z(upsizer_out_data[67]));
Q_AN02 U74 ( .A0(upsizer_out_valid), .A1(buffer[4]), .Z(upsizer_out_data[68]));
Q_AN02 U75 ( .A0(upsizer_out_valid), .A1(buffer[5]), .Z(upsizer_out_data[69]));
Q_AN02 U76 ( .A0(upsizer_out_valid), .A1(buffer[6]), .Z(upsizer_out_data[70]));
Q_AN02 U77 ( .A0(upsizer_out_valid), .A1(buffer[7]), .Z(upsizer_out_data[71]));
Q_AN02 U78 ( .A0(upsizer_out_valid), .A1(buffer[8]), .Z(upsizer_out_data[72]));
Q_AN02 U79 ( .A0(upsizer_out_valid), .A1(buffer[9]), .Z(upsizer_out_data[73]));
Q_AN02 U80 ( .A0(upsizer_out_valid), .A1(buffer[10]), .Z(upsizer_out_data[74]));
Q_AN02 U81 ( .A0(upsizer_out_valid), .A1(buffer[11]), .Z(upsizer_out_data[75]));
Q_AN02 U82 ( .A0(upsizer_out_valid), .A1(buffer[12]), .Z(upsizer_out_data[76]));
Q_AN02 U83 ( .A0(upsizer_out_valid), .A1(buffer[13]), .Z(upsizer_out_data[77]));
Q_AN02 U84 ( .A0(upsizer_out_valid), .A1(buffer[14]), .Z(upsizer_out_data[78]));
Q_AN02 U85 ( .A0(upsizer_out_valid), .A1(buffer[15]), .Z(upsizer_out_data[79]));
Q_AN02 U86 ( .A0(upsizer_out_valid), .A1(buffer[16]), .Z(upsizer_out_data[80]));
Q_AN02 U87 ( .A0(upsizer_out_valid), .A1(buffer[17]), .Z(upsizer_out_data[81]));
Q_AN02 U88 ( .A0(upsizer_out_valid), .A1(buffer[18]), .Z(upsizer_out_data[82]));
Q_AN02 U89 ( .A0(upsizer_out_valid), .A1(buffer[19]), .Z(upsizer_out_data[83]));
Q_AN02 U90 ( .A0(upsizer_out_valid), .A1(buffer[20]), .Z(upsizer_out_data[84]));
Q_AN02 U91 ( .A0(upsizer_out_valid), .A1(buffer[21]), .Z(upsizer_out_data[85]));
Q_AN02 U92 ( .A0(upsizer_out_valid), .A1(buffer[22]), .Z(upsizer_out_data[86]));
Q_AN02 U93 ( .A0(upsizer_out_valid), .A1(buffer[23]), .Z(upsizer_out_data[87]));
Q_AN02 U94 ( .A0(upsizer_out_valid), .A1(buffer[24]), .Z(upsizer_out_data[88]));
Q_AN02 U95 ( .A0(upsizer_out_valid), .A1(buffer[25]), .Z(upsizer_out_data[89]));
Q_AN02 U96 ( .A0(upsizer_out_valid), .A1(buffer[26]), .Z(upsizer_out_data[90]));
Q_AN02 U97 ( .A0(upsizer_out_valid), .A1(buffer[27]), .Z(upsizer_out_data[91]));
Q_AN02 U98 ( .A0(upsizer_out_valid), .A1(buffer[28]), .Z(upsizer_out_data[92]));
Q_AN02 U99 ( .A0(upsizer_out_valid), .A1(buffer[29]), .Z(upsizer_out_data[93]));
Q_AN02 U100 ( .A0(upsizer_out_valid), .A1(buffer[30]), .Z(upsizer_out_data[94]));
Q_AN02 U101 ( .A0(upsizer_out_valid), .A1(buffer[31]), .Z(upsizer_out_data[95]));
Q_AN02 U102 ( .A0(upsizer_out_valid), .A1(buffer[32]), .Z(upsizer_out_data[96]));
Q_AN02 U103 ( .A0(upsizer_out_valid), .A1(buffer[33]), .Z(upsizer_out_data[97]));
Q_AN02 U104 ( .A0(upsizer_out_valid), .A1(buffer[34]), .Z(upsizer_out_data[98]));
Q_AN02 U105 ( .A0(upsizer_out_valid), .A1(buffer[35]), .Z(upsizer_out_data[99]));
Q_AN02 U106 ( .A0(upsizer_out_valid), .A1(buffer[36]), .Z(upsizer_out_data[100]));
Q_AN02 U107 ( .A0(upsizer_out_valid), .A1(buffer[37]), .Z(upsizer_out_data[101]));
Q_AN02 U108 ( .A0(upsizer_out_valid), .A1(buffer[38]), .Z(upsizer_out_data[102]));
Q_AN02 U109 ( .A0(upsizer_out_valid), .A1(buffer[39]), .Z(upsizer_out_data[103]));
Q_AN02 U110 ( .A0(upsizer_out_valid), .A1(buffer[40]), .Z(upsizer_out_data[104]));
Q_AN02 U111 ( .A0(upsizer_out_valid), .A1(buffer[41]), .Z(upsizer_out_data[105]));
Q_AN02 U112 ( .A0(upsizer_out_valid), .A1(buffer[42]), .Z(upsizer_out_data[106]));
Q_AN02 U113 ( .A0(upsizer_out_valid), .A1(buffer[43]), .Z(upsizer_out_data[107]));
Q_AN02 U114 ( .A0(upsizer_out_valid), .A1(buffer[44]), .Z(upsizer_out_data[108]));
Q_AN02 U115 ( .A0(upsizer_out_valid), .A1(buffer[45]), .Z(upsizer_out_data[109]));
Q_AN02 U116 ( .A0(upsizer_out_valid), .A1(buffer[46]), .Z(upsizer_out_data[110]));
Q_AN02 U117 ( .A0(upsizer_out_valid), .A1(buffer[47]), .Z(upsizer_out_data[111]));
Q_AN02 U118 ( .A0(upsizer_out_valid), .A1(buffer[48]), .Z(upsizer_out_data[112]));
Q_AN02 U119 ( .A0(upsizer_out_valid), .A1(buffer[49]), .Z(upsizer_out_data[113]));
Q_AN02 U120 ( .A0(upsizer_out_valid), .A1(buffer[50]), .Z(upsizer_out_data[114]));
Q_AN02 U121 ( .A0(upsizer_out_valid), .A1(buffer[51]), .Z(upsizer_out_data[115]));
Q_AN02 U122 ( .A0(upsizer_out_valid), .A1(buffer[52]), .Z(upsizer_out_data[116]));
Q_AN02 U123 ( .A0(upsizer_out_valid), .A1(buffer[53]), .Z(upsizer_out_data[117]));
Q_AN02 U124 ( .A0(upsizer_out_valid), .A1(buffer[54]), .Z(upsizer_out_data[118]));
Q_AN02 U125 ( .A0(upsizer_out_valid), .A1(buffer[55]), .Z(upsizer_out_data[119]));
Q_AN02 U126 ( .A0(upsizer_out_valid), .A1(buffer[56]), .Z(upsizer_out_data[120]));
Q_AN02 U127 ( .A0(upsizer_out_valid), .A1(buffer[57]), .Z(upsizer_out_data[121]));
Q_AN02 U128 ( .A0(upsizer_out_valid), .A1(buffer[58]), .Z(upsizer_out_data[122]));
Q_AN02 U129 ( .A0(upsizer_out_valid), .A1(buffer[59]), .Z(upsizer_out_data[123]));
Q_AN02 U130 ( .A0(upsizer_out_valid), .A1(buffer[60]), .Z(upsizer_out_data[124]));
Q_AN02 U131 ( .A0(upsizer_out_valid), .A1(buffer[61]), .Z(upsizer_out_data[125]));
Q_AN02 U132 ( .A0(upsizer_out_valid), .A1(buffer[62]), .Z(upsizer_out_data[126]));
Q_AN02 U133 ( .A0(upsizer_out_valid), .A1(buffer[63]), .Z(upsizer_out_data[127]));
Q_AN02 U134 ( .A0(upsizer_out_valid), .A1(in_upsizer_eof), .Z(upsizer_out_eof));
Q_AN03 U135 ( .A0(n3), .A1(send_data), .A2(in_upsizer_valid), .Z(upsizer_out_valid));
Q_INV U136 ( .A(out_upsizer_stall), .Z(n3));
Q_FDP4EP send_data_REG  ( .CK(clk), .CE(in_upsizer_valid), .R(n4), .D(n1), .Q(send_data));
Q_INV U138 ( .A(rst_n), .Z(n4));
Q_INV U139 ( .A(send_data), .Z(n1));
Q_FDP4EP \buffer_REG[0] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[0]), .Q(buffer[0]));
Q_FDP4EP \buffer_REG[1] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[1]), .Q(buffer[1]));
Q_FDP4EP \buffer_REG[2] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[2]), .Q(buffer[2]));
Q_FDP4EP \buffer_REG[3] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[3]), .Q(buffer[3]));
Q_FDP4EP \buffer_REG[4] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[4]), .Q(buffer[4]));
Q_FDP4EP \buffer_REG[5] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[5]), .Q(buffer[5]));
Q_FDP4EP \buffer_REG[6] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[6]), .Q(buffer[6]));
Q_FDP4EP \buffer_REG[7] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[7]), .Q(buffer[7]));
Q_FDP4EP \buffer_REG[8] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[8]), .Q(buffer[8]));
Q_FDP4EP \buffer_REG[9] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[9]), .Q(buffer[9]));
Q_FDP4EP \buffer_REG[10] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[10]), .Q(buffer[10]));
Q_FDP4EP \buffer_REG[11] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[11]), .Q(buffer[11]));
Q_FDP4EP \buffer_REG[12] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[12]), .Q(buffer[12]));
Q_FDP4EP \buffer_REG[13] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[13]), .Q(buffer[13]));
Q_FDP4EP \buffer_REG[14] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[14]), .Q(buffer[14]));
Q_FDP4EP \buffer_REG[15] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[15]), .Q(buffer[15]));
Q_FDP4EP \buffer_REG[16] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[16]), .Q(buffer[16]));
Q_FDP4EP \buffer_REG[17] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[17]), .Q(buffer[17]));
Q_FDP4EP \buffer_REG[18] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[18]), .Q(buffer[18]));
Q_FDP4EP \buffer_REG[19] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[19]), .Q(buffer[19]));
Q_FDP4EP \buffer_REG[20] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[20]), .Q(buffer[20]));
Q_FDP4EP \buffer_REG[21] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[21]), .Q(buffer[21]));
Q_FDP4EP \buffer_REG[22] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[22]), .Q(buffer[22]));
Q_FDP4EP \buffer_REG[23] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[23]), .Q(buffer[23]));
Q_FDP4EP \buffer_REG[24] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[24]), .Q(buffer[24]));
Q_FDP4EP \buffer_REG[25] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[25]), .Q(buffer[25]));
Q_FDP4EP \buffer_REG[26] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[26]), .Q(buffer[26]));
Q_FDP4EP \buffer_REG[27] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[27]), .Q(buffer[27]));
Q_FDP4EP \buffer_REG[28] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[28]), .Q(buffer[28]));
Q_FDP4EP \buffer_REG[29] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[29]), .Q(buffer[29]));
Q_FDP4EP \buffer_REG[30] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[30]), .Q(buffer[30]));
Q_FDP4EP \buffer_REG[31] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[31]), .Q(buffer[31]));
Q_FDP4EP \buffer_REG[32] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[32]), .Q(buffer[32]));
Q_FDP4EP \buffer_REG[33] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[33]), .Q(buffer[33]));
Q_FDP4EP \buffer_REG[34] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[34]), .Q(buffer[34]));
Q_FDP4EP \buffer_REG[35] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[35]), .Q(buffer[35]));
Q_FDP4EP \buffer_REG[36] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[36]), .Q(buffer[36]));
Q_FDP4EP \buffer_REG[37] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[37]), .Q(buffer[37]));
Q_FDP4EP \buffer_REG[38] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[38]), .Q(buffer[38]));
Q_FDP4EP \buffer_REG[39] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[39]), .Q(buffer[39]));
Q_FDP4EP \buffer_REG[40] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[40]), .Q(buffer[40]));
Q_FDP4EP \buffer_REG[41] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[41]), .Q(buffer[41]));
Q_FDP4EP \buffer_REG[42] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[42]), .Q(buffer[42]));
Q_FDP4EP \buffer_REG[43] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[43]), .Q(buffer[43]));
Q_FDP4EP \buffer_REG[44] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[44]), .Q(buffer[44]));
Q_FDP4EP \buffer_REG[45] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[45]), .Q(buffer[45]));
Q_FDP4EP \buffer_REG[46] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[46]), .Q(buffer[46]));
Q_FDP4EP \buffer_REG[47] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[47]), .Q(buffer[47]));
Q_FDP4EP \buffer_REG[48] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[48]), .Q(buffer[48]));
Q_FDP4EP \buffer_REG[49] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[49]), .Q(buffer[49]));
Q_FDP4EP \buffer_REG[50] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[50]), .Q(buffer[50]));
Q_FDP4EP \buffer_REG[51] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[51]), .Q(buffer[51]));
Q_FDP4EP \buffer_REG[52] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[52]), .Q(buffer[52]));
Q_FDP4EP \buffer_REG[53] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[53]), .Q(buffer[53]));
Q_FDP4EP \buffer_REG[54] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[54]), .Q(buffer[54]));
Q_FDP4EP \buffer_REG[55] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[55]), .Q(buffer[55]));
Q_FDP4EP \buffer_REG[56] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[56]), .Q(buffer[56]));
Q_FDP4EP \buffer_REG[57] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[57]), .Q(buffer[57]));
Q_FDP4EP \buffer_REG[58] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[58]), .Q(buffer[58]));
Q_FDP4EP \buffer_REG[59] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[59]), .Q(buffer[59]));
Q_FDP4EP \buffer_REG[60] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[60]), .Q(buffer[60]));
Q_FDP4EP \buffer_REG[61] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[61]), .Q(buffer[61]));
Q_FDP4EP \buffer_REG[62] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[62]), .Q(buffer[62]));
Q_FDP4EP \buffer_REG[63] ( .CK(clk), .CE(n2), .R(n4), .D(in_upsizer_data[63]), .Q(buffer[63]));
endmodule
