
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module ixc_context_read_1024 ( rdata);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input [1023:0] rdata;
supply1 n1;
supply0 n2;
Q_NOT_TOUCH _zzqnthw ( .sig());
`ifdef CBV

reg [511:0] _zymem [0:1];
always @(n2 or rdata[511] or rdata[510] or rdata[509] or rdata[508]
 or rdata[507] or rdata[506] or rdata[505] or rdata[504] or rdata[503] or rdata[502] or rdata[501] or rdata[500]
 or rdata[499] or rdata[498] or rdata[497] or rdata[496] or rdata[495] or rdata[494] or rdata[493] or rdata[492]
 or rdata[491] or rdata[490] or rdata[489] or rdata[488] or rdata[487] or rdata[486] or rdata[485] or rdata[484]
 or rdata[483] or rdata[482] or rdata[481] or rdata[480] or rdata[479] or rdata[478] or rdata[477] or rdata[476]
 or rdata[475] or rdata[474] or rdata[473] or rdata[472] or rdata[471] or rdata[470] or rdata[469] or rdata[468]
 or rdata[467] or rdata[466] or rdata[465] or rdata[464] or rdata[463] or rdata[462] or rdata[461] or rdata[460]
 or rdata[459] or rdata[458] or rdata[457] or rdata[456] or rdata[455] or rdata[454] or rdata[453] or rdata[452]
 or rdata[451] or rdata[450] or rdata[449] or rdata[448] or rdata[447] or rdata[446] or rdata[445] or rdata[444]
 or rdata[443] or rdata[442] or rdata[441] or rdata[440] or rdata[439] or rdata[438] or rdata[437] or rdata[436]
 or rdata[435] or rdata[434] or rdata[433] or rdata[432] or rdata[431] or rdata[430] or rdata[429] or rdata[428]
 or rdata[427] or rdata[426] or rdata[425] or rdata[424] or rdata[423] or rdata[422] or rdata[421] or rdata[420]
 or rdata[419] or rdata[418] or rdata[417] or rdata[416] or rdata[415] or rdata[414] or rdata[413] or rdata[412]
 or rdata[411] or rdata[410] or rdata[409] or rdata[408] or rdata[407] or rdata[406] or rdata[405] or rdata[404]
 or rdata[403] or rdata[402] or rdata[401] or rdata[400] or rdata[399] or rdata[398] or rdata[397] or rdata[396]
 or rdata[395] or rdata[394] or rdata[393] or rdata[392] or rdata[391] or rdata[390] or rdata[389] or rdata[388]
 or rdata[387] or rdata[386] or rdata[385] or rdata[384] or rdata[383] or rdata[382] or rdata[381] or rdata[380]
 or rdata[379] or rdata[378] or rdata[377] or rdata[376] or rdata[375] or rdata[374] or rdata[373] or rdata[372]
 or rdata[371] or rdata[370] or rdata[369] or rdata[368] or rdata[367] or rdata[366] or rdata[365] or rdata[364]
 or rdata[363] or rdata[362] or rdata[361] or rdata[360] or rdata[359] or rdata[358] or rdata[357] or rdata[356]
 or rdata[355] or rdata[354] or rdata[353] or rdata[352] or rdata[351] or rdata[350] or rdata[349] or rdata[348]
 or rdata[347] or rdata[346] or rdata[345] or rdata[344] or rdata[343] or rdata[342] or rdata[341] or rdata[340]
 or rdata[339] or rdata[338] or rdata[337] or rdata[336] or rdata[335] or rdata[334] or rdata[333] or rdata[332]
 or rdata[331] or rdata[330] or rdata[329] or rdata[328] or rdata[327] or rdata[326] or rdata[325] or rdata[324]
 or rdata[323] or rdata[322] or rdata[321] or rdata[320] or rdata[319] or rdata[318] or rdata[317] or rdata[316]
 or rdata[315] or rdata[314] or rdata[313] or rdata[312] or rdata[311] or rdata[310] or rdata[309] or rdata[308]
 or rdata[307] or rdata[306] or rdata[305] or rdata[304] or rdata[303] or rdata[302] or rdata[301] or rdata[300]
 or rdata[299] or rdata[298] or rdata[297] or rdata[296] or rdata[295] or rdata[294] or rdata[293] or rdata[292]
 or rdata[291] or rdata[290] or rdata[289] or rdata[288] or rdata[287] or rdata[286] or rdata[285] or rdata[284]
 or rdata[283] or rdata[282] or rdata[281] or rdata[280] or rdata[279] or rdata[278] or rdata[277] or rdata[276]
 or rdata[275] or rdata[274] or rdata[273] or rdata[272] or rdata[271] or rdata[270] or rdata[269] or rdata[268]
 or rdata[267] or rdata[266] or rdata[265] or rdata[264] or rdata[263] or rdata[262] or rdata[261] or rdata[260]
 or rdata[259] or rdata[258] or rdata[257] or rdata[256] or rdata[255] or rdata[254] or rdata[253] or rdata[252]
 or rdata[251] or rdata[250] or rdata[249] or rdata[248] or rdata[247] or rdata[246] or rdata[245] or rdata[244]
 or rdata[243] or rdata[242] or rdata[241] or rdata[240] or rdata[239] or rdata[238] or rdata[237] or rdata[236]
 or rdata[235] or rdata[234] or rdata[233] or rdata[232] or rdata[231] or rdata[230] or rdata[229] or rdata[228]
 or rdata[227] or rdata[226] or rdata[225] or rdata[224] or rdata[223] or rdata[222] or rdata[221] or rdata[220]
 or rdata[219] or rdata[218] or rdata[217] or rdata[216] or rdata[215] or rdata[214] or rdata[213] or rdata[212]
 or rdata[211] or rdata[210] or rdata[209] or rdata[208] or rdata[207] or rdata[206] or rdata[205] or rdata[204]
 or rdata[203] or rdata[202] or rdata[201] or rdata[200] or rdata[199] or rdata[198] or rdata[197] or rdata[196]
 or rdata[195] or rdata[194] or rdata[193] or rdata[192] or rdata[191] or rdata[190] or rdata[189] or rdata[188]
 or rdata[187] or rdata[186] or rdata[185] or rdata[184] or rdata[183] or rdata[182] or rdata[181] or rdata[180]
 or rdata[179] or rdata[178] or rdata[177] or rdata[176] or rdata[175] or rdata[174] or rdata[173] or rdata[172]
 or rdata[171] or rdata[170] or rdata[169] or rdata[168] or rdata[167] or rdata[166] or rdata[165] or rdata[164]
 or rdata[163] or rdata[162] or rdata[161] or rdata[160] or rdata[159] or rdata[158] or rdata[157] or rdata[156]
 or rdata[155] or rdata[154] or rdata[153] or rdata[152] or rdata[151] or rdata[150] or rdata[149] or rdata[148]
 or rdata[147] or rdata[146] or rdata[145] or rdata[144] or rdata[143] or rdata[142] or rdata[141] or rdata[140]
 or rdata[139] or rdata[138] or rdata[137] or rdata[136] or rdata[135] or rdata[134] or rdata[133] or rdata[132]
 or rdata[131] or rdata[130] or rdata[129] or rdata[128] or rdata[127] or rdata[126] or rdata[125] or rdata[124]
 or rdata[123] or rdata[122] or rdata[121] or rdata[120] or rdata[119] or rdata[118] or rdata[117] or rdata[116]
 or rdata[115] or rdata[114] or rdata[113] or rdata[112] or rdata[111] or rdata[110] or rdata[109] or rdata[108]
 or rdata[107] or rdata[106] or rdata[105] or rdata[104] or rdata[103] or rdata[102] or rdata[101] or rdata[100]
 or rdata[99] or rdata[98] or rdata[97] or rdata[96] or rdata[95] or rdata[94] or rdata[93] or rdata[92]
 or rdata[91] or rdata[90] or rdata[89] or rdata[88] or rdata[87] or rdata[86] or rdata[85] or rdata[84]
 or rdata[83] or rdata[82] or rdata[81] or rdata[80] or rdata[79] or rdata[78] or rdata[77] or rdata[76]
 or rdata[75] or rdata[74] or rdata[73] or rdata[72] or rdata[71] or rdata[70] or rdata[69] or rdata[68]
 or rdata[67] or rdata[66] or rdata[65] or rdata[64] or rdata[63] or rdata[62] or rdata[61] or rdata[60]
 or rdata[59] or rdata[58] or rdata[57] or rdata[56] or rdata[55] or rdata[54] or rdata[53] or rdata[52]
 or rdata[51] or rdata[50] or rdata[49] or rdata[48] or rdata[47] or rdata[46] or rdata[45] or rdata[44]
 or rdata[43] or rdata[42] or rdata[41] or rdata[40] or rdata[39] or rdata[38] or rdata[37] or rdata[36]
 or rdata[35] or rdata[34] or rdata[33] or rdata[32] or rdata[31] or rdata[30] or rdata[29] or rdata[28]
 or rdata[27] or rdata[26] or rdata[25] or rdata[24] or rdata[23] or rdata[22] or rdata[21] or rdata[20]
 or rdata[19] or rdata[18] or rdata[17] or rdata[16] or rdata[15] or rdata[14] or rdata[13] or rdata[12]
 or rdata[11] or rdata[10] or rdata[9] or rdata[8] or rdata[7] or rdata[6] or rdata[5] or rdata[4]
 or rdata[3] or rdata[2] or rdata[1] or rdata[0] or n1 or rdata[1023] or rdata[1022] or rdata[1021]
 or rdata[1020] or rdata[1019] or rdata[1018] or rdata[1017] or rdata[1016] or rdata[1015] or rdata[1014] or rdata[1013]
 or rdata[1012] or rdata[1011] or rdata[1010] or rdata[1009] or rdata[1008] or rdata[1007] or rdata[1006] or rdata[1005]
 or rdata[1004] or rdata[1003] or rdata[1002] or rdata[1001] or rdata[1000] or rdata[999] or rdata[998] or rdata[997]
 or rdata[996] or rdata[995] or rdata[994] or rdata[993] or rdata[992] or rdata[991] or rdata[990] or rdata[989]
 or rdata[988] or rdata[987] or rdata[986] or rdata[985] or rdata[984] or rdata[983] or rdata[982] or rdata[981]
 or rdata[980] or rdata[979] or rdata[978] or rdata[977] or rdata[976] or rdata[975] or rdata[974] or rdata[973]
 or rdata[972] or rdata[971] or rdata[970] or rdata[969] or rdata[968] or rdata[967] or rdata[966] or rdata[965]
 or rdata[964] or rdata[963] or rdata[962] or rdata[961] or rdata[960] or rdata[959] or rdata[958] or rdata[957]
 or rdata[956] or rdata[955] or rdata[954] or rdata[953] or rdata[952] or rdata[951] or rdata[950] or rdata[949]
 or rdata[948] or rdata[947] or rdata[946] or rdata[945] or rdata[944] or rdata[943] or rdata[942] or rdata[941]
 or rdata[940] or rdata[939] or rdata[938] or rdata[937] or rdata[936] or rdata[935] or rdata[934] or rdata[933]
 or rdata[932] or rdata[931] or rdata[930] or rdata[929] or rdata[928] or rdata[927] or rdata[926] or rdata[925]
 or rdata[924] or rdata[923] or rdata[922] or rdata[921] or rdata[920] or rdata[919] or rdata[918] or rdata[917]
 or rdata[916] or rdata[915] or rdata[914] or rdata[913] or rdata[912] or rdata[911] or rdata[910] or rdata[909]
 or rdata[908] or rdata[907] or rdata[906] or rdata[905] or rdata[904] or rdata[903] or rdata[902] or rdata[901]
 or rdata[900] or rdata[899] or rdata[898] or rdata[897] or rdata[896] or rdata[895] or rdata[894] or rdata[893]
 or rdata[892] or rdata[891] or rdata[890] or rdata[889] or rdata[888] or rdata[887] or rdata[886] or rdata[885]
 or rdata[884] or rdata[883] or rdata[882] or rdata[881] or rdata[880] or rdata[879] or rdata[878] or rdata[877]
 or rdata[876] or rdata[875] or rdata[874] or rdata[873] or rdata[872] or rdata[871] or rdata[870] or rdata[869]
 or rdata[868] or rdata[867] or rdata[866] or rdata[865] or rdata[864] or rdata[863] or rdata[862] or rdata[861]
 or rdata[860] or rdata[859] or rdata[858] or rdata[857] or rdata[856] or rdata[855] or rdata[854] or rdata[853]
 or rdata[852] or rdata[851] or rdata[850] or rdata[849] or rdata[848] or rdata[847] or rdata[846] or rdata[845]
 or rdata[844] or rdata[843] or rdata[842] or rdata[841] or rdata[840] or rdata[839] or rdata[838] or rdata[837]
 or rdata[836] or rdata[835] or rdata[834] or rdata[833] or rdata[832] or rdata[831] or rdata[830] or rdata[829]
 or rdata[828] or rdata[827] or rdata[826] or rdata[825] or rdata[824] or rdata[823] or rdata[822] or rdata[821]
 or rdata[820] or rdata[819] or rdata[818] or rdata[817] or rdata[816] or rdata[815] or rdata[814] or rdata[813]
 or rdata[812] or rdata[811] or rdata[810] or rdata[809] or rdata[808] or rdata[807] or rdata[806] or rdata[805]
 or rdata[804] or rdata[803] or rdata[802] or rdata[801] or rdata[800] or rdata[799] or rdata[798] or rdata[797]
 or rdata[796] or rdata[795] or rdata[794] or rdata[793] or rdata[792] or rdata[791] or rdata[790] or rdata[789]
 or rdata[788] or rdata[787] or rdata[786] or rdata[785] or rdata[784] or rdata[783] or rdata[782] or rdata[781]
 or rdata[780] or rdata[779] or rdata[778] or rdata[777] or rdata[776] or rdata[775] or rdata[774] or rdata[773]
 or rdata[772] or rdata[771] or rdata[770] or rdata[769] or rdata[768] or rdata[767] or rdata[766] or rdata[765]
 or rdata[764] or rdata[763] or rdata[762] or rdata[761] or rdata[760] or rdata[759] or rdata[758] or rdata[757]
 or rdata[756] or rdata[755] or rdata[754] or rdata[753] or rdata[752] or rdata[751] or rdata[750] or rdata[749]
 or rdata[748] or rdata[747] or rdata[746] or rdata[745] or rdata[744] or rdata[743] or rdata[742] or rdata[741]
 or rdata[740] or rdata[739] or rdata[738] or rdata[737] or rdata[736] or rdata[735] or rdata[734] or rdata[733]
 or rdata[732] or rdata[731] or rdata[730] or rdata[729] or rdata[728] or rdata[727] or rdata[726] or rdata[725]
 or rdata[724] or rdata[723] or rdata[722] or rdata[721] or rdata[720] or rdata[719] or rdata[718] or rdata[717]
 or rdata[716] or rdata[715] or rdata[714] or rdata[713] or rdata[712] or rdata[711] or rdata[710] or rdata[709]
 or rdata[708] or rdata[707] or rdata[706] or rdata[705] or rdata[704] or rdata[703] or rdata[702] or rdata[701]
 or rdata[700] or rdata[699] or rdata[698] or rdata[697] or rdata[696] or rdata[695] or rdata[694] or rdata[693]
 or rdata[692] or rdata[691] or rdata[690] or rdata[689] or rdata[688] or rdata[687] or rdata[686] or rdata[685]
 or rdata[684] or rdata[683] or rdata[682] or rdata[681] or rdata[680] or rdata[679] or rdata[678] or rdata[677]
 or rdata[676] or rdata[675] or rdata[674] or rdata[673] or rdata[672] or rdata[671] or rdata[670] or rdata[669]
 or rdata[668] or rdata[667] or rdata[666] or rdata[665] or rdata[664] or rdata[663] or rdata[662] or rdata[661]
 or rdata[660] or rdata[659] or rdata[658] or rdata[657] or rdata[656] or rdata[655] or rdata[654] or rdata[653]
 or rdata[652] or rdata[651] or rdata[650] or rdata[649] or rdata[648] or rdata[647] or rdata[646] or rdata[645]
 or rdata[644] or rdata[643] or rdata[642] or rdata[641] or rdata[640] or rdata[639] or rdata[638] or rdata[637]
 or rdata[636] or rdata[635] or rdata[634] or rdata[633] or rdata[632] or rdata[631] or rdata[630] or rdata[629]
 or rdata[628] or rdata[627] or rdata[626] or rdata[625] or rdata[624] or rdata[623] or rdata[622] or rdata[621]
 or rdata[620] or rdata[619] or rdata[618] or rdata[617] or rdata[616] or rdata[615] or rdata[614] or rdata[613]
 or rdata[612] or rdata[611] or rdata[610] or rdata[609] or rdata[608] or rdata[607] or rdata[606] or rdata[605]
 or rdata[604] or rdata[603] or rdata[602] or rdata[601] or rdata[600] or rdata[599] or rdata[598] or rdata[597]
 or rdata[596] or rdata[595] or rdata[594] or rdata[593] or rdata[592] or rdata[591] or rdata[590] or rdata[589]
 or rdata[588] or rdata[587] or rdata[586] or rdata[585] or rdata[584] or rdata[583] or rdata[582] or rdata[581]
 or rdata[580] or rdata[579] or rdata[578] or rdata[577] or rdata[576] or rdata[575] or rdata[574] or rdata[573]
 or rdata[572] or rdata[571] or rdata[570] or rdata[569] or rdata[568] or rdata[567] or rdata[566] or rdata[565]
 or rdata[564] or rdata[563] or rdata[562] or rdata[561] or rdata[560] or rdata[559] or rdata[558] or rdata[557]
 or rdata[556] or rdata[555] or rdata[554] or rdata[553] or rdata[552] or rdata[551] or rdata[550] or rdata[549]
 or rdata[548] or rdata[547] or rdata[546] or rdata[545] or rdata[544] or rdata[543] or rdata[542] or rdata[541]
 or rdata[540] or rdata[539] or rdata[538] or rdata[537] or rdata[536] or rdata[535] or rdata[534] or rdata[533]
 or rdata[532] or rdata[531] or rdata[530] or rdata[529] or rdata[528] or rdata[527] or rdata[526] or rdata[525]
 or rdata[524] or rdata[523] or rdata[522] or rdata[521] or rdata[520] or rdata[519] or rdata[518] or rdata[517]
 or rdata[516] or rdata[515] or rdata[514] or rdata[513] or rdata[512])
#0 begin
if (n1)
_zymem[{n2}] =
{rdata[511], rdata[510], rdata[509], rdata[508], rdata[507],
 rdata[506], rdata[505], rdata[504], rdata[503], rdata[502], rdata[501], rdata[500], rdata[499],
 rdata[498], rdata[497], rdata[496], rdata[495], rdata[494], rdata[493], rdata[492], rdata[491],
 rdata[490], rdata[489], rdata[488], rdata[487], rdata[486], rdata[485], rdata[484], rdata[483],
 rdata[482], rdata[481], rdata[480], rdata[479], rdata[478], rdata[477], rdata[476], rdata[475],
 rdata[474], rdata[473], rdata[472], rdata[471], rdata[470], rdata[469], rdata[468], rdata[467],
 rdata[466], rdata[465], rdata[464], rdata[463], rdata[462], rdata[461], rdata[460], rdata[459],
 rdata[458], rdata[457], rdata[456], rdata[455], rdata[454], rdata[453], rdata[452], rdata[451],
 rdata[450], rdata[449], rdata[448], rdata[447], rdata[446], rdata[445], rdata[444], rdata[443],
 rdata[442], rdata[441], rdata[440], rdata[439], rdata[438], rdata[437], rdata[436], rdata[435],
 rdata[434], rdata[433], rdata[432], rdata[431], rdata[430], rdata[429], rdata[428], rdata[427],
 rdata[426], rdata[425], rdata[424], rdata[423], rdata[422], rdata[421], rdata[420], rdata[419],
 rdata[418], rdata[417], rdata[416], rdata[415], rdata[414], rdata[413], rdata[412], rdata[411],
 rdata[410], rdata[409], rdata[408], rdata[407], rdata[406], rdata[405], rdata[404], rdata[403],
 rdata[402], rdata[401], rdata[400], rdata[399], rdata[398], rdata[397], rdata[396], rdata[395],
 rdata[394], rdata[393], rdata[392], rdata[391], rdata[390], rdata[389], rdata[388], rdata[387],
 rdata[386], rdata[385], rdata[384], rdata[383], rdata[382], rdata[381], rdata[380], rdata[379],
 rdata[378], rdata[377], rdata[376], rdata[375], rdata[374], rdata[373], rdata[372], rdata[371],
 rdata[370], rdata[369], rdata[368], rdata[367], rdata[366], rdata[365], rdata[364], rdata[363],
 rdata[362], rdata[361], rdata[360], rdata[359], rdata[358], rdata[357], rdata[356], rdata[355],
 rdata[354], rdata[353], rdata[352], rdata[351], rdata[350], rdata[349], rdata[348], rdata[347],
 rdata[346], rdata[345], rdata[344], rdata[343], rdata[342], rdata[341], rdata[340], rdata[339],
 rdata[338], rdata[337], rdata[336], rdata[335], rdata[334], rdata[333], rdata[332], rdata[331],
 rdata[330], rdata[329], rdata[328], rdata[327], rdata[326], rdata[325], rdata[324], rdata[323],
 rdata[322], rdata[321], rdata[320], rdata[319], rdata[318], rdata[317], rdata[316], rdata[315],
 rdata[314], rdata[313], rdata[312], rdata[311], rdata[310], rdata[309], rdata[308], rdata[307],
 rdata[306], rdata[305], rdata[304], rdata[303], rdata[302], rdata[301], rdata[300], rdata[299],
 rdata[298], rdata[297], rdata[296], rdata[295], rdata[294], rdata[293], rdata[292], rdata[291],
 rdata[290], rdata[289], rdata[288], rdata[287], rdata[286], rdata[285], rdata[284], rdata[283],
 rdata[282], rdata[281], rdata[280], rdata[279], rdata[278], rdata[277], rdata[276], rdata[275],
 rdata[274], rdata[273], rdata[272], rdata[271], rdata[270], rdata[269], rdata[268], rdata[267],
 rdata[266], rdata[265], rdata[264], rdata[263], rdata[262], rdata[261], rdata[260], rdata[259],
 rdata[258], rdata[257], rdata[256], rdata[255], rdata[254], rdata[253], rdata[252], rdata[251],
 rdata[250], rdata[249], rdata[248], rdata[247], rdata[246], rdata[245], rdata[244], rdata[243],
 rdata[242], rdata[241], rdata[240], rdata[239], rdata[238], rdata[237], rdata[236], rdata[235],
 rdata[234], rdata[233], rdata[232], rdata[231], rdata[230], rdata[229], rdata[228], rdata[227],
 rdata[226], rdata[225], rdata[224], rdata[223], rdata[222], rdata[221], rdata[220], rdata[219],
 rdata[218], rdata[217], rdata[216], rdata[215], rdata[214], rdata[213], rdata[212], rdata[211],
 rdata[210], rdata[209], rdata[208], rdata[207], rdata[206], rdata[205], rdata[204], rdata[203],
 rdata[202], rdata[201], rdata[200], rdata[199], rdata[198], rdata[197], rdata[196], rdata[195],
 rdata[194], rdata[193], rdata[192], rdata[191], rdata[190], rdata[189], rdata[188], rdata[187],
 rdata[186], rdata[185], rdata[184], rdata[183], rdata[182], rdata[181], rdata[180], rdata[179],
 rdata[178], rdata[177], rdata[176], rdata[175], rdata[174], rdata[173], rdata[172], rdata[171],
 rdata[170], rdata[169], rdata[168], rdata[167], rdata[166], rdata[165], rdata[164], rdata[163],
 rdata[162], rdata[161], rdata[160], rdata[159], rdata[158], rdata[157], rdata[156], rdata[155],
 rdata[154], rdata[153], rdata[152], rdata[151], rdata[150], rdata[149], rdata[148], rdata[147],
 rdata[146], rdata[145], rdata[144], rdata[143], rdata[142], rdata[141], rdata[140], rdata[139],
 rdata[138], rdata[137], rdata[136], rdata[135], rdata[134], rdata[133], rdata[132], rdata[131],
 rdata[130], rdata[129], rdata[128], rdata[127], rdata[126], rdata[125], rdata[124], rdata[123],
 rdata[122], rdata[121], rdata[120], rdata[119], rdata[118], rdata[117], rdata[116], rdata[115],
 rdata[114], rdata[113], rdata[112], rdata[111], rdata[110], rdata[109], rdata[108], rdata[107],
 rdata[106], rdata[105], rdata[104], rdata[103], rdata[102], rdata[101], rdata[100], rdata[99],
 rdata[98], rdata[97], rdata[96], rdata[95], rdata[94], rdata[93], rdata[92], rdata[91],
 rdata[90], rdata[89], rdata[88], rdata[87], rdata[86], rdata[85], rdata[84], rdata[83],
 rdata[82], rdata[81], rdata[80], rdata[79], rdata[78], rdata[77], rdata[76], rdata[75],
 rdata[74], rdata[73], rdata[72], rdata[71], rdata[70], rdata[69], rdata[68], rdata[67],
 rdata[66], rdata[65], rdata[64], rdata[63], rdata[62], rdata[61], rdata[60], rdata[59],
 rdata[58], rdata[57], rdata[56], rdata[55], rdata[54], rdata[53], rdata[52], rdata[51],
 rdata[50], rdata[49], rdata[48], rdata[47], rdata[46], rdata[45], rdata[44], rdata[43],
 rdata[42], rdata[41], rdata[40], rdata[39], rdata[38], rdata[37], rdata[36], rdata[35],
 rdata[34], rdata[33], rdata[32], rdata[31], rdata[30], rdata[29], rdata[28], rdata[27],
 rdata[26], rdata[25], rdata[24], rdata[23], rdata[22], rdata[21], rdata[20], rdata[19],
 rdata[18], rdata[17], rdata[16], rdata[15], rdata[14], rdata[13], rdata[12], rdata[11],
 rdata[10], rdata[9], rdata[8], rdata[7], rdata[6], rdata[5], rdata[4], rdata[3],
 rdata[2], rdata[1], rdata[0]};
if (n1)
_zymem[{n1}] =
{rdata[1023], rdata[1022], rdata[1021], rdata[1020], rdata[1019],
 rdata[1018], rdata[1017], rdata[1016], rdata[1015], rdata[1014], rdata[1013], rdata[1012], rdata[1011],
 rdata[1010], rdata[1009], rdata[1008], rdata[1007], rdata[1006], rdata[1005], rdata[1004], rdata[1003],
 rdata[1002], rdata[1001], rdata[1000], rdata[999], rdata[998], rdata[997], rdata[996], rdata[995],
 rdata[994], rdata[993], rdata[992], rdata[991], rdata[990], rdata[989], rdata[988], rdata[987],
 rdata[986], rdata[985], rdata[984], rdata[983], rdata[982], rdata[981], rdata[980], rdata[979],
 rdata[978], rdata[977], rdata[976], rdata[975], rdata[974], rdata[973], rdata[972], rdata[971],
 rdata[970], rdata[969], rdata[968], rdata[967], rdata[966], rdata[965], rdata[964], rdata[963],
 rdata[962], rdata[961], rdata[960], rdata[959], rdata[958], rdata[957], rdata[956], rdata[955],
 rdata[954], rdata[953], rdata[952], rdata[951], rdata[950], rdata[949], rdata[948], rdata[947],
 rdata[946], rdata[945], rdata[944], rdata[943], rdata[942], rdata[941], rdata[940], rdata[939],
 rdata[938], rdata[937], rdata[936], rdata[935], rdata[934], rdata[933], rdata[932], rdata[931],
 rdata[930], rdata[929], rdata[928], rdata[927], rdata[926], rdata[925], rdata[924], rdata[923],
 rdata[922], rdata[921], rdata[920], rdata[919], rdata[918], rdata[917], rdata[916], rdata[915],
 rdata[914], rdata[913], rdata[912], rdata[911], rdata[910], rdata[909], rdata[908], rdata[907],
 rdata[906], rdata[905], rdata[904], rdata[903], rdata[902], rdata[901], rdata[900], rdata[899],
 rdata[898], rdata[897], rdata[896], rdata[895], rdata[894], rdata[893], rdata[892], rdata[891],
 rdata[890], rdata[889], rdata[888], rdata[887], rdata[886], rdata[885], rdata[884], rdata[883],
 rdata[882], rdata[881], rdata[880], rdata[879], rdata[878], rdata[877], rdata[876], rdata[875],
 rdata[874], rdata[873], rdata[872], rdata[871], rdata[870], rdata[869], rdata[868], rdata[867],
 rdata[866], rdata[865], rdata[864], rdata[863], rdata[862], rdata[861], rdata[860], rdata[859],
 rdata[858], rdata[857], rdata[856], rdata[855], rdata[854], rdata[853], rdata[852], rdata[851],
 rdata[850], rdata[849], rdata[848], rdata[847], rdata[846], rdata[845], rdata[844], rdata[843],
 rdata[842], rdata[841], rdata[840], rdata[839], rdata[838], rdata[837], rdata[836], rdata[835],
 rdata[834], rdata[833], rdata[832], rdata[831], rdata[830], rdata[829], rdata[828], rdata[827],
 rdata[826], rdata[825], rdata[824], rdata[823], rdata[822], rdata[821], rdata[820], rdata[819],
 rdata[818], rdata[817], rdata[816], rdata[815], rdata[814], rdata[813], rdata[812], rdata[811],
 rdata[810], rdata[809], rdata[808], rdata[807], rdata[806], rdata[805], rdata[804], rdata[803],
 rdata[802], rdata[801], rdata[800], rdata[799], rdata[798], rdata[797], rdata[796], rdata[795],
 rdata[794], rdata[793], rdata[792], rdata[791], rdata[790], rdata[789], rdata[788], rdata[787],
 rdata[786], rdata[785], rdata[784], rdata[783], rdata[782], rdata[781], rdata[780], rdata[779],
 rdata[778], rdata[777], rdata[776], rdata[775], rdata[774], rdata[773], rdata[772], rdata[771],
 rdata[770], rdata[769], rdata[768], rdata[767], rdata[766], rdata[765], rdata[764], rdata[763],
 rdata[762], rdata[761], rdata[760], rdata[759], rdata[758], rdata[757], rdata[756], rdata[755],
 rdata[754], rdata[753], rdata[752], rdata[751], rdata[750], rdata[749], rdata[748], rdata[747],
 rdata[746], rdata[745], rdata[744], rdata[743], rdata[742], rdata[741], rdata[740], rdata[739],
 rdata[738], rdata[737], rdata[736], rdata[735], rdata[734], rdata[733], rdata[732], rdata[731],
 rdata[730], rdata[729], rdata[728], rdata[727], rdata[726], rdata[725], rdata[724], rdata[723],
 rdata[722], rdata[721], rdata[720], rdata[719], rdata[718], rdata[717], rdata[716], rdata[715],
 rdata[714], rdata[713], rdata[712], rdata[711], rdata[710], rdata[709], rdata[708], rdata[707],
 rdata[706], rdata[705], rdata[704], rdata[703], rdata[702], rdata[701], rdata[700], rdata[699],
 rdata[698], rdata[697], rdata[696], rdata[695], rdata[694], rdata[693], rdata[692], rdata[691],
 rdata[690], rdata[689], rdata[688], rdata[687], rdata[686], rdata[685], rdata[684], rdata[683],
 rdata[682], rdata[681], rdata[680], rdata[679], rdata[678], rdata[677], rdata[676], rdata[675],
 rdata[674], rdata[673], rdata[672], rdata[671], rdata[670], rdata[669], rdata[668], rdata[667],
 rdata[666], rdata[665], rdata[664], rdata[663], rdata[662], rdata[661], rdata[660], rdata[659],
 rdata[658], rdata[657], rdata[656], rdata[655], rdata[654], rdata[653], rdata[652], rdata[651],
 rdata[650], rdata[649], rdata[648], rdata[647], rdata[646], rdata[645], rdata[644], rdata[643],
 rdata[642], rdata[641], rdata[640], rdata[639], rdata[638], rdata[637], rdata[636], rdata[635],
 rdata[634], rdata[633], rdata[632], rdata[631], rdata[630], rdata[629], rdata[628], rdata[627],
 rdata[626], rdata[625], rdata[624], rdata[623], rdata[622], rdata[621], rdata[620], rdata[619],
 rdata[618], rdata[617], rdata[616], rdata[615], rdata[614], rdata[613], rdata[612], rdata[611],
 rdata[610], rdata[609], rdata[608], rdata[607], rdata[606], rdata[605], rdata[604], rdata[603],
 rdata[602], rdata[601], rdata[600], rdata[599], rdata[598], rdata[597], rdata[596], rdata[595],
 rdata[594], rdata[593], rdata[592], rdata[591], rdata[590], rdata[589], rdata[588], rdata[587],
 rdata[586], rdata[585], rdata[584], rdata[583], rdata[582], rdata[581], rdata[580], rdata[579],
 rdata[578], rdata[577], rdata[576], rdata[575], rdata[574], rdata[573], rdata[572], rdata[571],
 rdata[570], rdata[569], rdata[568], rdata[567], rdata[566], rdata[565], rdata[564], rdata[563],
 rdata[562], rdata[561], rdata[560], rdata[559], rdata[558], rdata[557], rdata[556], rdata[555],
 rdata[554], rdata[553], rdata[552], rdata[551], rdata[550], rdata[549], rdata[548], rdata[547],
 rdata[546], rdata[545], rdata[544], rdata[543], rdata[542], rdata[541], rdata[540], rdata[539],
 rdata[538], rdata[537], rdata[536], rdata[535], rdata[534], rdata[533], rdata[532], rdata[531],
 rdata[530], rdata[529], rdata[528], rdata[527], rdata[526], rdata[525], rdata[524], rdata[523],
 rdata[522], rdata[521], rdata[520], rdata[519], rdata[518], rdata[517], rdata[516], rdata[515],
 rdata[514], rdata[513], rdata[512]};
end
`else

MPW2X512 _zymem ( .A0(n2), .DI511(rdata[511]), .DI510(rdata[510]), .DI509(rdata[509]), .DI508(rdata[508]), .DI507(rdata[507]),
 .DI506(rdata[506]), .DI505(rdata[505]), .DI504(rdata[504]), .DI503(rdata[503]), .DI502(rdata[502]), .DI501(rdata[501]), .DI500(rdata[500]), .DI499(rdata[499]),
 .DI498(rdata[498]), .DI497(rdata[497]), .DI496(rdata[496]), .DI495(rdata[495]), .DI494(rdata[494]), .DI493(rdata[493]), .DI492(rdata[492]), .DI491(rdata[491]),
 .DI490(rdata[490]), .DI489(rdata[489]), .DI488(rdata[488]), .DI487(rdata[487]), .DI486(rdata[486]), .DI485(rdata[485]), .DI484(rdata[484]), .DI483(rdata[483]),
 .DI482(rdata[482]), .DI481(rdata[481]), .DI480(rdata[480]), .DI479(rdata[479]), .DI478(rdata[478]), .DI477(rdata[477]), .DI476(rdata[476]), .DI475(rdata[475]),
 .DI474(rdata[474]), .DI473(rdata[473]), .DI472(rdata[472]), .DI471(rdata[471]), .DI470(rdata[470]), .DI469(rdata[469]), .DI468(rdata[468]), .DI467(rdata[467]),
 .DI466(rdata[466]), .DI465(rdata[465]), .DI464(rdata[464]), .DI463(rdata[463]), .DI462(rdata[462]), .DI461(rdata[461]), .DI460(rdata[460]), .DI459(rdata[459]),
 .DI458(rdata[458]), .DI457(rdata[457]), .DI456(rdata[456]), .DI455(rdata[455]), .DI454(rdata[454]), .DI453(rdata[453]), .DI452(rdata[452]), .DI451(rdata[451]),
 .DI450(rdata[450]), .DI449(rdata[449]), .DI448(rdata[448]), .DI447(rdata[447]), .DI446(rdata[446]), .DI445(rdata[445]), .DI444(rdata[444]), .DI443(rdata[443]),
 .DI442(rdata[442]), .DI441(rdata[441]), .DI440(rdata[440]), .DI439(rdata[439]), .DI438(rdata[438]), .DI437(rdata[437]), .DI436(rdata[436]), .DI435(rdata[435]),
 .DI434(rdata[434]), .DI433(rdata[433]), .DI432(rdata[432]), .DI431(rdata[431]), .DI430(rdata[430]), .DI429(rdata[429]), .DI428(rdata[428]), .DI427(rdata[427]),
 .DI426(rdata[426]), .DI425(rdata[425]), .DI424(rdata[424]), .DI423(rdata[423]), .DI422(rdata[422]), .DI421(rdata[421]), .DI420(rdata[420]), .DI419(rdata[419]),
 .DI418(rdata[418]), .DI417(rdata[417]), .DI416(rdata[416]), .DI415(rdata[415]), .DI414(rdata[414]), .DI413(rdata[413]), .DI412(rdata[412]), .DI411(rdata[411]),
 .DI410(rdata[410]), .DI409(rdata[409]), .DI408(rdata[408]), .DI407(rdata[407]), .DI406(rdata[406]), .DI405(rdata[405]), .DI404(rdata[404]), .DI403(rdata[403]),
 .DI402(rdata[402]), .DI401(rdata[401]), .DI400(rdata[400]), .DI399(rdata[399]), .DI398(rdata[398]), .DI397(rdata[397]), .DI396(rdata[396]), .DI395(rdata[395]),
 .DI394(rdata[394]), .DI393(rdata[393]), .DI392(rdata[392]), .DI391(rdata[391]), .DI390(rdata[390]), .DI389(rdata[389]), .DI388(rdata[388]), .DI387(rdata[387]),
 .DI386(rdata[386]), .DI385(rdata[385]), .DI384(rdata[384]), .DI383(rdata[383]), .DI382(rdata[382]), .DI381(rdata[381]), .DI380(rdata[380]), .DI379(rdata[379]),
 .DI378(rdata[378]), .DI377(rdata[377]), .DI376(rdata[376]), .DI375(rdata[375]), .DI374(rdata[374]), .DI373(rdata[373]), .DI372(rdata[372]), .DI371(rdata[371]),
 .DI370(rdata[370]), .DI369(rdata[369]), .DI368(rdata[368]), .DI367(rdata[367]), .DI366(rdata[366]), .DI365(rdata[365]), .DI364(rdata[364]), .DI363(rdata[363]),
 .DI362(rdata[362]), .DI361(rdata[361]), .DI360(rdata[360]), .DI359(rdata[359]), .DI358(rdata[358]), .DI357(rdata[357]), .DI356(rdata[356]), .DI355(rdata[355]),
 .DI354(rdata[354]), .DI353(rdata[353]), .DI352(rdata[352]), .DI351(rdata[351]), .DI350(rdata[350]), .DI349(rdata[349]), .DI348(rdata[348]), .DI347(rdata[347]),
 .DI346(rdata[346]), .DI345(rdata[345]), .DI344(rdata[344]), .DI343(rdata[343]), .DI342(rdata[342]), .DI341(rdata[341]), .DI340(rdata[340]), .DI339(rdata[339]),
 .DI338(rdata[338]), .DI337(rdata[337]), .DI336(rdata[336]), .DI335(rdata[335]), .DI334(rdata[334]), .DI333(rdata[333]), .DI332(rdata[332]), .DI331(rdata[331]),
 .DI330(rdata[330]), .DI329(rdata[329]), .DI328(rdata[328]), .DI327(rdata[327]), .DI326(rdata[326]), .DI325(rdata[325]), .DI324(rdata[324]), .DI323(rdata[323]),
 .DI322(rdata[322]), .DI321(rdata[321]), .DI320(rdata[320]), .DI319(rdata[319]), .DI318(rdata[318]), .DI317(rdata[317]), .DI316(rdata[316]), .DI315(rdata[315]),
 .DI314(rdata[314]), .DI313(rdata[313]), .DI312(rdata[312]), .DI311(rdata[311]), .DI310(rdata[310]), .DI309(rdata[309]), .DI308(rdata[308]), .DI307(rdata[307]),
 .DI306(rdata[306]), .DI305(rdata[305]), .DI304(rdata[304]), .DI303(rdata[303]), .DI302(rdata[302]), .DI301(rdata[301]), .DI300(rdata[300]), .DI299(rdata[299]),
 .DI298(rdata[298]), .DI297(rdata[297]), .DI296(rdata[296]), .DI295(rdata[295]), .DI294(rdata[294]), .DI293(rdata[293]), .DI292(rdata[292]), .DI291(rdata[291]),
 .DI290(rdata[290]), .DI289(rdata[289]), .DI288(rdata[288]), .DI287(rdata[287]), .DI286(rdata[286]), .DI285(rdata[285]), .DI284(rdata[284]), .DI283(rdata[283]),
 .DI282(rdata[282]), .DI281(rdata[281]), .DI280(rdata[280]), .DI279(rdata[279]), .DI278(rdata[278]), .DI277(rdata[277]), .DI276(rdata[276]), .DI275(rdata[275]),
 .DI274(rdata[274]), .DI273(rdata[273]), .DI272(rdata[272]), .DI271(rdata[271]), .DI270(rdata[270]), .DI269(rdata[269]), .DI268(rdata[268]), .DI267(rdata[267]),
 .DI266(rdata[266]), .DI265(rdata[265]), .DI264(rdata[264]), .DI263(rdata[263]), .DI262(rdata[262]), .DI261(rdata[261]), .DI260(rdata[260]), .DI259(rdata[259]),
 .DI258(rdata[258]), .DI257(rdata[257]), .DI256(rdata[256]), .DI255(rdata[255]), .DI254(rdata[254]), .DI253(rdata[253]), .DI252(rdata[252]), .DI251(rdata[251]),
 .DI250(rdata[250]), .DI249(rdata[249]), .DI248(rdata[248]), .DI247(rdata[247]), .DI246(rdata[246]), .DI245(rdata[245]), .DI244(rdata[244]), .DI243(rdata[243]),
 .DI242(rdata[242]), .DI241(rdata[241]), .DI240(rdata[240]), .DI239(rdata[239]), .DI238(rdata[238]), .DI237(rdata[237]), .DI236(rdata[236]), .DI235(rdata[235]),
 .DI234(rdata[234]), .DI233(rdata[233]), .DI232(rdata[232]), .DI231(rdata[231]), .DI230(rdata[230]), .DI229(rdata[229]), .DI228(rdata[228]), .DI227(rdata[227]),
 .DI226(rdata[226]), .DI225(rdata[225]), .DI224(rdata[224]), .DI223(rdata[223]), .DI222(rdata[222]), .DI221(rdata[221]), .DI220(rdata[220]), .DI219(rdata[219]),
 .DI218(rdata[218]), .DI217(rdata[217]), .DI216(rdata[216]), .DI215(rdata[215]), .DI214(rdata[214]), .DI213(rdata[213]), .DI212(rdata[212]), .DI211(rdata[211]),
 .DI210(rdata[210]), .DI209(rdata[209]), .DI208(rdata[208]), .DI207(rdata[207]), .DI206(rdata[206]), .DI205(rdata[205]), .DI204(rdata[204]), .DI203(rdata[203]),
 .DI202(rdata[202]), .DI201(rdata[201]), .DI200(rdata[200]), .DI199(rdata[199]), .DI198(rdata[198]), .DI197(rdata[197]), .DI196(rdata[196]), .DI195(rdata[195]),
 .DI194(rdata[194]), .DI193(rdata[193]), .DI192(rdata[192]), .DI191(rdata[191]), .DI190(rdata[190]), .DI189(rdata[189]), .DI188(rdata[188]), .DI187(rdata[187]),
 .DI186(rdata[186]), .DI185(rdata[185]), .DI184(rdata[184]), .DI183(rdata[183]), .DI182(rdata[182]), .DI181(rdata[181]), .DI180(rdata[180]), .DI179(rdata[179]),
 .DI178(rdata[178]), .DI177(rdata[177]), .DI176(rdata[176]), .DI175(rdata[175]), .DI174(rdata[174]), .DI173(rdata[173]), .DI172(rdata[172]), .DI171(rdata[171]),
 .DI170(rdata[170]), .DI169(rdata[169]), .DI168(rdata[168]), .DI167(rdata[167]), .DI166(rdata[166]), .DI165(rdata[165]), .DI164(rdata[164]), .DI163(rdata[163]),
 .DI162(rdata[162]), .DI161(rdata[161]), .DI160(rdata[160]), .DI159(rdata[159]), .DI158(rdata[158]), .DI157(rdata[157]), .DI156(rdata[156]), .DI155(rdata[155]),
 .DI154(rdata[154]), .DI153(rdata[153]), .DI152(rdata[152]), .DI151(rdata[151]), .DI150(rdata[150]), .DI149(rdata[149]), .DI148(rdata[148]), .DI147(rdata[147]),
 .DI146(rdata[146]), .DI145(rdata[145]), .DI144(rdata[144]), .DI143(rdata[143]), .DI142(rdata[142]), .DI141(rdata[141]), .DI140(rdata[140]), .DI139(rdata[139]),
 .DI138(rdata[138]), .DI137(rdata[137]), .DI136(rdata[136]), .DI135(rdata[135]), .DI134(rdata[134]), .DI133(rdata[133]), .DI132(rdata[132]), .DI131(rdata[131]),
 .DI130(rdata[130]), .DI129(rdata[129]), .DI128(rdata[128]), .DI127(rdata[127]), .DI126(rdata[126]), .DI125(rdata[125]), .DI124(rdata[124]), .DI123(rdata[123]),
 .DI122(rdata[122]), .DI121(rdata[121]), .DI120(rdata[120]), .DI119(rdata[119]), .DI118(rdata[118]), .DI117(rdata[117]), .DI116(rdata[116]), .DI115(rdata[115]),
 .DI114(rdata[114]), .DI113(rdata[113]), .DI112(rdata[112]), .DI111(rdata[111]), .DI110(rdata[110]), .DI109(rdata[109]), .DI108(rdata[108]), .DI107(rdata[107]),
 .DI106(rdata[106]), .DI105(rdata[105]), .DI104(rdata[104]), .DI103(rdata[103]), .DI102(rdata[102]), .DI101(rdata[101]), .DI100(rdata[100]), .DI99(rdata[99]),
 .DI98(rdata[98]), .DI97(rdata[97]), .DI96(rdata[96]), .DI95(rdata[95]), .DI94(rdata[94]), .DI93(rdata[93]), .DI92(rdata[92]), .DI91(rdata[91]),
 .DI90(rdata[90]), .DI89(rdata[89]), .DI88(rdata[88]), .DI87(rdata[87]), .DI86(rdata[86]), .DI85(rdata[85]), .DI84(rdata[84]), .DI83(rdata[83]),
 .DI82(rdata[82]), .DI81(rdata[81]), .DI80(rdata[80]), .DI79(rdata[79]), .DI78(rdata[78]), .DI77(rdata[77]), .DI76(rdata[76]), .DI75(rdata[75]),
 .DI74(rdata[74]), .DI73(rdata[73]), .DI72(rdata[72]), .DI71(rdata[71]), .DI70(rdata[70]), .DI69(rdata[69]), .DI68(rdata[68]), .DI67(rdata[67]),
 .DI66(rdata[66]), .DI65(rdata[65]), .DI64(rdata[64]), .DI63(rdata[63]), .DI62(rdata[62]), .DI61(rdata[61]), .DI60(rdata[60]), .DI59(rdata[59]),
 .DI58(rdata[58]), .DI57(rdata[57]), .DI56(rdata[56]), .DI55(rdata[55]), .DI54(rdata[54]), .DI53(rdata[53]), .DI52(rdata[52]), .DI51(rdata[51]),
 .DI50(rdata[50]), .DI49(rdata[49]), .DI48(rdata[48]), .DI47(rdata[47]), .DI46(rdata[46]), .DI45(rdata[45]), .DI44(rdata[44]), .DI43(rdata[43]),
 .DI42(rdata[42]), .DI41(rdata[41]), .DI40(rdata[40]), .DI39(rdata[39]), .DI38(rdata[38]), .DI37(rdata[37]), .DI36(rdata[36]), .DI35(rdata[35]),
 .DI34(rdata[34]), .DI33(rdata[33]), .DI32(rdata[32]), .DI31(rdata[31]), .DI30(rdata[30]), .DI29(rdata[29]), .DI28(rdata[28]), .DI27(rdata[27]),
 .DI26(rdata[26]), .DI25(rdata[25]), .DI24(rdata[24]), .DI23(rdata[23]), .DI22(rdata[22]), .DI21(rdata[21]), .DI20(rdata[20]), .DI19(rdata[19]),
 .DI18(rdata[18]), .DI17(rdata[17]), .DI16(rdata[16]), .DI15(rdata[15]), .DI14(rdata[14]), .DI13(rdata[13]), .DI12(rdata[12]), .DI11(rdata[11]),
 .DI10(rdata[10]), .DI9(rdata[9]), .DI8(rdata[8]), .DI7(rdata[7]), .DI6(rdata[6]), .DI5(rdata[5]), .DI4(rdata[4]), .DI3(rdata[3]),
 .DI2(rdata[2]), .DI1(rdata[1]), .DI0(rdata[0]), .WE(n1), .SYNC_IN(n2), .SYNC_OUT(n4));
// pragma CVASTRPROP INSTANCE "_zymem" HDL_MEMORY_DECL "1 511 0 0 1"
MPW2X512 U2 ( .A0(n1), .DI511(rdata[1023]), .DI510(rdata[1022]), .DI509(rdata[1021]), .DI508(rdata[1020]), .DI507(rdata[1019]),
 .DI506(rdata[1018]), .DI505(rdata[1017]), .DI504(rdata[1016]), .DI503(rdata[1015]), .DI502(rdata[1014]), .DI501(rdata[1013]), .DI500(rdata[1012]), .DI499(rdata[1011]),
 .DI498(rdata[1010]), .DI497(rdata[1009]), .DI496(rdata[1008]), .DI495(rdata[1007]), .DI494(rdata[1006]), .DI493(rdata[1005]), .DI492(rdata[1004]), .DI491(rdata[1003]),
 .DI490(rdata[1002]), .DI489(rdata[1001]), .DI488(rdata[1000]), .DI487(rdata[999]), .DI486(rdata[998]), .DI485(rdata[997]), .DI484(rdata[996]), .DI483(rdata[995]),
 .DI482(rdata[994]), .DI481(rdata[993]), .DI480(rdata[992]), .DI479(rdata[991]), .DI478(rdata[990]), .DI477(rdata[989]), .DI476(rdata[988]), .DI475(rdata[987]),
 .DI474(rdata[986]), .DI473(rdata[985]), .DI472(rdata[984]), .DI471(rdata[983]), .DI470(rdata[982]), .DI469(rdata[981]), .DI468(rdata[980]), .DI467(rdata[979]),
 .DI466(rdata[978]), .DI465(rdata[977]), .DI464(rdata[976]), .DI463(rdata[975]), .DI462(rdata[974]), .DI461(rdata[973]), .DI460(rdata[972]), .DI459(rdata[971]),
 .DI458(rdata[970]), .DI457(rdata[969]), .DI456(rdata[968]), .DI455(rdata[967]), .DI454(rdata[966]), .DI453(rdata[965]), .DI452(rdata[964]), .DI451(rdata[963]),
 .DI450(rdata[962]), .DI449(rdata[961]), .DI448(rdata[960]), .DI447(rdata[959]), .DI446(rdata[958]), .DI445(rdata[957]), .DI444(rdata[956]), .DI443(rdata[955]),
 .DI442(rdata[954]), .DI441(rdata[953]), .DI440(rdata[952]), .DI439(rdata[951]), .DI438(rdata[950]), .DI437(rdata[949]), .DI436(rdata[948]), .DI435(rdata[947]),
 .DI434(rdata[946]), .DI433(rdata[945]), .DI432(rdata[944]), .DI431(rdata[943]), .DI430(rdata[942]), .DI429(rdata[941]), .DI428(rdata[940]), .DI427(rdata[939]),
 .DI426(rdata[938]), .DI425(rdata[937]), .DI424(rdata[936]), .DI423(rdata[935]), .DI422(rdata[934]), .DI421(rdata[933]), .DI420(rdata[932]), .DI419(rdata[931]),
 .DI418(rdata[930]), .DI417(rdata[929]), .DI416(rdata[928]), .DI415(rdata[927]), .DI414(rdata[926]), .DI413(rdata[925]), .DI412(rdata[924]), .DI411(rdata[923]),
 .DI410(rdata[922]), .DI409(rdata[921]), .DI408(rdata[920]), .DI407(rdata[919]), .DI406(rdata[918]), .DI405(rdata[917]), .DI404(rdata[916]), .DI403(rdata[915]),
 .DI402(rdata[914]), .DI401(rdata[913]), .DI400(rdata[912]), .DI399(rdata[911]), .DI398(rdata[910]), .DI397(rdata[909]), .DI396(rdata[908]), .DI395(rdata[907]),
 .DI394(rdata[906]), .DI393(rdata[905]), .DI392(rdata[904]), .DI391(rdata[903]), .DI390(rdata[902]), .DI389(rdata[901]), .DI388(rdata[900]), .DI387(rdata[899]),
 .DI386(rdata[898]), .DI385(rdata[897]), .DI384(rdata[896]), .DI383(rdata[895]), .DI382(rdata[894]), .DI381(rdata[893]), .DI380(rdata[892]), .DI379(rdata[891]),
 .DI378(rdata[890]), .DI377(rdata[889]), .DI376(rdata[888]), .DI375(rdata[887]), .DI374(rdata[886]), .DI373(rdata[885]), .DI372(rdata[884]), .DI371(rdata[883]),
 .DI370(rdata[882]), .DI369(rdata[881]), .DI368(rdata[880]), .DI367(rdata[879]), .DI366(rdata[878]), .DI365(rdata[877]), .DI364(rdata[876]), .DI363(rdata[875]),
 .DI362(rdata[874]), .DI361(rdata[873]), .DI360(rdata[872]), .DI359(rdata[871]), .DI358(rdata[870]), .DI357(rdata[869]), .DI356(rdata[868]), .DI355(rdata[867]),
 .DI354(rdata[866]), .DI353(rdata[865]), .DI352(rdata[864]), .DI351(rdata[863]), .DI350(rdata[862]), .DI349(rdata[861]), .DI348(rdata[860]), .DI347(rdata[859]),
 .DI346(rdata[858]), .DI345(rdata[857]), .DI344(rdata[856]), .DI343(rdata[855]), .DI342(rdata[854]), .DI341(rdata[853]), .DI340(rdata[852]), .DI339(rdata[851]),
 .DI338(rdata[850]), .DI337(rdata[849]), .DI336(rdata[848]), .DI335(rdata[847]), .DI334(rdata[846]), .DI333(rdata[845]), .DI332(rdata[844]), .DI331(rdata[843]),
 .DI330(rdata[842]), .DI329(rdata[841]), .DI328(rdata[840]), .DI327(rdata[839]), .DI326(rdata[838]), .DI325(rdata[837]), .DI324(rdata[836]), .DI323(rdata[835]),
 .DI322(rdata[834]), .DI321(rdata[833]), .DI320(rdata[832]), .DI319(rdata[831]), .DI318(rdata[830]), .DI317(rdata[829]), .DI316(rdata[828]), .DI315(rdata[827]),
 .DI314(rdata[826]), .DI313(rdata[825]), .DI312(rdata[824]), .DI311(rdata[823]), .DI310(rdata[822]), .DI309(rdata[821]), .DI308(rdata[820]), .DI307(rdata[819]),
 .DI306(rdata[818]), .DI305(rdata[817]), .DI304(rdata[816]), .DI303(rdata[815]), .DI302(rdata[814]), .DI301(rdata[813]), .DI300(rdata[812]), .DI299(rdata[811]),
 .DI298(rdata[810]), .DI297(rdata[809]), .DI296(rdata[808]), .DI295(rdata[807]), .DI294(rdata[806]), .DI293(rdata[805]), .DI292(rdata[804]), .DI291(rdata[803]),
 .DI290(rdata[802]), .DI289(rdata[801]), .DI288(rdata[800]), .DI287(rdata[799]), .DI286(rdata[798]), .DI285(rdata[797]), .DI284(rdata[796]), .DI283(rdata[795]),
 .DI282(rdata[794]), .DI281(rdata[793]), .DI280(rdata[792]), .DI279(rdata[791]), .DI278(rdata[790]), .DI277(rdata[789]), .DI276(rdata[788]), .DI275(rdata[787]),
 .DI274(rdata[786]), .DI273(rdata[785]), .DI272(rdata[784]), .DI271(rdata[783]), .DI270(rdata[782]), .DI269(rdata[781]), .DI268(rdata[780]), .DI267(rdata[779]),
 .DI266(rdata[778]), .DI265(rdata[777]), .DI264(rdata[776]), .DI263(rdata[775]), .DI262(rdata[774]), .DI261(rdata[773]), .DI260(rdata[772]), .DI259(rdata[771]),
 .DI258(rdata[770]), .DI257(rdata[769]), .DI256(rdata[768]), .DI255(rdata[767]), .DI254(rdata[766]), .DI253(rdata[765]), .DI252(rdata[764]), .DI251(rdata[763]),
 .DI250(rdata[762]), .DI249(rdata[761]), .DI248(rdata[760]), .DI247(rdata[759]), .DI246(rdata[758]), .DI245(rdata[757]), .DI244(rdata[756]), .DI243(rdata[755]),
 .DI242(rdata[754]), .DI241(rdata[753]), .DI240(rdata[752]), .DI239(rdata[751]), .DI238(rdata[750]), .DI237(rdata[749]), .DI236(rdata[748]), .DI235(rdata[747]),
 .DI234(rdata[746]), .DI233(rdata[745]), .DI232(rdata[744]), .DI231(rdata[743]), .DI230(rdata[742]), .DI229(rdata[741]), .DI228(rdata[740]), .DI227(rdata[739]),
 .DI226(rdata[738]), .DI225(rdata[737]), .DI224(rdata[736]), .DI223(rdata[735]), .DI222(rdata[734]), .DI221(rdata[733]), .DI220(rdata[732]), .DI219(rdata[731]),
 .DI218(rdata[730]), .DI217(rdata[729]), .DI216(rdata[728]), .DI215(rdata[727]), .DI214(rdata[726]), .DI213(rdata[725]), .DI212(rdata[724]), .DI211(rdata[723]),
 .DI210(rdata[722]), .DI209(rdata[721]), .DI208(rdata[720]), .DI207(rdata[719]), .DI206(rdata[718]), .DI205(rdata[717]), .DI204(rdata[716]), .DI203(rdata[715]),
 .DI202(rdata[714]), .DI201(rdata[713]), .DI200(rdata[712]), .DI199(rdata[711]), .DI198(rdata[710]), .DI197(rdata[709]), .DI196(rdata[708]), .DI195(rdata[707]),
 .DI194(rdata[706]), .DI193(rdata[705]), .DI192(rdata[704]), .DI191(rdata[703]), .DI190(rdata[702]), .DI189(rdata[701]), .DI188(rdata[700]), .DI187(rdata[699]),
 .DI186(rdata[698]), .DI185(rdata[697]), .DI184(rdata[696]), .DI183(rdata[695]), .DI182(rdata[694]), .DI181(rdata[693]), .DI180(rdata[692]), .DI179(rdata[691]),
 .DI178(rdata[690]), .DI177(rdata[689]), .DI176(rdata[688]), .DI175(rdata[687]), .DI174(rdata[686]), .DI173(rdata[685]), .DI172(rdata[684]), .DI171(rdata[683]),
 .DI170(rdata[682]), .DI169(rdata[681]), .DI168(rdata[680]), .DI167(rdata[679]), .DI166(rdata[678]), .DI165(rdata[677]), .DI164(rdata[676]), .DI163(rdata[675]),
 .DI162(rdata[674]), .DI161(rdata[673]), .DI160(rdata[672]), .DI159(rdata[671]), .DI158(rdata[670]), .DI157(rdata[669]), .DI156(rdata[668]), .DI155(rdata[667]),
 .DI154(rdata[666]), .DI153(rdata[665]), .DI152(rdata[664]), .DI151(rdata[663]), .DI150(rdata[662]), .DI149(rdata[661]), .DI148(rdata[660]), .DI147(rdata[659]),
 .DI146(rdata[658]), .DI145(rdata[657]), .DI144(rdata[656]), .DI143(rdata[655]), .DI142(rdata[654]), .DI141(rdata[653]), .DI140(rdata[652]), .DI139(rdata[651]),
 .DI138(rdata[650]), .DI137(rdata[649]), .DI136(rdata[648]), .DI135(rdata[647]), .DI134(rdata[646]), .DI133(rdata[645]), .DI132(rdata[644]), .DI131(rdata[643]),
 .DI130(rdata[642]), .DI129(rdata[641]), .DI128(rdata[640]), .DI127(rdata[639]), .DI126(rdata[638]), .DI125(rdata[637]), .DI124(rdata[636]), .DI123(rdata[635]),
 .DI122(rdata[634]), .DI121(rdata[633]), .DI120(rdata[632]), .DI119(rdata[631]), .DI118(rdata[630]), .DI117(rdata[629]), .DI116(rdata[628]), .DI115(rdata[627]),
 .DI114(rdata[626]), .DI113(rdata[625]), .DI112(rdata[624]), .DI111(rdata[623]), .DI110(rdata[622]), .DI109(rdata[621]), .DI108(rdata[620]), .DI107(rdata[619]),
 .DI106(rdata[618]), .DI105(rdata[617]), .DI104(rdata[616]), .DI103(rdata[615]), .DI102(rdata[614]), .DI101(rdata[613]), .DI100(rdata[612]), .DI99(rdata[611]),
 .DI98(rdata[610]), .DI97(rdata[609]), .DI96(rdata[608]), .DI95(rdata[607]), .DI94(rdata[606]), .DI93(rdata[605]), .DI92(rdata[604]), .DI91(rdata[603]),
 .DI90(rdata[602]), .DI89(rdata[601]), .DI88(rdata[600]), .DI87(rdata[599]), .DI86(rdata[598]), .DI85(rdata[597]), .DI84(rdata[596]), .DI83(rdata[595]),
 .DI82(rdata[594]), .DI81(rdata[593]), .DI80(rdata[592]), .DI79(rdata[591]), .DI78(rdata[590]), .DI77(rdata[589]), .DI76(rdata[588]), .DI75(rdata[587]),
 .DI74(rdata[586]), .DI73(rdata[585]), .DI72(rdata[584]), .DI71(rdata[583]), .DI70(rdata[582]), .DI69(rdata[581]), .DI68(rdata[580]), .DI67(rdata[579]),
 .DI66(rdata[578]), .DI65(rdata[577]), .DI64(rdata[576]), .DI63(rdata[575]), .DI62(rdata[574]), .DI61(rdata[573]), .DI60(rdata[572]), .DI59(rdata[571]),
 .DI58(rdata[570]), .DI57(rdata[569]), .DI56(rdata[568]), .DI55(rdata[567]), .DI54(rdata[566]), .DI53(rdata[565]), .DI52(rdata[564]), .DI51(rdata[563]),
 .DI50(rdata[562]), .DI49(rdata[561]), .DI48(rdata[560]), .DI47(rdata[559]), .DI46(rdata[558]), .DI45(rdata[557]), .DI44(rdata[556]), .DI43(rdata[555]),
 .DI42(rdata[554]), .DI41(rdata[553]), .DI40(rdata[552]), .DI39(rdata[551]), .DI38(rdata[550]), .DI37(rdata[549]), .DI36(rdata[548]), .DI35(rdata[547]),
 .DI34(rdata[546]), .DI33(rdata[545]), .DI32(rdata[544]), .DI31(rdata[543]), .DI30(rdata[542]), .DI29(rdata[541]), .DI28(rdata[540]), .DI27(rdata[539]),
 .DI26(rdata[538]), .DI25(rdata[537]), .DI24(rdata[536]), .DI23(rdata[535]), .DI22(rdata[534]), .DI21(rdata[533]), .DI20(rdata[532]), .DI19(rdata[531]),
 .DI18(rdata[530]), .DI17(rdata[529]), .DI16(rdata[528]), .DI15(rdata[527]), .DI14(rdata[526]), .DI13(rdata[525]), .DI12(rdata[524]), .DI11(rdata[523]),
 .DI10(rdata[522]), .DI9(rdata[521]), .DI8(rdata[520]), .DI7(rdata[519]), .DI6(rdata[518]), .DI5(rdata[517]), .DI4(rdata[516]), .DI3(rdata[515]),
 .DI2(rdata[514]), .DI1(rdata[513]), .DI0(rdata[512]), .WE(n1), .SYNC_IN(n4), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "_zymem 1 511 0 0 1"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE CVAIUSNAMES_FORGEN_LABEL "genblk1"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "ixc_context_read"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW2X512_MPR2X512
`else
module MPW2X512( A0, DI511, DI510, DI509, DI508, DI507, DI506,
 DI505, DI504, DI503, DI502, DI501, DI500, DI499, DI498,
 DI497, DI496, DI495, DI494, DI493, DI492, DI491, DI490,
 DI489, DI488, DI487, DI486, DI485, DI484, DI483, DI482,
 DI481, DI480, DI479, DI478, DI477, DI476, DI475, DI474,
 DI473, DI472, DI471, DI470, DI469, DI468, DI467, DI466,
 DI465, DI464, DI463, DI462, DI461, DI460, DI459, DI458,
 DI457, DI456, DI455, DI454, DI453, DI452, DI451, DI450,
 DI449, DI448, DI447, DI446, DI445, DI444, DI443, DI442,
 DI441, DI440, DI439, DI438, DI437, DI436, DI435, DI434,
 DI433, DI432, DI431, DI430, DI429, DI428, DI427, DI426,
 DI425, DI424, DI423, DI422, DI421, DI420, DI419, DI418,
 DI417, DI416, DI415, DI414, DI413, DI412, DI411, DI410,
 DI409, DI408, DI407, DI406, DI405, DI404, DI403, DI402,
 DI401, DI400, DI399, DI398, DI397, DI396, DI395, DI394,
 DI393, DI392, DI391, DI390, DI389, DI388, DI387, DI386,
 DI385, DI384, DI383, DI382, DI381, DI380, DI379, DI378,
 DI377, DI376, DI375, DI374, DI373, DI372, DI371, DI370,
 DI369, DI368, DI367, DI366, DI365, DI364, DI363, DI362,
 DI361, DI360, DI359, DI358, DI357, DI356, DI355, DI354,
 DI353, DI352, DI351, DI350, DI349, DI348, DI347, DI346,
 DI345, DI344, DI343, DI342, DI341, DI340, DI339, DI338,
 DI337, DI336, DI335, DI334, DI333, DI332, DI331, DI330,
 DI329, DI328, DI327, DI326, DI325, DI324, DI323, DI322,
 DI321, DI320, DI319, DI318, DI317, DI316, DI315, DI314,
 DI313, DI312, DI311, DI310, DI309, DI308, DI307, DI306,
 DI305, DI304, DI303, DI302, DI301, DI300, DI299, DI298,
 DI297, DI296, DI295, DI294, DI293, DI292, DI291, DI290,
 DI289, DI288, DI287, DI286, DI285, DI284, DI283, DI282,
 DI281, DI280, DI279, DI278, DI277, DI276, DI275, DI274,
 DI273, DI272, DI271, DI270, DI269, DI268, DI267, DI266,
 DI265, DI264, DI263, DI262, DI261, DI260, DI259, DI258,
 DI257, DI256, DI255, DI254, DI253, DI252, DI251, DI250,
 DI249, DI248, DI247, DI246, DI245, DI244, DI243, DI242,
 DI241, DI240, DI239, DI238, DI237, DI236, DI235, DI234,
 DI233, DI232, DI231, DI230, DI229, DI228, DI227, DI226,
 DI225, DI224, DI223, DI222, DI221, DI220, DI219, DI218,
 DI217, DI216, DI215, DI214, DI213, DI212, DI211, DI210,
 DI209, DI208, DI207, DI206, DI205, DI204, DI203, DI202,
 DI201, DI200, DI199, DI198, DI197, DI196, DI195, DI194,
 DI193, DI192, DI191, DI190, DI189, DI188, DI187, DI186,
 DI185, DI184, DI183, DI182, DI181, DI180, DI179, DI178,
 DI177, DI176, DI175, DI174, DI173, DI172, DI171, DI170,
 DI169, DI168, DI167, DI166, DI165, DI164, DI163, DI162,
 DI161, DI160, DI159, DI158, DI157, DI156, DI155, DI154,
 DI153, DI152, DI151, DI150, DI149, DI148, DI147, DI146,
 DI145, DI144, DI143, DI142, DI141, DI140, DI139, DI138,
 DI137, DI136, DI135, DI134, DI133, DI132, DI131, DI130,
 DI129, DI128, DI127, DI126, DI125, DI124, DI123, DI122,
 DI121, DI120, DI119, DI118, DI117, DI116, DI115, DI114,
 DI113, DI112, DI111, DI110, DI109, DI108, DI107, DI106,
 DI105, DI104, DI103, DI102, DI101, DI100, DI99, DI98,
 DI97, DI96, DI95, DI94, DI93, DI92, DI91, DI90,
 DI89, DI88, DI87, DI86, DI85, DI84, DI83, DI82,
 DI81, DI80, DI79, DI78, DI77, DI76, DI75, DI74,
 DI73, DI72, DI71, DI70, DI69, DI68, DI67, DI66,
 DI65, DI64, DI63, DI62, DI61, DI60, DI59, DI58,
 DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42,
 DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34,
 DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26,
 DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18,
 DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2,
 DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A0, DI511, DI510, DI509, DI508, DI507, DI506, DI505,
 DI504, DI503, DI502, DI501, DI500, DI499, DI498, DI497, DI496, DI495,
 DI494, DI493, DI492, DI491, DI490, DI489, DI488, DI487, DI486, DI485,
 DI484, DI483, DI482, DI481, DI480, DI479, DI478, DI477, DI476, DI475,
 DI474, DI473, DI472, DI471, DI470, DI469, DI468, DI467, DI466, DI465,
 DI464, DI463, DI462, DI461, DI460, DI459, DI458, DI457, DI456, DI455,
 DI454, DI453, DI452, DI451, DI450, DI449, DI448, DI447, DI446, DI445,
 DI444, DI443, DI442, DI441, DI440, DI439, DI438, DI437, DI436, DI435,
 DI434, DI433, DI432, DI431, DI430, DI429, DI428, DI427, DI426, DI425,
 DI424, DI423, DI422, DI421, DI420, DI419, DI418, DI417, DI416, DI415,
 DI414, DI413, DI412, DI411, DI410, DI409, DI408, DI407, DI406, DI405,
 DI404, DI403, DI402, DI401, DI400, DI399, DI398, DI397, DI396, DI395,
 DI394, DI393, DI392, DI391, DI390, DI389, DI388, DI387, DI386, DI385,
 DI384, DI383, DI382, DI381, DI380, DI379, DI378, DI377, DI376, DI375,
 DI374, DI373, DI372, DI371, DI370, DI369, DI368, DI367, DI366, DI365,
 DI364, DI363, DI362, DI361, DI360, DI359, DI358, DI357, DI356, DI355,
 DI354, DI353, DI352, DI351, DI350, DI349, DI348, DI347, DI346, DI345,
 DI344, DI343, DI342, DI341, DI340, DI339, DI338, DI337, DI336, DI335,
 DI334, DI333, DI332, DI331, DI330, DI329, DI328, DI327, DI326, DI325,
 DI324, DI323, DI322, DI321, DI320, DI319, DI318, DI317, DI316, DI315,
 DI314, DI313, DI312, DI311, DI310, DI309, DI308, DI307, DI306, DI305,
 DI304, DI303, DI302, DI301, DI300, DI299, DI298, DI297, DI296, DI295,
 DI294, DI293, DI292, DI291, DI290, DI289, DI288, DI287, DI286, DI285,
 DI284, DI283, DI282, DI281, DI280, DI279, DI278, DI277, DI276, DI275,
 DI274, DI273, DI272, DI271, DI270, DI269, DI268, DI267, DI266, DI265,
 DI264, DI263, DI262, DI261, DI260, DI259, DI258, DI257, DI256, DI255,
 DI254, DI253, DI252, DI251, DI250, DI249, DI248, DI247, DI246, DI245,
 DI244, DI243, DI242, DI241, DI240, DI239, DI238, DI237, DI236, DI235,
 DI234, DI233, DI232, DI231, DI230, DI229, DI228, DI227, DI226, DI225,
 DI224, DI223, DI222, DI221, DI220, DI219, DI218, DI217, DI216, DI215,
 DI214, DI213, DI212, DI211, DI210, DI209, DI208, DI207, DI206, DI205,
 DI204, DI203, DI202, DI201, DI200, DI199, DI198, DI197, DI196, DI195,
 DI194, DI193, DI192, DI191, DI190, DI189, DI188, DI187, DI186, DI185,
 DI184, DI183, DI182, DI181, DI180, DI179, DI178, DI177, DI176, DI175,
 DI174, DI173, DI172, DI171, DI170, DI169, DI168, DI167, DI166, DI165,
 DI164, DI163, DI162, DI161, DI160, DI159, DI158, DI157, DI156, DI155,
 DI154, DI153, DI152, DI151, DI150, DI149, DI148, DI147, DI146, DI145,
 DI144, DI143, DI142, DI141, DI140, DI139, DI138, DI137, DI136, DI135,
 DI134, DI133, DI132, DI131, DI130, DI129, DI128, DI127, DI126, DI125,
 DI124, DI123, DI122, DI121, DI120, DI119, DI118, DI117, DI116, DI115,
 DI114, DI113, DI112, DI111, DI110, DI109, DI108, DI107, DI106, DI105,
 DI104, DI103, DI102, DI101, DI100, DI99, DI98, DI97, DI96, DI95,
 DI94, DI93, DI92, DI91, DI90, DI89, DI88, DI87, DI86, DI85,
 DI84, DI83, DI82, DI81, DI80, DI79, DI78, DI77, DI76, DI75,
 DI74, DI73, DI72, DI71, DI70, DI69, DI68, DI67, DI66, DI65,
 DI64, DI63, DI62, DI61, DI60, DI59, DI58, DI57, DI56, DI55,
 DI54, DI53, DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45,
 DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35,
 DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25,
 DI24, DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15,
 DI14, DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5,
 DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR2X512_
`else
module MPR2X512( A0, SYNC_IN, DO511, DO510, DO509, DO508, DO507,
 DO506, DO505, DO504, DO503, DO502, DO501, DO500, DO499,
 DO498, DO497, DO496, DO495, DO494, DO493, DO492, DO491,
 DO490, DO489, DO488, DO487, DO486, DO485, DO484, DO483,
 DO482, DO481, DO480, DO479, DO478, DO477, DO476, DO475,
 DO474, DO473, DO472, DO471, DO470, DO469, DO468, DO467,
 DO466, DO465, DO464, DO463, DO462, DO461, DO460, DO459,
 DO458, DO457, DO456, DO455, DO454, DO453, DO452, DO451,
 DO450, DO449, DO448, DO447, DO446, DO445, DO444, DO443,
 DO442, DO441, DO440, DO439, DO438, DO437, DO436, DO435,
 DO434, DO433, DO432, DO431, DO430, DO429, DO428, DO427,
 DO426, DO425, DO424, DO423, DO422, DO421, DO420, DO419,
 DO418, DO417, DO416, DO415, DO414, DO413, DO412, DO411,
 DO410, DO409, DO408, DO407, DO406, DO405, DO404, DO403,
 DO402, DO401, DO400, DO399, DO398, DO397, DO396, DO395,
 DO394, DO393, DO392, DO391, DO390, DO389, DO388, DO387,
 DO386, DO385, DO384, DO383, DO382, DO381, DO380, DO379,
 DO378, DO377, DO376, DO375, DO374, DO373, DO372, DO371,
 DO370, DO369, DO368, DO367, DO366, DO365, DO364, DO363,
 DO362, DO361, DO360, DO359, DO358, DO357, DO356, DO355,
 DO354, DO353, DO352, DO351, DO350, DO349, DO348, DO347,
 DO346, DO345, DO344, DO343, DO342, DO341, DO340, DO339,
 DO338, DO337, DO336, DO335, DO334, DO333, DO332, DO331,
 DO330, DO329, DO328, DO327, DO326, DO325, DO324, DO323,
 DO322, DO321, DO320, DO319, DO318, DO317, DO316, DO315,
 DO314, DO313, DO312, DO311, DO310, DO309, DO308, DO307,
 DO306, DO305, DO304, DO303, DO302, DO301, DO300, DO299,
 DO298, DO297, DO296, DO295, DO294, DO293, DO292, DO291,
 DO290, DO289, DO288, DO287, DO286, DO285, DO284, DO283,
 DO282, DO281, DO280, DO279, DO278, DO277, DO276, DO275,
 DO274, DO273, DO272, DO271, DO270, DO269, DO268, DO267,
 DO266, DO265, DO264, DO263, DO262, DO261, DO260, DO259,
 DO258, DO257, DO256, DO255, DO254, DO253, DO252, DO251,
 DO250, DO249, DO248, DO247, DO246, DO245, DO244, DO243,
 DO242, DO241, DO240, DO239, DO238, DO237, DO236, DO235,
 DO234, DO233, DO232, DO231, DO230, DO229, DO228, DO227,
 DO226, DO225, DO224, DO223, DO222, DO221, DO220, DO219,
 DO218, DO217, DO216, DO215, DO214, DO213, DO212, DO211,
 DO210, DO209, DO208, DO207, DO206, DO205, DO204, DO203,
 DO202, DO201, DO200, DO199, DO198, DO197, DO196, DO195,
 DO194, DO193, DO192, DO191, DO190, DO189, DO188, DO187,
 DO186, DO185, DO184, DO183, DO182, DO181, DO180, DO179,
 DO178, DO177, DO176, DO175, DO174, DO173, DO172, DO171,
 DO170, DO169, DO168, DO167, DO166, DO165, DO164, DO163,
 DO162, DO161, DO160, DO159, DO158, DO157, DO156, DO155,
 DO154, DO153, DO152, DO151, DO150, DO149, DO148, DO147,
 DO146, DO145, DO144, DO143, DO142, DO141, DO140, DO139,
 DO138, DO137, DO136, DO135, DO134, DO133, DO132, DO131,
 DO130, DO129, DO128, DO127, DO126, DO125, DO124, DO123,
 DO122, DO121, DO120, DO119, DO118, DO117, DO116, DO115,
 DO114, DO113, DO112, DO111, DO110, DO109, DO108, DO107,
 DO106, DO105, DO104, DO103, DO102, DO101, DO100, DO99,
 DO98, DO97, DO96, DO95, DO94, DO93, DO92, DO91,
 DO90, DO89, DO88, DO87, DO86, DO85, DO84, DO83,
 DO82, DO81, DO80, DO79, DO78, DO77, DO76, DO75,
 DO74, DO73, DO72, DO71, DO70, DO69, DO68, DO67,
 DO66, DO65, DO64, DO63, DO62, DO61, DO60, DO59,
 DO58, DO57, DO56, DO55, DO54, DO53, DO52, DO51,
 DO50, DO49, DO48, DO47, DO46, DO45, DO44, DO43,
 DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35,
 DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27,
 DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19,
 DO18, DO17, DO16, DO15, DO14, DO13, DO12, DO11,
 DO10, DO9, DO8, DO7, DO6, DO5, DO4, DO3,
 DO2, DO1, DO0, SYNC_OUT);
input  A0, SYNC_IN;
output  DO511, DO510, DO509, DO508, DO507, DO506, DO505, DO504,
 DO503, DO502, DO501, DO500, DO499, DO498, DO497, DO496, DO495, DO494,
 DO493, DO492, DO491, DO490, DO489, DO488, DO487, DO486, DO485, DO484,
 DO483, DO482, DO481, DO480, DO479, DO478, DO477, DO476, DO475, DO474,
 DO473, DO472, DO471, DO470, DO469, DO468, DO467, DO466, DO465, DO464,
 DO463, DO462, DO461, DO460, DO459, DO458, DO457, DO456, DO455, DO454,
 DO453, DO452, DO451, DO450, DO449, DO448, DO447, DO446, DO445, DO444,
 DO443, DO442, DO441, DO440, DO439, DO438, DO437, DO436, DO435, DO434,
 DO433, DO432, DO431, DO430, DO429, DO428, DO427, DO426, DO425, DO424,
 DO423, DO422, DO421, DO420, DO419, DO418, DO417, DO416, DO415, DO414,
 DO413, DO412, DO411, DO410, DO409, DO408, DO407, DO406, DO405, DO404,
 DO403, DO402, DO401, DO400, DO399, DO398, DO397, DO396, DO395, DO394,
 DO393, DO392, DO391, DO390, DO389, DO388, DO387, DO386, DO385, DO384,
 DO383, DO382, DO381, DO380, DO379, DO378, DO377, DO376, DO375, DO374,
 DO373, DO372, DO371, DO370, DO369, DO368, DO367, DO366, DO365, DO364,
 DO363, DO362, DO361, DO360, DO359, DO358, DO357, DO356, DO355, DO354,
 DO353, DO352, DO351, DO350, DO349, DO348, DO347, DO346, DO345, DO344,
 DO343, DO342, DO341, DO340, DO339, DO338, DO337, DO336, DO335, DO334,
 DO333, DO332, DO331, DO330, DO329, DO328, DO327, DO326, DO325, DO324,
 DO323, DO322, DO321, DO320, DO319, DO318, DO317, DO316, DO315, DO314,
 DO313, DO312, DO311, DO310, DO309, DO308, DO307, DO306, DO305, DO304,
 DO303, DO302, DO301, DO300, DO299, DO298, DO297, DO296, DO295, DO294,
 DO293, DO292, DO291, DO290, DO289, DO288, DO287, DO286, DO285, DO284,
 DO283, DO282, DO281, DO280, DO279, DO278, DO277, DO276, DO275, DO274,
 DO273, DO272, DO271, DO270, DO269, DO268, DO267, DO266, DO265, DO264,
 DO263, DO262, DO261, DO260, DO259, DO258, DO257, DO256, DO255, DO254,
 DO253, DO252, DO251, DO250, DO249, DO248, DO247, DO246, DO245, DO244,
 DO243, DO242, DO241, DO240, DO239, DO238, DO237, DO236, DO235, DO234,
 DO233, DO232, DO231, DO230, DO229, DO228, DO227, DO226, DO225, DO224,
 DO223, DO222, DO221, DO220, DO219, DO218, DO217, DO216, DO215, DO214,
 DO213, DO212, DO211, DO210, DO209, DO208, DO207, DO206, DO205, DO204,
 DO203, DO202, DO201, DO200, DO199, DO198, DO197, DO196, DO195, DO194,
 DO193, DO192, DO191, DO190, DO189, DO188, DO187, DO186, DO185, DO184,
 DO183, DO182, DO181, DO180, DO179, DO178, DO177, DO176, DO175, DO174,
 DO173, DO172, DO171, DO170, DO169, DO168, DO167, DO166, DO165, DO164,
 DO163, DO162, DO161, DO160, DO159, DO158, DO157, DO156, DO155, DO154,
 DO153, DO152, DO151, DO150, DO149, DO148, DO147, DO146, DO145, DO144,
 DO143, DO142, DO141, DO140, DO139, DO138, DO137, DO136, DO135, DO134,
 DO133, DO132, DO131, DO130, DO129, DO128, DO127, DO126, DO125, DO124,
 DO123, DO122, DO121, DO120, DO119, DO118, DO117, DO116, DO115, DO114,
 DO113, DO112, DO111, DO110, DO109, DO108, DO107, DO106, DO105, DO104,
 DO103, DO102, DO101, DO100, DO99, DO98, DO97, DO96, DO95, DO94,
 DO93, DO92, DO91, DO90, DO89, DO88, DO87, DO86, DO85, DO84,
 DO83, DO82, DO81, DO80, DO79, DO78, DO77, DO76, DO75, DO74,
 DO73, DO72, DO71, DO70, DO69, DO68, DO67, DO66, DO65, DO64,
 DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56, DO55, DO54,
 DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46, DO45, DO44,
 DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35, DO34,
 DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26, DO25, DO24,
 DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6, DO5, DO4,
 DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR2X512_
`endif
`define MPW2X512_MPR2X512
`endif
`endif
