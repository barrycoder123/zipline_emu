
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_kop_gcm ( set_gcm_tag_fail_int, gcm_cmdfifo_ack, 
	gcm_upsizer_stall, gcm_tag_data_out_ack, gcm_kdf_valid, gcm_kdf_eof, 
	gcm_kdf_data, gcm_status_data_in_valid, .gcm_status_data_in( {
	\gcm_status_data_in.tag_mismatch [0]} ), clk, rst_n, 
	cmdfifo_gcm_valid, .cmdfifo_gcm_cmd( {\cmdfifo_gcm_cmd.key0 [255], 
	\cmdfifo_gcm_cmd.key0 [254], \cmdfifo_gcm_cmd.key0 [253], 
	\cmdfifo_gcm_cmd.key0 [252], \cmdfifo_gcm_cmd.key0 [251], 
	\cmdfifo_gcm_cmd.key0 [250], \cmdfifo_gcm_cmd.key0 [249], 
	\cmdfifo_gcm_cmd.key0 [248], \cmdfifo_gcm_cmd.key0 [247], 
	\cmdfifo_gcm_cmd.key0 [246], \cmdfifo_gcm_cmd.key0 [245], 
	\cmdfifo_gcm_cmd.key0 [244], \cmdfifo_gcm_cmd.key0 [243], 
	\cmdfifo_gcm_cmd.key0 [242], \cmdfifo_gcm_cmd.key0 [241], 
	\cmdfifo_gcm_cmd.key0 [240], \cmdfifo_gcm_cmd.key0 [239], 
	\cmdfifo_gcm_cmd.key0 [238], \cmdfifo_gcm_cmd.key0 [237], 
	\cmdfifo_gcm_cmd.key0 [236], \cmdfifo_gcm_cmd.key0 [235], 
	\cmdfifo_gcm_cmd.key0 [234], \cmdfifo_gcm_cmd.key0 [233], 
	\cmdfifo_gcm_cmd.key0 [232], \cmdfifo_gcm_cmd.key0 [231], 
	\cmdfifo_gcm_cmd.key0 [230], \cmdfifo_gcm_cmd.key0 [229], 
	\cmdfifo_gcm_cmd.key0 [228], \cmdfifo_gcm_cmd.key0 [227], 
	\cmdfifo_gcm_cmd.key0 [226], \cmdfifo_gcm_cmd.key0 [225], 
	\cmdfifo_gcm_cmd.key0 [224], \cmdfifo_gcm_cmd.key0 [223], 
	\cmdfifo_gcm_cmd.key0 [222], \cmdfifo_gcm_cmd.key0 [221], 
	\cmdfifo_gcm_cmd.key0 [220], \cmdfifo_gcm_cmd.key0 [219], 
	\cmdfifo_gcm_cmd.key0 [218], \cmdfifo_gcm_cmd.key0 [217], 
	\cmdfifo_gcm_cmd.key0 [216], \cmdfifo_gcm_cmd.key0 [215], 
	\cmdfifo_gcm_cmd.key0 [214], \cmdfifo_gcm_cmd.key0 [213], 
	\cmdfifo_gcm_cmd.key0 [212], \cmdfifo_gcm_cmd.key0 [211], 
	\cmdfifo_gcm_cmd.key0 [210], \cmdfifo_gcm_cmd.key0 [209], 
	\cmdfifo_gcm_cmd.key0 [208], \cmdfifo_gcm_cmd.key0 [207], 
	\cmdfifo_gcm_cmd.key0 [206], \cmdfifo_gcm_cmd.key0 [205], 
	\cmdfifo_gcm_cmd.key0 [204], \cmdfifo_gcm_cmd.key0 [203], 
	\cmdfifo_gcm_cmd.key0 [202], \cmdfifo_gcm_cmd.key0 [201], 
	\cmdfifo_gcm_cmd.key0 [200], \cmdfifo_gcm_cmd.key0 [199], 
	\cmdfifo_gcm_cmd.key0 [198], \cmdfifo_gcm_cmd.key0 [197], 
	\cmdfifo_gcm_cmd.key0 [196], \cmdfifo_gcm_cmd.key0 [195], 
	\cmdfifo_gcm_cmd.key0 [194], \cmdfifo_gcm_cmd.key0 [193], 
	\cmdfifo_gcm_cmd.key0 [192], \cmdfifo_gcm_cmd.key0 [191], 
	\cmdfifo_gcm_cmd.key0 [190], \cmdfifo_gcm_cmd.key0 [189], 
	\cmdfifo_gcm_cmd.key0 [188], \cmdfifo_gcm_cmd.key0 [187], 
	\cmdfifo_gcm_cmd.key0 [186], \cmdfifo_gcm_cmd.key0 [185], 
	\cmdfifo_gcm_cmd.key0 [184], \cmdfifo_gcm_cmd.key0 [183], 
	\cmdfifo_gcm_cmd.key0 [182], \cmdfifo_gcm_cmd.key0 [181], 
	\cmdfifo_gcm_cmd.key0 [180], \cmdfifo_gcm_cmd.key0 [179], 
	\cmdfifo_gcm_cmd.key0 [178], \cmdfifo_gcm_cmd.key0 [177], 
	\cmdfifo_gcm_cmd.key0 [176], \cmdfifo_gcm_cmd.key0 [175], 
	\cmdfifo_gcm_cmd.key0 [174], \cmdfifo_gcm_cmd.key0 [173], 
	\cmdfifo_gcm_cmd.key0 [172], \cmdfifo_gcm_cmd.key0 [171], 
	\cmdfifo_gcm_cmd.key0 [170], \cmdfifo_gcm_cmd.key0 [169], 
	\cmdfifo_gcm_cmd.key0 [168], \cmdfifo_gcm_cmd.key0 [167], 
	\cmdfifo_gcm_cmd.key0 [166], \cmdfifo_gcm_cmd.key0 [165], 
	\cmdfifo_gcm_cmd.key0 [164], \cmdfifo_gcm_cmd.key0 [163], 
	\cmdfifo_gcm_cmd.key0 [162], \cmdfifo_gcm_cmd.key0 [161], 
	\cmdfifo_gcm_cmd.key0 [160], \cmdfifo_gcm_cmd.key0 [159], 
	\cmdfifo_gcm_cmd.key0 [158], \cmdfifo_gcm_cmd.key0 [157], 
	\cmdfifo_gcm_cmd.key0 [156], \cmdfifo_gcm_cmd.key0 [155], 
	\cmdfifo_gcm_cmd.key0 [154], \cmdfifo_gcm_cmd.key0 [153], 
	\cmdfifo_gcm_cmd.key0 [152], \cmdfifo_gcm_cmd.key0 [151], 
	\cmdfifo_gcm_cmd.key0 [150], \cmdfifo_gcm_cmd.key0 [149], 
	\cmdfifo_gcm_cmd.key0 [148], \cmdfifo_gcm_cmd.key0 [147], 
	\cmdfifo_gcm_cmd.key0 [146], \cmdfifo_gcm_cmd.key0 [145], 
	\cmdfifo_gcm_cmd.key0 [144], \cmdfifo_gcm_cmd.key0 [143], 
	\cmdfifo_gcm_cmd.key0 [142], \cmdfifo_gcm_cmd.key0 [141], 
	\cmdfifo_gcm_cmd.key0 [140], \cmdfifo_gcm_cmd.key0 [139], 
	\cmdfifo_gcm_cmd.key0 [138], \cmdfifo_gcm_cmd.key0 [137], 
	\cmdfifo_gcm_cmd.key0 [136], \cmdfifo_gcm_cmd.key0 [135], 
	\cmdfifo_gcm_cmd.key0 [134], \cmdfifo_gcm_cmd.key0 [133], 
	\cmdfifo_gcm_cmd.key0 [132], \cmdfifo_gcm_cmd.key0 [131], 
	\cmdfifo_gcm_cmd.key0 [130], \cmdfifo_gcm_cmd.key0 [129], 
	\cmdfifo_gcm_cmd.key0 [128], \cmdfifo_gcm_cmd.key0 [127], 
	\cmdfifo_gcm_cmd.key0 [126], \cmdfifo_gcm_cmd.key0 [125], 
	\cmdfifo_gcm_cmd.key0 [124], \cmdfifo_gcm_cmd.key0 [123], 
	\cmdfifo_gcm_cmd.key0 [122], \cmdfifo_gcm_cmd.key0 [121], 
	\cmdfifo_gcm_cmd.key0 [120], \cmdfifo_gcm_cmd.key0 [119], 
	\cmdfifo_gcm_cmd.key0 [118], \cmdfifo_gcm_cmd.key0 [117], 
	\cmdfifo_gcm_cmd.key0 [116], \cmdfifo_gcm_cmd.key0 [115], 
	\cmdfifo_gcm_cmd.key0 [114], \cmdfifo_gcm_cmd.key0 [113], 
	\cmdfifo_gcm_cmd.key0 [112], \cmdfifo_gcm_cmd.key0 [111], 
	\cmdfifo_gcm_cmd.key0 [110], \cmdfifo_gcm_cmd.key0 [109], 
	\cmdfifo_gcm_cmd.key0 [108], \cmdfifo_gcm_cmd.key0 [107], 
	\cmdfifo_gcm_cmd.key0 [106], \cmdfifo_gcm_cmd.key0 [105], 
	\cmdfifo_gcm_cmd.key0 [104], \cmdfifo_gcm_cmd.key0 [103], 
	\cmdfifo_gcm_cmd.key0 [102], \cmdfifo_gcm_cmd.key0 [101], 
	\cmdfifo_gcm_cmd.key0 [100], \cmdfifo_gcm_cmd.key0 [99], 
	\cmdfifo_gcm_cmd.key0 [98], \cmdfifo_gcm_cmd.key0 [97], 
	\cmdfifo_gcm_cmd.key0 [96], \cmdfifo_gcm_cmd.key0 [95], 
	\cmdfifo_gcm_cmd.key0 [94], \cmdfifo_gcm_cmd.key0 [93], 
	\cmdfifo_gcm_cmd.key0 [92], \cmdfifo_gcm_cmd.key0 [91], 
	\cmdfifo_gcm_cmd.key0 [90], \cmdfifo_gcm_cmd.key0 [89], 
	\cmdfifo_gcm_cmd.key0 [88], \cmdfifo_gcm_cmd.key0 [87], 
	\cmdfifo_gcm_cmd.key0 [86], \cmdfifo_gcm_cmd.key0 [85], 
	\cmdfifo_gcm_cmd.key0 [84], \cmdfifo_gcm_cmd.key0 [83], 
	\cmdfifo_gcm_cmd.key0 [82], \cmdfifo_gcm_cmd.key0 [81], 
	\cmdfifo_gcm_cmd.key0 [80], \cmdfifo_gcm_cmd.key0 [79], 
	\cmdfifo_gcm_cmd.key0 [78], \cmdfifo_gcm_cmd.key0 [77], 
	\cmdfifo_gcm_cmd.key0 [76], \cmdfifo_gcm_cmd.key0 [75], 
	\cmdfifo_gcm_cmd.key0 [74], \cmdfifo_gcm_cmd.key0 [73], 
	\cmdfifo_gcm_cmd.key0 [72], \cmdfifo_gcm_cmd.key0 [71], 
	\cmdfifo_gcm_cmd.key0 [70], \cmdfifo_gcm_cmd.key0 [69], 
	\cmdfifo_gcm_cmd.key0 [68], \cmdfifo_gcm_cmd.key0 [67], 
	\cmdfifo_gcm_cmd.key0 [66], \cmdfifo_gcm_cmd.key0 [65], 
	\cmdfifo_gcm_cmd.key0 [64], \cmdfifo_gcm_cmd.key0 [63], 
	\cmdfifo_gcm_cmd.key0 [62], \cmdfifo_gcm_cmd.key0 [61], 
	\cmdfifo_gcm_cmd.key0 [60], \cmdfifo_gcm_cmd.key0 [59], 
	\cmdfifo_gcm_cmd.key0 [58], \cmdfifo_gcm_cmd.key0 [57], 
	\cmdfifo_gcm_cmd.key0 [56], \cmdfifo_gcm_cmd.key0 [55], 
	\cmdfifo_gcm_cmd.key0 [54], \cmdfifo_gcm_cmd.key0 [53], 
	\cmdfifo_gcm_cmd.key0 [52], \cmdfifo_gcm_cmd.key0 [51], 
	\cmdfifo_gcm_cmd.key0 [50], \cmdfifo_gcm_cmd.key0 [49], 
	\cmdfifo_gcm_cmd.key0 [48], \cmdfifo_gcm_cmd.key0 [47], 
	\cmdfifo_gcm_cmd.key0 [46], \cmdfifo_gcm_cmd.key0 [45], 
	\cmdfifo_gcm_cmd.key0 [44], \cmdfifo_gcm_cmd.key0 [43], 
	\cmdfifo_gcm_cmd.key0 [42], \cmdfifo_gcm_cmd.key0 [41], 
	\cmdfifo_gcm_cmd.key0 [40], \cmdfifo_gcm_cmd.key0 [39], 
	\cmdfifo_gcm_cmd.key0 [38], \cmdfifo_gcm_cmd.key0 [37], 
	\cmdfifo_gcm_cmd.key0 [36], \cmdfifo_gcm_cmd.key0 [35], 
	\cmdfifo_gcm_cmd.key0 [34], \cmdfifo_gcm_cmd.key0 [33], 
	\cmdfifo_gcm_cmd.key0 [32], \cmdfifo_gcm_cmd.key0 [31], 
	\cmdfifo_gcm_cmd.key0 [30], \cmdfifo_gcm_cmd.key0 [29], 
	\cmdfifo_gcm_cmd.key0 [28], \cmdfifo_gcm_cmd.key0 [27], 
	\cmdfifo_gcm_cmd.key0 [26], \cmdfifo_gcm_cmd.key0 [25], 
	\cmdfifo_gcm_cmd.key0 [24], \cmdfifo_gcm_cmd.key0 [23], 
	\cmdfifo_gcm_cmd.key0 [22], \cmdfifo_gcm_cmd.key0 [21], 
	\cmdfifo_gcm_cmd.key0 [20], \cmdfifo_gcm_cmd.key0 [19], 
	\cmdfifo_gcm_cmd.key0 [18], \cmdfifo_gcm_cmd.key0 [17], 
	\cmdfifo_gcm_cmd.key0 [16], \cmdfifo_gcm_cmd.key0 [15], 
	\cmdfifo_gcm_cmd.key0 [14], \cmdfifo_gcm_cmd.key0 [13], 
	\cmdfifo_gcm_cmd.key0 [12], \cmdfifo_gcm_cmd.key0 [11], 
	\cmdfifo_gcm_cmd.key0 [10], \cmdfifo_gcm_cmd.key0 [9], 
	\cmdfifo_gcm_cmd.key0 [8], \cmdfifo_gcm_cmd.key0 [7], 
	\cmdfifo_gcm_cmd.key0 [6], \cmdfifo_gcm_cmd.key0 [5], 
	\cmdfifo_gcm_cmd.key0 [4], \cmdfifo_gcm_cmd.key0 [3], 
	\cmdfifo_gcm_cmd.key0 [2], \cmdfifo_gcm_cmd.key0 [1], 
	\cmdfifo_gcm_cmd.key0 [0], \cmdfifo_gcm_cmd.key1 [255], 
	\cmdfifo_gcm_cmd.key1 [254], \cmdfifo_gcm_cmd.key1 [253], 
	\cmdfifo_gcm_cmd.key1 [252], \cmdfifo_gcm_cmd.key1 [251], 
	\cmdfifo_gcm_cmd.key1 [250], \cmdfifo_gcm_cmd.key1 [249], 
	\cmdfifo_gcm_cmd.key1 [248], \cmdfifo_gcm_cmd.key1 [247], 
	\cmdfifo_gcm_cmd.key1 [246], \cmdfifo_gcm_cmd.key1 [245], 
	\cmdfifo_gcm_cmd.key1 [244], \cmdfifo_gcm_cmd.key1 [243], 
	\cmdfifo_gcm_cmd.key1 [242], \cmdfifo_gcm_cmd.key1 [241], 
	\cmdfifo_gcm_cmd.key1 [240], \cmdfifo_gcm_cmd.key1 [239], 
	\cmdfifo_gcm_cmd.key1 [238], \cmdfifo_gcm_cmd.key1 [237], 
	\cmdfifo_gcm_cmd.key1 [236], \cmdfifo_gcm_cmd.key1 [235], 
	\cmdfifo_gcm_cmd.key1 [234], \cmdfifo_gcm_cmd.key1 [233], 
	\cmdfifo_gcm_cmd.key1 [232], \cmdfifo_gcm_cmd.key1 [231], 
	\cmdfifo_gcm_cmd.key1 [230], \cmdfifo_gcm_cmd.key1 [229], 
	\cmdfifo_gcm_cmd.key1 [228], \cmdfifo_gcm_cmd.key1 [227], 
	\cmdfifo_gcm_cmd.key1 [226], \cmdfifo_gcm_cmd.key1 [225], 
	\cmdfifo_gcm_cmd.key1 [224], \cmdfifo_gcm_cmd.key1 [223], 
	\cmdfifo_gcm_cmd.key1 [222], \cmdfifo_gcm_cmd.key1 [221], 
	\cmdfifo_gcm_cmd.key1 [220], \cmdfifo_gcm_cmd.key1 [219], 
	\cmdfifo_gcm_cmd.key1 [218], \cmdfifo_gcm_cmd.key1 [217], 
	\cmdfifo_gcm_cmd.key1 [216], \cmdfifo_gcm_cmd.key1 [215], 
	\cmdfifo_gcm_cmd.key1 [214], \cmdfifo_gcm_cmd.key1 [213], 
	\cmdfifo_gcm_cmd.key1 [212], \cmdfifo_gcm_cmd.key1 [211], 
	\cmdfifo_gcm_cmd.key1 [210], \cmdfifo_gcm_cmd.key1 [209], 
	\cmdfifo_gcm_cmd.key1 [208], \cmdfifo_gcm_cmd.key1 [207], 
	\cmdfifo_gcm_cmd.key1 [206], \cmdfifo_gcm_cmd.key1 [205], 
	\cmdfifo_gcm_cmd.key1 [204], \cmdfifo_gcm_cmd.key1 [203], 
	\cmdfifo_gcm_cmd.key1 [202], \cmdfifo_gcm_cmd.key1 [201], 
	\cmdfifo_gcm_cmd.key1 [200], \cmdfifo_gcm_cmd.key1 [199], 
	\cmdfifo_gcm_cmd.key1 [198], \cmdfifo_gcm_cmd.key1 [197], 
	\cmdfifo_gcm_cmd.key1 [196], \cmdfifo_gcm_cmd.key1 [195], 
	\cmdfifo_gcm_cmd.key1 [194], \cmdfifo_gcm_cmd.key1 [193], 
	\cmdfifo_gcm_cmd.key1 [192], \cmdfifo_gcm_cmd.key1 [191], 
	\cmdfifo_gcm_cmd.key1 [190], \cmdfifo_gcm_cmd.key1 [189], 
	\cmdfifo_gcm_cmd.key1 [188], \cmdfifo_gcm_cmd.key1 [187], 
	\cmdfifo_gcm_cmd.key1 [186], \cmdfifo_gcm_cmd.key1 [185], 
	\cmdfifo_gcm_cmd.key1 [184], \cmdfifo_gcm_cmd.key1 [183], 
	\cmdfifo_gcm_cmd.key1 [182], \cmdfifo_gcm_cmd.key1 [181], 
	\cmdfifo_gcm_cmd.key1 [180], \cmdfifo_gcm_cmd.key1 [179], 
	\cmdfifo_gcm_cmd.key1 [178], \cmdfifo_gcm_cmd.key1 [177], 
	\cmdfifo_gcm_cmd.key1 [176], \cmdfifo_gcm_cmd.key1 [175], 
	\cmdfifo_gcm_cmd.key1 [174], \cmdfifo_gcm_cmd.key1 [173], 
	\cmdfifo_gcm_cmd.key1 [172], \cmdfifo_gcm_cmd.key1 [171], 
	\cmdfifo_gcm_cmd.key1 [170], \cmdfifo_gcm_cmd.key1 [169], 
	\cmdfifo_gcm_cmd.key1 [168], \cmdfifo_gcm_cmd.key1 [167], 
	\cmdfifo_gcm_cmd.key1 [166], \cmdfifo_gcm_cmd.key1 [165], 
	\cmdfifo_gcm_cmd.key1 [164], \cmdfifo_gcm_cmd.key1 [163], 
	\cmdfifo_gcm_cmd.key1 [162], \cmdfifo_gcm_cmd.key1 [161], 
	\cmdfifo_gcm_cmd.key1 [160], \cmdfifo_gcm_cmd.key1 [159], 
	\cmdfifo_gcm_cmd.key1 [158], \cmdfifo_gcm_cmd.key1 [157], 
	\cmdfifo_gcm_cmd.key1 [156], \cmdfifo_gcm_cmd.key1 [155], 
	\cmdfifo_gcm_cmd.key1 [154], \cmdfifo_gcm_cmd.key1 [153], 
	\cmdfifo_gcm_cmd.key1 [152], \cmdfifo_gcm_cmd.key1 [151], 
	\cmdfifo_gcm_cmd.key1 [150], \cmdfifo_gcm_cmd.key1 [149], 
	\cmdfifo_gcm_cmd.key1 [148], \cmdfifo_gcm_cmd.key1 [147], 
	\cmdfifo_gcm_cmd.key1 [146], \cmdfifo_gcm_cmd.key1 [145], 
	\cmdfifo_gcm_cmd.key1 [144], \cmdfifo_gcm_cmd.key1 [143], 
	\cmdfifo_gcm_cmd.key1 [142], \cmdfifo_gcm_cmd.key1 [141], 
	\cmdfifo_gcm_cmd.key1 [140], \cmdfifo_gcm_cmd.key1 [139], 
	\cmdfifo_gcm_cmd.key1 [138], \cmdfifo_gcm_cmd.key1 [137], 
	\cmdfifo_gcm_cmd.key1 [136], \cmdfifo_gcm_cmd.key1 [135], 
	\cmdfifo_gcm_cmd.key1 [134], \cmdfifo_gcm_cmd.key1 [133], 
	\cmdfifo_gcm_cmd.key1 [132], \cmdfifo_gcm_cmd.key1 [131], 
	\cmdfifo_gcm_cmd.key1 [130], \cmdfifo_gcm_cmd.key1 [129], 
	\cmdfifo_gcm_cmd.key1 [128], \cmdfifo_gcm_cmd.key1 [127], 
	\cmdfifo_gcm_cmd.key1 [126], \cmdfifo_gcm_cmd.key1 [125], 
	\cmdfifo_gcm_cmd.key1 [124], \cmdfifo_gcm_cmd.key1 [123], 
	\cmdfifo_gcm_cmd.key1 [122], \cmdfifo_gcm_cmd.key1 [121], 
	\cmdfifo_gcm_cmd.key1 [120], \cmdfifo_gcm_cmd.key1 [119], 
	\cmdfifo_gcm_cmd.key1 [118], \cmdfifo_gcm_cmd.key1 [117], 
	\cmdfifo_gcm_cmd.key1 [116], \cmdfifo_gcm_cmd.key1 [115], 
	\cmdfifo_gcm_cmd.key1 [114], \cmdfifo_gcm_cmd.key1 [113], 
	\cmdfifo_gcm_cmd.key1 [112], \cmdfifo_gcm_cmd.key1 [111], 
	\cmdfifo_gcm_cmd.key1 [110], \cmdfifo_gcm_cmd.key1 [109], 
	\cmdfifo_gcm_cmd.key1 [108], \cmdfifo_gcm_cmd.key1 [107], 
	\cmdfifo_gcm_cmd.key1 [106], \cmdfifo_gcm_cmd.key1 [105], 
	\cmdfifo_gcm_cmd.key1 [104], \cmdfifo_gcm_cmd.key1 [103], 
	\cmdfifo_gcm_cmd.key1 [102], \cmdfifo_gcm_cmd.key1 [101], 
	\cmdfifo_gcm_cmd.key1 [100], \cmdfifo_gcm_cmd.key1 [99], 
	\cmdfifo_gcm_cmd.key1 [98], \cmdfifo_gcm_cmd.key1 [97], 
	\cmdfifo_gcm_cmd.key1 [96], \cmdfifo_gcm_cmd.key1 [95], 
	\cmdfifo_gcm_cmd.key1 [94], \cmdfifo_gcm_cmd.key1 [93], 
	\cmdfifo_gcm_cmd.key1 [92], \cmdfifo_gcm_cmd.key1 [91], 
	\cmdfifo_gcm_cmd.key1 [90], \cmdfifo_gcm_cmd.key1 [89], 
	\cmdfifo_gcm_cmd.key1 [88], \cmdfifo_gcm_cmd.key1 [87], 
	\cmdfifo_gcm_cmd.key1 [86], \cmdfifo_gcm_cmd.key1 [85], 
	\cmdfifo_gcm_cmd.key1 [84], \cmdfifo_gcm_cmd.key1 [83], 
	\cmdfifo_gcm_cmd.key1 [82], \cmdfifo_gcm_cmd.key1 [81], 
	\cmdfifo_gcm_cmd.key1 [80], \cmdfifo_gcm_cmd.key1 [79], 
	\cmdfifo_gcm_cmd.key1 [78], \cmdfifo_gcm_cmd.key1 [77], 
	\cmdfifo_gcm_cmd.key1 [76], \cmdfifo_gcm_cmd.key1 [75], 
	\cmdfifo_gcm_cmd.key1 [74], \cmdfifo_gcm_cmd.key1 [73], 
	\cmdfifo_gcm_cmd.key1 [72], \cmdfifo_gcm_cmd.key1 [71], 
	\cmdfifo_gcm_cmd.key1 [70], \cmdfifo_gcm_cmd.key1 [69], 
	\cmdfifo_gcm_cmd.key1 [68], \cmdfifo_gcm_cmd.key1 [67], 
	\cmdfifo_gcm_cmd.key1 [66], \cmdfifo_gcm_cmd.key1 [65], 
	\cmdfifo_gcm_cmd.key1 [64], \cmdfifo_gcm_cmd.key1 [63], 
	\cmdfifo_gcm_cmd.key1 [62], \cmdfifo_gcm_cmd.key1 [61], 
	\cmdfifo_gcm_cmd.key1 [60], \cmdfifo_gcm_cmd.key1 [59], 
	\cmdfifo_gcm_cmd.key1 [58], \cmdfifo_gcm_cmd.key1 [57], 
	\cmdfifo_gcm_cmd.key1 [56], \cmdfifo_gcm_cmd.key1 [55], 
	\cmdfifo_gcm_cmd.key1 [54], \cmdfifo_gcm_cmd.key1 [53], 
	\cmdfifo_gcm_cmd.key1 [52], \cmdfifo_gcm_cmd.key1 [51], 
	\cmdfifo_gcm_cmd.key1 [50], \cmdfifo_gcm_cmd.key1 [49], 
	\cmdfifo_gcm_cmd.key1 [48], \cmdfifo_gcm_cmd.key1 [47], 
	\cmdfifo_gcm_cmd.key1 [46], \cmdfifo_gcm_cmd.key1 [45], 
	\cmdfifo_gcm_cmd.key1 [44], \cmdfifo_gcm_cmd.key1 [43], 
	\cmdfifo_gcm_cmd.key1 [42], \cmdfifo_gcm_cmd.key1 [41], 
	\cmdfifo_gcm_cmd.key1 [40], \cmdfifo_gcm_cmd.key1 [39], 
	\cmdfifo_gcm_cmd.key1 [38], \cmdfifo_gcm_cmd.key1 [37], 
	\cmdfifo_gcm_cmd.key1 [36], \cmdfifo_gcm_cmd.key1 [35], 
	\cmdfifo_gcm_cmd.key1 [34], \cmdfifo_gcm_cmd.key1 [33], 
	\cmdfifo_gcm_cmd.key1 [32], \cmdfifo_gcm_cmd.key1 [31], 
	\cmdfifo_gcm_cmd.key1 [30], \cmdfifo_gcm_cmd.key1 [29], 
	\cmdfifo_gcm_cmd.key1 [28], \cmdfifo_gcm_cmd.key1 [27], 
	\cmdfifo_gcm_cmd.key1 [26], \cmdfifo_gcm_cmd.key1 [25], 
	\cmdfifo_gcm_cmd.key1 [24], \cmdfifo_gcm_cmd.key1 [23], 
	\cmdfifo_gcm_cmd.key1 [22], \cmdfifo_gcm_cmd.key1 [21], 
	\cmdfifo_gcm_cmd.key1 [20], \cmdfifo_gcm_cmd.key1 [19], 
	\cmdfifo_gcm_cmd.key1 [18], \cmdfifo_gcm_cmd.key1 [17], 
	\cmdfifo_gcm_cmd.key1 [16], \cmdfifo_gcm_cmd.key1 [15], 
	\cmdfifo_gcm_cmd.key1 [14], \cmdfifo_gcm_cmd.key1 [13], 
	\cmdfifo_gcm_cmd.key1 [12], \cmdfifo_gcm_cmd.key1 [11], 
	\cmdfifo_gcm_cmd.key1 [10], \cmdfifo_gcm_cmd.key1 [9], 
	\cmdfifo_gcm_cmd.key1 [8], \cmdfifo_gcm_cmd.key1 [7], 
	\cmdfifo_gcm_cmd.key1 [6], \cmdfifo_gcm_cmd.key1 [5], 
	\cmdfifo_gcm_cmd.key1 [4], \cmdfifo_gcm_cmd.key1 [3], 
	\cmdfifo_gcm_cmd.key1 [2], \cmdfifo_gcm_cmd.key1 [1], 
	\cmdfifo_gcm_cmd.key1 [0], \cmdfifo_gcm_cmd.iv [95], 
	\cmdfifo_gcm_cmd.iv [94], \cmdfifo_gcm_cmd.iv [93], 
	\cmdfifo_gcm_cmd.iv [92], \cmdfifo_gcm_cmd.iv [91], 
	\cmdfifo_gcm_cmd.iv [90], \cmdfifo_gcm_cmd.iv [89], 
	\cmdfifo_gcm_cmd.iv [88], \cmdfifo_gcm_cmd.iv [87], 
	\cmdfifo_gcm_cmd.iv [86], \cmdfifo_gcm_cmd.iv [85], 
	\cmdfifo_gcm_cmd.iv [84], \cmdfifo_gcm_cmd.iv [83], 
	\cmdfifo_gcm_cmd.iv [82], \cmdfifo_gcm_cmd.iv [81], 
	\cmdfifo_gcm_cmd.iv [80], \cmdfifo_gcm_cmd.iv [79], 
	\cmdfifo_gcm_cmd.iv [78], \cmdfifo_gcm_cmd.iv [77], 
	\cmdfifo_gcm_cmd.iv [76], \cmdfifo_gcm_cmd.iv [75], 
	\cmdfifo_gcm_cmd.iv [74], \cmdfifo_gcm_cmd.iv [73], 
	\cmdfifo_gcm_cmd.iv [72], \cmdfifo_gcm_cmd.iv [71], 
	\cmdfifo_gcm_cmd.iv [70], \cmdfifo_gcm_cmd.iv [69], 
	\cmdfifo_gcm_cmd.iv [68], \cmdfifo_gcm_cmd.iv [67], 
	\cmdfifo_gcm_cmd.iv [66], \cmdfifo_gcm_cmd.iv [65], 
	\cmdfifo_gcm_cmd.iv [64], \cmdfifo_gcm_cmd.iv [63], 
	\cmdfifo_gcm_cmd.iv [62], \cmdfifo_gcm_cmd.iv [61], 
	\cmdfifo_gcm_cmd.iv [60], \cmdfifo_gcm_cmd.iv [59], 
	\cmdfifo_gcm_cmd.iv [58], \cmdfifo_gcm_cmd.iv [57], 
	\cmdfifo_gcm_cmd.iv [56], \cmdfifo_gcm_cmd.iv [55], 
	\cmdfifo_gcm_cmd.iv [54], \cmdfifo_gcm_cmd.iv [53], 
	\cmdfifo_gcm_cmd.iv [52], \cmdfifo_gcm_cmd.iv [51], 
	\cmdfifo_gcm_cmd.iv [50], \cmdfifo_gcm_cmd.iv [49], 
	\cmdfifo_gcm_cmd.iv [48], \cmdfifo_gcm_cmd.iv [47], 
	\cmdfifo_gcm_cmd.iv [46], \cmdfifo_gcm_cmd.iv [45], 
	\cmdfifo_gcm_cmd.iv [44], \cmdfifo_gcm_cmd.iv [43], 
	\cmdfifo_gcm_cmd.iv [42], \cmdfifo_gcm_cmd.iv [41], 
	\cmdfifo_gcm_cmd.iv [40], \cmdfifo_gcm_cmd.iv [39], 
	\cmdfifo_gcm_cmd.iv [38], \cmdfifo_gcm_cmd.iv [37], 
	\cmdfifo_gcm_cmd.iv [36], \cmdfifo_gcm_cmd.iv [35], 
	\cmdfifo_gcm_cmd.iv [34], \cmdfifo_gcm_cmd.iv [33], 
	\cmdfifo_gcm_cmd.iv [32], \cmdfifo_gcm_cmd.iv [31], 
	\cmdfifo_gcm_cmd.iv [30], \cmdfifo_gcm_cmd.iv [29], 
	\cmdfifo_gcm_cmd.iv [28], \cmdfifo_gcm_cmd.iv [27], 
	\cmdfifo_gcm_cmd.iv [26], \cmdfifo_gcm_cmd.iv [25], 
	\cmdfifo_gcm_cmd.iv [24], \cmdfifo_gcm_cmd.iv [23], 
	\cmdfifo_gcm_cmd.iv [22], \cmdfifo_gcm_cmd.iv [21], 
	\cmdfifo_gcm_cmd.iv [20], \cmdfifo_gcm_cmd.iv [19], 
	\cmdfifo_gcm_cmd.iv [18], \cmdfifo_gcm_cmd.iv [17], 
	\cmdfifo_gcm_cmd.iv [16], \cmdfifo_gcm_cmd.iv [15], 
	\cmdfifo_gcm_cmd.iv [14], \cmdfifo_gcm_cmd.iv [13], 
	\cmdfifo_gcm_cmd.iv [12], \cmdfifo_gcm_cmd.iv [11], 
	\cmdfifo_gcm_cmd.iv [10], \cmdfifo_gcm_cmd.iv [9], 
	\cmdfifo_gcm_cmd.iv [8], \cmdfifo_gcm_cmd.iv [7], 
	\cmdfifo_gcm_cmd.iv [6], \cmdfifo_gcm_cmd.iv [5], 
	\cmdfifo_gcm_cmd.iv [4], \cmdfifo_gcm_cmd.iv [3], 
	\cmdfifo_gcm_cmd.iv [2], \cmdfifo_gcm_cmd.iv [1], 
	\cmdfifo_gcm_cmd.iv [0], \cmdfifo_gcm_cmd.op [2], 
	\cmdfifo_gcm_cmd.op [1], \cmdfifo_gcm_cmd.op [0]} ), 
	upsizer_gcm_valid, upsizer_gcm_eof, upsizer_gcm_data, 
	gcm_tag_data_out, gcm_tag_data_out_valid, kdf_gcm_stall, 
	gcm_status_data_in_stall);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output set_gcm_tag_fail_int;
output gcm_cmdfifo_ack;
output gcm_upsizer_stall;
output gcm_tag_data_out_ack;
output gcm_kdf_valid;
output gcm_kdf_eof;
output [127:0] gcm_kdf_data;
output gcm_status_data_in_valid;
output [0:0] \gcm_status_data_in.tag_mismatch ;
wire [0:0] gcm_status_data_in;
input clk;
input rst_n;
input cmdfifo_gcm_valid;
input [255:0] \cmdfifo_gcm_cmd.key0 ;
input [255:0] \cmdfifo_gcm_cmd.key1 ;
input [95:0] \cmdfifo_gcm_cmd.iv ;
input [2:0] \cmdfifo_gcm_cmd.op ;
wire [610:0] cmdfifo_gcm_cmd;
input upsizer_gcm_valid;
input upsizer_gcm_eof;
input [127:0] upsizer_gcm_data;
input [95:0] gcm_tag_data_out;
input gcm_tag_data_out_valid;
input kdf_gcm_stall;
input gcm_status_data_in_stall;
wire ciph_in_stall;
wire key_in_stall;
wire [127:0] ciph_out;
wire ciph_out_vld;
wire fifo_in_stall;
wire fifo_out_vld;
wire _zy_simnet_gcm_cmdfifo_ack_0_w$;
wire _zy_simnet_gcm_upsizer_stall_1_w$;
wire _zy_simnet_gcm_tag_data_out_ack_2_w$;
wire _zy_simnet_gcm_kdf_valid_3_w$;
wire _zy_simnet_gcm_kdf_eof_4_w$;
wire [0:127] _zy_simnet_gcm_kdf_data_5_w$;
wire _zy_simnet_gcm_status_data_in_valid_6_w$;
wire _zy_simnet_gcm_status_data_in_7_w$;
wire _zy_simnet_cio_8;
wire _zy_simnet_cio_9;
wire _zy_simnet_cio_10;
wire [0:127] _zy_simnet_ciph_in_11_w$;
wire _zy_simnet_ciph_in_vld_12_w$;
wire _zy_simnet_ciph_in_last_13_w$;
wire _zy_simnet_cio_14;
wire [0:255] _zy_simnet_key_in_15_w$;
wire _zy_simnet_key_in_vld_16_w$;
wire _zy_simnet_ciph_out_stall_17_w$;
wire [0:131] _zy_simnet_fifo_out_18_w$;
wire _zy_simnet_dio_19;
wire _zy_simnet_dio_20;
wire [0:131] _zy_simnet_fifo_in_21_w$;
wire _zy_simnet_fifo_in_vld_22_w$;
wire _zy_simnet_fifo_out_ack_23_w$;
wire _zy_simnet_cio_24;
wire [2:0] cur_state;
wire [2:0] nxt_state;
wire [127:0] ciph_in;
wire ciph_in_vld;
wire ciph_in_last;
wire [255:0] key_in;
wire key_in_vld;
wire ciph_out_stall;
wire [131:0] fifo_in;
wire fifo_in_vld;
wire [131:0] fifo_out;
wire fifo_out_ack;
wire [127:0] iv_counter;
wire [1:0] beat_num;
wire stream_end;
wire ciph_fifo_in_stall;
wire combo_dek512;
wire nxt_combo_dek512;
wire [127:0] operand_X;
wire [127:0] operand_Y;
wire [127:0] mult_out;
wire [127:0] h_value;
wire [127:0] nxt_h_value;
wire [127:0] auth_tag;
wire [127:0] nxt_auth_tag;
supply1 n1;
supply0 n1648;
wire [2:0] \fifo_in.op ;
wire [127:0] \fifo_in.pt ;
wire [0:0] \fifo_in.eof ;
wire [2:0] \fifo_out.op ;
wire [127:0] \fifo_out.pt ;
wire [0:0] \fifo_out.eof ;
tran (gcm_status_data_in[0], \gcm_status_data_in.tag_mismatch [0]);
tran (cmdfifo_gcm_cmd[610], \cmdfifo_gcm_cmd.key0 [255]);
tran (cmdfifo_gcm_cmd[609], \cmdfifo_gcm_cmd.key0 [254]);
tran (cmdfifo_gcm_cmd[608], \cmdfifo_gcm_cmd.key0 [253]);
tran (cmdfifo_gcm_cmd[607], \cmdfifo_gcm_cmd.key0 [252]);
tran (cmdfifo_gcm_cmd[606], \cmdfifo_gcm_cmd.key0 [251]);
tran (cmdfifo_gcm_cmd[605], \cmdfifo_gcm_cmd.key0 [250]);
tran (cmdfifo_gcm_cmd[604], \cmdfifo_gcm_cmd.key0 [249]);
tran (cmdfifo_gcm_cmd[603], \cmdfifo_gcm_cmd.key0 [248]);
tran (cmdfifo_gcm_cmd[602], \cmdfifo_gcm_cmd.key0 [247]);
tran (cmdfifo_gcm_cmd[601], \cmdfifo_gcm_cmd.key0 [246]);
tran (cmdfifo_gcm_cmd[600], \cmdfifo_gcm_cmd.key0 [245]);
tran (cmdfifo_gcm_cmd[599], \cmdfifo_gcm_cmd.key0 [244]);
tran (cmdfifo_gcm_cmd[598], \cmdfifo_gcm_cmd.key0 [243]);
tran (cmdfifo_gcm_cmd[597], \cmdfifo_gcm_cmd.key0 [242]);
tran (cmdfifo_gcm_cmd[596], \cmdfifo_gcm_cmd.key0 [241]);
tran (cmdfifo_gcm_cmd[595], \cmdfifo_gcm_cmd.key0 [240]);
tran (cmdfifo_gcm_cmd[594], \cmdfifo_gcm_cmd.key0 [239]);
tran (cmdfifo_gcm_cmd[593], \cmdfifo_gcm_cmd.key0 [238]);
tran (cmdfifo_gcm_cmd[592], \cmdfifo_gcm_cmd.key0 [237]);
tran (cmdfifo_gcm_cmd[591], \cmdfifo_gcm_cmd.key0 [236]);
tran (cmdfifo_gcm_cmd[590], \cmdfifo_gcm_cmd.key0 [235]);
tran (cmdfifo_gcm_cmd[589], \cmdfifo_gcm_cmd.key0 [234]);
tran (cmdfifo_gcm_cmd[588], \cmdfifo_gcm_cmd.key0 [233]);
tran (cmdfifo_gcm_cmd[587], \cmdfifo_gcm_cmd.key0 [232]);
tran (cmdfifo_gcm_cmd[586], \cmdfifo_gcm_cmd.key0 [231]);
tran (cmdfifo_gcm_cmd[585], \cmdfifo_gcm_cmd.key0 [230]);
tran (cmdfifo_gcm_cmd[584], \cmdfifo_gcm_cmd.key0 [229]);
tran (cmdfifo_gcm_cmd[583], \cmdfifo_gcm_cmd.key0 [228]);
tran (cmdfifo_gcm_cmd[582], \cmdfifo_gcm_cmd.key0 [227]);
tran (cmdfifo_gcm_cmd[581], \cmdfifo_gcm_cmd.key0 [226]);
tran (cmdfifo_gcm_cmd[580], \cmdfifo_gcm_cmd.key0 [225]);
tran (cmdfifo_gcm_cmd[579], \cmdfifo_gcm_cmd.key0 [224]);
tran (cmdfifo_gcm_cmd[578], \cmdfifo_gcm_cmd.key0 [223]);
tran (cmdfifo_gcm_cmd[577], \cmdfifo_gcm_cmd.key0 [222]);
tran (cmdfifo_gcm_cmd[576], \cmdfifo_gcm_cmd.key0 [221]);
tran (cmdfifo_gcm_cmd[575], \cmdfifo_gcm_cmd.key0 [220]);
tran (cmdfifo_gcm_cmd[574], \cmdfifo_gcm_cmd.key0 [219]);
tran (cmdfifo_gcm_cmd[573], \cmdfifo_gcm_cmd.key0 [218]);
tran (cmdfifo_gcm_cmd[572], \cmdfifo_gcm_cmd.key0 [217]);
tran (cmdfifo_gcm_cmd[571], \cmdfifo_gcm_cmd.key0 [216]);
tran (cmdfifo_gcm_cmd[570], \cmdfifo_gcm_cmd.key0 [215]);
tran (cmdfifo_gcm_cmd[569], \cmdfifo_gcm_cmd.key0 [214]);
tran (cmdfifo_gcm_cmd[568], \cmdfifo_gcm_cmd.key0 [213]);
tran (cmdfifo_gcm_cmd[567], \cmdfifo_gcm_cmd.key0 [212]);
tran (cmdfifo_gcm_cmd[566], \cmdfifo_gcm_cmd.key0 [211]);
tran (cmdfifo_gcm_cmd[565], \cmdfifo_gcm_cmd.key0 [210]);
tran (cmdfifo_gcm_cmd[564], \cmdfifo_gcm_cmd.key0 [209]);
tran (cmdfifo_gcm_cmd[563], \cmdfifo_gcm_cmd.key0 [208]);
tran (cmdfifo_gcm_cmd[562], \cmdfifo_gcm_cmd.key0 [207]);
tran (cmdfifo_gcm_cmd[561], \cmdfifo_gcm_cmd.key0 [206]);
tran (cmdfifo_gcm_cmd[560], \cmdfifo_gcm_cmd.key0 [205]);
tran (cmdfifo_gcm_cmd[559], \cmdfifo_gcm_cmd.key0 [204]);
tran (cmdfifo_gcm_cmd[558], \cmdfifo_gcm_cmd.key0 [203]);
tran (cmdfifo_gcm_cmd[557], \cmdfifo_gcm_cmd.key0 [202]);
tran (cmdfifo_gcm_cmd[556], \cmdfifo_gcm_cmd.key0 [201]);
tran (cmdfifo_gcm_cmd[555], \cmdfifo_gcm_cmd.key0 [200]);
tran (cmdfifo_gcm_cmd[554], \cmdfifo_gcm_cmd.key0 [199]);
tran (cmdfifo_gcm_cmd[553], \cmdfifo_gcm_cmd.key0 [198]);
tran (cmdfifo_gcm_cmd[552], \cmdfifo_gcm_cmd.key0 [197]);
tran (cmdfifo_gcm_cmd[551], \cmdfifo_gcm_cmd.key0 [196]);
tran (cmdfifo_gcm_cmd[550], \cmdfifo_gcm_cmd.key0 [195]);
tran (cmdfifo_gcm_cmd[549], \cmdfifo_gcm_cmd.key0 [194]);
tran (cmdfifo_gcm_cmd[548], \cmdfifo_gcm_cmd.key0 [193]);
tran (cmdfifo_gcm_cmd[547], \cmdfifo_gcm_cmd.key0 [192]);
tran (cmdfifo_gcm_cmd[546], \cmdfifo_gcm_cmd.key0 [191]);
tran (cmdfifo_gcm_cmd[545], \cmdfifo_gcm_cmd.key0 [190]);
tran (cmdfifo_gcm_cmd[544], \cmdfifo_gcm_cmd.key0 [189]);
tran (cmdfifo_gcm_cmd[543], \cmdfifo_gcm_cmd.key0 [188]);
tran (cmdfifo_gcm_cmd[542], \cmdfifo_gcm_cmd.key0 [187]);
tran (cmdfifo_gcm_cmd[541], \cmdfifo_gcm_cmd.key0 [186]);
tran (cmdfifo_gcm_cmd[540], \cmdfifo_gcm_cmd.key0 [185]);
tran (cmdfifo_gcm_cmd[539], \cmdfifo_gcm_cmd.key0 [184]);
tran (cmdfifo_gcm_cmd[538], \cmdfifo_gcm_cmd.key0 [183]);
tran (cmdfifo_gcm_cmd[537], \cmdfifo_gcm_cmd.key0 [182]);
tran (cmdfifo_gcm_cmd[536], \cmdfifo_gcm_cmd.key0 [181]);
tran (cmdfifo_gcm_cmd[535], \cmdfifo_gcm_cmd.key0 [180]);
tran (cmdfifo_gcm_cmd[534], \cmdfifo_gcm_cmd.key0 [179]);
tran (cmdfifo_gcm_cmd[533], \cmdfifo_gcm_cmd.key0 [178]);
tran (cmdfifo_gcm_cmd[532], \cmdfifo_gcm_cmd.key0 [177]);
tran (cmdfifo_gcm_cmd[531], \cmdfifo_gcm_cmd.key0 [176]);
tran (cmdfifo_gcm_cmd[530], \cmdfifo_gcm_cmd.key0 [175]);
tran (cmdfifo_gcm_cmd[529], \cmdfifo_gcm_cmd.key0 [174]);
tran (cmdfifo_gcm_cmd[528], \cmdfifo_gcm_cmd.key0 [173]);
tran (cmdfifo_gcm_cmd[527], \cmdfifo_gcm_cmd.key0 [172]);
tran (cmdfifo_gcm_cmd[526], \cmdfifo_gcm_cmd.key0 [171]);
tran (cmdfifo_gcm_cmd[525], \cmdfifo_gcm_cmd.key0 [170]);
tran (cmdfifo_gcm_cmd[524], \cmdfifo_gcm_cmd.key0 [169]);
tran (cmdfifo_gcm_cmd[523], \cmdfifo_gcm_cmd.key0 [168]);
tran (cmdfifo_gcm_cmd[522], \cmdfifo_gcm_cmd.key0 [167]);
tran (cmdfifo_gcm_cmd[521], \cmdfifo_gcm_cmd.key0 [166]);
tran (cmdfifo_gcm_cmd[520], \cmdfifo_gcm_cmd.key0 [165]);
tran (cmdfifo_gcm_cmd[519], \cmdfifo_gcm_cmd.key0 [164]);
tran (cmdfifo_gcm_cmd[518], \cmdfifo_gcm_cmd.key0 [163]);
tran (cmdfifo_gcm_cmd[517], \cmdfifo_gcm_cmd.key0 [162]);
tran (cmdfifo_gcm_cmd[516], \cmdfifo_gcm_cmd.key0 [161]);
tran (cmdfifo_gcm_cmd[515], \cmdfifo_gcm_cmd.key0 [160]);
tran (cmdfifo_gcm_cmd[514], \cmdfifo_gcm_cmd.key0 [159]);
tran (cmdfifo_gcm_cmd[513], \cmdfifo_gcm_cmd.key0 [158]);
tran (cmdfifo_gcm_cmd[512], \cmdfifo_gcm_cmd.key0 [157]);
tran (cmdfifo_gcm_cmd[511], \cmdfifo_gcm_cmd.key0 [156]);
tran (cmdfifo_gcm_cmd[510], \cmdfifo_gcm_cmd.key0 [155]);
tran (cmdfifo_gcm_cmd[509], \cmdfifo_gcm_cmd.key0 [154]);
tran (cmdfifo_gcm_cmd[508], \cmdfifo_gcm_cmd.key0 [153]);
tran (cmdfifo_gcm_cmd[507], \cmdfifo_gcm_cmd.key0 [152]);
tran (cmdfifo_gcm_cmd[506], \cmdfifo_gcm_cmd.key0 [151]);
tran (cmdfifo_gcm_cmd[505], \cmdfifo_gcm_cmd.key0 [150]);
tran (cmdfifo_gcm_cmd[504], \cmdfifo_gcm_cmd.key0 [149]);
tran (cmdfifo_gcm_cmd[503], \cmdfifo_gcm_cmd.key0 [148]);
tran (cmdfifo_gcm_cmd[502], \cmdfifo_gcm_cmd.key0 [147]);
tran (cmdfifo_gcm_cmd[501], \cmdfifo_gcm_cmd.key0 [146]);
tran (cmdfifo_gcm_cmd[500], \cmdfifo_gcm_cmd.key0 [145]);
tran (cmdfifo_gcm_cmd[499], \cmdfifo_gcm_cmd.key0 [144]);
tran (cmdfifo_gcm_cmd[498], \cmdfifo_gcm_cmd.key0 [143]);
tran (cmdfifo_gcm_cmd[497], \cmdfifo_gcm_cmd.key0 [142]);
tran (cmdfifo_gcm_cmd[496], \cmdfifo_gcm_cmd.key0 [141]);
tran (cmdfifo_gcm_cmd[495], \cmdfifo_gcm_cmd.key0 [140]);
tran (cmdfifo_gcm_cmd[494], \cmdfifo_gcm_cmd.key0 [139]);
tran (cmdfifo_gcm_cmd[493], \cmdfifo_gcm_cmd.key0 [138]);
tran (cmdfifo_gcm_cmd[492], \cmdfifo_gcm_cmd.key0 [137]);
tran (cmdfifo_gcm_cmd[491], \cmdfifo_gcm_cmd.key0 [136]);
tran (cmdfifo_gcm_cmd[490], \cmdfifo_gcm_cmd.key0 [135]);
tran (cmdfifo_gcm_cmd[489], \cmdfifo_gcm_cmd.key0 [134]);
tran (cmdfifo_gcm_cmd[488], \cmdfifo_gcm_cmd.key0 [133]);
tran (cmdfifo_gcm_cmd[487], \cmdfifo_gcm_cmd.key0 [132]);
tran (cmdfifo_gcm_cmd[486], \cmdfifo_gcm_cmd.key0 [131]);
tran (cmdfifo_gcm_cmd[485], \cmdfifo_gcm_cmd.key0 [130]);
tran (cmdfifo_gcm_cmd[484], \cmdfifo_gcm_cmd.key0 [129]);
tran (cmdfifo_gcm_cmd[483], \cmdfifo_gcm_cmd.key0 [128]);
tran (cmdfifo_gcm_cmd[482], \cmdfifo_gcm_cmd.key0 [127]);
tran (cmdfifo_gcm_cmd[481], \cmdfifo_gcm_cmd.key0 [126]);
tran (cmdfifo_gcm_cmd[480], \cmdfifo_gcm_cmd.key0 [125]);
tran (cmdfifo_gcm_cmd[479], \cmdfifo_gcm_cmd.key0 [124]);
tran (cmdfifo_gcm_cmd[478], \cmdfifo_gcm_cmd.key0 [123]);
tran (cmdfifo_gcm_cmd[477], \cmdfifo_gcm_cmd.key0 [122]);
tran (cmdfifo_gcm_cmd[476], \cmdfifo_gcm_cmd.key0 [121]);
tran (cmdfifo_gcm_cmd[475], \cmdfifo_gcm_cmd.key0 [120]);
tran (cmdfifo_gcm_cmd[474], \cmdfifo_gcm_cmd.key0 [119]);
tran (cmdfifo_gcm_cmd[473], \cmdfifo_gcm_cmd.key0 [118]);
tran (cmdfifo_gcm_cmd[472], \cmdfifo_gcm_cmd.key0 [117]);
tran (cmdfifo_gcm_cmd[471], \cmdfifo_gcm_cmd.key0 [116]);
tran (cmdfifo_gcm_cmd[470], \cmdfifo_gcm_cmd.key0 [115]);
tran (cmdfifo_gcm_cmd[469], \cmdfifo_gcm_cmd.key0 [114]);
tran (cmdfifo_gcm_cmd[468], \cmdfifo_gcm_cmd.key0 [113]);
tran (cmdfifo_gcm_cmd[467], \cmdfifo_gcm_cmd.key0 [112]);
tran (cmdfifo_gcm_cmd[466], \cmdfifo_gcm_cmd.key0 [111]);
tran (cmdfifo_gcm_cmd[465], \cmdfifo_gcm_cmd.key0 [110]);
tran (cmdfifo_gcm_cmd[464], \cmdfifo_gcm_cmd.key0 [109]);
tran (cmdfifo_gcm_cmd[463], \cmdfifo_gcm_cmd.key0 [108]);
tran (cmdfifo_gcm_cmd[462], \cmdfifo_gcm_cmd.key0 [107]);
tran (cmdfifo_gcm_cmd[461], \cmdfifo_gcm_cmd.key0 [106]);
tran (cmdfifo_gcm_cmd[460], \cmdfifo_gcm_cmd.key0 [105]);
tran (cmdfifo_gcm_cmd[459], \cmdfifo_gcm_cmd.key0 [104]);
tran (cmdfifo_gcm_cmd[458], \cmdfifo_gcm_cmd.key0 [103]);
tran (cmdfifo_gcm_cmd[457], \cmdfifo_gcm_cmd.key0 [102]);
tran (cmdfifo_gcm_cmd[456], \cmdfifo_gcm_cmd.key0 [101]);
tran (cmdfifo_gcm_cmd[455], \cmdfifo_gcm_cmd.key0 [100]);
tran (cmdfifo_gcm_cmd[454], \cmdfifo_gcm_cmd.key0 [99]);
tran (cmdfifo_gcm_cmd[453], \cmdfifo_gcm_cmd.key0 [98]);
tran (cmdfifo_gcm_cmd[452], \cmdfifo_gcm_cmd.key0 [97]);
tran (cmdfifo_gcm_cmd[451], \cmdfifo_gcm_cmd.key0 [96]);
tran (cmdfifo_gcm_cmd[450], \cmdfifo_gcm_cmd.key0 [95]);
tran (cmdfifo_gcm_cmd[449], \cmdfifo_gcm_cmd.key0 [94]);
tran (cmdfifo_gcm_cmd[448], \cmdfifo_gcm_cmd.key0 [93]);
tran (cmdfifo_gcm_cmd[447], \cmdfifo_gcm_cmd.key0 [92]);
tran (cmdfifo_gcm_cmd[446], \cmdfifo_gcm_cmd.key0 [91]);
tran (cmdfifo_gcm_cmd[445], \cmdfifo_gcm_cmd.key0 [90]);
tran (cmdfifo_gcm_cmd[444], \cmdfifo_gcm_cmd.key0 [89]);
tran (cmdfifo_gcm_cmd[443], \cmdfifo_gcm_cmd.key0 [88]);
tran (cmdfifo_gcm_cmd[442], \cmdfifo_gcm_cmd.key0 [87]);
tran (cmdfifo_gcm_cmd[441], \cmdfifo_gcm_cmd.key0 [86]);
tran (cmdfifo_gcm_cmd[440], \cmdfifo_gcm_cmd.key0 [85]);
tran (cmdfifo_gcm_cmd[439], \cmdfifo_gcm_cmd.key0 [84]);
tran (cmdfifo_gcm_cmd[438], \cmdfifo_gcm_cmd.key0 [83]);
tran (cmdfifo_gcm_cmd[437], \cmdfifo_gcm_cmd.key0 [82]);
tran (cmdfifo_gcm_cmd[436], \cmdfifo_gcm_cmd.key0 [81]);
tran (cmdfifo_gcm_cmd[435], \cmdfifo_gcm_cmd.key0 [80]);
tran (cmdfifo_gcm_cmd[434], \cmdfifo_gcm_cmd.key0 [79]);
tran (cmdfifo_gcm_cmd[433], \cmdfifo_gcm_cmd.key0 [78]);
tran (cmdfifo_gcm_cmd[432], \cmdfifo_gcm_cmd.key0 [77]);
tran (cmdfifo_gcm_cmd[431], \cmdfifo_gcm_cmd.key0 [76]);
tran (cmdfifo_gcm_cmd[430], \cmdfifo_gcm_cmd.key0 [75]);
tran (cmdfifo_gcm_cmd[429], \cmdfifo_gcm_cmd.key0 [74]);
tran (cmdfifo_gcm_cmd[428], \cmdfifo_gcm_cmd.key0 [73]);
tran (cmdfifo_gcm_cmd[427], \cmdfifo_gcm_cmd.key0 [72]);
tran (cmdfifo_gcm_cmd[426], \cmdfifo_gcm_cmd.key0 [71]);
tran (cmdfifo_gcm_cmd[425], \cmdfifo_gcm_cmd.key0 [70]);
tran (cmdfifo_gcm_cmd[424], \cmdfifo_gcm_cmd.key0 [69]);
tran (cmdfifo_gcm_cmd[423], \cmdfifo_gcm_cmd.key0 [68]);
tran (cmdfifo_gcm_cmd[422], \cmdfifo_gcm_cmd.key0 [67]);
tran (cmdfifo_gcm_cmd[421], \cmdfifo_gcm_cmd.key0 [66]);
tran (cmdfifo_gcm_cmd[420], \cmdfifo_gcm_cmd.key0 [65]);
tran (cmdfifo_gcm_cmd[419], \cmdfifo_gcm_cmd.key0 [64]);
tran (cmdfifo_gcm_cmd[418], \cmdfifo_gcm_cmd.key0 [63]);
tran (cmdfifo_gcm_cmd[417], \cmdfifo_gcm_cmd.key0 [62]);
tran (cmdfifo_gcm_cmd[416], \cmdfifo_gcm_cmd.key0 [61]);
tran (cmdfifo_gcm_cmd[415], \cmdfifo_gcm_cmd.key0 [60]);
tran (cmdfifo_gcm_cmd[414], \cmdfifo_gcm_cmd.key0 [59]);
tran (cmdfifo_gcm_cmd[413], \cmdfifo_gcm_cmd.key0 [58]);
tran (cmdfifo_gcm_cmd[412], \cmdfifo_gcm_cmd.key0 [57]);
tran (cmdfifo_gcm_cmd[411], \cmdfifo_gcm_cmd.key0 [56]);
tran (cmdfifo_gcm_cmd[410], \cmdfifo_gcm_cmd.key0 [55]);
tran (cmdfifo_gcm_cmd[409], \cmdfifo_gcm_cmd.key0 [54]);
tran (cmdfifo_gcm_cmd[408], \cmdfifo_gcm_cmd.key0 [53]);
tran (cmdfifo_gcm_cmd[407], \cmdfifo_gcm_cmd.key0 [52]);
tran (cmdfifo_gcm_cmd[406], \cmdfifo_gcm_cmd.key0 [51]);
tran (cmdfifo_gcm_cmd[405], \cmdfifo_gcm_cmd.key0 [50]);
tran (cmdfifo_gcm_cmd[404], \cmdfifo_gcm_cmd.key0 [49]);
tran (cmdfifo_gcm_cmd[403], \cmdfifo_gcm_cmd.key0 [48]);
tran (cmdfifo_gcm_cmd[402], \cmdfifo_gcm_cmd.key0 [47]);
tran (cmdfifo_gcm_cmd[401], \cmdfifo_gcm_cmd.key0 [46]);
tran (cmdfifo_gcm_cmd[400], \cmdfifo_gcm_cmd.key0 [45]);
tran (cmdfifo_gcm_cmd[399], \cmdfifo_gcm_cmd.key0 [44]);
tran (cmdfifo_gcm_cmd[398], \cmdfifo_gcm_cmd.key0 [43]);
tran (cmdfifo_gcm_cmd[397], \cmdfifo_gcm_cmd.key0 [42]);
tran (cmdfifo_gcm_cmd[396], \cmdfifo_gcm_cmd.key0 [41]);
tran (cmdfifo_gcm_cmd[395], \cmdfifo_gcm_cmd.key0 [40]);
tran (cmdfifo_gcm_cmd[394], \cmdfifo_gcm_cmd.key0 [39]);
tran (cmdfifo_gcm_cmd[393], \cmdfifo_gcm_cmd.key0 [38]);
tran (cmdfifo_gcm_cmd[392], \cmdfifo_gcm_cmd.key0 [37]);
tran (cmdfifo_gcm_cmd[391], \cmdfifo_gcm_cmd.key0 [36]);
tran (cmdfifo_gcm_cmd[390], \cmdfifo_gcm_cmd.key0 [35]);
tran (cmdfifo_gcm_cmd[389], \cmdfifo_gcm_cmd.key0 [34]);
tran (cmdfifo_gcm_cmd[388], \cmdfifo_gcm_cmd.key0 [33]);
tran (cmdfifo_gcm_cmd[387], \cmdfifo_gcm_cmd.key0 [32]);
tran (cmdfifo_gcm_cmd[386], \cmdfifo_gcm_cmd.key0 [31]);
tran (cmdfifo_gcm_cmd[385], \cmdfifo_gcm_cmd.key0 [30]);
tran (cmdfifo_gcm_cmd[384], \cmdfifo_gcm_cmd.key0 [29]);
tran (cmdfifo_gcm_cmd[383], \cmdfifo_gcm_cmd.key0 [28]);
tran (cmdfifo_gcm_cmd[382], \cmdfifo_gcm_cmd.key0 [27]);
tran (cmdfifo_gcm_cmd[381], \cmdfifo_gcm_cmd.key0 [26]);
tran (cmdfifo_gcm_cmd[380], \cmdfifo_gcm_cmd.key0 [25]);
tran (cmdfifo_gcm_cmd[379], \cmdfifo_gcm_cmd.key0 [24]);
tran (cmdfifo_gcm_cmd[378], \cmdfifo_gcm_cmd.key0 [23]);
tran (cmdfifo_gcm_cmd[377], \cmdfifo_gcm_cmd.key0 [22]);
tran (cmdfifo_gcm_cmd[376], \cmdfifo_gcm_cmd.key0 [21]);
tran (cmdfifo_gcm_cmd[375], \cmdfifo_gcm_cmd.key0 [20]);
tran (cmdfifo_gcm_cmd[374], \cmdfifo_gcm_cmd.key0 [19]);
tran (cmdfifo_gcm_cmd[373], \cmdfifo_gcm_cmd.key0 [18]);
tran (cmdfifo_gcm_cmd[372], \cmdfifo_gcm_cmd.key0 [17]);
tran (cmdfifo_gcm_cmd[371], \cmdfifo_gcm_cmd.key0 [16]);
tran (cmdfifo_gcm_cmd[370], \cmdfifo_gcm_cmd.key0 [15]);
tran (cmdfifo_gcm_cmd[369], \cmdfifo_gcm_cmd.key0 [14]);
tran (cmdfifo_gcm_cmd[368], \cmdfifo_gcm_cmd.key0 [13]);
tran (cmdfifo_gcm_cmd[367], \cmdfifo_gcm_cmd.key0 [12]);
tran (cmdfifo_gcm_cmd[366], \cmdfifo_gcm_cmd.key0 [11]);
tran (cmdfifo_gcm_cmd[365], \cmdfifo_gcm_cmd.key0 [10]);
tran (cmdfifo_gcm_cmd[364], \cmdfifo_gcm_cmd.key0 [9]);
tran (cmdfifo_gcm_cmd[363], \cmdfifo_gcm_cmd.key0 [8]);
tran (cmdfifo_gcm_cmd[362], \cmdfifo_gcm_cmd.key0 [7]);
tran (cmdfifo_gcm_cmd[361], \cmdfifo_gcm_cmd.key0 [6]);
tran (cmdfifo_gcm_cmd[360], \cmdfifo_gcm_cmd.key0 [5]);
tran (cmdfifo_gcm_cmd[359], \cmdfifo_gcm_cmd.key0 [4]);
tran (cmdfifo_gcm_cmd[358], \cmdfifo_gcm_cmd.key0 [3]);
tran (cmdfifo_gcm_cmd[357], \cmdfifo_gcm_cmd.key0 [2]);
tran (cmdfifo_gcm_cmd[356], \cmdfifo_gcm_cmd.key0 [1]);
tran (cmdfifo_gcm_cmd[355], \cmdfifo_gcm_cmd.key0 [0]);
tran (cmdfifo_gcm_cmd[354], \cmdfifo_gcm_cmd.key1 [255]);
tran (cmdfifo_gcm_cmd[353], \cmdfifo_gcm_cmd.key1 [254]);
tran (cmdfifo_gcm_cmd[352], \cmdfifo_gcm_cmd.key1 [253]);
tran (cmdfifo_gcm_cmd[351], \cmdfifo_gcm_cmd.key1 [252]);
tran (cmdfifo_gcm_cmd[350], \cmdfifo_gcm_cmd.key1 [251]);
tran (cmdfifo_gcm_cmd[349], \cmdfifo_gcm_cmd.key1 [250]);
tran (cmdfifo_gcm_cmd[348], \cmdfifo_gcm_cmd.key1 [249]);
tran (cmdfifo_gcm_cmd[347], \cmdfifo_gcm_cmd.key1 [248]);
tran (cmdfifo_gcm_cmd[346], \cmdfifo_gcm_cmd.key1 [247]);
tran (cmdfifo_gcm_cmd[345], \cmdfifo_gcm_cmd.key1 [246]);
tran (cmdfifo_gcm_cmd[344], \cmdfifo_gcm_cmd.key1 [245]);
tran (cmdfifo_gcm_cmd[343], \cmdfifo_gcm_cmd.key1 [244]);
tran (cmdfifo_gcm_cmd[342], \cmdfifo_gcm_cmd.key1 [243]);
tran (cmdfifo_gcm_cmd[341], \cmdfifo_gcm_cmd.key1 [242]);
tran (cmdfifo_gcm_cmd[340], \cmdfifo_gcm_cmd.key1 [241]);
tran (cmdfifo_gcm_cmd[339], \cmdfifo_gcm_cmd.key1 [240]);
tran (cmdfifo_gcm_cmd[338], \cmdfifo_gcm_cmd.key1 [239]);
tran (cmdfifo_gcm_cmd[337], \cmdfifo_gcm_cmd.key1 [238]);
tran (cmdfifo_gcm_cmd[336], \cmdfifo_gcm_cmd.key1 [237]);
tran (cmdfifo_gcm_cmd[335], \cmdfifo_gcm_cmd.key1 [236]);
tran (cmdfifo_gcm_cmd[334], \cmdfifo_gcm_cmd.key1 [235]);
tran (cmdfifo_gcm_cmd[333], \cmdfifo_gcm_cmd.key1 [234]);
tran (cmdfifo_gcm_cmd[332], \cmdfifo_gcm_cmd.key1 [233]);
tran (cmdfifo_gcm_cmd[331], \cmdfifo_gcm_cmd.key1 [232]);
tran (cmdfifo_gcm_cmd[330], \cmdfifo_gcm_cmd.key1 [231]);
tran (cmdfifo_gcm_cmd[329], \cmdfifo_gcm_cmd.key1 [230]);
tran (cmdfifo_gcm_cmd[328], \cmdfifo_gcm_cmd.key1 [229]);
tran (cmdfifo_gcm_cmd[327], \cmdfifo_gcm_cmd.key1 [228]);
tran (cmdfifo_gcm_cmd[326], \cmdfifo_gcm_cmd.key1 [227]);
tran (cmdfifo_gcm_cmd[325], \cmdfifo_gcm_cmd.key1 [226]);
tran (cmdfifo_gcm_cmd[324], \cmdfifo_gcm_cmd.key1 [225]);
tran (cmdfifo_gcm_cmd[323], \cmdfifo_gcm_cmd.key1 [224]);
tran (cmdfifo_gcm_cmd[322], \cmdfifo_gcm_cmd.key1 [223]);
tran (cmdfifo_gcm_cmd[321], \cmdfifo_gcm_cmd.key1 [222]);
tran (cmdfifo_gcm_cmd[320], \cmdfifo_gcm_cmd.key1 [221]);
tran (cmdfifo_gcm_cmd[319], \cmdfifo_gcm_cmd.key1 [220]);
tran (cmdfifo_gcm_cmd[318], \cmdfifo_gcm_cmd.key1 [219]);
tran (cmdfifo_gcm_cmd[317], \cmdfifo_gcm_cmd.key1 [218]);
tran (cmdfifo_gcm_cmd[316], \cmdfifo_gcm_cmd.key1 [217]);
tran (cmdfifo_gcm_cmd[315], \cmdfifo_gcm_cmd.key1 [216]);
tran (cmdfifo_gcm_cmd[314], \cmdfifo_gcm_cmd.key1 [215]);
tran (cmdfifo_gcm_cmd[313], \cmdfifo_gcm_cmd.key1 [214]);
tran (cmdfifo_gcm_cmd[312], \cmdfifo_gcm_cmd.key1 [213]);
tran (cmdfifo_gcm_cmd[311], \cmdfifo_gcm_cmd.key1 [212]);
tran (cmdfifo_gcm_cmd[310], \cmdfifo_gcm_cmd.key1 [211]);
tran (cmdfifo_gcm_cmd[309], \cmdfifo_gcm_cmd.key1 [210]);
tran (cmdfifo_gcm_cmd[308], \cmdfifo_gcm_cmd.key1 [209]);
tran (cmdfifo_gcm_cmd[307], \cmdfifo_gcm_cmd.key1 [208]);
tran (cmdfifo_gcm_cmd[306], \cmdfifo_gcm_cmd.key1 [207]);
tran (cmdfifo_gcm_cmd[305], \cmdfifo_gcm_cmd.key1 [206]);
tran (cmdfifo_gcm_cmd[304], \cmdfifo_gcm_cmd.key1 [205]);
tran (cmdfifo_gcm_cmd[303], \cmdfifo_gcm_cmd.key1 [204]);
tran (cmdfifo_gcm_cmd[302], \cmdfifo_gcm_cmd.key1 [203]);
tran (cmdfifo_gcm_cmd[301], \cmdfifo_gcm_cmd.key1 [202]);
tran (cmdfifo_gcm_cmd[300], \cmdfifo_gcm_cmd.key1 [201]);
tran (cmdfifo_gcm_cmd[299], \cmdfifo_gcm_cmd.key1 [200]);
tran (cmdfifo_gcm_cmd[298], \cmdfifo_gcm_cmd.key1 [199]);
tran (cmdfifo_gcm_cmd[297], \cmdfifo_gcm_cmd.key1 [198]);
tran (cmdfifo_gcm_cmd[296], \cmdfifo_gcm_cmd.key1 [197]);
tran (cmdfifo_gcm_cmd[295], \cmdfifo_gcm_cmd.key1 [196]);
tran (cmdfifo_gcm_cmd[294], \cmdfifo_gcm_cmd.key1 [195]);
tran (cmdfifo_gcm_cmd[293], \cmdfifo_gcm_cmd.key1 [194]);
tran (cmdfifo_gcm_cmd[292], \cmdfifo_gcm_cmd.key1 [193]);
tran (cmdfifo_gcm_cmd[291], \cmdfifo_gcm_cmd.key1 [192]);
tran (cmdfifo_gcm_cmd[290], \cmdfifo_gcm_cmd.key1 [191]);
tran (cmdfifo_gcm_cmd[289], \cmdfifo_gcm_cmd.key1 [190]);
tran (cmdfifo_gcm_cmd[288], \cmdfifo_gcm_cmd.key1 [189]);
tran (cmdfifo_gcm_cmd[287], \cmdfifo_gcm_cmd.key1 [188]);
tran (cmdfifo_gcm_cmd[286], \cmdfifo_gcm_cmd.key1 [187]);
tran (cmdfifo_gcm_cmd[285], \cmdfifo_gcm_cmd.key1 [186]);
tran (cmdfifo_gcm_cmd[284], \cmdfifo_gcm_cmd.key1 [185]);
tran (cmdfifo_gcm_cmd[283], \cmdfifo_gcm_cmd.key1 [184]);
tran (cmdfifo_gcm_cmd[282], \cmdfifo_gcm_cmd.key1 [183]);
tran (cmdfifo_gcm_cmd[281], \cmdfifo_gcm_cmd.key1 [182]);
tran (cmdfifo_gcm_cmd[280], \cmdfifo_gcm_cmd.key1 [181]);
tran (cmdfifo_gcm_cmd[279], \cmdfifo_gcm_cmd.key1 [180]);
tran (cmdfifo_gcm_cmd[278], \cmdfifo_gcm_cmd.key1 [179]);
tran (cmdfifo_gcm_cmd[277], \cmdfifo_gcm_cmd.key1 [178]);
tran (cmdfifo_gcm_cmd[276], \cmdfifo_gcm_cmd.key1 [177]);
tran (cmdfifo_gcm_cmd[275], \cmdfifo_gcm_cmd.key1 [176]);
tran (cmdfifo_gcm_cmd[274], \cmdfifo_gcm_cmd.key1 [175]);
tran (cmdfifo_gcm_cmd[273], \cmdfifo_gcm_cmd.key1 [174]);
tran (cmdfifo_gcm_cmd[272], \cmdfifo_gcm_cmd.key1 [173]);
tran (cmdfifo_gcm_cmd[271], \cmdfifo_gcm_cmd.key1 [172]);
tran (cmdfifo_gcm_cmd[270], \cmdfifo_gcm_cmd.key1 [171]);
tran (cmdfifo_gcm_cmd[269], \cmdfifo_gcm_cmd.key1 [170]);
tran (cmdfifo_gcm_cmd[268], \cmdfifo_gcm_cmd.key1 [169]);
tran (cmdfifo_gcm_cmd[267], \cmdfifo_gcm_cmd.key1 [168]);
tran (cmdfifo_gcm_cmd[266], \cmdfifo_gcm_cmd.key1 [167]);
tran (cmdfifo_gcm_cmd[265], \cmdfifo_gcm_cmd.key1 [166]);
tran (cmdfifo_gcm_cmd[264], \cmdfifo_gcm_cmd.key1 [165]);
tran (cmdfifo_gcm_cmd[263], \cmdfifo_gcm_cmd.key1 [164]);
tran (cmdfifo_gcm_cmd[262], \cmdfifo_gcm_cmd.key1 [163]);
tran (cmdfifo_gcm_cmd[261], \cmdfifo_gcm_cmd.key1 [162]);
tran (cmdfifo_gcm_cmd[260], \cmdfifo_gcm_cmd.key1 [161]);
tran (cmdfifo_gcm_cmd[259], \cmdfifo_gcm_cmd.key1 [160]);
tran (cmdfifo_gcm_cmd[258], \cmdfifo_gcm_cmd.key1 [159]);
tran (cmdfifo_gcm_cmd[257], \cmdfifo_gcm_cmd.key1 [158]);
tran (cmdfifo_gcm_cmd[256], \cmdfifo_gcm_cmd.key1 [157]);
tran (cmdfifo_gcm_cmd[255], \cmdfifo_gcm_cmd.key1 [156]);
tran (cmdfifo_gcm_cmd[254], \cmdfifo_gcm_cmd.key1 [155]);
tran (cmdfifo_gcm_cmd[253], \cmdfifo_gcm_cmd.key1 [154]);
tran (cmdfifo_gcm_cmd[252], \cmdfifo_gcm_cmd.key1 [153]);
tran (cmdfifo_gcm_cmd[251], \cmdfifo_gcm_cmd.key1 [152]);
tran (cmdfifo_gcm_cmd[250], \cmdfifo_gcm_cmd.key1 [151]);
tran (cmdfifo_gcm_cmd[249], \cmdfifo_gcm_cmd.key1 [150]);
tran (cmdfifo_gcm_cmd[248], \cmdfifo_gcm_cmd.key1 [149]);
tran (cmdfifo_gcm_cmd[247], \cmdfifo_gcm_cmd.key1 [148]);
tran (cmdfifo_gcm_cmd[246], \cmdfifo_gcm_cmd.key1 [147]);
tran (cmdfifo_gcm_cmd[245], \cmdfifo_gcm_cmd.key1 [146]);
tran (cmdfifo_gcm_cmd[244], \cmdfifo_gcm_cmd.key1 [145]);
tran (cmdfifo_gcm_cmd[243], \cmdfifo_gcm_cmd.key1 [144]);
tran (cmdfifo_gcm_cmd[242], \cmdfifo_gcm_cmd.key1 [143]);
tran (cmdfifo_gcm_cmd[241], \cmdfifo_gcm_cmd.key1 [142]);
tran (cmdfifo_gcm_cmd[240], \cmdfifo_gcm_cmd.key1 [141]);
tran (cmdfifo_gcm_cmd[239], \cmdfifo_gcm_cmd.key1 [140]);
tran (cmdfifo_gcm_cmd[238], \cmdfifo_gcm_cmd.key1 [139]);
tran (cmdfifo_gcm_cmd[237], \cmdfifo_gcm_cmd.key1 [138]);
tran (cmdfifo_gcm_cmd[236], \cmdfifo_gcm_cmd.key1 [137]);
tran (cmdfifo_gcm_cmd[235], \cmdfifo_gcm_cmd.key1 [136]);
tran (cmdfifo_gcm_cmd[234], \cmdfifo_gcm_cmd.key1 [135]);
tran (cmdfifo_gcm_cmd[233], \cmdfifo_gcm_cmd.key1 [134]);
tran (cmdfifo_gcm_cmd[232], \cmdfifo_gcm_cmd.key1 [133]);
tran (cmdfifo_gcm_cmd[231], \cmdfifo_gcm_cmd.key1 [132]);
tran (cmdfifo_gcm_cmd[230], \cmdfifo_gcm_cmd.key1 [131]);
tran (cmdfifo_gcm_cmd[229], \cmdfifo_gcm_cmd.key1 [130]);
tran (cmdfifo_gcm_cmd[228], \cmdfifo_gcm_cmd.key1 [129]);
tran (cmdfifo_gcm_cmd[227], \cmdfifo_gcm_cmd.key1 [128]);
tran (cmdfifo_gcm_cmd[226], \cmdfifo_gcm_cmd.key1 [127]);
tran (cmdfifo_gcm_cmd[225], \cmdfifo_gcm_cmd.key1 [126]);
tran (cmdfifo_gcm_cmd[224], \cmdfifo_gcm_cmd.key1 [125]);
tran (cmdfifo_gcm_cmd[223], \cmdfifo_gcm_cmd.key1 [124]);
tran (cmdfifo_gcm_cmd[222], \cmdfifo_gcm_cmd.key1 [123]);
tran (cmdfifo_gcm_cmd[221], \cmdfifo_gcm_cmd.key1 [122]);
tran (cmdfifo_gcm_cmd[220], \cmdfifo_gcm_cmd.key1 [121]);
tran (cmdfifo_gcm_cmd[219], \cmdfifo_gcm_cmd.key1 [120]);
tran (cmdfifo_gcm_cmd[218], \cmdfifo_gcm_cmd.key1 [119]);
tran (cmdfifo_gcm_cmd[217], \cmdfifo_gcm_cmd.key1 [118]);
tran (cmdfifo_gcm_cmd[216], \cmdfifo_gcm_cmd.key1 [117]);
tran (cmdfifo_gcm_cmd[215], \cmdfifo_gcm_cmd.key1 [116]);
tran (cmdfifo_gcm_cmd[214], \cmdfifo_gcm_cmd.key1 [115]);
tran (cmdfifo_gcm_cmd[213], \cmdfifo_gcm_cmd.key1 [114]);
tran (cmdfifo_gcm_cmd[212], \cmdfifo_gcm_cmd.key1 [113]);
tran (cmdfifo_gcm_cmd[211], \cmdfifo_gcm_cmd.key1 [112]);
tran (cmdfifo_gcm_cmd[210], \cmdfifo_gcm_cmd.key1 [111]);
tran (cmdfifo_gcm_cmd[209], \cmdfifo_gcm_cmd.key1 [110]);
tran (cmdfifo_gcm_cmd[208], \cmdfifo_gcm_cmd.key1 [109]);
tran (cmdfifo_gcm_cmd[207], \cmdfifo_gcm_cmd.key1 [108]);
tran (cmdfifo_gcm_cmd[206], \cmdfifo_gcm_cmd.key1 [107]);
tran (cmdfifo_gcm_cmd[205], \cmdfifo_gcm_cmd.key1 [106]);
tran (cmdfifo_gcm_cmd[204], \cmdfifo_gcm_cmd.key1 [105]);
tran (cmdfifo_gcm_cmd[203], \cmdfifo_gcm_cmd.key1 [104]);
tran (cmdfifo_gcm_cmd[202], \cmdfifo_gcm_cmd.key1 [103]);
tran (cmdfifo_gcm_cmd[201], \cmdfifo_gcm_cmd.key1 [102]);
tran (cmdfifo_gcm_cmd[200], \cmdfifo_gcm_cmd.key1 [101]);
tran (cmdfifo_gcm_cmd[199], \cmdfifo_gcm_cmd.key1 [100]);
tran (cmdfifo_gcm_cmd[198], \cmdfifo_gcm_cmd.key1 [99]);
tran (cmdfifo_gcm_cmd[197], \cmdfifo_gcm_cmd.key1 [98]);
tran (cmdfifo_gcm_cmd[196], \cmdfifo_gcm_cmd.key1 [97]);
tran (cmdfifo_gcm_cmd[195], \cmdfifo_gcm_cmd.key1 [96]);
tran (cmdfifo_gcm_cmd[194], \cmdfifo_gcm_cmd.key1 [95]);
tran (cmdfifo_gcm_cmd[193], \cmdfifo_gcm_cmd.key1 [94]);
tran (cmdfifo_gcm_cmd[192], \cmdfifo_gcm_cmd.key1 [93]);
tran (cmdfifo_gcm_cmd[191], \cmdfifo_gcm_cmd.key1 [92]);
tran (cmdfifo_gcm_cmd[190], \cmdfifo_gcm_cmd.key1 [91]);
tran (cmdfifo_gcm_cmd[189], \cmdfifo_gcm_cmd.key1 [90]);
tran (cmdfifo_gcm_cmd[188], \cmdfifo_gcm_cmd.key1 [89]);
tran (cmdfifo_gcm_cmd[187], \cmdfifo_gcm_cmd.key1 [88]);
tran (cmdfifo_gcm_cmd[186], \cmdfifo_gcm_cmd.key1 [87]);
tran (cmdfifo_gcm_cmd[185], \cmdfifo_gcm_cmd.key1 [86]);
tran (cmdfifo_gcm_cmd[184], \cmdfifo_gcm_cmd.key1 [85]);
tran (cmdfifo_gcm_cmd[183], \cmdfifo_gcm_cmd.key1 [84]);
tran (cmdfifo_gcm_cmd[182], \cmdfifo_gcm_cmd.key1 [83]);
tran (cmdfifo_gcm_cmd[181], \cmdfifo_gcm_cmd.key1 [82]);
tran (cmdfifo_gcm_cmd[180], \cmdfifo_gcm_cmd.key1 [81]);
tran (cmdfifo_gcm_cmd[179], \cmdfifo_gcm_cmd.key1 [80]);
tran (cmdfifo_gcm_cmd[178], \cmdfifo_gcm_cmd.key1 [79]);
tran (cmdfifo_gcm_cmd[177], \cmdfifo_gcm_cmd.key1 [78]);
tran (cmdfifo_gcm_cmd[176], \cmdfifo_gcm_cmd.key1 [77]);
tran (cmdfifo_gcm_cmd[175], \cmdfifo_gcm_cmd.key1 [76]);
tran (cmdfifo_gcm_cmd[174], \cmdfifo_gcm_cmd.key1 [75]);
tran (cmdfifo_gcm_cmd[173], \cmdfifo_gcm_cmd.key1 [74]);
tran (cmdfifo_gcm_cmd[172], \cmdfifo_gcm_cmd.key1 [73]);
tran (cmdfifo_gcm_cmd[171], \cmdfifo_gcm_cmd.key1 [72]);
tran (cmdfifo_gcm_cmd[170], \cmdfifo_gcm_cmd.key1 [71]);
tran (cmdfifo_gcm_cmd[169], \cmdfifo_gcm_cmd.key1 [70]);
tran (cmdfifo_gcm_cmd[168], \cmdfifo_gcm_cmd.key1 [69]);
tran (cmdfifo_gcm_cmd[167], \cmdfifo_gcm_cmd.key1 [68]);
tran (cmdfifo_gcm_cmd[166], \cmdfifo_gcm_cmd.key1 [67]);
tran (cmdfifo_gcm_cmd[165], \cmdfifo_gcm_cmd.key1 [66]);
tran (cmdfifo_gcm_cmd[164], \cmdfifo_gcm_cmd.key1 [65]);
tran (cmdfifo_gcm_cmd[163], \cmdfifo_gcm_cmd.key1 [64]);
tran (cmdfifo_gcm_cmd[162], \cmdfifo_gcm_cmd.key1 [63]);
tran (cmdfifo_gcm_cmd[161], \cmdfifo_gcm_cmd.key1 [62]);
tran (cmdfifo_gcm_cmd[160], \cmdfifo_gcm_cmd.key1 [61]);
tran (cmdfifo_gcm_cmd[159], \cmdfifo_gcm_cmd.key1 [60]);
tran (cmdfifo_gcm_cmd[158], \cmdfifo_gcm_cmd.key1 [59]);
tran (cmdfifo_gcm_cmd[157], \cmdfifo_gcm_cmd.key1 [58]);
tran (cmdfifo_gcm_cmd[156], \cmdfifo_gcm_cmd.key1 [57]);
tran (cmdfifo_gcm_cmd[155], \cmdfifo_gcm_cmd.key1 [56]);
tran (cmdfifo_gcm_cmd[154], \cmdfifo_gcm_cmd.key1 [55]);
tran (cmdfifo_gcm_cmd[153], \cmdfifo_gcm_cmd.key1 [54]);
tran (cmdfifo_gcm_cmd[152], \cmdfifo_gcm_cmd.key1 [53]);
tran (cmdfifo_gcm_cmd[151], \cmdfifo_gcm_cmd.key1 [52]);
tran (cmdfifo_gcm_cmd[150], \cmdfifo_gcm_cmd.key1 [51]);
tran (cmdfifo_gcm_cmd[149], \cmdfifo_gcm_cmd.key1 [50]);
tran (cmdfifo_gcm_cmd[148], \cmdfifo_gcm_cmd.key1 [49]);
tran (cmdfifo_gcm_cmd[147], \cmdfifo_gcm_cmd.key1 [48]);
tran (cmdfifo_gcm_cmd[146], \cmdfifo_gcm_cmd.key1 [47]);
tran (cmdfifo_gcm_cmd[145], \cmdfifo_gcm_cmd.key1 [46]);
tran (cmdfifo_gcm_cmd[144], \cmdfifo_gcm_cmd.key1 [45]);
tran (cmdfifo_gcm_cmd[143], \cmdfifo_gcm_cmd.key1 [44]);
tran (cmdfifo_gcm_cmd[142], \cmdfifo_gcm_cmd.key1 [43]);
tran (cmdfifo_gcm_cmd[141], \cmdfifo_gcm_cmd.key1 [42]);
tran (cmdfifo_gcm_cmd[140], \cmdfifo_gcm_cmd.key1 [41]);
tran (cmdfifo_gcm_cmd[139], \cmdfifo_gcm_cmd.key1 [40]);
tran (cmdfifo_gcm_cmd[138], \cmdfifo_gcm_cmd.key1 [39]);
tran (cmdfifo_gcm_cmd[137], \cmdfifo_gcm_cmd.key1 [38]);
tran (cmdfifo_gcm_cmd[136], \cmdfifo_gcm_cmd.key1 [37]);
tran (cmdfifo_gcm_cmd[135], \cmdfifo_gcm_cmd.key1 [36]);
tran (cmdfifo_gcm_cmd[134], \cmdfifo_gcm_cmd.key1 [35]);
tran (cmdfifo_gcm_cmd[133], \cmdfifo_gcm_cmd.key1 [34]);
tran (cmdfifo_gcm_cmd[132], \cmdfifo_gcm_cmd.key1 [33]);
tran (cmdfifo_gcm_cmd[131], \cmdfifo_gcm_cmd.key1 [32]);
tran (cmdfifo_gcm_cmd[130], \cmdfifo_gcm_cmd.key1 [31]);
tran (cmdfifo_gcm_cmd[129], \cmdfifo_gcm_cmd.key1 [30]);
tran (cmdfifo_gcm_cmd[128], \cmdfifo_gcm_cmd.key1 [29]);
tran (cmdfifo_gcm_cmd[127], \cmdfifo_gcm_cmd.key1 [28]);
tran (cmdfifo_gcm_cmd[126], \cmdfifo_gcm_cmd.key1 [27]);
tran (cmdfifo_gcm_cmd[125], \cmdfifo_gcm_cmd.key1 [26]);
tran (cmdfifo_gcm_cmd[124], \cmdfifo_gcm_cmd.key1 [25]);
tran (cmdfifo_gcm_cmd[123], \cmdfifo_gcm_cmd.key1 [24]);
tran (cmdfifo_gcm_cmd[122], \cmdfifo_gcm_cmd.key1 [23]);
tran (cmdfifo_gcm_cmd[121], \cmdfifo_gcm_cmd.key1 [22]);
tran (cmdfifo_gcm_cmd[120], \cmdfifo_gcm_cmd.key1 [21]);
tran (cmdfifo_gcm_cmd[119], \cmdfifo_gcm_cmd.key1 [20]);
tran (cmdfifo_gcm_cmd[118], \cmdfifo_gcm_cmd.key1 [19]);
tran (cmdfifo_gcm_cmd[117], \cmdfifo_gcm_cmd.key1 [18]);
tran (cmdfifo_gcm_cmd[116], \cmdfifo_gcm_cmd.key1 [17]);
tran (cmdfifo_gcm_cmd[115], \cmdfifo_gcm_cmd.key1 [16]);
tran (cmdfifo_gcm_cmd[114], \cmdfifo_gcm_cmd.key1 [15]);
tran (cmdfifo_gcm_cmd[113], \cmdfifo_gcm_cmd.key1 [14]);
tran (cmdfifo_gcm_cmd[112], \cmdfifo_gcm_cmd.key1 [13]);
tran (cmdfifo_gcm_cmd[111], \cmdfifo_gcm_cmd.key1 [12]);
tran (cmdfifo_gcm_cmd[110], \cmdfifo_gcm_cmd.key1 [11]);
tran (cmdfifo_gcm_cmd[109], \cmdfifo_gcm_cmd.key1 [10]);
tran (cmdfifo_gcm_cmd[108], \cmdfifo_gcm_cmd.key1 [9]);
tran (cmdfifo_gcm_cmd[107], \cmdfifo_gcm_cmd.key1 [8]);
tran (cmdfifo_gcm_cmd[106], \cmdfifo_gcm_cmd.key1 [7]);
tran (cmdfifo_gcm_cmd[105], \cmdfifo_gcm_cmd.key1 [6]);
tran (cmdfifo_gcm_cmd[104], \cmdfifo_gcm_cmd.key1 [5]);
tran (cmdfifo_gcm_cmd[103], \cmdfifo_gcm_cmd.key1 [4]);
tran (cmdfifo_gcm_cmd[102], \cmdfifo_gcm_cmd.key1 [3]);
tran (cmdfifo_gcm_cmd[101], \cmdfifo_gcm_cmd.key1 [2]);
tran (cmdfifo_gcm_cmd[100], \cmdfifo_gcm_cmd.key1 [1]);
tran (cmdfifo_gcm_cmd[99], \cmdfifo_gcm_cmd.key1 [0]);
tran (cmdfifo_gcm_cmd[98], \cmdfifo_gcm_cmd.iv [95]);
tran (cmdfifo_gcm_cmd[97], \cmdfifo_gcm_cmd.iv [94]);
tran (cmdfifo_gcm_cmd[96], \cmdfifo_gcm_cmd.iv [93]);
tran (cmdfifo_gcm_cmd[95], \cmdfifo_gcm_cmd.iv [92]);
tran (cmdfifo_gcm_cmd[94], \cmdfifo_gcm_cmd.iv [91]);
tran (cmdfifo_gcm_cmd[93], \cmdfifo_gcm_cmd.iv [90]);
tran (cmdfifo_gcm_cmd[92], \cmdfifo_gcm_cmd.iv [89]);
tran (cmdfifo_gcm_cmd[91], \cmdfifo_gcm_cmd.iv [88]);
tran (cmdfifo_gcm_cmd[90], \cmdfifo_gcm_cmd.iv [87]);
tran (cmdfifo_gcm_cmd[89], \cmdfifo_gcm_cmd.iv [86]);
tran (cmdfifo_gcm_cmd[88], \cmdfifo_gcm_cmd.iv [85]);
tran (cmdfifo_gcm_cmd[87], \cmdfifo_gcm_cmd.iv [84]);
tran (cmdfifo_gcm_cmd[86], \cmdfifo_gcm_cmd.iv [83]);
tran (cmdfifo_gcm_cmd[85], \cmdfifo_gcm_cmd.iv [82]);
tran (cmdfifo_gcm_cmd[84], \cmdfifo_gcm_cmd.iv [81]);
tran (cmdfifo_gcm_cmd[83], \cmdfifo_gcm_cmd.iv [80]);
tran (cmdfifo_gcm_cmd[82], \cmdfifo_gcm_cmd.iv [79]);
tran (cmdfifo_gcm_cmd[81], \cmdfifo_gcm_cmd.iv [78]);
tran (cmdfifo_gcm_cmd[80], \cmdfifo_gcm_cmd.iv [77]);
tran (cmdfifo_gcm_cmd[79], \cmdfifo_gcm_cmd.iv [76]);
tran (cmdfifo_gcm_cmd[78], \cmdfifo_gcm_cmd.iv [75]);
tran (cmdfifo_gcm_cmd[77], \cmdfifo_gcm_cmd.iv [74]);
tran (cmdfifo_gcm_cmd[76], \cmdfifo_gcm_cmd.iv [73]);
tran (cmdfifo_gcm_cmd[75], \cmdfifo_gcm_cmd.iv [72]);
tran (cmdfifo_gcm_cmd[74], \cmdfifo_gcm_cmd.iv [71]);
tran (cmdfifo_gcm_cmd[73], \cmdfifo_gcm_cmd.iv [70]);
tran (cmdfifo_gcm_cmd[72], \cmdfifo_gcm_cmd.iv [69]);
tran (cmdfifo_gcm_cmd[71], \cmdfifo_gcm_cmd.iv [68]);
tran (cmdfifo_gcm_cmd[70], \cmdfifo_gcm_cmd.iv [67]);
tran (cmdfifo_gcm_cmd[69], \cmdfifo_gcm_cmd.iv [66]);
tran (cmdfifo_gcm_cmd[68], \cmdfifo_gcm_cmd.iv [65]);
tran (cmdfifo_gcm_cmd[67], \cmdfifo_gcm_cmd.iv [64]);
tran (cmdfifo_gcm_cmd[66], \cmdfifo_gcm_cmd.iv [63]);
tran (cmdfifo_gcm_cmd[65], \cmdfifo_gcm_cmd.iv [62]);
tran (cmdfifo_gcm_cmd[64], \cmdfifo_gcm_cmd.iv [61]);
tran (cmdfifo_gcm_cmd[63], \cmdfifo_gcm_cmd.iv [60]);
tran (cmdfifo_gcm_cmd[62], \cmdfifo_gcm_cmd.iv [59]);
tran (cmdfifo_gcm_cmd[61], \cmdfifo_gcm_cmd.iv [58]);
tran (cmdfifo_gcm_cmd[60], \cmdfifo_gcm_cmd.iv [57]);
tran (cmdfifo_gcm_cmd[59], \cmdfifo_gcm_cmd.iv [56]);
tran (cmdfifo_gcm_cmd[58], \cmdfifo_gcm_cmd.iv [55]);
tran (cmdfifo_gcm_cmd[57], \cmdfifo_gcm_cmd.iv [54]);
tran (cmdfifo_gcm_cmd[56], \cmdfifo_gcm_cmd.iv [53]);
tran (cmdfifo_gcm_cmd[55], \cmdfifo_gcm_cmd.iv [52]);
tran (cmdfifo_gcm_cmd[54], \cmdfifo_gcm_cmd.iv [51]);
tran (cmdfifo_gcm_cmd[53], \cmdfifo_gcm_cmd.iv [50]);
tran (cmdfifo_gcm_cmd[52], \cmdfifo_gcm_cmd.iv [49]);
tran (cmdfifo_gcm_cmd[51], \cmdfifo_gcm_cmd.iv [48]);
tran (cmdfifo_gcm_cmd[50], \cmdfifo_gcm_cmd.iv [47]);
tran (cmdfifo_gcm_cmd[49], \cmdfifo_gcm_cmd.iv [46]);
tran (cmdfifo_gcm_cmd[48], \cmdfifo_gcm_cmd.iv [45]);
tran (cmdfifo_gcm_cmd[47], \cmdfifo_gcm_cmd.iv [44]);
tran (cmdfifo_gcm_cmd[46], \cmdfifo_gcm_cmd.iv [43]);
tran (cmdfifo_gcm_cmd[45], \cmdfifo_gcm_cmd.iv [42]);
tran (cmdfifo_gcm_cmd[44], \cmdfifo_gcm_cmd.iv [41]);
tran (cmdfifo_gcm_cmd[43], \cmdfifo_gcm_cmd.iv [40]);
tran (cmdfifo_gcm_cmd[42], \cmdfifo_gcm_cmd.iv [39]);
tran (cmdfifo_gcm_cmd[41], \cmdfifo_gcm_cmd.iv [38]);
tran (cmdfifo_gcm_cmd[40], \cmdfifo_gcm_cmd.iv [37]);
tran (cmdfifo_gcm_cmd[39], \cmdfifo_gcm_cmd.iv [36]);
tran (cmdfifo_gcm_cmd[38], \cmdfifo_gcm_cmd.iv [35]);
tran (cmdfifo_gcm_cmd[37], \cmdfifo_gcm_cmd.iv [34]);
tran (cmdfifo_gcm_cmd[36], \cmdfifo_gcm_cmd.iv [33]);
tran (cmdfifo_gcm_cmd[35], \cmdfifo_gcm_cmd.iv [32]);
tran (cmdfifo_gcm_cmd[34], \cmdfifo_gcm_cmd.iv [31]);
tran (cmdfifo_gcm_cmd[33], \cmdfifo_gcm_cmd.iv [30]);
tran (cmdfifo_gcm_cmd[32], \cmdfifo_gcm_cmd.iv [29]);
tran (cmdfifo_gcm_cmd[31], \cmdfifo_gcm_cmd.iv [28]);
tran (cmdfifo_gcm_cmd[30], \cmdfifo_gcm_cmd.iv [27]);
tran (cmdfifo_gcm_cmd[29], \cmdfifo_gcm_cmd.iv [26]);
tran (cmdfifo_gcm_cmd[28], \cmdfifo_gcm_cmd.iv [25]);
tran (cmdfifo_gcm_cmd[27], \cmdfifo_gcm_cmd.iv [24]);
tran (cmdfifo_gcm_cmd[26], \cmdfifo_gcm_cmd.iv [23]);
tran (cmdfifo_gcm_cmd[25], \cmdfifo_gcm_cmd.iv [22]);
tran (cmdfifo_gcm_cmd[24], \cmdfifo_gcm_cmd.iv [21]);
tran (cmdfifo_gcm_cmd[23], \cmdfifo_gcm_cmd.iv [20]);
tran (cmdfifo_gcm_cmd[22], \cmdfifo_gcm_cmd.iv [19]);
tran (cmdfifo_gcm_cmd[21], \cmdfifo_gcm_cmd.iv [18]);
tran (cmdfifo_gcm_cmd[20], \cmdfifo_gcm_cmd.iv [17]);
tran (cmdfifo_gcm_cmd[19], \cmdfifo_gcm_cmd.iv [16]);
tran (cmdfifo_gcm_cmd[18], \cmdfifo_gcm_cmd.iv [15]);
tran (cmdfifo_gcm_cmd[17], \cmdfifo_gcm_cmd.iv [14]);
tran (cmdfifo_gcm_cmd[16], \cmdfifo_gcm_cmd.iv [13]);
tran (cmdfifo_gcm_cmd[15], \cmdfifo_gcm_cmd.iv [12]);
tran (cmdfifo_gcm_cmd[14], \cmdfifo_gcm_cmd.iv [11]);
tran (cmdfifo_gcm_cmd[13], \cmdfifo_gcm_cmd.iv [10]);
tran (cmdfifo_gcm_cmd[12], \cmdfifo_gcm_cmd.iv [9]);
tran (cmdfifo_gcm_cmd[11], \cmdfifo_gcm_cmd.iv [8]);
tran (cmdfifo_gcm_cmd[10], \cmdfifo_gcm_cmd.iv [7]);
tran (cmdfifo_gcm_cmd[9], \cmdfifo_gcm_cmd.iv [6]);
tran (cmdfifo_gcm_cmd[8], \cmdfifo_gcm_cmd.iv [5]);
tran (cmdfifo_gcm_cmd[7], \cmdfifo_gcm_cmd.iv [4]);
tran (cmdfifo_gcm_cmd[6], \cmdfifo_gcm_cmd.iv [3]);
tran (cmdfifo_gcm_cmd[5], \cmdfifo_gcm_cmd.iv [2]);
tran (cmdfifo_gcm_cmd[4], \cmdfifo_gcm_cmd.iv [1]);
tran (cmdfifo_gcm_cmd[3], \cmdfifo_gcm_cmd.iv [0]);
tran (cmdfifo_gcm_cmd[2], \cmdfifo_gcm_cmd.op [2]);
tran (cmdfifo_gcm_cmd[1], \cmdfifo_gcm_cmd.op [1]);
tran (cmdfifo_gcm_cmd[0], \cmdfifo_gcm_cmd.op [0]);
tran (fifo_in[130], \fifo_in.op [1]);
tran (fifo_in[0], \fifo_in.eof [0]);
tran (fifo_in[1], \fifo_in.pt [0]);
tran (fifo_in[2], \fifo_in.pt [1]);
tran (fifo_in[3], \fifo_in.pt [2]);
tran (fifo_in[4], \fifo_in.pt [3]);
tran (fifo_in[5], \fifo_in.pt [4]);
tran (fifo_in[6], \fifo_in.pt [5]);
tran (fifo_in[7], \fifo_in.pt [6]);
tran (fifo_in[8], \fifo_in.pt [7]);
tran (fifo_in[9], \fifo_in.pt [8]);
tran (fifo_in[10], \fifo_in.pt [9]);
tran (fifo_in[11], \fifo_in.pt [10]);
tran (fifo_in[12], \fifo_in.pt [11]);
tran (fifo_in[13], \fifo_in.pt [12]);
tran (fifo_in[14], \fifo_in.pt [13]);
tran (fifo_in[15], \fifo_in.pt [14]);
tran (fifo_in[16], \fifo_in.pt [15]);
tran (fifo_in[17], \fifo_in.pt [16]);
tran (fifo_in[18], \fifo_in.pt [17]);
tran (fifo_in[19], \fifo_in.pt [18]);
tran (fifo_in[20], \fifo_in.pt [19]);
tran (fifo_in[21], \fifo_in.pt [20]);
tran (fifo_in[22], \fifo_in.pt [21]);
tran (fifo_in[23], \fifo_in.pt [22]);
tran (fifo_in[24], \fifo_in.pt [23]);
tran (fifo_in[25], \fifo_in.pt [24]);
tran (fifo_in[26], \fifo_in.pt [25]);
tran (fifo_in[27], \fifo_in.pt [26]);
tran (fifo_in[28], \fifo_in.pt [27]);
tran (fifo_in[29], \fifo_in.pt [28]);
tran (fifo_in[30], \fifo_in.pt [29]);
tran (fifo_in[31], \fifo_in.pt [30]);
tran (fifo_in[32], \fifo_in.pt [31]);
tran (fifo_in[33], \fifo_in.pt [32]);
tran (fifo_in[34], \fifo_in.pt [33]);
tran (fifo_in[35], \fifo_in.pt [34]);
tran (fifo_in[36], \fifo_in.pt [35]);
tran (fifo_in[37], \fifo_in.pt [36]);
tran (fifo_in[38], \fifo_in.pt [37]);
tran (fifo_in[39], \fifo_in.pt [38]);
tran (fifo_in[40], \fifo_in.pt [39]);
tran (fifo_in[41], \fifo_in.pt [40]);
tran (fifo_in[42], \fifo_in.pt [41]);
tran (fifo_in[43], \fifo_in.pt [42]);
tran (fifo_in[44], \fifo_in.pt [43]);
tran (fifo_in[45], \fifo_in.pt [44]);
tran (fifo_in[46], \fifo_in.pt [45]);
tran (fifo_in[47], \fifo_in.pt [46]);
tran (fifo_in[48], \fifo_in.pt [47]);
tran (fifo_in[49], \fifo_in.pt [48]);
tran (fifo_in[50], \fifo_in.pt [49]);
tran (fifo_in[51], \fifo_in.pt [50]);
tran (fifo_in[52], \fifo_in.pt [51]);
tran (fifo_in[53], \fifo_in.pt [52]);
tran (fifo_in[54], \fifo_in.pt [53]);
tran (fifo_in[55], \fifo_in.pt [54]);
tran (fifo_in[56], \fifo_in.pt [55]);
tran (fifo_in[57], \fifo_in.pt [56]);
tran (fifo_in[58], \fifo_in.pt [57]);
tran (fifo_in[59], \fifo_in.pt [58]);
tran (fifo_in[60], \fifo_in.pt [59]);
tran (fifo_in[61], \fifo_in.pt [60]);
tran (fifo_in[62], \fifo_in.pt [61]);
tran (fifo_in[63], \fifo_in.pt [62]);
tran (fifo_in[64], \fifo_in.pt [63]);
tran (fifo_in[65], \fifo_in.pt [64]);
tran (fifo_in[66], \fifo_in.pt [65]);
tran (fifo_in[67], \fifo_in.pt [66]);
tran (fifo_in[68], \fifo_in.pt [67]);
tran (fifo_in[69], \fifo_in.pt [68]);
tran (fifo_in[70], \fifo_in.pt [69]);
tran (fifo_in[71], \fifo_in.pt [70]);
tran (fifo_in[72], \fifo_in.pt [71]);
tran (fifo_in[73], \fifo_in.pt [72]);
tran (fifo_in[74], \fifo_in.pt [73]);
tran (fifo_in[75], \fifo_in.pt [74]);
tran (fifo_in[76], \fifo_in.pt [75]);
tran (fifo_in[77], \fifo_in.pt [76]);
tran (fifo_in[78], \fifo_in.pt [77]);
tran (fifo_in[79], \fifo_in.pt [78]);
tran (fifo_in[80], \fifo_in.pt [79]);
tran (fifo_in[81], \fifo_in.pt [80]);
tran (fifo_in[82], \fifo_in.pt [81]);
tran (fifo_in[83], \fifo_in.pt [82]);
tran (fifo_in[84], \fifo_in.pt [83]);
tran (fifo_in[85], \fifo_in.pt [84]);
tran (fifo_in[86], \fifo_in.pt [85]);
tran (fifo_in[87], \fifo_in.pt [86]);
tran (fifo_in[88], \fifo_in.pt [87]);
tran (fifo_in[89], \fifo_in.pt [88]);
tran (fifo_in[90], \fifo_in.pt [89]);
tran (fifo_in[91], \fifo_in.pt [90]);
tran (fifo_in[92], \fifo_in.pt [91]);
tran (fifo_in[93], \fifo_in.pt [92]);
tran (fifo_in[94], \fifo_in.pt [93]);
tran (fifo_in[95], \fifo_in.pt [94]);
tran (fifo_in[96], \fifo_in.pt [95]);
tran (fifo_in[97], \fifo_in.pt [96]);
tran (fifo_in[98], \fifo_in.pt [97]);
tran (fifo_in[99], \fifo_in.pt [98]);
tran (fifo_in[100], \fifo_in.pt [99]);
tran (fifo_in[101], \fifo_in.pt [100]);
tran (fifo_in[102], \fifo_in.pt [101]);
tran (fifo_in[103], \fifo_in.pt [102]);
tran (fifo_in[104], \fifo_in.pt [103]);
tran (fifo_in[105], \fifo_in.pt [104]);
tran (fifo_in[106], \fifo_in.pt [105]);
tran (fifo_in[107], \fifo_in.pt [106]);
tran (fifo_in[108], \fifo_in.pt [107]);
tran (fifo_in[109], \fifo_in.pt [108]);
tran (fifo_in[110], \fifo_in.pt [109]);
tran (fifo_in[111], \fifo_in.pt [110]);
tran (fifo_in[112], \fifo_in.pt [111]);
tran (fifo_in[113], \fifo_in.pt [112]);
tran (fifo_in[114], \fifo_in.pt [113]);
tran (fifo_in[115], \fifo_in.pt [114]);
tran (fifo_in[116], \fifo_in.pt [115]);
tran (fifo_in[117], \fifo_in.pt [116]);
tran (fifo_in[118], \fifo_in.pt [117]);
tran (fifo_in[119], \fifo_in.pt [118]);
tran (fifo_in[120], \fifo_in.pt [119]);
tran (fifo_in[121], \fifo_in.pt [120]);
tran (fifo_in[122], \fifo_in.pt [121]);
tran (fifo_in[123], \fifo_in.pt [122]);
tran (fifo_in[124], \fifo_in.pt [123]);
tran (fifo_in[125], \fifo_in.pt [124]);
tran (fifo_in[126], \fifo_in.pt [125]);
tran (fifo_in[127], \fifo_in.pt [126]);
tran (fifo_in[128], \fifo_in.pt [127]);
tran (fifo_in[129], \fifo_in.op [0]);
tran (fifo_in[131], \fifo_in.op [2]);
tran (fifo_out[0], \fifo_out.eof [0]);
tran (fifo_out[1], \fifo_out.pt [0]);
tran (fifo_out[2], \fifo_out.pt [1]);
tran (fifo_out[3], \fifo_out.pt [2]);
tran (fifo_out[4], \fifo_out.pt [3]);
tran (fifo_out[5], \fifo_out.pt [4]);
tran (fifo_out[6], \fifo_out.pt [5]);
tran (fifo_out[7], \fifo_out.pt [6]);
tran (fifo_out[8], \fifo_out.pt [7]);
tran (fifo_out[9], \fifo_out.pt [8]);
tran (fifo_out[10], \fifo_out.pt [9]);
tran (fifo_out[11], \fifo_out.pt [10]);
tran (fifo_out[12], \fifo_out.pt [11]);
tran (fifo_out[13], \fifo_out.pt [12]);
tran (fifo_out[14], \fifo_out.pt [13]);
tran (fifo_out[15], \fifo_out.pt [14]);
tran (fifo_out[16], \fifo_out.pt [15]);
tran (fifo_out[17], \fifo_out.pt [16]);
tran (fifo_out[18], \fifo_out.pt [17]);
tran (fifo_out[19], \fifo_out.pt [18]);
tran (fifo_out[20], \fifo_out.pt [19]);
tran (fifo_out[21], \fifo_out.pt [20]);
tran (fifo_out[22], \fifo_out.pt [21]);
tran (fifo_out[23], \fifo_out.pt [22]);
tran (fifo_out[24], \fifo_out.pt [23]);
tran (fifo_out[25], \fifo_out.pt [24]);
tran (fifo_out[26], \fifo_out.pt [25]);
tran (fifo_out[27], \fifo_out.pt [26]);
tran (fifo_out[28], \fifo_out.pt [27]);
tran (fifo_out[29], \fifo_out.pt [28]);
tran (fifo_out[30], \fifo_out.pt [29]);
tran (fifo_out[31], \fifo_out.pt [30]);
tran (fifo_out[32], \fifo_out.pt [31]);
tran (fifo_out[33], \fifo_out.pt [32]);
tran (fifo_out[34], \fifo_out.pt [33]);
tran (fifo_out[35], \fifo_out.pt [34]);
tran (fifo_out[36], \fifo_out.pt [35]);
tran (fifo_out[37], \fifo_out.pt [36]);
tran (fifo_out[38], \fifo_out.pt [37]);
tran (fifo_out[39], \fifo_out.pt [38]);
tran (fifo_out[40], \fifo_out.pt [39]);
tran (fifo_out[41], \fifo_out.pt [40]);
tran (fifo_out[42], \fifo_out.pt [41]);
tran (fifo_out[43], \fifo_out.pt [42]);
tran (fifo_out[44], \fifo_out.pt [43]);
tran (fifo_out[45], \fifo_out.pt [44]);
tran (fifo_out[46], \fifo_out.pt [45]);
tran (fifo_out[47], \fifo_out.pt [46]);
tran (fifo_out[48], \fifo_out.pt [47]);
tran (fifo_out[49], \fifo_out.pt [48]);
tran (fifo_out[50], \fifo_out.pt [49]);
tran (fifo_out[51], \fifo_out.pt [50]);
tran (fifo_out[52], \fifo_out.pt [51]);
tran (fifo_out[53], \fifo_out.pt [52]);
tran (fifo_out[54], \fifo_out.pt [53]);
tran (fifo_out[55], \fifo_out.pt [54]);
tran (fifo_out[56], \fifo_out.pt [55]);
tran (fifo_out[57], \fifo_out.pt [56]);
tran (fifo_out[58], \fifo_out.pt [57]);
tran (fifo_out[59], \fifo_out.pt [58]);
tran (fifo_out[60], \fifo_out.pt [59]);
tran (fifo_out[61], \fifo_out.pt [60]);
tran (fifo_out[62], \fifo_out.pt [61]);
tran (fifo_out[63], \fifo_out.pt [62]);
tran (fifo_out[64], \fifo_out.pt [63]);
tran (fifo_out[65], \fifo_out.pt [64]);
tran (fifo_out[66], \fifo_out.pt [65]);
tran (fifo_out[67], \fifo_out.pt [66]);
tran (fifo_out[68], \fifo_out.pt [67]);
tran (fifo_out[69], \fifo_out.pt [68]);
tran (fifo_out[70], \fifo_out.pt [69]);
tran (fifo_out[71], \fifo_out.pt [70]);
tran (fifo_out[72], \fifo_out.pt [71]);
tran (fifo_out[73], \fifo_out.pt [72]);
tran (fifo_out[74], \fifo_out.pt [73]);
tran (fifo_out[75], \fifo_out.pt [74]);
tran (fifo_out[76], \fifo_out.pt [75]);
tran (fifo_out[77], \fifo_out.pt [76]);
tran (fifo_out[78], \fifo_out.pt [77]);
tran (fifo_out[79], \fifo_out.pt [78]);
tran (fifo_out[80], \fifo_out.pt [79]);
tran (fifo_out[81], \fifo_out.pt [80]);
tran (fifo_out[82], \fifo_out.pt [81]);
tran (fifo_out[83], \fifo_out.pt [82]);
tran (fifo_out[84], \fifo_out.pt [83]);
tran (fifo_out[85], \fifo_out.pt [84]);
tran (fifo_out[86], \fifo_out.pt [85]);
tran (fifo_out[87], \fifo_out.pt [86]);
tran (fifo_out[88], \fifo_out.pt [87]);
tran (fifo_out[89], \fifo_out.pt [88]);
tran (fifo_out[90], \fifo_out.pt [89]);
tran (fifo_out[91], \fifo_out.pt [90]);
tran (fifo_out[92], \fifo_out.pt [91]);
tran (fifo_out[93], \fifo_out.pt [92]);
tran (fifo_out[94], \fifo_out.pt [93]);
tran (fifo_out[95], \fifo_out.pt [94]);
tran (fifo_out[96], \fifo_out.pt [95]);
tran (fifo_out[97], \fifo_out.pt [96]);
tran (fifo_out[98], \fifo_out.pt [97]);
tran (fifo_out[99], \fifo_out.pt [98]);
tran (fifo_out[100], \fifo_out.pt [99]);
tran (fifo_out[101], \fifo_out.pt [100]);
tran (fifo_out[102], \fifo_out.pt [101]);
tran (fifo_out[103], \fifo_out.pt [102]);
tran (fifo_out[104], \fifo_out.pt [103]);
tran (fifo_out[105], \fifo_out.pt [104]);
tran (fifo_out[106], \fifo_out.pt [105]);
tran (fifo_out[107], \fifo_out.pt [106]);
tran (fifo_out[108], \fifo_out.pt [107]);
tran (fifo_out[109], \fifo_out.pt [108]);
tran (fifo_out[110], \fifo_out.pt [109]);
tran (fifo_out[111], \fifo_out.pt [110]);
tran (fifo_out[112], \fifo_out.pt [111]);
tran (fifo_out[113], \fifo_out.pt [112]);
tran (fifo_out[114], \fifo_out.pt [113]);
tran (fifo_out[115], \fifo_out.pt [114]);
tran (fifo_out[116], \fifo_out.pt [115]);
tran (fifo_out[117], \fifo_out.pt [116]);
tran (fifo_out[118], \fifo_out.pt [117]);
tran (fifo_out[119], \fifo_out.pt [118]);
tran (fifo_out[120], \fifo_out.pt [119]);
tran (fifo_out[121], \fifo_out.pt [120]);
tran (fifo_out[122], \fifo_out.pt [121]);
tran (fifo_out[123], \fifo_out.pt [122]);
tran (fifo_out[124], \fifo_out.pt [123]);
tran (fifo_out[125], \fifo_out.pt [124]);
tran (fifo_out[126], \fifo_out.pt [125]);
tran (fifo_out[127], \fifo_out.pt [126]);
tran (fifo_out[128], \fifo_out.pt [127]);
tran (fifo_out[129], \fifo_out.op [0]);
tran (fifo_out[130], \fifo_out.op [1]);
tran (fifo_out[131], \fifo_out.op [2]);
Q_BUF U0 ( .A(n1648), .Z(mult_out[127]));
Q_BUF U1 ( .A(n1648), .Z(mult_out[126]));
Q_BUF U2 ( .A(n1648), .Z(mult_out[125]));
Q_BUF U3 ( .A(n1648), .Z(mult_out[124]));
Q_BUF U4 ( .A(n1648), .Z(mult_out[123]));
Q_BUF U5 ( .A(n1648), .Z(mult_out[122]));
Q_BUF U6 ( .A(n1648), .Z(mult_out[121]));
Q_BUF U7 ( .A(n1648), .Z(mult_out[120]));
Q_BUF U8 ( .A(n1648), .Z(mult_out[119]));
Q_BUF U9 ( .A(n1648), .Z(mult_out[118]));
Q_BUF U10 ( .A(n1648), .Z(mult_out[117]));
Q_BUF U11 ( .A(n1648), .Z(mult_out[116]));
Q_BUF U12 ( .A(n1648), .Z(mult_out[115]));
Q_BUF U13 ( .A(n1648), .Z(mult_out[114]));
Q_BUF U14 ( .A(n1648), .Z(mult_out[113]));
Q_BUF U15 ( .A(n1648), .Z(mult_out[112]));
Q_BUF U16 ( .A(n1648), .Z(mult_out[111]));
Q_BUF U17 ( .A(n1648), .Z(mult_out[110]));
Q_BUF U18 ( .A(n1648), .Z(mult_out[109]));
Q_BUF U19 ( .A(n1648), .Z(mult_out[108]));
Q_BUF U20 ( .A(n1648), .Z(mult_out[107]));
Q_BUF U21 ( .A(n1648), .Z(mult_out[106]));
Q_BUF U22 ( .A(n1648), .Z(mult_out[105]));
Q_BUF U23 ( .A(n1648), .Z(mult_out[104]));
Q_BUF U24 ( .A(n1648), .Z(mult_out[103]));
Q_BUF U25 ( .A(n1648), .Z(mult_out[102]));
Q_BUF U26 ( .A(n1648), .Z(mult_out[101]));
Q_BUF U27 ( .A(n1648), .Z(mult_out[100]));
Q_BUF U28 ( .A(n1648), .Z(mult_out[99]));
Q_BUF U29 ( .A(n1648), .Z(mult_out[98]));
Q_BUF U30 ( .A(n1648), .Z(mult_out[97]));
Q_BUF U31 ( .A(n1648), .Z(mult_out[96]));
Q_BUF U32 ( .A(n1648), .Z(mult_out[95]));
Q_BUF U33 ( .A(n1648), .Z(mult_out[94]));
Q_BUF U34 ( .A(n1648), .Z(mult_out[93]));
Q_BUF U35 ( .A(n1648), .Z(mult_out[92]));
Q_BUF U36 ( .A(n1648), .Z(mult_out[91]));
Q_BUF U37 ( .A(n1648), .Z(mult_out[90]));
Q_BUF U38 ( .A(n1648), .Z(mult_out[89]));
Q_BUF U39 ( .A(n1648), .Z(mult_out[88]));
Q_BUF U40 ( .A(n1648), .Z(mult_out[87]));
Q_BUF U41 ( .A(n1648), .Z(mult_out[86]));
Q_BUF U42 ( .A(n1648), .Z(mult_out[85]));
Q_BUF U43 ( .A(n1648), .Z(mult_out[84]));
Q_BUF U44 ( .A(n1648), .Z(mult_out[83]));
Q_BUF U45 ( .A(n1648), .Z(mult_out[82]));
Q_BUF U46 ( .A(n1648), .Z(mult_out[81]));
Q_BUF U47 ( .A(n1648), .Z(mult_out[80]));
Q_BUF U48 ( .A(n1648), .Z(mult_out[79]));
Q_BUF U49 ( .A(n1648), .Z(mult_out[78]));
Q_BUF U50 ( .A(n1648), .Z(mult_out[77]));
Q_BUF U51 ( .A(n1648), .Z(mult_out[76]));
Q_BUF U52 ( .A(n1648), .Z(mult_out[75]));
Q_BUF U53 ( .A(n1648), .Z(mult_out[74]));
Q_BUF U54 ( .A(n1648), .Z(mult_out[73]));
Q_BUF U55 ( .A(n1648), .Z(mult_out[72]));
Q_BUF U56 ( .A(n1648), .Z(mult_out[71]));
Q_BUF U57 ( .A(n1648), .Z(mult_out[70]));
Q_BUF U58 ( .A(n1648), .Z(mult_out[69]));
Q_BUF U59 ( .A(n1648), .Z(mult_out[68]));
Q_BUF U60 ( .A(n1648), .Z(mult_out[67]));
Q_BUF U61 ( .A(n1648), .Z(mult_out[66]));
Q_BUF U62 ( .A(n1648), .Z(mult_out[65]));
Q_BUF U63 ( .A(n1648), .Z(mult_out[64]));
Q_BUF U64 ( .A(n1648), .Z(mult_out[63]));
Q_BUF U65 ( .A(n1648), .Z(mult_out[62]));
Q_BUF U66 ( .A(n1648), .Z(mult_out[61]));
Q_BUF U67 ( .A(n1648), .Z(mult_out[60]));
Q_BUF U68 ( .A(n1648), .Z(mult_out[59]));
Q_BUF U69 ( .A(n1648), .Z(mult_out[58]));
Q_BUF U70 ( .A(n1648), .Z(mult_out[57]));
Q_BUF U71 ( .A(n1648), .Z(mult_out[56]));
Q_BUF U72 ( .A(n1648), .Z(mult_out[55]));
Q_BUF U73 ( .A(n1648), .Z(mult_out[54]));
Q_BUF U74 ( .A(n1648), .Z(mult_out[53]));
Q_BUF U75 ( .A(n1648), .Z(mult_out[52]));
Q_BUF U76 ( .A(n1648), .Z(mult_out[51]));
Q_BUF U77 ( .A(n1648), .Z(mult_out[50]));
Q_BUF U78 ( .A(n1648), .Z(mult_out[49]));
Q_BUF U79 ( .A(n1648), .Z(mult_out[48]));
Q_BUF U80 ( .A(n1648), .Z(mult_out[47]));
Q_BUF U81 ( .A(n1648), .Z(mult_out[46]));
Q_BUF U82 ( .A(n1648), .Z(mult_out[45]));
Q_BUF U83 ( .A(n1648), .Z(mult_out[44]));
Q_BUF U84 ( .A(n1648), .Z(mult_out[43]));
Q_BUF U85 ( .A(n1648), .Z(mult_out[42]));
Q_BUF U86 ( .A(n1648), .Z(mult_out[41]));
Q_BUF U87 ( .A(n1648), .Z(mult_out[40]));
Q_BUF U88 ( .A(n1648), .Z(mult_out[39]));
Q_BUF U89 ( .A(n1648), .Z(mult_out[38]));
Q_BUF U90 ( .A(n1648), .Z(mult_out[37]));
Q_BUF U91 ( .A(n1648), .Z(mult_out[36]));
Q_BUF U92 ( .A(n1648), .Z(mult_out[35]));
Q_BUF U93 ( .A(n1648), .Z(mult_out[34]));
Q_BUF U94 ( .A(n1648), .Z(mult_out[33]));
Q_BUF U95 ( .A(n1648), .Z(mult_out[32]));
Q_BUF U96 ( .A(n1648), .Z(mult_out[31]));
Q_BUF U97 ( .A(n1648), .Z(mult_out[30]));
Q_BUF U98 ( .A(n1648), .Z(mult_out[29]));
Q_BUF U99 ( .A(n1648), .Z(mult_out[28]));
Q_BUF U100 ( .A(n1648), .Z(mult_out[27]));
Q_BUF U101 ( .A(n1648), .Z(mult_out[26]));
Q_BUF U102 ( .A(n1648), .Z(mult_out[25]));
Q_BUF U103 ( .A(n1648), .Z(mult_out[24]));
Q_BUF U104 ( .A(n1648), .Z(mult_out[23]));
Q_BUF U105 ( .A(n1648), .Z(mult_out[22]));
Q_BUF U106 ( .A(n1648), .Z(mult_out[21]));
Q_BUF U107 ( .A(n1648), .Z(mult_out[20]));
Q_BUF U108 ( .A(n1648), .Z(mult_out[19]));
Q_BUF U109 ( .A(n1648), .Z(mult_out[18]));
Q_BUF U110 ( .A(n1648), .Z(mult_out[17]));
Q_BUF U111 ( .A(n1648), .Z(mult_out[16]));
Q_BUF U112 ( .A(n1648), .Z(mult_out[15]));
Q_BUF U113 ( .A(n1648), .Z(mult_out[14]));
Q_BUF U114 ( .A(n1648), .Z(mult_out[13]));
Q_BUF U115 ( .A(n1648), .Z(mult_out[12]));
Q_BUF U116 ( .A(n1648), .Z(mult_out[11]));
Q_BUF U117 ( .A(n1648), .Z(mult_out[10]));
Q_BUF U118 ( .A(n1648), .Z(mult_out[9]));
Q_BUF U119 ( .A(n1648), .Z(mult_out[8]));
Q_BUF U120 ( .A(n1648), .Z(mult_out[7]));
Q_BUF U121 ( .A(n1648), .Z(mult_out[6]));
Q_BUF U122 ( .A(n1648), .Z(mult_out[5]));
Q_BUF U123 ( .A(n1648), .Z(mult_out[4]));
Q_BUF U124 ( .A(n1648), .Z(mult_out[3]));
Q_BUF U125 ( .A(n1648), .Z(mult_out[2]));
Q_BUF U126 ( .A(n1648), .Z(mult_out[1]));
Q_BUF U127 ( .A(n1648), .Z(mult_out[0]));
Q_BUF U128 ( .A(n1648), .Z(_zy_simnet_cio_8));
Q_BUF U129 ( .A(n1648), .Z(_zy_simnet_cio_9));
Q_BUF U130 ( .A(n1), .Z(_zy_simnet_cio_10));
Q_BUF U131 ( .A(n1), .Z(_zy_simnet_cio_14));
Q_BUF U132 ( .A(n1648), .Z(_zy_simnet_cio_24));
Q_BUF U133 ( .A(n1648), .Z(set_gcm_tag_fail_int));
Q_BUF U134 ( .A(fifo_in_vld), .Z(ciph_in_vld));
Q_ASSIGN U135 ( .B(ciph_out_vld), .A(fifo_out_ack));
Q_BUF U136 ( .A(h_value[127]), .Z(operand_Y[127]));
Q_BUF U137 ( .A(h_value[126]), .Z(operand_Y[126]));
Q_BUF U138 ( .A(h_value[125]), .Z(operand_Y[125]));
Q_BUF U139 ( .A(h_value[124]), .Z(operand_Y[124]));
Q_BUF U140 ( .A(h_value[123]), .Z(operand_Y[123]));
Q_BUF U141 ( .A(h_value[122]), .Z(operand_Y[122]));
Q_BUF U142 ( .A(h_value[121]), .Z(operand_Y[121]));
Q_BUF U143 ( .A(h_value[120]), .Z(operand_Y[120]));
Q_BUF U144 ( .A(h_value[119]), .Z(operand_Y[119]));
Q_BUF U145 ( .A(h_value[118]), .Z(operand_Y[118]));
Q_BUF U146 ( .A(h_value[117]), .Z(operand_Y[117]));
Q_BUF U147 ( .A(h_value[116]), .Z(operand_Y[116]));
Q_BUF U148 ( .A(h_value[115]), .Z(operand_Y[115]));
Q_BUF U149 ( .A(h_value[114]), .Z(operand_Y[114]));
Q_BUF U150 ( .A(h_value[113]), .Z(operand_Y[113]));
Q_BUF U151 ( .A(h_value[112]), .Z(operand_Y[112]));
Q_BUF U152 ( .A(h_value[111]), .Z(operand_Y[111]));
Q_BUF U153 ( .A(h_value[110]), .Z(operand_Y[110]));
Q_BUF U154 ( .A(h_value[109]), .Z(operand_Y[109]));
Q_BUF U155 ( .A(h_value[108]), .Z(operand_Y[108]));
Q_BUF U156 ( .A(h_value[107]), .Z(operand_Y[107]));
Q_BUF U157 ( .A(h_value[106]), .Z(operand_Y[106]));
Q_BUF U158 ( .A(h_value[105]), .Z(operand_Y[105]));
Q_BUF U159 ( .A(h_value[104]), .Z(operand_Y[104]));
Q_BUF U160 ( .A(h_value[103]), .Z(operand_Y[103]));
Q_BUF U161 ( .A(h_value[102]), .Z(operand_Y[102]));
Q_BUF U162 ( .A(h_value[101]), .Z(operand_Y[101]));
Q_BUF U163 ( .A(h_value[100]), .Z(operand_Y[100]));
Q_BUF U164 ( .A(h_value[99]), .Z(operand_Y[99]));
Q_BUF U165 ( .A(h_value[98]), .Z(operand_Y[98]));
Q_BUF U166 ( .A(h_value[97]), .Z(operand_Y[97]));
Q_BUF U167 ( .A(h_value[96]), .Z(operand_Y[96]));
Q_BUF U168 ( .A(h_value[95]), .Z(operand_Y[95]));
Q_BUF U169 ( .A(h_value[94]), .Z(operand_Y[94]));
Q_BUF U170 ( .A(h_value[93]), .Z(operand_Y[93]));
Q_BUF U171 ( .A(h_value[92]), .Z(operand_Y[92]));
Q_BUF U172 ( .A(h_value[91]), .Z(operand_Y[91]));
Q_BUF U173 ( .A(h_value[90]), .Z(operand_Y[90]));
Q_BUF U174 ( .A(h_value[89]), .Z(operand_Y[89]));
Q_BUF U175 ( .A(h_value[88]), .Z(operand_Y[88]));
Q_BUF U176 ( .A(h_value[87]), .Z(operand_Y[87]));
Q_BUF U177 ( .A(h_value[86]), .Z(operand_Y[86]));
Q_BUF U178 ( .A(h_value[85]), .Z(operand_Y[85]));
Q_BUF U179 ( .A(h_value[84]), .Z(operand_Y[84]));
Q_BUF U180 ( .A(h_value[83]), .Z(operand_Y[83]));
Q_BUF U181 ( .A(h_value[82]), .Z(operand_Y[82]));
Q_BUF U182 ( .A(h_value[81]), .Z(operand_Y[81]));
Q_BUF U183 ( .A(h_value[80]), .Z(operand_Y[80]));
Q_BUF U184 ( .A(h_value[79]), .Z(operand_Y[79]));
Q_BUF U185 ( .A(h_value[78]), .Z(operand_Y[78]));
Q_BUF U186 ( .A(h_value[77]), .Z(operand_Y[77]));
Q_BUF U187 ( .A(h_value[76]), .Z(operand_Y[76]));
Q_BUF U188 ( .A(h_value[75]), .Z(operand_Y[75]));
Q_BUF U189 ( .A(h_value[74]), .Z(operand_Y[74]));
Q_BUF U190 ( .A(h_value[73]), .Z(operand_Y[73]));
Q_BUF U191 ( .A(h_value[72]), .Z(operand_Y[72]));
Q_BUF U192 ( .A(h_value[71]), .Z(operand_Y[71]));
Q_BUF U193 ( .A(h_value[70]), .Z(operand_Y[70]));
Q_BUF U194 ( .A(h_value[69]), .Z(operand_Y[69]));
Q_BUF U195 ( .A(h_value[68]), .Z(operand_Y[68]));
Q_BUF U196 ( .A(h_value[67]), .Z(operand_Y[67]));
Q_BUF U197 ( .A(h_value[66]), .Z(operand_Y[66]));
Q_BUF U198 ( .A(h_value[65]), .Z(operand_Y[65]));
Q_BUF U199 ( .A(h_value[64]), .Z(operand_Y[64]));
Q_BUF U200 ( .A(h_value[63]), .Z(operand_Y[63]));
Q_BUF U201 ( .A(h_value[62]), .Z(operand_Y[62]));
Q_BUF U202 ( .A(h_value[61]), .Z(operand_Y[61]));
Q_BUF U203 ( .A(h_value[60]), .Z(operand_Y[60]));
Q_BUF U204 ( .A(h_value[59]), .Z(operand_Y[59]));
Q_BUF U205 ( .A(h_value[58]), .Z(operand_Y[58]));
Q_BUF U206 ( .A(h_value[57]), .Z(operand_Y[57]));
Q_BUF U207 ( .A(h_value[56]), .Z(operand_Y[56]));
Q_BUF U208 ( .A(h_value[55]), .Z(operand_Y[55]));
Q_BUF U209 ( .A(h_value[54]), .Z(operand_Y[54]));
Q_BUF U210 ( .A(h_value[53]), .Z(operand_Y[53]));
Q_BUF U211 ( .A(h_value[52]), .Z(operand_Y[52]));
Q_BUF U212 ( .A(h_value[51]), .Z(operand_Y[51]));
Q_BUF U213 ( .A(h_value[50]), .Z(operand_Y[50]));
Q_BUF U214 ( .A(h_value[49]), .Z(operand_Y[49]));
Q_BUF U215 ( .A(h_value[48]), .Z(operand_Y[48]));
Q_BUF U216 ( .A(h_value[47]), .Z(operand_Y[47]));
Q_BUF U217 ( .A(h_value[46]), .Z(operand_Y[46]));
Q_BUF U218 ( .A(h_value[45]), .Z(operand_Y[45]));
Q_BUF U219 ( .A(h_value[44]), .Z(operand_Y[44]));
Q_BUF U220 ( .A(h_value[43]), .Z(operand_Y[43]));
Q_BUF U221 ( .A(h_value[42]), .Z(operand_Y[42]));
Q_BUF U222 ( .A(h_value[41]), .Z(operand_Y[41]));
Q_BUF U223 ( .A(h_value[40]), .Z(operand_Y[40]));
Q_BUF U224 ( .A(h_value[39]), .Z(operand_Y[39]));
Q_BUF U225 ( .A(h_value[38]), .Z(operand_Y[38]));
Q_BUF U226 ( .A(h_value[37]), .Z(operand_Y[37]));
Q_BUF U227 ( .A(h_value[36]), .Z(operand_Y[36]));
Q_BUF U228 ( .A(h_value[35]), .Z(operand_Y[35]));
Q_BUF U229 ( .A(h_value[34]), .Z(operand_Y[34]));
Q_BUF U230 ( .A(h_value[33]), .Z(operand_Y[33]));
Q_BUF U231 ( .A(h_value[32]), .Z(operand_Y[32]));
Q_BUF U232 ( .A(h_value[31]), .Z(operand_Y[31]));
Q_BUF U233 ( .A(h_value[30]), .Z(operand_Y[30]));
Q_BUF U234 ( .A(h_value[29]), .Z(operand_Y[29]));
Q_BUF U235 ( .A(h_value[28]), .Z(operand_Y[28]));
Q_BUF U236 ( .A(h_value[27]), .Z(operand_Y[27]));
Q_BUF U237 ( .A(h_value[26]), .Z(operand_Y[26]));
Q_BUF U238 ( .A(h_value[25]), .Z(operand_Y[25]));
Q_BUF U239 ( .A(h_value[24]), .Z(operand_Y[24]));
Q_BUF U240 ( .A(h_value[23]), .Z(operand_Y[23]));
Q_BUF U241 ( .A(h_value[22]), .Z(operand_Y[22]));
Q_BUF U242 ( .A(h_value[21]), .Z(operand_Y[21]));
Q_BUF U243 ( .A(h_value[20]), .Z(operand_Y[20]));
Q_BUF U244 ( .A(h_value[19]), .Z(operand_Y[19]));
Q_BUF U245 ( .A(h_value[18]), .Z(operand_Y[18]));
Q_BUF U246 ( .A(h_value[17]), .Z(operand_Y[17]));
Q_BUF U247 ( .A(h_value[16]), .Z(operand_Y[16]));
Q_BUF U248 ( .A(h_value[15]), .Z(operand_Y[15]));
Q_BUF U249 ( .A(h_value[14]), .Z(operand_Y[14]));
Q_BUF U250 ( .A(h_value[13]), .Z(operand_Y[13]));
Q_BUF U251 ( .A(h_value[12]), .Z(operand_Y[12]));
Q_BUF U252 ( .A(h_value[11]), .Z(operand_Y[11]));
Q_BUF U253 ( .A(h_value[10]), .Z(operand_Y[10]));
Q_BUF U254 ( .A(h_value[9]), .Z(operand_Y[9]));
Q_BUF U255 ( .A(h_value[8]), .Z(operand_Y[8]));
Q_BUF U256 ( .A(h_value[7]), .Z(operand_Y[7]));
Q_BUF U257 ( .A(h_value[6]), .Z(operand_Y[6]));
Q_BUF U258 ( .A(h_value[5]), .Z(operand_Y[5]));
Q_BUF U259 ( .A(h_value[4]), .Z(operand_Y[4]));
Q_BUF U260 ( .A(h_value[3]), .Z(operand_Y[3]));
Q_BUF U261 ( .A(h_value[2]), .Z(operand_Y[2]));
Q_BUF U262 ( .A(h_value[1]), .Z(operand_Y[1]));
Q_BUF U263 ( .A(h_value[0]), .Z(operand_Y[0]));
Q_BUF U264 ( .A(n1648), .Z(gcm_status_data_in[0]));
Q_OR02 U265 ( .A0(n1222), .A1(n627), .Z(n2));
Q_OR02 U266 ( .A0(n560), .A1(n549), .Z(n3));
Q_INV U267 ( .A(fifo_out[129]), .Z(n24));
Q_INV U268 ( .A(fifo_out_vld), .Z(n9));
Q_OR02 U269 ( .A0(fifo_out[131]), .A1(n9), .Z(n20));
Q_OR02 U270 ( .A0(fifo_out[130]), .A1(n20), .Z(n14));
Q_INV U271 ( .A(ciph_out_vld), .Z(n21));
Q_OR02 U272 ( .A0(n21), .A1(n14), .Z(n18));
Q_INV U273 ( .A(fifo_out[130]), .Z(n10));
Q_OR02 U274 ( .A0(n10), .A1(n20), .Z(n15));
Q_OR02 U275 ( .A0(n21), .A1(n15), .Z(n23));
Q_ND02 U276 ( .A0(n11), .A1(n12), .Z(gcm_kdf_valid));
Q_OR02 U277 ( .A0(n24), .A1(n18), .Z(n11));
Q_OR02 U278 ( .A0(fifo_out[129]), .A1(n23), .Z(n12));
Q_INV U279 ( .A(n12), .Z(n4));
Q_ND02 U280 ( .A0(fifo_out[131]), .A1(fifo_out_vld), .Z(n13));
Q_OR02 U281 ( .A0(fifo_out[130]), .A1(n13), .Z(n17));
Q_NR02 U282 ( .A0(n21), .A1(n17), .Z(gcm_status_data_in_valid));
Q_MX02 U283 ( .S(fifo_out[129]), .A0(n15), .A1(n14), .Z(n16));
Q_INV U284 ( .A(n17), .Z(n5));
Q_INV U285 ( .A(n23), .Z(n6));
Q_OR02 U286 ( .A0(fifo_out[129]), .A1(n18), .Z(n19));
Q_OR03 U287 ( .A0(n21), .A1(n20), .A2(fifo_out[129]), .Z(n22));
Q_AN02 U288 ( .A0(n25), .A1(n22), .Z(n7));
Q_OR02 U289 ( .A0(n24), .A1(n23), .Z(n25));
Q_INV U290 ( .A(n25), .Z(n8));
Q_AN02 U291 ( .A0(gcm_kdf_valid), .A1(fifo_out[0]), .Z(gcm_kdf_eof));
Q_MX02 U292 ( .S(n11), .A0(fifo_out[128]), .A1(n26), .Z(gcm_kdf_data[127]));
Q_AN02 U293 ( .A0(n4), .A1(n411), .Z(n26));
Q_MX02 U294 ( .S(n11), .A0(fifo_out[127]), .A1(n27), .Z(gcm_kdf_data[126]));
Q_AN02 U295 ( .A0(n4), .A1(n412), .Z(n27));
Q_MX02 U296 ( .S(n11), .A0(fifo_out[126]), .A1(n28), .Z(gcm_kdf_data[125]));
Q_AN02 U297 ( .A0(n4), .A1(n413), .Z(n28));
Q_MX02 U298 ( .S(n11), .A0(fifo_out[125]), .A1(n29), .Z(gcm_kdf_data[124]));
Q_AN02 U299 ( .A0(n4), .A1(n414), .Z(n29));
Q_MX02 U300 ( .S(n11), .A0(fifo_out[124]), .A1(n30), .Z(gcm_kdf_data[123]));
Q_AN02 U301 ( .A0(n4), .A1(n415), .Z(n30));
Q_MX02 U302 ( .S(n11), .A0(fifo_out[123]), .A1(n31), .Z(gcm_kdf_data[122]));
Q_AN02 U303 ( .A0(n4), .A1(n416), .Z(n31));
Q_MX02 U304 ( .S(n11), .A0(fifo_out[122]), .A1(n32), .Z(gcm_kdf_data[121]));
Q_AN02 U305 ( .A0(n4), .A1(n417), .Z(n32));
Q_MX02 U306 ( .S(n11), .A0(fifo_out[121]), .A1(n33), .Z(gcm_kdf_data[120]));
Q_AN02 U307 ( .A0(n4), .A1(n418), .Z(n33));
Q_MX02 U308 ( .S(n11), .A0(fifo_out[120]), .A1(n34), .Z(gcm_kdf_data[119]));
Q_AN02 U309 ( .A0(n4), .A1(n419), .Z(n34));
Q_MX02 U310 ( .S(n11), .A0(fifo_out[119]), .A1(n35), .Z(gcm_kdf_data[118]));
Q_AN02 U311 ( .A0(n4), .A1(n420), .Z(n35));
Q_MX02 U312 ( .S(n11), .A0(fifo_out[118]), .A1(n36), .Z(gcm_kdf_data[117]));
Q_AN02 U313 ( .A0(n4), .A1(n421), .Z(n36));
Q_MX02 U314 ( .S(n11), .A0(fifo_out[117]), .A1(n37), .Z(gcm_kdf_data[116]));
Q_AN02 U315 ( .A0(n4), .A1(n422), .Z(n37));
Q_MX02 U316 ( .S(n11), .A0(fifo_out[116]), .A1(n38), .Z(gcm_kdf_data[115]));
Q_AN02 U317 ( .A0(n4), .A1(n423), .Z(n38));
Q_MX02 U318 ( .S(n11), .A0(fifo_out[115]), .A1(n39), .Z(gcm_kdf_data[114]));
Q_AN02 U319 ( .A0(n4), .A1(n424), .Z(n39));
Q_MX02 U320 ( .S(n11), .A0(fifo_out[114]), .A1(n40), .Z(gcm_kdf_data[113]));
Q_AN02 U321 ( .A0(n4), .A1(n425), .Z(n40));
Q_MX02 U322 ( .S(n11), .A0(fifo_out[113]), .A1(n41), .Z(gcm_kdf_data[112]));
Q_AN02 U323 ( .A0(n4), .A1(n426), .Z(n41));
Q_MX02 U324 ( .S(n11), .A0(fifo_out[112]), .A1(n42), .Z(gcm_kdf_data[111]));
Q_AN02 U325 ( .A0(n4), .A1(n427), .Z(n42));
Q_MX02 U326 ( .S(n11), .A0(fifo_out[111]), .A1(n43), .Z(gcm_kdf_data[110]));
Q_AN02 U327 ( .A0(n4), .A1(n428), .Z(n43));
Q_MX02 U328 ( .S(n11), .A0(fifo_out[110]), .A1(n44), .Z(gcm_kdf_data[109]));
Q_AN02 U329 ( .A0(n4), .A1(n429), .Z(n44));
Q_MX02 U330 ( .S(n11), .A0(fifo_out[109]), .A1(n45), .Z(gcm_kdf_data[108]));
Q_AN02 U331 ( .A0(n4), .A1(n430), .Z(n45));
Q_MX02 U332 ( .S(n11), .A0(fifo_out[108]), .A1(n46), .Z(gcm_kdf_data[107]));
Q_AN02 U333 ( .A0(n4), .A1(n431), .Z(n46));
Q_MX02 U334 ( .S(n11), .A0(fifo_out[107]), .A1(n47), .Z(gcm_kdf_data[106]));
Q_AN02 U335 ( .A0(n4), .A1(n432), .Z(n47));
Q_MX02 U336 ( .S(n11), .A0(fifo_out[106]), .A1(n48), .Z(gcm_kdf_data[105]));
Q_AN02 U337 ( .A0(n4), .A1(n433), .Z(n48));
Q_MX02 U338 ( .S(n11), .A0(fifo_out[105]), .A1(n49), .Z(gcm_kdf_data[104]));
Q_AN02 U339 ( .A0(n4), .A1(n434), .Z(n49));
Q_MX02 U340 ( .S(n11), .A0(fifo_out[104]), .A1(n50), .Z(gcm_kdf_data[103]));
Q_AN02 U341 ( .A0(n4), .A1(n435), .Z(n50));
Q_MX02 U342 ( .S(n11), .A0(fifo_out[103]), .A1(n51), .Z(gcm_kdf_data[102]));
Q_AN02 U343 ( .A0(n4), .A1(n436), .Z(n51));
Q_MX02 U344 ( .S(n11), .A0(fifo_out[102]), .A1(n52), .Z(gcm_kdf_data[101]));
Q_AN02 U345 ( .A0(n4), .A1(n437), .Z(n52));
Q_MX02 U346 ( .S(n11), .A0(fifo_out[101]), .A1(n53), .Z(gcm_kdf_data[100]));
Q_AN02 U347 ( .A0(n4), .A1(n438), .Z(n53));
Q_MX02 U348 ( .S(n11), .A0(fifo_out[100]), .A1(n54), .Z(gcm_kdf_data[99]));
Q_AN02 U349 ( .A0(n4), .A1(n439), .Z(n54));
Q_MX02 U350 ( .S(n11), .A0(fifo_out[99]), .A1(n55), .Z(gcm_kdf_data[98]));
Q_AN02 U351 ( .A0(n4), .A1(n440), .Z(n55));
Q_MX02 U352 ( .S(n11), .A0(fifo_out[98]), .A1(n56), .Z(gcm_kdf_data[97]));
Q_AN02 U353 ( .A0(n4), .A1(n441), .Z(n56));
Q_MX02 U354 ( .S(n11), .A0(fifo_out[97]), .A1(n57), .Z(gcm_kdf_data[96]));
Q_AN02 U355 ( .A0(n4), .A1(n442), .Z(n57));
Q_MX02 U356 ( .S(n11), .A0(fifo_out[96]), .A1(n58), .Z(gcm_kdf_data[95]));
Q_AN02 U357 ( .A0(n4), .A1(n443), .Z(n58));
Q_MX02 U358 ( .S(n11), .A0(fifo_out[95]), .A1(n59), .Z(gcm_kdf_data[94]));
Q_AN02 U359 ( .A0(n4), .A1(n444), .Z(n59));
Q_MX02 U360 ( .S(n11), .A0(fifo_out[94]), .A1(n60), .Z(gcm_kdf_data[93]));
Q_AN02 U361 ( .A0(n4), .A1(n445), .Z(n60));
Q_MX02 U362 ( .S(n11), .A0(fifo_out[93]), .A1(n61), .Z(gcm_kdf_data[92]));
Q_AN02 U363 ( .A0(n4), .A1(n446), .Z(n61));
Q_MX02 U364 ( .S(n11), .A0(fifo_out[92]), .A1(n62), .Z(gcm_kdf_data[91]));
Q_AN02 U365 ( .A0(n4), .A1(n447), .Z(n62));
Q_MX02 U366 ( .S(n11), .A0(fifo_out[91]), .A1(n63), .Z(gcm_kdf_data[90]));
Q_AN02 U367 ( .A0(n4), .A1(n448), .Z(n63));
Q_MX02 U368 ( .S(n11), .A0(fifo_out[90]), .A1(n64), .Z(gcm_kdf_data[89]));
Q_AN02 U369 ( .A0(n4), .A1(n449), .Z(n64));
Q_MX02 U370 ( .S(n11), .A0(fifo_out[89]), .A1(n65), .Z(gcm_kdf_data[88]));
Q_AN02 U371 ( .A0(n4), .A1(n450), .Z(n65));
Q_MX02 U372 ( .S(n11), .A0(fifo_out[88]), .A1(n66), .Z(gcm_kdf_data[87]));
Q_AN02 U373 ( .A0(n4), .A1(n451), .Z(n66));
Q_MX02 U374 ( .S(n11), .A0(fifo_out[87]), .A1(n67), .Z(gcm_kdf_data[86]));
Q_AN02 U375 ( .A0(n4), .A1(n452), .Z(n67));
Q_MX02 U376 ( .S(n11), .A0(fifo_out[86]), .A1(n68), .Z(gcm_kdf_data[85]));
Q_AN02 U377 ( .A0(n4), .A1(n453), .Z(n68));
Q_MX02 U378 ( .S(n11), .A0(fifo_out[85]), .A1(n69), .Z(gcm_kdf_data[84]));
Q_AN02 U379 ( .A0(n4), .A1(n454), .Z(n69));
Q_MX02 U380 ( .S(n11), .A0(fifo_out[84]), .A1(n70), .Z(gcm_kdf_data[83]));
Q_AN02 U381 ( .A0(n4), .A1(n455), .Z(n70));
Q_MX02 U382 ( .S(n11), .A0(fifo_out[83]), .A1(n71), .Z(gcm_kdf_data[82]));
Q_AN02 U383 ( .A0(n4), .A1(n456), .Z(n71));
Q_MX02 U384 ( .S(n11), .A0(fifo_out[82]), .A1(n72), .Z(gcm_kdf_data[81]));
Q_AN02 U385 ( .A0(n4), .A1(n457), .Z(n72));
Q_MX02 U386 ( .S(n11), .A0(fifo_out[81]), .A1(n73), .Z(gcm_kdf_data[80]));
Q_AN02 U387 ( .A0(n4), .A1(n458), .Z(n73));
Q_MX02 U388 ( .S(n11), .A0(fifo_out[80]), .A1(n74), .Z(gcm_kdf_data[79]));
Q_AN02 U389 ( .A0(n4), .A1(n459), .Z(n74));
Q_MX02 U390 ( .S(n11), .A0(fifo_out[79]), .A1(n75), .Z(gcm_kdf_data[78]));
Q_AN02 U391 ( .A0(n4), .A1(n460), .Z(n75));
Q_MX02 U392 ( .S(n11), .A0(fifo_out[78]), .A1(n76), .Z(gcm_kdf_data[77]));
Q_AN02 U393 ( .A0(n4), .A1(n461), .Z(n76));
Q_MX02 U394 ( .S(n11), .A0(fifo_out[77]), .A1(n77), .Z(gcm_kdf_data[76]));
Q_AN02 U395 ( .A0(n4), .A1(n462), .Z(n77));
Q_MX02 U396 ( .S(n11), .A0(fifo_out[76]), .A1(n78), .Z(gcm_kdf_data[75]));
Q_AN02 U397 ( .A0(n4), .A1(n463), .Z(n78));
Q_MX02 U398 ( .S(n11), .A0(fifo_out[75]), .A1(n79), .Z(gcm_kdf_data[74]));
Q_AN02 U399 ( .A0(n4), .A1(n464), .Z(n79));
Q_MX02 U400 ( .S(n11), .A0(fifo_out[74]), .A1(n80), .Z(gcm_kdf_data[73]));
Q_AN02 U401 ( .A0(n4), .A1(n465), .Z(n80));
Q_MX02 U402 ( .S(n11), .A0(fifo_out[73]), .A1(n81), .Z(gcm_kdf_data[72]));
Q_AN02 U403 ( .A0(n4), .A1(n466), .Z(n81));
Q_MX02 U404 ( .S(n11), .A0(fifo_out[72]), .A1(n82), .Z(gcm_kdf_data[71]));
Q_AN02 U405 ( .A0(n4), .A1(n467), .Z(n82));
Q_MX02 U406 ( .S(n11), .A0(fifo_out[71]), .A1(n83), .Z(gcm_kdf_data[70]));
Q_AN02 U407 ( .A0(n4), .A1(n468), .Z(n83));
Q_MX02 U408 ( .S(n11), .A0(fifo_out[70]), .A1(n84), .Z(gcm_kdf_data[69]));
Q_AN02 U409 ( .A0(n4), .A1(n469), .Z(n84));
Q_MX02 U410 ( .S(n11), .A0(fifo_out[69]), .A1(n85), .Z(gcm_kdf_data[68]));
Q_AN02 U411 ( .A0(n4), .A1(n470), .Z(n85));
Q_MX02 U412 ( .S(n11), .A0(fifo_out[68]), .A1(n86), .Z(gcm_kdf_data[67]));
Q_AN02 U413 ( .A0(n4), .A1(n471), .Z(n86));
Q_MX02 U414 ( .S(n11), .A0(fifo_out[67]), .A1(n87), .Z(gcm_kdf_data[66]));
Q_AN02 U415 ( .A0(n4), .A1(n472), .Z(n87));
Q_MX02 U416 ( .S(n11), .A0(fifo_out[66]), .A1(n88), .Z(gcm_kdf_data[65]));
Q_AN02 U417 ( .A0(n4), .A1(n473), .Z(n88));
Q_MX02 U418 ( .S(n11), .A0(fifo_out[65]), .A1(n89), .Z(gcm_kdf_data[64]));
Q_AN02 U419 ( .A0(n4), .A1(n474), .Z(n89));
Q_MX02 U420 ( .S(n11), .A0(fifo_out[64]), .A1(n90), .Z(gcm_kdf_data[63]));
Q_AN02 U421 ( .A0(n4), .A1(n475), .Z(n90));
Q_MX02 U422 ( .S(n11), .A0(fifo_out[63]), .A1(n91), .Z(gcm_kdf_data[62]));
Q_AN02 U423 ( .A0(n4), .A1(n476), .Z(n91));
Q_MX02 U424 ( .S(n11), .A0(fifo_out[62]), .A1(n92), .Z(gcm_kdf_data[61]));
Q_AN02 U425 ( .A0(n4), .A1(n477), .Z(n92));
Q_MX02 U426 ( .S(n11), .A0(fifo_out[61]), .A1(n93), .Z(gcm_kdf_data[60]));
Q_AN02 U427 ( .A0(n4), .A1(n478), .Z(n93));
Q_MX02 U428 ( .S(n11), .A0(fifo_out[60]), .A1(n94), .Z(gcm_kdf_data[59]));
Q_AN02 U429 ( .A0(n4), .A1(n479), .Z(n94));
Q_MX02 U430 ( .S(n11), .A0(fifo_out[59]), .A1(n95), .Z(gcm_kdf_data[58]));
Q_AN02 U431 ( .A0(n4), .A1(n480), .Z(n95));
Q_MX02 U432 ( .S(n11), .A0(fifo_out[58]), .A1(n96), .Z(gcm_kdf_data[57]));
Q_AN02 U433 ( .A0(n4), .A1(n481), .Z(n96));
Q_MX02 U434 ( .S(n11), .A0(fifo_out[57]), .A1(n97), .Z(gcm_kdf_data[56]));
Q_AN02 U435 ( .A0(n4), .A1(n482), .Z(n97));
Q_MX02 U436 ( .S(n11), .A0(fifo_out[56]), .A1(n98), .Z(gcm_kdf_data[55]));
Q_AN02 U437 ( .A0(n4), .A1(n483), .Z(n98));
Q_MX02 U438 ( .S(n11), .A0(fifo_out[55]), .A1(n99), .Z(gcm_kdf_data[54]));
Q_AN02 U439 ( .A0(n4), .A1(n484), .Z(n99));
Q_MX02 U440 ( .S(n11), .A0(fifo_out[54]), .A1(n100), .Z(gcm_kdf_data[53]));
Q_AN02 U441 ( .A0(n4), .A1(n485), .Z(n100));
Q_MX02 U442 ( .S(n11), .A0(fifo_out[53]), .A1(n101), .Z(gcm_kdf_data[52]));
Q_AN02 U443 ( .A0(n4), .A1(n486), .Z(n101));
Q_MX02 U444 ( .S(n11), .A0(fifo_out[52]), .A1(n102), .Z(gcm_kdf_data[51]));
Q_AN02 U445 ( .A0(n4), .A1(n487), .Z(n102));
Q_MX02 U446 ( .S(n11), .A0(fifo_out[51]), .A1(n103), .Z(gcm_kdf_data[50]));
Q_AN02 U447 ( .A0(n4), .A1(n488), .Z(n103));
Q_MX02 U448 ( .S(n11), .A0(fifo_out[50]), .A1(n104), .Z(gcm_kdf_data[49]));
Q_AN02 U449 ( .A0(n4), .A1(n489), .Z(n104));
Q_MX02 U450 ( .S(n11), .A0(fifo_out[49]), .A1(n105), .Z(gcm_kdf_data[48]));
Q_AN02 U451 ( .A0(n4), .A1(n490), .Z(n105));
Q_MX02 U452 ( .S(n11), .A0(fifo_out[48]), .A1(n106), .Z(gcm_kdf_data[47]));
Q_AN02 U453 ( .A0(n4), .A1(n491), .Z(n106));
Q_MX02 U454 ( .S(n11), .A0(fifo_out[47]), .A1(n107), .Z(gcm_kdf_data[46]));
Q_AN02 U455 ( .A0(n4), .A1(n492), .Z(n107));
Q_MX02 U456 ( .S(n11), .A0(fifo_out[46]), .A1(n108), .Z(gcm_kdf_data[45]));
Q_AN02 U457 ( .A0(n4), .A1(n493), .Z(n108));
Q_MX02 U458 ( .S(n11), .A0(fifo_out[45]), .A1(n109), .Z(gcm_kdf_data[44]));
Q_AN02 U459 ( .A0(n4), .A1(n494), .Z(n109));
Q_MX02 U460 ( .S(n11), .A0(fifo_out[44]), .A1(n110), .Z(gcm_kdf_data[43]));
Q_AN02 U461 ( .A0(n4), .A1(n495), .Z(n110));
Q_MX02 U462 ( .S(n11), .A0(fifo_out[43]), .A1(n111), .Z(gcm_kdf_data[42]));
Q_AN02 U463 ( .A0(n4), .A1(n496), .Z(n111));
Q_MX02 U464 ( .S(n11), .A0(fifo_out[42]), .A1(n112), .Z(gcm_kdf_data[41]));
Q_AN02 U465 ( .A0(n4), .A1(n497), .Z(n112));
Q_MX02 U466 ( .S(n11), .A0(fifo_out[41]), .A1(n113), .Z(gcm_kdf_data[40]));
Q_AN02 U467 ( .A0(n4), .A1(n498), .Z(n113));
Q_MX02 U468 ( .S(n11), .A0(fifo_out[40]), .A1(n114), .Z(gcm_kdf_data[39]));
Q_AN02 U469 ( .A0(n4), .A1(n499), .Z(n114));
Q_MX02 U470 ( .S(n11), .A0(fifo_out[39]), .A1(n115), .Z(gcm_kdf_data[38]));
Q_AN02 U471 ( .A0(n4), .A1(n500), .Z(n115));
Q_MX02 U472 ( .S(n11), .A0(fifo_out[38]), .A1(n116), .Z(gcm_kdf_data[37]));
Q_AN02 U473 ( .A0(n4), .A1(n501), .Z(n116));
Q_MX02 U474 ( .S(n11), .A0(fifo_out[37]), .A1(n117), .Z(gcm_kdf_data[36]));
Q_AN02 U475 ( .A0(n4), .A1(n502), .Z(n117));
Q_MX02 U476 ( .S(n11), .A0(fifo_out[36]), .A1(n118), .Z(gcm_kdf_data[35]));
Q_AN02 U477 ( .A0(n4), .A1(n503), .Z(n118));
Q_MX02 U478 ( .S(n11), .A0(fifo_out[35]), .A1(n119), .Z(gcm_kdf_data[34]));
Q_AN02 U479 ( .A0(n4), .A1(n504), .Z(n119));
Q_MX02 U480 ( .S(n11), .A0(fifo_out[34]), .A1(n120), .Z(gcm_kdf_data[33]));
Q_AN02 U481 ( .A0(n4), .A1(n505), .Z(n120));
Q_MX02 U482 ( .S(n11), .A0(fifo_out[33]), .A1(n121), .Z(gcm_kdf_data[32]));
Q_AN02 U483 ( .A0(n4), .A1(n506), .Z(n121));
Q_MX02 U484 ( .S(n11), .A0(fifo_out[32]), .A1(n122), .Z(gcm_kdf_data[31]));
Q_AN02 U485 ( .A0(n4), .A1(n507), .Z(n122));
Q_MX02 U486 ( .S(n11), .A0(fifo_out[31]), .A1(n123), .Z(gcm_kdf_data[30]));
Q_AN02 U487 ( .A0(n4), .A1(n508), .Z(n123));
Q_MX02 U488 ( .S(n11), .A0(fifo_out[30]), .A1(n124), .Z(gcm_kdf_data[29]));
Q_AN02 U489 ( .A0(n4), .A1(n509), .Z(n124));
Q_MX02 U490 ( .S(n11), .A0(fifo_out[29]), .A1(n125), .Z(gcm_kdf_data[28]));
Q_AN02 U491 ( .A0(n4), .A1(n510), .Z(n125));
Q_MX02 U492 ( .S(n11), .A0(fifo_out[28]), .A1(n126), .Z(gcm_kdf_data[27]));
Q_AN02 U493 ( .A0(n4), .A1(n511), .Z(n126));
Q_MX02 U494 ( .S(n11), .A0(fifo_out[27]), .A1(n127), .Z(gcm_kdf_data[26]));
Q_AN02 U495 ( .A0(n4), .A1(n512), .Z(n127));
Q_MX02 U496 ( .S(n11), .A0(fifo_out[26]), .A1(n128), .Z(gcm_kdf_data[25]));
Q_AN02 U497 ( .A0(n4), .A1(n513), .Z(n128));
Q_MX02 U498 ( .S(n11), .A0(fifo_out[25]), .A1(n129), .Z(gcm_kdf_data[24]));
Q_AN02 U499 ( .A0(n4), .A1(n514), .Z(n129));
Q_MX02 U500 ( .S(n11), .A0(fifo_out[24]), .A1(n130), .Z(gcm_kdf_data[23]));
Q_AN02 U501 ( .A0(n4), .A1(n515), .Z(n130));
Q_MX02 U502 ( .S(n11), .A0(fifo_out[23]), .A1(n131), .Z(gcm_kdf_data[22]));
Q_AN02 U503 ( .A0(n4), .A1(n516), .Z(n131));
Q_MX02 U504 ( .S(n11), .A0(fifo_out[22]), .A1(n132), .Z(gcm_kdf_data[21]));
Q_AN02 U505 ( .A0(n4), .A1(n517), .Z(n132));
Q_MX02 U506 ( .S(n11), .A0(fifo_out[21]), .A1(n133), .Z(gcm_kdf_data[20]));
Q_AN02 U507 ( .A0(n4), .A1(n518), .Z(n133));
Q_MX02 U508 ( .S(n11), .A0(fifo_out[20]), .A1(n134), .Z(gcm_kdf_data[19]));
Q_AN02 U509 ( .A0(n4), .A1(n519), .Z(n134));
Q_MX02 U510 ( .S(n11), .A0(fifo_out[19]), .A1(n135), .Z(gcm_kdf_data[18]));
Q_AN02 U511 ( .A0(n4), .A1(n520), .Z(n135));
Q_MX02 U512 ( .S(n11), .A0(fifo_out[18]), .A1(n136), .Z(gcm_kdf_data[17]));
Q_AN02 U513 ( .A0(n4), .A1(n521), .Z(n136));
Q_MX02 U514 ( .S(n11), .A0(fifo_out[17]), .A1(n137), .Z(gcm_kdf_data[16]));
Q_AN02 U515 ( .A0(n4), .A1(n522), .Z(n137));
Q_MX02 U516 ( .S(n11), .A0(fifo_out[16]), .A1(n138), .Z(gcm_kdf_data[15]));
Q_AN02 U517 ( .A0(n4), .A1(n523), .Z(n138));
Q_MX02 U518 ( .S(n11), .A0(fifo_out[15]), .A1(n139), .Z(gcm_kdf_data[14]));
Q_AN02 U519 ( .A0(n4), .A1(n524), .Z(n139));
Q_MX02 U520 ( .S(n11), .A0(fifo_out[14]), .A1(n140), .Z(gcm_kdf_data[13]));
Q_AN02 U521 ( .A0(n4), .A1(n525), .Z(n140));
Q_MX02 U522 ( .S(n11), .A0(fifo_out[13]), .A1(n141), .Z(gcm_kdf_data[12]));
Q_AN02 U523 ( .A0(n4), .A1(n526), .Z(n141));
Q_MX02 U524 ( .S(n11), .A0(fifo_out[12]), .A1(n142), .Z(gcm_kdf_data[11]));
Q_AN02 U525 ( .A0(n4), .A1(n527), .Z(n142));
Q_MX02 U526 ( .S(n11), .A0(fifo_out[11]), .A1(n143), .Z(gcm_kdf_data[10]));
Q_AN02 U527 ( .A0(n4), .A1(n528), .Z(n143));
Q_MX02 U528 ( .S(n11), .A0(fifo_out[10]), .A1(n144), .Z(gcm_kdf_data[9]));
Q_AN02 U529 ( .A0(n4), .A1(n529), .Z(n144));
Q_MX02 U530 ( .S(n11), .A0(fifo_out[9]), .A1(n145), .Z(gcm_kdf_data[8]));
Q_AN02 U531 ( .A0(n4), .A1(n530), .Z(n145));
Q_MX02 U532 ( .S(n11), .A0(fifo_out[8]), .A1(n146), .Z(gcm_kdf_data[7]));
Q_AN02 U533 ( .A0(n4), .A1(n531), .Z(n146));
Q_MX02 U534 ( .S(n11), .A0(fifo_out[7]), .A1(n147), .Z(gcm_kdf_data[6]));
Q_AN02 U535 ( .A0(n4), .A1(n532), .Z(n147));
Q_MX02 U536 ( .S(n11), .A0(fifo_out[6]), .A1(n148), .Z(gcm_kdf_data[5]));
Q_AN02 U537 ( .A0(n4), .A1(n533), .Z(n148));
Q_MX02 U538 ( .S(n11), .A0(fifo_out[5]), .A1(n149), .Z(gcm_kdf_data[4]));
Q_AN02 U539 ( .A0(n4), .A1(n534), .Z(n149));
Q_MX02 U540 ( .S(n11), .A0(fifo_out[4]), .A1(n150), .Z(gcm_kdf_data[3]));
Q_AN02 U541 ( .A0(n4), .A1(n535), .Z(n150));
Q_MX02 U542 ( .S(n11), .A0(fifo_out[3]), .A1(n151), .Z(gcm_kdf_data[2]));
Q_AN02 U543 ( .A0(n4), .A1(n536), .Z(n151));
Q_MX02 U544 ( .S(n11), .A0(fifo_out[2]), .A1(n152), .Z(gcm_kdf_data[1]));
Q_AN02 U545 ( .A0(n4), .A1(n537), .Z(n152));
Q_MX02 U546 ( .S(n11), .A0(fifo_out[1]), .A1(n153), .Z(gcm_kdf_data[0]));
Q_AN02 U547 ( .A0(n4), .A1(n538), .Z(n153));
Q_MX02 U548 ( .S(n16), .A0(kdf_gcm_stall), .A1(n154), .Z(ciph_out_stall));
Q_AN02 U549 ( .A0(n5), .A1(gcm_status_data_in_stall), .Z(n154));
Q_AN02 U550 ( .A0(n6), .A1(n283), .Z(operand_X[127]));
Q_AN02 U551 ( .A0(n6), .A1(n284), .Z(operand_X[126]));
Q_AN02 U552 ( .A0(n6), .A1(n285), .Z(operand_X[125]));
Q_AN02 U553 ( .A0(n6), .A1(n286), .Z(operand_X[124]));
Q_AN02 U554 ( .A0(n6), .A1(n287), .Z(operand_X[123]));
Q_AN02 U555 ( .A0(n6), .A1(n288), .Z(operand_X[122]));
Q_AN02 U556 ( .A0(n6), .A1(n289), .Z(operand_X[121]));
Q_AN02 U557 ( .A0(n6), .A1(n290), .Z(operand_X[120]));
Q_AN02 U558 ( .A0(n6), .A1(n291), .Z(operand_X[119]));
Q_AN02 U559 ( .A0(n6), .A1(n292), .Z(operand_X[118]));
Q_AN02 U560 ( .A0(n6), .A1(n293), .Z(operand_X[117]));
Q_AN02 U561 ( .A0(n6), .A1(n294), .Z(operand_X[116]));
Q_AN02 U562 ( .A0(n6), .A1(n295), .Z(operand_X[115]));
Q_AN02 U563 ( .A0(n6), .A1(n296), .Z(operand_X[114]));
Q_AN02 U564 ( .A0(n6), .A1(n297), .Z(operand_X[113]));
Q_AN02 U565 ( .A0(n6), .A1(n298), .Z(operand_X[112]));
Q_AN02 U566 ( .A0(n6), .A1(n299), .Z(operand_X[111]));
Q_AN02 U567 ( .A0(n6), .A1(n300), .Z(operand_X[110]));
Q_AN02 U568 ( .A0(n6), .A1(n301), .Z(operand_X[109]));
Q_AN02 U569 ( .A0(n6), .A1(n302), .Z(operand_X[108]));
Q_AN02 U570 ( .A0(n6), .A1(n303), .Z(operand_X[107]));
Q_AN02 U571 ( .A0(n6), .A1(n304), .Z(operand_X[106]));
Q_AN02 U572 ( .A0(n6), .A1(n305), .Z(operand_X[105]));
Q_AN02 U573 ( .A0(n6), .A1(n306), .Z(operand_X[104]));
Q_AN02 U574 ( .A0(n6), .A1(n307), .Z(operand_X[103]));
Q_AN02 U575 ( .A0(n6), .A1(n308), .Z(operand_X[102]));
Q_AN02 U576 ( .A0(n6), .A1(n309), .Z(operand_X[101]));
Q_AN02 U577 ( .A0(n6), .A1(n310), .Z(operand_X[100]));
Q_AN02 U578 ( .A0(n6), .A1(n311), .Z(operand_X[99]));
Q_AN02 U579 ( .A0(n6), .A1(n312), .Z(operand_X[98]));
Q_AN02 U580 ( .A0(n6), .A1(n313), .Z(operand_X[97]));
Q_AN02 U581 ( .A0(n6), .A1(n314), .Z(operand_X[96]));
Q_AN02 U582 ( .A0(n6), .A1(n315), .Z(operand_X[95]));
Q_AN02 U583 ( .A0(n6), .A1(n316), .Z(operand_X[94]));
Q_AN02 U584 ( .A0(n6), .A1(n317), .Z(operand_X[93]));
Q_AN02 U585 ( .A0(n6), .A1(n318), .Z(operand_X[92]));
Q_AN02 U586 ( .A0(n6), .A1(n319), .Z(operand_X[91]));
Q_AN02 U587 ( .A0(n6), .A1(n320), .Z(operand_X[90]));
Q_AN02 U588 ( .A0(n6), .A1(n321), .Z(operand_X[89]));
Q_AN02 U589 ( .A0(n6), .A1(n322), .Z(operand_X[88]));
Q_AN02 U590 ( .A0(n6), .A1(n323), .Z(operand_X[87]));
Q_AN02 U591 ( .A0(n6), .A1(n324), .Z(operand_X[86]));
Q_AN02 U592 ( .A0(n6), .A1(n325), .Z(operand_X[85]));
Q_AN02 U593 ( .A0(n6), .A1(n326), .Z(operand_X[84]));
Q_AN02 U594 ( .A0(n6), .A1(n327), .Z(operand_X[83]));
Q_AN02 U595 ( .A0(n6), .A1(n328), .Z(operand_X[82]));
Q_AN02 U596 ( .A0(n6), .A1(n329), .Z(operand_X[81]));
Q_AN02 U597 ( .A0(n6), .A1(n330), .Z(operand_X[80]));
Q_AN02 U598 ( .A0(n6), .A1(n331), .Z(operand_X[79]));
Q_AN02 U599 ( .A0(n6), .A1(n332), .Z(operand_X[78]));
Q_AN02 U600 ( .A0(n6), .A1(n333), .Z(operand_X[77]));
Q_AN02 U601 ( .A0(n6), .A1(n334), .Z(operand_X[76]));
Q_AN02 U602 ( .A0(n6), .A1(n335), .Z(operand_X[75]));
Q_AN02 U603 ( .A0(n6), .A1(n336), .Z(operand_X[74]));
Q_AN02 U604 ( .A0(n6), .A1(n337), .Z(operand_X[73]));
Q_AN02 U605 ( .A0(n6), .A1(n338), .Z(operand_X[72]));
Q_AN02 U606 ( .A0(n6), .A1(n339), .Z(operand_X[71]));
Q_AN02 U607 ( .A0(n6), .A1(n340), .Z(operand_X[70]));
Q_AN02 U608 ( .A0(n6), .A1(n341), .Z(operand_X[69]));
Q_AN02 U609 ( .A0(n6), .A1(n342), .Z(operand_X[68]));
Q_AN02 U610 ( .A0(n6), .A1(n343), .Z(operand_X[67]));
Q_AN02 U611 ( .A0(n6), .A1(n344), .Z(operand_X[66]));
Q_AN02 U612 ( .A0(n6), .A1(n345), .Z(operand_X[65]));
Q_AN02 U613 ( .A0(n6), .A1(n346), .Z(operand_X[64]));
Q_AN02 U614 ( .A0(n6), .A1(n347), .Z(operand_X[63]));
Q_AN02 U615 ( .A0(n6), .A1(n348), .Z(operand_X[62]));
Q_AN02 U616 ( .A0(n6), .A1(n349), .Z(operand_X[61]));
Q_AN02 U617 ( .A0(n6), .A1(n350), .Z(operand_X[60]));
Q_AN02 U618 ( .A0(n6), .A1(n351), .Z(operand_X[59]));
Q_AN02 U619 ( .A0(n6), .A1(n352), .Z(operand_X[58]));
Q_AN02 U620 ( .A0(n6), .A1(n353), .Z(operand_X[57]));
Q_AN02 U621 ( .A0(n6), .A1(n354), .Z(operand_X[56]));
Q_AN02 U622 ( .A0(n6), .A1(n355), .Z(operand_X[55]));
Q_AN02 U623 ( .A0(n6), .A1(n356), .Z(operand_X[54]));
Q_AN02 U624 ( .A0(n6), .A1(n357), .Z(operand_X[53]));
Q_AN02 U625 ( .A0(n6), .A1(n358), .Z(operand_X[52]));
Q_AN02 U626 ( .A0(n6), .A1(n359), .Z(operand_X[51]));
Q_AN02 U627 ( .A0(n6), .A1(n360), .Z(operand_X[50]));
Q_AN02 U628 ( .A0(n6), .A1(n361), .Z(operand_X[49]));
Q_AN02 U629 ( .A0(n6), .A1(n362), .Z(operand_X[48]));
Q_AN02 U630 ( .A0(n6), .A1(n363), .Z(operand_X[47]));
Q_AN02 U631 ( .A0(n6), .A1(n364), .Z(operand_X[46]));
Q_AN02 U632 ( .A0(n6), .A1(n365), .Z(operand_X[45]));
Q_AN02 U633 ( .A0(n6), .A1(n366), .Z(operand_X[44]));
Q_AN02 U634 ( .A0(n6), .A1(n367), .Z(operand_X[43]));
Q_AN02 U635 ( .A0(n6), .A1(n368), .Z(operand_X[42]));
Q_AN02 U636 ( .A0(n6), .A1(n369), .Z(operand_X[41]));
Q_AN02 U637 ( .A0(n6), .A1(n370), .Z(operand_X[40]));
Q_AN02 U638 ( .A0(n6), .A1(n371), .Z(operand_X[39]));
Q_AN02 U639 ( .A0(n6), .A1(n372), .Z(operand_X[38]));
Q_AN02 U640 ( .A0(n6), .A1(n373), .Z(operand_X[37]));
Q_AN02 U641 ( .A0(n6), .A1(n374), .Z(operand_X[36]));
Q_AN02 U642 ( .A0(n6), .A1(n375), .Z(operand_X[35]));
Q_AN02 U643 ( .A0(n6), .A1(n376), .Z(operand_X[34]));
Q_AN02 U644 ( .A0(n6), .A1(n377), .Z(operand_X[33]));
Q_AN02 U645 ( .A0(n6), .A1(n378), .Z(operand_X[32]));
Q_AN02 U646 ( .A0(n6), .A1(n379), .Z(operand_X[31]));
Q_AN02 U647 ( .A0(n6), .A1(n380), .Z(operand_X[30]));
Q_AN02 U648 ( .A0(n6), .A1(n381), .Z(operand_X[29]));
Q_AN02 U649 ( .A0(n6), .A1(n382), .Z(operand_X[28]));
Q_AN02 U650 ( .A0(n6), .A1(n383), .Z(operand_X[27]));
Q_AN02 U651 ( .A0(n6), .A1(n384), .Z(operand_X[26]));
Q_AN02 U652 ( .A0(n6), .A1(n385), .Z(operand_X[25]));
Q_AN02 U653 ( .A0(n6), .A1(n386), .Z(operand_X[24]));
Q_AN02 U654 ( .A0(n6), .A1(n387), .Z(operand_X[23]));
Q_AN02 U655 ( .A0(n6), .A1(n388), .Z(operand_X[22]));
Q_AN02 U656 ( .A0(n6), .A1(n389), .Z(operand_X[21]));
Q_AN02 U657 ( .A0(n6), .A1(n390), .Z(operand_X[20]));
Q_AN02 U658 ( .A0(n6), .A1(n391), .Z(operand_X[19]));
Q_AN02 U659 ( .A0(n6), .A1(n392), .Z(operand_X[18]));
Q_AN02 U660 ( .A0(n6), .A1(n393), .Z(operand_X[17]));
Q_AN02 U661 ( .A0(n6), .A1(n394), .Z(operand_X[16]));
Q_AN02 U662 ( .A0(n6), .A1(n395), .Z(operand_X[15]));
Q_AN02 U663 ( .A0(n6), .A1(n396), .Z(operand_X[14]));
Q_AN02 U664 ( .A0(n6), .A1(n397), .Z(operand_X[13]));
Q_AN02 U665 ( .A0(n6), .A1(n398), .Z(operand_X[12]));
Q_AN02 U666 ( .A0(n6), .A1(n399), .Z(operand_X[11]));
Q_AN02 U667 ( .A0(n6), .A1(n400), .Z(operand_X[10]));
Q_AN02 U668 ( .A0(n6), .A1(n401), .Z(operand_X[9]));
Q_AN02 U669 ( .A0(n6), .A1(n402), .Z(operand_X[8]));
Q_AN02 U670 ( .A0(n6), .A1(n403), .Z(operand_X[7]));
Q_AN02 U671 ( .A0(n6), .A1(n404), .Z(operand_X[6]));
Q_AN02 U672 ( .A0(n6), .A1(n405), .Z(operand_X[5]));
Q_AN02 U673 ( .A0(n6), .A1(n406), .Z(operand_X[4]));
Q_AN02 U674 ( .A0(n6), .A1(n407), .Z(operand_X[3]));
Q_AN02 U675 ( .A0(n6), .A1(n408), .Z(operand_X[2]));
Q_AN02 U676 ( .A0(n6), .A1(n409), .Z(operand_X[1]));
Q_AN02 U677 ( .A0(n6), .A1(n410), .Z(operand_X[0]));
Q_MX02 U678 ( .S(n19), .A0(ciph_out[127]), .A1(operand_Y[127]), .Z(nxt_h_value[127]));
Q_MX02 U679 ( .S(n19), .A0(ciph_out[126]), .A1(operand_Y[126]), .Z(nxt_h_value[126]));
Q_MX02 U680 ( .S(n19), .A0(ciph_out[125]), .A1(operand_Y[125]), .Z(nxt_h_value[125]));
Q_MX02 U681 ( .S(n19), .A0(ciph_out[124]), .A1(operand_Y[124]), .Z(nxt_h_value[124]));
Q_MX02 U682 ( .S(n19), .A0(ciph_out[123]), .A1(operand_Y[123]), .Z(nxt_h_value[123]));
Q_MX02 U683 ( .S(n19), .A0(ciph_out[122]), .A1(operand_Y[122]), .Z(nxt_h_value[122]));
Q_MX02 U684 ( .S(n19), .A0(ciph_out[121]), .A1(operand_Y[121]), .Z(nxt_h_value[121]));
Q_MX02 U685 ( .S(n19), .A0(ciph_out[120]), .A1(operand_Y[120]), .Z(nxt_h_value[120]));
Q_MX02 U686 ( .S(n19), .A0(ciph_out[119]), .A1(operand_Y[119]), .Z(nxt_h_value[119]));
Q_MX02 U687 ( .S(n19), .A0(ciph_out[118]), .A1(operand_Y[118]), .Z(nxt_h_value[118]));
Q_MX02 U688 ( .S(n19), .A0(ciph_out[117]), .A1(operand_Y[117]), .Z(nxt_h_value[117]));
Q_MX02 U689 ( .S(n19), .A0(ciph_out[116]), .A1(operand_Y[116]), .Z(nxt_h_value[116]));
Q_MX02 U690 ( .S(n19), .A0(ciph_out[115]), .A1(operand_Y[115]), .Z(nxt_h_value[115]));
Q_MX02 U691 ( .S(n19), .A0(ciph_out[114]), .A1(operand_Y[114]), .Z(nxt_h_value[114]));
Q_MX02 U692 ( .S(n19), .A0(ciph_out[113]), .A1(operand_Y[113]), .Z(nxt_h_value[113]));
Q_MX02 U693 ( .S(n19), .A0(ciph_out[112]), .A1(operand_Y[112]), .Z(nxt_h_value[112]));
Q_MX02 U694 ( .S(n19), .A0(ciph_out[111]), .A1(operand_Y[111]), .Z(nxt_h_value[111]));
Q_MX02 U695 ( .S(n19), .A0(ciph_out[110]), .A1(operand_Y[110]), .Z(nxt_h_value[110]));
Q_MX02 U696 ( .S(n19), .A0(ciph_out[109]), .A1(operand_Y[109]), .Z(nxt_h_value[109]));
Q_MX02 U697 ( .S(n19), .A0(ciph_out[108]), .A1(operand_Y[108]), .Z(nxt_h_value[108]));
Q_MX02 U698 ( .S(n19), .A0(ciph_out[107]), .A1(operand_Y[107]), .Z(nxt_h_value[107]));
Q_MX02 U699 ( .S(n19), .A0(ciph_out[106]), .A1(operand_Y[106]), .Z(nxt_h_value[106]));
Q_MX02 U700 ( .S(n19), .A0(ciph_out[105]), .A1(operand_Y[105]), .Z(nxt_h_value[105]));
Q_MX02 U701 ( .S(n19), .A0(ciph_out[104]), .A1(operand_Y[104]), .Z(nxt_h_value[104]));
Q_MX02 U702 ( .S(n19), .A0(ciph_out[103]), .A1(operand_Y[103]), .Z(nxt_h_value[103]));
Q_MX02 U703 ( .S(n19), .A0(ciph_out[102]), .A1(operand_Y[102]), .Z(nxt_h_value[102]));
Q_MX02 U704 ( .S(n19), .A0(ciph_out[101]), .A1(operand_Y[101]), .Z(nxt_h_value[101]));
Q_MX02 U705 ( .S(n19), .A0(ciph_out[100]), .A1(operand_Y[100]), .Z(nxt_h_value[100]));
Q_MX02 U706 ( .S(n19), .A0(ciph_out[99]), .A1(operand_Y[99]), .Z(nxt_h_value[99]));
Q_MX02 U707 ( .S(n19), .A0(ciph_out[98]), .A1(operand_Y[98]), .Z(nxt_h_value[98]));
Q_MX02 U708 ( .S(n19), .A0(ciph_out[97]), .A1(operand_Y[97]), .Z(nxt_h_value[97]));
Q_MX02 U709 ( .S(n19), .A0(ciph_out[96]), .A1(operand_Y[96]), .Z(nxt_h_value[96]));
Q_MX02 U710 ( .S(n19), .A0(ciph_out[95]), .A1(operand_Y[95]), .Z(nxt_h_value[95]));
Q_MX02 U711 ( .S(n19), .A0(ciph_out[94]), .A1(operand_Y[94]), .Z(nxt_h_value[94]));
Q_MX02 U712 ( .S(n19), .A0(ciph_out[93]), .A1(operand_Y[93]), .Z(nxt_h_value[93]));
Q_MX02 U713 ( .S(n19), .A0(ciph_out[92]), .A1(operand_Y[92]), .Z(nxt_h_value[92]));
Q_MX02 U714 ( .S(n19), .A0(ciph_out[91]), .A1(operand_Y[91]), .Z(nxt_h_value[91]));
Q_MX02 U715 ( .S(n19), .A0(ciph_out[90]), .A1(operand_Y[90]), .Z(nxt_h_value[90]));
Q_MX02 U716 ( .S(n19), .A0(ciph_out[89]), .A1(operand_Y[89]), .Z(nxt_h_value[89]));
Q_MX02 U717 ( .S(n19), .A0(ciph_out[88]), .A1(operand_Y[88]), .Z(nxt_h_value[88]));
Q_MX02 U718 ( .S(n19), .A0(ciph_out[87]), .A1(operand_Y[87]), .Z(nxt_h_value[87]));
Q_MX02 U719 ( .S(n19), .A0(ciph_out[86]), .A1(operand_Y[86]), .Z(nxt_h_value[86]));
Q_MX02 U720 ( .S(n19), .A0(ciph_out[85]), .A1(operand_Y[85]), .Z(nxt_h_value[85]));
Q_MX02 U721 ( .S(n19), .A0(ciph_out[84]), .A1(operand_Y[84]), .Z(nxt_h_value[84]));
Q_MX02 U722 ( .S(n19), .A0(ciph_out[83]), .A1(operand_Y[83]), .Z(nxt_h_value[83]));
Q_MX02 U723 ( .S(n19), .A0(ciph_out[82]), .A1(operand_Y[82]), .Z(nxt_h_value[82]));
Q_MX02 U724 ( .S(n19), .A0(ciph_out[81]), .A1(operand_Y[81]), .Z(nxt_h_value[81]));
Q_MX02 U725 ( .S(n19), .A0(ciph_out[80]), .A1(operand_Y[80]), .Z(nxt_h_value[80]));
Q_MX02 U726 ( .S(n19), .A0(ciph_out[79]), .A1(operand_Y[79]), .Z(nxt_h_value[79]));
Q_MX02 U727 ( .S(n19), .A0(ciph_out[78]), .A1(operand_Y[78]), .Z(nxt_h_value[78]));
Q_MX02 U728 ( .S(n19), .A0(ciph_out[77]), .A1(operand_Y[77]), .Z(nxt_h_value[77]));
Q_MX02 U729 ( .S(n19), .A0(ciph_out[76]), .A1(operand_Y[76]), .Z(nxt_h_value[76]));
Q_MX02 U730 ( .S(n19), .A0(ciph_out[75]), .A1(operand_Y[75]), .Z(nxt_h_value[75]));
Q_MX02 U731 ( .S(n19), .A0(ciph_out[74]), .A1(operand_Y[74]), .Z(nxt_h_value[74]));
Q_MX02 U732 ( .S(n19), .A0(ciph_out[73]), .A1(operand_Y[73]), .Z(nxt_h_value[73]));
Q_MX02 U733 ( .S(n19), .A0(ciph_out[72]), .A1(operand_Y[72]), .Z(nxt_h_value[72]));
Q_MX02 U734 ( .S(n19), .A0(ciph_out[71]), .A1(operand_Y[71]), .Z(nxt_h_value[71]));
Q_MX02 U735 ( .S(n19), .A0(ciph_out[70]), .A1(operand_Y[70]), .Z(nxt_h_value[70]));
Q_MX02 U736 ( .S(n19), .A0(ciph_out[69]), .A1(operand_Y[69]), .Z(nxt_h_value[69]));
Q_MX02 U737 ( .S(n19), .A0(ciph_out[68]), .A1(operand_Y[68]), .Z(nxt_h_value[68]));
Q_MX02 U738 ( .S(n19), .A0(ciph_out[67]), .A1(operand_Y[67]), .Z(nxt_h_value[67]));
Q_MX02 U739 ( .S(n19), .A0(ciph_out[66]), .A1(operand_Y[66]), .Z(nxt_h_value[66]));
Q_MX02 U740 ( .S(n19), .A0(ciph_out[65]), .A1(operand_Y[65]), .Z(nxt_h_value[65]));
Q_MX02 U741 ( .S(n19), .A0(ciph_out[64]), .A1(operand_Y[64]), .Z(nxt_h_value[64]));
Q_MX02 U742 ( .S(n19), .A0(ciph_out[63]), .A1(operand_Y[63]), .Z(nxt_h_value[63]));
Q_MX02 U743 ( .S(n19), .A0(ciph_out[62]), .A1(operand_Y[62]), .Z(nxt_h_value[62]));
Q_MX02 U744 ( .S(n19), .A0(ciph_out[61]), .A1(operand_Y[61]), .Z(nxt_h_value[61]));
Q_MX02 U745 ( .S(n19), .A0(ciph_out[60]), .A1(operand_Y[60]), .Z(nxt_h_value[60]));
Q_MX02 U746 ( .S(n19), .A0(ciph_out[59]), .A1(operand_Y[59]), .Z(nxt_h_value[59]));
Q_MX02 U747 ( .S(n19), .A0(ciph_out[58]), .A1(operand_Y[58]), .Z(nxt_h_value[58]));
Q_MX02 U748 ( .S(n19), .A0(ciph_out[57]), .A1(operand_Y[57]), .Z(nxt_h_value[57]));
Q_MX02 U749 ( .S(n19), .A0(ciph_out[56]), .A1(operand_Y[56]), .Z(nxt_h_value[56]));
Q_MX02 U750 ( .S(n19), .A0(ciph_out[55]), .A1(operand_Y[55]), .Z(nxt_h_value[55]));
Q_MX02 U751 ( .S(n19), .A0(ciph_out[54]), .A1(operand_Y[54]), .Z(nxt_h_value[54]));
Q_MX02 U752 ( .S(n19), .A0(ciph_out[53]), .A1(operand_Y[53]), .Z(nxt_h_value[53]));
Q_MX02 U753 ( .S(n19), .A0(ciph_out[52]), .A1(operand_Y[52]), .Z(nxt_h_value[52]));
Q_MX02 U754 ( .S(n19), .A0(ciph_out[51]), .A1(operand_Y[51]), .Z(nxt_h_value[51]));
Q_MX02 U755 ( .S(n19), .A0(ciph_out[50]), .A1(operand_Y[50]), .Z(nxt_h_value[50]));
Q_MX02 U756 ( .S(n19), .A0(ciph_out[49]), .A1(operand_Y[49]), .Z(nxt_h_value[49]));
Q_MX02 U757 ( .S(n19), .A0(ciph_out[48]), .A1(operand_Y[48]), .Z(nxt_h_value[48]));
Q_MX02 U758 ( .S(n19), .A0(ciph_out[47]), .A1(operand_Y[47]), .Z(nxt_h_value[47]));
Q_MX02 U759 ( .S(n19), .A0(ciph_out[46]), .A1(operand_Y[46]), .Z(nxt_h_value[46]));
Q_MX02 U760 ( .S(n19), .A0(ciph_out[45]), .A1(operand_Y[45]), .Z(nxt_h_value[45]));
Q_MX02 U761 ( .S(n19), .A0(ciph_out[44]), .A1(operand_Y[44]), .Z(nxt_h_value[44]));
Q_MX02 U762 ( .S(n19), .A0(ciph_out[43]), .A1(operand_Y[43]), .Z(nxt_h_value[43]));
Q_MX02 U763 ( .S(n19), .A0(ciph_out[42]), .A1(operand_Y[42]), .Z(nxt_h_value[42]));
Q_MX02 U764 ( .S(n19), .A0(ciph_out[41]), .A1(operand_Y[41]), .Z(nxt_h_value[41]));
Q_MX02 U765 ( .S(n19), .A0(ciph_out[40]), .A1(operand_Y[40]), .Z(nxt_h_value[40]));
Q_MX02 U766 ( .S(n19), .A0(ciph_out[39]), .A1(operand_Y[39]), .Z(nxt_h_value[39]));
Q_MX02 U767 ( .S(n19), .A0(ciph_out[38]), .A1(operand_Y[38]), .Z(nxt_h_value[38]));
Q_MX02 U768 ( .S(n19), .A0(ciph_out[37]), .A1(operand_Y[37]), .Z(nxt_h_value[37]));
Q_MX02 U769 ( .S(n19), .A0(ciph_out[36]), .A1(operand_Y[36]), .Z(nxt_h_value[36]));
Q_MX02 U770 ( .S(n19), .A0(ciph_out[35]), .A1(operand_Y[35]), .Z(nxt_h_value[35]));
Q_MX02 U771 ( .S(n19), .A0(ciph_out[34]), .A1(operand_Y[34]), .Z(nxt_h_value[34]));
Q_MX02 U772 ( .S(n19), .A0(ciph_out[33]), .A1(operand_Y[33]), .Z(nxt_h_value[33]));
Q_MX02 U773 ( .S(n19), .A0(ciph_out[32]), .A1(operand_Y[32]), .Z(nxt_h_value[32]));
Q_MX02 U774 ( .S(n19), .A0(ciph_out[31]), .A1(operand_Y[31]), .Z(nxt_h_value[31]));
Q_MX02 U775 ( .S(n19), .A0(ciph_out[30]), .A1(operand_Y[30]), .Z(nxt_h_value[30]));
Q_MX02 U776 ( .S(n19), .A0(ciph_out[29]), .A1(operand_Y[29]), .Z(nxt_h_value[29]));
Q_MX02 U777 ( .S(n19), .A0(ciph_out[28]), .A1(operand_Y[28]), .Z(nxt_h_value[28]));
Q_MX02 U778 ( .S(n19), .A0(ciph_out[27]), .A1(operand_Y[27]), .Z(nxt_h_value[27]));
Q_MX02 U779 ( .S(n19), .A0(ciph_out[26]), .A1(operand_Y[26]), .Z(nxt_h_value[26]));
Q_MX02 U780 ( .S(n19), .A0(ciph_out[25]), .A1(operand_Y[25]), .Z(nxt_h_value[25]));
Q_MX02 U781 ( .S(n19), .A0(ciph_out[24]), .A1(operand_Y[24]), .Z(nxt_h_value[24]));
Q_MX02 U782 ( .S(n19), .A0(ciph_out[23]), .A1(operand_Y[23]), .Z(nxt_h_value[23]));
Q_MX02 U783 ( .S(n19), .A0(ciph_out[22]), .A1(operand_Y[22]), .Z(nxt_h_value[22]));
Q_MX02 U784 ( .S(n19), .A0(ciph_out[21]), .A1(operand_Y[21]), .Z(nxt_h_value[21]));
Q_MX02 U785 ( .S(n19), .A0(ciph_out[20]), .A1(operand_Y[20]), .Z(nxt_h_value[20]));
Q_MX02 U786 ( .S(n19), .A0(ciph_out[19]), .A1(operand_Y[19]), .Z(nxt_h_value[19]));
Q_MX02 U787 ( .S(n19), .A0(ciph_out[18]), .A1(operand_Y[18]), .Z(nxt_h_value[18]));
Q_MX02 U788 ( .S(n19), .A0(ciph_out[17]), .A1(operand_Y[17]), .Z(nxt_h_value[17]));
Q_MX02 U789 ( .S(n19), .A0(ciph_out[16]), .A1(operand_Y[16]), .Z(nxt_h_value[16]));
Q_MX02 U790 ( .S(n19), .A0(ciph_out[15]), .A1(operand_Y[15]), .Z(nxt_h_value[15]));
Q_MX02 U791 ( .S(n19), .A0(ciph_out[14]), .A1(operand_Y[14]), .Z(nxt_h_value[14]));
Q_MX02 U792 ( .S(n19), .A0(ciph_out[13]), .A1(operand_Y[13]), .Z(nxt_h_value[13]));
Q_MX02 U793 ( .S(n19), .A0(ciph_out[12]), .A1(operand_Y[12]), .Z(nxt_h_value[12]));
Q_MX02 U794 ( .S(n19), .A0(ciph_out[11]), .A1(operand_Y[11]), .Z(nxt_h_value[11]));
Q_MX02 U795 ( .S(n19), .A0(ciph_out[10]), .A1(operand_Y[10]), .Z(nxt_h_value[10]));
Q_MX02 U796 ( .S(n19), .A0(ciph_out[9]), .A1(operand_Y[9]), .Z(nxt_h_value[9]));
Q_MX02 U797 ( .S(n19), .A0(ciph_out[8]), .A1(operand_Y[8]), .Z(nxt_h_value[8]));
Q_MX02 U798 ( .S(n19), .A0(ciph_out[7]), .A1(operand_Y[7]), .Z(nxt_h_value[7]));
Q_MX02 U799 ( .S(n19), .A0(ciph_out[6]), .A1(operand_Y[6]), .Z(nxt_h_value[6]));
Q_MX02 U800 ( .S(n19), .A0(ciph_out[5]), .A1(operand_Y[5]), .Z(nxt_h_value[5]));
Q_MX02 U801 ( .S(n19), .A0(ciph_out[4]), .A1(operand_Y[4]), .Z(nxt_h_value[4]));
Q_MX02 U802 ( .S(n19), .A0(ciph_out[3]), .A1(operand_Y[3]), .Z(nxt_h_value[3]));
Q_MX02 U803 ( .S(n19), .A0(ciph_out[2]), .A1(operand_Y[2]), .Z(nxt_h_value[2]));
Q_MX02 U804 ( .S(n19), .A0(ciph_out[1]), .A1(operand_Y[1]), .Z(nxt_h_value[1]));
Q_MX02 U805 ( .S(n19), .A0(ciph_out[0]), .A1(operand_Y[0]), .Z(nxt_h_value[0]));
Q_MX02 U806 ( .S(n7), .A0(n155), .A1(auth_tag[127]), .Z(nxt_auth_tag[127]));
Q_AN02 U807 ( .A0(n8), .A1(ciph_out[127]), .Z(n155));
Q_MX02 U808 ( .S(n7), .A0(n156), .A1(auth_tag[126]), .Z(nxt_auth_tag[126]));
Q_AN02 U809 ( .A0(n8), .A1(ciph_out[126]), .Z(n156));
Q_MX02 U810 ( .S(n7), .A0(n157), .A1(auth_tag[125]), .Z(nxt_auth_tag[125]));
Q_AN02 U811 ( .A0(n8), .A1(ciph_out[125]), .Z(n157));
Q_MX02 U812 ( .S(n7), .A0(n158), .A1(auth_tag[124]), .Z(nxt_auth_tag[124]));
Q_AN02 U813 ( .A0(n8), .A1(ciph_out[124]), .Z(n158));
Q_MX02 U814 ( .S(n7), .A0(n159), .A1(auth_tag[123]), .Z(nxt_auth_tag[123]));
Q_AN02 U815 ( .A0(n8), .A1(ciph_out[123]), .Z(n159));
Q_MX02 U816 ( .S(n7), .A0(n160), .A1(auth_tag[122]), .Z(nxt_auth_tag[122]));
Q_AN02 U817 ( .A0(n8), .A1(ciph_out[122]), .Z(n160));
Q_MX02 U818 ( .S(n7), .A0(n161), .A1(auth_tag[121]), .Z(nxt_auth_tag[121]));
Q_AN02 U819 ( .A0(n8), .A1(ciph_out[121]), .Z(n161));
Q_MX02 U820 ( .S(n7), .A0(n162), .A1(auth_tag[120]), .Z(nxt_auth_tag[120]));
Q_AN02 U821 ( .A0(n8), .A1(ciph_out[120]), .Z(n162));
Q_MX02 U822 ( .S(n7), .A0(n163), .A1(auth_tag[119]), .Z(nxt_auth_tag[119]));
Q_AN02 U823 ( .A0(n8), .A1(ciph_out[119]), .Z(n163));
Q_MX02 U824 ( .S(n7), .A0(n164), .A1(auth_tag[118]), .Z(nxt_auth_tag[118]));
Q_AN02 U825 ( .A0(n8), .A1(ciph_out[118]), .Z(n164));
Q_MX02 U826 ( .S(n7), .A0(n165), .A1(auth_tag[117]), .Z(nxt_auth_tag[117]));
Q_AN02 U827 ( .A0(n8), .A1(ciph_out[117]), .Z(n165));
Q_MX02 U828 ( .S(n7), .A0(n166), .A1(auth_tag[116]), .Z(nxt_auth_tag[116]));
Q_AN02 U829 ( .A0(n8), .A1(ciph_out[116]), .Z(n166));
Q_MX02 U830 ( .S(n7), .A0(n167), .A1(auth_tag[115]), .Z(nxt_auth_tag[115]));
Q_AN02 U831 ( .A0(n8), .A1(ciph_out[115]), .Z(n167));
Q_MX02 U832 ( .S(n7), .A0(n168), .A1(auth_tag[114]), .Z(nxt_auth_tag[114]));
Q_AN02 U833 ( .A0(n8), .A1(ciph_out[114]), .Z(n168));
Q_MX02 U834 ( .S(n7), .A0(n169), .A1(auth_tag[113]), .Z(nxt_auth_tag[113]));
Q_AN02 U835 ( .A0(n8), .A1(ciph_out[113]), .Z(n169));
Q_MX02 U836 ( .S(n7), .A0(n170), .A1(auth_tag[112]), .Z(nxt_auth_tag[112]));
Q_AN02 U837 ( .A0(n8), .A1(ciph_out[112]), .Z(n170));
Q_MX02 U838 ( .S(n7), .A0(n171), .A1(auth_tag[111]), .Z(nxt_auth_tag[111]));
Q_AN02 U839 ( .A0(n8), .A1(ciph_out[111]), .Z(n171));
Q_MX02 U840 ( .S(n7), .A0(n172), .A1(auth_tag[110]), .Z(nxt_auth_tag[110]));
Q_AN02 U841 ( .A0(n8), .A1(ciph_out[110]), .Z(n172));
Q_MX02 U842 ( .S(n7), .A0(n173), .A1(auth_tag[109]), .Z(nxt_auth_tag[109]));
Q_AN02 U843 ( .A0(n8), .A1(ciph_out[109]), .Z(n173));
Q_MX02 U844 ( .S(n7), .A0(n174), .A1(auth_tag[108]), .Z(nxt_auth_tag[108]));
Q_AN02 U845 ( .A0(n8), .A1(ciph_out[108]), .Z(n174));
Q_MX02 U846 ( .S(n7), .A0(n175), .A1(auth_tag[107]), .Z(nxt_auth_tag[107]));
Q_AN02 U847 ( .A0(n8), .A1(ciph_out[107]), .Z(n175));
Q_MX02 U848 ( .S(n7), .A0(n176), .A1(auth_tag[106]), .Z(nxt_auth_tag[106]));
Q_AN02 U849 ( .A0(n8), .A1(ciph_out[106]), .Z(n176));
Q_MX02 U850 ( .S(n7), .A0(n177), .A1(auth_tag[105]), .Z(nxt_auth_tag[105]));
Q_AN02 U851 ( .A0(n8), .A1(ciph_out[105]), .Z(n177));
Q_MX02 U852 ( .S(n7), .A0(n178), .A1(auth_tag[104]), .Z(nxt_auth_tag[104]));
Q_AN02 U853 ( .A0(n8), .A1(ciph_out[104]), .Z(n178));
Q_MX02 U854 ( .S(n7), .A0(n179), .A1(auth_tag[103]), .Z(nxt_auth_tag[103]));
Q_AN02 U855 ( .A0(n8), .A1(ciph_out[103]), .Z(n179));
Q_MX02 U856 ( .S(n7), .A0(n180), .A1(auth_tag[102]), .Z(nxt_auth_tag[102]));
Q_AN02 U857 ( .A0(n8), .A1(ciph_out[102]), .Z(n180));
Q_MX02 U858 ( .S(n7), .A0(n181), .A1(auth_tag[101]), .Z(nxt_auth_tag[101]));
Q_AN02 U859 ( .A0(n8), .A1(ciph_out[101]), .Z(n181));
Q_MX02 U860 ( .S(n7), .A0(n182), .A1(auth_tag[100]), .Z(nxt_auth_tag[100]));
Q_AN02 U861 ( .A0(n8), .A1(ciph_out[100]), .Z(n182));
Q_MX02 U862 ( .S(n7), .A0(n183), .A1(auth_tag[99]), .Z(nxt_auth_tag[99]));
Q_AN02 U863 ( .A0(n8), .A1(ciph_out[99]), .Z(n183));
Q_MX02 U864 ( .S(n7), .A0(n184), .A1(auth_tag[98]), .Z(nxt_auth_tag[98]));
Q_AN02 U865 ( .A0(n8), .A1(ciph_out[98]), .Z(n184));
Q_MX02 U866 ( .S(n7), .A0(n185), .A1(auth_tag[97]), .Z(nxt_auth_tag[97]));
Q_AN02 U867 ( .A0(n8), .A1(ciph_out[97]), .Z(n185));
Q_MX02 U868 ( .S(n7), .A0(n186), .A1(auth_tag[96]), .Z(nxt_auth_tag[96]));
Q_AN02 U869 ( .A0(n8), .A1(ciph_out[96]), .Z(n186));
Q_MX02 U870 ( .S(n7), .A0(n187), .A1(auth_tag[95]), .Z(nxt_auth_tag[95]));
Q_AN02 U871 ( .A0(n8), .A1(ciph_out[95]), .Z(n187));
Q_MX02 U872 ( .S(n7), .A0(n188), .A1(auth_tag[94]), .Z(nxt_auth_tag[94]));
Q_AN02 U873 ( .A0(n8), .A1(ciph_out[94]), .Z(n188));
Q_MX02 U874 ( .S(n7), .A0(n189), .A1(auth_tag[93]), .Z(nxt_auth_tag[93]));
Q_AN02 U875 ( .A0(n8), .A1(ciph_out[93]), .Z(n189));
Q_MX02 U876 ( .S(n7), .A0(n190), .A1(auth_tag[92]), .Z(nxt_auth_tag[92]));
Q_AN02 U877 ( .A0(n8), .A1(ciph_out[92]), .Z(n190));
Q_MX02 U878 ( .S(n7), .A0(n191), .A1(auth_tag[91]), .Z(nxt_auth_tag[91]));
Q_AN02 U879 ( .A0(n8), .A1(ciph_out[91]), .Z(n191));
Q_MX02 U880 ( .S(n7), .A0(n192), .A1(auth_tag[90]), .Z(nxt_auth_tag[90]));
Q_AN02 U881 ( .A0(n8), .A1(ciph_out[90]), .Z(n192));
Q_MX02 U882 ( .S(n7), .A0(n193), .A1(auth_tag[89]), .Z(nxt_auth_tag[89]));
Q_AN02 U883 ( .A0(n8), .A1(ciph_out[89]), .Z(n193));
Q_MX02 U884 ( .S(n7), .A0(n194), .A1(auth_tag[88]), .Z(nxt_auth_tag[88]));
Q_AN02 U885 ( .A0(n8), .A1(ciph_out[88]), .Z(n194));
Q_MX02 U886 ( .S(n7), .A0(n195), .A1(auth_tag[87]), .Z(nxt_auth_tag[87]));
Q_AN02 U887 ( .A0(n8), .A1(ciph_out[87]), .Z(n195));
Q_MX02 U888 ( .S(n7), .A0(n196), .A1(auth_tag[86]), .Z(nxt_auth_tag[86]));
Q_AN02 U889 ( .A0(n8), .A1(ciph_out[86]), .Z(n196));
Q_MX02 U890 ( .S(n7), .A0(n197), .A1(auth_tag[85]), .Z(nxt_auth_tag[85]));
Q_AN02 U891 ( .A0(n8), .A1(ciph_out[85]), .Z(n197));
Q_MX02 U892 ( .S(n7), .A0(n198), .A1(auth_tag[84]), .Z(nxt_auth_tag[84]));
Q_AN02 U893 ( .A0(n8), .A1(ciph_out[84]), .Z(n198));
Q_MX02 U894 ( .S(n7), .A0(n199), .A1(auth_tag[83]), .Z(nxt_auth_tag[83]));
Q_AN02 U895 ( .A0(n8), .A1(ciph_out[83]), .Z(n199));
Q_MX02 U896 ( .S(n7), .A0(n200), .A1(auth_tag[82]), .Z(nxt_auth_tag[82]));
Q_AN02 U897 ( .A0(n8), .A1(ciph_out[82]), .Z(n200));
Q_MX02 U898 ( .S(n7), .A0(n201), .A1(auth_tag[81]), .Z(nxt_auth_tag[81]));
Q_AN02 U899 ( .A0(n8), .A1(ciph_out[81]), .Z(n201));
Q_MX02 U900 ( .S(n7), .A0(n202), .A1(auth_tag[80]), .Z(nxt_auth_tag[80]));
Q_AN02 U901 ( .A0(n8), .A1(ciph_out[80]), .Z(n202));
Q_MX02 U902 ( .S(n7), .A0(n203), .A1(auth_tag[79]), .Z(nxt_auth_tag[79]));
Q_AN02 U903 ( .A0(n8), .A1(ciph_out[79]), .Z(n203));
Q_MX02 U904 ( .S(n7), .A0(n204), .A1(auth_tag[78]), .Z(nxt_auth_tag[78]));
Q_AN02 U905 ( .A0(n8), .A1(ciph_out[78]), .Z(n204));
Q_MX02 U906 ( .S(n7), .A0(n205), .A1(auth_tag[77]), .Z(nxt_auth_tag[77]));
Q_AN02 U907 ( .A0(n8), .A1(ciph_out[77]), .Z(n205));
Q_MX02 U908 ( .S(n7), .A0(n206), .A1(auth_tag[76]), .Z(nxt_auth_tag[76]));
Q_AN02 U909 ( .A0(n8), .A1(ciph_out[76]), .Z(n206));
Q_MX02 U910 ( .S(n7), .A0(n207), .A1(auth_tag[75]), .Z(nxt_auth_tag[75]));
Q_AN02 U911 ( .A0(n8), .A1(ciph_out[75]), .Z(n207));
Q_MX02 U912 ( .S(n7), .A0(n208), .A1(auth_tag[74]), .Z(nxt_auth_tag[74]));
Q_AN02 U913 ( .A0(n8), .A1(ciph_out[74]), .Z(n208));
Q_MX02 U914 ( .S(n7), .A0(n209), .A1(auth_tag[73]), .Z(nxt_auth_tag[73]));
Q_AN02 U915 ( .A0(n8), .A1(ciph_out[73]), .Z(n209));
Q_MX02 U916 ( .S(n7), .A0(n210), .A1(auth_tag[72]), .Z(nxt_auth_tag[72]));
Q_AN02 U917 ( .A0(n8), .A1(ciph_out[72]), .Z(n210));
Q_MX02 U918 ( .S(n7), .A0(n211), .A1(auth_tag[71]), .Z(nxt_auth_tag[71]));
Q_AN02 U919 ( .A0(n8), .A1(ciph_out[71]), .Z(n211));
Q_MX02 U920 ( .S(n7), .A0(n212), .A1(auth_tag[70]), .Z(nxt_auth_tag[70]));
Q_AN02 U921 ( .A0(n8), .A1(ciph_out[70]), .Z(n212));
Q_MX02 U922 ( .S(n7), .A0(n213), .A1(auth_tag[69]), .Z(nxt_auth_tag[69]));
Q_AN02 U923 ( .A0(n8), .A1(ciph_out[69]), .Z(n213));
Q_MX02 U924 ( .S(n7), .A0(n214), .A1(auth_tag[68]), .Z(nxt_auth_tag[68]));
Q_AN02 U925 ( .A0(n8), .A1(ciph_out[68]), .Z(n214));
Q_MX02 U926 ( .S(n7), .A0(n215), .A1(auth_tag[67]), .Z(nxt_auth_tag[67]));
Q_AN02 U927 ( .A0(n8), .A1(ciph_out[67]), .Z(n215));
Q_MX02 U928 ( .S(n7), .A0(n216), .A1(auth_tag[66]), .Z(nxt_auth_tag[66]));
Q_AN02 U929 ( .A0(n8), .A1(ciph_out[66]), .Z(n216));
Q_MX02 U930 ( .S(n7), .A0(n217), .A1(auth_tag[65]), .Z(nxt_auth_tag[65]));
Q_AN02 U931 ( .A0(n8), .A1(ciph_out[65]), .Z(n217));
Q_MX02 U932 ( .S(n7), .A0(n218), .A1(auth_tag[64]), .Z(nxt_auth_tag[64]));
Q_AN02 U933 ( .A0(n8), .A1(ciph_out[64]), .Z(n218));
Q_MX02 U934 ( .S(n7), .A0(n219), .A1(auth_tag[63]), .Z(nxt_auth_tag[63]));
Q_AN02 U935 ( .A0(n8), .A1(ciph_out[63]), .Z(n219));
Q_MX02 U936 ( .S(n7), .A0(n220), .A1(auth_tag[62]), .Z(nxt_auth_tag[62]));
Q_AN02 U937 ( .A0(n8), .A1(ciph_out[62]), .Z(n220));
Q_MX02 U938 ( .S(n7), .A0(n221), .A1(auth_tag[61]), .Z(nxt_auth_tag[61]));
Q_AN02 U939 ( .A0(n8), .A1(ciph_out[61]), .Z(n221));
Q_MX02 U940 ( .S(n7), .A0(n222), .A1(auth_tag[60]), .Z(nxt_auth_tag[60]));
Q_AN02 U941 ( .A0(n8), .A1(ciph_out[60]), .Z(n222));
Q_MX02 U942 ( .S(n7), .A0(n223), .A1(auth_tag[59]), .Z(nxt_auth_tag[59]));
Q_AN02 U943 ( .A0(n8), .A1(ciph_out[59]), .Z(n223));
Q_MX02 U944 ( .S(n7), .A0(n224), .A1(auth_tag[58]), .Z(nxt_auth_tag[58]));
Q_AN02 U945 ( .A0(n8), .A1(ciph_out[58]), .Z(n224));
Q_MX02 U946 ( .S(n7), .A0(n225), .A1(auth_tag[57]), .Z(nxt_auth_tag[57]));
Q_AN02 U947 ( .A0(n8), .A1(ciph_out[57]), .Z(n225));
Q_MX02 U948 ( .S(n7), .A0(n226), .A1(auth_tag[56]), .Z(nxt_auth_tag[56]));
Q_AN02 U949 ( .A0(n8), .A1(ciph_out[56]), .Z(n226));
Q_MX02 U950 ( .S(n7), .A0(n227), .A1(auth_tag[55]), .Z(nxt_auth_tag[55]));
Q_AN02 U951 ( .A0(n8), .A1(ciph_out[55]), .Z(n227));
Q_MX02 U952 ( .S(n7), .A0(n228), .A1(auth_tag[54]), .Z(nxt_auth_tag[54]));
Q_AN02 U953 ( .A0(n8), .A1(ciph_out[54]), .Z(n228));
Q_MX02 U954 ( .S(n7), .A0(n229), .A1(auth_tag[53]), .Z(nxt_auth_tag[53]));
Q_AN02 U955 ( .A0(n8), .A1(ciph_out[53]), .Z(n229));
Q_MX02 U956 ( .S(n7), .A0(n230), .A1(auth_tag[52]), .Z(nxt_auth_tag[52]));
Q_AN02 U957 ( .A0(n8), .A1(ciph_out[52]), .Z(n230));
Q_MX02 U958 ( .S(n7), .A0(n231), .A1(auth_tag[51]), .Z(nxt_auth_tag[51]));
Q_AN02 U959 ( .A0(n8), .A1(ciph_out[51]), .Z(n231));
Q_MX02 U960 ( .S(n7), .A0(n232), .A1(auth_tag[50]), .Z(nxt_auth_tag[50]));
Q_AN02 U961 ( .A0(n8), .A1(ciph_out[50]), .Z(n232));
Q_MX02 U962 ( .S(n7), .A0(n233), .A1(auth_tag[49]), .Z(nxt_auth_tag[49]));
Q_AN02 U963 ( .A0(n8), .A1(ciph_out[49]), .Z(n233));
Q_MX02 U964 ( .S(n7), .A0(n234), .A1(auth_tag[48]), .Z(nxt_auth_tag[48]));
Q_AN02 U965 ( .A0(n8), .A1(ciph_out[48]), .Z(n234));
Q_MX02 U966 ( .S(n7), .A0(n235), .A1(auth_tag[47]), .Z(nxt_auth_tag[47]));
Q_AN02 U967 ( .A0(n8), .A1(ciph_out[47]), .Z(n235));
Q_MX02 U968 ( .S(n7), .A0(n236), .A1(auth_tag[46]), .Z(nxt_auth_tag[46]));
Q_AN02 U969 ( .A0(n8), .A1(ciph_out[46]), .Z(n236));
Q_MX02 U970 ( .S(n7), .A0(n237), .A1(auth_tag[45]), .Z(nxt_auth_tag[45]));
Q_AN02 U971 ( .A0(n8), .A1(ciph_out[45]), .Z(n237));
Q_MX02 U972 ( .S(n7), .A0(n238), .A1(auth_tag[44]), .Z(nxt_auth_tag[44]));
Q_AN02 U973 ( .A0(n8), .A1(ciph_out[44]), .Z(n238));
Q_MX02 U974 ( .S(n7), .A0(n239), .A1(auth_tag[43]), .Z(nxt_auth_tag[43]));
Q_AN02 U975 ( .A0(n8), .A1(ciph_out[43]), .Z(n239));
Q_MX02 U976 ( .S(n7), .A0(n240), .A1(auth_tag[42]), .Z(nxt_auth_tag[42]));
Q_AN02 U977 ( .A0(n8), .A1(ciph_out[42]), .Z(n240));
Q_MX02 U978 ( .S(n7), .A0(n241), .A1(auth_tag[41]), .Z(nxt_auth_tag[41]));
Q_AN02 U979 ( .A0(n8), .A1(ciph_out[41]), .Z(n241));
Q_MX02 U980 ( .S(n7), .A0(n242), .A1(auth_tag[40]), .Z(nxt_auth_tag[40]));
Q_AN02 U981 ( .A0(n8), .A1(ciph_out[40]), .Z(n242));
Q_MX02 U982 ( .S(n7), .A0(n243), .A1(auth_tag[39]), .Z(nxt_auth_tag[39]));
Q_AN02 U983 ( .A0(n8), .A1(ciph_out[39]), .Z(n243));
Q_MX02 U984 ( .S(n7), .A0(n244), .A1(auth_tag[38]), .Z(nxt_auth_tag[38]));
Q_AN02 U985 ( .A0(n8), .A1(ciph_out[38]), .Z(n244));
Q_MX02 U986 ( .S(n7), .A0(n245), .A1(auth_tag[37]), .Z(nxt_auth_tag[37]));
Q_AN02 U987 ( .A0(n8), .A1(ciph_out[37]), .Z(n245));
Q_MX02 U988 ( .S(n7), .A0(n246), .A1(auth_tag[36]), .Z(nxt_auth_tag[36]));
Q_AN02 U989 ( .A0(n8), .A1(ciph_out[36]), .Z(n246));
Q_MX02 U990 ( .S(n7), .A0(n247), .A1(auth_tag[35]), .Z(nxt_auth_tag[35]));
Q_AN02 U991 ( .A0(n8), .A1(ciph_out[35]), .Z(n247));
Q_MX02 U992 ( .S(n7), .A0(n248), .A1(auth_tag[34]), .Z(nxt_auth_tag[34]));
Q_AN02 U993 ( .A0(n8), .A1(ciph_out[34]), .Z(n248));
Q_MX02 U994 ( .S(n7), .A0(n249), .A1(auth_tag[33]), .Z(nxt_auth_tag[33]));
Q_AN02 U995 ( .A0(n8), .A1(ciph_out[33]), .Z(n249));
Q_MX02 U996 ( .S(n7), .A0(n250), .A1(auth_tag[32]), .Z(nxt_auth_tag[32]));
Q_AN02 U997 ( .A0(n8), .A1(ciph_out[32]), .Z(n250));
Q_MX02 U998 ( .S(n7), .A0(n251), .A1(auth_tag[31]), .Z(nxt_auth_tag[31]));
Q_AN02 U999 ( .A0(n8), .A1(ciph_out[31]), .Z(n251));
Q_MX02 U1000 ( .S(n7), .A0(n252), .A1(auth_tag[30]), .Z(nxt_auth_tag[30]));
Q_AN02 U1001 ( .A0(n8), .A1(ciph_out[30]), .Z(n252));
Q_MX02 U1002 ( .S(n7), .A0(n253), .A1(auth_tag[29]), .Z(nxt_auth_tag[29]));
Q_AN02 U1003 ( .A0(n8), .A1(ciph_out[29]), .Z(n253));
Q_MX02 U1004 ( .S(n7), .A0(n254), .A1(auth_tag[28]), .Z(nxt_auth_tag[28]));
Q_AN02 U1005 ( .A0(n8), .A1(ciph_out[28]), .Z(n254));
Q_MX02 U1006 ( .S(n7), .A0(n255), .A1(auth_tag[27]), .Z(nxt_auth_tag[27]));
Q_AN02 U1007 ( .A0(n8), .A1(ciph_out[27]), .Z(n255));
Q_MX02 U1008 ( .S(n7), .A0(n256), .A1(auth_tag[26]), .Z(nxt_auth_tag[26]));
Q_AN02 U1009 ( .A0(n8), .A1(ciph_out[26]), .Z(n256));
Q_MX02 U1010 ( .S(n7), .A0(n257), .A1(auth_tag[25]), .Z(nxt_auth_tag[25]));
Q_AN02 U1011 ( .A0(n8), .A1(ciph_out[25]), .Z(n257));
Q_MX02 U1012 ( .S(n7), .A0(n258), .A1(auth_tag[24]), .Z(nxt_auth_tag[24]));
Q_AN02 U1013 ( .A0(n8), .A1(ciph_out[24]), .Z(n258));
Q_MX02 U1014 ( .S(n7), .A0(n259), .A1(auth_tag[23]), .Z(nxt_auth_tag[23]));
Q_AN02 U1015 ( .A0(n8), .A1(ciph_out[23]), .Z(n259));
Q_MX02 U1016 ( .S(n7), .A0(n260), .A1(auth_tag[22]), .Z(nxt_auth_tag[22]));
Q_AN02 U1017 ( .A0(n8), .A1(ciph_out[22]), .Z(n260));
Q_MX02 U1018 ( .S(n7), .A0(n261), .A1(auth_tag[21]), .Z(nxt_auth_tag[21]));
Q_AN02 U1019 ( .A0(n8), .A1(ciph_out[21]), .Z(n261));
Q_MX02 U1020 ( .S(n7), .A0(n262), .A1(auth_tag[20]), .Z(nxt_auth_tag[20]));
Q_AN02 U1021 ( .A0(n8), .A1(ciph_out[20]), .Z(n262));
Q_MX02 U1022 ( .S(n7), .A0(n263), .A1(auth_tag[19]), .Z(nxt_auth_tag[19]));
Q_AN02 U1023 ( .A0(n8), .A1(ciph_out[19]), .Z(n263));
Q_MX02 U1024 ( .S(n7), .A0(n264), .A1(auth_tag[18]), .Z(nxt_auth_tag[18]));
Q_AN02 U1025 ( .A0(n8), .A1(ciph_out[18]), .Z(n264));
Q_MX02 U1026 ( .S(n7), .A0(n265), .A1(auth_tag[17]), .Z(nxt_auth_tag[17]));
Q_AN02 U1027 ( .A0(n8), .A1(ciph_out[17]), .Z(n265));
Q_MX02 U1028 ( .S(n7), .A0(n266), .A1(auth_tag[16]), .Z(nxt_auth_tag[16]));
Q_AN02 U1029 ( .A0(n8), .A1(ciph_out[16]), .Z(n266));
Q_MX02 U1030 ( .S(n7), .A0(n267), .A1(auth_tag[15]), .Z(nxt_auth_tag[15]));
Q_AN02 U1031 ( .A0(n8), .A1(ciph_out[15]), .Z(n267));
Q_MX02 U1032 ( .S(n7), .A0(n268), .A1(auth_tag[14]), .Z(nxt_auth_tag[14]));
Q_AN02 U1033 ( .A0(n8), .A1(ciph_out[14]), .Z(n268));
Q_MX02 U1034 ( .S(n7), .A0(n269), .A1(auth_tag[13]), .Z(nxt_auth_tag[13]));
Q_AN02 U1035 ( .A0(n8), .A1(ciph_out[13]), .Z(n269));
Q_MX02 U1036 ( .S(n7), .A0(n270), .A1(auth_tag[12]), .Z(nxt_auth_tag[12]));
Q_AN02 U1037 ( .A0(n8), .A1(ciph_out[12]), .Z(n270));
Q_MX02 U1038 ( .S(n7), .A0(n271), .A1(auth_tag[11]), .Z(nxt_auth_tag[11]));
Q_AN02 U1039 ( .A0(n8), .A1(ciph_out[11]), .Z(n271));
Q_MX02 U1040 ( .S(n7), .A0(n272), .A1(auth_tag[10]), .Z(nxt_auth_tag[10]));
Q_AN02 U1041 ( .A0(n8), .A1(ciph_out[10]), .Z(n272));
Q_MX02 U1042 ( .S(n7), .A0(n273), .A1(auth_tag[9]), .Z(nxt_auth_tag[9]));
Q_AN02 U1043 ( .A0(n8), .A1(ciph_out[9]), .Z(n273));
Q_MX02 U1044 ( .S(n7), .A0(n274), .A1(auth_tag[8]), .Z(nxt_auth_tag[8]));
Q_AN02 U1045 ( .A0(n8), .A1(ciph_out[8]), .Z(n274));
Q_MX02 U1046 ( .S(n7), .A0(n275), .A1(auth_tag[7]), .Z(nxt_auth_tag[7]));
Q_AN02 U1047 ( .A0(n8), .A1(ciph_out[7]), .Z(n275));
Q_MX02 U1048 ( .S(n7), .A0(n276), .A1(auth_tag[6]), .Z(nxt_auth_tag[6]));
Q_AN02 U1049 ( .A0(n8), .A1(ciph_out[6]), .Z(n276));
Q_MX02 U1050 ( .S(n7), .A0(n277), .A1(auth_tag[5]), .Z(nxt_auth_tag[5]));
Q_AN02 U1051 ( .A0(n8), .A1(ciph_out[5]), .Z(n277));
Q_MX02 U1052 ( .S(n7), .A0(n278), .A1(auth_tag[4]), .Z(nxt_auth_tag[4]));
Q_AN02 U1053 ( .A0(n8), .A1(ciph_out[4]), .Z(n278));
Q_MX02 U1054 ( .S(n7), .A0(n279), .A1(auth_tag[3]), .Z(nxt_auth_tag[3]));
Q_AN02 U1055 ( .A0(n8), .A1(ciph_out[3]), .Z(n279));
Q_MX02 U1056 ( .S(n7), .A0(n280), .A1(auth_tag[2]), .Z(nxt_auth_tag[2]));
Q_AN02 U1057 ( .A0(n8), .A1(ciph_out[2]), .Z(n280));
Q_MX02 U1058 ( .S(n7), .A0(n281), .A1(auth_tag[1]), .Z(nxt_auth_tag[1]));
Q_AN02 U1059 ( .A0(n8), .A1(ciph_out[1]), .Z(n281));
Q_MX02 U1060 ( .S(n7), .A0(n282), .A1(auth_tag[0]), .Z(nxt_auth_tag[0]));
Q_AN02 U1061 ( .A0(n8), .A1(ciph_out[0]), .Z(n282));
Q_XOR2 U1062 ( .A0(fifo_out[128]), .A1(auth_tag[127]), .Z(n283));
Q_XOR2 U1063 ( .A0(fifo_out[127]), .A1(auth_tag[126]), .Z(n284));
Q_XOR2 U1064 ( .A0(fifo_out[126]), .A1(auth_tag[125]), .Z(n285));
Q_XOR2 U1065 ( .A0(fifo_out[125]), .A1(auth_tag[124]), .Z(n286));
Q_XOR2 U1066 ( .A0(fifo_out[124]), .A1(auth_tag[123]), .Z(n287));
Q_XOR2 U1067 ( .A0(fifo_out[123]), .A1(auth_tag[122]), .Z(n288));
Q_XOR2 U1068 ( .A0(fifo_out[122]), .A1(auth_tag[121]), .Z(n289));
Q_XOR2 U1069 ( .A0(fifo_out[121]), .A1(auth_tag[120]), .Z(n290));
Q_XOR2 U1070 ( .A0(fifo_out[120]), .A1(auth_tag[119]), .Z(n291));
Q_XOR2 U1071 ( .A0(fifo_out[119]), .A1(auth_tag[118]), .Z(n292));
Q_XOR2 U1072 ( .A0(fifo_out[118]), .A1(auth_tag[117]), .Z(n293));
Q_XOR2 U1073 ( .A0(fifo_out[117]), .A1(auth_tag[116]), .Z(n294));
Q_XOR2 U1074 ( .A0(fifo_out[116]), .A1(auth_tag[115]), .Z(n295));
Q_XOR2 U1075 ( .A0(fifo_out[115]), .A1(auth_tag[114]), .Z(n296));
Q_XOR2 U1076 ( .A0(fifo_out[114]), .A1(auth_tag[113]), .Z(n297));
Q_XOR2 U1077 ( .A0(fifo_out[113]), .A1(auth_tag[112]), .Z(n298));
Q_XOR2 U1078 ( .A0(fifo_out[112]), .A1(auth_tag[111]), .Z(n299));
Q_XOR2 U1079 ( .A0(fifo_out[111]), .A1(auth_tag[110]), .Z(n300));
Q_XOR2 U1080 ( .A0(fifo_out[110]), .A1(auth_tag[109]), .Z(n301));
Q_XOR2 U1081 ( .A0(fifo_out[109]), .A1(auth_tag[108]), .Z(n302));
Q_XOR2 U1082 ( .A0(fifo_out[108]), .A1(auth_tag[107]), .Z(n303));
Q_XOR2 U1083 ( .A0(fifo_out[107]), .A1(auth_tag[106]), .Z(n304));
Q_XOR2 U1084 ( .A0(fifo_out[106]), .A1(auth_tag[105]), .Z(n305));
Q_XOR2 U1085 ( .A0(fifo_out[105]), .A1(auth_tag[104]), .Z(n306));
Q_XOR2 U1086 ( .A0(fifo_out[104]), .A1(auth_tag[103]), .Z(n307));
Q_XOR2 U1087 ( .A0(fifo_out[103]), .A1(auth_tag[102]), .Z(n308));
Q_XOR2 U1088 ( .A0(fifo_out[102]), .A1(auth_tag[101]), .Z(n309));
Q_XOR2 U1089 ( .A0(fifo_out[101]), .A1(auth_tag[100]), .Z(n310));
Q_XOR2 U1090 ( .A0(fifo_out[100]), .A1(auth_tag[99]), .Z(n311));
Q_XOR2 U1091 ( .A0(fifo_out[99]), .A1(auth_tag[98]), .Z(n312));
Q_XOR2 U1092 ( .A0(fifo_out[98]), .A1(auth_tag[97]), .Z(n313));
Q_XOR2 U1093 ( .A0(fifo_out[97]), .A1(auth_tag[96]), .Z(n314));
Q_XOR2 U1094 ( .A0(fifo_out[96]), .A1(auth_tag[95]), .Z(n315));
Q_XOR2 U1095 ( .A0(fifo_out[95]), .A1(auth_tag[94]), .Z(n316));
Q_XOR2 U1096 ( .A0(fifo_out[94]), .A1(auth_tag[93]), .Z(n317));
Q_XOR2 U1097 ( .A0(fifo_out[93]), .A1(auth_tag[92]), .Z(n318));
Q_XOR2 U1098 ( .A0(fifo_out[92]), .A1(auth_tag[91]), .Z(n319));
Q_XOR2 U1099 ( .A0(fifo_out[91]), .A1(auth_tag[90]), .Z(n320));
Q_XOR2 U1100 ( .A0(fifo_out[90]), .A1(auth_tag[89]), .Z(n321));
Q_XOR2 U1101 ( .A0(fifo_out[89]), .A1(auth_tag[88]), .Z(n322));
Q_XOR2 U1102 ( .A0(fifo_out[88]), .A1(auth_tag[87]), .Z(n323));
Q_XOR2 U1103 ( .A0(fifo_out[87]), .A1(auth_tag[86]), .Z(n324));
Q_XOR2 U1104 ( .A0(fifo_out[86]), .A1(auth_tag[85]), .Z(n325));
Q_XOR2 U1105 ( .A0(fifo_out[85]), .A1(auth_tag[84]), .Z(n326));
Q_XOR2 U1106 ( .A0(fifo_out[84]), .A1(auth_tag[83]), .Z(n327));
Q_XOR2 U1107 ( .A0(fifo_out[83]), .A1(auth_tag[82]), .Z(n328));
Q_XOR2 U1108 ( .A0(fifo_out[82]), .A1(auth_tag[81]), .Z(n329));
Q_XOR2 U1109 ( .A0(fifo_out[81]), .A1(auth_tag[80]), .Z(n330));
Q_XOR2 U1110 ( .A0(fifo_out[80]), .A1(auth_tag[79]), .Z(n331));
Q_XOR2 U1111 ( .A0(fifo_out[79]), .A1(auth_tag[78]), .Z(n332));
Q_XOR2 U1112 ( .A0(fifo_out[78]), .A1(auth_tag[77]), .Z(n333));
Q_XOR2 U1113 ( .A0(fifo_out[77]), .A1(auth_tag[76]), .Z(n334));
Q_XOR2 U1114 ( .A0(fifo_out[76]), .A1(auth_tag[75]), .Z(n335));
Q_XOR2 U1115 ( .A0(fifo_out[75]), .A1(auth_tag[74]), .Z(n336));
Q_XOR2 U1116 ( .A0(fifo_out[74]), .A1(auth_tag[73]), .Z(n337));
Q_XOR2 U1117 ( .A0(fifo_out[73]), .A1(auth_tag[72]), .Z(n338));
Q_XOR2 U1118 ( .A0(fifo_out[72]), .A1(auth_tag[71]), .Z(n339));
Q_XOR2 U1119 ( .A0(fifo_out[71]), .A1(auth_tag[70]), .Z(n340));
Q_XOR2 U1120 ( .A0(fifo_out[70]), .A1(auth_tag[69]), .Z(n341));
Q_XOR2 U1121 ( .A0(fifo_out[69]), .A1(auth_tag[68]), .Z(n342));
Q_XOR2 U1122 ( .A0(fifo_out[68]), .A1(auth_tag[67]), .Z(n343));
Q_XOR2 U1123 ( .A0(fifo_out[67]), .A1(auth_tag[66]), .Z(n344));
Q_XOR2 U1124 ( .A0(fifo_out[66]), .A1(auth_tag[65]), .Z(n345));
Q_XOR2 U1125 ( .A0(fifo_out[65]), .A1(auth_tag[64]), .Z(n346));
Q_XOR2 U1126 ( .A0(fifo_out[64]), .A1(auth_tag[63]), .Z(n347));
Q_XOR2 U1127 ( .A0(fifo_out[63]), .A1(auth_tag[62]), .Z(n348));
Q_XOR2 U1128 ( .A0(fifo_out[62]), .A1(auth_tag[61]), .Z(n349));
Q_XOR2 U1129 ( .A0(fifo_out[61]), .A1(auth_tag[60]), .Z(n350));
Q_XOR2 U1130 ( .A0(fifo_out[60]), .A1(auth_tag[59]), .Z(n351));
Q_XOR2 U1131 ( .A0(fifo_out[59]), .A1(auth_tag[58]), .Z(n352));
Q_XOR2 U1132 ( .A0(fifo_out[58]), .A1(auth_tag[57]), .Z(n353));
Q_XOR2 U1133 ( .A0(fifo_out[57]), .A1(auth_tag[56]), .Z(n354));
Q_XOR2 U1134 ( .A0(fifo_out[56]), .A1(auth_tag[55]), .Z(n355));
Q_XOR2 U1135 ( .A0(fifo_out[55]), .A1(auth_tag[54]), .Z(n356));
Q_XOR2 U1136 ( .A0(fifo_out[54]), .A1(auth_tag[53]), .Z(n357));
Q_XOR2 U1137 ( .A0(fifo_out[53]), .A1(auth_tag[52]), .Z(n358));
Q_XOR2 U1138 ( .A0(fifo_out[52]), .A1(auth_tag[51]), .Z(n359));
Q_XOR2 U1139 ( .A0(fifo_out[51]), .A1(auth_tag[50]), .Z(n360));
Q_XOR2 U1140 ( .A0(fifo_out[50]), .A1(auth_tag[49]), .Z(n361));
Q_XOR2 U1141 ( .A0(fifo_out[49]), .A1(auth_tag[48]), .Z(n362));
Q_XOR2 U1142 ( .A0(fifo_out[48]), .A1(auth_tag[47]), .Z(n363));
Q_XOR2 U1143 ( .A0(fifo_out[47]), .A1(auth_tag[46]), .Z(n364));
Q_XOR2 U1144 ( .A0(fifo_out[46]), .A1(auth_tag[45]), .Z(n365));
Q_XOR2 U1145 ( .A0(fifo_out[45]), .A1(auth_tag[44]), .Z(n366));
Q_XOR2 U1146 ( .A0(fifo_out[44]), .A1(auth_tag[43]), .Z(n367));
Q_XOR2 U1147 ( .A0(fifo_out[43]), .A1(auth_tag[42]), .Z(n368));
Q_XOR2 U1148 ( .A0(fifo_out[42]), .A1(auth_tag[41]), .Z(n369));
Q_XOR2 U1149 ( .A0(fifo_out[41]), .A1(auth_tag[40]), .Z(n370));
Q_XOR2 U1150 ( .A0(fifo_out[40]), .A1(auth_tag[39]), .Z(n371));
Q_XOR2 U1151 ( .A0(fifo_out[39]), .A1(auth_tag[38]), .Z(n372));
Q_XOR2 U1152 ( .A0(fifo_out[38]), .A1(auth_tag[37]), .Z(n373));
Q_XOR2 U1153 ( .A0(fifo_out[37]), .A1(auth_tag[36]), .Z(n374));
Q_XOR2 U1154 ( .A0(fifo_out[36]), .A1(auth_tag[35]), .Z(n375));
Q_XOR2 U1155 ( .A0(fifo_out[35]), .A1(auth_tag[34]), .Z(n376));
Q_XOR2 U1156 ( .A0(fifo_out[34]), .A1(auth_tag[33]), .Z(n377));
Q_XOR2 U1157 ( .A0(fifo_out[33]), .A1(auth_tag[32]), .Z(n378));
Q_XOR2 U1158 ( .A0(fifo_out[32]), .A1(auth_tag[31]), .Z(n379));
Q_XOR2 U1159 ( .A0(fifo_out[31]), .A1(auth_tag[30]), .Z(n380));
Q_XOR2 U1160 ( .A0(fifo_out[30]), .A1(auth_tag[29]), .Z(n381));
Q_XOR2 U1161 ( .A0(fifo_out[29]), .A1(auth_tag[28]), .Z(n382));
Q_XOR2 U1162 ( .A0(fifo_out[28]), .A1(auth_tag[27]), .Z(n383));
Q_XOR2 U1163 ( .A0(fifo_out[27]), .A1(auth_tag[26]), .Z(n384));
Q_XOR2 U1164 ( .A0(fifo_out[26]), .A1(auth_tag[25]), .Z(n385));
Q_XOR2 U1165 ( .A0(fifo_out[25]), .A1(auth_tag[24]), .Z(n386));
Q_XOR2 U1166 ( .A0(fifo_out[24]), .A1(auth_tag[23]), .Z(n387));
Q_XOR2 U1167 ( .A0(fifo_out[23]), .A1(auth_tag[22]), .Z(n388));
Q_XOR2 U1168 ( .A0(fifo_out[22]), .A1(auth_tag[21]), .Z(n389));
Q_XOR2 U1169 ( .A0(fifo_out[21]), .A1(auth_tag[20]), .Z(n390));
Q_XOR2 U1170 ( .A0(fifo_out[20]), .A1(auth_tag[19]), .Z(n391));
Q_XOR2 U1171 ( .A0(fifo_out[19]), .A1(auth_tag[18]), .Z(n392));
Q_XOR2 U1172 ( .A0(fifo_out[18]), .A1(auth_tag[17]), .Z(n393));
Q_XOR2 U1173 ( .A0(fifo_out[17]), .A1(auth_tag[16]), .Z(n394));
Q_XOR2 U1174 ( .A0(fifo_out[16]), .A1(auth_tag[15]), .Z(n395));
Q_XOR2 U1175 ( .A0(fifo_out[15]), .A1(auth_tag[14]), .Z(n396));
Q_XOR2 U1176 ( .A0(fifo_out[14]), .A1(auth_tag[13]), .Z(n397));
Q_XOR2 U1177 ( .A0(fifo_out[13]), .A1(auth_tag[12]), .Z(n398));
Q_XOR2 U1178 ( .A0(fifo_out[12]), .A1(auth_tag[11]), .Z(n399));
Q_XOR2 U1179 ( .A0(fifo_out[11]), .A1(auth_tag[10]), .Z(n400));
Q_XOR2 U1180 ( .A0(fifo_out[10]), .A1(auth_tag[9]), .Z(n401));
Q_XOR2 U1181 ( .A0(fifo_out[9]), .A1(auth_tag[8]), .Z(n402));
Q_XOR2 U1182 ( .A0(fifo_out[8]), .A1(auth_tag[7]), .Z(n403));
Q_XOR2 U1183 ( .A0(fifo_out[7]), .A1(auth_tag[6]), .Z(n404));
Q_XOR2 U1184 ( .A0(fifo_out[6]), .A1(auth_tag[5]), .Z(n405));
Q_XOR2 U1185 ( .A0(fifo_out[5]), .A1(auth_tag[4]), .Z(n406));
Q_XOR2 U1186 ( .A0(fifo_out[4]), .A1(auth_tag[3]), .Z(n407));
Q_XOR2 U1187 ( .A0(fifo_out[3]), .A1(auth_tag[2]), .Z(n408));
Q_XOR2 U1188 ( .A0(fifo_out[2]), .A1(auth_tag[1]), .Z(n409));
Q_XOR2 U1189 ( .A0(fifo_out[1]), .A1(auth_tag[0]), .Z(n410));
Q_XOR2 U1190 ( .A0(fifo_out[128]), .A1(ciph_out[127]), .Z(n411));
Q_XOR2 U1191 ( .A0(fifo_out[127]), .A1(ciph_out[126]), .Z(n412));
Q_XOR2 U1192 ( .A0(fifo_out[126]), .A1(ciph_out[125]), .Z(n413));
Q_XOR2 U1193 ( .A0(fifo_out[125]), .A1(ciph_out[124]), .Z(n414));
Q_XOR2 U1194 ( .A0(fifo_out[124]), .A1(ciph_out[123]), .Z(n415));
Q_XOR2 U1195 ( .A0(fifo_out[123]), .A1(ciph_out[122]), .Z(n416));
Q_XOR2 U1196 ( .A0(fifo_out[122]), .A1(ciph_out[121]), .Z(n417));
Q_XOR2 U1197 ( .A0(fifo_out[121]), .A1(ciph_out[120]), .Z(n418));
Q_XOR2 U1198 ( .A0(fifo_out[120]), .A1(ciph_out[119]), .Z(n419));
Q_XOR2 U1199 ( .A0(fifo_out[119]), .A1(ciph_out[118]), .Z(n420));
Q_XOR2 U1200 ( .A0(fifo_out[118]), .A1(ciph_out[117]), .Z(n421));
Q_XOR2 U1201 ( .A0(fifo_out[117]), .A1(ciph_out[116]), .Z(n422));
Q_XOR2 U1202 ( .A0(fifo_out[116]), .A1(ciph_out[115]), .Z(n423));
Q_XOR2 U1203 ( .A0(fifo_out[115]), .A1(ciph_out[114]), .Z(n424));
Q_XOR2 U1204 ( .A0(fifo_out[114]), .A1(ciph_out[113]), .Z(n425));
Q_XOR2 U1205 ( .A0(fifo_out[113]), .A1(ciph_out[112]), .Z(n426));
Q_XOR2 U1206 ( .A0(fifo_out[112]), .A1(ciph_out[111]), .Z(n427));
Q_XOR2 U1207 ( .A0(fifo_out[111]), .A1(ciph_out[110]), .Z(n428));
Q_XOR2 U1208 ( .A0(fifo_out[110]), .A1(ciph_out[109]), .Z(n429));
Q_XOR2 U1209 ( .A0(fifo_out[109]), .A1(ciph_out[108]), .Z(n430));
Q_XOR2 U1210 ( .A0(fifo_out[108]), .A1(ciph_out[107]), .Z(n431));
Q_XOR2 U1211 ( .A0(fifo_out[107]), .A1(ciph_out[106]), .Z(n432));
Q_XOR2 U1212 ( .A0(fifo_out[106]), .A1(ciph_out[105]), .Z(n433));
Q_XOR2 U1213 ( .A0(fifo_out[105]), .A1(ciph_out[104]), .Z(n434));
Q_XOR2 U1214 ( .A0(fifo_out[104]), .A1(ciph_out[103]), .Z(n435));
Q_XOR2 U1215 ( .A0(fifo_out[103]), .A1(ciph_out[102]), .Z(n436));
Q_XOR2 U1216 ( .A0(fifo_out[102]), .A1(ciph_out[101]), .Z(n437));
Q_XOR2 U1217 ( .A0(fifo_out[101]), .A1(ciph_out[100]), .Z(n438));
Q_XOR2 U1218 ( .A0(fifo_out[100]), .A1(ciph_out[99]), .Z(n439));
Q_XOR2 U1219 ( .A0(fifo_out[99]), .A1(ciph_out[98]), .Z(n440));
Q_XOR2 U1220 ( .A0(fifo_out[98]), .A1(ciph_out[97]), .Z(n441));
Q_XOR2 U1221 ( .A0(fifo_out[97]), .A1(ciph_out[96]), .Z(n442));
Q_XOR2 U1222 ( .A0(fifo_out[96]), .A1(ciph_out[95]), .Z(n443));
Q_XOR2 U1223 ( .A0(fifo_out[95]), .A1(ciph_out[94]), .Z(n444));
Q_XOR2 U1224 ( .A0(fifo_out[94]), .A1(ciph_out[93]), .Z(n445));
Q_XOR2 U1225 ( .A0(fifo_out[93]), .A1(ciph_out[92]), .Z(n446));
Q_XOR2 U1226 ( .A0(fifo_out[92]), .A1(ciph_out[91]), .Z(n447));
Q_XOR2 U1227 ( .A0(fifo_out[91]), .A1(ciph_out[90]), .Z(n448));
Q_XOR2 U1228 ( .A0(fifo_out[90]), .A1(ciph_out[89]), .Z(n449));
Q_XOR2 U1229 ( .A0(fifo_out[89]), .A1(ciph_out[88]), .Z(n450));
Q_XOR2 U1230 ( .A0(fifo_out[88]), .A1(ciph_out[87]), .Z(n451));
Q_XOR2 U1231 ( .A0(fifo_out[87]), .A1(ciph_out[86]), .Z(n452));
Q_XOR2 U1232 ( .A0(fifo_out[86]), .A1(ciph_out[85]), .Z(n453));
Q_XOR2 U1233 ( .A0(fifo_out[85]), .A1(ciph_out[84]), .Z(n454));
Q_XOR2 U1234 ( .A0(fifo_out[84]), .A1(ciph_out[83]), .Z(n455));
Q_XOR2 U1235 ( .A0(fifo_out[83]), .A1(ciph_out[82]), .Z(n456));
Q_XOR2 U1236 ( .A0(fifo_out[82]), .A1(ciph_out[81]), .Z(n457));
Q_XOR2 U1237 ( .A0(fifo_out[81]), .A1(ciph_out[80]), .Z(n458));
Q_XOR2 U1238 ( .A0(fifo_out[80]), .A1(ciph_out[79]), .Z(n459));
Q_XOR2 U1239 ( .A0(fifo_out[79]), .A1(ciph_out[78]), .Z(n460));
Q_XOR2 U1240 ( .A0(fifo_out[78]), .A1(ciph_out[77]), .Z(n461));
Q_XOR2 U1241 ( .A0(fifo_out[77]), .A1(ciph_out[76]), .Z(n462));
Q_XOR2 U1242 ( .A0(fifo_out[76]), .A1(ciph_out[75]), .Z(n463));
Q_XOR2 U1243 ( .A0(fifo_out[75]), .A1(ciph_out[74]), .Z(n464));
Q_XOR2 U1244 ( .A0(fifo_out[74]), .A1(ciph_out[73]), .Z(n465));
Q_XOR2 U1245 ( .A0(fifo_out[73]), .A1(ciph_out[72]), .Z(n466));
Q_XOR2 U1246 ( .A0(fifo_out[72]), .A1(ciph_out[71]), .Z(n467));
Q_XOR2 U1247 ( .A0(fifo_out[71]), .A1(ciph_out[70]), .Z(n468));
Q_XOR2 U1248 ( .A0(fifo_out[70]), .A1(ciph_out[69]), .Z(n469));
Q_XOR2 U1249 ( .A0(fifo_out[69]), .A1(ciph_out[68]), .Z(n470));
Q_XOR2 U1250 ( .A0(fifo_out[68]), .A1(ciph_out[67]), .Z(n471));
Q_XOR2 U1251 ( .A0(fifo_out[67]), .A1(ciph_out[66]), .Z(n472));
Q_XOR2 U1252 ( .A0(fifo_out[66]), .A1(ciph_out[65]), .Z(n473));
Q_XOR2 U1253 ( .A0(fifo_out[65]), .A1(ciph_out[64]), .Z(n474));
Q_XOR2 U1254 ( .A0(fifo_out[64]), .A1(ciph_out[63]), .Z(n475));
Q_XOR2 U1255 ( .A0(fifo_out[63]), .A1(ciph_out[62]), .Z(n476));
Q_XOR2 U1256 ( .A0(fifo_out[62]), .A1(ciph_out[61]), .Z(n477));
Q_XOR2 U1257 ( .A0(fifo_out[61]), .A1(ciph_out[60]), .Z(n478));
Q_XOR2 U1258 ( .A0(fifo_out[60]), .A1(ciph_out[59]), .Z(n479));
Q_XOR2 U1259 ( .A0(fifo_out[59]), .A1(ciph_out[58]), .Z(n480));
Q_XOR2 U1260 ( .A0(fifo_out[58]), .A1(ciph_out[57]), .Z(n481));
Q_XOR2 U1261 ( .A0(fifo_out[57]), .A1(ciph_out[56]), .Z(n482));
Q_XOR2 U1262 ( .A0(fifo_out[56]), .A1(ciph_out[55]), .Z(n483));
Q_XOR2 U1263 ( .A0(fifo_out[55]), .A1(ciph_out[54]), .Z(n484));
Q_XOR2 U1264 ( .A0(fifo_out[54]), .A1(ciph_out[53]), .Z(n485));
Q_XOR2 U1265 ( .A0(fifo_out[53]), .A1(ciph_out[52]), .Z(n486));
Q_XOR2 U1266 ( .A0(fifo_out[52]), .A1(ciph_out[51]), .Z(n487));
Q_XOR2 U1267 ( .A0(fifo_out[51]), .A1(ciph_out[50]), .Z(n488));
Q_XOR2 U1268 ( .A0(fifo_out[50]), .A1(ciph_out[49]), .Z(n489));
Q_XOR2 U1269 ( .A0(fifo_out[49]), .A1(ciph_out[48]), .Z(n490));
Q_XOR2 U1270 ( .A0(fifo_out[48]), .A1(ciph_out[47]), .Z(n491));
Q_XOR2 U1271 ( .A0(fifo_out[47]), .A1(ciph_out[46]), .Z(n492));
Q_XOR2 U1272 ( .A0(fifo_out[46]), .A1(ciph_out[45]), .Z(n493));
Q_XOR2 U1273 ( .A0(fifo_out[45]), .A1(ciph_out[44]), .Z(n494));
Q_XOR2 U1274 ( .A0(fifo_out[44]), .A1(ciph_out[43]), .Z(n495));
Q_XOR2 U1275 ( .A0(fifo_out[43]), .A1(ciph_out[42]), .Z(n496));
Q_XOR2 U1276 ( .A0(fifo_out[42]), .A1(ciph_out[41]), .Z(n497));
Q_XOR2 U1277 ( .A0(fifo_out[41]), .A1(ciph_out[40]), .Z(n498));
Q_XOR2 U1278 ( .A0(fifo_out[40]), .A1(ciph_out[39]), .Z(n499));
Q_XOR2 U1279 ( .A0(fifo_out[39]), .A1(ciph_out[38]), .Z(n500));
Q_XOR2 U1280 ( .A0(fifo_out[38]), .A1(ciph_out[37]), .Z(n501));
Q_XOR2 U1281 ( .A0(fifo_out[37]), .A1(ciph_out[36]), .Z(n502));
Q_XOR2 U1282 ( .A0(fifo_out[36]), .A1(ciph_out[35]), .Z(n503));
Q_XOR2 U1283 ( .A0(fifo_out[35]), .A1(ciph_out[34]), .Z(n504));
Q_XOR2 U1284 ( .A0(fifo_out[34]), .A1(ciph_out[33]), .Z(n505));
Q_XOR2 U1285 ( .A0(fifo_out[33]), .A1(ciph_out[32]), .Z(n506));
Q_XOR2 U1286 ( .A0(fifo_out[32]), .A1(ciph_out[31]), .Z(n507));
Q_XOR2 U1287 ( .A0(fifo_out[31]), .A1(ciph_out[30]), .Z(n508));
Q_XOR2 U1288 ( .A0(fifo_out[30]), .A1(ciph_out[29]), .Z(n509));
Q_XOR2 U1289 ( .A0(fifo_out[29]), .A1(ciph_out[28]), .Z(n510));
Q_XOR2 U1290 ( .A0(fifo_out[28]), .A1(ciph_out[27]), .Z(n511));
Q_XOR2 U1291 ( .A0(fifo_out[27]), .A1(ciph_out[26]), .Z(n512));
Q_XOR2 U1292 ( .A0(fifo_out[26]), .A1(ciph_out[25]), .Z(n513));
Q_XOR2 U1293 ( .A0(fifo_out[25]), .A1(ciph_out[24]), .Z(n514));
Q_XOR2 U1294 ( .A0(fifo_out[24]), .A1(ciph_out[23]), .Z(n515));
Q_XOR2 U1295 ( .A0(fifo_out[23]), .A1(ciph_out[22]), .Z(n516));
Q_XOR2 U1296 ( .A0(fifo_out[22]), .A1(ciph_out[21]), .Z(n517));
Q_XOR2 U1297 ( .A0(fifo_out[21]), .A1(ciph_out[20]), .Z(n518));
Q_XOR2 U1298 ( .A0(fifo_out[20]), .A1(ciph_out[19]), .Z(n519));
Q_XOR2 U1299 ( .A0(fifo_out[19]), .A1(ciph_out[18]), .Z(n520));
Q_XOR2 U1300 ( .A0(fifo_out[18]), .A1(ciph_out[17]), .Z(n521));
Q_XOR2 U1301 ( .A0(fifo_out[17]), .A1(ciph_out[16]), .Z(n522));
Q_XOR2 U1302 ( .A0(fifo_out[16]), .A1(ciph_out[15]), .Z(n523));
Q_XOR2 U1303 ( .A0(fifo_out[15]), .A1(ciph_out[14]), .Z(n524));
Q_XOR2 U1304 ( .A0(fifo_out[14]), .A1(ciph_out[13]), .Z(n525));
Q_XOR2 U1305 ( .A0(fifo_out[13]), .A1(ciph_out[12]), .Z(n526));
Q_XOR2 U1306 ( .A0(fifo_out[12]), .A1(ciph_out[11]), .Z(n527));
Q_XOR2 U1307 ( .A0(fifo_out[11]), .A1(ciph_out[10]), .Z(n528));
Q_XOR2 U1308 ( .A0(fifo_out[10]), .A1(ciph_out[9]), .Z(n529));
Q_XOR2 U1309 ( .A0(fifo_out[9]), .A1(ciph_out[8]), .Z(n530));
Q_XOR2 U1310 ( .A0(fifo_out[8]), .A1(ciph_out[7]), .Z(n531));
Q_XOR2 U1311 ( .A0(fifo_out[7]), .A1(ciph_out[6]), .Z(n532));
Q_XOR2 U1312 ( .A0(fifo_out[6]), .A1(ciph_out[5]), .Z(n533));
Q_XOR2 U1313 ( .A0(fifo_out[5]), .A1(ciph_out[4]), .Z(n534));
Q_XOR2 U1314 ( .A0(fifo_out[4]), .A1(ciph_out[3]), .Z(n535));
Q_XOR2 U1315 ( .A0(fifo_out[3]), .A1(ciph_out[2]), .Z(n536));
Q_XOR2 U1316 ( .A0(fifo_out[2]), .A1(ciph_out[1]), .Z(n537));
Q_XOR2 U1317 ( .A0(fifo_out[1]), .A1(ciph_out[0]), .Z(n538));
Q_OR02 U1318 ( .A0(cmdfifo_gcm_cmd[1]), .A1(cmdfifo_gcm_cmd[2]), .Z(n580));
Q_ND02 U1319 ( .A0(upsizer_gcm_valid), .A1(n580), .Z(n552));
Q_OR02 U1320 ( .A0(n626), .A1(n552), .Z(n553));
Q_INV U1321 ( .A(cmdfifo_gcm_cmd[2]), .Z(n583));
Q_OA21 U1322 ( .A0(cmdfifo_gcm_cmd[1]), .A1(n583), .B0(cmdfifo_gcm_cmd[0]), .Z(n555));
Q_INV U1323 ( .A(cmdfifo_gcm_cmd[1]), .Z(n605));
Q_OA21 U1324 ( .A0(n605), .A1(cmdfifo_gcm_cmd[2]), .B0(n1224), .Z(n554));
Q_OR02 U1325 ( .A0(n555), .A1(n554), .Z(n624));
Q_INV U1326 ( .A(upsizer_gcm_valid), .Z(n620));
Q_OR03 U1327 ( .A0(n573), .A1(n624), .A2(n1237), .Z(n557));
Q_ND03 U1328 ( .A0(cur_state[0]), .A1(n540), .A2(cur_state[2]), .Z(n556));
Q_AN02 U1329 ( .A0(n557), .A1(n564), .Z(n558));
Q_INV U1330 ( .A(n558), .Z(n543));
Q_ND02 U1331 ( .A0(cur_state[2]), .A1(n540), .Z(n559));
Q_INV U1332 ( .A(n568), .Z(gcm_tag_data_out_ack));
Q_INV U1333 ( .A(n622), .Z(n549));
Q_OR02 U1334 ( .A0(n1243), .A1(ciph_fifo_in_stall), .Z(n618));
Q_NR02 U1335 ( .A0(n1649), .A1(n618), .Z(n560));
Q_AN02 U1336 ( .A0(ciph_fifo_in_stall), .A1(cur_state[0]), .Z(n566));
Q_NR02 U1337 ( .A0(upsizer_gcm_valid), .A1(cur_state[0]), .Z(n561));
Q_OR03 U1338 ( .A0(n566), .A1(n561), .A2(cur_state[2]), .Z(n570));
Q_OA21 U1339 ( .A0(n540), .A1(n1238), .B0(n1650), .Z(n562));
Q_INV U1340 ( .A(n562), .Z(n602));
Q_AN02 U1341 ( .A0(n571), .A1(n603), .Z(n563));
Q_INV U1342 ( .A(n563), .Z(fifo_in_vld));
Q_OR02 U1343 ( .A0(cur_state[1]), .A1(n556), .Z(n564));
Q_INV U1344 ( .A(n564), .Z(ciph_in_last));
Q_OR03 U1345 ( .A0(cur_state[0]), .A1(n541), .A2(cur_state[2]), .Z(n631));
Q_INV U1346 ( .A(n632), .Z(key_in_vld));
Q_OR03 U1347 ( .A0(n620), .A1(beat_num[1]), .A2(n624), .Z(n565));
Q_AO21 U1348 ( .A0(n565), .A1(n1243), .B0(n566), .Z(n567));
Q_OR03 U1349 ( .A0(cur_state[2]), .A1(n567), .A2(n1237), .Z(n569));
Q_OR02 U1350 ( .A0(n559), .A1(cur_state[1]), .Z(n568));
Q_AN02 U1351 ( .A0(n569), .A1(n568), .Z(n544));
Q_OR02 U1352 ( .A0(n1237), .A1(n570), .Z(n571));
Q_INV U1353 ( .A(n571), .Z(n545));
Q_MX02 U1354 ( .S(cmdfifo_gcm_cmd[0]), .A0(cmdfifo_gcm_cmd[2]), .A1(cmdfifo_gcm_cmd[1]), .Z(n628));
Q_MX02 U1355 ( .S(beat_num[1]), .A0(n628), .A1(n580), .Z(n572));
Q_OR02 U1356 ( .A0(cur_state[2]), .A1(n621), .Z(n573));
Q_OR02 U1357 ( .A0(n573), .A1(n572), .Z(n574));
Q_INV U1358 ( .A(n540), .Z(n616));
Q_OR03 U1359 ( .A0(n542), .A1(n616), .A2(n1243), .Z(n575));
Q_AN03 U1360 ( .A0(n575), .A1(n617), .A2(cur_state[2]), .Z(n577));
Q_AN02 U1361 ( .A0(n618), .A1(n1238), .Z(n576));
Q_OR02 U1362 ( .A0(n577), .A1(n576), .Z(n578));
Q_MX02 U1363 ( .S(cur_state[1]), .A0(n578), .A1(n574), .Z(n579));
Q_OR02 U1364 ( .A0(cmdfifo_gcm_cmd[0]), .A1(n580), .Z(n610));
Q_OA21 U1365 ( .A0(beat_num[0]), .A1(n610), .B0(beat_num[1]), .Z(n581));
Q_AO21 U1366 ( .A0(n610), .A1(n597), .B0(n581), .Z(n586));
Q_OR02 U1367 ( .A0(n622), .A1(n586), .Z(n582));
Q_INV U1368 ( .A(n582), .Z(n546));
Q_XOR2 U1369 ( .A0(cmdfifo_gcm_cmd[1]), .A1(n583), .Z(n591));
Q_ND02 U1370 ( .A0(n606), .A1(n592), .Z(n584));
Q_OR02 U1371 ( .A0(ciph_fifo_in_stall), .A1(n584), .Z(n585));
Q_ND02 U1372 ( .A0(upsizer_gcm_valid), .A1(n586), .Z(n587));
Q_MX02 U1373 ( .S(cur_state[0]), .A0(n587), .A1(n585), .Z(n588));
Q_OR03 U1374 ( .A0(cur_state[2]), .A1(n588), .A2(n1237), .Z(n589));
Q_ND02 U1375 ( .A0(n589), .A1(n603), .Z(n590));
Q_OR02 U1376 ( .A0(cmdfifo_gcm_cmd[0]), .A1(n591), .Z(n592));
Q_INV U1377 ( .A(n592), .Z(n593));
Q_OR02 U1378 ( .A0(ciph_fifo_in_stall), .A1(n593), .Z(n594));
Q_AN02 U1379 ( .A0(cmdfifo_gcm_cmd[2]), .A1(n1224), .Z(n595));
Q_OR02 U1380 ( .A0(n555), .A1(n595), .Z(n596));
Q_MX02 U1381 ( .S(beat_num[0]), .A0(n624), .A1(n596), .Z(n598));
Q_AO21 U1382 ( .A0(n598), .A1(n597), .B0(n581), .Z(n599));
Q_OR02 U1383 ( .A0(n620), .A1(n599), .Z(n600));
Q_MX02 U1384 ( .S(cur_state[0]), .A0(n600), .A1(n594), .Z(n601));
Q_OR03 U1385 ( .A0(cur_state[2]), .A1(n601), .A2(n1237), .Z(n604));
Q_OR02 U1386 ( .A0(n602), .A1(cur_state[1]), .Z(n603));
Q_AN02 U1387 ( .A0(n604), .A1(n603), .Z(n547));
Q_AO21 U1388 ( .A0(combo_dek512), .A1(cmdfifo_gcm_cmd[2]), .B0(n606), .Z(n607));
Q_ND02 U1389 ( .A0(cmdfifo_gcm_cmd[0]), .A1(cmdfifo_gcm_cmd[1]), .Z(n606));
Q_INV U1390 ( .A(n607), .Z(n608));
Q_OR02 U1391 ( .A0(ciph_fifo_in_stall), .A1(n608), .Z(n609));
Q_OA21 U1392 ( .A0(n611), .A1(n610), .B0(upsizer_gcm_valid), .Z(n612));
Q_INV U1393 ( .A(n612), .Z(n613));
Q_MX02 U1394 ( .S(cur_state[0]), .A0(n613), .A1(n609), .Z(n614));
Q_OR02 U1395 ( .A0(cur_state[2]), .A1(n614), .Z(n615));
Q_OR02 U1396 ( .A0(cur_state[0]), .A1(n616), .Z(n617));
Q_AO21 U1397 ( .A0(n617), .A1(cur_state[2]), .B0(n576), .Z(n619));
Q_MX02 U1398 ( .S(cur_state[1]), .A0(n619), .A1(n615), .Z(n548));
Q_OR02 U1399 ( .A0(cur_state[0]), .A1(n620), .Z(n621));
Q_OR02 U1400 ( .A0(n1649), .A1(n621), .Z(n622));
Q_OR02 U1401 ( .A0(n622), .A1(n628), .Z(n623));
Q_ND02 U1402 ( .A0(upsizer_gcm_valid), .A1(n624), .Z(n625));
Q_OR02 U1403 ( .A0(n1237), .A1(n630), .Z(n626));
Q_NR02 U1404 ( .A0(n626), .A1(n625), .Z(n627));
Q_ND03 U1405 ( .A0(upsizer_gcm_valid), .A1(n539), .A2(n628), .Z(n629));
Q_OR02 U1406 ( .A0(cur_state[2]), .A1(cur_state[0]), .Z(n630));
Q_OR03 U1407 ( .A0(n630), .A1(n629), .A2(n1237), .Z(n633));
Q_OR02 U1408 ( .A0(n631), .A1(cur_state[1]), .Z(n632));
Q_AN02 U1409 ( .A0(n633), .A1(n632), .Z(n550));
Q_INV U1410 ( .A(n633), .Z(n551));
Q_MX02 U1411 ( .S(n553), .A0(n634), .A1(n543), .Z(gcm_cmdfifo_ack));
Q_MX02 U1412 ( .S(n558), .A0(n1221), .A1(n539), .Z(n1220));
Q_OR02 U1413 ( .A0(n626), .A1(ciph_fifo_in_stall), .Z(gcm_upsizer_stall));
Q_AN02 U1414 ( .A0(n3), .A1(iv_counter[127]), .Z(ciph_in[127]));
Q_AN02 U1415 ( .A0(n3), .A1(iv_counter[126]), .Z(ciph_in[126]));
Q_AN02 U1416 ( .A0(n3), .A1(iv_counter[125]), .Z(ciph_in[125]));
Q_AN02 U1417 ( .A0(n3), .A1(iv_counter[124]), .Z(ciph_in[124]));
Q_AN02 U1418 ( .A0(n3), .A1(iv_counter[123]), .Z(ciph_in[123]));
Q_AN02 U1419 ( .A0(n3), .A1(iv_counter[122]), .Z(ciph_in[122]));
Q_AN02 U1420 ( .A0(n3), .A1(iv_counter[121]), .Z(ciph_in[121]));
Q_AN02 U1421 ( .A0(n3), .A1(iv_counter[120]), .Z(ciph_in[120]));
Q_AN02 U1422 ( .A0(n3), .A1(iv_counter[119]), .Z(ciph_in[119]));
Q_AN02 U1423 ( .A0(n3), .A1(iv_counter[118]), .Z(ciph_in[118]));
Q_AN02 U1424 ( .A0(n3), .A1(iv_counter[117]), .Z(ciph_in[117]));
Q_AN02 U1425 ( .A0(n3), .A1(iv_counter[116]), .Z(ciph_in[116]));
Q_AN02 U1426 ( .A0(n3), .A1(iv_counter[115]), .Z(ciph_in[115]));
Q_AN02 U1427 ( .A0(n3), .A1(iv_counter[114]), .Z(ciph_in[114]));
Q_AN02 U1428 ( .A0(n3), .A1(iv_counter[113]), .Z(ciph_in[113]));
Q_AN02 U1429 ( .A0(n3), .A1(iv_counter[112]), .Z(ciph_in[112]));
Q_AN02 U1430 ( .A0(n3), .A1(iv_counter[111]), .Z(ciph_in[111]));
Q_AN02 U1431 ( .A0(n3), .A1(iv_counter[110]), .Z(ciph_in[110]));
Q_AN02 U1432 ( .A0(n3), .A1(iv_counter[109]), .Z(ciph_in[109]));
Q_AN02 U1433 ( .A0(n3), .A1(iv_counter[108]), .Z(ciph_in[108]));
Q_AN02 U1434 ( .A0(n3), .A1(iv_counter[107]), .Z(ciph_in[107]));
Q_AN02 U1435 ( .A0(n3), .A1(iv_counter[106]), .Z(ciph_in[106]));
Q_AN02 U1436 ( .A0(n3), .A1(iv_counter[105]), .Z(ciph_in[105]));
Q_AN02 U1437 ( .A0(n3), .A1(iv_counter[104]), .Z(ciph_in[104]));
Q_AN02 U1438 ( .A0(n3), .A1(iv_counter[103]), .Z(ciph_in[103]));
Q_AN02 U1439 ( .A0(n3), .A1(iv_counter[102]), .Z(ciph_in[102]));
Q_AN02 U1440 ( .A0(n3), .A1(iv_counter[101]), .Z(ciph_in[101]));
Q_AN02 U1441 ( .A0(n3), .A1(iv_counter[100]), .Z(ciph_in[100]));
Q_AN02 U1442 ( .A0(n3), .A1(iv_counter[99]), .Z(ciph_in[99]));
Q_AN02 U1443 ( .A0(n3), .A1(iv_counter[98]), .Z(ciph_in[98]));
Q_AN02 U1444 ( .A0(n3), .A1(iv_counter[97]), .Z(ciph_in[97]));
Q_AN02 U1445 ( .A0(n3), .A1(iv_counter[96]), .Z(ciph_in[96]));
Q_AN02 U1446 ( .A0(n3), .A1(iv_counter[95]), .Z(ciph_in[95]));
Q_AN02 U1447 ( .A0(n3), .A1(iv_counter[94]), .Z(ciph_in[94]));
Q_AN02 U1448 ( .A0(n3), .A1(iv_counter[93]), .Z(ciph_in[93]));
Q_AN02 U1449 ( .A0(n3), .A1(iv_counter[92]), .Z(ciph_in[92]));
Q_AN02 U1450 ( .A0(n3), .A1(iv_counter[91]), .Z(ciph_in[91]));
Q_AN02 U1451 ( .A0(n3), .A1(iv_counter[90]), .Z(ciph_in[90]));
Q_AN02 U1452 ( .A0(n3), .A1(iv_counter[89]), .Z(ciph_in[89]));
Q_AN02 U1453 ( .A0(n3), .A1(iv_counter[88]), .Z(ciph_in[88]));
Q_AN02 U1454 ( .A0(n3), .A1(iv_counter[87]), .Z(ciph_in[87]));
Q_AN02 U1455 ( .A0(n3), .A1(iv_counter[86]), .Z(ciph_in[86]));
Q_AN02 U1456 ( .A0(n3), .A1(iv_counter[85]), .Z(ciph_in[85]));
Q_AN02 U1457 ( .A0(n3), .A1(iv_counter[84]), .Z(ciph_in[84]));
Q_AN02 U1458 ( .A0(n3), .A1(iv_counter[83]), .Z(ciph_in[83]));
Q_AN02 U1459 ( .A0(n3), .A1(iv_counter[82]), .Z(ciph_in[82]));
Q_AN02 U1460 ( .A0(n3), .A1(iv_counter[81]), .Z(ciph_in[81]));
Q_AN02 U1461 ( .A0(n3), .A1(iv_counter[80]), .Z(ciph_in[80]));
Q_AN02 U1462 ( .A0(n3), .A1(iv_counter[79]), .Z(ciph_in[79]));
Q_AN02 U1463 ( .A0(n3), .A1(iv_counter[78]), .Z(ciph_in[78]));
Q_AN02 U1464 ( .A0(n3), .A1(iv_counter[77]), .Z(ciph_in[77]));
Q_AN02 U1465 ( .A0(n3), .A1(iv_counter[76]), .Z(ciph_in[76]));
Q_AN02 U1466 ( .A0(n3), .A1(iv_counter[75]), .Z(ciph_in[75]));
Q_AN02 U1467 ( .A0(n3), .A1(iv_counter[74]), .Z(ciph_in[74]));
Q_AN02 U1468 ( .A0(n3), .A1(iv_counter[73]), .Z(ciph_in[73]));
Q_AN02 U1469 ( .A0(n3), .A1(iv_counter[72]), .Z(ciph_in[72]));
Q_AN02 U1470 ( .A0(n3), .A1(iv_counter[71]), .Z(ciph_in[71]));
Q_AN02 U1471 ( .A0(n3), .A1(iv_counter[70]), .Z(ciph_in[70]));
Q_AN02 U1472 ( .A0(n3), .A1(iv_counter[69]), .Z(ciph_in[69]));
Q_AN02 U1473 ( .A0(n3), .A1(iv_counter[68]), .Z(ciph_in[68]));
Q_AN02 U1474 ( .A0(n3), .A1(iv_counter[67]), .Z(ciph_in[67]));
Q_AN02 U1475 ( .A0(n3), .A1(iv_counter[66]), .Z(ciph_in[66]));
Q_AN02 U1476 ( .A0(n3), .A1(iv_counter[65]), .Z(ciph_in[65]));
Q_AN02 U1477 ( .A0(n3), .A1(iv_counter[64]), .Z(ciph_in[64]));
Q_AN02 U1478 ( .A0(n3), .A1(iv_counter[63]), .Z(ciph_in[63]));
Q_AN02 U1479 ( .A0(n3), .A1(iv_counter[62]), .Z(ciph_in[62]));
Q_AN02 U1480 ( .A0(n3), .A1(iv_counter[61]), .Z(ciph_in[61]));
Q_AN02 U1481 ( .A0(n3), .A1(iv_counter[60]), .Z(ciph_in[60]));
Q_AN02 U1482 ( .A0(n3), .A1(iv_counter[59]), .Z(ciph_in[59]));
Q_AN02 U1483 ( .A0(n3), .A1(iv_counter[58]), .Z(ciph_in[58]));
Q_AN02 U1484 ( .A0(n3), .A1(iv_counter[57]), .Z(ciph_in[57]));
Q_AN02 U1485 ( .A0(n3), .A1(iv_counter[56]), .Z(ciph_in[56]));
Q_AN02 U1486 ( .A0(n3), .A1(iv_counter[55]), .Z(ciph_in[55]));
Q_AN02 U1487 ( .A0(n3), .A1(iv_counter[54]), .Z(ciph_in[54]));
Q_AN02 U1488 ( .A0(n3), .A1(iv_counter[53]), .Z(ciph_in[53]));
Q_AN02 U1489 ( .A0(n3), .A1(iv_counter[52]), .Z(ciph_in[52]));
Q_AN02 U1490 ( .A0(n3), .A1(iv_counter[51]), .Z(ciph_in[51]));
Q_AN02 U1491 ( .A0(n3), .A1(iv_counter[50]), .Z(ciph_in[50]));
Q_AN02 U1492 ( .A0(n3), .A1(iv_counter[49]), .Z(ciph_in[49]));
Q_AN02 U1493 ( .A0(n3), .A1(iv_counter[48]), .Z(ciph_in[48]));
Q_AN02 U1494 ( .A0(n3), .A1(iv_counter[47]), .Z(ciph_in[47]));
Q_AN02 U1495 ( .A0(n3), .A1(iv_counter[46]), .Z(ciph_in[46]));
Q_AN02 U1496 ( .A0(n3), .A1(iv_counter[45]), .Z(ciph_in[45]));
Q_AN02 U1497 ( .A0(n3), .A1(iv_counter[44]), .Z(ciph_in[44]));
Q_AN02 U1498 ( .A0(n3), .A1(iv_counter[43]), .Z(ciph_in[43]));
Q_AN02 U1499 ( .A0(n3), .A1(iv_counter[42]), .Z(ciph_in[42]));
Q_AN02 U1500 ( .A0(n3), .A1(iv_counter[41]), .Z(ciph_in[41]));
Q_AN02 U1501 ( .A0(n3), .A1(iv_counter[40]), .Z(ciph_in[40]));
Q_AN02 U1502 ( .A0(n3), .A1(iv_counter[39]), .Z(ciph_in[39]));
Q_AN02 U1503 ( .A0(n3), .A1(iv_counter[38]), .Z(ciph_in[38]));
Q_AN02 U1504 ( .A0(n3), .A1(iv_counter[37]), .Z(ciph_in[37]));
Q_AN02 U1505 ( .A0(n3), .A1(iv_counter[36]), .Z(ciph_in[36]));
Q_AN02 U1506 ( .A0(n3), .A1(iv_counter[35]), .Z(ciph_in[35]));
Q_AN02 U1507 ( .A0(n3), .A1(iv_counter[34]), .Z(ciph_in[34]));
Q_AN02 U1508 ( .A0(n3), .A1(iv_counter[33]), .Z(ciph_in[33]));
Q_AN02 U1509 ( .A0(n3), .A1(iv_counter[32]), .Z(ciph_in[32]));
Q_AN02 U1510 ( .A0(n549), .A1(iv_counter[31]), .Z(ciph_in[31]));
Q_AN02 U1511 ( .A0(n549), .A1(iv_counter[30]), .Z(ciph_in[30]));
Q_AN02 U1512 ( .A0(n549), .A1(iv_counter[29]), .Z(ciph_in[29]));
Q_AN02 U1513 ( .A0(n549), .A1(iv_counter[28]), .Z(ciph_in[28]));
Q_AN02 U1514 ( .A0(n549), .A1(iv_counter[27]), .Z(ciph_in[27]));
Q_AN02 U1515 ( .A0(n549), .A1(iv_counter[26]), .Z(ciph_in[26]));
Q_AN02 U1516 ( .A0(n549), .A1(iv_counter[25]), .Z(ciph_in[25]));
Q_AN02 U1517 ( .A0(n549), .A1(iv_counter[24]), .Z(ciph_in[24]));
Q_AN02 U1518 ( .A0(n549), .A1(iv_counter[23]), .Z(ciph_in[23]));
Q_AN02 U1519 ( .A0(n549), .A1(iv_counter[22]), .Z(ciph_in[22]));
Q_AN02 U1520 ( .A0(n549), .A1(iv_counter[21]), .Z(ciph_in[21]));
Q_AN02 U1521 ( .A0(n549), .A1(iv_counter[20]), .Z(ciph_in[20]));
Q_AN02 U1522 ( .A0(n549), .A1(iv_counter[19]), .Z(ciph_in[19]));
Q_AN02 U1523 ( .A0(n549), .A1(iv_counter[18]), .Z(ciph_in[18]));
Q_AN02 U1524 ( .A0(n549), .A1(iv_counter[17]), .Z(ciph_in[17]));
Q_AN02 U1525 ( .A0(n549), .A1(iv_counter[16]), .Z(ciph_in[16]));
Q_AN02 U1526 ( .A0(n549), .A1(iv_counter[15]), .Z(ciph_in[15]));
Q_AN02 U1527 ( .A0(n549), .A1(iv_counter[14]), .Z(ciph_in[14]));
Q_AN02 U1528 ( .A0(n549), .A1(iv_counter[13]), .Z(ciph_in[13]));
Q_AN02 U1529 ( .A0(n549), .A1(iv_counter[12]), .Z(ciph_in[12]));
Q_AN02 U1530 ( .A0(n549), .A1(iv_counter[11]), .Z(ciph_in[11]));
Q_AN02 U1531 ( .A0(n549), .A1(iv_counter[10]), .Z(ciph_in[10]));
Q_AN02 U1532 ( .A0(n549), .A1(iv_counter[9]), .Z(ciph_in[9]));
Q_AN02 U1533 ( .A0(n549), .A1(iv_counter[8]), .Z(ciph_in[8]));
Q_AN02 U1534 ( .A0(n549), .A1(iv_counter[7]), .Z(ciph_in[7]));
Q_AN02 U1535 ( .A0(n549), .A1(iv_counter[6]), .Z(ciph_in[6]));
Q_AN02 U1536 ( .A0(n549), .A1(iv_counter[5]), .Z(ciph_in[5]));
Q_AN02 U1537 ( .A0(n549), .A1(iv_counter[4]), .Z(ciph_in[4]));
Q_AN02 U1538 ( .A0(n549), .A1(iv_counter[3]), .Z(ciph_in[3]));
Q_AN02 U1539 ( .A0(n549), .A1(iv_counter[2]), .Z(ciph_in[2]));
Q_AN02 U1540 ( .A0(n549), .A1(iv_counter[1]), .Z(ciph_in[1]));
Q_MX02 U1541 ( .S(n622), .A0(iv_counter[0]), .A1(n560), .Z(ciph_in[0]));
Q_AN02 U1542 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[354]), .Z(key_in[255]));
Q_AN02 U1543 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[353]), .Z(key_in[254]));
Q_AN02 U1544 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[352]), .Z(key_in[253]));
Q_AN02 U1545 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[351]), .Z(key_in[252]));
Q_AN02 U1546 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[350]), .Z(key_in[251]));
Q_AN02 U1547 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[349]), .Z(key_in[250]));
Q_AN02 U1548 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[348]), .Z(key_in[249]));
Q_AN02 U1549 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[347]), .Z(key_in[248]));
Q_AN02 U1550 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[346]), .Z(key_in[247]));
Q_AN02 U1551 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[345]), .Z(key_in[246]));
Q_AN02 U1552 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[344]), .Z(key_in[245]));
Q_AN02 U1553 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[343]), .Z(key_in[244]));
Q_AN02 U1554 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[342]), .Z(key_in[243]));
Q_AN02 U1555 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[341]), .Z(key_in[242]));
Q_AN02 U1556 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[340]), .Z(key_in[241]));
Q_AN02 U1557 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[339]), .Z(key_in[240]));
Q_AN02 U1558 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[338]), .Z(key_in[239]));
Q_AN02 U1559 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[337]), .Z(key_in[238]));
Q_AN02 U1560 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[336]), .Z(key_in[237]));
Q_AN02 U1561 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[335]), .Z(key_in[236]));
Q_AN02 U1562 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[334]), .Z(key_in[235]));
Q_AN02 U1563 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[333]), .Z(key_in[234]));
Q_AN02 U1564 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[332]), .Z(key_in[233]));
Q_AN02 U1565 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[331]), .Z(key_in[232]));
Q_AN02 U1566 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[330]), .Z(key_in[231]));
Q_AN02 U1567 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[329]), .Z(key_in[230]));
Q_AN02 U1568 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[328]), .Z(key_in[229]));
Q_AN02 U1569 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[327]), .Z(key_in[228]));
Q_AN02 U1570 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[326]), .Z(key_in[227]));
Q_AN02 U1571 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[325]), .Z(key_in[226]));
Q_AN02 U1572 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[324]), .Z(key_in[225]));
Q_AN02 U1573 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[323]), .Z(key_in[224]));
Q_AN02 U1574 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[322]), .Z(key_in[223]));
Q_AN02 U1575 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[321]), .Z(key_in[222]));
Q_AN02 U1576 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[320]), .Z(key_in[221]));
Q_AN02 U1577 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[319]), .Z(key_in[220]));
Q_AN02 U1578 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[318]), .Z(key_in[219]));
Q_AN02 U1579 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[317]), .Z(key_in[218]));
Q_AN02 U1580 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[316]), .Z(key_in[217]));
Q_AN02 U1581 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[315]), .Z(key_in[216]));
Q_AN02 U1582 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[314]), .Z(key_in[215]));
Q_AN02 U1583 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[313]), .Z(key_in[214]));
Q_AN02 U1584 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[312]), .Z(key_in[213]));
Q_AN02 U1585 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[311]), .Z(key_in[212]));
Q_AN02 U1586 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[310]), .Z(key_in[211]));
Q_AN02 U1587 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[309]), .Z(key_in[210]));
Q_AN02 U1588 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[308]), .Z(key_in[209]));
Q_AN02 U1589 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[307]), .Z(key_in[208]));
Q_AN02 U1590 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[306]), .Z(key_in[207]));
Q_AN02 U1591 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[305]), .Z(key_in[206]));
Q_AN02 U1592 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[304]), .Z(key_in[205]));
Q_AN02 U1593 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[303]), .Z(key_in[204]));
Q_AN02 U1594 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[302]), .Z(key_in[203]));
Q_AN02 U1595 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[301]), .Z(key_in[202]));
Q_AN02 U1596 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[300]), .Z(key_in[201]));
Q_AN02 U1597 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[299]), .Z(key_in[200]));
Q_AN02 U1598 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[298]), .Z(key_in[199]));
Q_AN02 U1599 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[297]), .Z(key_in[198]));
Q_AN02 U1600 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[296]), .Z(key_in[197]));
Q_AN02 U1601 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[295]), .Z(key_in[196]));
Q_AN02 U1602 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[294]), .Z(key_in[195]));
Q_AN02 U1603 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[293]), .Z(key_in[194]));
Q_AN02 U1604 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[292]), .Z(key_in[193]));
Q_AN02 U1605 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[291]), .Z(key_in[192]));
Q_AN02 U1606 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[290]), .Z(key_in[191]));
Q_AN02 U1607 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[289]), .Z(key_in[190]));
Q_AN02 U1608 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[288]), .Z(key_in[189]));
Q_AN02 U1609 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[287]), .Z(key_in[188]));
Q_AN02 U1610 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[286]), .Z(key_in[187]));
Q_AN02 U1611 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[285]), .Z(key_in[186]));
Q_AN02 U1612 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[284]), .Z(key_in[185]));
Q_AN02 U1613 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[283]), .Z(key_in[184]));
Q_AN02 U1614 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[282]), .Z(key_in[183]));
Q_AN02 U1615 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[281]), .Z(key_in[182]));
Q_AN02 U1616 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[280]), .Z(key_in[181]));
Q_AN02 U1617 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[279]), .Z(key_in[180]));
Q_AN02 U1618 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[278]), .Z(key_in[179]));
Q_AN02 U1619 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[277]), .Z(key_in[178]));
Q_AN02 U1620 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[276]), .Z(key_in[177]));
Q_AN02 U1621 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[275]), .Z(key_in[176]));
Q_AN02 U1622 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[274]), .Z(key_in[175]));
Q_AN02 U1623 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[273]), .Z(key_in[174]));
Q_AN02 U1624 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[272]), .Z(key_in[173]));
Q_AN02 U1625 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[271]), .Z(key_in[172]));
Q_AN02 U1626 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[270]), .Z(key_in[171]));
Q_AN02 U1627 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[269]), .Z(key_in[170]));
Q_AN02 U1628 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[268]), .Z(key_in[169]));
Q_AN02 U1629 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[267]), .Z(key_in[168]));
Q_AN02 U1630 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[266]), .Z(key_in[167]));
Q_AN02 U1631 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[265]), .Z(key_in[166]));
Q_AN02 U1632 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[264]), .Z(key_in[165]));
Q_AN02 U1633 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[263]), .Z(key_in[164]));
Q_AN02 U1634 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[262]), .Z(key_in[163]));
Q_AN02 U1635 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[261]), .Z(key_in[162]));
Q_AN02 U1636 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[260]), .Z(key_in[161]));
Q_AN02 U1637 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[259]), .Z(key_in[160]));
Q_AN02 U1638 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[258]), .Z(key_in[159]));
Q_AN02 U1639 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[257]), .Z(key_in[158]));
Q_AN02 U1640 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[256]), .Z(key_in[157]));
Q_AN02 U1641 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[255]), .Z(key_in[156]));
Q_AN02 U1642 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[254]), .Z(key_in[155]));
Q_AN02 U1643 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[253]), .Z(key_in[154]));
Q_AN02 U1644 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[252]), .Z(key_in[153]));
Q_AN02 U1645 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[251]), .Z(key_in[152]));
Q_AN02 U1646 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[250]), .Z(key_in[151]));
Q_AN02 U1647 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[249]), .Z(key_in[150]));
Q_AN02 U1648 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[248]), .Z(key_in[149]));
Q_AN02 U1649 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[247]), .Z(key_in[148]));
Q_AN02 U1650 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[246]), .Z(key_in[147]));
Q_AN02 U1651 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[245]), .Z(key_in[146]));
Q_AN02 U1652 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[244]), .Z(key_in[145]));
Q_AN02 U1653 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[243]), .Z(key_in[144]));
Q_AN02 U1654 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[242]), .Z(key_in[143]));
Q_AN02 U1655 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[241]), .Z(key_in[142]));
Q_AN02 U1656 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[240]), .Z(key_in[141]));
Q_AN02 U1657 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[239]), .Z(key_in[140]));
Q_AN02 U1658 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[238]), .Z(key_in[139]));
Q_AN02 U1659 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[237]), .Z(key_in[138]));
Q_AN02 U1660 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[236]), .Z(key_in[137]));
Q_AN02 U1661 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[235]), .Z(key_in[136]));
Q_AN02 U1662 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[234]), .Z(key_in[135]));
Q_AN02 U1663 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[233]), .Z(key_in[134]));
Q_AN02 U1664 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[232]), .Z(key_in[133]));
Q_AN02 U1665 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[231]), .Z(key_in[132]));
Q_AN02 U1666 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[230]), .Z(key_in[131]));
Q_AN02 U1667 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[229]), .Z(key_in[130]));
Q_AN02 U1668 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[228]), .Z(key_in[129]));
Q_AN02 U1669 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[227]), .Z(key_in[128]));
Q_AN02 U1670 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[226]), .Z(key_in[127]));
Q_AN02 U1671 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[225]), .Z(key_in[126]));
Q_AN02 U1672 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[224]), .Z(key_in[125]));
Q_AN02 U1673 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[223]), .Z(key_in[124]));
Q_AN02 U1674 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[222]), .Z(key_in[123]));
Q_AN02 U1675 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[221]), .Z(key_in[122]));
Q_AN02 U1676 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[220]), .Z(key_in[121]));
Q_AN02 U1677 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[219]), .Z(key_in[120]));
Q_AN02 U1678 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[218]), .Z(key_in[119]));
Q_AN02 U1679 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[217]), .Z(key_in[118]));
Q_AN02 U1680 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[216]), .Z(key_in[117]));
Q_AN02 U1681 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[215]), .Z(key_in[116]));
Q_AN02 U1682 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[214]), .Z(key_in[115]));
Q_AN02 U1683 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[213]), .Z(key_in[114]));
Q_AN02 U1684 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[212]), .Z(key_in[113]));
Q_AN02 U1685 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[211]), .Z(key_in[112]));
Q_AN02 U1686 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[210]), .Z(key_in[111]));
Q_AN02 U1687 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[209]), .Z(key_in[110]));
Q_AN02 U1688 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[208]), .Z(key_in[109]));
Q_AN02 U1689 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[207]), .Z(key_in[108]));
Q_AN02 U1690 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[206]), .Z(key_in[107]));
Q_AN02 U1691 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[205]), .Z(key_in[106]));
Q_AN02 U1692 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[204]), .Z(key_in[105]));
Q_AN02 U1693 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[203]), .Z(key_in[104]));
Q_AN02 U1694 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[202]), .Z(key_in[103]));
Q_AN02 U1695 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[201]), .Z(key_in[102]));
Q_AN02 U1696 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[200]), .Z(key_in[101]));
Q_AN02 U1697 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[199]), .Z(key_in[100]));
Q_AN02 U1698 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[198]), .Z(key_in[99]));
Q_AN02 U1699 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[197]), .Z(key_in[98]));
Q_AN02 U1700 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[196]), .Z(key_in[97]));
Q_AN02 U1701 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[195]), .Z(key_in[96]));
Q_AN02 U1702 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[194]), .Z(key_in[95]));
Q_AN02 U1703 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[193]), .Z(key_in[94]));
Q_AN02 U1704 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[192]), .Z(key_in[93]));
Q_AN02 U1705 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[191]), .Z(key_in[92]));
Q_AN02 U1706 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[190]), .Z(key_in[91]));
Q_AN02 U1707 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[189]), .Z(key_in[90]));
Q_AN02 U1708 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[188]), .Z(key_in[89]));
Q_AN02 U1709 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[187]), .Z(key_in[88]));
Q_AN02 U1710 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[186]), .Z(key_in[87]));
Q_AN02 U1711 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[185]), .Z(key_in[86]));
Q_AN02 U1712 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[184]), .Z(key_in[85]));
Q_AN02 U1713 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[183]), .Z(key_in[84]));
Q_AN02 U1714 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[182]), .Z(key_in[83]));
Q_AN02 U1715 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[181]), .Z(key_in[82]));
Q_AN02 U1716 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[180]), .Z(key_in[81]));
Q_AN02 U1717 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[179]), .Z(key_in[80]));
Q_AN02 U1718 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[178]), .Z(key_in[79]));
Q_AN02 U1719 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[177]), .Z(key_in[78]));
Q_AN02 U1720 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[176]), .Z(key_in[77]));
Q_AN02 U1721 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[175]), .Z(key_in[76]));
Q_AN02 U1722 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[174]), .Z(key_in[75]));
Q_AN02 U1723 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[173]), .Z(key_in[74]));
Q_AN02 U1724 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[172]), .Z(key_in[73]));
Q_AN02 U1725 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[171]), .Z(key_in[72]));
Q_AN02 U1726 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[170]), .Z(key_in[71]));
Q_AN02 U1727 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[169]), .Z(key_in[70]));
Q_AN02 U1728 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[168]), .Z(key_in[69]));
Q_AN02 U1729 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[167]), .Z(key_in[68]));
Q_AN02 U1730 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[166]), .Z(key_in[67]));
Q_AN02 U1731 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[165]), .Z(key_in[66]));
Q_AN02 U1732 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[164]), .Z(key_in[65]));
Q_AN02 U1733 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[163]), .Z(key_in[64]));
Q_AN02 U1734 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[162]), .Z(key_in[63]));
Q_AN02 U1735 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[161]), .Z(key_in[62]));
Q_AN02 U1736 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[160]), .Z(key_in[61]));
Q_AN02 U1737 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[159]), .Z(key_in[60]));
Q_AN02 U1738 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[158]), .Z(key_in[59]));
Q_AN02 U1739 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[157]), .Z(key_in[58]));
Q_AN02 U1740 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[156]), .Z(key_in[57]));
Q_AN02 U1741 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[155]), .Z(key_in[56]));
Q_AN02 U1742 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[154]), .Z(key_in[55]));
Q_AN02 U1743 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[153]), .Z(key_in[54]));
Q_AN02 U1744 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[152]), .Z(key_in[53]));
Q_AN02 U1745 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[151]), .Z(key_in[52]));
Q_AN02 U1746 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[150]), .Z(key_in[51]));
Q_AN02 U1747 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[149]), .Z(key_in[50]));
Q_AN02 U1748 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[148]), .Z(key_in[49]));
Q_AN02 U1749 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[147]), .Z(key_in[48]));
Q_AN02 U1750 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[146]), .Z(key_in[47]));
Q_AN02 U1751 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[145]), .Z(key_in[46]));
Q_AN02 U1752 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[144]), .Z(key_in[45]));
Q_AN02 U1753 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[143]), .Z(key_in[44]));
Q_AN02 U1754 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[142]), .Z(key_in[43]));
Q_AN02 U1755 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[141]), .Z(key_in[42]));
Q_AN02 U1756 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[140]), .Z(key_in[41]));
Q_AN02 U1757 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[139]), .Z(key_in[40]));
Q_AN02 U1758 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[138]), .Z(key_in[39]));
Q_AN02 U1759 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[137]), .Z(key_in[38]));
Q_AN02 U1760 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[136]), .Z(key_in[37]));
Q_AN02 U1761 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[135]), .Z(key_in[36]));
Q_AN02 U1762 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[134]), .Z(key_in[35]));
Q_AN02 U1763 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[133]), .Z(key_in[34]));
Q_AN02 U1764 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[132]), .Z(key_in[33]));
Q_AN02 U1765 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[131]), .Z(key_in[32]));
Q_AN02 U1766 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[130]), .Z(key_in[31]));
Q_AN02 U1767 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[129]), .Z(key_in[30]));
Q_AN02 U1768 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[128]), .Z(key_in[29]));
Q_AN02 U1769 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[127]), .Z(key_in[28]));
Q_AN02 U1770 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[126]), .Z(key_in[27]));
Q_AN02 U1771 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[125]), .Z(key_in[26]));
Q_AN02 U1772 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[124]), .Z(key_in[25]));
Q_AN02 U1773 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[123]), .Z(key_in[24]));
Q_AN02 U1774 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[122]), .Z(key_in[23]));
Q_AN02 U1775 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[121]), .Z(key_in[22]));
Q_AN02 U1776 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[120]), .Z(key_in[21]));
Q_AN02 U1777 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[119]), .Z(key_in[20]));
Q_AN02 U1778 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[118]), .Z(key_in[19]));
Q_AN02 U1779 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[117]), .Z(key_in[18]));
Q_AN02 U1780 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[116]), .Z(key_in[17]));
Q_AN02 U1781 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[115]), .Z(key_in[16]));
Q_AN02 U1782 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[114]), .Z(key_in[15]));
Q_AN02 U1783 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[113]), .Z(key_in[14]));
Q_AN02 U1784 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[112]), .Z(key_in[13]));
Q_AN02 U1785 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[111]), .Z(key_in[12]));
Q_AN02 U1786 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[110]), .Z(key_in[11]));
Q_AN02 U1787 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[109]), .Z(key_in[10]));
Q_AN02 U1788 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[108]), .Z(key_in[9]));
Q_AN02 U1789 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[107]), .Z(key_in[8]));
Q_AN02 U1790 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[106]), .Z(key_in[7]));
Q_AN02 U1791 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[105]), .Z(key_in[6]));
Q_AN02 U1792 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[104]), .Z(key_in[5]));
Q_AN02 U1793 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[103]), .Z(key_in[4]));
Q_AN02 U1794 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[102]), .Z(key_in[3]));
Q_AN02 U1795 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[101]), .Z(key_in[2]));
Q_AN02 U1796 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[100]), .Z(key_in[1]));
Q_AN02 U1797 ( .A0(key_in_vld), .A1(cmdfifo_gcm_cmd[99]), .Z(key_in[0]));
Q_AN02 U1798 ( .A0(n635), .A1(n571), .Z(fifo_in[131]));
Q_INV U1799 ( .A(n544), .Z(n635));
Q_AN02 U1800 ( .A0(n545), .A1(n579), .Z(fifo_in[130]));
Q_MX02 U1801 ( .S(n544), .A0(n636), .A1(n637), .Z(fifo_in[129]));
Q_ND02 U1802 ( .A0(n571), .A1(n579), .Z(n636));
Q_NR02 U1803 ( .A0(n571), .A1(n579), .Z(n637));
Q_MX02 U1804 ( .S(n582), .A0(n642), .A1(n638), .Z(fifo_in[128]));
Q_AN02 U1805 ( .A0(n590), .A1(n639), .Z(n638));
Q_MX02 U1806 ( .S(n547), .A0(n640), .A1(n641), .Z(n639));
Q_AN02 U1807 ( .A0(n548), .A1(gcm_tag_data_out[95]), .Z(n640));
Q_MX02 U1808 ( .S(n548), .A0(upsizer_gcm_data[127]), .A1(cmdfifo_gcm_cmd[226]), .Z(n641));
Q_MX03 U1809 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[354]), .A1(cmdfifo_gcm_cmd[482]), .A2(cmdfifo_gcm_cmd[610]), .Z(n642));
Q_MX02 U1810 ( .S(n582), .A0(n647), .A1(n643), .Z(fifo_in[127]));
Q_AN02 U1811 ( .A0(n590), .A1(n644), .Z(n643));
Q_MX02 U1812 ( .S(n547), .A0(n645), .A1(n646), .Z(n644));
Q_AN02 U1813 ( .A0(n548), .A1(gcm_tag_data_out[94]), .Z(n645));
Q_MX02 U1814 ( .S(n548), .A0(upsizer_gcm_data[126]), .A1(cmdfifo_gcm_cmd[225]), .Z(n646));
Q_MX03 U1815 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[353]), .A1(cmdfifo_gcm_cmd[481]), .A2(cmdfifo_gcm_cmd[609]), .Z(n647));
Q_MX02 U1816 ( .S(n582), .A0(n652), .A1(n648), .Z(fifo_in[126]));
Q_AN02 U1817 ( .A0(n590), .A1(n649), .Z(n648));
Q_MX02 U1818 ( .S(n547), .A0(n650), .A1(n651), .Z(n649));
Q_AN02 U1819 ( .A0(n548), .A1(gcm_tag_data_out[93]), .Z(n650));
Q_MX02 U1820 ( .S(n548), .A0(upsizer_gcm_data[125]), .A1(cmdfifo_gcm_cmd[224]), .Z(n651));
Q_MX03 U1821 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[352]), .A1(cmdfifo_gcm_cmd[480]), .A2(cmdfifo_gcm_cmd[608]), .Z(n652));
Q_MX02 U1822 ( .S(n582), .A0(n657), .A1(n653), .Z(fifo_in[125]));
Q_AN02 U1823 ( .A0(n590), .A1(n654), .Z(n653));
Q_MX02 U1824 ( .S(n547), .A0(n655), .A1(n656), .Z(n654));
Q_AN02 U1825 ( .A0(n548), .A1(gcm_tag_data_out[92]), .Z(n655));
Q_MX02 U1826 ( .S(n548), .A0(upsizer_gcm_data[124]), .A1(cmdfifo_gcm_cmd[223]), .Z(n656));
Q_MX03 U1827 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[351]), .A1(cmdfifo_gcm_cmd[479]), .A2(cmdfifo_gcm_cmd[607]), .Z(n657));
Q_MX02 U1828 ( .S(n582), .A0(n662), .A1(n658), .Z(fifo_in[124]));
Q_AN02 U1829 ( .A0(n590), .A1(n659), .Z(n658));
Q_MX02 U1830 ( .S(n547), .A0(n660), .A1(n661), .Z(n659));
Q_AN02 U1831 ( .A0(n548), .A1(gcm_tag_data_out[91]), .Z(n660));
Q_MX02 U1832 ( .S(n548), .A0(upsizer_gcm_data[123]), .A1(cmdfifo_gcm_cmd[222]), .Z(n661));
Q_MX03 U1833 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[350]), .A1(cmdfifo_gcm_cmd[478]), .A2(cmdfifo_gcm_cmd[606]), .Z(n662));
Q_MX02 U1834 ( .S(n582), .A0(n667), .A1(n663), .Z(fifo_in[123]));
Q_AN02 U1835 ( .A0(n590), .A1(n664), .Z(n663));
Q_MX02 U1836 ( .S(n547), .A0(n665), .A1(n666), .Z(n664));
Q_AN02 U1837 ( .A0(n548), .A1(gcm_tag_data_out[90]), .Z(n665));
Q_MX02 U1838 ( .S(n548), .A0(upsizer_gcm_data[122]), .A1(cmdfifo_gcm_cmd[221]), .Z(n666));
Q_MX03 U1839 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[349]), .A1(cmdfifo_gcm_cmd[477]), .A2(cmdfifo_gcm_cmd[605]), .Z(n667));
Q_MX02 U1840 ( .S(n582), .A0(n672), .A1(n668), .Z(fifo_in[122]));
Q_AN02 U1841 ( .A0(n590), .A1(n669), .Z(n668));
Q_MX02 U1842 ( .S(n547), .A0(n670), .A1(n671), .Z(n669));
Q_AN02 U1843 ( .A0(n548), .A1(gcm_tag_data_out[89]), .Z(n670));
Q_MX02 U1844 ( .S(n548), .A0(upsizer_gcm_data[121]), .A1(cmdfifo_gcm_cmd[220]), .Z(n671));
Q_MX03 U1845 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[348]), .A1(cmdfifo_gcm_cmd[476]), .A2(cmdfifo_gcm_cmd[604]), .Z(n672));
Q_MX02 U1846 ( .S(n582), .A0(n677), .A1(n673), .Z(fifo_in[121]));
Q_AN02 U1847 ( .A0(n590), .A1(n674), .Z(n673));
Q_MX02 U1848 ( .S(n547), .A0(n675), .A1(n676), .Z(n674));
Q_AN02 U1849 ( .A0(n548), .A1(gcm_tag_data_out[88]), .Z(n675));
Q_MX02 U1850 ( .S(n548), .A0(upsizer_gcm_data[120]), .A1(cmdfifo_gcm_cmd[219]), .Z(n676));
Q_MX03 U1851 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[347]), .A1(cmdfifo_gcm_cmd[475]), .A2(cmdfifo_gcm_cmd[603]), .Z(n677));
Q_MX02 U1852 ( .S(n582), .A0(n682), .A1(n678), .Z(fifo_in[120]));
Q_AN02 U1853 ( .A0(n590), .A1(n679), .Z(n678));
Q_MX02 U1854 ( .S(n547), .A0(n680), .A1(n681), .Z(n679));
Q_AN02 U1855 ( .A0(n548), .A1(gcm_tag_data_out[87]), .Z(n680));
Q_MX02 U1856 ( .S(n548), .A0(upsizer_gcm_data[119]), .A1(cmdfifo_gcm_cmd[218]), .Z(n681));
Q_MX03 U1857 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[346]), .A1(cmdfifo_gcm_cmd[474]), .A2(cmdfifo_gcm_cmd[602]), .Z(n682));
Q_MX02 U1858 ( .S(n582), .A0(n687), .A1(n683), .Z(fifo_in[119]));
Q_AN02 U1859 ( .A0(n590), .A1(n684), .Z(n683));
Q_MX02 U1860 ( .S(n547), .A0(n685), .A1(n686), .Z(n684));
Q_AN02 U1861 ( .A0(n548), .A1(gcm_tag_data_out[86]), .Z(n685));
Q_MX02 U1862 ( .S(n548), .A0(upsizer_gcm_data[118]), .A1(cmdfifo_gcm_cmd[217]), .Z(n686));
Q_MX03 U1863 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[345]), .A1(cmdfifo_gcm_cmd[473]), .A2(cmdfifo_gcm_cmd[601]), .Z(n687));
Q_MX02 U1864 ( .S(n582), .A0(n692), .A1(n688), .Z(fifo_in[118]));
Q_AN02 U1865 ( .A0(n590), .A1(n689), .Z(n688));
Q_MX02 U1866 ( .S(n547), .A0(n690), .A1(n691), .Z(n689));
Q_AN02 U1867 ( .A0(n548), .A1(gcm_tag_data_out[85]), .Z(n690));
Q_MX02 U1868 ( .S(n548), .A0(upsizer_gcm_data[117]), .A1(cmdfifo_gcm_cmd[216]), .Z(n691));
Q_MX03 U1869 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[344]), .A1(cmdfifo_gcm_cmd[472]), .A2(cmdfifo_gcm_cmd[600]), .Z(n692));
Q_MX02 U1870 ( .S(n582), .A0(n697), .A1(n693), .Z(fifo_in[117]));
Q_AN02 U1871 ( .A0(n590), .A1(n694), .Z(n693));
Q_MX02 U1872 ( .S(n547), .A0(n695), .A1(n696), .Z(n694));
Q_AN02 U1873 ( .A0(n548), .A1(gcm_tag_data_out[84]), .Z(n695));
Q_MX02 U1874 ( .S(n548), .A0(upsizer_gcm_data[116]), .A1(cmdfifo_gcm_cmd[215]), .Z(n696));
Q_MX03 U1875 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[343]), .A1(cmdfifo_gcm_cmd[471]), .A2(cmdfifo_gcm_cmd[599]), .Z(n697));
Q_MX02 U1876 ( .S(n582), .A0(n702), .A1(n698), .Z(fifo_in[116]));
Q_AN02 U1877 ( .A0(n590), .A1(n699), .Z(n698));
Q_MX02 U1878 ( .S(n547), .A0(n700), .A1(n701), .Z(n699));
Q_AN02 U1879 ( .A0(n548), .A1(gcm_tag_data_out[83]), .Z(n700));
Q_MX02 U1880 ( .S(n548), .A0(upsizer_gcm_data[115]), .A1(cmdfifo_gcm_cmd[214]), .Z(n701));
Q_MX03 U1881 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[342]), .A1(cmdfifo_gcm_cmd[470]), .A2(cmdfifo_gcm_cmd[598]), .Z(n702));
Q_MX02 U1882 ( .S(n582), .A0(n707), .A1(n703), .Z(fifo_in[115]));
Q_AN02 U1883 ( .A0(n590), .A1(n704), .Z(n703));
Q_MX02 U1884 ( .S(n547), .A0(n705), .A1(n706), .Z(n704));
Q_AN02 U1885 ( .A0(n548), .A1(gcm_tag_data_out[82]), .Z(n705));
Q_MX02 U1886 ( .S(n548), .A0(upsizer_gcm_data[114]), .A1(cmdfifo_gcm_cmd[213]), .Z(n706));
Q_MX03 U1887 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[341]), .A1(cmdfifo_gcm_cmd[469]), .A2(cmdfifo_gcm_cmd[597]), .Z(n707));
Q_MX02 U1888 ( .S(n582), .A0(n712), .A1(n708), .Z(fifo_in[114]));
Q_AN02 U1889 ( .A0(n590), .A1(n709), .Z(n708));
Q_MX02 U1890 ( .S(n547), .A0(n710), .A1(n711), .Z(n709));
Q_AN02 U1891 ( .A0(n548), .A1(gcm_tag_data_out[81]), .Z(n710));
Q_MX02 U1892 ( .S(n548), .A0(upsizer_gcm_data[113]), .A1(cmdfifo_gcm_cmd[212]), .Z(n711));
Q_MX03 U1893 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[340]), .A1(cmdfifo_gcm_cmd[468]), .A2(cmdfifo_gcm_cmd[596]), .Z(n712));
Q_MX02 U1894 ( .S(n582), .A0(n717), .A1(n713), .Z(fifo_in[113]));
Q_AN02 U1895 ( .A0(n590), .A1(n714), .Z(n713));
Q_MX02 U1896 ( .S(n547), .A0(n715), .A1(n716), .Z(n714));
Q_AN02 U1897 ( .A0(n548), .A1(gcm_tag_data_out[80]), .Z(n715));
Q_MX02 U1898 ( .S(n548), .A0(upsizer_gcm_data[112]), .A1(cmdfifo_gcm_cmd[211]), .Z(n716));
Q_MX03 U1899 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[339]), .A1(cmdfifo_gcm_cmd[467]), .A2(cmdfifo_gcm_cmd[595]), .Z(n717));
Q_MX02 U1900 ( .S(n582), .A0(n722), .A1(n718), .Z(fifo_in[112]));
Q_AN02 U1901 ( .A0(n590), .A1(n719), .Z(n718));
Q_MX02 U1902 ( .S(n547), .A0(n720), .A1(n721), .Z(n719));
Q_AN02 U1903 ( .A0(n548), .A1(gcm_tag_data_out[79]), .Z(n720));
Q_MX02 U1904 ( .S(n548), .A0(upsizer_gcm_data[111]), .A1(cmdfifo_gcm_cmd[210]), .Z(n721));
Q_MX03 U1905 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[338]), .A1(cmdfifo_gcm_cmd[466]), .A2(cmdfifo_gcm_cmd[594]), .Z(n722));
Q_MX02 U1906 ( .S(n582), .A0(n727), .A1(n723), .Z(fifo_in[111]));
Q_AN02 U1907 ( .A0(n590), .A1(n724), .Z(n723));
Q_MX02 U1908 ( .S(n547), .A0(n725), .A1(n726), .Z(n724));
Q_AN02 U1909 ( .A0(n548), .A1(gcm_tag_data_out[78]), .Z(n725));
Q_MX02 U1910 ( .S(n548), .A0(upsizer_gcm_data[110]), .A1(cmdfifo_gcm_cmd[209]), .Z(n726));
Q_MX03 U1911 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[337]), .A1(cmdfifo_gcm_cmd[465]), .A2(cmdfifo_gcm_cmd[593]), .Z(n727));
Q_MX02 U1912 ( .S(n582), .A0(n732), .A1(n728), .Z(fifo_in[110]));
Q_AN02 U1913 ( .A0(n590), .A1(n729), .Z(n728));
Q_MX02 U1914 ( .S(n547), .A0(n730), .A1(n731), .Z(n729));
Q_AN02 U1915 ( .A0(n548), .A1(gcm_tag_data_out[77]), .Z(n730));
Q_MX02 U1916 ( .S(n548), .A0(upsizer_gcm_data[109]), .A1(cmdfifo_gcm_cmd[208]), .Z(n731));
Q_MX03 U1917 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[336]), .A1(cmdfifo_gcm_cmd[464]), .A2(cmdfifo_gcm_cmd[592]), .Z(n732));
Q_MX02 U1918 ( .S(n582), .A0(n737), .A1(n733), .Z(fifo_in[109]));
Q_AN02 U1919 ( .A0(n590), .A1(n734), .Z(n733));
Q_MX02 U1920 ( .S(n547), .A0(n735), .A1(n736), .Z(n734));
Q_AN02 U1921 ( .A0(n548), .A1(gcm_tag_data_out[76]), .Z(n735));
Q_MX02 U1922 ( .S(n548), .A0(upsizer_gcm_data[108]), .A1(cmdfifo_gcm_cmd[207]), .Z(n736));
Q_MX03 U1923 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[335]), .A1(cmdfifo_gcm_cmd[463]), .A2(cmdfifo_gcm_cmd[591]), .Z(n737));
Q_MX02 U1924 ( .S(n582), .A0(n742), .A1(n738), .Z(fifo_in[108]));
Q_AN02 U1925 ( .A0(n590), .A1(n739), .Z(n738));
Q_MX02 U1926 ( .S(n547), .A0(n740), .A1(n741), .Z(n739));
Q_AN02 U1927 ( .A0(n548), .A1(gcm_tag_data_out[75]), .Z(n740));
Q_MX02 U1928 ( .S(n548), .A0(upsizer_gcm_data[107]), .A1(cmdfifo_gcm_cmd[206]), .Z(n741));
Q_MX03 U1929 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[334]), .A1(cmdfifo_gcm_cmd[462]), .A2(cmdfifo_gcm_cmd[590]), .Z(n742));
Q_MX02 U1930 ( .S(n582), .A0(n747), .A1(n743), .Z(fifo_in[107]));
Q_AN02 U1931 ( .A0(n590), .A1(n744), .Z(n743));
Q_MX02 U1932 ( .S(n547), .A0(n745), .A1(n746), .Z(n744));
Q_AN02 U1933 ( .A0(n548), .A1(gcm_tag_data_out[74]), .Z(n745));
Q_MX02 U1934 ( .S(n548), .A0(upsizer_gcm_data[106]), .A1(cmdfifo_gcm_cmd[205]), .Z(n746));
Q_MX03 U1935 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[333]), .A1(cmdfifo_gcm_cmd[461]), .A2(cmdfifo_gcm_cmd[589]), .Z(n747));
Q_MX02 U1936 ( .S(n582), .A0(n752), .A1(n748), .Z(fifo_in[106]));
Q_AN02 U1937 ( .A0(n590), .A1(n749), .Z(n748));
Q_MX02 U1938 ( .S(n547), .A0(n750), .A1(n751), .Z(n749));
Q_AN02 U1939 ( .A0(n548), .A1(gcm_tag_data_out[73]), .Z(n750));
Q_MX02 U1940 ( .S(n548), .A0(upsizer_gcm_data[105]), .A1(cmdfifo_gcm_cmd[204]), .Z(n751));
Q_MX03 U1941 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[332]), .A1(cmdfifo_gcm_cmd[460]), .A2(cmdfifo_gcm_cmd[588]), .Z(n752));
Q_MX02 U1942 ( .S(n582), .A0(n757), .A1(n753), .Z(fifo_in[105]));
Q_AN02 U1943 ( .A0(n590), .A1(n754), .Z(n753));
Q_MX02 U1944 ( .S(n547), .A0(n755), .A1(n756), .Z(n754));
Q_AN02 U1945 ( .A0(n548), .A1(gcm_tag_data_out[72]), .Z(n755));
Q_MX02 U1946 ( .S(n548), .A0(upsizer_gcm_data[104]), .A1(cmdfifo_gcm_cmd[203]), .Z(n756));
Q_MX03 U1947 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[331]), .A1(cmdfifo_gcm_cmd[459]), .A2(cmdfifo_gcm_cmd[587]), .Z(n757));
Q_MX02 U1948 ( .S(n582), .A0(n762), .A1(n758), .Z(fifo_in[104]));
Q_AN02 U1949 ( .A0(n590), .A1(n759), .Z(n758));
Q_MX02 U1950 ( .S(n547), .A0(n760), .A1(n761), .Z(n759));
Q_AN02 U1951 ( .A0(n548), .A1(gcm_tag_data_out[71]), .Z(n760));
Q_MX02 U1952 ( .S(n548), .A0(upsizer_gcm_data[103]), .A1(cmdfifo_gcm_cmd[202]), .Z(n761));
Q_MX03 U1953 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[330]), .A1(cmdfifo_gcm_cmd[458]), .A2(cmdfifo_gcm_cmd[586]), .Z(n762));
Q_MX02 U1954 ( .S(n582), .A0(n767), .A1(n763), .Z(fifo_in[103]));
Q_AN02 U1955 ( .A0(n590), .A1(n764), .Z(n763));
Q_MX02 U1956 ( .S(n547), .A0(n765), .A1(n766), .Z(n764));
Q_AN02 U1957 ( .A0(n548), .A1(gcm_tag_data_out[70]), .Z(n765));
Q_MX02 U1958 ( .S(n548), .A0(upsizer_gcm_data[102]), .A1(cmdfifo_gcm_cmd[201]), .Z(n766));
Q_MX03 U1959 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[329]), .A1(cmdfifo_gcm_cmd[457]), .A2(cmdfifo_gcm_cmd[585]), .Z(n767));
Q_MX02 U1960 ( .S(n582), .A0(n772), .A1(n768), .Z(fifo_in[102]));
Q_AN02 U1961 ( .A0(n590), .A1(n769), .Z(n768));
Q_MX02 U1962 ( .S(n547), .A0(n770), .A1(n771), .Z(n769));
Q_AN02 U1963 ( .A0(n548), .A1(gcm_tag_data_out[69]), .Z(n770));
Q_MX02 U1964 ( .S(n548), .A0(upsizer_gcm_data[101]), .A1(cmdfifo_gcm_cmd[200]), .Z(n771));
Q_MX03 U1965 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[328]), .A1(cmdfifo_gcm_cmd[456]), .A2(cmdfifo_gcm_cmd[584]), .Z(n772));
Q_MX02 U1966 ( .S(n582), .A0(n777), .A1(n773), .Z(fifo_in[101]));
Q_AN02 U1967 ( .A0(n590), .A1(n774), .Z(n773));
Q_MX02 U1968 ( .S(n547), .A0(n775), .A1(n776), .Z(n774));
Q_AN02 U1969 ( .A0(n548), .A1(gcm_tag_data_out[68]), .Z(n775));
Q_MX02 U1970 ( .S(n548), .A0(upsizer_gcm_data[100]), .A1(cmdfifo_gcm_cmd[199]), .Z(n776));
Q_MX03 U1971 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[327]), .A1(cmdfifo_gcm_cmd[455]), .A2(cmdfifo_gcm_cmd[583]), .Z(n777));
Q_MX02 U1972 ( .S(n582), .A0(n782), .A1(n778), .Z(fifo_in[100]));
Q_AN02 U1973 ( .A0(n590), .A1(n779), .Z(n778));
Q_MX02 U1974 ( .S(n547), .A0(n780), .A1(n781), .Z(n779));
Q_AN02 U1975 ( .A0(n548), .A1(gcm_tag_data_out[67]), .Z(n780));
Q_MX02 U1976 ( .S(n548), .A0(upsizer_gcm_data[99]), .A1(cmdfifo_gcm_cmd[198]), .Z(n781));
Q_MX03 U1977 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[326]), .A1(cmdfifo_gcm_cmd[454]), .A2(cmdfifo_gcm_cmd[582]), .Z(n782));
Q_MX02 U1978 ( .S(n582), .A0(n787), .A1(n783), .Z(fifo_in[99]));
Q_AN02 U1979 ( .A0(n590), .A1(n784), .Z(n783));
Q_MX02 U1980 ( .S(n547), .A0(n785), .A1(n786), .Z(n784));
Q_AN02 U1981 ( .A0(n548), .A1(gcm_tag_data_out[66]), .Z(n785));
Q_MX02 U1982 ( .S(n548), .A0(upsizer_gcm_data[98]), .A1(cmdfifo_gcm_cmd[197]), .Z(n786));
Q_MX03 U1983 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[325]), .A1(cmdfifo_gcm_cmd[453]), .A2(cmdfifo_gcm_cmd[581]), .Z(n787));
Q_MX02 U1984 ( .S(n582), .A0(n792), .A1(n788), .Z(fifo_in[98]));
Q_AN02 U1985 ( .A0(n590), .A1(n789), .Z(n788));
Q_MX02 U1986 ( .S(n547), .A0(n790), .A1(n791), .Z(n789));
Q_AN02 U1987 ( .A0(n548), .A1(gcm_tag_data_out[65]), .Z(n790));
Q_MX02 U1988 ( .S(n548), .A0(upsizer_gcm_data[97]), .A1(cmdfifo_gcm_cmd[196]), .Z(n791));
Q_MX03 U1989 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[324]), .A1(cmdfifo_gcm_cmd[452]), .A2(cmdfifo_gcm_cmd[580]), .Z(n792));
Q_MX02 U1990 ( .S(n582), .A0(n797), .A1(n793), .Z(fifo_in[97]));
Q_AN02 U1991 ( .A0(n590), .A1(n794), .Z(n793));
Q_MX02 U1992 ( .S(n547), .A0(n795), .A1(n796), .Z(n794));
Q_AN02 U1993 ( .A0(n548), .A1(gcm_tag_data_out[64]), .Z(n795));
Q_MX02 U1994 ( .S(n548), .A0(upsizer_gcm_data[96]), .A1(cmdfifo_gcm_cmd[195]), .Z(n796));
Q_MX03 U1995 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[323]), .A1(cmdfifo_gcm_cmd[451]), .A2(cmdfifo_gcm_cmd[579]), .Z(n797));
Q_MX02 U1996 ( .S(n582), .A0(n802), .A1(n798), .Z(fifo_in[96]));
Q_AN02 U1997 ( .A0(n590), .A1(n799), .Z(n798));
Q_MX02 U1998 ( .S(n547), .A0(n800), .A1(n801), .Z(n799));
Q_AN02 U1999 ( .A0(n548), .A1(gcm_tag_data_out[63]), .Z(n800));
Q_MX02 U2000 ( .S(n548), .A0(upsizer_gcm_data[95]), .A1(cmdfifo_gcm_cmd[194]), .Z(n801));
Q_MX03 U2001 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[322]), .A1(cmdfifo_gcm_cmd[450]), .A2(cmdfifo_gcm_cmd[578]), .Z(n802));
Q_MX02 U2002 ( .S(n582), .A0(n807), .A1(n803), .Z(fifo_in[95]));
Q_AN02 U2003 ( .A0(n590), .A1(n804), .Z(n803));
Q_MX02 U2004 ( .S(n547), .A0(n805), .A1(n806), .Z(n804));
Q_AN02 U2005 ( .A0(n548), .A1(gcm_tag_data_out[62]), .Z(n805));
Q_MX02 U2006 ( .S(n548), .A0(upsizer_gcm_data[94]), .A1(cmdfifo_gcm_cmd[193]), .Z(n806));
Q_MX03 U2007 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[321]), .A1(cmdfifo_gcm_cmd[449]), .A2(cmdfifo_gcm_cmd[577]), .Z(n807));
Q_MX02 U2008 ( .S(n582), .A0(n812), .A1(n808), .Z(fifo_in[94]));
Q_AN02 U2009 ( .A0(n590), .A1(n809), .Z(n808));
Q_MX02 U2010 ( .S(n547), .A0(n810), .A1(n811), .Z(n809));
Q_AN02 U2011 ( .A0(n548), .A1(gcm_tag_data_out[61]), .Z(n810));
Q_MX02 U2012 ( .S(n548), .A0(upsizer_gcm_data[93]), .A1(cmdfifo_gcm_cmd[192]), .Z(n811));
Q_MX03 U2013 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[320]), .A1(cmdfifo_gcm_cmd[448]), .A2(cmdfifo_gcm_cmd[576]), .Z(n812));
Q_MX02 U2014 ( .S(n582), .A0(n817), .A1(n813), .Z(fifo_in[93]));
Q_AN02 U2015 ( .A0(n590), .A1(n814), .Z(n813));
Q_MX02 U2016 ( .S(n547), .A0(n815), .A1(n816), .Z(n814));
Q_AN02 U2017 ( .A0(n548), .A1(gcm_tag_data_out[60]), .Z(n815));
Q_MX02 U2018 ( .S(n548), .A0(upsizer_gcm_data[92]), .A1(cmdfifo_gcm_cmd[191]), .Z(n816));
Q_MX03 U2019 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[319]), .A1(cmdfifo_gcm_cmd[447]), .A2(cmdfifo_gcm_cmd[575]), .Z(n817));
Q_MX02 U2020 ( .S(n582), .A0(n822), .A1(n818), .Z(fifo_in[92]));
Q_AN02 U2021 ( .A0(n590), .A1(n819), .Z(n818));
Q_MX02 U2022 ( .S(n547), .A0(n820), .A1(n821), .Z(n819));
Q_AN02 U2023 ( .A0(n548), .A1(gcm_tag_data_out[59]), .Z(n820));
Q_MX02 U2024 ( .S(n548), .A0(upsizer_gcm_data[91]), .A1(cmdfifo_gcm_cmd[190]), .Z(n821));
Q_MX03 U2025 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[318]), .A1(cmdfifo_gcm_cmd[446]), .A2(cmdfifo_gcm_cmd[574]), .Z(n822));
Q_MX02 U2026 ( .S(n582), .A0(n827), .A1(n823), .Z(fifo_in[91]));
Q_AN02 U2027 ( .A0(n590), .A1(n824), .Z(n823));
Q_MX02 U2028 ( .S(n547), .A0(n825), .A1(n826), .Z(n824));
Q_AN02 U2029 ( .A0(n548), .A1(gcm_tag_data_out[58]), .Z(n825));
Q_MX02 U2030 ( .S(n548), .A0(upsizer_gcm_data[90]), .A1(cmdfifo_gcm_cmd[189]), .Z(n826));
Q_MX03 U2031 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[317]), .A1(cmdfifo_gcm_cmd[445]), .A2(cmdfifo_gcm_cmd[573]), .Z(n827));
Q_MX02 U2032 ( .S(n582), .A0(n832), .A1(n828), .Z(fifo_in[90]));
Q_AN02 U2033 ( .A0(n590), .A1(n829), .Z(n828));
Q_MX02 U2034 ( .S(n547), .A0(n830), .A1(n831), .Z(n829));
Q_AN02 U2035 ( .A0(n548), .A1(gcm_tag_data_out[57]), .Z(n830));
Q_MX02 U2036 ( .S(n548), .A0(upsizer_gcm_data[89]), .A1(cmdfifo_gcm_cmd[188]), .Z(n831));
Q_MX03 U2037 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[316]), .A1(cmdfifo_gcm_cmd[444]), .A2(cmdfifo_gcm_cmd[572]), .Z(n832));
Q_MX02 U2038 ( .S(n582), .A0(n837), .A1(n833), .Z(fifo_in[89]));
Q_AN02 U2039 ( .A0(n590), .A1(n834), .Z(n833));
Q_MX02 U2040 ( .S(n547), .A0(n835), .A1(n836), .Z(n834));
Q_AN02 U2041 ( .A0(n548), .A1(gcm_tag_data_out[56]), .Z(n835));
Q_MX02 U2042 ( .S(n548), .A0(upsizer_gcm_data[88]), .A1(cmdfifo_gcm_cmd[187]), .Z(n836));
Q_MX03 U2043 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[315]), .A1(cmdfifo_gcm_cmd[443]), .A2(cmdfifo_gcm_cmd[571]), .Z(n837));
Q_MX02 U2044 ( .S(n582), .A0(n842), .A1(n838), .Z(fifo_in[88]));
Q_AN02 U2045 ( .A0(n590), .A1(n839), .Z(n838));
Q_MX02 U2046 ( .S(n547), .A0(n840), .A1(n841), .Z(n839));
Q_AN02 U2047 ( .A0(n548), .A1(gcm_tag_data_out[55]), .Z(n840));
Q_MX02 U2048 ( .S(n548), .A0(upsizer_gcm_data[87]), .A1(cmdfifo_gcm_cmd[186]), .Z(n841));
Q_MX03 U2049 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[314]), .A1(cmdfifo_gcm_cmd[442]), .A2(cmdfifo_gcm_cmd[570]), .Z(n842));
Q_MX02 U2050 ( .S(n582), .A0(n847), .A1(n843), .Z(fifo_in[87]));
Q_AN02 U2051 ( .A0(n590), .A1(n844), .Z(n843));
Q_MX02 U2052 ( .S(n547), .A0(n845), .A1(n846), .Z(n844));
Q_AN02 U2053 ( .A0(n548), .A1(gcm_tag_data_out[54]), .Z(n845));
Q_MX02 U2054 ( .S(n548), .A0(upsizer_gcm_data[86]), .A1(cmdfifo_gcm_cmd[185]), .Z(n846));
Q_MX03 U2055 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[313]), .A1(cmdfifo_gcm_cmd[441]), .A2(cmdfifo_gcm_cmd[569]), .Z(n847));
Q_MX02 U2056 ( .S(n582), .A0(n852), .A1(n848), .Z(fifo_in[86]));
Q_AN02 U2057 ( .A0(n590), .A1(n849), .Z(n848));
Q_MX02 U2058 ( .S(n547), .A0(n850), .A1(n851), .Z(n849));
Q_AN02 U2059 ( .A0(n548), .A1(gcm_tag_data_out[53]), .Z(n850));
Q_MX02 U2060 ( .S(n548), .A0(upsizer_gcm_data[85]), .A1(cmdfifo_gcm_cmd[184]), .Z(n851));
Q_MX03 U2061 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[312]), .A1(cmdfifo_gcm_cmd[440]), .A2(cmdfifo_gcm_cmd[568]), .Z(n852));
Q_MX02 U2062 ( .S(n582), .A0(n857), .A1(n853), .Z(fifo_in[85]));
Q_AN02 U2063 ( .A0(n590), .A1(n854), .Z(n853));
Q_MX02 U2064 ( .S(n547), .A0(n855), .A1(n856), .Z(n854));
Q_AN02 U2065 ( .A0(n548), .A1(gcm_tag_data_out[52]), .Z(n855));
Q_MX02 U2066 ( .S(n548), .A0(upsizer_gcm_data[84]), .A1(cmdfifo_gcm_cmd[183]), .Z(n856));
Q_MX03 U2067 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[311]), .A1(cmdfifo_gcm_cmd[439]), .A2(cmdfifo_gcm_cmd[567]), .Z(n857));
Q_MX02 U2068 ( .S(n582), .A0(n862), .A1(n858), .Z(fifo_in[84]));
Q_AN02 U2069 ( .A0(n590), .A1(n859), .Z(n858));
Q_MX02 U2070 ( .S(n547), .A0(n860), .A1(n861), .Z(n859));
Q_AN02 U2071 ( .A0(n548), .A1(gcm_tag_data_out[51]), .Z(n860));
Q_MX02 U2072 ( .S(n548), .A0(upsizer_gcm_data[83]), .A1(cmdfifo_gcm_cmd[182]), .Z(n861));
Q_MX03 U2073 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[310]), .A1(cmdfifo_gcm_cmd[438]), .A2(cmdfifo_gcm_cmd[566]), .Z(n862));
Q_MX02 U2074 ( .S(n582), .A0(n867), .A1(n863), .Z(fifo_in[83]));
Q_AN02 U2075 ( .A0(n590), .A1(n864), .Z(n863));
Q_MX02 U2076 ( .S(n547), .A0(n865), .A1(n866), .Z(n864));
Q_AN02 U2077 ( .A0(n548), .A1(gcm_tag_data_out[50]), .Z(n865));
Q_MX02 U2078 ( .S(n548), .A0(upsizer_gcm_data[82]), .A1(cmdfifo_gcm_cmd[181]), .Z(n866));
Q_MX03 U2079 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[309]), .A1(cmdfifo_gcm_cmd[437]), .A2(cmdfifo_gcm_cmd[565]), .Z(n867));
Q_MX02 U2080 ( .S(n582), .A0(n872), .A1(n868), .Z(fifo_in[82]));
Q_AN02 U2081 ( .A0(n590), .A1(n869), .Z(n868));
Q_MX02 U2082 ( .S(n547), .A0(n870), .A1(n871), .Z(n869));
Q_AN02 U2083 ( .A0(n548), .A1(gcm_tag_data_out[49]), .Z(n870));
Q_MX02 U2084 ( .S(n548), .A0(upsizer_gcm_data[81]), .A1(cmdfifo_gcm_cmd[180]), .Z(n871));
Q_MX03 U2085 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[308]), .A1(cmdfifo_gcm_cmd[436]), .A2(cmdfifo_gcm_cmd[564]), .Z(n872));
Q_MX02 U2086 ( .S(n582), .A0(n877), .A1(n873), .Z(fifo_in[81]));
Q_AN02 U2087 ( .A0(n590), .A1(n874), .Z(n873));
Q_MX02 U2088 ( .S(n547), .A0(n875), .A1(n876), .Z(n874));
Q_AN02 U2089 ( .A0(n548), .A1(gcm_tag_data_out[48]), .Z(n875));
Q_MX02 U2090 ( .S(n548), .A0(upsizer_gcm_data[80]), .A1(cmdfifo_gcm_cmd[179]), .Z(n876));
Q_MX03 U2091 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[307]), .A1(cmdfifo_gcm_cmd[435]), .A2(cmdfifo_gcm_cmd[563]), .Z(n877));
Q_MX02 U2092 ( .S(n582), .A0(n882), .A1(n878), .Z(fifo_in[80]));
Q_AN02 U2093 ( .A0(n590), .A1(n879), .Z(n878));
Q_MX02 U2094 ( .S(n547), .A0(n880), .A1(n881), .Z(n879));
Q_AN02 U2095 ( .A0(n548), .A1(gcm_tag_data_out[47]), .Z(n880));
Q_MX02 U2096 ( .S(n548), .A0(upsizer_gcm_data[79]), .A1(cmdfifo_gcm_cmd[178]), .Z(n881));
Q_MX03 U2097 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[306]), .A1(cmdfifo_gcm_cmd[434]), .A2(cmdfifo_gcm_cmd[562]), .Z(n882));
Q_MX02 U2098 ( .S(n582), .A0(n887), .A1(n883), .Z(fifo_in[79]));
Q_AN02 U2099 ( .A0(n590), .A1(n884), .Z(n883));
Q_MX02 U2100 ( .S(n547), .A0(n885), .A1(n886), .Z(n884));
Q_AN02 U2101 ( .A0(n548), .A1(gcm_tag_data_out[46]), .Z(n885));
Q_MX02 U2102 ( .S(n548), .A0(upsizer_gcm_data[78]), .A1(cmdfifo_gcm_cmd[177]), .Z(n886));
Q_MX03 U2103 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[305]), .A1(cmdfifo_gcm_cmd[433]), .A2(cmdfifo_gcm_cmd[561]), .Z(n887));
Q_MX02 U2104 ( .S(n582), .A0(n892), .A1(n888), .Z(fifo_in[78]));
Q_AN02 U2105 ( .A0(n590), .A1(n889), .Z(n888));
Q_MX02 U2106 ( .S(n547), .A0(n890), .A1(n891), .Z(n889));
Q_AN02 U2107 ( .A0(n548), .A1(gcm_tag_data_out[45]), .Z(n890));
Q_MX02 U2108 ( .S(n548), .A0(upsizer_gcm_data[77]), .A1(cmdfifo_gcm_cmd[176]), .Z(n891));
Q_MX03 U2109 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[304]), .A1(cmdfifo_gcm_cmd[432]), .A2(cmdfifo_gcm_cmd[560]), .Z(n892));
Q_MX02 U2110 ( .S(n582), .A0(n897), .A1(n893), .Z(fifo_in[77]));
Q_AN02 U2111 ( .A0(n590), .A1(n894), .Z(n893));
Q_MX02 U2112 ( .S(n547), .A0(n895), .A1(n896), .Z(n894));
Q_AN02 U2113 ( .A0(n548), .A1(gcm_tag_data_out[44]), .Z(n895));
Q_MX02 U2114 ( .S(n548), .A0(upsizer_gcm_data[76]), .A1(cmdfifo_gcm_cmd[175]), .Z(n896));
Q_MX03 U2115 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[303]), .A1(cmdfifo_gcm_cmd[431]), .A2(cmdfifo_gcm_cmd[559]), .Z(n897));
Q_MX02 U2116 ( .S(n582), .A0(n902), .A1(n898), .Z(fifo_in[76]));
Q_AN02 U2117 ( .A0(n590), .A1(n899), .Z(n898));
Q_MX02 U2118 ( .S(n547), .A0(n900), .A1(n901), .Z(n899));
Q_AN02 U2119 ( .A0(n548), .A1(gcm_tag_data_out[43]), .Z(n900));
Q_MX02 U2120 ( .S(n548), .A0(upsizer_gcm_data[75]), .A1(cmdfifo_gcm_cmd[174]), .Z(n901));
Q_MX03 U2121 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[302]), .A1(cmdfifo_gcm_cmd[430]), .A2(cmdfifo_gcm_cmd[558]), .Z(n902));
Q_MX02 U2122 ( .S(n582), .A0(n907), .A1(n903), .Z(fifo_in[75]));
Q_AN02 U2123 ( .A0(n590), .A1(n904), .Z(n903));
Q_MX02 U2124 ( .S(n547), .A0(n905), .A1(n906), .Z(n904));
Q_AN02 U2125 ( .A0(n548), .A1(gcm_tag_data_out[42]), .Z(n905));
Q_MX02 U2126 ( .S(n548), .A0(upsizer_gcm_data[74]), .A1(cmdfifo_gcm_cmd[173]), .Z(n906));
Q_MX03 U2127 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[301]), .A1(cmdfifo_gcm_cmd[429]), .A2(cmdfifo_gcm_cmd[557]), .Z(n907));
Q_MX02 U2128 ( .S(n582), .A0(n912), .A1(n908), .Z(fifo_in[74]));
Q_AN02 U2129 ( .A0(n590), .A1(n909), .Z(n908));
Q_MX02 U2130 ( .S(n547), .A0(n910), .A1(n911), .Z(n909));
Q_AN02 U2131 ( .A0(n548), .A1(gcm_tag_data_out[41]), .Z(n910));
Q_MX02 U2132 ( .S(n548), .A0(upsizer_gcm_data[73]), .A1(cmdfifo_gcm_cmd[172]), .Z(n911));
Q_MX03 U2133 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[300]), .A1(cmdfifo_gcm_cmd[428]), .A2(cmdfifo_gcm_cmd[556]), .Z(n912));
Q_MX02 U2134 ( .S(n582), .A0(n917), .A1(n913), .Z(fifo_in[73]));
Q_AN02 U2135 ( .A0(n590), .A1(n914), .Z(n913));
Q_MX02 U2136 ( .S(n547), .A0(n915), .A1(n916), .Z(n914));
Q_AN02 U2137 ( .A0(n548), .A1(gcm_tag_data_out[40]), .Z(n915));
Q_MX02 U2138 ( .S(n548), .A0(upsizer_gcm_data[72]), .A1(cmdfifo_gcm_cmd[171]), .Z(n916));
Q_MX03 U2139 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[299]), .A1(cmdfifo_gcm_cmd[427]), .A2(cmdfifo_gcm_cmd[555]), .Z(n917));
Q_MX02 U2140 ( .S(n582), .A0(n922), .A1(n918), .Z(fifo_in[72]));
Q_AN02 U2141 ( .A0(n590), .A1(n919), .Z(n918));
Q_MX02 U2142 ( .S(n547), .A0(n920), .A1(n921), .Z(n919));
Q_AN02 U2143 ( .A0(n548), .A1(gcm_tag_data_out[39]), .Z(n920));
Q_MX02 U2144 ( .S(n548), .A0(upsizer_gcm_data[71]), .A1(cmdfifo_gcm_cmd[170]), .Z(n921));
Q_MX03 U2145 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[298]), .A1(cmdfifo_gcm_cmd[426]), .A2(cmdfifo_gcm_cmd[554]), .Z(n922));
Q_MX02 U2146 ( .S(n582), .A0(n927), .A1(n923), .Z(fifo_in[71]));
Q_AN02 U2147 ( .A0(n590), .A1(n924), .Z(n923));
Q_MX02 U2148 ( .S(n547), .A0(n925), .A1(n926), .Z(n924));
Q_AN02 U2149 ( .A0(n548), .A1(gcm_tag_data_out[38]), .Z(n925));
Q_MX02 U2150 ( .S(n548), .A0(upsizer_gcm_data[70]), .A1(cmdfifo_gcm_cmd[169]), .Z(n926));
Q_MX03 U2151 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[297]), .A1(cmdfifo_gcm_cmd[425]), .A2(cmdfifo_gcm_cmd[553]), .Z(n927));
Q_MX02 U2152 ( .S(n582), .A0(n932), .A1(n928), .Z(fifo_in[70]));
Q_AN02 U2153 ( .A0(n590), .A1(n929), .Z(n928));
Q_MX02 U2154 ( .S(n547), .A0(n930), .A1(n931), .Z(n929));
Q_AN02 U2155 ( .A0(n548), .A1(gcm_tag_data_out[37]), .Z(n930));
Q_MX02 U2156 ( .S(n548), .A0(upsizer_gcm_data[69]), .A1(cmdfifo_gcm_cmd[168]), .Z(n931));
Q_MX03 U2157 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[296]), .A1(cmdfifo_gcm_cmd[424]), .A2(cmdfifo_gcm_cmd[552]), .Z(n932));
Q_MX02 U2158 ( .S(n582), .A0(n937), .A1(n933), .Z(fifo_in[69]));
Q_AN02 U2159 ( .A0(n590), .A1(n934), .Z(n933));
Q_MX02 U2160 ( .S(n547), .A0(n935), .A1(n936), .Z(n934));
Q_AN02 U2161 ( .A0(n548), .A1(gcm_tag_data_out[36]), .Z(n935));
Q_MX02 U2162 ( .S(n548), .A0(upsizer_gcm_data[68]), .A1(cmdfifo_gcm_cmd[167]), .Z(n936));
Q_MX03 U2163 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[295]), .A1(cmdfifo_gcm_cmd[423]), .A2(cmdfifo_gcm_cmd[551]), .Z(n937));
Q_MX02 U2164 ( .S(n582), .A0(n942), .A1(n938), .Z(fifo_in[68]));
Q_AN02 U2165 ( .A0(n590), .A1(n939), .Z(n938));
Q_MX02 U2166 ( .S(n547), .A0(n940), .A1(n941), .Z(n939));
Q_AN02 U2167 ( .A0(n548), .A1(gcm_tag_data_out[35]), .Z(n940));
Q_MX02 U2168 ( .S(n548), .A0(upsizer_gcm_data[67]), .A1(cmdfifo_gcm_cmd[166]), .Z(n941));
Q_MX03 U2169 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[294]), .A1(cmdfifo_gcm_cmd[422]), .A2(cmdfifo_gcm_cmd[550]), .Z(n942));
Q_MX02 U2170 ( .S(n582), .A0(n947), .A1(n943), .Z(fifo_in[67]));
Q_AN02 U2171 ( .A0(n590), .A1(n944), .Z(n943));
Q_MX02 U2172 ( .S(n547), .A0(n945), .A1(n946), .Z(n944));
Q_AN02 U2173 ( .A0(n548), .A1(gcm_tag_data_out[34]), .Z(n945));
Q_MX02 U2174 ( .S(n548), .A0(upsizer_gcm_data[66]), .A1(cmdfifo_gcm_cmd[165]), .Z(n946));
Q_MX03 U2175 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[293]), .A1(cmdfifo_gcm_cmd[421]), .A2(cmdfifo_gcm_cmd[549]), .Z(n947));
Q_MX02 U2176 ( .S(n582), .A0(n952), .A1(n948), .Z(fifo_in[66]));
Q_AN02 U2177 ( .A0(n590), .A1(n949), .Z(n948));
Q_MX02 U2178 ( .S(n547), .A0(n950), .A1(n951), .Z(n949));
Q_AN02 U2179 ( .A0(n548), .A1(gcm_tag_data_out[33]), .Z(n950));
Q_MX02 U2180 ( .S(n548), .A0(upsizer_gcm_data[65]), .A1(cmdfifo_gcm_cmd[164]), .Z(n951));
Q_MX03 U2181 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[292]), .A1(cmdfifo_gcm_cmd[420]), .A2(cmdfifo_gcm_cmd[548]), .Z(n952));
Q_MX02 U2182 ( .S(n582), .A0(n957), .A1(n953), .Z(fifo_in[65]));
Q_AN02 U2183 ( .A0(n590), .A1(n954), .Z(n953));
Q_MX02 U2184 ( .S(n547), .A0(n955), .A1(n956), .Z(n954));
Q_AN02 U2185 ( .A0(n548), .A1(gcm_tag_data_out[32]), .Z(n955));
Q_MX02 U2186 ( .S(n548), .A0(upsizer_gcm_data[64]), .A1(cmdfifo_gcm_cmd[163]), .Z(n956));
Q_MX03 U2187 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[291]), .A1(cmdfifo_gcm_cmd[419]), .A2(cmdfifo_gcm_cmd[547]), .Z(n957));
Q_MX02 U2188 ( .S(n582), .A0(n962), .A1(n958), .Z(fifo_in[64]));
Q_AN02 U2189 ( .A0(n590), .A1(n959), .Z(n958));
Q_MX02 U2190 ( .S(n547), .A0(n960), .A1(n961), .Z(n959));
Q_AN02 U2191 ( .A0(n548), .A1(gcm_tag_data_out[31]), .Z(n960));
Q_MX02 U2192 ( .S(n548), .A0(upsizer_gcm_data[63]), .A1(cmdfifo_gcm_cmd[162]), .Z(n961));
Q_MX03 U2193 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[290]), .A1(cmdfifo_gcm_cmd[418]), .A2(cmdfifo_gcm_cmd[546]), .Z(n962));
Q_MX02 U2194 ( .S(n582), .A0(n967), .A1(n963), .Z(fifo_in[63]));
Q_AN02 U2195 ( .A0(n590), .A1(n964), .Z(n963));
Q_MX02 U2196 ( .S(n547), .A0(n965), .A1(n966), .Z(n964));
Q_AN02 U2197 ( .A0(n548), .A1(gcm_tag_data_out[30]), .Z(n965));
Q_MX02 U2198 ( .S(n548), .A0(upsizer_gcm_data[62]), .A1(cmdfifo_gcm_cmd[161]), .Z(n966));
Q_MX03 U2199 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[289]), .A1(cmdfifo_gcm_cmd[417]), .A2(cmdfifo_gcm_cmd[545]), .Z(n967));
Q_MX02 U2200 ( .S(n582), .A0(n972), .A1(n968), .Z(fifo_in[62]));
Q_AN02 U2201 ( .A0(n590), .A1(n969), .Z(n968));
Q_MX02 U2202 ( .S(n547), .A0(n970), .A1(n971), .Z(n969));
Q_AN02 U2203 ( .A0(n548), .A1(gcm_tag_data_out[29]), .Z(n970));
Q_MX02 U2204 ( .S(n548), .A0(upsizer_gcm_data[61]), .A1(cmdfifo_gcm_cmd[160]), .Z(n971));
Q_MX03 U2205 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[288]), .A1(cmdfifo_gcm_cmd[416]), .A2(cmdfifo_gcm_cmd[544]), .Z(n972));
Q_MX02 U2206 ( .S(n582), .A0(n977), .A1(n973), .Z(fifo_in[61]));
Q_AN02 U2207 ( .A0(n590), .A1(n974), .Z(n973));
Q_MX02 U2208 ( .S(n547), .A0(n975), .A1(n976), .Z(n974));
Q_AN02 U2209 ( .A0(n548), .A1(gcm_tag_data_out[28]), .Z(n975));
Q_MX02 U2210 ( .S(n548), .A0(upsizer_gcm_data[60]), .A1(cmdfifo_gcm_cmd[159]), .Z(n976));
Q_MX03 U2211 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[287]), .A1(cmdfifo_gcm_cmd[415]), .A2(cmdfifo_gcm_cmd[543]), .Z(n977));
Q_MX02 U2212 ( .S(n582), .A0(n982), .A1(n978), .Z(fifo_in[60]));
Q_AN02 U2213 ( .A0(n590), .A1(n979), .Z(n978));
Q_MX02 U2214 ( .S(n547), .A0(n980), .A1(n981), .Z(n979));
Q_AN02 U2215 ( .A0(n548), .A1(gcm_tag_data_out[27]), .Z(n980));
Q_MX02 U2216 ( .S(n548), .A0(upsizer_gcm_data[59]), .A1(cmdfifo_gcm_cmd[158]), .Z(n981));
Q_MX03 U2217 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[286]), .A1(cmdfifo_gcm_cmd[414]), .A2(cmdfifo_gcm_cmd[542]), .Z(n982));
Q_MX02 U2218 ( .S(n582), .A0(n987), .A1(n983), .Z(fifo_in[59]));
Q_AN02 U2219 ( .A0(n590), .A1(n984), .Z(n983));
Q_MX02 U2220 ( .S(n547), .A0(n985), .A1(n986), .Z(n984));
Q_AN02 U2221 ( .A0(n548), .A1(gcm_tag_data_out[26]), .Z(n985));
Q_MX02 U2222 ( .S(n548), .A0(upsizer_gcm_data[58]), .A1(cmdfifo_gcm_cmd[157]), .Z(n986));
Q_MX03 U2223 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[285]), .A1(cmdfifo_gcm_cmd[413]), .A2(cmdfifo_gcm_cmd[541]), .Z(n987));
Q_MX02 U2224 ( .S(n582), .A0(n992), .A1(n988), .Z(fifo_in[58]));
Q_AN02 U2225 ( .A0(n590), .A1(n989), .Z(n988));
Q_MX02 U2226 ( .S(n547), .A0(n990), .A1(n991), .Z(n989));
Q_AN02 U2227 ( .A0(n548), .A1(gcm_tag_data_out[25]), .Z(n990));
Q_MX02 U2228 ( .S(n548), .A0(upsizer_gcm_data[57]), .A1(cmdfifo_gcm_cmd[156]), .Z(n991));
Q_MX03 U2229 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[284]), .A1(cmdfifo_gcm_cmd[412]), .A2(cmdfifo_gcm_cmd[540]), .Z(n992));
Q_MX02 U2230 ( .S(n582), .A0(n997), .A1(n993), .Z(fifo_in[57]));
Q_AN02 U2231 ( .A0(n590), .A1(n994), .Z(n993));
Q_MX02 U2232 ( .S(n547), .A0(n995), .A1(n996), .Z(n994));
Q_AN02 U2233 ( .A0(n548), .A1(gcm_tag_data_out[24]), .Z(n995));
Q_MX02 U2234 ( .S(n548), .A0(upsizer_gcm_data[56]), .A1(cmdfifo_gcm_cmd[155]), .Z(n996));
Q_MX03 U2235 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[283]), .A1(cmdfifo_gcm_cmd[411]), .A2(cmdfifo_gcm_cmd[539]), .Z(n997));
Q_MX02 U2236 ( .S(n582), .A0(n1002), .A1(n998), .Z(fifo_in[56]));
Q_AN02 U2237 ( .A0(n590), .A1(n999), .Z(n998));
Q_MX02 U2238 ( .S(n547), .A0(n1000), .A1(n1001), .Z(n999));
Q_AN02 U2239 ( .A0(n548), .A1(gcm_tag_data_out[23]), .Z(n1000));
Q_MX02 U2240 ( .S(n548), .A0(upsizer_gcm_data[55]), .A1(cmdfifo_gcm_cmd[154]), .Z(n1001));
Q_MX03 U2241 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[282]), .A1(cmdfifo_gcm_cmd[410]), .A2(cmdfifo_gcm_cmd[538]), .Z(n1002));
Q_MX02 U2242 ( .S(n582), .A0(n1007), .A1(n1003), .Z(fifo_in[55]));
Q_AN02 U2243 ( .A0(n590), .A1(n1004), .Z(n1003));
Q_MX02 U2244 ( .S(n547), .A0(n1005), .A1(n1006), .Z(n1004));
Q_AN02 U2245 ( .A0(n548), .A1(gcm_tag_data_out[22]), .Z(n1005));
Q_MX02 U2246 ( .S(n548), .A0(upsizer_gcm_data[54]), .A1(cmdfifo_gcm_cmd[153]), .Z(n1006));
Q_MX03 U2247 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[281]), .A1(cmdfifo_gcm_cmd[409]), .A2(cmdfifo_gcm_cmd[537]), .Z(n1007));
Q_MX02 U2248 ( .S(n582), .A0(n1012), .A1(n1008), .Z(fifo_in[54]));
Q_AN02 U2249 ( .A0(n590), .A1(n1009), .Z(n1008));
Q_MX02 U2250 ( .S(n547), .A0(n1010), .A1(n1011), .Z(n1009));
Q_AN02 U2251 ( .A0(n548), .A1(gcm_tag_data_out[21]), .Z(n1010));
Q_MX02 U2252 ( .S(n548), .A0(upsizer_gcm_data[53]), .A1(cmdfifo_gcm_cmd[152]), .Z(n1011));
Q_MX03 U2253 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[280]), .A1(cmdfifo_gcm_cmd[408]), .A2(cmdfifo_gcm_cmd[536]), .Z(n1012));
Q_MX02 U2254 ( .S(n582), .A0(n1017), .A1(n1013), .Z(fifo_in[53]));
Q_AN02 U2255 ( .A0(n590), .A1(n1014), .Z(n1013));
Q_MX02 U2256 ( .S(n547), .A0(n1015), .A1(n1016), .Z(n1014));
Q_AN02 U2257 ( .A0(n548), .A1(gcm_tag_data_out[20]), .Z(n1015));
Q_MX02 U2258 ( .S(n548), .A0(upsizer_gcm_data[52]), .A1(cmdfifo_gcm_cmd[151]), .Z(n1016));
Q_MX03 U2259 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[279]), .A1(cmdfifo_gcm_cmd[407]), .A2(cmdfifo_gcm_cmd[535]), .Z(n1017));
Q_MX02 U2260 ( .S(n582), .A0(n1022), .A1(n1018), .Z(fifo_in[52]));
Q_AN02 U2261 ( .A0(n590), .A1(n1019), .Z(n1018));
Q_MX02 U2262 ( .S(n547), .A0(n1020), .A1(n1021), .Z(n1019));
Q_AN02 U2263 ( .A0(n548), .A1(gcm_tag_data_out[19]), .Z(n1020));
Q_MX02 U2264 ( .S(n548), .A0(upsizer_gcm_data[51]), .A1(cmdfifo_gcm_cmd[150]), .Z(n1021));
Q_MX03 U2265 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[278]), .A1(cmdfifo_gcm_cmd[406]), .A2(cmdfifo_gcm_cmd[534]), .Z(n1022));
Q_MX02 U2266 ( .S(n582), .A0(n1027), .A1(n1023), .Z(fifo_in[51]));
Q_AN02 U2267 ( .A0(n590), .A1(n1024), .Z(n1023));
Q_MX02 U2268 ( .S(n547), .A0(n1025), .A1(n1026), .Z(n1024));
Q_AN02 U2269 ( .A0(n548), .A1(gcm_tag_data_out[18]), .Z(n1025));
Q_MX02 U2270 ( .S(n548), .A0(upsizer_gcm_data[50]), .A1(cmdfifo_gcm_cmd[149]), .Z(n1026));
Q_MX03 U2271 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[277]), .A1(cmdfifo_gcm_cmd[405]), .A2(cmdfifo_gcm_cmd[533]), .Z(n1027));
Q_MX02 U2272 ( .S(n582), .A0(n1032), .A1(n1028), .Z(fifo_in[50]));
Q_AN02 U2273 ( .A0(n590), .A1(n1029), .Z(n1028));
Q_MX02 U2274 ( .S(n547), .A0(n1030), .A1(n1031), .Z(n1029));
Q_AN02 U2275 ( .A0(n548), .A1(gcm_tag_data_out[17]), .Z(n1030));
Q_MX02 U2276 ( .S(n548), .A0(upsizer_gcm_data[49]), .A1(cmdfifo_gcm_cmd[148]), .Z(n1031));
Q_MX03 U2277 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[276]), .A1(cmdfifo_gcm_cmd[404]), .A2(cmdfifo_gcm_cmd[532]), .Z(n1032));
Q_MX02 U2278 ( .S(n582), .A0(n1037), .A1(n1033), .Z(fifo_in[49]));
Q_AN02 U2279 ( .A0(n590), .A1(n1034), .Z(n1033));
Q_MX02 U2280 ( .S(n547), .A0(n1035), .A1(n1036), .Z(n1034));
Q_AN02 U2281 ( .A0(n548), .A1(gcm_tag_data_out[16]), .Z(n1035));
Q_MX02 U2282 ( .S(n548), .A0(upsizer_gcm_data[48]), .A1(cmdfifo_gcm_cmd[147]), .Z(n1036));
Q_MX03 U2283 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[275]), .A1(cmdfifo_gcm_cmd[403]), .A2(cmdfifo_gcm_cmd[531]), .Z(n1037));
Q_MX02 U2284 ( .S(n582), .A0(n1042), .A1(n1038), .Z(fifo_in[48]));
Q_AN02 U2285 ( .A0(n590), .A1(n1039), .Z(n1038));
Q_MX02 U2286 ( .S(n547), .A0(n1040), .A1(n1041), .Z(n1039));
Q_AN02 U2287 ( .A0(n548), .A1(gcm_tag_data_out[15]), .Z(n1040));
Q_MX02 U2288 ( .S(n548), .A0(upsizer_gcm_data[47]), .A1(cmdfifo_gcm_cmd[146]), .Z(n1041));
Q_MX03 U2289 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[274]), .A1(cmdfifo_gcm_cmd[402]), .A2(cmdfifo_gcm_cmd[530]), .Z(n1042));
Q_MX02 U2290 ( .S(n582), .A0(n1047), .A1(n1043), .Z(fifo_in[47]));
Q_AN02 U2291 ( .A0(n590), .A1(n1044), .Z(n1043));
Q_MX02 U2292 ( .S(n547), .A0(n1045), .A1(n1046), .Z(n1044));
Q_AN02 U2293 ( .A0(n548), .A1(gcm_tag_data_out[14]), .Z(n1045));
Q_MX02 U2294 ( .S(n548), .A0(upsizer_gcm_data[46]), .A1(cmdfifo_gcm_cmd[145]), .Z(n1046));
Q_MX03 U2295 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[273]), .A1(cmdfifo_gcm_cmd[401]), .A2(cmdfifo_gcm_cmd[529]), .Z(n1047));
Q_MX02 U2296 ( .S(n582), .A0(n1052), .A1(n1048), .Z(fifo_in[46]));
Q_AN02 U2297 ( .A0(n590), .A1(n1049), .Z(n1048));
Q_MX02 U2298 ( .S(n547), .A0(n1050), .A1(n1051), .Z(n1049));
Q_AN02 U2299 ( .A0(n548), .A1(gcm_tag_data_out[13]), .Z(n1050));
Q_MX02 U2300 ( .S(n548), .A0(upsizer_gcm_data[45]), .A1(cmdfifo_gcm_cmd[144]), .Z(n1051));
Q_MX03 U2301 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[272]), .A1(cmdfifo_gcm_cmd[400]), .A2(cmdfifo_gcm_cmd[528]), .Z(n1052));
Q_MX02 U2302 ( .S(n582), .A0(n1057), .A1(n1053), .Z(fifo_in[45]));
Q_AN02 U2303 ( .A0(n590), .A1(n1054), .Z(n1053));
Q_MX02 U2304 ( .S(n547), .A0(n1055), .A1(n1056), .Z(n1054));
Q_AN02 U2305 ( .A0(n548), .A1(gcm_tag_data_out[12]), .Z(n1055));
Q_MX02 U2306 ( .S(n548), .A0(upsizer_gcm_data[44]), .A1(cmdfifo_gcm_cmd[143]), .Z(n1056));
Q_MX03 U2307 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[271]), .A1(cmdfifo_gcm_cmd[399]), .A2(cmdfifo_gcm_cmd[527]), .Z(n1057));
Q_MX02 U2308 ( .S(n582), .A0(n1062), .A1(n1058), .Z(fifo_in[44]));
Q_AN02 U2309 ( .A0(n590), .A1(n1059), .Z(n1058));
Q_MX02 U2310 ( .S(n547), .A0(n1060), .A1(n1061), .Z(n1059));
Q_AN02 U2311 ( .A0(n548), .A1(gcm_tag_data_out[11]), .Z(n1060));
Q_MX02 U2312 ( .S(n548), .A0(upsizer_gcm_data[43]), .A1(cmdfifo_gcm_cmd[142]), .Z(n1061));
Q_MX03 U2313 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[270]), .A1(cmdfifo_gcm_cmd[398]), .A2(cmdfifo_gcm_cmd[526]), .Z(n1062));
Q_MX02 U2314 ( .S(n582), .A0(n1067), .A1(n1063), .Z(fifo_in[43]));
Q_AN02 U2315 ( .A0(n590), .A1(n1064), .Z(n1063));
Q_MX02 U2316 ( .S(n547), .A0(n1065), .A1(n1066), .Z(n1064));
Q_AN02 U2317 ( .A0(n548), .A1(gcm_tag_data_out[10]), .Z(n1065));
Q_MX02 U2318 ( .S(n548), .A0(upsizer_gcm_data[42]), .A1(cmdfifo_gcm_cmd[141]), .Z(n1066));
Q_MX03 U2319 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[269]), .A1(cmdfifo_gcm_cmd[397]), .A2(cmdfifo_gcm_cmd[525]), .Z(n1067));
Q_MX02 U2320 ( .S(n582), .A0(n1072), .A1(n1068), .Z(fifo_in[42]));
Q_AN02 U2321 ( .A0(n590), .A1(n1069), .Z(n1068));
Q_MX02 U2322 ( .S(n547), .A0(n1070), .A1(n1071), .Z(n1069));
Q_AN02 U2323 ( .A0(n548), .A1(gcm_tag_data_out[9]), .Z(n1070));
Q_MX02 U2324 ( .S(n548), .A0(upsizer_gcm_data[41]), .A1(cmdfifo_gcm_cmd[140]), .Z(n1071));
Q_MX03 U2325 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[268]), .A1(cmdfifo_gcm_cmd[396]), .A2(cmdfifo_gcm_cmd[524]), .Z(n1072));
Q_MX02 U2326 ( .S(n582), .A0(n1077), .A1(n1073), .Z(fifo_in[41]));
Q_AN02 U2327 ( .A0(n590), .A1(n1074), .Z(n1073));
Q_MX02 U2328 ( .S(n547), .A0(n1075), .A1(n1076), .Z(n1074));
Q_AN02 U2329 ( .A0(n548), .A1(gcm_tag_data_out[8]), .Z(n1075));
Q_MX02 U2330 ( .S(n548), .A0(upsizer_gcm_data[40]), .A1(cmdfifo_gcm_cmd[139]), .Z(n1076));
Q_MX03 U2331 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[267]), .A1(cmdfifo_gcm_cmd[395]), .A2(cmdfifo_gcm_cmd[523]), .Z(n1077));
Q_MX02 U2332 ( .S(n582), .A0(n1082), .A1(n1078), .Z(fifo_in[40]));
Q_AN02 U2333 ( .A0(n590), .A1(n1079), .Z(n1078));
Q_MX02 U2334 ( .S(n547), .A0(n1080), .A1(n1081), .Z(n1079));
Q_AN02 U2335 ( .A0(n548), .A1(gcm_tag_data_out[7]), .Z(n1080));
Q_MX02 U2336 ( .S(n548), .A0(upsizer_gcm_data[39]), .A1(cmdfifo_gcm_cmd[138]), .Z(n1081));
Q_MX03 U2337 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[266]), .A1(cmdfifo_gcm_cmd[394]), .A2(cmdfifo_gcm_cmd[522]), .Z(n1082));
Q_MX02 U2338 ( .S(n582), .A0(n1087), .A1(n1083), .Z(fifo_in[39]));
Q_AN02 U2339 ( .A0(n590), .A1(n1084), .Z(n1083));
Q_MX02 U2340 ( .S(n547), .A0(n1085), .A1(n1086), .Z(n1084));
Q_AN02 U2341 ( .A0(n548), .A1(gcm_tag_data_out[6]), .Z(n1085));
Q_MX02 U2342 ( .S(n548), .A0(upsizer_gcm_data[38]), .A1(cmdfifo_gcm_cmd[137]), .Z(n1086));
Q_MX03 U2343 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[265]), .A1(cmdfifo_gcm_cmd[393]), .A2(cmdfifo_gcm_cmd[521]), .Z(n1087));
Q_MX02 U2344 ( .S(n582), .A0(n1092), .A1(n1088), .Z(fifo_in[38]));
Q_AN02 U2345 ( .A0(n590), .A1(n1089), .Z(n1088));
Q_MX02 U2346 ( .S(n547), .A0(n1090), .A1(n1091), .Z(n1089));
Q_AN02 U2347 ( .A0(n548), .A1(gcm_tag_data_out[5]), .Z(n1090));
Q_MX02 U2348 ( .S(n548), .A0(upsizer_gcm_data[37]), .A1(cmdfifo_gcm_cmd[136]), .Z(n1091));
Q_MX03 U2349 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[264]), .A1(cmdfifo_gcm_cmd[392]), .A2(cmdfifo_gcm_cmd[520]), .Z(n1092));
Q_MX02 U2350 ( .S(n582), .A0(n1097), .A1(n1093), .Z(fifo_in[37]));
Q_AN02 U2351 ( .A0(n590), .A1(n1094), .Z(n1093));
Q_MX02 U2352 ( .S(n547), .A0(n1095), .A1(n1096), .Z(n1094));
Q_AN02 U2353 ( .A0(n548), .A1(gcm_tag_data_out[4]), .Z(n1095));
Q_MX02 U2354 ( .S(n548), .A0(upsizer_gcm_data[36]), .A1(cmdfifo_gcm_cmd[135]), .Z(n1096));
Q_MX03 U2355 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[263]), .A1(cmdfifo_gcm_cmd[391]), .A2(cmdfifo_gcm_cmd[519]), .Z(n1097));
Q_MX02 U2356 ( .S(n582), .A0(n1102), .A1(n1098), .Z(fifo_in[36]));
Q_AN02 U2357 ( .A0(n590), .A1(n1099), .Z(n1098));
Q_MX02 U2358 ( .S(n547), .A0(n1100), .A1(n1101), .Z(n1099));
Q_AN02 U2359 ( .A0(n548), .A1(gcm_tag_data_out[3]), .Z(n1100));
Q_MX02 U2360 ( .S(n548), .A0(upsizer_gcm_data[35]), .A1(cmdfifo_gcm_cmd[134]), .Z(n1101));
Q_MX03 U2361 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[262]), .A1(cmdfifo_gcm_cmd[390]), .A2(cmdfifo_gcm_cmd[518]), .Z(n1102));
Q_MX02 U2362 ( .S(n582), .A0(n1107), .A1(n1103), .Z(fifo_in[35]));
Q_AN02 U2363 ( .A0(n590), .A1(n1104), .Z(n1103));
Q_MX02 U2364 ( .S(n547), .A0(n1105), .A1(n1106), .Z(n1104));
Q_AN02 U2365 ( .A0(n548), .A1(gcm_tag_data_out[2]), .Z(n1105));
Q_MX02 U2366 ( .S(n548), .A0(upsizer_gcm_data[34]), .A1(cmdfifo_gcm_cmd[133]), .Z(n1106));
Q_MX03 U2367 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[261]), .A1(cmdfifo_gcm_cmd[389]), .A2(cmdfifo_gcm_cmd[517]), .Z(n1107));
Q_MX02 U2368 ( .S(n582), .A0(n1112), .A1(n1108), .Z(fifo_in[34]));
Q_AN02 U2369 ( .A0(n590), .A1(n1109), .Z(n1108));
Q_MX02 U2370 ( .S(n547), .A0(n1110), .A1(n1111), .Z(n1109));
Q_AN02 U2371 ( .A0(n548), .A1(gcm_tag_data_out[1]), .Z(n1110));
Q_MX02 U2372 ( .S(n548), .A0(upsizer_gcm_data[33]), .A1(cmdfifo_gcm_cmd[132]), .Z(n1111));
Q_MX03 U2373 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[260]), .A1(cmdfifo_gcm_cmd[388]), .A2(cmdfifo_gcm_cmd[516]), .Z(n1112));
Q_MX02 U2374 ( .S(n582), .A0(n1117), .A1(n1113), .Z(fifo_in[33]));
Q_AN02 U2375 ( .A0(n590), .A1(n1114), .Z(n1113));
Q_MX02 U2376 ( .S(n547), .A0(n1115), .A1(n1116), .Z(n1114));
Q_AN02 U2377 ( .A0(n548), .A1(gcm_tag_data_out[0]), .Z(n1115));
Q_MX02 U2378 ( .S(n548), .A0(upsizer_gcm_data[32]), .A1(cmdfifo_gcm_cmd[131]), .Z(n1116));
Q_MX03 U2379 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[259]), .A1(cmdfifo_gcm_cmd[387]), .A2(cmdfifo_gcm_cmd[515]), .Z(n1117));
Q_MX02 U2380 ( .S(n582), .A0(n1120), .A1(n1118), .Z(fifo_in[32]));
Q_AN03 U2381 ( .A0(n547), .A1(n1119), .A2(n590), .Z(n1118));
Q_MX02 U2382 ( .S(n548), .A0(upsizer_gcm_data[31]), .A1(cmdfifo_gcm_cmd[130]), .Z(n1119));
Q_MX03 U2383 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[258]), .A1(cmdfifo_gcm_cmd[386]), .A2(cmdfifo_gcm_cmd[514]), .Z(n1120));
Q_MX02 U2384 ( .S(n582), .A0(n1123), .A1(n1121), .Z(fifo_in[31]));
Q_AN03 U2385 ( .A0(n547), .A1(n1122), .A2(n590), .Z(n1121));
Q_MX02 U2386 ( .S(n548), .A0(upsizer_gcm_data[30]), .A1(cmdfifo_gcm_cmd[129]), .Z(n1122));
Q_MX03 U2387 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[257]), .A1(cmdfifo_gcm_cmd[385]), .A2(cmdfifo_gcm_cmd[513]), .Z(n1123));
Q_MX02 U2388 ( .S(n582), .A0(n1126), .A1(n1124), .Z(fifo_in[30]));
Q_AN03 U2389 ( .A0(n547), .A1(n1125), .A2(n590), .Z(n1124));
Q_MX02 U2390 ( .S(n548), .A0(upsizer_gcm_data[29]), .A1(cmdfifo_gcm_cmd[128]), .Z(n1125));
Q_MX03 U2391 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[256]), .A1(cmdfifo_gcm_cmd[384]), .A2(cmdfifo_gcm_cmd[512]), .Z(n1126));
Q_MX02 U2392 ( .S(n582), .A0(n1129), .A1(n1127), .Z(fifo_in[29]));
Q_AN03 U2393 ( .A0(n547), .A1(n1128), .A2(n590), .Z(n1127));
Q_MX02 U2394 ( .S(n548), .A0(upsizer_gcm_data[28]), .A1(cmdfifo_gcm_cmd[127]), .Z(n1128));
Q_MX03 U2395 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[255]), .A1(cmdfifo_gcm_cmd[383]), .A2(cmdfifo_gcm_cmd[511]), .Z(n1129));
Q_MX02 U2396 ( .S(n582), .A0(n1132), .A1(n1130), .Z(fifo_in[28]));
Q_AN03 U2397 ( .A0(n547), .A1(n1131), .A2(n590), .Z(n1130));
Q_MX02 U2398 ( .S(n548), .A0(upsizer_gcm_data[27]), .A1(cmdfifo_gcm_cmd[126]), .Z(n1131));
Q_MX03 U2399 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[254]), .A1(cmdfifo_gcm_cmd[382]), .A2(cmdfifo_gcm_cmd[510]), .Z(n1132));
Q_MX02 U2400 ( .S(n582), .A0(n1135), .A1(n1133), .Z(fifo_in[27]));
Q_AN03 U2401 ( .A0(n547), .A1(n1134), .A2(n590), .Z(n1133));
Q_MX02 U2402 ( .S(n548), .A0(upsizer_gcm_data[26]), .A1(cmdfifo_gcm_cmd[125]), .Z(n1134));
Q_MX03 U2403 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[253]), .A1(cmdfifo_gcm_cmd[381]), .A2(cmdfifo_gcm_cmd[509]), .Z(n1135));
Q_MX02 U2404 ( .S(n582), .A0(n1138), .A1(n1136), .Z(fifo_in[26]));
Q_AN03 U2405 ( .A0(n547), .A1(n1137), .A2(n590), .Z(n1136));
Q_MX02 U2406 ( .S(n548), .A0(upsizer_gcm_data[25]), .A1(cmdfifo_gcm_cmd[124]), .Z(n1137));
Q_MX03 U2407 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[252]), .A1(cmdfifo_gcm_cmd[380]), .A2(cmdfifo_gcm_cmd[508]), .Z(n1138));
Q_MX02 U2408 ( .S(n582), .A0(n1141), .A1(n1139), .Z(fifo_in[25]));
Q_AN03 U2409 ( .A0(n547), .A1(n1140), .A2(n590), .Z(n1139));
Q_MX02 U2410 ( .S(n548), .A0(upsizer_gcm_data[24]), .A1(cmdfifo_gcm_cmd[123]), .Z(n1140));
Q_MX03 U2411 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[251]), .A1(cmdfifo_gcm_cmd[379]), .A2(cmdfifo_gcm_cmd[507]), .Z(n1141));
Q_MX02 U2412 ( .S(n582), .A0(n1144), .A1(n1142), .Z(fifo_in[24]));
Q_AN03 U2413 ( .A0(n547), .A1(n1143), .A2(n590), .Z(n1142));
Q_MX02 U2414 ( .S(n548), .A0(upsizer_gcm_data[23]), .A1(cmdfifo_gcm_cmd[122]), .Z(n1143));
Q_MX03 U2415 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[250]), .A1(cmdfifo_gcm_cmd[378]), .A2(cmdfifo_gcm_cmd[506]), .Z(n1144));
Q_MX02 U2416 ( .S(n582), .A0(n1147), .A1(n1145), .Z(fifo_in[23]));
Q_AN03 U2417 ( .A0(n547), .A1(n1146), .A2(n590), .Z(n1145));
Q_MX02 U2418 ( .S(n548), .A0(upsizer_gcm_data[22]), .A1(cmdfifo_gcm_cmd[121]), .Z(n1146));
Q_MX03 U2419 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[249]), .A1(cmdfifo_gcm_cmd[377]), .A2(cmdfifo_gcm_cmd[505]), .Z(n1147));
Q_MX02 U2420 ( .S(n582), .A0(n1150), .A1(n1148), .Z(fifo_in[22]));
Q_AN03 U2421 ( .A0(n547), .A1(n1149), .A2(n590), .Z(n1148));
Q_MX02 U2422 ( .S(n548), .A0(upsizer_gcm_data[21]), .A1(cmdfifo_gcm_cmd[120]), .Z(n1149));
Q_MX03 U2423 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[248]), .A1(cmdfifo_gcm_cmd[376]), .A2(cmdfifo_gcm_cmd[504]), .Z(n1150));
Q_MX02 U2424 ( .S(n582), .A0(n1153), .A1(n1151), .Z(fifo_in[21]));
Q_AN03 U2425 ( .A0(n547), .A1(n1152), .A2(n590), .Z(n1151));
Q_MX02 U2426 ( .S(n548), .A0(upsizer_gcm_data[20]), .A1(cmdfifo_gcm_cmd[119]), .Z(n1152));
Q_MX03 U2427 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[247]), .A1(cmdfifo_gcm_cmd[375]), .A2(cmdfifo_gcm_cmd[503]), .Z(n1153));
Q_MX02 U2428 ( .S(n582), .A0(n1156), .A1(n1154), .Z(fifo_in[20]));
Q_AN03 U2429 ( .A0(n547), .A1(n1155), .A2(n590), .Z(n1154));
Q_MX02 U2430 ( .S(n548), .A0(upsizer_gcm_data[19]), .A1(cmdfifo_gcm_cmd[118]), .Z(n1155));
Q_MX03 U2431 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[246]), .A1(cmdfifo_gcm_cmd[374]), .A2(cmdfifo_gcm_cmd[502]), .Z(n1156));
Q_MX02 U2432 ( .S(n582), .A0(n1159), .A1(n1157), .Z(fifo_in[19]));
Q_AN03 U2433 ( .A0(n547), .A1(n1158), .A2(n590), .Z(n1157));
Q_MX02 U2434 ( .S(n548), .A0(upsizer_gcm_data[18]), .A1(cmdfifo_gcm_cmd[117]), .Z(n1158));
Q_MX03 U2435 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[245]), .A1(cmdfifo_gcm_cmd[373]), .A2(cmdfifo_gcm_cmd[501]), .Z(n1159));
Q_MX02 U2436 ( .S(n582), .A0(n1162), .A1(n1160), .Z(fifo_in[18]));
Q_AN03 U2437 ( .A0(n547), .A1(n1161), .A2(n590), .Z(n1160));
Q_MX02 U2438 ( .S(n548), .A0(upsizer_gcm_data[17]), .A1(cmdfifo_gcm_cmd[116]), .Z(n1161));
Q_MX03 U2439 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[244]), .A1(cmdfifo_gcm_cmd[372]), .A2(cmdfifo_gcm_cmd[500]), .Z(n1162));
Q_MX02 U2440 ( .S(n582), .A0(n1165), .A1(n1163), .Z(fifo_in[17]));
Q_AN03 U2441 ( .A0(n547), .A1(n1164), .A2(n590), .Z(n1163));
Q_MX02 U2442 ( .S(n548), .A0(upsizer_gcm_data[16]), .A1(cmdfifo_gcm_cmd[115]), .Z(n1164));
Q_MX03 U2443 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[243]), .A1(cmdfifo_gcm_cmd[371]), .A2(cmdfifo_gcm_cmd[499]), .Z(n1165));
Q_MX02 U2444 ( .S(n582), .A0(n1168), .A1(n1166), .Z(fifo_in[16]));
Q_AN03 U2445 ( .A0(n547), .A1(n1167), .A2(n590), .Z(n1166));
Q_MX02 U2446 ( .S(n548), .A0(upsizer_gcm_data[15]), .A1(cmdfifo_gcm_cmd[114]), .Z(n1167));
Q_MX03 U2447 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[242]), .A1(cmdfifo_gcm_cmd[370]), .A2(cmdfifo_gcm_cmd[498]), .Z(n1168));
Q_MX02 U2448 ( .S(n582), .A0(n1171), .A1(n1169), .Z(fifo_in[15]));
Q_AN03 U2449 ( .A0(n547), .A1(n1170), .A2(n590), .Z(n1169));
Q_MX02 U2450 ( .S(n548), .A0(upsizer_gcm_data[14]), .A1(cmdfifo_gcm_cmd[113]), .Z(n1170));
Q_MX03 U2451 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[241]), .A1(cmdfifo_gcm_cmd[369]), .A2(cmdfifo_gcm_cmd[497]), .Z(n1171));
Q_MX02 U2452 ( .S(n582), .A0(n1174), .A1(n1172), .Z(fifo_in[14]));
Q_AN03 U2453 ( .A0(n547), .A1(n1173), .A2(n590), .Z(n1172));
Q_MX02 U2454 ( .S(n548), .A0(upsizer_gcm_data[13]), .A1(cmdfifo_gcm_cmd[112]), .Z(n1173));
Q_MX03 U2455 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[240]), .A1(cmdfifo_gcm_cmd[368]), .A2(cmdfifo_gcm_cmd[496]), .Z(n1174));
Q_MX02 U2456 ( .S(n582), .A0(n1177), .A1(n1175), .Z(fifo_in[13]));
Q_AN03 U2457 ( .A0(n547), .A1(n1176), .A2(n590), .Z(n1175));
Q_MX02 U2458 ( .S(n548), .A0(upsizer_gcm_data[12]), .A1(cmdfifo_gcm_cmd[111]), .Z(n1176));
Q_MX03 U2459 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[239]), .A1(cmdfifo_gcm_cmd[367]), .A2(cmdfifo_gcm_cmd[495]), .Z(n1177));
Q_MX02 U2460 ( .S(n582), .A0(n1180), .A1(n1178), .Z(fifo_in[12]));
Q_AN03 U2461 ( .A0(n547), .A1(n1179), .A2(n590), .Z(n1178));
Q_MX02 U2462 ( .S(n548), .A0(upsizer_gcm_data[11]), .A1(cmdfifo_gcm_cmd[110]), .Z(n1179));
Q_MX03 U2463 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[238]), .A1(cmdfifo_gcm_cmd[366]), .A2(cmdfifo_gcm_cmd[494]), .Z(n1180));
Q_MX02 U2464 ( .S(n582), .A0(n1183), .A1(n1181), .Z(fifo_in[11]));
Q_AN03 U2465 ( .A0(n547), .A1(n1182), .A2(n590), .Z(n1181));
Q_MX02 U2466 ( .S(n548), .A0(upsizer_gcm_data[10]), .A1(cmdfifo_gcm_cmd[109]), .Z(n1182));
Q_MX03 U2467 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[237]), .A1(cmdfifo_gcm_cmd[365]), .A2(cmdfifo_gcm_cmd[493]), .Z(n1183));
Q_MX03 U2468 ( .S0(n590), .S1(n546), .A0(n1184), .A1(n1185), .A2(n1187), .Z(fifo_in[10]));
Q_INV U2469 ( .A(n547), .Z(n1184));
Q_AN02 U2470 ( .A0(n547), .A1(n1186), .Z(n1185));
Q_MX02 U2471 ( .S(n548), .A0(upsizer_gcm_data[9]), .A1(cmdfifo_gcm_cmd[108]), .Z(n1186));
Q_MX03 U2472 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[236]), .A1(cmdfifo_gcm_cmd[364]), .A2(cmdfifo_gcm_cmd[492]), .Z(n1187));
Q_MX03 U2473 ( .S0(n590), .S1(n546), .A0(n1188), .A1(n1189), .A2(n1191), .Z(fifo_in[9]));
Q_INV U2474 ( .A(n548), .Z(n1188));
Q_AN02 U2475 ( .A0(n547), .A1(n1190), .Z(n1189));
Q_MX02 U2476 ( .S(n548), .A0(upsizer_gcm_data[8]), .A1(cmdfifo_gcm_cmd[107]), .Z(n1190));
Q_MX03 U2477 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[235]), .A1(cmdfifo_gcm_cmd[363]), .A2(cmdfifo_gcm_cmd[491]), .Z(n1191));
Q_MX02 U2478 ( .S(n582), .A0(n1194), .A1(n1192), .Z(fifo_in[8]));
Q_AN03 U2479 ( .A0(n547), .A1(n1193), .A2(n590), .Z(n1192));
Q_MX02 U2480 ( .S(n548), .A0(upsizer_gcm_data[7]), .A1(cmdfifo_gcm_cmd[106]), .Z(n1193));
Q_MX03 U2481 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[234]), .A1(cmdfifo_gcm_cmd[362]), .A2(cmdfifo_gcm_cmd[490]), .Z(n1194));
Q_MX02 U2482 ( .S(n582), .A0(n1197), .A1(n1195), .Z(fifo_in[7]));
Q_AN03 U2483 ( .A0(n547), .A1(n1196), .A2(n590), .Z(n1195));
Q_MX02 U2484 ( .S(n548), .A0(upsizer_gcm_data[6]), .A1(cmdfifo_gcm_cmd[105]), .Z(n1196));
Q_MX03 U2485 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[233]), .A1(cmdfifo_gcm_cmd[361]), .A2(cmdfifo_gcm_cmd[489]), .Z(n1197));
Q_MX02 U2486 ( .S(n582), .A0(n1200), .A1(n1198), .Z(fifo_in[6]));
Q_AN03 U2487 ( .A0(n547), .A1(n1199), .A2(n590), .Z(n1198));
Q_MX02 U2488 ( .S(n548), .A0(upsizer_gcm_data[5]), .A1(cmdfifo_gcm_cmd[104]), .Z(n1199));
Q_MX03 U2489 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[232]), .A1(cmdfifo_gcm_cmd[360]), .A2(cmdfifo_gcm_cmd[488]), .Z(n1200));
Q_MX02 U2490 ( .S(n582), .A0(n1203), .A1(n1201), .Z(fifo_in[5]));
Q_AN03 U2491 ( .A0(n547), .A1(n1202), .A2(n590), .Z(n1201));
Q_MX02 U2492 ( .S(n548), .A0(upsizer_gcm_data[4]), .A1(cmdfifo_gcm_cmd[103]), .Z(n1202));
Q_MX03 U2493 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[231]), .A1(cmdfifo_gcm_cmd[359]), .A2(cmdfifo_gcm_cmd[487]), .Z(n1203));
Q_MX02 U2494 ( .S(n582), .A0(n1206), .A1(n1204), .Z(fifo_in[4]));
Q_AN03 U2495 ( .A0(n547), .A1(n1205), .A2(n590), .Z(n1204));
Q_MX02 U2496 ( .S(n548), .A0(upsizer_gcm_data[3]), .A1(cmdfifo_gcm_cmd[102]), .Z(n1205));
Q_MX03 U2497 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[230]), .A1(cmdfifo_gcm_cmd[358]), .A2(cmdfifo_gcm_cmd[486]), .Z(n1206));
Q_MX02 U2498 ( .S(n582), .A0(n1209), .A1(n1207), .Z(fifo_in[3]));
Q_AN03 U2499 ( .A0(n547), .A1(n1208), .A2(n590), .Z(n1207));
Q_MX02 U2500 ( .S(n548), .A0(upsizer_gcm_data[2]), .A1(cmdfifo_gcm_cmd[101]), .Z(n1208));
Q_MX03 U2501 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[229]), .A1(cmdfifo_gcm_cmd[357]), .A2(cmdfifo_gcm_cmd[485]), .Z(n1209));
Q_MX02 U2502 ( .S(n582), .A0(n1212), .A1(n1210), .Z(fifo_in[2]));
Q_AN03 U2503 ( .A0(n547), .A1(n1211), .A2(n590), .Z(n1210));
Q_MX02 U2504 ( .S(n548), .A0(upsizer_gcm_data[1]), .A1(cmdfifo_gcm_cmd[100]), .Z(n1211));
Q_MX03 U2505 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[228]), .A1(cmdfifo_gcm_cmd[356]), .A2(cmdfifo_gcm_cmd[484]), .Z(n1212));
Q_MX02 U2506 ( .S(n582), .A0(n1215), .A1(n1213), .Z(fifo_in[1]));
Q_AN03 U2507 ( .A0(n547), .A1(n1214), .A2(n590), .Z(n1213));
Q_MX02 U2508 ( .S(n548), .A0(upsizer_gcm_data[0]), .A1(cmdfifo_gcm_cmd[99]), .Z(n1214));
Q_MX03 U2509 ( .S0(n548), .S1(n547), .A0(cmdfifo_gcm_cmd[227]), .A1(cmdfifo_gcm_cmd[355]), .A2(cmdfifo_gcm_cmd[483]), .Z(n1215));
Q_AN02 U2510 ( .A0(n549), .A1(upsizer_gcm_eof), .Z(fifo_in[0]));
Q_MX02 U2511 ( .S(n623), .A0(n1217), .A1(n1216), .Z(stream_end));
Q_MX02 U2512 ( .S(n550), .A0(n1218), .A1(combo_dek512), .Z(nxt_combo_dek512));
Q_AN02 U2513 ( .A0(n551), .A1(upsizer_gcm_eof), .Z(n1218));
Q_AN03 U2514 ( .A0(upsizer_gcm_eof), .A1(n1219), .A2(n627), .Z(n1216));
Q_INV U2515 ( .A(n539), .Z(n1219));
Q_AN02 U2516 ( .A0(n1220), .A1(upsizer_gcm_eof), .Z(n634));
Q_AN03 U2517 ( .A0(cmdfifo_gcm_cmd[0]), .A1(n605), .A2(cmdfifo_gcm_cmd[2]), .Z(n1221));
Q_AN02 U2518 ( .A0(upsizer_gcm_eof), .A1(n2), .Z(n1217));
Q_INV U2519 ( .A(n1221), .Z(n1222));
Q_XOR2 U2520 ( .A0(cmdfifo_gcm_cmd[1]), .A1(n595), .Z(n542));
Q_AN02 U2521 ( .A0(n1223), .A1(gcm_tag_data_out_valid), .Z(n540));
Q_INV U2522 ( .A(ciph_fifo_in_stall), .Z(n1223));
Q_AN03 U2523 ( .A0(n1224), .A1(cmdfifo_gcm_cmd[1]), .A2(cmdfifo_gcm_cmd[2]), .Z(n539));
Q_INV U2524 ( .A(cmdfifo_gcm_cmd[0]), .Z(n1224));
Q_ND02 U2525 ( .A0(cmdfifo_gcm_valid), .A1(n1225), .Z(n541));
Q_INV U2526 ( .A(key_in_stall), .Z(n1225));
Q_OR02 U2527 ( .A0(ciph_in_stall), .A1(fifo_in_stall), .Z(ciph_fifo_in_stall));
Q_AN02 U2528 ( .A0(n1238), .A1(cur_state[1]), .Z(n1245));
Q_AN03 U2529 ( .A0(cur_state[0]), .A1(n1230), .A2(n1245), .Z(n1231));
Q_INV U2530 ( .A(n1226), .Z(n1230));
Q_AN02 U2531 ( .A0(cur_state[2]), .A1(n1237), .Z(n1232));
Q_AO21 U2532 ( .A0(n1232), .A1(n1243), .B0(n1231), .Z(n1242));
Q_AO21 U2533 ( .A0(n1232), .A1(cur_state[0]), .B0(n1242), .Z(n1234));
Q_AN03 U2534 ( .A0(ciph_in_vld), .A1(n1226), .A2(cur_state[0]), .Z(n1233));
Q_OA21 U2535 ( .A0(n1233), .A1(n1244), .B0(n1245), .Z(n1235));
Q_AN02 U2536 ( .A0(n1234), .A1(ciph_in_vld), .Z(n1240));
Q_OR02 U2537 ( .A0(n1240), .A1(n1235), .Z(n1236));
Q_INV U2538 ( .A(n1236), .Z(n1227));
Q_AO21 U2539 ( .A0(cur_state[0]), .A1(ciph_in_vld), .B0(n1247), .Z(n1239));
Q_NR02 U2540 ( .A0(cur_state[0]), .A1(ciph_in_stall), .Z(n1247));
Q_NR02 U2541 ( .A0(cur_state[2]), .A1(cur_state[1]), .Z(n1248));
Q_AO21 U2542 ( .A0(n1239), .A1(n1248), .B0(n1240), .Z(n1241));
Q_INV U2543 ( .A(n1241), .Z(n1228));
Q_AO21 U2544 ( .A0(n1242), .A1(ciph_in_vld), .B0(n1249), .Z(n1229));
Q_AN02 U2545 ( .A0(n1243), .A1(stream_end), .Z(n1244));
Q_AO21 U2546 ( .A0(n1245), .A1(n1244), .B0(n1246), .Z(n1249));
Q_AN02 U2547 ( .A0(n1248), .A1(n1247), .Z(n1246));
Q_AO21 U2548 ( .A0(n1250), .A1(cur_state[0]), .B0(n1229), .Z(nxt_state[0]));
Q_AO21 U2549 ( .A0(n1250), .A1(cur_state[1]), .B0(n1255), .Z(nxt_state[1]));
Q_AO21 U2550 ( .A0(n1250), .A1(cur_state[2]), .B0(n1253), .Z(nxt_state[2]));
Q_NR02 U2551 ( .A0(n1241), .A1(n1236), .Z(n1250));
Q_XOR2 U2552 ( .A0(n1228), .A1(n1236), .Z(n1251));
Q_NR02 U2553 ( .A0(n1241), .A1(n1227), .Z(n1252));
Q_MX02 U2554 ( .S(n1229), .A0(n1252), .A1(n1251), .Z(n1253));
Q_NR02 U2555 ( .A0(n1228), .A1(n1236), .Z(n1254));
Q_MX02 U2556 ( .S(n1229), .A0(n1254), .A1(n1228), .Z(n1255));
Q_AN03 U2557 ( .A0(cmdfifo_gcm_cmd[0]), .A1(cmdfifo_gcm_cmd[1]), .A2(cmdfifo_gcm_cmd[2]), .Z(n1226));
Q_INV U2558 ( .A(upsizer_gcm_eof), .Z(n1256));
Q_AN02 U2559 ( .A0(n1256), .A1(n1259), .Z(n1257));
Q_NR02 U2560 ( .A0(upsizer_gcm_eof), .A1(beat_num[0]), .Z(n1258));
Q_XOR2 U2561 ( .A0(beat_num[1]), .A1(beat_num[0]), .Z(n1259));
Q_AN02 U2562 ( .A0(n1647), .A1(n1260), .Z(n1261));
Q_MX02 U2563 ( .S(n1647), .A0(cmdfifo_gcm_cmd[98]), .A1(n1391), .Z(n1262));
Q_MX02 U2564 ( .S(n1647), .A0(cmdfifo_gcm_cmd[97]), .A1(n1393), .Z(n1263));
Q_MX02 U2565 ( .S(n1647), .A0(cmdfifo_gcm_cmd[96]), .A1(n1395), .Z(n1264));
Q_MX02 U2566 ( .S(n1647), .A0(cmdfifo_gcm_cmd[95]), .A1(n1397), .Z(n1265));
Q_MX02 U2567 ( .S(n1647), .A0(cmdfifo_gcm_cmd[94]), .A1(n1399), .Z(n1266));
Q_MX02 U2568 ( .S(n1647), .A0(cmdfifo_gcm_cmd[93]), .A1(n1401), .Z(n1267));
Q_MX02 U2569 ( .S(n1647), .A0(cmdfifo_gcm_cmd[92]), .A1(n1403), .Z(n1268));
Q_MX02 U2570 ( .S(n1647), .A0(cmdfifo_gcm_cmd[91]), .A1(n1405), .Z(n1269));
Q_MX02 U2571 ( .S(n1647), .A0(cmdfifo_gcm_cmd[90]), .A1(n1407), .Z(n1270));
Q_MX02 U2572 ( .S(n1647), .A0(cmdfifo_gcm_cmd[89]), .A1(n1409), .Z(n1271));
Q_MX02 U2573 ( .S(n1647), .A0(cmdfifo_gcm_cmd[88]), .A1(n1411), .Z(n1272));
Q_MX02 U2574 ( .S(n1647), .A0(cmdfifo_gcm_cmd[87]), .A1(n1413), .Z(n1273));
Q_MX02 U2575 ( .S(n1647), .A0(cmdfifo_gcm_cmd[86]), .A1(n1415), .Z(n1274));
Q_MX02 U2576 ( .S(n1647), .A0(cmdfifo_gcm_cmd[85]), .A1(n1417), .Z(n1275));
Q_MX02 U2577 ( .S(n1647), .A0(cmdfifo_gcm_cmd[84]), .A1(n1419), .Z(n1276));
Q_MX02 U2578 ( .S(n1647), .A0(cmdfifo_gcm_cmd[83]), .A1(n1421), .Z(n1277));
Q_MX02 U2579 ( .S(n1647), .A0(cmdfifo_gcm_cmd[82]), .A1(n1423), .Z(n1278));
Q_MX02 U2580 ( .S(n1647), .A0(cmdfifo_gcm_cmd[81]), .A1(n1425), .Z(n1279));
Q_MX02 U2581 ( .S(n1647), .A0(cmdfifo_gcm_cmd[80]), .A1(n1427), .Z(n1280));
Q_MX02 U2582 ( .S(n1647), .A0(cmdfifo_gcm_cmd[79]), .A1(n1429), .Z(n1281));
Q_MX02 U2583 ( .S(n1647), .A0(cmdfifo_gcm_cmd[78]), .A1(n1431), .Z(n1282));
Q_MX02 U2584 ( .S(n1647), .A0(cmdfifo_gcm_cmd[77]), .A1(n1433), .Z(n1283));
Q_MX02 U2585 ( .S(n1647), .A0(cmdfifo_gcm_cmd[76]), .A1(n1435), .Z(n1284));
Q_MX02 U2586 ( .S(n1647), .A0(cmdfifo_gcm_cmd[75]), .A1(n1437), .Z(n1285));
Q_MX02 U2587 ( .S(n1647), .A0(cmdfifo_gcm_cmd[74]), .A1(n1439), .Z(n1286));
Q_MX02 U2588 ( .S(n1647), .A0(cmdfifo_gcm_cmd[73]), .A1(n1441), .Z(n1287));
Q_MX02 U2589 ( .S(n1647), .A0(cmdfifo_gcm_cmd[72]), .A1(n1443), .Z(n1288));
Q_MX02 U2590 ( .S(n1647), .A0(cmdfifo_gcm_cmd[71]), .A1(n1445), .Z(n1289));
Q_MX02 U2591 ( .S(n1647), .A0(cmdfifo_gcm_cmd[70]), .A1(n1447), .Z(n1290));
Q_MX02 U2592 ( .S(n1647), .A0(cmdfifo_gcm_cmd[69]), .A1(n1449), .Z(n1291));
Q_MX02 U2593 ( .S(n1647), .A0(cmdfifo_gcm_cmd[68]), .A1(n1451), .Z(n1292));
Q_MX02 U2594 ( .S(n1647), .A0(cmdfifo_gcm_cmd[67]), .A1(n1453), .Z(n1293));
Q_MX02 U2595 ( .S(n1647), .A0(cmdfifo_gcm_cmd[66]), .A1(n1455), .Z(n1294));
Q_MX02 U2596 ( .S(n1647), .A0(cmdfifo_gcm_cmd[65]), .A1(n1457), .Z(n1295));
Q_MX02 U2597 ( .S(n1647), .A0(cmdfifo_gcm_cmd[64]), .A1(n1459), .Z(n1296));
Q_MX02 U2598 ( .S(n1647), .A0(cmdfifo_gcm_cmd[63]), .A1(n1461), .Z(n1297));
Q_MX02 U2599 ( .S(n1647), .A0(cmdfifo_gcm_cmd[62]), .A1(n1463), .Z(n1298));
Q_MX02 U2600 ( .S(n1647), .A0(cmdfifo_gcm_cmd[61]), .A1(n1465), .Z(n1299));
Q_MX02 U2601 ( .S(n1647), .A0(cmdfifo_gcm_cmd[60]), .A1(n1467), .Z(n1300));
Q_MX02 U2602 ( .S(n1647), .A0(cmdfifo_gcm_cmd[59]), .A1(n1469), .Z(n1301));
Q_MX02 U2603 ( .S(n1647), .A0(cmdfifo_gcm_cmd[58]), .A1(n1471), .Z(n1302));
Q_MX02 U2604 ( .S(n1647), .A0(cmdfifo_gcm_cmd[57]), .A1(n1473), .Z(n1303));
Q_MX02 U2605 ( .S(n1647), .A0(cmdfifo_gcm_cmd[56]), .A1(n1475), .Z(n1304));
Q_MX02 U2606 ( .S(n1647), .A0(cmdfifo_gcm_cmd[55]), .A1(n1477), .Z(n1305));
Q_MX02 U2607 ( .S(n1647), .A0(cmdfifo_gcm_cmd[54]), .A1(n1479), .Z(n1306));
Q_MX02 U2608 ( .S(n1647), .A0(cmdfifo_gcm_cmd[53]), .A1(n1481), .Z(n1307));
Q_MX02 U2609 ( .S(n1647), .A0(cmdfifo_gcm_cmd[52]), .A1(n1483), .Z(n1308));
Q_MX02 U2610 ( .S(n1647), .A0(cmdfifo_gcm_cmd[51]), .A1(n1485), .Z(n1309));
Q_MX02 U2611 ( .S(n1647), .A0(cmdfifo_gcm_cmd[50]), .A1(n1487), .Z(n1310));
Q_MX02 U2612 ( .S(n1647), .A0(cmdfifo_gcm_cmd[49]), .A1(n1489), .Z(n1311));
Q_MX02 U2613 ( .S(n1647), .A0(cmdfifo_gcm_cmd[48]), .A1(n1491), .Z(n1312));
Q_MX02 U2614 ( .S(n1647), .A0(cmdfifo_gcm_cmd[47]), .A1(n1493), .Z(n1313));
Q_MX02 U2615 ( .S(n1647), .A0(cmdfifo_gcm_cmd[46]), .A1(n1495), .Z(n1314));
Q_MX02 U2616 ( .S(n1647), .A0(cmdfifo_gcm_cmd[45]), .A1(n1497), .Z(n1315));
Q_MX02 U2617 ( .S(n1647), .A0(cmdfifo_gcm_cmd[44]), .A1(n1499), .Z(n1316));
Q_MX02 U2618 ( .S(n1647), .A0(cmdfifo_gcm_cmd[43]), .A1(n1501), .Z(n1317));
Q_MX02 U2619 ( .S(n1647), .A0(cmdfifo_gcm_cmd[42]), .A1(n1503), .Z(n1318));
Q_MX02 U2620 ( .S(n1647), .A0(cmdfifo_gcm_cmd[41]), .A1(n1505), .Z(n1319));
Q_MX02 U2621 ( .S(n1647), .A0(cmdfifo_gcm_cmd[40]), .A1(n1507), .Z(n1320));
Q_MX02 U2622 ( .S(n1647), .A0(cmdfifo_gcm_cmd[39]), .A1(n1509), .Z(n1321));
Q_MX02 U2623 ( .S(n1647), .A0(cmdfifo_gcm_cmd[38]), .A1(n1511), .Z(n1322));
Q_MX02 U2624 ( .S(n1647), .A0(cmdfifo_gcm_cmd[37]), .A1(n1513), .Z(n1323));
Q_MX02 U2625 ( .S(n1647), .A0(cmdfifo_gcm_cmd[36]), .A1(n1515), .Z(n1324));
Q_MX02 U2626 ( .S(n1647), .A0(cmdfifo_gcm_cmd[35]), .A1(n1517), .Z(n1325));
Q_MX02 U2627 ( .S(n1647), .A0(cmdfifo_gcm_cmd[34]), .A1(n1519), .Z(n1326));
Q_MX02 U2628 ( .S(n1647), .A0(cmdfifo_gcm_cmd[33]), .A1(n1521), .Z(n1327));
Q_MX02 U2629 ( .S(n1647), .A0(cmdfifo_gcm_cmd[32]), .A1(n1523), .Z(n1328));
Q_MX02 U2630 ( .S(n1647), .A0(cmdfifo_gcm_cmd[31]), .A1(n1525), .Z(n1329));
Q_MX02 U2631 ( .S(n1647), .A0(cmdfifo_gcm_cmd[30]), .A1(n1527), .Z(n1330));
Q_MX02 U2632 ( .S(n1647), .A0(cmdfifo_gcm_cmd[29]), .A1(n1529), .Z(n1331));
Q_MX02 U2633 ( .S(n1647), .A0(cmdfifo_gcm_cmd[28]), .A1(n1531), .Z(n1332));
Q_MX02 U2634 ( .S(n1647), .A0(cmdfifo_gcm_cmd[27]), .A1(n1533), .Z(n1333));
Q_MX02 U2635 ( .S(n1647), .A0(cmdfifo_gcm_cmd[26]), .A1(n1535), .Z(n1334));
Q_MX02 U2636 ( .S(n1647), .A0(cmdfifo_gcm_cmd[25]), .A1(n1537), .Z(n1335));
Q_MX02 U2637 ( .S(n1647), .A0(cmdfifo_gcm_cmd[24]), .A1(n1539), .Z(n1336));
Q_MX02 U2638 ( .S(n1647), .A0(cmdfifo_gcm_cmd[23]), .A1(n1541), .Z(n1337));
Q_MX02 U2639 ( .S(n1647), .A0(cmdfifo_gcm_cmd[22]), .A1(n1543), .Z(n1338));
Q_MX02 U2640 ( .S(n1647), .A0(cmdfifo_gcm_cmd[21]), .A1(n1545), .Z(n1339));
Q_MX02 U2641 ( .S(n1647), .A0(cmdfifo_gcm_cmd[20]), .A1(n1547), .Z(n1340));
Q_MX02 U2642 ( .S(n1647), .A0(cmdfifo_gcm_cmd[19]), .A1(n1549), .Z(n1341));
Q_MX02 U2643 ( .S(n1647), .A0(cmdfifo_gcm_cmd[18]), .A1(n1551), .Z(n1342));
Q_MX02 U2644 ( .S(n1647), .A0(cmdfifo_gcm_cmd[17]), .A1(n1553), .Z(n1343));
Q_MX02 U2645 ( .S(n1647), .A0(cmdfifo_gcm_cmd[16]), .A1(n1555), .Z(n1344));
Q_MX02 U2646 ( .S(n1647), .A0(cmdfifo_gcm_cmd[15]), .A1(n1557), .Z(n1345));
Q_MX02 U2647 ( .S(n1647), .A0(cmdfifo_gcm_cmd[14]), .A1(n1559), .Z(n1346));
Q_MX02 U2648 ( .S(n1647), .A0(cmdfifo_gcm_cmd[13]), .A1(n1561), .Z(n1347));
Q_MX02 U2649 ( .S(n1647), .A0(cmdfifo_gcm_cmd[12]), .A1(n1563), .Z(n1348));
Q_MX02 U2650 ( .S(n1647), .A0(cmdfifo_gcm_cmd[11]), .A1(n1565), .Z(n1349));
Q_MX02 U2651 ( .S(n1647), .A0(cmdfifo_gcm_cmd[10]), .A1(n1567), .Z(n1350));
Q_MX02 U2652 ( .S(n1647), .A0(cmdfifo_gcm_cmd[9]), .A1(n1569), .Z(n1351));
Q_MX02 U2653 ( .S(n1647), .A0(cmdfifo_gcm_cmd[8]), .A1(n1571), .Z(n1352));
Q_MX02 U2654 ( .S(n1647), .A0(cmdfifo_gcm_cmd[7]), .A1(n1573), .Z(n1353));
Q_MX02 U2655 ( .S(n1647), .A0(cmdfifo_gcm_cmd[6]), .A1(n1575), .Z(n1354));
Q_MX02 U2656 ( .S(n1647), .A0(cmdfifo_gcm_cmd[5]), .A1(n1577), .Z(n1355));
Q_MX02 U2657 ( .S(n1647), .A0(cmdfifo_gcm_cmd[4]), .A1(n1579), .Z(n1356));
Q_MX02 U2658 ( .S(n1647), .A0(cmdfifo_gcm_cmd[3]), .A1(n1581), .Z(n1357));
Q_AN02 U2659 ( .A0(n1647), .A1(n1583), .Z(n1358));
Q_AN02 U2660 ( .A0(n1647), .A1(n1585), .Z(n1359));
Q_AN02 U2661 ( .A0(n1647), .A1(n1587), .Z(n1360));
Q_AN02 U2662 ( .A0(n1647), .A1(n1589), .Z(n1361));
Q_AN02 U2663 ( .A0(n1647), .A1(n1591), .Z(n1362));
Q_AN02 U2664 ( .A0(n1647), .A1(n1593), .Z(n1363));
Q_AN02 U2665 ( .A0(n1647), .A1(n1595), .Z(n1364));
Q_AN02 U2666 ( .A0(n1647), .A1(n1597), .Z(n1365));
Q_AN02 U2667 ( .A0(n1647), .A1(n1599), .Z(n1366));
Q_AN02 U2668 ( .A0(n1647), .A1(n1601), .Z(n1367));
Q_AN02 U2669 ( .A0(n1647), .A1(n1603), .Z(n1368));
Q_AN02 U2670 ( .A0(n1647), .A1(n1605), .Z(n1369));
Q_AN02 U2671 ( .A0(n1647), .A1(n1607), .Z(n1370));
Q_AN02 U2672 ( .A0(n1647), .A1(n1609), .Z(n1371));
Q_AN02 U2673 ( .A0(n1647), .A1(n1611), .Z(n1372));
Q_AN02 U2674 ( .A0(n1647), .A1(n1613), .Z(n1373));
Q_AN02 U2675 ( .A0(n1647), .A1(n1615), .Z(n1374));
Q_AN02 U2676 ( .A0(n1647), .A1(n1617), .Z(n1375));
Q_AN02 U2677 ( .A0(n1647), .A1(n1619), .Z(n1376));
Q_AN02 U2678 ( .A0(n1647), .A1(n1621), .Z(n1377));
Q_AN02 U2679 ( .A0(n1647), .A1(n1623), .Z(n1378));
Q_AN02 U2680 ( .A0(n1647), .A1(n1625), .Z(n1379));
Q_AN02 U2681 ( .A0(n1647), .A1(n1627), .Z(n1380));
Q_AN02 U2682 ( .A0(n1647), .A1(n1629), .Z(n1381));
Q_AN02 U2683 ( .A0(n1647), .A1(n1631), .Z(n1382));
Q_AN02 U2684 ( .A0(n1647), .A1(n1633), .Z(n1383));
Q_AN02 U2685 ( .A0(n1647), .A1(n1635), .Z(n1384));
Q_AN02 U2686 ( .A0(n1647), .A1(n1637), .Z(n1385));
Q_AN02 U2687 ( .A0(n1647), .A1(n1639), .Z(n1386));
Q_AN02 U2688 ( .A0(n1647), .A1(n1641), .Z(n1387));
Q_OR02 U2689 ( .A0(n1389), .A1(n1643), .Z(n1388));
Q_INV U2690 ( .A(n1647), .Z(n1389));
Q_AN02 U2691 ( .A0(n1647), .A1(n1644), .Z(n1390));
Q_XOR2 U2692 ( .A0(iv_counter[127]), .A1(n1392), .Z(n1391));
Q_AD01HF U2693 ( .A0(iv_counter[126]), .B0(n1394), .S(n1393), .CO(n1392));
Q_AD01HF U2694 ( .A0(iv_counter[125]), .B0(n1396), .S(n1395), .CO(n1394));
Q_AD01HF U2695 ( .A0(iv_counter[124]), .B0(n1398), .S(n1397), .CO(n1396));
Q_AD01HF U2696 ( .A0(iv_counter[123]), .B0(n1400), .S(n1399), .CO(n1398));
Q_AD01HF U2697 ( .A0(iv_counter[122]), .B0(n1402), .S(n1401), .CO(n1400));
Q_AD01HF U2698 ( .A0(iv_counter[121]), .B0(n1404), .S(n1403), .CO(n1402));
Q_AD01HF U2699 ( .A0(iv_counter[120]), .B0(n1406), .S(n1405), .CO(n1404));
Q_AD01HF U2700 ( .A0(iv_counter[119]), .B0(n1408), .S(n1407), .CO(n1406));
Q_AD01HF U2701 ( .A0(iv_counter[118]), .B0(n1410), .S(n1409), .CO(n1408));
Q_AD01HF U2702 ( .A0(iv_counter[117]), .B0(n1412), .S(n1411), .CO(n1410));
Q_AD01HF U2703 ( .A0(iv_counter[116]), .B0(n1414), .S(n1413), .CO(n1412));
Q_AD01HF U2704 ( .A0(iv_counter[115]), .B0(n1416), .S(n1415), .CO(n1414));
Q_AD01HF U2705 ( .A0(iv_counter[114]), .B0(n1418), .S(n1417), .CO(n1416));
Q_AD01HF U2706 ( .A0(iv_counter[113]), .B0(n1420), .S(n1419), .CO(n1418));
Q_AD01HF U2707 ( .A0(iv_counter[112]), .B0(n1422), .S(n1421), .CO(n1420));
Q_AD01HF U2708 ( .A0(iv_counter[111]), .B0(n1424), .S(n1423), .CO(n1422));
Q_AD01HF U2709 ( .A0(iv_counter[110]), .B0(n1426), .S(n1425), .CO(n1424));
Q_AD01HF U2710 ( .A0(iv_counter[109]), .B0(n1428), .S(n1427), .CO(n1426));
Q_AD01HF U2711 ( .A0(iv_counter[108]), .B0(n1430), .S(n1429), .CO(n1428));
Q_AD01HF U2712 ( .A0(iv_counter[107]), .B0(n1432), .S(n1431), .CO(n1430));
Q_AD01HF U2713 ( .A0(iv_counter[106]), .B0(n1434), .S(n1433), .CO(n1432));
Q_AD01HF U2714 ( .A0(iv_counter[105]), .B0(n1436), .S(n1435), .CO(n1434));
Q_AD01HF U2715 ( .A0(iv_counter[104]), .B0(n1438), .S(n1437), .CO(n1436));
Q_AD01HF U2716 ( .A0(iv_counter[103]), .B0(n1440), .S(n1439), .CO(n1438));
Q_AD01HF U2717 ( .A0(iv_counter[102]), .B0(n1442), .S(n1441), .CO(n1440));
Q_AD01HF U2718 ( .A0(iv_counter[101]), .B0(n1444), .S(n1443), .CO(n1442));
Q_AD01HF U2719 ( .A0(iv_counter[100]), .B0(n1446), .S(n1445), .CO(n1444));
Q_AD01HF U2720 ( .A0(iv_counter[99]), .B0(n1448), .S(n1447), .CO(n1446));
Q_AD01HF U2721 ( .A0(iv_counter[98]), .B0(n1450), .S(n1449), .CO(n1448));
Q_AD01HF U2722 ( .A0(iv_counter[97]), .B0(n1452), .S(n1451), .CO(n1450));
Q_AD01HF U2723 ( .A0(iv_counter[96]), .B0(n1454), .S(n1453), .CO(n1452));
Q_AD01HF U2724 ( .A0(iv_counter[95]), .B0(n1456), .S(n1455), .CO(n1454));
Q_AD01HF U2725 ( .A0(iv_counter[94]), .B0(n1458), .S(n1457), .CO(n1456));
Q_AD01HF U2726 ( .A0(iv_counter[93]), .B0(n1460), .S(n1459), .CO(n1458));
Q_AD01HF U2727 ( .A0(iv_counter[92]), .B0(n1462), .S(n1461), .CO(n1460));
Q_AD01HF U2728 ( .A0(iv_counter[91]), .B0(n1464), .S(n1463), .CO(n1462));
Q_AD01HF U2729 ( .A0(iv_counter[90]), .B0(n1466), .S(n1465), .CO(n1464));
Q_AD01HF U2730 ( .A0(iv_counter[89]), .B0(n1468), .S(n1467), .CO(n1466));
Q_AD01HF U2731 ( .A0(iv_counter[88]), .B0(n1470), .S(n1469), .CO(n1468));
Q_AD01HF U2732 ( .A0(iv_counter[87]), .B0(n1472), .S(n1471), .CO(n1470));
Q_AD01HF U2733 ( .A0(iv_counter[86]), .B0(n1474), .S(n1473), .CO(n1472));
Q_AD01HF U2734 ( .A0(iv_counter[85]), .B0(n1476), .S(n1475), .CO(n1474));
Q_AD01HF U2735 ( .A0(iv_counter[84]), .B0(n1478), .S(n1477), .CO(n1476));
Q_AD01HF U2736 ( .A0(iv_counter[83]), .B0(n1480), .S(n1479), .CO(n1478));
Q_AD01HF U2737 ( .A0(iv_counter[82]), .B0(n1482), .S(n1481), .CO(n1480));
Q_AD01HF U2738 ( .A0(iv_counter[81]), .B0(n1484), .S(n1483), .CO(n1482));
Q_AD01HF U2739 ( .A0(iv_counter[80]), .B0(n1486), .S(n1485), .CO(n1484));
Q_AD01HF U2740 ( .A0(iv_counter[79]), .B0(n1488), .S(n1487), .CO(n1486));
Q_AD01HF U2741 ( .A0(iv_counter[78]), .B0(n1490), .S(n1489), .CO(n1488));
Q_AD01HF U2742 ( .A0(iv_counter[77]), .B0(n1492), .S(n1491), .CO(n1490));
Q_AD01HF U2743 ( .A0(iv_counter[76]), .B0(n1494), .S(n1493), .CO(n1492));
Q_AD01HF U2744 ( .A0(iv_counter[75]), .B0(n1496), .S(n1495), .CO(n1494));
Q_AD01HF U2745 ( .A0(iv_counter[74]), .B0(n1498), .S(n1497), .CO(n1496));
Q_AD01HF U2746 ( .A0(iv_counter[73]), .B0(n1500), .S(n1499), .CO(n1498));
Q_AD01HF U2747 ( .A0(iv_counter[72]), .B0(n1502), .S(n1501), .CO(n1500));
Q_AD01HF U2748 ( .A0(iv_counter[71]), .B0(n1504), .S(n1503), .CO(n1502));
Q_AD01HF U2749 ( .A0(iv_counter[70]), .B0(n1506), .S(n1505), .CO(n1504));
Q_AD01HF U2750 ( .A0(iv_counter[69]), .B0(n1508), .S(n1507), .CO(n1506));
Q_AD01HF U2751 ( .A0(iv_counter[68]), .B0(n1510), .S(n1509), .CO(n1508));
Q_AD01HF U2752 ( .A0(iv_counter[67]), .B0(n1512), .S(n1511), .CO(n1510));
Q_AD01HF U2753 ( .A0(iv_counter[66]), .B0(n1514), .S(n1513), .CO(n1512));
Q_AD01HF U2754 ( .A0(iv_counter[65]), .B0(n1516), .S(n1515), .CO(n1514));
Q_AD01HF U2755 ( .A0(iv_counter[64]), .B0(n1518), .S(n1517), .CO(n1516));
Q_AD01HF U2756 ( .A0(iv_counter[63]), .B0(n1520), .S(n1519), .CO(n1518));
Q_AD01HF U2757 ( .A0(iv_counter[62]), .B0(n1522), .S(n1521), .CO(n1520));
Q_AD01HF U2758 ( .A0(iv_counter[61]), .B0(n1524), .S(n1523), .CO(n1522));
Q_AD01HF U2759 ( .A0(iv_counter[60]), .B0(n1526), .S(n1525), .CO(n1524));
Q_AD01HF U2760 ( .A0(iv_counter[59]), .B0(n1528), .S(n1527), .CO(n1526));
Q_AD01HF U2761 ( .A0(iv_counter[58]), .B0(n1530), .S(n1529), .CO(n1528));
Q_AD01HF U2762 ( .A0(iv_counter[57]), .B0(n1532), .S(n1531), .CO(n1530));
Q_AD01HF U2763 ( .A0(iv_counter[56]), .B0(n1534), .S(n1533), .CO(n1532));
Q_AD01HF U2764 ( .A0(iv_counter[55]), .B0(n1536), .S(n1535), .CO(n1534));
Q_AD01HF U2765 ( .A0(iv_counter[54]), .B0(n1538), .S(n1537), .CO(n1536));
Q_AD01HF U2766 ( .A0(iv_counter[53]), .B0(n1540), .S(n1539), .CO(n1538));
Q_AD01HF U2767 ( .A0(iv_counter[52]), .B0(n1542), .S(n1541), .CO(n1540));
Q_AD01HF U2768 ( .A0(iv_counter[51]), .B0(n1544), .S(n1543), .CO(n1542));
Q_AD01HF U2769 ( .A0(iv_counter[50]), .B0(n1546), .S(n1545), .CO(n1544));
Q_AD01HF U2770 ( .A0(iv_counter[49]), .B0(n1548), .S(n1547), .CO(n1546));
Q_AD01HF U2771 ( .A0(iv_counter[48]), .B0(n1550), .S(n1549), .CO(n1548));
Q_AD01HF U2772 ( .A0(iv_counter[47]), .B0(n1552), .S(n1551), .CO(n1550));
Q_AD01HF U2773 ( .A0(iv_counter[46]), .B0(n1554), .S(n1553), .CO(n1552));
Q_AD01HF U2774 ( .A0(iv_counter[45]), .B0(n1556), .S(n1555), .CO(n1554));
Q_AD01HF U2775 ( .A0(iv_counter[44]), .B0(n1558), .S(n1557), .CO(n1556));
Q_AD01HF U2776 ( .A0(iv_counter[43]), .B0(n1560), .S(n1559), .CO(n1558));
Q_AD01HF U2777 ( .A0(iv_counter[42]), .B0(n1562), .S(n1561), .CO(n1560));
Q_AD01HF U2778 ( .A0(iv_counter[41]), .B0(n1564), .S(n1563), .CO(n1562));
Q_AD01HF U2779 ( .A0(iv_counter[40]), .B0(n1566), .S(n1565), .CO(n1564));
Q_AD01HF U2780 ( .A0(iv_counter[39]), .B0(n1568), .S(n1567), .CO(n1566));
Q_AD01HF U2781 ( .A0(iv_counter[38]), .B0(n1570), .S(n1569), .CO(n1568));
Q_AD01HF U2782 ( .A0(iv_counter[37]), .B0(n1572), .S(n1571), .CO(n1570));
Q_AD01HF U2783 ( .A0(iv_counter[36]), .B0(n1574), .S(n1573), .CO(n1572));
Q_AD01HF U2784 ( .A0(iv_counter[35]), .B0(n1576), .S(n1575), .CO(n1574));
Q_AD01HF U2785 ( .A0(iv_counter[34]), .B0(n1578), .S(n1577), .CO(n1576));
Q_AD01HF U2786 ( .A0(iv_counter[33]), .B0(n1580), .S(n1579), .CO(n1578));
Q_AD01HF U2787 ( .A0(iv_counter[32]), .B0(n1582), .S(n1581), .CO(n1580));
Q_AD01HF U2788 ( .A0(iv_counter[31]), .B0(n1584), .S(n1583), .CO(n1582));
Q_AD01HF U2789 ( .A0(iv_counter[30]), .B0(n1586), .S(n1585), .CO(n1584));
Q_AD01HF U2790 ( .A0(iv_counter[29]), .B0(n1588), .S(n1587), .CO(n1586));
Q_AD01HF U2791 ( .A0(iv_counter[28]), .B0(n1590), .S(n1589), .CO(n1588));
Q_AD01HF U2792 ( .A0(iv_counter[27]), .B0(n1592), .S(n1591), .CO(n1590));
Q_AD01HF U2793 ( .A0(iv_counter[26]), .B0(n1594), .S(n1593), .CO(n1592));
Q_AD01HF U2794 ( .A0(iv_counter[25]), .B0(n1596), .S(n1595), .CO(n1594));
Q_AD01HF U2795 ( .A0(iv_counter[24]), .B0(n1598), .S(n1597), .CO(n1596));
Q_AD01HF U2796 ( .A0(iv_counter[23]), .B0(n1600), .S(n1599), .CO(n1598));
Q_AD01HF U2797 ( .A0(iv_counter[22]), .B0(n1602), .S(n1601), .CO(n1600));
Q_AD01HF U2798 ( .A0(iv_counter[21]), .B0(n1604), .S(n1603), .CO(n1602));
Q_AD01HF U2799 ( .A0(iv_counter[20]), .B0(n1606), .S(n1605), .CO(n1604));
Q_AD01HF U2800 ( .A0(iv_counter[19]), .B0(n1608), .S(n1607), .CO(n1606));
Q_AD01HF U2801 ( .A0(iv_counter[18]), .B0(n1610), .S(n1609), .CO(n1608));
Q_AD01HF U2802 ( .A0(iv_counter[17]), .B0(n1612), .S(n1611), .CO(n1610));
Q_AD01HF U2803 ( .A0(iv_counter[16]), .B0(n1614), .S(n1613), .CO(n1612));
Q_AD01HF U2804 ( .A0(iv_counter[15]), .B0(n1616), .S(n1615), .CO(n1614));
Q_AD01HF U2805 ( .A0(iv_counter[14]), .B0(n1618), .S(n1617), .CO(n1616));
Q_AD01HF U2806 ( .A0(iv_counter[13]), .B0(n1620), .S(n1619), .CO(n1618));
Q_AD01HF U2807 ( .A0(iv_counter[12]), .B0(n1622), .S(n1621), .CO(n1620));
Q_AD01HF U2808 ( .A0(iv_counter[11]), .B0(n1624), .S(n1623), .CO(n1622));
Q_AD01HF U2809 ( .A0(iv_counter[10]), .B0(n1626), .S(n1625), .CO(n1624));
Q_AD01HF U2810 ( .A0(iv_counter[9]), .B0(n1628), .S(n1627), .CO(n1626));
Q_AD01HF U2811 ( .A0(iv_counter[8]), .B0(n1630), .S(n1629), .CO(n1628));
Q_AD01HF U2812 ( .A0(iv_counter[7]), .B0(n1632), .S(n1631), .CO(n1630));
Q_AD01HF U2813 ( .A0(iv_counter[6]), .B0(n1634), .S(n1633), .CO(n1632));
Q_AD01HF U2814 ( .A0(iv_counter[5]), .B0(n1636), .S(n1635), .CO(n1634));
Q_AD01HF U2815 ( .A0(iv_counter[4]), .B0(n1638), .S(n1637), .CO(n1636));
Q_AD01HF U2816 ( .A0(iv_counter[3]), .B0(n1640), .S(n1639), .CO(n1638));
Q_AD01HF U2817 ( .A0(iv_counter[2]), .B0(n1642), .S(n1641), .CO(n1640));
Q_AD01HF U2818 ( .A0(iv_counter[1]), .B0(iv_counter[0]), .S(n1643), .CO(n1642));
Q_OR02 U2819 ( .A0(n563), .A1(n1645), .Z(n1260));
Q_OR03 U2820 ( .A0(fifo_in[129]), .A1(n1646), .A2(fifo_in[131]), .Z(n1645));
Q_INV U2821 ( .A(fifo_in[130]), .Z(n1646));
Q_OR03 U2822 ( .A0(cur_state[0]), .A1(cur_state[1]), .A2(cur_state[2]), .Z(n1647));
Q_FDP1 \cur_state_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_state[2]), .Q(cur_state[2]), .QN(n1238));
Q_FDP1 \cur_state_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_state[1]), .Q(cur_state[1]), .QN(n1237));
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN(n1243));
Q_FDP1 \h_value_REG[127] ( .CK(clk), .R(rst_n), .D(nxt_h_value[127]), .Q(h_value[127]), .QN( ));
Q_FDP1 \h_value_REG[126] ( .CK(clk), .R(rst_n), .D(nxt_h_value[126]), .Q(h_value[126]), .QN( ));
Q_FDP1 \h_value_REG[125] ( .CK(clk), .R(rst_n), .D(nxt_h_value[125]), .Q(h_value[125]), .QN( ));
Q_FDP1 \h_value_REG[124] ( .CK(clk), .R(rst_n), .D(nxt_h_value[124]), .Q(h_value[124]), .QN( ));
Q_FDP1 \h_value_REG[123] ( .CK(clk), .R(rst_n), .D(nxt_h_value[123]), .Q(h_value[123]), .QN( ));
Q_FDP1 \h_value_REG[122] ( .CK(clk), .R(rst_n), .D(nxt_h_value[122]), .Q(h_value[122]), .QN( ));
Q_FDP1 \h_value_REG[121] ( .CK(clk), .R(rst_n), .D(nxt_h_value[121]), .Q(h_value[121]), .QN( ));
Q_FDP1 \h_value_REG[120] ( .CK(clk), .R(rst_n), .D(nxt_h_value[120]), .Q(h_value[120]), .QN( ));
Q_FDP1 \h_value_REG[119] ( .CK(clk), .R(rst_n), .D(nxt_h_value[119]), .Q(h_value[119]), .QN( ));
Q_FDP1 \h_value_REG[118] ( .CK(clk), .R(rst_n), .D(nxt_h_value[118]), .Q(h_value[118]), .QN( ));
Q_FDP1 \h_value_REG[117] ( .CK(clk), .R(rst_n), .D(nxt_h_value[117]), .Q(h_value[117]), .QN( ));
Q_FDP1 \h_value_REG[116] ( .CK(clk), .R(rst_n), .D(nxt_h_value[116]), .Q(h_value[116]), .QN( ));
Q_FDP1 \h_value_REG[115] ( .CK(clk), .R(rst_n), .D(nxt_h_value[115]), .Q(h_value[115]), .QN( ));
Q_FDP1 \h_value_REG[114] ( .CK(clk), .R(rst_n), .D(nxt_h_value[114]), .Q(h_value[114]), .QN( ));
Q_FDP1 \h_value_REG[113] ( .CK(clk), .R(rst_n), .D(nxt_h_value[113]), .Q(h_value[113]), .QN( ));
Q_FDP1 \h_value_REG[112] ( .CK(clk), .R(rst_n), .D(nxt_h_value[112]), .Q(h_value[112]), .QN( ));
Q_FDP1 \h_value_REG[111] ( .CK(clk), .R(rst_n), .D(nxt_h_value[111]), .Q(h_value[111]), .QN( ));
Q_FDP1 \h_value_REG[110] ( .CK(clk), .R(rst_n), .D(nxt_h_value[110]), .Q(h_value[110]), .QN( ));
Q_FDP1 \h_value_REG[109] ( .CK(clk), .R(rst_n), .D(nxt_h_value[109]), .Q(h_value[109]), .QN( ));
Q_FDP1 \h_value_REG[108] ( .CK(clk), .R(rst_n), .D(nxt_h_value[108]), .Q(h_value[108]), .QN( ));
Q_FDP1 \h_value_REG[107] ( .CK(clk), .R(rst_n), .D(nxt_h_value[107]), .Q(h_value[107]), .QN( ));
Q_FDP1 \h_value_REG[106] ( .CK(clk), .R(rst_n), .D(nxt_h_value[106]), .Q(h_value[106]), .QN( ));
Q_FDP1 \h_value_REG[105] ( .CK(clk), .R(rst_n), .D(nxt_h_value[105]), .Q(h_value[105]), .QN( ));
Q_FDP1 \h_value_REG[104] ( .CK(clk), .R(rst_n), .D(nxt_h_value[104]), .Q(h_value[104]), .QN( ));
Q_FDP1 \h_value_REG[103] ( .CK(clk), .R(rst_n), .D(nxt_h_value[103]), .Q(h_value[103]), .QN( ));
Q_FDP1 \h_value_REG[102] ( .CK(clk), .R(rst_n), .D(nxt_h_value[102]), .Q(h_value[102]), .QN( ));
Q_FDP1 \h_value_REG[101] ( .CK(clk), .R(rst_n), .D(nxt_h_value[101]), .Q(h_value[101]), .QN( ));
Q_FDP1 \h_value_REG[100] ( .CK(clk), .R(rst_n), .D(nxt_h_value[100]), .Q(h_value[100]), .QN( ));
Q_FDP1 \h_value_REG[99] ( .CK(clk), .R(rst_n), .D(nxt_h_value[99]), .Q(h_value[99]), .QN( ));
Q_FDP1 \h_value_REG[98] ( .CK(clk), .R(rst_n), .D(nxt_h_value[98]), .Q(h_value[98]), .QN( ));
Q_FDP1 \h_value_REG[97] ( .CK(clk), .R(rst_n), .D(nxt_h_value[97]), .Q(h_value[97]), .QN( ));
Q_FDP1 \h_value_REG[96] ( .CK(clk), .R(rst_n), .D(nxt_h_value[96]), .Q(h_value[96]), .QN( ));
Q_FDP1 \h_value_REG[95] ( .CK(clk), .R(rst_n), .D(nxt_h_value[95]), .Q(h_value[95]), .QN( ));
Q_FDP1 \h_value_REG[94] ( .CK(clk), .R(rst_n), .D(nxt_h_value[94]), .Q(h_value[94]), .QN( ));
Q_FDP1 \h_value_REG[93] ( .CK(clk), .R(rst_n), .D(nxt_h_value[93]), .Q(h_value[93]), .QN( ));
Q_FDP1 \h_value_REG[92] ( .CK(clk), .R(rst_n), .D(nxt_h_value[92]), .Q(h_value[92]), .QN( ));
Q_FDP1 \h_value_REG[91] ( .CK(clk), .R(rst_n), .D(nxt_h_value[91]), .Q(h_value[91]), .QN( ));
Q_FDP1 \h_value_REG[90] ( .CK(clk), .R(rst_n), .D(nxt_h_value[90]), .Q(h_value[90]), .QN( ));
Q_FDP1 \h_value_REG[89] ( .CK(clk), .R(rst_n), .D(nxt_h_value[89]), .Q(h_value[89]), .QN( ));
Q_FDP1 \h_value_REG[88] ( .CK(clk), .R(rst_n), .D(nxt_h_value[88]), .Q(h_value[88]), .QN( ));
Q_FDP1 \h_value_REG[87] ( .CK(clk), .R(rst_n), .D(nxt_h_value[87]), .Q(h_value[87]), .QN( ));
Q_FDP1 \h_value_REG[86] ( .CK(clk), .R(rst_n), .D(nxt_h_value[86]), .Q(h_value[86]), .QN( ));
Q_FDP1 \h_value_REG[85] ( .CK(clk), .R(rst_n), .D(nxt_h_value[85]), .Q(h_value[85]), .QN( ));
Q_FDP1 \h_value_REG[84] ( .CK(clk), .R(rst_n), .D(nxt_h_value[84]), .Q(h_value[84]), .QN( ));
Q_FDP1 \h_value_REG[83] ( .CK(clk), .R(rst_n), .D(nxt_h_value[83]), .Q(h_value[83]), .QN( ));
Q_FDP1 \h_value_REG[82] ( .CK(clk), .R(rst_n), .D(nxt_h_value[82]), .Q(h_value[82]), .QN( ));
Q_FDP1 \h_value_REG[81] ( .CK(clk), .R(rst_n), .D(nxt_h_value[81]), .Q(h_value[81]), .QN( ));
Q_FDP1 \h_value_REG[80] ( .CK(clk), .R(rst_n), .D(nxt_h_value[80]), .Q(h_value[80]), .QN( ));
Q_FDP1 \h_value_REG[79] ( .CK(clk), .R(rst_n), .D(nxt_h_value[79]), .Q(h_value[79]), .QN( ));
Q_FDP1 \h_value_REG[78] ( .CK(clk), .R(rst_n), .D(nxt_h_value[78]), .Q(h_value[78]), .QN( ));
Q_FDP1 \h_value_REG[77] ( .CK(clk), .R(rst_n), .D(nxt_h_value[77]), .Q(h_value[77]), .QN( ));
Q_FDP1 \h_value_REG[76] ( .CK(clk), .R(rst_n), .D(nxt_h_value[76]), .Q(h_value[76]), .QN( ));
Q_FDP1 \h_value_REG[75] ( .CK(clk), .R(rst_n), .D(nxt_h_value[75]), .Q(h_value[75]), .QN( ));
Q_FDP1 \h_value_REG[74] ( .CK(clk), .R(rst_n), .D(nxt_h_value[74]), .Q(h_value[74]), .QN( ));
Q_FDP1 \h_value_REG[73] ( .CK(clk), .R(rst_n), .D(nxt_h_value[73]), .Q(h_value[73]), .QN( ));
Q_FDP1 \h_value_REG[72] ( .CK(clk), .R(rst_n), .D(nxt_h_value[72]), .Q(h_value[72]), .QN( ));
Q_FDP1 \h_value_REG[71] ( .CK(clk), .R(rst_n), .D(nxt_h_value[71]), .Q(h_value[71]), .QN( ));
Q_FDP1 \h_value_REG[70] ( .CK(clk), .R(rst_n), .D(nxt_h_value[70]), .Q(h_value[70]), .QN( ));
Q_FDP1 \h_value_REG[69] ( .CK(clk), .R(rst_n), .D(nxt_h_value[69]), .Q(h_value[69]), .QN( ));
Q_FDP1 \h_value_REG[68] ( .CK(clk), .R(rst_n), .D(nxt_h_value[68]), .Q(h_value[68]), .QN( ));
Q_FDP1 \h_value_REG[67] ( .CK(clk), .R(rst_n), .D(nxt_h_value[67]), .Q(h_value[67]), .QN( ));
Q_FDP1 \h_value_REG[66] ( .CK(clk), .R(rst_n), .D(nxt_h_value[66]), .Q(h_value[66]), .QN( ));
Q_FDP1 \h_value_REG[65] ( .CK(clk), .R(rst_n), .D(nxt_h_value[65]), .Q(h_value[65]), .QN( ));
Q_FDP1 \h_value_REG[64] ( .CK(clk), .R(rst_n), .D(nxt_h_value[64]), .Q(h_value[64]), .QN( ));
Q_FDP1 \h_value_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_h_value[63]), .Q(h_value[63]), .QN( ));
Q_FDP1 \h_value_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_h_value[62]), .Q(h_value[62]), .QN( ));
Q_FDP1 \h_value_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_h_value[61]), .Q(h_value[61]), .QN( ));
Q_FDP1 \h_value_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_h_value[60]), .Q(h_value[60]), .QN( ));
Q_FDP1 \h_value_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_h_value[59]), .Q(h_value[59]), .QN( ));
Q_FDP1 \h_value_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_h_value[58]), .Q(h_value[58]), .QN( ));
Q_FDP1 \h_value_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_h_value[57]), .Q(h_value[57]), .QN( ));
Q_FDP1 \h_value_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_h_value[56]), .Q(h_value[56]), .QN( ));
Q_FDP1 \h_value_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_h_value[55]), .Q(h_value[55]), .QN( ));
Q_FDP1 \h_value_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_h_value[54]), .Q(h_value[54]), .QN( ));
Q_FDP1 \h_value_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_h_value[53]), .Q(h_value[53]), .QN( ));
Q_FDP1 \h_value_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_h_value[52]), .Q(h_value[52]), .QN( ));
Q_FDP1 \h_value_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_h_value[51]), .Q(h_value[51]), .QN( ));
Q_FDP1 \h_value_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_h_value[50]), .Q(h_value[50]), .QN( ));
Q_FDP1 \h_value_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_h_value[49]), .Q(h_value[49]), .QN( ));
Q_FDP1 \h_value_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_h_value[48]), .Q(h_value[48]), .QN( ));
Q_FDP1 \h_value_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_h_value[47]), .Q(h_value[47]), .QN( ));
Q_FDP1 \h_value_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_h_value[46]), .Q(h_value[46]), .QN( ));
Q_FDP1 \h_value_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_h_value[45]), .Q(h_value[45]), .QN( ));
Q_FDP1 \h_value_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_h_value[44]), .Q(h_value[44]), .QN( ));
Q_FDP1 \h_value_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_h_value[43]), .Q(h_value[43]), .QN( ));
Q_FDP1 \h_value_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_h_value[42]), .Q(h_value[42]), .QN( ));
Q_FDP1 \h_value_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_h_value[41]), .Q(h_value[41]), .QN( ));
Q_FDP1 \h_value_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_h_value[40]), .Q(h_value[40]), .QN( ));
Q_FDP1 \h_value_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_h_value[39]), .Q(h_value[39]), .QN( ));
Q_FDP1 \h_value_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_h_value[38]), .Q(h_value[38]), .QN( ));
Q_FDP1 \h_value_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_h_value[37]), .Q(h_value[37]), .QN( ));
Q_FDP1 \h_value_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_h_value[36]), .Q(h_value[36]), .QN( ));
Q_FDP1 \h_value_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_h_value[35]), .Q(h_value[35]), .QN( ));
Q_FDP1 \h_value_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_h_value[34]), .Q(h_value[34]), .QN( ));
Q_FDP1 \h_value_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_h_value[33]), .Q(h_value[33]), .QN( ));
Q_FDP1 \h_value_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_h_value[32]), .Q(h_value[32]), .QN( ));
Q_FDP1 \h_value_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_h_value[31]), .Q(h_value[31]), .QN( ));
Q_FDP1 \h_value_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_h_value[30]), .Q(h_value[30]), .QN( ));
Q_FDP1 \h_value_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_h_value[29]), .Q(h_value[29]), .QN( ));
Q_FDP1 \h_value_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_h_value[28]), .Q(h_value[28]), .QN( ));
Q_FDP1 \h_value_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_h_value[27]), .Q(h_value[27]), .QN( ));
Q_FDP1 \h_value_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_h_value[26]), .Q(h_value[26]), .QN( ));
Q_FDP1 \h_value_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_h_value[25]), .Q(h_value[25]), .QN( ));
Q_FDP1 \h_value_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_h_value[24]), .Q(h_value[24]), .QN( ));
Q_FDP1 \h_value_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_h_value[23]), .Q(h_value[23]), .QN( ));
Q_FDP1 \h_value_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_h_value[22]), .Q(h_value[22]), .QN( ));
Q_FDP1 \h_value_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_h_value[21]), .Q(h_value[21]), .QN( ));
Q_FDP1 \h_value_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_h_value[20]), .Q(h_value[20]), .QN( ));
Q_FDP1 \h_value_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_h_value[19]), .Q(h_value[19]), .QN( ));
Q_FDP1 \h_value_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_h_value[18]), .Q(h_value[18]), .QN( ));
Q_FDP1 \h_value_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_h_value[17]), .Q(h_value[17]), .QN( ));
Q_FDP1 \h_value_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_h_value[16]), .Q(h_value[16]), .QN( ));
Q_FDP1 \h_value_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_h_value[15]), .Q(h_value[15]), .QN( ));
Q_FDP1 \h_value_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_h_value[14]), .Q(h_value[14]), .QN( ));
Q_FDP1 \h_value_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_h_value[13]), .Q(h_value[13]), .QN( ));
Q_FDP1 \h_value_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_h_value[12]), .Q(h_value[12]), .QN( ));
Q_FDP1 \h_value_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_h_value[11]), .Q(h_value[11]), .QN( ));
Q_FDP1 \h_value_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_h_value[10]), .Q(h_value[10]), .QN( ));
Q_FDP1 \h_value_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_h_value[9]), .Q(h_value[9]), .QN( ));
Q_FDP1 \h_value_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_h_value[8]), .Q(h_value[8]), .QN( ));
Q_FDP1 \h_value_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_h_value[7]), .Q(h_value[7]), .QN( ));
Q_FDP1 \h_value_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_h_value[6]), .Q(h_value[6]), .QN( ));
Q_FDP1 \h_value_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_h_value[5]), .Q(h_value[5]), .QN( ));
Q_FDP1 \h_value_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_h_value[4]), .Q(h_value[4]), .QN( ));
Q_FDP1 \h_value_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_h_value[3]), .Q(h_value[3]), .QN( ));
Q_FDP1 \h_value_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_h_value[2]), .Q(h_value[2]), .QN( ));
Q_FDP1 \h_value_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_h_value[1]), .Q(h_value[1]), .QN( ));
Q_FDP1 \h_value_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_h_value[0]), .Q(h_value[0]), .QN( ));
Q_FDP1 \auth_tag_REG[127] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[127]), .Q(auth_tag[127]), .QN( ));
Q_FDP1 \auth_tag_REG[126] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[126]), .Q(auth_tag[126]), .QN( ));
Q_FDP1 \auth_tag_REG[125] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[125]), .Q(auth_tag[125]), .QN( ));
Q_FDP1 \auth_tag_REG[124] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[124]), .Q(auth_tag[124]), .QN( ));
Q_FDP1 \auth_tag_REG[123] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[123]), .Q(auth_tag[123]), .QN( ));
Q_FDP1 \auth_tag_REG[122] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[122]), .Q(auth_tag[122]), .QN( ));
Q_FDP1 \auth_tag_REG[121] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[121]), .Q(auth_tag[121]), .QN( ));
Q_FDP1 \auth_tag_REG[120] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[120]), .Q(auth_tag[120]), .QN( ));
Q_FDP1 \auth_tag_REG[119] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[119]), .Q(auth_tag[119]), .QN( ));
Q_FDP1 \auth_tag_REG[118] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[118]), .Q(auth_tag[118]), .QN( ));
Q_FDP1 \auth_tag_REG[117] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[117]), .Q(auth_tag[117]), .QN( ));
Q_FDP1 \auth_tag_REG[116] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[116]), .Q(auth_tag[116]), .QN( ));
Q_FDP1 \auth_tag_REG[115] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[115]), .Q(auth_tag[115]), .QN( ));
Q_FDP1 \auth_tag_REG[114] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[114]), .Q(auth_tag[114]), .QN( ));
Q_FDP1 \auth_tag_REG[113] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[113]), .Q(auth_tag[113]), .QN( ));
Q_FDP1 \auth_tag_REG[112] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[112]), .Q(auth_tag[112]), .QN( ));
Q_FDP1 \auth_tag_REG[111] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[111]), .Q(auth_tag[111]), .QN( ));
Q_FDP1 \auth_tag_REG[110] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[110]), .Q(auth_tag[110]), .QN( ));
Q_FDP1 \auth_tag_REG[109] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[109]), .Q(auth_tag[109]), .QN( ));
Q_FDP1 \auth_tag_REG[108] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[108]), .Q(auth_tag[108]), .QN( ));
Q_FDP1 \auth_tag_REG[107] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[107]), .Q(auth_tag[107]), .QN( ));
Q_FDP1 \auth_tag_REG[106] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[106]), .Q(auth_tag[106]), .QN( ));
Q_FDP1 \auth_tag_REG[105] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[105]), .Q(auth_tag[105]), .QN( ));
Q_FDP1 \auth_tag_REG[104] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[104]), .Q(auth_tag[104]), .QN( ));
Q_FDP1 \auth_tag_REG[103] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[103]), .Q(auth_tag[103]), .QN( ));
Q_FDP1 \auth_tag_REG[102] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[102]), .Q(auth_tag[102]), .QN( ));
Q_FDP1 \auth_tag_REG[101] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[101]), .Q(auth_tag[101]), .QN( ));
Q_FDP1 \auth_tag_REG[100] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[100]), .Q(auth_tag[100]), .QN( ));
Q_FDP1 \auth_tag_REG[99] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[99]), .Q(auth_tag[99]), .QN( ));
Q_FDP1 \auth_tag_REG[98] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[98]), .Q(auth_tag[98]), .QN( ));
Q_FDP1 \auth_tag_REG[97] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[97]), .Q(auth_tag[97]), .QN( ));
Q_FDP1 \auth_tag_REG[96] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[96]), .Q(auth_tag[96]), .QN( ));
Q_FDP1 \auth_tag_REG[95] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[95]), .Q(auth_tag[95]), .QN( ));
Q_FDP1 \auth_tag_REG[94] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[94]), .Q(auth_tag[94]), .QN( ));
Q_FDP1 \auth_tag_REG[93] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[93]), .Q(auth_tag[93]), .QN( ));
Q_FDP1 \auth_tag_REG[92] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[92]), .Q(auth_tag[92]), .QN( ));
Q_FDP1 \auth_tag_REG[91] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[91]), .Q(auth_tag[91]), .QN( ));
Q_FDP1 \auth_tag_REG[90] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[90]), .Q(auth_tag[90]), .QN( ));
Q_FDP1 \auth_tag_REG[89] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[89]), .Q(auth_tag[89]), .QN( ));
Q_FDP1 \auth_tag_REG[88] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[88]), .Q(auth_tag[88]), .QN( ));
Q_FDP1 \auth_tag_REG[87] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[87]), .Q(auth_tag[87]), .QN( ));
Q_FDP1 \auth_tag_REG[86] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[86]), .Q(auth_tag[86]), .QN( ));
Q_FDP1 \auth_tag_REG[85] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[85]), .Q(auth_tag[85]), .QN( ));
Q_FDP1 \auth_tag_REG[84] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[84]), .Q(auth_tag[84]), .QN( ));
Q_FDP1 \auth_tag_REG[83] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[83]), .Q(auth_tag[83]), .QN( ));
Q_FDP1 \auth_tag_REG[82] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[82]), .Q(auth_tag[82]), .QN( ));
Q_FDP1 \auth_tag_REG[81] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[81]), .Q(auth_tag[81]), .QN( ));
Q_FDP1 \auth_tag_REG[80] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[80]), .Q(auth_tag[80]), .QN( ));
Q_FDP1 \auth_tag_REG[79] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[79]), .Q(auth_tag[79]), .QN( ));
Q_FDP1 \auth_tag_REG[78] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[78]), .Q(auth_tag[78]), .QN( ));
Q_FDP1 \auth_tag_REG[77] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[77]), .Q(auth_tag[77]), .QN( ));
Q_FDP1 \auth_tag_REG[76] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[76]), .Q(auth_tag[76]), .QN( ));
Q_FDP1 \auth_tag_REG[75] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[75]), .Q(auth_tag[75]), .QN( ));
Q_FDP1 \auth_tag_REG[74] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[74]), .Q(auth_tag[74]), .QN( ));
Q_FDP1 \auth_tag_REG[73] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[73]), .Q(auth_tag[73]), .QN( ));
Q_FDP1 \auth_tag_REG[72] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[72]), .Q(auth_tag[72]), .QN( ));
Q_FDP1 \auth_tag_REG[71] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[71]), .Q(auth_tag[71]), .QN( ));
Q_FDP1 \auth_tag_REG[70] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[70]), .Q(auth_tag[70]), .QN( ));
Q_FDP1 \auth_tag_REG[69] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[69]), .Q(auth_tag[69]), .QN( ));
Q_FDP1 \auth_tag_REG[68] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[68]), .Q(auth_tag[68]), .QN( ));
Q_FDP1 \auth_tag_REG[67] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[67]), .Q(auth_tag[67]), .QN( ));
Q_FDP1 \auth_tag_REG[66] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[66]), .Q(auth_tag[66]), .QN( ));
Q_FDP1 \auth_tag_REG[65] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[65]), .Q(auth_tag[65]), .QN( ));
Q_FDP1 \auth_tag_REG[64] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[64]), .Q(auth_tag[64]), .QN( ));
Q_FDP1 \auth_tag_REG[63] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[63]), .Q(auth_tag[63]), .QN( ));
Q_FDP1 \auth_tag_REG[62] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[62]), .Q(auth_tag[62]), .QN( ));
Q_FDP1 \auth_tag_REG[61] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[61]), .Q(auth_tag[61]), .QN( ));
Q_FDP1 \auth_tag_REG[60] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[60]), .Q(auth_tag[60]), .QN( ));
Q_FDP1 \auth_tag_REG[59] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[59]), .Q(auth_tag[59]), .QN( ));
Q_FDP1 \auth_tag_REG[58] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[58]), .Q(auth_tag[58]), .QN( ));
Q_FDP1 \auth_tag_REG[57] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[57]), .Q(auth_tag[57]), .QN( ));
Q_FDP1 \auth_tag_REG[56] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[56]), .Q(auth_tag[56]), .QN( ));
Q_FDP1 \auth_tag_REG[55] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[55]), .Q(auth_tag[55]), .QN( ));
Q_FDP1 \auth_tag_REG[54] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[54]), .Q(auth_tag[54]), .QN( ));
Q_FDP1 \auth_tag_REG[53] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[53]), .Q(auth_tag[53]), .QN( ));
Q_FDP1 \auth_tag_REG[52] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[52]), .Q(auth_tag[52]), .QN( ));
Q_FDP1 \auth_tag_REG[51] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[51]), .Q(auth_tag[51]), .QN( ));
Q_FDP1 \auth_tag_REG[50] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[50]), .Q(auth_tag[50]), .QN( ));
Q_FDP1 \auth_tag_REG[49] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[49]), .Q(auth_tag[49]), .QN( ));
Q_FDP1 \auth_tag_REG[48] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[48]), .Q(auth_tag[48]), .QN( ));
Q_FDP1 \auth_tag_REG[47] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[47]), .Q(auth_tag[47]), .QN( ));
Q_FDP1 \auth_tag_REG[46] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[46]), .Q(auth_tag[46]), .QN( ));
Q_FDP1 \auth_tag_REG[45] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[45]), .Q(auth_tag[45]), .QN( ));
Q_FDP1 \auth_tag_REG[44] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[44]), .Q(auth_tag[44]), .QN( ));
Q_FDP1 \auth_tag_REG[43] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[43]), .Q(auth_tag[43]), .QN( ));
Q_FDP1 \auth_tag_REG[42] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[42]), .Q(auth_tag[42]), .QN( ));
Q_FDP1 \auth_tag_REG[41] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[41]), .Q(auth_tag[41]), .QN( ));
Q_FDP1 \auth_tag_REG[40] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[40]), .Q(auth_tag[40]), .QN( ));
Q_FDP1 \auth_tag_REG[39] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[39]), .Q(auth_tag[39]), .QN( ));
Q_FDP1 \auth_tag_REG[38] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[38]), .Q(auth_tag[38]), .QN( ));
Q_FDP1 \auth_tag_REG[37] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[37]), .Q(auth_tag[37]), .QN( ));
Q_FDP1 \auth_tag_REG[36] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[36]), .Q(auth_tag[36]), .QN( ));
Q_FDP1 \auth_tag_REG[35] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[35]), .Q(auth_tag[35]), .QN( ));
Q_FDP1 \auth_tag_REG[34] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[34]), .Q(auth_tag[34]), .QN( ));
Q_FDP1 \auth_tag_REG[33] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[33]), .Q(auth_tag[33]), .QN( ));
Q_FDP1 \auth_tag_REG[32] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[32]), .Q(auth_tag[32]), .QN( ));
Q_FDP1 \auth_tag_REG[31] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[31]), .Q(auth_tag[31]), .QN( ));
Q_FDP1 \auth_tag_REG[30] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[30]), .Q(auth_tag[30]), .QN( ));
Q_FDP1 \auth_tag_REG[29] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[29]), .Q(auth_tag[29]), .QN( ));
Q_FDP1 \auth_tag_REG[28] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[28]), .Q(auth_tag[28]), .QN( ));
Q_FDP1 \auth_tag_REG[27] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[27]), .Q(auth_tag[27]), .QN( ));
Q_FDP1 \auth_tag_REG[26] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[26]), .Q(auth_tag[26]), .QN( ));
Q_FDP1 \auth_tag_REG[25] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[25]), .Q(auth_tag[25]), .QN( ));
Q_FDP1 \auth_tag_REG[24] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[24]), .Q(auth_tag[24]), .QN( ));
Q_FDP1 \auth_tag_REG[23] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[23]), .Q(auth_tag[23]), .QN( ));
Q_FDP1 \auth_tag_REG[22] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[22]), .Q(auth_tag[22]), .QN( ));
Q_FDP1 \auth_tag_REG[21] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[21]), .Q(auth_tag[21]), .QN( ));
Q_FDP1 \auth_tag_REG[20] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[20]), .Q(auth_tag[20]), .QN( ));
Q_FDP1 \auth_tag_REG[19] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[19]), .Q(auth_tag[19]), .QN( ));
Q_FDP1 \auth_tag_REG[18] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[18]), .Q(auth_tag[18]), .QN( ));
Q_FDP1 \auth_tag_REG[17] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[17]), .Q(auth_tag[17]), .QN( ));
Q_FDP1 \auth_tag_REG[16] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[16]), .Q(auth_tag[16]), .QN( ));
Q_FDP1 \auth_tag_REG[15] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[15]), .Q(auth_tag[15]), .QN( ));
Q_FDP1 \auth_tag_REG[14] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[14]), .Q(auth_tag[14]), .QN( ));
Q_FDP1 \auth_tag_REG[13] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[13]), .Q(auth_tag[13]), .QN( ));
Q_FDP1 \auth_tag_REG[12] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[12]), .Q(auth_tag[12]), .QN( ));
Q_FDP1 \auth_tag_REG[11] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[11]), .Q(auth_tag[11]), .QN( ));
Q_FDP1 \auth_tag_REG[10] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[10]), .Q(auth_tag[10]), .QN( ));
Q_FDP1 \auth_tag_REG[9] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[9]), .Q(auth_tag[9]), .QN( ));
Q_FDP1 \auth_tag_REG[8] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[8]), .Q(auth_tag[8]), .QN( ));
Q_FDP1 \auth_tag_REG[7] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[7]), .Q(auth_tag[7]), .QN( ));
Q_FDP1 \auth_tag_REG[6] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[6]), .Q(auth_tag[6]), .QN( ));
Q_FDP1 \auth_tag_REG[5] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[5]), .Q(auth_tag[5]), .QN( ));
Q_FDP1 \auth_tag_REG[4] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[4]), .Q(auth_tag[4]), .QN( ));
Q_FDP1 \auth_tag_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[3]), .Q(auth_tag[3]), .QN( ));
Q_FDP1 \auth_tag_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[2]), .Q(auth_tag[2]), .QN( ));
Q_FDP1 \auth_tag_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[1]), .Q(auth_tag[1]), .QN( ));
Q_FDP1 \auth_tag_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_auth_tag[0]), .Q(auth_tag[0]), .QN( ));
Q_FDP1 combo_dek512_REG  ( .CK(clk), .R(rst_n), .D(nxt_combo_dek512), .Q(combo_dek512), .QN( ));
ixc_assign _zz_strnp_0 ( _zy_simnet_gcm_cmdfifo_ack_0_w$, gcm_cmdfifo_ack);
ixc_assign _zz_strnp_1 ( _zy_simnet_gcm_upsizer_stall_1_w$, gcm_upsizer_stall);
ixc_assign _zz_strnp_2 ( _zy_simnet_gcm_tag_data_out_ack_2_w$, 
	gcm_tag_data_out_ack);
ixc_assign _zz_strnp_3 ( _zy_simnet_gcm_kdf_valid_3_w$, gcm_kdf_valid);
ixc_assign _zz_strnp_4 ( _zy_simnet_gcm_kdf_eof_4_w$, gcm_kdf_eof);
ixc_assign_128 _zz_strnp_5 ( _zy_simnet_gcm_kdf_data_5_w$[0:127], 
	gcm_kdf_data[127:0]);
ixc_assign _zz_strnp_6 ( _zy_simnet_gcm_status_data_in_valid_6_w$, 
	gcm_status_data_in_valid);
ixc_assign _zz_strnp_7 ( _zy_simnet_gcm_status_data_in_7_w$, n1648);
ixc_assign_128 _zz_strnp_8 ( _zy_simnet_ciph_in_11_w$[0:127], ciph_in[127:0]);
ixc_assign _zz_strnp_9 ( _zy_simnet_ciph_in_vld_12_w$, ciph_in_vld);
ixc_assign _zz_strnp_10 ( _zy_simnet_ciph_in_last_13_w$, ciph_in_last);
ixc_assign_256 _zz_strnp_11 ( _zy_simnet_key_in_15_w$[0:255], key_in[255:0]);
ixc_assign _zz_strnp_12 ( _zy_simnet_key_in_vld_16_w$, key_in_vld);
ixc_assign _zz_strnp_13 ( _zy_simnet_ciph_out_stall_17_w$, ciph_out_stall);
ixc_assign_132 _zz_strnp_14 ( fifo_out[131:0], 
	_zy_simnet_fifo_out_18_w$[0:131]);
ixc_assign_132 _zz_strnp_15 ( _zy_simnet_fifo_in_21_w$[0:131], fifo_in[131:0]);
ixc_assign _zz_strnp_16 ( _zy_simnet_fifo_in_vld_22_w$, ciph_in_vld);
ixc_assign _zz_strnp_17 ( _zy_simnet_fifo_out_ack_23_w$, ciph_out_vld);
AesSecIStub AesSecI ( .AesCiphOutR( ciph_out[127:0]), .AesCiphOutVldR( 
	ciph_out_vld), .KeyInitStall( key_in_stall), .CiphInStall( 
	ciph_in_stall), .Aes128( _zy_simnet_cio_8), .Aes192( 
	_zy_simnet_cio_9), .Aes256( _zy_simnet_cio_10), .CiphIn( 
	_zy_simnet_ciph_in_11_w$[0:127]), .CiphInVldR( 
	_zy_simnet_ciph_in_vld_12_w$), .CiphInLastR( 
	_zy_simnet_ciph_in_last_13_w$), .EncryptEn( _zy_simnet_cio_14), 
	.KeyIn( _zy_simnet_key_in_15_w$[0:255]), .KeyInitVldR( 
	_zy_simnet_key_in_vld_16_w$), .AesCiphOutStall( 
	_zy_simnet_ciph_out_stall_17_w$), .clk( clk), .rst_n( rst_n));
cr_kme_fifo_xcm55 bypass_fifo ( .fifo_in_stall( fifo_in_stall), .fifo_out( 
	_zy_simnet_fifo_out_18_w$[0:131]), .fifo_out_valid( fifo_out_vld), 
	.fifo_overflow( _zy_simnet_dio_19), .fifo_underflow( 
	_zy_simnet_dio_20), .clk( clk), .rst_n( rst_n), .fifo_in( 
	_zy_simnet_fifo_in_21_w$[0:131]), .fifo_in_valid( 
	_zy_simnet_fifo_in_vld_22_w$), .fifo_out_ack( 
	_zy_simnet_fifo_out_ack_23_w$), .fifo_in_stall_override( 
	_zy_simnet_cio_24));
Q_INV U3103 ( .A(n1245), .Z(n1649));
Q_INV U3104 ( .A(n576), .Z(n1650));
Q_INV U3105 ( .A(n1261), .Z(n1651));
Q_FDP4EP \iv_counter_REG[127] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1262), .Q(iv_counter[127]));
Q_INV U3107 ( .A(rst_n), .Z(n1652));
Q_FDP4EP \iv_counter_REG[126] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1263), .Q(iv_counter[126]));
Q_FDP4EP \iv_counter_REG[125] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1264), .Q(iv_counter[125]));
Q_FDP4EP \iv_counter_REG[124] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1265), .Q(iv_counter[124]));
Q_FDP4EP \iv_counter_REG[123] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1266), .Q(iv_counter[123]));
Q_FDP4EP \iv_counter_REG[122] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1267), .Q(iv_counter[122]));
Q_FDP4EP \iv_counter_REG[121] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1268), .Q(iv_counter[121]));
Q_FDP4EP \iv_counter_REG[120] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1269), .Q(iv_counter[120]));
Q_FDP4EP \iv_counter_REG[119] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1270), .Q(iv_counter[119]));
Q_FDP4EP \iv_counter_REG[118] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1271), .Q(iv_counter[118]));
Q_FDP4EP \iv_counter_REG[117] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1272), .Q(iv_counter[117]));
Q_FDP4EP \iv_counter_REG[116] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1273), .Q(iv_counter[116]));
Q_FDP4EP \iv_counter_REG[115] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1274), .Q(iv_counter[115]));
Q_FDP4EP \iv_counter_REG[114] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1275), .Q(iv_counter[114]));
Q_FDP4EP \iv_counter_REG[113] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1276), .Q(iv_counter[113]));
Q_FDP4EP \iv_counter_REG[112] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1277), .Q(iv_counter[112]));
Q_FDP4EP \iv_counter_REG[111] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1278), .Q(iv_counter[111]));
Q_FDP4EP \iv_counter_REG[110] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1279), .Q(iv_counter[110]));
Q_FDP4EP \iv_counter_REG[109] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1280), .Q(iv_counter[109]));
Q_FDP4EP \iv_counter_REG[108] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1281), .Q(iv_counter[108]));
Q_FDP4EP \iv_counter_REG[107] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1282), .Q(iv_counter[107]));
Q_FDP4EP \iv_counter_REG[106] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1283), .Q(iv_counter[106]));
Q_FDP4EP \iv_counter_REG[105] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1284), .Q(iv_counter[105]));
Q_FDP4EP \iv_counter_REG[104] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1285), .Q(iv_counter[104]));
Q_FDP4EP \iv_counter_REG[103] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1286), .Q(iv_counter[103]));
Q_FDP4EP \iv_counter_REG[102] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1287), .Q(iv_counter[102]));
Q_FDP4EP \iv_counter_REG[101] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1288), .Q(iv_counter[101]));
Q_FDP4EP \iv_counter_REG[100] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1289), .Q(iv_counter[100]));
Q_FDP4EP \iv_counter_REG[99] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1290), .Q(iv_counter[99]));
Q_FDP4EP \iv_counter_REG[98] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1291), .Q(iv_counter[98]));
Q_FDP4EP \iv_counter_REG[97] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1292), .Q(iv_counter[97]));
Q_FDP4EP \iv_counter_REG[96] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1293), .Q(iv_counter[96]));
Q_FDP4EP \iv_counter_REG[95] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1294), .Q(iv_counter[95]));
Q_FDP4EP \iv_counter_REG[94] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1295), .Q(iv_counter[94]));
Q_FDP4EP \iv_counter_REG[93] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1296), .Q(iv_counter[93]));
Q_FDP4EP \iv_counter_REG[92] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1297), .Q(iv_counter[92]));
Q_FDP4EP \iv_counter_REG[91] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1298), .Q(iv_counter[91]));
Q_FDP4EP \iv_counter_REG[90] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1299), .Q(iv_counter[90]));
Q_FDP4EP \iv_counter_REG[89] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1300), .Q(iv_counter[89]));
Q_FDP4EP \iv_counter_REG[88] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1301), .Q(iv_counter[88]));
Q_FDP4EP \iv_counter_REG[87] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1302), .Q(iv_counter[87]));
Q_FDP4EP \iv_counter_REG[86] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1303), .Q(iv_counter[86]));
Q_FDP4EP \iv_counter_REG[85] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1304), .Q(iv_counter[85]));
Q_FDP4EP \iv_counter_REG[84] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1305), .Q(iv_counter[84]));
Q_FDP4EP \iv_counter_REG[83] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1306), .Q(iv_counter[83]));
Q_FDP4EP \iv_counter_REG[82] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1307), .Q(iv_counter[82]));
Q_FDP4EP \iv_counter_REG[81] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1308), .Q(iv_counter[81]));
Q_FDP4EP \iv_counter_REG[80] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1309), .Q(iv_counter[80]));
Q_FDP4EP \iv_counter_REG[79] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1310), .Q(iv_counter[79]));
Q_FDP4EP \iv_counter_REG[78] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1311), .Q(iv_counter[78]));
Q_FDP4EP \iv_counter_REG[77] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1312), .Q(iv_counter[77]));
Q_FDP4EP \iv_counter_REG[76] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1313), .Q(iv_counter[76]));
Q_FDP4EP \iv_counter_REG[75] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1314), .Q(iv_counter[75]));
Q_FDP4EP \iv_counter_REG[74] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1315), .Q(iv_counter[74]));
Q_FDP4EP \iv_counter_REG[73] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1316), .Q(iv_counter[73]));
Q_FDP4EP \iv_counter_REG[72] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1317), .Q(iv_counter[72]));
Q_FDP4EP \iv_counter_REG[71] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1318), .Q(iv_counter[71]));
Q_FDP4EP \iv_counter_REG[70] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1319), .Q(iv_counter[70]));
Q_FDP4EP \iv_counter_REG[69] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1320), .Q(iv_counter[69]));
Q_FDP4EP \iv_counter_REG[68] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1321), .Q(iv_counter[68]));
Q_FDP4EP \iv_counter_REG[67] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1322), .Q(iv_counter[67]));
Q_FDP4EP \iv_counter_REG[66] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1323), .Q(iv_counter[66]));
Q_FDP4EP \iv_counter_REG[65] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1324), .Q(iv_counter[65]));
Q_FDP4EP \iv_counter_REG[64] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1325), .Q(iv_counter[64]));
Q_FDP4EP \iv_counter_REG[63] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1326), .Q(iv_counter[63]));
Q_FDP4EP \iv_counter_REG[62] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1327), .Q(iv_counter[62]));
Q_FDP4EP \iv_counter_REG[61] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1328), .Q(iv_counter[61]));
Q_FDP4EP \iv_counter_REG[60] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1329), .Q(iv_counter[60]));
Q_FDP4EP \iv_counter_REG[59] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1330), .Q(iv_counter[59]));
Q_FDP4EP \iv_counter_REG[58] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1331), .Q(iv_counter[58]));
Q_FDP4EP \iv_counter_REG[57] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1332), .Q(iv_counter[57]));
Q_FDP4EP \iv_counter_REG[56] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1333), .Q(iv_counter[56]));
Q_FDP4EP \iv_counter_REG[55] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1334), .Q(iv_counter[55]));
Q_FDP4EP \iv_counter_REG[54] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1335), .Q(iv_counter[54]));
Q_FDP4EP \iv_counter_REG[53] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1336), .Q(iv_counter[53]));
Q_FDP4EP \iv_counter_REG[52] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1337), .Q(iv_counter[52]));
Q_FDP4EP \iv_counter_REG[51] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1338), .Q(iv_counter[51]));
Q_FDP4EP \iv_counter_REG[50] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1339), .Q(iv_counter[50]));
Q_FDP4EP \iv_counter_REG[49] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1340), .Q(iv_counter[49]));
Q_FDP4EP \iv_counter_REG[48] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1341), .Q(iv_counter[48]));
Q_FDP4EP \iv_counter_REG[47] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1342), .Q(iv_counter[47]));
Q_FDP4EP \iv_counter_REG[46] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1343), .Q(iv_counter[46]));
Q_FDP4EP \iv_counter_REG[45] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1344), .Q(iv_counter[45]));
Q_FDP4EP \iv_counter_REG[44] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1345), .Q(iv_counter[44]));
Q_FDP4EP \iv_counter_REG[43] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1346), .Q(iv_counter[43]));
Q_FDP4EP \iv_counter_REG[42] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1347), .Q(iv_counter[42]));
Q_FDP4EP \iv_counter_REG[41] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1348), .Q(iv_counter[41]));
Q_FDP4EP \iv_counter_REG[40] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1349), .Q(iv_counter[40]));
Q_FDP4EP \iv_counter_REG[39] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1350), .Q(iv_counter[39]));
Q_FDP4EP \iv_counter_REG[38] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1351), .Q(iv_counter[38]));
Q_FDP4EP \iv_counter_REG[37] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1352), .Q(iv_counter[37]));
Q_FDP4EP \iv_counter_REG[36] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1353), .Q(iv_counter[36]));
Q_FDP4EP \iv_counter_REG[35] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1354), .Q(iv_counter[35]));
Q_FDP4EP \iv_counter_REG[34] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1355), .Q(iv_counter[34]));
Q_FDP4EP \iv_counter_REG[33] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1356), .Q(iv_counter[33]));
Q_FDP4EP \iv_counter_REG[32] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1357), .Q(iv_counter[32]));
Q_FDP4EP \iv_counter_REG[31] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1358), .Q(iv_counter[31]));
Q_FDP4EP \iv_counter_REG[30] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1359), .Q(iv_counter[30]));
Q_FDP4EP \iv_counter_REG[29] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1360), .Q(iv_counter[29]));
Q_FDP4EP \iv_counter_REG[28] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1361), .Q(iv_counter[28]));
Q_FDP4EP \iv_counter_REG[27] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1362), .Q(iv_counter[27]));
Q_FDP4EP \iv_counter_REG[26] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1363), .Q(iv_counter[26]));
Q_FDP4EP \iv_counter_REG[25] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1364), .Q(iv_counter[25]));
Q_FDP4EP \iv_counter_REG[24] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1365), .Q(iv_counter[24]));
Q_FDP4EP \iv_counter_REG[23] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1366), .Q(iv_counter[23]));
Q_FDP4EP \iv_counter_REG[22] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1367), .Q(iv_counter[22]));
Q_FDP4EP \iv_counter_REG[21] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1368), .Q(iv_counter[21]));
Q_FDP4EP \iv_counter_REG[20] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1369), .Q(iv_counter[20]));
Q_FDP4EP \iv_counter_REG[19] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1370), .Q(iv_counter[19]));
Q_FDP4EP \iv_counter_REG[18] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1371), .Q(iv_counter[18]));
Q_FDP4EP \iv_counter_REG[17] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1372), .Q(iv_counter[17]));
Q_FDP4EP \iv_counter_REG[16] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1373), .Q(iv_counter[16]));
Q_FDP4EP \iv_counter_REG[15] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1374), .Q(iv_counter[15]));
Q_FDP4EP \iv_counter_REG[14] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1375), .Q(iv_counter[14]));
Q_FDP4EP \iv_counter_REG[13] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1376), .Q(iv_counter[13]));
Q_FDP4EP \iv_counter_REG[12] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1377), .Q(iv_counter[12]));
Q_FDP4EP \iv_counter_REG[11] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1378), .Q(iv_counter[11]));
Q_FDP4EP \iv_counter_REG[10] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1379), .Q(iv_counter[10]));
Q_FDP4EP \iv_counter_REG[9] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1380), .Q(iv_counter[9]));
Q_FDP4EP \iv_counter_REG[8] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1381), .Q(iv_counter[8]));
Q_FDP4EP \iv_counter_REG[7] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1382), .Q(iv_counter[7]));
Q_FDP4EP \iv_counter_REG[6] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1383), .Q(iv_counter[6]));
Q_FDP4EP \iv_counter_REG[5] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1384), .Q(iv_counter[5]));
Q_FDP4EP \iv_counter_REG[4] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1385), .Q(iv_counter[4]));
Q_FDP4EP \iv_counter_REG[3] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1386), .Q(iv_counter[3]));
Q_FDP4EP \iv_counter_REG[2] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1387), .Q(iv_counter[2]));
Q_FDP4EP \iv_counter_REG[1] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1388), .Q(iv_counter[1]));
Q_FDP4EP \iv_counter_REG[0] ( .CK(clk), .CE(n1651), .R(n1652), .D(n1390), .Q(iv_counter[0]));
Q_INV U3235 ( .A(iv_counter[0]), .Z(n1644));
Q_FDP4EP \beat_num_REG[1] ( .CK(clk), .CE(upsizer_gcm_valid), .R(n1652), .D(n1257), .Q(beat_num[1]));
Q_INV U3237 ( .A(beat_num[1]), .Z(n597));
Q_FDP4EP \beat_num_REG[0] ( .CK(clk), .CE(upsizer_gcm_valid), .R(n1652), .D(n1258), .Q(beat_num[0]));
Q_INV U3239 ( .A(beat_num[0]), .Z(n611));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\gcm_status_data_in.tag_mismatch  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\cmdfifo_gcm_cmd.key0  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\cmdfifo_gcm_cmd.key1  (1,0) 1 255 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\cmdfifo_gcm_cmd.iv  (1,0) 1 95 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\cmdfifo_gcm_cmd.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\fifo_in.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\fifo_in.pt  (1,0) 1 127 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\fifo_in.eof  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\fifo_out.op  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\fifo_out.pt  (1,0) 1 127 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\fifo_out.eof  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "11"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "gcm_status_data_in 1 \gcm_status_data_in.tag_mismatch "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "cmdfifo_gcm_cmd 4 \cmdfifo_gcm_cmd.key0  \cmdfifo_gcm_cmd.key1  \cmdfifo_gcm_cmd.iv  \cmdfifo_gcm_cmd.op "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "fifo_in 3 \fifo_in.op  \fifo_in.pt  \fifo_in.eof "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "fifo_out 3 \fifo_out.op  \fifo_out.pt  \fifo_out.eof "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "4"
endmodule
