library ieee, quickturn ;
use ieee.std_logic_1164.all ;
use quickturn.verilog.all ;
entity ixcEcmHold is
  attribute _2_state_: integer;
  attribute upf_always_on : integer;
  attribute upf_always_on of ixcEcmHold: entity is 1 ;
  attribute _2_state_ of ixcEcmHold: entity is 1 ;
end ixcEcmHold ;
