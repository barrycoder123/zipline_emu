
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_regfile_glue ( ckv_cmnd_op, ckv_cmnd_addr, ckv_wr_dat, 
	.ckv_ia_capability( {\ckv_ia_capability.r.part0 [19], 
	\ckv_ia_capability.r.part0 [18], \ckv_ia_capability.r.part0 [17], 
	\ckv_ia_capability.r.part0 [16], \ckv_ia_capability.r.part0 [15], 
	\ckv_ia_capability.r.part0 [14], \ckv_ia_capability.r.part0 [13], 
	\ckv_ia_capability.r.part0 [12], \ckv_ia_capability.r.part0 [11], 
	\ckv_ia_capability.r.part0 [10], \ckv_ia_capability.r.part0 [9], 
	\ckv_ia_capability.r.part0 [8], \ckv_ia_capability.r.part0 [7], 
	\ckv_ia_capability.r.part0 [6], \ckv_ia_capability.r.part0 [5], 
	\ckv_ia_capability.r.part0 [4], \ckv_ia_capability.r.part0 [3], 
	\ckv_ia_capability.r.part0 [2], \ckv_ia_capability.r.part0 [1], 
	\ckv_ia_capability.r.part0 [0]} ), ckv_ia_rdata_part0, 
	ckv_ia_rdata_part1, .ckv_ia_status( {\ckv_ia_status.r.part0 [22], 
	\ckv_ia_status.r.part0 [21], \ckv_ia_status.r.part0 [20], 
	\ckv_ia_status.r.part0 [19], \ckv_ia_status.r.part0 [18], 
	\ckv_ia_status.r.part0 [17], \ckv_ia_status.r.part0 [16], 
	\ckv_ia_status.r.part0 [15], \ckv_ia_status.r.part0 [14], 
	\ckv_ia_status.r.part0 [13], \ckv_ia_status.r.part0 [12], 
	\ckv_ia_status.r.part0 [11], \ckv_ia_status.r.part0 [10], 
	\ckv_ia_status.r.part0 [9], \ckv_ia_status.r.part0 [8], 
	\ckv_ia_status.r.part0 [7], \ckv_ia_status.r.part0 [6], 
	\ckv_ia_status.r.part0 [5], \ckv_ia_status.r.part0 [4], 
	\ckv_ia_status.r.part0 [3], \ckv_ia_status.r.part0 [2], 
	\ckv_ia_status.r.part0 [1], \ckv_ia_status.r.part0 [0]} ), 
	kim_cmnd_op, kim_cmnd_addr, kim_wr_dat, .kim_ia_capability( {
	\kim_ia_capability.r.part0 [19], \kim_ia_capability.r.part0 [18], 
	\kim_ia_capability.r.part0 [17], \kim_ia_capability.r.part0 [16], 
	\kim_ia_capability.r.part0 [15], \kim_ia_capability.r.part0 [14], 
	\kim_ia_capability.r.part0 [13], \kim_ia_capability.r.part0 [12], 
	\kim_ia_capability.r.part0 [11], \kim_ia_capability.r.part0 [10], 
	\kim_ia_capability.r.part0 [9], \kim_ia_capability.r.part0 [8], 
	\kim_ia_capability.r.part0 [7], \kim_ia_capability.r.part0 [6], 
	\kim_ia_capability.r.part0 [5], \kim_ia_capability.r.part0 [4], 
	\kim_ia_capability.r.part0 [3], \kim_ia_capability.r.part0 [2], 
	\kim_ia_capability.r.part0 [1], \kim_ia_capability.r.part0 [0]} ), 
	kim_ia_rdata_part0, kim_ia_rdata_part1, .kim_ia_status( {
	\kim_ia_status.r.part0 [21], \kim_ia_status.r.part0 [20], 
	\kim_ia_status.r.part0 [19], \kim_ia_status.r.part0 [18], 
	\kim_ia_status.r.part0 [17], \kim_ia_status.r.part0 [16], 
	\kim_ia_status.r.part0 [15], \kim_ia_status.r.part0 [14], 
	\kim_ia_status.r.part0 [13], \kim_ia_status.r.part0 [12], 
	\kim_ia_status.r.part0 [11], \kim_ia_status.r.part0 [10], 
	\kim_ia_status.r.part0 [9], \kim_ia_status.r.part0 [8], 
	\kim_ia_status.r.part0 [7], \kim_ia_status.r.part0 [6], 
	\kim_ia_status.r.part0 [5], \kim_ia_status.r.part0 [4], 
	\kim_ia_status.r.part0 [3], \kim_ia_status.r.part0 [2], 
	\kim_ia_status.r.part0 [1], \kim_ia_status.r.part0 [0]} ), 
	engine_sticky_status, disable_ckv_kim_ism_reads, send_kme_ib_beat, 
	debug_kme_ib_tvalid, debug_kme_ib_tlast, debug_kme_ib_tid, 
	debug_kme_ib_tstrb, debug_kme_ib_tuser, debug_kme_ib_tdata, 
	.kme_cceip0_ob_out( {\kme_cceip0_ob_out.tvalid , 
	\kme_cceip0_ob_out.tlast , \kme_cceip0_ob_out.tid [0], 
	\kme_cceip0_ob_out.tstrb [7], \kme_cceip0_ob_out.tstrb [6], 
	\kme_cceip0_ob_out.tstrb [5], \kme_cceip0_ob_out.tstrb [4], 
	\kme_cceip0_ob_out.tstrb [3], \kme_cceip0_ob_out.tstrb [2], 
	\kme_cceip0_ob_out.tstrb [1], \kme_cceip0_ob_out.tstrb [0], 
	\kme_cceip0_ob_out.tuser [7], \kme_cceip0_ob_out.tuser [6], 
	\kme_cceip0_ob_out.tuser [5], \kme_cceip0_ob_out.tuser [4], 
	\kme_cceip0_ob_out.tuser [3], \kme_cceip0_ob_out.tuser [2], 
	\kme_cceip0_ob_out.tuser [1], \kme_cceip0_ob_out.tuser [0], 
	\kme_cceip0_ob_out.tdata [63], \kme_cceip0_ob_out.tdata [62], 
	\kme_cceip0_ob_out.tdata [61], \kme_cceip0_ob_out.tdata [60], 
	\kme_cceip0_ob_out.tdata [59], \kme_cceip0_ob_out.tdata [58], 
	\kme_cceip0_ob_out.tdata [57], \kme_cceip0_ob_out.tdata [56], 
	\kme_cceip0_ob_out.tdata [55], \kme_cceip0_ob_out.tdata [54], 
	\kme_cceip0_ob_out.tdata [53], \kme_cceip0_ob_out.tdata [52], 
	\kme_cceip0_ob_out.tdata [51], \kme_cceip0_ob_out.tdata [50], 
	\kme_cceip0_ob_out.tdata [49], \kme_cceip0_ob_out.tdata [48], 
	\kme_cceip0_ob_out.tdata [47], \kme_cceip0_ob_out.tdata [46], 
	\kme_cceip0_ob_out.tdata [45], \kme_cceip0_ob_out.tdata [44], 
	\kme_cceip0_ob_out.tdata [43], \kme_cceip0_ob_out.tdata [42], 
	\kme_cceip0_ob_out.tdata [41], \kme_cceip0_ob_out.tdata [40], 
	\kme_cceip0_ob_out.tdata [39], \kme_cceip0_ob_out.tdata [38], 
	\kme_cceip0_ob_out.tdata [37], \kme_cceip0_ob_out.tdata [36], 
	\kme_cceip0_ob_out.tdata [35], \kme_cceip0_ob_out.tdata [34], 
	\kme_cceip0_ob_out.tdata [33], \kme_cceip0_ob_out.tdata [32], 
	\kme_cceip0_ob_out.tdata [31], \kme_cceip0_ob_out.tdata [30], 
	\kme_cceip0_ob_out.tdata [29], \kme_cceip0_ob_out.tdata [28], 
	\kme_cceip0_ob_out.tdata [27], \kme_cceip0_ob_out.tdata [26], 
	\kme_cceip0_ob_out.tdata [25], \kme_cceip0_ob_out.tdata [24], 
	\kme_cceip0_ob_out.tdata [23], \kme_cceip0_ob_out.tdata [22], 
	\kme_cceip0_ob_out.tdata [21], \kme_cceip0_ob_out.tdata [20], 
	\kme_cceip0_ob_out.tdata [19], \kme_cceip0_ob_out.tdata [18], 
	\kme_cceip0_ob_out.tdata [17], \kme_cceip0_ob_out.tdata [16], 
	\kme_cceip0_ob_out.tdata [15], \kme_cceip0_ob_out.tdata [14], 
	\kme_cceip0_ob_out.tdata [13], \kme_cceip0_ob_out.tdata [12], 
	\kme_cceip0_ob_out.tdata [11], \kme_cceip0_ob_out.tdata [10], 
	\kme_cceip0_ob_out.tdata [9], \kme_cceip0_ob_out.tdata [8], 
	\kme_cceip0_ob_out.tdata [7], \kme_cceip0_ob_out.tdata [6], 
	\kme_cceip0_ob_out.tdata [5], \kme_cceip0_ob_out.tdata [4], 
	\kme_cceip0_ob_out.tdata [3], \kme_cceip0_ob_out.tdata [2], 
	\kme_cceip0_ob_out.tdata [1], \kme_cceip0_ob_out.tdata [0]} ), 
	.kme_cceip1_ob_out( {\kme_cceip1_ob_out.tvalid , 
	\kme_cceip1_ob_out.tlast , \kme_cceip1_ob_out.tid [0], 
	\kme_cceip1_ob_out.tstrb [7], \kme_cceip1_ob_out.tstrb [6], 
	\kme_cceip1_ob_out.tstrb [5], \kme_cceip1_ob_out.tstrb [4], 
	\kme_cceip1_ob_out.tstrb [3], \kme_cceip1_ob_out.tstrb [2], 
	\kme_cceip1_ob_out.tstrb [1], \kme_cceip1_ob_out.tstrb [0], 
	\kme_cceip1_ob_out.tuser [7], \kme_cceip1_ob_out.tuser [6], 
	\kme_cceip1_ob_out.tuser [5], \kme_cceip1_ob_out.tuser [4], 
	\kme_cceip1_ob_out.tuser [3], \kme_cceip1_ob_out.tuser [2], 
	\kme_cceip1_ob_out.tuser [1], \kme_cceip1_ob_out.tuser [0], 
	\kme_cceip1_ob_out.tdata [63], \kme_cceip1_ob_out.tdata [62], 
	\kme_cceip1_ob_out.tdata [61], \kme_cceip1_ob_out.tdata [60], 
	\kme_cceip1_ob_out.tdata [59], \kme_cceip1_ob_out.tdata [58], 
	\kme_cceip1_ob_out.tdata [57], \kme_cceip1_ob_out.tdata [56], 
	\kme_cceip1_ob_out.tdata [55], \kme_cceip1_ob_out.tdata [54], 
	\kme_cceip1_ob_out.tdata [53], \kme_cceip1_ob_out.tdata [52], 
	\kme_cceip1_ob_out.tdata [51], \kme_cceip1_ob_out.tdata [50], 
	\kme_cceip1_ob_out.tdata [49], \kme_cceip1_ob_out.tdata [48], 
	\kme_cceip1_ob_out.tdata [47], \kme_cceip1_ob_out.tdata [46], 
	\kme_cceip1_ob_out.tdata [45], \kme_cceip1_ob_out.tdata [44], 
	\kme_cceip1_ob_out.tdata [43], \kme_cceip1_ob_out.tdata [42], 
	\kme_cceip1_ob_out.tdata [41], \kme_cceip1_ob_out.tdata [40], 
	\kme_cceip1_ob_out.tdata [39], \kme_cceip1_ob_out.tdata [38], 
	\kme_cceip1_ob_out.tdata [37], \kme_cceip1_ob_out.tdata [36], 
	\kme_cceip1_ob_out.tdata [35], \kme_cceip1_ob_out.tdata [34], 
	\kme_cceip1_ob_out.tdata [33], \kme_cceip1_ob_out.tdata [32], 
	\kme_cceip1_ob_out.tdata [31], \kme_cceip1_ob_out.tdata [30], 
	\kme_cceip1_ob_out.tdata [29], \kme_cceip1_ob_out.tdata [28], 
	\kme_cceip1_ob_out.tdata [27], \kme_cceip1_ob_out.tdata [26], 
	\kme_cceip1_ob_out.tdata [25], \kme_cceip1_ob_out.tdata [24], 
	\kme_cceip1_ob_out.tdata [23], \kme_cceip1_ob_out.tdata [22], 
	\kme_cceip1_ob_out.tdata [21], \kme_cceip1_ob_out.tdata [20], 
	\kme_cceip1_ob_out.tdata [19], \kme_cceip1_ob_out.tdata [18], 
	\kme_cceip1_ob_out.tdata [17], \kme_cceip1_ob_out.tdata [16], 
	\kme_cceip1_ob_out.tdata [15], \kme_cceip1_ob_out.tdata [14], 
	\kme_cceip1_ob_out.tdata [13], \kme_cceip1_ob_out.tdata [12], 
	\kme_cceip1_ob_out.tdata [11], \kme_cceip1_ob_out.tdata [10], 
	\kme_cceip1_ob_out.tdata [9], \kme_cceip1_ob_out.tdata [8], 
	\kme_cceip1_ob_out.tdata [7], \kme_cceip1_ob_out.tdata [6], 
	\kme_cceip1_ob_out.tdata [5], \kme_cceip1_ob_out.tdata [4], 
	\kme_cceip1_ob_out.tdata [3], \kme_cceip1_ob_out.tdata [2], 
	\kme_cceip1_ob_out.tdata [1], \kme_cceip1_ob_out.tdata [0]} ), 
	.kme_cceip2_ob_out( {\kme_cceip2_ob_out.tvalid , 
	\kme_cceip2_ob_out.tlast , \kme_cceip2_ob_out.tid [0], 
	\kme_cceip2_ob_out.tstrb [7], \kme_cceip2_ob_out.tstrb [6], 
	\kme_cceip2_ob_out.tstrb [5], \kme_cceip2_ob_out.tstrb [4], 
	\kme_cceip2_ob_out.tstrb [3], \kme_cceip2_ob_out.tstrb [2], 
	\kme_cceip2_ob_out.tstrb [1], \kme_cceip2_ob_out.tstrb [0], 
	\kme_cceip2_ob_out.tuser [7], \kme_cceip2_ob_out.tuser [6], 
	\kme_cceip2_ob_out.tuser [5], \kme_cceip2_ob_out.tuser [4], 
	\kme_cceip2_ob_out.tuser [3], \kme_cceip2_ob_out.tuser [2], 
	\kme_cceip2_ob_out.tuser [1], \kme_cceip2_ob_out.tuser [0], 
	\kme_cceip2_ob_out.tdata [63], \kme_cceip2_ob_out.tdata [62], 
	\kme_cceip2_ob_out.tdata [61], \kme_cceip2_ob_out.tdata [60], 
	\kme_cceip2_ob_out.tdata [59], \kme_cceip2_ob_out.tdata [58], 
	\kme_cceip2_ob_out.tdata [57], \kme_cceip2_ob_out.tdata [56], 
	\kme_cceip2_ob_out.tdata [55], \kme_cceip2_ob_out.tdata [54], 
	\kme_cceip2_ob_out.tdata [53], \kme_cceip2_ob_out.tdata [52], 
	\kme_cceip2_ob_out.tdata [51], \kme_cceip2_ob_out.tdata [50], 
	\kme_cceip2_ob_out.tdata [49], \kme_cceip2_ob_out.tdata [48], 
	\kme_cceip2_ob_out.tdata [47], \kme_cceip2_ob_out.tdata [46], 
	\kme_cceip2_ob_out.tdata [45], \kme_cceip2_ob_out.tdata [44], 
	\kme_cceip2_ob_out.tdata [43], \kme_cceip2_ob_out.tdata [42], 
	\kme_cceip2_ob_out.tdata [41], \kme_cceip2_ob_out.tdata [40], 
	\kme_cceip2_ob_out.tdata [39], \kme_cceip2_ob_out.tdata [38], 
	\kme_cceip2_ob_out.tdata [37], \kme_cceip2_ob_out.tdata [36], 
	\kme_cceip2_ob_out.tdata [35], \kme_cceip2_ob_out.tdata [34], 
	\kme_cceip2_ob_out.tdata [33], \kme_cceip2_ob_out.tdata [32], 
	\kme_cceip2_ob_out.tdata [31], \kme_cceip2_ob_out.tdata [30], 
	\kme_cceip2_ob_out.tdata [29], \kme_cceip2_ob_out.tdata [28], 
	\kme_cceip2_ob_out.tdata [27], \kme_cceip2_ob_out.tdata [26], 
	\kme_cceip2_ob_out.tdata [25], \kme_cceip2_ob_out.tdata [24], 
	\kme_cceip2_ob_out.tdata [23], \kme_cceip2_ob_out.tdata [22], 
	\kme_cceip2_ob_out.tdata [21], \kme_cceip2_ob_out.tdata [20], 
	\kme_cceip2_ob_out.tdata [19], \kme_cceip2_ob_out.tdata [18], 
	\kme_cceip2_ob_out.tdata [17], \kme_cceip2_ob_out.tdata [16], 
	\kme_cceip2_ob_out.tdata [15], \kme_cceip2_ob_out.tdata [14], 
	\kme_cceip2_ob_out.tdata [13], \kme_cceip2_ob_out.tdata [12], 
	\kme_cceip2_ob_out.tdata [11], \kme_cceip2_ob_out.tdata [10], 
	\kme_cceip2_ob_out.tdata [9], \kme_cceip2_ob_out.tdata [8], 
	\kme_cceip2_ob_out.tdata [7], \kme_cceip2_ob_out.tdata [6], 
	\kme_cceip2_ob_out.tdata [5], \kme_cceip2_ob_out.tdata [4], 
	\kme_cceip2_ob_out.tdata [3], \kme_cceip2_ob_out.tdata [2], 
	\kme_cceip2_ob_out.tdata [1], \kme_cceip2_ob_out.tdata [0]} ), 
	.kme_cceip3_ob_out( {\kme_cceip3_ob_out.tvalid , 
	\kme_cceip3_ob_out.tlast , \kme_cceip3_ob_out.tid [0], 
	\kme_cceip3_ob_out.tstrb [7], \kme_cceip3_ob_out.tstrb [6], 
	\kme_cceip3_ob_out.tstrb [5], \kme_cceip3_ob_out.tstrb [4], 
	\kme_cceip3_ob_out.tstrb [3], \kme_cceip3_ob_out.tstrb [2], 
	\kme_cceip3_ob_out.tstrb [1], \kme_cceip3_ob_out.tstrb [0], 
	\kme_cceip3_ob_out.tuser [7], \kme_cceip3_ob_out.tuser [6], 
	\kme_cceip3_ob_out.tuser [5], \kme_cceip3_ob_out.tuser [4], 
	\kme_cceip3_ob_out.tuser [3], \kme_cceip3_ob_out.tuser [2], 
	\kme_cceip3_ob_out.tuser [1], \kme_cceip3_ob_out.tuser [0], 
	\kme_cceip3_ob_out.tdata [63], \kme_cceip3_ob_out.tdata [62], 
	\kme_cceip3_ob_out.tdata [61], \kme_cceip3_ob_out.tdata [60], 
	\kme_cceip3_ob_out.tdata [59], \kme_cceip3_ob_out.tdata [58], 
	\kme_cceip3_ob_out.tdata [57], \kme_cceip3_ob_out.tdata [56], 
	\kme_cceip3_ob_out.tdata [55], \kme_cceip3_ob_out.tdata [54], 
	\kme_cceip3_ob_out.tdata [53], \kme_cceip3_ob_out.tdata [52], 
	\kme_cceip3_ob_out.tdata [51], \kme_cceip3_ob_out.tdata [50], 
	\kme_cceip3_ob_out.tdata [49], \kme_cceip3_ob_out.tdata [48], 
	\kme_cceip3_ob_out.tdata [47], \kme_cceip3_ob_out.tdata [46], 
	\kme_cceip3_ob_out.tdata [45], \kme_cceip3_ob_out.tdata [44], 
	\kme_cceip3_ob_out.tdata [43], \kme_cceip3_ob_out.tdata [42], 
	\kme_cceip3_ob_out.tdata [41], \kme_cceip3_ob_out.tdata [40], 
	\kme_cceip3_ob_out.tdata [39], \kme_cceip3_ob_out.tdata [38], 
	\kme_cceip3_ob_out.tdata [37], \kme_cceip3_ob_out.tdata [36], 
	\kme_cceip3_ob_out.tdata [35], \kme_cceip3_ob_out.tdata [34], 
	\kme_cceip3_ob_out.tdata [33], \kme_cceip3_ob_out.tdata [32], 
	\kme_cceip3_ob_out.tdata [31], \kme_cceip3_ob_out.tdata [30], 
	\kme_cceip3_ob_out.tdata [29], \kme_cceip3_ob_out.tdata [28], 
	\kme_cceip3_ob_out.tdata [27], \kme_cceip3_ob_out.tdata [26], 
	\kme_cceip3_ob_out.tdata [25], \kme_cceip3_ob_out.tdata [24], 
	\kme_cceip3_ob_out.tdata [23], \kme_cceip3_ob_out.tdata [22], 
	\kme_cceip3_ob_out.tdata [21], \kme_cceip3_ob_out.tdata [20], 
	\kme_cceip3_ob_out.tdata [19], \kme_cceip3_ob_out.tdata [18], 
	\kme_cceip3_ob_out.tdata [17], \kme_cceip3_ob_out.tdata [16], 
	\kme_cceip3_ob_out.tdata [15], \kme_cceip3_ob_out.tdata [14], 
	\kme_cceip3_ob_out.tdata [13], \kme_cceip3_ob_out.tdata [12], 
	\kme_cceip3_ob_out.tdata [11], \kme_cceip3_ob_out.tdata [10], 
	\kme_cceip3_ob_out.tdata [9], \kme_cceip3_ob_out.tdata [8], 
	\kme_cceip3_ob_out.tdata [7], \kme_cceip3_ob_out.tdata [6], 
	\kme_cceip3_ob_out.tdata [5], \kme_cceip3_ob_out.tdata [4], 
	\kme_cceip3_ob_out.tdata [3], \kme_cceip3_ob_out.tdata [2], 
	\kme_cceip3_ob_out.tdata [1], \kme_cceip3_ob_out.tdata [0]} ), 
	.kme_cddip0_ob_out( {\kme_cddip0_ob_out.tvalid , 
	\kme_cddip0_ob_out.tlast , \kme_cddip0_ob_out.tid [0], 
	\kme_cddip0_ob_out.tstrb [7], \kme_cddip0_ob_out.tstrb [6], 
	\kme_cddip0_ob_out.tstrb [5], \kme_cddip0_ob_out.tstrb [4], 
	\kme_cddip0_ob_out.tstrb [3], \kme_cddip0_ob_out.tstrb [2], 
	\kme_cddip0_ob_out.tstrb [1], \kme_cddip0_ob_out.tstrb [0], 
	\kme_cddip0_ob_out.tuser [7], \kme_cddip0_ob_out.tuser [6], 
	\kme_cddip0_ob_out.tuser [5], \kme_cddip0_ob_out.tuser [4], 
	\kme_cddip0_ob_out.tuser [3], \kme_cddip0_ob_out.tuser [2], 
	\kme_cddip0_ob_out.tuser [1], \kme_cddip0_ob_out.tuser [0], 
	\kme_cddip0_ob_out.tdata [63], \kme_cddip0_ob_out.tdata [62], 
	\kme_cddip0_ob_out.tdata [61], \kme_cddip0_ob_out.tdata [60], 
	\kme_cddip0_ob_out.tdata [59], \kme_cddip0_ob_out.tdata [58], 
	\kme_cddip0_ob_out.tdata [57], \kme_cddip0_ob_out.tdata [56], 
	\kme_cddip0_ob_out.tdata [55], \kme_cddip0_ob_out.tdata [54], 
	\kme_cddip0_ob_out.tdata [53], \kme_cddip0_ob_out.tdata [52], 
	\kme_cddip0_ob_out.tdata [51], \kme_cddip0_ob_out.tdata [50], 
	\kme_cddip0_ob_out.tdata [49], \kme_cddip0_ob_out.tdata [48], 
	\kme_cddip0_ob_out.tdata [47], \kme_cddip0_ob_out.tdata [46], 
	\kme_cddip0_ob_out.tdata [45], \kme_cddip0_ob_out.tdata [44], 
	\kme_cddip0_ob_out.tdata [43], \kme_cddip0_ob_out.tdata [42], 
	\kme_cddip0_ob_out.tdata [41], \kme_cddip0_ob_out.tdata [40], 
	\kme_cddip0_ob_out.tdata [39], \kme_cddip0_ob_out.tdata [38], 
	\kme_cddip0_ob_out.tdata [37], \kme_cddip0_ob_out.tdata [36], 
	\kme_cddip0_ob_out.tdata [35], \kme_cddip0_ob_out.tdata [34], 
	\kme_cddip0_ob_out.tdata [33], \kme_cddip0_ob_out.tdata [32], 
	\kme_cddip0_ob_out.tdata [31], \kme_cddip0_ob_out.tdata [30], 
	\kme_cddip0_ob_out.tdata [29], \kme_cddip0_ob_out.tdata [28], 
	\kme_cddip0_ob_out.tdata [27], \kme_cddip0_ob_out.tdata [26], 
	\kme_cddip0_ob_out.tdata [25], \kme_cddip0_ob_out.tdata [24], 
	\kme_cddip0_ob_out.tdata [23], \kme_cddip0_ob_out.tdata [22], 
	\kme_cddip0_ob_out.tdata [21], \kme_cddip0_ob_out.tdata [20], 
	\kme_cddip0_ob_out.tdata [19], \kme_cddip0_ob_out.tdata [18], 
	\kme_cddip0_ob_out.tdata [17], \kme_cddip0_ob_out.tdata [16], 
	\kme_cddip0_ob_out.tdata [15], \kme_cddip0_ob_out.tdata [14], 
	\kme_cddip0_ob_out.tdata [13], \kme_cddip0_ob_out.tdata [12], 
	\kme_cddip0_ob_out.tdata [11], \kme_cddip0_ob_out.tdata [10], 
	\kme_cddip0_ob_out.tdata [9], \kme_cddip0_ob_out.tdata [8], 
	\kme_cddip0_ob_out.tdata [7], \kme_cddip0_ob_out.tdata [6], 
	\kme_cddip0_ob_out.tdata [5], \kme_cddip0_ob_out.tdata [4], 
	\kme_cddip0_ob_out.tdata [3], \kme_cddip0_ob_out.tdata [2], 
	\kme_cddip0_ob_out.tdata [1], \kme_cddip0_ob_out.tdata [0]} ), 
	.kme_cddip1_ob_out( {\kme_cddip1_ob_out.tvalid , 
	\kme_cddip1_ob_out.tlast , \kme_cddip1_ob_out.tid [0], 
	\kme_cddip1_ob_out.tstrb [7], \kme_cddip1_ob_out.tstrb [6], 
	\kme_cddip1_ob_out.tstrb [5], \kme_cddip1_ob_out.tstrb [4], 
	\kme_cddip1_ob_out.tstrb [3], \kme_cddip1_ob_out.tstrb [2], 
	\kme_cddip1_ob_out.tstrb [1], \kme_cddip1_ob_out.tstrb [0], 
	\kme_cddip1_ob_out.tuser [7], \kme_cddip1_ob_out.tuser [6], 
	\kme_cddip1_ob_out.tuser [5], \kme_cddip1_ob_out.tuser [4], 
	\kme_cddip1_ob_out.tuser [3], \kme_cddip1_ob_out.tuser [2], 
	\kme_cddip1_ob_out.tuser [1], \kme_cddip1_ob_out.tuser [0], 
	\kme_cddip1_ob_out.tdata [63], \kme_cddip1_ob_out.tdata [62], 
	\kme_cddip1_ob_out.tdata [61], \kme_cddip1_ob_out.tdata [60], 
	\kme_cddip1_ob_out.tdata [59], \kme_cddip1_ob_out.tdata [58], 
	\kme_cddip1_ob_out.tdata [57], \kme_cddip1_ob_out.tdata [56], 
	\kme_cddip1_ob_out.tdata [55], \kme_cddip1_ob_out.tdata [54], 
	\kme_cddip1_ob_out.tdata [53], \kme_cddip1_ob_out.tdata [52], 
	\kme_cddip1_ob_out.tdata [51], \kme_cddip1_ob_out.tdata [50], 
	\kme_cddip1_ob_out.tdata [49], \kme_cddip1_ob_out.tdata [48], 
	\kme_cddip1_ob_out.tdata [47], \kme_cddip1_ob_out.tdata [46], 
	\kme_cddip1_ob_out.tdata [45], \kme_cddip1_ob_out.tdata [44], 
	\kme_cddip1_ob_out.tdata [43], \kme_cddip1_ob_out.tdata [42], 
	\kme_cddip1_ob_out.tdata [41], \kme_cddip1_ob_out.tdata [40], 
	\kme_cddip1_ob_out.tdata [39], \kme_cddip1_ob_out.tdata [38], 
	\kme_cddip1_ob_out.tdata [37], \kme_cddip1_ob_out.tdata [36], 
	\kme_cddip1_ob_out.tdata [35], \kme_cddip1_ob_out.tdata [34], 
	\kme_cddip1_ob_out.tdata [33], \kme_cddip1_ob_out.tdata [32], 
	\kme_cddip1_ob_out.tdata [31], \kme_cddip1_ob_out.tdata [30], 
	\kme_cddip1_ob_out.tdata [29], \kme_cddip1_ob_out.tdata [28], 
	\kme_cddip1_ob_out.tdata [27], \kme_cddip1_ob_out.tdata [26], 
	\kme_cddip1_ob_out.tdata [25], \kme_cddip1_ob_out.tdata [24], 
	\kme_cddip1_ob_out.tdata [23], \kme_cddip1_ob_out.tdata [22], 
	\kme_cddip1_ob_out.tdata [21], \kme_cddip1_ob_out.tdata [20], 
	\kme_cddip1_ob_out.tdata [19], \kme_cddip1_ob_out.tdata [18], 
	\kme_cddip1_ob_out.tdata [17], \kme_cddip1_ob_out.tdata [16], 
	\kme_cddip1_ob_out.tdata [15], \kme_cddip1_ob_out.tdata [14], 
	\kme_cddip1_ob_out.tdata [13], \kme_cddip1_ob_out.tdata [12], 
	\kme_cddip1_ob_out.tdata [11], \kme_cddip1_ob_out.tdata [10], 
	\kme_cddip1_ob_out.tdata [9], \kme_cddip1_ob_out.tdata [8], 
	\kme_cddip1_ob_out.tdata [7], \kme_cddip1_ob_out.tdata [6], 
	\kme_cddip1_ob_out.tdata [5], \kme_cddip1_ob_out.tdata [4], 
	\kme_cddip1_ob_out.tdata [3], \kme_cddip1_ob_out.tdata [2], 
	\kme_cddip1_ob_out.tdata [1], \kme_cddip1_ob_out.tdata [0]} ), 
	.kme_cddip2_ob_out( {\kme_cddip2_ob_out.tvalid , 
	\kme_cddip2_ob_out.tlast , \kme_cddip2_ob_out.tid [0], 
	\kme_cddip2_ob_out.tstrb [7], \kme_cddip2_ob_out.tstrb [6], 
	\kme_cddip2_ob_out.tstrb [5], \kme_cddip2_ob_out.tstrb [4], 
	\kme_cddip2_ob_out.tstrb [3], \kme_cddip2_ob_out.tstrb [2], 
	\kme_cddip2_ob_out.tstrb [1], \kme_cddip2_ob_out.tstrb [0], 
	\kme_cddip2_ob_out.tuser [7], \kme_cddip2_ob_out.tuser [6], 
	\kme_cddip2_ob_out.tuser [5], \kme_cddip2_ob_out.tuser [4], 
	\kme_cddip2_ob_out.tuser [3], \kme_cddip2_ob_out.tuser [2], 
	\kme_cddip2_ob_out.tuser [1], \kme_cddip2_ob_out.tuser [0], 
	\kme_cddip2_ob_out.tdata [63], \kme_cddip2_ob_out.tdata [62], 
	\kme_cddip2_ob_out.tdata [61], \kme_cddip2_ob_out.tdata [60], 
	\kme_cddip2_ob_out.tdata [59], \kme_cddip2_ob_out.tdata [58], 
	\kme_cddip2_ob_out.tdata [57], \kme_cddip2_ob_out.tdata [56], 
	\kme_cddip2_ob_out.tdata [55], \kme_cddip2_ob_out.tdata [54], 
	\kme_cddip2_ob_out.tdata [53], \kme_cddip2_ob_out.tdata [52], 
	\kme_cddip2_ob_out.tdata [51], \kme_cddip2_ob_out.tdata [50], 
	\kme_cddip2_ob_out.tdata [49], \kme_cddip2_ob_out.tdata [48], 
	\kme_cddip2_ob_out.tdata [47], \kme_cddip2_ob_out.tdata [46], 
	\kme_cddip2_ob_out.tdata [45], \kme_cddip2_ob_out.tdata [44], 
	\kme_cddip2_ob_out.tdata [43], \kme_cddip2_ob_out.tdata [42], 
	\kme_cddip2_ob_out.tdata [41], \kme_cddip2_ob_out.tdata [40], 
	\kme_cddip2_ob_out.tdata [39], \kme_cddip2_ob_out.tdata [38], 
	\kme_cddip2_ob_out.tdata [37], \kme_cddip2_ob_out.tdata [36], 
	\kme_cddip2_ob_out.tdata [35], \kme_cddip2_ob_out.tdata [34], 
	\kme_cddip2_ob_out.tdata [33], \kme_cddip2_ob_out.tdata [32], 
	\kme_cddip2_ob_out.tdata [31], \kme_cddip2_ob_out.tdata [30], 
	\kme_cddip2_ob_out.tdata [29], \kme_cddip2_ob_out.tdata [28], 
	\kme_cddip2_ob_out.tdata [27], \kme_cddip2_ob_out.tdata [26], 
	\kme_cddip2_ob_out.tdata [25], \kme_cddip2_ob_out.tdata [24], 
	\kme_cddip2_ob_out.tdata [23], \kme_cddip2_ob_out.tdata [22], 
	\kme_cddip2_ob_out.tdata [21], \kme_cddip2_ob_out.tdata [20], 
	\kme_cddip2_ob_out.tdata [19], \kme_cddip2_ob_out.tdata [18], 
	\kme_cddip2_ob_out.tdata [17], \kme_cddip2_ob_out.tdata [16], 
	\kme_cddip2_ob_out.tdata [15], \kme_cddip2_ob_out.tdata [14], 
	\kme_cddip2_ob_out.tdata [13], \kme_cddip2_ob_out.tdata [12], 
	\kme_cddip2_ob_out.tdata [11], \kme_cddip2_ob_out.tdata [10], 
	\kme_cddip2_ob_out.tdata [9], \kme_cddip2_ob_out.tdata [8], 
	\kme_cddip2_ob_out.tdata [7], \kme_cddip2_ob_out.tdata [6], 
	\kme_cddip2_ob_out.tdata [5], \kme_cddip2_ob_out.tdata [4], 
	\kme_cddip2_ob_out.tdata [3], \kme_cddip2_ob_out.tdata [2], 
	\kme_cddip2_ob_out.tdata [1], \kme_cddip2_ob_out.tdata [0]} ), 
	.kme_cddip3_ob_out( {\kme_cddip3_ob_out.tvalid , 
	\kme_cddip3_ob_out.tlast , \kme_cddip3_ob_out.tid [0], 
	\kme_cddip3_ob_out.tstrb [7], \kme_cddip3_ob_out.tstrb [6], 
	\kme_cddip3_ob_out.tstrb [5], \kme_cddip3_ob_out.tstrb [4], 
	\kme_cddip3_ob_out.tstrb [3], \kme_cddip3_ob_out.tstrb [2], 
	\kme_cddip3_ob_out.tstrb [1], \kme_cddip3_ob_out.tstrb [0], 
	\kme_cddip3_ob_out.tuser [7], \kme_cddip3_ob_out.tuser [6], 
	\kme_cddip3_ob_out.tuser [5], \kme_cddip3_ob_out.tuser [4], 
	\kme_cddip3_ob_out.tuser [3], \kme_cddip3_ob_out.tuser [2], 
	\kme_cddip3_ob_out.tuser [1], \kme_cddip3_ob_out.tuser [0], 
	\kme_cddip3_ob_out.tdata [63], \kme_cddip3_ob_out.tdata [62], 
	\kme_cddip3_ob_out.tdata [61], \kme_cddip3_ob_out.tdata [60], 
	\kme_cddip3_ob_out.tdata [59], \kme_cddip3_ob_out.tdata [58], 
	\kme_cddip3_ob_out.tdata [57], \kme_cddip3_ob_out.tdata [56], 
	\kme_cddip3_ob_out.tdata [55], \kme_cddip3_ob_out.tdata [54], 
	\kme_cddip3_ob_out.tdata [53], \kme_cddip3_ob_out.tdata [52], 
	\kme_cddip3_ob_out.tdata [51], \kme_cddip3_ob_out.tdata [50], 
	\kme_cddip3_ob_out.tdata [49], \kme_cddip3_ob_out.tdata [48], 
	\kme_cddip3_ob_out.tdata [47], \kme_cddip3_ob_out.tdata [46], 
	\kme_cddip3_ob_out.tdata [45], \kme_cddip3_ob_out.tdata [44], 
	\kme_cddip3_ob_out.tdata [43], \kme_cddip3_ob_out.tdata [42], 
	\kme_cddip3_ob_out.tdata [41], \kme_cddip3_ob_out.tdata [40], 
	\kme_cddip3_ob_out.tdata [39], \kme_cddip3_ob_out.tdata [38], 
	\kme_cddip3_ob_out.tdata [37], \kme_cddip3_ob_out.tdata [36], 
	\kme_cddip3_ob_out.tdata [35], \kme_cddip3_ob_out.tdata [34], 
	\kme_cddip3_ob_out.tdata [33], \kme_cddip3_ob_out.tdata [32], 
	\kme_cddip3_ob_out.tdata [31], \kme_cddip3_ob_out.tdata [30], 
	\kme_cddip3_ob_out.tdata [29], \kme_cddip3_ob_out.tdata [28], 
	\kme_cddip3_ob_out.tdata [27], \kme_cddip3_ob_out.tdata [26], 
	\kme_cddip3_ob_out.tdata [25], \kme_cddip3_ob_out.tdata [24], 
	\kme_cddip3_ob_out.tdata [23], \kme_cddip3_ob_out.tdata [22], 
	\kme_cddip3_ob_out.tdata [21], \kme_cddip3_ob_out.tdata [20], 
	\kme_cddip3_ob_out.tdata [19], \kme_cddip3_ob_out.tdata [18], 
	\kme_cddip3_ob_out.tdata [17], \kme_cddip3_ob_out.tdata [16], 
	\kme_cddip3_ob_out.tdata [15], \kme_cddip3_ob_out.tdata [14], 
	\kme_cddip3_ob_out.tdata [13], \kme_cddip3_ob_out.tdata [12], 
	\kme_cddip3_ob_out.tdata [11], \kme_cddip3_ob_out.tdata [10], 
	\kme_cddip3_ob_out.tdata [9], \kme_cddip3_ob_out.tdata [8], 
	\kme_cddip3_ob_out.tdata [7], \kme_cddip3_ob_out.tdata [6], 
	\kme_cddip3_ob_out.tdata [5], \kme_cddip3_ob_out.tdata [4], 
	\kme_cddip3_ob_out.tdata [3], \kme_cddip3_ob_out.tdata [2], 
	\kme_cddip3_ob_out.tdata [1], \kme_cddip3_ob_out.tdata [0]} ), 
	cceip_encrypt_bimc_isync, cceip_encrypt_bimc_idat, 
	cceip_validate_bimc_isync, cceip_validate_bimc_idat, 
	cddip_decrypt_bimc_isync, cddip_decrypt_bimc_idat, axi_bimc_isync, 
	axi_bimc_idat, axi_term_bimc_isync, axi_term_bimc_idat, clk, rst_n, 
	ckv_stat_code, ckv_stat_datawords, ckv_stat_addr, 
	ckv_capability_type, ckv_capability_lst, ckv_rd_dat, .o_ckv_ia_config( {
	\o_ckv_ia_config.r.part0 [18], \o_ckv_ia_config.r.part0 [17], 
	\o_ckv_ia_config.r.part0 [16], \o_ckv_ia_config.r.part0 [15], 
	\o_ckv_ia_config.r.part0 [14], \o_ckv_ia_config.r.part0 [13], 
	\o_ckv_ia_config.r.part0 [12], \o_ckv_ia_config.r.part0 [11], 
	\o_ckv_ia_config.r.part0 [10], \o_ckv_ia_config.r.part0 [9], 
	\o_ckv_ia_config.r.part0 [8], \o_ckv_ia_config.r.part0 [7], 
	\o_ckv_ia_config.r.part0 [6], \o_ckv_ia_config.r.part0 [5], 
	\o_ckv_ia_config.r.part0 [4], \o_ckv_ia_config.r.part0 [3], 
	\o_ckv_ia_config.r.part0 [2], \o_ckv_ia_config.r.part0 [1], 
	\o_ckv_ia_config.r.part0 [0]} ), o_ckv_ia_wdata_part0, 
	o_ckv_ia_wdata_part1, kim_stat_code, kim_stat_datawords, 
	kim_stat_addr, kim_capability_type, kim_capability_lst, kim_rd_dat, 
	.o_kim_ia_config( {\o_kim_ia_config.r.part0 [17], 
	\o_kim_ia_config.r.part0 [16], \o_kim_ia_config.r.part0 [15], 
	\o_kim_ia_config.r.part0 [14], \o_kim_ia_config.r.part0 [13], 
	\o_kim_ia_config.r.part0 [12], \o_kim_ia_config.r.part0 [11], 
	\o_kim_ia_config.r.part0 [10], \o_kim_ia_config.r.part0 [9], 
	\o_kim_ia_config.r.part0 [8], \o_kim_ia_config.r.part0 [7], 
	\o_kim_ia_config.r.part0 [6], \o_kim_ia_config.r.part0 [5], 
	\o_kim_ia_config.r.part0 [4], \o_kim_ia_config.r.part0 [3], 
	\o_kim_ia_config.r.part0 [2], \o_kim_ia_config.r.part0 [1], 
	\o_kim_ia_config.r.part0 [0]} ), o_kim_ia_wdata_part0, 
	o_kim_ia_wdata_part1, set_rsm_is_backpressuring, wr_stb, wr_data, 
	reg_addr, o_engine_sticky_status, o_disable_ckv_kim_ism_reads, 
	o_send_kme_ib_beat, .cceip0_out_ia_wdata( {
	\cceip0_out_ia_wdata.r.part2 [31], \cceip0_out_ia_wdata.r.part2 [30], 
	\cceip0_out_ia_wdata.r.part2 [29], \cceip0_out_ia_wdata.r.part2 [28], 
	\cceip0_out_ia_wdata.r.part2 [27], \cceip0_out_ia_wdata.r.part2 [26], 
	\cceip0_out_ia_wdata.r.part2 [25], \cceip0_out_ia_wdata.r.part2 [24], 
	\cceip0_out_ia_wdata.r.part2 [23], \cceip0_out_ia_wdata.r.part2 [22], 
	\cceip0_out_ia_wdata.r.part2 [21], \cceip0_out_ia_wdata.r.part2 [20], 
	\cceip0_out_ia_wdata.r.part2 [19], \cceip0_out_ia_wdata.r.part2 [18], 
	\cceip0_out_ia_wdata.r.part2 [17], \cceip0_out_ia_wdata.r.part2 [16], 
	\cceip0_out_ia_wdata.r.part2 [15], \cceip0_out_ia_wdata.r.part2 [14], 
	\cceip0_out_ia_wdata.r.part2 [13], \cceip0_out_ia_wdata.r.part2 [12], 
	\cceip0_out_ia_wdata.r.part2 [11], \cceip0_out_ia_wdata.r.part2 [10], 
	\cceip0_out_ia_wdata.r.part2 [9], \cceip0_out_ia_wdata.r.part2 [8], 
	\cceip0_out_ia_wdata.r.part2 [7], \cceip0_out_ia_wdata.r.part2 [6], 
	\cceip0_out_ia_wdata.r.part2 [5], \cceip0_out_ia_wdata.r.part2 [4], 
	\cceip0_out_ia_wdata.r.part2 [3], \cceip0_out_ia_wdata.r.part2 [2], 
	\cceip0_out_ia_wdata.r.part2 [1], \cceip0_out_ia_wdata.r.part2 [0], 
	\cceip0_out_ia_wdata.r.part1 [31], \cceip0_out_ia_wdata.r.part1 [30], 
	\cceip0_out_ia_wdata.r.part1 [29], \cceip0_out_ia_wdata.r.part1 [28], 
	\cceip0_out_ia_wdata.r.part1 [27], \cceip0_out_ia_wdata.r.part1 [26], 
	\cceip0_out_ia_wdata.r.part1 [25], \cceip0_out_ia_wdata.r.part1 [24], 
	\cceip0_out_ia_wdata.r.part1 [23], \cceip0_out_ia_wdata.r.part1 [22], 
	\cceip0_out_ia_wdata.r.part1 [21], \cceip0_out_ia_wdata.r.part1 [20], 
	\cceip0_out_ia_wdata.r.part1 [19], \cceip0_out_ia_wdata.r.part1 [18], 
	\cceip0_out_ia_wdata.r.part1 [17], \cceip0_out_ia_wdata.r.part1 [16], 
	\cceip0_out_ia_wdata.r.part1 [15], \cceip0_out_ia_wdata.r.part1 [14], 
	\cceip0_out_ia_wdata.r.part1 [13], \cceip0_out_ia_wdata.r.part1 [12], 
	\cceip0_out_ia_wdata.r.part1 [11], \cceip0_out_ia_wdata.r.part1 [10], 
	\cceip0_out_ia_wdata.r.part1 [9], \cceip0_out_ia_wdata.r.part1 [8], 
	\cceip0_out_ia_wdata.r.part1 [7], \cceip0_out_ia_wdata.r.part1 [6], 
	\cceip0_out_ia_wdata.r.part1 [5], \cceip0_out_ia_wdata.r.part1 [4], 
	\cceip0_out_ia_wdata.r.part1 [3], \cceip0_out_ia_wdata.r.part1 [2], 
	\cceip0_out_ia_wdata.r.part1 [1], \cceip0_out_ia_wdata.r.part1 [0], 
	\cceip0_out_ia_wdata.r.part0 [31], \cceip0_out_ia_wdata.r.part0 [30], 
	\cceip0_out_ia_wdata.r.part0 [29], \cceip0_out_ia_wdata.r.part0 [28], 
	\cceip0_out_ia_wdata.r.part0 [27], \cceip0_out_ia_wdata.r.part0 [26], 
	\cceip0_out_ia_wdata.r.part0 [25], \cceip0_out_ia_wdata.r.part0 [24], 
	\cceip0_out_ia_wdata.r.part0 [23], \cceip0_out_ia_wdata.r.part0 [22], 
	\cceip0_out_ia_wdata.r.part0 [21], \cceip0_out_ia_wdata.r.part0 [20], 
	\cceip0_out_ia_wdata.r.part0 [19], \cceip0_out_ia_wdata.r.part0 [18], 
	\cceip0_out_ia_wdata.r.part0 [17], \cceip0_out_ia_wdata.r.part0 [16], 
	\cceip0_out_ia_wdata.r.part0 [15], \cceip0_out_ia_wdata.r.part0 [14], 
	\cceip0_out_ia_wdata.r.part0 [13], \cceip0_out_ia_wdata.r.part0 [12], 
	\cceip0_out_ia_wdata.r.part0 [11], \cceip0_out_ia_wdata.r.part0 [10], 
	\cceip0_out_ia_wdata.r.part0 [9], \cceip0_out_ia_wdata.r.part0 [8], 
	\cceip0_out_ia_wdata.r.part0 [7], \cceip0_out_ia_wdata.r.part0 [6], 
	\cceip0_out_ia_wdata.r.part0 [5], \cceip0_out_ia_wdata.r.part0 [4], 
	\cceip0_out_ia_wdata.r.part0 [3], \cceip0_out_ia_wdata.r.part0 [2], 
	\cceip0_out_ia_wdata.r.part0 [1], \cceip0_out_ia_wdata.r.part0 [0]} ), 
	debug_kme_ib_tready, .tready_override( {
	\tready_override.r.part0 [8], \tready_override.r.part0 [7], 
	\tready_override.r.part0 [6], \tready_override.r.part0 [5], 
	\tready_override.r.part0 [4], \tready_override.r.part0 [3], 
	\tready_override.r.part0 [2], \tready_override.r.part0 [1], 
	\tready_override.r.part0 [0]} ), .kme_cceip0_ob_out_post( {
	\kme_cceip0_ob_out_post.tvalid , \kme_cceip0_ob_out_post.tlast , 
	\kme_cceip0_ob_out_post.tid [0], \kme_cceip0_ob_out_post.tstrb [7], 
	\kme_cceip0_ob_out_post.tstrb [6], \kme_cceip0_ob_out_post.tstrb [5], 
	\kme_cceip0_ob_out_post.tstrb [4], \kme_cceip0_ob_out_post.tstrb [3], 
	\kme_cceip0_ob_out_post.tstrb [2], \kme_cceip0_ob_out_post.tstrb [1], 
	\kme_cceip0_ob_out_post.tstrb [0], \kme_cceip0_ob_out_post.tuser [7], 
	\kme_cceip0_ob_out_post.tuser [6], \kme_cceip0_ob_out_post.tuser [5], 
	\kme_cceip0_ob_out_post.tuser [4], \kme_cceip0_ob_out_post.tuser [3], 
	\kme_cceip0_ob_out_post.tuser [2], \kme_cceip0_ob_out_post.tuser [1], 
	\kme_cceip0_ob_out_post.tuser [0], 
	\kme_cceip0_ob_out_post.tdata [63], 
	\kme_cceip0_ob_out_post.tdata [62], 
	\kme_cceip0_ob_out_post.tdata [61], 
	\kme_cceip0_ob_out_post.tdata [60], 
	\kme_cceip0_ob_out_post.tdata [59], 
	\kme_cceip0_ob_out_post.tdata [58], 
	\kme_cceip0_ob_out_post.tdata [57], 
	\kme_cceip0_ob_out_post.tdata [56], 
	\kme_cceip0_ob_out_post.tdata [55], 
	\kme_cceip0_ob_out_post.tdata [54], 
	\kme_cceip0_ob_out_post.tdata [53], 
	\kme_cceip0_ob_out_post.tdata [52], 
	\kme_cceip0_ob_out_post.tdata [51], 
	\kme_cceip0_ob_out_post.tdata [50], 
	\kme_cceip0_ob_out_post.tdata [49], 
	\kme_cceip0_ob_out_post.tdata [48], 
	\kme_cceip0_ob_out_post.tdata [47], 
	\kme_cceip0_ob_out_post.tdata [46], 
	\kme_cceip0_ob_out_post.tdata [45], 
	\kme_cceip0_ob_out_post.tdata [44], 
	\kme_cceip0_ob_out_post.tdata [43], 
	\kme_cceip0_ob_out_post.tdata [42], 
	\kme_cceip0_ob_out_post.tdata [41], 
	\kme_cceip0_ob_out_post.tdata [40], 
	\kme_cceip0_ob_out_post.tdata [39], 
	\kme_cceip0_ob_out_post.tdata [38], 
	\kme_cceip0_ob_out_post.tdata [37], 
	\kme_cceip0_ob_out_post.tdata [36], 
	\kme_cceip0_ob_out_post.tdata [35], 
	\kme_cceip0_ob_out_post.tdata [34], 
	\kme_cceip0_ob_out_post.tdata [33], 
	\kme_cceip0_ob_out_post.tdata [32], 
	\kme_cceip0_ob_out_post.tdata [31], 
	\kme_cceip0_ob_out_post.tdata [30], 
	\kme_cceip0_ob_out_post.tdata [29], 
	\kme_cceip0_ob_out_post.tdata [28], 
	\kme_cceip0_ob_out_post.tdata [27], 
	\kme_cceip0_ob_out_post.tdata [26], 
	\kme_cceip0_ob_out_post.tdata [25], 
	\kme_cceip0_ob_out_post.tdata [24], 
	\kme_cceip0_ob_out_post.tdata [23], 
	\kme_cceip0_ob_out_post.tdata [22], 
	\kme_cceip0_ob_out_post.tdata [21], 
	\kme_cceip0_ob_out_post.tdata [20], 
	\kme_cceip0_ob_out_post.tdata [19], 
	\kme_cceip0_ob_out_post.tdata [18], 
	\kme_cceip0_ob_out_post.tdata [17], 
	\kme_cceip0_ob_out_post.tdata [16], 
	\kme_cceip0_ob_out_post.tdata [15], 
	\kme_cceip0_ob_out_post.tdata [14], 
	\kme_cceip0_ob_out_post.tdata [13], 
	\kme_cceip0_ob_out_post.tdata [12], 
	\kme_cceip0_ob_out_post.tdata [11], 
	\kme_cceip0_ob_out_post.tdata [10], 
	\kme_cceip0_ob_out_post.tdata [9], \kme_cceip0_ob_out_post.tdata [8], 
	\kme_cceip0_ob_out_post.tdata [7], \kme_cceip0_ob_out_post.tdata [6], 
	\kme_cceip0_ob_out_post.tdata [5], \kme_cceip0_ob_out_post.tdata [4], 
	\kme_cceip0_ob_out_post.tdata [3], \kme_cceip0_ob_out_post.tdata [2], 
	\kme_cceip0_ob_out_post.tdata [1], \kme_cceip0_ob_out_post.tdata [0]} ), 
	.kme_cceip1_ob_out_post( {\kme_cceip1_ob_out_post.tvalid , 
	\kme_cceip1_ob_out_post.tlast , \kme_cceip1_ob_out_post.tid [0], 
	\kme_cceip1_ob_out_post.tstrb [7], \kme_cceip1_ob_out_post.tstrb [6], 
	\kme_cceip1_ob_out_post.tstrb [5], \kme_cceip1_ob_out_post.tstrb [4], 
	\kme_cceip1_ob_out_post.tstrb [3], \kme_cceip1_ob_out_post.tstrb [2], 
	\kme_cceip1_ob_out_post.tstrb [1], \kme_cceip1_ob_out_post.tstrb [0], 
	\kme_cceip1_ob_out_post.tuser [7], \kme_cceip1_ob_out_post.tuser [6], 
	\kme_cceip1_ob_out_post.tuser [5], \kme_cceip1_ob_out_post.tuser [4], 
	\kme_cceip1_ob_out_post.tuser [3], \kme_cceip1_ob_out_post.tuser [2], 
	\kme_cceip1_ob_out_post.tuser [1], \kme_cceip1_ob_out_post.tuser [0], 
	\kme_cceip1_ob_out_post.tdata [63], 
	\kme_cceip1_ob_out_post.tdata [62], 
	\kme_cceip1_ob_out_post.tdata [61], 
	\kme_cceip1_ob_out_post.tdata [60], 
	\kme_cceip1_ob_out_post.tdata [59], 
	\kme_cceip1_ob_out_post.tdata [58], 
	\kme_cceip1_ob_out_post.tdata [57], 
	\kme_cceip1_ob_out_post.tdata [56], 
	\kme_cceip1_ob_out_post.tdata [55], 
	\kme_cceip1_ob_out_post.tdata [54], 
	\kme_cceip1_ob_out_post.tdata [53], 
	\kme_cceip1_ob_out_post.tdata [52], 
	\kme_cceip1_ob_out_post.tdata [51], 
	\kme_cceip1_ob_out_post.tdata [50], 
	\kme_cceip1_ob_out_post.tdata [49], 
	\kme_cceip1_ob_out_post.tdata [48], 
	\kme_cceip1_ob_out_post.tdata [47], 
	\kme_cceip1_ob_out_post.tdata [46], 
	\kme_cceip1_ob_out_post.tdata [45], 
	\kme_cceip1_ob_out_post.tdata [44], 
	\kme_cceip1_ob_out_post.tdata [43], 
	\kme_cceip1_ob_out_post.tdata [42], 
	\kme_cceip1_ob_out_post.tdata [41], 
	\kme_cceip1_ob_out_post.tdata [40], 
	\kme_cceip1_ob_out_post.tdata [39], 
	\kme_cceip1_ob_out_post.tdata [38], 
	\kme_cceip1_ob_out_post.tdata [37], 
	\kme_cceip1_ob_out_post.tdata [36], 
	\kme_cceip1_ob_out_post.tdata [35], 
	\kme_cceip1_ob_out_post.tdata [34], 
	\kme_cceip1_ob_out_post.tdata [33], 
	\kme_cceip1_ob_out_post.tdata [32], 
	\kme_cceip1_ob_out_post.tdata [31], 
	\kme_cceip1_ob_out_post.tdata [30], 
	\kme_cceip1_ob_out_post.tdata [29], 
	\kme_cceip1_ob_out_post.tdata [28], 
	\kme_cceip1_ob_out_post.tdata [27], 
	\kme_cceip1_ob_out_post.tdata [26], 
	\kme_cceip1_ob_out_post.tdata [25], 
	\kme_cceip1_ob_out_post.tdata [24], 
	\kme_cceip1_ob_out_post.tdata [23], 
	\kme_cceip1_ob_out_post.tdata [22], 
	\kme_cceip1_ob_out_post.tdata [21], 
	\kme_cceip1_ob_out_post.tdata [20], 
	\kme_cceip1_ob_out_post.tdata [19], 
	\kme_cceip1_ob_out_post.tdata [18], 
	\kme_cceip1_ob_out_post.tdata [17], 
	\kme_cceip1_ob_out_post.tdata [16], 
	\kme_cceip1_ob_out_post.tdata [15], 
	\kme_cceip1_ob_out_post.tdata [14], 
	\kme_cceip1_ob_out_post.tdata [13], 
	\kme_cceip1_ob_out_post.tdata [12], 
	\kme_cceip1_ob_out_post.tdata [11], 
	\kme_cceip1_ob_out_post.tdata [10], 
	\kme_cceip1_ob_out_post.tdata [9], \kme_cceip1_ob_out_post.tdata [8], 
	\kme_cceip1_ob_out_post.tdata [7], \kme_cceip1_ob_out_post.tdata [6], 
	\kme_cceip1_ob_out_post.tdata [5], \kme_cceip1_ob_out_post.tdata [4], 
	\kme_cceip1_ob_out_post.tdata [3], \kme_cceip1_ob_out_post.tdata [2], 
	\kme_cceip1_ob_out_post.tdata [1], \kme_cceip1_ob_out_post.tdata [0]} ), 
	.kme_cceip2_ob_out_post( {\kme_cceip2_ob_out_post.tvalid , 
	\kme_cceip2_ob_out_post.tlast , \kme_cceip2_ob_out_post.tid [0], 
	\kme_cceip2_ob_out_post.tstrb [7], \kme_cceip2_ob_out_post.tstrb [6], 
	\kme_cceip2_ob_out_post.tstrb [5], \kme_cceip2_ob_out_post.tstrb [4], 
	\kme_cceip2_ob_out_post.tstrb [3], \kme_cceip2_ob_out_post.tstrb [2], 
	\kme_cceip2_ob_out_post.tstrb [1], \kme_cceip2_ob_out_post.tstrb [0], 
	\kme_cceip2_ob_out_post.tuser [7], \kme_cceip2_ob_out_post.tuser [6], 
	\kme_cceip2_ob_out_post.tuser [5], \kme_cceip2_ob_out_post.tuser [4], 
	\kme_cceip2_ob_out_post.tuser [3], \kme_cceip2_ob_out_post.tuser [2], 
	\kme_cceip2_ob_out_post.tuser [1], \kme_cceip2_ob_out_post.tuser [0], 
	\kme_cceip2_ob_out_post.tdata [63], 
	\kme_cceip2_ob_out_post.tdata [62], 
	\kme_cceip2_ob_out_post.tdata [61], 
	\kme_cceip2_ob_out_post.tdata [60], 
	\kme_cceip2_ob_out_post.tdata [59], 
	\kme_cceip2_ob_out_post.tdata [58], 
	\kme_cceip2_ob_out_post.tdata [57], 
	\kme_cceip2_ob_out_post.tdata [56], 
	\kme_cceip2_ob_out_post.tdata [55], 
	\kme_cceip2_ob_out_post.tdata [54], 
	\kme_cceip2_ob_out_post.tdata [53], 
	\kme_cceip2_ob_out_post.tdata [52], 
	\kme_cceip2_ob_out_post.tdata [51], 
	\kme_cceip2_ob_out_post.tdata [50], 
	\kme_cceip2_ob_out_post.tdata [49], 
	\kme_cceip2_ob_out_post.tdata [48], 
	\kme_cceip2_ob_out_post.tdata [47], 
	\kme_cceip2_ob_out_post.tdata [46], 
	\kme_cceip2_ob_out_post.tdata [45], 
	\kme_cceip2_ob_out_post.tdata [44], 
	\kme_cceip2_ob_out_post.tdata [43], 
	\kme_cceip2_ob_out_post.tdata [42], 
	\kme_cceip2_ob_out_post.tdata [41], 
	\kme_cceip2_ob_out_post.tdata [40], 
	\kme_cceip2_ob_out_post.tdata [39], 
	\kme_cceip2_ob_out_post.tdata [38], 
	\kme_cceip2_ob_out_post.tdata [37], 
	\kme_cceip2_ob_out_post.tdata [36], 
	\kme_cceip2_ob_out_post.tdata [35], 
	\kme_cceip2_ob_out_post.tdata [34], 
	\kme_cceip2_ob_out_post.tdata [33], 
	\kme_cceip2_ob_out_post.tdata [32], 
	\kme_cceip2_ob_out_post.tdata [31], 
	\kme_cceip2_ob_out_post.tdata [30], 
	\kme_cceip2_ob_out_post.tdata [29], 
	\kme_cceip2_ob_out_post.tdata [28], 
	\kme_cceip2_ob_out_post.tdata [27], 
	\kme_cceip2_ob_out_post.tdata [26], 
	\kme_cceip2_ob_out_post.tdata [25], 
	\kme_cceip2_ob_out_post.tdata [24], 
	\kme_cceip2_ob_out_post.tdata [23], 
	\kme_cceip2_ob_out_post.tdata [22], 
	\kme_cceip2_ob_out_post.tdata [21], 
	\kme_cceip2_ob_out_post.tdata [20], 
	\kme_cceip2_ob_out_post.tdata [19], 
	\kme_cceip2_ob_out_post.tdata [18], 
	\kme_cceip2_ob_out_post.tdata [17], 
	\kme_cceip2_ob_out_post.tdata [16], 
	\kme_cceip2_ob_out_post.tdata [15], 
	\kme_cceip2_ob_out_post.tdata [14], 
	\kme_cceip2_ob_out_post.tdata [13], 
	\kme_cceip2_ob_out_post.tdata [12], 
	\kme_cceip2_ob_out_post.tdata [11], 
	\kme_cceip2_ob_out_post.tdata [10], 
	\kme_cceip2_ob_out_post.tdata [9], \kme_cceip2_ob_out_post.tdata [8], 
	\kme_cceip2_ob_out_post.tdata [7], \kme_cceip2_ob_out_post.tdata [6], 
	\kme_cceip2_ob_out_post.tdata [5], \kme_cceip2_ob_out_post.tdata [4], 
	\kme_cceip2_ob_out_post.tdata [3], \kme_cceip2_ob_out_post.tdata [2], 
	\kme_cceip2_ob_out_post.tdata [1], \kme_cceip2_ob_out_post.tdata [0]} ), 
	.kme_cceip3_ob_out_post( {\kme_cceip3_ob_out_post.tvalid , 
	\kme_cceip3_ob_out_post.tlast , \kme_cceip3_ob_out_post.tid [0], 
	\kme_cceip3_ob_out_post.tstrb [7], \kme_cceip3_ob_out_post.tstrb [6], 
	\kme_cceip3_ob_out_post.tstrb [5], \kme_cceip3_ob_out_post.tstrb [4], 
	\kme_cceip3_ob_out_post.tstrb [3], \kme_cceip3_ob_out_post.tstrb [2], 
	\kme_cceip3_ob_out_post.tstrb [1], \kme_cceip3_ob_out_post.tstrb [0], 
	\kme_cceip3_ob_out_post.tuser [7], \kme_cceip3_ob_out_post.tuser [6], 
	\kme_cceip3_ob_out_post.tuser [5], \kme_cceip3_ob_out_post.tuser [4], 
	\kme_cceip3_ob_out_post.tuser [3], \kme_cceip3_ob_out_post.tuser [2], 
	\kme_cceip3_ob_out_post.tuser [1], \kme_cceip3_ob_out_post.tuser [0], 
	\kme_cceip3_ob_out_post.tdata [63], 
	\kme_cceip3_ob_out_post.tdata [62], 
	\kme_cceip3_ob_out_post.tdata [61], 
	\kme_cceip3_ob_out_post.tdata [60], 
	\kme_cceip3_ob_out_post.tdata [59], 
	\kme_cceip3_ob_out_post.tdata [58], 
	\kme_cceip3_ob_out_post.tdata [57], 
	\kme_cceip3_ob_out_post.tdata [56], 
	\kme_cceip3_ob_out_post.tdata [55], 
	\kme_cceip3_ob_out_post.tdata [54], 
	\kme_cceip3_ob_out_post.tdata [53], 
	\kme_cceip3_ob_out_post.tdata [52], 
	\kme_cceip3_ob_out_post.tdata [51], 
	\kme_cceip3_ob_out_post.tdata [50], 
	\kme_cceip3_ob_out_post.tdata [49], 
	\kme_cceip3_ob_out_post.tdata [48], 
	\kme_cceip3_ob_out_post.tdata [47], 
	\kme_cceip3_ob_out_post.tdata [46], 
	\kme_cceip3_ob_out_post.tdata [45], 
	\kme_cceip3_ob_out_post.tdata [44], 
	\kme_cceip3_ob_out_post.tdata [43], 
	\kme_cceip3_ob_out_post.tdata [42], 
	\kme_cceip3_ob_out_post.tdata [41], 
	\kme_cceip3_ob_out_post.tdata [40], 
	\kme_cceip3_ob_out_post.tdata [39], 
	\kme_cceip3_ob_out_post.tdata [38], 
	\kme_cceip3_ob_out_post.tdata [37], 
	\kme_cceip3_ob_out_post.tdata [36], 
	\kme_cceip3_ob_out_post.tdata [35], 
	\kme_cceip3_ob_out_post.tdata [34], 
	\kme_cceip3_ob_out_post.tdata [33], 
	\kme_cceip3_ob_out_post.tdata [32], 
	\kme_cceip3_ob_out_post.tdata [31], 
	\kme_cceip3_ob_out_post.tdata [30], 
	\kme_cceip3_ob_out_post.tdata [29], 
	\kme_cceip3_ob_out_post.tdata [28], 
	\kme_cceip3_ob_out_post.tdata [27], 
	\kme_cceip3_ob_out_post.tdata [26], 
	\kme_cceip3_ob_out_post.tdata [25], 
	\kme_cceip3_ob_out_post.tdata [24], 
	\kme_cceip3_ob_out_post.tdata [23], 
	\kme_cceip3_ob_out_post.tdata [22], 
	\kme_cceip3_ob_out_post.tdata [21], 
	\kme_cceip3_ob_out_post.tdata [20], 
	\kme_cceip3_ob_out_post.tdata [19], 
	\kme_cceip3_ob_out_post.tdata [18], 
	\kme_cceip3_ob_out_post.tdata [17], 
	\kme_cceip3_ob_out_post.tdata [16], 
	\kme_cceip3_ob_out_post.tdata [15], 
	\kme_cceip3_ob_out_post.tdata [14], 
	\kme_cceip3_ob_out_post.tdata [13], 
	\kme_cceip3_ob_out_post.tdata [12], 
	\kme_cceip3_ob_out_post.tdata [11], 
	\kme_cceip3_ob_out_post.tdata [10], 
	\kme_cceip3_ob_out_post.tdata [9], \kme_cceip3_ob_out_post.tdata [8], 
	\kme_cceip3_ob_out_post.tdata [7], \kme_cceip3_ob_out_post.tdata [6], 
	\kme_cceip3_ob_out_post.tdata [5], \kme_cceip3_ob_out_post.tdata [4], 
	\kme_cceip3_ob_out_post.tdata [3], \kme_cceip3_ob_out_post.tdata [2], 
	\kme_cceip3_ob_out_post.tdata [1], \kme_cceip3_ob_out_post.tdata [0]} ), 
	.kme_cddip0_ob_out_post( {\kme_cddip0_ob_out_post.tvalid , 
	\kme_cddip0_ob_out_post.tlast , \kme_cddip0_ob_out_post.tid [0], 
	\kme_cddip0_ob_out_post.tstrb [7], \kme_cddip0_ob_out_post.tstrb [6], 
	\kme_cddip0_ob_out_post.tstrb [5], \kme_cddip0_ob_out_post.tstrb [4], 
	\kme_cddip0_ob_out_post.tstrb [3], \kme_cddip0_ob_out_post.tstrb [2], 
	\kme_cddip0_ob_out_post.tstrb [1], \kme_cddip0_ob_out_post.tstrb [0], 
	\kme_cddip0_ob_out_post.tuser [7], \kme_cddip0_ob_out_post.tuser [6], 
	\kme_cddip0_ob_out_post.tuser [5], \kme_cddip0_ob_out_post.tuser [4], 
	\kme_cddip0_ob_out_post.tuser [3], \kme_cddip0_ob_out_post.tuser [2], 
	\kme_cddip0_ob_out_post.tuser [1], \kme_cddip0_ob_out_post.tuser [0], 
	\kme_cddip0_ob_out_post.tdata [63], 
	\kme_cddip0_ob_out_post.tdata [62], 
	\kme_cddip0_ob_out_post.tdata [61], 
	\kme_cddip0_ob_out_post.tdata [60], 
	\kme_cddip0_ob_out_post.tdata [59], 
	\kme_cddip0_ob_out_post.tdata [58], 
	\kme_cddip0_ob_out_post.tdata [57], 
	\kme_cddip0_ob_out_post.tdata [56], 
	\kme_cddip0_ob_out_post.tdata [55], 
	\kme_cddip0_ob_out_post.tdata [54], 
	\kme_cddip0_ob_out_post.tdata [53], 
	\kme_cddip0_ob_out_post.tdata [52], 
	\kme_cddip0_ob_out_post.tdata [51], 
	\kme_cddip0_ob_out_post.tdata [50], 
	\kme_cddip0_ob_out_post.tdata [49], 
	\kme_cddip0_ob_out_post.tdata [48], 
	\kme_cddip0_ob_out_post.tdata [47], 
	\kme_cddip0_ob_out_post.tdata [46], 
	\kme_cddip0_ob_out_post.tdata [45], 
	\kme_cddip0_ob_out_post.tdata [44], 
	\kme_cddip0_ob_out_post.tdata [43], 
	\kme_cddip0_ob_out_post.tdata [42], 
	\kme_cddip0_ob_out_post.tdata [41], 
	\kme_cddip0_ob_out_post.tdata [40], 
	\kme_cddip0_ob_out_post.tdata [39], 
	\kme_cddip0_ob_out_post.tdata [38], 
	\kme_cddip0_ob_out_post.tdata [37], 
	\kme_cddip0_ob_out_post.tdata [36], 
	\kme_cddip0_ob_out_post.tdata [35], 
	\kme_cddip0_ob_out_post.tdata [34], 
	\kme_cddip0_ob_out_post.tdata [33], 
	\kme_cddip0_ob_out_post.tdata [32], 
	\kme_cddip0_ob_out_post.tdata [31], 
	\kme_cddip0_ob_out_post.tdata [30], 
	\kme_cddip0_ob_out_post.tdata [29], 
	\kme_cddip0_ob_out_post.tdata [28], 
	\kme_cddip0_ob_out_post.tdata [27], 
	\kme_cddip0_ob_out_post.tdata [26], 
	\kme_cddip0_ob_out_post.tdata [25], 
	\kme_cddip0_ob_out_post.tdata [24], 
	\kme_cddip0_ob_out_post.tdata [23], 
	\kme_cddip0_ob_out_post.tdata [22], 
	\kme_cddip0_ob_out_post.tdata [21], 
	\kme_cddip0_ob_out_post.tdata [20], 
	\kme_cddip0_ob_out_post.tdata [19], 
	\kme_cddip0_ob_out_post.tdata [18], 
	\kme_cddip0_ob_out_post.tdata [17], 
	\kme_cddip0_ob_out_post.tdata [16], 
	\kme_cddip0_ob_out_post.tdata [15], 
	\kme_cddip0_ob_out_post.tdata [14], 
	\kme_cddip0_ob_out_post.tdata [13], 
	\kme_cddip0_ob_out_post.tdata [12], 
	\kme_cddip0_ob_out_post.tdata [11], 
	\kme_cddip0_ob_out_post.tdata [10], 
	\kme_cddip0_ob_out_post.tdata [9], \kme_cddip0_ob_out_post.tdata [8], 
	\kme_cddip0_ob_out_post.tdata [7], \kme_cddip0_ob_out_post.tdata [6], 
	\kme_cddip0_ob_out_post.tdata [5], \kme_cddip0_ob_out_post.tdata [4], 
	\kme_cddip0_ob_out_post.tdata [3], \kme_cddip0_ob_out_post.tdata [2], 
	\kme_cddip0_ob_out_post.tdata [1], \kme_cddip0_ob_out_post.tdata [0]} ), 
	.kme_cddip1_ob_out_post( {\kme_cddip1_ob_out_post.tvalid , 
	\kme_cddip1_ob_out_post.tlast , \kme_cddip1_ob_out_post.tid [0], 
	\kme_cddip1_ob_out_post.tstrb [7], \kme_cddip1_ob_out_post.tstrb [6], 
	\kme_cddip1_ob_out_post.tstrb [5], \kme_cddip1_ob_out_post.tstrb [4], 
	\kme_cddip1_ob_out_post.tstrb [3], \kme_cddip1_ob_out_post.tstrb [2], 
	\kme_cddip1_ob_out_post.tstrb [1], \kme_cddip1_ob_out_post.tstrb [0], 
	\kme_cddip1_ob_out_post.tuser [7], \kme_cddip1_ob_out_post.tuser [6], 
	\kme_cddip1_ob_out_post.tuser [5], \kme_cddip1_ob_out_post.tuser [4], 
	\kme_cddip1_ob_out_post.tuser [3], \kme_cddip1_ob_out_post.tuser [2], 
	\kme_cddip1_ob_out_post.tuser [1], \kme_cddip1_ob_out_post.tuser [0], 
	\kme_cddip1_ob_out_post.tdata [63], 
	\kme_cddip1_ob_out_post.tdata [62], 
	\kme_cddip1_ob_out_post.tdata [61], 
	\kme_cddip1_ob_out_post.tdata [60], 
	\kme_cddip1_ob_out_post.tdata [59], 
	\kme_cddip1_ob_out_post.tdata [58], 
	\kme_cddip1_ob_out_post.tdata [57], 
	\kme_cddip1_ob_out_post.tdata [56], 
	\kme_cddip1_ob_out_post.tdata [55], 
	\kme_cddip1_ob_out_post.tdata [54], 
	\kme_cddip1_ob_out_post.tdata [53], 
	\kme_cddip1_ob_out_post.tdata [52], 
	\kme_cddip1_ob_out_post.tdata [51], 
	\kme_cddip1_ob_out_post.tdata [50], 
	\kme_cddip1_ob_out_post.tdata [49], 
	\kme_cddip1_ob_out_post.tdata [48], 
	\kme_cddip1_ob_out_post.tdata [47], 
	\kme_cddip1_ob_out_post.tdata [46], 
	\kme_cddip1_ob_out_post.tdata [45], 
	\kme_cddip1_ob_out_post.tdata [44], 
	\kme_cddip1_ob_out_post.tdata [43], 
	\kme_cddip1_ob_out_post.tdata [42], 
	\kme_cddip1_ob_out_post.tdata [41], 
	\kme_cddip1_ob_out_post.tdata [40], 
	\kme_cddip1_ob_out_post.tdata [39], 
	\kme_cddip1_ob_out_post.tdata [38], 
	\kme_cddip1_ob_out_post.tdata [37], 
	\kme_cddip1_ob_out_post.tdata [36], 
	\kme_cddip1_ob_out_post.tdata [35], 
	\kme_cddip1_ob_out_post.tdata [34], 
	\kme_cddip1_ob_out_post.tdata [33], 
	\kme_cddip1_ob_out_post.tdata [32], 
	\kme_cddip1_ob_out_post.tdata [31], 
	\kme_cddip1_ob_out_post.tdata [30], 
	\kme_cddip1_ob_out_post.tdata [29], 
	\kme_cddip1_ob_out_post.tdata [28], 
	\kme_cddip1_ob_out_post.tdata [27], 
	\kme_cddip1_ob_out_post.tdata [26], 
	\kme_cddip1_ob_out_post.tdata [25], 
	\kme_cddip1_ob_out_post.tdata [24], 
	\kme_cddip1_ob_out_post.tdata [23], 
	\kme_cddip1_ob_out_post.tdata [22], 
	\kme_cddip1_ob_out_post.tdata [21], 
	\kme_cddip1_ob_out_post.tdata [20], 
	\kme_cddip1_ob_out_post.tdata [19], 
	\kme_cddip1_ob_out_post.tdata [18], 
	\kme_cddip1_ob_out_post.tdata [17], 
	\kme_cddip1_ob_out_post.tdata [16], 
	\kme_cddip1_ob_out_post.tdata [15], 
	\kme_cddip1_ob_out_post.tdata [14], 
	\kme_cddip1_ob_out_post.tdata [13], 
	\kme_cddip1_ob_out_post.tdata [12], 
	\kme_cddip1_ob_out_post.tdata [11], 
	\kme_cddip1_ob_out_post.tdata [10], 
	\kme_cddip1_ob_out_post.tdata [9], \kme_cddip1_ob_out_post.tdata [8], 
	\kme_cddip1_ob_out_post.tdata [7], \kme_cddip1_ob_out_post.tdata [6], 
	\kme_cddip1_ob_out_post.tdata [5], \kme_cddip1_ob_out_post.tdata [4], 
	\kme_cddip1_ob_out_post.tdata [3], \kme_cddip1_ob_out_post.tdata [2], 
	\kme_cddip1_ob_out_post.tdata [1], \kme_cddip1_ob_out_post.tdata [0]} ), 
	.kme_cddip2_ob_out_post( {\kme_cddip2_ob_out_post.tvalid , 
	\kme_cddip2_ob_out_post.tlast , \kme_cddip2_ob_out_post.tid [0], 
	\kme_cddip2_ob_out_post.tstrb [7], \kme_cddip2_ob_out_post.tstrb [6], 
	\kme_cddip2_ob_out_post.tstrb [5], \kme_cddip2_ob_out_post.tstrb [4], 
	\kme_cddip2_ob_out_post.tstrb [3], \kme_cddip2_ob_out_post.tstrb [2], 
	\kme_cddip2_ob_out_post.tstrb [1], \kme_cddip2_ob_out_post.tstrb [0], 
	\kme_cddip2_ob_out_post.tuser [7], \kme_cddip2_ob_out_post.tuser [6], 
	\kme_cddip2_ob_out_post.tuser [5], \kme_cddip2_ob_out_post.tuser [4], 
	\kme_cddip2_ob_out_post.tuser [3], \kme_cddip2_ob_out_post.tuser [2], 
	\kme_cddip2_ob_out_post.tuser [1], \kme_cddip2_ob_out_post.tuser [0], 
	\kme_cddip2_ob_out_post.tdata [63], 
	\kme_cddip2_ob_out_post.tdata [62], 
	\kme_cddip2_ob_out_post.tdata [61], 
	\kme_cddip2_ob_out_post.tdata [60], 
	\kme_cddip2_ob_out_post.tdata [59], 
	\kme_cddip2_ob_out_post.tdata [58], 
	\kme_cddip2_ob_out_post.tdata [57], 
	\kme_cddip2_ob_out_post.tdata [56], 
	\kme_cddip2_ob_out_post.tdata [55], 
	\kme_cddip2_ob_out_post.tdata [54], 
	\kme_cddip2_ob_out_post.tdata [53], 
	\kme_cddip2_ob_out_post.tdata [52], 
	\kme_cddip2_ob_out_post.tdata [51], 
	\kme_cddip2_ob_out_post.tdata [50], 
	\kme_cddip2_ob_out_post.tdata [49], 
	\kme_cddip2_ob_out_post.tdata [48], 
	\kme_cddip2_ob_out_post.tdata [47], 
	\kme_cddip2_ob_out_post.tdata [46], 
	\kme_cddip2_ob_out_post.tdata [45], 
	\kme_cddip2_ob_out_post.tdata [44], 
	\kme_cddip2_ob_out_post.tdata [43], 
	\kme_cddip2_ob_out_post.tdata [42], 
	\kme_cddip2_ob_out_post.tdata [41], 
	\kme_cddip2_ob_out_post.tdata [40], 
	\kme_cddip2_ob_out_post.tdata [39], 
	\kme_cddip2_ob_out_post.tdata [38], 
	\kme_cddip2_ob_out_post.tdata [37], 
	\kme_cddip2_ob_out_post.tdata [36], 
	\kme_cddip2_ob_out_post.tdata [35], 
	\kme_cddip2_ob_out_post.tdata [34], 
	\kme_cddip2_ob_out_post.tdata [33], 
	\kme_cddip2_ob_out_post.tdata [32], 
	\kme_cddip2_ob_out_post.tdata [31], 
	\kme_cddip2_ob_out_post.tdata [30], 
	\kme_cddip2_ob_out_post.tdata [29], 
	\kme_cddip2_ob_out_post.tdata [28], 
	\kme_cddip2_ob_out_post.tdata [27], 
	\kme_cddip2_ob_out_post.tdata [26], 
	\kme_cddip2_ob_out_post.tdata [25], 
	\kme_cddip2_ob_out_post.tdata [24], 
	\kme_cddip2_ob_out_post.tdata [23], 
	\kme_cddip2_ob_out_post.tdata [22], 
	\kme_cddip2_ob_out_post.tdata [21], 
	\kme_cddip2_ob_out_post.tdata [20], 
	\kme_cddip2_ob_out_post.tdata [19], 
	\kme_cddip2_ob_out_post.tdata [18], 
	\kme_cddip2_ob_out_post.tdata [17], 
	\kme_cddip2_ob_out_post.tdata [16], 
	\kme_cddip2_ob_out_post.tdata [15], 
	\kme_cddip2_ob_out_post.tdata [14], 
	\kme_cddip2_ob_out_post.tdata [13], 
	\kme_cddip2_ob_out_post.tdata [12], 
	\kme_cddip2_ob_out_post.tdata [11], 
	\kme_cddip2_ob_out_post.tdata [10], 
	\kme_cddip2_ob_out_post.tdata [9], \kme_cddip2_ob_out_post.tdata [8], 
	\kme_cddip2_ob_out_post.tdata [7], \kme_cddip2_ob_out_post.tdata [6], 
	\kme_cddip2_ob_out_post.tdata [5], \kme_cddip2_ob_out_post.tdata [4], 
	\kme_cddip2_ob_out_post.tdata [3], \kme_cddip2_ob_out_post.tdata [2], 
	\kme_cddip2_ob_out_post.tdata [1], \kme_cddip2_ob_out_post.tdata [0]} ), 
	.kme_cddip3_ob_out_post( {\kme_cddip3_ob_out_post.tvalid , 
	\kme_cddip3_ob_out_post.tlast , \kme_cddip3_ob_out_post.tid [0], 
	\kme_cddip3_ob_out_post.tstrb [7], \kme_cddip3_ob_out_post.tstrb [6], 
	\kme_cddip3_ob_out_post.tstrb [5], \kme_cddip3_ob_out_post.tstrb [4], 
	\kme_cddip3_ob_out_post.tstrb [3], \kme_cddip3_ob_out_post.tstrb [2], 
	\kme_cddip3_ob_out_post.tstrb [1], \kme_cddip3_ob_out_post.tstrb [0], 
	\kme_cddip3_ob_out_post.tuser [7], \kme_cddip3_ob_out_post.tuser [6], 
	\kme_cddip3_ob_out_post.tuser [5], \kme_cddip3_ob_out_post.tuser [4], 
	\kme_cddip3_ob_out_post.tuser [3], \kme_cddip3_ob_out_post.tuser [2], 
	\kme_cddip3_ob_out_post.tuser [1], \kme_cddip3_ob_out_post.tuser [0], 
	\kme_cddip3_ob_out_post.tdata [63], 
	\kme_cddip3_ob_out_post.tdata [62], 
	\kme_cddip3_ob_out_post.tdata [61], 
	\kme_cddip3_ob_out_post.tdata [60], 
	\kme_cddip3_ob_out_post.tdata [59], 
	\kme_cddip3_ob_out_post.tdata [58], 
	\kme_cddip3_ob_out_post.tdata [57], 
	\kme_cddip3_ob_out_post.tdata [56], 
	\kme_cddip3_ob_out_post.tdata [55], 
	\kme_cddip3_ob_out_post.tdata [54], 
	\kme_cddip3_ob_out_post.tdata [53], 
	\kme_cddip3_ob_out_post.tdata [52], 
	\kme_cddip3_ob_out_post.tdata [51], 
	\kme_cddip3_ob_out_post.tdata [50], 
	\kme_cddip3_ob_out_post.tdata [49], 
	\kme_cddip3_ob_out_post.tdata [48], 
	\kme_cddip3_ob_out_post.tdata [47], 
	\kme_cddip3_ob_out_post.tdata [46], 
	\kme_cddip3_ob_out_post.tdata [45], 
	\kme_cddip3_ob_out_post.tdata [44], 
	\kme_cddip3_ob_out_post.tdata [43], 
	\kme_cddip3_ob_out_post.tdata [42], 
	\kme_cddip3_ob_out_post.tdata [41], 
	\kme_cddip3_ob_out_post.tdata [40], 
	\kme_cddip3_ob_out_post.tdata [39], 
	\kme_cddip3_ob_out_post.tdata [38], 
	\kme_cddip3_ob_out_post.tdata [37], 
	\kme_cddip3_ob_out_post.tdata [36], 
	\kme_cddip3_ob_out_post.tdata [35], 
	\kme_cddip3_ob_out_post.tdata [34], 
	\kme_cddip3_ob_out_post.tdata [33], 
	\kme_cddip3_ob_out_post.tdata [32], 
	\kme_cddip3_ob_out_post.tdata [31], 
	\kme_cddip3_ob_out_post.tdata [30], 
	\kme_cddip3_ob_out_post.tdata [29], 
	\kme_cddip3_ob_out_post.tdata [28], 
	\kme_cddip3_ob_out_post.tdata [27], 
	\kme_cddip3_ob_out_post.tdata [26], 
	\kme_cddip3_ob_out_post.tdata [25], 
	\kme_cddip3_ob_out_post.tdata [24], 
	\kme_cddip3_ob_out_post.tdata [23], 
	\kme_cddip3_ob_out_post.tdata [22], 
	\kme_cddip3_ob_out_post.tdata [21], 
	\kme_cddip3_ob_out_post.tdata [20], 
	\kme_cddip3_ob_out_post.tdata [19], 
	\kme_cddip3_ob_out_post.tdata [18], 
	\kme_cddip3_ob_out_post.tdata [17], 
	\kme_cddip3_ob_out_post.tdata [16], 
	\kme_cddip3_ob_out_post.tdata [15], 
	\kme_cddip3_ob_out_post.tdata [14], 
	\kme_cddip3_ob_out_post.tdata [13], 
	\kme_cddip3_ob_out_post.tdata [12], 
	\kme_cddip3_ob_out_post.tdata [11], 
	\kme_cddip3_ob_out_post.tdata [10], 
	\kme_cddip3_ob_out_post.tdata [9], \kme_cddip3_ob_out_post.tdata [8], 
	\kme_cddip3_ob_out_post.tdata [7], \kme_cddip3_ob_out_post.tdata [6], 
	\kme_cddip3_ob_out_post.tdata [5], \kme_cddip3_ob_out_post.tdata [4], 
	\kme_cddip3_ob_out_post.tdata [3], \kme_cddip3_ob_out_post.tdata [2], 
	\kme_cddip3_ob_out_post.tdata [1], \kme_cddip3_ob_out_post.tdata [0]} ), 
	cddip3_ism_osync, cddip3_ism_odat, cceip_encrypt_bimc_osync, 
	cceip_encrypt_bimc_odat, cceip_validate_bimc_osync, 
	cceip_validate_bimc_odat, cddip_decrypt_bimc_osync, 
	cddip_decrypt_bimc_odat, axi_bimc_osync, axi_bimc_odat);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [3:0] ckv_cmnd_op;
output [14:0] ckv_cmnd_addr;
output [63:0] ckv_wr_dat;
output [19:0] \ckv_ia_capability.r.part0 ;
wire [3:0] \ckv_ia_capability.f.mem_type ;
wire \ckv_ia_capability.f.ack_error ;
wire \ckv_ia_capability.f.sim_tmo ;
wire [3:0] \ckv_ia_capability.f.reserved_op ;
wire \ckv_ia_capability.f.compare ;
wire \ckv_ia_capability.f.set_init_start ;
wire \ckv_ia_capability.f.initialize_inc ;
wire \ckv_ia_capability.f.initialize ;
wire \ckv_ia_capability.f.reset ;
wire \ckv_ia_capability.f.disabled ;
wire \ckv_ia_capability.f.enable ;
wire \ckv_ia_capability.f.write ;
wire \ckv_ia_capability.f.read ;
wire \ckv_ia_capability.f.nop ;
wire [19:0] ckv_ia_capability;
output [31:0] ckv_ia_rdata_part0;
output [31:0] ckv_ia_rdata_part1;
output [22:0] \ckv_ia_status.r.part0 ;
wire [2:0] \ckv_ia_status.f.code ;
wire [4:0] \ckv_ia_status.f.datawords ;
wire [14:0] \ckv_ia_status.f.addr ;
wire [22:0] ckv_ia_status;
output [3:0] kim_cmnd_op;
output [13:0] kim_cmnd_addr;
output [37:0] kim_wr_dat;
output [19:0] \kim_ia_capability.r.part0 ;
wire [3:0] \kim_ia_capability.f.mem_type ;
wire \kim_ia_capability.f.ack_error ;
wire \kim_ia_capability.f.sim_tmo ;
wire [3:0] \kim_ia_capability.f.reserved_op ;
wire \kim_ia_capability.f.compare ;
wire \kim_ia_capability.f.set_init_start ;
wire \kim_ia_capability.f.initialize_inc ;
wire \kim_ia_capability.f.initialize ;
wire \kim_ia_capability.f.reset ;
wire \kim_ia_capability.f.disabled ;
wire \kim_ia_capability.f.enable ;
wire \kim_ia_capability.f.write ;
wire \kim_ia_capability.f.read ;
wire \kim_ia_capability.f.nop ;
wire [19:0] kim_ia_capability;
output [20:0] kim_ia_rdata_part0;
output [16:0] kim_ia_rdata_part1;
output [21:0] \kim_ia_status.r.part0 ;
wire [2:0] \kim_ia_status.f.code ;
wire [4:0] \kim_ia_status.f.datawords ;
wire [13:0] \kim_ia_status.f.addr ;
wire [21:0] kim_ia_status;
output [7:0] engine_sticky_status;
output disable_ckv_kim_ism_reads;
output send_kme_ib_beat;
output debug_kme_ib_tvalid;
output debug_kme_ib_tlast;
output [0:0] debug_kme_ib_tid;
output [7:0] debug_kme_ib_tstrb;
output [7:0] debug_kme_ib_tuser;
output [63:0] debug_kme_ib_tdata;
output \kme_cceip0_ob_out.tvalid ;
output \kme_cceip0_ob_out.tlast ;
output [0:0] \kme_cceip0_ob_out.tid ;
output [7:0] \kme_cceip0_ob_out.tstrb ;
output [7:0] \kme_cceip0_ob_out.tuser ;
output [63:0] \kme_cceip0_ob_out.tdata ;
wire [82:0] kme_cceip0_ob_out;
output \kme_cceip1_ob_out.tvalid ;
output \kme_cceip1_ob_out.tlast ;
output [0:0] \kme_cceip1_ob_out.tid ;
output [7:0] \kme_cceip1_ob_out.tstrb ;
output [7:0] \kme_cceip1_ob_out.tuser ;
output [63:0] \kme_cceip1_ob_out.tdata ;
wire [82:0] kme_cceip1_ob_out;
output \kme_cceip2_ob_out.tvalid ;
output \kme_cceip2_ob_out.tlast ;
output [0:0] \kme_cceip2_ob_out.tid ;
output [7:0] \kme_cceip2_ob_out.tstrb ;
output [7:0] \kme_cceip2_ob_out.tuser ;
output [63:0] \kme_cceip2_ob_out.tdata ;
wire [82:0] kme_cceip2_ob_out;
output \kme_cceip3_ob_out.tvalid ;
output \kme_cceip3_ob_out.tlast ;
output [0:0] \kme_cceip3_ob_out.tid ;
output [7:0] \kme_cceip3_ob_out.tstrb ;
output [7:0] \kme_cceip3_ob_out.tuser ;
output [63:0] \kme_cceip3_ob_out.tdata ;
wire [82:0] kme_cceip3_ob_out;
output \kme_cddip0_ob_out.tvalid ;
output \kme_cddip0_ob_out.tlast ;
output [0:0] \kme_cddip0_ob_out.tid ;
output [7:0] \kme_cddip0_ob_out.tstrb ;
output [7:0] \kme_cddip0_ob_out.tuser ;
output [63:0] \kme_cddip0_ob_out.tdata ;
wire [82:0] kme_cddip0_ob_out;
output \kme_cddip1_ob_out.tvalid ;
output \kme_cddip1_ob_out.tlast ;
output [0:0] \kme_cddip1_ob_out.tid ;
output [7:0] \kme_cddip1_ob_out.tstrb ;
output [7:0] \kme_cddip1_ob_out.tuser ;
output [63:0] \kme_cddip1_ob_out.tdata ;
wire [82:0] kme_cddip1_ob_out;
output \kme_cddip2_ob_out.tvalid ;
output \kme_cddip2_ob_out.tlast ;
output [0:0] \kme_cddip2_ob_out.tid ;
output [7:0] \kme_cddip2_ob_out.tstrb ;
output [7:0] \kme_cddip2_ob_out.tuser ;
output [63:0] \kme_cddip2_ob_out.tdata ;
wire [82:0] kme_cddip2_ob_out;
output \kme_cddip3_ob_out.tvalid ;
output \kme_cddip3_ob_out.tlast ;
output [0:0] \kme_cddip3_ob_out.tid ;
output [7:0] \kme_cddip3_ob_out.tstrb ;
output [7:0] \kme_cddip3_ob_out.tuser ;
output [63:0] \kme_cddip3_ob_out.tdata ;
wire [82:0] kme_cddip3_ob_out;
output cceip_encrypt_bimc_isync;
output cceip_encrypt_bimc_idat;
output cceip_validate_bimc_isync;
output cceip_validate_bimc_idat;
output cddip_decrypt_bimc_isync;
output cddip_decrypt_bimc_idat;
output axi_bimc_isync;
output axi_bimc_idat;
output axi_term_bimc_isync;
output axi_term_bimc_idat;
input clk;
input rst_n;
input [2:0] ckv_stat_code;
input [4:0] ckv_stat_datawords;
input [14:0] ckv_stat_addr;
input [3:0] ckv_capability_type;
input [15:0] ckv_capability_lst;
input [63:0] ckv_rd_dat;
input [18:0] \o_ckv_ia_config.r.part0 ;
wire [3:0] \o_ckv_ia_config.f.op ;
wire [14:0] \o_ckv_ia_config.f.addr ;
wire [18:0] o_ckv_ia_config;
input [31:0] o_ckv_ia_wdata_part0;
input [31:0] o_ckv_ia_wdata_part1;
input [2:0] kim_stat_code;
input [4:0] kim_stat_datawords;
input [13:0] kim_stat_addr;
input [3:0] kim_capability_type;
input [15:0] kim_capability_lst;
input [37:0] kim_rd_dat;
input [17:0] \o_kim_ia_config.r.part0 ;
wire [3:0] \o_kim_ia_config.f.op ;
wire [13:0] \o_kim_ia_config.f.addr ;
wire [17:0] o_kim_ia_config;
input [20:0] o_kim_ia_wdata_part0;
input [16:0] o_kim_ia_wdata_part1;
input [7:0] set_rsm_is_backpressuring;
input wr_stb;
input [31:0] wr_data;
input [10:0] reg_addr;
input [7:0] o_engine_sticky_status;
input o_disable_ckv_kim_ism_reads;
input o_send_kme_ib_beat;
input [31:0] \cceip0_out_ia_wdata.r.part2 ;
input [31:0] \cceip0_out_ia_wdata.r.part1 ;
input [31:0] \cceip0_out_ia_wdata.r.part0 ;
wire [31:0] \cceip0_out_ia_wdata.f.tdata_hi ;
wire [31:0] \cceip0_out_ia_wdata.f.tdata_lo ;
wire \cceip0_out_ia_wdata.f.eob ;
wire [7:0] \cceip0_out_ia_wdata.f.bytes_vld ;
wire [7:0] \cceip0_out_ia_wdata.f.unused1 ;
wire \cceip0_out_ia_wdata.f.tid ;
wire [7:0] \cceip0_out_ia_wdata.f.tuser ;
wire [5:0] \cceip0_out_ia_wdata.f.unused0 ;
wire [95:0] cceip0_out_ia_wdata;
input debug_kme_ib_tready;
input [8:0] \tready_override.r.part0 ;
wire \tready_override.f.txc_tready_override ;
wire \tready_override.f.engine_7_tready_override ;
wire \tready_override.f.engine_6_tready_override ;
wire \tready_override.f.engine_5_tready_override ;
wire \tready_override.f.engine_4_tready_override ;
wire \tready_override.f.engine_3_tready_override ;
wire \tready_override.f.engine_2_tready_override ;
wire \tready_override.f.engine_1_tready_override ;
wire \tready_override.f.engine_0_tready_override ;
wire [8:0] tready_override;
input \kme_cceip0_ob_out_post.tvalid ;
input \kme_cceip0_ob_out_post.tlast ;
input [0:0] \kme_cceip0_ob_out_post.tid ;
input [7:0] \kme_cceip0_ob_out_post.tstrb ;
input [7:0] \kme_cceip0_ob_out_post.tuser ;
input [63:0] \kme_cceip0_ob_out_post.tdata ;
wire [82:0] kme_cceip0_ob_out_post;
input \kme_cceip1_ob_out_post.tvalid ;
input \kme_cceip1_ob_out_post.tlast ;
input [0:0] \kme_cceip1_ob_out_post.tid ;
input [7:0] \kme_cceip1_ob_out_post.tstrb ;
input [7:0] \kme_cceip1_ob_out_post.tuser ;
input [63:0] \kme_cceip1_ob_out_post.tdata ;
wire [82:0] kme_cceip1_ob_out_post;
input \kme_cceip2_ob_out_post.tvalid ;
input \kme_cceip2_ob_out_post.tlast ;
input [0:0] \kme_cceip2_ob_out_post.tid ;
input [7:0] \kme_cceip2_ob_out_post.tstrb ;
input [7:0] \kme_cceip2_ob_out_post.tuser ;
input [63:0] \kme_cceip2_ob_out_post.tdata ;
wire [82:0] kme_cceip2_ob_out_post;
input \kme_cceip3_ob_out_post.tvalid ;
input \kme_cceip3_ob_out_post.tlast ;
input [0:0] \kme_cceip3_ob_out_post.tid ;
input [7:0] \kme_cceip3_ob_out_post.tstrb ;
input [7:0] \kme_cceip3_ob_out_post.tuser ;
input [63:0] \kme_cceip3_ob_out_post.tdata ;
wire [82:0] kme_cceip3_ob_out_post;
input \kme_cddip0_ob_out_post.tvalid ;
input \kme_cddip0_ob_out_post.tlast ;
input [0:0] \kme_cddip0_ob_out_post.tid ;
input [7:0] \kme_cddip0_ob_out_post.tstrb ;
input [7:0] \kme_cddip0_ob_out_post.tuser ;
input [63:0] \kme_cddip0_ob_out_post.tdata ;
wire [82:0] kme_cddip0_ob_out_post;
input \kme_cddip1_ob_out_post.tvalid ;
input \kme_cddip1_ob_out_post.tlast ;
input [0:0] \kme_cddip1_ob_out_post.tid ;
input [7:0] \kme_cddip1_ob_out_post.tstrb ;
input [7:0] \kme_cddip1_ob_out_post.tuser ;
input [63:0] \kme_cddip1_ob_out_post.tdata ;
wire [82:0] kme_cddip1_ob_out_post;
input \kme_cddip2_ob_out_post.tvalid ;
input \kme_cddip2_ob_out_post.tlast ;
input [0:0] \kme_cddip2_ob_out_post.tid ;
input [7:0] \kme_cddip2_ob_out_post.tstrb ;
input [7:0] \kme_cddip2_ob_out_post.tuser ;
input [63:0] \kme_cddip2_ob_out_post.tdata ;
wire [82:0] kme_cddip2_ob_out_post;
input \kme_cddip3_ob_out_post.tvalid ;
input \kme_cddip3_ob_out_post.tlast ;
input [0:0] \kme_cddip3_ob_out_post.tid ;
input [7:0] \kme_cddip3_ob_out_post.tstrb ;
input [7:0] \kme_cddip3_ob_out_post.tuser ;
input [63:0] \kme_cddip3_ob_out_post.tdata ;
wire [82:0] kme_cddip3_ob_out_post;
input cddip3_ism_osync;
input cddip3_ism_odat;
input cceip_encrypt_bimc_osync;
input cceip_encrypt_bimc_odat;
input cceip_validate_bimc_osync;
input cceip_validate_bimc_odat;
input cddip_decrypt_bimc_osync;
input cddip_decrypt_bimc_odat;
input axi_bimc_osync;
input axi_bimc_odat;
wire [0:19] _zy_simnet_ckv_ia_capability_0_w$;
wire [0:22] _zy_simnet_ckv_ia_status_1_w$;
wire [0:19] _zy_simnet_kim_ia_capability_2_w$;
wire [0:21] _zy_simnet_kim_ia_status_3_w$;
wire [0:7] _zy_simnet_engine_sticky_status_4_w$;
wire _zy_simnet_disable_ckv_kim_ism_reads_5_w$;
wire _zy_simnet_send_kme_ib_beat_6_w$;
wire _zy_simnet_debug_kme_ib_tvalid_7_w$;
wire _zy_simnet_debug_kme_ib_tlast_8_w$;
wire _zy_simnet_debug_kme_ib_tid_9_w$;
wire [0:7] _zy_simnet_debug_kme_ib_tstrb_10_w$;
wire [0:7] _zy_simnet_debug_kme_ib_tuser_11_w$;
wire [0:63] _zy_simnet_debug_kme_ib_tdata_12_w$;
wire [0:82] _zy_simnet_kme_cceip0_ob_out_13_w$;
wire [0:82] _zy_simnet_kme_cceip1_ob_out_14_w$;
wire [0:82] _zy_simnet_kme_cceip2_ob_out_15_w$;
wire [0:82] _zy_simnet_kme_cceip3_ob_out_16_w$;
wire [0:82] _zy_simnet_kme_cddip0_ob_out_17_w$;
wire [0:82] _zy_simnet_kme_cddip1_ob_out_18_w$;
wire [0:82] _zy_simnet_kme_cddip2_ob_out_19_w$;
wire [0:82] _zy_simnet_kme_cddip3_ob_out_20_w$;
wire [31:0] i;
tran (ckv_ia_capability[19], \ckv_ia_capability.r.part0 [19]);
tran (ckv_ia_capability[19], \ckv_ia_capability.f.mem_type [3]);
tran (ckv_ia_capability[18], \ckv_ia_capability.r.part0 [18]);
tran (ckv_ia_capability[18], \ckv_ia_capability.f.mem_type [2]);
tran (ckv_ia_capability[17], \ckv_ia_capability.r.part0 [17]);
tran (ckv_ia_capability[17], \ckv_ia_capability.f.mem_type [1]);
tran (ckv_ia_capability[16], \ckv_ia_capability.r.part0 [16]);
tran (ckv_ia_capability[16], \ckv_ia_capability.f.mem_type [0]);
tran (ckv_ia_capability[15], \ckv_ia_capability.r.part0 [15]);
tran (ckv_ia_capability[15], \ckv_ia_capability.f.ack_error );
tran (ckv_ia_capability[14], \ckv_ia_capability.r.part0 [14]);
tran (ckv_ia_capability[14], \ckv_ia_capability.f.sim_tmo );
tran (ckv_ia_capability[13], \ckv_ia_capability.r.part0 [13]);
tran (ckv_ia_capability[13], \ckv_ia_capability.f.reserved_op [3]);
tran (ckv_ia_capability[12], \ckv_ia_capability.r.part0 [12]);
tran (ckv_ia_capability[12], \ckv_ia_capability.f.reserved_op [2]);
tran (ckv_ia_capability[11], \ckv_ia_capability.r.part0 [11]);
tran (ckv_ia_capability[11], \ckv_ia_capability.f.reserved_op [1]);
tran (ckv_ia_capability[10], \ckv_ia_capability.r.part0 [10]);
tran (ckv_ia_capability[10], \ckv_ia_capability.f.reserved_op [0]);
tran (ckv_ia_capability[9], \ckv_ia_capability.r.part0 [9]);
tran (ckv_ia_capability[9], \ckv_ia_capability.f.compare );
tran (ckv_ia_capability[8], \ckv_ia_capability.r.part0 [8]);
tran (ckv_ia_capability[8], \ckv_ia_capability.f.set_init_start );
tran (ckv_ia_capability[7], \ckv_ia_capability.r.part0 [7]);
tran (ckv_ia_capability[7], \ckv_ia_capability.f.initialize_inc );
tran (ckv_ia_capability[6], \ckv_ia_capability.r.part0 [6]);
tran (ckv_ia_capability[6], \ckv_ia_capability.f.initialize );
tran (ckv_ia_capability[5], \ckv_ia_capability.r.part0 [5]);
tran (ckv_ia_capability[5], \ckv_ia_capability.f.reset );
tran (ckv_ia_capability[4], \ckv_ia_capability.r.part0 [4]);
tran (ckv_ia_capability[4], \ckv_ia_capability.f.disabled );
tran (ckv_ia_capability[3], \ckv_ia_capability.r.part0 [3]);
tran (ckv_ia_capability[3], \ckv_ia_capability.f.enable );
tran (ckv_ia_capability[2], \ckv_ia_capability.r.part0 [2]);
tran (ckv_ia_capability[2], \ckv_ia_capability.f.write );
tran (ckv_ia_capability[1], \ckv_ia_capability.r.part0 [1]);
tran (ckv_ia_capability[1], \ckv_ia_capability.f.read );
tran (ckv_ia_capability[0], \ckv_ia_capability.r.part0 [0]);
tran (ckv_ia_capability[0], \ckv_ia_capability.f.nop );
tran (ckv_ia_status[22], \ckv_ia_status.r.part0 [22]);
tran (ckv_ia_status[22], \ckv_ia_status.f.code [2]);
tran (ckv_ia_status[21], \ckv_ia_status.r.part0 [21]);
tran (ckv_ia_status[21], \ckv_ia_status.f.code [1]);
tran (ckv_ia_status[20], \ckv_ia_status.r.part0 [20]);
tran (ckv_ia_status[20], \ckv_ia_status.f.code [0]);
tran (ckv_ia_status[19], \ckv_ia_status.r.part0 [19]);
tran (ckv_ia_status[19], \ckv_ia_status.f.datawords [4]);
tran (ckv_ia_status[18], \ckv_ia_status.r.part0 [18]);
tran (ckv_ia_status[18], \ckv_ia_status.f.datawords [3]);
tran (ckv_ia_status[17], \ckv_ia_status.r.part0 [17]);
tran (ckv_ia_status[17], \ckv_ia_status.f.datawords [2]);
tran (ckv_ia_status[16], \ckv_ia_status.r.part0 [16]);
tran (ckv_ia_status[16], \ckv_ia_status.f.datawords [1]);
tran (ckv_ia_status[15], \ckv_ia_status.r.part0 [15]);
tran (ckv_ia_status[15], \ckv_ia_status.f.datawords [0]);
tran (ckv_ia_status[14], \ckv_ia_status.r.part0 [14]);
tran (ckv_ia_status[14], \ckv_ia_status.f.addr [14]);
tran (ckv_ia_status[13], \ckv_ia_status.r.part0 [13]);
tran (ckv_ia_status[13], \ckv_ia_status.f.addr [13]);
tran (ckv_ia_status[12], \ckv_ia_status.r.part0 [12]);
tran (ckv_ia_status[12], \ckv_ia_status.f.addr [12]);
tran (ckv_ia_status[11], \ckv_ia_status.r.part0 [11]);
tran (ckv_ia_status[11], \ckv_ia_status.f.addr [11]);
tran (ckv_ia_status[10], \ckv_ia_status.r.part0 [10]);
tran (ckv_ia_status[10], \ckv_ia_status.f.addr [10]);
tran (ckv_ia_status[9], \ckv_ia_status.r.part0 [9]);
tran (ckv_ia_status[9], \ckv_ia_status.f.addr [9]);
tran (ckv_ia_status[8], \ckv_ia_status.r.part0 [8]);
tran (ckv_ia_status[8], \ckv_ia_status.f.addr [8]);
tran (ckv_ia_status[7], \ckv_ia_status.r.part0 [7]);
tran (ckv_ia_status[7], \ckv_ia_status.f.addr [7]);
tran (ckv_ia_status[6], \ckv_ia_status.r.part0 [6]);
tran (ckv_ia_status[6], \ckv_ia_status.f.addr [6]);
tran (ckv_ia_status[5], \ckv_ia_status.r.part0 [5]);
tran (ckv_ia_status[5], \ckv_ia_status.f.addr [5]);
tran (ckv_ia_status[4], \ckv_ia_status.r.part0 [4]);
tran (ckv_ia_status[4], \ckv_ia_status.f.addr [4]);
tran (ckv_ia_status[3], \ckv_ia_status.r.part0 [3]);
tran (ckv_ia_status[3], \ckv_ia_status.f.addr [3]);
tran (ckv_ia_status[2], \ckv_ia_status.r.part0 [2]);
tran (ckv_ia_status[2], \ckv_ia_status.f.addr [2]);
tran (ckv_ia_status[1], \ckv_ia_status.r.part0 [1]);
tran (ckv_ia_status[1], \ckv_ia_status.f.addr [1]);
tran (ckv_ia_status[0], \ckv_ia_status.r.part0 [0]);
tran (ckv_ia_status[0], \ckv_ia_status.f.addr [0]);
tran (kim_ia_capability[19], \kim_ia_capability.r.part0 [19]);
tran (kim_ia_capability[19], \kim_ia_capability.f.mem_type [3]);
tran (kim_ia_capability[18], \kim_ia_capability.r.part0 [18]);
tran (kim_ia_capability[18], \kim_ia_capability.f.mem_type [2]);
tran (kim_ia_capability[17], \kim_ia_capability.r.part0 [17]);
tran (kim_ia_capability[17], \kim_ia_capability.f.mem_type [1]);
tran (kim_ia_capability[16], \kim_ia_capability.r.part0 [16]);
tran (kim_ia_capability[16], \kim_ia_capability.f.mem_type [0]);
tran (kim_ia_capability[15], \kim_ia_capability.r.part0 [15]);
tran (kim_ia_capability[15], \kim_ia_capability.f.ack_error );
tran (kim_ia_capability[14], \kim_ia_capability.r.part0 [14]);
tran (kim_ia_capability[14], \kim_ia_capability.f.sim_tmo );
tran (kim_ia_capability[13], \kim_ia_capability.r.part0 [13]);
tran (kim_ia_capability[13], \kim_ia_capability.f.reserved_op [3]);
tran (kim_ia_capability[12], \kim_ia_capability.r.part0 [12]);
tran (kim_ia_capability[12], \kim_ia_capability.f.reserved_op [2]);
tran (kim_ia_capability[11], \kim_ia_capability.r.part0 [11]);
tran (kim_ia_capability[11], \kim_ia_capability.f.reserved_op [1]);
tran (kim_ia_capability[10], \kim_ia_capability.r.part0 [10]);
tran (kim_ia_capability[10], \kim_ia_capability.f.reserved_op [0]);
tran (kim_ia_capability[9], \kim_ia_capability.r.part0 [9]);
tran (kim_ia_capability[9], \kim_ia_capability.f.compare );
tran (kim_ia_capability[8], \kim_ia_capability.r.part0 [8]);
tran (kim_ia_capability[8], \kim_ia_capability.f.set_init_start );
tran (kim_ia_capability[7], \kim_ia_capability.r.part0 [7]);
tran (kim_ia_capability[7], \kim_ia_capability.f.initialize_inc );
tran (kim_ia_capability[6], \kim_ia_capability.r.part0 [6]);
tran (kim_ia_capability[6], \kim_ia_capability.f.initialize );
tran (kim_ia_capability[5], \kim_ia_capability.r.part0 [5]);
tran (kim_ia_capability[5], \kim_ia_capability.f.reset );
tran (kim_ia_capability[4], \kim_ia_capability.r.part0 [4]);
tran (kim_ia_capability[4], \kim_ia_capability.f.disabled );
tran (kim_ia_capability[3], \kim_ia_capability.r.part0 [3]);
tran (kim_ia_capability[3], \kim_ia_capability.f.enable );
tran (kim_ia_capability[2], \kim_ia_capability.r.part0 [2]);
tran (kim_ia_capability[2], \kim_ia_capability.f.write );
tran (kim_ia_capability[1], \kim_ia_capability.r.part0 [1]);
tran (kim_ia_capability[1], \kim_ia_capability.f.read );
tran (kim_ia_capability[0], \kim_ia_capability.r.part0 [0]);
tran (kim_ia_capability[0], \kim_ia_capability.f.nop );
tran (kim_ia_status[21], \kim_ia_status.r.part0 [21]);
tran (kim_ia_status[21], \kim_ia_status.f.code [2]);
tran (kim_ia_status[20], \kim_ia_status.r.part0 [20]);
tran (kim_ia_status[20], \kim_ia_status.f.code [1]);
tran (kim_ia_status[19], \kim_ia_status.r.part0 [19]);
tran (kim_ia_status[19], \kim_ia_status.f.code [0]);
tran (kim_ia_status[18], \kim_ia_status.r.part0 [18]);
tran (kim_ia_status[18], \kim_ia_status.f.datawords [4]);
tran (kim_ia_status[17], \kim_ia_status.r.part0 [17]);
tran (kim_ia_status[17], \kim_ia_status.f.datawords [3]);
tran (kim_ia_status[16], \kim_ia_status.r.part0 [16]);
tran (kim_ia_status[16], \kim_ia_status.f.datawords [2]);
tran (kim_ia_status[15], \kim_ia_status.r.part0 [15]);
tran (kim_ia_status[15], \kim_ia_status.f.datawords [1]);
tran (kim_ia_status[14], \kim_ia_status.r.part0 [14]);
tran (kim_ia_status[14], \kim_ia_status.f.datawords [0]);
tran (kim_ia_status[13], \kim_ia_status.r.part0 [13]);
tran (kim_ia_status[13], \kim_ia_status.f.addr [13]);
tran (kim_ia_status[12], \kim_ia_status.r.part0 [12]);
tran (kim_ia_status[12], \kim_ia_status.f.addr [12]);
tran (kim_ia_status[11], \kim_ia_status.r.part0 [11]);
tran (kim_ia_status[11], \kim_ia_status.f.addr [11]);
tran (kim_ia_status[10], \kim_ia_status.r.part0 [10]);
tran (kim_ia_status[10], \kim_ia_status.f.addr [10]);
tran (kim_ia_status[9], \kim_ia_status.r.part0 [9]);
tran (kim_ia_status[9], \kim_ia_status.f.addr [9]);
tran (kim_ia_status[8], \kim_ia_status.r.part0 [8]);
tran (kim_ia_status[8], \kim_ia_status.f.addr [8]);
tran (kim_ia_status[7], \kim_ia_status.r.part0 [7]);
tran (kim_ia_status[7], \kim_ia_status.f.addr [7]);
tran (kim_ia_status[6], \kim_ia_status.r.part0 [6]);
tran (kim_ia_status[6], \kim_ia_status.f.addr [6]);
tran (kim_ia_status[5], \kim_ia_status.r.part0 [5]);
tran (kim_ia_status[5], \kim_ia_status.f.addr [5]);
tran (kim_ia_status[4], \kim_ia_status.r.part0 [4]);
tran (kim_ia_status[4], \kim_ia_status.f.addr [4]);
tran (kim_ia_status[3], \kim_ia_status.r.part0 [3]);
tran (kim_ia_status[3], \kim_ia_status.f.addr [3]);
tran (kim_ia_status[2], \kim_ia_status.r.part0 [2]);
tran (kim_ia_status[2], \kim_ia_status.f.addr [2]);
tran (kim_ia_status[1], \kim_ia_status.r.part0 [1]);
tran (kim_ia_status[1], \kim_ia_status.f.addr [1]);
tran (kim_ia_status[0], \kim_ia_status.r.part0 [0]);
tran (kim_ia_status[0], \kim_ia_status.f.addr [0]);
tran (kme_cceip0_ob_out[82], \kme_cceip0_ob_out.tvalid );
tran (kme_cceip0_ob_out[81], \kme_cceip0_ob_out.tlast );
tran (kme_cceip0_ob_out[80], \kme_cceip0_ob_out.tid [0]);
tran (kme_cceip0_ob_out[79], \kme_cceip0_ob_out.tstrb [7]);
tran (kme_cceip0_ob_out[78], \kme_cceip0_ob_out.tstrb [6]);
tran (kme_cceip0_ob_out[77], \kme_cceip0_ob_out.tstrb [5]);
tran (kme_cceip0_ob_out[76], \kme_cceip0_ob_out.tstrb [4]);
tran (kme_cceip0_ob_out[75], \kme_cceip0_ob_out.tstrb [3]);
tran (kme_cceip0_ob_out[74], \kme_cceip0_ob_out.tstrb [2]);
tran (kme_cceip0_ob_out[73], \kme_cceip0_ob_out.tstrb [1]);
tran (kme_cceip0_ob_out[72], \kme_cceip0_ob_out.tstrb [0]);
tran (kme_cceip0_ob_out[71], \kme_cceip0_ob_out.tuser [7]);
tran (kme_cceip0_ob_out[70], \kme_cceip0_ob_out.tuser [6]);
tran (kme_cceip0_ob_out[69], \kme_cceip0_ob_out.tuser [5]);
tran (kme_cceip0_ob_out[68], \kme_cceip0_ob_out.tuser [4]);
tran (kme_cceip0_ob_out[67], \kme_cceip0_ob_out.tuser [3]);
tran (kme_cceip0_ob_out[66], \kme_cceip0_ob_out.tuser [2]);
tran (kme_cceip0_ob_out[65], \kme_cceip0_ob_out.tuser [1]);
tran (kme_cceip0_ob_out[64], \kme_cceip0_ob_out.tuser [0]);
tran (kme_cceip0_ob_out[63], \kme_cceip0_ob_out.tdata [63]);
tran (kme_cceip0_ob_out[62], \kme_cceip0_ob_out.tdata [62]);
tran (kme_cceip0_ob_out[61], \kme_cceip0_ob_out.tdata [61]);
tran (kme_cceip0_ob_out[60], \kme_cceip0_ob_out.tdata [60]);
tran (kme_cceip0_ob_out[59], \kme_cceip0_ob_out.tdata [59]);
tran (kme_cceip0_ob_out[58], \kme_cceip0_ob_out.tdata [58]);
tran (kme_cceip0_ob_out[57], \kme_cceip0_ob_out.tdata [57]);
tran (kme_cceip0_ob_out[56], \kme_cceip0_ob_out.tdata [56]);
tran (kme_cceip0_ob_out[55], \kme_cceip0_ob_out.tdata [55]);
tran (kme_cceip0_ob_out[54], \kme_cceip0_ob_out.tdata [54]);
tran (kme_cceip0_ob_out[53], \kme_cceip0_ob_out.tdata [53]);
tran (kme_cceip0_ob_out[52], \kme_cceip0_ob_out.tdata [52]);
tran (kme_cceip0_ob_out[51], \kme_cceip0_ob_out.tdata [51]);
tran (kme_cceip0_ob_out[50], \kme_cceip0_ob_out.tdata [50]);
tran (kme_cceip0_ob_out[49], \kme_cceip0_ob_out.tdata [49]);
tran (kme_cceip0_ob_out[48], \kme_cceip0_ob_out.tdata [48]);
tran (kme_cceip0_ob_out[47], \kme_cceip0_ob_out.tdata [47]);
tran (kme_cceip0_ob_out[46], \kme_cceip0_ob_out.tdata [46]);
tran (kme_cceip0_ob_out[45], \kme_cceip0_ob_out.tdata [45]);
tran (kme_cceip0_ob_out[44], \kme_cceip0_ob_out.tdata [44]);
tran (kme_cceip0_ob_out[43], \kme_cceip0_ob_out.tdata [43]);
tran (kme_cceip0_ob_out[42], \kme_cceip0_ob_out.tdata [42]);
tran (kme_cceip0_ob_out[41], \kme_cceip0_ob_out.tdata [41]);
tran (kme_cceip0_ob_out[40], \kme_cceip0_ob_out.tdata [40]);
tran (kme_cceip0_ob_out[39], \kme_cceip0_ob_out.tdata [39]);
tran (kme_cceip0_ob_out[38], \kme_cceip0_ob_out.tdata [38]);
tran (kme_cceip0_ob_out[37], \kme_cceip0_ob_out.tdata [37]);
tran (kme_cceip0_ob_out[36], \kme_cceip0_ob_out.tdata [36]);
tran (kme_cceip0_ob_out[35], \kme_cceip0_ob_out.tdata [35]);
tran (kme_cceip0_ob_out[34], \kme_cceip0_ob_out.tdata [34]);
tran (kme_cceip0_ob_out[33], \kme_cceip0_ob_out.tdata [33]);
tran (kme_cceip0_ob_out[32], \kme_cceip0_ob_out.tdata [32]);
tran (kme_cceip0_ob_out[31], \kme_cceip0_ob_out.tdata [31]);
tran (kme_cceip0_ob_out[30], \kme_cceip0_ob_out.tdata [30]);
tran (kme_cceip0_ob_out[29], \kme_cceip0_ob_out.tdata [29]);
tran (kme_cceip0_ob_out[28], \kme_cceip0_ob_out.tdata [28]);
tran (kme_cceip0_ob_out[27], \kme_cceip0_ob_out.tdata [27]);
tran (kme_cceip0_ob_out[26], \kme_cceip0_ob_out.tdata [26]);
tran (kme_cceip0_ob_out[25], \kme_cceip0_ob_out.tdata [25]);
tran (kme_cceip0_ob_out[24], \kme_cceip0_ob_out.tdata [24]);
tran (kme_cceip0_ob_out[23], \kme_cceip0_ob_out.tdata [23]);
tran (kme_cceip0_ob_out[22], \kme_cceip0_ob_out.tdata [22]);
tran (kme_cceip0_ob_out[21], \kme_cceip0_ob_out.tdata [21]);
tran (kme_cceip0_ob_out[20], \kme_cceip0_ob_out.tdata [20]);
tran (kme_cceip0_ob_out[19], \kme_cceip0_ob_out.tdata [19]);
tran (kme_cceip0_ob_out[18], \kme_cceip0_ob_out.tdata [18]);
tran (kme_cceip0_ob_out[17], \kme_cceip0_ob_out.tdata [17]);
tran (kme_cceip0_ob_out[16], \kme_cceip0_ob_out.tdata [16]);
tran (kme_cceip0_ob_out[15], \kme_cceip0_ob_out.tdata [15]);
tran (kme_cceip0_ob_out[14], \kme_cceip0_ob_out.tdata [14]);
tran (kme_cceip0_ob_out[13], \kme_cceip0_ob_out.tdata [13]);
tran (kme_cceip0_ob_out[12], \kme_cceip0_ob_out.tdata [12]);
tran (kme_cceip0_ob_out[11], \kme_cceip0_ob_out.tdata [11]);
tran (kme_cceip0_ob_out[10], \kme_cceip0_ob_out.tdata [10]);
tran (kme_cceip0_ob_out[9], \kme_cceip0_ob_out.tdata [9]);
tran (kme_cceip0_ob_out[8], \kme_cceip0_ob_out.tdata [8]);
tran (kme_cceip0_ob_out[7], \kme_cceip0_ob_out.tdata [7]);
tran (kme_cceip0_ob_out[6], \kme_cceip0_ob_out.tdata [6]);
tran (kme_cceip0_ob_out[5], \kme_cceip0_ob_out.tdata [5]);
tran (kme_cceip0_ob_out[4], \kme_cceip0_ob_out.tdata [4]);
tran (kme_cceip0_ob_out[3], \kme_cceip0_ob_out.tdata [3]);
tran (kme_cceip0_ob_out[2], \kme_cceip0_ob_out.tdata [2]);
tran (kme_cceip0_ob_out[1], \kme_cceip0_ob_out.tdata [1]);
tran (kme_cceip0_ob_out[0], \kme_cceip0_ob_out.tdata [0]);
tran (kme_cceip1_ob_out[82], \kme_cceip1_ob_out.tvalid );
tran (kme_cceip1_ob_out[81], \kme_cceip1_ob_out.tlast );
tran (kme_cceip1_ob_out[80], \kme_cceip1_ob_out.tid [0]);
tran (kme_cceip1_ob_out[79], \kme_cceip1_ob_out.tstrb [7]);
tran (kme_cceip1_ob_out[78], \kme_cceip1_ob_out.tstrb [6]);
tran (kme_cceip1_ob_out[77], \kme_cceip1_ob_out.tstrb [5]);
tran (kme_cceip1_ob_out[76], \kme_cceip1_ob_out.tstrb [4]);
tran (kme_cceip1_ob_out[75], \kme_cceip1_ob_out.tstrb [3]);
tran (kme_cceip1_ob_out[74], \kme_cceip1_ob_out.tstrb [2]);
tran (kme_cceip1_ob_out[73], \kme_cceip1_ob_out.tstrb [1]);
tran (kme_cceip1_ob_out[72], \kme_cceip1_ob_out.tstrb [0]);
tran (kme_cceip1_ob_out[71], \kme_cceip1_ob_out.tuser [7]);
tran (kme_cceip1_ob_out[70], \kme_cceip1_ob_out.tuser [6]);
tran (kme_cceip1_ob_out[69], \kme_cceip1_ob_out.tuser [5]);
tran (kme_cceip1_ob_out[68], \kme_cceip1_ob_out.tuser [4]);
tran (kme_cceip1_ob_out[67], \kme_cceip1_ob_out.tuser [3]);
tran (kme_cceip1_ob_out[66], \kme_cceip1_ob_out.tuser [2]);
tran (kme_cceip1_ob_out[65], \kme_cceip1_ob_out.tuser [1]);
tran (kme_cceip1_ob_out[64], \kme_cceip1_ob_out.tuser [0]);
tran (kme_cceip1_ob_out[63], \kme_cceip1_ob_out.tdata [63]);
tran (kme_cceip1_ob_out[62], \kme_cceip1_ob_out.tdata [62]);
tran (kme_cceip1_ob_out[61], \kme_cceip1_ob_out.tdata [61]);
tran (kme_cceip1_ob_out[60], \kme_cceip1_ob_out.tdata [60]);
tran (kme_cceip1_ob_out[59], \kme_cceip1_ob_out.tdata [59]);
tran (kme_cceip1_ob_out[58], \kme_cceip1_ob_out.tdata [58]);
tran (kme_cceip1_ob_out[57], \kme_cceip1_ob_out.tdata [57]);
tran (kme_cceip1_ob_out[56], \kme_cceip1_ob_out.tdata [56]);
tran (kme_cceip1_ob_out[55], \kme_cceip1_ob_out.tdata [55]);
tran (kme_cceip1_ob_out[54], \kme_cceip1_ob_out.tdata [54]);
tran (kme_cceip1_ob_out[53], \kme_cceip1_ob_out.tdata [53]);
tran (kme_cceip1_ob_out[52], \kme_cceip1_ob_out.tdata [52]);
tran (kme_cceip1_ob_out[51], \kme_cceip1_ob_out.tdata [51]);
tran (kme_cceip1_ob_out[50], \kme_cceip1_ob_out.tdata [50]);
tran (kme_cceip1_ob_out[49], \kme_cceip1_ob_out.tdata [49]);
tran (kme_cceip1_ob_out[48], \kme_cceip1_ob_out.tdata [48]);
tran (kme_cceip1_ob_out[47], \kme_cceip1_ob_out.tdata [47]);
tran (kme_cceip1_ob_out[46], \kme_cceip1_ob_out.tdata [46]);
tran (kme_cceip1_ob_out[45], \kme_cceip1_ob_out.tdata [45]);
tran (kme_cceip1_ob_out[44], \kme_cceip1_ob_out.tdata [44]);
tran (kme_cceip1_ob_out[43], \kme_cceip1_ob_out.tdata [43]);
tran (kme_cceip1_ob_out[42], \kme_cceip1_ob_out.tdata [42]);
tran (kme_cceip1_ob_out[41], \kme_cceip1_ob_out.tdata [41]);
tran (kme_cceip1_ob_out[40], \kme_cceip1_ob_out.tdata [40]);
tran (kme_cceip1_ob_out[39], \kme_cceip1_ob_out.tdata [39]);
tran (kme_cceip1_ob_out[38], \kme_cceip1_ob_out.tdata [38]);
tran (kme_cceip1_ob_out[37], \kme_cceip1_ob_out.tdata [37]);
tran (kme_cceip1_ob_out[36], \kme_cceip1_ob_out.tdata [36]);
tran (kme_cceip1_ob_out[35], \kme_cceip1_ob_out.tdata [35]);
tran (kme_cceip1_ob_out[34], \kme_cceip1_ob_out.tdata [34]);
tran (kme_cceip1_ob_out[33], \kme_cceip1_ob_out.tdata [33]);
tran (kme_cceip1_ob_out[32], \kme_cceip1_ob_out.tdata [32]);
tran (kme_cceip1_ob_out[31], \kme_cceip1_ob_out.tdata [31]);
tran (kme_cceip1_ob_out[30], \kme_cceip1_ob_out.tdata [30]);
tran (kme_cceip1_ob_out[29], \kme_cceip1_ob_out.tdata [29]);
tran (kme_cceip1_ob_out[28], \kme_cceip1_ob_out.tdata [28]);
tran (kme_cceip1_ob_out[27], \kme_cceip1_ob_out.tdata [27]);
tran (kme_cceip1_ob_out[26], \kme_cceip1_ob_out.tdata [26]);
tran (kme_cceip1_ob_out[25], \kme_cceip1_ob_out.tdata [25]);
tran (kme_cceip1_ob_out[24], \kme_cceip1_ob_out.tdata [24]);
tran (kme_cceip1_ob_out[23], \kme_cceip1_ob_out.tdata [23]);
tran (kme_cceip1_ob_out[22], \kme_cceip1_ob_out.tdata [22]);
tran (kme_cceip1_ob_out[21], \kme_cceip1_ob_out.tdata [21]);
tran (kme_cceip1_ob_out[20], \kme_cceip1_ob_out.tdata [20]);
tran (kme_cceip1_ob_out[19], \kme_cceip1_ob_out.tdata [19]);
tran (kme_cceip1_ob_out[18], \kme_cceip1_ob_out.tdata [18]);
tran (kme_cceip1_ob_out[17], \kme_cceip1_ob_out.tdata [17]);
tran (kme_cceip1_ob_out[16], \kme_cceip1_ob_out.tdata [16]);
tran (kme_cceip1_ob_out[15], \kme_cceip1_ob_out.tdata [15]);
tran (kme_cceip1_ob_out[14], \kme_cceip1_ob_out.tdata [14]);
tran (kme_cceip1_ob_out[13], \kme_cceip1_ob_out.tdata [13]);
tran (kme_cceip1_ob_out[12], \kme_cceip1_ob_out.tdata [12]);
tran (kme_cceip1_ob_out[11], \kme_cceip1_ob_out.tdata [11]);
tran (kme_cceip1_ob_out[10], \kme_cceip1_ob_out.tdata [10]);
tran (kme_cceip1_ob_out[9], \kme_cceip1_ob_out.tdata [9]);
tran (kme_cceip1_ob_out[8], \kme_cceip1_ob_out.tdata [8]);
tran (kme_cceip1_ob_out[7], \kme_cceip1_ob_out.tdata [7]);
tran (kme_cceip1_ob_out[6], \kme_cceip1_ob_out.tdata [6]);
tran (kme_cceip1_ob_out[5], \kme_cceip1_ob_out.tdata [5]);
tran (kme_cceip1_ob_out[4], \kme_cceip1_ob_out.tdata [4]);
tran (kme_cceip1_ob_out[3], \kme_cceip1_ob_out.tdata [3]);
tran (kme_cceip1_ob_out[2], \kme_cceip1_ob_out.tdata [2]);
tran (kme_cceip1_ob_out[1], \kme_cceip1_ob_out.tdata [1]);
tran (kme_cceip1_ob_out[0], \kme_cceip1_ob_out.tdata [0]);
tran (kme_cceip2_ob_out[82], \kme_cceip2_ob_out.tvalid );
tran (kme_cceip2_ob_out[81], \kme_cceip2_ob_out.tlast );
tran (kme_cceip2_ob_out[80], \kme_cceip2_ob_out.tid [0]);
tran (kme_cceip2_ob_out[79], \kme_cceip2_ob_out.tstrb [7]);
tran (kme_cceip2_ob_out[78], \kme_cceip2_ob_out.tstrb [6]);
tran (kme_cceip2_ob_out[77], \kme_cceip2_ob_out.tstrb [5]);
tran (kme_cceip2_ob_out[76], \kme_cceip2_ob_out.tstrb [4]);
tran (kme_cceip2_ob_out[75], \kme_cceip2_ob_out.tstrb [3]);
tran (kme_cceip2_ob_out[74], \kme_cceip2_ob_out.tstrb [2]);
tran (kme_cceip2_ob_out[73], \kme_cceip2_ob_out.tstrb [1]);
tran (kme_cceip2_ob_out[72], \kme_cceip2_ob_out.tstrb [0]);
tran (kme_cceip2_ob_out[71], \kme_cceip2_ob_out.tuser [7]);
tran (kme_cceip2_ob_out[70], \kme_cceip2_ob_out.tuser [6]);
tran (kme_cceip2_ob_out[69], \kme_cceip2_ob_out.tuser [5]);
tran (kme_cceip2_ob_out[68], \kme_cceip2_ob_out.tuser [4]);
tran (kme_cceip2_ob_out[67], \kme_cceip2_ob_out.tuser [3]);
tran (kme_cceip2_ob_out[66], \kme_cceip2_ob_out.tuser [2]);
tran (kme_cceip2_ob_out[65], \kme_cceip2_ob_out.tuser [1]);
tran (kme_cceip2_ob_out[64], \kme_cceip2_ob_out.tuser [0]);
tran (kme_cceip2_ob_out[63], \kme_cceip2_ob_out.tdata [63]);
tran (kme_cceip2_ob_out[62], \kme_cceip2_ob_out.tdata [62]);
tran (kme_cceip2_ob_out[61], \kme_cceip2_ob_out.tdata [61]);
tran (kme_cceip2_ob_out[60], \kme_cceip2_ob_out.tdata [60]);
tran (kme_cceip2_ob_out[59], \kme_cceip2_ob_out.tdata [59]);
tran (kme_cceip2_ob_out[58], \kme_cceip2_ob_out.tdata [58]);
tran (kme_cceip2_ob_out[57], \kme_cceip2_ob_out.tdata [57]);
tran (kme_cceip2_ob_out[56], \kme_cceip2_ob_out.tdata [56]);
tran (kme_cceip2_ob_out[55], \kme_cceip2_ob_out.tdata [55]);
tran (kme_cceip2_ob_out[54], \kme_cceip2_ob_out.tdata [54]);
tran (kme_cceip2_ob_out[53], \kme_cceip2_ob_out.tdata [53]);
tran (kme_cceip2_ob_out[52], \kme_cceip2_ob_out.tdata [52]);
tran (kme_cceip2_ob_out[51], \kme_cceip2_ob_out.tdata [51]);
tran (kme_cceip2_ob_out[50], \kme_cceip2_ob_out.tdata [50]);
tran (kme_cceip2_ob_out[49], \kme_cceip2_ob_out.tdata [49]);
tran (kme_cceip2_ob_out[48], \kme_cceip2_ob_out.tdata [48]);
tran (kme_cceip2_ob_out[47], \kme_cceip2_ob_out.tdata [47]);
tran (kme_cceip2_ob_out[46], \kme_cceip2_ob_out.tdata [46]);
tran (kme_cceip2_ob_out[45], \kme_cceip2_ob_out.tdata [45]);
tran (kme_cceip2_ob_out[44], \kme_cceip2_ob_out.tdata [44]);
tran (kme_cceip2_ob_out[43], \kme_cceip2_ob_out.tdata [43]);
tran (kme_cceip2_ob_out[42], \kme_cceip2_ob_out.tdata [42]);
tran (kme_cceip2_ob_out[41], \kme_cceip2_ob_out.tdata [41]);
tran (kme_cceip2_ob_out[40], \kme_cceip2_ob_out.tdata [40]);
tran (kme_cceip2_ob_out[39], \kme_cceip2_ob_out.tdata [39]);
tran (kme_cceip2_ob_out[38], \kme_cceip2_ob_out.tdata [38]);
tran (kme_cceip2_ob_out[37], \kme_cceip2_ob_out.tdata [37]);
tran (kme_cceip2_ob_out[36], \kme_cceip2_ob_out.tdata [36]);
tran (kme_cceip2_ob_out[35], \kme_cceip2_ob_out.tdata [35]);
tran (kme_cceip2_ob_out[34], \kme_cceip2_ob_out.tdata [34]);
tran (kme_cceip2_ob_out[33], \kme_cceip2_ob_out.tdata [33]);
tran (kme_cceip2_ob_out[32], \kme_cceip2_ob_out.tdata [32]);
tran (kme_cceip2_ob_out[31], \kme_cceip2_ob_out.tdata [31]);
tran (kme_cceip2_ob_out[30], \kme_cceip2_ob_out.tdata [30]);
tran (kme_cceip2_ob_out[29], \kme_cceip2_ob_out.tdata [29]);
tran (kme_cceip2_ob_out[28], \kme_cceip2_ob_out.tdata [28]);
tran (kme_cceip2_ob_out[27], \kme_cceip2_ob_out.tdata [27]);
tran (kme_cceip2_ob_out[26], \kme_cceip2_ob_out.tdata [26]);
tran (kme_cceip2_ob_out[25], \kme_cceip2_ob_out.tdata [25]);
tran (kme_cceip2_ob_out[24], \kme_cceip2_ob_out.tdata [24]);
tran (kme_cceip2_ob_out[23], \kme_cceip2_ob_out.tdata [23]);
tran (kme_cceip2_ob_out[22], \kme_cceip2_ob_out.tdata [22]);
tran (kme_cceip2_ob_out[21], \kme_cceip2_ob_out.tdata [21]);
tran (kme_cceip2_ob_out[20], \kme_cceip2_ob_out.tdata [20]);
tran (kme_cceip2_ob_out[19], \kme_cceip2_ob_out.tdata [19]);
tran (kme_cceip2_ob_out[18], \kme_cceip2_ob_out.tdata [18]);
tran (kme_cceip2_ob_out[17], \kme_cceip2_ob_out.tdata [17]);
tran (kme_cceip2_ob_out[16], \kme_cceip2_ob_out.tdata [16]);
tran (kme_cceip2_ob_out[15], \kme_cceip2_ob_out.tdata [15]);
tran (kme_cceip2_ob_out[14], \kme_cceip2_ob_out.tdata [14]);
tran (kme_cceip2_ob_out[13], \kme_cceip2_ob_out.tdata [13]);
tran (kme_cceip2_ob_out[12], \kme_cceip2_ob_out.tdata [12]);
tran (kme_cceip2_ob_out[11], \kme_cceip2_ob_out.tdata [11]);
tran (kme_cceip2_ob_out[10], \kme_cceip2_ob_out.tdata [10]);
tran (kme_cceip2_ob_out[9], \kme_cceip2_ob_out.tdata [9]);
tran (kme_cceip2_ob_out[8], \kme_cceip2_ob_out.tdata [8]);
tran (kme_cceip2_ob_out[7], \kme_cceip2_ob_out.tdata [7]);
tran (kme_cceip2_ob_out[6], \kme_cceip2_ob_out.tdata [6]);
tran (kme_cceip2_ob_out[5], \kme_cceip2_ob_out.tdata [5]);
tran (kme_cceip2_ob_out[4], \kme_cceip2_ob_out.tdata [4]);
tran (kme_cceip2_ob_out[3], \kme_cceip2_ob_out.tdata [3]);
tran (kme_cceip2_ob_out[2], \kme_cceip2_ob_out.tdata [2]);
tran (kme_cceip2_ob_out[1], \kme_cceip2_ob_out.tdata [1]);
tran (kme_cceip2_ob_out[0], \kme_cceip2_ob_out.tdata [0]);
tran (kme_cceip3_ob_out[82], \kme_cceip3_ob_out.tvalid );
tran (kme_cceip3_ob_out[81], \kme_cceip3_ob_out.tlast );
tran (kme_cceip3_ob_out[80], \kme_cceip3_ob_out.tid [0]);
tran (kme_cceip3_ob_out[79], \kme_cceip3_ob_out.tstrb [7]);
tran (kme_cceip3_ob_out[78], \kme_cceip3_ob_out.tstrb [6]);
tran (kme_cceip3_ob_out[77], \kme_cceip3_ob_out.tstrb [5]);
tran (kme_cceip3_ob_out[76], \kme_cceip3_ob_out.tstrb [4]);
tran (kme_cceip3_ob_out[75], \kme_cceip3_ob_out.tstrb [3]);
tran (kme_cceip3_ob_out[74], \kme_cceip3_ob_out.tstrb [2]);
tran (kme_cceip3_ob_out[73], \kme_cceip3_ob_out.tstrb [1]);
tran (kme_cceip3_ob_out[72], \kme_cceip3_ob_out.tstrb [0]);
tran (kme_cceip3_ob_out[71], \kme_cceip3_ob_out.tuser [7]);
tran (kme_cceip3_ob_out[70], \kme_cceip3_ob_out.tuser [6]);
tran (kme_cceip3_ob_out[69], \kme_cceip3_ob_out.tuser [5]);
tran (kme_cceip3_ob_out[68], \kme_cceip3_ob_out.tuser [4]);
tran (kme_cceip3_ob_out[67], \kme_cceip3_ob_out.tuser [3]);
tran (kme_cceip3_ob_out[66], \kme_cceip3_ob_out.tuser [2]);
tran (kme_cceip3_ob_out[65], \kme_cceip3_ob_out.tuser [1]);
tran (kme_cceip3_ob_out[64], \kme_cceip3_ob_out.tuser [0]);
tran (kme_cceip3_ob_out[63], \kme_cceip3_ob_out.tdata [63]);
tran (kme_cceip3_ob_out[62], \kme_cceip3_ob_out.tdata [62]);
tran (kme_cceip3_ob_out[61], \kme_cceip3_ob_out.tdata [61]);
tran (kme_cceip3_ob_out[60], \kme_cceip3_ob_out.tdata [60]);
tran (kme_cceip3_ob_out[59], \kme_cceip3_ob_out.tdata [59]);
tran (kme_cceip3_ob_out[58], \kme_cceip3_ob_out.tdata [58]);
tran (kme_cceip3_ob_out[57], \kme_cceip3_ob_out.tdata [57]);
tran (kme_cceip3_ob_out[56], \kme_cceip3_ob_out.tdata [56]);
tran (kme_cceip3_ob_out[55], \kme_cceip3_ob_out.tdata [55]);
tran (kme_cceip3_ob_out[54], \kme_cceip3_ob_out.tdata [54]);
tran (kme_cceip3_ob_out[53], \kme_cceip3_ob_out.tdata [53]);
tran (kme_cceip3_ob_out[52], \kme_cceip3_ob_out.tdata [52]);
tran (kme_cceip3_ob_out[51], \kme_cceip3_ob_out.tdata [51]);
tran (kme_cceip3_ob_out[50], \kme_cceip3_ob_out.tdata [50]);
tran (kme_cceip3_ob_out[49], \kme_cceip3_ob_out.tdata [49]);
tran (kme_cceip3_ob_out[48], \kme_cceip3_ob_out.tdata [48]);
tran (kme_cceip3_ob_out[47], \kme_cceip3_ob_out.tdata [47]);
tran (kme_cceip3_ob_out[46], \kme_cceip3_ob_out.tdata [46]);
tran (kme_cceip3_ob_out[45], \kme_cceip3_ob_out.tdata [45]);
tran (kme_cceip3_ob_out[44], \kme_cceip3_ob_out.tdata [44]);
tran (kme_cceip3_ob_out[43], \kme_cceip3_ob_out.tdata [43]);
tran (kme_cceip3_ob_out[42], \kme_cceip3_ob_out.tdata [42]);
tran (kme_cceip3_ob_out[41], \kme_cceip3_ob_out.tdata [41]);
tran (kme_cceip3_ob_out[40], \kme_cceip3_ob_out.tdata [40]);
tran (kme_cceip3_ob_out[39], \kme_cceip3_ob_out.tdata [39]);
tran (kme_cceip3_ob_out[38], \kme_cceip3_ob_out.tdata [38]);
tran (kme_cceip3_ob_out[37], \kme_cceip3_ob_out.tdata [37]);
tran (kme_cceip3_ob_out[36], \kme_cceip3_ob_out.tdata [36]);
tran (kme_cceip3_ob_out[35], \kme_cceip3_ob_out.tdata [35]);
tran (kme_cceip3_ob_out[34], \kme_cceip3_ob_out.tdata [34]);
tran (kme_cceip3_ob_out[33], \kme_cceip3_ob_out.tdata [33]);
tran (kme_cceip3_ob_out[32], \kme_cceip3_ob_out.tdata [32]);
tran (kme_cceip3_ob_out[31], \kme_cceip3_ob_out.tdata [31]);
tran (kme_cceip3_ob_out[30], \kme_cceip3_ob_out.tdata [30]);
tran (kme_cceip3_ob_out[29], \kme_cceip3_ob_out.tdata [29]);
tran (kme_cceip3_ob_out[28], \kme_cceip3_ob_out.tdata [28]);
tran (kme_cceip3_ob_out[27], \kme_cceip3_ob_out.tdata [27]);
tran (kme_cceip3_ob_out[26], \kme_cceip3_ob_out.tdata [26]);
tran (kme_cceip3_ob_out[25], \kme_cceip3_ob_out.tdata [25]);
tran (kme_cceip3_ob_out[24], \kme_cceip3_ob_out.tdata [24]);
tran (kme_cceip3_ob_out[23], \kme_cceip3_ob_out.tdata [23]);
tran (kme_cceip3_ob_out[22], \kme_cceip3_ob_out.tdata [22]);
tran (kme_cceip3_ob_out[21], \kme_cceip3_ob_out.tdata [21]);
tran (kme_cceip3_ob_out[20], \kme_cceip3_ob_out.tdata [20]);
tran (kme_cceip3_ob_out[19], \kme_cceip3_ob_out.tdata [19]);
tran (kme_cceip3_ob_out[18], \kme_cceip3_ob_out.tdata [18]);
tran (kme_cceip3_ob_out[17], \kme_cceip3_ob_out.tdata [17]);
tran (kme_cceip3_ob_out[16], \kme_cceip3_ob_out.tdata [16]);
tran (kme_cceip3_ob_out[15], \kme_cceip3_ob_out.tdata [15]);
tran (kme_cceip3_ob_out[14], \kme_cceip3_ob_out.tdata [14]);
tran (kme_cceip3_ob_out[13], \kme_cceip3_ob_out.tdata [13]);
tran (kme_cceip3_ob_out[12], \kme_cceip3_ob_out.tdata [12]);
tran (kme_cceip3_ob_out[11], \kme_cceip3_ob_out.tdata [11]);
tran (kme_cceip3_ob_out[10], \kme_cceip3_ob_out.tdata [10]);
tran (kme_cceip3_ob_out[9], \kme_cceip3_ob_out.tdata [9]);
tran (kme_cceip3_ob_out[8], \kme_cceip3_ob_out.tdata [8]);
tran (kme_cceip3_ob_out[7], \kme_cceip3_ob_out.tdata [7]);
tran (kme_cceip3_ob_out[6], \kme_cceip3_ob_out.tdata [6]);
tran (kme_cceip3_ob_out[5], \kme_cceip3_ob_out.tdata [5]);
tran (kme_cceip3_ob_out[4], \kme_cceip3_ob_out.tdata [4]);
tran (kme_cceip3_ob_out[3], \kme_cceip3_ob_out.tdata [3]);
tran (kme_cceip3_ob_out[2], \kme_cceip3_ob_out.tdata [2]);
tran (kme_cceip3_ob_out[1], \kme_cceip3_ob_out.tdata [1]);
tran (kme_cceip3_ob_out[0], \kme_cceip3_ob_out.tdata [0]);
tran (kme_cddip0_ob_out[82], \kme_cddip0_ob_out.tvalid );
tran (kme_cddip0_ob_out[81], \kme_cddip0_ob_out.tlast );
tran (kme_cddip0_ob_out[80], \kme_cddip0_ob_out.tid [0]);
tran (kme_cddip0_ob_out[79], \kme_cddip0_ob_out.tstrb [7]);
tran (kme_cddip0_ob_out[78], \kme_cddip0_ob_out.tstrb [6]);
tran (kme_cddip0_ob_out[77], \kme_cddip0_ob_out.tstrb [5]);
tran (kme_cddip0_ob_out[76], \kme_cddip0_ob_out.tstrb [4]);
tran (kme_cddip0_ob_out[75], \kme_cddip0_ob_out.tstrb [3]);
tran (kme_cddip0_ob_out[74], \kme_cddip0_ob_out.tstrb [2]);
tran (kme_cddip0_ob_out[73], \kme_cddip0_ob_out.tstrb [1]);
tran (kme_cddip0_ob_out[72], \kme_cddip0_ob_out.tstrb [0]);
tran (kme_cddip0_ob_out[71], \kme_cddip0_ob_out.tuser [7]);
tran (kme_cddip0_ob_out[70], \kme_cddip0_ob_out.tuser [6]);
tran (kme_cddip0_ob_out[69], \kme_cddip0_ob_out.tuser [5]);
tran (kme_cddip0_ob_out[68], \kme_cddip0_ob_out.tuser [4]);
tran (kme_cddip0_ob_out[67], \kme_cddip0_ob_out.tuser [3]);
tran (kme_cddip0_ob_out[66], \kme_cddip0_ob_out.tuser [2]);
tran (kme_cddip0_ob_out[65], \kme_cddip0_ob_out.tuser [1]);
tran (kme_cddip0_ob_out[64], \kme_cddip0_ob_out.tuser [0]);
tran (kme_cddip0_ob_out[63], \kme_cddip0_ob_out.tdata [63]);
tran (kme_cddip0_ob_out[62], \kme_cddip0_ob_out.tdata [62]);
tran (kme_cddip0_ob_out[61], \kme_cddip0_ob_out.tdata [61]);
tran (kme_cddip0_ob_out[60], \kme_cddip0_ob_out.tdata [60]);
tran (kme_cddip0_ob_out[59], \kme_cddip0_ob_out.tdata [59]);
tran (kme_cddip0_ob_out[58], \kme_cddip0_ob_out.tdata [58]);
tran (kme_cddip0_ob_out[57], \kme_cddip0_ob_out.tdata [57]);
tran (kme_cddip0_ob_out[56], \kme_cddip0_ob_out.tdata [56]);
tran (kme_cddip0_ob_out[55], \kme_cddip0_ob_out.tdata [55]);
tran (kme_cddip0_ob_out[54], \kme_cddip0_ob_out.tdata [54]);
tran (kme_cddip0_ob_out[53], \kme_cddip0_ob_out.tdata [53]);
tran (kme_cddip0_ob_out[52], \kme_cddip0_ob_out.tdata [52]);
tran (kme_cddip0_ob_out[51], \kme_cddip0_ob_out.tdata [51]);
tran (kme_cddip0_ob_out[50], \kme_cddip0_ob_out.tdata [50]);
tran (kme_cddip0_ob_out[49], \kme_cddip0_ob_out.tdata [49]);
tran (kme_cddip0_ob_out[48], \kme_cddip0_ob_out.tdata [48]);
tran (kme_cddip0_ob_out[47], \kme_cddip0_ob_out.tdata [47]);
tran (kme_cddip0_ob_out[46], \kme_cddip0_ob_out.tdata [46]);
tran (kme_cddip0_ob_out[45], \kme_cddip0_ob_out.tdata [45]);
tran (kme_cddip0_ob_out[44], \kme_cddip0_ob_out.tdata [44]);
tran (kme_cddip0_ob_out[43], \kme_cddip0_ob_out.tdata [43]);
tran (kme_cddip0_ob_out[42], \kme_cddip0_ob_out.tdata [42]);
tran (kme_cddip0_ob_out[41], \kme_cddip0_ob_out.tdata [41]);
tran (kme_cddip0_ob_out[40], \kme_cddip0_ob_out.tdata [40]);
tran (kme_cddip0_ob_out[39], \kme_cddip0_ob_out.tdata [39]);
tran (kme_cddip0_ob_out[38], \kme_cddip0_ob_out.tdata [38]);
tran (kme_cddip0_ob_out[37], \kme_cddip0_ob_out.tdata [37]);
tran (kme_cddip0_ob_out[36], \kme_cddip0_ob_out.tdata [36]);
tran (kme_cddip0_ob_out[35], \kme_cddip0_ob_out.tdata [35]);
tran (kme_cddip0_ob_out[34], \kme_cddip0_ob_out.tdata [34]);
tran (kme_cddip0_ob_out[33], \kme_cddip0_ob_out.tdata [33]);
tran (kme_cddip0_ob_out[32], \kme_cddip0_ob_out.tdata [32]);
tran (kme_cddip0_ob_out[31], \kme_cddip0_ob_out.tdata [31]);
tran (kme_cddip0_ob_out[30], \kme_cddip0_ob_out.tdata [30]);
tran (kme_cddip0_ob_out[29], \kme_cddip0_ob_out.tdata [29]);
tran (kme_cddip0_ob_out[28], \kme_cddip0_ob_out.tdata [28]);
tran (kme_cddip0_ob_out[27], \kme_cddip0_ob_out.tdata [27]);
tran (kme_cddip0_ob_out[26], \kme_cddip0_ob_out.tdata [26]);
tran (kme_cddip0_ob_out[25], \kme_cddip0_ob_out.tdata [25]);
tran (kme_cddip0_ob_out[24], \kme_cddip0_ob_out.tdata [24]);
tran (kme_cddip0_ob_out[23], \kme_cddip0_ob_out.tdata [23]);
tran (kme_cddip0_ob_out[22], \kme_cddip0_ob_out.tdata [22]);
tran (kme_cddip0_ob_out[21], \kme_cddip0_ob_out.tdata [21]);
tran (kme_cddip0_ob_out[20], \kme_cddip0_ob_out.tdata [20]);
tran (kme_cddip0_ob_out[19], \kme_cddip0_ob_out.tdata [19]);
tran (kme_cddip0_ob_out[18], \kme_cddip0_ob_out.tdata [18]);
tran (kme_cddip0_ob_out[17], \kme_cddip0_ob_out.tdata [17]);
tran (kme_cddip0_ob_out[16], \kme_cddip0_ob_out.tdata [16]);
tran (kme_cddip0_ob_out[15], \kme_cddip0_ob_out.tdata [15]);
tran (kme_cddip0_ob_out[14], \kme_cddip0_ob_out.tdata [14]);
tran (kme_cddip0_ob_out[13], \kme_cddip0_ob_out.tdata [13]);
tran (kme_cddip0_ob_out[12], \kme_cddip0_ob_out.tdata [12]);
tran (kme_cddip0_ob_out[11], \kme_cddip0_ob_out.tdata [11]);
tran (kme_cddip0_ob_out[10], \kme_cddip0_ob_out.tdata [10]);
tran (kme_cddip0_ob_out[9], \kme_cddip0_ob_out.tdata [9]);
tran (kme_cddip0_ob_out[8], \kme_cddip0_ob_out.tdata [8]);
tran (kme_cddip0_ob_out[7], \kme_cddip0_ob_out.tdata [7]);
tran (kme_cddip0_ob_out[6], \kme_cddip0_ob_out.tdata [6]);
tran (kme_cddip0_ob_out[5], \kme_cddip0_ob_out.tdata [5]);
tran (kme_cddip0_ob_out[4], \kme_cddip0_ob_out.tdata [4]);
tran (kme_cddip0_ob_out[3], \kme_cddip0_ob_out.tdata [3]);
tran (kme_cddip0_ob_out[2], \kme_cddip0_ob_out.tdata [2]);
tran (kme_cddip0_ob_out[1], \kme_cddip0_ob_out.tdata [1]);
tran (kme_cddip0_ob_out[0], \kme_cddip0_ob_out.tdata [0]);
tran (kme_cddip1_ob_out[82], \kme_cddip1_ob_out.tvalid );
tran (kme_cddip1_ob_out[81], \kme_cddip1_ob_out.tlast );
tran (kme_cddip1_ob_out[80], \kme_cddip1_ob_out.tid [0]);
tran (kme_cddip1_ob_out[79], \kme_cddip1_ob_out.tstrb [7]);
tran (kme_cddip1_ob_out[78], \kme_cddip1_ob_out.tstrb [6]);
tran (kme_cddip1_ob_out[77], \kme_cddip1_ob_out.tstrb [5]);
tran (kme_cddip1_ob_out[76], \kme_cddip1_ob_out.tstrb [4]);
tran (kme_cddip1_ob_out[75], \kme_cddip1_ob_out.tstrb [3]);
tran (kme_cddip1_ob_out[74], \kme_cddip1_ob_out.tstrb [2]);
tran (kme_cddip1_ob_out[73], \kme_cddip1_ob_out.tstrb [1]);
tran (kme_cddip1_ob_out[72], \kme_cddip1_ob_out.tstrb [0]);
tran (kme_cddip1_ob_out[71], \kme_cddip1_ob_out.tuser [7]);
tran (kme_cddip1_ob_out[70], \kme_cddip1_ob_out.tuser [6]);
tran (kme_cddip1_ob_out[69], \kme_cddip1_ob_out.tuser [5]);
tran (kme_cddip1_ob_out[68], \kme_cddip1_ob_out.tuser [4]);
tran (kme_cddip1_ob_out[67], \kme_cddip1_ob_out.tuser [3]);
tran (kme_cddip1_ob_out[66], \kme_cddip1_ob_out.tuser [2]);
tran (kme_cddip1_ob_out[65], \kme_cddip1_ob_out.tuser [1]);
tran (kme_cddip1_ob_out[64], \kme_cddip1_ob_out.tuser [0]);
tran (kme_cddip1_ob_out[63], \kme_cddip1_ob_out.tdata [63]);
tran (kme_cddip1_ob_out[62], \kme_cddip1_ob_out.tdata [62]);
tran (kme_cddip1_ob_out[61], \kme_cddip1_ob_out.tdata [61]);
tran (kme_cddip1_ob_out[60], \kme_cddip1_ob_out.tdata [60]);
tran (kme_cddip1_ob_out[59], \kme_cddip1_ob_out.tdata [59]);
tran (kme_cddip1_ob_out[58], \kme_cddip1_ob_out.tdata [58]);
tran (kme_cddip1_ob_out[57], \kme_cddip1_ob_out.tdata [57]);
tran (kme_cddip1_ob_out[56], \kme_cddip1_ob_out.tdata [56]);
tran (kme_cddip1_ob_out[55], \kme_cddip1_ob_out.tdata [55]);
tran (kme_cddip1_ob_out[54], \kme_cddip1_ob_out.tdata [54]);
tran (kme_cddip1_ob_out[53], \kme_cddip1_ob_out.tdata [53]);
tran (kme_cddip1_ob_out[52], \kme_cddip1_ob_out.tdata [52]);
tran (kme_cddip1_ob_out[51], \kme_cddip1_ob_out.tdata [51]);
tran (kme_cddip1_ob_out[50], \kme_cddip1_ob_out.tdata [50]);
tran (kme_cddip1_ob_out[49], \kme_cddip1_ob_out.tdata [49]);
tran (kme_cddip1_ob_out[48], \kme_cddip1_ob_out.tdata [48]);
tran (kme_cddip1_ob_out[47], \kme_cddip1_ob_out.tdata [47]);
tran (kme_cddip1_ob_out[46], \kme_cddip1_ob_out.tdata [46]);
tran (kme_cddip1_ob_out[45], \kme_cddip1_ob_out.tdata [45]);
tran (kme_cddip1_ob_out[44], \kme_cddip1_ob_out.tdata [44]);
tran (kme_cddip1_ob_out[43], \kme_cddip1_ob_out.tdata [43]);
tran (kme_cddip1_ob_out[42], \kme_cddip1_ob_out.tdata [42]);
tran (kme_cddip1_ob_out[41], \kme_cddip1_ob_out.tdata [41]);
tran (kme_cddip1_ob_out[40], \kme_cddip1_ob_out.tdata [40]);
tran (kme_cddip1_ob_out[39], \kme_cddip1_ob_out.tdata [39]);
tran (kme_cddip1_ob_out[38], \kme_cddip1_ob_out.tdata [38]);
tran (kme_cddip1_ob_out[37], \kme_cddip1_ob_out.tdata [37]);
tran (kme_cddip1_ob_out[36], \kme_cddip1_ob_out.tdata [36]);
tran (kme_cddip1_ob_out[35], \kme_cddip1_ob_out.tdata [35]);
tran (kme_cddip1_ob_out[34], \kme_cddip1_ob_out.tdata [34]);
tran (kme_cddip1_ob_out[33], \kme_cddip1_ob_out.tdata [33]);
tran (kme_cddip1_ob_out[32], \kme_cddip1_ob_out.tdata [32]);
tran (kme_cddip1_ob_out[31], \kme_cddip1_ob_out.tdata [31]);
tran (kme_cddip1_ob_out[30], \kme_cddip1_ob_out.tdata [30]);
tran (kme_cddip1_ob_out[29], \kme_cddip1_ob_out.tdata [29]);
tran (kme_cddip1_ob_out[28], \kme_cddip1_ob_out.tdata [28]);
tran (kme_cddip1_ob_out[27], \kme_cddip1_ob_out.tdata [27]);
tran (kme_cddip1_ob_out[26], \kme_cddip1_ob_out.tdata [26]);
tran (kme_cddip1_ob_out[25], \kme_cddip1_ob_out.tdata [25]);
tran (kme_cddip1_ob_out[24], \kme_cddip1_ob_out.tdata [24]);
tran (kme_cddip1_ob_out[23], \kme_cddip1_ob_out.tdata [23]);
tran (kme_cddip1_ob_out[22], \kme_cddip1_ob_out.tdata [22]);
tran (kme_cddip1_ob_out[21], \kme_cddip1_ob_out.tdata [21]);
tran (kme_cddip1_ob_out[20], \kme_cddip1_ob_out.tdata [20]);
tran (kme_cddip1_ob_out[19], \kme_cddip1_ob_out.tdata [19]);
tran (kme_cddip1_ob_out[18], \kme_cddip1_ob_out.tdata [18]);
tran (kme_cddip1_ob_out[17], \kme_cddip1_ob_out.tdata [17]);
tran (kme_cddip1_ob_out[16], \kme_cddip1_ob_out.tdata [16]);
tran (kme_cddip1_ob_out[15], \kme_cddip1_ob_out.tdata [15]);
tran (kme_cddip1_ob_out[14], \kme_cddip1_ob_out.tdata [14]);
tran (kme_cddip1_ob_out[13], \kme_cddip1_ob_out.tdata [13]);
tran (kme_cddip1_ob_out[12], \kme_cddip1_ob_out.tdata [12]);
tran (kme_cddip1_ob_out[11], \kme_cddip1_ob_out.tdata [11]);
tran (kme_cddip1_ob_out[10], \kme_cddip1_ob_out.tdata [10]);
tran (kme_cddip1_ob_out[9], \kme_cddip1_ob_out.tdata [9]);
tran (kme_cddip1_ob_out[8], \kme_cddip1_ob_out.tdata [8]);
tran (kme_cddip1_ob_out[7], \kme_cddip1_ob_out.tdata [7]);
tran (kme_cddip1_ob_out[6], \kme_cddip1_ob_out.tdata [6]);
tran (kme_cddip1_ob_out[5], \kme_cddip1_ob_out.tdata [5]);
tran (kme_cddip1_ob_out[4], \kme_cddip1_ob_out.tdata [4]);
tran (kme_cddip1_ob_out[3], \kme_cddip1_ob_out.tdata [3]);
tran (kme_cddip1_ob_out[2], \kme_cddip1_ob_out.tdata [2]);
tran (kme_cddip1_ob_out[1], \kme_cddip1_ob_out.tdata [1]);
tran (kme_cddip1_ob_out[0], \kme_cddip1_ob_out.tdata [0]);
tran (kme_cddip2_ob_out[82], \kme_cddip2_ob_out.tvalid );
tran (kme_cddip2_ob_out[81], \kme_cddip2_ob_out.tlast );
tran (kme_cddip2_ob_out[80], \kme_cddip2_ob_out.tid [0]);
tran (kme_cddip2_ob_out[79], \kme_cddip2_ob_out.tstrb [7]);
tran (kme_cddip2_ob_out[78], \kme_cddip2_ob_out.tstrb [6]);
tran (kme_cddip2_ob_out[77], \kme_cddip2_ob_out.tstrb [5]);
tran (kme_cddip2_ob_out[76], \kme_cddip2_ob_out.tstrb [4]);
tran (kme_cddip2_ob_out[75], \kme_cddip2_ob_out.tstrb [3]);
tran (kme_cddip2_ob_out[74], \kme_cddip2_ob_out.tstrb [2]);
tran (kme_cddip2_ob_out[73], \kme_cddip2_ob_out.tstrb [1]);
tran (kme_cddip2_ob_out[72], \kme_cddip2_ob_out.tstrb [0]);
tran (kme_cddip2_ob_out[71], \kme_cddip2_ob_out.tuser [7]);
tran (kme_cddip2_ob_out[70], \kme_cddip2_ob_out.tuser [6]);
tran (kme_cddip2_ob_out[69], \kme_cddip2_ob_out.tuser [5]);
tran (kme_cddip2_ob_out[68], \kme_cddip2_ob_out.tuser [4]);
tran (kme_cddip2_ob_out[67], \kme_cddip2_ob_out.tuser [3]);
tran (kme_cddip2_ob_out[66], \kme_cddip2_ob_out.tuser [2]);
tran (kme_cddip2_ob_out[65], \kme_cddip2_ob_out.tuser [1]);
tran (kme_cddip2_ob_out[64], \kme_cddip2_ob_out.tuser [0]);
tran (kme_cddip2_ob_out[63], \kme_cddip2_ob_out.tdata [63]);
tran (kme_cddip2_ob_out[62], \kme_cddip2_ob_out.tdata [62]);
tran (kme_cddip2_ob_out[61], \kme_cddip2_ob_out.tdata [61]);
tran (kme_cddip2_ob_out[60], \kme_cddip2_ob_out.tdata [60]);
tran (kme_cddip2_ob_out[59], \kme_cddip2_ob_out.tdata [59]);
tran (kme_cddip2_ob_out[58], \kme_cddip2_ob_out.tdata [58]);
tran (kme_cddip2_ob_out[57], \kme_cddip2_ob_out.tdata [57]);
tran (kme_cddip2_ob_out[56], \kme_cddip2_ob_out.tdata [56]);
tran (kme_cddip2_ob_out[55], \kme_cddip2_ob_out.tdata [55]);
tran (kme_cddip2_ob_out[54], \kme_cddip2_ob_out.tdata [54]);
tran (kme_cddip2_ob_out[53], \kme_cddip2_ob_out.tdata [53]);
tran (kme_cddip2_ob_out[52], \kme_cddip2_ob_out.tdata [52]);
tran (kme_cddip2_ob_out[51], \kme_cddip2_ob_out.tdata [51]);
tran (kme_cddip2_ob_out[50], \kme_cddip2_ob_out.tdata [50]);
tran (kme_cddip2_ob_out[49], \kme_cddip2_ob_out.tdata [49]);
tran (kme_cddip2_ob_out[48], \kme_cddip2_ob_out.tdata [48]);
tran (kme_cddip2_ob_out[47], \kme_cddip2_ob_out.tdata [47]);
tran (kme_cddip2_ob_out[46], \kme_cddip2_ob_out.tdata [46]);
tran (kme_cddip2_ob_out[45], \kme_cddip2_ob_out.tdata [45]);
tran (kme_cddip2_ob_out[44], \kme_cddip2_ob_out.tdata [44]);
tran (kme_cddip2_ob_out[43], \kme_cddip2_ob_out.tdata [43]);
tran (kme_cddip2_ob_out[42], \kme_cddip2_ob_out.tdata [42]);
tran (kme_cddip2_ob_out[41], \kme_cddip2_ob_out.tdata [41]);
tran (kme_cddip2_ob_out[40], \kme_cddip2_ob_out.tdata [40]);
tran (kme_cddip2_ob_out[39], \kme_cddip2_ob_out.tdata [39]);
tran (kme_cddip2_ob_out[38], \kme_cddip2_ob_out.tdata [38]);
tran (kme_cddip2_ob_out[37], \kme_cddip2_ob_out.tdata [37]);
tran (kme_cddip2_ob_out[36], \kme_cddip2_ob_out.tdata [36]);
tran (kme_cddip2_ob_out[35], \kme_cddip2_ob_out.tdata [35]);
tran (kme_cddip2_ob_out[34], \kme_cddip2_ob_out.tdata [34]);
tran (kme_cddip2_ob_out[33], \kme_cddip2_ob_out.tdata [33]);
tran (kme_cddip2_ob_out[32], \kme_cddip2_ob_out.tdata [32]);
tran (kme_cddip2_ob_out[31], \kme_cddip2_ob_out.tdata [31]);
tran (kme_cddip2_ob_out[30], \kme_cddip2_ob_out.tdata [30]);
tran (kme_cddip2_ob_out[29], \kme_cddip2_ob_out.tdata [29]);
tran (kme_cddip2_ob_out[28], \kme_cddip2_ob_out.tdata [28]);
tran (kme_cddip2_ob_out[27], \kme_cddip2_ob_out.tdata [27]);
tran (kme_cddip2_ob_out[26], \kme_cddip2_ob_out.tdata [26]);
tran (kme_cddip2_ob_out[25], \kme_cddip2_ob_out.tdata [25]);
tran (kme_cddip2_ob_out[24], \kme_cddip2_ob_out.tdata [24]);
tran (kme_cddip2_ob_out[23], \kme_cddip2_ob_out.tdata [23]);
tran (kme_cddip2_ob_out[22], \kme_cddip2_ob_out.tdata [22]);
tran (kme_cddip2_ob_out[21], \kme_cddip2_ob_out.tdata [21]);
tran (kme_cddip2_ob_out[20], \kme_cddip2_ob_out.tdata [20]);
tran (kme_cddip2_ob_out[19], \kme_cddip2_ob_out.tdata [19]);
tran (kme_cddip2_ob_out[18], \kme_cddip2_ob_out.tdata [18]);
tran (kme_cddip2_ob_out[17], \kme_cddip2_ob_out.tdata [17]);
tran (kme_cddip2_ob_out[16], \kme_cddip2_ob_out.tdata [16]);
tran (kme_cddip2_ob_out[15], \kme_cddip2_ob_out.tdata [15]);
tran (kme_cddip2_ob_out[14], \kme_cddip2_ob_out.tdata [14]);
tran (kme_cddip2_ob_out[13], \kme_cddip2_ob_out.tdata [13]);
tran (kme_cddip2_ob_out[12], \kme_cddip2_ob_out.tdata [12]);
tran (kme_cddip2_ob_out[11], \kme_cddip2_ob_out.tdata [11]);
tran (kme_cddip2_ob_out[10], \kme_cddip2_ob_out.tdata [10]);
tran (kme_cddip2_ob_out[9], \kme_cddip2_ob_out.tdata [9]);
tran (kme_cddip2_ob_out[8], \kme_cddip2_ob_out.tdata [8]);
tran (kme_cddip2_ob_out[7], \kme_cddip2_ob_out.tdata [7]);
tran (kme_cddip2_ob_out[6], \kme_cddip2_ob_out.tdata [6]);
tran (kme_cddip2_ob_out[5], \kme_cddip2_ob_out.tdata [5]);
tran (kme_cddip2_ob_out[4], \kme_cddip2_ob_out.tdata [4]);
tran (kme_cddip2_ob_out[3], \kme_cddip2_ob_out.tdata [3]);
tran (kme_cddip2_ob_out[2], \kme_cddip2_ob_out.tdata [2]);
tran (kme_cddip2_ob_out[1], \kme_cddip2_ob_out.tdata [1]);
tran (kme_cddip2_ob_out[0], \kme_cddip2_ob_out.tdata [0]);
tran (kme_cddip3_ob_out[82], \kme_cddip3_ob_out.tvalid );
tran (kme_cddip3_ob_out[81], \kme_cddip3_ob_out.tlast );
tran (kme_cddip3_ob_out[80], \kme_cddip3_ob_out.tid [0]);
tran (kme_cddip3_ob_out[79], \kme_cddip3_ob_out.tstrb [7]);
tran (kme_cddip3_ob_out[78], \kme_cddip3_ob_out.tstrb [6]);
tran (kme_cddip3_ob_out[77], \kme_cddip3_ob_out.tstrb [5]);
tran (kme_cddip3_ob_out[76], \kme_cddip3_ob_out.tstrb [4]);
tran (kme_cddip3_ob_out[75], \kme_cddip3_ob_out.tstrb [3]);
tran (kme_cddip3_ob_out[74], \kme_cddip3_ob_out.tstrb [2]);
tran (kme_cddip3_ob_out[73], \kme_cddip3_ob_out.tstrb [1]);
tran (kme_cddip3_ob_out[72], \kme_cddip3_ob_out.tstrb [0]);
tran (kme_cddip3_ob_out[71], \kme_cddip3_ob_out.tuser [7]);
tran (kme_cddip3_ob_out[70], \kme_cddip3_ob_out.tuser [6]);
tran (kme_cddip3_ob_out[69], \kme_cddip3_ob_out.tuser [5]);
tran (kme_cddip3_ob_out[68], \kme_cddip3_ob_out.tuser [4]);
tran (kme_cddip3_ob_out[67], \kme_cddip3_ob_out.tuser [3]);
tran (kme_cddip3_ob_out[66], \kme_cddip3_ob_out.tuser [2]);
tran (kme_cddip3_ob_out[65], \kme_cddip3_ob_out.tuser [1]);
tran (kme_cddip3_ob_out[64], \kme_cddip3_ob_out.tuser [0]);
tran (kme_cddip3_ob_out[63], \kme_cddip3_ob_out.tdata [63]);
tran (kme_cddip3_ob_out[62], \kme_cddip3_ob_out.tdata [62]);
tran (kme_cddip3_ob_out[61], \kme_cddip3_ob_out.tdata [61]);
tran (kme_cddip3_ob_out[60], \kme_cddip3_ob_out.tdata [60]);
tran (kme_cddip3_ob_out[59], \kme_cddip3_ob_out.tdata [59]);
tran (kme_cddip3_ob_out[58], \kme_cddip3_ob_out.tdata [58]);
tran (kme_cddip3_ob_out[57], \kme_cddip3_ob_out.tdata [57]);
tran (kme_cddip3_ob_out[56], \kme_cddip3_ob_out.tdata [56]);
tran (kme_cddip3_ob_out[55], \kme_cddip3_ob_out.tdata [55]);
tran (kme_cddip3_ob_out[54], \kme_cddip3_ob_out.tdata [54]);
tran (kme_cddip3_ob_out[53], \kme_cddip3_ob_out.tdata [53]);
tran (kme_cddip3_ob_out[52], \kme_cddip3_ob_out.tdata [52]);
tran (kme_cddip3_ob_out[51], \kme_cddip3_ob_out.tdata [51]);
tran (kme_cddip3_ob_out[50], \kme_cddip3_ob_out.tdata [50]);
tran (kme_cddip3_ob_out[49], \kme_cddip3_ob_out.tdata [49]);
tran (kme_cddip3_ob_out[48], \kme_cddip3_ob_out.tdata [48]);
tran (kme_cddip3_ob_out[47], \kme_cddip3_ob_out.tdata [47]);
tran (kme_cddip3_ob_out[46], \kme_cddip3_ob_out.tdata [46]);
tran (kme_cddip3_ob_out[45], \kme_cddip3_ob_out.tdata [45]);
tran (kme_cddip3_ob_out[44], \kme_cddip3_ob_out.tdata [44]);
tran (kme_cddip3_ob_out[43], \kme_cddip3_ob_out.tdata [43]);
tran (kme_cddip3_ob_out[42], \kme_cddip3_ob_out.tdata [42]);
tran (kme_cddip3_ob_out[41], \kme_cddip3_ob_out.tdata [41]);
tran (kme_cddip3_ob_out[40], \kme_cddip3_ob_out.tdata [40]);
tran (kme_cddip3_ob_out[39], \kme_cddip3_ob_out.tdata [39]);
tran (kme_cddip3_ob_out[38], \kme_cddip3_ob_out.tdata [38]);
tran (kme_cddip3_ob_out[37], \kme_cddip3_ob_out.tdata [37]);
tran (kme_cddip3_ob_out[36], \kme_cddip3_ob_out.tdata [36]);
tran (kme_cddip3_ob_out[35], \kme_cddip3_ob_out.tdata [35]);
tran (kme_cddip3_ob_out[34], \kme_cddip3_ob_out.tdata [34]);
tran (kme_cddip3_ob_out[33], \kme_cddip3_ob_out.tdata [33]);
tran (kme_cddip3_ob_out[32], \kme_cddip3_ob_out.tdata [32]);
tran (kme_cddip3_ob_out[31], \kme_cddip3_ob_out.tdata [31]);
tran (kme_cddip3_ob_out[30], \kme_cddip3_ob_out.tdata [30]);
tran (kme_cddip3_ob_out[29], \kme_cddip3_ob_out.tdata [29]);
tran (kme_cddip3_ob_out[28], \kme_cddip3_ob_out.tdata [28]);
tran (kme_cddip3_ob_out[27], \kme_cddip3_ob_out.tdata [27]);
tran (kme_cddip3_ob_out[26], \kme_cddip3_ob_out.tdata [26]);
tran (kme_cddip3_ob_out[25], \kme_cddip3_ob_out.tdata [25]);
tran (kme_cddip3_ob_out[24], \kme_cddip3_ob_out.tdata [24]);
tran (kme_cddip3_ob_out[23], \kme_cddip3_ob_out.tdata [23]);
tran (kme_cddip3_ob_out[22], \kme_cddip3_ob_out.tdata [22]);
tran (kme_cddip3_ob_out[21], \kme_cddip3_ob_out.tdata [21]);
tran (kme_cddip3_ob_out[20], \kme_cddip3_ob_out.tdata [20]);
tran (kme_cddip3_ob_out[19], \kme_cddip3_ob_out.tdata [19]);
tran (kme_cddip3_ob_out[18], \kme_cddip3_ob_out.tdata [18]);
tran (kme_cddip3_ob_out[17], \kme_cddip3_ob_out.tdata [17]);
tran (kme_cddip3_ob_out[16], \kme_cddip3_ob_out.tdata [16]);
tran (kme_cddip3_ob_out[15], \kme_cddip3_ob_out.tdata [15]);
tran (kme_cddip3_ob_out[14], \kme_cddip3_ob_out.tdata [14]);
tran (kme_cddip3_ob_out[13], \kme_cddip3_ob_out.tdata [13]);
tran (kme_cddip3_ob_out[12], \kme_cddip3_ob_out.tdata [12]);
tran (kme_cddip3_ob_out[11], \kme_cddip3_ob_out.tdata [11]);
tran (kme_cddip3_ob_out[10], \kme_cddip3_ob_out.tdata [10]);
tran (kme_cddip3_ob_out[9], \kme_cddip3_ob_out.tdata [9]);
tran (kme_cddip3_ob_out[8], \kme_cddip3_ob_out.tdata [8]);
tran (kme_cddip3_ob_out[7], \kme_cddip3_ob_out.tdata [7]);
tran (kme_cddip3_ob_out[6], \kme_cddip3_ob_out.tdata [6]);
tran (kme_cddip3_ob_out[5], \kme_cddip3_ob_out.tdata [5]);
tran (kme_cddip3_ob_out[4], \kme_cddip3_ob_out.tdata [4]);
tran (kme_cddip3_ob_out[3], \kme_cddip3_ob_out.tdata [3]);
tran (kme_cddip3_ob_out[2], \kme_cddip3_ob_out.tdata [2]);
tran (kme_cddip3_ob_out[1], \kme_cddip3_ob_out.tdata [1]);
tran (kme_cddip3_ob_out[0], \kme_cddip3_ob_out.tdata [0]);
tran (o_ckv_ia_config[18], \o_ckv_ia_config.r.part0 [18]);
tran (o_ckv_ia_config[18], \o_ckv_ia_config.f.op [3]);
tran (o_ckv_ia_config[17], \o_ckv_ia_config.r.part0 [17]);
tran (o_ckv_ia_config[17], \o_ckv_ia_config.f.op [2]);
tran (o_ckv_ia_config[16], \o_ckv_ia_config.r.part0 [16]);
tran (o_ckv_ia_config[16], \o_ckv_ia_config.f.op [1]);
tran (o_ckv_ia_config[15], \o_ckv_ia_config.r.part0 [15]);
tran (o_ckv_ia_config[15], \o_ckv_ia_config.f.op [0]);
tran (o_ckv_ia_config[14], \o_ckv_ia_config.r.part0 [14]);
tran (o_ckv_ia_config[14], \o_ckv_ia_config.f.addr [14]);
tran (o_ckv_ia_config[13], \o_ckv_ia_config.r.part0 [13]);
tran (o_ckv_ia_config[13], \o_ckv_ia_config.f.addr [13]);
tran (o_ckv_ia_config[12], \o_ckv_ia_config.r.part0 [12]);
tran (o_ckv_ia_config[12], \o_ckv_ia_config.f.addr [12]);
tran (o_ckv_ia_config[11], \o_ckv_ia_config.r.part0 [11]);
tran (o_ckv_ia_config[11], \o_ckv_ia_config.f.addr [11]);
tran (o_ckv_ia_config[10], \o_ckv_ia_config.r.part0 [10]);
tran (o_ckv_ia_config[10], \o_ckv_ia_config.f.addr [10]);
tran (o_ckv_ia_config[9], \o_ckv_ia_config.r.part0 [9]);
tran (o_ckv_ia_config[9], \o_ckv_ia_config.f.addr [9]);
tran (o_ckv_ia_config[8], \o_ckv_ia_config.r.part0 [8]);
tran (o_ckv_ia_config[8], \o_ckv_ia_config.f.addr [8]);
tran (o_ckv_ia_config[7], \o_ckv_ia_config.r.part0 [7]);
tran (o_ckv_ia_config[7], \o_ckv_ia_config.f.addr [7]);
tran (o_ckv_ia_config[6], \o_ckv_ia_config.r.part0 [6]);
tran (o_ckv_ia_config[6], \o_ckv_ia_config.f.addr [6]);
tran (o_ckv_ia_config[5], \o_ckv_ia_config.r.part0 [5]);
tran (o_ckv_ia_config[5], \o_ckv_ia_config.f.addr [5]);
tran (o_ckv_ia_config[4], \o_ckv_ia_config.r.part0 [4]);
tran (o_ckv_ia_config[4], \o_ckv_ia_config.f.addr [4]);
tran (o_ckv_ia_config[3], \o_ckv_ia_config.r.part0 [3]);
tran (o_ckv_ia_config[3], \o_ckv_ia_config.f.addr [3]);
tran (o_ckv_ia_config[2], \o_ckv_ia_config.r.part0 [2]);
tran (o_ckv_ia_config[2], \o_ckv_ia_config.f.addr [2]);
tran (o_ckv_ia_config[1], \o_ckv_ia_config.r.part0 [1]);
tran (o_ckv_ia_config[1], \o_ckv_ia_config.f.addr [1]);
tran (o_ckv_ia_config[0], \o_ckv_ia_config.r.part0 [0]);
tran (o_ckv_ia_config[0], \o_ckv_ia_config.f.addr [0]);
tran (o_kim_ia_config[17], \o_kim_ia_config.r.part0 [17]);
tran (o_kim_ia_config[17], \o_kim_ia_config.f.op [3]);
tran (o_kim_ia_config[16], \o_kim_ia_config.r.part0 [16]);
tran (o_kim_ia_config[16], \o_kim_ia_config.f.op [2]);
tran (o_kim_ia_config[15], \o_kim_ia_config.r.part0 [15]);
tran (o_kim_ia_config[15], \o_kim_ia_config.f.op [1]);
tran (o_kim_ia_config[14], \o_kim_ia_config.r.part0 [14]);
tran (o_kim_ia_config[14], \o_kim_ia_config.f.op [0]);
tran (o_kim_ia_config[13], \o_kim_ia_config.r.part0 [13]);
tran (o_kim_ia_config[13], \o_kim_ia_config.f.addr [13]);
tran (o_kim_ia_config[12], \o_kim_ia_config.r.part0 [12]);
tran (o_kim_ia_config[12], \o_kim_ia_config.f.addr [12]);
tran (o_kim_ia_config[11], \o_kim_ia_config.r.part0 [11]);
tran (o_kim_ia_config[11], \o_kim_ia_config.f.addr [11]);
tran (o_kim_ia_config[10], \o_kim_ia_config.r.part0 [10]);
tran (o_kim_ia_config[10], \o_kim_ia_config.f.addr [10]);
tran (o_kim_ia_config[9], \o_kim_ia_config.r.part0 [9]);
tran (o_kim_ia_config[9], \o_kim_ia_config.f.addr [9]);
tran (o_kim_ia_config[8], \o_kim_ia_config.r.part0 [8]);
tran (o_kim_ia_config[8], \o_kim_ia_config.f.addr [8]);
tran (o_kim_ia_config[7], \o_kim_ia_config.r.part0 [7]);
tran (o_kim_ia_config[7], \o_kim_ia_config.f.addr [7]);
tran (o_kim_ia_config[6], \o_kim_ia_config.r.part0 [6]);
tran (o_kim_ia_config[6], \o_kim_ia_config.f.addr [6]);
tran (o_kim_ia_config[5], \o_kim_ia_config.r.part0 [5]);
tran (o_kim_ia_config[5], \o_kim_ia_config.f.addr [5]);
tran (o_kim_ia_config[4], \o_kim_ia_config.r.part0 [4]);
tran (o_kim_ia_config[4], \o_kim_ia_config.f.addr [4]);
tran (o_kim_ia_config[3], \o_kim_ia_config.r.part0 [3]);
tran (o_kim_ia_config[3], \o_kim_ia_config.f.addr [3]);
tran (o_kim_ia_config[2], \o_kim_ia_config.r.part0 [2]);
tran (o_kim_ia_config[2], \o_kim_ia_config.f.addr [2]);
tran (o_kim_ia_config[1], \o_kim_ia_config.r.part0 [1]);
tran (o_kim_ia_config[1], \o_kim_ia_config.f.addr [1]);
tran (o_kim_ia_config[0], \o_kim_ia_config.r.part0 [0]);
tran (o_kim_ia_config[0], \o_kim_ia_config.f.addr [0]);
tran (cceip0_out_ia_wdata[95], \cceip0_out_ia_wdata.r.part2 [31]);
tran (cceip0_out_ia_wdata[95], \cceip0_out_ia_wdata.f.tdata_hi [31]);
tran (cceip0_out_ia_wdata[94], \cceip0_out_ia_wdata.r.part2 [30]);
tran (cceip0_out_ia_wdata[94], \cceip0_out_ia_wdata.f.tdata_hi [30]);
tran (cceip0_out_ia_wdata[93], \cceip0_out_ia_wdata.r.part2 [29]);
tran (cceip0_out_ia_wdata[93], \cceip0_out_ia_wdata.f.tdata_hi [29]);
tran (cceip0_out_ia_wdata[92], \cceip0_out_ia_wdata.r.part2 [28]);
tran (cceip0_out_ia_wdata[92], \cceip0_out_ia_wdata.f.tdata_hi [28]);
tran (cceip0_out_ia_wdata[91], \cceip0_out_ia_wdata.r.part2 [27]);
tran (cceip0_out_ia_wdata[91], \cceip0_out_ia_wdata.f.tdata_hi [27]);
tran (cceip0_out_ia_wdata[90], \cceip0_out_ia_wdata.r.part2 [26]);
tran (cceip0_out_ia_wdata[90], \cceip0_out_ia_wdata.f.tdata_hi [26]);
tran (cceip0_out_ia_wdata[89], \cceip0_out_ia_wdata.r.part2 [25]);
tran (cceip0_out_ia_wdata[89], \cceip0_out_ia_wdata.f.tdata_hi [25]);
tran (cceip0_out_ia_wdata[88], \cceip0_out_ia_wdata.r.part2 [24]);
tran (cceip0_out_ia_wdata[88], \cceip0_out_ia_wdata.f.tdata_hi [24]);
tran (cceip0_out_ia_wdata[87], \cceip0_out_ia_wdata.r.part2 [23]);
tran (cceip0_out_ia_wdata[87], \cceip0_out_ia_wdata.f.tdata_hi [23]);
tran (cceip0_out_ia_wdata[86], \cceip0_out_ia_wdata.r.part2 [22]);
tran (cceip0_out_ia_wdata[86], \cceip0_out_ia_wdata.f.tdata_hi [22]);
tran (cceip0_out_ia_wdata[85], \cceip0_out_ia_wdata.r.part2 [21]);
tran (cceip0_out_ia_wdata[85], \cceip0_out_ia_wdata.f.tdata_hi [21]);
tran (cceip0_out_ia_wdata[84], \cceip0_out_ia_wdata.r.part2 [20]);
tran (cceip0_out_ia_wdata[84], \cceip0_out_ia_wdata.f.tdata_hi [20]);
tran (cceip0_out_ia_wdata[83], \cceip0_out_ia_wdata.r.part2 [19]);
tran (cceip0_out_ia_wdata[83], \cceip0_out_ia_wdata.f.tdata_hi [19]);
tran (cceip0_out_ia_wdata[82], \cceip0_out_ia_wdata.r.part2 [18]);
tran (cceip0_out_ia_wdata[82], \cceip0_out_ia_wdata.f.tdata_hi [18]);
tran (cceip0_out_ia_wdata[81], \cceip0_out_ia_wdata.r.part2 [17]);
tran (cceip0_out_ia_wdata[81], \cceip0_out_ia_wdata.f.tdata_hi [17]);
tran (cceip0_out_ia_wdata[80], \cceip0_out_ia_wdata.r.part2 [16]);
tran (cceip0_out_ia_wdata[80], \cceip0_out_ia_wdata.f.tdata_hi [16]);
tran (cceip0_out_ia_wdata[79], \cceip0_out_ia_wdata.r.part2 [15]);
tran (cceip0_out_ia_wdata[79], \cceip0_out_ia_wdata.f.tdata_hi [15]);
tran (cceip0_out_ia_wdata[78], \cceip0_out_ia_wdata.r.part2 [14]);
tran (cceip0_out_ia_wdata[78], \cceip0_out_ia_wdata.f.tdata_hi [14]);
tran (cceip0_out_ia_wdata[77], \cceip0_out_ia_wdata.r.part2 [13]);
tran (cceip0_out_ia_wdata[77], \cceip0_out_ia_wdata.f.tdata_hi [13]);
tran (cceip0_out_ia_wdata[76], \cceip0_out_ia_wdata.r.part2 [12]);
tran (cceip0_out_ia_wdata[76], \cceip0_out_ia_wdata.f.tdata_hi [12]);
tran (cceip0_out_ia_wdata[75], \cceip0_out_ia_wdata.r.part2 [11]);
tran (cceip0_out_ia_wdata[75], \cceip0_out_ia_wdata.f.tdata_hi [11]);
tran (cceip0_out_ia_wdata[74], \cceip0_out_ia_wdata.r.part2 [10]);
tran (cceip0_out_ia_wdata[74], \cceip0_out_ia_wdata.f.tdata_hi [10]);
tran (cceip0_out_ia_wdata[73], \cceip0_out_ia_wdata.r.part2 [9]);
tran (cceip0_out_ia_wdata[73], \cceip0_out_ia_wdata.f.tdata_hi [9]);
tran (cceip0_out_ia_wdata[72], \cceip0_out_ia_wdata.r.part2 [8]);
tran (cceip0_out_ia_wdata[72], \cceip0_out_ia_wdata.f.tdata_hi [8]);
tran (cceip0_out_ia_wdata[71], \cceip0_out_ia_wdata.r.part2 [7]);
tran (cceip0_out_ia_wdata[71], \cceip0_out_ia_wdata.f.tdata_hi [7]);
tran (cceip0_out_ia_wdata[70], \cceip0_out_ia_wdata.r.part2 [6]);
tran (cceip0_out_ia_wdata[70], \cceip0_out_ia_wdata.f.tdata_hi [6]);
tran (cceip0_out_ia_wdata[69], \cceip0_out_ia_wdata.r.part2 [5]);
tran (cceip0_out_ia_wdata[69], \cceip0_out_ia_wdata.f.tdata_hi [5]);
tran (cceip0_out_ia_wdata[68], \cceip0_out_ia_wdata.r.part2 [4]);
tran (cceip0_out_ia_wdata[68], \cceip0_out_ia_wdata.f.tdata_hi [4]);
tran (cceip0_out_ia_wdata[67], \cceip0_out_ia_wdata.r.part2 [3]);
tran (cceip0_out_ia_wdata[67], \cceip0_out_ia_wdata.f.tdata_hi [3]);
tran (cceip0_out_ia_wdata[66], \cceip0_out_ia_wdata.r.part2 [2]);
tran (cceip0_out_ia_wdata[66], \cceip0_out_ia_wdata.f.tdata_hi [2]);
tran (cceip0_out_ia_wdata[65], \cceip0_out_ia_wdata.r.part2 [1]);
tran (cceip0_out_ia_wdata[65], \cceip0_out_ia_wdata.f.tdata_hi [1]);
tran (cceip0_out_ia_wdata[64], \cceip0_out_ia_wdata.r.part2 [0]);
tran (cceip0_out_ia_wdata[64], \cceip0_out_ia_wdata.f.tdata_hi [0]);
tran (cceip0_out_ia_wdata[63], \cceip0_out_ia_wdata.r.part1 [31]);
tran (cceip0_out_ia_wdata[63], \cceip0_out_ia_wdata.f.tdata_lo [31]);
tran (cceip0_out_ia_wdata[62], \cceip0_out_ia_wdata.r.part1 [30]);
tran (cceip0_out_ia_wdata[62], \cceip0_out_ia_wdata.f.tdata_lo [30]);
tran (cceip0_out_ia_wdata[61], \cceip0_out_ia_wdata.r.part1 [29]);
tran (cceip0_out_ia_wdata[61], \cceip0_out_ia_wdata.f.tdata_lo [29]);
tran (cceip0_out_ia_wdata[60], \cceip0_out_ia_wdata.r.part1 [28]);
tran (cceip0_out_ia_wdata[60], \cceip0_out_ia_wdata.f.tdata_lo [28]);
tran (cceip0_out_ia_wdata[59], \cceip0_out_ia_wdata.r.part1 [27]);
tran (cceip0_out_ia_wdata[59], \cceip0_out_ia_wdata.f.tdata_lo [27]);
tran (cceip0_out_ia_wdata[58], \cceip0_out_ia_wdata.r.part1 [26]);
tran (cceip0_out_ia_wdata[58], \cceip0_out_ia_wdata.f.tdata_lo [26]);
tran (cceip0_out_ia_wdata[57], \cceip0_out_ia_wdata.r.part1 [25]);
tran (cceip0_out_ia_wdata[57], \cceip0_out_ia_wdata.f.tdata_lo [25]);
tran (cceip0_out_ia_wdata[56], \cceip0_out_ia_wdata.r.part1 [24]);
tran (cceip0_out_ia_wdata[56], \cceip0_out_ia_wdata.f.tdata_lo [24]);
tran (cceip0_out_ia_wdata[55], \cceip0_out_ia_wdata.r.part1 [23]);
tran (cceip0_out_ia_wdata[55], \cceip0_out_ia_wdata.f.tdata_lo [23]);
tran (cceip0_out_ia_wdata[54], \cceip0_out_ia_wdata.r.part1 [22]);
tran (cceip0_out_ia_wdata[54], \cceip0_out_ia_wdata.f.tdata_lo [22]);
tran (cceip0_out_ia_wdata[53], \cceip0_out_ia_wdata.r.part1 [21]);
tran (cceip0_out_ia_wdata[53], \cceip0_out_ia_wdata.f.tdata_lo [21]);
tran (cceip0_out_ia_wdata[52], \cceip0_out_ia_wdata.r.part1 [20]);
tran (cceip0_out_ia_wdata[52], \cceip0_out_ia_wdata.f.tdata_lo [20]);
tran (cceip0_out_ia_wdata[51], \cceip0_out_ia_wdata.r.part1 [19]);
tran (cceip0_out_ia_wdata[51], \cceip0_out_ia_wdata.f.tdata_lo [19]);
tran (cceip0_out_ia_wdata[50], \cceip0_out_ia_wdata.r.part1 [18]);
tran (cceip0_out_ia_wdata[50], \cceip0_out_ia_wdata.f.tdata_lo [18]);
tran (cceip0_out_ia_wdata[49], \cceip0_out_ia_wdata.r.part1 [17]);
tran (cceip0_out_ia_wdata[49], \cceip0_out_ia_wdata.f.tdata_lo [17]);
tran (cceip0_out_ia_wdata[48], \cceip0_out_ia_wdata.r.part1 [16]);
tran (cceip0_out_ia_wdata[48], \cceip0_out_ia_wdata.f.tdata_lo [16]);
tran (cceip0_out_ia_wdata[47], \cceip0_out_ia_wdata.r.part1 [15]);
tran (cceip0_out_ia_wdata[47], \cceip0_out_ia_wdata.f.tdata_lo [15]);
tran (cceip0_out_ia_wdata[46], \cceip0_out_ia_wdata.r.part1 [14]);
tran (cceip0_out_ia_wdata[46], \cceip0_out_ia_wdata.f.tdata_lo [14]);
tran (cceip0_out_ia_wdata[45], \cceip0_out_ia_wdata.r.part1 [13]);
tran (cceip0_out_ia_wdata[45], \cceip0_out_ia_wdata.f.tdata_lo [13]);
tran (cceip0_out_ia_wdata[44], \cceip0_out_ia_wdata.r.part1 [12]);
tran (cceip0_out_ia_wdata[44], \cceip0_out_ia_wdata.f.tdata_lo [12]);
tran (cceip0_out_ia_wdata[43], \cceip0_out_ia_wdata.r.part1 [11]);
tran (cceip0_out_ia_wdata[43], \cceip0_out_ia_wdata.f.tdata_lo [11]);
tran (cceip0_out_ia_wdata[42], \cceip0_out_ia_wdata.r.part1 [10]);
tran (cceip0_out_ia_wdata[42], \cceip0_out_ia_wdata.f.tdata_lo [10]);
tran (cceip0_out_ia_wdata[41], \cceip0_out_ia_wdata.r.part1 [9]);
tran (cceip0_out_ia_wdata[41], \cceip0_out_ia_wdata.f.tdata_lo [9]);
tran (cceip0_out_ia_wdata[40], \cceip0_out_ia_wdata.r.part1 [8]);
tran (cceip0_out_ia_wdata[40], \cceip0_out_ia_wdata.f.tdata_lo [8]);
tran (cceip0_out_ia_wdata[39], \cceip0_out_ia_wdata.r.part1 [7]);
tran (cceip0_out_ia_wdata[39], \cceip0_out_ia_wdata.f.tdata_lo [7]);
tran (cceip0_out_ia_wdata[38], \cceip0_out_ia_wdata.r.part1 [6]);
tran (cceip0_out_ia_wdata[38], \cceip0_out_ia_wdata.f.tdata_lo [6]);
tran (cceip0_out_ia_wdata[37], \cceip0_out_ia_wdata.r.part1 [5]);
tran (cceip0_out_ia_wdata[37], \cceip0_out_ia_wdata.f.tdata_lo [5]);
tran (cceip0_out_ia_wdata[36], \cceip0_out_ia_wdata.r.part1 [4]);
tran (cceip0_out_ia_wdata[36], \cceip0_out_ia_wdata.f.tdata_lo [4]);
tran (cceip0_out_ia_wdata[35], \cceip0_out_ia_wdata.r.part1 [3]);
tran (cceip0_out_ia_wdata[35], \cceip0_out_ia_wdata.f.tdata_lo [3]);
tran (cceip0_out_ia_wdata[34], \cceip0_out_ia_wdata.r.part1 [2]);
tran (cceip0_out_ia_wdata[34], \cceip0_out_ia_wdata.f.tdata_lo [2]);
tran (cceip0_out_ia_wdata[33], \cceip0_out_ia_wdata.r.part1 [1]);
tran (cceip0_out_ia_wdata[33], \cceip0_out_ia_wdata.f.tdata_lo [1]);
tran (cceip0_out_ia_wdata[32], \cceip0_out_ia_wdata.r.part1 [0]);
tran (cceip0_out_ia_wdata[32], \cceip0_out_ia_wdata.f.tdata_lo [0]);
tran (cceip0_out_ia_wdata[31], \cceip0_out_ia_wdata.r.part0 [31]);
tran (cceip0_out_ia_wdata[31], \cceip0_out_ia_wdata.f.eob );
tran (cceip0_out_ia_wdata[30], \cceip0_out_ia_wdata.r.part0 [30]);
tran (cceip0_out_ia_wdata[30], \cceip0_out_ia_wdata.f.bytes_vld [7]);
tran (cceip0_out_ia_wdata[29], \cceip0_out_ia_wdata.r.part0 [29]);
tran (cceip0_out_ia_wdata[29], \cceip0_out_ia_wdata.f.bytes_vld [6]);
tran (cceip0_out_ia_wdata[28], \cceip0_out_ia_wdata.r.part0 [28]);
tran (cceip0_out_ia_wdata[28], \cceip0_out_ia_wdata.f.bytes_vld [5]);
tran (cceip0_out_ia_wdata[27], \cceip0_out_ia_wdata.r.part0 [27]);
tran (cceip0_out_ia_wdata[27], \cceip0_out_ia_wdata.f.bytes_vld [4]);
tran (cceip0_out_ia_wdata[26], \cceip0_out_ia_wdata.r.part0 [26]);
tran (cceip0_out_ia_wdata[26], \cceip0_out_ia_wdata.f.bytes_vld [3]);
tran (cceip0_out_ia_wdata[25], \cceip0_out_ia_wdata.r.part0 [25]);
tran (cceip0_out_ia_wdata[25], \cceip0_out_ia_wdata.f.bytes_vld [2]);
tran (cceip0_out_ia_wdata[24], \cceip0_out_ia_wdata.r.part0 [24]);
tran (cceip0_out_ia_wdata[24], \cceip0_out_ia_wdata.f.bytes_vld [1]);
tran (cceip0_out_ia_wdata[23], \cceip0_out_ia_wdata.r.part0 [23]);
tran (cceip0_out_ia_wdata[23], \cceip0_out_ia_wdata.f.bytes_vld [0]);
tran (cceip0_out_ia_wdata[22], \cceip0_out_ia_wdata.r.part0 [22]);
tran (cceip0_out_ia_wdata[22], \cceip0_out_ia_wdata.f.unused1 [7]);
tran (cceip0_out_ia_wdata[21], \cceip0_out_ia_wdata.r.part0 [21]);
tran (cceip0_out_ia_wdata[21], \cceip0_out_ia_wdata.f.unused1 [6]);
tran (cceip0_out_ia_wdata[20], \cceip0_out_ia_wdata.r.part0 [20]);
tran (cceip0_out_ia_wdata[20], \cceip0_out_ia_wdata.f.unused1 [5]);
tran (cceip0_out_ia_wdata[19], \cceip0_out_ia_wdata.r.part0 [19]);
tran (cceip0_out_ia_wdata[19], \cceip0_out_ia_wdata.f.unused1 [4]);
tran (cceip0_out_ia_wdata[18], \cceip0_out_ia_wdata.r.part0 [18]);
tran (cceip0_out_ia_wdata[18], \cceip0_out_ia_wdata.f.unused1 [3]);
tran (cceip0_out_ia_wdata[17], \cceip0_out_ia_wdata.r.part0 [17]);
tran (cceip0_out_ia_wdata[17], \cceip0_out_ia_wdata.f.unused1 [2]);
tran (cceip0_out_ia_wdata[16], \cceip0_out_ia_wdata.r.part0 [16]);
tran (cceip0_out_ia_wdata[16], \cceip0_out_ia_wdata.f.unused1 [1]);
tran (cceip0_out_ia_wdata[15], \cceip0_out_ia_wdata.r.part0 [15]);
tran (cceip0_out_ia_wdata[15], \cceip0_out_ia_wdata.f.unused1 [0]);
tran (cceip0_out_ia_wdata[14], \cceip0_out_ia_wdata.r.part0 [14]);
tran (cceip0_out_ia_wdata[14], \cceip0_out_ia_wdata.f.tid );
tran (cceip0_out_ia_wdata[13], \cceip0_out_ia_wdata.r.part0 [13]);
tran (cceip0_out_ia_wdata[13], \cceip0_out_ia_wdata.f.tuser [7]);
tran (cceip0_out_ia_wdata[12], \cceip0_out_ia_wdata.r.part0 [12]);
tran (cceip0_out_ia_wdata[12], \cceip0_out_ia_wdata.f.tuser [6]);
tran (cceip0_out_ia_wdata[11], \cceip0_out_ia_wdata.r.part0 [11]);
tran (cceip0_out_ia_wdata[11], \cceip0_out_ia_wdata.f.tuser [5]);
tran (cceip0_out_ia_wdata[10], \cceip0_out_ia_wdata.r.part0 [10]);
tran (cceip0_out_ia_wdata[10], \cceip0_out_ia_wdata.f.tuser [4]);
tran (cceip0_out_ia_wdata[9], \cceip0_out_ia_wdata.r.part0 [9]);
tran (cceip0_out_ia_wdata[9], \cceip0_out_ia_wdata.f.tuser [3]);
tran (cceip0_out_ia_wdata[8], \cceip0_out_ia_wdata.r.part0 [8]);
tran (cceip0_out_ia_wdata[8], \cceip0_out_ia_wdata.f.tuser [2]);
tran (cceip0_out_ia_wdata[7], \cceip0_out_ia_wdata.r.part0 [7]);
tran (cceip0_out_ia_wdata[7], \cceip0_out_ia_wdata.f.tuser [1]);
tran (cceip0_out_ia_wdata[6], \cceip0_out_ia_wdata.r.part0 [6]);
tran (cceip0_out_ia_wdata[6], \cceip0_out_ia_wdata.f.tuser [0]);
tran (cceip0_out_ia_wdata[5], \cceip0_out_ia_wdata.r.part0 [5]);
tran (cceip0_out_ia_wdata[5], \cceip0_out_ia_wdata.f.unused0 [5]);
tran (cceip0_out_ia_wdata[4], \cceip0_out_ia_wdata.r.part0 [4]);
tran (cceip0_out_ia_wdata[4], \cceip0_out_ia_wdata.f.unused0 [4]);
tran (cceip0_out_ia_wdata[3], \cceip0_out_ia_wdata.r.part0 [3]);
tran (cceip0_out_ia_wdata[3], \cceip0_out_ia_wdata.f.unused0 [3]);
tran (cceip0_out_ia_wdata[2], \cceip0_out_ia_wdata.r.part0 [2]);
tran (cceip0_out_ia_wdata[2], \cceip0_out_ia_wdata.f.unused0 [2]);
tran (cceip0_out_ia_wdata[1], \cceip0_out_ia_wdata.r.part0 [1]);
tran (cceip0_out_ia_wdata[1], \cceip0_out_ia_wdata.f.unused0 [1]);
tran (cceip0_out_ia_wdata[0], \cceip0_out_ia_wdata.r.part0 [0]);
tran (cceip0_out_ia_wdata[0], \cceip0_out_ia_wdata.f.unused0 [0]);
tran (tready_override[8], \tready_override.r.part0 [8]);
tran (tready_override[8], \tready_override.f.txc_tready_override );
tran (tready_override[7], \tready_override.r.part0 [7]);
tran (tready_override[7], \tready_override.f.engine_7_tready_override );
tran (tready_override[6], \tready_override.r.part0 [6]);
tran (tready_override[6], \tready_override.f.engine_6_tready_override );
tran (tready_override[5], \tready_override.r.part0 [5]);
tran (tready_override[5], \tready_override.f.engine_5_tready_override );
tran (tready_override[4], \tready_override.r.part0 [4]);
tran (tready_override[4], \tready_override.f.engine_4_tready_override );
tran (tready_override[3], \tready_override.r.part0 [3]);
tran (tready_override[3], \tready_override.f.engine_3_tready_override );
tran (tready_override[2], \tready_override.r.part0 [2]);
tran (tready_override[2], \tready_override.f.engine_2_tready_override );
tran (tready_override[1], \tready_override.r.part0 [1]);
tran (tready_override[1], \tready_override.f.engine_1_tready_override );
tran (tready_override[0], \tready_override.r.part0 [0]);
tran (tready_override[0], \tready_override.f.engine_0_tready_override );
tran (kme_cceip0_ob_out_post[82], \kme_cceip0_ob_out_post.tvalid );
tran (kme_cceip0_ob_out_post[81], \kme_cceip0_ob_out_post.tlast );
tran (kme_cceip0_ob_out_post[80], \kme_cceip0_ob_out_post.tid [0]);
tran (kme_cceip0_ob_out_post[79], \kme_cceip0_ob_out_post.tstrb [7]);
tran (kme_cceip0_ob_out_post[78], \kme_cceip0_ob_out_post.tstrb [6]);
tran (kme_cceip0_ob_out_post[77], \kme_cceip0_ob_out_post.tstrb [5]);
tran (kme_cceip0_ob_out_post[76], \kme_cceip0_ob_out_post.tstrb [4]);
tran (kme_cceip0_ob_out_post[75], \kme_cceip0_ob_out_post.tstrb [3]);
tran (kme_cceip0_ob_out_post[74], \kme_cceip0_ob_out_post.tstrb [2]);
tran (kme_cceip0_ob_out_post[73], \kme_cceip0_ob_out_post.tstrb [1]);
tran (kme_cceip0_ob_out_post[72], \kme_cceip0_ob_out_post.tstrb [0]);
tran (kme_cceip0_ob_out_post[71], \kme_cceip0_ob_out_post.tuser [7]);
tran (kme_cceip0_ob_out_post[70], \kme_cceip0_ob_out_post.tuser [6]);
tran (kme_cceip0_ob_out_post[69], \kme_cceip0_ob_out_post.tuser [5]);
tran (kme_cceip0_ob_out_post[68], \kme_cceip0_ob_out_post.tuser [4]);
tran (kme_cceip0_ob_out_post[67], \kme_cceip0_ob_out_post.tuser [3]);
tran (kme_cceip0_ob_out_post[66], \kme_cceip0_ob_out_post.tuser [2]);
tran (kme_cceip0_ob_out_post[65], \kme_cceip0_ob_out_post.tuser [1]);
tran (kme_cceip0_ob_out_post[64], \kme_cceip0_ob_out_post.tuser [0]);
tran (kme_cceip0_ob_out_post[63], \kme_cceip0_ob_out_post.tdata [63]);
tran (kme_cceip0_ob_out_post[62], \kme_cceip0_ob_out_post.tdata [62]);
tran (kme_cceip0_ob_out_post[61], \kme_cceip0_ob_out_post.tdata [61]);
tran (kme_cceip0_ob_out_post[60], \kme_cceip0_ob_out_post.tdata [60]);
tran (kme_cceip0_ob_out_post[59], \kme_cceip0_ob_out_post.tdata [59]);
tran (kme_cceip0_ob_out_post[58], \kme_cceip0_ob_out_post.tdata [58]);
tran (kme_cceip0_ob_out_post[57], \kme_cceip0_ob_out_post.tdata [57]);
tran (kme_cceip0_ob_out_post[56], \kme_cceip0_ob_out_post.tdata [56]);
tran (kme_cceip0_ob_out_post[55], \kme_cceip0_ob_out_post.tdata [55]);
tran (kme_cceip0_ob_out_post[54], \kme_cceip0_ob_out_post.tdata [54]);
tran (kme_cceip0_ob_out_post[53], \kme_cceip0_ob_out_post.tdata [53]);
tran (kme_cceip0_ob_out_post[52], \kme_cceip0_ob_out_post.tdata [52]);
tran (kme_cceip0_ob_out_post[51], \kme_cceip0_ob_out_post.tdata [51]);
tran (kme_cceip0_ob_out_post[50], \kme_cceip0_ob_out_post.tdata [50]);
tran (kme_cceip0_ob_out_post[49], \kme_cceip0_ob_out_post.tdata [49]);
tran (kme_cceip0_ob_out_post[48], \kme_cceip0_ob_out_post.tdata [48]);
tran (kme_cceip0_ob_out_post[47], \kme_cceip0_ob_out_post.tdata [47]);
tran (kme_cceip0_ob_out_post[46], \kme_cceip0_ob_out_post.tdata [46]);
tran (kme_cceip0_ob_out_post[45], \kme_cceip0_ob_out_post.tdata [45]);
tran (kme_cceip0_ob_out_post[44], \kme_cceip0_ob_out_post.tdata [44]);
tran (kme_cceip0_ob_out_post[43], \kme_cceip0_ob_out_post.tdata [43]);
tran (kme_cceip0_ob_out_post[42], \kme_cceip0_ob_out_post.tdata [42]);
tran (kme_cceip0_ob_out_post[41], \kme_cceip0_ob_out_post.tdata [41]);
tran (kme_cceip0_ob_out_post[40], \kme_cceip0_ob_out_post.tdata [40]);
tran (kme_cceip0_ob_out_post[39], \kme_cceip0_ob_out_post.tdata [39]);
tran (kme_cceip0_ob_out_post[38], \kme_cceip0_ob_out_post.tdata [38]);
tran (kme_cceip0_ob_out_post[37], \kme_cceip0_ob_out_post.tdata [37]);
tran (kme_cceip0_ob_out_post[36], \kme_cceip0_ob_out_post.tdata [36]);
tran (kme_cceip0_ob_out_post[35], \kme_cceip0_ob_out_post.tdata [35]);
tran (kme_cceip0_ob_out_post[34], \kme_cceip0_ob_out_post.tdata [34]);
tran (kme_cceip0_ob_out_post[33], \kme_cceip0_ob_out_post.tdata [33]);
tran (kme_cceip0_ob_out_post[32], \kme_cceip0_ob_out_post.tdata [32]);
tran (kme_cceip0_ob_out_post[31], \kme_cceip0_ob_out_post.tdata [31]);
tran (kme_cceip0_ob_out_post[30], \kme_cceip0_ob_out_post.tdata [30]);
tran (kme_cceip0_ob_out_post[29], \kme_cceip0_ob_out_post.tdata [29]);
tran (kme_cceip0_ob_out_post[28], \kme_cceip0_ob_out_post.tdata [28]);
tran (kme_cceip0_ob_out_post[27], \kme_cceip0_ob_out_post.tdata [27]);
tran (kme_cceip0_ob_out_post[26], \kme_cceip0_ob_out_post.tdata [26]);
tran (kme_cceip0_ob_out_post[25], \kme_cceip0_ob_out_post.tdata [25]);
tran (kme_cceip0_ob_out_post[24], \kme_cceip0_ob_out_post.tdata [24]);
tran (kme_cceip0_ob_out_post[23], \kme_cceip0_ob_out_post.tdata [23]);
tran (kme_cceip0_ob_out_post[22], \kme_cceip0_ob_out_post.tdata [22]);
tran (kme_cceip0_ob_out_post[21], \kme_cceip0_ob_out_post.tdata [21]);
tran (kme_cceip0_ob_out_post[20], \kme_cceip0_ob_out_post.tdata [20]);
tran (kme_cceip0_ob_out_post[19], \kme_cceip0_ob_out_post.tdata [19]);
tran (kme_cceip0_ob_out_post[18], \kme_cceip0_ob_out_post.tdata [18]);
tran (kme_cceip0_ob_out_post[17], \kme_cceip0_ob_out_post.tdata [17]);
tran (kme_cceip0_ob_out_post[16], \kme_cceip0_ob_out_post.tdata [16]);
tran (kme_cceip0_ob_out_post[15], \kme_cceip0_ob_out_post.tdata [15]);
tran (kme_cceip0_ob_out_post[14], \kme_cceip0_ob_out_post.tdata [14]);
tran (kme_cceip0_ob_out_post[13], \kme_cceip0_ob_out_post.tdata [13]);
tran (kme_cceip0_ob_out_post[12], \kme_cceip0_ob_out_post.tdata [12]);
tran (kme_cceip0_ob_out_post[11], \kme_cceip0_ob_out_post.tdata [11]);
tran (kme_cceip0_ob_out_post[10], \kme_cceip0_ob_out_post.tdata [10]);
tran (kme_cceip0_ob_out_post[9], \kme_cceip0_ob_out_post.tdata [9]);
tran (kme_cceip0_ob_out_post[8], \kme_cceip0_ob_out_post.tdata [8]);
tran (kme_cceip0_ob_out_post[7], \kme_cceip0_ob_out_post.tdata [7]);
tran (kme_cceip0_ob_out_post[6], \kme_cceip0_ob_out_post.tdata [6]);
tran (kme_cceip0_ob_out_post[5], \kme_cceip0_ob_out_post.tdata [5]);
tran (kme_cceip0_ob_out_post[4], \kme_cceip0_ob_out_post.tdata [4]);
tran (kme_cceip0_ob_out_post[3], \kme_cceip0_ob_out_post.tdata [3]);
tran (kme_cceip0_ob_out_post[2], \kme_cceip0_ob_out_post.tdata [2]);
tran (kme_cceip0_ob_out_post[1], \kme_cceip0_ob_out_post.tdata [1]);
tran (kme_cceip0_ob_out_post[0], \kme_cceip0_ob_out_post.tdata [0]);
tran (kme_cceip1_ob_out_post[82], \kme_cceip1_ob_out_post.tvalid );
tran (kme_cceip1_ob_out_post[81], \kme_cceip1_ob_out_post.tlast );
tran (kme_cceip1_ob_out_post[80], \kme_cceip1_ob_out_post.tid [0]);
tran (kme_cceip1_ob_out_post[79], \kme_cceip1_ob_out_post.tstrb [7]);
tran (kme_cceip1_ob_out_post[78], \kme_cceip1_ob_out_post.tstrb [6]);
tran (kme_cceip1_ob_out_post[77], \kme_cceip1_ob_out_post.tstrb [5]);
tran (kme_cceip1_ob_out_post[76], \kme_cceip1_ob_out_post.tstrb [4]);
tran (kme_cceip1_ob_out_post[75], \kme_cceip1_ob_out_post.tstrb [3]);
tran (kme_cceip1_ob_out_post[74], \kme_cceip1_ob_out_post.tstrb [2]);
tran (kme_cceip1_ob_out_post[73], \kme_cceip1_ob_out_post.tstrb [1]);
tran (kme_cceip1_ob_out_post[72], \kme_cceip1_ob_out_post.tstrb [0]);
tran (kme_cceip1_ob_out_post[71], \kme_cceip1_ob_out_post.tuser [7]);
tran (kme_cceip1_ob_out_post[70], \kme_cceip1_ob_out_post.tuser [6]);
tran (kme_cceip1_ob_out_post[69], \kme_cceip1_ob_out_post.tuser [5]);
tran (kme_cceip1_ob_out_post[68], \kme_cceip1_ob_out_post.tuser [4]);
tran (kme_cceip1_ob_out_post[67], \kme_cceip1_ob_out_post.tuser [3]);
tran (kme_cceip1_ob_out_post[66], \kme_cceip1_ob_out_post.tuser [2]);
tran (kme_cceip1_ob_out_post[65], \kme_cceip1_ob_out_post.tuser [1]);
tran (kme_cceip1_ob_out_post[64], \kme_cceip1_ob_out_post.tuser [0]);
tran (kme_cceip1_ob_out_post[63], \kme_cceip1_ob_out_post.tdata [63]);
tran (kme_cceip1_ob_out_post[62], \kme_cceip1_ob_out_post.tdata [62]);
tran (kme_cceip1_ob_out_post[61], \kme_cceip1_ob_out_post.tdata [61]);
tran (kme_cceip1_ob_out_post[60], \kme_cceip1_ob_out_post.tdata [60]);
tran (kme_cceip1_ob_out_post[59], \kme_cceip1_ob_out_post.tdata [59]);
tran (kme_cceip1_ob_out_post[58], \kme_cceip1_ob_out_post.tdata [58]);
tran (kme_cceip1_ob_out_post[57], \kme_cceip1_ob_out_post.tdata [57]);
tran (kme_cceip1_ob_out_post[56], \kme_cceip1_ob_out_post.tdata [56]);
tran (kme_cceip1_ob_out_post[55], \kme_cceip1_ob_out_post.tdata [55]);
tran (kme_cceip1_ob_out_post[54], \kme_cceip1_ob_out_post.tdata [54]);
tran (kme_cceip1_ob_out_post[53], \kme_cceip1_ob_out_post.tdata [53]);
tran (kme_cceip1_ob_out_post[52], \kme_cceip1_ob_out_post.tdata [52]);
tran (kme_cceip1_ob_out_post[51], \kme_cceip1_ob_out_post.tdata [51]);
tran (kme_cceip1_ob_out_post[50], \kme_cceip1_ob_out_post.tdata [50]);
tran (kme_cceip1_ob_out_post[49], \kme_cceip1_ob_out_post.tdata [49]);
tran (kme_cceip1_ob_out_post[48], \kme_cceip1_ob_out_post.tdata [48]);
tran (kme_cceip1_ob_out_post[47], \kme_cceip1_ob_out_post.tdata [47]);
tran (kme_cceip1_ob_out_post[46], \kme_cceip1_ob_out_post.tdata [46]);
tran (kme_cceip1_ob_out_post[45], \kme_cceip1_ob_out_post.tdata [45]);
tran (kme_cceip1_ob_out_post[44], \kme_cceip1_ob_out_post.tdata [44]);
tran (kme_cceip1_ob_out_post[43], \kme_cceip1_ob_out_post.tdata [43]);
tran (kme_cceip1_ob_out_post[42], \kme_cceip1_ob_out_post.tdata [42]);
tran (kme_cceip1_ob_out_post[41], \kme_cceip1_ob_out_post.tdata [41]);
tran (kme_cceip1_ob_out_post[40], \kme_cceip1_ob_out_post.tdata [40]);
tran (kme_cceip1_ob_out_post[39], \kme_cceip1_ob_out_post.tdata [39]);
tran (kme_cceip1_ob_out_post[38], \kme_cceip1_ob_out_post.tdata [38]);
tran (kme_cceip1_ob_out_post[37], \kme_cceip1_ob_out_post.tdata [37]);
tran (kme_cceip1_ob_out_post[36], \kme_cceip1_ob_out_post.tdata [36]);
tran (kme_cceip1_ob_out_post[35], \kme_cceip1_ob_out_post.tdata [35]);
tran (kme_cceip1_ob_out_post[34], \kme_cceip1_ob_out_post.tdata [34]);
tran (kme_cceip1_ob_out_post[33], \kme_cceip1_ob_out_post.tdata [33]);
tran (kme_cceip1_ob_out_post[32], \kme_cceip1_ob_out_post.tdata [32]);
tran (kme_cceip1_ob_out_post[31], \kme_cceip1_ob_out_post.tdata [31]);
tran (kme_cceip1_ob_out_post[30], \kme_cceip1_ob_out_post.tdata [30]);
tran (kme_cceip1_ob_out_post[29], \kme_cceip1_ob_out_post.tdata [29]);
tran (kme_cceip1_ob_out_post[28], \kme_cceip1_ob_out_post.tdata [28]);
tran (kme_cceip1_ob_out_post[27], \kme_cceip1_ob_out_post.tdata [27]);
tran (kme_cceip1_ob_out_post[26], \kme_cceip1_ob_out_post.tdata [26]);
tran (kme_cceip1_ob_out_post[25], \kme_cceip1_ob_out_post.tdata [25]);
tran (kme_cceip1_ob_out_post[24], \kme_cceip1_ob_out_post.tdata [24]);
tran (kme_cceip1_ob_out_post[23], \kme_cceip1_ob_out_post.tdata [23]);
tran (kme_cceip1_ob_out_post[22], \kme_cceip1_ob_out_post.tdata [22]);
tran (kme_cceip1_ob_out_post[21], \kme_cceip1_ob_out_post.tdata [21]);
tran (kme_cceip1_ob_out_post[20], \kme_cceip1_ob_out_post.tdata [20]);
tran (kme_cceip1_ob_out_post[19], \kme_cceip1_ob_out_post.tdata [19]);
tran (kme_cceip1_ob_out_post[18], \kme_cceip1_ob_out_post.tdata [18]);
tran (kme_cceip1_ob_out_post[17], \kme_cceip1_ob_out_post.tdata [17]);
tran (kme_cceip1_ob_out_post[16], \kme_cceip1_ob_out_post.tdata [16]);
tran (kme_cceip1_ob_out_post[15], \kme_cceip1_ob_out_post.tdata [15]);
tran (kme_cceip1_ob_out_post[14], \kme_cceip1_ob_out_post.tdata [14]);
tran (kme_cceip1_ob_out_post[13], \kme_cceip1_ob_out_post.tdata [13]);
tran (kme_cceip1_ob_out_post[12], \kme_cceip1_ob_out_post.tdata [12]);
tran (kme_cceip1_ob_out_post[11], \kme_cceip1_ob_out_post.tdata [11]);
tran (kme_cceip1_ob_out_post[10], \kme_cceip1_ob_out_post.tdata [10]);
tran (kme_cceip1_ob_out_post[9], \kme_cceip1_ob_out_post.tdata [9]);
tran (kme_cceip1_ob_out_post[8], \kme_cceip1_ob_out_post.tdata [8]);
tran (kme_cceip1_ob_out_post[7], \kme_cceip1_ob_out_post.tdata [7]);
tran (kme_cceip1_ob_out_post[6], \kme_cceip1_ob_out_post.tdata [6]);
tran (kme_cceip1_ob_out_post[5], \kme_cceip1_ob_out_post.tdata [5]);
tran (kme_cceip1_ob_out_post[4], \kme_cceip1_ob_out_post.tdata [4]);
tran (kme_cceip1_ob_out_post[3], \kme_cceip1_ob_out_post.tdata [3]);
tran (kme_cceip1_ob_out_post[2], \kme_cceip1_ob_out_post.tdata [2]);
tran (kme_cceip1_ob_out_post[1], \kme_cceip1_ob_out_post.tdata [1]);
tran (kme_cceip1_ob_out_post[0], \kme_cceip1_ob_out_post.tdata [0]);
tran (kme_cceip2_ob_out_post[82], \kme_cceip2_ob_out_post.tvalid );
tran (kme_cceip2_ob_out_post[81], \kme_cceip2_ob_out_post.tlast );
tran (kme_cceip2_ob_out_post[80], \kme_cceip2_ob_out_post.tid [0]);
tran (kme_cceip2_ob_out_post[79], \kme_cceip2_ob_out_post.tstrb [7]);
tran (kme_cceip2_ob_out_post[78], \kme_cceip2_ob_out_post.tstrb [6]);
tran (kme_cceip2_ob_out_post[77], \kme_cceip2_ob_out_post.tstrb [5]);
tran (kme_cceip2_ob_out_post[76], \kme_cceip2_ob_out_post.tstrb [4]);
tran (kme_cceip2_ob_out_post[75], \kme_cceip2_ob_out_post.tstrb [3]);
tran (kme_cceip2_ob_out_post[74], \kme_cceip2_ob_out_post.tstrb [2]);
tran (kme_cceip2_ob_out_post[73], \kme_cceip2_ob_out_post.tstrb [1]);
tran (kme_cceip2_ob_out_post[72], \kme_cceip2_ob_out_post.tstrb [0]);
tran (kme_cceip2_ob_out_post[71], \kme_cceip2_ob_out_post.tuser [7]);
tran (kme_cceip2_ob_out_post[70], \kme_cceip2_ob_out_post.tuser [6]);
tran (kme_cceip2_ob_out_post[69], \kme_cceip2_ob_out_post.tuser [5]);
tran (kme_cceip2_ob_out_post[68], \kme_cceip2_ob_out_post.tuser [4]);
tran (kme_cceip2_ob_out_post[67], \kme_cceip2_ob_out_post.tuser [3]);
tran (kme_cceip2_ob_out_post[66], \kme_cceip2_ob_out_post.tuser [2]);
tran (kme_cceip2_ob_out_post[65], \kme_cceip2_ob_out_post.tuser [1]);
tran (kme_cceip2_ob_out_post[64], \kme_cceip2_ob_out_post.tuser [0]);
tran (kme_cceip2_ob_out_post[63], \kme_cceip2_ob_out_post.tdata [63]);
tran (kme_cceip2_ob_out_post[62], \kme_cceip2_ob_out_post.tdata [62]);
tran (kme_cceip2_ob_out_post[61], \kme_cceip2_ob_out_post.tdata [61]);
tran (kme_cceip2_ob_out_post[60], \kme_cceip2_ob_out_post.tdata [60]);
tran (kme_cceip2_ob_out_post[59], \kme_cceip2_ob_out_post.tdata [59]);
tran (kme_cceip2_ob_out_post[58], \kme_cceip2_ob_out_post.tdata [58]);
tran (kme_cceip2_ob_out_post[57], \kme_cceip2_ob_out_post.tdata [57]);
tran (kme_cceip2_ob_out_post[56], \kme_cceip2_ob_out_post.tdata [56]);
tran (kme_cceip2_ob_out_post[55], \kme_cceip2_ob_out_post.tdata [55]);
tran (kme_cceip2_ob_out_post[54], \kme_cceip2_ob_out_post.tdata [54]);
tran (kme_cceip2_ob_out_post[53], \kme_cceip2_ob_out_post.tdata [53]);
tran (kme_cceip2_ob_out_post[52], \kme_cceip2_ob_out_post.tdata [52]);
tran (kme_cceip2_ob_out_post[51], \kme_cceip2_ob_out_post.tdata [51]);
tran (kme_cceip2_ob_out_post[50], \kme_cceip2_ob_out_post.tdata [50]);
tran (kme_cceip2_ob_out_post[49], \kme_cceip2_ob_out_post.tdata [49]);
tran (kme_cceip2_ob_out_post[48], \kme_cceip2_ob_out_post.tdata [48]);
tran (kme_cceip2_ob_out_post[47], \kme_cceip2_ob_out_post.tdata [47]);
tran (kme_cceip2_ob_out_post[46], \kme_cceip2_ob_out_post.tdata [46]);
tran (kme_cceip2_ob_out_post[45], \kme_cceip2_ob_out_post.tdata [45]);
tran (kme_cceip2_ob_out_post[44], \kme_cceip2_ob_out_post.tdata [44]);
tran (kme_cceip2_ob_out_post[43], \kme_cceip2_ob_out_post.tdata [43]);
tran (kme_cceip2_ob_out_post[42], \kme_cceip2_ob_out_post.tdata [42]);
tran (kme_cceip2_ob_out_post[41], \kme_cceip2_ob_out_post.tdata [41]);
tran (kme_cceip2_ob_out_post[40], \kme_cceip2_ob_out_post.tdata [40]);
tran (kme_cceip2_ob_out_post[39], \kme_cceip2_ob_out_post.tdata [39]);
tran (kme_cceip2_ob_out_post[38], \kme_cceip2_ob_out_post.tdata [38]);
tran (kme_cceip2_ob_out_post[37], \kme_cceip2_ob_out_post.tdata [37]);
tran (kme_cceip2_ob_out_post[36], \kme_cceip2_ob_out_post.tdata [36]);
tran (kme_cceip2_ob_out_post[35], \kme_cceip2_ob_out_post.tdata [35]);
tran (kme_cceip2_ob_out_post[34], \kme_cceip2_ob_out_post.tdata [34]);
tran (kme_cceip2_ob_out_post[33], \kme_cceip2_ob_out_post.tdata [33]);
tran (kme_cceip2_ob_out_post[32], \kme_cceip2_ob_out_post.tdata [32]);
tran (kme_cceip2_ob_out_post[31], \kme_cceip2_ob_out_post.tdata [31]);
tran (kme_cceip2_ob_out_post[30], \kme_cceip2_ob_out_post.tdata [30]);
tran (kme_cceip2_ob_out_post[29], \kme_cceip2_ob_out_post.tdata [29]);
tran (kme_cceip2_ob_out_post[28], \kme_cceip2_ob_out_post.tdata [28]);
tran (kme_cceip2_ob_out_post[27], \kme_cceip2_ob_out_post.tdata [27]);
tran (kme_cceip2_ob_out_post[26], \kme_cceip2_ob_out_post.tdata [26]);
tran (kme_cceip2_ob_out_post[25], \kme_cceip2_ob_out_post.tdata [25]);
tran (kme_cceip2_ob_out_post[24], \kme_cceip2_ob_out_post.tdata [24]);
tran (kme_cceip2_ob_out_post[23], \kme_cceip2_ob_out_post.tdata [23]);
tran (kme_cceip2_ob_out_post[22], \kme_cceip2_ob_out_post.tdata [22]);
tran (kme_cceip2_ob_out_post[21], \kme_cceip2_ob_out_post.tdata [21]);
tran (kme_cceip2_ob_out_post[20], \kme_cceip2_ob_out_post.tdata [20]);
tran (kme_cceip2_ob_out_post[19], \kme_cceip2_ob_out_post.tdata [19]);
tran (kme_cceip2_ob_out_post[18], \kme_cceip2_ob_out_post.tdata [18]);
tran (kme_cceip2_ob_out_post[17], \kme_cceip2_ob_out_post.tdata [17]);
tran (kme_cceip2_ob_out_post[16], \kme_cceip2_ob_out_post.tdata [16]);
tran (kme_cceip2_ob_out_post[15], \kme_cceip2_ob_out_post.tdata [15]);
tran (kme_cceip2_ob_out_post[14], \kme_cceip2_ob_out_post.tdata [14]);
tran (kme_cceip2_ob_out_post[13], \kme_cceip2_ob_out_post.tdata [13]);
tran (kme_cceip2_ob_out_post[12], \kme_cceip2_ob_out_post.tdata [12]);
tran (kme_cceip2_ob_out_post[11], \kme_cceip2_ob_out_post.tdata [11]);
tran (kme_cceip2_ob_out_post[10], \kme_cceip2_ob_out_post.tdata [10]);
tran (kme_cceip2_ob_out_post[9], \kme_cceip2_ob_out_post.tdata [9]);
tran (kme_cceip2_ob_out_post[8], \kme_cceip2_ob_out_post.tdata [8]);
tran (kme_cceip2_ob_out_post[7], \kme_cceip2_ob_out_post.tdata [7]);
tran (kme_cceip2_ob_out_post[6], \kme_cceip2_ob_out_post.tdata [6]);
tran (kme_cceip2_ob_out_post[5], \kme_cceip2_ob_out_post.tdata [5]);
tran (kme_cceip2_ob_out_post[4], \kme_cceip2_ob_out_post.tdata [4]);
tran (kme_cceip2_ob_out_post[3], \kme_cceip2_ob_out_post.tdata [3]);
tran (kme_cceip2_ob_out_post[2], \kme_cceip2_ob_out_post.tdata [2]);
tran (kme_cceip2_ob_out_post[1], \kme_cceip2_ob_out_post.tdata [1]);
tran (kme_cceip2_ob_out_post[0], \kme_cceip2_ob_out_post.tdata [0]);
tran (kme_cceip3_ob_out_post[82], \kme_cceip3_ob_out_post.tvalid );
tran (kme_cceip3_ob_out_post[81], \kme_cceip3_ob_out_post.tlast );
tran (kme_cceip3_ob_out_post[80], \kme_cceip3_ob_out_post.tid [0]);
tran (kme_cceip3_ob_out_post[79], \kme_cceip3_ob_out_post.tstrb [7]);
tran (kme_cceip3_ob_out_post[78], \kme_cceip3_ob_out_post.tstrb [6]);
tran (kme_cceip3_ob_out_post[77], \kme_cceip3_ob_out_post.tstrb [5]);
tran (kme_cceip3_ob_out_post[76], \kme_cceip3_ob_out_post.tstrb [4]);
tran (kme_cceip3_ob_out_post[75], \kme_cceip3_ob_out_post.tstrb [3]);
tran (kme_cceip3_ob_out_post[74], \kme_cceip3_ob_out_post.tstrb [2]);
tran (kme_cceip3_ob_out_post[73], \kme_cceip3_ob_out_post.tstrb [1]);
tran (kme_cceip3_ob_out_post[72], \kme_cceip3_ob_out_post.tstrb [0]);
tran (kme_cceip3_ob_out_post[71], \kme_cceip3_ob_out_post.tuser [7]);
tran (kme_cceip3_ob_out_post[70], \kme_cceip3_ob_out_post.tuser [6]);
tran (kme_cceip3_ob_out_post[69], \kme_cceip3_ob_out_post.tuser [5]);
tran (kme_cceip3_ob_out_post[68], \kme_cceip3_ob_out_post.tuser [4]);
tran (kme_cceip3_ob_out_post[67], \kme_cceip3_ob_out_post.tuser [3]);
tran (kme_cceip3_ob_out_post[66], \kme_cceip3_ob_out_post.tuser [2]);
tran (kme_cceip3_ob_out_post[65], \kme_cceip3_ob_out_post.tuser [1]);
tran (kme_cceip3_ob_out_post[64], \kme_cceip3_ob_out_post.tuser [0]);
tran (kme_cceip3_ob_out_post[63], \kme_cceip3_ob_out_post.tdata [63]);
tran (kme_cceip3_ob_out_post[62], \kme_cceip3_ob_out_post.tdata [62]);
tran (kme_cceip3_ob_out_post[61], \kme_cceip3_ob_out_post.tdata [61]);
tran (kme_cceip3_ob_out_post[60], \kme_cceip3_ob_out_post.tdata [60]);
tran (kme_cceip3_ob_out_post[59], \kme_cceip3_ob_out_post.tdata [59]);
tran (kme_cceip3_ob_out_post[58], \kme_cceip3_ob_out_post.tdata [58]);
tran (kme_cceip3_ob_out_post[57], \kme_cceip3_ob_out_post.tdata [57]);
tran (kme_cceip3_ob_out_post[56], \kme_cceip3_ob_out_post.tdata [56]);
tran (kme_cceip3_ob_out_post[55], \kme_cceip3_ob_out_post.tdata [55]);
tran (kme_cceip3_ob_out_post[54], \kme_cceip3_ob_out_post.tdata [54]);
tran (kme_cceip3_ob_out_post[53], \kme_cceip3_ob_out_post.tdata [53]);
tran (kme_cceip3_ob_out_post[52], \kme_cceip3_ob_out_post.tdata [52]);
tran (kme_cceip3_ob_out_post[51], \kme_cceip3_ob_out_post.tdata [51]);
tran (kme_cceip3_ob_out_post[50], \kme_cceip3_ob_out_post.tdata [50]);
tran (kme_cceip3_ob_out_post[49], \kme_cceip3_ob_out_post.tdata [49]);
tran (kme_cceip3_ob_out_post[48], \kme_cceip3_ob_out_post.tdata [48]);
tran (kme_cceip3_ob_out_post[47], \kme_cceip3_ob_out_post.tdata [47]);
tran (kme_cceip3_ob_out_post[46], \kme_cceip3_ob_out_post.tdata [46]);
tran (kme_cceip3_ob_out_post[45], \kme_cceip3_ob_out_post.tdata [45]);
tran (kme_cceip3_ob_out_post[44], \kme_cceip3_ob_out_post.tdata [44]);
tran (kme_cceip3_ob_out_post[43], \kme_cceip3_ob_out_post.tdata [43]);
tran (kme_cceip3_ob_out_post[42], \kme_cceip3_ob_out_post.tdata [42]);
tran (kme_cceip3_ob_out_post[41], \kme_cceip3_ob_out_post.tdata [41]);
tran (kme_cceip3_ob_out_post[40], \kme_cceip3_ob_out_post.tdata [40]);
tran (kme_cceip3_ob_out_post[39], \kme_cceip3_ob_out_post.tdata [39]);
tran (kme_cceip3_ob_out_post[38], \kme_cceip3_ob_out_post.tdata [38]);
tran (kme_cceip3_ob_out_post[37], \kme_cceip3_ob_out_post.tdata [37]);
tran (kme_cceip3_ob_out_post[36], \kme_cceip3_ob_out_post.tdata [36]);
tran (kme_cceip3_ob_out_post[35], \kme_cceip3_ob_out_post.tdata [35]);
tran (kme_cceip3_ob_out_post[34], \kme_cceip3_ob_out_post.tdata [34]);
tran (kme_cceip3_ob_out_post[33], \kme_cceip3_ob_out_post.tdata [33]);
tran (kme_cceip3_ob_out_post[32], \kme_cceip3_ob_out_post.tdata [32]);
tran (kme_cceip3_ob_out_post[31], \kme_cceip3_ob_out_post.tdata [31]);
tran (kme_cceip3_ob_out_post[30], \kme_cceip3_ob_out_post.tdata [30]);
tran (kme_cceip3_ob_out_post[29], \kme_cceip3_ob_out_post.tdata [29]);
tran (kme_cceip3_ob_out_post[28], \kme_cceip3_ob_out_post.tdata [28]);
tran (kme_cceip3_ob_out_post[27], \kme_cceip3_ob_out_post.tdata [27]);
tran (kme_cceip3_ob_out_post[26], \kme_cceip3_ob_out_post.tdata [26]);
tran (kme_cceip3_ob_out_post[25], \kme_cceip3_ob_out_post.tdata [25]);
tran (kme_cceip3_ob_out_post[24], \kme_cceip3_ob_out_post.tdata [24]);
tran (kme_cceip3_ob_out_post[23], \kme_cceip3_ob_out_post.tdata [23]);
tran (kme_cceip3_ob_out_post[22], \kme_cceip3_ob_out_post.tdata [22]);
tran (kme_cceip3_ob_out_post[21], \kme_cceip3_ob_out_post.tdata [21]);
tran (kme_cceip3_ob_out_post[20], \kme_cceip3_ob_out_post.tdata [20]);
tran (kme_cceip3_ob_out_post[19], \kme_cceip3_ob_out_post.tdata [19]);
tran (kme_cceip3_ob_out_post[18], \kme_cceip3_ob_out_post.tdata [18]);
tran (kme_cceip3_ob_out_post[17], \kme_cceip3_ob_out_post.tdata [17]);
tran (kme_cceip3_ob_out_post[16], \kme_cceip3_ob_out_post.tdata [16]);
tran (kme_cceip3_ob_out_post[15], \kme_cceip3_ob_out_post.tdata [15]);
tran (kme_cceip3_ob_out_post[14], \kme_cceip3_ob_out_post.tdata [14]);
tran (kme_cceip3_ob_out_post[13], \kme_cceip3_ob_out_post.tdata [13]);
tran (kme_cceip3_ob_out_post[12], \kme_cceip3_ob_out_post.tdata [12]);
tran (kme_cceip3_ob_out_post[11], \kme_cceip3_ob_out_post.tdata [11]);
tran (kme_cceip3_ob_out_post[10], \kme_cceip3_ob_out_post.tdata [10]);
tran (kme_cceip3_ob_out_post[9], \kme_cceip3_ob_out_post.tdata [9]);
tran (kme_cceip3_ob_out_post[8], \kme_cceip3_ob_out_post.tdata [8]);
tran (kme_cceip3_ob_out_post[7], \kme_cceip3_ob_out_post.tdata [7]);
tran (kme_cceip3_ob_out_post[6], \kme_cceip3_ob_out_post.tdata [6]);
tran (kme_cceip3_ob_out_post[5], \kme_cceip3_ob_out_post.tdata [5]);
tran (kme_cceip3_ob_out_post[4], \kme_cceip3_ob_out_post.tdata [4]);
tran (kme_cceip3_ob_out_post[3], \kme_cceip3_ob_out_post.tdata [3]);
tran (kme_cceip3_ob_out_post[2], \kme_cceip3_ob_out_post.tdata [2]);
tran (kme_cceip3_ob_out_post[1], \kme_cceip3_ob_out_post.tdata [1]);
tran (kme_cceip3_ob_out_post[0], \kme_cceip3_ob_out_post.tdata [0]);
tran (kme_cddip0_ob_out_post[82], \kme_cddip0_ob_out_post.tvalid );
tran (kme_cddip0_ob_out_post[81], \kme_cddip0_ob_out_post.tlast );
tran (kme_cddip0_ob_out_post[80], \kme_cddip0_ob_out_post.tid [0]);
tran (kme_cddip0_ob_out_post[79], \kme_cddip0_ob_out_post.tstrb [7]);
tran (kme_cddip0_ob_out_post[78], \kme_cddip0_ob_out_post.tstrb [6]);
tran (kme_cddip0_ob_out_post[77], \kme_cddip0_ob_out_post.tstrb [5]);
tran (kme_cddip0_ob_out_post[76], \kme_cddip0_ob_out_post.tstrb [4]);
tran (kme_cddip0_ob_out_post[75], \kme_cddip0_ob_out_post.tstrb [3]);
tran (kme_cddip0_ob_out_post[74], \kme_cddip0_ob_out_post.tstrb [2]);
tran (kme_cddip0_ob_out_post[73], \kme_cddip0_ob_out_post.tstrb [1]);
tran (kme_cddip0_ob_out_post[72], \kme_cddip0_ob_out_post.tstrb [0]);
tran (kme_cddip0_ob_out_post[71], \kme_cddip0_ob_out_post.tuser [7]);
tran (kme_cddip0_ob_out_post[70], \kme_cddip0_ob_out_post.tuser [6]);
tran (kme_cddip0_ob_out_post[69], \kme_cddip0_ob_out_post.tuser [5]);
tran (kme_cddip0_ob_out_post[68], \kme_cddip0_ob_out_post.tuser [4]);
tran (kme_cddip0_ob_out_post[67], \kme_cddip0_ob_out_post.tuser [3]);
tran (kme_cddip0_ob_out_post[66], \kme_cddip0_ob_out_post.tuser [2]);
tran (kme_cddip0_ob_out_post[65], \kme_cddip0_ob_out_post.tuser [1]);
tran (kme_cddip0_ob_out_post[64], \kme_cddip0_ob_out_post.tuser [0]);
tran (kme_cddip0_ob_out_post[63], \kme_cddip0_ob_out_post.tdata [63]);
tran (kme_cddip0_ob_out_post[62], \kme_cddip0_ob_out_post.tdata [62]);
tran (kme_cddip0_ob_out_post[61], \kme_cddip0_ob_out_post.tdata [61]);
tran (kme_cddip0_ob_out_post[60], \kme_cddip0_ob_out_post.tdata [60]);
tran (kme_cddip0_ob_out_post[59], \kme_cddip0_ob_out_post.tdata [59]);
tran (kme_cddip0_ob_out_post[58], \kme_cddip0_ob_out_post.tdata [58]);
tran (kme_cddip0_ob_out_post[57], \kme_cddip0_ob_out_post.tdata [57]);
tran (kme_cddip0_ob_out_post[56], \kme_cddip0_ob_out_post.tdata [56]);
tran (kme_cddip0_ob_out_post[55], \kme_cddip0_ob_out_post.tdata [55]);
tran (kme_cddip0_ob_out_post[54], \kme_cddip0_ob_out_post.tdata [54]);
tran (kme_cddip0_ob_out_post[53], \kme_cddip0_ob_out_post.tdata [53]);
tran (kme_cddip0_ob_out_post[52], \kme_cddip0_ob_out_post.tdata [52]);
tran (kme_cddip0_ob_out_post[51], \kme_cddip0_ob_out_post.tdata [51]);
tran (kme_cddip0_ob_out_post[50], \kme_cddip0_ob_out_post.tdata [50]);
tran (kme_cddip0_ob_out_post[49], \kme_cddip0_ob_out_post.tdata [49]);
tran (kme_cddip0_ob_out_post[48], \kme_cddip0_ob_out_post.tdata [48]);
tran (kme_cddip0_ob_out_post[47], \kme_cddip0_ob_out_post.tdata [47]);
tran (kme_cddip0_ob_out_post[46], \kme_cddip0_ob_out_post.tdata [46]);
tran (kme_cddip0_ob_out_post[45], \kme_cddip0_ob_out_post.tdata [45]);
tran (kme_cddip0_ob_out_post[44], \kme_cddip0_ob_out_post.tdata [44]);
tran (kme_cddip0_ob_out_post[43], \kme_cddip0_ob_out_post.tdata [43]);
tran (kme_cddip0_ob_out_post[42], \kme_cddip0_ob_out_post.tdata [42]);
tran (kme_cddip0_ob_out_post[41], \kme_cddip0_ob_out_post.tdata [41]);
tran (kme_cddip0_ob_out_post[40], \kme_cddip0_ob_out_post.tdata [40]);
tran (kme_cddip0_ob_out_post[39], \kme_cddip0_ob_out_post.tdata [39]);
tran (kme_cddip0_ob_out_post[38], \kme_cddip0_ob_out_post.tdata [38]);
tran (kme_cddip0_ob_out_post[37], \kme_cddip0_ob_out_post.tdata [37]);
tran (kme_cddip0_ob_out_post[36], \kme_cddip0_ob_out_post.tdata [36]);
tran (kme_cddip0_ob_out_post[35], \kme_cddip0_ob_out_post.tdata [35]);
tran (kme_cddip0_ob_out_post[34], \kme_cddip0_ob_out_post.tdata [34]);
tran (kme_cddip0_ob_out_post[33], \kme_cddip0_ob_out_post.tdata [33]);
tran (kme_cddip0_ob_out_post[32], \kme_cddip0_ob_out_post.tdata [32]);
tran (kme_cddip0_ob_out_post[31], \kme_cddip0_ob_out_post.tdata [31]);
tran (kme_cddip0_ob_out_post[30], \kme_cddip0_ob_out_post.tdata [30]);
tran (kme_cddip0_ob_out_post[29], \kme_cddip0_ob_out_post.tdata [29]);
tran (kme_cddip0_ob_out_post[28], \kme_cddip0_ob_out_post.tdata [28]);
tran (kme_cddip0_ob_out_post[27], \kme_cddip0_ob_out_post.tdata [27]);
tran (kme_cddip0_ob_out_post[26], \kme_cddip0_ob_out_post.tdata [26]);
tran (kme_cddip0_ob_out_post[25], \kme_cddip0_ob_out_post.tdata [25]);
tran (kme_cddip0_ob_out_post[24], \kme_cddip0_ob_out_post.tdata [24]);
tran (kme_cddip0_ob_out_post[23], \kme_cddip0_ob_out_post.tdata [23]);
tran (kme_cddip0_ob_out_post[22], \kme_cddip0_ob_out_post.tdata [22]);
tran (kme_cddip0_ob_out_post[21], \kme_cddip0_ob_out_post.tdata [21]);
tran (kme_cddip0_ob_out_post[20], \kme_cddip0_ob_out_post.tdata [20]);
tran (kme_cddip0_ob_out_post[19], \kme_cddip0_ob_out_post.tdata [19]);
tran (kme_cddip0_ob_out_post[18], \kme_cddip0_ob_out_post.tdata [18]);
tran (kme_cddip0_ob_out_post[17], \kme_cddip0_ob_out_post.tdata [17]);
tran (kme_cddip0_ob_out_post[16], \kme_cddip0_ob_out_post.tdata [16]);
tran (kme_cddip0_ob_out_post[15], \kme_cddip0_ob_out_post.tdata [15]);
tran (kme_cddip0_ob_out_post[14], \kme_cddip0_ob_out_post.tdata [14]);
tran (kme_cddip0_ob_out_post[13], \kme_cddip0_ob_out_post.tdata [13]);
tran (kme_cddip0_ob_out_post[12], \kme_cddip0_ob_out_post.tdata [12]);
tran (kme_cddip0_ob_out_post[11], \kme_cddip0_ob_out_post.tdata [11]);
tran (kme_cddip0_ob_out_post[10], \kme_cddip0_ob_out_post.tdata [10]);
tran (kme_cddip0_ob_out_post[9], \kme_cddip0_ob_out_post.tdata [9]);
tran (kme_cddip0_ob_out_post[8], \kme_cddip0_ob_out_post.tdata [8]);
tran (kme_cddip0_ob_out_post[7], \kme_cddip0_ob_out_post.tdata [7]);
tran (kme_cddip0_ob_out_post[6], \kme_cddip0_ob_out_post.tdata [6]);
tran (kme_cddip0_ob_out_post[5], \kme_cddip0_ob_out_post.tdata [5]);
tran (kme_cddip0_ob_out_post[4], \kme_cddip0_ob_out_post.tdata [4]);
tran (kme_cddip0_ob_out_post[3], \kme_cddip0_ob_out_post.tdata [3]);
tran (kme_cddip0_ob_out_post[2], \kme_cddip0_ob_out_post.tdata [2]);
tran (kme_cddip0_ob_out_post[1], \kme_cddip0_ob_out_post.tdata [1]);
tran (kme_cddip0_ob_out_post[0], \kme_cddip0_ob_out_post.tdata [0]);
tran (kme_cddip1_ob_out_post[82], \kme_cddip1_ob_out_post.tvalid );
tran (kme_cddip1_ob_out_post[81], \kme_cddip1_ob_out_post.tlast );
tran (kme_cddip1_ob_out_post[80], \kme_cddip1_ob_out_post.tid [0]);
tran (kme_cddip1_ob_out_post[79], \kme_cddip1_ob_out_post.tstrb [7]);
tran (kme_cddip1_ob_out_post[78], \kme_cddip1_ob_out_post.tstrb [6]);
tran (kme_cddip1_ob_out_post[77], \kme_cddip1_ob_out_post.tstrb [5]);
tran (kme_cddip1_ob_out_post[76], \kme_cddip1_ob_out_post.tstrb [4]);
tran (kme_cddip1_ob_out_post[75], \kme_cddip1_ob_out_post.tstrb [3]);
tran (kme_cddip1_ob_out_post[74], \kme_cddip1_ob_out_post.tstrb [2]);
tran (kme_cddip1_ob_out_post[73], \kme_cddip1_ob_out_post.tstrb [1]);
tran (kme_cddip1_ob_out_post[72], \kme_cddip1_ob_out_post.tstrb [0]);
tran (kme_cddip1_ob_out_post[71], \kme_cddip1_ob_out_post.tuser [7]);
tran (kme_cddip1_ob_out_post[70], \kme_cddip1_ob_out_post.tuser [6]);
tran (kme_cddip1_ob_out_post[69], \kme_cddip1_ob_out_post.tuser [5]);
tran (kme_cddip1_ob_out_post[68], \kme_cddip1_ob_out_post.tuser [4]);
tran (kme_cddip1_ob_out_post[67], \kme_cddip1_ob_out_post.tuser [3]);
tran (kme_cddip1_ob_out_post[66], \kme_cddip1_ob_out_post.tuser [2]);
tran (kme_cddip1_ob_out_post[65], \kme_cddip1_ob_out_post.tuser [1]);
tran (kme_cddip1_ob_out_post[64], \kme_cddip1_ob_out_post.tuser [0]);
tran (kme_cddip1_ob_out_post[63], \kme_cddip1_ob_out_post.tdata [63]);
tran (kme_cddip1_ob_out_post[62], \kme_cddip1_ob_out_post.tdata [62]);
tran (kme_cddip1_ob_out_post[61], \kme_cddip1_ob_out_post.tdata [61]);
tran (kme_cddip1_ob_out_post[60], \kme_cddip1_ob_out_post.tdata [60]);
tran (kme_cddip1_ob_out_post[59], \kme_cddip1_ob_out_post.tdata [59]);
tran (kme_cddip1_ob_out_post[58], \kme_cddip1_ob_out_post.tdata [58]);
tran (kme_cddip1_ob_out_post[57], \kme_cddip1_ob_out_post.tdata [57]);
tran (kme_cddip1_ob_out_post[56], \kme_cddip1_ob_out_post.tdata [56]);
tran (kme_cddip1_ob_out_post[55], \kme_cddip1_ob_out_post.tdata [55]);
tran (kme_cddip1_ob_out_post[54], \kme_cddip1_ob_out_post.tdata [54]);
tran (kme_cddip1_ob_out_post[53], \kme_cddip1_ob_out_post.tdata [53]);
tran (kme_cddip1_ob_out_post[52], \kme_cddip1_ob_out_post.tdata [52]);
tran (kme_cddip1_ob_out_post[51], \kme_cddip1_ob_out_post.tdata [51]);
tran (kme_cddip1_ob_out_post[50], \kme_cddip1_ob_out_post.tdata [50]);
tran (kme_cddip1_ob_out_post[49], \kme_cddip1_ob_out_post.tdata [49]);
tran (kme_cddip1_ob_out_post[48], \kme_cddip1_ob_out_post.tdata [48]);
tran (kme_cddip1_ob_out_post[47], \kme_cddip1_ob_out_post.tdata [47]);
tran (kme_cddip1_ob_out_post[46], \kme_cddip1_ob_out_post.tdata [46]);
tran (kme_cddip1_ob_out_post[45], \kme_cddip1_ob_out_post.tdata [45]);
tran (kme_cddip1_ob_out_post[44], \kme_cddip1_ob_out_post.tdata [44]);
tran (kme_cddip1_ob_out_post[43], \kme_cddip1_ob_out_post.tdata [43]);
tran (kme_cddip1_ob_out_post[42], \kme_cddip1_ob_out_post.tdata [42]);
tran (kme_cddip1_ob_out_post[41], \kme_cddip1_ob_out_post.tdata [41]);
tran (kme_cddip1_ob_out_post[40], \kme_cddip1_ob_out_post.tdata [40]);
tran (kme_cddip1_ob_out_post[39], \kme_cddip1_ob_out_post.tdata [39]);
tran (kme_cddip1_ob_out_post[38], \kme_cddip1_ob_out_post.tdata [38]);
tran (kme_cddip1_ob_out_post[37], \kme_cddip1_ob_out_post.tdata [37]);
tran (kme_cddip1_ob_out_post[36], \kme_cddip1_ob_out_post.tdata [36]);
tran (kme_cddip1_ob_out_post[35], \kme_cddip1_ob_out_post.tdata [35]);
tran (kme_cddip1_ob_out_post[34], \kme_cddip1_ob_out_post.tdata [34]);
tran (kme_cddip1_ob_out_post[33], \kme_cddip1_ob_out_post.tdata [33]);
tran (kme_cddip1_ob_out_post[32], \kme_cddip1_ob_out_post.tdata [32]);
tran (kme_cddip1_ob_out_post[31], \kme_cddip1_ob_out_post.tdata [31]);
tran (kme_cddip1_ob_out_post[30], \kme_cddip1_ob_out_post.tdata [30]);
tran (kme_cddip1_ob_out_post[29], \kme_cddip1_ob_out_post.tdata [29]);
tran (kme_cddip1_ob_out_post[28], \kme_cddip1_ob_out_post.tdata [28]);
tran (kme_cddip1_ob_out_post[27], \kme_cddip1_ob_out_post.tdata [27]);
tran (kme_cddip1_ob_out_post[26], \kme_cddip1_ob_out_post.tdata [26]);
tran (kme_cddip1_ob_out_post[25], \kme_cddip1_ob_out_post.tdata [25]);
tran (kme_cddip1_ob_out_post[24], \kme_cddip1_ob_out_post.tdata [24]);
tran (kme_cddip1_ob_out_post[23], \kme_cddip1_ob_out_post.tdata [23]);
tran (kme_cddip1_ob_out_post[22], \kme_cddip1_ob_out_post.tdata [22]);
tran (kme_cddip1_ob_out_post[21], \kme_cddip1_ob_out_post.tdata [21]);
tran (kme_cddip1_ob_out_post[20], \kme_cddip1_ob_out_post.tdata [20]);
tran (kme_cddip1_ob_out_post[19], \kme_cddip1_ob_out_post.tdata [19]);
tran (kme_cddip1_ob_out_post[18], \kme_cddip1_ob_out_post.tdata [18]);
tran (kme_cddip1_ob_out_post[17], \kme_cddip1_ob_out_post.tdata [17]);
tran (kme_cddip1_ob_out_post[16], \kme_cddip1_ob_out_post.tdata [16]);
tran (kme_cddip1_ob_out_post[15], \kme_cddip1_ob_out_post.tdata [15]);
tran (kme_cddip1_ob_out_post[14], \kme_cddip1_ob_out_post.tdata [14]);
tran (kme_cddip1_ob_out_post[13], \kme_cddip1_ob_out_post.tdata [13]);
tran (kme_cddip1_ob_out_post[12], \kme_cddip1_ob_out_post.tdata [12]);
tran (kme_cddip1_ob_out_post[11], \kme_cddip1_ob_out_post.tdata [11]);
tran (kme_cddip1_ob_out_post[10], \kme_cddip1_ob_out_post.tdata [10]);
tran (kme_cddip1_ob_out_post[9], \kme_cddip1_ob_out_post.tdata [9]);
tran (kme_cddip1_ob_out_post[8], \kme_cddip1_ob_out_post.tdata [8]);
tran (kme_cddip1_ob_out_post[7], \kme_cddip1_ob_out_post.tdata [7]);
tran (kme_cddip1_ob_out_post[6], \kme_cddip1_ob_out_post.tdata [6]);
tran (kme_cddip1_ob_out_post[5], \kme_cddip1_ob_out_post.tdata [5]);
tran (kme_cddip1_ob_out_post[4], \kme_cddip1_ob_out_post.tdata [4]);
tran (kme_cddip1_ob_out_post[3], \kme_cddip1_ob_out_post.tdata [3]);
tran (kme_cddip1_ob_out_post[2], \kme_cddip1_ob_out_post.tdata [2]);
tran (kme_cddip1_ob_out_post[1], \kme_cddip1_ob_out_post.tdata [1]);
tran (kme_cddip1_ob_out_post[0], \kme_cddip1_ob_out_post.tdata [0]);
tran (kme_cddip2_ob_out_post[82], \kme_cddip2_ob_out_post.tvalid );
tran (kme_cddip2_ob_out_post[81], \kme_cddip2_ob_out_post.tlast );
tran (kme_cddip2_ob_out_post[80], \kme_cddip2_ob_out_post.tid [0]);
tran (kme_cddip2_ob_out_post[79], \kme_cddip2_ob_out_post.tstrb [7]);
tran (kme_cddip2_ob_out_post[78], \kme_cddip2_ob_out_post.tstrb [6]);
tran (kme_cddip2_ob_out_post[77], \kme_cddip2_ob_out_post.tstrb [5]);
tran (kme_cddip2_ob_out_post[76], \kme_cddip2_ob_out_post.tstrb [4]);
tran (kme_cddip2_ob_out_post[75], \kme_cddip2_ob_out_post.tstrb [3]);
tran (kme_cddip2_ob_out_post[74], \kme_cddip2_ob_out_post.tstrb [2]);
tran (kme_cddip2_ob_out_post[73], \kme_cddip2_ob_out_post.tstrb [1]);
tran (kme_cddip2_ob_out_post[72], \kme_cddip2_ob_out_post.tstrb [0]);
tran (kme_cddip2_ob_out_post[71], \kme_cddip2_ob_out_post.tuser [7]);
tran (kme_cddip2_ob_out_post[70], \kme_cddip2_ob_out_post.tuser [6]);
tran (kme_cddip2_ob_out_post[69], \kme_cddip2_ob_out_post.tuser [5]);
tran (kme_cddip2_ob_out_post[68], \kme_cddip2_ob_out_post.tuser [4]);
tran (kme_cddip2_ob_out_post[67], \kme_cddip2_ob_out_post.tuser [3]);
tran (kme_cddip2_ob_out_post[66], \kme_cddip2_ob_out_post.tuser [2]);
tran (kme_cddip2_ob_out_post[65], \kme_cddip2_ob_out_post.tuser [1]);
tran (kme_cddip2_ob_out_post[64], \kme_cddip2_ob_out_post.tuser [0]);
tran (kme_cddip2_ob_out_post[63], \kme_cddip2_ob_out_post.tdata [63]);
tran (kme_cddip2_ob_out_post[62], \kme_cddip2_ob_out_post.tdata [62]);
tran (kme_cddip2_ob_out_post[61], \kme_cddip2_ob_out_post.tdata [61]);
tran (kme_cddip2_ob_out_post[60], \kme_cddip2_ob_out_post.tdata [60]);
tran (kme_cddip2_ob_out_post[59], \kme_cddip2_ob_out_post.tdata [59]);
tran (kme_cddip2_ob_out_post[58], \kme_cddip2_ob_out_post.tdata [58]);
tran (kme_cddip2_ob_out_post[57], \kme_cddip2_ob_out_post.tdata [57]);
tran (kme_cddip2_ob_out_post[56], \kme_cddip2_ob_out_post.tdata [56]);
tran (kme_cddip2_ob_out_post[55], \kme_cddip2_ob_out_post.tdata [55]);
tran (kme_cddip2_ob_out_post[54], \kme_cddip2_ob_out_post.tdata [54]);
tran (kme_cddip2_ob_out_post[53], \kme_cddip2_ob_out_post.tdata [53]);
tran (kme_cddip2_ob_out_post[52], \kme_cddip2_ob_out_post.tdata [52]);
tran (kme_cddip2_ob_out_post[51], \kme_cddip2_ob_out_post.tdata [51]);
tran (kme_cddip2_ob_out_post[50], \kme_cddip2_ob_out_post.tdata [50]);
tran (kme_cddip2_ob_out_post[49], \kme_cddip2_ob_out_post.tdata [49]);
tran (kme_cddip2_ob_out_post[48], \kme_cddip2_ob_out_post.tdata [48]);
tran (kme_cddip2_ob_out_post[47], \kme_cddip2_ob_out_post.tdata [47]);
tran (kme_cddip2_ob_out_post[46], \kme_cddip2_ob_out_post.tdata [46]);
tran (kme_cddip2_ob_out_post[45], \kme_cddip2_ob_out_post.tdata [45]);
tran (kme_cddip2_ob_out_post[44], \kme_cddip2_ob_out_post.tdata [44]);
tran (kme_cddip2_ob_out_post[43], \kme_cddip2_ob_out_post.tdata [43]);
tran (kme_cddip2_ob_out_post[42], \kme_cddip2_ob_out_post.tdata [42]);
tran (kme_cddip2_ob_out_post[41], \kme_cddip2_ob_out_post.tdata [41]);
tran (kme_cddip2_ob_out_post[40], \kme_cddip2_ob_out_post.tdata [40]);
tran (kme_cddip2_ob_out_post[39], \kme_cddip2_ob_out_post.tdata [39]);
tran (kme_cddip2_ob_out_post[38], \kme_cddip2_ob_out_post.tdata [38]);
tran (kme_cddip2_ob_out_post[37], \kme_cddip2_ob_out_post.tdata [37]);
tran (kme_cddip2_ob_out_post[36], \kme_cddip2_ob_out_post.tdata [36]);
tran (kme_cddip2_ob_out_post[35], \kme_cddip2_ob_out_post.tdata [35]);
tran (kme_cddip2_ob_out_post[34], \kme_cddip2_ob_out_post.tdata [34]);
tran (kme_cddip2_ob_out_post[33], \kme_cddip2_ob_out_post.tdata [33]);
tran (kme_cddip2_ob_out_post[32], \kme_cddip2_ob_out_post.tdata [32]);
tran (kme_cddip2_ob_out_post[31], \kme_cddip2_ob_out_post.tdata [31]);
tran (kme_cddip2_ob_out_post[30], \kme_cddip2_ob_out_post.tdata [30]);
tran (kme_cddip2_ob_out_post[29], \kme_cddip2_ob_out_post.tdata [29]);
tran (kme_cddip2_ob_out_post[28], \kme_cddip2_ob_out_post.tdata [28]);
tran (kme_cddip2_ob_out_post[27], \kme_cddip2_ob_out_post.tdata [27]);
tran (kme_cddip2_ob_out_post[26], \kme_cddip2_ob_out_post.tdata [26]);
tran (kme_cddip2_ob_out_post[25], \kme_cddip2_ob_out_post.tdata [25]);
tran (kme_cddip2_ob_out_post[24], \kme_cddip2_ob_out_post.tdata [24]);
tran (kme_cddip2_ob_out_post[23], \kme_cddip2_ob_out_post.tdata [23]);
tran (kme_cddip2_ob_out_post[22], \kme_cddip2_ob_out_post.tdata [22]);
tran (kme_cddip2_ob_out_post[21], \kme_cddip2_ob_out_post.tdata [21]);
tran (kme_cddip2_ob_out_post[20], \kme_cddip2_ob_out_post.tdata [20]);
tran (kme_cddip2_ob_out_post[19], \kme_cddip2_ob_out_post.tdata [19]);
tran (kme_cddip2_ob_out_post[18], \kme_cddip2_ob_out_post.tdata [18]);
tran (kme_cddip2_ob_out_post[17], \kme_cddip2_ob_out_post.tdata [17]);
tran (kme_cddip2_ob_out_post[16], \kme_cddip2_ob_out_post.tdata [16]);
tran (kme_cddip2_ob_out_post[15], \kme_cddip2_ob_out_post.tdata [15]);
tran (kme_cddip2_ob_out_post[14], \kme_cddip2_ob_out_post.tdata [14]);
tran (kme_cddip2_ob_out_post[13], \kme_cddip2_ob_out_post.tdata [13]);
tran (kme_cddip2_ob_out_post[12], \kme_cddip2_ob_out_post.tdata [12]);
tran (kme_cddip2_ob_out_post[11], \kme_cddip2_ob_out_post.tdata [11]);
tran (kme_cddip2_ob_out_post[10], \kme_cddip2_ob_out_post.tdata [10]);
tran (kme_cddip2_ob_out_post[9], \kme_cddip2_ob_out_post.tdata [9]);
tran (kme_cddip2_ob_out_post[8], \kme_cddip2_ob_out_post.tdata [8]);
tran (kme_cddip2_ob_out_post[7], \kme_cddip2_ob_out_post.tdata [7]);
tran (kme_cddip2_ob_out_post[6], \kme_cddip2_ob_out_post.tdata [6]);
tran (kme_cddip2_ob_out_post[5], \kme_cddip2_ob_out_post.tdata [5]);
tran (kme_cddip2_ob_out_post[4], \kme_cddip2_ob_out_post.tdata [4]);
tran (kme_cddip2_ob_out_post[3], \kme_cddip2_ob_out_post.tdata [3]);
tran (kme_cddip2_ob_out_post[2], \kme_cddip2_ob_out_post.tdata [2]);
tran (kme_cddip2_ob_out_post[1], \kme_cddip2_ob_out_post.tdata [1]);
tran (kme_cddip2_ob_out_post[0], \kme_cddip2_ob_out_post.tdata [0]);
tran (kme_cddip3_ob_out_post[82], \kme_cddip3_ob_out_post.tvalid );
tran (kme_cddip3_ob_out_post[81], \kme_cddip3_ob_out_post.tlast );
tran (kme_cddip3_ob_out_post[80], \kme_cddip3_ob_out_post.tid [0]);
tran (kme_cddip3_ob_out_post[79], \kme_cddip3_ob_out_post.tstrb [7]);
tran (kme_cddip3_ob_out_post[78], \kme_cddip3_ob_out_post.tstrb [6]);
tran (kme_cddip3_ob_out_post[77], \kme_cddip3_ob_out_post.tstrb [5]);
tran (kme_cddip3_ob_out_post[76], \kme_cddip3_ob_out_post.tstrb [4]);
tran (kme_cddip3_ob_out_post[75], \kme_cddip3_ob_out_post.tstrb [3]);
tran (kme_cddip3_ob_out_post[74], \kme_cddip3_ob_out_post.tstrb [2]);
tran (kme_cddip3_ob_out_post[73], \kme_cddip3_ob_out_post.tstrb [1]);
tran (kme_cddip3_ob_out_post[72], \kme_cddip3_ob_out_post.tstrb [0]);
tran (kme_cddip3_ob_out_post[71], \kme_cddip3_ob_out_post.tuser [7]);
tran (kme_cddip3_ob_out_post[70], \kme_cddip3_ob_out_post.tuser [6]);
tran (kme_cddip3_ob_out_post[69], \kme_cddip3_ob_out_post.tuser [5]);
tran (kme_cddip3_ob_out_post[68], \kme_cddip3_ob_out_post.tuser [4]);
tran (kme_cddip3_ob_out_post[67], \kme_cddip3_ob_out_post.tuser [3]);
tran (kme_cddip3_ob_out_post[66], \kme_cddip3_ob_out_post.tuser [2]);
tran (kme_cddip3_ob_out_post[65], \kme_cddip3_ob_out_post.tuser [1]);
tran (kme_cddip3_ob_out_post[64], \kme_cddip3_ob_out_post.tuser [0]);
tran (kme_cddip3_ob_out_post[63], \kme_cddip3_ob_out_post.tdata [63]);
tran (kme_cddip3_ob_out_post[62], \kme_cddip3_ob_out_post.tdata [62]);
tran (kme_cddip3_ob_out_post[61], \kme_cddip3_ob_out_post.tdata [61]);
tran (kme_cddip3_ob_out_post[60], \kme_cddip3_ob_out_post.tdata [60]);
tran (kme_cddip3_ob_out_post[59], \kme_cddip3_ob_out_post.tdata [59]);
tran (kme_cddip3_ob_out_post[58], \kme_cddip3_ob_out_post.tdata [58]);
tran (kme_cddip3_ob_out_post[57], \kme_cddip3_ob_out_post.tdata [57]);
tran (kme_cddip3_ob_out_post[56], \kme_cddip3_ob_out_post.tdata [56]);
tran (kme_cddip3_ob_out_post[55], \kme_cddip3_ob_out_post.tdata [55]);
tran (kme_cddip3_ob_out_post[54], \kme_cddip3_ob_out_post.tdata [54]);
tran (kme_cddip3_ob_out_post[53], \kme_cddip3_ob_out_post.tdata [53]);
tran (kme_cddip3_ob_out_post[52], \kme_cddip3_ob_out_post.tdata [52]);
tran (kme_cddip3_ob_out_post[51], \kme_cddip3_ob_out_post.tdata [51]);
tran (kme_cddip3_ob_out_post[50], \kme_cddip3_ob_out_post.tdata [50]);
tran (kme_cddip3_ob_out_post[49], \kme_cddip3_ob_out_post.tdata [49]);
tran (kme_cddip3_ob_out_post[48], \kme_cddip3_ob_out_post.tdata [48]);
tran (kme_cddip3_ob_out_post[47], \kme_cddip3_ob_out_post.tdata [47]);
tran (kme_cddip3_ob_out_post[46], \kme_cddip3_ob_out_post.tdata [46]);
tran (kme_cddip3_ob_out_post[45], \kme_cddip3_ob_out_post.tdata [45]);
tran (kme_cddip3_ob_out_post[44], \kme_cddip3_ob_out_post.tdata [44]);
tran (kme_cddip3_ob_out_post[43], \kme_cddip3_ob_out_post.tdata [43]);
tran (kme_cddip3_ob_out_post[42], \kme_cddip3_ob_out_post.tdata [42]);
tran (kme_cddip3_ob_out_post[41], \kme_cddip3_ob_out_post.tdata [41]);
tran (kme_cddip3_ob_out_post[40], \kme_cddip3_ob_out_post.tdata [40]);
tran (kme_cddip3_ob_out_post[39], \kme_cddip3_ob_out_post.tdata [39]);
tran (kme_cddip3_ob_out_post[38], \kme_cddip3_ob_out_post.tdata [38]);
tran (kme_cddip3_ob_out_post[37], \kme_cddip3_ob_out_post.tdata [37]);
tran (kme_cddip3_ob_out_post[36], \kme_cddip3_ob_out_post.tdata [36]);
tran (kme_cddip3_ob_out_post[35], \kme_cddip3_ob_out_post.tdata [35]);
tran (kme_cddip3_ob_out_post[34], \kme_cddip3_ob_out_post.tdata [34]);
tran (kme_cddip3_ob_out_post[33], \kme_cddip3_ob_out_post.tdata [33]);
tran (kme_cddip3_ob_out_post[32], \kme_cddip3_ob_out_post.tdata [32]);
tran (kme_cddip3_ob_out_post[31], \kme_cddip3_ob_out_post.tdata [31]);
tran (kme_cddip3_ob_out_post[30], \kme_cddip3_ob_out_post.tdata [30]);
tran (kme_cddip3_ob_out_post[29], \kme_cddip3_ob_out_post.tdata [29]);
tran (kme_cddip3_ob_out_post[28], \kme_cddip3_ob_out_post.tdata [28]);
tran (kme_cddip3_ob_out_post[27], \kme_cddip3_ob_out_post.tdata [27]);
tran (kme_cddip3_ob_out_post[26], \kme_cddip3_ob_out_post.tdata [26]);
tran (kme_cddip3_ob_out_post[25], \kme_cddip3_ob_out_post.tdata [25]);
tran (kme_cddip3_ob_out_post[24], \kme_cddip3_ob_out_post.tdata [24]);
tran (kme_cddip3_ob_out_post[23], \kme_cddip3_ob_out_post.tdata [23]);
tran (kme_cddip3_ob_out_post[22], \kme_cddip3_ob_out_post.tdata [22]);
tran (kme_cddip3_ob_out_post[21], \kme_cddip3_ob_out_post.tdata [21]);
tran (kme_cddip3_ob_out_post[20], \kme_cddip3_ob_out_post.tdata [20]);
tran (kme_cddip3_ob_out_post[19], \kme_cddip3_ob_out_post.tdata [19]);
tran (kme_cddip3_ob_out_post[18], \kme_cddip3_ob_out_post.tdata [18]);
tran (kme_cddip3_ob_out_post[17], \kme_cddip3_ob_out_post.tdata [17]);
tran (kme_cddip3_ob_out_post[16], \kme_cddip3_ob_out_post.tdata [16]);
tran (kme_cddip3_ob_out_post[15], \kme_cddip3_ob_out_post.tdata [15]);
tran (kme_cddip3_ob_out_post[14], \kme_cddip3_ob_out_post.tdata [14]);
tran (kme_cddip3_ob_out_post[13], \kme_cddip3_ob_out_post.tdata [13]);
tran (kme_cddip3_ob_out_post[12], \kme_cddip3_ob_out_post.tdata [12]);
tran (kme_cddip3_ob_out_post[11], \kme_cddip3_ob_out_post.tdata [11]);
tran (kme_cddip3_ob_out_post[10], \kme_cddip3_ob_out_post.tdata [10]);
tran (kme_cddip3_ob_out_post[9], \kme_cddip3_ob_out_post.tdata [9]);
tran (kme_cddip3_ob_out_post[8], \kme_cddip3_ob_out_post.tdata [8]);
tran (kme_cddip3_ob_out_post[7], \kme_cddip3_ob_out_post.tdata [7]);
tran (kme_cddip3_ob_out_post[6], \kme_cddip3_ob_out_post.tdata [6]);
tran (kme_cddip3_ob_out_post[5], \kme_cddip3_ob_out_post.tdata [5]);
tran (kme_cddip3_ob_out_post[4], \kme_cddip3_ob_out_post.tdata [4]);
tran (kme_cddip3_ob_out_post[3], \kme_cddip3_ob_out_post.tdata [3]);
tran (kme_cddip3_ob_out_post[2], \kme_cddip3_ob_out_post.tdata [2]);
tran (kme_cddip3_ob_out_post[1], \kme_cddip3_ob_out_post.tdata [1]);
tran (kme_cddip3_ob_out_post[0], \kme_cddip3_ob_out_post.tdata [0]);
Q_BUF U0 ( .A(send_kme_ib_beat), .Z(debug_kme_ib_tvalid));
Q_ASSIGN U1 ( .B(kme_cceip0_ob_out_post[81]), .A(kme_cceip0_ob_out[81]));
Q_ASSIGN U2 ( .B(kme_cceip0_ob_out_post[80]), .A(kme_cceip0_ob_out[80]));
Q_ASSIGN U3 ( .B(kme_cceip0_ob_out_post[79]), .A(kme_cceip0_ob_out[79]));
Q_ASSIGN U4 ( .B(kme_cceip0_ob_out_post[78]), .A(kme_cceip0_ob_out[78]));
Q_ASSIGN U5 ( .B(kme_cceip0_ob_out_post[77]), .A(kme_cceip0_ob_out[77]));
Q_ASSIGN U6 ( .B(kme_cceip0_ob_out_post[76]), .A(kme_cceip0_ob_out[76]));
Q_ASSIGN U7 ( .B(kme_cceip0_ob_out_post[75]), .A(kme_cceip0_ob_out[75]));
Q_ASSIGN U8 ( .B(kme_cceip0_ob_out_post[74]), .A(kme_cceip0_ob_out[74]));
Q_ASSIGN U9 ( .B(kme_cceip0_ob_out_post[73]), .A(kme_cceip0_ob_out[73]));
Q_ASSIGN U10 ( .B(kme_cceip0_ob_out_post[72]), .A(kme_cceip0_ob_out[72]));
Q_ASSIGN U11 ( .B(kme_cceip0_ob_out_post[71]), .A(kme_cceip0_ob_out[71]));
Q_ASSIGN U12 ( .B(kme_cceip0_ob_out_post[70]), .A(kme_cceip0_ob_out[70]));
Q_ASSIGN U13 ( .B(kme_cceip0_ob_out_post[69]), .A(kme_cceip0_ob_out[69]));
Q_ASSIGN U14 ( .B(kme_cceip0_ob_out_post[68]), .A(kme_cceip0_ob_out[68]));
Q_ASSIGN U15 ( .B(kme_cceip0_ob_out_post[67]), .A(kme_cceip0_ob_out[67]));
Q_ASSIGN U16 ( .B(kme_cceip0_ob_out_post[66]), .A(kme_cceip0_ob_out[66]));
Q_ASSIGN U17 ( .B(kme_cceip0_ob_out_post[65]), .A(kme_cceip0_ob_out[65]));
Q_ASSIGN U18 ( .B(kme_cceip0_ob_out_post[64]), .A(kme_cceip0_ob_out[64]));
Q_ASSIGN U19 ( .B(kme_cceip0_ob_out_post[63]), .A(kme_cceip0_ob_out[63]));
Q_ASSIGN U20 ( .B(kme_cceip0_ob_out_post[62]), .A(kme_cceip0_ob_out[62]));
Q_ASSIGN U21 ( .B(kme_cceip0_ob_out_post[61]), .A(kme_cceip0_ob_out[61]));
Q_ASSIGN U22 ( .B(kme_cceip0_ob_out_post[60]), .A(kme_cceip0_ob_out[60]));
Q_ASSIGN U23 ( .B(kme_cceip0_ob_out_post[59]), .A(kme_cceip0_ob_out[59]));
Q_ASSIGN U24 ( .B(kme_cceip0_ob_out_post[58]), .A(kme_cceip0_ob_out[58]));
Q_ASSIGN U25 ( .B(kme_cceip0_ob_out_post[57]), .A(kme_cceip0_ob_out[57]));
Q_ASSIGN U26 ( .B(kme_cceip0_ob_out_post[56]), .A(kme_cceip0_ob_out[56]));
Q_ASSIGN U27 ( .B(kme_cceip0_ob_out_post[55]), .A(kme_cceip0_ob_out[55]));
Q_ASSIGN U28 ( .B(kme_cceip0_ob_out_post[54]), .A(kme_cceip0_ob_out[54]));
Q_ASSIGN U29 ( .B(kme_cceip0_ob_out_post[53]), .A(kme_cceip0_ob_out[53]));
Q_ASSIGN U30 ( .B(kme_cceip0_ob_out_post[52]), .A(kme_cceip0_ob_out[52]));
Q_ASSIGN U31 ( .B(kme_cceip0_ob_out_post[51]), .A(kme_cceip0_ob_out[51]));
Q_ASSIGN U32 ( .B(kme_cceip0_ob_out_post[50]), .A(kme_cceip0_ob_out[50]));
Q_ASSIGN U33 ( .B(kme_cceip0_ob_out_post[49]), .A(kme_cceip0_ob_out[49]));
Q_ASSIGN U34 ( .B(kme_cceip0_ob_out_post[48]), .A(kme_cceip0_ob_out[48]));
Q_ASSIGN U35 ( .B(kme_cceip0_ob_out_post[47]), .A(kme_cceip0_ob_out[47]));
Q_ASSIGN U36 ( .B(kme_cceip0_ob_out_post[46]), .A(kme_cceip0_ob_out[46]));
Q_ASSIGN U37 ( .B(kme_cceip0_ob_out_post[45]), .A(kme_cceip0_ob_out[45]));
Q_ASSIGN U38 ( .B(kme_cceip0_ob_out_post[44]), .A(kme_cceip0_ob_out[44]));
Q_ASSIGN U39 ( .B(kme_cceip0_ob_out_post[43]), .A(kme_cceip0_ob_out[43]));
Q_ASSIGN U40 ( .B(kme_cceip0_ob_out_post[42]), .A(kme_cceip0_ob_out[42]));
Q_ASSIGN U41 ( .B(kme_cceip0_ob_out_post[41]), .A(kme_cceip0_ob_out[41]));
Q_ASSIGN U42 ( .B(kme_cceip0_ob_out_post[40]), .A(kme_cceip0_ob_out[40]));
Q_ASSIGN U43 ( .B(kme_cceip0_ob_out_post[39]), .A(kme_cceip0_ob_out[39]));
Q_ASSIGN U44 ( .B(kme_cceip0_ob_out_post[38]), .A(kme_cceip0_ob_out[38]));
Q_ASSIGN U45 ( .B(kme_cceip0_ob_out_post[37]), .A(kme_cceip0_ob_out[37]));
Q_ASSIGN U46 ( .B(kme_cceip0_ob_out_post[36]), .A(kme_cceip0_ob_out[36]));
Q_ASSIGN U47 ( .B(kme_cceip0_ob_out_post[35]), .A(kme_cceip0_ob_out[35]));
Q_ASSIGN U48 ( .B(kme_cceip0_ob_out_post[34]), .A(kme_cceip0_ob_out[34]));
Q_ASSIGN U49 ( .B(kme_cceip0_ob_out_post[33]), .A(kme_cceip0_ob_out[33]));
Q_ASSIGN U50 ( .B(kme_cceip0_ob_out_post[32]), .A(kme_cceip0_ob_out[32]));
Q_ASSIGN U51 ( .B(kme_cceip0_ob_out_post[31]), .A(kme_cceip0_ob_out[31]));
Q_ASSIGN U52 ( .B(kme_cceip0_ob_out_post[30]), .A(kme_cceip0_ob_out[30]));
Q_ASSIGN U53 ( .B(kme_cceip0_ob_out_post[29]), .A(kme_cceip0_ob_out[29]));
Q_ASSIGN U54 ( .B(kme_cceip0_ob_out_post[28]), .A(kme_cceip0_ob_out[28]));
Q_ASSIGN U55 ( .B(kme_cceip0_ob_out_post[27]), .A(kme_cceip0_ob_out[27]));
Q_ASSIGN U56 ( .B(kme_cceip0_ob_out_post[26]), .A(kme_cceip0_ob_out[26]));
Q_ASSIGN U57 ( .B(kme_cceip0_ob_out_post[25]), .A(kme_cceip0_ob_out[25]));
Q_ASSIGN U58 ( .B(kme_cceip0_ob_out_post[24]), .A(kme_cceip0_ob_out[24]));
Q_ASSIGN U59 ( .B(kme_cceip0_ob_out_post[23]), .A(kme_cceip0_ob_out[23]));
Q_ASSIGN U60 ( .B(kme_cceip0_ob_out_post[22]), .A(kme_cceip0_ob_out[22]));
Q_ASSIGN U61 ( .B(kme_cceip0_ob_out_post[21]), .A(kme_cceip0_ob_out[21]));
Q_ASSIGN U62 ( .B(kme_cceip0_ob_out_post[20]), .A(kme_cceip0_ob_out[20]));
Q_ASSIGN U63 ( .B(kme_cceip0_ob_out_post[19]), .A(kme_cceip0_ob_out[19]));
Q_ASSIGN U64 ( .B(kme_cceip0_ob_out_post[18]), .A(kme_cceip0_ob_out[18]));
Q_ASSIGN U65 ( .B(kme_cceip0_ob_out_post[17]), .A(kme_cceip0_ob_out[17]));
Q_ASSIGN U66 ( .B(kme_cceip0_ob_out_post[16]), .A(kme_cceip0_ob_out[16]));
Q_ASSIGN U67 ( .B(kme_cceip0_ob_out_post[15]), .A(kme_cceip0_ob_out[15]));
Q_ASSIGN U68 ( .B(kme_cceip0_ob_out_post[14]), .A(kme_cceip0_ob_out[14]));
Q_ASSIGN U69 ( .B(kme_cceip0_ob_out_post[13]), .A(kme_cceip0_ob_out[13]));
Q_ASSIGN U70 ( .B(kme_cceip0_ob_out_post[12]), .A(kme_cceip0_ob_out[12]));
Q_ASSIGN U71 ( .B(kme_cceip0_ob_out_post[11]), .A(kme_cceip0_ob_out[11]));
Q_ASSIGN U72 ( .B(kme_cceip0_ob_out_post[10]), .A(kme_cceip0_ob_out[10]));
Q_ASSIGN U73 ( .B(kme_cceip0_ob_out_post[9]), .A(kme_cceip0_ob_out[9]));
Q_ASSIGN U74 ( .B(kme_cceip0_ob_out_post[8]), .A(kme_cceip0_ob_out[8]));
Q_ASSIGN U75 ( .B(kme_cceip0_ob_out_post[7]), .A(kme_cceip0_ob_out[7]));
Q_ASSIGN U76 ( .B(kme_cceip0_ob_out_post[6]), .A(kme_cceip0_ob_out[6]));
Q_ASSIGN U77 ( .B(kme_cceip0_ob_out_post[5]), .A(kme_cceip0_ob_out[5]));
Q_ASSIGN U78 ( .B(kme_cceip0_ob_out_post[4]), .A(kme_cceip0_ob_out[4]));
Q_ASSIGN U79 ( .B(kme_cceip0_ob_out_post[3]), .A(kme_cceip0_ob_out[3]));
Q_ASSIGN U80 ( .B(kme_cceip0_ob_out_post[2]), .A(kme_cceip0_ob_out[2]));
Q_ASSIGN U81 ( .B(kme_cceip0_ob_out_post[1]), .A(kme_cceip0_ob_out[1]));
Q_ASSIGN U82 ( .B(kme_cceip0_ob_out_post[0]), .A(kme_cceip0_ob_out[0]));
Q_ASSIGN U83 ( .B(kme_cceip1_ob_out_post[81]), .A(kme_cceip1_ob_out[81]));
Q_ASSIGN U84 ( .B(kme_cceip1_ob_out_post[80]), .A(kme_cceip1_ob_out[80]));
Q_ASSIGN U85 ( .B(kme_cceip1_ob_out_post[79]), .A(kme_cceip1_ob_out[79]));
Q_ASSIGN U86 ( .B(kme_cceip1_ob_out_post[78]), .A(kme_cceip1_ob_out[78]));
Q_ASSIGN U87 ( .B(kme_cceip1_ob_out_post[77]), .A(kme_cceip1_ob_out[77]));
Q_ASSIGN U88 ( .B(kme_cceip1_ob_out_post[76]), .A(kme_cceip1_ob_out[76]));
Q_ASSIGN U89 ( .B(kme_cceip1_ob_out_post[75]), .A(kme_cceip1_ob_out[75]));
Q_ASSIGN U90 ( .B(kme_cceip1_ob_out_post[74]), .A(kme_cceip1_ob_out[74]));
Q_ASSIGN U91 ( .B(kme_cceip1_ob_out_post[73]), .A(kme_cceip1_ob_out[73]));
Q_ASSIGN U92 ( .B(kme_cceip1_ob_out_post[72]), .A(kme_cceip1_ob_out[72]));
Q_ASSIGN U93 ( .B(kme_cceip1_ob_out_post[71]), .A(kme_cceip1_ob_out[71]));
Q_ASSIGN U94 ( .B(kme_cceip1_ob_out_post[70]), .A(kme_cceip1_ob_out[70]));
Q_ASSIGN U95 ( .B(kme_cceip1_ob_out_post[69]), .A(kme_cceip1_ob_out[69]));
Q_ASSIGN U96 ( .B(kme_cceip1_ob_out_post[68]), .A(kme_cceip1_ob_out[68]));
Q_ASSIGN U97 ( .B(kme_cceip1_ob_out_post[67]), .A(kme_cceip1_ob_out[67]));
Q_ASSIGN U98 ( .B(kme_cceip1_ob_out_post[66]), .A(kme_cceip1_ob_out[66]));
Q_ASSIGN U99 ( .B(kme_cceip1_ob_out_post[65]), .A(kme_cceip1_ob_out[65]));
Q_ASSIGN U100 ( .B(kme_cceip1_ob_out_post[64]), .A(kme_cceip1_ob_out[64]));
Q_ASSIGN U101 ( .B(kme_cceip1_ob_out_post[63]), .A(kme_cceip1_ob_out[63]));
Q_ASSIGN U102 ( .B(kme_cceip1_ob_out_post[62]), .A(kme_cceip1_ob_out[62]));
Q_ASSIGN U103 ( .B(kme_cceip1_ob_out_post[61]), .A(kme_cceip1_ob_out[61]));
Q_ASSIGN U104 ( .B(kme_cceip1_ob_out_post[60]), .A(kme_cceip1_ob_out[60]));
Q_ASSIGN U105 ( .B(kme_cceip1_ob_out_post[59]), .A(kme_cceip1_ob_out[59]));
Q_ASSIGN U106 ( .B(kme_cceip1_ob_out_post[58]), .A(kme_cceip1_ob_out[58]));
Q_ASSIGN U107 ( .B(kme_cceip1_ob_out_post[57]), .A(kme_cceip1_ob_out[57]));
Q_ASSIGN U108 ( .B(kme_cceip1_ob_out_post[56]), .A(kme_cceip1_ob_out[56]));
Q_ASSIGN U109 ( .B(kme_cceip1_ob_out_post[55]), .A(kme_cceip1_ob_out[55]));
Q_ASSIGN U110 ( .B(kme_cceip1_ob_out_post[54]), .A(kme_cceip1_ob_out[54]));
Q_ASSIGN U111 ( .B(kme_cceip1_ob_out_post[53]), .A(kme_cceip1_ob_out[53]));
Q_ASSIGN U112 ( .B(kme_cceip1_ob_out_post[52]), .A(kme_cceip1_ob_out[52]));
Q_ASSIGN U113 ( .B(kme_cceip1_ob_out_post[51]), .A(kme_cceip1_ob_out[51]));
Q_ASSIGN U114 ( .B(kme_cceip1_ob_out_post[50]), .A(kme_cceip1_ob_out[50]));
Q_ASSIGN U115 ( .B(kme_cceip1_ob_out_post[49]), .A(kme_cceip1_ob_out[49]));
Q_ASSIGN U116 ( .B(kme_cceip1_ob_out_post[48]), .A(kme_cceip1_ob_out[48]));
Q_ASSIGN U117 ( .B(kme_cceip1_ob_out_post[47]), .A(kme_cceip1_ob_out[47]));
Q_ASSIGN U118 ( .B(kme_cceip1_ob_out_post[46]), .A(kme_cceip1_ob_out[46]));
Q_ASSIGN U119 ( .B(kme_cceip1_ob_out_post[45]), .A(kme_cceip1_ob_out[45]));
Q_ASSIGN U120 ( .B(kme_cceip1_ob_out_post[44]), .A(kme_cceip1_ob_out[44]));
Q_ASSIGN U121 ( .B(kme_cceip1_ob_out_post[43]), .A(kme_cceip1_ob_out[43]));
Q_ASSIGN U122 ( .B(kme_cceip1_ob_out_post[42]), .A(kme_cceip1_ob_out[42]));
Q_ASSIGN U123 ( .B(kme_cceip1_ob_out_post[41]), .A(kme_cceip1_ob_out[41]));
Q_ASSIGN U124 ( .B(kme_cceip1_ob_out_post[40]), .A(kme_cceip1_ob_out[40]));
Q_ASSIGN U125 ( .B(kme_cceip1_ob_out_post[39]), .A(kme_cceip1_ob_out[39]));
Q_ASSIGN U126 ( .B(kme_cceip1_ob_out_post[38]), .A(kme_cceip1_ob_out[38]));
Q_ASSIGN U127 ( .B(kme_cceip1_ob_out_post[37]), .A(kme_cceip1_ob_out[37]));
Q_ASSIGN U128 ( .B(kme_cceip1_ob_out_post[36]), .A(kme_cceip1_ob_out[36]));
Q_ASSIGN U129 ( .B(kme_cceip1_ob_out_post[35]), .A(kme_cceip1_ob_out[35]));
Q_ASSIGN U130 ( .B(kme_cceip1_ob_out_post[34]), .A(kme_cceip1_ob_out[34]));
Q_ASSIGN U131 ( .B(kme_cceip1_ob_out_post[33]), .A(kme_cceip1_ob_out[33]));
Q_ASSIGN U132 ( .B(kme_cceip1_ob_out_post[32]), .A(kme_cceip1_ob_out[32]));
Q_ASSIGN U133 ( .B(kme_cceip1_ob_out_post[31]), .A(kme_cceip1_ob_out[31]));
Q_ASSIGN U134 ( .B(kme_cceip1_ob_out_post[30]), .A(kme_cceip1_ob_out[30]));
Q_ASSIGN U135 ( .B(kme_cceip1_ob_out_post[29]), .A(kme_cceip1_ob_out[29]));
Q_ASSIGN U136 ( .B(kme_cceip1_ob_out_post[28]), .A(kme_cceip1_ob_out[28]));
Q_ASSIGN U137 ( .B(kme_cceip1_ob_out_post[27]), .A(kme_cceip1_ob_out[27]));
Q_ASSIGN U138 ( .B(kme_cceip1_ob_out_post[26]), .A(kme_cceip1_ob_out[26]));
Q_ASSIGN U139 ( .B(kme_cceip1_ob_out_post[25]), .A(kme_cceip1_ob_out[25]));
Q_ASSIGN U140 ( .B(kme_cceip1_ob_out_post[24]), .A(kme_cceip1_ob_out[24]));
Q_ASSIGN U141 ( .B(kme_cceip1_ob_out_post[23]), .A(kme_cceip1_ob_out[23]));
Q_ASSIGN U142 ( .B(kme_cceip1_ob_out_post[22]), .A(kme_cceip1_ob_out[22]));
Q_ASSIGN U143 ( .B(kme_cceip1_ob_out_post[21]), .A(kme_cceip1_ob_out[21]));
Q_ASSIGN U144 ( .B(kme_cceip1_ob_out_post[20]), .A(kme_cceip1_ob_out[20]));
Q_ASSIGN U145 ( .B(kme_cceip1_ob_out_post[19]), .A(kme_cceip1_ob_out[19]));
Q_ASSIGN U146 ( .B(kme_cceip1_ob_out_post[18]), .A(kme_cceip1_ob_out[18]));
Q_ASSIGN U147 ( .B(kme_cceip1_ob_out_post[17]), .A(kme_cceip1_ob_out[17]));
Q_ASSIGN U148 ( .B(kme_cceip1_ob_out_post[16]), .A(kme_cceip1_ob_out[16]));
Q_ASSIGN U149 ( .B(kme_cceip1_ob_out_post[15]), .A(kme_cceip1_ob_out[15]));
Q_ASSIGN U150 ( .B(kme_cceip1_ob_out_post[14]), .A(kme_cceip1_ob_out[14]));
Q_ASSIGN U151 ( .B(kme_cceip1_ob_out_post[13]), .A(kme_cceip1_ob_out[13]));
Q_ASSIGN U152 ( .B(kme_cceip1_ob_out_post[12]), .A(kme_cceip1_ob_out[12]));
Q_ASSIGN U153 ( .B(kme_cceip1_ob_out_post[11]), .A(kme_cceip1_ob_out[11]));
Q_ASSIGN U154 ( .B(kme_cceip1_ob_out_post[10]), .A(kme_cceip1_ob_out[10]));
Q_ASSIGN U155 ( .B(kme_cceip1_ob_out_post[9]), .A(kme_cceip1_ob_out[9]));
Q_ASSIGN U156 ( .B(kme_cceip1_ob_out_post[8]), .A(kme_cceip1_ob_out[8]));
Q_ASSIGN U157 ( .B(kme_cceip1_ob_out_post[7]), .A(kme_cceip1_ob_out[7]));
Q_ASSIGN U158 ( .B(kme_cceip1_ob_out_post[6]), .A(kme_cceip1_ob_out[6]));
Q_ASSIGN U159 ( .B(kme_cceip1_ob_out_post[5]), .A(kme_cceip1_ob_out[5]));
Q_ASSIGN U160 ( .B(kme_cceip1_ob_out_post[4]), .A(kme_cceip1_ob_out[4]));
Q_ASSIGN U161 ( .B(kme_cceip1_ob_out_post[3]), .A(kme_cceip1_ob_out[3]));
Q_ASSIGN U162 ( .B(kme_cceip1_ob_out_post[2]), .A(kme_cceip1_ob_out[2]));
Q_ASSIGN U163 ( .B(kme_cceip1_ob_out_post[1]), .A(kme_cceip1_ob_out[1]));
Q_ASSIGN U164 ( .B(kme_cceip1_ob_out_post[0]), .A(kme_cceip1_ob_out[0]));
Q_ASSIGN U165 ( .B(kme_cceip2_ob_out_post[81]), .A(kme_cceip2_ob_out[81]));
Q_ASSIGN U166 ( .B(kme_cceip2_ob_out_post[80]), .A(kme_cceip2_ob_out[80]));
Q_ASSIGN U167 ( .B(kme_cceip2_ob_out_post[79]), .A(kme_cceip2_ob_out[79]));
Q_ASSIGN U168 ( .B(kme_cceip2_ob_out_post[78]), .A(kme_cceip2_ob_out[78]));
Q_ASSIGN U169 ( .B(kme_cceip2_ob_out_post[77]), .A(kme_cceip2_ob_out[77]));
Q_ASSIGN U170 ( .B(kme_cceip2_ob_out_post[76]), .A(kme_cceip2_ob_out[76]));
Q_ASSIGN U171 ( .B(kme_cceip2_ob_out_post[75]), .A(kme_cceip2_ob_out[75]));
Q_ASSIGN U172 ( .B(kme_cceip2_ob_out_post[74]), .A(kme_cceip2_ob_out[74]));
Q_ASSIGN U173 ( .B(kme_cceip2_ob_out_post[73]), .A(kme_cceip2_ob_out[73]));
Q_ASSIGN U174 ( .B(kme_cceip2_ob_out_post[72]), .A(kme_cceip2_ob_out[72]));
Q_ASSIGN U175 ( .B(kme_cceip2_ob_out_post[71]), .A(kme_cceip2_ob_out[71]));
Q_ASSIGN U176 ( .B(kme_cceip2_ob_out_post[70]), .A(kme_cceip2_ob_out[70]));
Q_ASSIGN U177 ( .B(kme_cceip2_ob_out_post[69]), .A(kme_cceip2_ob_out[69]));
Q_ASSIGN U178 ( .B(kme_cceip2_ob_out_post[68]), .A(kme_cceip2_ob_out[68]));
Q_ASSIGN U179 ( .B(kme_cceip2_ob_out_post[67]), .A(kme_cceip2_ob_out[67]));
Q_ASSIGN U180 ( .B(kme_cceip2_ob_out_post[66]), .A(kme_cceip2_ob_out[66]));
Q_ASSIGN U181 ( .B(kme_cceip2_ob_out_post[65]), .A(kme_cceip2_ob_out[65]));
Q_ASSIGN U182 ( .B(kme_cceip2_ob_out_post[64]), .A(kme_cceip2_ob_out[64]));
Q_ASSIGN U183 ( .B(kme_cceip2_ob_out_post[63]), .A(kme_cceip2_ob_out[63]));
Q_ASSIGN U184 ( .B(kme_cceip2_ob_out_post[62]), .A(kme_cceip2_ob_out[62]));
Q_ASSIGN U185 ( .B(kme_cceip2_ob_out_post[61]), .A(kme_cceip2_ob_out[61]));
Q_ASSIGN U186 ( .B(kme_cceip2_ob_out_post[60]), .A(kme_cceip2_ob_out[60]));
Q_ASSIGN U187 ( .B(kme_cceip2_ob_out_post[59]), .A(kme_cceip2_ob_out[59]));
Q_ASSIGN U188 ( .B(kme_cceip2_ob_out_post[58]), .A(kme_cceip2_ob_out[58]));
Q_ASSIGN U189 ( .B(kme_cceip2_ob_out_post[57]), .A(kme_cceip2_ob_out[57]));
Q_ASSIGN U190 ( .B(kme_cceip2_ob_out_post[56]), .A(kme_cceip2_ob_out[56]));
Q_ASSIGN U191 ( .B(kme_cceip2_ob_out_post[55]), .A(kme_cceip2_ob_out[55]));
Q_ASSIGN U192 ( .B(kme_cceip2_ob_out_post[54]), .A(kme_cceip2_ob_out[54]));
Q_ASSIGN U193 ( .B(kme_cceip2_ob_out_post[53]), .A(kme_cceip2_ob_out[53]));
Q_ASSIGN U194 ( .B(kme_cceip2_ob_out_post[52]), .A(kme_cceip2_ob_out[52]));
Q_ASSIGN U195 ( .B(kme_cceip2_ob_out_post[51]), .A(kme_cceip2_ob_out[51]));
Q_ASSIGN U196 ( .B(kme_cceip2_ob_out_post[50]), .A(kme_cceip2_ob_out[50]));
Q_ASSIGN U197 ( .B(kme_cceip2_ob_out_post[49]), .A(kme_cceip2_ob_out[49]));
Q_ASSIGN U198 ( .B(kme_cceip2_ob_out_post[48]), .A(kme_cceip2_ob_out[48]));
Q_ASSIGN U199 ( .B(kme_cceip2_ob_out_post[47]), .A(kme_cceip2_ob_out[47]));
Q_ASSIGN U200 ( .B(kme_cceip2_ob_out_post[46]), .A(kme_cceip2_ob_out[46]));
Q_ASSIGN U201 ( .B(kme_cceip2_ob_out_post[45]), .A(kme_cceip2_ob_out[45]));
Q_ASSIGN U202 ( .B(kme_cceip2_ob_out_post[44]), .A(kme_cceip2_ob_out[44]));
Q_ASSIGN U203 ( .B(kme_cceip2_ob_out_post[43]), .A(kme_cceip2_ob_out[43]));
Q_ASSIGN U204 ( .B(kme_cceip2_ob_out_post[42]), .A(kme_cceip2_ob_out[42]));
Q_ASSIGN U205 ( .B(kme_cceip2_ob_out_post[41]), .A(kme_cceip2_ob_out[41]));
Q_ASSIGN U206 ( .B(kme_cceip2_ob_out_post[40]), .A(kme_cceip2_ob_out[40]));
Q_ASSIGN U207 ( .B(kme_cceip2_ob_out_post[39]), .A(kme_cceip2_ob_out[39]));
Q_ASSIGN U208 ( .B(kme_cceip2_ob_out_post[38]), .A(kme_cceip2_ob_out[38]));
Q_ASSIGN U209 ( .B(kme_cceip2_ob_out_post[37]), .A(kme_cceip2_ob_out[37]));
Q_ASSIGN U210 ( .B(kme_cceip2_ob_out_post[36]), .A(kme_cceip2_ob_out[36]));
Q_ASSIGN U211 ( .B(kme_cceip2_ob_out_post[35]), .A(kme_cceip2_ob_out[35]));
Q_ASSIGN U212 ( .B(kme_cceip2_ob_out_post[34]), .A(kme_cceip2_ob_out[34]));
Q_ASSIGN U213 ( .B(kme_cceip2_ob_out_post[33]), .A(kme_cceip2_ob_out[33]));
Q_ASSIGN U214 ( .B(kme_cceip2_ob_out_post[32]), .A(kme_cceip2_ob_out[32]));
Q_ASSIGN U215 ( .B(kme_cceip2_ob_out_post[31]), .A(kme_cceip2_ob_out[31]));
Q_ASSIGN U216 ( .B(kme_cceip2_ob_out_post[30]), .A(kme_cceip2_ob_out[30]));
Q_ASSIGN U217 ( .B(kme_cceip2_ob_out_post[29]), .A(kme_cceip2_ob_out[29]));
Q_ASSIGN U218 ( .B(kme_cceip2_ob_out_post[28]), .A(kme_cceip2_ob_out[28]));
Q_ASSIGN U219 ( .B(kme_cceip2_ob_out_post[27]), .A(kme_cceip2_ob_out[27]));
Q_ASSIGN U220 ( .B(kme_cceip2_ob_out_post[26]), .A(kme_cceip2_ob_out[26]));
Q_ASSIGN U221 ( .B(kme_cceip2_ob_out_post[25]), .A(kme_cceip2_ob_out[25]));
Q_ASSIGN U222 ( .B(kme_cceip2_ob_out_post[24]), .A(kme_cceip2_ob_out[24]));
Q_ASSIGN U223 ( .B(kme_cceip2_ob_out_post[23]), .A(kme_cceip2_ob_out[23]));
Q_ASSIGN U224 ( .B(kme_cceip2_ob_out_post[22]), .A(kme_cceip2_ob_out[22]));
Q_ASSIGN U225 ( .B(kme_cceip2_ob_out_post[21]), .A(kme_cceip2_ob_out[21]));
Q_ASSIGN U226 ( .B(kme_cceip2_ob_out_post[20]), .A(kme_cceip2_ob_out[20]));
Q_ASSIGN U227 ( .B(kme_cceip2_ob_out_post[19]), .A(kme_cceip2_ob_out[19]));
Q_ASSIGN U228 ( .B(kme_cceip2_ob_out_post[18]), .A(kme_cceip2_ob_out[18]));
Q_ASSIGN U229 ( .B(kme_cceip2_ob_out_post[17]), .A(kme_cceip2_ob_out[17]));
Q_ASSIGN U230 ( .B(kme_cceip2_ob_out_post[16]), .A(kme_cceip2_ob_out[16]));
Q_ASSIGN U231 ( .B(kme_cceip2_ob_out_post[15]), .A(kme_cceip2_ob_out[15]));
Q_ASSIGN U232 ( .B(kme_cceip2_ob_out_post[14]), .A(kme_cceip2_ob_out[14]));
Q_ASSIGN U233 ( .B(kme_cceip2_ob_out_post[13]), .A(kme_cceip2_ob_out[13]));
Q_ASSIGN U234 ( .B(kme_cceip2_ob_out_post[12]), .A(kme_cceip2_ob_out[12]));
Q_ASSIGN U235 ( .B(kme_cceip2_ob_out_post[11]), .A(kme_cceip2_ob_out[11]));
Q_ASSIGN U236 ( .B(kme_cceip2_ob_out_post[10]), .A(kme_cceip2_ob_out[10]));
Q_ASSIGN U237 ( .B(kme_cceip2_ob_out_post[9]), .A(kme_cceip2_ob_out[9]));
Q_ASSIGN U238 ( .B(kme_cceip2_ob_out_post[8]), .A(kme_cceip2_ob_out[8]));
Q_ASSIGN U239 ( .B(kme_cceip2_ob_out_post[7]), .A(kme_cceip2_ob_out[7]));
Q_ASSIGN U240 ( .B(kme_cceip2_ob_out_post[6]), .A(kme_cceip2_ob_out[6]));
Q_ASSIGN U241 ( .B(kme_cceip2_ob_out_post[5]), .A(kme_cceip2_ob_out[5]));
Q_ASSIGN U242 ( .B(kme_cceip2_ob_out_post[4]), .A(kme_cceip2_ob_out[4]));
Q_ASSIGN U243 ( .B(kme_cceip2_ob_out_post[3]), .A(kme_cceip2_ob_out[3]));
Q_ASSIGN U244 ( .B(kme_cceip2_ob_out_post[2]), .A(kme_cceip2_ob_out[2]));
Q_ASSIGN U245 ( .B(kme_cceip2_ob_out_post[1]), .A(kme_cceip2_ob_out[1]));
Q_ASSIGN U246 ( .B(kme_cceip2_ob_out_post[0]), .A(kme_cceip2_ob_out[0]));
Q_ASSIGN U247 ( .B(kme_cceip3_ob_out_post[81]), .A(kme_cceip3_ob_out[81]));
Q_ASSIGN U248 ( .B(kme_cceip3_ob_out_post[80]), .A(kme_cceip3_ob_out[80]));
Q_ASSIGN U249 ( .B(kme_cceip3_ob_out_post[79]), .A(kme_cceip3_ob_out[79]));
Q_ASSIGN U250 ( .B(kme_cceip3_ob_out_post[78]), .A(kme_cceip3_ob_out[78]));
Q_ASSIGN U251 ( .B(kme_cceip3_ob_out_post[77]), .A(kme_cceip3_ob_out[77]));
Q_ASSIGN U252 ( .B(kme_cceip3_ob_out_post[76]), .A(kme_cceip3_ob_out[76]));
Q_ASSIGN U253 ( .B(kme_cceip3_ob_out_post[75]), .A(kme_cceip3_ob_out[75]));
Q_ASSIGN U254 ( .B(kme_cceip3_ob_out_post[74]), .A(kme_cceip3_ob_out[74]));
Q_ASSIGN U255 ( .B(kme_cceip3_ob_out_post[73]), .A(kme_cceip3_ob_out[73]));
Q_ASSIGN U256 ( .B(kme_cceip3_ob_out_post[72]), .A(kme_cceip3_ob_out[72]));
Q_ASSIGN U257 ( .B(kme_cceip3_ob_out_post[71]), .A(kme_cceip3_ob_out[71]));
Q_ASSIGN U258 ( .B(kme_cceip3_ob_out_post[70]), .A(kme_cceip3_ob_out[70]));
Q_ASSIGN U259 ( .B(kme_cceip3_ob_out_post[69]), .A(kme_cceip3_ob_out[69]));
Q_ASSIGN U260 ( .B(kme_cceip3_ob_out_post[68]), .A(kme_cceip3_ob_out[68]));
Q_ASSIGN U261 ( .B(kme_cceip3_ob_out_post[67]), .A(kme_cceip3_ob_out[67]));
Q_ASSIGN U262 ( .B(kme_cceip3_ob_out_post[66]), .A(kme_cceip3_ob_out[66]));
Q_ASSIGN U263 ( .B(kme_cceip3_ob_out_post[65]), .A(kme_cceip3_ob_out[65]));
Q_ASSIGN U264 ( .B(kme_cceip3_ob_out_post[64]), .A(kme_cceip3_ob_out[64]));
Q_ASSIGN U265 ( .B(kme_cceip3_ob_out_post[63]), .A(kme_cceip3_ob_out[63]));
Q_ASSIGN U266 ( .B(kme_cceip3_ob_out_post[62]), .A(kme_cceip3_ob_out[62]));
Q_ASSIGN U267 ( .B(kme_cceip3_ob_out_post[61]), .A(kme_cceip3_ob_out[61]));
Q_ASSIGN U268 ( .B(kme_cceip3_ob_out_post[60]), .A(kme_cceip3_ob_out[60]));
Q_ASSIGN U269 ( .B(kme_cceip3_ob_out_post[59]), .A(kme_cceip3_ob_out[59]));
Q_ASSIGN U270 ( .B(kme_cceip3_ob_out_post[58]), .A(kme_cceip3_ob_out[58]));
Q_ASSIGN U271 ( .B(kme_cceip3_ob_out_post[57]), .A(kme_cceip3_ob_out[57]));
Q_ASSIGN U272 ( .B(kme_cceip3_ob_out_post[56]), .A(kme_cceip3_ob_out[56]));
Q_ASSIGN U273 ( .B(kme_cceip3_ob_out_post[55]), .A(kme_cceip3_ob_out[55]));
Q_ASSIGN U274 ( .B(kme_cceip3_ob_out_post[54]), .A(kme_cceip3_ob_out[54]));
Q_ASSIGN U275 ( .B(kme_cceip3_ob_out_post[53]), .A(kme_cceip3_ob_out[53]));
Q_ASSIGN U276 ( .B(kme_cceip3_ob_out_post[52]), .A(kme_cceip3_ob_out[52]));
Q_ASSIGN U277 ( .B(kme_cceip3_ob_out_post[51]), .A(kme_cceip3_ob_out[51]));
Q_ASSIGN U278 ( .B(kme_cceip3_ob_out_post[50]), .A(kme_cceip3_ob_out[50]));
Q_ASSIGN U279 ( .B(kme_cceip3_ob_out_post[49]), .A(kme_cceip3_ob_out[49]));
Q_ASSIGN U280 ( .B(kme_cceip3_ob_out_post[48]), .A(kme_cceip3_ob_out[48]));
Q_ASSIGN U281 ( .B(kme_cceip3_ob_out_post[47]), .A(kme_cceip3_ob_out[47]));
Q_ASSIGN U282 ( .B(kme_cceip3_ob_out_post[46]), .A(kme_cceip3_ob_out[46]));
Q_ASSIGN U283 ( .B(kme_cceip3_ob_out_post[45]), .A(kme_cceip3_ob_out[45]));
Q_ASSIGN U284 ( .B(kme_cceip3_ob_out_post[44]), .A(kme_cceip3_ob_out[44]));
Q_ASSIGN U285 ( .B(kme_cceip3_ob_out_post[43]), .A(kme_cceip3_ob_out[43]));
Q_ASSIGN U286 ( .B(kme_cceip3_ob_out_post[42]), .A(kme_cceip3_ob_out[42]));
Q_ASSIGN U287 ( .B(kme_cceip3_ob_out_post[41]), .A(kme_cceip3_ob_out[41]));
Q_ASSIGN U288 ( .B(kme_cceip3_ob_out_post[40]), .A(kme_cceip3_ob_out[40]));
Q_ASSIGN U289 ( .B(kme_cceip3_ob_out_post[39]), .A(kme_cceip3_ob_out[39]));
Q_ASSIGN U290 ( .B(kme_cceip3_ob_out_post[38]), .A(kme_cceip3_ob_out[38]));
Q_ASSIGN U291 ( .B(kme_cceip3_ob_out_post[37]), .A(kme_cceip3_ob_out[37]));
Q_ASSIGN U292 ( .B(kme_cceip3_ob_out_post[36]), .A(kme_cceip3_ob_out[36]));
Q_ASSIGN U293 ( .B(kme_cceip3_ob_out_post[35]), .A(kme_cceip3_ob_out[35]));
Q_ASSIGN U294 ( .B(kme_cceip3_ob_out_post[34]), .A(kme_cceip3_ob_out[34]));
Q_ASSIGN U295 ( .B(kme_cceip3_ob_out_post[33]), .A(kme_cceip3_ob_out[33]));
Q_ASSIGN U296 ( .B(kme_cceip3_ob_out_post[32]), .A(kme_cceip3_ob_out[32]));
Q_ASSIGN U297 ( .B(kme_cceip3_ob_out_post[31]), .A(kme_cceip3_ob_out[31]));
Q_ASSIGN U298 ( .B(kme_cceip3_ob_out_post[30]), .A(kme_cceip3_ob_out[30]));
Q_ASSIGN U299 ( .B(kme_cceip3_ob_out_post[29]), .A(kme_cceip3_ob_out[29]));
Q_ASSIGN U300 ( .B(kme_cceip3_ob_out_post[28]), .A(kme_cceip3_ob_out[28]));
Q_ASSIGN U301 ( .B(kme_cceip3_ob_out_post[27]), .A(kme_cceip3_ob_out[27]));
Q_ASSIGN U302 ( .B(kme_cceip3_ob_out_post[26]), .A(kme_cceip3_ob_out[26]));
Q_ASSIGN U303 ( .B(kme_cceip3_ob_out_post[25]), .A(kme_cceip3_ob_out[25]));
Q_ASSIGN U304 ( .B(kme_cceip3_ob_out_post[24]), .A(kme_cceip3_ob_out[24]));
Q_ASSIGN U305 ( .B(kme_cceip3_ob_out_post[23]), .A(kme_cceip3_ob_out[23]));
Q_ASSIGN U306 ( .B(kme_cceip3_ob_out_post[22]), .A(kme_cceip3_ob_out[22]));
Q_ASSIGN U307 ( .B(kme_cceip3_ob_out_post[21]), .A(kme_cceip3_ob_out[21]));
Q_ASSIGN U308 ( .B(kme_cceip3_ob_out_post[20]), .A(kme_cceip3_ob_out[20]));
Q_ASSIGN U309 ( .B(kme_cceip3_ob_out_post[19]), .A(kme_cceip3_ob_out[19]));
Q_ASSIGN U310 ( .B(kme_cceip3_ob_out_post[18]), .A(kme_cceip3_ob_out[18]));
Q_ASSIGN U311 ( .B(kme_cceip3_ob_out_post[17]), .A(kme_cceip3_ob_out[17]));
Q_ASSIGN U312 ( .B(kme_cceip3_ob_out_post[16]), .A(kme_cceip3_ob_out[16]));
Q_ASSIGN U313 ( .B(kme_cceip3_ob_out_post[15]), .A(kme_cceip3_ob_out[15]));
Q_ASSIGN U314 ( .B(kme_cceip3_ob_out_post[14]), .A(kme_cceip3_ob_out[14]));
Q_ASSIGN U315 ( .B(kme_cceip3_ob_out_post[13]), .A(kme_cceip3_ob_out[13]));
Q_ASSIGN U316 ( .B(kme_cceip3_ob_out_post[12]), .A(kme_cceip3_ob_out[12]));
Q_ASSIGN U317 ( .B(kme_cceip3_ob_out_post[11]), .A(kme_cceip3_ob_out[11]));
Q_ASSIGN U318 ( .B(kme_cceip3_ob_out_post[10]), .A(kme_cceip3_ob_out[10]));
Q_ASSIGN U319 ( .B(kme_cceip3_ob_out_post[9]), .A(kme_cceip3_ob_out[9]));
Q_ASSIGN U320 ( .B(kme_cceip3_ob_out_post[8]), .A(kme_cceip3_ob_out[8]));
Q_ASSIGN U321 ( .B(kme_cceip3_ob_out_post[7]), .A(kme_cceip3_ob_out[7]));
Q_ASSIGN U322 ( .B(kme_cceip3_ob_out_post[6]), .A(kme_cceip3_ob_out[6]));
Q_ASSIGN U323 ( .B(kme_cceip3_ob_out_post[5]), .A(kme_cceip3_ob_out[5]));
Q_ASSIGN U324 ( .B(kme_cceip3_ob_out_post[4]), .A(kme_cceip3_ob_out[4]));
Q_ASSIGN U325 ( .B(kme_cceip3_ob_out_post[3]), .A(kme_cceip3_ob_out[3]));
Q_ASSIGN U326 ( .B(kme_cceip3_ob_out_post[2]), .A(kme_cceip3_ob_out[2]));
Q_ASSIGN U327 ( .B(kme_cceip3_ob_out_post[1]), .A(kme_cceip3_ob_out[1]));
Q_ASSIGN U328 ( .B(kme_cceip3_ob_out_post[0]), .A(kme_cceip3_ob_out[0]));
Q_ASSIGN U329 ( .B(kme_cddip0_ob_out_post[81]), .A(kme_cddip0_ob_out[81]));
Q_ASSIGN U330 ( .B(kme_cddip0_ob_out_post[80]), .A(kme_cddip0_ob_out[80]));
Q_ASSIGN U331 ( .B(kme_cddip0_ob_out_post[79]), .A(kme_cddip0_ob_out[79]));
Q_ASSIGN U332 ( .B(kme_cddip0_ob_out_post[78]), .A(kme_cddip0_ob_out[78]));
Q_ASSIGN U333 ( .B(kme_cddip0_ob_out_post[77]), .A(kme_cddip0_ob_out[77]));
Q_ASSIGN U334 ( .B(kme_cddip0_ob_out_post[76]), .A(kme_cddip0_ob_out[76]));
Q_ASSIGN U335 ( .B(kme_cddip0_ob_out_post[75]), .A(kme_cddip0_ob_out[75]));
Q_ASSIGN U336 ( .B(kme_cddip0_ob_out_post[74]), .A(kme_cddip0_ob_out[74]));
Q_ASSIGN U337 ( .B(kme_cddip0_ob_out_post[73]), .A(kme_cddip0_ob_out[73]));
Q_ASSIGN U338 ( .B(kme_cddip0_ob_out_post[72]), .A(kme_cddip0_ob_out[72]));
Q_ASSIGN U339 ( .B(kme_cddip0_ob_out_post[71]), .A(kme_cddip0_ob_out[71]));
Q_ASSIGN U340 ( .B(kme_cddip0_ob_out_post[70]), .A(kme_cddip0_ob_out[70]));
Q_ASSIGN U341 ( .B(kme_cddip0_ob_out_post[69]), .A(kme_cddip0_ob_out[69]));
Q_ASSIGN U342 ( .B(kme_cddip0_ob_out_post[68]), .A(kme_cddip0_ob_out[68]));
Q_ASSIGN U343 ( .B(kme_cddip0_ob_out_post[67]), .A(kme_cddip0_ob_out[67]));
Q_ASSIGN U344 ( .B(kme_cddip0_ob_out_post[66]), .A(kme_cddip0_ob_out[66]));
Q_ASSIGN U345 ( .B(kme_cddip0_ob_out_post[65]), .A(kme_cddip0_ob_out[65]));
Q_ASSIGN U346 ( .B(kme_cddip0_ob_out_post[64]), .A(kme_cddip0_ob_out[64]));
Q_ASSIGN U347 ( .B(kme_cddip0_ob_out_post[63]), .A(kme_cddip0_ob_out[63]));
Q_ASSIGN U348 ( .B(kme_cddip0_ob_out_post[62]), .A(kme_cddip0_ob_out[62]));
Q_ASSIGN U349 ( .B(kme_cddip0_ob_out_post[61]), .A(kme_cddip0_ob_out[61]));
Q_ASSIGN U350 ( .B(kme_cddip0_ob_out_post[60]), .A(kme_cddip0_ob_out[60]));
Q_ASSIGN U351 ( .B(kme_cddip0_ob_out_post[59]), .A(kme_cddip0_ob_out[59]));
Q_ASSIGN U352 ( .B(kme_cddip0_ob_out_post[58]), .A(kme_cddip0_ob_out[58]));
Q_ASSIGN U353 ( .B(kme_cddip0_ob_out_post[57]), .A(kme_cddip0_ob_out[57]));
Q_ASSIGN U354 ( .B(kme_cddip0_ob_out_post[56]), .A(kme_cddip0_ob_out[56]));
Q_ASSIGN U355 ( .B(kme_cddip0_ob_out_post[55]), .A(kme_cddip0_ob_out[55]));
Q_ASSIGN U356 ( .B(kme_cddip0_ob_out_post[54]), .A(kme_cddip0_ob_out[54]));
Q_ASSIGN U357 ( .B(kme_cddip0_ob_out_post[53]), .A(kme_cddip0_ob_out[53]));
Q_ASSIGN U358 ( .B(kme_cddip0_ob_out_post[52]), .A(kme_cddip0_ob_out[52]));
Q_ASSIGN U359 ( .B(kme_cddip0_ob_out_post[51]), .A(kme_cddip0_ob_out[51]));
Q_ASSIGN U360 ( .B(kme_cddip0_ob_out_post[50]), .A(kme_cddip0_ob_out[50]));
Q_ASSIGN U361 ( .B(kme_cddip0_ob_out_post[49]), .A(kme_cddip0_ob_out[49]));
Q_ASSIGN U362 ( .B(kme_cddip0_ob_out_post[48]), .A(kme_cddip0_ob_out[48]));
Q_ASSIGN U363 ( .B(kme_cddip0_ob_out_post[47]), .A(kme_cddip0_ob_out[47]));
Q_ASSIGN U364 ( .B(kme_cddip0_ob_out_post[46]), .A(kme_cddip0_ob_out[46]));
Q_ASSIGN U365 ( .B(kme_cddip0_ob_out_post[45]), .A(kme_cddip0_ob_out[45]));
Q_ASSIGN U366 ( .B(kme_cddip0_ob_out_post[44]), .A(kme_cddip0_ob_out[44]));
Q_ASSIGN U367 ( .B(kme_cddip0_ob_out_post[43]), .A(kme_cddip0_ob_out[43]));
Q_ASSIGN U368 ( .B(kme_cddip0_ob_out_post[42]), .A(kme_cddip0_ob_out[42]));
Q_ASSIGN U369 ( .B(kme_cddip0_ob_out_post[41]), .A(kme_cddip0_ob_out[41]));
Q_ASSIGN U370 ( .B(kme_cddip0_ob_out_post[40]), .A(kme_cddip0_ob_out[40]));
Q_ASSIGN U371 ( .B(kme_cddip0_ob_out_post[39]), .A(kme_cddip0_ob_out[39]));
Q_ASSIGN U372 ( .B(kme_cddip0_ob_out_post[38]), .A(kme_cddip0_ob_out[38]));
Q_ASSIGN U373 ( .B(kme_cddip0_ob_out_post[37]), .A(kme_cddip0_ob_out[37]));
Q_ASSIGN U374 ( .B(kme_cddip0_ob_out_post[36]), .A(kme_cddip0_ob_out[36]));
Q_ASSIGN U375 ( .B(kme_cddip0_ob_out_post[35]), .A(kme_cddip0_ob_out[35]));
Q_ASSIGN U376 ( .B(kme_cddip0_ob_out_post[34]), .A(kme_cddip0_ob_out[34]));
Q_ASSIGN U377 ( .B(kme_cddip0_ob_out_post[33]), .A(kme_cddip0_ob_out[33]));
Q_ASSIGN U378 ( .B(kme_cddip0_ob_out_post[32]), .A(kme_cddip0_ob_out[32]));
Q_ASSIGN U379 ( .B(kme_cddip0_ob_out_post[31]), .A(kme_cddip0_ob_out[31]));
Q_ASSIGN U380 ( .B(kme_cddip0_ob_out_post[30]), .A(kme_cddip0_ob_out[30]));
Q_ASSIGN U381 ( .B(kme_cddip0_ob_out_post[29]), .A(kme_cddip0_ob_out[29]));
Q_ASSIGN U382 ( .B(kme_cddip0_ob_out_post[28]), .A(kme_cddip0_ob_out[28]));
Q_ASSIGN U383 ( .B(kme_cddip0_ob_out_post[27]), .A(kme_cddip0_ob_out[27]));
Q_ASSIGN U384 ( .B(kme_cddip0_ob_out_post[26]), .A(kme_cddip0_ob_out[26]));
Q_ASSIGN U385 ( .B(kme_cddip0_ob_out_post[25]), .A(kme_cddip0_ob_out[25]));
Q_ASSIGN U386 ( .B(kme_cddip0_ob_out_post[24]), .A(kme_cddip0_ob_out[24]));
Q_ASSIGN U387 ( .B(kme_cddip0_ob_out_post[23]), .A(kme_cddip0_ob_out[23]));
Q_ASSIGN U388 ( .B(kme_cddip0_ob_out_post[22]), .A(kme_cddip0_ob_out[22]));
Q_ASSIGN U389 ( .B(kme_cddip0_ob_out_post[21]), .A(kme_cddip0_ob_out[21]));
Q_ASSIGN U390 ( .B(kme_cddip0_ob_out_post[20]), .A(kme_cddip0_ob_out[20]));
Q_ASSIGN U391 ( .B(kme_cddip0_ob_out_post[19]), .A(kme_cddip0_ob_out[19]));
Q_ASSIGN U392 ( .B(kme_cddip0_ob_out_post[18]), .A(kme_cddip0_ob_out[18]));
Q_ASSIGN U393 ( .B(kme_cddip0_ob_out_post[17]), .A(kme_cddip0_ob_out[17]));
Q_ASSIGN U394 ( .B(kme_cddip0_ob_out_post[16]), .A(kme_cddip0_ob_out[16]));
Q_ASSIGN U395 ( .B(kme_cddip0_ob_out_post[15]), .A(kme_cddip0_ob_out[15]));
Q_ASSIGN U396 ( .B(kme_cddip0_ob_out_post[14]), .A(kme_cddip0_ob_out[14]));
Q_ASSIGN U397 ( .B(kme_cddip0_ob_out_post[13]), .A(kme_cddip0_ob_out[13]));
Q_ASSIGN U398 ( .B(kme_cddip0_ob_out_post[12]), .A(kme_cddip0_ob_out[12]));
Q_ASSIGN U399 ( .B(kme_cddip0_ob_out_post[11]), .A(kme_cddip0_ob_out[11]));
Q_ASSIGN U400 ( .B(kme_cddip0_ob_out_post[10]), .A(kme_cddip0_ob_out[10]));
Q_ASSIGN U401 ( .B(kme_cddip0_ob_out_post[9]), .A(kme_cddip0_ob_out[9]));
Q_ASSIGN U402 ( .B(kme_cddip0_ob_out_post[8]), .A(kme_cddip0_ob_out[8]));
Q_ASSIGN U403 ( .B(kme_cddip0_ob_out_post[7]), .A(kme_cddip0_ob_out[7]));
Q_ASSIGN U404 ( .B(kme_cddip0_ob_out_post[6]), .A(kme_cddip0_ob_out[6]));
Q_ASSIGN U405 ( .B(kme_cddip0_ob_out_post[5]), .A(kme_cddip0_ob_out[5]));
Q_ASSIGN U406 ( .B(kme_cddip0_ob_out_post[4]), .A(kme_cddip0_ob_out[4]));
Q_ASSIGN U407 ( .B(kme_cddip0_ob_out_post[3]), .A(kme_cddip0_ob_out[3]));
Q_ASSIGN U408 ( .B(kme_cddip0_ob_out_post[2]), .A(kme_cddip0_ob_out[2]));
Q_ASSIGN U409 ( .B(kme_cddip0_ob_out_post[1]), .A(kme_cddip0_ob_out[1]));
Q_ASSIGN U410 ( .B(kme_cddip0_ob_out_post[0]), .A(kme_cddip0_ob_out[0]));
Q_ASSIGN U411 ( .B(kme_cddip1_ob_out_post[81]), .A(kme_cddip1_ob_out[81]));
Q_ASSIGN U412 ( .B(kme_cddip1_ob_out_post[80]), .A(kme_cddip1_ob_out[80]));
Q_ASSIGN U413 ( .B(kme_cddip1_ob_out_post[79]), .A(kme_cddip1_ob_out[79]));
Q_ASSIGN U414 ( .B(kme_cddip1_ob_out_post[78]), .A(kme_cddip1_ob_out[78]));
Q_ASSIGN U415 ( .B(kme_cddip1_ob_out_post[77]), .A(kme_cddip1_ob_out[77]));
Q_ASSIGN U416 ( .B(kme_cddip1_ob_out_post[76]), .A(kme_cddip1_ob_out[76]));
Q_ASSIGN U417 ( .B(kme_cddip1_ob_out_post[75]), .A(kme_cddip1_ob_out[75]));
Q_ASSIGN U418 ( .B(kme_cddip1_ob_out_post[74]), .A(kme_cddip1_ob_out[74]));
Q_ASSIGN U419 ( .B(kme_cddip1_ob_out_post[73]), .A(kme_cddip1_ob_out[73]));
Q_ASSIGN U420 ( .B(kme_cddip1_ob_out_post[72]), .A(kme_cddip1_ob_out[72]));
Q_ASSIGN U421 ( .B(kme_cddip1_ob_out_post[71]), .A(kme_cddip1_ob_out[71]));
Q_ASSIGN U422 ( .B(kme_cddip1_ob_out_post[70]), .A(kme_cddip1_ob_out[70]));
Q_ASSIGN U423 ( .B(kme_cddip1_ob_out_post[69]), .A(kme_cddip1_ob_out[69]));
Q_ASSIGN U424 ( .B(kme_cddip1_ob_out_post[68]), .A(kme_cddip1_ob_out[68]));
Q_ASSIGN U425 ( .B(kme_cddip1_ob_out_post[67]), .A(kme_cddip1_ob_out[67]));
Q_ASSIGN U426 ( .B(kme_cddip1_ob_out_post[66]), .A(kme_cddip1_ob_out[66]));
Q_ASSIGN U427 ( .B(kme_cddip1_ob_out_post[65]), .A(kme_cddip1_ob_out[65]));
Q_ASSIGN U428 ( .B(kme_cddip1_ob_out_post[64]), .A(kme_cddip1_ob_out[64]));
Q_ASSIGN U429 ( .B(kme_cddip1_ob_out_post[63]), .A(kme_cddip1_ob_out[63]));
Q_ASSIGN U430 ( .B(kme_cddip1_ob_out_post[62]), .A(kme_cddip1_ob_out[62]));
Q_ASSIGN U431 ( .B(kme_cddip1_ob_out_post[61]), .A(kme_cddip1_ob_out[61]));
Q_ASSIGN U432 ( .B(kme_cddip1_ob_out_post[60]), .A(kme_cddip1_ob_out[60]));
Q_ASSIGN U433 ( .B(kme_cddip1_ob_out_post[59]), .A(kme_cddip1_ob_out[59]));
Q_ASSIGN U434 ( .B(kme_cddip1_ob_out_post[58]), .A(kme_cddip1_ob_out[58]));
Q_ASSIGN U435 ( .B(kme_cddip1_ob_out_post[57]), .A(kme_cddip1_ob_out[57]));
Q_ASSIGN U436 ( .B(kme_cddip1_ob_out_post[56]), .A(kme_cddip1_ob_out[56]));
Q_ASSIGN U437 ( .B(kme_cddip1_ob_out_post[55]), .A(kme_cddip1_ob_out[55]));
Q_ASSIGN U438 ( .B(kme_cddip1_ob_out_post[54]), .A(kme_cddip1_ob_out[54]));
Q_ASSIGN U439 ( .B(kme_cddip1_ob_out_post[53]), .A(kme_cddip1_ob_out[53]));
Q_ASSIGN U440 ( .B(kme_cddip1_ob_out_post[52]), .A(kme_cddip1_ob_out[52]));
Q_ASSIGN U441 ( .B(kme_cddip1_ob_out_post[51]), .A(kme_cddip1_ob_out[51]));
Q_ASSIGN U442 ( .B(kme_cddip1_ob_out_post[50]), .A(kme_cddip1_ob_out[50]));
Q_ASSIGN U443 ( .B(kme_cddip1_ob_out_post[49]), .A(kme_cddip1_ob_out[49]));
Q_ASSIGN U444 ( .B(kme_cddip1_ob_out_post[48]), .A(kme_cddip1_ob_out[48]));
Q_ASSIGN U445 ( .B(kme_cddip1_ob_out_post[47]), .A(kme_cddip1_ob_out[47]));
Q_ASSIGN U446 ( .B(kme_cddip1_ob_out_post[46]), .A(kme_cddip1_ob_out[46]));
Q_ASSIGN U447 ( .B(kme_cddip1_ob_out_post[45]), .A(kme_cddip1_ob_out[45]));
Q_ASSIGN U448 ( .B(kme_cddip1_ob_out_post[44]), .A(kme_cddip1_ob_out[44]));
Q_ASSIGN U449 ( .B(kme_cddip1_ob_out_post[43]), .A(kme_cddip1_ob_out[43]));
Q_ASSIGN U450 ( .B(kme_cddip1_ob_out_post[42]), .A(kme_cddip1_ob_out[42]));
Q_ASSIGN U451 ( .B(kme_cddip1_ob_out_post[41]), .A(kme_cddip1_ob_out[41]));
Q_ASSIGN U452 ( .B(kme_cddip1_ob_out_post[40]), .A(kme_cddip1_ob_out[40]));
Q_ASSIGN U453 ( .B(kme_cddip1_ob_out_post[39]), .A(kme_cddip1_ob_out[39]));
Q_ASSIGN U454 ( .B(kme_cddip1_ob_out_post[38]), .A(kme_cddip1_ob_out[38]));
Q_ASSIGN U455 ( .B(kme_cddip1_ob_out_post[37]), .A(kme_cddip1_ob_out[37]));
Q_ASSIGN U456 ( .B(kme_cddip1_ob_out_post[36]), .A(kme_cddip1_ob_out[36]));
Q_ASSIGN U457 ( .B(kme_cddip1_ob_out_post[35]), .A(kme_cddip1_ob_out[35]));
Q_ASSIGN U458 ( .B(kme_cddip1_ob_out_post[34]), .A(kme_cddip1_ob_out[34]));
Q_ASSIGN U459 ( .B(kme_cddip1_ob_out_post[33]), .A(kme_cddip1_ob_out[33]));
Q_ASSIGN U460 ( .B(kme_cddip1_ob_out_post[32]), .A(kme_cddip1_ob_out[32]));
Q_ASSIGN U461 ( .B(kme_cddip1_ob_out_post[31]), .A(kme_cddip1_ob_out[31]));
Q_ASSIGN U462 ( .B(kme_cddip1_ob_out_post[30]), .A(kme_cddip1_ob_out[30]));
Q_ASSIGN U463 ( .B(kme_cddip1_ob_out_post[29]), .A(kme_cddip1_ob_out[29]));
Q_ASSIGN U464 ( .B(kme_cddip1_ob_out_post[28]), .A(kme_cddip1_ob_out[28]));
Q_ASSIGN U465 ( .B(kme_cddip1_ob_out_post[27]), .A(kme_cddip1_ob_out[27]));
Q_ASSIGN U466 ( .B(kme_cddip1_ob_out_post[26]), .A(kme_cddip1_ob_out[26]));
Q_ASSIGN U467 ( .B(kme_cddip1_ob_out_post[25]), .A(kme_cddip1_ob_out[25]));
Q_ASSIGN U468 ( .B(kme_cddip1_ob_out_post[24]), .A(kme_cddip1_ob_out[24]));
Q_ASSIGN U469 ( .B(kme_cddip1_ob_out_post[23]), .A(kme_cddip1_ob_out[23]));
Q_ASSIGN U470 ( .B(kme_cddip1_ob_out_post[22]), .A(kme_cddip1_ob_out[22]));
Q_ASSIGN U471 ( .B(kme_cddip1_ob_out_post[21]), .A(kme_cddip1_ob_out[21]));
Q_ASSIGN U472 ( .B(kme_cddip1_ob_out_post[20]), .A(kme_cddip1_ob_out[20]));
Q_ASSIGN U473 ( .B(kme_cddip1_ob_out_post[19]), .A(kme_cddip1_ob_out[19]));
Q_ASSIGN U474 ( .B(kme_cddip1_ob_out_post[18]), .A(kme_cddip1_ob_out[18]));
Q_ASSIGN U475 ( .B(kme_cddip1_ob_out_post[17]), .A(kme_cddip1_ob_out[17]));
Q_ASSIGN U476 ( .B(kme_cddip1_ob_out_post[16]), .A(kme_cddip1_ob_out[16]));
Q_ASSIGN U477 ( .B(kme_cddip1_ob_out_post[15]), .A(kme_cddip1_ob_out[15]));
Q_ASSIGN U478 ( .B(kme_cddip1_ob_out_post[14]), .A(kme_cddip1_ob_out[14]));
Q_ASSIGN U479 ( .B(kme_cddip1_ob_out_post[13]), .A(kme_cddip1_ob_out[13]));
Q_ASSIGN U480 ( .B(kme_cddip1_ob_out_post[12]), .A(kme_cddip1_ob_out[12]));
Q_ASSIGN U481 ( .B(kme_cddip1_ob_out_post[11]), .A(kme_cddip1_ob_out[11]));
Q_ASSIGN U482 ( .B(kme_cddip1_ob_out_post[10]), .A(kme_cddip1_ob_out[10]));
Q_ASSIGN U483 ( .B(kme_cddip1_ob_out_post[9]), .A(kme_cddip1_ob_out[9]));
Q_ASSIGN U484 ( .B(kme_cddip1_ob_out_post[8]), .A(kme_cddip1_ob_out[8]));
Q_ASSIGN U485 ( .B(kme_cddip1_ob_out_post[7]), .A(kme_cddip1_ob_out[7]));
Q_ASSIGN U486 ( .B(kme_cddip1_ob_out_post[6]), .A(kme_cddip1_ob_out[6]));
Q_ASSIGN U487 ( .B(kme_cddip1_ob_out_post[5]), .A(kme_cddip1_ob_out[5]));
Q_ASSIGN U488 ( .B(kme_cddip1_ob_out_post[4]), .A(kme_cddip1_ob_out[4]));
Q_ASSIGN U489 ( .B(kme_cddip1_ob_out_post[3]), .A(kme_cddip1_ob_out[3]));
Q_ASSIGN U490 ( .B(kme_cddip1_ob_out_post[2]), .A(kme_cddip1_ob_out[2]));
Q_ASSIGN U491 ( .B(kme_cddip1_ob_out_post[1]), .A(kme_cddip1_ob_out[1]));
Q_ASSIGN U492 ( .B(kme_cddip1_ob_out_post[0]), .A(kme_cddip1_ob_out[0]));
Q_ASSIGN U493 ( .B(kme_cddip2_ob_out_post[81]), .A(kme_cddip2_ob_out[81]));
Q_ASSIGN U494 ( .B(kme_cddip2_ob_out_post[80]), .A(kme_cddip2_ob_out[80]));
Q_ASSIGN U495 ( .B(kme_cddip2_ob_out_post[79]), .A(kme_cddip2_ob_out[79]));
Q_ASSIGN U496 ( .B(kme_cddip2_ob_out_post[78]), .A(kme_cddip2_ob_out[78]));
Q_ASSIGN U497 ( .B(kme_cddip2_ob_out_post[77]), .A(kme_cddip2_ob_out[77]));
Q_ASSIGN U498 ( .B(kme_cddip2_ob_out_post[76]), .A(kme_cddip2_ob_out[76]));
Q_ASSIGN U499 ( .B(kme_cddip2_ob_out_post[75]), .A(kme_cddip2_ob_out[75]));
Q_ASSIGN U500 ( .B(kme_cddip2_ob_out_post[74]), .A(kme_cddip2_ob_out[74]));
Q_ASSIGN U501 ( .B(kme_cddip2_ob_out_post[73]), .A(kme_cddip2_ob_out[73]));
Q_ASSIGN U502 ( .B(kme_cddip2_ob_out_post[72]), .A(kme_cddip2_ob_out[72]));
Q_ASSIGN U503 ( .B(kme_cddip2_ob_out_post[71]), .A(kme_cddip2_ob_out[71]));
Q_ASSIGN U504 ( .B(kme_cddip2_ob_out_post[70]), .A(kme_cddip2_ob_out[70]));
Q_ASSIGN U505 ( .B(kme_cddip2_ob_out_post[69]), .A(kme_cddip2_ob_out[69]));
Q_ASSIGN U506 ( .B(kme_cddip2_ob_out_post[68]), .A(kme_cddip2_ob_out[68]));
Q_ASSIGN U507 ( .B(kme_cddip2_ob_out_post[67]), .A(kme_cddip2_ob_out[67]));
Q_ASSIGN U508 ( .B(kme_cddip2_ob_out_post[66]), .A(kme_cddip2_ob_out[66]));
Q_ASSIGN U509 ( .B(kme_cddip2_ob_out_post[65]), .A(kme_cddip2_ob_out[65]));
Q_ASSIGN U510 ( .B(kme_cddip2_ob_out_post[64]), .A(kme_cddip2_ob_out[64]));
Q_ASSIGN U511 ( .B(kme_cddip2_ob_out_post[63]), .A(kme_cddip2_ob_out[63]));
Q_ASSIGN U512 ( .B(kme_cddip2_ob_out_post[62]), .A(kme_cddip2_ob_out[62]));
Q_ASSIGN U513 ( .B(kme_cddip2_ob_out_post[61]), .A(kme_cddip2_ob_out[61]));
Q_ASSIGN U514 ( .B(kme_cddip2_ob_out_post[60]), .A(kme_cddip2_ob_out[60]));
Q_ASSIGN U515 ( .B(kme_cddip2_ob_out_post[59]), .A(kme_cddip2_ob_out[59]));
Q_ASSIGN U516 ( .B(kme_cddip2_ob_out_post[58]), .A(kme_cddip2_ob_out[58]));
Q_ASSIGN U517 ( .B(kme_cddip2_ob_out_post[57]), .A(kme_cddip2_ob_out[57]));
Q_ASSIGN U518 ( .B(kme_cddip2_ob_out_post[56]), .A(kme_cddip2_ob_out[56]));
Q_ASSIGN U519 ( .B(kme_cddip2_ob_out_post[55]), .A(kme_cddip2_ob_out[55]));
Q_ASSIGN U520 ( .B(kme_cddip2_ob_out_post[54]), .A(kme_cddip2_ob_out[54]));
Q_ASSIGN U521 ( .B(kme_cddip2_ob_out_post[53]), .A(kme_cddip2_ob_out[53]));
Q_ASSIGN U522 ( .B(kme_cddip2_ob_out_post[52]), .A(kme_cddip2_ob_out[52]));
Q_ASSIGN U523 ( .B(kme_cddip2_ob_out_post[51]), .A(kme_cddip2_ob_out[51]));
Q_ASSIGN U524 ( .B(kme_cddip2_ob_out_post[50]), .A(kme_cddip2_ob_out[50]));
Q_ASSIGN U525 ( .B(kme_cddip2_ob_out_post[49]), .A(kme_cddip2_ob_out[49]));
Q_ASSIGN U526 ( .B(kme_cddip2_ob_out_post[48]), .A(kme_cddip2_ob_out[48]));
Q_ASSIGN U527 ( .B(kme_cddip2_ob_out_post[47]), .A(kme_cddip2_ob_out[47]));
Q_ASSIGN U528 ( .B(kme_cddip2_ob_out_post[46]), .A(kme_cddip2_ob_out[46]));
Q_ASSIGN U529 ( .B(kme_cddip2_ob_out_post[45]), .A(kme_cddip2_ob_out[45]));
Q_ASSIGN U530 ( .B(kme_cddip2_ob_out_post[44]), .A(kme_cddip2_ob_out[44]));
Q_ASSIGN U531 ( .B(kme_cddip2_ob_out_post[43]), .A(kme_cddip2_ob_out[43]));
Q_ASSIGN U532 ( .B(kme_cddip2_ob_out_post[42]), .A(kme_cddip2_ob_out[42]));
Q_ASSIGN U533 ( .B(kme_cddip2_ob_out_post[41]), .A(kme_cddip2_ob_out[41]));
Q_ASSIGN U534 ( .B(kme_cddip2_ob_out_post[40]), .A(kme_cddip2_ob_out[40]));
Q_ASSIGN U535 ( .B(kme_cddip2_ob_out_post[39]), .A(kme_cddip2_ob_out[39]));
Q_ASSIGN U536 ( .B(kme_cddip2_ob_out_post[38]), .A(kme_cddip2_ob_out[38]));
Q_ASSIGN U537 ( .B(kme_cddip2_ob_out_post[37]), .A(kme_cddip2_ob_out[37]));
Q_ASSIGN U538 ( .B(kme_cddip2_ob_out_post[36]), .A(kme_cddip2_ob_out[36]));
Q_ASSIGN U539 ( .B(kme_cddip2_ob_out_post[35]), .A(kme_cddip2_ob_out[35]));
Q_ASSIGN U540 ( .B(kme_cddip2_ob_out_post[34]), .A(kme_cddip2_ob_out[34]));
Q_ASSIGN U541 ( .B(kme_cddip2_ob_out_post[33]), .A(kme_cddip2_ob_out[33]));
Q_ASSIGN U542 ( .B(kme_cddip2_ob_out_post[32]), .A(kme_cddip2_ob_out[32]));
Q_ASSIGN U543 ( .B(kme_cddip2_ob_out_post[31]), .A(kme_cddip2_ob_out[31]));
Q_ASSIGN U544 ( .B(kme_cddip2_ob_out_post[30]), .A(kme_cddip2_ob_out[30]));
Q_ASSIGN U545 ( .B(kme_cddip2_ob_out_post[29]), .A(kme_cddip2_ob_out[29]));
Q_ASSIGN U546 ( .B(kme_cddip2_ob_out_post[28]), .A(kme_cddip2_ob_out[28]));
Q_ASSIGN U547 ( .B(kme_cddip2_ob_out_post[27]), .A(kme_cddip2_ob_out[27]));
Q_ASSIGN U548 ( .B(kme_cddip2_ob_out_post[26]), .A(kme_cddip2_ob_out[26]));
Q_ASSIGN U549 ( .B(kme_cddip2_ob_out_post[25]), .A(kme_cddip2_ob_out[25]));
Q_ASSIGN U550 ( .B(kme_cddip2_ob_out_post[24]), .A(kme_cddip2_ob_out[24]));
Q_ASSIGN U551 ( .B(kme_cddip2_ob_out_post[23]), .A(kme_cddip2_ob_out[23]));
Q_ASSIGN U552 ( .B(kme_cddip2_ob_out_post[22]), .A(kme_cddip2_ob_out[22]));
Q_ASSIGN U553 ( .B(kme_cddip2_ob_out_post[21]), .A(kme_cddip2_ob_out[21]));
Q_ASSIGN U554 ( .B(kme_cddip2_ob_out_post[20]), .A(kme_cddip2_ob_out[20]));
Q_ASSIGN U555 ( .B(kme_cddip2_ob_out_post[19]), .A(kme_cddip2_ob_out[19]));
Q_ASSIGN U556 ( .B(kme_cddip2_ob_out_post[18]), .A(kme_cddip2_ob_out[18]));
Q_ASSIGN U557 ( .B(kme_cddip2_ob_out_post[17]), .A(kme_cddip2_ob_out[17]));
Q_ASSIGN U558 ( .B(kme_cddip2_ob_out_post[16]), .A(kme_cddip2_ob_out[16]));
Q_ASSIGN U559 ( .B(kme_cddip2_ob_out_post[15]), .A(kme_cddip2_ob_out[15]));
Q_ASSIGN U560 ( .B(kme_cddip2_ob_out_post[14]), .A(kme_cddip2_ob_out[14]));
Q_ASSIGN U561 ( .B(kme_cddip2_ob_out_post[13]), .A(kme_cddip2_ob_out[13]));
Q_ASSIGN U562 ( .B(kme_cddip2_ob_out_post[12]), .A(kme_cddip2_ob_out[12]));
Q_ASSIGN U563 ( .B(kme_cddip2_ob_out_post[11]), .A(kme_cddip2_ob_out[11]));
Q_ASSIGN U564 ( .B(kme_cddip2_ob_out_post[10]), .A(kme_cddip2_ob_out[10]));
Q_ASSIGN U565 ( .B(kme_cddip2_ob_out_post[9]), .A(kme_cddip2_ob_out[9]));
Q_ASSIGN U566 ( .B(kme_cddip2_ob_out_post[8]), .A(kme_cddip2_ob_out[8]));
Q_ASSIGN U567 ( .B(kme_cddip2_ob_out_post[7]), .A(kme_cddip2_ob_out[7]));
Q_ASSIGN U568 ( .B(kme_cddip2_ob_out_post[6]), .A(kme_cddip2_ob_out[6]));
Q_ASSIGN U569 ( .B(kme_cddip2_ob_out_post[5]), .A(kme_cddip2_ob_out[5]));
Q_ASSIGN U570 ( .B(kme_cddip2_ob_out_post[4]), .A(kme_cddip2_ob_out[4]));
Q_ASSIGN U571 ( .B(kme_cddip2_ob_out_post[3]), .A(kme_cddip2_ob_out[3]));
Q_ASSIGN U572 ( .B(kme_cddip2_ob_out_post[2]), .A(kme_cddip2_ob_out[2]));
Q_ASSIGN U573 ( .B(kme_cddip2_ob_out_post[1]), .A(kme_cddip2_ob_out[1]));
Q_ASSIGN U574 ( .B(kme_cddip2_ob_out_post[0]), .A(kme_cddip2_ob_out[0]));
Q_ASSIGN U575 ( .B(kme_cddip3_ob_out_post[81]), .A(kme_cddip3_ob_out[81]));
Q_ASSIGN U576 ( .B(kme_cddip3_ob_out_post[80]), .A(kme_cddip3_ob_out[80]));
Q_ASSIGN U577 ( .B(kme_cddip3_ob_out_post[79]), .A(kme_cddip3_ob_out[79]));
Q_ASSIGN U578 ( .B(kme_cddip3_ob_out_post[78]), .A(kme_cddip3_ob_out[78]));
Q_ASSIGN U579 ( .B(kme_cddip3_ob_out_post[77]), .A(kme_cddip3_ob_out[77]));
Q_ASSIGN U580 ( .B(kme_cddip3_ob_out_post[76]), .A(kme_cddip3_ob_out[76]));
Q_ASSIGN U581 ( .B(kme_cddip3_ob_out_post[75]), .A(kme_cddip3_ob_out[75]));
Q_ASSIGN U582 ( .B(kme_cddip3_ob_out_post[74]), .A(kme_cddip3_ob_out[74]));
Q_ASSIGN U583 ( .B(kme_cddip3_ob_out_post[73]), .A(kme_cddip3_ob_out[73]));
Q_ASSIGN U584 ( .B(kme_cddip3_ob_out_post[72]), .A(kme_cddip3_ob_out[72]));
Q_ASSIGN U585 ( .B(kme_cddip3_ob_out_post[71]), .A(kme_cddip3_ob_out[71]));
Q_ASSIGN U586 ( .B(kme_cddip3_ob_out_post[70]), .A(kme_cddip3_ob_out[70]));
Q_ASSIGN U587 ( .B(kme_cddip3_ob_out_post[69]), .A(kme_cddip3_ob_out[69]));
Q_ASSIGN U588 ( .B(kme_cddip3_ob_out_post[68]), .A(kme_cddip3_ob_out[68]));
Q_ASSIGN U589 ( .B(kme_cddip3_ob_out_post[67]), .A(kme_cddip3_ob_out[67]));
Q_ASSIGN U590 ( .B(kme_cddip3_ob_out_post[66]), .A(kme_cddip3_ob_out[66]));
Q_ASSIGN U591 ( .B(kme_cddip3_ob_out_post[65]), .A(kme_cddip3_ob_out[65]));
Q_ASSIGN U592 ( .B(kme_cddip3_ob_out_post[64]), .A(kme_cddip3_ob_out[64]));
Q_ASSIGN U593 ( .B(kme_cddip3_ob_out_post[63]), .A(kme_cddip3_ob_out[63]));
Q_ASSIGN U594 ( .B(kme_cddip3_ob_out_post[62]), .A(kme_cddip3_ob_out[62]));
Q_ASSIGN U595 ( .B(kme_cddip3_ob_out_post[61]), .A(kme_cddip3_ob_out[61]));
Q_ASSIGN U596 ( .B(kme_cddip3_ob_out_post[60]), .A(kme_cddip3_ob_out[60]));
Q_ASSIGN U597 ( .B(kme_cddip3_ob_out_post[59]), .A(kme_cddip3_ob_out[59]));
Q_ASSIGN U598 ( .B(kme_cddip3_ob_out_post[58]), .A(kme_cddip3_ob_out[58]));
Q_ASSIGN U599 ( .B(kme_cddip3_ob_out_post[57]), .A(kme_cddip3_ob_out[57]));
Q_ASSIGN U600 ( .B(kme_cddip3_ob_out_post[56]), .A(kme_cddip3_ob_out[56]));
Q_ASSIGN U601 ( .B(kme_cddip3_ob_out_post[55]), .A(kme_cddip3_ob_out[55]));
Q_ASSIGN U602 ( .B(kme_cddip3_ob_out_post[54]), .A(kme_cddip3_ob_out[54]));
Q_ASSIGN U603 ( .B(kme_cddip3_ob_out_post[53]), .A(kme_cddip3_ob_out[53]));
Q_ASSIGN U604 ( .B(kme_cddip3_ob_out_post[52]), .A(kme_cddip3_ob_out[52]));
Q_ASSIGN U605 ( .B(kme_cddip3_ob_out_post[51]), .A(kme_cddip3_ob_out[51]));
Q_ASSIGN U606 ( .B(kme_cddip3_ob_out_post[50]), .A(kme_cddip3_ob_out[50]));
Q_ASSIGN U607 ( .B(kme_cddip3_ob_out_post[49]), .A(kme_cddip3_ob_out[49]));
Q_ASSIGN U608 ( .B(kme_cddip3_ob_out_post[48]), .A(kme_cddip3_ob_out[48]));
Q_ASSIGN U609 ( .B(kme_cddip3_ob_out_post[47]), .A(kme_cddip3_ob_out[47]));
Q_ASSIGN U610 ( .B(kme_cddip3_ob_out_post[46]), .A(kme_cddip3_ob_out[46]));
Q_ASSIGN U611 ( .B(kme_cddip3_ob_out_post[45]), .A(kme_cddip3_ob_out[45]));
Q_ASSIGN U612 ( .B(kme_cddip3_ob_out_post[44]), .A(kme_cddip3_ob_out[44]));
Q_ASSIGN U613 ( .B(kme_cddip3_ob_out_post[43]), .A(kme_cddip3_ob_out[43]));
Q_ASSIGN U614 ( .B(kme_cddip3_ob_out_post[42]), .A(kme_cddip3_ob_out[42]));
Q_ASSIGN U615 ( .B(kme_cddip3_ob_out_post[41]), .A(kme_cddip3_ob_out[41]));
Q_ASSIGN U616 ( .B(kme_cddip3_ob_out_post[40]), .A(kme_cddip3_ob_out[40]));
Q_ASSIGN U617 ( .B(kme_cddip3_ob_out_post[39]), .A(kme_cddip3_ob_out[39]));
Q_ASSIGN U618 ( .B(kme_cddip3_ob_out_post[38]), .A(kme_cddip3_ob_out[38]));
Q_ASSIGN U619 ( .B(kme_cddip3_ob_out_post[37]), .A(kme_cddip3_ob_out[37]));
Q_ASSIGN U620 ( .B(kme_cddip3_ob_out_post[36]), .A(kme_cddip3_ob_out[36]));
Q_ASSIGN U621 ( .B(kme_cddip3_ob_out_post[35]), .A(kme_cddip3_ob_out[35]));
Q_ASSIGN U622 ( .B(kme_cddip3_ob_out_post[34]), .A(kme_cddip3_ob_out[34]));
Q_ASSIGN U623 ( .B(kme_cddip3_ob_out_post[33]), .A(kme_cddip3_ob_out[33]));
Q_ASSIGN U624 ( .B(kme_cddip3_ob_out_post[32]), .A(kme_cddip3_ob_out[32]));
Q_ASSIGN U625 ( .B(kme_cddip3_ob_out_post[31]), .A(kme_cddip3_ob_out[31]));
Q_ASSIGN U626 ( .B(kme_cddip3_ob_out_post[30]), .A(kme_cddip3_ob_out[30]));
Q_ASSIGN U627 ( .B(kme_cddip3_ob_out_post[29]), .A(kme_cddip3_ob_out[29]));
Q_ASSIGN U628 ( .B(kme_cddip3_ob_out_post[28]), .A(kme_cddip3_ob_out[28]));
Q_ASSIGN U629 ( .B(kme_cddip3_ob_out_post[27]), .A(kme_cddip3_ob_out[27]));
Q_ASSIGN U630 ( .B(kme_cddip3_ob_out_post[26]), .A(kme_cddip3_ob_out[26]));
Q_ASSIGN U631 ( .B(kme_cddip3_ob_out_post[25]), .A(kme_cddip3_ob_out[25]));
Q_ASSIGN U632 ( .B(kme_cddip3_ob_out_post[24]), .A(kme_cddip3_ob_out[24]));
Q_ASSIGN U633 ( .B(kme_cddip3_ob_out_post[23]), .A(kme_cddip3_ob_out[23]));
Q_ASSIGN U634 ( .B(kme_cddip3_ob_out_post[22]), .A(kme_cddip3_ob_out[22]));
Q_ASSIGN U635 ( .B(kme_cddip3_ob_out_post[21]), .A(kme_cddip3_ob_out[21]));
Q_ASSIGN U636 ( .B(kme_cddip3_ob_out_post[20]), .A(kme_cddip3_ob_out[20]));
Q_ASSIGN U637 ( .B(kme_cddip3_ob_out_post[19]), .A(kme_cddip3_ob_out[19]));
Q_ASSIGN U638 ( .B(kme_cddip3_ob_out_post[18]), .A(kme_cddip3_ob_out[18]));
Q_ASSIGN U639 ( .B(kme_cddip3_ob_out_post[17]), .A(kme_cddip3_ob_out[17]));
Q_ASSIGN U640 ( .B(kme_cddip3_ob_out_post[16]), .A(kme_cddip3_ob_out[16]));
Q_ASSIGN U641 ( .B(kme_cddip3_ob_out_post[15]), .A(kme_cddip3_ob_out[15]));
Q_ASSIGN U642 ( .B(kme_cddip3_ob_out_post[14]), .A(kme_cddip3_ob_out[14]));
Q_ASSIGN U643 ( .B(kme_cddip3_ob_out_post[13]), .A(kme_cddip3_ob_out[13]));
Q_ASSIGN U644 ( .B(kme_cddip3_ob_out_post[12]), .A(kme_cddip3_ob_out[12]));
Q_ASSIGN U645 ( .B(kme_cddip3_ob_out_post[11]), .A(kme_cddip3_ob_out[11]));
Q_ASSIGN U646 ( .B(kme_cddip3_ob_out_post[10]), .A(kme_cddip3_ob_out[10]));
Q_ASSIGN U647 ( .B(kme_cddip3_ob_out_post[9]), .A(kme_cddip3_ob_out[9]));
Q_ASSIGN U648 ( .B(kme_cddip3_ob_out_post[8]), .A(kme_cddip3_ob_out[8]));
Q_ASSIGN U649 ( .B(kme_cddip3_ob_out_post[7]), .A(kme_cddip3_ob_out[7]));
Q_ASSIGN U650 ( .B(kme_cddip3_ob_out_post[6]), .A(kme_cddip3_ob_out[6]));
Q_ASSIGN U651 ( .B(kme_cddip3_ob_out_post[5]), .A(kme_cddip3_ob_out[5]));
Q_ASSIGN U652 ( .B(kme_cddip3_ob_out_post[4]), .A(kme_cddip3_ob_out[4]));
Q_ASSIGN U653 ( .B(kme_cddip3_ob_out_post[3]), .A(kme_cddip3_ob_out[3]));
Q_ASSIGN U654 ( .B(kme_cddip3_ob_out_post[2]), .A(kme_cddip3_ob_out[2]));
Q_ASSIGN U655 ( .B(kme_cddip3_ob_out_post[1]), .A(kme_cddip3_ob_out[1]));
Q_ASSIGN U656 ( .B(kme_cddip3_ob_out_post[0]), .A(kme_cddip3_ob_out[0]));
Q_INV U657 ( .A(tready_override[0]), .Z(n1));
Q_INV U658 ( .A(tready_override[1]), .Z(n2));
Q_INV U659 ( .A(tready_override[2]), .Z(n3));
Q_INV U660 ( .A(tready_override[3]), .Z(n4));
Q_INV U661 ( .A(tready_override[4]), .Z(n5));
Q_INV U662 ( .A(tready_override[5]), .Z(n6));
Q_INV U663 ( .A(tready_override[6]), .Z(n7));
Q_INV U664 ( .A(tready_override[7]), .Z(n8));
Q_AN02 U665 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[31]), .Z(debug_kme_ib_tlast));
Q_AN02 U666 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[14]), .Z(debug_kme_ib_tid[0]));
Q_AN02 U667 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[30]), .Z(debug_kme_ib_tstrb[7]));
Q_AN02 U668 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[29]), .Z(debug_kme_ib_tstrb[6]));
Q_AN02 U669 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[28]), .Z(debug_kme_ib_tstrb[5]));
Q_AN02 U670 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[27]), .Z(debug_kme_ib_tstrb[4]));
Q_AN02 U671 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[26]), .Z(debug_kme_ib_tstrb[3]));
Q_AN02 U672 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[25]), .Z(debug_kme_ib_tstrb[2]));
Q_AN02 U673 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[24]), .Z(debug_kme_ib_tstrb[1]));
Q_AN02 U674 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[23]), .Z(debug_kme_ib_tstrb[0]));
Q_AN02 U675 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[13]), .Z(debug_kme_ib_tuser[7]));
Q_AN02 U676 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[12]), .Z(debug_kme_ib_tuser[6]));
Q_AN02 U677 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[11]), .Z(debug_kme_ib_tuser[5]));
Q_AN02 U678 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[10]), .Z(debug_kme_ib_tuser[4]));
Q_AN02 U679 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[9]), .Z(debug_kme_ib_tuser[3]));
Q_AN02 U680 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[8]), .Z(debug_kme_ib_tuser[2]));
Q_AN02 U681 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[7]), .Z(debug_kme_ib_tuser[1]));
Q_AN02 U682 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[6]), .Z(debug_kme_ib_tuser[0]));
Q_AN02 U683 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[95]), .Z(debug_kme_ib_tdata[63]));
Q_AN02 U684 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[94]), .Z(debug_kme_ib_tdata[62]));
Q_AN02 U685 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[93]), .Z(debug_kme_ib_tdata[61]));
Q_AN02 U686 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[92]), .Z(debug_kme_ib_tdata[60]));
Q_AN02 U687 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[91]), .Z(debug_kme_ib_tdata[59]));
Q_AN02 U688 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[90]), .Z(debug_kme_ib_tdata[58]));
Q_AN02 U689 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[89]), .Z(debug_kme_ib_tdata[57]));
Q_AN02 U690 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[88]), .Z(debug_kme_ib_tdata[56]));
Q_AN02 U691 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[87]), .Z(debug_kme_ib_tdata[55]));
Q_AN02 U692 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[86]), .Z(debug_kme_ib_tdata[54]));
Q_AN02 U693 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[85]), .Z(debug_kme_ib_tdata[53]));
Q_AN02 U694 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[84]), .Z(debug_kme_ib_tdata[52]));
Q_AN02 U695 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[83]), .Z(debug_kme_ib_tdata[51]));
Q_AN02 U696 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[82]), .Z(debug_kme_ib_tdata[50]));
Q_AN02 U697 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[81]), .Z(debug_kme_ib_tdata[49]));
Q_AN02 U698 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[80]), .Z(debug_kme_ib_tdata[48]));
Q_AN02 U699 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[79]), .Z(debug_kme_ib_tdata[47]));
Q_AN02 U700 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[78]), .Z(debug_kme_ib_tdata[46]));
Q_AN02 U701 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[77]), .Z(debug_kme_ib_tdata[45]));
Q_AN02 U702 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[76]), .Z(debug_kme_ib_tdata[44]));
Q_AN02 U703 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[75]), .Z(debug_kme_ib_tdata[43]));
Q_AN02 U704 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[74]), .Z(debug_kme_ib_tdata[42]));
Q_AN02 U705 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[73]), .Z(debug_kme_ib_tdata[41]));
Q_AN02 U706 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[72]), .Z(debug_kme_ib_tdata[40]));
Q_AN02 U707 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[71]), .Z(debug_kme_ib_tdata[39]));
Q_AN02 U708 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[70]), .Z(debug_kme_ib_tdata[38]));
Q_AN02 U709 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[69]), .Z(debug_kme_ib_tdata[37]));
Q_AN02 U710 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[68]), .Z(debug_kme_ib_tdata[36]));
Q_AN02 U711 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[67]), .Z(debug_kme_ib_tdata[35]));
Q_AN02 U712 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[66]), .Z(debug_kme_ib_tdata[34]));
Q_AN02 U713 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[65]), .Z(debug_kme_ib_tdata[33]));
Q_AN02 U714 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[64]), .Z(debug_kme_ib_tdata[32]));
Q_AN02 U715 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[63]), .Z(debug_kme_ib_tdata[31]));
Q_AN02 U716 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[62]), .Z(debug_kme_ib_tdata[30]));
Q_AN02 U717 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[61]), .Z(debug_kme_ib_tdata[29]));
Q_AN02 U718 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[60]), .Z(debug_kme_ib_tdata[28]));
Q_AN02 U719 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[59]), .Z(debug_kme_ib_tdata[27]));
Q_AN02 U720 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[58]), .Z(debug_kme_ib_tdata[26]));
Q_AN02 U721 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[57]), .Z(debug_kme_ib_tdata[25]));
Q_AN02 U722 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[56]), .Z(debug_kme_ib_tdata[24]));
Q_AN02 U723 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[55]), .Z(debug_kme_ib_tdata[23]));
Q_AN02 U724 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[54]), .Z(debug_kme_ib_tdata[22]));
Q_AN02 U725 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[53]), .Z(debug_kme_ib_tdata[21]));
Q_AN02 U726 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[52]), .Z(debug_kme_ib_tdata[20]));
Q_AN02 U727 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[51]), .Z(debug_kme_ib_tdata[19]));
Q_AN02 U728 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[50]), .Z(debug_kme_ib_tdata[18]));
Q_AN02 U729 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[49]), .Z(debug_kme_ib_tdata[17]));
Q_AN02 U730 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[48]), .Z(debug_kme_ib_tdata[16]));
Q_AN02 U731 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[47]), .Z(debug_kme_ib_tdata[15]));
Q_AN02 U732 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[46]), .Z(debug_kme_ib_tdata[14]));
Q_AN02 U733 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[45]), .Z(debug_kme_ib_tdata[13]));
Q_AN02 U734 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[44]), .Z(debug_kme_ib_tdata[12]));
Q_AN02 U735 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[43]), .Z(debug_kme_ib_tdata[11]));
Q_AN02 U736 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[42]), .Z(debug_kme_ib_tdata[10]));
Q_AN02 U737 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[41]), .Z(debug_kme_ib_tdata[9]));
Q_AN02 U738 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[40]), .Z(debug_kme_ib_tdata[8]));
Q_AN02 U739 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[39]), .Z(debug_kme_ib_tdata[7]));
Q_AN02 U740 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[38]), .Z(debug_kme_ib_tdata[6]));
Q_AN02 U741 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[37]), .Z(debug_kme_ib_tdata[5]));
Q_AN02 U742 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[36]), .Z(debug_kme_ib_tdata[4]));
Q_AN02 U743 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[35]), .Z(debug_kme_ib_tdata[3]));
Q_AN02 U744 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[34]), .Z(debug_kme_ib_tdata[2]));
Q_AN02 U745 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[33]), .Z(debug_kme_ib_tdata[1]));
Q_AN02 U746 ( .A0(send_kme_ib_beat), .A1(cceip0_out_ia_wdata[32]), .Z(debug_kme_ib_tdata[0]));
Q_AN02 U747 ( .A0(n1), .A1(kme_cceip0_ob_out_post[82]), .Z(kme_cceip0_ob_out[82]));
Q_AN02 U748 ( .A0(n2), .A1(kme_cceip1_ob_out_post[82]), .Z(kme_cceip1_ob_out[82]));
Q_AN02 U749 ( .A0(n3), .A1(kme_cceip2_ob_out_post[82]), .Z(kme_cceip2_ob_out[82]));
Q_AN02 U750 ( .A0(n4), .A1(kme_cceip3_ob_out_post[82]), .Z(kme_cceip3_ob_out[82]));
Q_AN02 U751 ( .A0(n5), .A1(kme_cddip0_ob_out_post[82]), .Z(kme_cddip0_ob_out[82]));
Q_AN02 U752 ( .A0(n6), .A1(kme_cddip1_ob_out_post[82]), .Z(kme_cddip1_ob_out[82]));
Q_AN02 U753 ( .A0(n7), .A1(kme_cddip2_ob_out_post[82]), .Z(kme_cddip2_ob_out[82]));
Q_AN02 U754 ( .A0(n8), .A1(kme_cddip3_ob_out_post[82]), .Z(kme_cddip3_ob_out[82]));
Q_NR02 U755 ( .A0(send_kme_ib_beat), .A1(n9), .Z(n11));
Q_INV U756 ( .A(debug_kme_ib_tready), .Z(n10));
Q_AO21 U757 ( .A0(send_kme_ib_beat), .A1(n10), .B0(n11), .Z(n12));
Q_AO21 U758 ( .A0(n13), .A1(wr_data[1]), .B0(disable_ckv_kim_ism_reads), .Z(n20));
Q_AN02 U759 ( .A0(n13), .A1(wr_data[0]), .Z(n9));
Q_AN02 U760 ( .A0(wr_stb), .A1(n14), .Z(n13));
Q_NR03 U761 ( .A0(n17), .A1(n16), .A2(n15), .Z(n14));
Q_OR03 U762 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n18), .Z(n15));
Q_OR03 U763 ( .A0(reg_addr[4]), .A1(n19), .A2(reg_addr[2]), .Z(n16));
Q_OR03 U764 ( .A0(reg_addr[7]), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n17));
Q_OR03 U765 ( .A0(reg_addr[10]), .A1(reg_addr[9]), .A2(reg_addr[8]), .Z(n18));
Q_INV U766 ( .A(reg_addr[3]), .Z(n19));
Q_FDP1 disable_ckv_kim_ism_reads_REG  ( .CK(clk), .R(rst_n), .D(n20), .Q(disable_ckv_kim_ism_reads), .QN(n55));
Q_INV U768 ( .A(n28), .Z(n36));
Q_NR02 U769 ( .A0(n28), .A1(set_rsm_is_backpressuring[0]), .Z(n37));
Q_INV U770 ( .A(n27), .Z(n35));
Q_NR02 U771 ( .A0(n27), .A1(set_rsm_is_backpressuring[1]), .Z(n38));
Q_INV U772 ( .A(n26), .Z(n34));
Q_NR02 U773 ( .A0(n26), .A1(set_rsm_is_backpressuring[2]), .Z(n39));
Q_INV U774 ( .A(n25), .Z(n33));
Q_NR02 U775 ( .A0(n25), .A1(set_rsm_is_backpressuring[3]), .Z(n40));
Q_INV U776 ( .A(n24), .Z(n32));
Q_NR02 U777 ( .A0(n24), .A1(set_rsm_is_backpressuring[4]), .Z(n41));
Q_INV U778 ( .A(n23), .Z(n31));
Q_NR02 U779 ( .A0(n23), .A1(set_rsm_is_backpressuring[5]), .Z(n42));
Q_INV U780 ( .A(n22), .Z(n30));
Q_NR02 U781 ( .A0(n22), .A1(set_rsm_is_backpressuring[6]), .Z(n43));
Q_INV U782 ( .A(n21), .Z(n29));
Q_NR02 U783 ( .A0(n21), .A1(set_rsm_is_backpressuring[7]), .Z(n44));
Q_AN02 U784 ( .A0(n45), .A1(wr_data[7]), .Z(n21));
Q_AN02 U785 ( .A0(n45), .A1(wr_data[6]), .Z(n22));
Q_AN02 U786 ( .A0(n45), .A1(wr_data[5]), .Z(n23));
Q_AN02 U787 ( .A0(n45), .A1(wr_data[4]), .Z(n24));
Q_AN02 U788 ( .A0(n45), .A1(wr_data[3]), .Z(n25));
Q_AN02 U789 ( .A0(n45), .A1(wr_data[2]), .Z(n26));
Q_AN02 U790 ( .A0(n45), .A1(wr_data[1]), .Z(n27));
Q_AN02 U791 ( .A0(n45), .A1(wr_data[0]), .Z(n28));
Q_AN02 U792 ( .A0(wr_stb), .A1(n46), .Z(n45));
Q_NR03 U793 ( .A0(n49), .A1(n48), .A2(n47), .Z(n46));
Q_OR03 U794 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n50), .Z(n47));
Q_OR03 U795 ( .A0(reg_addr[4]), .A1(reg_addr[3]), .A2(n54), .Z(n48));
Q_OR03 U796 ( .A0(n53), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n49));
Q_OR03 U797 ( .A0(reg_addr[10]), .A1(n51), .A2(n52), .Z(n50));
Q_INV U798 ( .A(reg_addr[9]), .Z(n51));
Q_INV U799 ( .A(reg_addr[8]), .Z(n52));
Q_INV U800 ( .A(reg_addr[7]), .Z(n53));
Q_INV U801 ( .A(reg_addr[2]), .Z(n54));
Q_AN02 U802 ( .A0(n55), .A1(kim_rd_dat[37]), .Z(kim_ia_rdata_part0[20]));
Q_AN02 U803 ( .A0(n55), .A1(kim_rd_dat[36]), .Z(kim_ia_rdata_part0[19]));
Q_AN02 U804 ( .A0(n55), .A1(kim_rd_dat[35]), .Z(kim_ia_rdata_part0[18]));
Q_AN02 U805 ( .A0(n55), .A1(kim_rd_dat[34]), .Z(kim_ia_rdata_part0[17]));
Q_AN02 U806 ( .A0(n55), .A1(kim_rd_dat[33]), .Z(kim_ia_rdata_part0[16]));
Q_AN02 U807 ( .A0(n55), .A1(kim_rd_dat[32]), .Z(kim_ia_rdata_part0[15]));
Q_AN02 U808 ( .A0(n55), .A1(kim_rd_dat[31]), .Z(kim_ia_rdata_part0[14]));
Q_AN02 U809 ( .A0(n55), .A1(kim_rd_dat[30]), .Z(kim_ia_rdata_part0[13]));
Q_AN02 U810 ( .A0(n55), .A1(kim_rd_dat[29]), .Z(kim_ia_rdata_part0[12]));
Q_AN02 U811 ( .A0(n55), .A1(kim_rd_dat[28]), .Z(kim_ia_rdata_part0[11]));
Q_AN02 U812 ( .A0(n55), .A1(kim_rd_dat[27]), .Z(kim_ia_rdata_part0[10]));
Q_AN02 U813 ( .A0(n55), .A1(kim_rd_dat[26]), .Z(kim_ia_rdata_part0[9]));
Q_AN02 U814 ( .A0(n55), .A1(kim_rd_dat[25]), .Z(kim_ia_rdata_part0[8]));
Q_AN02 U815 ( .A0(n55), .A1(kim_rd_dat[24]), .Z(kim_ia_rdata_part0[7]));
Q_AN02 U816 ( .A0(n55), .A1(kim_rd_dat[23]), .Z(kim_ia_rdata_part0[6]));
Q_AN02 U817 ( .A0(n55), .A1(kim_rd_dat[22]), .Z(kim_ia_rdata_part0[5]));
Q_AN02 U818 ( .A0(n55), .A1(kim_rd_dat[21]), .Z(kim_ia_rdata_part0[4]));
Q_AN02 U819 ( .A0(n55), .A1(kim_rd_dat[20]), .Z(kim_ia_rdata_part0[3]));
Q_AN02 U820 ( .A0(n55), .A1(kim_rd_dat[19]), .Z(kim_ia_rdata_part0[2]));
Q_AN02 U821 ( .A0(n55), .A1(kim_rd_dat[18]), .Z(kim_ia_rdata_part0[1]));
Q_AN02 U822 ( .A0(n55), .A1(kim_rd_dat[17]), .Z(kim_ia_rdata_part0[0]));
Q_AN02 U823 ( .A0(n55), .A1(kim_rd_dat[16]), .Z(kim_ia_rdata_part1[16]));
Q_AN02 U824 ( .A0(n55), .A1(kim_rd_dat[15]), .Z(kim_ia_rdata_part1[15]));
Q_AN02 U825 ( .A0(n55), .A1(kim_rd_dat[14]), .Z(kim_ia_rdata_part1[14]));
Q_AN02 U826 ( .A0(n55), .A1(kim_rd_dat[13]), .Z(kim_ia_rdata_part1[13]));
Q_AN02 U827 ( .A0(n55), .A1(kim_rd_dat[12]), .Z(kim_ia_rdata_part1[12]));
Q_AN02 U828 ( .A0(n55), .A1(kim_rd_dat[11]), .Z(kim_ia_rdata_part1[11]));
Q_AN02 U829 ( .A0(n55), .A1(kim_rd_dat[10]), .Z(kim_ia_rdata_part1[10]));
Q_AN02 U830 ( .A0(n55), .A1(kim_rd_dat[9]), .Z(kim_ia_rdata_part1[9]));
Q_AN02 U831 ( .A0(n55), .A1(kim_rd_dat[8]), .Z(kim_ia_rdata_part1[8]));
Q_AN02 U832 ( .A0(n55), .A1(kim_rd_dat[7]), .Z(kim_ia_rdata_part1[7]));
Q_AN02 U833 ( .A0(n55), .A1(kim_rd_dat[6]), .Z(kim_ia_rdata_part1[6]));
Q_AN02 U834 ( .A0(n55), .A1(kim_rd_dat[5]), .Z(kim_ia_rdata_part1[5]));
Q_AN02 U835 ( .A0(n55), .A1(kim_rd_dat[4]), .Z(kim_ia_rdata_part1[4]));
Q_AN02 U836 ( .A0(n55), .A1(kim_rd_dat[3]), .Z(kim_ia_rdata_part1[3]));
Q_AN02 U837 ( .A0(n55), .A1(kim_rd_dat[2]), .Z(kim_ia_rdata_part1[2]));
Q_AN02 U838 ( .A0(n55), .A1(kim_rd_dat[1]), .Z(kim_ia_rdata_part1[1]));
Q_AN02 U839 ( .A0(n55), .A1(kim_rd_dat[0]), .Z(kim_ia_rdata_part1[0]));
Q_AN02 U840 ( .A0(n55), .A1(ckv_rd_dat[63]), .Z(ckv_ia_rdata_part1[31]));
Q_AN02 U841 ( .A0(n55), .A1(ckv_rd_dat[62]), .Z(ckv_ia_rdata_part1[30]));
Q_AN02 U842 ( .A0(n55), .A1(ckv_rd_dat[61]), .Z(ckv_ia_rdata_part1[29]));
Q_AN02 U843 ( .A0(n55), .A1(ckv_rd_dat[60]), .Z(ckv_ia_rdata_part1[28]));
Q_AN02 U844 ( .A0(n55), .A1(ckv_rd_dat[59]), .Z(ckv_ia_rdata_part1[27]));
Q_AN02 U845 ( .A0(n55), .A1(ckv_rd_dat[58]), .Z(ckv_ia_rdata_part1[26]));
Q_AN02 U846 ( .A0(n55), .A1(ckv_rd_dat[57]), .Z(ckv_ia_rdata_part1[25]));
Q_AN02 U847 ( .A0(n55), .A1(ckv_rd_dat[56]), .Z(ckv_ia_rdata_part1[24]));
Q_AN02 U848 ( .A0(n55), .A1(ckv_rd_dat[55]), .Z(ckv_ia_rdata_part1[23]));
Q_AN02 U849 ( .A0(n55), .A1(ckv_rd_dat[54]), .Z(ckv_ia_rdata_part1[22]));
Q_AN02 U850 ( .A0(n55), .A1(ckv_rd_dat[53]), .Z(ckv_ia_rdata_part1[21]));
Q_AN02 U851 ( .A0(n55), .A1(ckv_rd_dat[52]), .Z(ckv_ia_rdata_part1[20]));
Q_AN02 U852 ( .A0(n55), .A1(ckv_rd_dat[51]), .Z(ckv_ia_rdata_part1[19]));
Q_AN02 U853 ( .A0(n55), .A1(ckv_rd_dat[50]), .Z(ckv_ia_rdata_part1[18]));
Q_AN02 U854 ( .A0(n55), .A1(ckv_rd_dat[49]), .Z(ckv_ia_rdata_part1[17]));
Q_AN02 U855 ( .A0(n55), .A1(ckv_rd_dat[48]), .Z(ckv_ia_rdata_part1[16]));
Q_AN02 U856 ( .A0(n55), .A1(ckv_rd_dat[47]), .Z(ckv_ia_rdata_part1[15]));
Q_AN02 U857 ( .A0(n55), .A1(ckv_rd_dat[46]), .Z(ckv_ia_rdata_part1[14]));
Q_AN02 U858 ( .A0(n55), .A1(ckv_rd_dat[45]), .Z(ckv_ia_rdata_part1[13]));
Q_AN02 U859 ( .A0(n55), .A1(ckv_rd_dat[44]), .Z(ckv_ia_rdata_part1[12]));
Q_AN02 U860 ( .A0(n55), .A1(ckv_rd_dat[43]), .Z(ckv_ia_rdata_part1[11]));
Q_AN02 U861 ( .A0(n55), .A1(ckv_rd_dat[42]), .Z(ckv_ia_rdata_part1[10]));
Q_AN02 U862 ( .A0(n55), .A1(ckv_rd_dat[41]), .Z(ckv_ia_rdata_part1[9]));
Q_AN02 U863 ( .A0(n55), .A1(ckv_rd_dat[40]), .Z(ckv_ia_rdata_part1[8]));
Q_AN02 U864 ( .A0(n55), .A1(ckv_rd_dat[39]), .Z(ckv_ia_rdata_part1[7]));
Q_AN02 U865 ( .A0(n55), .A1(ckv_rd_dat[38]), .Z(ckv_ia_rdata_part1[6]));
Q_AN02 U866 ( .A0(n55), .A1(ckv_rd_dat[37]), .Z(ckv_ia_rdata_part1[5]));
Q_AN02 U867 ( .A0(n55), .A1(ckv_rd_dat[36]), .Z(ckv_ia_rdata_part1[4]));
Q_AN02 U868 ( .A0(n55), .A1(ckv_rd_dat[35]), .Z(ckv_ia_rdata_part1[3]));
Q_AN02 U869 ( .A0(n55), .A1(ckv_rd_dat[34]), .Z(ckv_ia_rdata_part1[2]));
Q_AN02 U870 ( .A0(n55), .A1(ckv_rd_dat[33]), .Z(ckv_ia_rdata_part1[1]));
Q_AN02 U871 ( .A0(n55), .A1(ckv_rd_dat[32]), .Z(ckv_ia_rdata_part1[0]));
Q_AN02 U872 ( .A0(n55), .A1(ckv_rd_dat[31]), .Z(ckv_ia_rdata_part0[31]));
Q_AN02 U873 ( .A0(n55), .A1(ckv_rd_dat[30]), .Z(ckv_ia_rdata_part0[30]));
Q_AN02 U874 ( .A0(n55), .A1(ckv_rd_dat[29]), .Z(ckv_ia_rdata_part0[29]));
Q_AN02 U875 ( .A0(n55), .A1(ckv_rd_dat[28]), .Z(ckv_ia_rdata_part0[28]));
Q_AN02 U876 ( .A0(n55), .A1(ckv_rd_dat[27]), .Z(ckv_ia_rdata_part0[27]));
Q_AN02 U877 ( .A0(n55), .A1(ckv_rd_dat[26]), .Z(ckv_ia_rdata_part0[26]));
Q_AN02 U878 ( .A0(n55), .A1(ckv_rd_dat[25]), .Z(ckv_ia_rdata_part0[25]));
Q_AN02 U879 ( .A0(n55), .A1(ckv_rd_dat[24]), .Z(ckv_ia_rdata_part0[24]));
Q_AN02 U880 ( .A0(n55), .A1(ckv_rd_dat[23]), .Z(ckv_ia_rdata_part0[23]));
Q_AN02 U881 ( .A0(n55), .A1(ckv_rd_dat[22]), .Z(ckv_ia_rdata_part0[22]));
Q_AN02 U882 ( .A0(n55), .A1(ckv_rd_dat[21]), .Z(ckv_ia_rdata_part0[21]));
Q_AN02 U883 ( .A0(n55), .A1(ckv_rd_dat[20]), .Z(ckv_ia_rdata_part0[20]));
Q_AN02 U884 ( .A0(n55), .A1(ckv_rd_dat[19]), .Z(ckv_ia_rdata_part0[19]));
Q_AN02 U885 ( .A0(n55), .A1(ckv_rd_dat[18]), .Z(ckv_ia_rdata_part0[18]));
Q_AN02 U886 ( .A0(n55), .A1(ckv_rd_dat[17]), .Z(ckv_ia_rdata_part0[17]));
Q_AN02 U887 ( .A0(n55), .A1(ckv_rd_dat[16]), .Z(ckv_ia_rdata_part0[16]));
Q_AN02 U888 ( .A0(n55), .A1(ckv_rd_dat[15]), .Z(ckv_ia_rdata_part0[15]));
Q_AN02 U889 ( .A0(n55), .A1(ckv_rd_dat[14]), .Z(ckv_ia_rdata_part0[14]));
Q_AN02 U890 ( .A0(n55), .A1(ckv_rd_dat[13]), .Z(ckv_ia_rdata_part0[13]));
Q_AN02 U891 ( .A0(n55), .A1(ckv_rd_dat[12]), .Z(ckv_ia_rdata_part0[12]));
Q_AN02 U892 ( .A0(n55), .A1(ckv_rd_dat[11]), .Z(ckv_ia_rdata_part0[11]));
Q_AN02 U893 ( .A0(n55), .A1(ckv_rd_dat[10]), .Z(ckv_ia_rdata_part0[10]));
Q_AN02 U894 ( .A0(n55), .A1(ckv_rd_dat[9]), .Z(ckv_ia_rdata_part0[9]));
Q_AN02 U895 ( .A0(n55), .A1(ckv_rd_dat[8]), .Z(ckv_ia_rdata_part0[8]));
Q_AN02 U896 ( .A0(n55), .A1(ckv_rd_dat[7]), .Z(ckv_ia_rdata_part0[7]));
Q_AN02 U897 ( .A0(n55), .A1(ckv_rd_dat[6]), .Z(ckv_ia_rdata_part0[6]));
Q_AN02 U898 ( .A0(n55), .A1(ckv_rd_dat[5]), .Z(ckv_ia_rdata_part0[5]));
Q_AN02 U899 ( .A0(n55), .A1(ckv_rd_dat[4]), .Z(ckv_ia_rdata_part0[4]));
Q_AN02 U900 ( .A0(n55), .A1(ckv_rd_dat[3]), .Z(ckv_ia_rdata_part0[3]));
Q_AN02 U901 ( .A0(n55), .A1(ckv_rd_dat[2]), .Z(ckv_ia_rdata_part0[2]));
Q_AN02 U902 ( .A0(n55), .A1(ckv_rd_dat[1]), .Z(ckv_ia_rdata_part0[1]));
Q_AN02 U903 ( .A0(n55), .A1(ckv_rd_dat[0]), .Z(ckv_ia_rdata_part0[0]));
ixc_assign_4 _zz_strnp_0 ( ckv_cmnd_op[3:0], o_ckv_ia_config[18:15]);
ixc_assign_15 _zz_strnp_1 ( ckv_cmnd_addr[14:0], o_ckv_ia_config[14:0]);
ixc_assign_20 _zz_strnp_2 ( ckv_ia_capability[19:0], { 
	ckv_capability_type[3], ckv_capability_type[2], 
	ckv_capability_type[1], ckv_capability_type[0], 
	ckv_capability_lst[15], ckv_capability_lst[14], 
	ckv_capability_lst[13], ckv_capability_lst[12], 
	ckv_capability_lst[11], ckv_capability_lst[10], 
	ckv_capability_lst[9], ckv_capability_lst[8], ckv_capability_lst[7], 
	ckv_capability_lst[6], ckv_capability_lst[5], ckv_capability_lst[4], 
	ckv_capability_lst[3], ckv_capability_lst[2], ckv_capability_lst[1], 
	ckv_capability_lst[0]});
ixc_assign_3 _zz_strnp_3 ( ckv_ia_status[22:20], ckv_stat_code[2:0]);
ixc_assign_5 _zz_strnp_4 ( ckv_ia_status[19:15], ckv_stat_datawords[4:0]);
ixc_assign_15 _zz_strnp_5 ( ckv_ia_status[14:0], ckv_stat_addr[14:0]);
ixc_assign_64 _zz_strnp_6 ( ckv_wr_dat[63:0], { o_ckv_ia_wdata_part1[31], 
	o_ckv_ia_wdata_part1[30], o_ckv_ia_wdata_part1[29], 
	o_ckv_ia_wdata_part1[28], o_ckv_ia_wdata_part1[27], 
	o_ckv_ia_wdata_part1[26], o_ckv_ia_wdata_part1[25], 
	o_ckv_ia_wdata_part1[24], o_ckv_ia_wdata_part1[23], 
	o_ckv_ia_wdata_part1[22], o_ckv_ia_wdata_part1[21], 
	o_ckv_ia_wdata_part1[20], o_ckv_ia_wdata_part1[19], 
	o_ckv_ia_wdata_part1[18], o_ckv_ia_wdata_part1[17], 
	o_ckv_ia_wdata_part1[16], o_ckv_ia_wdata_part1[15], 
	o_ckv_ia_wdata_part1[14], o_ckv_ia_wdata_part1[13], 
	o_ckv_ia_wdata_part1[12], o_ckv_ia_wdata_part1[11], 
	o_ckv_ia_wdata_part1[10], o_ckv_ia_wdata_part1[9], 
	o_ckv_ia_wdata_part1[8], o_ckv_ia_wdata_part1[7], 
	o_ckv_ia_wdata_part1[6], o_ckv_ia_wdata_part1[5], 
	o_ckv_ia_wdata_part1[4], o_ckv_ia_wdata_part1[3], 
	o_ckv_ia_wdata_part1[2], o_ckv_ia_wdata_part1[1], 
	o_ckv_ia_wdata_part1[0], o_ckv_ia_wdata_part0[31], 
	o_ckv_ia_wdata_part0[30], o_ckv_ia_wdata_part0[29], 
	o_ckv_ia_wdata_part0[28], o_ckv_ia_wdata_part0[27], 
	o_ckv_ia_wdata_part0[26], o_ckv_ia_wdata_part0[25], 
	o_ckv_ia_wdata_part0[24], o_ckv_ia_wdata_part0[23], 
	o_ckv_ia_wdata_part0[22], o_ckv_ia_wdata_part0[21], 
	o_ckv_ia_wdata_part0[20], o_ckv_ia_wdata_part0[19], 
	o_ckv_ia_wdata_part0[18], o_ckv_ia_wdata_part0[17], 
	o_ckv_ia_wdata_part0[16], o_ckv_ia_wdata_part0[15], 
	o_ckv_ia_wdata_part0[14], o_ckv_ia_wdata_part0[13], 
	o_ckv_ia_wdata_part0[12], o_ckv_ia_wdata_part0[11], 
	o_ckv_ia_wdata_part0[10], o_ckv_ia_wdata_part0[9], 
	o_ckv_ia_wdata_part0[8], o_ckv_ia_wdata_part0[7], 
	o_ckv_ia_wdata_part0[6], o_ckv_ia_wdata_part0[5], 
	o_ckv_ia_wdata_part0[4], o_ckv_ia_wdata_part0[3], 
	o_ckv_ia_wdata_part0[2], o_ckv_ia_wdata_part0[1], 
	o_ckv_ia_wdata_part0[0]});
ixc_assign_4 _zz_strnp_7 ( kim_cmnd_op[3:0], o_kim_ia_config[17:14]);
ixc_assign_14 _zz_strnp_8 ( kim_cmnd_addr[13:0], o_kim_ia_config[13:0]);
ixc_assign_20 _zz_strnp_9 ( kim_ia_capability[19:0], { 
	kim_capability_type[3], kim_capability_type[2], 
	kim_capability_type[1], kim_capability_type[0], 
	kim_capability_lst[15], kim_capability_lst[14], 
	kim_capability_lst[13], kim_capability_lst[12], 
	kim_capability_lst[11], kim_capability_lst[10], 
	kim_capability_lst[9], kim_capability_lst[8], kim_capability_lst[7], 
	kim_capability_lst[6], kim_capability_lst[5], kim_capability_lst[4], 
	kim_capability_lst[3], kim_capability_lst[2], kim_capability_lst[1], 
	kim_capability_lst[0]});
ixc_assign_3 _zz_strnp_10 ( kim_ia_status[21:19], kim_stat_code[2:0]);
ixc_assign_5 _zz_strnp_11 ( kim_ia_status[18:14], kim_stat_datawords[4:0]);
ixc_assign_14 _zz_strnp_12 ( kim_ia_status[13:0], kim_stat_addr[13:0]);
ixc_assign_38 _zz_strnp_13 ( kim_wr_dat[37:0], { o_kim_ia_wdata_part0[20], 
	o_kim_ia_wdata_part0[19], o_kim_ia_wdata_part0[18], 
	o_kim_ia_wdata_part0[17], o_kim_ia_wdata_part0[16], 
	o_kim_ia_wdata_part0[15], o_kim_ia_wdata_part0[14], 
	o_kim_ia_wdata_part0[13], o_kim_ia_wdata_part0[12], 
	o_kim_ia_wdata_part0[11], o_kim_ia_wdata_part0[10], 
	o_kim_ia_wdata_part0[9], o_kim_ia_wdata_part0[8], 
	o_kim_ia_wdata_part0[7], o_kim_ia_wdata_part0[6], 
	o_kim_ia_wdata_part0[5], o_kim_ia_wdata_part0[4], 
	o_kim_ia_wdata_part0[3], o_kim_ia_wdata_part0[2], 
	o_kim_ia_wdata_part0[1], o_kim_ia_wdata_part0[0], 
	o_kim_ia_wdata_part1[16], o_kim_ia_wdata_part1[15], 
	o_kim_ia_wdata_part1[14], o_kim_ia_wdata_part1[13], 
	o_kim_ia_wdata_part1[12], o_kim_ia_wdata_part1[11], 
	o_kim_ia_wdata_part1[10], o_kim_ia_wdata_part1[9], 
	o_kim_ia_wdata_part1[8], o_kim_ia_wdata_part1[7], 
	o_kim_ia_wdata_part1[6], o_kim_ia_wdata_part1[5], 
	o_kim_ia_wdata_part1[4], o_kim_ia_wdata_part1[3], 
	o_kim_ia_wdata_part1[2], o_kim_ia_wdata_part1[1], 
	o_kim_ia_wdata_part1[0]});
ixc_assign _zz_strnp_14 ( cceip_encrypt_bimc_isync, cddip3_ism_osync);
ixc_assign _zz_strnp_15 ( cceip_encrypt_bimc_idat, cddip3_ism_odat);
ixc_assign _zz_strnp_16 ( cceip_validate_bimc_isync, cceip_encrypt_bimc_osync);
ixc_assign _zz_strnp_17 ( cceip_validate_bimc_idat, cceip_encrypt_bimc_odat);
ixc_assign _zz_strnp_18 ( cddip_decrypt_bimc_isync, cceip_validate_bimc_osync);
ixc_assign _zz_strnp_19 ( cddip_decrypt_bimc_idat, cceip_validate_bimc_odat);
ixc_assign _zz_strnp_20 ( axi_bimc_isync, cddip_decrypt_bimc_osync);
ixc_assign _zz_strnp_21 ( axi_bimc_idat, cddip_decrypt_bimc_odat);
ixc_assign _zz_strnp_22 ( axi_term_bimc_isync, axi_bimc_osync);
ixc_assign _zz_strnp_23 ( axi_term_bimc_idat, axi_bimc_odat);
ixc_assign_20 _zz_strnp_24 ( _zy_simnet_ckv_ia_capability_0_w$[0:19], 
	ckv_ia_capability[19:0]);
ixc_assign_23 _zz_strnp_25 ( _zy_simnet_ckv_ia_status_1_w$[0:22], 
	ckv_ia_status[22:0]);
ixc_assign_20 _zz_strnp_26 ( _zy_simnet_kim_ia_capability_2_w$[0:19], 
	kim_ia_capability[19:0]);
ixc_assign_22 _zz_strnp_27 ( _zy_simnet_kim_ia_status_3_w$[0:21], 
	kim_ia_status[21:0]);
ixc_assign_8 _zz_strnp_28 ( _zy_simnet_engine_sticky_status_4_w$[0:7], 
	engine_sticky_status[7:0]);
ixc_assign _zz_strnp_29 ( _zy_simnet_disable_ckv_kim_ism_reads_5_w$, 
	disable_ckv_kim_ism_reads);
ixc_assign _zz_strnp_30 ( _zy_simnet_send_kme_ib_beat_6_w$, send_kme_ib_beat);
ixc_assign _zz_strnp_31 ( _zy_simnet_debug_kme_ib_tvalid_7_w$, 
	send_kme_ib_beat);
ixc_assign _zz_strnp_32 ( _zy_simnet_debug_kme_ib_tlast_8_w$, 
	debug_kme_ib_tlast);
ixc_assign _zz_strnp_33 ( _zy_simnet_debug_kme_ib_tid_9_w$, 
	debug_kme_ib_tid[0]);
ixc_assign_8 _zz_strnp_34 ( _zy_simnet_debug_kme_ib_tstrb_10_w$[0:7], 
	debug_kme_ib_tstrb[7:0]);
ixc_assign_8 _zz_strnp_35 ( _zy_simnet_debug_kme_ib_tuser_11_w$[0:7], 
	debug_kme_ib_tuser[7:0]);
ixc_assign_64 _zz_strnp_36 ( _zy_simnet_debug_kme_ib_tdata_12_w$[0:63], 
	debug_kme_ib_tdata[63:0]);
ixc_assign_83 _zz_strnp_37 ( _zy_simnet_kme_cceip0_ob_out_13_w$[0:82], { 
	kme_cceip0_ob_out[82], kme_cceip0_ob_out_post[81], 
	kme_cceip0_ob_out_post[80], kme_cceip0_ob_out_post[79], 
	kme_cceip0_ob_out_post[78], kme_cceip0_ob_out_post[77], 
	kme_cceip0_ob_out_post[76], kme_cceip0_ob_out_post[75], 
	kme_cceip0_ob_out_post[74], kme_cceip0_ob_out_post[73], 
	kme_cceip0_ob_out_post[72], kme_cceip0_ob_out_post[71], 
	kme_cceip0_ob_out_post[70], kme_cceip0_ob_out_post[69], 
	kme_cceip0_ob_out_post[68], kme_cceip0_ob_out_post[67], 
	kme_cceip0_ob_out_post[66], kme_cceip0_ob_out_post[65], 
	kme_cceip0_ob_out_post[64], kme_cceip0_ob_out_post[63], 
	kme_cceip0_ob_out_post[62], kme_cceip0_ob_out_post[61], 
	kme_cceip0_ob_out_post[60], kme_cceip0_ob_out_post[59], 
	kme_cceip0_ob_out_post[58], kme_cceip0_ob_out_post[57], 
	kme_cceip0_ob_out_post[56], kme_cceip0_ob_out_post[55], 
	kme_cceip0_ob_out_post[54], kme_cceip0_ob_out_post[53], 
	kme_cceip0_ob_out_post[52], kme_cceip0_ob_out_post[51], 
	kme_cceip0_ob_out_post[50], kme_cceip0_ob_out_post[49], 
	kme_cceip0_ob_out_post[48], kme_cceip0_ob_out_post[47], 
	kme_cceip0_ob_out_post[46], kme_cceip0_ob_out_post[45], 
	kme_cceip0_ob_out_post[44], kme_cceip0_ob_out_post[43], 
	kme_cceip0_ob_out_post[42], kme_cceip0_ob_out_post[41], 
	kme_cceip0_ob_out_post[40], kme_cceip0_ob_out_post[39], 
	kme_cceip0_ob_out_post[38], kme_cceip0_ob_out_post[37], 
	kme_cceip0_ob_out_post[36], kme_cceip0_ob_out_post[35], 
	kme_cceip0_ob_out_post[34], kme_cceip0_ob_out_post[33], 
	kme_cceip0_ob_out_post[32], kme_cceip0_ob_out_post[31], 
	kme_cceip0_ob_out_post[30], kme_cceip0_ob_out_post[29], 
	kme_cceip0_ob_out_post[28], kme_cceip0_ob_out_post[27], 
	kme_cceip0_ob_out_post[26], kme_cceip0_ob_out_post[25], 
	kme_cceip0_ob_out_post[24], kme_cceip0_ob_out_post[23], 
	kme_cceip0_ob_out_post[22], kme_cceip0_ob_out_post[21], 
	kme_cceip0_ob_out_post[20], kme_cceip0_ob_out_post[19], 
	kme_cceip0_ob_out_post[18], kme_cceip0_ob_out_post[17], 
	kme_cceip0_ob_out_post[16], kme_cceip0_ob_out_post[15], 
	kme_cceip0_ob_out_post[14], kme_cceip0_ob_out_post[13], 
	kme_cceip0_ob_out_post[12], kme_cceip0_ob_out_post[11], 
	kme_cceip0_ob_out_post[10], kme_cceip0_ob_out_post[9], 
	kme_cceip0_ob_out_post[8], kme_cceip0_ob_out_post[7], 
	kme_cceip0_ob_out_post[6], kme_cceip0_ob_out_post[5], 
	kme_cceip0_ob_out_post[4], kme_cceip0_ob_out_post[3], 
	kme_cceip0_ob_out_post[2], kme_cceip0_ob_out_post[1], 
	kme_cceip0_ob_out_post[0]});
ixc_assign_83 _zz_strnp_38 ( _zy_simnet_kme_cceip1_ob_out_14_w$[0:82], { 
	kme_cceip1_ob_out[82], kme_cceip1_ob_out_post[81], 
	kme_cceip1_ob_out_post[80], kme_cceip1_ob_out_post[79], 
	kme_cceip1_ob_out_post[78], kme_cceip1_ob_out_post[77], 
	kme_cceip1_ob_out_post[76], kme_cceip1_ob_out_post[75], 
	kme_cceip1_ob_out_post[74], kme_cceip1_ob_out_post[73], 
	kme_cceip1_ob_out_post[72], kme_cceip1_ob_out_post[71], 
	kme_cceip1_ob_out_post[70], kme_cceip1_ob_out_post[69], 
	kme_cceip1_ob_out_post[68], kme_cceip1_ob_out_post[67], 
	kme_cceip1_ob_out_post[66], kme_cceip1_ob_out_post[65], 
	kme_cceip1_ob_out_post[64], kme_cceip1_ob_out_post[63], 
	kme_cceip1_ob_out_post[62], kme_cceip1_ob_out_post[61], 
	kme_cceip1_ob_out_post[60], kme_cceip1_ob_out_post[59], 
	kme_cceip1_ob_out_post[58], kme_cceip1_ob_out_post[57], 
	kme_cceip1_ob_out_post[56], kme_cceip1_ob_out_post[55], 
	kme_cceip1_ob_out_post[54], kme_cceip1_ob_out_post[53], 
	kme_cceip1_ob_out_post[52], kme_cceip1_ob_out_post[51], 
	kme_cceip1_ob_out_post[50], kme_cceip1_ob_out_post[49], 
	kme_cceip1_ob_out_post[48], kme_cceip1_ob_out_post[47], 
	kme_cceip1_ob_out_post[46], kme_cceip1_ob_out_post[45], 
	kme_cceip1_ob_out_post[44], kme_cceip1_ob_out_post[43], 
	kme_cceip1_ob_out_post[42], kme_cceip1_ob_out_post[41], 
	kme_cceip1_ob_out_post[40], kme_cceip1_ob_out_post[39], 
	kme_cceip1_ob_out_post[38], kme_cceip1_ob_out_post[37], 
	kme_cceip1_ob_out_post[36], kme_cceip1_ob_out_post[35], 
	kme_cceip1_ob_out_post[34], kme_cceip1_ob_out_post[33], 
	kme_cceip1_ob_out_post[32], kme_cceip1_ob_out_post[31], 
	kme_cceip1_ob_out_post[30], kme_cceip1_ob_out_post[29], 
	kme_cceip1_ob_out_post[28], kme_cceip1_ob_out_post[27], 
	kme_cceip1_ob_out_post[26], kme_cceip1_ob_out_post[25], 
	kme_cceip1_ob_out_post[24], kme_cceip1_ob_out_post[23], 
	kme_cceip1_ob_out_post[22], kme_cceip1_ob_out_post[21], 
	kme_cceip1_ob_out_post[20], kme_cceip1_ob_out_post[19], 
	kme_cceip1_ob_out_post[18], kme_cceip1_ob_out_post[17], 
	kme_cceip1_ob_out_post[16], kme_cceip1_ob_out_post[15], 
	kme_cceip1_ob_out_post[14], kme_cceip1_ob_out_post[13], 
	kme_cceip1_ob_out_post[12], kme_cceip1_ob_out_post[11], 
	kme_cceip1_ob_out_post[10], kme_cceip1_ob_out_post[9], 
	kme_cceip1_ob_out_post[8], kme_cceip1_ob_out_post[7], 
	kme_cceip1_ob_out_post[6], kme_cceip1_ob_out_post[5], 
	kme_cceip1_ob_out_post[4], kme_cceip1_ob_out_post[3], 
	kme_cceip1_ob_out_post[2], kme_cceip1_ob_out_post[1], 
	kme_cceip1_ob_out_post[0]});
ixc_assign_83 _zz_strnp_39 ( _zy_simnet_kme_cceip2_ob_out_15_w$[0:82], { 
	kme_cceip2_ob_out[82], kme_cceip2_ob_out_post[81], 
	kme_cceip2_ob_out_post[80], kme_cceip2_ob_out_post[79], 
	kme_cceip2_ob_out_post[78], kme_cceip2_ob_out_post[77], 
	kme_cceip2_ob_out_post[76], kme_cceip2_ob_out_post[75], 
	kme_cceip2_ob_out_post[74], kme_cceip2_ob_out_post[73], 
	kme_cceip2_ob_out_post[72], kme_cceip2_ob_out_post[71], 
	kme_cceip2_ob_out_post[70], kme_cceip2_ob_out_post[69], 
	kme_cceip2_ob_out_post[68], kme_cceip2_ob_out_post[67], 
	kme_cceip2_ob_out_post[66], kme_cceip2_ob_out_post[65], 
	kme_cceip2_ob_out_post[64], kme_cceip2_ob_out_post[63], 
	kme_cceip2_ob_out_post[62], kme_cceip2_ob_out_post[61], 
	kme_cceip2_ob_out_post[60], kme_cceip2_ob_out_post[59], 
	kme_cceip2_ob_out_post[58], kme_cceip2_ob_out_post[57], 
	kme_cceip2_ob_out_post[56], kme_cceip2_ob_out_post[55], 
	kme_cceip2_ob_out_post[54], kme_cceip2_ob_out_post[53], 
	kme_cceip2_ob_out_post[52], kme_cceip2_ob_out_post[51], 
	kme_cceip2_ob_out_post[50], kme_cceip2_ob_out_post[49], 
	kme_cceip2_ob_out_post[48], kme_cceip2_ob_out_post[47], 
	kme_cceip2_ob_out_post[46], kme_cceip2_ob_out_post[45], 
	kme_cceip2_ob_out_post[44], kme_cceip2_ob_out_post[43], 
	kme_cceip2_ob_out_post[42], kme_cceip2_ob_out_post[41], 
	kme_cceip2_ob_out_post[40], kme_cceip2_ob_out_post[39], 
	kme_cceip2_ob_out_post[38], kme_cceip2_ob_out_post[37], 
	kme_cceip2_ob_out_post[36], kme_cceip2_ob_out_post[35], 
	kme_cceip2_ob_out_post[34], kme_cceip2_ob_out_post[33], 
	kme_cceip2_ob_out_post[32], kme_cceip2_ob_out_post[31], 
	kme_cceip2_ob_out_post[30], kme_cceip2_ob_out_post[29], 
	kme_cceip2_ob_out_post[28], kme_cceip2_ob_out_post[27], 
	kme_cceip2_ob_out_post[26], kme_cceip2_ob_out_post[25], 
	kme_cceip2_ob_out_post[24], kme_cceip2_ob_out_post[23], 
	kme_cceip2_ob_out_post[22], kme_cceip2_ob_out_post[21], 
	kme_cceip2_ob_out_post[20], kme_cceip2_ob_out_post[19], 
	kme_cceip2_ob_out_post[18], kme_cceip2_ob_out_post[17], 
	kme_cceip2_ob_out_post[16], kme_cceip2_ob_out_post[15], 
	kme_cceip2_ob_out_post[14], kme_cceip2_ob_out_post[13], 
	kme_cceip2_ob_out_post[12], kme_cceip2_ob_out_post[11], 
	kme_cceip2_ob_out_post[10], kme_cceip2_ob_out_post[9], 
	kme_cceip2_ob_out_post[8], kme_cceip2_ob_out_post[7], 
	kme_cceip2_ob_out_post[6], kme_cceip2_ob_out_post[5], 
	kme_cceip2_ob_out_post[4], kme_cceip2_ob_out_post[3], 
	kme_cceip2_ob_out_post[2], kme_cceip2_ob_out_post[1], 
	kme_cceip2_ob_out_post[0]});
ixc_assign_83 _zz_strnp_40 ( _zy_simnet_kme_cceip3_ob_out_16_w$[0:82], { 
	kme_cceip3_ob_out[82], kme_cceip3_ob_out_post[81], 
	kme_cceip3_ob_out_post[80], kme_cceip3_ob_out_post[79], 
	kme_cceip3_ob_out_post[78], kme_cceip3_ob_out_post[77], 
	kme_cceip3_ob_out_post[76], kme_cceip3_ob_out_post[75], 
	kme_cceip3_ob_out_post[74], kme_cceip3_ob_out_post[73], 
	kme_cceip3_ob_out_post[72], kme_cceip3_ob_out_post[71], 
	kme_cceip3_ob_out_post[70], kme_cceip3_ob_out_post[69], 
	kme_cceip3_ob_out_post[68], kme_cceip3_ob_out_post[67], 
	kme_cceip3_ob_out_post[66], kme_cceip3_ob_out_post[65], 
	kme_cceip3_ob_out_post[64], kme_cceip3_ob_out_post[63], 
	kme_cceip3_ob_out_post[62], kme_cceip3_ob_out_post[61], 
	kme_cceip3_ob_out_post[60], kme_cceip3_ob_out_post[59], 
	kme_cceip3_ob_out_post[58], kme_cceip3_ob_out_post[57], 
	kme_cceip3_ob_out_post[56], kme_cceip3_ob_out_post[55], 
	kme_cceip3_ob_out_post[54], kme_cceip3_ob_out_post[53], 
	kme_cceip3_ob_out_post[52], kme_cceip3_ob_out_post[51], 
	kme_cceip3_ob_out_post[50], kme_cceip3_ob_out_post[49], 
	kme_cceip3_ob_out_post[48], kme_cceip3_ob_out_post[47], 
	kme_cceip3_ob_out_post[46], kme_cceip3_ob_out_post[45], 
	kme_cceip3_ob_out_post[44], kme_cceip3_ob_out_post[43], 
	kme_cceip3_ob_out_post[42], kme_cceip3_ob_out_post[41], 
	kme_cceip3_ob_out_post[40], kme_cceip3_ob_out_post[39], 
	kme_cceip3_ob_out_post[38], kme_cceip3_ob_out_post[37], 
	kme_cceip3_ob_out_post[36], kme_cceip3_ob_out_post[35], 
	kme_cceip3_ob_out_post[34], kme_cceip3_ob_out_post[33], 
	kme_cceip3_ob_out_post[32], kme_cceip3_ob_out_post[31], 
	kme_cceip3_ob_out_post[30], kme_cceip3_ob_out_post[29], 
	kme_cceip3_ob_out_post[28], kme_cceip3_ob_out_post[27], 
	kme_cceip3_ob_out_post[26], kme_cceip3_ob_out_post[25], 
	kme_cceip3_ob_out_post[24], kme_cceip3_ob_out_post[23], 
	kme_cceip3_ob_out_post[22], kme_cceip3_ob_out_post[21], 
	kme_cceip3_ob_out_post[20], kme_cceip3_ob_out_post[19], 
	kme_cceip3_ob_out_post[18], kme_cceip3_ob_out_post[17], 
	kme_cceip3_ob_out_post[16], kme_cceip3_ob_out_post[15], 
	kme_cceip3_ob_out_post[14], kme_cceip3_ob_out_post[13], 
	kme_cceip3_ob_out_post[12], kme_cceip3_ob_out_post[11], 
	kme_cceip3_ob_out_post[10], kme_cceip3_ob_out_post[9], 
	kme_cceip3_ob_out_post[8], kme_cceip3_ob_out_post[7], 
	kme_cceip3_ob_out_post[6], kme_cceip3_ob_out_post[5], 
	kme_cceip3_ob_out_post[4], kme_cceip3_ob_out_post[3], 
	kme_cceip3_ob_out_post[2], kme_cceip3_ob_out_post[1], 
	kme_cceip3_ob_out_post[0]});
ixc_assign_83 _zz_strnp_41 ( _zy_simnet_kme_cddip0_ob_out_17_w$[0:82], { 
	kme_cddip0_ob_out[82], kme_cddip0_ob_out_post[81], 
	kme_cddip0_ob_out_post[80], kme_cddip0_ob_out_post[79], 
	kme_cddip0_ob_out_post[78], kme_cddip0_ob_out_post[77], 
	kme_cddip0_ob_out_post[76], kme_cddip0_ob_out_post[75], 
	kme_cddip0_ob_out_post[74], kme_cddip0_ob_out_post[73], 
	kme_cddip0_ob_out_post[72], kme_cddip0_ob_out_post[71], 
	kme_cddip0_ob_out_post[70], kme_cddip0_ob_out_post[69], 
	kme_cddip0_ob_out_post[68], kme_cddip0_ob_out_post[67], 
	kme_cddip0_ob_out_post[66], kme_cddip0_ob_out_post[65], 
	kme_cddip0_ob_out_post[64], kme_cddip0_ob_out_post[63], 
	kme_cddip0_ob_out_post[62], kme_cddip0_ob_out_post[61], 
	kme_cddip0_ob_out_post[60], kme_cddip0_ob_out_post[59], 
	kme_cddip0_ob_out_post[58], kme_cddip0_ob_out_post[57], 
	kme_cddip0_ob_out_post[56], kme_cddip0_ob_out_post[55], 
	kme_cddip0_ob_out_post[54], kme_cddip0_ob_out_post[53], 
	kme_cddip0_ob_out_post[52], kme_cddip0_ob_out_post[51], 
	kme_cddip0_ob_out_post[50], kme_cddip0_ob_out_post[49], 
	kme_cddip0_ob_out_post[48], kme_cddip0_ob_out_post[47], 
	kme_cddip0_ob_out_post[46], kme_cddip0_ob_out_post[45], 
	kme_cddip0_ob_out_post[44], kme_cddip0_ob_out_post[43], 
	kme_cddip0_ob_out_post[42], kme_cddip0_ob_out_post[41], 
	kme_cddip0_ob_out_post[40], kme_cddip0_ob_out_post[39], 
	kme_cddip0_ob_out_post[38], kme_cddip0_ob_out_post[37], 
	kme_cddip0_ob_out_post[36], kme_cddip0_ob_out_post[35], 
	kme_cddip0_ob_out_post[34], kme_cddip0_ob_out_post[33], 
	kme_cddip0_ob_out_post[32], kme_cddip0_ob_out_post[31], 
	kme_cddip0_ob_out_post[30], kme_cddip0_ob_out_post[29], 
	kme_cddip0_ob_out_post[28], kme_cddip0_ob_out_post[27], 
	kme_cddip0_ob_out_post[26], kme_cddip0_ob_out_post[25], 
	kme_cddip0_ob_out_post[24], kme_cddip0_ob_out_post[23], 
	kme_cddip0_ob_out_post[22], kme_cddip0_ob_out_post[21], 
	kme_cddip0_ob_out_post[20], kme_cddip0_ob_out_post[19], 
	kme_cddip0_ob_out_post[18], kme_cddip0_ob_out_post[17], 
	kme_cddip0_ob_out_post[16], kme_cddip0_ob_out_post[15], 
	kme_cddip0_ob_out_post[14], kme_cddip0_ob_out_post[13], 
	kme_cddip0_ob_out_post[12], kme_cddip0_ob_out_post[11], 
	kme_cddip0_ob_out_post[10], kme_cddip0_ob_out_post[9], 
	kme_cddip0_ob_out_post[8], kme_cddip0_ob_out_post[7], 
	kme_cddip0_ob_out_post[6], kme_cddip0_ob_out_post[5], 
	kme_cddip0_ob_out_post[4], kme_cddip0_ob_out_post[3], 
	kme_cddip0_ob_out_post[2], kme_cddip0_ob_out_post[1], 
	kme_cddip0_ob_out_post[0]});
ixc_assign_83 _zz_strnp_42 ( _zy_simnet_kme_cddip1_ob_out_18_w$[0:82], { 
	kme_cddip1_ob_out[82], kme_cddip1_ob_out_post[81], 
	kme_cddip1_ob_out_post[80], kme_cddip1_ob_out_post[79], 
	kme_cddip1_ob_out_post[78], kme_cddip1_ob_out_post[77], 
	kme_cddip1_ob_out_post[76], kme_cddip1_ob_out_post[75], 
	kme_cddip1_ob_out_post[74], kme_cddip1_ob_out_post[73], 
	kme_cddip1_ob_out_post[72], kme_cddip1_ob_out_post[71], 
	kme_cddip1_ob_out_post[70], kme_cddip1_ob_out_post[69], 
	kme_cddip1_ob_out_post[68], kme_cddip1_ob_out_post[67], 
	kme_cddip1_ob_out_post[66], kme_cddip1_ob_out_post[65], 
	kme_cddip1_ob_out_post[64], kme_cddip1_ob_out_post[63], 
	kme_cddip1_ob_out_post[62], kme_cddip1_ob_out_post[61], 
	kme_cddip1_ob_out_post[60], kme_cddip1_ob_out_post[59], 
	kme_cddip1_ob_out_post[58], kme_cddip1_ob_out_post[57], 
	kme_cddip1_ob_out_post[56], kme_cddip1_ob_out_post[55], 
	kme_cddip1_ob_out_post[54], kme_cddip1_ob_out_post[53], 
	kme_cddip1_ob_out_post[52], kme_cddip1_ob_out_post[51], 
	kme_cddip1_ob_out_post[50], kme_cddip1_ob_out_post[49], 
	kme_cddip1_ob_out_post[48], kme_cddip1_ob_out_post[47], 
	kme_cddip1_ob_out_post[46], kme_cddip1_ob_out_post[45], 
	kme_cddip1_ob_out_post[44], kme_cddip1_ob_out_post[43], 
	kme_cddip1_ob_out_post[42], kme_cddip1_ob_out_post[41], 
	kme_cddip1_ob_out_post[40], kme_cddip1_ob_out_post[39], 
	kme_cddip1_ob_out_post[38], kme_cddip1_ob_out_post[37], 
	kme_cddip1_ob_out_post[36], kme_cddip1_ob_out_post[35], 
	kme_cddip1_ob_out_post[34], kme_cddip1_ob_out_post[33], 
	kme_cddip1_ob_out_post[32], kme_cddip1_ob_out_post[31], 
	kme_cddip1_ob_out_post[30], kme_cddip1_ob_out_post[29], 
	kme_cddip1_ob_out_post[28], kme_cddip1_ob_out_post[27], 
	kme_cddip1_ob_out_post[26], kme_cddip1_ob_out_post[25], 
	kme_cddip1_ob_out_post[24], kme_cddip1_ob_out_post[23], 
	kme_cddip1_ob_out_post[22], kme_cddip1_ob_out_post[21], 
	kme_cddip1_ob_out_post[20], kme_cddip1_ob_out_post[19], 
	kme_cddip1_ob_out_post[18], kme_cddip1_ob_out_post[17], 
	kme_cddip1_ob_out_post[16], kme_cddip1_ob_out_post[15], 
	kme_cddip1_ob_out_post[14], kme_cddip1_ob_out_post[13], 
	kme_cddip1_ob_out_post[12], kme_cddip1_ob_out_post[11], 
	kme_cddip1_ob_out_post[10], kme_cddip1_ob_out_post[9], 
	kme_cddip1_ob_out_post[8], kme_cddip1_ob_out_post[7], 
	kme_cddip1_ob_out_post[6], kme_cddip1_ob_out_post[5], 
	kme_cddip1_ob_out_post[4], kme_cddip1_ob_out_post[3], 
	kme_cddip1_ob_out_post[2], kme_cddip1_ob_out_post[1], 
	kme_cddip1_ob_out_post[0]});
ixc_assign_83 _zz_strnp_43 ( _zy_simnet_kme_cddip2_ob_out_19_w$[0:82], { 
	kme_cddip2_ob_out[82], kme_cddip2_ob_out_post[81], 
	kme_cddip2_ob_out_post[80], kme_cddip2_ob_out_post[79], 
	kme_cddip2_ob_out_post[78], kme_cddip2_ob_out_post[77], 
	kme_cddip2_ob_out_post[76], kme_cddip2_ob_out_post[75], 
	kme_cddip2_ob_out_post[74], kme_cddip2_ob_out_post[73], 
	kme_cddip2_ob_out_post[72], kme_cddip2_ob_out_post[71], 
	kme_cddip2_ob_out_post[70], kme_cddip2_ob_out_post[69], 
	kme_cddip2_ob_out_post[68], kme_cddip2_ob_out_post[67], 
	kme_cddip2_ob_out_post[66], kme_cddip2_ob_out_post[65], 
	kme_cddip2_ob_out_post[64], kme_cddip2_ob_out_post[63], 
	kme_cddip2_ob_out_post[62], kme_cddip2_ob_out_post[61], 
	kme_cddip2_ob_out_post[60], kme_cddip2_ob_out_post[59], 
	kme_cddip2_ob_out_post[58], kme_cddip2_ob_out_post[57], 
	kme_cddip2_ob_out_post[56], kme_cddip2_ob_out_post[55], 
	kme_cddip2_ob_out_post[54], kme_cddip2_ob_out_post[53], 
	kme_cddip2_ob_out_post[52], kme_cddip2_ob_out_post[51], 
	kme_cddip2_ob_out_post[50], kme_cddip2_ob_out_post[49], 
	kme_cddip2_ob_out_post[48], kme_cddip2_ob_out_post[47], 
	kme_cddip2_ob_out_post[46], kme_cddip2_ob_out_post[45], 
	kme_cddip2_ob_out_post[44], kme_cddip2_ob_out_post[43], 
	kme_cddip2_ob_out_post[42], kme_cddip2_ob_out_post[41], 
	kme_cddip2_ob_out_post[40], kme_cddip2_ob_out_post[39], 
	kme_cddip2_ob_out_post[38], kme_cddip2_ob_out_post[37], 
	kme_cddip2_ob_out_post[36], kme_cddip2_ob_out_post[35], 
	kme_cddip2_ob_out_post[34], kme_cddip2_ob_out_post[33], 
	kme_cddip2_ob_out_post[32], kme_cddip2_ob_out_post[31], 
	kme_cddip2_ob_out_post[30], kme_cddip2_ob_out_post[29], 
	kme_cddip2_ob_out_post[28], kme_cddip2_ob_out_post[27], 
	kme_cddip2_ob_out_post[26], kme_cddip2_ob_out_post[25], 
	kme_cddip2_ob_out_post[24], kme_cddip2_ob_out_post[23], 
	kme_cddip2_ob_out_post[22], kme_cddip2_ob_out_post[21], 
	kme_cddip2_ob_out_post[20], kme_cddip2_ob_out_post[19], 
	kme_cddip2_ob_out_post[18], kme_cddip2_ob_out_post[17], 
	kme_cddip2_ob_out_post[16], kme_cddip2_ob_out_post[15], 
	kme_cddip2_ob_out_post[14], kme_cddip2_ob_out_post[13], 
	kme_cddip2_ob_out_post[12], kme_cddip2_ob_out_post[11], 
	kme_cddip2_ob_out_post[10], kme_cddip2_ob_out_post[9], 
	kme_cddip2_ob_out_post[8], kme_cddip2_ob_out_post[7], 
	kme_cddip2_ob_out_post[6], kme_cddip2_ob_out_post[5], 
	kme_cddip2_ob_out_post[4], kme_cddip2_ob_out_post[3], 
	kme_cddip2_ob_out_post[2], kme_cddip2_ob_out_post[1], 
	kme_cddip2_ob_out_post[0]});
ixc_assign_83 _zz_strnp_44 ( _zy_simnet_kme_cddip3_ob_out_20_w$[0:82], { 
	kme_cddip3_ob_out[82], kme_cddip3_ob_out_post[81], 
	kme_cddip3_ob_out_post[80], kme_cddip3_ob_out_post[79], 
	kme_cddip3_ob_out_post[78], kme_cddip3_ob_out_post[77], 
	kme_cddip3_ob_out_post[76], kme_cddip3_ob_out_post[75], 
	kme_cddip3_ob_out_post[74], kme_cddip3_ob_out_post[73], 
	kme_cddip3_ob_out_post[72], kme_cddip3_ob_out_post[71], 
	kme_cddip3_ob_out_post[70], kme_cddip3_ob_out_post[69], 
	kme_cddip3_ob_out_post[68], kme_cddip3_ob_out_post[67], 
	kme_cddip3_ob_out_post[66], kme_cddip3_ob_out_post[65], 
	kme_cddip3_ob_out_post[64], kme_cddip3_ob_out_post[63], 
	kme_cddip3_ob_out_post[62], kme_cddip3_ob_out_post[61], 
	kme_cddip3_ob_out_post[60], kme_cddip3_ob_out_post[59], 
	kme_cddip3_ob_out_post[58], kme_cddip3_ob_out_post[57], 
	kme_cddip3_ob_out_post[56], kme_cddip3_ob_out_post[55], 
	kme_cddip3_ob_out_post[54], kme_cddip3_ob_out_post[53], 
	kme_cddip3_ob_out_post[52], kme_cddip3_ob_out_post[51], 
	kme_cddip3_ob_out_post[50], kme_cddip3_ob_out_post[49], 
	kme_cddip3_ob_out_post[48], kme_cddip3_ob_out_post[47], 
	kme_cddip3_ob_out_post[46], kme_cddip3_ob_out_post[45], 
	kme_cddip3_ob_out_post[44], kme_cddip3_ob_out_post[43], 
	kme_cddip3_ob_out_post[42], kme_cddip3_ob_out_post[41], 
	kme_cddip3_ob_out_post[40], kme_cddip3_ob_out_post[39], 
	kme_cddip3_ob_out_post[38], kme_cddip3_ob_out_post[37], 
	kme_cddip3_ob_out_post[36], kme_cddip3_ob_out_post[35], 
	kme_cddip3_ob_out_post[34], kme_cddip3_ob_out_post[33], 
	kme_cddip3_ob_out_post[32], kme_cddip3_ob_out_post[31], 
	kme_cddip3_ob_out_post[30], kme_cddip3_ob_out_post[29], 
	kme_cddip3_ob_out_post[28], kme_cddip3_ob_out_post[27], 
	kme_cddip3_ob_out_post[26], kme_cddip3_ob_out_post[25], 
	kme_cddip3_ob_out_post[24], kme_cddip3_ob_out_post[23], 
	kme_cddip3_ob_out_post[22], kme_cddip3_ob_out_post[21], 
	kme_cddip3_ob_out_post[20], kme_cddip3_ob_out_post[19], 
	kme_cddip3_ob_out_post[18], kme_cddip3_ob_out_post[17], 
	kme_cddip3_ob_out_post[16], kme_cddip3_ob_out_post[15], 
	kme_cddip3_ob_out_post[14], kme_cddip3_ob_out_post[13], 
	kme_cddip3_ob_out_post[12], kme_cddip3_ob_out_post[11], 
	kme_cddip3_ob_out_post[10], kme_cddip3_ob_out_post[9], 
	kme_cddip3_ob_out_post[8], kme_cddip3_ob_out_post[7], 
	kme_cddip3_ob_out_post[6], kme_cddip3_ob_out_post[5], 
	kme_cddip3_ob_out_post[4], kme_cddip3_ob_out_post[3], 
	kme_cddip3_ob_out_post[2], kme_cddip3_ob_out_post[1], 
	kme_cddip3_ob_out_post[0]});
Q_INV U949 ( .A(n44), .Z(n56));
Q_FDP4EP \engine_sticky_status_REG[7] ( .CK(clk), .CE(n56), .R(n57), .D(n29), .Q(engine_sticky_status[7]));
Q_INV U951 ( .A(rst_n), .Z(n57));
Q_INV U952 ( .A(n43), .Z(n58));
Q_FDP4EP \engine_sticky_status_REG[6] ( .CK(clk), .CE(n58), .R(n57), .D(n30), .Q(engine_sticky_status[6]));
Q_INV U954 ( .A(n42), .Z(n59));
Q_FDP4EP \engine_sticky_status_REG[5] ( .CK(clk), .CE(n59), .R(n57), .D(n31), .Q(engine_sticky_status[5]));
Q_INV U956 ( .A(n41), .Z(n60));
Q_FDP4EP \engine_sticky_status_REG[4] ( .CK(clk), .CE(n60), .R(n57), .D(n32), .Q(engine_sticky_status[4]));
Q_INV U958 ( .A(n40), .Z(n61));
Q_FDP4EP \engine_sticky_status_REG[3] ( .CK(clk), .CE(n61), .R(n57), .D(n33), .Q(engine_sticky_status[3]));
Q_INV U960 ( .A(n39), .Z(n62));
Q_FDP4EP \engine_sticky_status_REG[2] ( .CK(clk), .CE(n62), .R(n57), .D(n34), .Q(engine_sticky_status[2]));
Q_INV U962 ( .A(n38), .Z(n63));
Q_FDP4EP \engine_sticky_status_REG[1] ( .CK(clk), .CE(n63), .R(n57), .D(n35), .Q(engine_sticky_status[1]));
Q_INV U964 ( .A(n37), .Z(n64));
Q_FDP4EP \engine_sticky_status_REG[0] ( .CK(clk), .CE(n64), .R(n57), .D(n36), .Q(engine_sticky_status[0]));
Q_INV U966 ( .A(n12), .Z(n65));
Q_INV U967 ( .A(send_kme_ib_beat), .Z(n66));
Q_FDP4EP send_kme_ib_beat_REG  ( .CK(clk), .CE(n65), .R(n57), .D(n66), .Q(send_kme_ib_beat));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "\ckv_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "\ckv_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m3 "\ckv_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m4 "\ckv_ia_status.r.part0  (1,0) 1 22 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m5 "\ckv_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m6 "\ckv_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m7 "\ckv_ia_status.f.addr  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m8 "\kim_ia_capability.r.part0  (1,0) 1 19 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m9 "\kim_ia_capability.f.mem_type  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m10 "\kim_ia_capability.f.reserved_op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m11 "\kim_ia_status.r.part0  (1,0) 1 21 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m12 "\kim_ia_status.f.code  (1,0) 1 2 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m13 "\kim_ia_status.f.datawords  (1,0) 1 4 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m14 "\kim_ia_status.f.addr  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m15 "\kme_cceip0_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m16 "\kme_cceip0_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m17 "\kme_cceip0_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m18 "\kme_cceip0_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m19 "\kme_cceip1_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m20 "\kme_cceip1_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m21 "\kme_cceip1_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m22 "\kme_cceip1_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m23 "\kme_cceip2_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m24 "\kme_cceip2_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m25 "\kme_cceip2_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m26 "\kme_cceip2_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m27 "\kme_cceip3_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m28 "\kme_cceip3_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m29 "\kme_cceip3_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m30 "\kme_cceip3_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m31 "\kme_cddip0_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m32 "\kme_cddip0_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m33 "\kme_cddip0_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m34 "\kme_cddip0_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m35 "\kme_cddip1_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m36 "\kme_cddip1_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m37 "\kme_cddip1_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m38 "\kme_cddip1_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m39 "\kme_cddip2_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m40 "\kme_cddip2_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m41 "\kme_cddip2_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m42 "\kme_cddip2_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m43 "\kme_cddip3_ob_out.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m44 "\kme_cddip3_ob_out.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m45 "\kme_cddip3_ob_out.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m46 "\kme_cddip3_ob_out.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m47 "\o_ckv_ia_config.r.part0  (1,0) 1 18 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m48 "\o_ckv_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m49 "\o_ckv_ia_config.f.addr  (1,0) 1 14 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m50 "\o_kim_ia_config.r.part0  (1,0) 1 17 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m51 "\o_kim_ia_config.f.op  (1,0) 1 3 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m52 "\o_kim_ia_config.f.addr  (1,0) 1 13 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m53 "\cceip0_out_ia_wdata.r.part2  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m54 "\cceip0_out_ia_wdata.r.part1  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m55 "\cceip0_out_ia_wdata.r.part0  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m56 "\cceip0_out_ia_wdata.f.tdata_hi  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m57 "\cceip0_out_ia_wdata.f.tdata_lo  (1,0) 1 31 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m58 "\cceip0_out_ia_wdata.f.bytes_vld  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m59 "\cceip0_out_ia_wdata.f.unused1  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m60 "\cceip0_out_ia_wdata.f.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m61 "\cceip0_out_ia_wdata.f.unused0  (1,0) 1 5 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m62 "\tready_override.r.part0  (1,0) 1 8 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m63 "\kme_cceip0_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m64 "\kme_cceip0_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m65 "\kme_cceip0_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m66 "\kme_cceip0_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m67 "\kme_cceip1_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m68 "\kme_cceip1_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m69 "\kme_cceip1_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m70 "\kme_cceip1_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m71 "\kme_cceip2_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m72 "\kme_cceip2_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m73 "\kme_cceip2_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m74 "\kme_cceip2_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m75 "\kme_cceip3_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m76 "\kme_cceip3_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m77 "\kme_cceip3_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m78 "\kme_cceip3_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m79 "\kme_cddip0_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m80 "\kme_cddip0_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m81 "\kme_cddip0_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m82 "\kme_cddip0_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m83 "\kme_cddip1_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m84 "\kme_cddip1_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m85 "\kme_cddip1_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m86 "\kme_cddip1_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m87 "\kme_cddip2_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m88 "\kme_cddip2_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m89 "\kme_cddip2_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m90 "\kme_cddip2_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m91 "\kme_cddip3_ob_out_post.tid  (1,0) 1 0 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m92 "\kme_cddip3_ob_out_post.tstrb  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m93 "\kme_cddip3_ob_out_post.tuser  (1,0) 1 7 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m94 "\kme_cddip3_ob_out_post.tdata  (1,0) 1 63 0 -2147483648 -2147483648"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "94"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r1 "ckv_ia_capability 2 \ckv_ia_capability.r  { \ckv_ia_capability.r.part0  } \ckv_ia_capability.f  { \ckv_ia_capability.f.mem_type  \ckv_ia_capability.f.ack_error  \ckv_ia_capability.f.sim_tmo  \ckv_ia_capability.f.reserved_op  \ckv_ia_capability.f.compare  \ckv_ia_capability.f.set_init_start  \ckv_ia_capability.f.initialize_inc  \ckv_ia_capability.f.initialize  \ckv_ia_capability.f.reset  \ckv_ia_capability.f.disabled  \ckv_ia_capability.f.enable  \ckv_ia_capability.f.write  \ckv_ia_capability.f.read  \ckv_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r2 "ckv_ia_status 2 \ckv_ia_status.r  { \ckv_ia_status.r.part0  } \ckv_ia_status.f  { \ckv_ia_status.f.code  \ckv_ia_status.f.datawords  \ckv_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r3 "kim_ia_capability 2 \kim_ia_capability.r  { \kim_ia_capability.r.part0  } \kim_ia_capability.f  { \kim_ia_capability.f.mem_type  \kim_ia_capability.f.ack_error  \kim_ia_capability.f.sim_tmo  \kim_ia_capability.f.reserved_op  \kim_ia_capability.f.compare  \kim_ia_capability.f.set_init_start  \kim_ia_capability.f.initialize_inc  \kim_ia_capability.f.initialize  \kim_ia_capability.f.reset  \kim_ia_capability.f.disabled  \kim_ia_capability.f.enable  \kim_ia_capability.f.write  \kim_ia_capability.f.read  \kim_ia_capability.f.nop  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r4 "kim_ia_status 2 \kim_ia_status.r  { \kim_ia_status.r.part0  } \kim_ia_status.f  { \kim_ia_status.f.code  \kim_ia_status.f.datawords  \kim_ia_status.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r1 "kme_cceip0_ob_out 6 \kme_cceip0_ob_out.tvalid  \kme_cceip0_ob_out.tlast  \kme_cceip0_ob_out.tid  \kme_cceip0_ob_out.tstrb  \kme_cceip0_ob_out.tuser  \kme_cceip0_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r2 "kme_cceip1_ob_out 6 \kme_cceip1_ob_out.tvalid  \kme_cceip1_ob_out.tlast  \kme_cceip1_ob_out.tid  \kme_cceip1_ob_out.tstrb  \kme_cceip1_ob_out.tuser  \kme_cceip1_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r3 "kme_cceip2_ob_out 6 \kme_cceip2_ob_out.tvalid  \kme_cceip2_ob_out.tlast  \kme_cceip2_ob_out.tid  \kme_cceip2_ob_out.tstrb  \kme_cceip2_ob_out.tuser  \kme_cceip2_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r4 "kme_cceip3_ob_out 6 \kme_cceip3_ob_out.tvalid  \kme_cceip3_ob_out.tlast  \kme_cceip3_ob_out.tid  \kme_cceip3_ob_out.tstrb  \kme_cceip3_ob_out.tuser  \kme_cceip3_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r5 "kme_cddip0_ob_out 6 \kme_cddip0_ob_out.tvalid  \kme_cddip0_ob_out.tlast  \kme_cddip0_ob_out.tid  \kme_cddip0_ob_out.tstrb  \kme_cddip0_ob_out.tuser  \kme_cddip0_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r6 "kme_cddip1_ob_out 6 \kme_cddip1_ob_out.tvalid  \kme_cddip1_ob_out.tlast  \kme_cddip1_ob_out.tid  \kme_cddip1_ob_out.tstrb  \kme_cddip1_ob_out.tuser  \kme_cddip1_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r7 "kme_cddip2_ob_out 6 \kme_cddip2_ob_out.tvalid  \kme_cddip2_ob_out.tlast  \kme_cddip2_ob_out.tid  \kme_cddip2_ob_out.tstrb  \kme_cddip2_ob_out.tuser  \kme_cddip2_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r8 "kme_cddip3_ob_out 6 \kme_cddip3_ob_out.tvalid  \kme_cddip3_ob_out.tlast  \kme_cddip3_ob_out.tid  \kme_cddip3_ob_out.tstrb  \kme_cddip3_ob_out.tuser  \kme_cddip3_ob_out.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r5 "o_ckv_ia_config 2 \o_ckv_ia_config.r  { \o_ckv_ia_config.r.part0  } \o_ckv_ia_config.f  { \o_ckv_ia_config.f.op  \o_ckv_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r6 "o_kim_ia_config 2 \o_kim_ia_config.r  { \o_kim_ia_config.r.part0  } \o_kim_ia_config.f  { \o_kim_ia_config.f.op  \o_kim_ia_config.f.addr  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r7 "cceip0_out_ia_wdata 2 \cceip0_out_ia_wdata.r  { \cceip0_out_ia_wdata.r.part2  \cceip0_out_ia_wdata.r.part1  \cceip0_out_ia_wdata.r.part0  } \cceip0_out_ia_wdata.f  { \cceip0_out_ia_wdata.f.tdata_hi  \cceip0_out_ia_wdata.f.tdata_lo  \cceip0_out_ia_wdata.f.eob  \cceip0_out_ia_wdata.f.bytes_vld  \cceip0_out_ia_wdata.f.unused1  \cceip0_out_ia_wdata.f.tid  \cceip0_out_ia_wdata.f.tuser  \cceip0_out_ia_wdata.f.unused0  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_r8 "tready_override 2 \tready_override.r  { \tready_override.r.part0  } \tready_override.f  { \tready_override.f.txc_tready_override  \tready_override.f.engine_7_tready_override  \tready_override.f.engine_6_tready_override  \tready_override.f.engine_5_tready_override  \tready_override.f.engine_4_tready_override  \tready_override.f.engine_3_tready_override  \tready_override.f.engine_2_tready_override  \tready_override.f.engine_1_tready_override  \tready_override.f.engine_0_tready_override  }"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r9 "kme_cceip0_ob_out_post 6 \kme_cceip0_ob_out_post.tvalid  \kme_cceip0_ob_out_post.tlast  \kme_cceip0_ob_out_post.tid  \kme_cceip0_ob_out_post.tstrb  \kme_cceip0_ob_out_post.tuser  \kme_cceip0_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r10 "kme_cceip1_ob_out_post 6 \kme_cceip1_ob_out_post.tvalid  \kme_cceip1_ob_out_post.tlast  \kme_cceip1_ob_out_post.tid  \kme_cceip1_ob_out_post.tstrb  \kme_cceip1_ob_out_post.tuser  \kme_cceip1_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r11 "kme_cceip2_ob_out_post 6 \kme_cceip2_ob_out_post.tvalid  \kme_cceip2_ob_out_post.tlast  \kme_cceip2_ob_out_post.tid  \kme_cceip2_ob_out_post.tstrb  \kme_cceip2_ob_out_post.tuser  \kme_cceip2_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r12 "kme_cceip3_ob_out_post 6 \kme_cceip3_ob_out_post.tvalid  \kme_cceip3_ob_out_post.tlast  \kme_cceip3_ob_out_post.tid  \kme_cceip3_ob_out_post.tstrb  \kme_cceip3_ob_out_post.tuser  \kme_cceip3_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r13 "kme_cddip0_ob_out_post 6 \kme_cddip0_ob_out_post.tvalid  \kme_cddip0_ob_out_post.tlast  \kme_cddip0_ob_out_post.tid  \kme_cddip0_ob_out_post.tstrb  \kme_cddip0_ob_out_post.tuser  \kme_cddip0_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r14 "kme_cddip1_ob_out_post 6 \kme_cddip1_ob_out_post.tvalid  \kme_cddip1_ob_out_post.tlast  \kme_cddip1_ob_out_post.tid  \kme_cddip1_ob_out_post.tstrb  \kme_cddip1_ob_out_post.tuser  \kme_cddip1_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r15 "kme_cddip2_ob_out_post 6 \kme_cddip2_ob_out_post.tvalid  \kme_cddip2_ob_out_post.tlast  \kme_cddip2_ob_out_post.tid  \kme_cddip2_ob_out_post.tstrb  \kme_cddip2_ob_out_post.tuser  \kme_cddip2_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_r16 "kme_cddip3_ob_out_post 6 \kme_cddip3_ob_out_post.tvalid  \kme_cddip3_ob_out_post.tlast  \kme_cddip3_ob_out_post.tid  \kme_cddip3_ob_out_post.tstrb  \kme_cddip3_ob_out_post.tuser  \kme_cddip3_ob_out_post.tdata "
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_NUM "16"
// pragma CVASTRPROP MODULE HDLICE HDL_RECORD_PACKED_UNION_NUM "8"
endmodule
