
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module bimc_master ( bimc_ecc_error, bimc_interrupt, bimc_odat, bimc_osync, 
	bimc_rst_n, clk, rst_n, bimc_idat, bimc_isync, o_bimc_monitor_mask, 
	o_bimc_ecc_uncorrectable_error_cnt, o_bimc_ecc_correctable_error_cnt, 
	o_bimc_parity_error_cnt, o_bimc_global_config, o_bimc_eccpar_debug, 
	o_bimc_cmd2, o_bimc_cmd1, o_bimc_cmd0, o_bimc_rxcmd2, o_bimc_rxrsp2, 
	o_bimc_pollrsp2, o_bimc_dbgcmd2, i_bimc_monitor, 
	i_bimc_ecc_uncorrectable_error_cnt, i_bimc_ecc_correctable_error_cnt, 
	i_bimc_parity_error_cnt, i_bimc_global_config, i_bimc_memid, 
	i_bimc_eccpar_debug, i_bimc_cmd2, i_bimc_rxcmd2, i_bimc_rxcmd1, 
	i_bimc_rxcmd0, i_bimc_rxrsp2, i_bimc_rxrsp1, i_bimc_rxrsp0, 
	i_bimc_pollrsp2, i_bimc_pollrsp1, i_bimc_pollrsp0, i_bimc_dbgcmd2, 
	i_bimc_dbgcmd1, i_bimc_dbgcmd0);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output bimc_ecc_error;
output bimc_interrupt;
output bimc_odat;
output bimc_osync;
output bimc_rst_n;
input clk;
input rst_n;
input bimc_idat;
input bimc_isync;
input [6:0] o_bimc_monitor_mask;
input [31:0] o_bimc_ecc_uncorrectable_error_cnt;
input [31:0] o_bimc_ecc_correctable_error_cnt;
input [31:0] o_bimc_parity_error_cnt;
input [31:0] o_bimc_global_config;
input [28:0] o_bimc_eccpar_debug;
input [10:0] o_bimc_cmd2;
input [31:0] o_bimc_cmd1;
input [31:0] o_bimc_cmd0;
input [9:0] o_bimc_rxcmd2;
input [9:0] o_bimc_rxrsp2;
input [9:0] o_bimc_pollrsp2;
input [9:0] o_bimc_dbgcmd2;
output [6:0] i_bimc_monitor;
output [31:0] i_bimc_ecc_uncorrectable_error_cnt;
output [31:0] i_bimc_ecc_correctable_error_cnt;
output [31:0] i_bimc_parity_error_cnt;
output [31:0] i_bimc_global_config;
output [11:0] i_bimc_memid;
output [28:0] i_bimc_eccpar_debug;
output [10:0] i_bimc_cmd2;
output [9:0] i_bimc_rxcmd2;
output [31:0] i_bimc_rxcmd1;
output [31:0] i_bimc_rxcmd0;
output [9:0] i_bimc_rxrsp2;
output [31:0] i_bimc_rxrsp1;
output [31:0] i_bimc_rxrsp0;
output [9:0] i_bimc_pollrsp2;
output [31:0] i_bimc_pollrsp1;
output [31:0] i_bimc_pollrsp0;
output [9:0] i_bimc_dbgcmd2;
output [31:0] i_bimc_dbgcmd1;
output [31:0] i_bimc_dbgcmd0;
wire [1:0] bimc_eccpar_debug_eccpar_corrupt;
wire [1:0] bimc_eccpar_debug_eccpar_disable;
wire [3:0] bimc_eccpar_debug_jabber_off;
wire [11:0] bimc_eccpar_debug_memaddr;
wire [3:0] bimc_eccpar_debug_memtype;
wire bimc_eccpar_debug_write_notify_ev;
wire bimc_global_config_poll_ecc_par_error;
wire [25:0] bimc_global_config_poll_ecc_par_timer;
wire bimc_global_config_mem_wr_init;
wire [31:0] bimc_cmd0_data;
wire [15:0] bimc_cmd1_addr;
wire [11:0] bimc_cmd1_mem;
wire [3:0] bimc_cmd1_memtype;
wire [7:0] bimc_cmd2_opcode;
wire bimc_cmd2_write_notify_ev;
wire bimc_ecc_error_c;
wire bimc_interrupt_c;
wire bimc_global_config_soft_reset;
wire [71:0] rcv_dat;
wire rcv_resp;
wire rcv_frm;
wire rcv_chk;
wire [3:0] bm_type;
wire [7:0] bm_op;
wire [11:0] bm_mem;
wire [15:0] bm_addr;
wire [31:0] bm_dat;
wire new_frame;
wire [103:0] rstate_text;
wire [72:0] cputx_frame;
wire [95:0] tstate_text;
wire _zy_simnet_bimc_ecc_error_0_w$;
wire _zy_simnet_bimc_interrupt_1_w$;
wire _zy_simnet_bimc_odat_2_w$;
wire _zy_simnet_bimc_osync_3_w$;
wire _zy_simnet_bimc_rst_n_4_w$;
wire bimc_monitor_uncorrectable_ecc_error_din;
wire bimc_monitor_correctable_ecc_error_din;
wire bimc_monitor_parity_error_din;
wire bimc_monitor_bimc_chain_rcv_error_din;
wire bimc_monitor_rcv_invalid_opcode_din;
wire bimc_monitor_unanswered_read_din;
wire bimc_ecc_uncorrectable_error_cnt_uncorrectable_ecc_en;
wire bimc_ecc_correctable_error_cnt_correctable_ecc_en;
wire bimc_parity_error_cnt_parity_errors_en;
wire debug_write_en;
wire [11:0] number_of_memories;
wire bimc_eccpar_debug_send;
wire [2:0] r_bimc_eccpar_debug_write_notify_ev;
wire bimc_eccpar_debug_sent_din;
wire bimc_eccpar_debug_sent;
wire bimc_cmd2_send;
wire [2:0] r_bimc_cmd2_write_notify_ev;
wire bimc_cmd2_sent_din;
wire bimc_rxrsp2_rxflag_din;
wire [31:0] bimc_rxrsp0_data_din;
wire [31:0] bimc_rxrsp1_data_din;
wire [7:0] bimc_rxrsp2_data_din;
wire bimc_pollrsp2_rxflag_din;
wire [31:0] bimc_pollrsp0_data_din;
wire [31:0] bimc_pollrsp1_data_din;
wire [7:0] bimc_pollrsp2_data_din;
wire bimc_rxcmd2_rxflag_din;
wire [31:0] bimc_rxcmd0_data_din;
wire [15:0] bimc_rxcmd1_addr_din;
wire [11:0] bimc_rxcmd1_mem_din;
wire [3:0] bimc_rxcmd1_memtype_din;
wire [7:0] bimc_rxcmd2_opcode_din;
wire bimc_dbgcmd2_rxflag_din;
wire [31:0] bimc_dbgcmd0_data_din;
wire [15:0] bimc_dbgcmd1_addr_din;
wire [11:0] bimc_dbgcmd1_mem_din;
wire [3:0] bimc_dbgcmd1_memtype_din;
wire [7:0] bimc_dbgcmd2_opcode_din;
wire bimc_cmd2_sent;
wire [31:0] bimc_ecc_uncorrectable_error_cnt;
wire [31:0] bimc_ecc_correctable_error_cnt;
wire [31:0] bimc_parity_error_cnt;
wire [71:0] bimc_rdat;
wire [71:0] bimc_dat;
wire bimc_frm;
wire bimc_chk;
wire [3:0] rx_type;
wire [7:0] rx_op;
wire [11:0] rx_mem;
wire [15:0] rx_addr;
wire [31:0] rx_dat;
wire rx_resp;
wire rx_frm;
wire [1:0] rx_chk;
wire bm_resp;
wire [6:0] bm_cnt;
wire [3:0] rstate;
wire [3:0] nxt_rstate;
wire [3:0] tstate;
wire [3:0] nxt_tstate;
wire bimc_global_config_bimc_mem_init_done_din;
wire [6:0] sync_cnt;
wire cmd_cnt;
wire mem_wr_init_dly;
wire mem_wr_init_ev;
wire eccpar_debug_ev;
wire cpu_transmit_ev;
wire [72:0] reg_send;
wire [72:0] r_reg_send;
wire [3:0] cputx_type;
wire [7:0] cputx_op;
wire [11:0] cputx_mem;
wire [15:0] cputx_addr;
wire [31:0] cputx_dat;
wire auto_poll_ecc_par_ev;
wire [25:0] poll_ecc_par_timer;
supply1 n1;
supply0 n2;
supply0 n1318;
Q_BUF U0 ( .A(n2), .Z(rstate_text[4]));
Q_BUF U1 ( .A(n1), .Z(rstate_text[2]));
Q_BUF U2 ( .A(n2), .Z(tstate_text[7]));
Q_BUF U3 ( .A(n1), .Z(tstate_text[2]));
Q_BUF U4 ( .A(n2), .Z(i_bimc_monitor[3]));
Q_BUF U5 ( .A(n1), .Z(tstate_text[6]));
Q_BUF U6 ( .A(n1), .Z(tstate_text[14]));
Q_BUF U7 ( .A(n1), .Z(tstate_text[22]));
Q_BUF U8 ( .A(n2), .Z(tstate_text[15]));
Q_BUF U9 ( .A(n2), .Z(tstate_text[23]));
Q_BUF U10 ( .A(n2), .Z(tstate_text[31]));
Q_BUF U11 ( .A(n2), .Z(tstate_text[39]));
Q_BUF U12 ( .A(n2), .Z(tstate_text[47]));
Q_BUF U13 ( .A(n2), .Z(tstate_text[55]));
Q_BUF U14 ( .A(n2), .Z(tstate_text[57]));
Q_BUF U15 ( .A(n2), .Z(tstate_text[59]));
Q_BUF U16 ( .A(n2), .Z(tstate_text[63]));
Q_BUF U17 ( .A(n2), .Z(tstate_text[65]));
Q_BUF U18 ( .A(n2), .Z(tstate_text[71]));
Q_BUF U19 ( .A(n2), .Z(tstate_text[74]));
Q_BUF U20 ( .A(n2), .Z(tstate_text[75]));
Q_BUF U21 ( .A(n2), .Z(tstate_text[76]));
Q_BUF U22 ( .A(n2), .Z(tstate_text[79]));
Q_BUF U23 ( .A(n2), .Z(tstate_text[82]));
Q_BUF U24 ( .A(n2), .Z(tstate_text[83]));
Q_BUF U25 ( .A(n2), .Z(tstate_text[84]));
Q_BUF U26 ( .A(n2), .Z(tstate_text[87]));
Q_BUF U27 ( .A(n2), .Z(tstate_text[89]));
Q_BUF U28 ( .A(n2), .Z(tstate_text[91]));
Q_BUF U29 ( .A(n2), .Z(tstate_text[92]));
Q_BUF U30 ( .A(n2), .Z(tstate_text[95]));
Q_BUF U31 ( .A(n1), .Z(rstate_text[6]));
Q_BUF U32 ( .A(n1), .Z(rstate_text[10]));
Q_BUF U33 ( .A(n1), .Z(rstate_text[14]));
Q_BUF U34 ( .A(n1), .Z(rstate_text[22]));
Q_BUF U35 ( .A(n1), .Z(rstate_text[30]));
Q_BUF U36 ( .A(n2), .Z(rstate_text[7]));
Q_BUF U37 ( .A(n2), .Z(rstate_text[15]));
Q_BUF U38 ( .A(n2), .Z(rstate_text[20]));
Q_BUF U39 ( .A(n2), .Z(rstate_text[23]));
Q_BUF U40 ( .A(n2), .Z(rstate_text[31]));
Q_BUF U41 ( .A(n2), .Z(rstate_text[39]));
Q_BUF U42 ( .A(n2), .Z(rstate_text[47]));
Q_BUF U43 ( .A(n2), .Z(rstate_text[55]));
Q_BUF U44 ( .A(n2), .Z(rstate_text[63]));
Q_BUF U45 ( .A(n2), .Z(rstate_text[71]));
Q_BUF U46 ( .A(n2), .Z(rstate_text[79]));
Q_BUF U47 ( .A(n2), .Z(rstate_text[87]));
Q_BUF U48 ( .A(n2), .Z(rstate_text[95]));
Q_BUF U49 ( .A(n2), .Z(rstate_text[96]));
Q_BUF U50 ( .A(n2), .Z(rstate_text[98]));
Q_BUF U51 ( .A(n2), .Z(rstate_text[99]));
Q_BUF U52 ( .A(n2), .Z(rstate_text[103]));
Q_BUF U53 ( .A(rstate_text[100]), .Z(rstate_text[102]));
Q_BUF U54 ( .A(rstate_text[90]), .Z(rstate_text[100]));
Q_BUF U55 ( .A(rstate_text[88]), .Z(rstate_text[90]));
Q_BUF U56 ( .A(rstate_text[65]), .Z(rstate_text[88]));
Q_BUF U57 ( .A(rstate_text[64]), .Z(rstate_text[65]));
Q_BUF U58 ( .A(rstate_text[84]), .Z(rstate_text[97]));
Q_BUF U59 ( .A(rstate_text[86]), .Z(rstate_text[94]));
Q_BUF U60 ( .A(rstate_text[78]), .Z(rstate_text[86]));
Q_BUF U61 ( .A(rstate_text[70]), .Z(rstate_text[78]));
Q_BUF U62 ( .A(rstate_text[58]), .Z(rstate_text[70]));
Q_BUF U63 ( .A(rstate_text[85]), .Z(rstate_text[93]));
Q_BUF U64 ( .A(rstate_text[77]), .Z(rstate_text[85]));
Q_BUF U65 ( .A(rstate_text[69]), .Z(rstate_text[77]));
Q_BUF U66 ( .A(rstate_text[28]), .Z(rstate_text[92]));
Q_BUF U67 ( .A(rstate_text[68]), .Z(rstate_text[89]));
Q_BUF U68 ( .A(rstate_text[75]), .Z(rstate_text[83]));
Q_BUF U69 ( .A(rstate_text[74]), .Z(rstate_text[75]));
Q_BUF U70 ( .A(rstate_text[59]), .Z(rstate_text[80]));
Q_BUF U71 ( .A(rstate_text[72]), .Z(rstate_text[73]));
Q_BUF U72 ( .A(rstate_text[66]), .Z(rstate_text[67]));
Q_BUF U73 ( .A(rstate_text[46]), .Z(rstate_text[54]));
Q_BUF U74 ( .A(rstate_text[38]), .Z(rstate_text[46]));
Q_BUF U75 ( .A(rstate_text[16]), .Z(rstate_text[26]));
Q_BUF U76 ( .A(tstate_text[90]), .Z(tstate_text[94]));
Q_BUF U77 ( .A(tstate_text[88]), .Z(tstate_text[90]));
Q_BUF U78 ( .A(tstate_text[86]), .Z(tstate_text[88]));
Q_BUF U79 ( .A(tstate_text[81]), .Z(tstate_text[86]));
Q_BUF U80 ( .A(tstate_text[80]), .Z(tstate_text[81]));
Q_BUF U81 ( .A(tstate_text[78]), .Z(tstate_text[80]));
Q_BUF U82 ( .A(tstate_text[73]), .Z(tstate_text[78]));
Q_BUF U83 ( .A(tstate_text[72]), .Z(tstate_text[73]));
Q_BUF U84 ( .A(tstate_text[68]), .Z(tstate_text[72]));
Q_BUF U85 ( .A(tstate_text[49]), .Z(tstate_text[68]));
Q_BUF U86 ( .A(tstate_text[85]), .Z(tstate_text[93]));
Q_BUF U87 ( .A(tstate_text[77]), .Z(tstate_text[85]));
Q_BUF U88 ( .A(tstate_text[66]), .Z(tstate_text[67]));
Q_BUF U89 ( .A(tstate_text[64]), .Z(tstate_text[66]));
Q_BUF U90 ( .A(tstate_text[58]), .Z(tstate_text[64]));
Q_BUF U91 ( .A(tstate_text[53]), .Z(tstate_text[61]));
Q_BUF U92 ( .A(tstate_text[44]), .Z(tstate_text[56]));
Q_BUF U93 ( .A(tstate_text[29]), .Z(tstate_text[37]));
Q_BUF U94 ( .A(rstate_text[45]), .Z(rstate_text[53]));
Q_BUF U95 ( .A(rstate_text[37]), .Z(rstate_text[45]));
Q_BUF U96 ( .A(rstate_text[29]), .Z(rstate_text[37]));
Q_BUF U97 ( .A(rstate_text[21]), .Z(rstate_text[29]));
Q_BUF U98 ( .A(rstate_text[13]), .Z(rstate_text[21]));
Q_BUF U99 ( .A(rstate_text[5]), .Z(rstate_text[13]));
Q_BUF U100 ( .A(rstate_text[8]), .Z(rstate_text[25]));
Q_BUF U101 ( .A(rstate_text[1]), .Z(rstate_text[12]));
Q_BUF U102 ( .A(tstate_text[1]), .Z(tstate_text[43]));
Q_BUF U103 ( .A(tstate_text[13]), .Z(tstate_text[21]));
Q_BUF U104 ( .A(tstate_text[5]), .Z(tstate_text[13]));
Q_AN02 U105 ( .A0(n987), .A1(rx_resp), .Z(n3));
Q_AN02 U106 ( .A0(rx_resp), .A1(rx_frm), .Z(n4));
Q_INV U107 ( .A(n1232), .Z(n5));
Q_INV U108 ( .A(n1222), .Z(n6));
Q_INV U109 ( .A(n1288), .Z(n7));
Q_INV U110 ( .A(n763), .Z(n8));
Q_INV U111 ( .A(n1225), .Z(n9));
Q_INV U112 ( .A(n1227), .Z(n10));
Q_OR03 U113 ( .A0(tstate[3]), .A1(n1221), .A2(n6), .Z(n22));
Q_ND02 U114 ( .A0(n182), .A1(n22), .Z(n13));
Q_OR02 U115 ( .A0(tstate[1]), .A1(n141), .Z(n26));
Q_OR02 U116 ( .A0(tstate[3]), .A1(n26), .Z(n24));
Q_NR03 U117 ( .A0(n1212), .A1(tstate[2]), .A2(n24), .Z(n23));
Q_OR02 U118 ( .A0(n19), .A1(n23), .Z(n14));
Q_NR02 U119 ( .A0(n6), .A1(n24), .Z(n25));
Q_OR02 U120 ( .A0(n18), .A1(n25), .Z(n15));
Q_NR03 U121 ( .A0(n5), .A1(n26), .A2(tstate[0]), .Z(n27));
Q_OR02 U122 ( .A0(n17), .A1(n27), .Z(n16));
Q_INV U123 ( .A(n12), .Z(n21));
Q_FDP1 \poll_ecc_par_timer_REG[0] ( .CK(clk), .R(rst_n), .D(n54), .Q(poll_ecc_par_timer[0]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[1] ( .CK(clk), .R(rst_n), .D(n53), .Q(poll_ecc_par_timer[1]), .QN(n195));
Q_FDP1 \poll_ecc_par_timer_REG[2] ( .CK(clk), .R(rst_n), .D(n52), .Q(poll_ecc_par_timer[2]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[3] ( .CK(clk), .R(rst_n), .D(n51), .Q(poll_ecc_par_timer[3]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[4] ( .CK(clk), .R(rst_n), .D(n50), .Q(poll_ecc_par_timer[4]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[5] ( .CK(clk), .R(rst_n), .D(n49), .Q(poll_ecc_par_timer[5]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[6] ( .CK(clk), .R(rst_n), .D(n48), .Q(poll_ecc_par_timer[6]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[7] ( .CK(clk), .R(rst_n), .D(n47), .Q(poll_ecc_par_timer[7]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[8] ( .CK(clk), .R(rst_n), .D(n46), .Q(poll_ecc_par_timer[8]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[9] ( .CK(clk), .R(rst_n), .D(n45), .Q(poll_ecc_par_timer[9]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[10] ( .CK(clk), .R(rst_n), .D(n44), .Q(poll_ecc_par_timer[10]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[11] ( .CK(clk), .R(rst_n), .D(n43), .Q(poll_ecc_par_timer[11]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[12] ( .CK(clk), .R(rst_n), .D(n42), .Q(poll_ecc_par_timer[12]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[13] ( .CK(clk), .R(rst_n), .D(n41), .Q(poll_ecc_par_timer[13]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[14] ( .CK(clk), .R(rst_n), .D(n40), .Q(poll_ecc_par_timer[14]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[15] ( .CK(clk), .R(rst_n), .D(n39), .Q(poll_ecc_par_timer[15]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[16] ( .CK(clk), .R(rst_n), .D(n38), .Q(poll_ecc_par_timer[16]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[17] ( .CK(clk), .R(rst_n), .D(n37), .Q(poll_ecc_par_timer[17]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[18] ( .CK(clk), .R(rst_n), .D(n36), .Q(poll_ecc_par_timer[18]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[19] ( .CK(clk), .R(rst_n), .D(n35), .Q(poll_ecc_par_timer[19]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[20] ( .CK(clk), .R(rst_n), .D(n34), .Q(poll_ecc_par_timer[20]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[21] ( .CK(clk), .R(rst_n), .D(n33), .Q(poll_ecc_par_timer[21]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[22] ( .CK(clk), .R(rst_n), .D(n32), .Q(poll_ecc_par_timer[22]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[23] ( .CK(clk), .R(rst_n), .D(n31), .Q(poll_ecc_par_timer[23]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[24] ( .CK(clk), .R(rst_n), .D(n30), .Q(poll_ecc_par_timer[24]), .QN( ));
Q_FDP1 \poll_ecc_par_timer_REG[25] ( .CK(clk), .R(rst_n), .D(n29), .Q(poll_ecc_par_timer[25]), .QN( ));
Q_XOR2 U150 ( .A0(n108), .A1(cmd_cnt), .Z(n28));
Q_FDP2 cmd_cnt_REG  ( .CK(clk), .S(rst_n), .D(n28), .Q(cmd_cnt), .QN(n756));
Q_FDP2 \sync_cnt_REG[0] ( .CK(clk), .S(rst_n), .D(n111), .Q(sync_cnt[0]), .QN(n725));
Q_FDP1 \sync_cnt_REG[1] ( .CK(clk), .R(rst_n), .D(n110), .Q(sync_cnt[1]), .QN( ));
Q_FDP1 \sync_cnt_REG[2] ( .CK(clk), .R(rst_n), .D(n109), .Q(sync_cnt[2]), .QN( ));
Q_FDP1 \sync_cnt_REG[3] ( .CK(clk), .R(rst_n), .D(n107), .Q(sync_cnt[3]), .QN(n768));
Q_FDP1 \sync_cnt_REG[4] ( .CK(clk), .R(rst_n), .D(n106), .Q(sync_cnt[4]), .QN( ));
Q_FDP1 \sync_cnt_REG[5] ( .CK(clk), .R(rst_n), .D(n105), .Q(sync_cnt[5]), .QN( ));
Q_FDP1 \sync_cnt_REG[6] ( .CK(clk), .R(rst_n), .D(n104), .Q(sync_cnt[6]), .QN(n766));
Q_FDP1 bimc_cmd2_sent_din_REG  ( .CK(clk), .R(rst_n), .D(n135), .Q(bimc_cmd2_sent_din), .QN( ));
Q_FDP1 \r_bimc_cmd2_write_notify_ev_REG[0] ( .CK(clk), .R(rst_n), .D(bimc_cmd2_write_notify_ev), .Q(r_bimc_cmd2_write_notify_ev[0]), .QN( ));
Q_FDP1 \r_bimc_cmd2_write_notify_ev_REG[1] ( .CK(clk), .R(rst_n), .D(r_bimc_cmd2_write_notify_ev[0]), .Q(r_bimc_cmd2_write_notify_ev[1]), .QN( ));
Q_FDP1 \r_bimc_cmd2_write_notify_ev_REG[2] ( .CK(clk), .R(rst_n), .D(r_bimc_cmd2_write_notify_ev[1]), .Q(r_bimc_cmd2_write_notify_ev[2]), .QN( ));
Q_FDP1 bimc_eccpar_debug_sent_din_REG  ( .CK(clk), .R(rst_n), .D(n136), .Q(bimc_eccpar_debug_sent_din), .QN( ));
Q_FDP1 \r_bimc_eccpar_debug_write_notify_ev_REG[0] ( .CK(clk), .R(rst_n), .D(bimc_eccpar_debug_write_notify_ev), .Q(r_bimc_eccpar_debug_write_notify_ev[0]), .QN( ));
Q_FDP1 \r_bimc_eccpar_debug_write_notify_ev_REG[1] ( .CK(clk), .R(rst_n), .D(r_bimc_eccpar_debug_write_notify_ev[0]), .Q(r_bimc_eccpar_debug_write_notify_ev[1]), .QN( ));
Q_FDP1 \r_bimc_eccpar_debug_write_notify_ev_REG[2] ( .CK(clk), .R(rst_n), .D(r_bimc_eccpar_debug_write_notify_ev[1]), .Q(r_bimc_eccpar_debug_write_notify_ev[2]), .QN( ));
Q_FDP1 bimc_rst_n_REG  ( .CK(clk), .R(rst_n), .D(n199), .Q(bimc_rst_n), .QN(n765));
Q_FDP1 bimc_osync_REG  ( .CK(clk), .R(rst_n), .D(n138), .Q(bimc_osync), .QN( ));
Q_FDP1 bimc_odat_REG  ( .CK(clk), .R(rst_n), .D(n123), .Q(bimc_odat), .QN( ));
Q_AN02 U170 ( .A0(n21), .A1(n55), .Z(n29));
Q_AN02 U171 ( .A0(n21), .A1(n57), .Z(n30));
Q_AN02 U172 ( .A0(n21), .A1(n59), .Z(n31));
Q_AN02 U173 ( .A0(n21), .A1(n61), .Z(n32));
Q_AN02 U174 ( .A0(n21), .A1(n63), .Z(n33));
Q_AN02 U175 ( .A0(n21), .A1(n65), .Z(n34));
Q_AN02 U176 ( .A0(n21), .A1(n67), .Z(n35));
Q_AN02 U177 ( .A0(n21), .A1(n69), .Z(n36));
Q_AN02 U178 ( .A0(n21), .A1(n71), .Z(n37));
Q_AN02 U179 ( .A0(n21), .A1(n73), .Z(n38));
Q_AN02 U180 ( .A0(n21), .A1(n75), .Z(n39));
Q_AN02 U181 ( .A0(n21), .A1(n77), .Z(n40));
Q_AN02 U182 ( .A0(n21), .A1(n79), .Z(n41));
Q_AN02 U183 ( .A0(n21), .A1(n81), .Z(n42));
Q_AN02 U184 ( .A0(n21), .A1(n83), .Z(n43));
Q_AN02 U185 ( .A0(n21), .A1(n85), .Z(n44));
Q_AN02 U186 ( .A0(n21), .A1(n87), .Z(n45));
Q_AN02 U187 ( .A0(n21), .A1(n89), .Z(n46));
Q_AN02 U188 ( .A0(n21), .A1(n91), .Z(n47));
Q_AN02 U189 ( .A0(n21), .A1(n93), .Z(n48));
Q_AN02 U190 ( .A0(n21), .A1(n95), .Z(n49));
Q_AN02 U191 ( .A0(n21), .A1(n97), .Z(n50));
Q_AN02 U192 ( .A0(n21), .A1(n99), .Z(n51));
Q_AN02 U193 ( .A0(n21), .A1(n101), .Z(n52));
Q_AN02 U194 ( .A0(n21), .A1(n103), .Z(n53));
Q_NR02 U195 ( .A0(n12), .A1(poll_ecc_par_timer[0]), .Z(n54));
Q_XOR2 U196 ( .A0(poll_ecc_par_timer[25]), .A1(n56), .Z(n55));
Q_AD01HF U197 ( .A0(poll_ecc_par_timer[24]), .B0(n58), .S(n57), .CO(n56));
Q_AD01HF U198 ( .A0(poll_ecc_par_timer[23]), .B0(n60), .S(n59), .CO(n58));
Q_AD01HF U199 ( .A0(poll_ecc_par_timer[22]), .B0(n62), .S(n61), .CO(n60));
Q_AD01HF U200 ( .A0(poll_ecc_par_timer[21]), .B0(n64), .S(n63), .CO(n62));
Q_AD01HF U201 ( .A0(poll_ecc_par_timer[20]), .B0(n66), .S(n65), .CO(n64));
Q_AD01HF U202 ( .A0(poll_ecc_par_timer[19]), .B0(n68), .S(n67), .CO(n66));
Q_AD01HF U203 ( .A0(poll_ecc_par_timer[18]), .B0(n70), .S(n69), .CO(n68));
Q_AD01HF U204 ( .A0(poll_ecc_par_timer[17]), .B0(n72), .S(n71), .CO(n70));
Q_AD01HF U205 ( .A0(poll_ecc_par_timer[16]), .B0(n74), .S(n73), .CO(n72));
Q_AD01HF U206 ( .A0(poll_ecc_par_timer[15]), .B0(n76), .S(n75), .CO(n74));
Q_AD01HF U207 ( .A0(poll_ecc_par_timer[14]), .B0(n78), .S(n77), .CO(n76));
Q_AD01HF U208 ( .A0(poll_ecc_par_timer[13]), .B0(n80), .S(n79), .CO(n78));
Q_AD01HF U209 ( .A0(poll_ecc_par_timer[12]), .B0(n82), .S(n81), .CO(n80));
Q_AD01HF U210 ( .A0(poll_ecc_par_timer[11]), .B0(n84), .S(n83), .CO(n82));
Q_AD01HF U211 ( .A0(poll_ecc_par_timer[10]), .B0(n86), .S(n85), .CO(n84));
Q_AD01HF U212 ( .A0(poll_ecc_par_timer[9]), .B0(n88), .S(n87), .CO(n86));
Q_AD01HF U213 ( .A0(poll_ecc_par_timer[8]), .B0(n90), .S(n89), .CO(n88));
Q_AD01HF U214 ( .A0(poll_ecc_par_timer[7]), .B0(n92), .S(n91), .CO(n90));
Q_AD01HF U215 ( .A0(poll_ecc_par_timer[6]), .B0(n94), .S(n93), .CO(n92));
Q_AD01HF U216 ( .A0(poll_ecc_par_timer[5]), .B0(n96), .S(n95), .CO(n94));
Q_AD01HF U217 ( .A0(poll_ecc_par_timer[4]), .B0(n98), .S(n97), .CO(n96));
Q_AD01HF U218 ( .A0(poll_ecc_par_timer[3]), .B0(n100), .S(n99), .CO(n98));
Q_AD01HF U219 ( .A0(poll_ecc_par_timer[2]), .B0(n102), .S(n101), .CO(n100));
Q_AD01HF U220 ( .A0(poll_ecc_par_timer[1]), .B0(poll_ecc_par_timer[0]), .S(n103), .CO(n102));
Q_OR02 U221 ( .A0(n108), .A1(n112), .Z(n104));
Q_AN02 U222 ( .A0(n196), .A1(n114), .Z(n105));
Q_AN02 U223 ( .A0(n196), .A1(n116), .Z(n106));
Q_OR02 U224 ( .A0(n108), .A1(n118), .Z(n107));
Q_INV U225 ( .A(n196), .Z(n108));
Q_AN02 U226 ( .A0(n196), .A1(n120), .Z(n109));
Q_AN02 U227 ( .A0(n196), .A1(n122), .Z(n110));
Q_AN02 U228 ( .A0(n196), .A1(n725), .Z(n111));
Q_XNR2 U229 ( .A0(sync_cnt[6]), .A1(n113), .Z(n112));
Q_OR02 U230 ( .A0(sync_cnt[5]), .A1(n115), .Z(n113));
Q_XNR2 U231 ( .A0(sync_cnt[5]), .A1(n115), .Z(n114));
Q_OR02 U232 ( .A0(sync_cnt[4]), .A1(n117), .Z(n115));
Q_XNR2 U233 ( .A0(sync_cnt[4]), .A1(n117), .Z(n116));
Q_OR02 U234 ( .A0(sync_cnt[3]), .A1(n119), .Z(n117));
Q_XNR2 U235 ( .A0(sync_cnt[3]), .A1(n119), .Z(n118));
Q_OR02 U236 ( .A0(sync_cnt[2]), .A1(n121), .Z(n119));
Q_XNR2 U237 ( .A0(sync_cnt[2]), .A1(n121), .Z(n120));
Q_OR02 U238 ( .A0(sync_cnt[1]), .A1(sync_cnt[0]), .Z(n121));
Q_XNR2 U239 ( .A0(sync_cnt[1]), .A1(sync_cnt[0]), .Z(n122));
Q_MX02 U240 ( .S(sync_cnt[6]), .A0(n124), .A1(n133), .Z(n123));
Q_MX08 U241 ( .S0(sync_cnt[3]), .S1(sync_cnt[4]), .S2(sync_cnt[5]), .A0(n125), .A1(n126), .A2(n127), .A3(n128), .A4(n129), .A5(n130), .A6(n131), .A7(n132), .Z(n124));
Q_MX08 U242 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[0]), .A1(reg_send[1]), .A2(reg_send[2]), .A3(reg_send[3]), .A4(reg_send[4]), .A5(reg_send[5]), .A6(reg_send[6]), .A7(reg_send[7]), .Z(n125));
Q_MX08 U243 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[8]), .A1(reg_send[9]), .A2(reg_send[10]), .A3(reg_send[11]), .A4(reg_send[12]), .A5(reg_send[13]), .A6(reg_send[14]), .A7(reg_send[15]), .Z(n126));
Q_MX08 U244 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[16]), .A1(reg_send[17]), .A2(reg_send[18]), .A3(reg_send[19]), .A4(reg_send[20]), .A5(reg_send[21]), .A6(reg_send[22]), .A7(reg_send[23]), .Z(n127));
Q_MX08 U245 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[24]), .A1(reg_send[25]), .A2(reg_send[26]), .A3(reg_send[27]), .A4(reg_send[28]), .A5(reg_send[29]), .A6(reg_send[30]), .A7(reg_send[31]), .Z(n128));
Q_MX08 U246 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[32]), .A1(reg_send[33]), .A2(reg_send[34]), .A3(reg_send[35]), .A4(reg_send[36]), .A5(reg_send[37]), .A6(reg_send[38]), .A7(reg_send[39]), .Z(n129));
Q_MX08 U247 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[40]), .A1(reg_send[41]), .A2(reg_send[42]), .A3(reg_send[43]), .A4(reg_send[44]), .A5(reg_send[45]), .A6(reg_send[46]), .A7(reg_send[47]), .Z(n130));
Q_MX08 U248 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[48]), .A1(reg_send[49]), .A2(reg_send[50]), .A3(reg_send[51]), .A4(reg_send[52]), .A5(reg_send[53]), .A6(reg_send[54]), .A7(reg_send[55]), .Z(n131));
Q_MX08 U249 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[56]), .A1(reg_send[57]), .A2(reg_send[58]), .A3(reg_send[59]), .A4(reg_send[60]), .A5(reg_send[61]), .A6(reg_send[62]), .A7(reg_send[63]), .Z(n132));
Q_MX02 U250 ( .S(sync_cnt[3]), .A0(n134), .A1(reg_send[72]), .Z(n133));
Q_MX08 U251 ( .S0(sync_cnt[0]), .S1(sync_cnt[1]), .S2(sync_cnt[2]), .A0(reg_send[64]), .A1(reg_send[65]), .A2(reg_send[66]), .A3(reg_send[67]), .A4(reg_send[68]), .A5(reg_send[69]), .A6(reg_send[70]), .A7(reg_send[71]), .Z(n134));
Q_NR03 U252 ( .A0(n1212), .A1(n1165), .A2(n141), .Z(n135));
Q_AN03 U253 ( .A0(tstate[0]), .A1(n137), .A2(n11), .Z(n136));
Q_AN03 U254 ( .A0(n1196), .A1(tstate[2]), .A2(n1221), .Z(n137));
Q_NR03 U255 ( .A0(sync_cnt[0]), .A1(n140), .A2(n139), .Z(n138));
Q_OR03 U256 ( .A0(n768), .A1(sync_cnt[2]), .A2(sync_cnt[1]), .Z(n139));
Q_OR03 U257 ( .A0(n766), .A1(sync_cnt[5]), .A2(sync_cnt[4]), .Z(n140));
Q_AN02 U258 ( .A0(r_bimc_cmd2_write_notify_ev[2]), .A1(bimc_cmd2_send), .Z(n19));
Q_AN02 U259 ( .A0(r_bimc_eccpar_debug_write_notify_ev[2]), .A1(bimc_eccpar_debug_send), .Z(n18));
Q_INV U260 ( .A(n141), .Z(n11));
Q_OR03 U261 ( .A0(n725), .A1(n198), .A2(n197), .Z(n141));
Q_AN02 U262 ( .A0(n142), .A1(bimc_global_config_mem_wr_init), .Z(n17));
Q_INV U263 ( .A(bimc_global_config_poll_ecc_par_error), .Z(n143));
Q_AO21 U264 ( .A0(n145), .A1(n144), .B0(n143), .Z(n12));
Q_AN03 U265 ( .A0(n148), .A1(n147), .A2(n146), .Z(n144));
Q_AN03 U266 ( .A0(n151), .A1(n150), .A2(n149), .Z(n145));
Q_AN03 U267 ( .A0(n154), .A1(n153), .A2(n152), .Z(n146));
Q_AN03 U268 ( .A0(n180), .A1(n181), .A2(n155), .Z(n147));
Q_AN03 U269 ( .A0(n177), .A1(n178), .A2(n179), .Z(n148));
Q_AN03 U270 ( .A0(n174), .A1(n175), .A2(n176), .Z(n149));
Q_AN03 U271 ( .A0(n171), .A1(n172), .A2(n173), .Z(n150));
Q_AN03 U272 ( .A0(n168), .A1(n169), .A2(n170), .Z(n151));
Q_AN03 U273 ( .A0(n165), .A1(n166), .A2(n167), .Z(n152));
Q_AN03 U274 ( .A0(n162), .A1(n163), .A2(n164), .Z(n153));
Q_AN03 U275 ( .A0(n159), .A1(n160), .A2(n161), .Z(n154));
Q_AN03 U276 ( .A0(n156), .A1(n157), .A2(n158), .Z(n155));
Q_XNR2 U277 ( .A0(poll_ecc_par_timer[25]), .A1(bimc_global_config_poll_ecc_par_timer[25]), .Z(n156));
Q_XNR2 U278 ( .A0(poll_ecc_par_timer[24]), .A1(bimc_global_config_poll_ecc_par_timer[24]), .Z(n157));
Q_XNR2 U279 ( .A0(poll_ecc_par_timer[23]), .A1(bimc_global_config_poll_ecc_par_timer[23]), .Z(n158));
Q_XNR2 U280 ( .A0(poll_ecc_par_timer[22]), .A1(bimc_global_config_poll_ecc_par_timer[22]), .Z(n159));
Q_XNR2 U281 ( .A0(poll_ecc_par_timer[21]), .A1(bimc_global_config_poll_ecc_par_timer[21]), .Z(n160));
Q_XNR2 U282 ( .A0(poll_ecc_par_timer[20]), .A1(bimc_global_config_poll_ecc_par_timer[20]), .Z(n161));
Q_XNR2 U283 ( .A0(poll_ecc_par_timer[19]), .A1(bimc_global_config_poll_ecc_par_timer[19]), .Z(n162));
Q_XNR2 U284 ( .A0(poll_ecc_par_timer[18]), .A1(bimc_global_config_poll_ecc_par_timer[18]), .Z(n163));
Q_XNR2 U285 ( .A0(poll_ecc_par_timer[17]), .A1(bimc_global_config_poll_ecc_par_timer[17]), .Z(n164));
Q_XNR2 U286 ( .A0(poll_ecc_par_timer[16]), .A1(bimc_global_config_poll_ecc_par_timer[16]), .Z(n165));
Q_XNR2 U287 ( .A0(poll_ecc_par_timer[15]), .A1(bimc_global_config_poll_ecc_par_timer[15]), .Z(n166));
Q_XNR2 U288 ( .A0(poll_ecc_par_timer[14]), .A1(bimc_global_config_poll_ecc_par_timer[14]), .Z(n167));
Q_XNR2 U289 ( .A0(poll_ecc_par_timer[13]), .A1(bimc_global_config_poll_ecc_par_timer[13]), .Z(n168));
Q_XNR2 U290 ( .A0(poll_ecc_par_timer[12]), .A1(bimc_global_config_poll_ecc_par_timer[12]), .Z(n169));
Q_XNR2 U291 ( .A0(poll_ecc_par_timer[11]), .A1(bimc_global_config_poll_ecc_par_timer[11]), .Z(n170));
Q_XNR2 U292 ( .A0(poll_ecc_par_timer[10]), .A1(bimc_global_config_poll_ecc_par_timer[10]), .Z(n171));
Q_XNR2 U293 ( .A0(poll_ecc_par_timer[9]), .A1(bimc_global_config_poll_ecc_par_timer[9]), .Z(n172));
Q_XNR2 U294 ( .A0(poll_ecc_par_timer[8]), .A1(bimc_global_config_poll_ecc_par_timer[8]), .Z(n173));
Q_XNR2 U295 ( .A0(poll_ecc_par_timer[7]), .A1(bimc_global_config_poll_ecc_par_timer[7]), .Z(n174));
Q_XNR2 U296 ( .A0(poll_ecc_par_timer[6]), .A1(bimc_global_config_poll_ecc_par_timer[6]), .Z(n175));
Q_XNR2 U297 ( .A0(poll_ecc_par_timer[5]), .A1(bimc_global_config_poll_ecc_par_timer[5]), .Z(n176));
Q_XNR2 U298 ( .A0(poll_ecc_par_timer[4]), .A1(bimc_global_config_poll_ecc_par_timer[4]), .Z(n177));
Q_XNR2 U299 ( .A0(poll_ecc_par_timer[3]), .A1(bimc_global_config_poll_ecc_par_timer[3]), .Z(n178));
Q_XNR2 U300 ( .A0(poll_ecc_par_timer[2]), .A1(bimc_global_config_poll_ecc_par_timer[2]), .Z(n179));
Q_XNR2 U301 ( .A0(poll_ecc_par_timer[1]), .A1(bimc_global_config_poll_ecc_par_timer[1]), .Z(n180));
Q_XNR2 U302 ( .A0(poll_ecc_par_timer[0]), .A1(bimc_global_config_poll_ecc_par_timer[0]), .Z(n181));
Q_INV U303 ( .A(n182), .Z(n20));
Q_OR02 U304 ( .A0(n184), .A1(n183), .Z(n182));
Q_OR03 U305 ( .A0(n187), .A1(n186), .A2(n185), .Z(n183));
Q_OR03 U306 ( .A0(n190), .A1(n189), .A2(n188), .Z(n184));
Q_OR03 U307 ( .A0(n193), .A1(n192), .A2(n191), .Z(n185));
Q_OR03 U308 ( .A0(n195), .A1(poll_ecc_par_timer[0]), .A2(n194), .Z(n186));
Q_OR03 U309 ( .A0(poll_ecc_par_timer[4]), .A1(poll_ecc_par_timer[3]), .A2(poll_ecc_par_timer[2]), .Z(n187));
Q_OR03 U310 ( .A0(poll_ecc_par_timer[7]), .A1(poll_ecc_par_timer[6]), .A2(poll_ecc_par_timer[5]), .Z(n188));
Q_OR03 U311 ( .A0(poll_ecc_par_timer[10]), .A1(poll_ecc_par_timer[9]), .A2(poll_ecc_par_timer[8]), .Z(n189));
Q_OR03 U312 ( .A0(poll_ecc_par_timer[13]), .A1(poll_ecc_par_timer[12]), .A2(poll_ecc_par_timer[11]), .Z(n190));
Q_OR03 U313 ( .A0(poll_ecc_par_timer[16]), .A1(poll_ecc_par_timer[15]), .A2(poll_ecc_par_timer[14]), .Z(n191));
Q_OR03 U314 ( .A0(poll_ecc_par_timer[19]), .A1(poll_ecc_par_timer[18]), .A2(poll_ecc_par_timer[17]), .Z(n192));
Q_OR03 U315 ( .A0(poll_ecc_par_timer[22]), .A1(poll_ecc_par_timer[21]), .A2(poll_ecc_par_timer[20]), .Z(n193));
Q_OR03 U316 ( .A0(poll_ecc_par_timer[25]), .A1(poll_ecc_par_timer[24]), .A2(poll_ecc_par_timer[23]), .Z(n194));
Q_OR03 U317 ( .A0(sync_cnt[0]), .A1(n198), .A2(n197), .Z(n196));
Q_OR03 U318 ( .A0(sync_cnt[3]), .A1(sync_cnt[2]), .A2(sync_cnt[1]), .Z(n197));
Q_OR03 U319 ( .A0(sync_cnt[6]), .A1(sync_cnt[5]), .A2(sync_cnt[4]), .Z(n198));
Q_INV U320 ( .A(bimc_global_config_soft_reset), .Z(n199));
Q_FDP1 \r_reg_send_REG[0] ( .CK(clk), .R(rst_n), .D(reg_send[0]), .Q(r_reg_send[0]), .QN( ));
Q_FDP1 \r_reg_send_REG[1] ( .CK(clk), .R(rst_n), .D(reg_send[1]), .Q(r_reg_send[1]), .QN( ));
Q_FDP1 \r_reg_send_REG[2] ( .CK(clk), .R(rst_n), .D(reg_send[2]), .Q(r_reg_send[2]), .QN( ));
Q_FDP1 \r_reg_send_REG[3] ( .CK(clk), .R(rst_n), .D(reg_send[3]), .Q(r_reg_send[3]), .QN( ));
Q_FDP1 \r_reg_send_REG[4] ( .CK(clk), .R(rst_n), .D(reg_send[4]), .Q(r_reg_send[4]), .QN( ));
Q_FDP1 \r_reg_send_REG[5] ( .CK(clk), .R(rst_n), .D(reg_send[5]), .Q(r_reg_send[5]), .QN( ));
Q_FDP1 \r_reg_send_REG[6] ( .CK(clk), .R(rst_n), .D(reg_send[6]), .Q(r_reg_send[6]), .QN( ));
Q_FDP1 \r_reg_send_REG[7] ( .CK(clk), .R(rst_n), .D(reg_send[7]), .Q(r_reg_send[7]), .QN( ));
Q_FDP1 \r_reg_send_REG[8] ( .CK(clk), .R(rst_n), .D(reg_send[8]), .Q(r_reg_send[8]), .QN( ));
Q_FDP1 \r_reg_send_REG[9] ( .CK(clk), .R(rst_n), .D(reg_send[9]), .Q(r_reg_send[9]), .QN( ));
Q_FDP1 \r_reg_send_REG[10] ( .CK(clk), .R(rst_n), .D(reg_send[10]), .Q(r_reg_send[10]), .QN( ));
Q_FDP1 \r_reg_send_REG[11] ( .CK(clk), .R(rst_n), .D(reg_send[11]), .Q(r_reg_send[11]), .QN( ));
Q_FDP1 \r_reg_send_REG[12] ( .CK(clk), .R(rst_n), .D(reg_send[12]), .Q(r_reg_send[12]), .QN( ));
Q_FDP1 \r_reg_send_REG[13] ( .CK(clk), .R(rst_n), .D(reg_send[13]), .Q(r_reg_send[13]), .QN( ));
Q_FDP1 \r_reg_send_REG[14] ( .CK(clk), .R(rst_n), .D(reg_send[14]), .Q(r_reg_send[14]), .QN( ));
Q_FDP1 \r_reg_send_REG[15] ( .CK(clk), .R(rst_n), .D(reg_send[15]), .Q(r_reg_send[15]), .QN( ));
Q_FDP1 \r_reg_send_REG[16] ( .CK(clk), .R(rst_n), .D(reg_send[16]), .Q(r_reg_send[16]), .QN( ));
Q_FDP1 \r_reg_send_REG[17] ( .CK(clk), .R(rst_n), .D(reg_send[17]), .Q(r_reg_send[17]), .QN( ));
Q_FDP1 \r_reg_send_REG[18] ( .CK(clk), .R(rst_n), .D(reg_send[18]), .Q(r_reg_send[18]), .QN( ));
Q_FDP1 \r_reg_send_REG[19] ( .CK(clk), .R(rst_n), .D(reg_send[19]), .Q(r_reg_send[19]), .QN( ));
Q_FDP1 \r_reg_send_REG[20] ( .CK(clk), .R(rst_n), .D(reg_send[20]), .Q(r_reg_send[20]), .QN( ));
Q_FDP1 \r_reg_send_REG[21] ( .CK(clk), .R(rst_n), .D(reg_send[21]), .Q(r_reg_send[21]), .QN( ));
Q_FDP1 \r_reg_send_REG[22] ( .CK(clk), .R(rst_n), .D(reg_send[22]), .Q(r_reg_send[22]), .QN( ));
Q_FDP1 \r_reg_send_REG[23] ( .CK(clk), .R(rst_n), .D(reg_send[23]), .Q(r_reg_send[23]), .QN( ));
Q_FDP1 \r_reg_send_REG[24] ( .CK(clk), .R(rst_n), .D(reg_send[24]), .Q(r_reg_send[24]), .QN( ));
Q_FDP1 \r_reg_send_REG[25] ( .CK(clk), .R(rst_n), .D(reg_send[25]), .Q(r_reg_send[25]), .QN( ));
Q_FDP1 \r_reg_send_REG[26] ( .CK(clk), .R(rst_n), .D(reg_send[26]), .Q(r_reg_send[26]), .QN( ));
Q_FDP1 \r_reg_send_REG[27] ( .CK(clk), .R(rst_n), .D(reg_send[27]), .Q(r_reg_send[27]), .QN( ));
Q_FDP1 \r_reg_send_REG[28] ( .CK(clk), .R(rst_n), .D(reg_send[28]), .Q(r_reg_send[28]), .QN( ));
Q_FDP1 \r_reg_send_REG[29] ( .CK(clk), .R(rst_n), .D(reg_send[29]), .Q(r_reg_send[29]), .QN( ));
Q_FDP1 \r_reg_send_REG[30] ( .CK(clk), .R(rst_n), .D(reg_send[30]), .Q(r_reg_send[30]), .QN( ));
Q_FDP1 \r_reg_send_REG[31] ( .CK(clk), .R(rst_n), .D(reg_send[31]), .Q(r_reg_send[31]), .QN( ));
Q_FDP1 \r_reg_send_REG[32] ( .CK(clk), .R(rst_n), .D(reg_send[32]), .Q(r_reg_send[32]), .QN( ));
Q_FDP1 \r_reg_send_REG[33] ( .CK(clk), .R(rst_n), .D(reg_send[33]), .Q(r_reg_send[33]), .QN( ));
Q_FDP1 \r_reg_send_REG[34] ( .CK(clk), .R(rst_n), .D(reg_send[34]), .Q(r_reg_send[34]), .QN( ));
Q_FDP1 \r_reg_send_REG[35] ( .CK(clk), .R(rst_n), .D(reg_send[35]), .Q(r_reg_send[35]), .QN( ));
Q_FDP1 \r_reg_send_REG[36] ( .CK(clk), .R(rst_n), .D(reg_send[36]), .Q(r_reg_send[36]), .QN( ));
Q_FDP1 \r_reg_send_REG[37] ( .CK(clk), .R(rst_n), .D(reg_send[37]), .Q(r_reg_send[37]), .QN( ));
Q_FDP1 \r_reg_send_REG[38] ( .CK(clk), .R(rst_n), .D(reg_send[38]), .Q(r_reg_send[38]), .QN( ));
Q_FDP1 \r_reg_send_REG[39] ( .CK(clk), .R(rst_n), .D(reg_send[39]), .Q(r_reg_send[39]), .QN( ));
Q_FDP1 \r_reg_send_REG[40] ( .CK(clk), .R(rst_n), .D(reg_send[40]), .Q(r_reg_send[40]), .QN( ));
Q_FDP1 \r_reg_send_REG[41] ( .CK(clk), .R(rst_n), .D(reg_send[41]), .Q(r_reg_send[41]), .QN( ));
Q_FDP1 \r_reg_send_REG[42] ( .CK(clk), .R(rst_n), .D(reg_send[42]), .Q(r_reg_send[42]), .QN( ));
Q_FDP1 \r_reg_send_REG[43] ( .CK(clk), .R(rst_n), .D(reg_send[43]), .Q(r_reg_send[43]), .QN( ));
Q_FDP1 \r_reg_send_REG[44] ( .CK(clk), .R(rst_n), .D(reg_send[44]), .Q(r_reg_send[44]), .QN( ));
Q_FDP1 \r_reg_send_REG[45] ( .CK(clk), .R(rst_n), .D(reg_send[45]), .Q(r_reg_send[45]), .QN( ));
Q_FDP1 \r_reg_send_REG[46] ( .CK(clk), .R(rst_n), .D(reg_send[46]), .Q(r_reg_send[46]), .QN( ));
Q_FDP1 \r_reg_send_REG[47] ( .CK(clk), .R(rst_n), .D(reg_send[47]), .Q(r_reg_send[47]), .QN( ));
Q_FDP1 \r_reg_send_REG[48] ( .CK(clk), .R(rst_n), .D(reg_send[48]), .Q(r_reg_send[48]), .QN( ));
Q_FDP1 \r_reg_send_REG[49] ( .CK(clk), .R(rst_n), .D(reg_send[49]), .Q(r_reg_send[49]), .QN( ));
Q_FDP1 \r_reg_send_REG[50] ( .CK(clk), .R(rst_n), .D(reg_send[50]), .Q(r_reg_send[50]), .QN( ));
Q_FDP1 \r_reg_send_REG[51] ( .CK(clk), .R(rst_n), .D(reg_send[51]), .Q(r_reg_send[51]), .QN( ));
Q_FDP1 \r_reg_send_REG[52] ( .CK(clk), .R(rst_n), .D(reg_send[52]), .Q(r_reg_send[52]), .QN( ));
Q_FDP1 \r_reg_send_REG[53] ( .CK(clk), .R(rst_n), .D(reg_send[53]), .Q(r_reg_send[53]), .QN( ));
Q_FDP1 \r_reg_send_REG[54] ( .CK(clk), .R(rst_n), .D(reg_send[54]), .Q(r_reg_send[54]), .QN( ));
Q_FDP1 \r_reg_send_REG[55] ( .CK(clk), .R(rst_n), .D(reg_send[55]), .Q(r_reg_send[55]), .QN( ));
Q_FDP1 \r_reg_send_REG[56] ( .CK(clk), .R(rst_n), .D(reg_send[56]), .Q(r_reg_send[56]), .QN( ));
Q_FDP1 \r_reg_send_REG[57] ( .CK(clk), .R(rst_n), .D(reg_send[57]), .Q(r_reg_send[57]), .QN( ));
Q_FDP1 \r_reg_send_REG[58] ( .CK(clk), .R(rst_n), .D(reg_send[58]), .Q(r_reg_send[58]), .QN( ));
Q_FDP1 \r_reg_send_REG[59] ( .CK(clk), .R(rst_n), .D(reg_send[59]), .Q(r_reg_send[59]), .QN( ));
Q_FDP1 \r_reg_send_REG[60] ( .CK(clk), .R(rst_n), .D(reg_send[60]), .Q(r_reg_send[60]), .QN( ));
Q_FDP1 \r_reg_send_REG[61] ( .CK(clk), .R(rst_n), .D(reg_send[61]), .Q(r_reg_send[61]), .QN( ));
Q_FDP1 \r_reg_send_REG[62] ( .CK(clk), .R(rst_n), .D(reg_send[62]), .Q(r_reg_send[62]), .QN( ));
Q_FDP1 \r_reg_send_REG[63] ( .CK(clk), .R(rst_n), .D(reg_send[63]), .Q(r_reg_send[63]), .QN( ));
Q_FDP1 \r_reg_send_REG[64] ( .CK(clk), .R(rst_n), .D(reg_send[64]), .Q(r_reg_send[64]), .QN( ));
Q_FDP1 \r_reg_send_REG[65] ( .CK(clk), .R(rst_n), .D(reg_send[65]), .Q(r_reg_send[65]), .QN( ));
Q_FDP1 \r_reg_send_REG[66] ( .CK(clk), .R(rst_n), .D(reg_send[66]), .Q(r_reg_send[66]), .QN( ));
Q_FDP1 \r_reg_send_REG[67] ( .CK(clk), .R(rst_n), .D(reg_send[67]), .Q(r_reg_send[67]), .QN( ));
Q_FDP1 \r_reg_send_REG[68] ( .CK(clk), .R(rst_n), .D(reg_send[68]), .Q(r_reg_send[68]), .QN( ));
Q_FDP1 \r_reg_send_REG[69] ( .CK(clk), .R(rst_n), .D(reg_send[69]), .Q(r_reg_send[69]), .QN( ));
Q_FDP1 \r_reg_send_REG[70] ( .CK(clk), .R(rst_n), .D(reg_send[70]), .Q(r_reg_send[70]), .QN( ));
Q_FDP1 \r_reg_send_REG[71] ( .CK(clk), .R(rst_n), .D(reg_send[71]), .Q(r_reg_send[71]), .QN( ));
Q_FDP1 \r_reg_send_REG[72] ( .CK(clk), .R(rst_n), .D(reg_send[72]), .Q(r_reg_send[72]), .QN( ));
Q_FDP1 mem_wr_init_dly_REG  ( .CK(clk), .R(rst_n), .D(bimc_global_config_mem_wr_init), .Q(mem_wr_init_dly), .QN(n142));
Q_FDP1 \tstate_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_tstate[0]), .Q(tstate[0]), .QN(n1212));
Q_FDP1 \tstate_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_tstate[1]), .Q(tstate[1]), .QN(n1221));
Q_FDP1 \tstate_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_tstate[2]), .Q(tstate[2]), .QN(n1201));
Q_FDP1 \tstate_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_tstate[3]), .Q(tstate[3]), .QN(n1196));
Q_FDP1 bimc_cmd2_send_REG  ( .CK(clk), .R(rst_n), .D(o_bimc_cmd2[8]), .Q(bimc_cmd2_send), .QN(n1317));
Q_FDP1 bimc_eccpar_debug_send_REG  ( .CK(clk), .R(rst_n), .D(o_bimc_eccpar_debug[22]), .Q(bimc_eccpar_debug_send), .QN(n1316));
Q_FDP1 bimc_interrupt_REG  ( .CK(clk), .R(rst_n), .D(bimc_interrupt_c), .Q(bimc_interrupt), .QN( ));
Q_FDP1 bimc_ecc_error_REG  ( .CK(clk), .R(rst_n), .D(bimc_ecc_error_c), .Q(bimc_ecc_error), .QN( ));
Q_INV U403 ( .A(o_bimc_eccpar_debug[28]), .Z(n205));
Q_NR02 U404 ( .A0(o_bimc_eccpar_debug[28]), .A1(bimc_eccpar_debug_sent_din), .Z(n202));
Q_AN02 U405 ( .A0(n205), .A1(bimc_eccpar_debug_sent_din), .Z(n203));
Q_INV U406 ( .A(o_bimc_cmd2[10]), .Z(n204));
Q_FDP1 \bimc_parity_error_cnt_REG[0] ( .CK(clk), .R(rst_n), .D(n270), .Q(bimc_parity_error_cnt[0]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[1] ( .CK(clk), .R(rst_n), .D(n269), .Q(bimc_parity_error_cnt[1]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[2] ( .CK(clk), .R(rst_n), .D(n268), .Q(bimc_parity_error_cnt[2]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[3] ( .CK(clk), .R(rst_n), .D(n267), .Q(bimc_parity_error_cnt[3]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[4] ( .CK(clk), .R(rst_n), .D(n266), .Q(bimc_parity_error_cnt[4]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[5] ( .CK(clk), .R(rst_n), .D(n265), .Q(bimc_parity_error_cnt[5]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[6] ( .CK(clk), .R(rst_n), .D(n264), .Q(bimc_parity_error_cnt[6]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[7] ( .CK(clk), .R(rst_n), .D(n263), .Q(bimc_parity_error_cnt[7]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[8] ( .CK(clk), .R(rst_n), .D(n262), .Q(bimc_parity_error_cnt[8]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[9] ( .CK(clk), .R(rst_n), .D(n261), .Q(bimc_parity_error_cnt[9]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[10] ( .CK(clk), .R(rst_n), .D(n260), .Q(bimc_parity_error_cnt[10]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[11] ( .CK(clk), .R(rst_n), .D(n259), .Q(bimc_parity_error_cnt[11]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[12] ( .CK(clk), .R(rst_n), .D(n258), .Q(bimc_parity_error_cnt[12]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[13] ( .CK(clk), .R(rst_n), .D(n257), .Q(bimc_parity_error_cnt[13]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[14] ( .CK(clk), .R(rst_n), .D(n256), .Q(bimc_parity_error_cnt[14]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[15] ( .CK(clk), .R(rst_n), .D(n255), .Q(bimc_parity_error_cnt[15]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[16] ( .CK(clk), .R(rst_n), .D(n254), .Q(bimc_parity_error_cnt[16]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[17] ( .CK(clk), .R(rst_n), .D(n253), .Q(bimc_parity_error_cnt[17]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[18] ( .CK(clk), .R(rst_n), .D(n252), .Q(bimc_parity_error_cnt[18]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[19] ( .CK(clk), .R(rst_n), .D(n251), .Q(bimc_parity_error_cnt[19]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[20] ( .CK(clk), .R(rst_n), .D(n250), .Q(bimc_parity_error_cnt[20]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[21] ( .CK(clk), .R(rst_n), .D(n249), .Q(bimc_parity_error_cnt[21]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[22] ( .CK(clk), .R(rst_n), .D(n248), .Q(bimc_parity_error_cnt[22]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[23] ( .CK(clk), .R(rst_n), .D(n247), .Q(bimc_parity_error_cnt[23]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[24] ( .CK(clk), .R(rst_n), .D(n246), .Q(bimc_parity_error_cnt[24]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[25] ( .CK(clk), .R(rst_n), .D(n245), .Q(bimc_parity_error_cnt[25]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[26] ( .CK(clk), .R(rst_n), .D(n244), .Q(bimc_parity_error_cnt[26]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[27] ( .CK(clk), .R(rst_n), .D(n243), .Q(bimc_parity_error_cnt[27]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[28] ( .CK(clk), .R(rst_n), .D(n242), .Q(bimc_parity_error_cnt[28]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[29] ( .CK(clk), .R(rst_n), .D(n241), .Q(bimc_parity_error_cnt[29]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[30] ( .CK(clk), .R(rst_n), .D(n240), .Q(bimc_parity_error_cnt[30]), .QN( ));
Q_FDP1 \bimc_parity_error_cnt_REG[31] ( .CK(clk), .R(rst_n), .D(n239), .Q(bimc_parity_error_cnt[31]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[0] ( .CK(clk), .R(rst_n), .D(n429), .Q(bimc_ecc_correctable_error_cnt[0]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[1] ( .CK(clk), .R(rst_n), .D(n428), .Q(bimc_ecc_correctable_error_cnt[1]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[2] ( .CK(clk), .R(rst_n), .D(n427), .Q(bimc_ecc_correctable_error_cnt[2]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[3] ( .CK(clk), .R(rst_n), .D(n426), .Q(bimc_ecc_correctable_error_cnt[3]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[4] ( .CK(clk), .R(rst_n), .D(n425), .Q(bimc_ecc_correctable_error_cnt[4]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[5] ( .CK(clk), .R(rst_n), .D(n424), .Q(bimc_ecc_correctable_error_cnt[5]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[6] ( .CK(clk), .R(rst_n), .D(n423), .Q(bimc_ecc_correctable_error_cnt[6]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[7] ( .CK(clk), .R(rst_n), .D(n422), .Q(bimc_ecc_correctable_error_cnt[7]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[8] ( .CK(clk), .R(rst_n), .D(n421), .Q(bimc_ecc_correctable_error_cnt[8]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[9] ( .CK(clk), .R(rst_n), .D(n420), .Q(bimc_ecc_correctable_error_cnt[9]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[10] ( .CK(clk), .R(rst_n), .D(n419), .Q(bimc_ecc_correctable_error_cnt[10]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[11] ( .CK(clk), .R(rst_n), .D(n418), .Q(bimc_ecc_correctable_error_cnt[11]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[12] ( .CK(clk), .R(rst_n), .D(n417), .Q(bimc_ecc_correctable_error_cnt[12]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[13] ( .CK(clk), .R(rst_n), .D(n416), .Q(bimc_ecc_correctable_error_cnt[13]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[14] ( .CK(clk), .R(rst_n), .D(n415), .Q(bimc_ecc_correctable_error_cnt[14]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[15] ( .CK(clk), .R(rst_n), .D(n414), .Q(bimc_ecc_correctable_error_cnt[15]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[16] ( .CK(clk), .R(rst_n), .D(n413), .Q(bimc_ecc_correctable_error_cnt[16]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[17] ( .CK(clk), .R(rst_n), .D(n412), .Q(bimc_ecc_correctable_error_cnt[17]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[18] ( .CK(clk), .R(rst_n), .D(n411), .Q(bimc_ecc_correctable_error_cnt[18]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[19] ( .CK(clk), .R(rst_n), .D(n410), .Q(bimc_ecc_correctable_error_cnt[19]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[20] ( .CK(clk), .R(rst_n), .D(n409), .Q(bimc_ecc_correctable_error_cnt[20]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[21] ( .CK(clk), .R(rst_n), .D(n408), .Q(bimc_ecc_correctable_error_cnt[21]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[22] ( .CK(clk), .R(rst_n), .D(n407), .Q(bimc_ecc_correctable_error_cnt[22]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[23] ( .CK(clk), .R(rst_n), .D(n406), .Q(bimc_ecc_correctable_error_cnt[23]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[24] ( .CK(clk), .R(rst_n), .D(n405), .Q(bimc_ecc_correctable_error_cnt[24]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[25] ( .CK(clk), .R(rst_n), .D(n404), .Q(bimc_ecc_correctable_error_cnt[25]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[26] ( .CK(clk), .R(rst_n), .D(n403), .Q(bimc_ecc_correctable_error_cnt[26]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[27] ( .CK(clk), .R(rst_n), .D(n402), .Q(bimc_ecc_correctable_error_cnt[27]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[28] ( .CK(clk), .R(rst_n), .D(n401), .Q(bimc_ecc_correctable_error_cnt[28]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[29] ( .CK(clk), .R(rst_n), .D(n400), .Q(bimc_ecc_correctable_error_cnt[29]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[30] ( .CK(clk), .R(rst_n), .D(n399), .Q(bimc_ecc_correctable_error_cnt[30]), .QN( ));
Q_FDP1 \bimc_ecc_correctable_error_cnt_REG[31] ( .CK(clk), .R(rst_n), .D(n398), .Q(bimc_ecc_correctable_error_cnt[31]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[0] ( .CK(clk), .R(rst_n), .D(n238), .Q(bimc_ecc_uncorrectable_error_cnt[0]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[1] ( .CK(clk), .R(rst_n), .D(n237), .Q(bimc_ecc_uncorrectable_error_cnt[1]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[2] ( .CK(clk), .R(rst_n), .D(n236), .Q(bimc_ecc_uncorrectable_error_cnt[2]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[3] ( .CK(clk), .R(rst_n), .D(n235), .Q(bimc_ecc_uncorrectable_error_cnt[3]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[4] ( .CK(clk), .R(rst_n), .D(n234), .Q(bimc_ecc_uncorrectable_error_cnt[4]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[5] ( .CK(clk), .R(rst_n), .D(n233), .Q(bimc_ecc_uncorrectable_error_cnt[5]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[6] ( .CK(clk), .R(rst_n), .D(n232), .Q(bimc_ecc_uncorrectable_error_cnt[6]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[7] ( .CK(clk), .R(rst_n), .D(n231), .Q(bimc_ecc_uncorrectable_error_cnt[7]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[8] ( .CK(clk), .R(rst_n), .D(n230), .Q(bimc_ecc_uncorrectable_error_cnt[8]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[9] ( .CK(clk), .R(rst_n), .D(n229), .Q(bimc_ecc_uncorrectable_error_cnt[9]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[10] ( .CK(clk), .R(rst_n), .D(n228), .Q(bimc_ecc_uncorrectable_error_cnt[10]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[11] ( .CK(clk), .R(rst_n), .D(n227), .Q(bimc_ecc_uncorrectable_error_cnt[11]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[12] ( .CK(clk), .R(rst_n), .D(n226), .Q(bimc_ecc_uncorrectable_error_cnt[12]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[13] ( .CK(clk), .R(rst_n), .D(n225), .Q(bimc_ecc_uncorrectable_error_cnt[13]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[14] ( .CK(clk), .R(rst_n), .D(n224), .Q(bimc_ecc_uncorrectable_error_cnt[14]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[15] ( .CK(clk), .R(rst_n), .D(n223), .Q(bimc_ecc_uncorrectable_error_cnt[15]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[16] ( .CK(clk), .R(rst_n), .D(n222), .Q(bimc_ecc_uncorrectable_error_cnt[16]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[17] ( .CK(clk), .R(rst_n), .D(n221), .Q(bimc_ecc_uncorrectable_error_cnt[17]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[18] ( .CK(clk), .R(rst_n), .D(n220), .Q(bimc_ecc_uncorrectable_error_cnt[18]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[19] ( .CK(clk), .R(rst_n), .D(n219), .Q(bimc_ecc_uncorrectable_error_cnt[19]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[20] ( .CK(clk), .R(rst_n), .D(n218), .Q(bimc_ecc_uncorrectable_error_cnt[20]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[21] ( .CK(clk), .R(rst_n), .D(n217), .Q(bimc_ecc_uncorrectable_error_cnt[21]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[22] ( .CK(clk), .R(rst_n), .D(n216), .Q(bimc_ecc_uncorrectable_error_cnt[22]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[23] ( .CK(clk), .R(rst_n), .D(n215), .Q(bimc_ecc_uncorrectable_error_cnt[23]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[24] ( .CK(clk), .R(rst_n), .D(n214), .Q(bimc_ecc_uncorrectable_error_cnt[24]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[25] ( .CK(clk), .R(rst_n), .D(n213), .Q(bimc_ecc_uncorrectable_error_cnt[25]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[26] ( .CK(clk), .R(rst_n), .D(n212), .Q(bimc_ecc_uncorrectable_error_cnt[26]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[27] ( .CK(clk), .R(rst_n), .D(n211), .Q(bimc_ecc_uncorrectable_error_cnt[27]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[28] ( .CK(clk), .R(rst_n), .D(n210), .Q(bimc_ecc_uncorrectable_error_cnt[28]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[29] ( .CK(clk), .R(rst_n), .D(n209), .Q(bimc_ecc_uncorrectable_error_cnt[29]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[30] ( .CK(clk), .R(rst_n), .D(n208), .Q(bimc_ecc_uncorrectable_error_cnt[30]), .QN( ));
Q_FDP1 \bimc_ecc_uncorrectable_error_cnt_REG[31] ( .CK(clk), .R(rst_n), .D(n207), .Q(bimc_ecc_uncorrectable_error_cnt[31]), .QN( ));
Q_FDP1 bimc_cmd2_sent_REG  ( .CK(clk), .R(rst_n), .D(n684), .Q(bimc_cmd2_sent), .QN( ));
Q_FDP1 bimc_eccpar_debug_sent_REG  ( .CK(clk), .R(rst_n), .D(n206), .Q(bimc_eccpar_debug_sent), .QN( ));
Q_MX02 U505 ( .S(n202), .A0(n203), .A1(i_bimc_eccpar_debug[23]), .Z(n206));
Q_AN02 U506 ( .A0(n1026), .A1(n557), .Z(n207));
Q_AN02 U507 ( .A0(n1026), .A1(n558), .Z(n208));
Q_AN02 U508 ( .A0(n1026), .A1(n559), .Z(n209));
Q_AN02 U509 ( .A0(n1026), .A1(n560), .Z(n210));
Q_AN02 U510 ( .A0(n1026), .A1(n561), .Z(n211));
Q_AN02 U511 ( .A0(n1026), .A1(n562), .Z(n212));
Q_AN02 U512 ( .A0(n1026), .A1(n563), .Z(n213));
Q_AN02 U513 ( .A0(n1026), .A1(n564), .Z(n214));
Q_AN02 U514 ( .A0(n1026), .A1(n565), .Z(n215));
Q_AN02 U515 ( .A0(n1026), .A1(n566), .Z(n216));
Q_AN02 U516 ( .A0(n1026), .A1(n567), .Z(n217));
Q_AN02 U517 ( .A0(n1026), .A1(n568), .Z(n218));
Q_AN02 U518 ( .A0(n1026), .A1(n569), .Z(n219));
Q_AN02 U519 ( .A0(n1026), .A1(n570), .Z(n220));
Q_AN02 U520 ( .A0(n1026), .A1(n571), .Z(n221));
Q_AN02 U521 ( .A0(n1026), .A1(n572), .Z(n222));
Q_AN02 U522 ( .A0(n1026), .A1(n573), .Z(n223));
Q_AN02 U523 ( .A0(n1026), .A1(n574), .Z(n224));
Q_AN02 U524 ( .A0(n1026), .A1(n575), .Z(n225));
Q_AN02 U525 ( .A0(n1026), .A1(n576), .Z(n226));
Q_AN02 U526 ( .A0(n1026), .A1(n577), .Z(n227));
Q_AN02 U527 ( .A0(n1026), .A1(n578), .Z(n228));
Q_AN02 U528 ( .A0(n1026), .A1(n579), .Z(n229));
Q_AN02 U529 ( .A0(n1026), .A1(n580), .Z(n230));
Q_AN02 U530 ( .A0(n1026), .A1(n581), .Z(n231));
Q_AN02 U531 ( .A0(n1026), .A1(n582), .Z(n232));
Q_AN02 U532 ( .A0(n1026), .A1(n583), .Z(n233));
Q_AN02 U533 ( .A0(n1026), .A1(n584), .Z(n234));
Q_AN02 U534 ( .A0(n1026), .A1(n585), .Z(n235));
Q_AN02 U535 ( .A0(n1026), .A1(n586), .Z(n236));
Q_AN02 U536 ( .A0(n1026), .A1(n587), .Z(n237));
Q_AN02 U537 ( .A0(n1026), .A1(n588), .Z(n238));
Q_AN02 U538 ( .A0(n1028), .A1(n271), .Z(n239));
Q_AN02 U539 ( .A0(n1028), .A1(n272), .Z(n240));
Q_AN02 U540 ( .A0(n1028), .A1(n273), .Z(n241));
Q_AN02 U541 ( .A0(n1028), .A1(n274), .Z(n242));
Q_AN02 U542 ( .A0(n1028), .A1(n275), .Z(n243));
Q_AN02 U543 ( .A0(n1028), .A1(n276), .Z(n244));
Q_AN02 U544 ( .A0(n1028), .A1(n277), .Z(n245));
Q_AN02 U545 ( .A0(n1028), .A1(n278), .Z(n246));
Q_AN02 U546 ( .A0(n1028), .A1(n279), .Z(n247));
Q_AN02 U547 ( .A0(n1028), .A1(n280), .Z(n248));
Q_AN02 U548 ( .A0(n1028), .A1(n281), .Z(n249));
Q_AN02 U549 ( .A0(n1028), .A1(n282), .Z(n250));
Q_AN02 U550 ( .A0(n1028), .A1(n283), .Z(n251));
Q_AN02 U551 ( .A0(n1028), .A1(n284), .Z(n252));
Q_AN02 U552 ( .A0(n1028), .A1(n285), .Z(n253));
Q_AN02 U553 ( .A0(n1028), .A1(n286), .Z(n254));
Q_AN02 U554 ( .A0(n1028), .A1(n287), .Z(n255));
Q_AN02 U555 ( .A0(n1028), .A1(n288), .Z(n256));
Q_AN02 U556 ( .A0(n1028), .A1(n289), .Z(n257));
Q_AN02 U557 ( .A0(n1028), .A1(n290), .Z(n258));
Q_AN02 U558 ( .A0(n1028), .A1(n291), .Z(n259));
Q_AN02 U559 ( .A0(n1028), .A1(n292), .Z(n260));
Q_AN02 U560 ( .A0(n1028), .A1(n293), .Z(n261));
Q_AN02 U561 ( .A0(n1028), .A1(n294), .Z(n262));
Q_AN02 U562 ( .A0(n1028), .A1(n295), .Z(n263));
Q_AN02 U563 ( .A0(n1028), .A1(n296), .Z(n264));
Q_AN02 U564 ( .A0(n1028), .A1(n297), .Z(n265));
Q_AN02 U565 ( .A0(n1028), .A1(n298), .Z(n266));
Q_AN02 U566 ( .A0(n1028), .A1(n299), .Z(n267));
Q_AN02 U567 ( .A0(n1028), .A1(n300), .Z(n268));
Q_AN02 U568 ( .A0(n1028), .A1(n301), .Z(n269));
Q_AN02 U569 ( .A0(n1028), .A1(n302), .Z(n270));
Q_MX02 U570 ( .S(debug_write_en), .A0(n303), .A1(o_bimc_parity_error_cnt[31]), .Z(n271));
Q_MX02 U571 ( .S(debug_write_en), .A0(n304), .A1(o_bimc_parity_error_cnt[30]), .Z(n272));
Q_MX02 U572 ( .S(debug_write_en), .A0(n305), .A1(o_bimc_parity_error_cnt[29]), .Z(n273));
Q_MX02 U573 ( .S(debug_write_en), .A0(n306), .A1(o_bimc_parity_error_cnt[28]), .Z(n274));
Q_MX02 U574 ( .S(debug_write_en), .A0(n307), .A1(o_bimc_parity_error_cnt[27]), .Z(n275));
Q_MX02 U575 ( .S(debug_write_en), .A0(n308), .A1(o_bimc_parity_error_cnt[26]), .Z(n276));
Q_MX02 U576 ( .S(debug_write_en), .A0(n309), .A1(o_bimc_parity_error_cnt[25]), .Z(n277));
Q_MX02 U577 ( .S(debug_write_en), .A0(n310), .A1(o_bimc_parity_error_cnt[24]), .Z(n278));
Q_MX02 U578 ( .S(debug_write_en), .A0(n311), .A1(o_bimc_parity_error_cnt[23]), .Z(n279));
Q_MX02 U579 ( .S(debug_write_en), .A0(n312), .A1(o_bimc_parity_error_cnt[22]), .Z(n280));
Q_MX02 U580 ( .S(debug_write_en), .A0(n313), .A1(o_bimc_parity_error_cnt[21]), .Z(n281));
Q_MX02 U581 ( .S(debug_write_en), .A0(n314), .A1(o_bimc_parity_error_cnt[20]), .Z(n282));
Q_MX02 U582 ( .S(debug_write_en), .A0(n315), .A1(o_bimc_parity_error_cnt[19]), .Z(n283));
Q_MX02 U583 ( .S(debug_write_en), .A0(n316), .A1(o_bimc_parity_error_cnt[18]), .Z(n284));
Q_MX02 U584 ( .S(debug_write_en), .A0(n317), .A1(o_bimc_parity_error_cnt[17]), .Z(n285));
Q_MX02 U585 ( .S(debug_write_en), .A0(n318), .A1(o_bimc_parity_error_cnt[16]), .Z(n286));
Q_MX02 U586 ( .S(debug_write_en), .A0(n319), .A1(o_bimc_parity_error_cnt[15]), .Z(n287));
Q_MX02 U587 ( .S(debug_write_en), .A0(n320), .A1(o_bimc_parity_error_cnt[14]), .Z(n288));
Q_MX02 U588 ( .S(debug_write_en), .A0(n321), .A1(o_bimc_parity_error_cnt[13]), .Z(n289));
Q_MX02 U589 ( .S(debug_write_en), .A0(n322), .A1(o_bimc_parity_error_cnt[12]), .Z(n290));
Q_MX02 U590 ( .S(debug_write_en), .A0(n323), .A1(o_bimc_parity_error_cnt[11]), .Z(n291));
Q_MX02 U591 ( .S(debug_write_en), .A0(n324), .A1(o_bimc_parity_error_cnt[10]), .Z(n292));
Q_MX02 U592 ( .S(debug_write_en), .A0(n325), .A1(o_bimc_parity_error_cnt[9]), .Z(n293));
Q_MX02 U593 ( .S(debug_write_en), .A0(n326), .A1(o_bimc_parity_error_cnt[8]), .Z(n294));
Q_MX02 U594 ( .S(debug_write_en), .A0(n327), .A1(o_bimc_parity_error_cnt[7]), .Z(n295));
Q_MX02 U595 ( .S(debug_write_en), .A0(n328), .A1(o_bimc_parity_error_cnt[6]), .Z(n296));
Q_MX02 U596 ( .S(debug_write_en), .A0(n329), .A1(o_bimc_parity_error_cnt[5]), .Z(n297));
Q_MX02 U597 ( .S(debug_write_en), .A0(n330), .A1(o_bimc_parity_error_cnt[4]), .Z(n298));
Q_MX02 U598 ( .S(debug_write_en), .A0(n331), .A1(o_bimc_parity_error_cnt[3]), .Z(n299));
Q_MX02 U599 ( .S(debug_write_en), .A0(n332), .A1(o_bimc_parity_error_cnt[2]), .Z(n300));
Q_MX02 U600 ( .S(debug_write_en), .A0(n333), .A1(o_bimc_parity_error_cnt[1]), .Z(n301));
Q_MX02 U601 ( .S(debug_write_en), .A0(n334), .A1(o_bimc_parity_error_cnt[0]), .Z(n302));
Q_OR02 U602 ( .A0(n200), .A1(n335), .Z(n303));
Q_OR02 U603 ( .A0(n200), .A1(n337), .Z(n304));
Q_OR02 U604 ( .A0(n200), .A1(n339), .Z(n305));
Q_OR02 U605 ( .A0(n200), .A1(n341), .Z(n306));
Q_OR02 U606 ( .A0(n200), .A1(n343), .Z(n307));
Q_OR02 U607 ( .A0(n200), .A1(n345), .Z(n308));
Q_OR02 U608 ( .A0(n200), .A1(n347), .Z(n309));
Q_OR02 U609 ( .A0(n200), .A1(n349), .Z(n310));
Q_OR02 U610 ( .A0(n200), .A1(n351), .Z(n311));
Q_OR02 U611 ( .A0(n200), .A1(n353), .Z(n312));
Q_OR02 U612 ( .A0(n200), .A1(n355), .Z(n313));
Q_OR02 U613 ( .A0(n200), .A1(n357), .Z(n314));
Q_OR02 U614 ( .A0(n200), .A1(n359), .Z(n315));
Q_OR02 U615 ( .A0(n200), .A1(n361), .Z(n316));
Q_OR02 U616 ( .A0(n200), .A1(n363), .Z(n317));
Q_OR02 U617 ( .A0(n200), .A1(n365), .Z(n318));
Q_OR02 U618 ( .A0(n200), .A1(n367), .Z(n319));
Q_OR02 U619 ( .A0(n200), .A1(n369), .Z(n320));
Q_OR02 U620 ( .A0(n200), .A1(n371), .Z(n321));
Q_OR02 U621 ( .A0(n200), .A1(n373), .Z(n322));
Q_OR02 U622 ( .A0(n200), .A1(n375), .Z(n323));
Q_OR02 U623 ( .A0(n200), .A1(n377), .Z(n324));
Q_OR02 U624 ( .A0(n200), .A1(n379), .Z(n325));
Q_OR02 U625 ( .A0(n200), .A1(n381), .Z(n326));
Q_OR02 U626 ( .A0(n200), .A1(n383), .Z(n327));
Q_OR02 U627 ( .A0(n200), .A1(n385), .Z(n328));
Q_OR02 U628 ( .A0(n200), .A1(n387), .Z(n329));
Q_OR02 U629 ( .A0(n200), .A1(n389), .Z(n330));
Q_OR02 U630 ( .A0(n200), .A1(n391), .Z(n331));
Q_OR02 U631 ( .A0(n200), .A1(n393), .Z(n332));
Q_OR02 U632 ( .A0(n200), .A1(n395), .Z(n333));
Q_OR02 U633 ( .A0(n200), .A1(n397), .Z(n334));
Q_XOR2 U634 ( .A0(i_bimc_parity_error_cnt[31]), .A1(n336), .Z(n335));
Q_AD01HF U635 ( .A0(i_bimc_parity_error_cnt[30]), .B0(n338), .S(n337), .CO(n336));
Q_AD01HF U636 ( .A0(i_bimc_parity_error_cnt[29]), .B0(n340), .S(n339), .CO(n338));
Q_AD01HF U637 ( .A0(i_bimc_parity_error_cnt[28]), .B0(n342), .S(n341), .CO(n340));
Q_AD01HF U638 ( .A0(i_bimc_parity_error_cnt[27]), .B0(n344), .S(n343), .CO(n342));
Q_AD01HF U639 ( .A0(i_bimc_parity_error_cnt[26]), .B0(n346), .S(n345), .CO(n344));
Q_AD01HF U640 ( .A0(i_bimc_parity_error_cnt[25]), .B0(n348), .S(n347), .CO(n346));
Q_AD01HF U641 ( .A0(i_bimc_parity_error_cnt[24]), .B0(n350), .S(n349), .CO(n348));
Q_AD01HF U642 ( .A0(i_bimc_parity_error_cnt[23]), .B0(n352), .S(n351), .CO(n350));
Q_AD01HF U643 ( .A0(i_bimc_parity_error_cnt[22]), .B0(n354), .S(n353), .CO(n352));
Q_AD01HF U644 ( .A0(i_bimc_parity_error_cnt[21]), .B0(n356), .S(n355), .CO(n354));
Q_AD01HF U645 ( .A0(i_bimc_parity_error_cnt[20]), .B0(n358), .S(n357), .CO(n356));
Q_AD01HF U646 ( .A0(i_bimc_parity_error_cnt[19]), .B0(n360), .S(n359), .CO(n358));
Q_AD01HF U647 ( .A0(i_bimc_parity_error_cnt[18]), .B0(n362), .S(n361), .CO(n360));
Q_AD01HF U648 ( .A0(i_bimc_parity_error_cnt[17]), .B0(n364), .S(n363), .CO(n362));
Q_AD01HF U649 ( .A0(i_bimc_parity_error_cnt[16]), .B0(n366), .S(n365), .CO(n364));
Q_AD01HF U650 ( .A0(i_bimc_parity_error_cnt[15]), .B0(n368), .S(n367), .CO(n366));
Q_AD01HF U651 ( .A0(i_bimc_parity_error_cnt[14]), .B0(n370), .S(n369), .CO(n368));
Q_AD01HF U652 ( .A0(i_bimc_parity_error_cnt[13]), .B0(n372), .S(n371), .CO(n370));
Q_AD01HF U653 ( .A0(i_bimc_parity_error_cnt[12]), .B0(n374), .S(n373), .CO(n372));
Q_AD01HF U654 ( .A0(i_bimc_parity_error_cnt[11]), .B0(n376), .S(n375), .CO(n374));
Q_AD01HF U655 ( .A0(i_bimc_parity_error_cnt[10]), .B0(n378), .S(n377), .CO(n376));
Q_AD01HF U656 ( .A0(i_bimc_parity_error_cnt[9]), .B0(n380), .S(n379), .CO(n378));
Q_AD01HF U657 ( .A0(i_bimc_parity_error_cnt[8]), .B0(n382), .S(n381), .CO(n380));
Q_AD01HF U658 ( .A0(i_bimc_parity_error_cnt[7]), .B0(n384), .S(n383), .CO(n382));
Q_AD01HF U659 ( .A0(i_bimc_parity_error_cnt[6]), .B0(n386), .S(n385), .CO(n384));
Q_AD01HF U660 ( .A0(i_bimc_parity_error_cnt[5]), .B0(n388), .S(n387), .CO(n386));
Q_AD01HF U661 ( .A0(i_bimc_parity_error_cnt[4]), .B0(n390), .S(n389), .CO(n388));
Q_AD01HF U662 ( .A0(i_bimc_parity_error_cnt[3]), .B0(n392), .S(n391), .CO(n390));
Q_AD01HF U663 ( .A0(i_bimc_parity_error_cnt[2]), .B0(n394), .S(n393), .CO(n392));
Q_AD01HF U664 ( .A0(i_bimc_parity_error_cnt[1]), .B0(n396), .S(n395), .CO(n394));
Q_AD01HF U665 ( .A0(i_bimc_parity_error_cnt[0]), .B0(bimc_parity_error_cnt_parity_errors_en), .S(n397), .CO(n396));
Q_AN02 U666 ( .A0(n1027), .A1(n430), .Z(n398));
Q_AN02 U667 ( .A0(n1027), .A1(n431), .Z(n399));
Q_AN02 U668 ( .A0(n1027), .A1(n432), .Z(n400));
Q_AN02 U669 ( .A0(n1027), .A1(n433), .Z(n401));
Q_AN02 U670 ( .A0(n1027), .A1(n434), .Z(n402));
Q_AN02 U671 ( .A0(n1027), .A1(n435), .Z(n403));
Q_AN02 U672 ( .A0(n1027), .A1(n436), .Z(n404));
Q_AN02 U673 ( .A0(n1027), .A1(n437), .Z(n405));
Q_AN02 U674 ( .A0(n1027), .A1(n438), .Z(n406));
Q_AN02 U675 ( .A0(n1027), .A1(n439), .Z(n407));
Q_AN02 U676 ( .A0(n1027), .A1(n440), .Z(n408));
Q_AN02 U677 ( .A0(n1027), .A1(n441), .Z(n409));
Q_AN02 U678 ( .A0(n1027), .A1(n442), .Z(n410));
Q_AN02 U679 ( .A0(n1027), .A1(n443), .Z(n411));
Q_AN02 U680 ( .A0(n1027), .A1(n444), .Z(n412));
Q_AN02 U681 ( .A0(n1027), .A1(n445), .Z(n413));
Q_AN02 U682 ( .A0(n1027), .A1(n446), .Z(n414));
Q_AN02 U683 ( .A0(n1027), .A1(n447), .Z(n415));
Q_AN02 U684 ( .A0(n1027), .A1(n448), .Z(n416));
Q_AN02 U685 ( .A0(n1027), .A1(n449), .Z(n417));
Q_AN02 U686 ( .A0(n1027), .A1(n450), .Z(n418));
Q_AN02 U687 ( .A0(n1027), .A1(n451), .Z(n419));
Q_AN02 U688 ( .A0(n1027), .A1(n452), .Z(n420));
Q_AN02 U689 ( .A0(n1027), .A1(n453), .Z(n421));
Q_AN02 U690 ( .A0(n1027), .A1(n454), .Z(n422));
Q_AN02 U691 ( .A0(n1027), .A1(n455), .Z(n423));
Q_AN02 U692 ( .A0(n1027), .A1(n456), .Z(n424));
Q_AN02 U693 ( .A0(n1027), .A1(n457), .Z(n425));
Q_AN02 U694 ( .A0(n1027), .A1(n458), .Z(n426));
Q_AN02 U695 ( .A0(n1027), .A1(n459), .Z(n427));
Q_AN02 U696 ( .A0(n1027), .A1(n460), .Z(n428));
Q_AN02 U697 ( .A0(n1027), .A1(n461), .Z(n429));
Q_MX02 U698 ( .S(debug_write_en), .A0(n462), .A1(o_bimc_ecc_correctable_error_cnt[31]), .Z(n430));
Q_MX02 U699 ( .S(debug_write_en), .A0(n463), .A1(o_bimc_ecc_correctable_error_cnt[30]), .Z(n431));
Q_MX02 U700 ( .S(debug_write_en), .A0(n464), .A1(o_bimc_ecc_correctable_error_cnt[29]), .Z(n432));
Q_MX02 U701 ( .S(debug_write_en), .A0(n465), .A1(o_bimc_ecc_correctable_error_cnt[28]), .Z(n433));
Q_MX02 U702 ( .S(debug_write_en), .A0(n466), .A1(o_bimc_ecc_correctable_error_cnt[27]), .Z(n434));
Q_MX02 U703 ( .S(debug_write_en), .A0(n467), .A1(o_bimc_ecc_correctable_error_cnt[26]), .Z(n435));
Q_MX02 U704 ( .S(debug_write_en), .A0(n468), .A1(o_bimc_ecc_correctable_error_cnt[25]), .Z(n436));
Q_MX02 U705 ( .S(debug_write_en), .A0(n469), .A1(o_bimc_ecc_correctable_error_cnt[24]), .Z(n437));
Q_MX02 U706 ( .S(debug_write_en), .A0(n470), .A1(o_bimc_ecc_correctable_error_cnt[23]), .Z(n438));
Q_MX02 U707 ( .S(debug_write_en), .A0(n471), .A1(o_bimc_ecc_correctable_error_cnt[22]), .Z(n439));
Q_MX02 U708 ( .S(debug_write_en), .A0(n472), .A1(o_bimc_ecc_correctable_error_cnt[21]), .Z(n440));
Q_MX02 U709 ( .S(debug_write_en), .A0(n473), .A1(o_bimc_ecc_correctable_error_cnt[20]), .Z(n441));
Q_MX02 U710 ( .S(debug_write_en), .A0(n474), .A1(o_bimc_ecc_correctable_error_cnt[19]), .Z(n442));
Q_MX02 U711 ( .S(debug_write_en), .A0(n475), .A1(o_bimc_ecc_correctable_error_cnt[18]), .Z(n443));
Q_MX02 U712 ( .S(debug_write_en), .A0(n476), .A1(o_bimc_ecc_correctable_error_cnt[17]), .Z(n444));
Q_MX02 U713 ( .S(debug_write_en), .A0(n477), .A1(o_bimc_ecc_correctable_error_cnt[16]), .Z(n445));
Q_MX02 U714 ( .S(debug_write_en), .A0(n478), .A1(o_bimc_ecc_correctable_error_cnt[15]), .Z(n446));
Q_MX02 U715 ( .S(debug_write_en), .A0(n479), .A1(o_bimc_ecc_correctable_error_cnt[14]), .Z(n447));
Q_MX02 U716 ( .S(debug_write_en), .A0(n480), .A1(o_bimc_ecc_correctable_error_cnt[13]), .Z(n448));
Q_MX02 U717 ( .S(debug_write_en), .A0(n481), .A1(o_bimc_ecc_correctable_error_cnt[12]), .Z(n449));
Q_MX02 U718 ( .S(debug_write_en), .A0(n482), .A1(o_bimc_ecc_correctable_error_cnt[11]), .Z(n450));
Q_MX02 U719 ( .S(debug_write_en), .A0(n483), .A1(o_bimc_ecc_correctable_error_cnt[10]), .Z(n451));
Q_MX02 U720 ( .S(debug_write_en), .A0(n484), .A1(o_bimc_ecc_correctable_error_cnt[9]), .Z(n452));
Q_MX02 U721 ( .S(debug_write_en), .A0(n485), .A1(o_bimc_ecc_correctable_error_cnt[8]), .Z(n453));
Q_MX02 U722 ( .S(debug_write_en), .A0(n486), .A1(o_bimc_ecc_correctable_error_cnt[7]), .Z(n454));
Q_MX02 U723 ( .S(debug_write_en), .A0(n487), .A1(o_bimc_ecc_correctable_error_cnt[6]), .Z(n455));
Q_MX02 U724 ( .S(debug_write_en), .A0(n488), .A1(o_bimc_ecc_correctable_error_cnt[5]), .Z(n456));
Q_MX02 U725 ( .S(debug_write_en), .A0(n489), .A1(o_bimc_ecc_correctable_error_cnt[4]), .Z(n457));
Q_MX02 U726 ( .S(debug_write_en), .A0(n490), .A1(o_bimc_ecc_correctable_error_cnt[3]), .Z(n458));
Q_MX02 U727 ( .S(debug_write_en), .A0(n491), .A1(o_bimc_ecc_correctable_error_cnt[2]), .Z(n459));
Q_MX02 U728 ( .S(debug_write_en), .A0(n492), .A1(o_bimc_ecc_correctable_error_cnt[1]), .Z(n460));
Q_MX02 U729 ( .S(debug_write_en), .A0(n493), .A1(o_bimc_ecc_correctable_error_cnt[0]), .Z(n461));
Q_OR02 U730 ( .A0(n201), .A1(n494), .Z(n462));
Q_OR02 U731 ( .A0(n201), .A1(n496), .Z(n463));
Q_OR02 U732 ( .A0(n201), .A1(n498), .Z(n464));
Q_OR02 U733 ( .A0(n201), .A1(n500), .Z(n465));
Q_OR02 U734 ( .A0(n201), .A1(n502), .Z(n466));
Q_OR02 U735 ( .A0(n201), .A1(n504), .Z(n467));
Q_OR02 U736 ( .A0(n201), .A1(n506), .Z(n468));
Q_OR02 U737 ( .A0(n201), .A1(n508), .Z(n469));
Q_OR02 U738 ( .A0(n201), .A1(n510), .Z(n470));
Q_OR02 U739 ( .A0(n201), .A1(n512), .Z(n471));
Q_OR02 U740 ( .A0(n201), .A1(n514), .Z(n472));
Q_OR02 U741 ( .A0(n201), .A1(n516), .Z(n473));
Q_OR02 U742 ( .A0(n201), .A1(n518), .Z(n474));
Q_OR02 U743 ( .A0(n201), .A1(n520), .Z(n475));
Q_OR02 U744 ( .A0(n201), .A1(n522), .Z(n476));
Q_OR02 U745 ( .A0(n201), .A1(n524), .Z(n477));
Q_OR02 U746 ( .A0(n201), .A1(n526), .Z(n478));
Q_OR02 U747 ( .A0(n201), .A1(n528), .Z(n479));
Q_OR02 U748 ( .A0(n201), .A1(n530), .Z(n480));
Q_OR02 U749 ( .A0(n201), .A1(n532), .Z(n481));
Q_OR02 U750 ( .A0(n201), .A1(n534), .Z(n482));
Q_OR02 U751 ( .A0(n201), .A1(n536), .Z(n483));
Q_OR02 U752 ( .A0(n201), .A1(n538), .Z(n484));
Q_OR02 U753 ( .A0(n201), .A1(n540), .Z(n485));
Q_OR02 U754 ( .A0(n201), .A1(n542), .Z(n486));
Q_OR02 U755 ( .A0(n201), .A1(n544), .Z(n487));
Q_OR02 U756 ( .A0(n201), .A1(n546), .Z(n488));
Q_OR02 U757 ( .A0(n201), .A1(n548), .Z(n489));
Q_OR02 U758 ( .A0(n201), .A1(n550), .Z(n490));
Q_OR02 U759 ( .A0(n201), .A1(n552), .Z(n491));
Q_OR02 U760 ( .A0(n201), .A1(n554), .Z(n492));
Q_OR02 U761 ( .A0(n201), .A1(n556), .Z(n493));
Q_XOR2 U762 ( .A0(i_bimc_ecc_correctable_error_cnt[31]), .A1(n495), .Z(n494));
Q_AD01HF U763 ( .A0(i_bimc_ecc_correctable_error_cnt[30]), .B0(n497), .S(n496), .CO(n495));
Q_AD01HF U764 ( .A0(i_bimc_ecc_correctable_error_cnt[29]), .B0(n499), .S(n498), .CO(n497));
Q_AD01HF U765 ( .A0(i_bimc_ecc_correctable_error_cnt[28]), .B0(n501), .S(n500), .CO(n499));
Q_AD01HF U766 ( .A0(i_bimc_ecc_correctable_error_cnt[27]), .B0(n503), .S(n502), .CO(n501));
Q_AD01HF U767 ( .A0(i_bimc_ecc_correctable_error_cnt[26]), .B0(n505), .S(n504), .CO(n503));
Q_AD01HF U768 ( .A0(i_bimc_ecc_correctable_error_cnt[25]), .B0(n507), .S(n506), .CO(n505));
Q_AD01HF U769 ( .A0(i_bimc_ecc_correctable_error_cnt[24]), .B0(n509), .S(n508), .CO(n507));
Q_AD01HF U770 ( .A0(i_bimc_ecc_correctable_error_cnt[23]), .B0(n511), .S(n510), .CO(n509));
Q_AD01HF U771 ( .A0(i_bimc_ecc_correctable_error_cnt[22]), .B0(n513), .S(n512), .CO(n511));
Q_AD01HF U772 ( .A0(i_bimc_ecc_correctable_error_cnt[21]), .B0(n515), .S(n514), .CO(n513));
Q_AD01HF U773 ( .A0(i_bimc_ecc_correctable_error_cnt[20]), .B0(n517), .S(n516), .CO(n515));
Q_AD01HF U774 ( .A0(i_bimc_ecc_correctable_error_cnt[19]), .B0(n519), .S(n518), .CO(n517));
Q_AD01HF U775 ( .A0(i_bimc_ecc_correctable_error_cnt[18]), .B0(n521), .S(n520), .CO(n519));
Q_AD01HF U776 ( .A0(i_bimc_ecc_correctable_error_cnt[17]), .B0(n523), .S(n522), .CO(n521));
Q_AD01HF U777 ( .A0(i_bimc_ecc_correctable_error_cnt[16]), .B0(n525), .S(n524), .CO(n523));
Q_AD01HF U778 ( .A0(i_bimc_ecc_correctable_error_cnt[15]), .B0(n527), .S(n526), .CO(n525));
Q_AD01HF U779 ( .A0(i_bimc_ecc_correctable_error_cnt[14]), .B0(n529), .S(n528), .CO(n527));
Q_AD01HF U780 ( .A0(i_bimc_ecc_correctable_error_cnt[13]), .B0(n531), .S(n530), .CO(n529));
Q_AD01HF U781 ( .A0(i_bimc_ecc_correctable_error_cnt[12]), .B0(n533), .S(n532), .CO(n531));
Q_AD01HF U782 ( .A0(i_bimc_ecc_correctable_error_cnt[11]), .B0(n535), .S(n534), .CO(n533));
Q_AD01HF U783 ( .A0(i_bimc_ecc_correctable_error_cnt[10]), .B0(n537), .S(n536), .CO(n535));
Q_AD01HF U784 ( .A0(i_bimc_ecc_correctable_error_cnt[9]), .B0(n539), .S(n538), .CO(n537));
Q_AD01HF U785 ( .A0(i_bimc_ecc_correctable_error_cnt[8]), .B0(n541), .S(n540), .CO(n539));
Q_AD01HF U786 ( .A0(i_bimc_ecc_correctable_error_cnt[7]), .B0(n543), .S(n542), .CO(n541));
Q_AD01HF U787 ( .A0(i_bimc_ecc_correctable_error_cnt[6]), .B0(n545), .S(n544), .CO(n543));
Q_AD01HF U788 ( .A0(i_bimc_ecc_correctable_error_cnt[5]), .B0(n547), .S(n546), .CO(n545));
Q_AD01HF U789 ( .A0(i_bimc_ecc_correctable_error_cnt[4]), .B0(n549), .S(n548), .CO(n547));
Q_AD01HF U790 ( .A0(i_bimc_ecc_correctable_error_cnt[3]), .B0(n551), .S(n550), .CO(n549));
Q_AD01HF U791 ( .A0(i_bimc_ecc_correctable_error_cnt[2]), .B0(n553), .S(n552), .CO(n551));
Q_AD01HF U792 ( .A0(i_bimc_ecc_correctable_error_cnt[1]), .B0(n555), .S(n554), .CO(n553));
Q_AD01HF U793 ( .A0(i_bimc_ecc_correctable_error_cnt[0]), .B0(bimc_ecc_correctable_error_cnt_correctable_ecc_en), .S(n556), .CO(n555));
Q_MX02 U794 ( .S(debug_write_en), .A0(n589), .A1(o_bimc_ecc_uncorrectable_error_cnt[31]), .Z(n557));
Q_MX02 U795 ( .S(debug_write_en), .A0(n590), .A1(o_bimc_ecc_uncorrectable_error_cnt[30]), .Z(n558));
Q_MX02 U796 ( .S(debug_write_en), .A0(n591), .A1(o_bimc_ecc_uncorrectable_error_cnt[29]), .Z(n559));
Q_MX02 U797 ( .S(debug_write_en), .A0(n592), .A1(o_bimc_ecc_uncorrectable_error_cnt[28]), .Z(n560));
Q_MX02 U798 ( .S(debug_write_en), .A0(n593), .A1(o_bimc_ecc_uncorrectable_error_cnt[27]), .Z(n561));
Q_MX02 U799 ( .S(debug_write_en), .A0(n594), .A1(o_bimc_ecc_uncorrectable_error_cnt[26]), .Z(n562));
Q_MX02 U800 ( .S(debug_write_en), .A0(n595), .A1(o_bimc_ecc_uncorrectable_error_cnt[25]), .Z(n563));
Q_MX02 U801 ( .S(debug_write_en), .A0(n596), .A1(o_bimc_ecc_uncorrectable_error_cnt[24]), .Z(n564));
Q_MX02 U802 ( .S(debug_write_en), .A0(n597), .A1(o_bimc_ecc_uncorrectable_error_cnt[23]), .Z(n565));
Q_MX02 U803 ( .S(debug_write_en), .A0(n598), .A1(o_bimc_ecc_uncorrectable_error_cnt[22]), .Z(n566));
Q_MX02 U804 ( .S(debug_write_en), .A0(n599), .A1(o_bimc_ecc_uncorrectable_error_cnt[21]), .Z(n567));
Q_MX02 U805 ( .S(debug_write_en), .A0(n600), .A1(o_bimc_ecc_uncorrectable_error_cnt[20]), .Z(n568));
Q_MX02 U806 ( .S(debug_write_en), .A0(n601), .A1(o_bimc_ecc_uncorrectable_error_cnt[19]), .Z(n569));
Q_MX02 U807 ( .S(debug_write_en), .A0(n602), .A1(o_bimc_ecc_uncorrectable_error_cnt[18]), .Z(n570));
Q_MX02 U808 ( .S(debug_write_en), .A0(n603), .A1(o_bimc_ecc_uncorrectable_error_cnt[17]), .Z(n571));
Q_MX02 U809 ( .S(debug_write_en), .A0(n604), .A1(o_bimc_ecc_uncorrectable_error_cnt[16]), .Z(n572));
Q_MX02 U810 ( .S(debug_write_en), .A0(n605), .A1(o_bimc_ecc_uncorrectable_error_cnt[15]), .Z(n573));
Q_MX02 U811 ( .S(debug_write_en), .A0(n606), .A1(o_bimc_ecc_uncorrectable_error_cnt[14]), .Z(n574));
Q_MX02 U812 ( .S(debug_write_en), .A0(n607), .A1(o_bimc_ecc_uncorrectable_error_cnt[13]), .Z(n575));
Q_MX02 U813 ( .S(debug_write_en), .A0(n608), .A1(o_bimc_ecc_uncorrectable_error_cnt[12]), .Z(n576));
Q_MX02 U814 ( .S(debug_write_en), .A0(n609), .A1(o_bimc_ecc_uncorrectable_error_cnt[11]), .Z(n577));
Q_MX02 U815 ( .S(debug_write_en), .A0(n610), .A1(o_bimc_ecc_uncorrectable_error_cnt[10]), .Z(n578));
Q_MX02 U816 ( .S(debug_write_en), .A0(n611), .A1(o_bimc_ecc_uncorrectable_error_cnt[9]), .Z(n579));
Q_MX02 U817 ( .S(debug_write_en), .A0(n612), .A1(o_bimc_ecc_uncorrectable_error_cnt[8]), .Z(n580));
Q_MX02 U818 ( .S(debug_write_en), .A0(n613), .A1(o_bimc_ecc_uncorrectable_error_cnt[7]), .Z(n581));
Q_MX02 U819 ( .S(debug_write_en), .A0(n614), .A1(o_bimc_ecc_uncorrectable_error_cnt[6]), .Z(n582));
Q_MX02 U820 ( .S(debug_write_en), .A0(n615), .A1(o_bimc_ecc_uncorrectable_error_cnt[5]), .Z(n583));
Q_MX02 U821 ( .S(debug_write_en), .A0(n616), .A1(o_bimc_ecc_uncorrectable_error_cnt[4]), .Z(n584));
Q_MX02 U822 ( .S(debug_write_en), .A0(n617), .A1(o_bimc_ecc_uncorrectable_error_cnt[3]), .Z(n585));
Q_MX02 U823 ( .S(debug_write_en), .A0(n618), .A1(o_bimc_ecc_uncorrectable_error_cnt[2]), .Z(n586));
Q_MX02 U824 ( .S(debug_write_en), .A0(n619), .A1(o_bimc_ecc_uncorrectable_error_cnt[1]), .Z(n587));
Q_MX02 U825 ( .S(debug_write_en), .A0(n620), .A1(o_bimc_ecc_uncorrectable_error_cnt[0]), .Z(n588));
Q_OR02 U826 ( .A0(n201), .A1(n621), .Z(n589));
Q_OR02 U827 ( .A0(n201), .A1(n623), .Z(n590));
Q_OR02 U828 ( .A0(n201), .A1(n625), .Z(n591));
Q_OR02 U829 ( .A0(n201), .A1(n627), .Z(n592));
Q_OR02 U830 ( .A0(n201), .A1(n629), .Z(n593));
Q_OR02 U831 ( .A0(n201), .A1(n631), .Z(n594));
Q_OR02 U832 ( .A0(n201), .A1(n633), .Z(n595));
Q_OR02 U833 ( .A0(n201), .A1(n635), .Z(n596));
Q_OR02 U834 ( .A0(n201), .A1(n637), .Z(n597));
Q_OR02 U835 ( .A0(n201), .A1(n639), .Z(n598));
Q_OR02 U836 ( .A0(n201), .A1(n641), .Z(n599));
Q_OR02 U837 ( .A0(n201), .A1(n643), .Z(n600));
Q_OR02 U838 ( .A0(n201), .A1(n645), .Z(n601));
Q_OR02 U839 ( .A0(n201), .A1(n647), .Z(n602));
Q_OR02 U840 ( .A0(n201), .A1(n649), .Z(n603));
Q_OR02 U841 ( .A0(n201), .A1(n651), .Z(n604));
Q_OR02 U842 ( .A0(n201), .A1(n653), .Z(n605));
Q_OR02 U843 ( .A0(n201), .A1(n655), .Z(n606));
Q_OR02 U844 ( .A0(n201), .A1(n657), .Z(n607));
Q_OR02 U845 ( .A0(n201), .A1(n659), .Z(n608));
Q_OR02 U846 ( .A0(n201), .A1(n661), .Z(n609));
Q_OR02 U847 ( .A0(n201), .A1(n663), .Z(n610));
Q_OR02 U848 ( .A0(n201), .A1(n665), .Z(n611));
Q_OR02 U849 ( .A0(n201), .A1(n667), .Z(n612));
Q_OR02 U850 ( .A0(n201), .A1(n669), .Z(n613));
Q_OR02 U851 ( .A0(n201), .A1(n671), .Z(n614));
Q_OR02 U852 ( .A0(n201), .A1(n673), .Z(n615));
Q_OR02 U853 ( .A0(n201), .A1(n675), .Z(n616));
Q_OR02 U854 ( .A0(n201), .A1(n677), .Z(n617));
Q_OR02 U855 ( .A0(n201), .A1(n679), .Z(n618));
Q_OR02 U856 ( .A0(n201), .A1(n681), .Z(n619));
Q_OR02 U857 ( .A0(n201), .A1(n683), .Z(n620));
Q_XOR2 U858 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[31]), .A1(n622), .Z(n621));
Q_AD01HF U859 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[30]), .B0(n624), .S(n623), .CO(n622));
Q_AD01HF U860 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[29]), .B0(n626), .S(n625), .CO(n624));
Q_AD01HF U861 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[28]), .B0(n628), .S(n627), .CO(n626));
Q_AD01HF U862 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[27]), .B0(n630), .S(n629), .CO(n628));
Q_AD01HF U863 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[26]), .B0(n632), .S(n631), .CO(n630));
Q_AD01HF U864 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[25]), .B0(n634), .S(n633), .CO(n632));
Q_AD01HF U865 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[24]), .B0(n636), .S(n635), .CO(n634));
Q_AD01HF U866 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[23]), .B0(n638), .S(n637), .CO(n636));
Q_AD01HF U867 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[22]), .B0(n640), .S(n639), .CO(n638));
Q_AD01HF U868 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[21]), .B0(n642), .S(n641), .CO(n640));
Q_AD01HF U869 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[20]), .B0(n644), .S(n643), .CO(n642));
Q_AD01HF U870 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[19]), .B0(n646), .S(n645), .CO(n644));
Q_AD01HF U871 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[18]), .B0(n648), .S(n647), .CO(n646));
Q_AD01HF U872 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[17]), .B0(n650), .S(n649), .CO(n648));
Q_AD01HF U873 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[16]), .B0(n652), .S(n651), .CO(n650));
Q_AD01HF U874 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[15]), .B0(n654), .S(n653), .CO(n652));
Q_AD01HF U875 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[14]), .B0(n656), .S(n655), .CO(n654));
Q_AD01HF U876 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[13]), .B0(n658), .S(n657), .CO(n656));
Q_AD01HF U877 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[12]), .B0(n660), .S(n659), .CO(n658));
Q_AD01HF U878 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[11]), .B0(n662), .S(n661), .CO(n660));
Q_AD01HF U879 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[10]), .B0(n664), .S(n663), .CO(n662));
Q_AD01HF U880 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[9]), .B0(n666), .S(n665), .CO(n664));
Q_AD01HF U881 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[8]), .B0(n668), .S(n667), .CO(n666));
Q_AD01HF U882 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[7]), .B0(n670), .S(n669), .CO(n668));
Q_AD01HF U883 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[6]), .B0(n672), .S(n671), .CO(n670));
Q_AD01HF U884 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[5]), .B0(n674), .S(n673), .CO(n672));
Q_AD01HF U885 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[4]), .B0(n676), .S(n675), .CO(n674));
Q_AD01HF U886 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[3]), .B0(n678), .S(n677), .CO(n676));
Q_AD01HF U887 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[2]), .B0(n680), .S(n679), .CO(n678));
Q_AD01HF U888 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[1]), .B0(n682), .S(n681), .CO(n680));
Q_AD01HF U889 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[0]), .B0(bimc_ecc_uncorrectable_error_cnt_uncorrectable_ecc_en), .S(n683), .CO(n682));
Q_OA21 U890 ( .A0(bimc_cmd2_sent_din), .A1(i_bimc_cmd2[9]), .B0(n204), .Z(n684));
Q_AN02 U891 ( .A0(n686), .A1(n685), .Z(n200));
Q_AN03 U892 ( .A0(n689), .A1(n688), .A2(n687), .Z(n685));
Q_AN03 U893 ( .A0(n692), .A1(n691), .A2(n690), .Z(n686));
Q_AN03 U894 ( .A0(n695), .A1(n694), .A2(n693), .Z(n687));
Q_AN03 U895 ( .A0(n698), .A1(n697), .A2(n696), .Z(n688));
Q_AN03 U896 ( .A0(i_bimc_parity_error_cnt[1]), .A1(i_bimc_parity_error_cnt[0]), .A2(n699), .Z(n689));
Q_AN03 U897 ( .A0(i_bimc_parity_error_cnt[4]), .A1(i_bimc_parity_error_cnt[3]), .A2(i_bimc_parity_error_cnt[2]), .Z(n690));
Q_AN03 U898 ( .A0(i_bimc_parity_error_cnt[7]), .A1(i_bimc_parity_error_cnt[6]), .A2(i_bimc_parity_error_cnt[5]), .Z(n691));
Q_AN03 U899 ( .A0(i_bimc_parity_error_cnt[10]), .A1(i_bimc_parity_error_cnt[9]), .A2(i_bimc_parity_error_cnt[8]), .Z(n692));
Q_AN03 U900 ( .A0(i_bimc_parity_error_cnt[13]), .A1(i_bimc_parity_error_cnt[12]), .A2(i_bimc_parity_error_cnt[11]), .Z(n693));
Q_AN03 U901 ( .A0(i_bimc_parity_error_cnt[16]), .A1(i_bimc_parity_error_cnt[15]), .A2(i_bimc_parity_error_cnt[14]), .Z(n694));
Q_AN03 U902 ( .A0(i_bimc_parity_error_cnt[19]), .A1(i_bimc_parity_error_cnt[18]), .A2(i_bimc_parity_error_cnt[17]), .Z(n695));
Q_AN03 U903 ( .A0(i_bimc_parity_error_cnt[22]), .A1(i_bimc_parity_error_cnt[21]), .A2(i_bimc_parity_error_cnt[20]), .Z(n696));
Q_AN03 U904 ( .A0(i_bimc_parity_error_cnt[25]), .A1(i_bimc_parity_error_cnt[24]), .A2(i_bimc_parity_error_cnt[23]), .Z(n697));
Q_AN03 U905 ( .A0(i_bimc_parity_error_cnt[28]), .A1(i_bimc_parity_error_cnt[27]), .A2(i_bimc_parity_error_cnt[26]), .Z(n698));
Q_AN03 U906 ( .A0(i_bimc_parity_error_cnt[31]), .A1(i_bimc_parity_error_cnt[30]), .A2(i_bimc_parity_error_cnt[29]), .Z(n699));
Q_AN02 U907 ( .A0(n701), .A1(n700), .Z(n201));
Q_AN03 U908 ( .A0(n704), .A1(n703), .A2(n702), .Z(n700));
Q_AN03 U909 ( .A0(n707), .A1(n706), .A2(n705), .Z(n701));
Q_AN03 U910 ( .A0(n710), .A1(n709), .A2(n708), .Z(n702));
Q_AN03 U911 ( .A0(n713), .A1(n712), .A2(n711), .Z(n703));
Q_AN03 U912 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[1]), .A1(i_bimc_ecc_uncorrectable_error_cnt[0]), .A2(n714), .Z(n704));
Q_AN03 U913 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[4]), .A1(i_bimc_ecc_uncorrectable_error_cnt[3]), .A2(i_bimc_ecc_uncorrectable_error_cnt[2]), .Z(n705));
Q_AN03 U914 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[7]), .A1(i_bimc_ecc_uncorrectable_error_cnt[6]), .A2(i_bimc_ecc_uncorrectable_error_cnt[5]), .Z(n706));
Q_AN03 U915 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[10]), .A1(i_bimc_ecc_uncorrectable_error_cnt[9]), .A2(i_bimc_ecc_uncorrectable_error_cnt[8]), .Z(n707));
Q_AN03 U916 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[13]), .A1(i_bimc_ecc_uncorrectable_error_cnt[12]), .A2(i_bimc_ecc_uncorrectable_error_cnt[11]), .Z(n708));
Q_AN03 U917 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[16]), .A1(i_bimc_ecc_uncorrectable_error_cnt[15]), .A2(i_bimc_ecc_uncorrectable_error_cnt[14]), .Z(n709));
Q_AN03 U918 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[19]), .A1(i_bimc_ecc_uncorrectable_error_cnt[18]), .A2(i_bimc_ecc_uncorrectable_error_cnt[17]), .Z(n710));
Q_AN03 U919 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[22]), .A1(i_bimc_ecc_uncorrectable_error_cnt[21]), .A2(i_bimc_ecc_uncorrectable_error_cnt[20]), .Z(n711));
Q_AN03 U920 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[25]), .A1(i_bimc_ecc_uncorrectable_error_cnt[24]), .A2(i_bimc_ecc_uncorrectable_error_cnt[23]), .Z(n712));
Q_AN03 U921 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[28]), .A1(i_bimc_ecc_uncorrectable_error_cnt[27]), .A2(i_bimc_ecc_uncorrectable_error_cnt[26]), .Z(n713));
Q_AN03 U922 ( .A0(i_bimc_ecc_uncorrectable_error_cnt[31]), .A1(i_bimc_ecc_uncorrectable_error_cnt[30]), .A2(i_bimc_ecc_uncorrectable_error_cnt[29]), .Z(n714));
Q_XNR2 U923 ( .A0(tstate[0]), .A1(n1221), .Z(n722));
Q_OR02 U924 ( .A0(tstate[2]), .A1(n722), .Z(n723));
Q_INV U925 ( .A(n778), .Z(n724));
Q_MX02 U926 ( .S(tstate[3]), .A0(n724), .A1(n723), .Z(n715));
Q_OR02 U927 ( .A0(n725), .A1(sync_cnt[1]), .Z(n726));
Q_OR02 U928 ( .A0(sync_cnt[2]), .A1(sync_cnt[6]), .Z(n727));
Q_OR03 U929 ( .A0(n727), .A1(n726), .A2(n761), .Z(n787));
Q_OR03 U930 ( .A0(sync_cnt[4]), .A1(sync_cnt[3]), .A2(sync_cnt[5]), .Z(n761));
Q_NR02 U931 ( .A0(tstate[1]), .A1(n787), .Z(n728));
Q_OR02 U932 ( .A0(n728), .A1(tstate[0]), .Z(n729));
Q_ND02 U933 ( .A0(n9), .A1(n729), .Z(n730));
Q_OR03 U934 ( .A0(tstate[2]), .A1(n730), .A2(n1196), .Z(n780));
Q_OR02 U935 ( .A0(n1212), .A1(n787), .Z(n731));
Q_INV U936 ( .A(n754), .Z(n732));
Q_OR02 U937 ( .A0(n755), .A1(n732), .Z(n733));
Q_OR03 U938 ( .A0(n743), .A1(n758), .A2(n733), .Z(n734));
Q_OA21 U939 ( .A0(n770), .A1(n734), .B0(tstate[1]), .Z(n735));
Q_MX03 U940 ( .S0(tstate[0]), .S1(tstate[2]), .A0(n773), .A1(n735), .A2(n731), .Z(n736));
Q_OA21 U941 ( .A0(n736), .A1(tstate[3]), .B0(n780), .Z(n737));
Q_INV U942 ( .A(n737), .Z(n716));
Q_INV U943 ( .A(n787), .Z(n790));
Q_MX02 U944 ( .S(tstate[0]), .A0(n763), .A1(n773), .Z(n738));
Q_INV U945 ( .A(n738), .Z(n739));
Q_OR03 U946 ( .A0(tstate[2]), .A1(n739), .A2(n1196), .Z(n794));
Q_AO21 U947 ( .A0(tstate[0]), .A1(n773), .B0(n1201), .Z(n784));
Q_NR02 U948 ( .A0(auto_poll_ecc_par_ev), .A1(mem_wr_init_ev), .Z(n740));
Q_OA21 U949 ( .A0(cpu_transmit_ev), .A1(n740), .B0(bimc_rst_n), .Z(n744));
Q_OR02 U950 ( .A0(n758), .A1(n755), .Z(n741));
Q_OR03 U951 ( .A0(n742), .A1(n741), .A2(n744), .Z(n745));
Q_OR02 U952 ( .A0(sync_cnt[3]), .A1(sync_cnt[2]), .Z(n743));
Q_OR02 U953 ( .A0(sync_cnt[4]), .A1(n743), .Z(n742));
Q_OR02 U954 ( .A0(n1221), .A1(sync_cnt[5]), .Z(n746));
Q_OR03 U955 ( .A0(n746), .A1(n745), .A2(n1212), .Z(n747));
Q_ND02 U956 ( .A0(n747), .A1(n10), .Z(n748));
Q_OR02 U957 ( .A0(n748), .A1(tstate[2]), .Z(n749));
Q_ND02 U958 ( .A0(n784), .A1(n749), .Z(n750));
Q_OA21 U959 ( .A0(n750), .A1(tstate[3]), .B0(n794), .Z(n751));
Q_INV U960 ( .A(n751), .Z(n717));
Q_OR02 U961 ( .A0(tstate[0]), .A1(n1201), .Z(n778));
Q_OA21 U962 ( .A0(mem_wr_init_ev), .A1(n752), .B0(n753), .Z(n759));
Q_OR02 U963 ( .A0(n765), .A1(cpu_transmit_ev), .Z(n754));
Q_OR02 U964 ( .A0(n755), .A1(n754), .Z(n757));
Q_OR02 U965 ( .A0(n756), .A1(sync_cnt[1]), .Z(n755));
Q_OR02 U966 ( .A0(sync_cnt[6]), .A1(sync_cnt[0]), .Z(n758));
Q_OR03 U967 ( .A0(sync_cnt[2]), .A1(n758), .A2(n757), .Z(n760));
Q_OR03 U968 ( .A0(n760), .A1(n759), .A2(n761), .Z(n762));
Q_AO21 U969 ( .A0(n762), .A1(tstate[1]), .B0(n763), .Z(n764));
Q_AN02 U970 ( .A0(n787), .A1(n1221), .Z(n763));
Q_AN02 U971 ( .A0(n787), .A1(tstate[1]), .Z(n773));
Q_OR02 U972 ( .A0(sync_cnt[1]), .A1(n765), .Z(n767));
Q_OR03 U973 ( .A0(n766), .A1(sync_cnt[0]), .A2(n767), .Z(n771));
Q_OR02 U974 ( .A0(n768), .A1(sync_cnt[2]), .Z(n769));
Q_OR03 U975 ( .A0(n770), .A1(n769), .A2(n771), .Z(n772));
Q_OR02 U976 ( .A0(sync_cnt[5]), .A1(sync_cnt[4]), .Z(n770));
Q_AO21 U977 ( .A0(n772), .A1(n1221), .B0(n773), .Z(n774));
Q_MX02 U978 ( .S(tstate[0]), .A0(n774), .A1(n764), .Z(n775));
Q_INV U979 ( .A(n775), .Z(n776));
Q_OR02 U980 ( .A0(n776), .A1(tstate[2]), .Z(n777));
Q_ND02 U981 ( .A0(n778), .A1(n777), .Z(n779));
Q_OA21 U982 ( .A0(n779), .A1(tstate[3]), .B0(n780), .Z(n781));
Q_INV U983 ( .A(n781), .Z(n718));
Q_OR02 U984 ( .A0(n1221), .A1(n787), .Z(n782));
Q_AO21 U985 ( .A0(n1212), .A1(n782), .B0(tstate[2]), .Z(n783));
Q_ND02 U986 ( .A0(n784), .A1(n783), .Z(n785));
Q_OA21 U987 ( .A0(n785), .A1(tstate[3]), .B0(n794), .Z(n719));
Q_OR03 U988 ( .A0(tstate[2]), .A1(tstate[0]), .A2(n8), .Z(n786));
Q_ND02 U989 ( .A0(n1222), .A1(n787), .Z(n788));
Q_MX02 U990 ( .S(tstate[3]), .A0(n788), .A1(n786), .Z(n720));
Q_OR03 U991 ( .A0(n1212), .A1(n789), .A2(n790), .Z(n791));
Q_ND02 U992 ( .A0(tstate[0]), .A1(n763), .Z(n792));
Q_MX02 U993 ( .S(tstate[2]), .A0(n792), .A1(n791), .Z(n793));
Q_OA21 U994 ( .A0(n793), .A1(tstate[3]), .B0(n794), .Z(n721));
Q_AO21 U995 ( .A0(n715), .A1(tstate[0]), .B0(n802), .Z(nxt_tstate[0]));
Q_AO21 U996 ( .A0(n715), .A1(tstate[1]), .B0(n800), .Z(nxt_tstate[1]));
Q_AO21 U997 ( .A0(n715), .A1(tstate[2]), .B0(n796), .Z(nxt_tstate[2]));
Q_AN02 U998 ( .A0(n715), .A1(tstate[3]), .Z(n795));
Q_XOR2 U999 ( .A0(n718), .A1(n737), .Z(n797));
Q_AO21 U1000 ( .A0(n717), .A1(n797), .B0(n795), .Z(nxt_tstate[3]));
Q_NR02 U1001 ( .A0(n781), .A1(n716), .Z(n796));
Q_OR02 U1002 ( .A0(n797), .A1(n717), .Z(n798));
Q_ND02 U1003 ( .A0(n803), .A1(n798), .Z(n799));
Q_NR02 U1004 ( .A0(n715), .A1(n799), .Z(n800));
Q_OR02 U1005 ( .A0(n718), .A1(n751), .Z(n803));
Q_ND02 U1006 ( .A0(n781), .A1(n737), .Z(n801));
Q_OA21 U1007 ( .A0(n801), .A1(n717), .B0(n803), .Z(n802));
Q_AN03 U1008 ( .A0(n720), .A1(n804), .A2(n719), .Z(reg_send[72]));
Q_MX02 U1009 ( .S(n721), .A0(cputx_frame[72]), .A1(r_reg_send[72]), .Z(n804));
Q_MX02 U1010 ( .S(n719), .A0(n867), .A1(n805), .Z(reg_send[71]));
Q_MX02 U1011 ( .S(n720), .A0(n806), .A1(n807), .Z(n805));
Q_OR02 U1012 ( .A0(n721), .A1(bimc_eccpar_debug_memtype[3]), .Z(n806));
Q_MX02 U1013 ( .S(n721), .A0(cputx_frame[71]), .A1(r_reg_send[71]), .Z(n807));
Q_MX02 U1014 ( .S(n719), .A0(n867), .A1(n808), .Z(reg_send[70]));
Q_MX02 U1015 ( .S(n720), .A0(n809), .A1(n810), .Z(n808));
Q_OR02 U1016 ( .A0(n721), .A1(bimc_eccpar_debug_memtype[2]), .Z(n809));
Q_MX02 U1017 ( .S(n721), .A0(cputx_frame[70]), .A1(r_reg_send[70]), .Z(n810));
Q_MX02 U1018 ( .S(n719), .A0(n867), .A1(n811), .Z(reg_send[69]));
Q_MX02 U1019 ( .S(n720), .A0(n812), .A1(n813), .Z(n811));
Q_OR02 U1020 ( .A0(n721), .A1(bimc_eccpar_debug_memtype[1]), .Z(n812));
Q_MX02 U1021 ( .S(n721), .A0(cputx_frame[69]), .A1(r_reg_send[69]), .Z(n813));
Q_MX02 U1022 ( .S(n719), .A0(n867), .A1(n814), .Z(reg_send[68]));
Q_MX02 U1023 ( .S(n720), .A0(n815), .A1(n816), .Z(n814));
Q_OR02 U1024 ( .A0(n721), .A1(bimc_eccpar_debug_memtype[0]), .Z(n815));
Q_MX02 U1025 ( .S(n721), .A0(cputx_frame[68]), .A1(r_reg_send[68]), .Z(n816));
Q_MX02 U1026 ( .S(n719), .A0(n827), .A1(n817), .Z(reg_send[67]));
Q_AN02 U1027 ( .A0(n720), .A1(n818), .Z(n817));
Q_MX02 U1028 ( .S(n721), .A0(cputx_frame[67]), .A1(r_reg_send[67]), .Z(n818));
Q_MX02 U1029 ( .S(n719), .A0(n827), .A1(n819), .Z(reg_send[66]));
Q_AN02 U1030 ( .A0(n720), .A1(n820), .Z(n819));
Q_MX02 U1031 ( .S(n721), .A0(cputx_frame[66]), .A1(r_reg_send[66]), .Z(n820));
Q_MX02 U1032 ( .S(n719), .A0(n827), .A1(n821), .Z(reg_send[65]));
Q_AN02 U1033 ( .A0(n720), .A1(n822), .Z(n821));
Q_MX02 U1034 ( .S(n721), .A0(cputx_frame[65]), .A1(r_reg_send[65]), .Z(n822));
Q_MX02 U1035 ( .S(n719), .A0(n827), .A1(n823), .Z(reg_send[64]));
Q_AN02 U1036 ( .A0(n720), .A1(n824), .Z(n823));
Q_MX02 U1037 ( .S(n721), .A0(cputx_frame[64]), .A1(r_reg_send[64]), .Z(n824));
Q_MX02 U1038 ( .S(n719), .A0(n827), .A1(n825), .Z(reg_send[63]));
Q_AN02 U1039 ( .A0(n720), .A1(n826), .Z(n825));
Q_MX02 U1040 ( .S(n721), .A0(cputx_frame[63]), .A1(r_reg_send[63]), .Z(n826));
Q_MX02 U1041 ( .S(n719), .A0(n827), .A1(n828), .Z(reg_send[62]));
Q_NR02 U1042 ( .A0(n720), .A1(n721), .Z(n827));
Q_AN02 U1043 ( .A0(n720), .A1(n829), .Z(n828));
Q_MX02 U1044 ( .S(n721), .A0(cputx_frame[62]), .A1(r_reg_send[62]), .Z(n829));
Q_MX02 U1045 ( .S(n719), .A0(n867), .A1(n830), .Z(reg_send[61]));
Q_OR02 U1046 ( .A0(n916), .A1(n831), .Z(n830));
Q_MX02 U1047 ( .S(n721), .A0(cputx_frame[61]), .A1(r_reg_send[61]), .Z(n831));
Q_MX02 U1048 ( .S(n719), .A0(n916), .A1(n832), .Z(reg_send[60]));
Q_AN02 U1049 ( .A0(n720), .A1(n833), .Z(n832));
Q_MX02 U1050 ( .S(n721), .A0(cputx_frame[60]), .A1(r_reg_send[60]), .Z(n833));
Q_MX02 U1051 ( .S(n719), .A0(n867), .A1(n834), .Z(reg_send[59]));
Q_MX02 U1052 ( .S(n720), .A0(n835), .A1(n836), .Z(n834));
Q_AN02 U1053 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[11]), .Z(n835));
Q_MX02 U1054 ( .S(n721), .A0(cputx_frame[59]), .A1(r_reg_send[59]), .Z(n836));
Q_MX02 U1055 ( .S(n719), .A0(n867), .A1(n837), .Z(reg_send[58]));
Q_MX02 U1056 ( .S(n720), .A0(n838), .A1(n839), .Z(n837));
Q_AN02 U1057 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[10]), .Z(n838));
Q_MX02 U1058 ( .S(n721), .A0(cputx_frame[58]), .A1(r_reg_send[58]), .Z(n839));
Q_MX02 U1059 ( .S(n719), .A0(n867), .A1(n840), .Z(reg_send[57]));
Q_MX02 U1060 ( .S(n720), .A0(n841), .A1(n842), .Z(n840));
Q_AN02 U1061 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[9]), .Z(n841));
Q_MX02 U1062 ( .S(n721), .A0(cputx_frame[57]), .A1(r_reg_send[57]), .Z(n842));
Q_MX02 U1063 ( .S(n719), .A0(n867), .A1(n843), .Z(reg_send[56]));
Q_MX02 U1064 ( .S(n720), .A0(n844), .A1(n845), .Z(n843));
Q_AN02 U1065 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[8]), .Z(n844));
Q_MX02 U1066 ( .S(n721), .A0(cputx_frame[56]), .A1(r_reg_send[56]), .Z(n845));
Q_MX02 U1067 ( .S(n719), .A0(n867), .A1(n846), .Z(reg_send[55]));
Q_MX02 U1068 ( .S(n720), .A0(n847), .A1(n848), .Z(n846));
Q_AN02 U1069 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[7]), .Z(n847));
Q_MX02 U1070 ( .S(n721), .A0(cputx_frame[55]), .A1(r_reg_send[55]), .Z(n848));
Q_MX02 U1071 ( .S(n719), .A0(n867), .A1(n849), .Z(reg_send[54]));
Q_MX02 U1072 ( .S(n720), .A0(n850), .A1(n851), .Z(n849));
Q_AN02 U1073 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[6]), .Z(n850));
Q_MX02 U1074 ( .S(n721), .A0(cputx_frame[54]), .A1(r_reg_send[54]), .Z(n851));
Q_MX02 U1075 ( .S(n719), .A0(n867), .A1(n852), .Z(reg_send[53]));
Q_MX02 U1076 ( .S(n720), .A0(n853), .A1(n854), .Z(n852));
Q_AN02 U1077 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[5]), .Z(n853));
Q_MX02 U1078 ( .S(n721), .A0(cputx_frame[53]), .A1(r_reg_send[53]), .Z(n854));
Q_MX02 U1079 ( .S(n719), .A0(n867), .A1(n855), .Z(reg_send[52]));
Q_MX02 U1080 ( .S(n720), .A0(n856), .A1(n857), .Z(n855));
Q_AN02 U1081 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[4]), .Z(n856));
Q_MX02 U1082 ( .S(n721), .A0(cputx_frame[52]), .A1(r_reg_send[52]), .Z(n857));
Q_MX02 U1083 ( .S(n719), .A0(n867), .A1(n858), .Z(reg_send[51]));
Q_MX02 U1084 ( .S(n720), .A0(n859), .A1(n860), .Z(n858));
Q_AN02 U1085 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[3]), .Z(n859));
Q_MX02 U1086 ( .S(n721), .A0(cputx_frame[51]), .A1(r_reg_send[51]), .Z(n860));
Q_MX02 U1087 ( .S(n719), .A0(n867), .A1(n861), .Z(reg_send[50]));
Q_MX02 U1088 ( .S(n720), .A0(n862), .A1(n863), .Z(n861));
Q_AN02 U1089 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[2]), .Z(n862));
Q_MX02 U1090 ( .S(n721), .A0(cputx_frame[50]), .A1(r_reg_send[50]), .Z(n863));
Q_MX02 U1091 ( .S(n719), .A0(n867), .A1(n864), .Z(reg_send[49]));
Q_MX02 U1092 ( .S(n720), .A0(n865), .A1(n866), .Z(n864));
Q_AN02 U1093 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[1]), .Z(n865));
Q_MX02 U1094 ( .S(n721), .A0(cputx_frame[49]), .A1(r_reg_send[49]), .Z(n866));
Q_MX02 U1095 ( .S(n719), .A0(n867), .A1(n868), .Z(reg_send[48]));
Q_ND02 U1096 ( .A0(n720), .A1(n721), .Z(n867));
Q_MX02 U1097 ( .S(n720), .A0(n869), .A1(n870), .Z(n868));
Q_AN02 U1098 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[0]), .Z(n869));
Q_MX02 U1099 ( .S(n721), .A0(cputx_frame[48]), .A1(r_reg_send[48]), .Z(n870));
Q_MX02 U1100 ( .S(n719), .A0(n909), .A1(n871), .Z(reg_send[47]));
Q_AN02 U1101 ( .A0(n720), .A1(n872), .Z(n871));
Q_MX02 U1102 ( .S(n721), .A0(cputx_frame[47]), .A1(r_reg_send[47]), .Z(n872));
Q_MX02 U1103 ( .S(n719), .A0(n909), .A1(n873), .Z(reg_send[46]));
Q_AN02 U1104 ( .A0(n720), .A1(n874), .Z(n873));
Q_MX02 U1105 ( .S(n721), .A0(cputx_frame[46]), .A1(r_reg_send[46]), .Z(n874));
Q_MX02 U1106 ( .S(n719), .A0(n909), .A1(n875), .Z(reg_send[45]));
Q_AN02 U1107 ( .A0(n720), .A1(n876), .Z(n875));
Q_MX02 U1108 ( .S(n721), .A0(cputx_frame[45]), .A1(r_reg_send[45]), .Z(n876));
Q_MX02 U1109 ( .S(n719), .A0(n909), .A1(n877), .Z(reg_send[44]));
Q_AN02 U1110 ( .A0(n720), .A1(n878), .Z(n877));
Q_MX02 U1111 ( .S(n721), .A0(cputx_frame[44]), .A1(r_reg_send[44]), .Z(n878));
Q_MX02 U1112 ( .S(n719), .A0(n909), .A1(n879), .Z(reg_send[43]));
Q_MX02 U1113 ( .S(n720), .A0(n880), .A1(n881), .Z(n879));
Q_AN02 U1114 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[11]), .Z(n880));
Q_MX02 U1115 ( .S(n721), .A0(cputx_frame[43]), .A1(r_reg_send[43]), .Z(n881));
Q_MX02 U1116 ( .S(n719), .A0(n909), .A1(n882), .Z(reg_send[42]));
Q_MX02 U1117 ( .S(n720), .A0(n883), .A1(n884), .Z(n882));
Q_AN02 U1118 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[10]), .Z(n883));
Q_MX02 U1119 ( .S(n721), .A0(cputx_frame[42]), .A1(r_reg_send[42]), .Z(n884));
Q_MX02 U1120 ( .S(n719), .A0(n909), .A1(n885), .Z(reg_send[41]));
Q_MX02 U1121 ( .S(n720), .A0(n886), .A1(n887), .Z(n885));
Q_AN02 U1122 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[9]), .Z(n886));
Q_MX02 U1123 ( .S(n721), .A0(cputx_frame[41]), .A1(r_reg_send[41]), .Z(n887));
Q_MX02 U1124 ( .S(n719), .A0(n909), .A1(n888), .Z(reg_send[40]));
Q_MX02 U1125 ( .S(n720), .A0(n889), .A1(n890), .Z(n888));
Q_AN02 U1126 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[8]), .Z(n889));
Q_MX02 U1127 ( .S(n721), .A0(cputx_frame[40]), .A1(r_reg_send[40]), .Z(n890));
Q_MX02 U1128 ( .S(n719), .A0(n909), .A1(n891), .Z(reg_send[39]));
Q_MX02 U1129 ( .S(n720), .A0(n892), .A1(n893), .Z(n891));
Q_AN02 U1130 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[7]), .Z(n892));
Q_MX02 U1131 ( .S(n721), .A0(cputx_frame[39]), .A1(r_reg_send[39]), .Z(n893));
Q_MX02 U1132 ( .S(n719), .A0(n909), .A1(n894), .Z(reg_send[38]));
Q_MX02 U1133 ( .S(n720), .A0(n895), .A1(n896), .Z(n894));
Q_AN02 U1134 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[6]), .Z(n895));
Q_MX02 U1135 ( .S(n721), .A0(cputx_frame[38]), .A1(r_reg_send[38]), .Z(n896));
Q_MX02 U1136 ( .S(n719), .A0(n909), .A1(n897), .Z(reg_send[37]));
Q_MX02 U1137 ( .S(n720), .A0(n898), .A1(n899), .Z(n897));
Q_AN02 U1138 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[5]), .Z(n898));
Q_MX02 U1139 ( .S(n721), .A0(cputx_frame[37]), .A1(r_reg_send[37]), .Z(n899));
Q_MX02 U1140 ( .S(n719), .A0(n909), .A1(n900), .Z(reg_send[36]));
Q_MX02 U1141 ( .S(n720), .A0(n901), .A1(n902), .Z(n900));
Q_AN02 U1142 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[4]), .Z(n901));
Q_MX02 U1143 ( .S(n721), .A0(cputx_frame[36]), .A1(r_reg_send[36]), .Z(n902));
Q_MX02 U1144 ( .S(n719), .A0(n916), .A1(n903), .Z(reg_send[35]));
Q_MX02 U1145 ( .S(n720), .A0(n904), .A1(n905), .Z(n903));
Q_OR02 U1146 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[3]), .Z(n904));
Q_MX02 U1147 ( .S(n721), .A0(cputx_frame[35]), .A1(r_reg_send[35]), .Z(n905));
Q_MX02 U1148 ( .S(n719), .A0(n909), .A1(n906), .Z(reg_send[34]));
Q_MX02 U1149 ( .S(n720), .A0(n907), .A1(n908), .Z(n906));
Q_AN02 U1150 ( .A0(n721), .A1(bimc_eccpar_debug_memaddr[2]), .Z(n907));
Q_MX02 U1151 ( .S(n721), .A0(cputx_frame[34]), .A1(r_reg_send[34]), .Z(n908));
Q_MX02 U1152 ( .S(n719), .A0(n909), .A1(n910), .Z(reg_send[33]));
Q_AN02 U1153 ( .A0(n916), .A1(n721), .Z(n909));
Q_MX02 U1154 ( .S(n720), .A0(n911), .A1(n912), .Z(n910));
Q_OR02 U1155 ( .A0(n956), .A1(bimc_eccpar_debug_memaddr[1]), .Z(n911));
Q_MX02 U1156 ( .S(n721), .A0(cputx_frame[33]), .A1(r_reg_send[33]), .Z(n912));
Q_MX02 U1157 ( .S(n721), .A0(n913), .A1(n915), .Z(reg_send[32]));
Q_OA21 U1158 ( .A0(n914), .A1(cputx_frame[32]), .B0(n720), .Z(n913));
Q_INV U1159 ( .A(n719), .Z(n914));
Q_MX02 U1160 ( .S(n719), .A0(n916), .A1(n917), .Z(n915));
Q_INV U1161 ( .A(n720), .Z(n916));
Q_MX02 U1162 ( .S(n720), .A0(bimc_eccpar_debug_memaddr[0]), .A1(r_reg_send[32]), .Z(n917));
Q_AN03 U1163 ( .A0(n720), .A1(n918), .A2(n719), .Z(reg_send[31]));
Q_MX02 U1164 ( .S(n721), .A0(cputx_frame[31]), .A1(r_reg_send[31]), .Z(n918));
Q_AN03 U1165 ( .A0(n720), .A1(n919), .A2(n719), .Z(reg_send[30]));
Q_MX02 U1166 ( .S(n721), .A0(cputx_frame[30]), .A1(r_reg_send[30]), .Z(n919));
Q_AN03 U1167 ( .A0(n720), .A1(n920), .A2(n719), .Z(reg_send[29]));
Q_MX02 U1168 ( .S(n721), .A0(cputx_frame[29]), .A1(r_reg_send[29]), .Z(n920));
Q_AN03 U1169 ( .A0(n720), .A1(n921), .A2(n719), .Z(reg_send[28]));
Q_MX02 U1170 ( .S(n721), .A0(cputx_frame[28]), .A1(r_reg_send[28]), .Z(n921));
Q_AN02 U1171 ( .A0(n719), .A1(n922), .Z(reg_send[27]));
Q_MX02 U1172 ( .S(n720), .A0(bimc_eccpar_debug_jabber_off[3]), .A1(n923), .Z(n922));
Q_MX02 U1173 ( .S(n721), .A0(cputx_frame[27]), .A1(r_reg_send[27]), .Z(n923));
Q_AN02 U1174 ( .A0(n719), .A1(n924), .Z(reg_send[26]));
Q_MX02 U1175 ( .S(n720), .A0(bimc_eccpar_debug_jabber_off[2]), .A1(n925), .Z(n924));
Q_MX02 U1176 ( .S(n721), .A0(cputx_frame[26]), .A1(r_reg_send[26]), .Z(n925));
Q_AN02 U1177 ( .A0(n719), .A1(n926), .Z(reg_send[25]));
Q_MX02 U1178 ( .S(n720), .A0(bimc_eccpar_debug_jabber_off[1]), .A1(n927), .Z(n926));
Q_MX02 U1179 ( .S(n721), .A0(cputx_frame[25]), .A1(r_reg_send[25]), .Z(n927));
Q_AN02 U1180 ( .A0(n719), .A1(n928), .Z(reg_send[24]));
Q_MX02 U1181 ( .S(n720), .A0(bimc_eccpar_debug_jabber_off[0]), .A1(n929), .Z(n928));
Q_MX02 U1182 ( .S(n721), .A0(cputx_frame[24]), .A1(r_reg_send[24]), .Z(n929));
Q_AN03 U1183 ( .A0(n720), .A1(n930), .A2(n719), .Z(reg_send[23]));
Q_MX02 U1184 ( .S(n721), .A0(cputx_frame[23]), .A1(r_reg_send[23]), .Z(n930));
Q_AN03 U1185 ( .A0(n720), .A1(n931), .A2(n719), .Z(reg_send[22]));
Q_MX02 U1186 ( .S(n721), .A0(cputx_frame[22]), .A1(r_reg_send[22]), .Z(n931));
Q_AN03 U1187 ( .A0(n720), .A1(n932), .A2(n719), .Z(reg_send[21]));
Q_MX02 U1188 ( .S(n721), .A0(cputx_frame[21]), .A1(r_reg_send[21]), .Z(n932));
Q_AN03 U1189 ( .A0(n720), .A1(n933), .A2(n719), .Z(reg_send[20]));
Q_MX02 U1190 ( .S(n721), .A0(cputx_frame[20]), .A1(r_reg_send[20]), .Z(n933));
Q_AN03 U1191 ( .A0(n720), .A1(n934), .A2(n719), .Z(reg_send[19]));
Q_MX02 U1192 ( .S(n721), .A0(cputx_frame[19]), .A1(r_reg_send[19]), .Z(n934));
Q_AN03 U1193 ( .A0(n720), .A1(n935), .A2(n719), .Z(reg_send[18]));
Q_MX02 U1194 ( .S(n721), .A0(cputx_frame[18]), .A1(r_reg_send[18]), .Z(n935));
Q_AN03 U1195 ( .A0(n720), .A1(n936), .A2(n719), .Z(reg_send[17]));
Q_MX02 U1196 ( .S(n721), .A0(cputx_frame[17]), .A1(r_reg_send[17]), .Z(n936));
Q_AN03 U1197 ( .A0(n720), .A1(n937), .A2(n719), .Z(reg_send[16]));
Q_MX02 U1198 ( .S(n721), .A0(cputx_frame[16]), .A1(r_reg_send[16]), .Z(n937));
Q_AN03 U1199 ( .A0(n720), .A1(n938), .A2(n719), .Z(reg_send[15]));
Q_MX02 U1200 ( .S(n721), .A0(cputx_frame[15]), .A1(r_reg_send[15]), .Z(n938));
Q_AN03 U1201 ( .A0(n720), .A1(n939), .A2(n719), .Z(reg_send[14]));
Q_MX02 U1202 ( .S(n721), .A0(cputx_frame[14]), .A1(r_reg_send[14]), .Z(n939));
Q_AN03 U1203 ( .A0(n720), .A1(n940), .A2(n719), .Z(reg_send[13]));
Q_MX02 U1204 ( .S(n721), .A0(cputx_frame[13]), .A1(r_reg_send[13]), .Z(n940));
Q_AN03 U1205 ( .A0(n720), .A1(n941), .A2(n719), .Z(reg_send[12]));
Q_MX02 U1206 ( .S(n721), .A0(cputx_frame[12]), .A1(r_reg_send[12]), .Z(n941));
Q_AN03 U1207 ( .A0(n720), .A1(n942), .A2(n719), .Z(reg_send[11]));
Q_MX02 U1208 ( .S(n721), .A0(cputx_frame[11]), .A1(r_reg_send[11]), .Z(n942));
Q_AN03 U1209 ( .A0(n720), .A1(n943), .A2(n719), .Z(reg_send[10]));
Q_MX02 U1210 ( .S(n721), .A0(cputx_frame[10]), .A1(r_reg_send[10]), .Z(n943));
Q_AN03 U1211 ( .A0(n720), .A1(n944), .A2(n719), .Z(reg_send[9]));
Q_MX02 U1212 ( .S(n721), .A0(cputx_frame[9]), .A1(r_reg_send[9]), .Z(n944));
Q_AN03 U1213 ( .A0(n720), .A1(n945), .A2(n719), .Z(reg_send[8]));
Q_MX02 U1214 ( .S(n721), .A0(cputx_frame[8]), .A1(r_reg_send[8]), .Z(n945));
Q_AN03 U1215 ( .A0(n720), .A1(n946), .A2(n719), .Z(reg_send[7]));
Q_MX02 U1216 ( .S(n721), .A0(cputx_frame[7]), .A1(r_reg_send[7]), .Z(n946));
Q_AN03 U1217 ( .A0(n720), .A1(n947), .A2(n719), .Z(reg_send[6]));
Q_MX02 U1218 ( .S(n721), .A0(cputx_frame[6]), .A1(r_reg_send[6]), .Z(n947));
Q_AN03 U1219 ( .A0(n720), .A1(n948), .A2(n719), .Z(reg_send[5]));
Q_MX02 U1220 ( .S(n721), .A0(cputx_frame[5]), .A1(r_reg_send[5]), .Z(n948));
Q_AN03 U1221 ( .A0(n720), .A1(n949), .A2(n719), .Z(reg_send[4]));
Q_MX02 U1222 ( .S(n721), .A0(cputx_frame[4]), .A1(r_reg_send[4]), .Z(n949));
Q_AN02 U1223 ( .A0(n719), .A1(n950), .Z(reg_send[3]));
Q_MX02 U1224 ( .S(n720), .A0(bimc_eccpar_debug_eccpar_corrupt[1]), .A1(n951), .Z(n950));
Q_MX02 U1225 ( .S(n721), .A0(cputx_frame[3]), .A1(r_reg_send[3]), .Z(n951));
Q_AN02 U1226 ( .A0(n719), .A1(n952), .Z(reg_send[2]));
Q_MX02 U1227 ( .S(n720), .A0(bimc_eccpar_debug_eccpar_corrupt[0]), .A1(n953), .Z(n952));
Q_MX02 U1228 ( .S(n721), .A0(cputx_frame[2]), .A1(r_reg_send[2]), .Z(n953));
Q_AN02 U1229 ( .A0(n719), .A1(n954), .Z(reg_send[1]));
Q_MX02 U1230 ( .S(n720), .A0(bimc_eccpar_debug_eccpar_disable[1]), .A1(n955), .Z(n954));
Q_MX02 U1231 ( .S(n721), .A0(cputx_frame[1]), .A1(r_reg_send[1]), .Z(n955));
Q_MX02 U1232 ( .S(n719), .A0(n956), .A1(n957), .Z(reg_send[0]));
Q_INV U1233 ( .A(n721), .Z(n956));
Q_MX02 U1234 ( .S(n720), .A0(bimc_eccpar_debug_eccpar_disable[0]), .A1(n958), .Z(n957));
Q_MX02 U1235 ( .S(n721), .A0(cputx_frame[0]), .A1(r_reg_send[0]), .Z(n958));
Q_AO21 U1236 ( .A0(bimc_eccpar_debug_memtype[0]), .A1(n959), .B0(tstate[1]), .Z(n789));
Q_AN03 U1237 ( .A0(bimc_eccpar_debug_memtype[3]), .A1(bimc_eccpar_debug_memtype[2]), .A2(bimc_eccpar_debug_memtype[1]), .Z(n959));
Q_ND03 U1238 ( .A0(rx_frm), .A1(new_frame), .A2(n1257), .Z(n970));
Q_OR02 U1239 ( .A0(n7), .A1(n970), .Z(n963));
Q_OR02 U1240 ( .A0(rx_op[5]), .A1(rx_op[6]), .Z(n964));
Q_OR02 U1241 ( .A0(rx_op[7]), .A1(n1137), .Z(n965));
Q_OR03 U1242 ( .A0(n965), .A1(n964), .A2(n1135), .Z(n986));
Q_OR02 U1243 ( .A0(n1057), .A1(n986), .Z(n987));
Q_OR02 U1244 ( .A0(n1261), .A1(n987), .Z(n966));
Q_XNR2 U1245 ( .A0(rx_chk[0]), .A1(rx_chk[1]), .Z(n977));
Q_NR02 U1246 ( .A0(n4), .A1(n977), .Z(n967));
Q_OR02 U1247 ( .A0(rstate[0]), .A1(n967), .Z(n973));
Q_INV U1248 ( .A(n973), .Z(n968));
Q_MX02 U1249 ( .S(rstate[1]), .A0(n968), .A1(n966), .Z(n969));
Q_MX03 U1250 ( .S0(rstate[2]), .S1(rstate[3]), .A0(n970), .A1(n969), .A2(n981), .Z(n960));
Q_INV U1251 ( .A(n977), .Z(new_frame));
Q_NR02 U1252 ( .A0(rstate[0]), .A1(new_frame), .Z(n971));
Q_OR02 U1253 ( .A0(n981), .A1(n971), .Z(n972));
Q_OR02 U1254 ( .A0(rstate[1]), .A1(n973), .Z(n974));
Q_MX02 U1255 ( .S(rstate[0]), .A0(n979), .A1(n986), .Z(n975));
Q_OR02 U1256 ( .A0(n1289), .A1(n975), .Z(n976));
Q_MX03 U1257 ( .S0(rstate[2]), .S1(rstate[3]), .A0(n976), .A1(n974), .A2(n972), .Z(n961));
Q_ND02 U1258 ( .A0(rx_frm), .A1(rx_resp), .Z(n978));
Q_OR02 U1259 ( .A0(n978), .A1(n977), .Z(n979));
Q_OR02 U1260 ( .A0(rstate[0]), .A1(n979), .Z(n980));
Q_INV U1261 ( .A(n980), .Z(n983));
Q_OR02 U1262 ( .A0(rstate[2]), .A1(rstate[1]), .Z(n981));
Q_OR02 U1263 ( .A0(n981), .A1(n983), .Z(n982));
Q_NR02 U1264 ( .A0(n980), .A1(rstate[1]), .Z(n984));
Q_OR02 U1265 ( .A0(n1284), .A1(n984), .Z(n985));
Q_NR03 U1266 ( .A0(n977), .A1(n3), .A2(n1154), .Z(n988));
Q_MX02 U1267 ( .S(rstate[0]), .A0(n988), .A1(n986), .Z(n989));
Q_AO21 U1268 ( .A0(n989), .A1(rstate[1]), .B0(n1299), .Z(n990));
Q_MX02 U1269 ( .S(rstate[2]), .A0(n990), .A1(n985), .Z(n991));
Q_INV U1270 ( .A(n991), .Z(n992));
Q_MX02 U1271 ( .S(rstate[3]), .A0(n992), .A1(n982), .Z(n962));
Q_INV U1272 ( .A(n961), .Z(n1003));
Q_OR02 U1273 ( .A0(n962), .A1(n960), .Z(n1002));
Q_INV U1274 ( .A(n998), .Z(n993));
Q_AN02 U1275 ( .A0(n1001), .A1(n993), .Z(n994));
Q_XOR2 U1276 ( .A0(n963), .A1(n994), .Z(nxt_rstate[3]));
Q_INV U1277 ( .A(n1004), .Z(n995));
Q_INV U1278 ( .A(n962), .Z(n996));
Q_OR02 U1279 ( .A0(n996), .A1(n960), .Z(n997));
Q_AO21 U1280 ( .A0(n997), .A1(n961), .B0(n998), .Z(n999));
Q_NR02 U1281 ( .A0(n960), .A1(n961), .Z(n998));
Q_MX02 U1282 ( .S(n963), .A0(n995), .A1(n999), .Z(n1000));
Q_INV U1283 ( .A(n1000), .Z(nxt_rstate[2]));
Q_OR02 U1284 ( .A0(n1003), .A1(n1002), .Z(n1001));
Q_AO21 U1285 ( .A0(n962), .A1(n961), .B0(n1004), .Z(n1005));
Q_NR02 U1286 ( .A0(n1002), .A1(n961), .Z(n1004));
Q_MX02 U1287 ( .S(n963), .A0(n1001), .A1(n1005), .Z(nxt_rstate[1]));
Q_XNR2 U1288 ( .A0(n962), .A1(n960), .Z(n1006));
Q_OR02 U1289 ( .A0(n961), .A1(n1006), .Z(n1007));
Q_ND02 U1290 ( .A0(n963), .A1(n1007), .Z(nxt_rstate[0]));
Q_OR02 U1291 ( .A0(n1013), .A1(n1008), .Z(n1014));
Q_OR02 U1292 ( .A0(rx_op[4]), .A1(rx_op[2]), .Z(n1036));
Q_OR03 U1293 ( .A0(rx_op[6]), .A1(rx_op[7]), .A2(n1036), .Z(n1037));
Q_OR03 U1294 ( .A0(rx_op[3]), .A1(rx_op[5]), .A2(n1037), .Z(n1053));
Q_OR03 U1295 ( .A0(rx_op[1]), .A1(rx_op[0]), .A2(n1053), .Z(n1048));
Q_INV U1296 ( .A(n1048), .Z(n1038));
Q_OR02 U1297 ( .A0(rstate[2]), .A1(n1038), .Z(n1044));
Q_OR03 U1298 ( .A0(rstate[1]), .A1(rstate[3]), .A2(n1044), .Z(n1040));
Q_NR03 U1299 ( .A0(bimc_dbgcmd2_rxflag_din), .A1(n1261), .A2(n1040), .Z(n1039));
Q_NR02 U1300 ( .A0(rstate[0]), .A1(n1040), .Z(n1041));
Q_OR02 U1301 ( .A0(o_bimc_dbgcmd2[9]), .A1(n1041), .Z(n1015));
Q_OR02 U1302 ( .A0(bimc_rxcmd2_rxflag_din), .A1(rstate[2]), .Z(n1042));
Q_NR03 U1303 ( .A0(n1061), .A1(n1042), .A2(n1261), .Z(n1043));
Q_AO21 U1304 ( .A0(n1278), .A1(n1256), .B0(o_bimc_rxcmd2[9]), .Z(n1016));
Q_OR02 U1305 ( .A0(n1253), .A1(n1044), .Z(n1046));
Q_NR03 U1306 ( .A0(bimc_pollrsp2_rxflag_din), .A1(n1298), .A2(n1046), .Z(n1045));
Q_NR02 U1307 ( .A0(n1308), .A1(n1046), .Z(n1047));
Q_OR02 U1308 ( .A0(o_bimc_pollrsp2[9]), .A1(n1047), .Z(n1017));
Q_ND02 U1309 ( .A0(rstate[2]), .A1(n1048), .Z(n1049));
Q_OR02 U1310 ( .A0(rstate[3]), .A1(n1049), .Z(n1051));
Q_NR03 U1311 ( .A0(bimc_rxrsp2_rxflag_din), .A1(n1298), .A2(n1051), .Z(n1050));
Q_NR02 U1312 ( .A0(n1308), .A1(n1051), .Z(n1052));
Q_OR02 U1313 ( .A0(o_bimc_rxrsp2[9]), .A1(n1052), .Z(n1018));
Q_OR02 U1314 ( .A0(n1137), .A1(n1053), .Z(n1056));
Q_OR02 U1315 ( .A0(rx_op[1]), .A1(n1056), .Z(n1059));
Q_ND02 U1316 ( .A0(n1299), .A1(n1288), .Z(n1054));
Q_NR02 U1317 ( .A0(n1054), .A1(n1059), .Z(n1055));
Q_OR02 U1318 ( .A0(o_bimc_monitor_mask[6]), .A1(n1055), .Z(n1020));
Q_OR02 U1319 ( .A0(n1057), .A1(n1056), .Z(n1058));
Q_MX02 U1320 ( .S(rstate[2]), .A0(n1059), .A1(n1058), .Z(n1060));
Q_INV U1321 ( .A(n1060), .Z(n1062));
Q_OR02 U1322 ( .A0(n1289), .A1(rstate[3]), .Z(n1061));
Q_NR03 U1323 ( .A0(n1261), .A1(n1061), .A2(n1062), .Z(n1063));
Q_OR02 U1324 ( .A0(o_bimc_monitor_mask[5]), .A1(n1063), .Z(n1021));
Q_OR02 U1325 ( .A0(n1012), .A1(o_bimc_monitor_mask[4]), .Z(n1022));
Q_OR02 U1326 ( .A0(n1010), .A1(o_bimc_monitor_mask[2]), .Z(n1023));
Q_OR02 U1327 ( .A0(n1011), .A1(o_bimc_monitor_mask[1]), .Z(n1024));
Q_OR02 U1328 ( .A0(n1009), .A1(o_bimc_monitor_mask[0]), .Z(n1025));
Q_INV U1329 ( .A(o_bimc_monitor_mask[0]), .Z(n1026));
Q_INV U1330 ( .A(o_bimc_monitor_mask[1]), .Z(n1027));
Q_INV U1331 ( .A(o_bimc_monitor_mask[2]), .Z(n1028));
Q_INV U1332 ( .A(o_bimc_monitor_mask[4]), .Z(n1029));
Q_INV U1333 ( .A(o_bimc_monitor_mask[5]), .Z(n1030));
Q_INV U1334 ( .A(o_bimc_monitor_mask[6]), .Z(n1031));
Q_INV U1335 ( .A(o_bimc_rxrsp2[9]), .Z(n1032));
Q_INV U1336 ( .A(o_bimc_pollrsp2[9]), .Z(n1033));
Q_INV U1337 ( .A(o_bimc_rxcmd2[9]), .Z(n1034));
Q_INV U1338 ( .A(o_bimc_dbgcmd2[9]), .Z(n1035));
Q_FDP1 \rx_chk_REG[0] ( .CK(clk), .R(rst_n), .D(rcv_chk), .Q(rx_chk[0]), .QN( ));
Q_FDP1 \rx_chk_REG[1] ( .CK(clk), .R(rst_n), .D(rx_chk[0]), .Q(rx_chk[1]), .QN( ));
Q_FDP1 bimc_parity_error_cnt_parity_errors_en_REG  ( .CK(clk), .R(rst_n), .D(n1010), .Q(bimc_parity_error_cnt_parity_errors_en), .QN( ));
Q_FDP1 bimc_ecc_correctable_error_cnt_correctable_ecc_en_REG  ( .CK(clk), .R(rst_n), .D(n1011), .Q(bimc_ecc_correctable_error_cnt_correctable_ecc_en), .QN( ));
Q_FDP1 bimc_ecc_uncorrectable_error_cnt_uncorrectable_ecc_en_REG  ( .CK(clk), .R(rst_n), .D(n1009), .Q(bimc_ecc_uncorrectable_error_cnt_uncorrectable_ecc_en), .QN( ));
Q_XNR2 U1344 ( .A0(rx_dat[11]), .A1(n1065), .Z(n1064));
Q_OR02 U1345 ( .A0(rx_dat[10]), .A1(n1067), .Z(n1065));
Q_XNR2 U1346 ( .A0(rx_dat[10]), .A1(n1067), .Z(n1066));
Q_OR02 U1347 ( .A0(rx_dat[9]), .A1(n1069), .Z(n1067));
Q_XNR2 U1348 ( .A0(rx_dat[9]), .A1(n1069), .Z(n1068));
Q_OR02 U1349 ( .A0(rx_dat[8]), .A1(n1071), .Z(n1069));
Q_XNR2 U1350 ( .A0(rx_dat[8]), .A1(n1071), .Z(n1070));
Q_OR02 U1351 ( .A0(rx_dat[7]), .A1(n1073), .Z(n1071));
Q_XNR2 U1352 ( .A0(rx_dat[7]), .A1(n1073), .Z(n1072));
Q_OR02 U1353 ( .A0(rx_dat[6]), .A1(n1075), .Z(n1073));
Q_XNR2 U1354 ( .A0(rx_dat[6]), .A1(n1075), .Z(n1074));
Q_OR02 U1355 ( .A0(rx_dat[5]), .A1(n1077), .Z(n1075));
Q_XNR2 U1356 ( .A0(rx_dat[5]), .A1(n1077), .Z(n1076));
Q_OR02 U1357 ( .A0(rx_dat[4]), .A1(n1079), .Z(n1077));
Q_XNR2 U1358 ( .A0(rx_dat[4]), .A1(n1079), .Z(n1078));
Q_OR02 U1359 ( .A0(rx_dat[3]), .A1(n1081), .Z(n1079));
Q_XNR2 U1360 ( .A0(rx_dat[3]), .A1(n1081), .Z(n1080));
Q_OR02 U1361 ( .A0(rx_dat[2]), .A1(n1083), .Z(n1081));
Q_XNR2 U1362 ( .A0(rx_dat[2]), .A1(n1083), .Z(n1082));
Q_OR02 U1363 ( .A0(rx_dat[1]), .A1(rx_dat[0]), .Z(n1083));
Q_XNR2 U1364 ( .A0(rx_dat[1]), .A1(rx_dat[0]), .Z(n1084));
Q_NR03 U1365 ( .A0(n1087), .A1(n1086), .A2(n1166), .Z(n1019));
Q_OR03 U1366 ( .A0(n1090), .A1(n1089), .A2(n1088), .Z(n1086));
Q_OR03 U1367 ( .A0(n1093), .A1(n1092), .A2(n1091), .Z(n1087));
Q_OR03 U1368 ( .A0(n1146), .A1(n1095), .A2(n1094), .Z(n1088));
Q_OR03 U1369 ( .A0(n1098), .A1(n1097), .A2(n1096), .Z(n1089));
Q_OR03 U1370 ( .A0(n1101), .A1(n1100), .A2(n1099), .Z(n1090));
Q_OR03 U1371 ( .A0(n1161), .A1(n1103), .A2(n1102), .Z(n1091));
Q_OR03 U1372 ( .A0(rx_addr[3]), .A1(rx_addr[2]), .A2(rx_addr[1]), .Z(n1092));
Q_OR03 U1373 ( .A0(rx_addr[6]), .A1(rx_addr[5]), .A2(rx_addr[4]), .Z(n1093));
Q_OR03 U1374 ( .A0(rx_addr[9]), .A1(rx_addr[8]), .A2(rx_addr[7]), .Z(n1094));
Q_OR03 U1375 ( .A0(rx_addr[12]), .A1(rx_addr[11]), .A2(rx_addr[10]), .Z(n1095));
Q_ND03 U1376 ( .A0(rx_mem[2]), .A1(rx_mem[1]), .A2(rx_mem[0]), .Z(n1096));
Q_ND03 U1377 ( .A0(rx_mem[5]), .A1(rx_mem[4]), .A2(rx_mem[3]), .Z(n1097));
Q_ND03 U1378 ( .A0(rx_mem[8]), .A1(rx_mem[7]), .A2(rx_mem[6]), .Z(n1098));
Q_ND03 U1379 ( .A0(rx_mem[11]), .A1(rx_mem[10]), .A2(rx_mem[9]), .Z(n1099));
Q_OR03 U1380 ( .A0(rx_op[2]), .A1(n1057), .A2(rx_op[0]), .Z(n1100));
Q_OR03 U1381 ( .A0(rx_op[5]), .A1(rx_op[4]), .A2(rx_op[3]), .Z(n1101));
Q_OR03 U1382 ( .A0(n1104), .A1(rx_op[7]), .A2(rx_op[6]), .Z(n1102));
Q_ND03 U1383 ( .A0(rx_type[3]), .A1(rx_type[2]), .A2(rx_type[1]), .Z(n1103));
Q_AN03 U1384 ( .A0(n1132), .A1(n1121), .A2(n1105), .Z(n1010));
Q_OR02 U1385 ( .A0(n1107), .A1(n1106), .Z(n1105));
Q_OR03 U1386 ( .A0(n1110), .A1(n1109), .A2(n1108), .Z(n1106));
Q_OR03 U1387 ( .A0(n1113), .A1(n1112), .A2(n1111), .Z(n1107));
Q_OR03 U1388 ( .A0(n1116), .A1(n1115), .A2(n1114), .Z(n1108));
Q_OR03 U1389 ( .A0(n1119), .A1(n1118), .A2(n1117), .Z(n1109));
Q_OR03 U1390 ( .A0(rx_dat[1]), .A1(rx_dat[0]), .A2(n1120), .Z(n1110));
Q_OR03 U1391 ( .A0(rx_dat[4]), .A1(rx_dat[3]), .A2(rx_dat[2]), .Z(n1111));
Q_OR03 U1392 ( .A0(rx_dat[7]), .A1(rx_dat[6]), .A2(rx_dat[5]), .Z(n1112));
Q_OR03 U1393 ( .A0(rx_dat[10]), .A1(rx_dat[9]), .A2(rx_dat[8]), .Z(n1113));
Q_OR03 U1394 ( .A0(rx_dat[13]), .A1(rx_dat[12]), .A2(rx_dat[11]), .Z(n1114));
Q_OR03 U1395 ( .A0(rx_dat[16]), .A1(rx_dat[15]), .A2(rx_dat[14]), .Z(n1115));
Q_OR03 U1396 ( .A0(rx_dat[19]), .A1(rx_dat[18]), .A2(rx_dat[17]), .Z(n1116));
Q_OR03 U1397 ( .A0(rx_dat[22]), .A1(rx_dat[21]), .A2(rx_dat[20]), .Z(n1117));
Q_OR03 U1398 ( .A0(rx_dat[25]), .A1(rx_dat[24]), .A2(rx_dat[23]), .Z(n1118));
Q_OR03 U1399 ( .A0(rx_dat[28]), .A1(rx_dat[27]), .A2(rx_dat[26]), .Z(n1119));
Q_OR03 U1400 ( .A0(rx_dat[31]), .A1(rx_dat[30]), .A2(rx_dat[29]), .Z(n1120));
Q_NR02 U1401 ( .A0(n1123), .A1(n1122), .Z(n1121));
Q_OR03 U1402 ( .A0(n1126), .A1(n1125), .A2(n1124), .Z(n1122));
Q_OR03 U1403 ( .A0(rx_addr[0]), .A1(n1146), .A2(n1127), .Z(n1123));
Q_OR03 U1404 ( .A0(rx_addr[3]), .A1(n1153), .A2(rx_addr[1]), .Z(n1124));
Q_OR03 U1405 ( .A0(rx_addr[6]), .A1(n1129), .A2(rx_addr[4]), .Z(n1125));
Q_OR03 U1406 ( .A0(rx_addr[9]), .A1(n1128), .A2(n1150), .Z(n1126));
Q_OR03 U1407 ( .A0(rx_addr[12]), .A1(n1147), .A2(rx_addr[10]), .Z(n1127));
Q_AN03 U1408 ( .A0(n1132), .A1(n1139), .A2(n1130), .Z(n1009));
Q_AN02 U1409 ( .A0(rx_dat[2]), .A1(rx_dat[0]), .Z(n1130));
Q_AN03 U1410 ( .A0(n1132), .A1(n1139), .A2(n1131), .Z(n1011));
Q_AN02 U1411 ( .A0(rx_dat[0]), .A1(rx_dat[1]), .Z(n1131));
Q_NR02 U1412 ( .A0(n1135), .A1(n1134), .Z(n1133));
Q_OR03 U1413 ( .A0(n1057), .A1(n1137), .A2(n1136), .Z(n1134));
Q_OR03 U1414 ( .A0(rx_op[4]), .A1(rx_op[3]), .A2(rx_op[2]), .Z(n1135));
Q_OR03 U1415 ( .A0(rx_op[7]), .A1(rx_op[6]), .A2(rx_op[5]), .Z(n1136));
Q_AN03 U1416 ( .A0(rstate[0]), .A1(n1138), .A2(n1133), .Z(n1132));
Q_AN03 U1417 ( .A0(rstate[3]), .A1(n1260), .A2(n1289), .Z(n1138));
Q_NR02 U1418 ( .A0(n1141), .A1(n1140), .Z(n1139));
Q_OR03 U1419 ( .A0(n1144), .A1(n1143), .A2(n1142), .Z(n1140));
Q_OR03 U1420 ( .A0(rx_addr[0]), .A1(n1146), .A2(n1145), .Z(n1141));
Q_OR03 U1421 ( .A0(n1152), .A1(n1153), .A2(rx_addr[1]), .Z(n1142));
Q_OR03 U1422 ( .A0(n1151), .A1(rx_addr[5]), .A2(rx_addr[4]), .Z(n1143));
Q_OR03 U1423 ( .A0(n1149), .A1(rx_addr[8]), .A2(n1150), .Z(n1144));
Q_OR03 U1424 ( .A0(rx_addr[12]), .A1(n1147), .A2(n1148), .Z(n1145));
Q_OR03 U1425 ( .A0(rx_addr[15]), .A1(rx_addr[14]), .A2(rx_addr[13]), .Z(n1146));
Q_NR03 U1426 ( .A0(n1157), .A1(rx_frm), .A2(n977), .Z(n1012));
Q_XOR2 U1427 ( .A0(rstate[2]), .A1(n1253), .Z(n1155));
Q_MX02 U1428 ( .S(rstate[1]), .A0(n1155), .A1(n7), .Z(n1156));
Q_OR02 U1429 ( .A0(rstate[0]), .A1(n1156), .Z(n1157));
Q_NR03 U1430 ( .A0(n1166), .A1(n1162), .A2(n1158), .Z(n1013));
Q_OR02 U1431 ( .A0(n1160), .A1(n1159), .Z(n1158));
Q_OR03 U1432 ( .A0(n1094), .A1(n1093), .A2(n1092), .Z(n1159));
Q_OR03 U1433 ( .A0(n1161), .A1(n1146), .A2(n1095), .Z(n1160));
Q_OR02 U1434 ( .A0(n1135), .A1(n1163), .Z(n1162));
Q_OR03 U1435 ( .A0(n1057), .A1(rx_op[0]), .A2(n1136), .Z(n1163));
Q_INV U1436 ( .A(n1164), .Z(n1008));
Q_OR02 U1437 ( .A0(tstate[0]), .A1(n1165), .Z(n1164));
Q_OR03 U1438 ( .A0(tstate[3]), .A1(tstate[2]), .A2(tstate[1]), .Z(n1165));
Q_OR02 U1439 ( .A0(n1261), .A1(n1167), .Z(n1166));
Q_OR03 U1440 ( .A0(rstate[3]), .A1(rstate[2]), .A2(rstate[1]), .Z(n1167));
Q_FDP1 \rstate_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_rstate[0]), .Q(rstate[0]), .QN(n1261));
Q_FDP2 \rstate_REG[1] ( .CK(clk), .S(rst_n), .D(nxt_rstate[1]), .Q(rstate[1]), .QN(n1289));
Q_FDP1 \rstate_REG[2] ( .CK(clk), .R(rst_n), .D(nxt_rstate[2]), .Q(rstate[2]), .QN(n1260));
Q_FDP1 \rstate_REG[3] ( .CK(clk), .R(rst_n), .D(nxt_rstate[3]), .Q(rstate[3]), .QN(n1253));
Q_FDP1 rx_frm_REG  ( .CK(clk), .R(rst_n), .D(rcv_frm), .Q(rx_frm), .QN(n1154));
Q_FDP1 rx_resp_REG  ( .CK(clk), .R(rst_n), .D(rcv_resp), .Q(rx_resp), .QN( ));
Q_FDP1 \rx_dat_REG[0] ( .CK(clk), .R(rst_n), .D(rcv_dat[0]), .Q(rx_dat[0]), .QN(n1085));
Q_FDP1 \rx_dat_REG[1] ( .CK(clk), .R(rst_n), .D(rcv_dat[1]), .Q(rx_dat[1]), .QN( ));
Q_FDP1 \rx_dat_REG[2] ( .CK(clk), .R(rst_n), .D(rcv_dat[2]), .Q(rx_dat[2]), .QN( ));
Q_FDP1 \rx_dat_REG[3] ( .CK(clk), .R(rst_n), .D(rcv_dat[3]), .Q(rx_dat[3]), .QN( ));
Q_FDP1 \rx_dat_REG[4] ( .CK(clk), .R(rst_n), .D(rcv_dat[4]), .Q(rx_dat[4]), .QN( ));
Q_FDP1 \rx_dat_REG[5] ( .CK(clk), .R(rst_n), .D(rcv_dat[5]), .Q(rx_dat[5]), .QN( ));
Q_FDP1 \rx_dat_REG[6] ( .CK(clk), .R(rst_n), .D(rcv_dat[6]), .Q(rx_dat[6]), .QN( ));
Q_FDP1 \rx_dat_REG[7] ( .CK(clk), .R(rst_n), .D(rcv_dat[7]), .Q(rx_dat[7]), .QN( ));
Q_FDP1 \rx_dat_REG[8] ( .CK(clk), .R(rst_n), .D(rcv_dat[8]), .Q(rx_dat[8]), .QN( ));
Q_FDP1 \rx_dat_REG[9] ( .CK(clk), .R(rst_n), .D(rcv_dat[9]), .Q(rx_dat[9]), .QN( ));
Q_FDP1 \rx_dat_REG[10] ( .CK(clk), .R(rst_n), .D(rcv_dat[10]), .Q(rx_dat[10]), .QN( ));
Q_FDP1 \rx_dat_REG[11] ( .CK(clk), .R(rst_n), .D(rcv_dat[11]), .Q(rx_dat[11]), .QN( ));
Q_FDP1 \rx_dat_REG[12] ( .CK(clk), .R(rst_n), .D(rcv_dat[12]), .Q(rx_dat[12]), .QN( ));
Q_FDP1 \rx_dat_REG[13] ( .CK(clk), .R(rst_n), .D(rcv_dat[13]), .Q(rx_dat[13]), .QN( ));
Q_FDP1 \rx_dat_REG[14] ( .CK(clk), .R(rst_n), .D(rcv_dat[14]), .Q(rx_dat[14]), .QN( ));
Q_FDP1 \rx_dat_REG[15] ( .CK(clk), .R(rst_n), .D(rcv_dat[15]), .Q(rx_dat[15]), .QN( ));
Q_FDP1 \rx_dat_REG[16] ( .CK(clk), .R(rst_n), .D(rcv_dat[16]), .Q(rx_dat[16]), .QN( ));
Q_FDP1 \rx_dat_REG[17] ( .CK(clk), .R(rst_n), .D(rcv_dat[17]), .Q(rx_dat[17]), .QN( ));
Q_FDP1 \rx_dat_REG[18] ( .CK(clk), .R(rst_n), .D(rcv_dat[18]), .Q(rx_dat[18]), .QN( ));
Q_FDP1 \rx_dat_REG[19] ( .CK(clk), .R(rst_n), .D(rcv_dat[19]), .Q(rx_dat[19]), .QN( ));
Q_FDP1 \rx_dat_REG[20] ( .CK(clk), .R(rst_n), .D(rcv_dat[20]), .Q(rx_dat[20]), .QN( ));
Q_FDP1 \rx_dat_REG[21] ( .CK(clk), .R(rst_n), .D(rcv_dat[21]), .Q(rx_dat[21]), .QN( ));
Q_FDP1 \rx_dat_REG[22] ( .CK(clk), .R(rst_n), .D(rcv_dat[22]), .Q(rx_dat[22]), .QN( ));
Q_FDP1 \rx_dat_REG[23] ( .CK(clk), .R(rst_n), .D(rcv_dat[23]), .Q(rx_dat[23]), .QN( ));
Q_FDP1 \rx_dat_REG[24] ( .CK(clk), .R(rst_n), .D(rcv_dat[24]), .Q(rx_dat[24]), .QN( ));
Q_FDP1 \rx_dat_REG[25] ( .CK(clk), .R(rst_n), .D(rcv_dat[25]), .Q(rx_dat[25]), .QN( ));
Q_FDP1 \rx_dat_REG[26] ( .CK(clk), .R(rst_n), .D(rcv_dat[26]), .Q(rx_dat[26]), .QN( ));
Q_FDP1 \rx_dat_REG[27] ( .CK(clk), .R(rst_n), .D(rcv_dat[27]), .Q(rx_dat[27]), .QN( ));
Q_FDP1 \rx_dat_REG[28] ( .CK(clk), .R(rst_n), .D(rcv_dat[28]), .Q(rx_dat[28]), .QN( ));
Q_FDP1 \rx_dat_REG[29] ( .CK(clk), .R(rst_n), .D(rcv_dat[29]), .Q(rx_dat[29]), .QN( ));
Q_FDP1 \rx_dat_REG[30] ( .CK(clk), .R(rst_n), .D(rcv_dat[30]), .Q(rx_dat[30]), .QN( ));
Q_FDP1 \rx_dat_REG[31] ( .CK(clk), .R(rst_n), .D(rcv_dat[31]), .Q(rx_dat[31]), .QN( ));
Q_FDP1 \rx_addr_REG[0] ( .CK(clk), .R(rst_n), .D(rcv_dat[32]), .Q(rx_addr[0]), .QN(n1161));
Q_FDP1 \rx_addr_REG[1] ( .CK(clk), .R(rst_n), .D(rcv_dat[33]), .Q(rx_addr[1]), .QN( ));
Q_FDP1 \rx_addr_REG[2] ( .CK(clk), .R(rst_n), .D(rcv_dat[34]), .Q(rx_addr[2]), .QN(n1153));
Q_FDP1 \rx_addr_REG[3] ( .CK(clk), .R(rst_n), .D(rcv_dat[35]), .Q(rx_addr[3]), .QN(n1152));
Q_FDP1 \rx_addr_REG[4] ( .CK(clk), .R(rst_n), .D(rcv_dat[36]), .Q(rx_addr[4]), .QN( ));
Q_FDP1 \rx_addr_REG[5] ( .CK(clk), .R(rst_n), .D(rcv_dat[37]), .Q(rx_addr[5]), .QN(n1129));
Q_FDP1 \rx_addr_REG[6] ( .CK(clk), .R(rst_n), .D(rcv_dat[38]), .Q(rx_addr[6]), .QN(n1151));
Q_FDP1 \rx_addr_REG[7] ( .CK(clk), .R(rst_n), .D(rcv_dat[39]), .Q(rx_addr[7]), .QN(n1150));
Q_FDP1 \rx_addr_REG[8] ( .CK(clk), .R(rst_n), .D(rcv_dat[40]), .Q(rx_addr[8]), .QN(n1128));
Q_FDP1 \rx_addr_REG[9] ( .CK(clk), .R(rst_n), .D(rcv_dat[41]), .Q(rx_addr[9]), .QN(n1149));
Q_FDP1 \rx_addr_REG[10] ( .CK(clk), .R(rst_n), .D(rcv_dat[42]), .Q(rx_addr[10]), .QN(n1148));
Q_FDP1 \rx_addr_REG[11] ( .CK(clk), .R(rst_n), .D(rcv_dat[43]), .Q(rx_addr[11]), .QN(n1147));
Q_FDP1 \rx_addr_REG[12] ( .CK(clk), .R(rst_n), .D(rcv_dat[44]), .Q(rx_addr[12]), .QN( ));
Q_FDP1 \rx_addr_REG[13] ( .CK(clk), .R(rst_n), .D(rcv_dat[45]), .Q(rx_addr[13]), .QN( ));
Q_FDP1 \rx_addr_REG[14] ( .CK(clk), .R(rst_n), .D(rcv_dat[46]), .Q(rx_addr[14]), .QN( ));
Q_FDP1 \rx_addr_REG[15] ( .CK(clk), .R(rst_n), .D(rcv_dat[47]), .Q(rx_addr[15]), .QN( ));
Q_FDP1 \rx_mem_REG[0] ( .CK(clk), .R(rst_n), .D(rcv_dat[48]), .Q(rx_mem[0]), .QN( ));
Q_FDP1 \rx_mem_REG[1] ( .CK(clk), .R(rst_n), .D(rcv_dat[49]), .Q(rx_mem[1]), .QN( ));
Q_FDP1 \rx_mem_REG[2] ( .CK(clk), .R(rst_n), .D(rcv_dat[50]), .Q(rx_mem[2]), .QN( ));
Q_FDP1 \rx_mem_REG[3] ( .CK(clk), .R(rst_n), .D(rcv_dat[51]), .Q(rx_mem[3]), .QN( ));
Q_FDP1 \rx_mem_REG[4] ( .CK(clk), .R(rst_n), .D(rcv_dat[52]), .Q(rx_mem[4]), .QN( ));
Q_FDP1 \rx_mem_REG[5] ( .CK(clk), .R(rst_n), .D(rcv_dat[53]), .Q(rx_mem[5]), .QN( ));
Q_FDP1 \rx_mem_REG[6] ( .CK(clk), .R(rst_n), .D(rcv_dat[54]), .Q(rx_mem[6]), .QN( ));
Q_FDP1 \rx_mem_REG[7] ( .CK(clk), .R(rst_n), .D(rcv_dat[55]), .Q(rx_mem[7]), .QN( ));
Q_FDP1 \rx_mem_REG[8] ( .CK(clk), .R(rst_n), .D(rcv_dat[56]), .Q(rx_mem[8]), .QN( ));
Q_FDP1 \rx_mem_REG[9] ( .CK(clk), .R(rst_n), .D(rcv_dat[57]), .Q(rx_mem[9]), .QN( ));
Q_FDP1 \rx_mem_REG[10] ( .CK(clk), .R(rst_n), .D(rcv_dat[58]), .Q(rx_mem[10]), .QN( ));
Q_FDP1 \rx_mem_REG[11] ( .CK(clk), .R(rst_n), .D(rcv_dat[59]), .Q(rx_mem[11]), .QN( ));
Q_FDP1 \rx_op_REG[0] ( .CK(clk), .R(rst_n), .D(rcv_dat[60]), .Q(rx_op[0]), .QN(n1137));
Q_FDP1 \rx_op_REG[1] ( .CK(clk), .R(rst_n), .D(rcv_dat[61]), .Q(rx_op[1]), .QN(n1057));
Q_FDP1 \rx_op_REG[2] ( .CK(clk), .R(rst_n), .D(rcv_dat[62]), .Q(rx_op[2]), .QN( ));
Q_FDP1 \rx_op_REG[3] ( .CK(clk), .R(rst_n), .D(rcv_dat[63]), .Q(rx_op[3]), .QN( ));
Q_FDP1 \rx_op_REG[4] ( .CK(clk), .R(rst_n), .D(rcv_dat[64]), .Q(rx_op[4]), .QN( ));
Q_FDP1 \rx_op_REG[5] ( .CK(clk), .R(rst_n), .D(rcv_dat[65]), .Q(rx_op[5]), .QN( ));
Q_FDP1 \rx_op_REG[6] ( .CK(clk), .R(rst_n), .D(rcv_dat[66]), .Q(rx_op[6]), .QN( ));
Q_FDP1 \rx_op_REG[7] ( .CK(clk), .R(rst_n), .D(rcv_dat[67]), .Q(rx_op[7]), .QN( ));
Q_FDP1 \rx_type_REG[0] ( .CK(clk), .R(rst_n), .D(rcv_dat[68]), .Q(rx_type[0]), .QN(n1104));
Q_FDP1 \rx_type_REG[1] ( .CK(clk), .R(rst_n), .D(rcv_dat[69]), .Q(rx_type[1]), .QN( ));
Q_FDP1 \rx_type_REG[2] ( .CK(clk), .R(rst_n), .D(rcv_dat[70]), .Q(rx_type[2]), .QN( ));
Q_FDP1 \rx_type_REG[3] ( .CK(clk), .R(rst_n), .D(rcv_dat[71]), .Q(rx_type[3]), .QN( ));
Q_INV U1519 ( .A(bimc_isync), .Z(n1169));
Q_FDP1 \bm_cnt_REG[0] ( .CK(clk), .R(rst_n), .D(n1176), .Q(bm_cnt[0]), .QN(n1188));
Q_FDP1 \bm_cnt_REG[1] ( .CK(clk), .R(rst_n), .D(n1175), .Q(bm_cnt[1]), .QN( ));
Q_FDP2 \bm_cnt_REG[2] ( .CK(clk), .S(rst_n), .D(n1174), .Q(bm_cnt[2]), .QN( ));
Q_FDP2 \bm_cnt_REG[3] ( .CK(clk), .S(rst_n), .D(n1173), .Q(bm_cnt[3]), .QN(n1193));
Q_FDP2 \bm_cnt_REG[4] ( .CK(clk), .S(rst_n), .D(n1172), .Q(bm_cnt[4]), .QN( ));
Q_FDP2 \bm_cnt_REG[5] ( .CK(clk), .S(rst_n), .D(n1171), .Q(bm_cnt[5]), .QN( ));
Q_FDP2 \bm_cnt_REG[6] ( .CK(clk), .S(rst_n), .D(n1170), .Q(bm_cnt[6]), .QN(n1192));
Q_FDP1 \bimc_rdat_REG[0] ( .CK(clk), .R(rst_n), .D(bimc_idat), .Q(bimc_rdat[0]), .QN( ));
Q_FDP1 \bimc_rdat_REG[1] ( .CK(clk), .R(rst_n), .D(bimc_rdat[0]), .Q(bimc_rdat[1]), .QN( ));
Q_FDP1 \bimc_rdat_REG[2] ( .CK(clk), .R(rst_n), .D(bimc_rdat[1]), .Q(bimc_rdat[2]), .QN( ));
Q_FDP1 \bimc_rdat_REG[3] ( .CK(clk), .R(rst_n), .D(bimc_rdat[2]), .Q(bimc_rdat[3]), .QN( ));
Q_FDP1 \bimc_rdat_REG[4] ( .CK(clk), .R(rst_n), .D(bimc_rdat[3]), .Q(bimc_rdat[4]), .QN( ));
Q_FDP1 \bimc_rdat_REG[5] ( .CK(clk), .R(rst_n), .D(bimc_rdat[4]), .Q(bimc_rdat[5]), .QN( ));
Q_FDP1 \bimc_rdat_REG[6] ( .CK(clk), .R(rst_n), .D(bimc_rdat[5]), .Q(bimc_rdat[6]), .QN( ));
Q_FDP1 \bimc_rdat_REG[7] ( .CK(clk), .R(rst_n), .D(bimc_rdat[6]), .Q(bimc_rdat[7]), .QN( ));
Q_FDP1 \bimc_rdat_REG[8] ( .CK(clk), .R(rst_n), .D(bimc_rdat[7]), .Q(bimc_rdat[8]), .QN( ));
Q_FDP1 \bimc_rdat_REG[9] ( .CK(clk), .R(rst_n), .D(bimc_rdat[8]), .Q(bimc_rdat[9]), .QN( ));
Q_FDP1 \bimc_rdat_REG[10] ( .CK(clk), .R(rst_n), .D(bimc_rdat[9]), .Q(bimc_rdat[10]), .QN( ));
Q_FDP1 \bimc_rdat_REG[11] ( .CK(clk), .R(rst_n), .D(bimc_rdat[10]), .Q(bimc_rdat[11]), .QN( ));
Q_FDP1 \bimc_rdat_REG[12] ( .CK(clk), .R(rst_n), .D(bimc_rdat[11]), .Q(bimc_rdat[12]), .QN( ));
Q_FDP1 \bimc_rdat_REG[13] ( .CK(clk), .R(rst_n), .D(bimc_rdat[12]), .Q(bimc_rdat[13]), .QN( ));
Q_FDP1 \bimc_rdat_REG[14] ( .CK(clk), .R(rst_n), .D(bimc_rdat[13]), .Q(bimc_rdat[14]), .QN( ));
Q_FDP1 \bimc_rdat_REG[15] ( .CK(clk), .R(rst_n), .D(bimc_rdat[14]), .Q(bimc_rdat[15]), .QN( ));
Q_FDP1 \bimc_rdat_REG[16] ( .CK(clk), .R(rst_n), .D(bimc_rdat[15]), .Q(bimc_rdat[16]), .QN( ));
Q_FDP1 \bimc_rdat_REG[17] ( .CK(clk), .R(rst_n), .D(bimc_rdat[16]), .Q(bimc_rdat[17]), .QN( ));
Q_FDP1 \bimc_rdat_REG[18] ( .CK(clk), .R(rst_n), .D(bimc_rdat[17]), .Q(bimc_rdat[18]), .QN( ));
Q_FDP1 \bimc_rdat_REG[19] ( .CK(clk), .R(rst_n), .D(bimc_rdat[18]), .Q(bimc_rdat[19]), .QN( ));
Q_FDP1 \bimc_rdat_REG[20] ( .CK(clk), .R(rst_n), .D(bimc_rdat[19]), .Q(bimc_rdat[20]), .QN( ));
Q_FDP1 \bimc_rdat_REG[21] ( .CK(clk), .R(rst_n), .D(bimc_rdat[20]), .Q(bimc_rdat[21]), .QN( ));
Q_FDP1 \bimc_rdat_REG[22] ( .CK(clk), .R(rst_n), .D(bimc_rdat[21]), .Q(bimc_rdat[22]), .QN( ));
Q_FDP1 \bimc_rdat_REG[23] ( .CK(clk), .R(rst_n), .D(bimc_rdat[22]), .Q(bimc_rdat[23]), .QN( ));
Q_FDP1 \bimc_rdat_REG[24] ( .CK(clk), .R(rst_n), .D(bimc_rdat[23]), .Q(bimc_rdat[24]), .QN( ));
Q_FDP1 \bimc_rdat_REG[25] ( .CK(clk), .R(rst_n), .D(bimc_rdat[24]), .Q(bimc_rdat[25]), .QN( ));
Q_FDP1 \bimc_rdat_REG[26] ( .CK(clk), .R(rst_n), .D(bimc_rdat[25]), .Q(bimc_rdat[26]), .QN( ));
Q_FDP1 \bimc_rdat_REG[27] ( .CK(clk), .R(rst_n), .D(bimc_rdat[26]), .Q(bimc_rdat[27]), .QN( ));
Q_FDP1 \bimc_rdat_REG[28] ( .CK(clk), .R(rst_n), .D(bimc_rdat[27]), .Q(bimc_rdat[28]), .QN( ));
Q_FDP1 \bimc_rdat_REG[29] ( .CK(clk), .R(rst_n), .D(bimc_rdat[28]), .Q(bimc_rdat[29]), .QN( ));
Q_FDP1 \bimc_rdat_REG[30] ( .CK(clk), .R(rst_n), .D(bimc_rdat[29]), .Q(bimc_rdat[30]), .QN( ));
Q_FDP1 \bimc_rdat_REG[31] ( .CK(clk), .R(rst_n), .D(bimc_rdat[30]), .Q(bimc_rdat[31]), .QN( ));
Q_FDP1 \bimc_rdat_REG[32] ( .CK(clk), .R(rst_n), .D(bimc_rdat[31]), .Q(bimc_rdat[32]), .QN( ));
Q_FDP1 \bimc_rdat_REG[33] ( .CK(clk), .R(rst_n), .D(bimc_rdat[32]), .Q(bimc_rdat[33]), .QN( ));
Q_FDP1 \bimc_rdat_REG[34] ( .CK(clk), .R(rst_n), .D(bimc_rdat[33]), .Q(bimc_rdat[34]), .QN( ));
Q_FDP1 \bimc_rdat_REG[35] ( .CK(clk), .R(rst_n), .D(bimc_rdat[34]), .Q(bimc_rdat[35]), .QN( ));
Q_FDP1 \bimc_rdat_REG[36] ( .CK(clk), .R(rst_n), .D(bimc_rdat[35]), .Q(bimc_rdat[36]), .QN( ));
Q_FDP1 \bimc_rdat_REG[37] ( .CK(clk), .R(rst_n), .D(bimc_rdat[36]), .Q(bimc_rdat[37]), .QN( ));
Q_FDP1 \bimc_rdat_REG[38] ( .CK(clk), .R(rst_n), .D(bimc_rdat[37]), .Q(bimc_rdat[38]), .QN( ));
Q_FDP1 \bimc_rdat_REG[39] ( .CK(clk), .R(rst_n), .D(bimc_rdat[38]), .Q(bimc_rdat[39]), .QN( ));
Q_FDP1 \bimc_rdat_REG[40] ( .CK(clk), .R(rst_n), .D(bimc_rdat[39]), .Q(bimc_rdat[40]), .QN( ));
Q_FDP1 \bimc_rdat_REG[41] ( .CK(clk), .R(rst_n), .D(bimc_rdat[40]), .Q(bimc_rdat[41]), .QN( ));
Q_FDP1 \bimc_rdat_REG[42] ( .CK(clk), .R(rst_n), .D(bimc_rdat[41]), .Q(bimc_rdat[42]), .QN( ));
Q_FDP1 \bimc_rdat_REG[43] ( .CK(clk), .R(rst_n), .D(bimc_rdat[42]), .Q(bimc_rdat[43]), .QN( ));
Q_FDP1 \bimc_rdat_REG[44] ( .CK(clk), .R(rst_n), .D(bimc_rdat[43]), .Q(bimc_rdat[44]), .QN( ));
Q_FDP1 \bimc_rdat_REG[45] ( .CK(clk), .R(rst_n), .D(bimc_rdat[44]), .Q(bimc_rdat[45]), .QN( ));
Q_FDP1 \bimc_rdat_REG[46] ( .CK(clk), .R(rst_n), .D(bimc_rdat[45]), .Q(bimc_rdat[46]), .QN( ));
Q_FDP1 \bimc_rdat_REG[47] ( .CK(clk), .R(rst_n), .D(bimc_rdat[46]), .Q(bimc_rdat[47]), .QN( ));
Q_FDP1 \bimc_rdat_REG[48] ( .CK(clk), .R(rst_n), .D(bimc_rdat[47]), .Q(bimc_rdat[48]), .QN( ));
Q_FDP1 \bimc_rdat_REG[49] ( .CK(clk), .R(rst_n), .D(bimc_rdat[48]), .Q(bimc_rdat[49]), .QN( ));
Q_FDP1 \bimc_rdat_REG[50] ( .CK(clk), .R(rst_n), .D(bimc_rdat[49]), .Q(bimc_rdat[50]), .QN( ));
Q_FDP1 \bimc_rdat_REG[51] ( .CK(clk), .R(rst_n), .D(bimc_rdat[50]), .Q(bimc_rdat[51]), .QN( ));
Q_FDP1 \bimc_rdat_REG[52] ( .CK(clk), .R(rst_n), .D(bimc_rdat[51]), .Q(bimc_rdat[52]), .QN( ));
Q_FDP1 \bimc_rdat_REG[53] ( .CK(clk), .R(rst_n), .D(bimc_rdat[52]), .Q(bimc_rdat[53]), .QN( ));
Q_FDP1 \bimc_rdat_REG[54] ( .CK(clk), .R(rst_n), .D(bimc_rdat[53]), .Q(bimc_rdat[54]), .QN( ));
Q_FDP1 \bimc_rdat_REG[55] ( .CK(clk), .R(rst_n), .D(bimc_rdat[54]), .Q(bimc_rdat[55]), .QN( ));
Q_FDP1 \bimc_rdat_REG[56] ( .CK(clk), .R(rst_n), .D(bimc_rdat[55]), .Q(bimc_rdat[56]), .QN( ));
Q_FDP1 \bimc_rdat_REG[57] ( .CK(clk), .R(rst_n), .D(bimc_rdat[56]), .Q(bimc_rdat[57]), .QN( ));
Q_FDP1 \bimc_rdat_REG[58] ( .CK(clk), .R(rst_n), .D(bimc_rdat[57]), .Q(bimc_rdat[58]), .QN( ));
Q_FDP1 \bimc_rdat_REG[59] ( .CK(clk), .R(rst_n), .D(bimc_rdat[58]), .Q(bimc_rdat[59]), .QN( ));
Q_FDP1 \bimc_rdat_REG[60] ( .CK(clk), .R(rst_n), .D(bimc_rdat[59]), .Q(bimc_rdat[60]), .QN( ));
Q_FDP1 \bimc_rdat_REG[61] ( .CK(clk), .R(rst_n), .D(bimc_rdat[60]), .Q(bimc_rdat[61]), .QN( ));
Q_FDP1 \bimc_rdat_REG[62] ( .CK(clk), .R(rst_n), .D(bimc_rdat[61]), .Q(bimc_rdat[62]), .QN( ));
Q_FDP1 \bimc_rdat_REG[63] ( .CK(clk), .R(rst_n), .D(bimc_rdat[62]), .Q(bimc_rdat[63]), .QN( ));
Q_FDP1 \bimc_rdat_REG[64] ( .CK(clk), .R(rst_n), .D(bimc_rdat[63]), .Q(bimc_rdat[64]), .QN( ));
Q_FDP1 \bimc_rdat_REG[65] ( .CK(clk), .R(rst_n), .D(bimc_rdat[64]), .Q(bimc_rdat[65]), .QN( ));
Q_FDP1 \bimc_rdat_REG[66] ( .CK(clk), .R(rst_n), .D(bimc_rdat[65]), .Q(bimc_rdat[66]), .QN( ));
Q_FDP1 \bimc_rdat_REG[67] ( .CK(clk), .R(rst_n), .D(bimc_rdat[66]), .Q(bimc_rdat[67]), .QN( ));
Q_FDP1 \bimc_rdat_REG[68] ( .CK(clk), .R(rst_n), .D(bimc_rdat[67]), .Q(bimc_rdat[68]), .QN( ));
Q_FDP1 \bimc_rdat_REG[69] ( .CK(clk), .R(rst_n), .D(bimc_rdat[68]), .Q(bimc_rdat[69]), .QN( ));
Q_FDP1 \bimc_rdat_REG[70] ( .CK(clk), .R(rst_n), .D(bimc_rdat[69]), .Q(bimc_rdat[70]), .QN( ));
Q_FDP1 \bimc_rdat_REG[71] ( .CK(clk), .R(rst_n), .D(bimc_rdat[70]), .Q(bimc_rdat[71]), .QN( ));
Q_OA21 U1599 ( .A0(n1168), .A1(n1177), .B0(n1169), .Z(n1170));
Q_OA21 U1600 ( .A0(n1168), .A1(n1179), .B0(n1169), .Z(n1171));
Q_OA21 U1601 ( .A0(n1168), .A1(n1181), .B0(n1169), .Z(n1172));
Q_OA21 U1602 ( .A0(n1168), .A1(n1183), .B0(n1169), .Z(n1173));
Q_OA21 U1603 ( .A0(n1168), .A1(n1185), .B0(n1169), .Z(n1174));
Q_OA21 U1604 ( .A0(n1168), .A1(n1187), .B0(n1169), .Z(n1175));
Q_OA21 U1605 ( .A0(n1168), .A1(n1188), .B0(n1169), .Z(n1176));
Q_XOR2 U1606 ( .A0(bm_cnt[6]), .A1(n1178), .Z(n1177));
Q_AD01HF U1607 ( .A0(bm_cnt[5]), .B0(n1180), .S(n1179), .CO(n1178));
Q_AD01HF U1608 ( .A0(bm_cnt[4]), .B0(n1182), .S(n1181), .CO(n1180));
Q_AD01HF U1609 ( .A0(bm_cnt[3]), .B0(n1184), .S(n1183), .CO(n1182));
Q_AD01HF U1610 ( .A0(bm_cnt[2]), .B0(n1186), .S(n1185), .CO(n1184));
Q_AD01HF U1611 ( .A0(bm_cnt[1]), .B0(bm_cnt[0]), .S(n1187), .CO(n1186));
Q_NR03 U1612 ( .A0(bm_cnt[0]), .A1(n1191), .A2(n1190), .Z(n1189));
Q_OR03 U1613 ( .A0(n1193), .A1(bm_cnt[2]), .A2(bm_cnt[1]), .Z(n1190));
Q_OR03 U1614 ( .A0(n1192), .A1(bm_cnt[5]), .A2(bm_cnt[4]), .Z(n1191));
Q_AN03 U1615 ( .A0(bm_cnt[0]), .A1(n1195), .A2(n1194), .Z(n1168));
Q_AN03 U1616 ( .A0(bm_cnt[3]), .A1(bm_cnt[2]), .A2(bm_cnt[1]), .Z(n1194));
Q_AN03 U1617 ( .A0(bm_cnt[6]), .A1(bm_cnt[5]), .A2(bm_cnt[4]), .Z(n1195));
Q_OA21 U1618 ( .A0(n1197), .A1(n1198), .B0(n1196), .Z(tstate_text[0]));
Q_NR02 U1619 ( .A0(n1199), .A1(n1200), .Z(tstate_text[3]));
Q_OA21 U1620 ( .A0(n1202), .A1(n1203), .B0(n1201), .Z(tstate_text[4]));
Q_INV U1621 ( .A(n1204), .Z(tstate_text[8]));
Q_OA21 U1622 ( .A0(n1197), .A1(n1205), .B0(n1196), .Z(n1204));
Q_AN02 U1623 ( .A0(n1206), .A1(n1201), .Z(n1197));
Q_NR02 U1624 ( .A0(n1199), .A1(tstate_text[62]), .Z(tstate_text[9]));
Q_ND02 U1625 ( .A0(n1201), .A1(n1207), .Z(tstate_text[10]));
Q_AO21 U1626 ( .A0(n1208), .A1(tstate[0]), .B0(n1203), .Z(n1207));
Q_AO21 U1627 ( .A0(tstate[3]), .A1(tstate[1]), .B0(n1202), .Z(n1208));
Q_AO21 U1628 ( .A0(n1210), .A1(n1211), .B0(n1209), .Z(tstate_text[11]));
Q_INV U1629 ( .A(n1213), .Z(tstate_text[12]));
Q_AO21 U1630 ( .A0(n1215), .A1(n1201), .B0(n1214), .Z(n1213));
Q_AO21 U1631 ( .A0(n1196), .A1(n1217), .B0(n1216), .Z(n1215));
Q_NR02 U1632 ( .A0(n1218), .A1(n1200), .Z(tstate_text[16]));
Q_INV U1633 ( .A(n1218), .Z(tstate_text[17]));
Q_AN02 U1634 ( .A0(n1219), .A1(n1217), .Z(n1218));
Q_INV U1635 ( .A(n1220), .Z(tstate_text[18]));
Q_NR02 U1636 ( .A0(tstate[3]), .A1(tstate[1]), .Z(n1202));
Q_OA21 U1637 ( .A0(n1201), .A1(n1222), .B0(n1202), .Z(n1220));
Q_AN02 U1638 ( .A0(tstate[2]), .A1(tstate[0]), .Z(n1222));
Q_INV U1639 ( .A(n1223), .Z(tstate_text[19]));
Q_OA21 U1640 ( .A0(n1224), .A1(n1198), .B0(n1196), .Z(n1223));
Q_AN02 U1641 ( .A0(tstate[2]), .A1(n1225), .Z(n1198));
Q_NR02 U1642 ( .A0(n1205), .A1(tstate[2]), .Z(n1224));
Q_AN02 U1643 ( .A0(n1219), .A1(n1227), .Z(tstate_text[20]));
Q_NR02 U1644 ( .A0(n1228), .A1(tstate_text[62]), .Z(tstate_text[5]));
Q_AO21 U1645 ( .A0(n1219), .A1(n1212), .B0(n1200), .Z(tstate_text[24]));
Q_NR02 U1646 ( .A0(n1199), .A1(tstate_text[56]), .Z(tstate_text[25]));
Q_NR02 U1647 ( .A0(n1229), .A1(n1214), .Z(tstate_text[26]));
Q_NR02 U1648 ( .A0(n1228), .A1(n1230), .Z(tstate_text[27]));
Q_AN02 U1649 ( .A0(n1231), .A1(n1201), .Z(n1228));
Q_AO21 U1650 ( .A0(n1196), .A1(n1225), .B0(n1216), .Z(n1231));
Q_OA21 U1651 ( .A0(n1232), .A1(n1196), .B0(n1205), .Z(tstate_text[28]));
Q_ND02 U1652 ( .A0(n1219), .A1(n1225), .Z(tstate_text[30]));
Q_NR02 U1653 ( .A0(n1233), .A1(tstate_text[70]), .Z(tstate_text[32]));
Q_NR02 U1654 ( .A0(n1234), .A1(tstate_text[94]), .Z(tstate_text[33]));
Q_OA21 U1655 ( .A0(n1235), .A1(n1236), .B0(n1201), .Z(n1234));
Q_AN02 U1656 ( .A0(tstate[0]), .A1(n1237), .Z(tstate_text[34]));
Q_AO21 U1657 ( .A0(n1232), .A1(tstate[1]), .B0(n1238), .Z(n1237));
Q_NR02 U1658 ( .A0(n1199), .A1(tstate_text[70]), .Z(tstate_text[35]));
Q_OA21 U1659 ( .A0(n1216), .A1(n1239), .B0(n1201), .Z(tstate_text[36]));
Q_INV U1660 ( .A(n1240), .Z(tstate_text[29]));
Q_AO21 U1661 ( .A0(n1216), .A1(n1201), .B0(tstate_text[62]), .Z(n1240));
Q_INV U1662 ( .A(n1229), .Z(tstate_text[38]));
Q_AN02 U1663 ( .A0(n1219), .A1(n1206), .Z(n1229));
Q_OR02 U1664 ( .A0(n1241), .A1(n1200), .Z(tstate_text[40]));
Q_OR02 U1665 ( .A0(tstate_text[67]), .A1(n1242), .Z(n1200));
Q_NR02 U1666 ( .A0(n1199), .A1(n1243), .Z(tstate_text[41]));
Q_INV U1667 ( .A(n1244), .Z(tstate_text[42]));
Q_OA21 U1668 ( .A0(n1245), .A1(n1246), .B0(n1201), .Z(n1244));
Q_NR02 U1669 ( .A0(n1199), .A1(n1209), .Z(tstate_text[1]));
Q_OR02 U1670 ( .A0(n1214), .A1(tstate_text[60]), .Z(n1209));
Q_NR02 U1671 ( .A0(n1241), .A1(tstate_text[62]), .Z(tstate_text[45]));
Q_AN02 U1672 ( .A0(n1232), .A1(n1205), .Z(n1241));
Q_INV U1673 ( .A(n1233), .Z(tstate_text[46]));
Q_AN02 U1674 ( .A0(n1219), .A1(n1226), .Z(n1233));
Q_INV U1675 ( .A(n1205), .Z(n1226));
Q_NR02 U1676 ( .A0(n1199), .A1(tstate_text[94]), .Z(tstate_text[48]));
Q_NR02 U1677 ( .A0(n1199), .A1(n1242), .Z(tstate_text[50]));
Q_AN02 U1678 ( .A0(n1201), .A1(n1203), .Z(tstate_text[51]));
Q_INV U1679 ( .A(n1247), .Z(tstate_text[52]));
Q_OA21 U1680 ( .A0(n1245), .A1(n1203), .B0(n1201), .Z(n1247));
Q_OR02 U1681 ( .A0(n1239), .A1(n1246), .Z(n1203));
Q_AN02 U1682 ( .A0(n1196), .A1(n1205), .Z(n1246));
Q_AN02 U1683 ( .A0(tstate[3]), .A1(n1227), .Z(n1239));
Q_INV U1684 ( .A(n1199), .Z(tstate_text[54]));
Q_AN02 U1685 ( .A0(n1201), .A1(n1245), .Z(n1199));
Q_OR02 U1686 ( .A0(n1216), .A1(n1236), .Z(n1245));
Q_AN02 U1687 ( .A0(n1206), .A1(n1196), .Z(n1236));
Q_OR02 U1688 ( .A0(n1225), .A1(n1217), .Z(n1206));
Q_AN02 U1689 ( .A0(tstate[1]), .A1(n1212), .Z(n1217));
Q_AN02 U1690 ( .A0(tstate[3]), .A1(n1205), .Z(n1235));
Q_AO21 U1691 ( .A0(n1196), .A1(n1227), .B0(n1235), .Z(n1216));
Q_OR02 U1692 ( .A0(n1214), .A1(tstate_text[94]), .Z(tstate_text[44]));
Q_AN02 U1693 ( .A0(n1219), .A1(n1205), .Z(tstate_text[60]));
Q_NR02 U1694 ( .A0(tstate[3]), .A1(tstate[2]), .Z(n1219));
Q_INV U1695 ( .A(tstate_text[62]), .Z(tstate_text[53]));
Q_OR02 U1696 ( .A0(n1214), .A1(n1242), .Z(tstate_text[62]));
Q_AN03 U1697 ( .A0(n1196), .A1(tstate[0]), .A2(n1248), .Z(n1242));
Q_AO21 U1698 ( .A0(tstate[2]), .A1(n1221), .B0(n1211), .Z(n1248));
Q_AN02 U1699 ( .A0(n1201), .A1(tstate[1]), .Z(n1211));
Q_OR02 U1700 ( .A0(n1243), .A1(tstate_text[67]), .Z(n1214));
Q_AN02 U1701 ( .A0(n1238), .A1(n1205), .Z(n1243));
Q_AN02 U1702 ( .A0(tstate[1]), .A1(tstate[0]), .Z(n1205));
Q_AN02 U1703 ( .A0(n1232), .A1(n1227), .Z(tstate_text[58]));
Q_NR02 U1704 ( .A0(tstate[1]), .A1(tstate[0]), .Z(n1227));
Q_INV U1705 ( .A(tstate_text[70]), .Z(tstate_text[69]));
Q_AN02 U1706 ( .A0(n1221), .A1(n1249), .Z(tstate_text[70]));
Q_AN02 U1707 ( .A0(n1238), .A1(tstate[0]), .Z(n1230));
Q_AO21 U1708 ( .A0(n1232), .A1(n1212), .B0(n1230), .Z(n1249));
Q_AN02 U1709 ( .A0(tstate[3]), .A1(n1201), .Z(n1232));
Q_INV U1710 ( .A(tstate_text[94]), .Z(tstate_text[77]));
Q_AN02 U1711 ( .A0(n1238), .A1(n1225), .Z(tstate_text[49]));
Q_AN02 U1712 ( .A0(n1221), .A1(tstate[0]), .Z(n1225));
Q_AN02 U1713 ( .A0(n1196), .A1(tstate[2]), .Z(n1238));
Q_OR02 U1714 ( .A0(n1250), .A1(n1251), .Z(rstate_text[0]));
Q_AO21 U1715 ( .A0(n1252), .A1(n1253), .B0(n1254), .Z(n1251));
Q_AO21 U1716 ( .A0(n1256), .A1(n1257), .B0(n1255), .Z(n1250));
Q_OR02 U1717 ( .A0(n1258), .A1(n1259), .Z(n1252));
Q_NR02 U1718 ( .A0(rstate[2]), .A1(rstate[0]), .Z(n1258));
Q_INV U1719 ( .A(rstate_text[11]), .Z(rstate_text[3]));
Q_NR02 U1720 ( .A0(n1262), .A1(n1263), .Z(rstate_text[9]));
Q_OR02 U1721 ( .A0(n1264), .A1(n1265), .Z(rstate_text[11]));
Q_OR03 U1722 ( .A0(n1266), .A1(n1267), .A2(n1254), .Z(n1265));
Q_OA21 U1723 ( .A0(n1260), .A1(n1268), .B0(n1253), .Z(n1264));
Q_NR02 U1724 ( .A0(n1269), .A1(n1270), .Z(rstate_text[1]));
Q_NR02 U1725 ( .A0(n1271), .A1(n1255), .Z(rstate_text[17]));
Q_OA21 U1726 ( .A0(n1272), .A1(n1259), .B0(n1253), .Z(n1271));
Q_ND02 U1727 ( .A0(n1273), .A1(n1274), .Z(rstate_text[18]));
Q_INV U1728 ( .A(n1259), .Z(n1274));
Q_NR03 U1729 ( .A0(n1276), .A1(n1267), .A2(n1275), .Z(rstate_text[19]));
Q_AN02 U1730 ( .A0(n1277), .A1(n1278), .Z(n1267));
Q_OA21 U1731 ( .A0(n1279), .A1(n1268), .B0(n1253), .Z(n1275));
Q_OR02 U1732 ( .A0(n1280), .A1(n1263), .Z(rstate_text[24]));
Q_OA21 U1733 ( .A0(n1279), .A1(n1259), .B0(n1253), .Z(n1280));
Q_NR02 U1734 ( .A0(n1281), .A1(n1282), .Z(rstate_text[8]));
Q_OA21 U1735 ( .A0(n1283), .A1(n1268), .B0(n1253), .Z(n1281));
Q_NR02 U1736 ( .A0(n1284), .A1(rstate[2]), .Z(n1283));
Q_INV U1737 ( .A(n1285), .Z(rstate_text[16]));
Q_OA21 U1738 ( .A0(n1262), .A1(n1255), .B0(n1261), .Z(n1285));
Q_ND02 U1739 ( .A0(n1261), .A1(n1286), .Z(rstate_text[27]));
Q_MX02 U1740 ( .S(rstate[1]), .A0(n1288), .A1(n1287), .Z(n1286));
Q_OR02 U1741 ( .A0(n1256), .A1(n1277), .Z(n1287));
Q_NR02 U1742 ( .A0(n1290), .A1(n1291), .Z(rstate_text[32]));
Q_INV U1743 ( .A(n1292), .Z(rstate_text[33]));
Q_OA21 U1744 ( .A0(n1279), .A1(n1293), .B0(n1253), .Z(n1292));
Q_NR02 U1745 ( .A0(n1278), .A1(rstate[2]), .Z(n1279));
Q_OR02 U1746 ( .A0(n1294), .A1(n1282), .Z(rstate_text[34]));
Q_NR02 U1747 ( .A0(n1295), .A1(n1291), .Z(rstate_text[35]));
Q_AO21 U1748 ( .A0(n1253), .A1(n1278), .B0(n1270), .Z(rstate_text[36]));
Q_OR02 U1749 ( .A0(rstate[3]), .A1(rstate[0]), .Z(rstate_text[41]));
Q_OA21 U1750 ( .A0(n1260), .A1(n1259), .B0(n1253), .Z(n1269));
Q_NR02 U1751 ( .A0(n1295), .A1(n1270), .Z(rstate_text[42]));
Q_NR02 U1752 ( .A0(n1296), .A1(n1270), .Z(rstate_text[43]));
Q_OA21 U1753 ( .A0(n1297), .A1(n1259), .B0(n1253), .Z(n1296));
Q_NR02 U1754 ( .A0(n1299), .A1(rstate[2]), .Z(n1297));
Q_INV U1755 ( .A(n1299), .Z(n1298));
Q_OR02 U1756 ( .A0(rstate_text[73]), .A1(n1270), .Z(rstate_text[44]));
Q_NR02 U1757 ( .A0(n1295), .A1(rstate_text[91]), .Z(rstate_text[48]));
Q_OA21 U1758 ( .A0(n1300), .A1(n1293), .B0(n1253), .Z(n1295));
Q_OR02 U1759 ( .A0(rstate_text[40]), .A1(n1282), .Z(rstate_text[49]));
Q_AN02 U1760 ( .A0(n1301), .A1(n1253), .Z(rstate_text[40]));
Q_AO21 U1761 ( .A0(n1260), .A1(rstate[0]), .B0(n1259), .Z(n1301));
Q_NR02 U1762 ( .A0(n1302), .A1(n1282), .Z(rstate_text[50]));
Q_AN02 U1763 ( .A0(n1303), .A1(n1261), .Z(n1282));
Q_AO21 U1764 ( .A0(n1277), .A1(rstate[1]), .B0(n1304), .Z(n1303));
Q_OA21 U1765 ( .A0(n1272), .A1(n1268), .B0(n1253), .Z(n1302));
Q_AN02 U1766 ( .A0(rstate[2]), .A1(n1278), .Z(n1268));
Q_NR02 U1767 ( .A0(n1306), .A1(rstate[2]), .Z(n1272));
Q_NR02 U1768 ( .A0(n1305), .A1(n1291), .Z(rstate_text[52]));
Q_OA21 U1769 ( .A0(n1260), .A1(n1293), .B0(n1253), .Z(n1305));
Q_NR02 U1770 ( .A0(n1294), .A1(n1270), .Z(rstate_text[5]));
Q_OA21 U1771 ( .A0(n1307), .A1(n1259), .B0(n1253), .Z(n1294));
Q_NR02 U1772 ( .A0(n1257), .A1(rstate[2]), .Z(n1307));
Q_INV U1773 ( .A(n1257), .Z(n1308));
Q_INV U1774 ( .A(n1290), .Z(rstate_text[38]));
Q_AN02 U1775 ( .A0(n1288), .A1(n1257), .Z(n1290));
Q_NR02 U1776 ( .A0(rstate[3]), .A1(rstate[2]), .Z(n1288));
Q_OR02 U1777 ( .A0(rstate_text[51]), .A1(rstate_text[83]), .Z(rstate_text[56]));
Q_OA21 U1778 ( .A0(n1309), .A1(n1293), .B0(n1253), .Z(rstate_text[51]));
Q_AN02 U1779 ( .A0(rstate[2]), .A1(n1299), .Z(n1293));
Q_OR02 U1780 ( .A0(n1310), .A1(rstate_text[60]), .Z(rstate_text[57]));
Q_AO21 U1781 ( .A0(n1277), .A1(n1299), .B0(n1266), .Z(rstate_text[60]));
Q_AN02 U1782 ( .A0(n1289), .A1(rstate[0]), .Z(n1299));
Q_INV U1783 ( .A(rstate_text[62]), .Z(rstate_text[61]));
Q_OR02 U1784 ( .A0(n1310), .A1(n1270), .Z(rstate_text[62]));
Q_OR02 U1785 ( .A0(n1304), .A1(n1254), .Z(n1270));
Q_OA21 U1786 ( .A0(n1309), .A1(n1259), .B0(n1253), .Z(n1310));
Q_AN02 U1787 ( .A0(n1306), .A1(n1260), .Z(n1309));
Q_OR02 U1788 ( .A0(n1278), .A1(n1284), .Z(n1306));
Q_OR02 U1789 ( .A0(rstate_text[97]), .A1(rstate_text[83]), .Z(rstate_text[66]));
Q_OR02 U1790 ( .A0(rstate_text[76]), .A1(n1291), .Z(rstate_text[59]));
Q_OR02 U1791 ( .A0(rstate_text[97]), .A1(n1291), .Z(rstate_text[81]));
Q_AN02 U1792 ( .A0(n1304), .A1(rstate[0]), .Z(n1291));
Q_OR02 U1793 ( .A0(rstate_text[73]), .A1(rstate_text[83]), .Z(rstate_text[82]));
Q_OR02 U1794 ( .A0(rstate_text[73]), .A1(rstate_text[91]), .Z(rstate_text[68]));
Q_AN02 U1795 ( .A0(n1311), .A1(n1273), .Z(rstate_text[72]));
Q_AN02 U1796 ( .A0(n1253), .A1(rstate[0]), .Z(n1273));
Q_AN02 U1797 ( .A0(n1277), .A1(n1261), .Z(rstate_text[91]));
Q_OA21 U1798 ( .A0(n1262), .A1(n1304), .B0(rstate[0]), .Z(rstate_text[28]));
Q_AN02 U1799 ( .A0(n1311), .A1(n1253), .Z(n1262));
Q_OR02 U1800 ( .A0(n1266), .A1(n1255), .Z(n1304));
Q_AN02 U1801 ( .A0(n1256), .A1(rstate[1]), .Z(n1266));
Q_OR02 U1802 ( .A0(n1300), .A1(n1259), .Z(n1311));
Q_AN02 U1803 ( .A0(n1260), .A1(rstate[1]), .Z(n1300));
Q_INV U1804 ( .A(rstate_text[94]), .Z(rstate_text[69]));
Q_OR02 U1805 ( .A0(rstate_text[76]), .A1(rstate_text[83]), .Z(rstate_text[58]));
Q_AN02 U1806 ( .A0(n1312), .A1(n1253), .Z(rstate_text[76]));
Q_OR02 U1807 ( .A0(n1263), .A1(n1254), .Z(rstate_text[74]));
Q_AN02 U1808 ( .A0(n1277), .A1(n1257), .Z(n1254));
Q_AN02 U1809 ( .A0(rstate[1]), .A1(n1261), .Z(n1257));
Q_OR02 U1810 ( .A0(n1276), .A1(n1255), .Z(n1263));
Q_AN02 U1811 ( .A0(n1277), .A1(n1289), .Z(n1255));
Q_AN02 U1812 ( .A0(n1256), .A1(n1284), .Z(n1276));
Q_AN02 U1813 ( .A0(rstate[2]), .A1(n1289), .Z(n1259));
Q_AO21 U1814 ( .A0(n1260), .A1(n1284), .B0(n1259), .Z(n1312));
Q_AN02 U1815 ( .A0(rstate[1]), .A1(rstate[0]), .Z(n1284));
Q_AN02 U1816 ( .A0(n1256), .A1(n1278), .Z(rstate_text[84]));
Q_NR02 U1817 ( .A0(rstate[1]), .A1(rstate[0]), .Z(n1278));
Q_INV U1818 ( .A(rstate_text[102]), .Z(rstate_text[101]));
Q_AN02 U1819 ( .A0(n1261), .A1(n1313), .Z(rstate_text[64]));
Q_AN02 U1820 ( .A0(rstate[3]), .A1(n1260), .Z(n1277));
Q_AO21 U1821 ( .A0(n1256), .A1(n1289), .B0(n1277), .Z(n1313));
Q_AN02 U1822 ( .A0(n1253), .A1(rstate[2]), .Z(n1256));
ixc_assign_4 _zz_strnp_0 ( bm_type[3:0], bimc_dat[71:68]);
ixc_assign_8 _zz_strnp_1 ( bm_op[7:0], bimc_dat[67:60]);
ixc_assign_12 _zz_strnp_2 ( bm_mem[11:0], bimc_dat[59:48]);
ixc_assign_16 _zz_strnp_3 ( bm_addr[15:0], bimc_dat[47:32]);
ixc_assign_32 _zz_strnp_4 ( bm_dat[31:0], bimc_dat[31:0]);
ixc_assign _zz_strnp_5 ( rcv_chk, bimc_chk);
ixc_assign _zz_strnp_6 ( rcv_frm, bimc_frm);
ixc_assign _zz_strnp_7 ( rcv_resp, bm_resp);
ixc_assign_72 _zz_strnp_8 ( rcv_dat[71:0], bimc_dat[71:0]);
ixc_assign_73 _zz_strnp_9 ( cputx_frame[72:0], { n1318, cputx_type[3], 
	cputx_type[2], cputx_type[1], cputx_type[0], cputx_op[7], 
	cputx_op[6], cputx_op[5], cputx_op[4], cputx_op[3], cputx_op[2], 
	cputx_op[1], cputx_op[0], cputx_mem[11], cputx_mem[10], cputx_mem[9], 
	cputx_mem[8], cputx_mem[7], cputx_mem[6], cputx_mem[5], cputx_mem[4], 
	cputx_mem[3], cputx_mem[2], cputx_mem[1], cputx_mem[0], 
	cputx_addr[15], cputx_addr[14], cputx_addr[13], cputx_addr[12], 
	cputx_addr[11], cputx_addr[10], cputx_addr[9], cputx_addr[8], 
	cputx_addr[7], cputx_addr[6], cputx_addr[5], cputx_addr[4], 
	cputx_addr[3], cputx_addr[2], cputx_addr[1], cputx_addr[0], 
	cputx_dat[31], cputx_dat[30], cputx_dat[29], cputx_dat[28], 
	cputx_dat[27], cputx_dat[26], cputx_dat[25], cputx_dat[24], 
	cputx_dat[23], cputx_dat[22], cputx_dat[21], cputx_dat[20], 
	cputx_dat[19], cputx_dat[18], cputx_dat[17], cputx_dat[16], 
	cputx_dat[15], cputx_dat[14], cputx_dat[13], cputx_dat[12], 
	cputx_dat[11], cputx_dat[10], cputx_dat[9], cputx_dat[8], 
	cputx_dat[7], cputx_dat[6], cputx_dat[5], cputx_dat[4], cputx_dat[3], 
	cputx_dat[2], cputx_dat[1], cputx_dat[0]});
ixc_assign_32 _zz_strnp_10 ( bimc_cmd0_data[31:0], o_bimc_cmd0[31:0]);
ixc_assign_16 _zz_strnp_11 ( bimc_cmd1_addr[15:0], o_bimc_cmd1[15:0]);
ixc_assign_12 _zz_strnp_12 ( bimc_cmd1_mem[11:0], o_bimc_cmd1[27:16]);
ixc_assign_4 _zz_strnp_13 ( bimc_cmd1_memtype[3:0], o_bimc_cmd1[31:28]);
ixc_assign_8 _zz_strnp_14 ( bimc_cmd2_opcode[7:0], o_bimc_cmd2[7:0]);
Q_AN02 U1838 ( .A0(o_bimc_cmd2[8]), .A1(n1317), .Z(bimc_cmd2_write_notify_ev));
ixc_assign_2 _zz_strnp_15 ( bimc_eccpar_debug_eccpar_corrupt[1:0], 
	o_bimc_eccpar_debug[17:16]);
ixc_assign_2 _zz_strnp_16 ( bimc_eccpar_debug_eccpar_disable[1:0], 
	o_bimc_eccpar_debug[21:20]);
ixc_assign_4 _zz_strnp_17 ( bimc_eccpar_debug_jabber_off[3:0], 
	o_bimc_eccpar_debug[27:24]);
ixc_assign_12 _zz_strnp_18 ( bimc_eccpar_debug_memaddr[11:0], 
	o_bimc_eccpar_debug[11:0]);
ixc_assign_4 _zz_strnp_19 ( bimc_eccpar_debug_memtype[3:0], 
	o_bimc_eccpar_debug[15:12]);
Q_AN02 U1844 ( .A0(o_bimc_eccpar_debug[22]), .A1(n1316), .Z(bimc_eccpar_debug_write_notify_ev));
ixc_assign _zz_strnp_20 ( bimc_global_config_mem_wr_init, 
	o_bimc_global_config[3]);
ixc_assign _zz_strnp_21 ( bimc_global_config_poll_ecc_par_error, 
	o_bimc_global_config[4]);
ixc_assign_26 _zz_strnp_22 ( bimc_global_config_poll_ecc_par_timer[25:0], 
	o_bimc_global_config[31:6]);
ixc_assign _zz_strnp_23 ( bimc_global_config_soft_reset, 
	o_bimc_global_config[0]);
Q_OR03 U1849 ( .A0(bimc_monitor_uncorrectable_ecc_error_din), .A1(bimc_monitor_correctable_ecc_error_din), .A2(bimc_monitor_parity_error_din), .Z(bimc_ecc_error_c));
ixc_assign _zz_strnp_24 ( debug_write_en, o_bimc_global_config[5]);
ixc_assign_2 _zz_strnp_25 ( i_bimc_global_config[1:0], 
	o_bimc_global_config[1:0]);
ixc_assign _zz_strnp_26 ( i_bimc_global_config[2], 
	bimc_global_config_bimc_mem_init_done_din);
ixc_assign_2 _zz_strnp_27 ( i_bimc_global_config[4:3], 
	o_bimc_global_config[4:3]);
ixc_assign _zz_strnp_28 ( i_bimc_global_config[5], debug_write_en);
ixc_assign_26 _zz_strnp_29 ( i_bimc_global_config[31:6], 
	o_bimc_global_config[31:6]);
ixc_assign _zz_strnp_30 ( i_bimc_cmd2[9], bimc_cmd2_sent);
ixc_assign_8 _zz_strnp_31 ( i_bimc_cmd2[7:0], o_bimc_cmd2[7:0]);
ixc_assign _zz_strnp_32 ( i_bimc_cmd2[8], o_bimc_cmd2[8]);
ixc_assign _zz_strnp_33 ( i_bimc_cmd2[10], o_bimc_cmd2[10]);
ixc_assign_23 _zz_strnp_34 ( i_bimc_eccpar_debug[22:0], 
	o_bimc_eccpar_debug[22:0]);
ixc_assign _zz_strnp_35 ( i_bimc_eccpar_debug[23], bimc_eccpar_debug_sent);
ixc_assign_5 _zz_strnp_36 ( i_bimc_eccpar_debug[28:24], 
	o_bimc_eccpar_debug[28:24]);
ixc_assign _zz_strnp_37 ( i_bimc_monitor[0], 
	bimc_monitor_uncorrectable_ecc_error_din);
ixc_assign _zz_strnp_38 ( i_bimc_monitor[1], 
	bimc_monitor_correctable_ecc_error_din);
ixc_assign _zz_strnp_39 ( i_bimc_monitor[2], bimc_monitor_parity_error_din);
ixc_assign _zz_strnp_40 ( i_bimc_monitor[4], 
	bimc_monitor_bimc_chain_rcv_error_din);
ixc_assign _zz_strnp_41 ( i_bimc_monitor[5], 
	bimc_monitor_rcv_invalid_opcode_din);
ixc_assign _zz_strnp_42 ( i_bimc_monitor[6], bimc_monitor_unanswered_read_din);
ixc_assign_32 _zz_strnp_43 ( i_bimc_ecc_uncorrectable_error_cnt[31:0], 
	bimc_ecc_uncorrectable_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_44 ( i_bimc_ecc_correctable_error_cnt[31:0], 
	bimc_ecc_correctable_error_cnt[31:0]);
ixc_assign_32 _zz_strnp_45 ( i_bimc_parity_error_cnt[31:0], 
	bimc_parity_error_cnt[31:0]);
ixc_assign_12 _zz_strnp_46 ( i_bimc_memid[11:0], number_of_memories[11:0]);
ixc_assign_32 _zz_strnp_47 ( i_bimc_rxcmd0[31:0], 
	bimc_rxcmd0_data_din[31:0]);
ixc_assign_16 _zz_strnp_48 ( i_bimc_rxcmd1[15:0], 
	bimc_rxcmd1_addr_din[15:0]);
ixc_assign_12 _zz_strnp_49 ( i_bimc_rxcmd1[27:16], bimc_rxcmd1_mem_din[11:0]);
ixc_assign_4 _zz_strnp_50 ( i_bimc_rxcmd1[31:28], 
	bimc_rxcmd1_memtype_din[3:0]);
ixc_assign_8 _zz_strnp_51 ( i_bimc_rxcmd2[7:0], bimc_rxcmd2_opcode_din[7:0]);
ixc_assign _zz_strnp_52 ( i_bimc_rxcmd2[8], bimc_rxcmd2_rxflag_din);
ixc_assign _zz_strnp_53 ( i_bimc_rxcmd2[9], o_bimc_rxcmd2[9]);
ixc_assign_32 _zz_strnp_54 ( i_bimc_dbgcmd0[31:0], 
	bimc_dbgcmd0_data_din[31:0]);
ixc_assign_16 _zz_strnp_55 ( i_bimc_dbgcmd1[15:0], 
	bimc_dbgcmd1_addr_din[15:0]);
ixc_assign_12 _zz_strnp_56 ( i_bimc_dbgcmd1[27:16], 
	bimc_dbgcmd1_mem_din[11:0]);
ixc_assign_4 _zz_strnp_57 ( i_bimc_dbgcmd1[31:28], 
	bimc_dbgcmd1_memtype_din[3:0]);
ixc_assign_8 _zz_strnp_58 ( i_bimc_dbgcmd2[7:0], bimc_dbgcmd2_opcode_din[7:0]);
ixc_assign _zz_strnp_59 ( i_bimc_dbgcmd2[8], bimc_dbgcmd2_rxflag_din);
ixc_assign _zz_strnp_60 ( i_bimc_dbgcmd2[9], o_bimc_dbgcmd2[9]);
ixc_assign_32 _zz_strnp_61 ( i_bimc_rxrsp0[31:0], 
	bimc_rxrsp0_data_din[31:0]);
ixc_assign_32 _zz_strnp_62 ( i_bimc_rxrsp1[31:0], 
	bimc_rxrsp1_data_din[31:0]);
ixc_assign_8 _zz_strnp_63 ( i_bimc_rxrsp2[7:0], bimc_rxrsp2_data_din[7:0]);
ixc_assign _zz_strnp_64 ( i_bimc_rxrsp2[8], bimc_rxrsp2_rxflag_din);
ixc_assign _zz_strnp_65 ( i_bimc_rxrsp2[9], o_bimc_rxrsp2[9]);
ixc_assign_32 _zz_strnp_66 ( i_bimc_pollrsp0[31:0], 
	bimc_pollrsp0_data_din[31:0]);
ixc_assign_32 _zz_strnp_67 ( i_bimc_pollrsp1[31:0], 
	bimc_pollrsp1_data_din[31:0]);
ixc_assign_8 _zz_strnp_68 ( i_bimc_pollrsp2[7:0], bimc_pollrsp2_data_din[7:0]);
ixc_assign _zz_strnp_69 ( i_bimc_pollrsp2[8], bimc_pollrsp2_rxflag_din);
ixc_assign _zz_strnp_70 ( i_bimc_pollrsp2[9], o_bimc_pollrsp2[9]);
ixc_assign _zz_strnp_71 ( _zy_simnet_bimc_ecc_error_0_w$, bimc_ecc_error);
ixc_assign _zz_strnp_72 ( _zy_simnet_bimc_interrupt_1_w$, bimc_interrupt);
ixc_assign _zz_strnp_73 ( _zy_simnet_bimc_odat_2_w$, bimc_odat);
ixc_assign _zz_strnp_74 ( _zy_simnet_bimc_osync_3_w$, bimc_osync);
ixc_assign _zz_strnp_75 ( _zy_simnet_bimc_rst_n_4_w$, bimc_rst_n);
Q_OR03 U1902 ( .A0(i_bimc_monitor[6]), .A1(i_bimc_monitor[5]), .A2(i_bimc_monitor[4]), .Z(n1315));
Q_OR03 U1903 ( .A0(i_bimc_monitor[2]), .A1(i_bimc_monitor[1]), .A2(i_bimc_monitor[0]), .Z(n1314));
Q_OR02 U1904 ( .A0(n1315), .A1(n1314), .Z(bimc_interrupt_c));
Q_XOR2 U1905 ( .A0(tstate[3]), .A1(n1212), .Z(n1210));
Q_FDP4EP \bimc_dat_REG[71] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[71]), .Q(bimc_dat[71]));
Q_INV U1907 ( .A(rst_n), .Z(n1319));
Q_FDP4EP \bimc_dat_REG[70] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[70]), .Q(bimc_dat[70]));
Q_FDP4EP \bimc_dat_REG[69] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[69]), .Q(bimc_dat[69]));
Q_FDP4EP \bimc_dat_REG[68] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[68]), .Q(bimc_dat[68]));
Q_FDP4EP \bimc_dat_REG[67] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[67]), .Q(bimc_dat[67]));
Q_FDP4EP \bimc_dat_REG[66] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[66]), .Q(bimc_dat[66]));
Q_FDP4EP \bimc_dat_REG[65] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[65]), .Q(bimc_dat[65]));
Q_FDP4EP \bimc_dat_REG[64] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[64]), .Q(bimc_dat[64]));
Q_FDP4EP \bimc_dat_REG[63] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[63]), .Q(bimc_dat[63]));
Q_FDP4EP \bimc_dat_REG[62] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[62]), .Q(bimc_dat[62]));
Q_FDP4EP \bimc_dat_REG[61] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[61]), .Q(bimc_dat[61]));
Q_FDP4EP \bimc_dat_REG[60] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[60]), .Q(bimc_dat[60]));
Q_FDP4EP \bimc_dat_REG[59] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[59]), .Q(bimc_dat[59]));
Q_FDP4EP \bimc_dat_REG[58] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[58]), .Q(bimc_dat[58]));
Q_FDP4EP \bimc_dat_REG[57] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[57]), .Q(bimc_dat[57]));
Q_FDP4EP \bimc_dat_REG[56] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[56]), .Q(bimc_dat[56]));
Q_FDP4EP \bimc_dat_REG[55] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[55]), .Q(bimc_dat[55]));
Q_FDP4EP \bimc_dat_REG[54] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[54]), .Q(bimc_dat[54]));
Q_FDP4EP \bimc_dat_REG[53] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[53]), .Q(bimc_dat[53]));
Q_FDP4EP \bimc_dat_REG[52] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[52]), .Q(bimc_dat[52]));
Q_FDP4EP \bimc_dat_REG[51] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[51]), .Q(bimc_dat[51]));
Q_FDP4EP \bimc_dat_REG[50] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[50]), .Q(bimc_dat[50]));
Q_FDP4EP \bimc_dat_REG[49] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[49]), .Q(bimc_dat[49]));
Q_FDP4EP \bimc_dat_REG[48] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[48]), .Q(bimc_dat[48]));
Q_FDP4EP \bimc_dat_REG[47] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[47]), .Q(bimc_dat[47]));
Q_FDP4EP \bimc_dat_REG[46] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[46]), .Q(bimc_dat[46]));
Q_FDP4EP \bimc_dat_REG[45] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[45]), .Q(bimc_dat[45]));
Q_FDP4EP \bimc_dat_REG[44] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[44]), .Q(bimc_dat[44]));
Q_FDP4EP \bimc_dat_REG[43] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[43]), .Q(bimc_dat[43]));
Q_FDP4EP \bimc_dat_REG[42] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[42]), .Q(bimc_dat[42]));
Q_FDP4EP \bimc_dat_REG[41] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[41]), .Q(bimc_dat[41]));
Q_FDP4EP \bimc_dat_REG[40] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[40]), .Q(bimc_dat[40]));
Q_FDP4EP \bimc_dat_REG[39] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[39]), .Q(bimc_dat[39]));
Q_FDP4EP \bimc_dat_REG[38] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[38]), .Q(bimc_dat[38]));
Q_FDP4EP \bimc_dat_REG[37] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[37]), .Q(bimc_dat[37]));
Q_FDP4EP \bimc_dat_REG[36] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[36]), .Q(bimc_dat[36]));
Q_FDP4EP \bimc_dat_REG[35] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[35]), .Q(bimc_dat[35]));
Q_FDP4EP \bimc_dat_REG[34] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[34]), .Q(bimc_dat[34]));
Q_FDP4EP \bimc_dat_REG[33] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[33]), .Q(bimc_dat[33]));
Q_FDP4EP \bimc_dat_REG[32] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[32]), .Q(bimc_dat[32]));
Q_FDP4EP \bimc_dat_REG[31] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[31]), .Q(bimc_dat[31]));
Q_FDP4EP \bimc_dat_REG[30] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[30]), .Q(bimc_dat[30]));
Q_FDP4EP \bimc_dat_REG[29] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[29]), .Q(bimc_dat[29]));
Q_FDP4EP \bimc_dat_REG[28] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[28]), .Q(bimc_dat[28]));
Q_FDP4EP \bimc_dat_REG[27] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[27]), .Q(bimc_dat[27]));
Q_FDP4EP \bimc_dat_REG[26] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[26]), .Q(bimc_dat[26]));
Q_FDP4EP \bimc_dat_REG[25] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[25]), .Q(bimc_dat[25]));
Q_FDP4EP \bimc_dat_REG[24] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[24]), .Q(bimc_dat[24]));
Q_FDP4EP \bimc_dat_REG[23] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[23]), .Q(bimc_dat[23]));
Q_FDP4EP \bimc_dat_REG[22] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[22]), .Q(bimc_dat[22]));
Q_FDP4EP \bimc_dat_REG[21] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[21]), .Q(bimc_dat[21]));
Q_FDP4EP \bimc_dat_REG[20] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[20]), .Q(bimc_dat[20]));
Q_FDP4EP \bimc_dat_REG[19] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[19]), .Q(bimc_dat[19]));
Q_FDP4EP \bimc_dat_REG[18] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[18]), .Q(bimc_dat[18]));
Q_FDP4EP \bimc_dat_REG[17] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[17]), .Q(bimc_dat[17]));
Q_FDP4EP \bimc_dat_REG[16] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[16]), .Q(bimc_dat[16]));
Q_FDP4EP \bimc_dat_REG[15] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[15]), .Q(bimc_dat[15]));
Q_FDP4EP \bimc_dat_REG[14] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[14]), .Q(bimc_dat[14]));
Q_FDP4EP \bimc_dat_REG[13] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[13]), .Q(bimc_dat[13]));
Q_FDP4EP \bimc_dat_REG[12] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[12]), .Q(bimc_dat[12]));
Q_FDP4EP \bimc_dat_REG[11] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[11]), .Q(bimc_dat[11]));
Q_FDP4EP \bimc_dat_REG[10] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[10]), .Q(bimc_dat[10]));
Q_FDP4EP \bimc_dat_REG[9] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[9]), .Q(bimc_dat[9]));
Q_FDP4EP \bimc_dat_REG[8] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[8]), .Q(bimc_dat[8]));
Q_FDP4EP \bimc_dat_REG[7] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[7]), .Q(bimc_dat[7]));
Q_FDP4EP \bimc_dat_REG[6] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[6]), .Q(bimc_dat[6]));
Q_FDP4EP \bimc_dat_REG[5] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[5]), .Q(bimc_dat[5]));
Q_FDP4EP \bimc_dat_REG[4] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[4]), .Q(bimc_dat[4]));
Q_FDP4EP \bimc_dat_REG[3] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[3]), .Q(bimc_dat[3]));
Q_FDP4EP \bimc_dat_REG[2] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[2]), .Q(bimc_dat[2]));
Q_FDP4EP \bimc_dat_REG[1] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[1]), .Q(bimc_dat[1]));
Q_FDP4EP \bimc_dat_REG[0] ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_rdat[0]), .Q(bimc_dat[0]));
Q_FDP4EP bm_resp_REG  ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(bimc_idat), .Q(bm_resp));
Q_FDP4EP bimc_frm_REG  ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(n1189), .Q(bimc_frm));
Q_INV U1981 ( .A(bimc_chk), .Z(n1320));
Q_FDP4EP bimc_chk_REG  ( .CK(clk), .CE(bimc_isync), .R(n1319), .D(n1320), .Q(bimc_chk));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[31] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[31]), .Q(bimc_rxrsp0_data_din[31]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[30] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[30]), .Q(bimc_rxrsp0_data_din[30]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[29] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[29]), .Q(bimc_rxrsp0_data_din[29]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[28] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[28]), .Q(bimc_rxrsp0_data_din[28]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[27] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[27]), .Q(bimc_rxrsp0_data_din[27]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[26] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[26]), .Q(bimc_rxrsp0_data_din[26]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[25] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[25]), .Q(bimc_rxrsp0_data_din[25]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[24] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[24]), .Q(bimc_rxrsp0_data_din[24]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[23] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[23]), .Q(bimc_rxrsp0_data_din[23]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[22] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[22]), .Q(bimc_rxrsp0_data_din[22]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[21] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[21]), .Q(bimc_rxrsp0_data_din[21]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[20] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[20]), .Q(bimc_rxrsp0_data_din[20]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[19] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[19]), .Q(bimc_rxrsp0_data_din[19]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[18] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[18]), .Q(bimc_rxrsp0_data_din[18]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[17] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[17]), .Q(bimc_rxrsp0_data_din[17]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[16] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[16]), .Q(bimc_rxrsp0_data_din[16]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[15] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[15]), .Q(bimc_rxrsp0_data_din[15]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[14] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[14]), .Q(bimc_rxrsp0_data_din[14]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[13] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[13]), .Q(bimc_rxrsp0_data_din[13]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[12] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[12]), .Q(bimc_rxrsp0_data_din[12]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[11] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[11]), .Q(bimc_rxrsp0_data_din[11]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[10] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[10]), .Q(bimc_rxrsp0_data_din[10]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[9] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[9]), .Q(bimc_rxrsp0_data_din[9]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[8] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[8]), .Q(bimc_rxrsp0_data_din[8]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[7] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[7]), .Q(bimc_rxrsp0_data_din[7]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[6] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[6]), .Q(bimc_rxrsp0_data_din[6]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[5] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[5]), .Q(bimc_rxrsp0_data_din[5]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[4] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[4]), .Q(bimc_rxrsp0_data_din[4]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[3] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[3]), .Q(bimc_rxrsp0_data_din[3]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[2] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[2]), .Q(bimc_rxrsp0_data_din[2]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[1] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[1]), .Q(bimc_rxrsp0_data_din[1]));
Q_FDP4EP \bimc_rxrsp0_data_din_REG[0] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_dat[0]), .Q(bimc_rxrsp0_data_din[0]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[7] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[7]), .Q(bimc_rxrsp2_data_din[7]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[6] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[6]), .Q(bimc_rxrsp2_data_din[6]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[5] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[5]), .Q(bimc_rxrsp2_data_din[5]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[4] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[4]), .Q(bimc_rxrsp2_data_din[4]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[3] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[3]), .Q(bimc_rxrsp2_data_din[3]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[2] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[2]), .Q(bimc_rxrsp2_data_din[2]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[1] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[1]), .Q(bimc_rxrsp2_data_din[1]));
Q_FDP4EP \bimc_rxrsp2_data_din_REG[0] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_op[0]), .Q(bimc_rxrsp2_data_din[0]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[31] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[31]), .Q(bimc_pollrsp0_data_din[31]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[30] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[30]), .Q(bimc_pollrsp0_data_din[30]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[29] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[29]), .Q(bimc_pollrsp0_data_din[29]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[28] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[28]), .Q(bimc_pollrsp0_data_din[28]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[27] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[27]), .Q(bimc_pollrsp0_data_din[27]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[26] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[26]), .Q(bimc_pollrsp0_data_din[26]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[25] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[25]), .Q(bimc_pollrsp0_data_din[25]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[24] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[24]), .Q(bimc_pollrsp0_data_din[24]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[23] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[23]), .Q(bimc_pollrsp0_data_din[23]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[22] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[22]), .Q(bimc_pollrsp0_data_din[22]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[21] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[21]), .Q(bimc_pollrsp0_data_din[21]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[20] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[20]), .Q(bimc_pollrsp0_data_din[20]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[19] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[19]), .Q(bimc_pollrsp0_data_din[19]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[18] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[18]), .Q(bimc_pollrsp0_data_din[18]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[17] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[17]), .Q(bimc_pollrsp0_data_din[17]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[16] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[16]), .Q(bimc_pollrsp0_data_din[16]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[15] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[15]), .Q(bimc_pollrsp0_data_din[15]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[14] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[14]), .Q(bimc_pollrsp0_data_din[14]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[13] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[13]), .Q(bimc_pollrsp0_data_din[13]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[12] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[12]), .Q(bimc_pollrsp0_data_din[12]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[11] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[11]), .Q(bimc_pollrsp0_data_din[11]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[10] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[10]), .Q(bimc_pollrsp0_data_din[10]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[9] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[9]), .Q(bimc_pollrsp0_data_din[9]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[8] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[8]), .Q(bimc_pollrsp0_data_din[8]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[7] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[7]), .Q(bimc_pollrsp0_data_din[7]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[6] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[6]), .Q(bimc_pollrsp0_data_din[6]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[5] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[5]), .Q(bimc_pollrsp0_data_din[5]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[4] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[4]), .Q(bimc_pollrsp0_data_din[4]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[3] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[3]), .Q(bimc_pollrsp0_data_din[3]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[2] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[2]), .Q(bimc_pollrsp0_data_din[2]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[1] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[1]), .Q(bimc_pollrsp0_data_din[1]));
Q_FDP4EP \bimc_pollrsp0_data_din_REG[0] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_dat[0]), .Q(bimc_pollrsp0_data_din[0]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[7] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[7]), .Q(bimc_pollrsp2_data_din[7]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[6] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[6]), .Q(bimc_pollrsp2_data_din[6]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[5] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[5]), .Q(bimc_pollrsp2_data_din[5]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[4] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[4]), .Q(bimc_pollrsp2_data_din[4]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[3] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[3]), .Q(bimc_pollrsp2_data_din[3]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[2] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[2]), .Q(bimc_pollrsp2_data_din[2]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[1] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[1]), .Q(bimc_pollrsp2_data_din[1]));
Q_FDP4EP \bimc_pollrsp2_data_din_REG[0] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_op[0]), .Q(bimc_pollrsp2_data_din[0]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[31] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[31]), .Q(bimc_rxcmd0_data_din[31]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[30] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[30]), .Q(bimc_rxcmd0_data_din[30]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[29] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[29]), .Q(bimc_rxcmd0_data_din[29]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[28] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[28]), .Q(bimc_rxcmd0_data_din[28]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[27] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[27]), .Q(bimc_rxcmd0_data_din[27]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[26] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[26]), .Q(bimc_rxcmd0_data_din[26]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[25] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[25]), .Q(bimc_rxcmd0_data_din[25]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[24] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[24]), .Q(bimc_rxcmd0_data_din[24]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[23] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[23]), .Q(bimc_rxcmd0_data_din[23]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[22] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[22]), .Q(bimc_rxcmd0_data_din[22]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[21] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[21]), .Q(bimc_rxcmd0_data_din[21]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[20] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[20]), .Q(bimc_rxcmd0_data_din[20]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[19] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[19]), .Q(bimc_rxcmd0_data_din[19]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[18] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[18]), .Q(bimc_rxcmd0_data_din[18]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[17] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[17]), .Q(bimc_rxcmd0_data_din[17]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[16] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[16]), .Q(bimc_rxcmd0_data_din[16]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[15] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[15]), .Q(bimc_rxcmd0_data_din[15]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[14] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[14]), .Q(bimc_rxcmd0_data_din[14]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[13] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[13]), .Q(bimc_rxcmd0_data_din[13]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[12] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[12]), .Q(bimc_rxcmd0_data_din[12]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[11] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[11]), .Q(bimc_rxcmd0_data_din[11]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[10] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[10]), .Q(bimc_rxcmd0_data_din[10]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[9] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[9]), .Q(bimc_rxcmd0_data_din[9]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[8] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[8]), .Q(bimc_rxcmd0_data_din[8]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[7] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[7]), .Q(bimc_rxcmd0_data_din[7]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[6] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[6]), .Q(bimc_rxcmd0_data_din[6]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[5] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[5]), .Q(bimc_rxcmd0_data_din[5]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[4] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[4]), .Q(bimc_rxcmd0_data_din[4]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[3] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[3]), .Q(bimc_rxcmd0_data_din[3]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[2] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[2]), .Q(bimc_rxcmd0_data_din[2]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[1] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[1]), .Q(bimc_rxcmd0_data_din[1]));
Q_FDP4EP \bimc_rxcmd0_data_din_REG[0] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_dat[0]), .Q(bimc_rxcmd0_data_din[0]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[15] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[15]), .Q(bimc_rxcmd1_addr_din[15]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[14] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[14]), .Q(bimc_rxcmd1_addr_din[14]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[13] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[13]), .Q(bimc_rxcmd1_addr_din[13]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[12] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[12]), .Q(bimc_rxcmd1_addr_din[12]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[11] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[11]), .Q(bimc_rxcmd1_addr_din[11]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[10] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[10]), .Q(bimc_rxcmd1_addr_din[10]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[9] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[9]), .Q(bimc_rxcmd1_addr_din[9]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[8] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[8]), .Q(bimc_rxcmd1_addr_din[8]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[7] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[7]), .Q(bimc_rxcmd1_addr_din[7]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[6] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[6]), .Q(bimc_rxcmd1_addr_din[6]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[5] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[5]), .Q(bimc_rxcmd1_addr_din[5]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[4] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[4]), .Q(bimc_rxcmd1_addr_din[4]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[3] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[3]), .Q(bimc_rxcmd1_addr_din[3]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[2] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[2]), .Q(bimc_rxcmd1_addr_din[2]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[1] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[1]), .Q(bimc_rxcmd1_addr_din[1]));
Q_FDP4EP \bimc_rxcmd1_addr_din_REG[0] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_addr[0]), .Q(bimc_rxcmd1_addr_din[0]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[11] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[11]), .Q(bimc_rxcmd1_mem_din[11]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[10] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[10]), .Q(bimc_rxcmd1_mem_din[10]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[9] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[9]), .Q(bimc_rxcmd1_mem_din[9]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[8] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[8]), .Q(bimc_rxcmd1_mem_din[8]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[7] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[7]), .Q(bimc_rxcmd1_mem_din[7]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[6] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[6]), .Q(bimc_rxcmd1_mem_din[6]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[5] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[5]), .Q(bimc_rxcmd1_mem_din[5]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[4] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[4]), .Q(bimc_rxcmd1_mem_din[4]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[3] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[3]), .Q(bimc_rxcmd1_mem_din[3]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[2] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[2]), .Q(bimc_rxcmd1_mem_din[2]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[1] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[1]), .Q(bimc_rxcmd1_mem_din[1]));
Q_FDP4EP \bimc_rxcmd1_mem_din_REG[0] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_mem[0]), .Q(bimc_rxcmd1_mem_din[0]));
Q_FDP4EP \bimc_rxcmd1_memtype_din_REG[3] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_type[3]), .Q(bimc_rxcmd1_memtype_din[3]));
Q_FDP4EP \bimc_rxcmd1_memtype_din_REG[2] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_type[2]), .Q(bimc_rxcmd1_memtype_din[2]));
Q_FDP4EP \bimc_rxcmd1_memtype_din_REG[1] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_type[1]), .Q(bimc_rxcmd1_memtype_din[1]));
Q_FDP4EP \bimc_rxcmd1_memtype_din_REG[0] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_type[0]), .Q(bimc_rxcmd1_memtype_din[0]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[7] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[7]), .Q(bimc_rxcmd2_opcode_din[7]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[6] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[6]), .Q(bimc_rxcmd2_opcode_din[6]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[5] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[5]), .Q(bimc_rxcmd2_opcode_din[5]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[4] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[4]), .Q(bimc_rxcmd2_opcode_din[4]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[3] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[3]), .Q(bimc_rxcmd2_opcode_din[3]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[2] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[2]), .Q(bimc_rxcmd2_opcode_din[2]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[1] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[1]), .Q(bimc_rxcmd2_opcode_din[1]));
Q_FDP4EP \bimc_rxcmd2_opcode_din_REG[0] ( .CK(clk), .CE(n1043), .R(n1319), .D(rx_op[0]), .Q(bimc_rxcmd2_opcode_din[0]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[31] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[31]), .Q(bimc_dbgcmd0_data_din[31]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[30] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[30]), .Q(bimc_dbgcmd0_data_din[30]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[29] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[29]), .Q(bimc_dbgcmd0_data_din[29]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[28] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[28]), .Q(bimc_dbgcmd0_data_din[28]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[27] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[27]), .Q(bimc_dbgcmd0_data_din[27]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[26] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[26]), .Q(bimc_dbgcmd0_data_din[26]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[25] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[25]), .Q(bimc_dbgcmd0_data_din[25]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[24] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[24]), .Q(bimc_dbgcmd0_data_din[24]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[23] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[23]), .Q(bimc_dbgcmd0_data_din[23]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[22] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[22]), .Q(bimc_dbgcmd0_data_din[22]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[21] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[21]), .Q(bimc_dbgcmd0_data_din[21]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[20] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[20]), .Q(bimc_dbgcmd0_data_din[20]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[19] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[19]), .Q(bimc_dbgcmd0_data_din[19]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[18] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[18]), .Q(bimc_dbgcmd0_data_din[18]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[17] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[17]), .Q(bimc_dbgcmd0_data_din[17]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[16] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[16]), .Q(bimc_dbgcmd0_data_din[16]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[15] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[15]), .Q(bimc_dbgcmd0_data_din[15]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[14] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[14]), .Q(bimc_dbgcmd0_data_din[14]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[13] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[13]), .Q(bimc_dbgcmd0_data_din[13]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[12] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[12]), .Q(bimc_dbgcmd0_data_din[12]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[11] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[11]), .Q(bimc_dbgcmd0_data_din[11]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[10] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[10]), .Q(bimc_dbgcmd0_data_din[10]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[9] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[9]), .Q(bimc_dbgcmd0_data_din[9]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[8] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[8]), .Q(bimc_dbgcmd0_data_din[8]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[7] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[7]), .Q(bimc_dbgcmd0_data_din[7]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[6] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[6]), .Q(bimc_dbgcmd0_data_din[6]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[5] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[5]), .Q(bimc_dbgcmd0_data_din[5]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[4] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[4]), .Q(bimc_dbgcmd0_data_din[4]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[3] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[3]), .Q(bimc_dbgcmd0_data_din[3]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[2] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[2]), .Q(bimc_dbgcmd0_data_din[2]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[1] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[1]), .Q(bimc_dbgcmd0_data_din[1]));
Q_FDP4EP \bimc_dbgcmd0_data_din_REG[0] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_dat[0]), .Q(bimc_dbgcmd0_data_din[0]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[15] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[15]), .Q(bimc_dbgcmd1_addr_din[15]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[14] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[14]), .Q(bimc_dbgcmd1_addr_din[14]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[13] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[13]), .Q(bimc_dbgcmd1_addr_din[13]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[12] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[12]), .Q(bimc_dbgcmd1_addr_din[12]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[11] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[11]), .Q(bimc_dbgcmd1_addr_din[11]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[10] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[10]), .Q(bimc_dbgcmd1_addr_din[10]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[9] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[9]), .Q(bimc_dbgcmd1_addr_din[9]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[8] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[8]), .Q(bimc_dbgcmd1_addr_din[8]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[7] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[7]), .Q(bimc_dbgcmd1_addr_din[7]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[6] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[6]), .Q(bimc_dbgcmd1_addr_din[6]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[5] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[5]), .Q(bimc_dbgcmd1_addr_din[5]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[4] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[4]), .Q(bimc_dbgcmd1_addr_din[4]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[3] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[3]), .Q(bimc_dbgcmd1_addr_din[3]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[2] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[2]), .Q(bimc_dbgcmd1_addr_din[2]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[1] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[1]), .Q(bimc_dbgcmd1_addr_din[1]));
Q_FDP4EP \bimc_dbgcmd1_addr_din_REG[0] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_addr[0]), .Q(bimc_dbgcmd1_addr_din[0]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[11] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[11]), .Q(bimc_dbgcmd1_mem_din[11]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[10] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[10]), .Q(bimc_dbgcmd1_mem_din[10]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[9] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[9]), .Q(bimc_dbgcmd1_mem_din[9]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[8] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[8]), .Q(bimc_dbgcmd1_mem_din[8]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[7] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[7]), .Q(bimc_dbgcmd1_mem_din[7]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[6] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[6]), .Q(bimc_dbgcmd1_mem_din[6]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[5] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[5]), .Q(bimc_dbgcmd1_mem_din[5]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[4] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[4]), .Q(bimc_dbgcmd1_mem_din[4]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[3] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[3]), .Q(bimc_dbgcmd1_mem_din[3]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[2] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[2]), .Q(bimc_dbgcmd1_mem_din[2]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[1] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[1]), .Q(bimc_dbgcmd1_mem_din[1]));
Q_FDP4EP \bimc_dbgcmd1_mem_din_REG[0] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_mem[0]), .Q(bimc_dbgcmd1_mem_din[0]));
Q_FDP4EP \bimc_dbgcmd1_memtype_din_REG[3] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_type[3]), .Q(bimc_dbgcmd1_memtype_din[3]));
Q_FDP4EP \bimc_dbgcmd1_memtype_din_REG[2] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_type[2]), .Q(bimc_dbgcmd1_memtype_din[2]));
Q_FDP4EP \bimc_dbgcmd1_memtype_din_REG[1] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_type[1]), .Q(bimc_dbgcmd1_memtype_din[1]));
Q_FDP4EP \bimc_dbgcmd1_memtype_din_REG[0] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_type[0]), .Q(bimc_dbgcmd1_memtype_din[0]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[7] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[7]), .Q(bimc_dbgcmd2_opcode_din[7]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[6] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[6]), .Q(bimc_dbgcmd2_opcode_din[6]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[5] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[5]), .Q(bimc_dbgcmd2_opcode_din[5]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[4] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[4]), .Q(bimc_dbgcmd2_opcode_din[4]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[3] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[3]), .Q(bimc_dbgcmd2_opcode_din[3]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[2] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[2]), .Q(bimc_dbgcmd2_opcode_din[2]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[1] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[1]), .Q(bimc_dbgcmd2_opcode_din[1]));
Q_FDP4EP \bimc_dbgcmd2_opcode_din_REG[0] ( .CK(clk), .CE(n1039), .R(n1319), .D(rx_op[0]), .Q(bimc_dbgcmd2_opcode_din[0]));
Q_FDP4EP \number_of_memories_REG[11] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1064), .Q(number_of_memories[11]));
Q_FDP4EP \number_of_memories_REG[10] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1066), .Q(number_of_memories[10]));
Q_FDP4EP \number_of_memories_REG[9] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1068), .Q(number_of_memories[9]));
Q_FDP4EP \number_of_memories_REG[8] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1070), .Q(number_of_memories[8]));
Q_FDP4EP \number_of_memories_REG[7] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1072), .Q(number_of_memories[7]));
Q_FDP4EP \number_of_memories_REG[6] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1074), .Q(number_of_memories[6]));
Q_FDP4EP \number_of_memories_REG[5] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1076), .Q(number_of_memories[5]));
Q_FDP4EP \number_of_memories_REG[4] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1078), .Q(number_of_memories[4]));
Q_FDP4EP \number_of_memories_REG[3] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1080), .Q(number_of_memories[3]));
Q_FDP4EP \number_of_memories_REG[2] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1082), .Q(number_of_memories[2]));
Q_FDP4EP \number_of_memories_REG[1] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1084), .Q(number_of_memories[1]));
Q_FDP4EP \number_of_memories_REG[0] ( .CK(clk), .CE(n1019), .R(n1319), .D(n1085), .Q(number_of_memories[0]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[31] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_type[3]), .Q(bimc_rxrsp1_data_din[31]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[30] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_type[2]), .Q(bimc_rxrsp1_data_din[30]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[29] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_type[1]), .Q(bimc_rxrsp1_data_din[29]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[28] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_type[0]), .Q(bimc_rxrsp1_data_din[28]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[27] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[11]), .Q(bimc_rxrsp1_data_din[27]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[26] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[10]), .Q(bimc_rxrsp1_data_din[26]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[25] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[9]), .Q(bimc_rxrsp1_data_din[25]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[24] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[8]), .Q(bimc_rxrsp1_data_din[24]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[23] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[7]), .Q(bimc_rxrsp1_data_din[23]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[22] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[6]), .Q(bimc_rxrsp1_data_din[22]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[21] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[5]), .Q(bimc_rxrsp1_data_din[21]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[20] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[4]), .Q(bimc_rxrsp1_data_din[20]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[19] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[3]), .Q(bimc_rxrsp1_data_din[19]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[18] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[2]), .Q(bimc_rxrsp1_data_din[18]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[17] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[1]), .Q(bimc_rxrsp1_data_din[17]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[16] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_mem[0]), .Q(bimc_rxrsp1_data_din[16]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[15] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[15]), .Q(bimc_rxrsp1_data_din[15]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[14] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[14]), .Q(bimc_rxrsp1_data_din[14]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[13] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[13]), .Q(bimc_rxrsp1_data_din[13]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[12] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[12]), .Q(bimc_rxrsp1_data_din[12]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[11] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[11]), .Q(bimc_rxrsp1_data_din[11]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[10] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[10]), .Q(bimc_rxrsp1_data_din[10]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[9] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[9]), .Q(bimc_rxrsp1_data_din[9]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[8] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[8]), .Q(bimc_rxrsp1_data_din[8]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[7] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[7]), .Q(bimc_rxrsp1_data_din[7]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[6] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[6]), .Q(bimc_rxrsp1_data_din[6]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[5] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[5]), .Q(bimc_rxrsp1_data_din[5]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[4] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[4]), .Q(bimc_rxrsp1_data_din[4]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[3] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[3]), .Q(bimc_rxrsp1_data_din[3]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[2] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[2]), .Q(bimc_rxrsp1_data_din[2]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[1] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[1]), .Q(bimc_rxrsp1_data_din[1]));
Q_FDP4EP \bimc_rxrsp1_data_din_REG[0] ( .CK(clk), .CE(n1050), .R(n1319), .D(rx_addr[0]), .Q(bimc_rxrsp1_data_din[0]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[31] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_type[3]), .Q(bimc_pollrsp1_data_din[31]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[30] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_type[2]), .Q(bimc_pollrsp1_data_din[30]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[29] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_type[1]), .Q(bimc_pollrsp1_data_din[29]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[28] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_type[0]), .Q(bimc_pollrsp1_data_din[28]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[27] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[11]), .Q(bimc_pollrsp1_data_din[27]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[26] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[10]), .Q(bimc_pollrsp1_data_din[26]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[25] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[9]), .Q(bimc_pollrsp1_data_din[25]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[24] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[8]), .Q(bimc_pollrsp1_data_din[24]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[23] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[7]), .Q(bimc_pollrsp1_data_din[23]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[22] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[6]), .Q(bimc_pollrsp1_data_din[22]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[21] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[5]), .Q(bimc_pollrsp1_data_din[21]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[20] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[4]), .Q(bimc_pollrsp1_data_din[20]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[19] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[3]), .Q(bimc_pollrsp1_data_din[19]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[18] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[2]), .Q(bimc_pollrsp1_data_din[18]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[17] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[1]), .Q(bimc_pollrsp1_data_din[17]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[16] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_mem[0]), .Q(bimc_pollrsp1_data_din[16]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[15] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[15]), .Q(bimc_pollrsp1_data_din[15]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[14] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[14]), .Q(bimc_pollrsp1_data_din[14]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[13] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[13]), .Q(bimc_pollrsp1_data_din[13]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[12] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[12]), .Q(bimc_pollrsp1_data_din[12]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[11] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[11]), .Q(bimc_pollrsp1_data_din[11]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[10] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[10]), .Q(bimc_pollrsp1_data_din[10]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[9] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[9]), .Q(bimc_pollrsp1_data_din[9]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[8] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[8]), .Q(bimc_pollrsp1_data_din[8]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[7] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[7]), .Q(bimc_pollrsp1_data_din[7]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[6] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[6]), .Q(bimc_pollrsp1_data_din[6]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[5] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[5]), .Q(bimc_pollrsp1_data_din[5]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[4] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[4]), .Q(bimc_pollrsp1_data_din[4]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[3] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[3]), .Q(bimc_pollrsp1_data_din[3]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[2] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[2]), .Q(bimc_pollrsp1_data_din[2]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[1] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[1]), .Q(bimc_pollrsp1_data_din[1]));
Q_FDP4EP \bimc_pollrsp1_data_din_REG[0] ( .CK(clk), .CE(n1045), .R(n1319), .D(rx_addr[0]), .Q(bimc_pollrsp1_data_din[0]));
Q_FDP4EP bimc_monitor_uncorrectable_ecc_error_din_REG  ( .CK(clk), .CE(n1025), .R(n1319), .D(n1026), .Q(bimc_monitor_uncorrectable_ecc_error_din));
Q_FDP4EP bimc_monitor_correctable_ecc_error_din_REG  ( .CK(clk), .CE(n1024), .R(n1319), .D(n1027), .Q(bimc_monitor_correctable_ecc_error_din));
Q_FDP4EP bimc_monitor_parity_error_din_REG  ( .CK(clk), .CE(n1023), .R(n1319), .D(n1028), .Q(bimc_monitor_parity_error_din));
Q_FDP4EP bimc_monitor_bimc_chain_rcv_error_din_REG  ( .CK(clk), .CE(n1022), .R(n1319), .D(n1029), .Q(bimc_monitor_bimc_chain_rcv_error_din));
Q_FDP4EP bimc_monitor_rcv_invalid_opcode_din_REG  ( .CK(clk), .CE(n1021), .R(n1319), .D(n1030), .Q(bimc_monitor_rcv_invalid_opcode_din));
Q_FDP4EP bimc_monitor_unanswered_read_din_REG  ( .CK(clk), .CE(n1020), .R(n1319), .D(n1031), .Q(bimc_monitor_unanswered_read_din));
Q_FDP4EP bimc_rxrsp2_rxflag_din_REG  ( .CK(clk), .CE(n1018), .R(n1319), .D(n1032), .Q(bimc_rxrsp2_rxflag_din));
Q_FDP4EP bimc_pollrsp2_rxflag_din_REG  ( .CK(clk), .CE(n1017), .R(n1319), .D(n1033), .Q(bimc_pollrsp2_rxflag_din));
Q_FDP4EP bimc_rxcmd2_rxflag_din_REG  ( .CK(clk), .CE(n1016), .R(n1319), .D(n1034), .Q(bimc_rxcmd2_rxflag_din));
Q_FDP4EP bimc_dbgcmd2_rxflag_din_REG  ( .CK(clk), .CE(n1015), .R(n1319), .D(n1035), .Q(bimc_dbgcmd2_rxflag_din));
Q_FDP4EP bimc_global_config_bimc_mem_init_done_din_REG  ( .CK(clk), .CE(n1014), .R(n1319), .D(n1164), .Q(bimc_global_config_bimc_mem_init_done_din));
Q_FDP4EP \cputx_type_REG[3] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_memtype[3]), .Q(cputx_type[3]));
Q_FDP4EP \cputx_type_REG[2] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_memtype[2]), .Q(cputx_type[2]));
Q_FDP4EP \cputx_type_REG[1] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_memtype[1]), .Q(cputx_type[1]));
Q_FDP4EP \cputx_type_REG[0] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_memtype[0]), .Q(cputx_type[0]));
Q_FDP4EP \cputx_op_REG[7] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[7]), .Q(cputx_op[7]));
Q_FDP4EP \cputx_op_REG[6] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[6]), .Q(cputx_op[6]));
Q_FDP4EP \cputx_op_REG[5] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[5]), .Q(cputx_op[5]));
Q_FDP4EP \cputx_op_REG[4] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[4]), .Q(cputx_op[4]));
Q_FDP4EP \cputx_op_REG[3] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[3]), .Q(cputx_op[3]));
Q_FDP4EP \cputx_op_REG[2] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[2]), .Q(cputx_op[2]));
Q_FDP4EP \cputx_op_REG[1] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[1]), .Q(cputx_op[1]));
Q_FDP4EP \cputx_op_REG[0] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd2_opcode[0]), .Q(cputx_op[0]));
Q_FDP4EP \cputx_mem_REG[11] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[11]), .Q(cputx_mem[11]));
Q_FDP4EP \cputx_mem_REG[10] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[10]), .Q(cputx_mem[10]));
Q_FDP4EP \cputx_mem_REG[9] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[9]), .Q(cputx_mem[9]));
Q_FDP4EP \cputx_mem_REG[8] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[8]), .Q(cputx_mem[8]));
Q_FDP4EP \cputx_mem_REG[7] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[7]), .Q(cputx_mem[7]));
Q_FDP4EP \cputx_mem_REG[6] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[6]), .Q(cputx_mem[6]));
Q_FDP4EP \cputx_mem_REG[5] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[5]), .Q(cputx_mem[5]));
Q_FDP4EP \cputx_mem_REG[4] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[4]), .Q(cputx_mem[4]));
Q_FDP4EP \cputx_mem_REG[3] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[3]), .Q(cputx_mem[3]));
Q_FDP4EP \cputx_mem_REG[2] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[2]), .Q(cputx_mem[2]));
Q_FDP4EP \cputx_mem_REG[1] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[1]), .Q(cputx_mem[1]));
Q_FDP4EP \cputx_mem_REG[0] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_mem[0]), .Q(cputx_mem[0]));
Q_FDP4EP \cputx_addr_REG[15] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[15]), .Q(cputx_addr[15]));
Q_FDP4EP \cputx_addr_REG[14] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[14]), .Q(cputx_addr[14]));
Q_FDP4EP \cputx_addr_REG[13] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[13]), .Q(cputx_addr[13]));
Q_FDP4EP \cputx_addr_REG[12] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[12]), .Q(cputx_addr[12]));
Q_FDP4EP \cputx_addr_REG[11] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[11]), .Q(cputx_addr[11]));
Q_FDP4EP \cputx_addr_REG[10] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[10]), .Q(cputx_addr[10]));
Q_FDP4EP \cputx_addr_REG[9] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[9]), .Q(cputx_addr[9]));
Q_FDP4EP \cputx_addr_REG[8] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[8]), .Q(cputx_addr[8]));
Q_FDP4EP \cputx_addr_REG[7] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[7]), .Q(cputx_addr[7]));
Q_FDP4EP \cputx_addr_REG[6] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[6]), .Q(cputx_addr[6]));
Q_FDP4EP \cputx_addr_REG[5] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[5]), .Q(cputx_addr[5]));
Q_FDP4EP \cputx_addr_REG[4] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[4]), .Q(cputx_addr[4]));
Q_FDP4EP \cputx_addr_REG[3] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[3]), .Q(cputx_addr[3]));
Q_FDP4EP \cputx_addr_REG[2] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[2]), .Q(cputx_addr[2]));
Q_FDP4EP \cputx_addr_REG[1] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[1]), .Q(cputx_addr[1]));
Q_FDP4EP \cputx_addr_REG[0] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd1_addr[0]), .Q(cputx_addr[0]));
Q_FDP4EP \cputx_dat_REG[31] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[31]), .Q(cputx_dat[31]));
Q_FDP4EP \cputx_dat_REG[30] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[30]), .Q(cputx_dat[30]));
Q_FDP4EP \cputx_dat_REG[29] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[29]), .Q(cputx_dat[29]));
Q_FDP4EP \cputx_dat_REG[28] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[28]), .Q(cputx_dat[28]));
Q_FDP4EP \cputx_dat_REG[27] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[27]), .Q(cputx_dat[27]));
Q_FDP4EP \cputx_dat_REG[26] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[26]), .Q(cputx_dat[26]));
Q_FDP4EP \cputx_dat_REG[25] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[25]), .Q(cputx_dat[25]));
Q_FDP4EP \cputx_dat_REG[24] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[24]), .Q(cputx_dat[24]));
Q_FDP4EP \cputx_dat_REG[23] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[23]), .Q(cputx_dat[23]));
Q_FDP4EP \cputx_dat_REG[22] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[22]), .Q(cputx_dat[22]));
Q_FDP4EP \cputx_dat_REG[21] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[21]), .Q(cputx_dat[21]));
Q_FDP4EP \cputx_dat_REG[20] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[20]), .Q(cputx_dat[20]));
Q_FDP4EP \cputx_dat_REG[19] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[19]), .Q(cputx_dat[19]));
Q_FDP4EP \cputx_dat_REG[18] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[18]), .Q(cputx_dat[18]));
Q_FDP4EP \cputx_dat_REG[17] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[17]), .Q(cputx_dat[17]));
Q_FDP4EP \cputx_dat_REG[16] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[16]), .Q(cputx_dat[16]));
Q_FDP4EP \cputx_dat_REG[15] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[15]), .Q(cputx_dat[15]));
Q_FDP4EP \cputx_dat_REG[14] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[14]), .Q(cputx_dat[14]));
Q_FDP4EP \cputx_dat_REG[13] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[13]), .Q(cputx_dat[13]));
Q_FDP4EP \cputx_dat_REG[12] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[12]), .Q(cputx_dat[12]));
Q_FDP4EP \cputx_dat_REG[11] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[11]), .Q(cputx_dat[11]));
Q_FDP4EP \cputx_dat_REG[10] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[10]), .Q(cputx_dat[10]));
Q_FDP4EP \cputx_dat_REG[9] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[9]), .Q(cputx_dat[9]));
Q_FDP4EP \cputx_dat_REG[8] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[8]), .Q(cputx_dat[8]));
Q_FDP4EP \cputx_dat_REG[7] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[7]), .Q(cputx_dat[7]));
Q_FDP4EP \cputx_dat_REG[6] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[6]), .Q(cputx_dat[6]));
Q_FDP4EP \cputx_dat_REG[5] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[5]), .Q(cputx_dat[5]));
Q_FDP4EP \cputx_dat_REG[4] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[4]), .Q(cputx_dat[4]));
Q_FDP4EP \cputx_dat_REG[3] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[3]), .Q(cputx_dat[3]));
Q_FDP4EP \cputx_dat_REG[2] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[2]), .Q(cputx_dat[2]));
Q_FDP4EP \cputx_dat_REG[1] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[1]), .Q(cputx_dat[1]));
Q_FDP4EP \cputx_dat_REG[0] ( .CK(clk), .CE(n19), .R(n1319), .D(bimc_cmd0_data[0]), .Q(cputx_dat[0]));
Q_FDP4EP mem_wr_init_ev_REG  ( .CK(clk), .CE(n16), .R(n1319), .D(n17), .Q(mem_wr_init_ev));
Q_FDP4EP eccpar_debug_ev_REG  ( .CK(clk), .CE(n15), .R(n1319), .D(n18), .Q(eccpar_debug_ev));
Q_INV U2368 ( .A(eccpar_debug_ev), .Z(n752));
Q_FDP4EP cpu_transmit_ev_REG  ( .CK(clk), .CE(n14), .R(n1319), .D(n19), .Q(cpu_transmit_ev));
Q_FDP4EP auto_poll_ecc_par_ev_REG  ( .CK(clk), .CE(n13), .R(n1319), .D(n20), .Q(auto_poll_ecc_par_ev));
Q_INV U2371 ( .A(auto_poll_ecc_par_ev), .Z(n753));
endmodule
