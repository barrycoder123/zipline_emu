architecture module of ixc_sfifo_bind_22_2 is

begin
end module;
