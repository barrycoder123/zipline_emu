
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module IXC_SV_SCG_GFIFO_VXE_64 ( scgGFreq);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output scgGFreq;
wire fclk;
wire GFreq;
wire [19:0] GFcbid;
wire [11:0] GFlen;
wire [511:0] GFidata;
wire GFtsReq;
wire [63:0] timeStampPkt;
`_2_ wire GFtsAdd;
`_2_ wire [11:0] argLen;
`_2_ wire [543:0] xdata;
`_2_ wire [63:0] wrtCnt;
`_2_ wire [63:0] wrtCntD;
`_2_ wire [16:0] ofifoAddr0;
`_2_ wire [16:0] ofifoAddr0N;
`_2_ wire [16:0] ofifoAddr1;
`_2_ wire [16:0] ofifoAddr2;
`_2_ wire [16:0] ofifoAddr3;
`_2_ wire [16:0] ofifoAddr4;
`_2_ wire [16:0] ofifoAddr5;
`_2_ wire [16:0] ofifoAddr6;
`_2_ wire [16:0] ofifoAddr7;
`_2_ wire [16:0] ofifoAddr8;
`_2_ wire [16:0] ofifoAddr1N;
`_2_ wire [16:0] ofifoAddr2N;
`_2_ wire [16:0] ofifoAddr3N;
`_2_ wire [16:0] ofifoAddr4N;
`_2_ wire [16:0] ofifoAddr5N;
`_2_ wire [16:0] ofifoAddr6N;
`_2_ wire [16:0] ofifoAddr7N;
`_2_ wire [16:0] ofifoAddr8N;
`_2_ wire [575:0] ofifoData;
`_2_ wire [575:0] ofifoDataN;
`_2_ wire [5:0] writeLen;
`_2_ wire reqD;
`_2_ wire [4:0] oFill;
`_2_ wire [4:0] oFillN;
`_2_ wire [16:0] ofifoWptr;
`_2_ wire [16:0] ofifoWptrN;
`_2_ wire [9:0] index;
supply0 n3317;
supply1 n3318;
Q_BUF U0 ( .A(n3317), .Z(index[5]));
Q_BUF U1 ( .A(n3317), .Z(index[4]));
Q_BUF U2 ( .A(n3317), .Z(index[3]));
Q_BUF U3 ( .A(n3317), .Z(index[2]));
Q_BUF U4 ( .A(n3317), .Z(index[1]));
Q_BUF U5 ( .A(n3317), .Z(index[0]));
Q_BUF U6 ( .A(n3318), .Z(timeStampPkt[31]));
Q_BUF U7 ( .A(ofifoAddr5N[1]), .Z(ofifoAddr1N[1]));
Q_BUF U8 ( .A(ofifoWptr[16]), .Z(ofifoAddr0N[16]));
Q_BUF U9 ( .A(ofifoWptr[15]), .Z(ofifoAddr0N[15]));
Q_BUF U10 ( .A(ofifoWptr[14]), .Z(ofifoAddr0N[14]));
Q_BUF U11 ( .A(ofifoWptr[13]), .Z(ofifoAddr0N[13]));
Q_BUF U12 ( .A(ofifoWptr[12]), .Z(ofifoAddr0N[12]));
Q_BUF U13 ( .A(ofifoWptr[11]), .Z(ofifoAddr0N[11]));
Q_BUF U14 ( .A(ofifoWptr[10]), .Z(ofifoAddr0N[10]));
Q_BUF U15 ( .A(ofifoWptr[9]), .Z(ofifoAddr0N[9]));
Q_BUF U16 ( .A(ofifoWptr[8]), .Z(ofifoAddr0N[8]));
Q_BUF U17 ( .A(ofifoWptr[7]), .Z(ofifoAddr0N[7]));
Q_BUF U18 ( .A(ofifoWptr[6]), .Z(ofifoAddr0N[6]));
Q_BUF U19 ( .A(ofifoWptr[5]), .Z(ofifoAddr0N[5]));
Q_BUF U20 ( .A(ofifoWptr[4]), .Z(ofifoAddr0N[4]));
Q_BUF U21 ( .A(ofifoWptr[3]), .Z(ofifoAddr0N[3]));
Q_BUF U22 ( .A(ofifoAddr5N[0]), .Z(ofifoAddr7N[0]));
Q_BUF U23 ( .A(ofifoAddr3N[0]), .Z(ofifoAddr5N[0]));
Q_BUF U24 ( .A(ofifoAddr1N[0]), .Z(ofifoAddr3N[0]));
Q_BUF U25 ( .A(ofifoAddr2N[1]), .Z(ofifoAddr6N[1]));
Q_BUF U26 ( .A(ofifoAddr3N[1]), .Z(ofifoAddr7N[1]));
Q_BUF U27 ( .A(ofifoAddr8N[2]), .Z(ofifoAddr0N[2]));
Q_BUF U28 ( .A(ofifoWptr[2]), .Z(ofifoAddr8N[2]));
Q_BUF U29 ( .A(ofifoAddr4N[1]), .Z(ofifoAddr0N[1]));
Q_BUF U30 ( .A(ofifoAddr8N[1]), .Z(ofifoAddr4N[1]));
Q_BUF U31 ( .A(ofifoWptr[1]), .Z(ofifoAddr8N[1]));
Q_BUF U32 ( .A(ofifoAddr2N[0]), .Z(ofifoAddr0N[0]));
Q_BUF U33 ( .A(ofifoAddr4N[0]), .Z(ofifoAddr2N[0]));
Q_BUF U34 ( .A(ofifoAddr6N[0]), .Z(ofifoAddr4N[0]));
Q_BUF U35 ( .A(ofifoAddr8N[0]), .Z(ofifoAddr6N[0]));
Q_BUF U36 ( .A(ofifoWptr[0]), .Z(ofifoAddr8N[0]));
Q_ASSIGN U37 ( .B(xc_top.ixcSimTime[55]), .A(timeStampPkt[63]));
Q_ASSIGN U38 ( .B(xc_top.ixcSimTime[54]), .A(timeStampPkt[62]));
Q_ASSIGN U39 ( .B(xc_top.ixcSimTime[53]), .A(timeStampPkt[61]));
Q_ASSIGN U40 ( .B(xc_top.ixcSimTime[52]), .A(timeStampPkt[60]));
Q_ASSIGN U41 ( .B(xc_top.ixcSimTime[51]), .A(timeStampPkt[59]));
Q_ASSIGN U42 ( .B(xc_top.ixcSimTime[50]), .A(timeStampPkt[58]));
Q_ASSIGN U43 ( .B(xc_top.ixcSimTime[49]), .A(timeStampPkt[57]));
Q_ASSIGN U44 ( .B(xc_top.ixcSimTime[48]), .A(timeStampPkt[56]));
Q_ASSIGN U45 ( .B(xc_top.ixcSimTime[47]), .A(timeStampPkt[55]));
Q_ASSIGN U46 ( .B(xc_top.ixcSimTime[46]), .A(timeStampPkt[54]));
Q_ASSIGN U47 ( .B(xc_top.ixcSimTime[45]), .A(timeStampPkt[53]));
Q_ASSIGN U48 ( .B(xc_top.ixcSimTime[44]), .A(timeStampPkt[52]));
Q_ASSIGN U49 ( .B(xc_top.ixcSimTime[43]), .A(timeStampPkt[51]));
Q_ASSIGN U50 ( .B(xc_top.ixcSimTime[42]), .A(timeStampPkt[50]));
Q_ASSIGN U51 ( .B(xc_top.ixcSimTime[41]), .A(timeStampPkt[49]));
Q_ASSIGN U52 ( .B(xc_top.ixcSimTime[40]), .A(timeStampPkt[48]));
Q_ASSIGN U53 ( .B(xc_top.ixcSimTime[39]), .A(timeStampPkt[47]));
Q_ASSIGN U54 ( .B(xc_top.ixcSimTime[38]), .A(timeStampPkt[46]));
Q_ASSIGN U55 ( .B(xc_top.ixcSimTime[37]), .A(timeStampPkt[45]));
Q_ASSIGN U56 ( .B(xc_top.ixcSimTime[36]), .A(timeStampPkt[44]));
Q_ASSIGN U57 ( .B(xc_top.ixcSimTime[35]), .A(timeStampPkt[43]));
Q_ASSIGN U58 ( .B(xc_top.ixcSimTime[34]), .A(timeStampPkt[42]));
Q_ASSIGN U59 ( .B(xc_top.ixcSimTime[33]), .A(timeStampPkt[41]));
Q_ASSIGN U60 ( .B(xc_top.ixcSimTime[32]), .A(timeStampPkt[40]));
Q_ASSIGN U61 ( .B(xc_top.ixcSimTime[31]), .A(timeStampPkt[39]));
Q_ASSIGN U62 ( .B(xc_top.ixcSimTime[30]), .A(timeStampPkt[38]));
Q_ASSIGN U63 ( .B(xc_top.ixcSimTime[29]), .A(timeStampPkt[37]));
Q_ASSIGN U64 ( .B(xc_top.ixcSimTime[28]), .A(timeStampPkt[36]));
Q_ASSIGN U65 ( .B(xc_top.ixcSimTime[27]), .A(timeStampPkt[35]));
Q_ASSIGN U66 ( .B(xc_top.ixcSimTime[26]), .A(timeStampPkt[34]));
Q_ASSIGN U67 ( .B(xc_top.ixcSimTime[25]), .A(timeStampPkt[33]));
Q_ASSIGN U68 ( .B(xc_top.ixcSimTime[24]), .A(timeStampPkt[32]));
Q_ASSIGN U69 ( .B(xc_top.ixcSimTime[23]), .A(timeStampPkt[23]));
Q_ASSIGN U70 ( .B(xc_top.ixcSimTime[22]), .A(timeStampPkt[22]));
Q_ASSIGN U71 ( .B(xc_top.ixcSimTime[21]), .A(timeStampPkt[21]));
Q_ASSIGN U72 ( .B(xc_top.ixcSimTime[20]), .A(timeStampPkt[20]));
Q_ASSIGN U73 ( .B(xc_top.ixcSimTime[19]), .A(timeStampPkt[19]));
Q_ASSIGN U74 ( .B(xc_top.ixcSimTime[18]), .A(timeStampPkt[18]));
Q_ASSIGN U75 ( .B(xc_top.ixcSimTime[17]), .A(timeStampPkt[17]));
Q_ASSIGN U76 ( .B(xc_top.ixcSimTime[16]), .A(timeStampPkt[16]));
Q_ASSIGN U77 ( .B(xc_top.ixcSimTime[15]), .A(timeStampPkt[15]));
Q_ASSIGN U78 ( .B(xc_top.ixcSimTime[14]), .A(timeStampPkt[14]));
Q_ASSIGN U79 ( .B(xc_top.ixcSimTime[13]), .A(timeStampPkt[13]));
Q_ASSIGN U80 ( .B(xc_top.ixcSimTime[12]), .A(timeStampPkt[12]));
Q_ASSIGN U81 ( .B(xc_top.ixcSimTime[11]), .A(timeStampPkt[11]));
Q_ASSIGN U82 ( .B(xc_top.ixcSimTime[10]), .A(timeStampPkt[10]));
Q_ASSIGN U83 ( .B(xc_top.ixcSimTime[9]), .A(timeStampPkt[9]));
Q_ASSIGN U84 ( .B(xc_top.ixcSimTime[8]), .A(timeStampPkt[8]));
Q_ASSIGN U85 ( .B(xc_top.ixcSimTime[7]), .A(timeStampPkt[7]));
Q_ASSIGN U86 ( .B(xc_top.ixcSimTime[6]), .A(timeStampPkt[6]));
Q_ASSIGN U87 ( .B(xc_top.ixcSimTime[5]), .A(timeStampPkt[5]));
Q_ASSIGN U88 ( .B(xc_top.ixcSimTime[4]), .A(timeStampPkt[4]));
Q_ASSIGN U89 ( .B(xc_top.ixcSimTime[3]), .A(timeStampPkt[3]));
Q_ASSIGN U90 ( .B(xc_top.ixcSimTime[2]), .A(timeStampPkt[2]));
Q_ASSIGN U91 ( .B(xc_top.ixcSimTime[1]), .A(timeStampPkt[1]));
Q_ASSIGN U92 ( .B(xc_top.ixcSimTime[0]), .A(timeStampPkt[0]));
Q_INV U93 ( .A(n97), .Z(n3347));
Q_INV U94 ( .A(n113), .Z(n3346));
Q_INV U95 ( .A(n98), .Z(n3345));
Q_INV U96 ( .A(ofifoAddr7N[2]), .Z(ofifoAddr3N[2]));
Q_INV U97 ( .A(ofifoAddr5N[2]), .Z(ofifoAddr1N[2]));
Q_INV U98 ( .A(n79), .Z(n3344));
Q_INV U99 ( .A(n80), .Z(n3343));
Q_INV U100 ( .A(n81), .Z(n3342));
Q_INV U101 ( .A(n82), .Z(n3341));
Q_INV U102 ( .A(ofifoAddr6N[2]), .Z(ofifoAddr2N[2]));
Q_INV U103 ( .A(ofifoAddr7N[1]), .Z(ofifoAddr5N[1]));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_XOR2 U105 ( .A0(n3320), .A1(n3319), .Z(timeStampPkt[24]));
Q_XOR3 U106 ( .A0(timeStampPkt[1]), .A1(timeStampPkt[0]), .A2(n3321), .Z(n3319));
Q_XOR3 U107 ( .A0(timeStampPkt[4]), .A1(timeStampPkt[3]), .A2(timeStampPkt[2]), .Z(n3320));
Q_XOR3 U108 ( .A0(timeStampPkt[7]), .A1(timeStampPkt[6]), .A2(timeStampPkt[5]), .Z(n3321));
Q_XOR2 U109 ( .A0(n3323), .A1(n3322), .Z(timeStampPkt[25]));
Q_XOR3 U110 ( .A0(timeStampPkt[9]), .A1(timeStampPkt[8]), .A2(n3324), .Z(n3322));
Q_XOR3 U111 ( .A0(timeStampPkt[12]), .A1(timeStampPkt[11]), .A2(timeStampPkt[10]), .Z(n3323));
Q_XOR3 U112 ( .A0(timeStampPkt[15]), .A1(timeStampPkt[14]), .A2(timeStampPkt[13]), .Z(n3324));
Q_XOR2 U113 ( .A0(n3326), .A1(n3325), .Z(timeStampPkt[26]));
Q_XOR3 U114 ( .A0(timeStampPkt[17]), .A1(timeStampPkt[16]), .A2(n3327), .Z(n3325));
Q_XOR3 U115 ( .A0(timeStampPkt[20]), .A1(timeStampPkt[19]), .A2(timeStampPkt[18]), .Z(n3326));
Q_XOR3 U116 ( .A0(timeStampPkt[23]), .A1(timeStampPkt[22]), .A2(timeStampPkt[21]), .Z(n3327));
Q_XOR2 U117 ( .A0(n3329), .A1(n3328), .Z(timeStampPkt[27]));
Q_XOR3 U118 ( .A0(timeStampPkt[33]), .A1(timeStampPkt[32]), .A2(n3330), .Z(n3328));
Q_XOR3 U119 ( .A0(timeStampPkt[36]), .A1(timeStampPkt[35]), .A2(timeStampPkt[34]), .Z(n3329));
Q_XOR3 U120 ( .A0(timeStampPkt[39]), .A1(timeStampPkt[38]), .A2(timeStampPkt[37]), .Z(n3330));
Q_XOR2 U121 ( .A0(n3332), .A1(n3331), .Z(timeStampPkt[28]));
Q_XOR3 U122 ( .A0(timeStampPkt[41]), .A1(timeStampPkt[40]), .A2(n3333), .Z(n3331));
Q_XOR3 U123 ( .A0(timeStampPkt[44]), .A1(timeStampPkt[43]), .A2(timeStampPkt[42]), .Z(n3332));
Q_XOR3 U124 ( .A0(timeStampPkt[47]), .A1(timeStampPkt[46]), .A2(timeStampPkt[45]), .Z(n3333));
Q_XOR2 U125 ( .A0(n3335), .A1(n3334), .Z(timeStampPkt[29]));
Q_XOR3 U126 ( .A0(timeStampPkt[49]), .A1(timeStampPkt[48]), .A2(n3336), .Z(n3334));
Q_XOR3 U127 ( .A0(timeStampPkt[52]), .A1(timeStampPkt[51]), .A2(timeStampPkt[50]), .Z(n3335));
Q_XOR3 U128 ( .A0(timeStampPkt[55]), .A1(timeStampPkt[54]), .A2(timeStampPkt[53]), .Z(n3336));
Q_XOR2 U129 ( .A0(n3338), .A1(n3337), .Z(timeStampPkt[30]));
Q_XOR3 U130 ( .A0(timeStampPkt[57]), .A1(timeStampPkt[56]), .A2(n3339), .Z(n3337));
Q_XOR3 U131 ( .A0(timeStampPkt[60]), .A1(timeStampPkt[59]), .A2(timeStampPkt[58]), .Z(n3338));
Q_XOR3 U132 ( .A0(timeStampPkt[63]), .A1(timeStampPkt[62]), .A2(timeStampPkt[61]), .Z(n3339));
ixc_assign _zz_strnp_0 ( scgGFreq, GFreq);
Q_RDN U134 ( .Z(GFtsReq));
Q_RDN U135 ( .Z(GFidata[0]));
Q_RDN U136 ( .Z(GFidata[1]));
Q_RDN U137 ( .Z(GFidata[2]));
Q_RDN U138 ( .Z(GFidata[3]));
Q_RDN U139 ( .Z(GFidata[4]));
Q_RDN U140 ( .Z(GFidata[5]));
Q_RDN U141 ( .Z(GFidata[6]));
Q_RDN U142 ( .Z(GFidata[7]));
Q_RDN U143 ( .Z(GFidata[8]));
Q_RDN U144 ( .Z(GFidata[9]));
Q_RDN U145 ( .Z(GFidata[10]));
Q_RDN U146 ( .Z(GFidata[11]));
Q_RDN U147 ( .Z(GFidata[12]));
Q_RDN U148 ( .Z(GFidata[13]));
Q_RDN U149 ( .Z(GFidata[14]));
Q_RDN U150 ( .Z(GFidata[15]));
Q_RDN U151 ( .Z(GFidata[16]));
Q_RDN U152 ( .Z(GFidata[17]));
Q_RDN U153 ( .Z(GFidata[18]));
Q_RDN U154 ( .Z(GFidata[19]));
Q_RDN U155 ( .Z(GFidata[20]));
Q_RDN U156 ( .Z(GFidata[21]));
Q_RDN U157 ( .Z(GFidata[22]));
Q_RDN U158 ( .Z(GFidata[23]));
Q_RDN U159 ( .Z(GFidata[24]));
Q_RDN U160 ( .Z(GFidata[25]));
Q_RDN U161 ( .Z(GFidata[26]));
Q_RDN U162 ( .Z(GFidata[27]));
Q_RDN U163 ( .Z(GFidata[28]));
Q_RDN U164 ( .Z(GFidata[29]));
Q_RDN U165 ( .Z(GFidata[30]));
Q_RDN U166 ( .Z(GFidata[31]));
Q_RDN U167 ( .Z(GFidata[32]));
Q_RDN U168 ( .Z(GFidata[33]));
Q_RDN U169 ( .Z(GFidata[34]));
Q_RDN U170 ( .Z(GFidata[35]));
Q_RDN U171 ( .Z(GFidata[36]));
Q_RDN U172 ( .Z(GFidata[37]));
Q_RDN U173 ( .Z(GFidata[38]));
Q_RDN U174 ( .Z(GFidata[39]));
Q_RDN U175 ( .Z(GFidata[40]));
Q_RDN U176 ( .Z(GFidata[41]));
Q_RDN U177 ( .Z(GFidata[42]));
Q_RDN U178 ( .Z(GFidata[43]));
Q_RDN U179 ( .Z(GFidata[44]));
Q_RDN U180 ( .Z(GFidata[45]));
Q_RDN U181 ( .Z(GFidata[46]));
Q_RDN U182 ( .Z(GFidata[47]));
Q_RDN U183 ( .Z(GFidata[48]));
Q_RDN U184 ( .Z(GFidata[49]));
Q_RDN U185 ( .Z(GFidata[50]));
Q_RDN U186 ( .Z(GFidata[51]));
Q_RDN U187 ( .Z(GFidata[52]));
Q_RDN U188 ( .Z(GFidata[53]));
Q_RDN U189 ( .Z(GFidata[54]));
Q_RDN U190 ( .Z(GFidata[55]));
Q_RDN U191 ( .Z(GFidata[56]));
Q_RDN U192 ( .Z(GFidata[57]));
Q_RDN U193 ( .Z(GFidata[58]));
Q_RDN U194 ( .Z(GFidata[59]));
Q_RDN U195 ( .Z(GFidata[60]));
Q_RDN U196 ( .Z(GFidata[61]));
Q_RDN U197 ( .Z(GFidata[62]));
Q_RDN U198 ( .Z(GFidata[63]));
Q_RDN U199 ( .Z(GFidata[64]));
Q_RDN U200 ( .Z(GFidata[65]));
Q_RDN U201 ( .Z(GFidata[66]));
Q_RDN U202 ( .Z(GFidata[67]));
Q_RDN U203 ( .Z(GFidata[68]));
Q_RDN U204 ( .Z(GFidata[69]));
Q_RDN U205 ( .Z(GFidata[70]));
Q_RDN U206 ( .Z(GFidata[71]));
Q_RDN U207 ( .Z(GFidata[72]));
Q_RDN U208 ( .Z(GFidata[73]));
Q_RDN U209 ( .Z(GFidata[74]));
Q_RDN U210 ( .Z(GFidata[75]));
Q_RDN U211 ( .Z(GFidata[76]));
Q_RDN U212 ( .Z(GFidata[77]));
Q_RDN U213 ( .Z(GFidata[78]));
Q_RDN U214 ( .Z(GFidata[79]));
Q_RDN U215 ( .Z(GFidata[80]));
Q_RDN U216 ( .Z(GFidata[81]));
Q_RDN U217 ( .Z(GFidata[82]));
Q_RDN U218 ( .Z(GFidata[83]));
Q_RDN U219 ( .Z(GFidata[84]));
Q_RDN U220 ( .Z(GFidata[85]));
Q_RDN U221 ( .Z(GFidata[86]));
Q_RDN U222 ( .Z(GFidata[87]));
Q_RDN U223 ( .Z(GFidata[88]));
Q_RDN U224 ( .Z(GFidata[89]));
Q_RDN U225 ( .Z(GFidata[90]));
Q_RDN U226 ( .Z(GFidata[91]));
Q_RDN U227 ( .Z(GFidata[92]));
Q_RDN U228 ( .Z(GFidata[93]));
Q_RDN U229 ( .Z(GFidata[94]));
Q_RDN U230 ( .Z(GFidata[95]));
Q_RDN U231 ( .Z(GFidata[96]));
Q_RDN U232 ( .Z(GFidata[97]));
Q_RDN U233 ( .Z(GFidata[98]));
Q_RDN U234 ( .Z(GFidata[99]));
Q_RDN U235 ( .Z(GFidata[100]));
Q_RDN U236 ( .Z(GFidata[101]));
Q_RDN U237 ( .Z(GFidata[102]));
Q_RDN U238 ( .Z(GFidata[103]));
Q_RDN U239 ( .Z(GFidata[104]));
Q_RDN U240 ( .Z(GFidata[105]));
Q_RDN U241 ( .Z(GFidata[106]));
Q_RDN U242 ( .Z(GFidata[107]));
Q_RDN U243 ( .Z(GFidata[108]));
Q_RDN U244 ( .Z(GFidata[109]));
Q_RDN U245 ( .Z(GFidata[110]));
Q_RDN U246 ( .Z(GFidata[111]));
Q_RDN U247 ( .Z(GFidata[112]));
Q_RDN U248 ( .Z(GFidata[113]));
Q_RDN U249 ( .Z(GFidata[114]));
Q_RDN U250 ( .Z(GFidata[115]));
Q_RDN U251 ( .Z(GFidata[116]));
Q_RDN U252 ( .Z(GFidata[117]));
Q_RDN U253 ( .Z(GFidata[118]));
Q_RDN U254 ( .Z(GFidata[119]));
Q_RDN U255 ( .Z(GFidata[120]));
Q_RDN U256 ( .Z(GFidata[121]));
Q_RDN U257 ( .Z(GFidata[122]));
Q_RDN U258 ( .Z(GFidata[123]));
Q_RDN U259 ( .Z(GFidata[124]));
Q_RDN U260 ( .Z(GFidata[125]));
Q_RDN U261 ( .Z(GFidata[126]));
Q_RDN U262 ( .Z(GFidata[127]));
Q_RDN U263 ( .Z(GFidata[128]));
Q_RDN U264 ( .Z(GFidata[129]));
Q_RDN U265 ( .Z(GFidata[130]));
Q_RDN U266 ( .Z(GFidata[131]));
Q_RDN U267 ( .Z(GFidata[132]));
Q_RDN U268 ( .Z(GFidata[133]));
Q_RDN U269 ( .Z(GFidata[134]));
Q_RDN U270 ( .Z(GFidata[135]));
Q_RDN U271 ( .Z(GFidata[136]));
Q_RDN U272 ( .Z(GFidata[137]));
Q_RDN U273 ( .Z(GFidata[138]));
Q_RDN U274 ( .Z(GFidata[139]));
Q_RDN U275 ( .Z(GFidata[140]));
Q_RDN U276 ( .Z(GFidata[141]));
Q_RDN U277 ( .Z(GFidata[142]));
Q_RDN U278 ( .Z(GFidata[143]));
Q_RDN U279 ( .Z(GFidata[144]));
Q_RDN U280 ( .Z(GFidata[145]));
Q_RDN U281 ( .Z(GFidata[146]));
Q_RDN U282 ( .Z(GFidata[147]));
Q_RDN U283 ( .Z(GFidata[148]));
Q_RDN U284 ( .Z(GFidata[149]));
Q_RDN U285 ( .Z(GFidata[150]));
Q_RDN U286 ( .Z(GFidata[151]));
Q_RDN U287 ( .Z(GFidata[152]));
Q_RDN U288 ( .Z(GFidata[153]));
Q_RDN U289 ( .Z(GFidata[154]));
Q_RDN U290 ( .Z(GFidata[155]));
Q_RDN U291 ( .Z(GFidata[156]));
Q_RDN U292 ( .Z(GFidata[157]));
Q_RDN U293 ( .Z(GFidata[158]));
Q_RDN U294 ( .Z(GFidata[159]));
Q_RDN U295 ( .Z(GFidata[160]));
Q_RDN U296 ( .Z(GFidata[161]));
Q_RDN U297 ( .Z(GFidata[162]));
Q_RDN U298 ( .Z(GFidata[163]));
Q_RDN U299 ( .Z(GFidata[164]));
Q_RDN U300 ( .Z(GFidata[165]));
Q_RDN U301 ( .Z(GFidata[166]));
Q_RDN U302 ( .Z(GFidata[167]));
Q_RDN U303 ( .Z(GFidata[168]));
Q_RDN U304 ( .Z(GFidata[169]));
Q_RDN U305 ( .Z(GFidata[170]));
Q_RDN U306 ( .Z(GFidata[171]));
Q_RDN U307 ( .Z(GFidata[172]));
Q_RDN U308 ( .Z(GFidata[173]));
Q_RDN U309 ( .Z(GFidata[174]));
Q_RDN U310 ( .Z(GFidata[175]));
Q_RDN U311 ( .Z(GFidata[176]));
Q_RDN U312 ( .Z(GFidata[177]));
Q_RDN U313 ( .Z(GFidata[178]));
Q_RDN U314 ( .Z(GFidata[179]));
Q_RDN U315 ( .Z(GFidata[180]));
Q_RDN U316 ( .Z(GFidata[181]));
Q_RDN U317 ( .Z(GFidata[182]));
Q_RDN U318 ( .Z(GFidata[183]));
Q_RDN U319 ( .Z(GFidata[184]));
Q_RDN U320 ( .Z(GFidata[185]));
Q_RDN U321 ( .Z(GFidata[186]));
Q_RDN U322 ( .Z(GFidata[187]));
Q_RDN U323 ( .Z(GFidata[188]));
Q_RDN U324 ( .Z(GFidata[189]));
Q_RDN U325 ( .Z(GFidata[190]));
Q_RDN U326 ( .Z(GFidata[191]));
Q_RDN U327 ( .Z(GFidata[192]));
Q_RDN U328 ( .Z(GFidata[193]));
Q_RDN U329 ( .Z(GFidata[194]));
Q_RDN U330 ( .Z(GFidata[195]));
Q_RDN U331 ( .Z(GFidata[196]));
Q_RDN U332 ( .Z(GFidata[197]));
Q_RDN U333 ( .Z(GFidata[198]));
Q_RDN U334 ( .Z(GFidata[199]));
Q_RDN U335 ( .Z(GFidata[200]));
Q_RDN U336 ( .Z(GFidata[201]));
Q_RDN U337 ( .Z(GFidata[202]));
Q_RDN U338 ( .Z(GFidata[203]));
Q_RDN U339 ( .Z(GFidata[204]));
Q_RDN U340 ( .Z(GFidata[205]));
Q_RDN U341 ( .Z(GFidata[206]));
Q_RDN U342 ( .Z(GFidata[207]));
Q_RDN U343 ( .Z(GFidata[208]));
Q_RDN U344 ( .Z(GFidata[209]));
Q_RDN U345 ( .Z(GFidata[210]));
Q_RDN U346 ( .Z(GFidata[211]));
Q_RDN U347 ( .Z(GFidata[212]));
Q_RDN U348 ( .Z(GFidata[213]));
Q_RDN U349 ( .Z(GFidata[214]));
Q_RDN U350 ( .Z(GFidata[215]));
Q_RDN U351 ( .Z(GFidata[216]));
Q_RDN U352 ( .Z(GFidata[217]));
Q_RDN U353 ( .Z(GFidata[218]));
Q_RDN U354 ( .Z(GFidata[219]));
Q_RDN U355 ( .Z(GFidata[220]));
Q_RDN U356 ( .Z(GFidata[221]));
Q_RDN U357 ( .Z(GFidata[222]));
Q_RDN U358 ( .Z(GFidata[223]));
Q_RDN U359 ( .Z(GFidata[224]));
Q_RDN U360 ( .Z(GFidata[225]));
Q_RDN U361 ( .Z(GFidata[226]));
Q_RDN U362 ( .Z(GFidata[227]));
Q_RDN U363 ( .Z(GFidata[228]));
Q_RDN U364 ( .Z(GFidata[229]));
Q_RDN U365 ( .Z(GFidata[230]));
Q_RDN U366 ( .Z(GFidata[231]));
Q_RDN U367 ( .Z(GFidata[232]));
Q_RDN U368 ( .Z(GFidata[233]));
Q_RDN U369 ( .Z(GFidata[234]));
Q_RDN U370 ( .Z(GFidata[235]));
Q_RDN U371 ( .Z(GFidata[236]));
Q_RDN U372 ( .Z(GFidata[237]));
Q_RDN U373 ( .Z(GFidata[238]));
Q_RDN U374 ( .Z(GFidata[239]));
Q_RDN U375 ( .Z(GFidata[240]));
Q_RDN U376 ( .Z(GFidata[241]));
Q_RDN U377 ( .Z(GFidata[242]));
Q_RDN U378 ( .Z(GFidata[243]));
Q_RDN U379 ( .Z(GFidata[244]));
Q_RDN U380 ( .Z(GFidata[245]));
Q_RDN U381 ( .Z(GFidata[246]));
Q_RDN U382 ( .Z(GFidata[247]));
Q_RDN U383 ( .Z(GFidata[248]));
Q_RDN U384 ( .Z(GFidata[249]));
Q_RDN U385 ( .Z(GFidata[250]));
Q_RDN U386 ( .Z(GFidata[251]));
Q_RDN U387 ( .Z(GFidata[252]));
Q_RDN U388 ( .Z(GFidata[253]));
Q_RDN U389 ( .Z(GFidata[254]));
Q_RDN U390 ( .Z(GFidata[255]));
Q_RDN U391 ( .Z(GFidata[256]));
Q_RDN U392 ( .Z(GFidata[257]));
Q_RDN U393 ( .Z(GFidata[258]));
Q_RDN U394 ( .Z(GFidata[259]));
Q_RDN U395 ( .Z(GFidata[260]));
Q_RDN U396 ( .Z(GFidata[261]));
Q_RDN U397 ( .Z(GFidata[262]));
Q_RDN U398 ( .Z(GFidata[263]));
Q_RDN U399 ( .Z(GFidata[264]));
Q_RDN U400 ( .Z(GFidata[265]));
Q_RDN U401 ( .Z(GFidata[266]));
Q_RDN U402 ( .Z(GFidata[267]));
Q_RDN U403 ( .Z(GFidata[268]));
Q_RDN U404 ( .Z(GFidata[269]));
Q_RDN U405 ( .Z(GFidata[270]));
Q_RDN U406 ( .Z(GFidata[271]));
Q_RDN U407 ( .Z(GFidata[272]));
Q_RDN U408 ( .Z(GFidata[273]));
Q_RDN U409 ( .Z(GFidata[274]));
Q_RDN U410 ( .Z(GFidata[275]));
Q_RDN U411 ( .Z(GFidata[276]));
Q_RDN U412 ( .Z(GFidata[277]));
Q_RDN U413 ( .Z(GFidata[278]));
Q_RDN U414 ( .Z(GFidata[279]));
Q_RDN U415 ( .Z(GFidata[280]));
Q_RDN U416 ( .Z(GFidata[281]));
Q_RDN U417 ( .Z(GFidata[282]));
Q_RDN U418 ( .Z(GFidata[283]));
Q_RDN U419 ( .Z(GFidata[284]));
Q_RDN U420 ( .Z(GFidata[285]));
Q_RDN U421 ( .Z(GFidata[286]));
Q_RDN U422 ( .Z(GFidata[287]));
Q_RDN U423 ( .Z(GFidata[288]));
Q_RDN U424 ( .Z(GFidata[289]));
Q_RDN U425 ( .Z(GFidata[290]));
Q_RDN U426 ( .Z(GFidata[291]));
Q_RDN U427 ( .Z(GFidata[292]));
Q_RDN U428 ( .Z(GFidata[293]));
Q_RDN U429 ( .Z(GFidata[294]));
Q_RDN U430 ( .Z(GFidata[295]));
Q_RDN U431 ( .Z(GFidata[296]));
Q_RDN U432 ( .Z(GFidata[297]));
Q_RDN U433 ( .Z(GFidata[298]));
Q_RDN U434 ( .Z(GFidata[299]));
Q_RDN U435 ( .Z(GFidata[300]));
Q_RDN U436 ( .Z(GFidata[301]));
Q_RDN U437 ( .Z(GFidata[302]));
Q_RDN U438 ( .Z(GFidata[303]));
Q_RDN U439 ( .Z(GFidata[304]));
Q_RDN U440 ( .Z(GFidata[305]));
Q_RDN U441 ( .Z(GFidata[306]));
Q_RDN U442 ( .Z(GFidata[307]));
Q_RDN U443 ( .Z(GFidata[308]));
Q_RDN U444 ( .Z(GFidata[309]));
Q_RDN U445 ( .Z(GFidata[310]));
Q_RDN U446 ( .Z(GFidata[311]));
Q_RDN U447 ( .Z(GFidata[312]));
Q_RDN U448 ( .Z(GFidata[313]));
Q_RDN U449 ( .Z(GFidata[314]));
Q_RDN U450 ( .Z(GFidata[315]));
Q_RDN U451 ( .Z(GFidata[316]));
Q_RDN U452 ( .Z(GFidata[317]));
Q_RDN U453 ( .Z(GFidata[318]));
Q_RDN U454 ( .Z(GFidata[319]));
Q_RDN U455 ( .Z(GFidata[320]));
Q_RDN U456 ( .Z(GFidata[321]));
Q_RDN U457 ( .Z(GFidata[322]));
Q_RDN U458 ( .Z(GFidata[323]));
Q_RDN U459 ( .Z(GFidata[324]));
Q_RDN U460 ( .Z(GFidata[325]));
Q_RDN U461 ( .Z(GFidata[326]));
Q_RDN U462 ( .Z(GFidata[327]));
Q_RDN U463 ( .Z(GFidata[328]));
Q_RDN U464 ( .Z(GFidata[329]));
Q_RDN U465 ( .Z(GFidata[330]));
Q_RDN U466 ( .Z(GFidata[331]));
Q_RDN U467 ( .Z(GFidata[332]));
Q_RDN U468 ( .Z(GFidata[333]));
Q_RDN U469 ( .Z(GFidata[334]));
Q_RDN U470 ( .Z(GFidata[335]));
Q_RDN U471 ( .Z(GFidata[336]));
Q_RDN U472 ( .Z(GFidata[337]));
Q_RDN U473 ( .Z(GFidata[338]));
Q_RDN U474 ( .Z(GFidata[339]));
Q_RDN U475 ( .Z(GFidata[340]));
Q_RDN U476 ( .Z(GFidata[341]));
Q_RDN U477 ( .Z(GFidata[342]));
Q_RDN U478 ( .Z(GFidata[343]));
Q_RDN U479 ( .Z(GFidata[344]));
Q_RDN U480 ( .Z(GFidata[345]));
Q_RDN U481 ( .Z(GFidata[346]));
Q_RDN U482 ( .Z(GFidata[347]));
Q_RDN U483 ( .Z(GFidata[348]));
Q_RDN U484 ( .Z(GFidata[349]));
Q_RDN U485 ( .Z(GFidata[350]));
Q_RDN U486 ( .Z(GFidata[351]));
Q_RDN U487 ( .Z(GFidata[352]));
Q_RDN U488 ( .Z(GFidata[353]));
Q_RDN U489 ( .Z(GFidata[354]));
Q_RDN U490 ( .Z(GFidata[355]));
Q_RDN U491 ( .Z(GFidata[356]));
Q_RDN U492 ( .Z(GFidata[357]));
Q_RDN U493 ( .Z(GFidata[358]));
Q_RDN U494 ( .Z(GFidata[359]));
Q_RDN U495 ( .Z(GFidata[360]));
Q_RDN U496 ( .Z(GFidata[361]));
Q_RDN U497 ( .Z(GFidata[362]));
Q_RDN U498 ( .Z(GFidata[363]));
Q_RDN U499 ( .Z(GFidata[364]));
Q_RDN U500 ( .Z(GFidata[365]));
Q_RDN U501 ( .Z(GFidata[366]));
Q_RDN U502 ( .Z(GFidata[367]));
Q_RDN U503 ( .Z(GFidata[368]));
Q_RDN U504 ( .Z(GFidata[369]));
Q_RDN U505 ( .Z(GFidata[370]));
Q_RDN U506 ( .Z(GFidata[371]));
Q_RDN U507 ( .Z(GFidata[372]));
Q_RDN U508 ( .Z(GFidata[373]));
Q_RDN U509 ( .Z(GFidata[374]));
Q_RDN U510 ( .Z(GFidata[375]));
Q_RDN U511 ( .Z(GFidata[376]));
Q_RDN U512 ( .Z(GFidata[377]));
Q_RDN U513 ( .Z(GFidata[378]));
Q_RDN U514 ( .Z(GFidata[379]));
Q_RDN U515 ( .Z(GFidata[380]));
Q_RDN U516 ( .Z(GFidata[381]));
Q_RDN U517 ( .Z(GFidata[382]));
Q_RDN U518 ( .Z(GFidata[383]));
Q_RDN U519 ( .Z(GFidata[384]));
Q_RDN U520 ( .Z(GFidata[385]));
Q_RDN U521 ( .Z(GFidata[386]));
Q_RDN U522 ( .Z(GFidata[387]));
Q_RDN U523 ( .Z(GFidata[388]));
Q_RDN U524 ( .Z(GFidata[389]));
Q_RDN U525 ( .Z(GFidata[390]));
Q_RDN U526 ( .Z(GFidata[391]));
Q_RDN U527 ( .Z(GFidata[392]));
Q_RDN U528 ( .Z(GFidata[393]));
Q_RDN U529 ( .Z(GFidata[394]));
Q_RDN U530 ( .Z(GFidata[395]));
Q_RDN U531 ( .Z(GFidata[396]));
Q_RDN U532 ( .Z(GFidata[397]));
Q_RDN U533 ( .Z(GFidata[398]));
Q_RDN U534 ( .Z(GFidata[399]));
Q_RDN U535 ( .Z(GFidata[400]));
Q_RDN U536 ( .Z(GFidata[401]));
Q_RDN U537 ( .Z(GFidata[402]));
Q_RDN U538 ( .Z(GFidata[403]));
Q_RDN U539 ( .Z(GFidata[404]));
Q_RDN U540 ( .Z(GFidata[405]));
Q_RDN U541 ( .Z(GFidata[406]));
Q_RDN U542 ( .Z(GFidata[407]));
Q_RDN U543 ( .Z(GFidata[408]));
Q_RDN U544 ( .Z(GFidata[409]));
Q_RDN U545 ( .Z(GFidata[410]));
Q_RDN U546 ( .Z(GFidata[411]));
Q_RDN U547 ( .Z(GFidata[412]));
Q_RDN U548 ( .Z(GFidata[413]));
Q_RDN U549 ( .Z(GFidata[414]));
Q_RDN U550 ( .Z(GFidata[415]));
Q_RDN U551 ( .Z(GFidata[416]));
Q_RDN U552 ( .Z(GFidata[417]));
Q_RDN U553 ( .Z(GFidata[418]));
Q_RDN U554 ( .Z(GFidata[419]));
Q_RDN U555 ( .Z(GFidata[420]));
Q_RDN U556 ( .Z(GFidata[421]));
Q_RDN U557 ( .Z(GFidata[422]));
Q_RDN U558 ( .Z(GFidata[423]));
Q_RDN U559 ( .Z(GFidata[424]));
Q_RDN U560 ( .Z(GFidata[425]));
Q_RDN U561 ( .Z(GFidata[426]));
Q_RDN U562 ( .Z(GFidata[427]));
Q_RDN U563 ( .Z(GFidata[428]));
Q_RDN U564 ( .Z(GFidata[429]));
Q_RDN U565 ( .Z(GFidata[430]));
Q_RDN U566 ( .Z(GFidata[431]));
Q_RDN U567 ( .Z(GFidata[432]));
Q_RDN U568 ( .Z(GFidata[433]));
Q_RDN U569 ( .Z(GFidata[434]));
Q_RDN U570 ( .Z(GFidata[435]));
Q_RDN U571 ( .Z(GFidata[436]));
Q_RDN U572 ( .Z(GFidata[437]));
Q_RDN U573 ( .Z(GFidata[438]));
Q_RDN U574 ( .Z(GFidata[439]));
Q_RDN U575 ( .Z(GFidata[440]));
Q_RDN U576 ( .Z(GFidata[441]));
Q_RDN U577 ( .Z(GFidata[442]));
Q_RDN U578 ( .Z(GFidata[443]));
Q_RDN U579 ( .Z(GFidata[444]));
Q_RDN U580 ( .Z(GFidata[445]));
Q_RDN U581 ( .Z(GFidata[446]));
Q_RDN U582 ( .Z(GFidata[447]));
Q_RDN U583 ( .Z(GFidata[448]));
Q_RDN U584 ( .Z(GFidata[449]));
Q_RDN U585 ( .Z(GFidata[450]));
Q_RDN U586 ( .Z(GFidata[451]));
Q_RDN U587 ( .Z(GFidata[452]));
Q_RDN U588 ( .Z(GFidata[453]));
Q_RDN U589 ( .Z(GFidata[454]));
Q_RDN U590 ( .Z(GFidata[455]));
Q_RDN U591 ( .Z(GFidata[456]));
Q_RDN U592 ( .Z(GFidata[457]));
Q_RDN U593 ( .Z(GFidata[458]));
Q_RDN U594 ( .Z(GFidata[459]));
Q_RDN U595 ( .Z(GFidata[460]));
Q_RDN U596 ( .Z(GFidata[461]));
Q_RDN U597 ( .Z(GFidata[462]));
Q_RDN U598 ( .Z(GFidata[463]));
Q_RDN U599 ( .Z(GFidata[464]));
Q_RDN U600 ( .Z(GFidata[465]));
Q_RDN U601 ( .Z(GFidata[466]));
Q_RDN U602 ( .Z(GFidata[467]));
Q_RDN U603 ( .Z(GFidata[468]));
Q_RDN U604 ( .Z(GFidata[469]));
Q_RDN U605 ( .Z(GFidata[470]));
Q_RDN U606 ( .Z(GFidata[471]));
Q_RDN U607 ( .Z(GFidata[472]));
Q_RDN U608 ( .Z(GFidata[473]));
Q_RDN U609 ( .Z(GFidata[474]));
Q_RDN U610 ( .Z(GFidata[475]));
Q_RDN U611 ( .Z(GFidata[476]));
Q_RDN U612 ( .Z(GFidata[477]));
Q_RDN U613 ( .Z(GFidata[478]));
Q_RDN U614 ( .Z(GFidata[479]));
Q_RDN U615 ( .Z(GFidata[480]));
Q_RDN U616 ( .Z(GFidata[481]));
Q_RDN U617 ( .Z(GFidata[482]));
Q_RDN U618 ( .Z(GFidata[483]));
Q_RDN U619 ( .Z(GFidata[484]));
Q_RDN U620 ( .Z(GFidata[485]));
Q_RDN U621 ( .Z(GFidata[486]));
Q_RDN U622 ( .Z(GFidata[487]));
Q_RDN U623 ( .Z(GFidata[488]));
Q_RDN U624 ( .Z(GFidata[489]));
Q_RDN U625 ( .Z(GFidata[490]));
Q_RDN U626 ( .Z(GFidata[491]));
Q_RDN U627 ( .Z(GFidata[492]));
Q_RDN U628 ( .Z(GFidata[493]));
Q_RDN U629 ( .Z(GFidata[494]));
Q_RDN U630 ( .Z(GFidata[495]));
Q_RDN U631 ( .Z(GFidata[496]));
Q_RDN U632 ( .Z(GFidata[497]));
Q_RDN U633 ( .Z(GFidata[498]));
Q_RDN U634 ( .Z(GFidata[499]));
Q_RDN U635 ( .Z(GFidata[500]));
Q_RDN U636 ( .Z(GFidata[501]));
Q_RDN U637 ( .Z(GFidata[502]));
Q_RDN U638 ( .Z(GFidata[503]));
Q_RDN U639 ( .Z(GFidata[504]));
Q_RDN U640 ( .Z(GFidata[505]));
Q_RDN U641 ( .Z(GFidata[506]));
Q_RDN U642 ( .Z(GFidata[507]));
Q_RDN U643 ( .Z(GFidata[508]));
Q_RDN U644 ( .Z(GFidata[509]));
Q_RDN U645 ( .Z(GFidata[510]));
Q_RDN U646 ( .Z(GFidata[511]));
Q_RDN U647 ( .Z(GFlen[0]));
Q_RDN U648 ( .Z(GFlen[1]));
Q_RDN U649 ( .Z(GFlen[2]));
Q_RDN U650 ( .Z(GFlen[3]));
Q_RDN U651 ( .Z(GFlen[4]));
Q_RDN U652 ( .Z(GFlen[5]));
Q_RDN U653 ( .Z(GFlen[6]));
Q_RDN U654 ( .Z(GFlen[7]));
Q_RDN U655 ( .Z(GFlen[8]));
Q_RDN U656 ( .Z(GFlen[9]));
Q_RDN U657 ( .Z(GFlen[10]));
Q_RDN U658 ( .Z(GFlen[11]));
Q_RDN U659 ( .Z(GFcbid[0]));
Q_RDN U660 ( .Z(GFcbid[1]));
Q_RDN U661 ( .Z(GFcbid[2]));
Q_RDN U662 ( .Z(GFcbid[3]));
Q_RDN U663 ( .Z(GFcbid[4]));
Q_RDN U664 ( .Z(GFcbid[5]));
Q_RDN U665 ( .Z(GFcbid[6]));
Q_RDN U666 ( .Z(GFcbid[7]));
Q_RDN U667 ( .Z(GFcbid[8]));
Q_RDN U668 ( .Z(GFcbid[9]));
Q_RDN U669 ( .Z(GFcbid[10]));
Q_RDN U670 ( .Z(GFcbid[11]));
Q_RDN U671 ( .Z(GFcbid[12]));
Q_RDN U672 ( .Z(GFcbid[13]));
Q_RDN U673 ( .Z(GFcbid[14]));
Q_RDN U674 ( .Z(GFcbid[15]));
Q_RDN U675 ( .Z(GFcbid[16]));
Q_RDN U676 ( .Z(GFcbid[17]));
Q_RDN U677 ( .Z(GFcbid[18]));
Q_RDN U678 ( .Z(GFcbid[19]));
Q_BUFZP U679 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[0]));
Q_BUFZP U680 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[1]));
Q_BUFZP U681 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[2]));
Q_BUFZP U682 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[3]));
Q_BUFZP U683 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[4]));
Q_BUFZP U684 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[5]));
Q_BUFZP U685 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[6]));
Q_BUFZP U686 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[7]));
Q_BUFZP U687 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[8]));
Q_BUFZP U688 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[9]));
Q_BUFZP U689 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[10]));
Q_BUFZP U690 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[11]));
Q_BUFZP U691 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[12]));
Q_BUFZP U692 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[13]));
Q_BUFZP U693 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[14]));
Q_BUFZP U694 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[15]));
Q_BUFZP U695 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[16]));
Q_BUFZP U696 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[17]));
Q_BUFZP U697 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[18]));
Q_BUFZP U698 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[19]));
Q_BUFZP U699 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[20]));
Q_BUFZP U700 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[21]));
Q_BUFZP U701 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[22]));
Q_BUFZP U702 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[23]));
Q_BUFZP U703 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[24]));
Q_BUFZP U704 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[25]));
Q_BUFZP U705 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[26]));
Q_BUFZP U706 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[27]));
Q_BUFZP U707 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[28]));
Q_BUFZP U708 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[29]));
Q_BUFZP U709 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[30]));
Q_BUFZP U710 ( .OE(GFtsAdd), .A(n3317), .Z(GFidata[31]));
Q_BUFZP U711 ( .OE(GFtsAdd), .A(n3317), .Z(GFcbid[0]));
Q_BUFZP U712 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[1]));
Q_BUFZP U713 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[2]));
Q_BUFZP U714 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[3]));
Q_BUFZP U715 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[4]));
Q_BUFZP U716 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[5]));
Q_BUFZP U717 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[6]));
Q_BUFZP U718 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[7]));
Q_BUFZP U719 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[8]));
Q_BUFZP U720 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[9]));
Q_BUFZP U721 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[10]));
Q_BUFZP U722 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[11]));
Q_BUFZP U723 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[12]));
Q_BUFZP U724 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[13]));
Q_BUFZP U725 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[14]));
Q_BUFZP U726 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[15]));
Q_BUFZP U727 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[16]));
Q_BUFZP U728 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[17]));
Q_BUFZP U729 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[18]));
Q_BUFZP U730 ( .OE(GFtsAdd), .A(n3318), .Z(GFcbid[19]));
Q_BUFZP U731 ( .OE(GFtsAdd), .A(n3318), .Z(GFlen[0]));
Q_BUFZP U732 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[1]));
Q_BUFZP U733 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[2]));
Q_BUFZP U734 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[3]));
Q_BUFZP U735 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[4]));
Q_BUFZP U736 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[5]));
Q_BUFZP U737 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[6]));
Q_BUFZP U738 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[7]));
Q_BUFZP U739 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[8]));
Q_BUFZP U740 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[9]));
Q_BUFZP U741 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[10]));
Q_BUFZP U742 ( .OE(GFtsAdd), .A(n3317), .Z(GFlen[11]));
Q_INV U743 ( .A(ofifoAddr0N[0]), .Z(ofifoAddr1N[0]));
Q_AD01HF U744 ( .A0(ofifoAddr0N[3]), .B0(n3316), .S(ofifoAddr1N[3]), .CO(n3315));
Q_AD01HF U745 ( .A0(ofifoAddr0N[4]), .B0(n3315), .S(ofifoAddr1N[4]), .CO(n3314));
Q_AD01HF U746 ( .A0(ofifoAddr0N[5]), .B0(n3314), .S(ofifoAddr1N[5]), .CO(n3313));
Q_AD01HF U747 ( .A0(ofifoAddr0N[6]), .B0(n3313), .S(ofifoAddr1N[6]), .CO(n3312));
Q_AD01HF U748 ( .A0(ofifoAddr0N[7]), .B0(n3312), .S(ofifoAddr1N[7]), .CO(n3311));
Q_AD01HF U749 ( .A0(ofifoAddr0N[8]), .B0(n3311), .S(ofifoAddr1N[8]), .CO(n3310));
Q_AD01HF U750 ( .A0(ofifoAddr0N[9]), .B0(n3310), .S(ofifoAddr1N[9]), .CO(n3309));
Q_AD01HF U751 ( .A0(ofifoAddr0N[10]), .B0(n3309), .S(ofifoAddr1N[10]), .CO(n3308));
Q_AD01HF U752 ( .A0(ofifoAddr0N[11]), .B0(n3308), .S(ofifoAddr1N[11]), .CO(n3307));
Q_AD01HF U753 ( .A0(ofifoAddr0N[12]), .B0(n3307), .S(ofifoAddr1N[12]), .CO(n3306));
Q_AD01HF U754 ( .A0(ofifoAddr0N[13]), .B0(n3306), .S(ofifoAddr1N[13]), .CO(n3305));
Q_AD01HF U755 ( .A0(ofifoAddr0N[14]), .B0(n3305), .S(ofifoAddr1N[14]), .CO(n3304));
Q_AD01HF U756 ( .A0(ofifoAddr0N[15]), .B0(n3304), .S(ofifoAddr1N[15]), .CO(n3303));
Q_XOR2 U757 ( .A0(ofifoAddr0N[16]), .A1(n3303), .Z(ofifoAddr1N[16]));
Q_INV U758 ( .A(ofifoAddr0N[1]), .Z(ofifoAddr2N[1]));
Q_AD01HF U759 ( .A0(ofifoAddr0N[3]), .B0(n3302), .S(ofifoAddr2N[3]), .CO(n3301));
Q_AD01HF U760 ( .A0(ofifoAddr0N[4]), .B0(n3301), .S(ofifoAddr2N[4]), .CO(n3300));
Q_AD01HF U761 ( .A0(ofifoAddr0N[5]), .B0(n3300), .S(ofifoAddr2N[5]), .CO(n3299));
Q_AD01HF U762 ( .A0(ofifoAddr0N[6]), .B0(n3299), .S(ofifoAddr2N[6]), .CO(n3298));
Q_AD01HF U763 ( .A0(ofifoAddr0N[7]), .B0(n3298), .S(ofifoAddr2N[7]), .CO(n3297));
Q_AD01HF U764 ( .A0(ofifoAddr0N[8]), .B0(n3297), .S(ofifoAddr2N[8]), .CO(n3296));
Q_AD01HF U765 ( .A0(ofifoAddr0N[9]), .B0(n3296), .S(ofifoAddr2N[9]), .CO(n3295));
Q_AD01HF U766 ( .A0(ofifoAddr0N[10]), .B0(n3295), .S(ofifoAddr2N[10]), .CO(n3294));
Q_AD01HF U767 ( .A0(ofifoAddr0N[11]), .B0(n3294), .S(ofifoAddr2N[11]), .CO(n3293));
Q_AD01HF U768 ( .A0(ofifoAddr0N[12]), .B0(n3293), .S(ofifoAddr2N[12]), .CO(n3292));
Q_AD01HF U769 ( .A0(ofifoAddr0N[13]), .B0(n3292), .S(ofifoAddr2N[13]), .CO(n3291));
Q_AD01HF U770 ( .A0(ofifoAddr0N[14]), .B0(n3291), .S(ofifoAddr2N[14]), .CO(n3290));
Q_AD01HF U771 ( .A0(ofifoAddr0N[15]), .B0(n3290), .S(ofifoAddr2N[15]), .CO(n3289));
Q_XOR2 U772 ( .A0(ofifoAddr0N[16]), .A1(n3289), .Z(ofifoAddr2N[16]));
Q_AD01HF U773 ( .A0(ofifoAddr0N[3]), .B0(n3288), .S(ofifoAddr3N[3]), .CO(n3287));
Q_AD01HF U774 ( .A0(ofifoAddr0N[4]), .B0(n3287), .S(ofifoAddr3N[4]), .CO(n3286));
Q_AD01HF U775 ( .A0(ofifoAddr0N[5]), .B0(n3286), .S(ofifoAddr3N[5]), .CO(n3285));
Q_AD01HF U776 ( .A0(ofifoAddr0N[6]), .B0(n3285), .S(ofifoAddr3N[6]), .CO(n3284));
Q_AD01HF U777 ( .A0(ofifoAddr0N[7]), .B0(n3284), .S(ofifoAddr3N[7]), .CO(n3283));
Q_AD01HF U778 ( .A0(ofifoAddr0N[8]), .B0(n3283), .S(ofifoAddr3N[8]), .CO(n3282));
Q_AD01HF U779 ( .A0(ofifoAddr0N[9]), .B0(n3282), .S(ofifoAddr3N[9]), .CO(n3281));
Q_AD01HF U780 ( .A0(ofifoAddr0N[10]), .B0(n3281), .S(ofifoAddr3N[10]), .CO(n3280));
Q_AD01HF U781 ( .A0(ofifoAddr0N[11]), .B0(n3280), .S(ofifoAddr3N[11]), .CO(n3279));
Q_AD01HF U782 ( .A0(ofifoAddr0N[12]), .B0(n3279), .S(ofifoAddr3N[12]), .CO(n3278));
Q_AD01HF U783 ( .A0(ofifoAddr0N[13]), .B0(n3278), .S(ofifoAddr3N[13]), .CO(n3277));
Q_AD01HF U784 ( .A0(ofifoAddr0N[14]), .B0(n3277), .S(ofifoAddr3N[14]), .CO(n3276));
Q_AD01HF U785 ( .A0(ofifoAddr0N[15]), .B0(n3276), .S(ofifoAddr3N[15]), .CO(n3275));
Q_XOR2 U786 ( .A0(ofifoAddr0N[16]), .A1(n3275), .Z(ofifoAddr3N[16]));
Q_INV U787 ( .A(ofifoAddr0N[2]), .Z(ofifoAddr4N[2]));
Q_AD01HF U788 ( .A0(ofifoAddr0N[3]), .B0(ofifoAddr0N[2]), .S(ofifoAddr4N[3]), .CO(n3274));
Q_AD01HF U789 ( .A0(ofifoAddr0N[4]), .B0(n3274), .S(ofifoAddr4N[4]), .CO(n3273));
Q_AD01HF U790 ( .A0(ofifoAddr0N[5]), .B0(n3273), .S(ofifoAddr4N[5]), .CO(n3272));
Q_AD01HF U791 ( .A0(ofifoAddr0N[6]), .B0(n3272), .S(ofifoAddr4N[6]), .CO(n3271));
Q_AD01HF U792 ( .A0(ofifoAddr0N[7]), .B0(n3271), .S(ofifoAddr4N[7]), .CO(n3270));
Q_AD01HF U793 ( .A0(ofifoAddr0N[8]), .B0(n3270), .S(ofifoAddr4N[8]), .CO(n3269));
Q_AD01HF U794 ( .A0(ofifoAddr0N[9]), .B0(n3269), .S(ofifoAddr4N[9]), .CO(n3268));
Q_AD01HF U795 ( .A0(ofifoAddr0N[10]), .B0(n3268), .S(ofifoAddr4N[10]), .CO(n3267));
Q_AD01HF U796 ( .A0(ofifoAddr0N[11]), .B0(n3267), .S(ofifoAddr4N[11]), .CO(n3266));
Q_AD01HF U797 ( .A0(ofifoAddr0N[12]), .B0(n3266), .S(ofifoAddr4N[12]), .CO(n3265));
Q_AD01HF U798 ( .A0(ofifoAddr0N[13]), .B0(n3265), .S(ofifoAddr4N[13]), .CO(n3264));
Q_AD01HF U799 ( .A0(ofifoAddr0N[14]), .B0(n3264), .S(ofifoAddr4N[14]), .CO(n3263));
Q_AD01HF U800 ( .A0(ofifoAddr0N[15]), .B0(n3263), .S(ofifoAddr4N[15]), .CO(n3262));
Q_XOR2 U801 ( .A0(ofifoAddr0N[16]), .A1(n3262), .Z(ofifoAddr4N[16]));
Q_XNR2 U802 ( .A0(ofifoAddr0N[2]), .A1(n3261), .Z(ofifoAddr5N[2]));
Q_OR02 U803 ( .A0(ofifoAddr0N[2]), .A1(n3261), .Z(n3260));
Q_AD01HF U804 ( .A0(ofifoAddr0N[3]), .B0(n3260), .S(ofifoAddr5N[3]), .CO(n3259));
Q_AD01HF U805 ( .A0(ofifoAddr0N[4]), .B0(n3259), .S(ofifoAddr5N[4]), .CO(n3258));
Q_AD01HF U806 ( .A0(ofifoAddr0N[5]), .B0(n3258), .S(ofifoAddr5N[5]), .CO(n3257));
Q_AD01HF U807 ( .A0(ofifoAddr0N[6]), .B0(n3257), .S(ofifoAddr5N[6]), .CO(n3256));
Q_AD01HF U808 ( .A0(ofifoAddr0N[7]), .B0(n3256), .S(ofifoAddr5N[7]), .CO(n3255));
Q_AD01HF U809 ( .A0(ofifoAddr0N[8]), .B0(n3255), .S(ofifoAddr5N[8]), .CO(n3254));
Q_AD01HF U810 ( .A0(ofifoAddr0N[9]), .B0(n3254), .S(ofifoAddr5N[9]), .CO(n3253));
Q_AD01HF U811 ( .A0(ofifoAddr0N[10]), .B0(n3253), .S(ofifoAddr5N[10]), .CO(n3252));
Q_AD01HF U812 ( .A0(ofifoAddr0N[11]), .B0(n3252), .S(ofifoAddr5N[11]), .CO(n3251));
Q_AD01HF U813 ( .A0(ofifoAddr0N[12]), .B0(n3251), .S(ofifoAddr5N[12]), .CO(n3250));
Q_AD01HF U814 ( .A0(ofifoAddr0N[13]), .B0(n3250), .S(ofifoAddr5N[13]), .CO(n3249));
Q_AD01HF U815 ( .A0(ofifoAddr0N[14]), .B0(n3249), .S(ofifoAddr5N[14]), .CO(n3248));
Q_AD01HF U816 ( .A0(ofifoAddr0N[15]), .B0(n3248), .S(ofifoAddr5N[15]), .CO(n3247));
Q_XOR2 U817 ( .A0(ofifoAddr0N[16]), .A1(n3247), .Z(ofifoAddr5N[16]));
Q_XNR2 U818 ( .A0(ofifoAddr0N[2]), .A1(ofifoAddr0N[1]), .Z(ofifoAddr6N[2]));
Q_OR02 U819 ( .A0(ofifoAddr0N[2]), .A1(ofifoAddr0N[1]), .Z(n3246));
Q_AD01HF U820 ( .A0(ofifoAddr0N[3]), .B0(n3246), .S(ofifoAddr6N[3]), .CO(n3245));
Q_AD01HF U821 ( .A0(ofifoAddr0N[4]), .B0(n3245), .S(ofifoAddr6N[4]), .CO(n3244));
Q_AD01HF U822 ( .A0(ofifoAddr0N[5]), .B0(n3244), .S(ofifoAddr6N[5]), .CO(n3243));
Q_AD01HF U823 ( .A0(ofifoAddr0N[6]), .B0(n3243), .S(ofifoAddr6N[6]), .CO(n3242));
Q_AD01HF U824 ( .A0(ofifoAddr0N[7]), .B0(n3242), .S(ofifoAddr6N[7]), .CO(n3241));
Q_AD01HF U825 ( .A0(ofifoAddr0N[8]), .B0(n3241), .S(ofifoAddr6N[8]), .CO(n3240));
Q_AD01HF U826 ( .A0(ofifoAddr0N[9]), .B0(n3240), .S(ofifoAddr6N[9]), .CO(n3239));
Q_AD01HF U827 ( .A0(ofifoAddr0N[10]), .B0(n3239), .S(ofifoAddr6N[10]), .CO(n3238));
Q_AD01HF U828 ( .A0(ofifoAddr0N[11]), .B0(n3238), .S(ofifoAddr6N[11]), .CO(n3237));
Q_AD01HF U829 ( .A0(ofifoAddr0N[12]), .B0(n3237), .S(ofifoAddr6N[12]), .CO(n3236));
Q_AD01HF U830 ( .A0(ofifoAddr0N[13]), .B0(n3236), .S(ofifoAddr6N[13]), .CO(n3235));
Q_AD01HF U831 ( .A0(ofifoAddr0N[14]), .B0(n3235), .S(ofifoAddr6N[14]), .CO(n3234));
Q_AD01HF U832 ( .A0(ofifoAddr0N[15]), .B0(n3234), .S(ofifoAddr6N[15]), .CO(n3233));
Q_XOR2 U833 ( .A0(ofifoAddr0N[16]), .A1(n3233), .Z(ofifoAddr6N[16]));
Q_XNR2 U834 ( .A0(ofifoAddr0N[1]), .A1(ofifoAddr0N[0]), .Z(ofifoAddr3N[1]));
Q_OR02 U835 ( .A0(ofifoAddr0N[1]), .A1(ofifoAddr0N[0]), .Z(n3232));
Q_XNR2 U836 ( .A0(ofifoAddr0N[2]), .A1(n3232), .Z(ofifoAddr7N[2]));
Q_OR02 U837 ( .A0(ofifoAddr0N[2]), .A1(n3232), .Z(n3231));
Q_AD01HF U838 ( .A0(ofifoAddr0N[3]), .B0(n3231), .S(ofifoAddr7N[3]), .CO(n3230));
Q_AD01HF U839 ( .A0(ofifoAddr0N[4]), .B0(n3230), .S(ofifoAddr7N[4]), .CO(n3229));
Q_AD01HF U840 ( .A0(ofifoAddr0N[5]), .B0(n3229), .S(ofifoAddr7N[5]), .CO(n3228));
Q_AD01HF U841 ( .A0(ofifoAddr0N[6]), .B0(n3228), .S(ofifoAddr7N[6]), .CO(n3227));
Q_AD01HF U842 ( .A0(ofifoAddr0N[7]), .B0(n3227), .S(ofifoAddr7N[7]), .CO(n3226));
Q_AD01HF U843 ( .A0(ofifoAddr0N[8]), .B0(n3226), .S(ofifoAddr7N[8]), .CO(n3225));
Q_AD01HF U844 ( .A0(ofifoAddr0N[9]), .B0(n3225), .S(ofifoAddr7N[9]), .CO(n3224));
Q_AD01HF U845 ( .A0(ofifoAddr0N[10]), .B0(n3224), .S(ofifoAddr7N[10]), .CO(n3223));
Q_AD01HF U846 ( .A0(ofifoAddr0N[11]), .B0(n3223), .S(ofifoAddr7N[11]), .CO(n3222));
Q_AD01HF U847 ( .A0(ofifoAddr0N[12]), .B0(n3222), .S(ofifoAddr7N[12]), .CO(n3221));
Q_AD01HF U848 ( .A0(ofifoAddr0N[13]), .B0(n3221), .S(ofifoAddr7N[13]), .CO(n3220));
Q_AD01HF U849 ( .A0(ofifoAddr0N[14]), .B0(n3220), .S(ofifoAddr7N[14]), .CO(n3219));
Q_AD01HF U850 ( .A0(ofifoAddr0N[15]), .B0(n3219), .S(ofifoAddr7N[15]), .CO(n3218));
Q_XOR2 U851 ( .A0(ofifoAddr0N[16]), .A1(n3218), .Z(ofifoAddr7N[16]));
Q_INV U852 ( .A(ofifoAddr0N[3]), .Z(ofifoAddr8N[3]));
Q_AD01HF U853 ( .A0(ofifoAddr0N[4]), .B0(ofifoAddr0N[3]), .S(ofifoAddr8N[4]), .CO(n3217));
Q_AD01HF U854 ( .A0(ofifoAddr0N[5]), .B0(n3217), .S(ofifoAddr8N[5]), .CO(n3216));
Q_AD01HF U855 ( .A0(ofifoAddr0N[6]), .B0(n3216), .S(ofifoAddr8N[6]), .CO(n3215));
Q_AD01HF U856 ( .A0(ofifoAddr0N[7]), .B0(n3215), .S(ofifoAddr8N[7]), .CO(n3214));
Q_AD01HF U857 ( .A0(ofifoAddr0N[8]), .B0(n3214), .S(ofifoAddr8N[8]), .CO(n3213));
Q_AD01HF U858 ( .A0(ofifoAddr0N[9]), .B0(n3213), .S(ofifoAddr8N[9]), .CO(n3212));
Q_AD01HF U859 ( .A0(ofifoAddr0N[10]), .B0(n3212), .S(ofifoAddr8N[10]), .CO(n3211));
Q_AD01HF U860 ( .A0(ofifoAddr0N[11]), .B0(n3211), .S(ofifoAddr8N[11]), .CO(n3210));
Q_AD01HF U861 ( .A0(ofifoAddr0N[12]), .B0(n3210), .S(ofifoAddr8N[12]), .CO(n3209));
Q_AD01HF U862 ( .A0(ofifoAddr0N[13]), .B0(n3209), .S(ofifoAddr8N[13]), .CO(n3208));
Q_AD01HF U863 ( .A0(ofifoAddr0N[14]), .B0(n3208), .S(ofifoAddr8N[14]), .CO(n3207));
Q_AD01HF U864 ( .A0(ofifoAddr0N[15]), .B0(n3207), .S(ofifoAddr8N[15]), .CO(n3206));
Q_XOR2 U865 ( .A0(ofifoAddr0N[16]), .A1(n3206), .Z(ofifoAddr8N[16]));
Q_AN02 U866 ( .A0(n2642), .A1(oFill[1]), .Z(index[6]));
Q_AN02 U867 ( .A0(n2642), .A1(oFill[2]), .Z(index[7]));
Q_AN02 U868 ( .A0(n2642), .A1(oFill[3]), .Z(index[8]));
Q_AN02 U869 ( .A0(n2642), .A1(oFill[4]), .Z(index[9]));
Q_AD01HF U870 ( .A0(oFill[0]), .B0(writeLen[0]), .S(oFillN[0]), .CO(n3205));
Q_AD01HF U871 ( .A0(writeLen[1]), .B0(n3205), .S(oFillN[1]), .CO(n3204));
Q_AD01HF U872 ( .A0(writeLen[2]), .B0(n3204), .S(oFillN[2]), .CO(n3203));
Q_AD01HF U873 ( .A0(writeLen[3]), .B0(n3203), .S(oFillN[3]), .CO(n3202));
Q_AD01HF U874 ( .A0(ofifoAddr0N[0]), .B0(oFillN[1]), .S(ofifoWptrN[0]), .CO(n3201));
Q_AD01 U875 ( .CI(oFillN[2]), .A0(ofifoAddr0N[1]), .B0(n3201), .S(ofifoWptrN[1]), .CO(n3200));
Q_AD02 U876 ( .CI(n3200), .A0(ofifoAddr0N[2]), .A1(ofifoAddr0N[3]), .B0(oFillN[3]), .B1(oFillN[4]), .S0(ofifoWptrN[2]), .S1(ofifoWptrN[3]), .CO(n3199));
Q_AD01HF U877 ( .A0(ofifoAddr0N[4]), .B0(n3199), .S(ofifoWptrN[4]), .CO(n3198));
Q_AD01HF U878 ( .A0(ofifoAddr0N[5]), .B0(n3198), .S(ofifoWptrN[5]), .CO(n3197));
Q_AD01HF U879 ( .A0(ofifoAddr0N[6]), .B0(n3197), .S(ofifoWptrN[6]), .CO(n3196));
Q_AD01HF U880 ( .A0(ofifoAddr0N[7]), .B0(n3196), .S(ofifoWptrN[7]), .CO(n3195));
Q_AD01HF U881 ( .A0(ofifoAddr0N[8]), .B0(n3195), .S(ofifoWptrN[8]), .CO(n3194));
Q_AD01HF U882 ( .A0(ofifoAddr0N[9]), .B0(n3194), .S(ofifoWptrN[9]), .CO(n3193));
Q_AD01HF U883 ( .A0(ofifoAddr0N[10]), .B0(n3193), .S(ofifoWptrN[10]), .CO(n3192));
Q_AD01HF U884 ( .A0(ofifoAddr0N[11]), .B0(n3192), .S(ofifoWptrN[11]), .CO(n3191));
Q_AD01HF U885 ( .A0(ofifoAddr0N[12]), .B0(n3191), .S(ofifoWptrN[12]), .CO(n3190));
Q_AD01HF U886 ( .A0(ofifoAddr0N[13]), .B0(n3190), .S(ofifoWptrN[13]), .CO(n3189));
Q_AD01HF U887 ( .A0(ofifoAddr0N[14]), .B0(n3189), .S(ofifoWptrN[14]), .CO(n3188));
Q_AD01HF U888 ( .A0(ofifoAddr0N[15]), .B0(n3188), .S(ofifoWptrN[15]), .CO(n3187));
Q_XOR2 U889 ( .A0(ofifoAddr0N[16]), .A1(n3187), .Z(ofifoWptrN[16]));
Q_AN02 U890 ( .A0(n2641), .A1(xdata[0]), .Z(n3186));
Q_MX02 U891 ( .S(n2642), .A0(n3186), .A1(n63), .Z(ofifoDataN[0]));
Q_AN02 U892 ( .A0(n2641), .A1(xdata[1]), .Z(n3185));
Q_MX02 U893 ( .S(n2642), .A0(n3185), .A1(n61), .Z(ofifoDataN[1]));
Q_AN02 U894 ( .A0(n2641), .A1(xdata[2]), .Z(n3184));
Q_MX02 U895 ( .S(n2642), .A0(n3184), .A1(n59), .Z(ofifoDataN[2]));
Q_AN02 U896 ( .A0(n2641), .A1(xdata[3]), .Z(n3183));
Q_MX02 U897 ( .S(n2642), .A0(n3183), .A1(n57), .Z(ofifoDataN[3]));
Q_AN02 U898 ( .A0(n2641), .A1(xdata[4]), .Z(n3182));
Q_MX02 U899 ( .S(n2642), .A0(n3182), .A1(n55), .Z(ofifoDataN[4]));
Q_AN02 U900 ( .A0(n2641), .A1(xdata[5]), .Z(n3181));
Q_MX02 U901 ( .S(n2642), .A0(n3181), .A1(n53), .Z(ofifoDataN[5]));
Q_AN02 U902 ( .A0(n2641), .A1(xdata[6]), .Z(n3180));
Q_MX02 U903 ( .S(n2642), .A0(n3180), .A1(n51), .Z(ofifoDataN[6]));
Q_AN02 U904 ( .A0(n2641), .A1(xdata[7]), .Z(n3179));
Q_MX02 U905 ( .S(n2642), .A0(n3179), .A1(n49), .Z(ofifoDataN[7]));
Q_AN02 U906 ( .A0(n2641), .A1(xdata[8]), .Z(n3178));
Q_MX02 U907 ( .S(n2642), .A0(n3178), .A1(n47), .Z(ofifoDataN[8]));
Q_AN02 U908 ( .A0(n2641), .A1(xdata[9]), .Z(n3177));
Q_MX02 U909 ( .S(n2642), .A0(n3177), .A1(n45), .Z(ofifoDataN[9]));
Q_AN02 U910 ( .A0(n2641), .A1(xdata[10]), .Z(n3176));
Q_MX02 U911 ( .S(n2642), .A0(n3176), .A1(n43), .Z(ofifoDataN[10]));
Q_AN02 U912 ( .A0(n2641), .A1(xdata[11]), .Z(n3175));
Q_MX02 U913 ( .S(n2642), .A0(n3175), .A1(n41), .Z(ofifoDataN[11]));
Q_AN02 U914 ( .A0(n2641), .A1(xdata[12]), .Z(n3174));
Q_MX02 U915 ( .S(n2642), .A0(n3174), .A1(n39), .Z(ofifoDataN[12]));
Q_AN02 U916 ( .A0(n2641), .A1(xdata[13]), .Z(n3173));
Q_MX02 U917 ( .S(n2642), .A0(n3173), .A1(n37), .Z(ofifoDataN[13]));
Q_AN02 U918 ( .A0(n2641), .A1(xdata[14]), .Z(n3172));
Q_MX02 U919 ( .S(n2642), .A0(n3172), .A1(n35), .Z(ofifoDataN[14]));
Q_AN02 U920 ( .A0(n2641), .A1(xdata[15]), .Z(n3171));
Q_MX02 U921 ( .S(n2642), .A0(n3171), .A1(n33), .Z(ofifoDataN[15]));
Q_AN02 U922 ( .A0(n2641), .A1(xdata[16]), .Z(n3170));
Q_MX02 U923 ( .S(n2642), .A0(n3170), .A1(n31), .Z(ofifoDataN[16]));
Q_AN02 U924 ( .A0(n2641), .A1(xdata[17]), .Z(n3169));
Q_MX02 U925 ( .S(n2642), .A0(n3169), .A1(n29), .Z(ofifoDataN[17]));
Q_AN02 U926 ( .A0(n2641), .A1(xdata[18]), .Z(n3168));
Q_MX02 U927 ( .S(n2642), .A0(n3168), .A1(n27), .Z(ofifoDataN[18]));
Q_AN02 U928 ( .A0(n2641), .A1(xdata[19]), .Z(n3167));
Q_MX02 U929 ( .S(n2642), .A0(n3167), .A1(n25), .Z(ofifoDataN[19]));
Q_AN02 U930 ( .A0(n2641), .A1(xdata[20]), .Z(n3166));
Q_MX02 U931 ( .S(n2642), .A0(n3166), .A1(n23), .Z(ofifoDataN[20]));
Q_AN02 U932 ( .A0(n2641), .A1(xdata[21]), .Z(n3165));
Q_MX02 U933 ( .S(n2642), .A0(n3165), .A1(n21), .Z(ofifoDataN[21]));
Q_AN02 U934 ( .A0(n2641), .A1(xdata[22]), .Z(n3164));
Q_MX02 U935 ( .S(n2642), .A0(n3164), .A1(n19), .Z(ofifoDataN[22]));
Q_AN02 U936 ( .A0(n2641), .A1(xdata[23]), .Z(n3163));
Q_MX02 U937 ( .S(n2642), .A0(n3163), .A1(n17), .Z(ofifoDataN[23]));
Q_AN02 U938 ( .A0(n2641), .A1(xdata[24]), .Z(n3162));
Q_MX02 U939 ( .S(n2642), .A0(n3162), .A1(n15), .Z(ofifoDataN[24]));
Q_AN02 U940 ( .A0(n2641), .A1(xdata[25]), .Z(n3161));
Q_MX02 U941 ( .S(n2642), .A0(n3161), .A1(n13), .Z(ofifoDataN[25]));
Q_AN02 U942 ( .A0(n2641), .A1(xdata[26]), .Z(n3160));
Q_MX02 U943 ( .S(n2642), .A0(n3160), .A1(n11), .Z(ofifoDataN[26]));
Q_AN02 U944 ( .A0(n2641), .A1(xdata[27]), .Z(n3159));
Q_MX02 U945 ( .S(n2642), .A0(n3159), .A1(n9), .Z(ofifoDataN[27]));
Q_AN02 U946 ( .A0(n2641), .A1(xdata[28]), .Z(n3158));
Q_MX02 U947 ( .S(n2642), .A0(n3158), .A1(n7), .Z(ofifoDataN[28]));
Q_AN02 U948 ( .A0(n2641), .A1(xdata[29]), .Z(n3157));
Q_MX02 U949 ( .S(n2642), .A0(n3157), .A1(n5), .Z(ofifoDataN[29]));
Q_AN02 U950 ( .A0(n2641), .A1(xdata[30]), .Z(n3156));
Q_MX02 U951 ( .S(n2642), .A0(n3156), .A1(n3), .Z(ofifoDataN[30]));
Q_AN02 U952 ( .A0(n2641), .A1(xdata[31]), .Z(n3155));
Q_MX02 U953 ( .S(n2642), .A0(n3155), .A1(n1), .Z(ofifoDataN[31]));
Q_AN02 U954 ( .A0(n2641), .A1(xdata[32]), .Z(n3154));
Q_MX02 U955 ( .S(n2642), .A0(n3154), .A1(xdata[0]), .Z(ofifoDataN[32]));
Q_AN02 U956 ( .A0(n2641), .A1(xdata[33]), .Z(n3153));
Q_MX02 U957 ( .S(n2642), .A0(n3153), .A1(xdata[1]), .Z(ofifoDataN[33]));
Q_AN02 U958 ( .A0(n2641), .A1(xdata[34]), .Z(n3152));
Q_MX02 U959 ( .S(n2642), .A0(n3152), .A1(xdata[2]), .Z(ofifoDataN[34]));
Q_AN02 U960 ( .A0(n2641), .A1(xdata[35]), .Z(n3151));
Q_MX02 U961 ( .S(n2642), .A0(n3151), .A1(xdata[3]), .Z(ofifoDataN[35]));
Q_AN02 U962 ( .A0(n2641), .A1(xdata[36]), .Z(n3150));
Q_MX02 U963 ( .S(n2642), .A0(n3150), .A1(xdata[4]), .Z(ofifoDataN[36]));
Q_AN02 U964 ( .A0(n2641), .A1(xdata[37]), .Z(n3149));
Q_MX02 U965 ( .S(n2642), .A0(n3149), .A1(xdata[5]), .Z(ofifoDataN[37]));
Q_AN02 U966 ( .A0(n2641), .A1(xdata[38]), .Z(n3148));
Q_MX02 U967 ( .S(n2642), .A0(n3148), .A1(xdata[6]), .Z(ofifoDataN[38]));
Q_AN02 U968 ( .A0(n2641), .A1(xdata[39]), .Z(n3147));
Q_MX02 U969 ( .S(n2642), .A0(n3147), .A1(xdata[7]), .Z(ofifoDataN[39]));
Q_AN02 U970 ( .A0(n2641), .A1(xdata[40]), .Z(n3146));
Q_MX02 U971 ( .S(n2642), .A0(n3146), .A1(xdata[8]), .Z(ofifoDataN[40]));
Q_AN02 U972 ( .A0(n2641), .A1(xdata[41]), .Z(n3145));
Q_MX02 U973 ( .S(n2642), .A0(n3145), .A1(xdata[9]), .Z(ofifoDataN[41]));
Q_AN02 U974 ( .A0(n2641), .A1(xdata[42]), .Z(n3144));
Q_MX02 U975 ( .S(n2642), .A0(n3144), .A1(xdata[10]), .Z(ofifoDataN[42]));
Q_AN02 U976 ( .A0(n2641), .A1(xdata[43]), .Z(n3143));
Q_MX02 U977 ( .S(n2642), .A0(n3143), .A1(xdata[11]), .Z(ofifoDataN[43]));
Q_AN02 U978 ( .A0(n2641), .A1(xdata[44]), .Z(n3142));
Q_MX02 U979 ( .S(n2642), .A0(n3142), .A1(xdata[12]), .Z(ofifoDataN[44]));
Q_AN02 U980 ( .A0(n2641), .A1(xdata[45]), .Z(n3141));
Q_MX02 U981 ( .S(n2642), .A0(n3141), .A1(xdata[13]), .Z(ofifoDataN[45]));
Q_AN02 U982 ( .A0(n2641), .A1(xdata[46]), .Z(n3140));
Q_MX02 U983 ( .S(n2642), .A0(n3140), .A1(xdata[14]), .Z(ofifoDataN[46]));
Q_AN02 U984 ( .A0(n2641), .A1(xdata[47]), .Z(n3139));
Q_MX02 U985 ( .S(n2642), .A0(n3139), .A1(xdata[15]), .Z(ofifoDataN[47]));
Q_AN02 U986 ( .A0(n2641), .A1(xdata[48]), .Z(n3138));
Q_MX02 U987 ( .S(n2642), .A0(n3138), .A1(xdata[16]), .Z(ofifoDataN[48]));
Q_AN02 U988 ( .A0(n2641), .A1(xdata[49]), .Z(n3137));
Q_MX02 U989 ( .S(n2642), .A0(n3137), .A1(xdata[17]), .Z(ofifoDataN[49]));
Q_AN02 U990 ( .A0(n2641), .A1(xdata[50]), .Z(n3136));
Q_MX02 U991 ( .S(n2642), .A0(n3136), .A1(xdata[18]), .Z(ofifoDataN[50]));
Q_AN02 U992 ( .A0(n2641), .A1(xdata[51]), .Z(n3135));
Q_MX02 U993 ( .S(n2642), .A0(n3135), .A1(xdata[19]), .Z(ofifoDataN[51]));
Q_AN02 U994 ( .A0(n2641), .A1(xdata[52]), .Z(n3134));
Q_MX02 U995 ( .S(n2642), .A0(n3134), .A1(xdata[20]), .Z(ofifoDataN[52]));
Q_AN02 U996 ( .A0(n2641), .A1(xdata[53]), .Z(n3133));
Q_MX02 U997 ( .S(n2642), .A0(n3133), .A1(xdata[21]), .Z(ofifoDataN[53]));
Q_AN02 U998 ( .A0(n2641), .A1(xdata[54]), .Z(n3132));
Q_MX02 U999 ( .S(n2642), .A0(n3132), .A1(xdata[22]), .Z(ofifoDataN[54]));
Q_AN02 U1000 ( .A0(n2641), .A1(xdata[55]), .Z(n3131));
Q_MX02 U1001 ( .S(n2642), .A0(n3131), .A1(xdata[23]), .Z(ofifoDataN[55]));
Q_AN02 U1002 ( .A0(n2641), .A1(xdata[56]), .Z(n3130));
Q_MX02 U1003 ( .S(n2642), .A0(n3130), .A1(xdata[24]), .Z(ofifoDataN[56]));
Q_AN02 U1004 ( .A0(n2641), .A1(xdata[57]), .Z(n3129));
Q_MX02 U1005 ( .S(n2642), .A0(n3129), .A1(xdata[25]), .Z(ofifoDataN[57]));
Q_AN02 U1006 ( .A0(n2641), .A1(xdata[58]), .Z(n3128));
Q_MX02 U1007 ( .S(n2642), .A0(n3128), .A1(xdata[26]), .Z(ofifoDataN[58]));
Q_AN02 U1008 ( .A0(n2641), .A1(xdata[59]), .Z(n3127));
Q_MX02 U1009 ( .S(n2642), .A0(n3127), .A1(xdata[27]), .Z(ofifoDataN[59]));
Q_AN02 U1010 ( .A0(n2641), .A1(xdata[60]), .Z(n3126));
Q_MX02 U1011 ( .S(n2642), .A0(n3126), .A1(xdata[28]), .Z(ofifoDataN[60]));
Q_AN02 U1012 ( .A0(n2641), .A1(xdata[61]), .Z(n3125));
Q_MX02 U1013 ( .S(n2642), .A0(n3125), .A1(xdata[29]), .Z(ofifoDataN[61]));
Q_AN02 U1014 ( .A0(n2641), .A1(xdata[62]), .Z(n3124));
Q_MX02 U1015 ( .S(n2642), .A0(n3124), .A1(xdata[30]), .Z(ofifoDataN[62]));
Q_AN02 U1016 ( .A0(n2641), .A1(xdata[63]), .Z(n3123));
Q_MX02 U1017 ( .S(n2642), .A0(n3123), .A1(xdata[31]), .Z(ofifoDataN[63]));
Q_AN02 U1018 ( .A0(n2641), .A1(xdata[64]), .Z(n3122));
Q_MX02 U1019 ( .S(n2642), .A0(n3122), .A1(xdata[32]), .Z(ofifoDataN[64]));
Q_AN02 U1020 ( .A0(n2641), .A1(xdata[65]), .Z(n3121));
Q_MX02 U1021 ( .S(n2642), .A0(n3121), .A1(xdata[33]), .Z(ofifoDataN[65]));
Q_AN02 U1022 ( .A0(n2641), .A1(xdata[66]), .Z(n3120));
Q_MX02 U1023 ( .S(n2642), .A0(n3120), .A1(xdata[34]), .Z(ofifoDataN[66]));
Q_AN02 U1024 ( .A0(n2641), .A1(xdata[67]), .Z(n3119));
Q_MX02 U1025 ( .S(n2642), .A0(n3119), .A1(xdata[35]), .Z(ofifoDataN[67]));
Q_AN02 U1026 ( .A0(n2641), .A1(xdata[68]), .Z(n3118));
Q_MX02 U1027 ( .S(n2642), .A0(n3118), .A1(xdata[36]), .Z(ofifoDataN[68]));
Q_AN02 U1028 ( .A0(n2641), .A1(xdata[69]), .Z(n3117));
Q_MX02 U1029 ( .S(n2642), .A0(n3117), .A1(xdata[37]), .Z(ofifoDataN[69]));
Q_AN02 U1030 ( .A0(n2641), .A1(xdata[70]), .Z(n3116));
Q_MX02 U1031 ( .S(n2642), .A0(n3116), .A1(xdata[38]), .Z(ofifoDataN[70]));
Q_AN02 U1032 ( .A0(n2641), .A1(xdata[71]), .Z(n3115));
Q_MX02 U1033 ( .S(n2642), .A0(n3115), .A1(xdata[39]), .Z(ofifoDataN[71]));
Q_AN02 U1034 ( .A0(n2641), .A1(xdata[72]), .Z(n3114));
Q_MX02 U1035 ( .S(n2642), .A0(n3114), .A1(xdata[40]), .Z(ofifoDataN[72]));
Q_AN02 U1036 ( .A0(n2641), .A1(xdata[73]), .Z(n3113));
Q_MX02 U1037 ( .S(n2642), .A0(n3113), .A1(xdata[41]), .Z(ofifoDataN[73]));
Q_AN02 U1038 ( .A0(n2641), .A1(xdata[74]), .Z(n3112));
Q_MX02 U1039 ( .S(n2642), .A0(n3112), .A1(xdata[42]), .Z(ofifoDataN[74]));
Q_AN02 U1040 ( .A0(n2641), .A1(xdata[75]), .Z(n3111));
Q_MX02 U1041 ( .S(n2642), .A0(n3111), .A1(xdata[43]), .Z(ofifoDataN[75]));
Q_AN02 U1042 ( .A0(n2641), .A1(xdata[76]), .Z(n3110));
Q_MX02 U1043 ( .S(n2642), .A0(n3110), .A1(xdata[44]), .Z(ofifoDataN[76]));
Q_AN02 U1044 ( .A0(n2641), .A1(xdata[77]), .Z(n3109));
Q_MX02 U1045 ( .S(n2642), .A0(n3109), .A1(xdata[45]), .Z(ofifoDataN[77]));
Q_AN02 U1046 ( .A0(n2641), .A1(xdata[78]), .Z(n3108));
Q_MX02 U1047 ( .S(n2642), .A0(n3108), .A1(xdata[46]), .Z(ofifoDataN[78]));
Q_AN02 U1048 ( .A0(n2641), .A1(xdata[79]), .Z(n3107));
Q_MX02 U1049 ( .S(n2642), .A0(n3107), .A1(xdata[47]), .Z(ofifoDataN[79]));
Q_AN02 U1050 ( .A0(n2641), .A1(xdata[80]), .Z(n3106));
Q_MX02 U1051 ( .S(n2642), .A0(n3106), .A1(xdata[48]), .Z(ofifoDataN[80]));
Q_AN02 U1052 ( .A0(n2641), .A1(xdata[81]), .Z(n3105));
Q_MX02 U1053 ( .S(n2642), .A0(n3105), .A1(xdata[49]), .Z(ofifoDataN[81]));
Q_AN02 U1054 ( .A0(n2641), .A1(xdata[82]), .Z(n3104));
Q_MX02 U1055 ( .S(n2642), .A0(n3104), .A1(xdata[50]), .Z(ofifoDataN[82]));
Q_AN02 U1056 ( .A0(n2641), .A1(xdata[83]), .Z(n3103));
Q_MX02 U1057 ( .S(n2642), .A0(n3103), .A1(xdata[51]), .Z(ofifoDataN[83]));
Q_AN02 U1058 ( .A0(n2641), .A1(xdata[84]), .Z(n3102));
Q_MX02 U1059 ( .S(n2642), .A0(n3102), .A1(xdata[52]), .Z(ofifoDataN[84]));
Q_AN02 U1060 ( .A0(n2641), .A1(xdata[85]), .Z(n3101));
Q_MX02 U1061 ( .S(n2642), .A0(n3101), .A1(xdata[53]), .Z(ofifoDataN[85]));
Q_AN02 U1062 ( .A0(n2641), .A1(xdata[86]), .Z(n3100));
Q_MX02 U1063 ( .S(n2642), .A0(n3100), .A1(xdata[54]), .Z(ofifoDataN[86]));
Q_AN02 U1064 ( .A0(n2641), .A1(xdata[87]), .Z(n3099));
Q_MX02 U1065 ( .S(n2642), .A0(n3099), .A1(xdata[55]), .Z(ofifoDataN[87]));
Q_AN02 U1066 ( .A0(n2641), .A1(xdata[88]), .Z(n3098));
Q_MX02 U1067 ( .S(n2642), .A0(n3098), .A1(xdata[56]), .Z(ofifoDataN[88]));
Q_AN02 U1068 ( .A0(n2641), .A1(xdata[89]), .Z(n3097));
Q_MX02 U1069 ( .S(n2642), .A0(n3097), .A1(xdata[57]), .Z(ofifoDataN[89]));
Q_AN02 U1070 ( .A0(n2641), .A1(xdata[90]), .Z(n3096));
Q_MX02 U1071 ( .S(n2642), .A0(n3096), .A1(xdata[58]), .Z(ofifoDataN[90]));
Q_AN02 U1072 ( .A0(n2641), .A1(xdata[91]), .Z(n3095));
Q_MX02 U1073 ( .S(n2642), .A0(n3095), .A1(xdata[59]), .Z(ofifoDataN[91]));
Q_AN02 U1074 ( .A0(n2641), .A1(xdata[92]), .Z(n3094));
Q_MX02 U1075 ( .S(n2642), .A0(n3094), .A1(xdata[60]), .Z(ofifoDataN[92]));
Q_AN02 U1076 ( .A0(n2641), .A1(xdata[93]), .Z(n3093));
Q_MX02 U1077 ( .S(n2642), .A0(n3093), .A1(xdata[61]), .Z(ofifoDataN[93]));
Q_AN02 U1078 ( .A0(n2641), .A1(xdata[94]), .Z(n3092));
Q_MX02 U1079 ( .S(n2642), .A0(n3092), .A1(xdata[62]), .Z(ofifoDataN[94]));
Q_AN02 U1080 ( .A0(n2641), .A1(xdata[95]), .Z(n3091));
Q_MX02 U1081 ( .S(n2642), .A0(n3091), .A1(xdata[63]), .Z(ofifoDataN[95]));
Q_AN02 U1082 ( .A0(n2641), .A1(xdata[96]), .Z(n3090));
Q_MX02 U1083 ( .S(n2642), .A0(n3090), .A1(xdata[64]), .Z(ofifoDataN[96]));
Q_AN02 U1084 ( .A0(n2641), .A1(xdata[97]), .Z(n3089));
Q_MX02 U1085 ( .S(n2642), .A0(n3089), .A1(xdata[65]), .Z(ofifoDataN[97]));
Q_AN02 U1086 ( .A0(n2641), .A1(xdata[98]), .Z(n3088));
Q_MX02 U1087 ( .S(n2642), .A0(n3088), .A1(xdata[66]), .Z(ofifoDataN[98]));
Q_AN02 U1088 ( .A0(n2641), .A1(xdata[99]), .Z(n3087));
Q_MX02 U1089 ( .S(n2642), .A0(n3087), .A1(xdata[67]), .Z(ofifoDataN[99]));
Q_AN02 U1090 ( .A0(n2641), .A1(xdata[100]), .Z(n3086));
Q_MX02 U1091 ( .S(n2642), .A0(n3086), .A1(xdata[68]), .Z(ofifoDataN[100]));
Q_AN02 U1092 ( .A0(n2641), .A1(xdata[101]), .Z(n3085));
Q_MX02 U1093 ( .S(n2642), .A0(n3085), .A1(xdata[69]), .Z(ofifoDataN[101]));
Q_AN02 U1094 ( .A0(n2641), .A1(xdata[102]), .Z(n3084));
Q_MX02 U1095 ( .S(n2642), .A0(n3084), .A1(xdata[70]), .Z(ofifoDataN[102]));
Q_AN02 U1096 ( .A0(n2641), .A1(xdata[103]), .Z(n3083));
Q_MX02 U1097 ( .S(n2642), .A0(n3083), .A1(xdata[71]), .Z(ofifoDataN[103]));
Q_AN02 U1098 ( .A0(n2641), .A1(xdata[104]), .Z(n3082));
Q_MX02 U1099 ( .S(n2642), .A0(n3082), .A1(xdata[72]), .Z(ofifoDataN[104]));
Q_AN02 U1100 ( .A0(n2641), .A1(xdata[105]), .Z(n3081));
Q_MX02 U1101 ( .S(n2642), .A0(n3081), .A1(xdata[73]), .Z(ofifoDataN[105]));
Q_AN02 U1102 ( .A0(n2641), .A1(xdata[106]), .Z(n3080));
Q_MX02 U1103 ( .S(n2642), .A0(n3080), .A1(xdata[74]), .Z(ofifoDataN[106]));
Q_AN02 U1104 ( .A0(n2641), .A1(xdata[107]), .Z(n3079));
Q_MX02 U1105 ( .S(n2642), .A0(n3079), .A1(xdata[75]), .Z(ofifoDataN[107]));
Q_AN02 U1106 ( .A0(n2641), .A1(xdata[108]), .Z(n3078));
Q_MX02 U1107 ( .S(n2642), .A0(n3078), .A1(xdata[76]), .Z(ofifoDataN[108]));
Q_AN02 U1108 ( .A0(n2641), .A1(xdata[109]), .Z(n3077));
Q_MX02 U1109 ( .S(n2642), .A0(n3077), .A1(xdata[77]), .Z(ofifoDataN[109]));
Q_AN02 U1110 ( .A0(n2641), .A1(xdata[110]), .Z(n3076));
Q_MX02 U1111 ( .S(n2642), .A0(n3076), .A1(xdata[78]), .Z(ofifoDataN[110]));
Q_AN02 U1112 ( .A0(n2641), .A1(xdata[111]), .Z(n3075));
Q_MX02 U1113 ( .S(n2642), .A0(n3075), .A1(xdata[79]), .Z(ofifoDataN[111]));
Q_AN02 U1114 ( .A0(n2641), .A1(xdata[112]), .Z(n3074));
Q_MX02 U1115 ( .S(n2642), .A0(n3074), .A1(xdata[80]), .Z(ofifoDataN[112]));
Q_AN02 U1116 ( .A0(n2641), .A1(xdata[113]), .Z(n3073));
Q_MX02 U1117 ( .S(n2642), .A0(n3073), .A1(xdata[81]), .Z(ofifoDataN[113]));
Q_AN02 U1118 ( .A0(n2641), .A1(xdata[114]), .Z(n3072));
Q_MX02 U1119 ( .S(n2642), .A0(n3072), .A1(xdata[82]), .Z(ofifoDataN[114]));
Q_AN02 U1120 ( .A0(n2641), .A1(xdata[115]), .Z(n3071));
Q_MX02 U1121 ( .S(n2642), .A0(n3071), .A1(xdata[83]), .Z(ofifoDataN[115]));
Q_AN02 U1122 ( .A0(n2641), .A1(xdata[116]), .Z(n3070));
Q_MX02 U1123 ( .S(n2642), .A0(n3070), .A1(xdata[84]), .Z(ofifoDataN[116]));
Q_AN02 U1124 ( .A0(n2641), .A1(xdata[117]), .Z(n3069));
Q_MX02 U1125 ( .S(n2642), .A0(n3069), .A1(xdata[85]), .Z(ofifoDataN[117]));
Q_AN02 U1126 ( .A0(n2641), .A1(xdata[118]), .Z(n3068));
Q_MX02 U1127 ( .S(n2642), .A0(n3068), .A1(xdata[86]), .Z(ofifoDataN[118]));
Q_AN02 U1128 ( .A0(n2641), .A1(xdata[119]), .Z(n3067));
Q_MX02 U1129 ( .S(n2642), .A0(n3067), .A1(xdata[87]), .Z(ofifoDataN[119]));
Q_AN02 U1130 ( .A0(n2641), .A1(xdata[120]), .Z(n3066));
Q_MX02 U1131 ( .S(n2642), .A0(n3066), .A1(xdata[88]), .Z(ofifoDataN[120]));
Q_AN02 U1132 ( .A0(n2641), .A1(xdata[121]), .Z(n3065));
Q_MX02 U1133 ( .S(n2642), .A0(n3065), .A1(xdata[89]), .Z(ofifoDataN[121]));
Q_AN02 U1134 ( .A0(n2641), .A1(xdata[122]), .Z(n3064));
Q_MX02 U1135 ( .S(n2642), .A0(n3064), .A1(xdata[90]), .Z(ofifoDataN[122]));
Q_AN02 U1136 ( .A0(n2641), .A1(xdata[123]), .Z(n3063));
Q_MX02 U1137 ( .S(n2642), .A0(n3063), .A1(xdata[91]), .Z(ofifoDataN[123]));
Q_AN02 U1138 ( .A0(n2641), .A1(xdata[124]), .Z(n3062));
Q_MX02 U1139 ( .S(n2642), .A0(n3062), .A1(xdata[92]), .Z(ofifoDataN[124]));
Q_AN02 U1140 ( .A0(n2641), .A1(xdata[125]), .Z(n3061));
Q_MX02 U1141 ( .S(n2642), .A0(n3061), .A1(xdata[93]), .Z(ofifoDataN[125]));
Q_AN02 U1142 ( .A0(n2641), .A1(xdata[126]), .Z(n3060));
Q_MX02 U1143 ( .S(n2642), .A0(n3060), .A1(xdata[94]), .Z(ofifoDataN[126]));
Q_AN02 U1144 ( .A0(n2641), .A1(xdata[127]), .Z(n3059));
Q_MX02 U1145 ( .S(n2642), .A0(n3059), .A1(xdata[95]), .Z(ofifoDataN[127]));
Q_AN02 U1146 ( .A0(n2641), .A1(xdata[128]), .Z(n3058));
Q_MX02 U1147 ( .S(n2642), .A0(n3058), .A1(xdata[96]), .Z(ofifoDataN[128]));
Q_AN02 U1148 ( .A0(n2641), .A1(xdata[129]), .Z(n3057));
Q_MX02 U1149 ( .S(n2642), .A0(n3057), .A1(xdata[97]), .Z(ofifoDataN[129]));
Q_AN02 U1150 ( .A0(n2641), .A1(xdata[130]), .Z(n3056));
Q_MX02 U1151 ( .S(n2642), .A0(n3056), .A1(xdata[98]), .Z(ofifoDataN[130]));
Q_AN02 U1152 ( .A0(n2641), .A1(xdata[131]), .Z(n3055));
Q_MX02 U1153 ( .S(n2642), .A0(n3055), .A1(xdata[99]), .Z(ofifoDataN[131]));
Q_AN02 U1154 ( .A0(n2641), .A1(xdata[132]), .Z(n3054));
Q_MX02 U1155 ( .S(n2642), .A0(n3054), .A1(xdata[100]), .Z(ofifoDataN[132]));
Q_AN02 U1156 ( .A0(n2641), .A1(xdata[133]), .Z(n3053));
Q_MX02 U1157 ( .S(n2642), .A0(n3053), .A1(xdata[101]), .Z(ofifoDataN[133]));
Q_AN02 U1158 ( .A0(n2641), .A1(xdata[134]), .Z(n3052));
Q_MX02 U1159 ( .S(n2642), .A0(n3052), .A1(xdata[102]), .Z(ofifoDataN[134]));
Q_AN02 U1160 ( .A0(n2641), .A1(xdata[135]), .Z(n3051));
Q_MX02 U1161 ( .S(n2642), .A0(n3051), .A1(xdata[103]), .Z(ofifoDataN[135]));
Q_AN02 U1162 ( .A0(n2641), .A1(xdata[136]), .Z(n3050));
Q_MX02 U1163 ( .S(n2642), .A0(n3050), .A1(xdata[104]), .Z(ofifoDataN[136]));
Q_AN02 U1164 ( .A0(n2641), .A1(xdata[137]), .Z(n3049));
Q_MX02 U1165 ( .S(n2642), .A0(n3049), .A1(xdata[105]), .Z(ofifoDataN[137]));
Q_AN02 U1166 ( .A0(n2641), .A1(xdata[138]), .Z(n3048));
Q_MX02 U1167 ( .S(n2642), .A0(n3048), .A1(xdata[106]), .Z(ofifoDataN[138]));
Q_AN02 U1168 ( .A0(n2641), .A1(xdata[139]), .Z(n3047));
Q_MX02 U1169 ( .S(n2642), .A0(n3047), .A1(xdata[107]), .Z(ofifoDataN[139]));
Q_AN02 U1170 ( .A0(n2641), .A1(xdata[140]), .Z(n3046));
Q_MX02 U1171 ( .S(n2642), .A0(n3046), .A1(xdata[108]), .Z(ofifoDataN[140]));
Q_AN02 U1172 ( .A0(n2641), .A1(xdata[141]), .Z(n3045));
Q_MX02 U1173 ( .S(n2642), .A0(n3045), .A1(xdata[109]), .Z(ofifoDataN[141]));
Q_AN02 U1174 ( .A0(n2641), .A1(xdata[142]), .Z(n3044));
Q_MX02 U1175 ( .S(n2642), .A0(n3044), .A1(xdata[110]), .Z(ofifoDataN[142]));
Q_AN02 U1176 ( .A0(n2641), .A1(xdata[143]), .Z(n3043));
Q_MX02 U1177 ( .S(n2642), .A0(n3043), .A1(xdata[111]), .Z(ofifoDataN[143]));
Q_AN02 U1178 ( .A0(n2641), .A1(xdata[144]), .Z(n3042));
Q_MX02 U1179 ( .S(n2642), .A0(n3042), .A1(xdata[112]), .Z(ofifoDataN[144]));
Q_AN02 U1180 ( .A0(n2641), .A1(xdata[145]), .Z(n3041));
Q_MX02 U1181 ( .S(n2642), .A0(n3041), .A1(xdata[113]), .Z(ofifoDataN[145]));
Q_AN02 U1182 ( .A0(n2641), .A1(xdata[146]), .Z(n3040));
Q_MX02 U1183 ( .S(n2642), .A0(n3040), .A1(xdata[114]), .Z(ofifoDataN[146]));
Q_AN02 U1184 ( .A0(n2641), .A1(xdata[147]), .Z(n3039));
Q_MX02 U1185 ( .S(n2642), .A0(n3039), .A1(xdata[115]), .Z(ofifoDataN[147]));
Q_AN02 U1186 ( .A0(n2641), .A1(xdata[148]), .Z(n3038));
Q_MX02 U1187 ( .S(n2642), .A0(n3038), .A1(xdata[116]), .Z(ofifoDataN[148]));
Q_AN02 U1188 ( .A0(n2641), .A1(xdata[149]), .Z(n3037));
Q_MX02 U1189 ( .S(n2642), .A0(n3037), .A1(xdata[117]), .Z(ofifoDataN[149]));
Q_AN02 U1190 ( .A0(n2641), .A1(xdata[150]), .Z(n3036));
Q_MX02 U1191 ( .S(n2642), .A0(n3036), .A1(xdata[118]), .Z(ofifoDataN[150]));
Q_AN02 U1192 ( .A0(n2641), .A1(xdata[151]), .Z(n3035));
Q_MX02 U1193 ( .S(n2642), .A0(n3035), .A1(xdata[119]), .Z(ofifoDataN[151]));
Q_AN02 U1194 ( .A0(n2641), .A1(xdata[152]), .Z(n3034));
Q_MX02 U1195 ( .S(n2642), .A0(n3034), .A1(xdata[120]), .Z(ofifoDataN[152]));
Q_AN02 U1196 ( .A0(n2641), .A1(xdata[153]), .Z(n3033));
Q_MX02 U1197 ( .S(n2642), .A0(n3033), .A1(xdata[121]), .Z(ofifoDataN[153]));
Q_AN02 U1198 ( .A0(n2641), .A1(xdata[154]), .Z(n3032));
Q_MX02 U1199 ( .S(n2642), .A0(n3032), .A1(xdata[122]), .Z(ofifoDataN[154]));
Q_AN02 U1200 ( .A0(n2641), .A1(xdata[155]), .Z(n3031));
Q_MX02 U1201 ( .S(n2642), .A0(n3031), .A1(xdata[123]), .Z(ofifoDataN[155]));
Q_AN02 U1202 ( .A0(n2641), .A1(xdata[156]), .Z(n3030));
Q_MX02 U1203 ( .S(n2642), .A0(n3030), .A1(xdata[124]), .Z(ofifoDataN[156]));
Q_AN02 U1204 ( .A0(n2641), .A1(xdata[157]), .Z(n3029));
Q_MX02 U1205 ( .S(n2642), .A0(n3029), .A1(xdata[125]), .Z(ofifoDataN[157]));
Q_AN02 U1206 ( .A0(n2641), .A1(xdata[158]), .Z(n3028));
Q_MX02 U1207 ( .S(n2642), .A0(n3028), .A1(xdata[126]), .Z(ofifoDataN[158]));
Q_AN02 U1208 ( .A0(n2641), .A1(xdata[159]), .Z(n3027));
Q_MX02 U1209 ( .S(n2642), .A0(n3027), .A1(xdata[127]), .Z(ofifoDataN[159]));
Q_AN02 U1210 ( .A0(n2641), .A1(xdata[160]), .Z(n3026));
Q_MX02 U1211 ( .S(n2642), .A0(n3026), .A1(xdata[128]), .Z(ofifoDataN[160]));
Q_AN02 U1212 ( .A0(n2641), .A1(xdata[161]), .Z(n3025));
Q_MX02 U1213 ( .S(n2642), .A0(n3025), .A1(xdata[129]), .Z(ofifoDataN[161]));
Q_AN02 U1214 ( .A0(n2641), .A1(xdata[162]), .Z(n3024));
Q_MX02 U1215 ( .S(n2642), .A0(n3024), .A1(xdata[130]), .Z(ofifoDataN[162]));
Q_AN02 U1216 ( .A0(n2641), .A1(xdata[163]), .Z(n3023));
Q_MX02 U1217 ( .S(n2642), .A0(n3023), .A1(xdata[131]), .Z(ofifoDataN[163]));
Q_AN02 U1218 ( .A0(n2641), .A1(xdata[164]), .Z(n3022));
Q_MX02 U1219 ( .S(n2642), .A0(n3022), .A1(xdata[132]), .Z(ofifoDataN[164]));
Q_AN02 U1220 ( .A0(n2641), .A1(xdata[165]), .Z(n3021));
Q_MX02 U1221 ( .S(n2642), .A0(n3021), .A1(xdata[133]), .Z(ofifoDataN[165]));
Q_AN02 U1222 ( .A0(n2641), .A1(xdata[166]), .Z(n3020));
Q_MX02 U1223 ( .S(n2642), .A0(n3020), .A1(xdata[134]), .Z(ofifoDataN[166]));
Q_AN02 U1224 ( .A0(n2641), .A1(xdata[167]), .Z(n3019));
Q_MX02 U1225 ( .S(n2642), .A0(n3019), .A1(xdata[135]), .Z(ofifoDataN[167]));
Q_AN02 U1226 ( .A0(n2641), .A1(xdata[168]), .Z(n3018));
Q_MX02 U1227 ( .S(n2642), .A0(n3018), .A1(xdata[136]), .Z(ofifoDataN[168]));
Q_AN02 U1228 ( .A0(n2641), .A1(xdata[169]), .Z(n3017));
Q_MX02 U1229 ( .S(n2642), .A0(n3017), .A1(xdata[137]), .Z(ofifoDataN[169]));
Q_AN02 U1230 ( .A0(n2641), .A1(xdata[170]), .Z(n3016));
Q_MX02 U1231 ( .S(n2642), .A0(n3016), .A1(xdata[138]), .Z(ofifoDataN[170]));
Q_AN02 U1232 ( .A0(n2641), .A1(xdata[171]), .Z(n3015));
Q_MX02 U1233 ( .S(n2642), .A0(n3015), .A1(xdata[139]), .Z(ofifoDataN[171]));
Q_AN02 U1234 ( .A0(n2641), .A1(xdata[172]), .Z(n3014));
Q_MX02 U1235 ( .S(n2642), .A0(n3014), .A1(xdata[140]), .Z(ofifoDataN[172]));
Q_AN02 U1236 ( .A0(n2641), .A1(xdata[173]), .Z(n3013));
Q_MX02 U1237 ( .S(n2642), .A0(n3013), .A1(xdata[141]), .Z(ofifoDataN[173]));
Q_AN02 U1238 ( .A0(n2641), .A1(xdata[174]), .Z(n3012));
Q_MX02 U1239 ( .S(n2642), .A0(n3012), .A1(xdata[142]), .Z(ofifoDataN[174]));
Q_AN02 U1240 ( .A0(n2641), .A1(xdata[175]), .Z(n3011));
Q_MX02 U1241 ( .S(n2642), .A0(n3011), .A1(xdata[143]), .Z(ofifoDataN[175]));
Q_AN02 U1242 ( .A0(n2641), .A1(xdata[176]), .Z(n3010));
Q_MX02 U1243 ( .S(n2642), .A0(n3010), .A1(xdata[144]), .Z(ofifoDataN[176]));
Q_AN02 U1244 ( .A0(n2641), .A1(xdata[177]), .Z(n3009));
Q_MX02 U1245 ( .S(n2642), .A0(n3009), .A1(xdata[145]), .Z(ofifoDataN[177]));
Q_AN02 U1246 ( .A0(n2641), .A1(xdata[178]), .Z(n3008));
Q_MX02 U1247 ( .S(n2642), .A0(n3008), .A1(xdata[146]), .Z(ofifoDataN[178]));
Q_AN02 U1248 ( .A0(n2641), .A1(xdata[179]), .Z(n3007));
Q_MX02 U1249 ( .S(n2642), .A0(n3007), .A1(xdata[147]), .Z(ofifoDataN[179]));
Q_AN02 U1250 ( .A0(n2641), .A1(xdata[180]), .Z(n3006));
Q_MX02 U1251 ( .S(n2642), .A0(n3006), .A1(xdata[148]), .Z(ofifoDataN[180]));
Q_AN02 U1252 ( .A0(n2641), .A1(xdata[181]), .Z(n3005));
Q_MX02 U1253 ( .S(n2642), .A0(n3005), .A1(xdata[149]), .Z(ofifoDataN[181]));
Q_AN02 U1254 ( .A0(n2641), .A1(xdata[182]), .Z(n3004));
Q_MX02 U1255 ( .S(n2642), .A0(n3004), .A1(xdata[150]), .Z(ofifoDataN[182]));
Q_AN02 U1256 ( .A0(n2641), .A1(xdata[183]), .Z(n3003));
Q_MX02 U1257 ( .S(n2642), .A0(n3003), .A1(xdata[151]), .Z(ofifoDataN[183]));
Q_AN02 U1258 ( .A0(n2641), .A1(xdata[184]), .Z(n3002));
Q_MX02 U1259 ( .S(n2642), .A0(n3002), .A1(xdata[152]), .Z(ofifoDataN[184]));
Q_AN02 U1260 ( .A0(n2641), .A1(xdata[185]), .Z(n3001));
Q_MX02 U1261 ( .S(n2642), .A0(n3001), .A1(xdata[153]), .Z(ofifoDataN[185]));
Q_AN02 U1262 ( .A0(n2641), .A1(xdata[186]), .Z(n3000));
Q_MX02 U1263 ( .S(n2642), .A0(n3000), .A1(xdata[154]), .Z(ofifoDataN[186]));
Q_AN02 U1264 ( .A0(n2641), .A1(xdata[187]), .Z(n2999));
Q_MX02 U1265 ( .S(n2642), .A0(n2999), .A1(xdata[155]), .Z(ofifoDataN[187]));
Q_AN02 U1266 ( .A0(n2641), .A1(xdata[188]), .Z(n2998));
Q_MX02 U1267 ( .S(n2642), .A0(n2998), .A1(xdata[156]), .Z(ofifoDataN[188]));
Q_AN02 U1268 ( .A0(n2641), .A1(xdata[189]), .Z(n2997));
Q_MX02 U1269 ( .S(n2642), .A0(n2997), .A1(xdata[157]), .Z(ofifoDataN[189]));
Q_AN02 U1270 ( .A0(n2641), .A1(xdata[190]), .Z(n2996));
Q_MX02 U1271 ( .S(n2642), .A0(n2996), .A1(xdata[158]), .Z(ofifoDataN[190]));
Q_AN02 U1272 ( .A0(n2641), .A1(xdata[191]), .Z(n2995));
Q_MX02 U1273 ( .S(n2642), .A0(n2995), .A1(xdata[159]), .Z(ofifoDataN[191]));
Q_AN02 U1274 ( .A0(n2641), .A1(xdata[192]), .Z(n2994));
Q_MX02 U1275 ( .S(n2642), .A0(n2994), .A1(xdata[160]), .Z(ofifoDataN[192]));
Q_AN02 U1276 ( .A0(n2641), .A1(xdata[193]), .Z(n2993));
Q_MX02 U1277 ( .S(n2642), .A0(n2993), .A1(xdata[161]), .Z(ofifoDataN[193]));
Q_AN02 U1278 ( .A0(n2641), .A1(xdata[194]), .Z(n2992));
Q_MX02 U1279 ( .S(n2642), .A0(n2992), .A1(xdata[162]), .Z(ofifoDataN[194]));
Q_AN02 U1280 ( .A0(n2641), .A1(xdata[195]), .Z(n2991));
Q_MX02 U1281 ( .S(n2642), .A0(n2991), .A1(xdata[163]), .Z(ofifoDataN[195]));
Q_AN02 U1282 ( .A0(n2641), .A1(xdata[196]), .Z(n2990));
Q_MX02 U1283 ( .S(n2642), .A0(n2990), .A1(xdata[164]), .Z(ofifoDataN[196]));
Q_AN02 U1284 ( .A0(n2641), .A1(xdata[197]), .Z(n2989));
Q_MX02 U1285 ( .S(n2642), .A0(n2989), .A1(xdata[165]), .Z(ofifoDataN[197]));
Q_AN02 U1286 ( .A0(n2641), .A1(xdata[198]), .Z(n2988));
Q_MX02 U1287 ( .S(n2642), .A0(n2988), .A1(xdata[166]), .Z(ofifoDataN[198]));
Q_AN02 U1288 ( .A0(n2641), .A1(xdata[199]), .Z(n2987));
Q_MX02 U1289 ( .S(n2642), .A0(n2987), .A1(xdata[167]), .Z(ofifoDataN[199]));
Q_AN02 U1290 ( .A0(n2641), .A1(xdata[200]), .Z(n2986));
Q_MX02 U1291 ( .S(n2642), .A0(n2986), .A1(xdata[168]), .Z(ofifoDataN[200]));
Q_AN02 U1292 ( .A0(n2641), .A1(xdata[201]), .Z(n2985));
Q_MX02 U1293 ( .S(n2642), .A0(n2985), .A1(xdata[169]), .Z(ofifoDataN[201]));
Q_AN02 U1294 ( .A0(n2641), .A1(xdata[202]), .Z(n2984));
Q_MX02 U1295 ( .S(n2642), .A0(n2984), .A1(xdata[170]), .Z(ofifoDataN[202]));
Q_AN02 U1296 ( .A0(n2641), .A1(xdata[203]), .Z(n2983));
Q_MX02 U1297 ( .S(n2642), .A0(n2983), .A1(xdata[171]), .Z(ofifoDataN[203]));
Q_AN02 U1298 ( .A0(n2641), .A1(xdata[204]), .Z(n2982));
Q_MX02 U1299 ( .S(n2642), .A0(n2982), .A1(xdata[172]), .Z(ofifoDataN[204]));
Q_AN02 U1300 ( .A0(n2641), .A1(xdata[205]), .Z(n2981));
Q_MX02 U1301 ( .S(n2642), .A0(n2981), .A1(xdata[173]), .Z(ofifoDataN[205]));
Q_AN02 U1302 ( .A0(n2641), .A1(xdata[206]), .Z(n2980));
Q_MX02 U1303 ( .S(n2642), .A0(n2980), .A1(xdata[174]), .Z(ofifoDataN[206]));
Q_AN02 U1304 ( .A0(n2641), .A1(xdata[207]), .Z(n2979));
Q_MX02 U1305 ( .S(n2642), .A0(n2979), .A1(xdata[175]), .Z(ofifoDataN[207]));
Q_AN02 U1306 ( .A0(n2641), .A1(xdata[208]), .Z(n2978));
Q_MX02 U1307 ( .S(n2642), .A0(n2978), .A1(xdata[176]), .Z(ofifoDataN[208]));
Q_AN02 U1308 ( .A0(n2641), .A1(xdata[209]), .Z(n2977));
Q_MX02 U1309 ( .S(n2642), .A0(n2977), .A1(xdata[177]), .Z(ofifoDataN[209]));
Q_AN02 U1310 ( .A0(n2641), .A1(xdata[210]), .Z(n2976));
Q_MX02 U1311 ( .S(n2642), .A0(n2976), .A1(xdata[178]), .Z(ofifoDataN[210]));
Q_AN02 U1312 ( .A0(n2641), .A1(xdata[211]), .Z(n2975));
Q_MX02 U1313 ( .S(n2642), .A0(n2975), .A1(xdata[179]), .Z(ofifoDataN[211]));
Q_AN02 U1314 ( .A0(n2641), .A1(xdata[212]), .Z(n2974));
Q_MX02 U1315 ( .S(n2642), .A0(n2974), .A1(xdata[180]), .Z(ofifoDataN[212]));
Q_AN02 U1316 ( .A0(n2641), .A1(xdata[213]), .Z(n2973));
Q_MX02 U1317 ( .S(n2642), .A0(n2973), .A1(xdata[181]), .Z(ofifoDataN[213]));
Q_AN02 U1318 ( .A0(n2641), .A1(xdata[214]), .Z(n2972));
Q_MX02 U1319 ( .S(n2642), .A0(n2972), .A1(xdata[182]), .Z(ofifoDataN[214]));
Q_AN02 U1320 ( .A0(n2641), .A1(xdata[215]), .Z(n2971));
Q_MX02 U1321 ( .S(n2642), .A0(n2971), .A1(xdata[183]), .Z(ofifoDataN[215]));
Q_AN02 U1322 ( .A0(n2641), .A1(xdata[216]), .Z(n2970));
Q_MX02 U1323 ( .S(n2642), .A0(n2970), .A1(xdata[184]), .Z(ofifoDataN[216]));
Q_AN02 U1324 ( .A0(n2641), .A1(xdata[217]), .Z(n2969));
Q_MX02 U1325 ( .S(n2642), .A0(n2969), .A1(xdata[185]), .Z(ofifoDataN[217]));
Q_AN02 U1326 ( .A0(n2641), .A1(xdata[218]), .Z(n2968));
Q_MX02 U1327 ( .S(n2642), .A0(n2968), .A1(xdata[186]), .Z(ofifoDataN[218]));
Q_AN02 U1328 ( .A0(n2641), .A1(xdata[219]), .Z(n2967));
Q_MX02 U1329 ( .S(n2642), .A0(n2967), .A1(xdata[187]), .Z(ofifoDataN[219]));
Q_AN02 U1330 ( .A0(n2641), .A1(xdata[220]), .Z(n2966));
Q_MX02 U1331 ( .S(n2642), .A0(n2966), .A1(xdata[188]), .Z(ofifoDataN[220]));
Q_AN02 U1332 ( .A0(n2641), .A1(xdata[221]), .Z(n2965));
Q_MX02 U1333 ( .S(n2642), .A0(n2965), .A1(xdata[189]), .Z(ofifoDataN[221]));
Q_AN02 U1334 ( .A0(n2641), .A1(xdata[222]), .Z(n2964));
Q_MX02 U1335 ( .S(n2642), .A0(n2964), .A1(xdata[190]), .Z(ofifoDataN[222]));
Q_AN02 U1336 ( .A0(n2641), .A1(xdata[223]), .Z(n2963));
Q_MX02 U1337 ( .S(n2642), .A0(n2963), .A1(xdata[191]), .Z(ofifoDataN[223]));
Q_AN02 U1338 ( .A0(n2641), .A1(xdata[224]), .Z(n2962));
Q_MX02 U1339 ( .S(n2642), .A0(n2962), .A1(xdata[192]), .Z(ofifoDataN[224]));
Q_AN02 U1340 ( .A0(n2641), .A1(xdata[225]), .Z(n2961));
Q_MX02 U1341 ( .S(n2642), .A0(n2961), .A1(xdata[193]), .Z(ofifoDataN[225]));
Q_AN02 U1342 ( .A0(n2641), .A1(xdata[226]), .Z(n2960));
Q_MX02 U1343 ( .S(n2642), .A0(n2960), .A1(xdata[194]), .Z(ofifoDataN[226]));
Q_AN02 U1344 ( .A0(n2641), .A1(xdata[227]), .Z(n2959));
Q_MX02 U1345 ( .S(n2642), .A0(n2959), .A1(xdata[195]), .Z(ofifoDataN[227]));
Q_AN02 U1346 ( .A0(n2641), .A1(xdata[228]), .Z(n2958));
Q_MX02 U1347 ( .S(n2642), .A0(n2958), .A1(xdata[196]), .Z(ofifoDataN[228]));
Q_AN02 U1348 ( .A0(n2641), .A1(xdata[229]), .Z(n2957));
Q_MX02 U1349 ( .S(n2642), .A0(n2957), .A1(xdata[197]), .Z(ofifoDataN[229]));
Q_AN02 U1350 ( .A0(n2641), .A1(xdata[230]), .Z(n2956));
Q_MX02 U1351 ( .S(n2642), .A0(n2956), .A1(xdata[198]), .Z(ofifoDataN[230]));
Q_AN02 U1352 ( .A0(n2641), .A1(xdata[231]), .Z(n2955));
Q_MX02 U1353 ( .S(n2642), .A0(n2955), .A1(xdata[199]), .Z(ofifoDataN[231]));
Q_AN02 U1354 ( .A0(n2641), .A1(xdata[232]), .Z(n2954));
Q_MX02 U1355 ( .S(n2642), .A0(n2954), .A1(xdata[200]), .Z(ofifoDataN[232]));
Q_AN02 U1356 ( .A0(n2641), .A1(xdata[233]), .Z(n2953));
Q_MX02 U1357 ( .S(n2642), .A0(n2953), .A1(xdata[201]), .Z(ofifoDataN[233]));
Q_AN02 U1358 ( .A0(n2641), .A1(xdata[234]), .Z(n2952));
Q_MX02 U1359 ( .S(n2642), .A0(n2952), .A1(xdata[202]), .Z(ofifoDataN[234]));
Q_AN02 U1360 ( .A0(n2641), .A1(xdata[235]), .Z(n2951));
Q_MX02 U1361 ( .S(n2642), .A0(n2951), .A1(xdata[203]), .Z(ofifoDataN[235]));
Q_AN02 U1362 ( .A0(n2641), .A1(xdata[236]), .Z(n2950));
Q_MX02 U1363 ( .S(n2642), .A0(n2950), .A1(xdata[204]), .Z(ofifoDataN[236]));
Q_AN02 U1364 ( .A0(n2641), .A1(xdata[237]), .Z(n2949));
Q_MX02 U1365 ( .S(n2642), .A0(n2949), .A1(xdata[205]), .Z(ofifoDataN[237]));
Q_AN02 U1366 ( .A0(n2641), .A1(xdata[238]), .Z(n2948));
Q_MX02 U1367 ( .S(n2642), .A0(n2948), .A1(xdata[206]), .Z(ofifoDataN[238]));
Q_AN02 U1368 ( .A0(n2641), .A1(xdata[239]), .Z(n2947));
Q_MX02 U1369 ( .S(n2642), .A0(n2947), .A1(xdata[207]), .Z(ofifoDataN[239]));
Q_AN02 U1370 ( .A0(n2641), .A1(xdata[240]), .Z(n2946));
Q_MX02 U1371 ( .S(n2642), .A0(n2946), .A1(xdata[208]), .Z(ofifoDataN[240]));
Q_AN02 U1372 ( .A0(n2641), .A1(xdata[241]), .Z(n2945));
Q_MX02 U1373 ( .S(n2642), .A0(n2945), .A1(xdata[209]), .Z(ofifoDataN[241]));
Q_AN02 U1374 ( .A0(n2641), .A1(xdata[242]), .Z(n2944));
Q_MX02 U1375 ( .S(n2642), .A0(n2944), .A1(xdata[210]), .Z(ofifoDataN[242]));
Q_AN02 U1376 ( .A0(n2641), .A1(xdata[243]), .Z(n2943));
Q_MX02 U1377 ( .S(n2642), .A0(n2943), .A1(xdata[211]), .Z(ofifoDataN[243]));
Q_AN02 U1378 ( .A0(n2641), .A1(xdata[244]), .Z(n2942));
Q_MX02 U1379 ( .S(n2642), .A0(n2942), .A1(xdata[212]), .Z(ofifoDataN[244]));
Q_AN02 U1380 ( .A0(n2641), .A1(xdata[245]), .Z(n2941));
Q_MX02 U1381 ( .S(n2642), .A0(n2941), .A1(xdata[213]), .Z(ofifoDataN[245]));
Q_AN02 U1382 ( .A0(n2641), .A1(xdata[246]), .Z(n2940));
Q_MX02 U1383 ( .S(n2642), .A0(n2940), .A1(xdata[214]), .Z(ofifoDataN[246]));
Q_AN02 U1384 ( .A0(n2641), .A1(xdata[247]), .Z(n2939));
Q_MX02 U1385 ( .S(n2642), .A0(n2939), .A1(xdata[215]), .Z(ofifoDataN[247]));
Q_AN02 U1386 ( .A0(n2641), .A1(xdata[248]), .Z(n2938));
Q_MX02 U1387 ( .S(n2642), .A0(n2938), .A1(xdata[216]), .Z(ofifoDataN[248]));
Q_AN02 U1388 ( .A0(n2641), .A1(xdata[249]), .Z(n2937));
Q_MX02 U1389 ( .S(n2642), .A0(n2937), .A1(xdata[217]), .Z(ofifoDataN[249]));
Q_AN02 U1390 ( .A0(n2641), .A1(xdata[250]), .Z(n2936));
Q_MX02 U1391 ( .S(n2642), .A0(n2936), .A1(xdata[218]), .Z(ofifoDataN[250]));
Q_AN02 U1392 ( .A0(n2641), .A1(xdata[251]), .Z(n2935));
Q_MX02 U1393 ( .S(n2642), .A0(n2935), .A1(xdata[219]), .Z(ofifoDataN[251]));
Q_AN02 U1394 ( .A0(n2641), .A1(xdata[252]), .Z(n2934));
Q_MX02 U1395 ( .S(n2642), .A0(n2934), .A1(xdata[220]), .Z(ofifoDataN[252]));
Q_AN02 U1396 ( .A0(n2641), .A1(xdata[253]), .Z(n2933));
Q_MX02 U1397 ( .S(n2642), .A0(n2933), .A1(xdata[221]), .Z(ofifoDataN[253]));
Q_AN02 U1398 ( .A0(n2641), .A1(xdata[254]), .Z(n2932));
Q_MX02 U1399 ( .S(n2642), .A0(n2932), .A1(xdata[222]), .Z(ofifoDataN[254]));
Q_AN02 U1400 ( .A0(n2641), .A1(xdata[255]), .Z(n2931));
Q_MX02 U1401 ( .S(n2642), .A0(n2931), .A1(xdata[223]), .Z(ofifoDataN[255]));
Q_AN02 U1402 ( .A0(n2641), .A1(xdata[256]), .Z(n2930));
Q_MX02 U1403 ( .S(n2642), .A0(n2930), .A1(xdata[224]), .Z(ofifoDataN[256]));
Q_AN02 U1404 ( .A0(n2641), .A1(xdata[257]), .Z(n2929));
Q_MX02 U1405 ( .S(n2642), .A0(n2929), .A1(xdata[225]), .Z(ofifoDataN[257]));
Q_AN02 U1406 ( .A0(n2641), .A1(xdata[258]), .Z(n2928));
Q_MX02 U1407 ( .S(n2642), .A0(n2928), .A1(xdata[226]), .Z(ofifoDataN[258]));
Q_AN02 U1408 ( .A0(n2641), .A1(xdata[259]), .Z(n2927));
Q_MX02 U1409 ( .S(n2642), .A0(n2927), .A1(xdata[227]), .Z(ofifoDataN[259]));
Q_AN02 U1410 ( .A0(n2641), .A1(xdata[260]), .Z(n2926));
Q_MX02 U1411 ( .S(n2642), .A0(n2926), .A1(xdata[228]), .Z(ofifoDataN[260]));
Q_AN02 U1412 ( .A0(n2641), .A1(xdata[261]), .Z(n2925));
Q_MX02 U1413 ( .S(n2642), .A0(n2925), .A1(xdata[229]), .Z(ofifoDataN[261]));
Q_AN02 U1414 ( .A0(n2641), .A1(xdata[262]), .Z(n2924));
Q_MX02 U1415 ( .S(n2642), .A0(n2924), .A1(xdata[230]), .Z(ofifoDataN[262]));
Q_AN02 U1416 ( .A0(n2641), .A1(xdata[263]), .Z(n2923));
Q_MX02 U1417 ( .S(n2642), .A0(n2923), .A1(xdata[231]), .Z(ofifoDataN[263]));
Q_AN02 U1418 ( .A0(n2641), .A1(xdata[264]), .Z(n2922));
Q_MX02 U1419 ( .S(n2642), .A0(n2922), .A1(xdata[232]), .Z(ofifoDataN[264]));
Q_AN02 U1420 ( .A0(n2641), .A1(xdata[265]), .Z(n2921));
Q_MX02 U1421 ( .S(n2642), .A0(n2921), .A1(xdata[233]), .Z(ofifoDataN[265]));
Q_AN02 U1422 ( .A0(n2641), .A1(xdata[266]), .Z(n2920));
Q_MX02 U1423 ( .S(n2642), .A0(n2920), .A1(xdata[234]), .Z(ofifoDataN[266]));
Q_AN02 U1424 ( .A0(n2641), .A1(xdata[267]), .Z(n2919));
Q_MX02 U1425 ( .S(n2642), .A0(n2919), .A1(xdata[235]), .Z(ofifoDataN[267]));
Q_AN02 U1426 ( .A0(n2641), .A1(xdata[268]), .Z(n2918));
Q_MX02 U1427 ( .S(n2642), .A0(n2918), .A1(xdata[236]), .Z(ofifoDataN[268]));
Q_AN02 U1428 ( .A0(n2641), .A1(xdata[269]), .Z(n2917));
Q_MX02 U1429 ( .S(n2642), .A0(n2917), .A1(xdata[237]), .Z(ofifoDataN[269]));
Q_AN02 U1430 ( .A0(n2641), .A1(xdata[270]), .Z(n2916));
Q_MX02 U1431 ( .S(n2642), .A0(n2916), .A1(xdata[238]), .Z(ofifoDataN[270]));
Q_AN02 U1432 ( .A0(n2641), .A1(xdata[271]), .Z(n2915));
Q_MX02 U1433 ( .S(n2642), .A0(n2915), .A1(xdata[239]), .Z(ofifoDataN[271]));
Q_AN02 U1434 ( .A0(n2641), .A1(xdata[272]), .Z(n2914));
Q_MX02 U1435 ( .S(n2642), .A0(n2914), .A1(xdata[240]), .Z(ofifoDataN[272]));
Q_AN02 U1436 ( .A0(n2641), .A1(xdata[273]), .Z(n2913));
Q_MX02 U1437 ( .S(n2642), .A0(n2913), .A1(xdata[241]), .Z(ofifoDataN[273]));
Q_AN02 U1438 ( .A0(n2641), .A1(xdata[274]), .Z(n2912));
Q_MX02 U1439 ( .S(n2642), .A0(n2912), .A1(xdata[242]), .Z(ofifoDataN[274]));
Q_AN02 U1440 ( .A0(n2641), .A1(xdata[275]), .Z(n2911));
Q_MX02 U1441 ( .S(n2642), .A0(n2911), .A1(xdata[243]), .Z(ofifoDataN[275]));
Q_AN02 U1442 ( .A0(n2641), .A1(xdata[276]), .Z(n2910));
Q_MX02 U1443 ( .S(n2642), .A0(n2910), .A1(xdata[244]), .Z(ofifoDataN[276]));
Q_AN02 U1444 ( .A0(n2641), .A1(xdata[277]), .Z(n2909));
Q_MX02 U1445 ( .S(n2642), .A0(n2909), .A1(xdata[245]), .Z(ofifoDataN[277]));
Q_AN02 U1446 ( .A0(n2641), .A1(xdata[278]), .Z(n2908));
Q_MX02 U1447 ( .S(n2642), .A0(n2908), .A1(xdata[246]), .Z(ofifoDataN[278]));
Q_AN02 U1448 ( .A0(n2641), .A1(xdata[279]), .Z(n2907));
Q_MX02 U1449 ( .S(n2642), .A0(n2907), .A1(xdata[247]), .Z(ofifoDataN[279]));
Q_AN02 U1450 ( .A0(n2641), .A1(xdata[280]), .Z(n2906));
Q_MX02 U1451 ( .S(n2642), .A0(n2906), .A1(xdata[248]), .Z(ofifoDataN[280]));
Q_AN02 U1452 ( .A0(n2641), .A1(xdata[281]), .Z(n2905));
Q_MX02 U1453 ( .S(n2642), .A0(n2905), .A1(xdata[249]), .Z(ofifoDataN[281]));
Q_AN02 U1454 ( .A0(n2641), .A1(xdata[282]), .Z(n2904));
Q_MX02 U1455 ( .S(n2642), .A0(n2904), .A1(xdata[250]), .Z(ofifoDataN[282]));
Q_AN02 U1456 ( .A0(n2641), .A1(xdata[283]), .Z(n2903));
Q_MX02 U1457 ( .S(n2642), .A0(n2903), .A1(xdata[251]), .Z(ofifoDataN[283]));
Q_AN02 U1458 ( .A0(n2641), .A1(xdata[284]), .Z(n2902));
Q_MX02 U1459 ( .S(n2642), .A0(n2902), .A1(xdata[252]), .Z(ofifoDataN[284]));
Q_AN02 U1460 ( .A0(n2641), .A1(xdata[285]), .Z(n2901));
Q_MX02 U1461 ( .S(n2642), .A0(n2901), .A1(xdata[253]), .Z(ofifoDataN[285]));
Q_AN02 U1462 ( .A0(n2641), .A1(xdata[286]), .Z(n2900));
Q_MX02 U1463 ( .S(n2642), .A0(n2900), .A1(xdata[254]), .Z(ofifoDataN[286]));
Q_AN02 U1464 ( .A0(n2641), .A1(xdata[287]), .Z(n2899));
Q_MX02 U1465 ( .S(n2642), .A0(n2899), .A1(xdata[255]), .Z(ofifoDataN[287]));
Q_AN02 U1466 ( .A0(n2641), .A1(xdata[288]), .Z(n2898));
Q_MX02 U1467 ( .S(n2642), .A0(n2898), .A1(xdata[256]), .Z(ofifoDataN[288]));
Q_AN02 U1468 ( .A0(n2641), .A1(xdata[289]), .Z(n2897));
Q_MX02 U1469 ( .S(n2642), .A0(n2897), .A1(xdata[257]), .Z(ofifoDataN[289]));
Q_AN02 U1470 ( .A0(n2641), .A1(xdata[290]), .Z(n2896));
Q_MX02 U1471 ( .S(n2642), .A0(n2896), .A1(xdata[258]), .Z(ofifoDataN[290]));
Q_AN02 U1472 ( .A0(n2641), .A1(xdata[291]), .Z(n2895));
Q_MX02 U1473 ( .S(n2642), .A0(n2895), .A1(xdata[259]), .Z(ofifoDataN[291]));
Q_AN02 U1474 ( .A0(n2641), .A1(xdata[292]), .Z(n2894));
Q_MX02 U1475 ( .S(n2642), .A0(n2894), .A1(xdata[260]), .Z(ofifoDataN[292]));
Q_AN02 U1476 ( .A0(n2641), .A1(xdata[293]), .Z(n2893));
Q_MX02 U1477 ( .S(n2642), .A0(n2893), .A1(xdata[261]), .Z(ofifoDataN[293]));
Q_AN02 U1478 ( .A0(n2641), .A1(xdata[294]), .Z(n2892));
Q_MX02 U1479 ( .S(n2642), .A0(n2892), .A1(xdata[262]), .Z(ofifoDataN[294]));
Q_AN02 U1480 ( .A0(n2641), .A1(xdata[295]), .Z(n2891));
Q_MX02 U1481 ( .S(n2642), .A0(n2891), .A1(xdata[263]), .Z(ofifoDataN[295]));
Q_AN02 U1482 ( .A0(n2641), .A1(xdata[296]), .Z(n2890));
Q_MX02 U1483 ( .S(n2642), .A0(n2890), .A1(xdata[264]), .Z(ofifoDataN[296]));
Q_AN02 U1484 ( .A0(n2641), .A1(xdata[297]), .Z(n2889));
Q_MX02 U1485 ( .S(n2642), .A0(n2889), .A1(xdata[265]), .Z(ofifoDataN[297]));
Q_AN02 U1486 ( .A0(n2641), .A1(xdata[298]), .Z(n2888));
Q_MX02 U1487 ( .S(n2642), .A0(n2888), .A1(xdata[266]), .Z(ofifoDataN[298]));
Q_AN02 U1488 ( .A0(n2641), .A1(xdata[299]), .Z(n2887));
Q_MX02 U1489 ( .S(n2642), .A0(n2887), .A1(xdata[267]), .Z(ofifoDataN[299]));
Q_AN02 U1490 ( .A0(n2641), .A1(xdata[300]), .Z(n2886));
Q_MX02 U1491 ( .S(n2642), .A0(n2886), .A1(xdata[268]), .Z(ofifoDataN[300]));
Q_AN02 U1492 ( .A0(n2641), .A1(xdata[301]), .Z(n2885));
Q_MX02 U1493 ( .S(n2642), .A0(n2885), .A1(xdata[269]), .Z(ofifoDataN[301]));
Q_AN02 U1494 ( .A0(n2641), .A1(xdata[302]), .Z(n2884));
Q_MX02 U1495 ( .S(n2642), .A0(n2884), .A1(xdata[270]), .Z(ofifoDataN[302]));
Q_AN02 U1496 ( .A0(n2641), .A1(xdata[303]), .Z(n2883));
Q_MX02 U1497 ( .S(n2642), .A0(n2883), .A1(xdata[271]), .Z(ofifoDataN[303]));
Q_AN02 U1498 ( .A0(n2641), .A1(xdata[304]), .Z(n2882));
Q_MX02 U1499 ( .S(n2642), .A0(n2882), .A1(xdata[272]), .Z(ofifoDataN[304]));
Q_AN02 U1500 ( .A0(n2641), .A1(xdata[305]), .Z(n2881));
Q_MX02 U1501 ( .S(n2642), .A0(n2881), .A1(xdata[273]), .Z(ofifoDataN[305]));
Q_AN02 U1502 ( .A0(n2641), .A1(xdata[306]), .Z(n2880));
Q_MX02 U1503 ( .S(n2642), .A0(n2880), .A1(xdata[274]), .Z(ofifoDataN[306]));
Q_AN02 U1504 ( .A0(n2641), .A1(xdata[307]), .Z(n2879));
Q_MX02 U1505 ( .S(n2642), .A0(n2879), .A1(xdata[275]), .Z(ofifoDataN[307]));
Q_AN02 U1506 ( .A0(n2641), .A1(xdata[308]), .Z(n2878));
Q_MX02 U1507 ( .S(n2642), .A0(n2878), .A1(xdata[276]), .Z(ofifoDataN[308]));
Q_AN02 U1508 ( .A0(n2641), .A1(xdata[309]), .Z(n2877));
Q_MX02 U1509 ( .S(n2642), .A0(n2877), .A1(xdata[277]), .Z(ofifoDataN[309]));
Q_AN02 U1510 ( .A0(n2641), .A1(xdata[310]), .Z(n2876));
Q_MX02 U1511 ( .S(n2642), .A0(n2876), .A1(xdata[278]), .Z(ofifoDataN[310]));
Q_AN02 U1512 ( .A0(n2641), .A1(xdata[311]), .Z(n2875));
Q_MX02 U1513 ( .S(n2642), .A0(n2875), .A1(xdata[279]), .Z(ofifoDataN[311]));
Q_AN02 U1514 ( .A0(n2641), .A1(xdata[312]), .Z(n2874));
Q_MX02 U1515 ( .S(n2642), .A0(n2874), .A1(xdata[280]), .Z(ofifoDataN[312]));
Q_AN02 U1516 ( .A0(n2641), .A1(xdata[313]), .Z(n2873));
Q_MX02 U1517 ( .S(n2642), .A0(n2873), .A1(xdata[281]), .Z(ofifoDataN[313]));
Q_AN02 U1518 ( .A0(n2641), .A1(xdata[314]), .Z(n2872));
Q_MX02 U1519 ( .S(n2642), .A0(n2872), .A1(xdata[282]), .Z(ofifoDataN[314]));
Q_AN02 U1520 ( .A0(n2641), .A1(xdata[315]), .Z(n2871));
Q_MX02 U1521 ( .S(n2642), .A0(n2871), .A1(xdata[283]), .Z(ofifoDataN[315]));
Q_AN02 U1522 ( .A0(n2641), .A1(xdata[316]), .Z(n2870));
Q_MX02 U1523 ( .S(n2642), .A0(n2870), .A1(xdata[284]), .Z(ofifoDataN[316]));
Q_AN02 U1524 ( .A0(n2641), .A1(xdata[317]), .Z(n2869));
Q_MX02 U1525 ( .S(n2642), .A0(n2869), .A1(xdata[285]), .Z(ofifoDataN[317]));
Q_AN02 U1526 ( .A0(n2641), .A1(xdata[318]), .Z(n2868));
Q_MX02 U1527 ( .S(n2642), .A0(n2868), .A1(xdata[286]), .Z(ofifoDataN[318]));
Q_AN02 U1528 ( .A0(n2641), .A1(xdata[319]), .Z(n2867));
Q_MX02 U1529 ( .S(n2642), .A0(n2867), .A1(xdata[287]), .Z(ofifoDataN[319]));
Q_AN02 U1530 ( .A0(n2641), .A1(xdata[320]), .Z(n2866));
Q_MX02 U1531 ( .S(n2642), .A0(n2866), .A1(xdata[288]), .Z(ofifoDataN[320]));
Q_AN02 U1532 ( .A0(n2641), .A1(xdata[321]), .Z(n2865));
Q_MX02 U1533 ( .S(n2642), .A0(n2865), .A1(xdata[289]), .Z(ofifoDataN[321]));
Q_AN02 U1534 ( .A0(n2641), .A1(xdata[322]), .Z(n2864));
Q_MX02 U1535 ( .S(n2642), .A0(n2864), .A1(xdata[290]), .Z(ofifoDataN[322]));
Q_AN02 U1536 ( .A0(n2641), .A1(xdata[323]), .Z(n2863));
Q_MX02 U1537 ( .S(n2642), .A0(n2863), .A1(xdata[291]), .Z(ofifoDataN[323]));
Q_AN02 U1538 ( .A0(n2641), .A1(xdata[324]), .Z(n2862));
Q_MX02 U1539 ( .S(n2642), .A0(n2862), .A1(xdata[292]), .Z(ofifoDataN[324]));
Q_AN02 U1540 ( .A0(n2641), .A1(xdata[325]), .Z(n2861));
Q_MX02 U1541 ( .S(n2642), .A0(n2861), .A1(xdata[293]), .Z(ofifoDataN[325]));
Q_AN02 U1542 ( .A0(n2641), .A1(xdata[326]), .Z(n2860));
Q_MX02 U1543 ( .S(n2642), .A0(n2860), .A1(xdata[294]), .Z(ofifoDataN[326]));
Q_AN02 U1544 ( .A0(n2641), .A1(xdata[327]), .Z(n2859));
Q_MX02 U1545 ( .S(n2642), .A0(n2859), .A1(xdata[295]), .Z(ofifoDataN[327]));
Q_AN02 U1546 ( .A0(n2641), .A1(xdata[328]), .Z(n2858));
Q_MX02 U1547 ( .S(n2642), .A0(n2858), .A1(xdata[296]), .Z(ofifoDataN[328]));
Q_AN02 U1548 ( .A0(n2641), .A1(xdata[329]), .Z(n2857));
Q_MX02 U1549 ( .S(n2642), .A0(n2857), .A1(xdata[297]), .Z(ofifoDataN[329]));
Q_AN02 U1550 ( .A0(n2641), .A1(xdata[330]), .Z(n2856));
Q_MX02 U1551 ( .S(n2642), .A0(n2856), .A1(xdata[298]), .Z(ofifoDataN[330]));
Q_AN02 U1552 ( .A0(n2641), .A1(xdata[331]), .Z(n2855));
Q_MX02 U1553 ( .S(n2642), .A0(n2855), .A1(xdata[299]), .Z(ofifoDataN[331]));
Q_AN02 U1554 ( .A0(n2641), .A1(xdata[332]), .Z(n2854));
Q_MX02 U1555 ( .S(n2642), .A0(n2854), .A1(xdata[300]), .Z(ofifoDataN[332]));
Q_AN02 U1556 ( .A0(n2641), .A1(xdata[333]), .Z(n2853));
Q_MX02 U1557 ( .S(n2642), .A0(n2853), .A1(xdata[301]), .Z(ofifoDataN[333]));
Q_AN02 U1558 ( .A0(n2641), .A1(xdata[334]), .Z(n2852));
Q_MX02 U1559 ( .S(n2642), .A0(n2852), .A1(xdata[302]), .Z(ofifoDataN[334]));
Q_AN02 U1560 ( .A0(n2641), .A1(xdata[335]), .Z(n2851));
Q_MX02 U1561 ( .S(n2642), .A0(n2851), .A1(xdata[303]), .Z(ofifoDataN[335]));
Q_AN02 U1562 ( .A0(n2641), .A1(xdata[336]), .Z(n2850));
Q_MX02 U1563 ( .S(n2642), .A0(n2850), .A1(xdata[304]), .Z(ofifoDataN[336]));
Q_AN02 U1564 ( .A0(n2641), .A1(xdata[337]), .Z(n2849));
Q_MX02 U1565 ( .S(n2642), .A0(n2849), .A1(xdata[305]), .Z(ofifoDataN[337]));
Q_AN02 U1566 ( .A0(n2641), .A1(xdata[338]), .Z(n2848));
Q_MX02 U1567 ( .S(n2642), .A0(n2848), .A1(xdata[306]), .Z(ofifoDataN[338]));
Q_AN02 U1568 ( .A0(n2641), .A1(xdata[339]), .Z(n2847));
Q_MX02 U1569 ( .S(n2642), .A0(n2847), .A1(xdata[307]), .Z(ofifoDataN[339]));
Q_AN02 U1570 ( .A0(n2641), .A1(xdata[340]), .Z(n2846));
Q_MX02 U1571 ( .S(n2642), .A0(n2846), .A1(xdata[308]), .Z(ofifoDataN[340]));
Q_AN02 U1572 ( .A0(n2641), .A1(xdata[341]), .Z(n2845));
Q_MX02 U1573 ( .S(n2642), .A0(n2845), .A1(xdata[309]), .Z(ofifoDataN[341]));
Q_AN02 U1574 ( .A0(n2641), .A1(xdata[342]), .Z(n2844));
Q_MX02 U1575 ( .S(n2642), .A0(n2844), .A1(xdata[310]), .Z(ofifoDataN[342]));
Q_AN02 U1576 ( .A0(n2641), .A1(xdata[343]), .Z(n2843));
Q_MX02 U1577 ( .S(n2642), .A0(n2843), .A1(xdata[311]), .Z(ofifoDataN[343]));
Q_AN02 U1578 ( .A0(n2641), .A1(xdata[344]), .Z(n2842));
Q_MX02 U1579 ( .S(n2642), .A0(n2842), .A1(xdata[312]), .Z(ofifoDataN[344]));
Q_AN02 U1580 ( .A0(n2641), .A1(xdata[345]), .Z(n2841));
Q_MX02 U1581 ( .S(n2642), .A0(n2841), .A1(xdata[313]), .Z(ofifoDataN[345]));
Q_AN02 U1582 ( .A0(n2641), .A1(xdata[346]), .Z(n2840));
Q_MX02 U1583 ( .S(n2642), .A0(n2840), .A1(xdata[314]), .Z(ofifoDataN[346]));
Q_AN02 U1584 ( .A0(n2641), .A1(xdata[347]), .Z(n2839));
Q_MX02 U1585 ( .S(n2642), .A0(n2839), .A1(xdata[315]), .Z(ofifoDataN[347]));
Q_AN02 U1586 ( .A0(n2641), .A1(xdata[348]), .Z(n2838));
Q_MX02 U1587 ( .S(n2642), .A0(n2838), .A1(xdata[316]), .Z(ofifoDataN[348]));
Q_AN02 U1588 ( .A0(n2641), .A1(xdata[349]), .Z(n2837));
Q_MX02 U1589 ( .S(n2642), .A0(n2837), .A1(xdata[317]), .Z(ofifoDataN[349]));
Q_AN02 U1590 ( .A0(n2641), .A1(xdata[350]), .Z(n2836));
Q_MX02 U1591 ( .S(n2642), .A0(n2836), .A1(xdata[318]), .Z(ofifoDataN[350]));
Q_AN02 U1592 ( .A0(n2641), .A1(xdata[351]), .Z(n2835));
Q_MX02 U1593 ( .S(n2642), .A0(n2835), .A1(xdata[319]), .Z(ofifoDataN[351]));
Q_AN02 U1594 ( .A0(n2641), .A1(xdata[352]), .Z(n2834));
Q_MX02 U1595 ( .S(n2642), .A0(n2834), .A1(xdata[320]), .Z(ofifoDataN[352]));
Q_AN02 U1596 ( .A0(n2641), .A1(xdata[353]), .Z(n2833));
Q_MX02 U1597 ( .S(n2642), .A0(n2833), .A1(xdata[321]), .Z(ofifoDataN[353]));
Q_AN02 U1598 ( .A0(n2641), .A1(xdata[354]), .Z(n2832));
Q_MX02 U1599 ( .S(n2642), .A0(n2832), .A1(xdata[322]), .Z(ofifoDataN[354]));
Q_AN02 U1600 ( .A0(n2641), .A1(xdata[355]), .Z(n2831));
Q_MX02 U1601 ( .S(n2642), .A0(n2831), .A1(xdata[323]), .Z(ofifoDataN[355]));
Q_AN02 U1602 ( .A0(n2641), .A1(xdata[356]), .Z(n2830));
Q_MX02 U1603 ( .S(n2642), .A0(n2830), .A1(xdata[324]), .Z(ofifoDataN[356]));
Q_AN02 U1604 ( .A0(n2641), .A1(xdata[357]), .Z(n2829));
Q_MX02 U1605 ( .S(n2642), .A0(n2829), .A1(xdata[325]), .Z(ofifoDataN[357]));
Q_AN02 U1606 ( .A0(n2641), .A1(xdata[358]), .Z(n2828));
Q_MX02 U1607 ( .S(n2642), .A0(n2828), .A1(xdata[326]), .Z(ofifoDataN[358]));
Q_AN02 U1608 ( .A0(n2641), .A1(xdata[359]), .Z(n2827));
Q_MX02 U1609 ( .S(n2642), .A0(n2827), .A1(xdata[327]), .Z(ofifoDataN[359]));
Q_AN02 U1610 ( .A0(n2641), .A1(xdata[360]), .Z(n2826));
Q_MX02 U1611 ( .S(n2642), .A0(n2826), .A1(xdata[328]), .Z(ofifoDataN[360]));
Q_AN02 U1612 ( .A0(n2641), .A1(xdata[361]), .Z(n2825));
Q_MX02 U1613 ( .S(n2642), .A0(n2825), .A1(xdata[329]), .Z(ofifoDataN[361]));
Q_AN02 U1614 ( .A0(n2641), .A1(xdata[362]), .Z(n2824));
Q_MX02 U1615 ( .S(n2642), .A0(n2824), .A1(xdata[330]), .Z(ofifoDataN[362]));
Q_AN02 U1616 ( .A0(n2641), .A1(xdata[363]), .Z(n2823));
Q_MX02 U1617 ( .S(n2642), .A0(n2823), .A1(xdata[331]), .Z(ofifoDataN[363]));
Q_AN02 U1618 ( .A0(n2641), .A1(xdata[364]), .Z(n2822));
Q_MX02 U1619 ( .S(n2642), .A0(n2822), .A1(xdata[332]), .Z(ofifoDataN[364]));
Q_AN02 U1620 ( .A0(n2641), .A1(xdata[365]), .Z(n2821));
Q_MX02 U1621 ( .S(n2642), .A0(n2821), .A1(xdata[333]), .Z(ofifoDataN[365]));
Q_AN02 U1622 ( .A0(n2641), .A1(xdata[366]), .Z(n2820));
Q_MX02 U1623 ( .S(n2642), .A0(n2820), .A1(xdata[334]), .Z(ofifoDataN[366]));
Q_AN02 U1624 ( .A0(n2641), .A1(xdata[367]), .Z(n2819));
Q_MX02 U1625 ( .S(n2642), .A0(n2819), .A1(xdata[335]), .Z(ofifoDataN[367]));
Q_AN02 U1626 ( .A0(n2641), .A1(xdata[368]), .Z(n2818));
Q_MX02 U1627 ( .S(n2642), .A0(n2818), .A1(xdata[336]), .Z(ofifoDataN[368]));
Q_AN02 U1628 ( .A0(n2641), .A1(xdata[369]), .Z(n2817));
Q_MX02 U1629 ( .S(n2642), .A0(n2817), .A1(xdata[337]), .Z(ofifoDataN[369]));
Q_AN02 U1630 ( .A0(n2641), .A1(xdata[370]), .Z(n2816));
Q_MX02 U1631 ( .S(n2642), .A0(n2816), .A1(xdata[338]), .Z(ofifoDataN[370]));
Q_AN02 U1632 ( .A0(n2641), .A1(xdata[371]), .Z(n2815));
Q_MX02 U1633 ( .S(n2642), .A0(n2815), .A1(xdata[339]), .Z(ofifoDataN[371]));
Q_AN02 U1634 ( .A0(n2641), .A1(xdata[372]), .Z(n2814));
Q_MX02 U1635 ( .S(n2642), .A0(n2814), .A1(xdata[340]), .Z(ofifoDataN[372]));
Q_AN02 U1636 ( .A0(n2641), .A1(xdata[373]), .Z(n2813));
Q_MX02 U1637 ( .S(n2642), .A0(n2813), .A1(xdata[341]), .Z(ofifoDataN[373]));
Q_AN02 U1638 ( .A0(n2641), .A1(xdata[374]), .Z(n2812));
Q_MX02 U1639 ( .S(n2642), .A0(n2812), .A1(xdata[342]), .Z(ofifoDataN[374]));
Q_AN02 U1640 ( .A0(n2641), .A1(xdata[375]), .Z(n2811));
Q_MX02 U1641 ( .S(n2642), .A0(n2811), .A1(xdata[343]), .Z(ofifoDataN[375]));
Q_AN02 U1642 ( .A0(n2641), .A1(xdata[376]), .Z(n2810));
Q_MX02 U1643 ( .S(n2642), .A0(n2810), .A1(xdata[344]), .Z(ofifoDataN[376]));
Q_AN02 U1644 ( .A0(n2641), .A1(xdata[377]), .Z(n2809));
Q_MX02 U1645 ( .S(n2642), .A0(n2809), .A1(xdata[345]), .Z(ofifoDataN[377]));
Q_AN02 U1646 ( .A0(n2641), .A1(xdata[378]), .Z(n2808));
Q_MX02 U1647 ( .S(n2642), .A0(n2808), .A1(xdata[346]), .Z(ofifoDataN[378]));
Q_AN02 U1648 ( .A0(n2641), .A1(xdata[379]), .Z(n2807));
Q_MX02 U1649 ( .S(n2642), .A0(n2807), .A1(xdata[347]), .Z(ofifoDataN[379]));
Q_AN02 U1650 ( .A0(n2641), .A1(xdata[380]), .Z(n2806));
Q_MX02 U1651 ( .S(n2642), .A0(n2806), .A1(xdata[348]), .Z(ofifoDataN[380]));
Q_AN02 U1652 ( .A0(n2641), .A1(xdata[381]), .Z(n2805));
Q_MX02 U1653 ( .S(n2642), .A0(n2805), .A1(xdata[349]), .Z(ofifoDataN[381]));
Q_AN02 U1654 ( .A0(n2641), .A1(xdata[382]), .Z(n2804));
Q_MX02 U1655 ( .S(n2642), .A0(n2804), .A1(xdata[350]), .Z(ofifoDataN[382]));
Q_AN02 U1656 ( .A0(n2641), .A1(xdata[383]), .Z(n2803));
Q_MX02 U1657 ( .S(n2642), .A0(n2803), .A1(xdata[351]), .Z(ofifoDataN[383]));
Q_AN02 U1658 ( .A0(n2641), .A1(xdata[384]), .Z(n2802));
Q_MX02 U1659 ( .S(n2642), .A0(n2802), .A1(xdata[352]), .Z(ofifoDataN[384]));
Q_AN02 U1660 ( .A0(n2641), .A1(xdata[385]), .Z(n2801));
Q_MX02 U1661 ( .S(n2642), .A0(n2801), .A1(xdata[353]), .Z(ofifoDataN[385]));
Q_AN02 U1662 ( .A0(n2641), .A1(xdata[386]), .Z(n2800));
Q_MX02 U1663 ( .S(n2642), .A0(n2800), .A1(xdata[354]), .Z(ofifoDataN[386]));
Q_AN02 U1664 ( .A0(n2641), .A1(xdata[387]), .Z(n2799));
Q_MX02 U1665 ( .S(n2642), .A0(n2799), .A1(xdata[355]), .Z(ofifoDataN[387]));
Q_AN02 U1666 ( .A0(n2641), .A1(xdata[388]), .Z(n2798));
Q_MX02 U1667 ( .S(n2642), .A0(n2798), .A1(xdata[356]), .Z(ofifoDataN[388]));
Q_AN02 U1668 ( .A0(n2641), .A1(xdata[389]), .Z(n2797));
Q_MX02 U1669 ( .S(n2642), .A0(n2797), .A1(xdata[357]), .Z(ofifoDataN[389]));
Q_AN02 U1670 ( .A0(n2641), .A1(xdata[390]), .Z(n2796));
Q_MX02 U1671 ( .S(n2642), .A0(n2796), .A1(xdata[358]), .Z(ofifoDataN[390]));
Q_AN02 U1672 ( .A0(n2641), .A1(xdata[391]), .Z(n2795));
Q_MX02 U1673 ( .S(n2642), .A0(n2795), .A1(xdata[359]), .Z(ofifoDataN[391]));
Q_AN02 U1674 ( .A0(n2641), .A1(xdata[392]), .Z(n2794));
Q_MX02 U1675 ( .S(n2642), .A0(n2794), .A1(xdata[360]), .Z(ofifoDataN[392]));
Q_AN02 U1676 ( .A0(n2641), .A1(xdata[393]), .Z(n2793));
Q_MX02 U1677 ( .S(n2642), .A0(n2793), .A1(xdata[361]), .Z(ofifoDataN[393]));
Q_AN02 U1678 ( .A0(n2641), .A1(xdata[394]), .Z(n2792));
Q_MX02 U1679 ( .S(n2642), .A0(n2792), .A1(xdata[362]), .Z(ofifoDataN[394]));
Q_AN02 U1680 ( .A0(n2641), .A1(xdata[395]), .Z(n2791));
Q_MX02 U1681 ( .S(n2642), .A0(n2791), .A1(xdata[363]), .Z(ofifoDataN[395]));
Q_AN02 U1682 ( .A0(n2641), .A1(xdata[396]), .Z(n2790));
Q_MX02 U1683 ( .S(n2642), .A0(n2790), .A1(xdata[364]), .Z(ofifoDataN[396]));
Q_AN02 U1684 ( .A0(n2641), .A1(xdata[397]), .Z(n2789));
Q_MX02 U1685 ( .S(n2642), .A0(n2789), .A1(xdata[365]), .Z(ofifoDataN[397]));
Q_AN02 U1686 ( .A0(n2641), .A1(xdata[398]), .Z(n2788));
Q_MX02 U1687 ( .S(n2642), .A0(n2788), .A1(xdata[366]), .Z(ofifoDataN[398]));
Q_AN02 U1688 ( .A0(n2641), .A1(xdata[399]), .Z(n2787));
Q_MX02 U1689 ( .S(n2642), .A0(n2787), .A1(xdata[367]), .Z(ofifoDataN[399]));
Q_AN02 U1690 ( .A0(n2641), .A1(xdata[400]), .Z(n2786));
Q_MX02 U1691 ( .S(n2642), .A0(n2786), .A1(xdata[368]), .Z(ofifoDataN[400]));
Q_AN02 U1692 ( .A0(n2641), .A1(xdata[401]), .Z(n2785));
Q_MX02 U1693 ( .S(n2642), .A0(n2785), .A1(xdata[369]), .Z(ofifoDataN[401]));
Q_AN02 U1694 ( .A0(n2641), .A1(xdata[402]), .Z(n2784));
Q_MX02 U1695 ( .S(n2642), .A0(n2784), .A1(xdata[370]), .Z(ofifoDataN[402]));
Q_AN02 U1696 ( .A0(n2641), .A1(xdata[403]), .Z(n2783));
Q_MX02 U1697 ( .S(n2642), .A0(n2783), .A1(xdata[371]), .Z(ofifoDataN[403]));
Q_AN02 U1698 ( .A0(n2641), .A1(xdata[404]), .Z(n2782));
Q_MX02 U1699 ( .S(n2642), .A0(n2782), .A1(xdata[372]), .Z(ofifoDataN[404]));
Q_AN02 U1700 ( .A0(n2641), .A1(xdata[405]), .Z(n2781));
Q_MX02 U1701 ( .S(n2642), .A0(n2781), .A1(xdata[373]), .Z(ofifoDataN[405]));
Q_AN02 U1702 ( .A0(n2641), .A1(xdata[406]), .Z(n2780));
Q_MX02 U1703 ( .S(n2642), .A0(n2780), .A1(xdata[374]), .Z(ofifoDataN[406]));
Q_AN02 U1704 ( .A0(n2641), .A1(xdata[407]), .Z(n2779));
Q_MX02 U1705 ( .S(n2642), .A0(n2779), .A1(xdata[375]), .Z(ofifoDataN[407]));
Q_AN02 U1706 ( .A0(n2641), .A1(xdata[408]), .Z(n2778));
Q_MX02 U1707 ( .S(n2642), .A0(n2778), .A1(xdata[376]), .Z(ofifoDataN[408]));
Q_AN02 U1708 ( .A0(n2641), .A1(xdata[409]), .Z(n2777));
Q_MX02 U1709 ( .S(n2642), .A0(n2777), .A1(xdata[377]), .Z(ofifoDataN[409]));
Q_AN02 U1710 ( .A0(n2641), .A1(xdata[410]), .Z(n2776));
Q_MX02 U1711 ( .S(n2642), .A0(n2776), .A1(xdata[378]), .Z(ofifoDataN[410]));
Q_AN02 U1712 ( .A0(n2641), .A1(xdata[411]), .Z(n2775));
Q_MX02 U1713 ( .S(n2642), .A0(n2775), .A1(xdata[379]), .Z(ofifoDataN[411]));
Q_AN02 U1714 ( .A0(n2641), .A1(xdata[412]), .Z(n2774));
Q_MX02 U1715 ( .S(n2642), .A0(n2774), .A1(xdata[380]), .Z(ofifoDataN[412]));
Q_AN02 U1716 ( .A0(n2641), .A1(xdata[413]), .Z(n2773));
Q_MX02 U1717 ( .S(n2642), .A0(n2773), .A1(xdata[381]), .Z(ofifoDataN[413]));
Q_AN02 U1718 ( .A0(n2641), .A1(xdata[414]), .Z(n2772));
Q_MX02 U1719 ( .S(n2642), .A0(n2772), .A1(xdata[382]), .Z(ofifoDataN[414]));
Q_AN02 U1720 ( .A0(n2641), .A1(xdata[415]), .Z(n2771));
Q_MX02 U1721 ( .S(n2642), .A0(n2771), .A1(xdata[383]), .Z(ofifoDataN[415]));
Q_AN02 U1722 ( .A0(n2641), .A1(xdata[416]), .Z(n2770));
Q_MX02 U1723 ( .S(n2642), .A0(n2770), .A1(xdata[384]), .Z(ofifoDataN[416]));
Q_AN02 U1724 ( .A0(n2641), .A1(xdata[417]), .Z(n2769));
Q_MX02 U1725 ( .S(n2642), .A0(n2769), .A1(xdata[385]), .Z(ofifoDataN[417]));
Q_AN02 U1726 ( .A0(n2641), .A1(xdata[418]), .Z(n2768));
Q_MX02 U1727 ( .S(n2642), .A0(n2768), .A1(xdata[386]), .Z(ofifoDataN[418]));
Q_AN02 U1728 ( .A0(n2641), .A1(xdata[419]), .Z(n2767));
Q_MX02 U1729 ( .S(n2642), .A0(n2767), .A1(xdata[387]), .Z(ofifoDataN[419]));
Q_AN02 U1730 ( .A0(n2641), .A1(xdata[420]), .Z(n2766));
Q_MX02 U1731 ( .S(n2642), .A0(n2766), .A1(xdata[388]), .Z(ofifoDataN[420]));
Q_AN02 U1732 ( .A0(n2641), .A1(xdata[421]), .Z(n2765));
Q_MX02 U1733 ( .S(n2642), .A0(n2765), .A1(xdata[389]), .Z(ofifoDataN[421]));
Q_AN02 U1734 ( .A0(n2641), .A1(xdata[422]), .Z(n2764));
Q_MX02 U1735 ( .S(n2642), .A0(n2764), .A1(xdata[390]), .Z(ofifoDataN[422]));
Q_AN02 U1736 ( .A0(n2641), .A1(xdata[423]), .Z(n2763));
Q_MX02 U1737 ( .S(n2642), .A0(n2763), .A1(xdata[391]), .Z(ofifoDataN[423]));
Q_AN02 U1738 ( .A0(n2641), .A1(xdata[424]), .Z(n2762));
Q_MX02 U1739 ( .S(n2642), .A0(n2762), .A1(xdata[392]), .Z(ofifoDataN[424]));
Q_AN02 U1740 ( .A0(n2641), .A1(xdata[425]), .Z(n2761));
Q_MX02 U1741 ( .S(n2642), .A0(n2761), .A1(xdata[393]), .Z(ofifoDataN[425]));
Q_AN02 U1742 ( .A0(n2641), .A1(xdata[426]), .Z(n2760));
Q_MX02 U1743 ( .S(n2642), .A0(n2760), .A1(xdata[394]), .Z(ofifoDataN[426]));
Q_AN02 U1744 ( .A0(n2641), .A1(xdata[427]), .Z(n2759));
Q_MX02 U1745 ( .S(n2642), .A0(n2759), .A1(xdata[395]), .Z(ofifoDataN[427]));
Q_AN02 U1746 ( .A0(n2641), .A1(xdata[428]), .Z(n2758));
Q_MX02 U1747 ( .S(n2642), .A0(n2758), .A1(xdata[396]), .Z(ofifoDataN[428]));
Q_AN02 U1748 ( .A0(n2641), .A1(xdata[429]), .Z(n2757));
Q_MX02 U1749 ( .S(n2642), .A0(n2757), .A1(xdata[397]), .Z(ofifoDataN[429]));
Q_AN02 U1750 ( .A0(n2641), .A1(xdata[430]), .Z(n2756));
Q_MX02 U1751 ( .S(n2642), .A0(n2756), .A1(xdata[398]), .Z(ofifoDataN[430]));
Q_AN02 U1752 ( .A0(n2641), .A1(xdata[431]), .Z(n2755));
Q_MX02 U1753 ( .S(n2642), .A0(n2755), .A1(xdata[399]), .Z(ofifoDataN[431]));
Q_AN02 U1754 ( .A0(n2641), .A1(xdata[432]), .Z(n2754));
Q_MX02 U1755 ( .S(n2642), .A0(n2754), .A1(xdata[400]), .Z(ofifoDataN[432]));
Q_AN02 U1756 ( .A0(n2641), .A1(xdata[433]), .Z(n2753));
Q_MX02 U1757 ( .S(n2642), .A0(n2753), .A1(xdata[401]), .Z(ofifoDataN[433]));
Q_AN02 U1758 ( .A0(n2641), .A1(xdata[434]), .Z(n2752));
Q_MX02 U1759 ( .S(n2642), .A0(n2752), .A1(xdata[402]), .Z(ofifoDataN[434]));
Q_AN02 U1760 ( .A0(n2641), .A1(xdata[435]), .Z(n2751));
Q_MX02 U1761 ( .S(n2642), .A0(n2751), .A1(xdata[403]), .Z(ofifoDataN[435]));
Q_AN02 U1762 ( .A0(n2641), .A1(xdata[436]), .Z(n2750));
Q_MX02 U1763 ( .S(n2642), .A0(n2750), .A1(xdata[404]), .Z(ofifoDataN[436]));
Q_AN02 U1764 ( .A0(n2641), .A1(xdata[437]), .Z(n2749));
Q_MX02 U1765 ( .S(n2642), .A0(n2749), .A1(xdata[405]), .Z(ofifoDataN[437]));
Q_AN02 U1766 ( .A0(n2641), .A1(xdata[438]), .Z(n2748));
Q_MX02 U1767 ( .S(n2642), .A0(n2748), .A1(xdata[406]), .Z(ofifoDataN[438]));
Q_AN02 U1768 ( .A0(n2641), .A1(xdata[439]), .Z(n2747));
Q_MX02 U1769 ( .S(n2642), .A0(n2747), .A1(xdata[407]), .Z(ofifoDataN[439]));
Q_AN02 U1770 ( .A0(n2641), .A1(xdata[440]), .Z(n2746));
Q_MX02 U1771 ( .S(n2642), .A0(n2746), .A1(xdata[408]), .Z(ofifoDataN[440]));
Q_AN02 U1772 ( .A0(n2641), .A1(xdata[441]), .Z(n2745));
Q_MX02 U1773 ( .S(n2642), .A0(n2745), .A1(xdata[409]), .Z(ofifoDataN[441]));
Q_AN02 U1774 ( .A0(n2641), .A1(xdata[442]), .Z(n2744));
Q_MX02 U1775 ( .S(n2642), .A0(n2744), .A1(xdata[410]), .Z(ofifoDataN[442]));
Q_AN02 U1776 ( .A0(n2641), .A1(xdata[443]), .Z(n2743));
Q_MX02 U1777 ( .S(n2642), .A0(n2743), .A1(xdata[411]), .Z(ofifoDataN[443]));
Q_AN02 U1778 ( .A0(n2641), .A1(xdata[444]), .Z(n2742));
Q_MX02 U1779 ( .S(n2642), .A0(n2742), .A1(xdata[412]), .Z(ofifoDataN[444]));
Q_AN02 U1780 ( .A0(n2641), .A1(xdata[445]), .Z(n2741));
Q_MX02 U1781 ( .S(n2642), .A0(n2741), .A1(xdata[413]), .Z(ofifoDataN[445]));
Q_AN02 U1782 ( .A0(n2641), .A1(xdata[446]), .Z(n2740));
Q_MX02 U1783 ( .S(n2642), .A0(n2740), .A1(xdata[414]), .Z(ofifoDataN[446]));
Q_AN02 U1784 ( .A0(n2641), .A1(xdata[447]), .Z(n2739));
Q_MX02 U1785 ( .S(n2642), .A0(n2739), .A1(xdata[415]), .Z(ofifoDataN[447]));
Q_AN02 U1786 ( .A0(n2641), .A1(xdata[448]), .Z(n2738));
Q_MX02 U1787 ( .S(n2642), .A0(n2738), .A1(xdata[416]), .Z(ofifoDataN[448]));
Q_AN02 U1788 ( .A0(n2641), .A1(xdata[449]), .Z(n2737));
Q_MX02 U1789 ( .S(n2642), .A0(n2737), .A1(xdata[417]), .Z(ofifoDataN[449]));
Q_AN02 U1790 ( .A0(n2641), .A1(xdata[450]), .Z(n2736));
Q_MX02 U1791 ( .S(n2642), .A0(n2736), .A1(xdata[418]), .Z(ofifoDataN[450]));
Q_AN02 U1792 ( .A0(n2641), .A1(xdata[451]), .Z(n2735));
Q_MX02 U1793 ( .S(n2642), .A0(n2735), .A1(xdata[419]), .Z(ofifoDataN[451]));
Q_AN02 U1794 ( .A0(n2641), .A1(xdata[452]), .Z(n2734));
Q_MX02 U1795 ( .S(n2642), .A0(n2734), .A1(xdata[420]), .Z(ofifoDataN[452]));
Q_AN02 U1796 ( .A0(n2641), .A1(xdata[453]), .Z(n2733));
Q_MX02 U1797 ( .S(n2642), .A0(n2733), .A1(xdata[421]), .Z(ofifoDataN[453]));
Q_AN02 U1798 ( .A0(n2641), .A1(xdata[454]), .Z(n2732));
Q_MX02 U1799 ( .S(n2642), .A0(n2732), .A1(xdata[422]), .Z(ofifoDataN[454]));
Q_AN02 U1800 ( .A0(n2641), .A1(xdata[455]), .Z(n2731));
Q_MX02 U1801 ( .S(n2642), .A0(n2731), .A1(xdata[423]), .Z(ofifoDataN[455]));
Q_AN02 U1802 ( .A0(n2641), .A1(xdata[456]), .Z(n2730));
Q_MX02 U1803 ( .S(n2642), .A0(n2730), .A1(xdata[424]), .Z(ofifoDataN[456]));
Q_AN02 U1804 ( .A0(n2641), .A1(xdata[457]), .Z(n2729));
Q_MX02 U1805 ( .S(n2642), .A0(n2729), .A1(xdata[425]), .Z(ofifoDataN[457]));
Q_AN02 U1806 ( .A0(n2641), .A1(xdata[458]), .Z(n2728));
Q_MX02 U1807 ( .S(n2642), .A0(n2728), .A1(xdata[426]), .Z(ofifoDataN[458]));
Q_AN02 U1808 ( .A0(n2641), .A1(xdata[459]), .Z(n2727));
Q_MX02 U1809 ( .S(n2642), .A0(n2727), .A1(xdata[427]), .Z(ofifoDataN[459]));
Q_AN02 U1810 ( .A0(n2641), .A1(xdata[460]), .Z(n2726));
Q_MX02 U1811 ( .S(n2642), .A0(n2726), .A1(xdata[428]), .Z(ofifoDataN[460]));
Q_AN02 U1812 ( .A0(n2641), .A1(xdata[461]), .Z(n2725));
Q_MX02 U1813 ( .S(n2642), .A0(n2725), .A1(xdata[429]), .Z(ofifoDataN[461]));
Q_AN02 U1814 ( .A0(n2641), .A1(xdata[462]), .Z(n2724));
Q_MX02 U1815 ( .S(n2642), .A0(n2724), .A1(xdata[430]), .Z(ofifoDataN[462]));
Q_AN02 U1816 ( .A0(n2641), .A1(xdata[463]), .Z(n2723));
Q_MX02 U1817 ( .S(n2642), .A0(n2723), .A1(xdata[431]), .Z(ofifoDataN[463]));
Q_AN02 U1818 ( .A0(n2641), .A1(xdata[464]), .Z(n2722));
Q_MX02 U1819 ( .S(n2642), .A0(n2722), .A1(xdata[432]), .Z(ofifoDataN[464]));
Q_AN02 U1820 ( .A0(n2641), .A1(xdata[465]), .Z(n2721));
Q_MX02 U1821 ( .S(n2642), .A0(n2721), .A1(xdata[433]), .Z(ofifoDataN[465]));
Q_AN02 U1822 ( .A0(n2641), .A1(xdata[466]), .Z(n2720));
Q_MX02 U1823 ( .S(n2642), .A0(n2720), .A1(xdata[434]), .Z(ofifoDataN[466]));
Q_AN02 U1824 ( .A0(n2641), .A1(xdata[467]), .Z(n2719));
Q_MX02 U1825 ( .S(n2642), .A0(n2719), .A1(xdata[435]), .Z(ofifoDataN[467]));
Q_AN02 U1826 ( .A0(n2641), .A1(xdata[468]), .Z(n2718));
Q_MX02 U1827 ( .S(n2642), .A0(n2718), .A1(xdata[436]), .Z(ofifoDataN[468]));
Q_AN02 U1828 ( .A0(n2641), .A1(xdata[469]), .Z(n2717));
Q_MX02 U1829 ( .S(n2642), .A0(n2717), .A1(xdata[437]), .Z(ofifoDataN[469]));
Q_AN02 U1830 ( .A0(n2641), .A1(xdata[470]), .Z(n2716));
Q_MX02 U1831 ( .S(n2642), .A0(n2716), .A1(xdata[438]), .Z(ofifoDataN[470]));
Q_AN02 U1832 ( .A0(n2641), .A1(xdata[471]), .Z(n2715));
Q_MX02 U1833 ( .S(n2642), .A0(n2715), .A1(xdata[439]), .Z(ofifoDataN[471]));
Q_AN02 U1834 ( .A0(n2641), .A1(xdata[472]), .Z(n2714));
Q_MX02 U1835 ( .S(n2642), .A0(n2714), .A1(xdata[440]), .Z(ofifoDataN[472]));
Q_AN02 U1836 ( .A0(n2641), .A1(xdata[473]), .Z(n2713));
Q_MX02 U1837 ( .S(n2642), .A0(n2713), .A1(xdata[441]), .Z(ofifoDataN[473]));
Q_AN02 U1838 ( .A0(n2641), .A1(xdata[474]), .Z(n2712));
Q_MX02 U1839 ( .S(n2642), .A0(n2712), .A1(xdata[442]), .Z(ofifoDataN[474]));
Q_AN02 U1840 ( .A0(n2641), .A1(xdata[475]), .Z(n2711));
Q_MX02 U1841 ( .S(n2642), .A0(n2711), .A1(xdata[443]), .Z(ofifoDataN[475]));
Q_AN02 U1842 ( .A0(n2641), .A1(xdata[476]), .Z(n2710));
Q_MX02 U1843 ( .S(n2642), .A0(n2710), .A1(xdata[444]), .Z(ofifoDataN[476]));
Q_AN02 U1844 ( .A0(n2641), .A1(xdata[477]), .Z(n2709));
Q_MX02 U1845 ( .S(n2642), .A0(n2709), .A1(xdata[445]), .Z(ofifoDataN[477]));
Q_AN02 U1846 ( .A0(n2641), .A1(xdata[478]), .Z(n2708));
Q_MX02 U1847 ( .S(n2642), .A0(n2708), .A1(xdata[446]), .Z(ofifoDataN[478]));
Q_AN02 U1848 ( .A0(n2641), .A1(xdata[479]), .Z(n2707));
Q_MX02 U1849 ( .S(n2642), .A0(n2707), .A1(xdata[447]), .Z(ofifoDataN[479]));
Q_AN02 U1850 ( .A0(n2641), .A1(xdata[480]), .Z(n2706));
Q_MX02 U1851 ( .S(n2642), .A0(n2706), .A1(xdata[448]), .Z(ofifoDataN[480]));
Q_AN02 U1852 ( .A0(n2641), .A1(xdata[481]), .Z(n2705));
Q_MX02 U1853 ( .S(n2642), .A0(n2705), .A1(xdata[449]), .Z(ofifoDataN[481]));
Q_AN02 U1854 ( .A0(n2641), .A1(xdata[482]), .Z(n2704));
Q_MX02 U1855 ( .S(n2642), .A0(n2704), .A1(xdata[450]), .Z(ofifoDataN[482]));
Q_AN02 U1856 ( .A0(n2641), .A1(xdata[483]), .Z(n2703));
Q_MX02 U1857 ( .S(n2642), .A0(n2703), .A1(xdata[451]), .Z(ofifoDataN[483]));
Q_AN02 U1858 ( .A0(n2641), .A1(xdata[484]), .Z(n2702));
Q_MX02 U1859 ( .S(n2642), .A0(n2702), .A1(xdata[452]), .Z(ofifoDataN[484]));
Q_AN02 U1860 ( .A0(n2641), .A1(xdata[485]), .Z(n2701));
Q_MX02 U1861 ( .S(n2642), .A0(n2701), .A1(xdata[453]), .Z(ofifoDataN[485]));
Q_AN02 U1862 ( .A0(n2641), .A1(xdata[486]), .Z(n2700));
Q_MX02 U1863 ( .S(n2642), .A0(n2700), .A1(xdata[454]), .Z(ofifoDataN[486]));
Q_AN02 U1864 ( .A0(n2641), .A1(xdata[487]), .Z(n2699));
Q_MX02 U1865 ( .S(n2642), .A0(n2699), .A1(xdata[455]), .Z(ofifoDataN[487]));
Q_AN02 U1866 ( .A0(n2641), .A1(xdata[488]), .Z(n2698));
Q_MX02 U1867 ( .S(n2642), .A0(n2698), .A1(xdata[456]), .Z(ofifoDataN[488]));
Q_AN02 U1868 ( .A0(n2641), .A1(xdata[489]), .Z(n2697));
Q_MX02 U1869 ( .S(n2642), .A0(n2697), .A1(xdata[457]), .Z(ofifoDataN[489]));
Q_AN02 U1870 ( .A0(n2641), .A1(xdata[490]), .Z(n2696));
Q_MX02 U1871 ( .S(n2642), .A0(n2696), .A1(xdata[458]), .Z(ofifoDataN[490]));
Q_AN02 U1872 ( .A0(n2641), .A1(xdata[491]), .Z(n2695));
Q_MX02 U1873 ( .S(n2642), .A0(n2695), .A1(xdata[459]), .Z(ofifoDataN[491]));
Q_AN02 U1874 ( .A0(n2641), .A1(xdata[492]), .Z(n2694));
Q_MX02 U1875 ( .S(n2642), .A0(n2694), .A1(xdata[460]), .Z(ofifoDataN[492]));
Q_AN02 U1876 ( .A0(n2641), .A1(xdata[493]), .Z(n2693));
Q_MX02 U1877 ( .S(n2642), .A0(n2693), .A1(xdata[461]), .Z(ofifoDataN[493]));
Q_AN02 U1878 ( .A0(n2641), .A1(xdata[494]), .Z(n2692));
Q_MX02 U1879 ( .S(n2642), .A0(n2692), .A1(xdata[462]), .Z(ofifoDataN[494]));
Q_AN02 U1880 ( .A0(n2641), .A1(xdata[495]), .Z(n2691));
Q_MX02 U1881 ( .S(n2642), .A0(n2691), .A1(xdata[463]), .Z(ofifoDataN[495]));
Q_AN02 U1882 ( .A0(n2641), .A1(xdata[496]), .Z(n2690));
Q_MX02 U1883 ( .S(n2642), .A0(n2690), .A1(xdata[464]), .Z(ofifoDataN[496]));
Q_AN02 U1884 ( .A0(n2641), .A1(xdata[497]), .Z(n2689));
Q_MX02 U1885 ( .S(n2642), .A0(n2689), .A1(xdata[465]), .Z(ofifoDataN[497]));
Q_AN02 U1886 ( .A0(n2641), .A1(xdata[498]), .Z(n2688));
Q_MX02 U1887 ( .S(n2642), .A0(n2688), .A1(xdata[466]), .Z(ofifoDataN[498]));
Q_AN02 U1888 ( .A0(n2641), .A1(xdata[499]), .Z(n2687));
Q_MX02 U1889 ( .S(n2642), .A0(n2687), .A1(xdata[467]), .Z(ofifoDataN[499]));
Q_AN02 U1890 ( .A0(n2641), .A1(xdata[500]), .Z(n2686));
Q_MX02 U1891 ( .S(n2642), .A0(n2686), .A1(xdata[468]), .Z(ofifoDataN[500]));
Q_AN02 U1892 ( .A0(n2641), .A1(xdata[501]), .Z(n2685));
Q_MX02 U1893 ( .S(n2642), .A0(n2685), .A1(xdata[469]), .Z(ofifoDataN[501]));
Q_AN02 U1894 ( .A0(n2641), .A1(xdata[502]), .Z(n2684));
Q_MX02 U1895 ( .S(n2642), .A0(n2684), .A1(xdata[470]), .Z(ofifoDataN[502]));
Q_AN02 U1896 ( .A0(n2641), .A1(xdata[503]), .Z(n2683));
Q_MX02 U1897 ( .S(n2642), .A0(n2683), .A1(xdata[471]), .Z(ofifoDataN[503]));
Q_AN02 U1898 ( .A0(n2641), .A1(xdata[504]), .Z(n2682));
Q_MX02 U1899 ( .S(n2642), .A0(n2682), .A1(xdata[472]), .Z(ofifoDataN[504]));
Q_AN02 U1900 ( .A0(n2641), .A1(xdata[505]), .Z(n2681));
Q_MX02 U1901 ( .S(n2642), .A0(n2681), .A1(xdata[473]), .Z(ofifoDataN[505]));
Q_AN02 U1902 ( .A0(n2641), .A1(xdata[506]), .Z(n2680));
Q_MX02 U1903 ( .S(n2642), .A0(n2680), .A1(xdata[474]), .Z(ofifoDataN[506]));
Q_AN02 U1904 ( .A0(n2641), .A1(xdata[507]), .Z(n2679));
Q_MX02 U1905 ( .S(n2642), .A0(n2679), .A1(xdata[475]), .Z(ofifoDataN[507]));
Q_AN02 U1906 ( .A0(n2641), .A1(xdata[508]), .Z(n2678));
Q_MX02 U1907 ( .S(n2642), .A0(n2678), .A1(xdata[476]), .Z(ofifoDataN[508]));
Q_AN02 U1908 ( .A0(n2641), .A1(xdata[509]), .Z(n2677));
Q_MX02 U1909 ( .S(n2642), .A0(n2677), .A1(xdata[477]), .Z(ofifoDataN[509]));
Q_AN02 U1910 ( .A0(n2641), .A1(xdata[510]), .Z(n2676));
Q_MX02 U1911 ( .S(n2642), .A0(n2676), .A1(xdata[478]), .Z(ofifoDataN[510]));
Q_AN02 U1912 ( .A0(n2641), .A1(xdata[511]), .Z(n2675));
Q_MX02 U1913 ( .S(n2642), .A0(n2675), .A1(xdata[479]), .Z(ofifoDataN[511]));
Q_AN02 U1914 ( .A0(n2641), .A1(xdata[512]), .Z(n2674));
Q_MX02 U1915 ( .S(n2642), .A0(n2674), .A1(xdata[480]), .Z(ofifoDataN[512]));
Q_AN02 U1916 ( .A0(n2641), .A1(xdata[513]), .Z(n2673));
Q_MX02 U1917 ( .S(n2642), .A0(n2673), .A1(xdata[481]), .Z(ofifoDataN[513]));
Q_AN02 U1918 ( .A0(n2641), .A1(xdata[514]), .Z(n2672));
Q_MX02 U1919 ( .S(n2642), .A0(n2672), .A1(xdata[482]), .Z(ofifoDataN[514]));
Q_AN02 U1920 ( .A0(n2641), .A1(xdata[515]), .Z(n2671));
Q_MX02 U1921 ( .S(n2642), .A0(n2671), .A1(xdata[483]), .Z(ofifoDataN[515]));
Q_AN02 U1922 ( .A0(n2641), .A1(xdata[516]), .Z(n2670));
Q_MX02 U1923 ( .S(n2642), .A0(n2670), .A1(xdata[484]), .Z(ofifoDataN[516]));
Q_AN02 U1924 ( .A0(n2641), .A1(xdata[517]), .Z(n2669));
Q_MX02 U1925 ( .S(n2642), .A0(n2669), .A1(xdata[485]), .Z(ofifoDataN[517]));
Q_AN02 U1926 ( .A0(n2641), .A1(xdata[518]), .Z(n2668));
Q_MX02 U1927 ( .S(n2642), .A0(n2668), .A1(xdata[486]), .Z(ofifoDataN[518]));
Q_AN02 U1928 ( .A0(n2641), .A1(xdata[519]), .Z(n2667));
Q_MX02 U1929 ( .S(n2642), .A0(n2667), .A1(xdata[487]), .Z(ofifoDataN[519]));
Q_AN02 U1930 ( .A0(n2641), .A1(xdata[520]), .Z(n2666));
Q_MX02 U1931 ( .S(n2642), .A0(n2666), .A1(xdata[488]), .Z(ofifoDataN[520]));
Q_AN02 U1932 ( .A0(n2641), .A1(xdata[521]), .Z(n2665));
Q_MX02 U1933 ( .S(n2642), .A0(n2665), .A1(xdata[489]), .Z(ofifoDataN[521]));
Q_AN02 U1934 ( .A0(n2641), .A1(xdata[522]), .Z(n2664));
Q_MX02 U1935 ( .S(n2642), .A0(n2664), .A1(xdata[490]), .Z(ofifoDataN[522]));
Q_AN02 U1936 ( .A0(n2641), .A1(xdata[523]), .Z(n2663));
Q_MX02 U1937 ( .S(n2642), .A0(n2663), .A1(xdata[491]), .Z(ofifoDataN[523]));
Q_AN02 U1938 ( .A0(n2641), .A1(xdata[524]), .Z(n2662));
Q_MX02 U1939 ( .S(n2642), .A0(n2662), .A1(xdata[492]), .Z(ofifoDataN[524]));
Q_AN02 U1940 ( .A0(n2641), .A1(xdata[525]), .Z(n2661));
Q_MX02 U1941 ( .S(n2642), .A0(n2661), .A1(xdata[493]), .Z(ofifoDataN[525]));
Q_AN02 U1942 ( .A0(n2641), .A1(xdata[526]), .Z(n2660));
Q_MX02 U1943 ( .S(n2642), .A0(n2660), .A1(xdata[494]), .Z(ofifoDataN[526]));
Q_AN02 U1944 ( .A0(n2641), .A1(xdata[527]), .Z(n2659));
Q_MX02 U1945 ( .S(n2642), .A0(n2659), .A1(xdata[495]), .Z(ofifoDataN[527]));
Q_AN02 U1946 ( .A0(n2641), .A1(xdata[528]), .Z(n2658));
Q_MX02 U1947 ( .S(n2642), .A0(n2658), .A1(xdata[496]), .Z(ofifoDataN[528]));
Q_AN02 U1948 ( .A0(n2641), .A1(xdata[529]), .Z(n2657));
Q_MX02 U1949 ( .S(n2642), .A0(n2657), .A1(xdata[497]), .Z(ofifoDataN[529]));
Q_AN02 U1950 ( .A0(n2641), .A1(xdata[530]), .Z(n2656));
Q_MX02 U1951 ( .S(n2642), .A0(n2656), .A1(xdata[498]), .Z(ofifoDataN[530]));
Q_AN02 U1952 ( .A0(n2641), .A1(xdata[531]), .Z(n2655));
Q_MX02 U1953 ( .S(n2642), .A0(n2655), .A1(xdata[499]), .Z(ofifoDataN[531]));
Q_AN02 U1954 ( .A0(n2641), .A1(xdata[532]), .Z(n2654));
Q_MX02 U1955 ( .S(n2642), .A0(n2654), .A1(xdata[500]), .Z(ofifoDataN[532]));
Q_AN02 U1956 ( .A0(n2641), .A1(xdata[533]), .Z(n2653));
Q_MX02 U1957 ( .S(n2642), .A0(n2653), .A1(xdata[501]), .Z(ofifoDataN[533]));
Q_AN02 U1958 ( .A0(n2641), .A1(xdata[534]), .Z(n2652));
Q_MX02 U1959 ( .S(n2642), .A0(n2652), .A1(xdata[502]), .Z(ofifoDataN[534]));
Q_AN02 U1960 ( .A0(n2641), .A1(xdata[535]), .Z(n2651));
Q_MX02 U1961 ( .S(n2642), .A0(n2651), .A1(xdata[503]), .Z(ofifoDataN[535]));
Q_AN02 U1962 ( .A0(n2641), .A1(xdata[536]), .Z(n2650));
Q_MX02 U1963 ( .S(n2642), .A0(n2650), .A1(xdata[504]), .Z(ofifoDataN[536]));
Q_AN02 U1964 ( .A0(n2641), .A1(xdata[537]), .Z(n2649));
Q_MX02 U1965 ( .S(n2642), .A0(n2649), .A1(xdata[505]), .Z(ofifoDataN[537]));
Q_AN02 U1966 ( .A0(n2641), .A1(xdata[538]), .Z(n2648));
Q_MX02 U1967 ( .S(n2642), .A0(n2648), .A1(xdata[506]), .Z(ofifoDataN[538]));
Q_AN02 U1968 ( .A0(n2641), .A1(xdata[539]), .Z(n2647));
Q_MX02 U1969 ( .S(n2642), .A0(n2647), .A1(xdata[507]), .Z(ofifoDataN[539]));
Q_AN02 U1970 ( .A0(n2641), .A1(xdata[540]), .Z(n2646));
Q_MX02 U1971 ( .S(n2642), .A0(n2646), .A1(xdata[508]), .Z(ofifoDataN[540]));
Q_AN02 U1972 ( .A0(n2641), .A1(xdata[541]), .Z(n2645));
Q_MX02 U1973 ( .S(n2642), .A0(n2645), .A1(xdata[509]), .Z(ofifoDataN[541]));
Q_AN02 U1974 ( .A0(n2641), .A1(xdata[542]), .Z(n2644));
Q_MX02 U1975 ( .S(n2642), .A0(n2644), .A1(xdata[510]), .Z(ofifoDataN[542]));
Q_AN02 U1976 ( .A0(n2641), .A1(xdata[543]), .Z(n2643));
Q_MX02 U1977 ( .S(n2642), .A0(n2643), .A1(xdata[511]), .Z(ofifoDataN[543]));
Q_AN02 U1978 ( .A0(n2642), .A1(xdata[512]), .Z(ofifoDataN[544]));
Q_AN02 U1979 ( .A0(n2642), .A1(xdata[513]), .Z(ofifoDataN[545]));
Q_AN02 U1980 ( .A0(n2642), .A1(xdata[514]), .Z(ofifoDataN[546]));
Q_AN02 U1981 ( .A0(n2642), .A1(xdata[515]), .Z(ofifoDataN[547]));
Q_AN02 U1982 ( .A0(n2642), .A1(xdata[516]), .Z(ofifoDataN[548]));
Q_AN02 U1983 ( .A0(n2642), .A1(xdata[517]), .Z(ofifoDataN[549]));
Q_AN02 U1984 ( .A0(n2642), .A1(xdata[518]), .Z(ofifoDataN[550]));
Q_AN02 U1985 ( .A0(n2642), .A1(xdata[519]), .Z(ofifoDataN[551]));
Q_AN02 U1986 ( .A0(n2642), .A1(xdata[520]), .Z(ofifoDataN[552]));
Q_AN02 U1987 ( .A0(n2642), .A1(xdata[521]), .Z(ofifoDataN[553]));
Q_AN02 U1988 ( .A0(n2642), .A1(xdata[522]), .Z(ofifoDataN[554]));
Q_AN02 U1989 ( .A0(n2642), .A1(xdata[523]), .Z(ofifoDataN[555]));
Q_AN02 U1990 ( .A0(n2642), .A1(xdata[524]), .Z(ofifoDataN[556]));
Q_AN02 U1991 ( .A0(n2642), .A1(xdata[525]), .Z(ofifoDataN[557]));
Q_AN02 U1992 ( .A0(n2642), .A1(xdata[526]), .Z(ofifoDataN[558]));
Q_AN02 U1993 ( .A0(n2642), .A1(xdata[527]), .Z(ofifoDataN[559]));
Q_AN02 U1994 ( .A0(n2642), .A1(xdata[528]), .Z(ofifoDataN[560]));
Q_AN02 U1995 ( .A0(n2642), .A1(xdata[529]), .Z(ofifoDataN[561]));
Q_AN02 U1996 ( .A0(n2642), .A1(xdata[530]), .Z(ofifoDataN[562]));
Q_AN02 U1997 ( .A0(n2642), .A1(xdata[531]), .Z(ofifoDataN[563]));
Q_AN02 U1998 ( .A0(n2642), .A1(xdata[532]), .Z(ofifoDataN[564]));
Q_AN02 U1999 ( .A0(n2642), .A1(xdata[533]), .Z(ofifoDataN[565]));
Q_AN02 U2000 ( .A0(n2642), .A1(xdata[534]), .Z(ofifoDataN[566]));
Q_AN02 U2001 ( .A0(n2642), .A1(xdata[535]), .Z(ofifoDataN[567]));
Q_AN02 U2002 ( .A0(n2642), .A1(xdata[536]), .Z(ofifoDataN[568]));
Q_AN02 U2003 ( .A0(n2642), .A1(xdata[537]), .Z(ofifoDataN[569]));
Q_AN02 U2004 ( .A0(n2642), .A1(xdata[538]), .Z(ofifoDataN[570]));
Q_AN02 U2005 ( .A0(n2642), .A1(xdata[539]), .Z(ofifoDataN[571]));
Q_AN02 U2006 ( .A0(n2642), .A1(xdata[540]), .Z(ofifoDataN[572]));
Q_AN02 U2007 ( .A0(n2642), .A1(xdata[541]), .Z(ofifoDataN[573]));
Q_AN02 U2008 ( .A0(n2642), .A1(xdata[542]), .Z(ofifoDataN[574]));
Q_AN02 U2009 ( .A0(n2642), .A1(xdata[543]), .Z(ofifoDataN[575]));
Q_NR02 U2010 ( .A0(xc_top.GFReset), .A1(oFill[0]), .Z(n2641));
Q_AN02 U2011 ( .A0(n65), .A1(oFill[0]), .Z(n2642));
Q_AN03 U2012 ( .A0(GFreq), .A1(n2640), .A2(GFtsReq), .Z(GFtsAdd));
Q_INV U2013 ( .A(reqD), .Z(n2640));
Q_FDP0UA U2014 ( .D(wrtCnt[0]), .QTFCLK( ), .Q(wrtCntD[0]));
Q_FDP0UA U2015 ( .D(wrtCnt[1]), .QTFCLK( ), .Q(wrtCntD[1]));
Q_FDP0UA U2016 ( .D(wrtCnt[2]), .QTFCLK( ), .Q(wrtCntD[2]));
Q_FDP0UA U2017 ( .D(wrtCnt[3]), .QTFCLK( ), .Q(wrtCntD[3]));
Q_FDP0UA U2018 ( .D(wrtCnt[4]), .QTFCLK( ), .Q(wrtCntD[4]));
Q_FDP0UA U2019 ( .D(wrtCnt[5]), .QTFCLK( ), .Q(wrtCntD[5]));
Q_FDP0UA U2020 ( .D(wrtCnt[6]), .QTFCLK( ), .Q(wrtCntD[6]));
Q_FDP0UA U2021 ( .D(wrtCnt[7]), .QTFCLK( ), .Q(wrtCntD[7]));
Q_FDP0UA U2022 ( .D(wrtCnt[8]), .QTFCLK( ), .Q(wrtCntD[8]));
Q_FDP0UA U2023 ( .D(wrtCnt[9]), .QTFCLK( ), .Q(wrtCntD[9]));
Q_FDP0UA U2024 ( .D(wrtCnt[10]), .QTFCLK( ), .Q(wrtCntD[10]));
Q_FDP0UA U2025 ( .D(wrtCnt[11]), .QTFCLK( ), .Q(wrtCntD[11]));
Q_FDP0UA U2026 ( .D(wrtCnt[12]), .QTFCLK( ), .Q(wrtCntD[12]));
Q_FDP0UA U2027 ( .D(wrtCnt[13]), .QTFCLK( ), .Q(wrtCntD[13]));
Q_FDP0UA U2028 ( .D(wrtCnt[14]), .QTFCLK( ), .Q(wrtCntD[14]));
Q_FDP0UA U2029 ( .D(wrtCnt[15]), .QTFCLK( ), .Q(wrtCntD[15]));
Q_FDP0UA U2030 ( .D(wrtCnt[16]), .QTFCLK( ), .Q(wrtCntD[16]));
Q_FDP0UA U2031 ( .D(wrtCnt[17]), .QTFCLK( ), .Q(wrtCntD[17]));
Q_FDP0UA U2032 ( .D(wrtCnt[18]), .QTFCLK( ), .Q(wrtCntD[18]));
Q_FDP0UA U2033 ( .D(wrtCnt[19]), .QTFCLK( ), .Q(wrtCntD[19]));
Q_FDP0UA U2034 ( .D(wrtCnt[20]), .QTFCLK( ), .Q(wrtCntD[20]));
Q_FDP0UA U2035 ( .D(wrtCnt[21]), .QTFCLK( ), .Q(wrtCntD[21]));
Q_FDP0UA U2036 ( .D(wrtCnt[22]), .QTFCLK( ), .Q(wrtCntD[22]));
Q_FDP0UA U2037 ( .D(wrtCnt[23]), .QTFCLK( ), .Q(wrtCntD[23]));
Q_FDP0UA U2038 ( .D(wrtCnt[24]), .QTFCLK( ), .Q(wrtCntD[24]));
Q_FDP0UA U2039 ( .D(wrtCnt[25]), .QTFCLK( ), .Q(wrtCntD[25]));
Q_FDP0UA U2040 ( .D(wrtCnt[26]), .QTFCLK( ), .Q(wrtCntD[26]));
Q_FDP0UA U2041 ( .D(wrtCnt[27]), .QTFCLK( ), .Q(wrtCntD[27]));
Q_FDP0UA U2042 ( .D(wrtCnt[28]), .QTFCLK( ), .Q(wrtCntD[28]));
Q_FDP0UA U2043 ( .D(wrtCnt[29]), .QTFCLK( ), .Q(wrtCntD[29]));
Q_FDP0UA U2044 ( .D(wrtCnt[30]), .QTFCLK( ), .Q(wrtCntD[30]));
Q_FDP0UA U2045 ( .D(wrtCnt[31]), .QTFCLK( ), .Q(wrtCntD[31]));
Q_FDP0UA U2046 ( .D(wrtCnt[32]), .QTFCLK( ), .Q(wrtCntD[32]));
Q_FDP0UA U2047 ( .D(wrtCnt[33]), .QTFCLK( ), .Q(wrtCntD[33]));
Q_FDP0UA U2048 ( .D(wrtCnt[34]), .QTFCLK( ), .Q(wrtCntD[34]));
Q_FDP0UA U2049 ( .D(wrtCnt[35]), .QTFCLK( ), .Q(wrtCntD[35]));
Q_FDP0UA U2050 ( .D(wrtCnt[36]), .QTFCLK( ), .Q(wrtCntD[36]));
Q_FDP0UA U2051 ( .D(wrtCnt[37]), .QTFCLK( ), .Q(wrtCntD[37]));
Q_FDP0UA U2052 ( .D(wrtCnt[38]), .QTFCLK( ), .Q(wrtCntD[38]));
Q_FDP0UA U2053 ( .D(wrtCnt[39]), .QTFCLK( ), .Q(wrtCntD[39]));
Q_FDP0UA U2054 ( .D(wrtCnt[40]), .QTFCLK( ), .Q(wrtCntD[40]));
Q_FDP0UA U2055 ( .D(wrtCnt[41]), .QTFCLK( ), .Q(wrtCntD[41]));
Q_FDP0UA U2056 ( .D(wrtCnt[42]), .QTFCLK( ), .Q(wrtCntD[42]));
Q_FDP0UA U2057 ( .D(wrtCnt[43]), .QTFCLK( ), .Q(wrtCntD[43]));
Q_FDP0UA U2058 ( .D(wrtCnt[44]), .QTFCLK( ), .Q(wrtCntD[44]));
Q_FDP0UA U2059 ( .D(wrtCnt[45]), .QTFCLK( ), .Q(wrtCntD[45]));
Q_FDP0UA U2060 ( .D(wrtCnt[46]), .QTFCLK( ), .Q(wrtCntD[46]));
Q_FDP0UA U2061 ( .D(wrtCnt[47]), .QTFCLK( ), .Q(wrtCntD[47]));
Q_FDP0UA U2062 ( .D(wrtCnt[48]), .QTFCLK( ), .Q(wrtCntD[48]));
Q_FDP0UA U2063 ( .D(wrtCnt[49]), .QTFCLK( ), .Q(wrtCntD[49]));
Q_FDP0UA U2064 ( .D(wrtCnt[50]), .QTFCLK( ), .Q(wrtCntD[50]));
Q_FDP0UA U2065 ( .D(wrtCnt[51]), .QTFCLK( ), .Q(wrtCntD[51]));
Q_FDP0UA U2066 ( .D(wrtCnt[52]), .QTFCLK( ), .Q(wrtCntD[52]));
Q_FDP0UA U2067 ( .D(wrtCnt[53]), .QTFCLK( ), .Q(wrtCntD[53]));
Q_FDP0UA U2068 ( .D(wrtCnt[54]), .QTFCLK( ), .Q(wrtCntD[54]));
Q_FDP0UA U2069 ( .D(wrtCnt[55]), .QTFCLK( ), .Q(wrtCntD[55]));
Q_FDP0UA U2070 ( .D(wrtCnt[56]), .QTFCLK( ), .Q(wrtCntD[56]));
Q_FDP0UA U2071 ( .D(wrtCnt[57]), .QTFCLK( ), .Q(wrtCntD[57]));
Q_FDP0UA U2072 ( .D(wrtCnt[58]), .QTFCLK( ), .Q(wrtCntD[58]));
Q_FDP0UA U2073 ( .D(wrtCnt[59]), .QTFCLK( ), .Q(wrtCntD[59]));
Q_FDP0UA U2074 ( .D(wrtCnt[60]), .QTFCLK( ), .Q(wrtCntD[60]));
Q_FDP0UA U2075 ( .D(wrtCnt[61]), .QTFCLK( ), .Q(wrtCntD[61]));
Q_FDP0UA U2076 ( .D(wrtCnt[62]), .QTFCLK( ), .Q(wrtCntD[62]));
Q_FDP0UA U2077 ( .D(wrtCnt[63]), .QTFCLK( ), .Q(wrtCntD[63]));
Q_FDP0UA U2078 ( .D(n2638), .QTFCLK( ), .Q(reqD));
Q_AN02 U2079 ( .A0(n65), .A1(GFreq), .Z(n2638));
Q_OA21 U2080 ( .A0(reqD), .A1(GFtsAdd), .B0(n2637), .Z(n784));
Q_INV U2081 ( .A(xc_top.GFLock1), .Z(n2637));
Q_INV U2082 ( .A(GFcbid[0]), .Z(n2636));
Q_AN03 U2083 ( .A0(GFcbid[19]), .A1(GFcbid[18]), .A2(GFcbid[17]), .Z(n2635));
Q_AN03 U2084 ( .A0(GFcbid[16]), .A1(GFcbid[15]), .A2(GFcbid[14]), .Z(n2634));
Q_AN03 U2085 ( .A0(GFcbid[13]), .A1(GFcbid[12]), .A2(GFcbid[11]), .Z(n2633));
Q_AN03 U2086 ( .A0(GFcbid[10]), .A1(GFcbid[9]), .A2(GFcbid[8]), .Z(n2632));
Q_AN03 U2087 ( .A0(GFcbid[7]), .A1(GFcbid[6]), .A2(GFcbid[5]), .Z(n2631));
Q_AN03 U2088 ( .A0(GFcbid[4]), .A1(GFcbid[3]), .A2(GFcbid[2]), .Z(n2630));
Q_AN03 U2089 ( .A0(GFcbid[1]), .A1(n2636), .A2(n2635), .Z(n2629));
Q_AN03 U2090 ( .A0(n2634), .A1(n2633), .A2(n2632), .Z(n2628));
Q_AN03 U2091 ( .A0(n2631), .A1(n2630), .A2(n2629), .Z(n2627));
Q_AN02 U2092 ( .A0(n2628), .A1(n2627), .Z(n788));
Q_OR02 U2093 ( .A0(GFlen[9]), .A1(GFlen[8]), .Z(n2626));
Q_OR03 U2094 ( .A0(GFlen[11]), .A1(GFlen[10]), .A2(n2626), .Z(n2625));
Q_OR03 U2095 ( .A0(GFlen[7]), .A1(GFlen[6]), .A2(GFlen[5]), .Z(n2624));
Q_OR02 U2096 ( .A0(GFlen[1]), .A1(GFlen[0]), .Z(n2623));
Q_OR02 U2097 ( .A0(GFlen[3]), .A1(GFlen[2]), .Z(n2622));
Q_OA21 U2098 ( .A0(n2622), .A1(n2623), .B0(GFlen[4]), .Z(n2621));
Q_OR03 U2099 ( .A0(n2625), .A1(n2624), .A2(n2621), .Z(n783));
Q_INV U2100 ( .A(n788), .Z(n2619));
Q_AN02 U2101 ( .A0(n2619), .A1(GFidata[32]), .Z(n2618));
Q_AN02 U2102 ( .A0(n2619), .A1(GFidata[33]), .Z(n2617));
Q_AN02 U2103 ( .A0(n2619), .A1(GFidata[34]), .Z(n2616));
Q_AN02 U2104 ( .A0(n2619), .A1(GFidata[35]), .Z(n2615));
Q_AN02 U2105 ( .A0(n2619), .A1(GFidata[36]), .Z(n2614));
Q_AN02 U2106 ( .A0(n2619), .A1(GFidata[37]), .Z(n2613));
Q_AN02 U2107 ( .A0(n2619), .A1(GFidata[38]), .Z(n2612));
Q_AN02 U2108 ( .A0(n2619), .A1(GFidata[39]), .Z(n2611));
Q_AN02 U2109 ( .A0(n2619), .A1(GFidata[40]), .Z(n2610));
Q_AN02 U2110 ( .A0(n2619), .A1(GFidata[41]), .Z(n2609));
Q_AN02 U2111 ( .A0(n2619), .A1(GFidata[42]), .Z(n2608));
Q_AN02 U2112 ( .A0(n2619), .A1(GFidata[43]), .Z(n2607));
Q_AN02 U2113 ( .A0(n2619), .A1(GFidata[44]), .Z(n2606));
Q_AN02 U2114 ( .A0(n2619), .A1(GFidata[45]), .Z(n2605));
Q_AN02 U2115 ( .A0(n2619), .A1(GFidata[46]), .Z(n2604));
Q_AN02 U2116 ( .A0(n2619), .A1(GFidata[47]), .Z(n2603));
Q_AN02 U2117 ( .A0(n2619), .A1(GFidata[48]), .Z(n2602));
Q_AN02 U2118 ( .A0(n2619), .A1(GFidata[49]), .Z(n2601));
Q_AN02 U2119 ( .A0(n2619), .A1(GFidata[50]), .Z(n2600));
Q_AN02 U2120 ( .A0(n2619), .A1(GFidata[51]), .Z(n2599));
Q_AN02 U2121 ( .A0(n2619), .A1(GFidata[52]), .Z(n2598));
Q_AN02 U2122 ( .A0(n2619), .A1(GFidata[53]), .Z(n2597));
Q_AN02 U2123 ( .A0(n2619), .A1(GFidata[54]), .Z(n2596));
Q_AN02 U2124 ( .A0(n2619), .A1(GFidata[55]), .Z(n2595));
Q_AN02 U2125 ( .A0(n2619), .A1(GFidata[56]), .Z(n2594));
Q_AN02 U2126 ( .A0(n2619), .A1(GFidata[57]), .Z(n2593));
Q_AN02 U2127 ( .A0(n2619), .A1(GFidata[58]), .Z(n2592));
Q_AN02 U2128 ( .A0(n2619), .A1(GFidata[59]), .Z(n2591));
Q_AN02 U2129 ( .A0(n2619), .A1(GFidata[60]), .Z(n2590));
Q_AN02 U2130 ( .A0(n2619), .A1(GFidata[61]), .Z(n2589));
Q_AN02 U2131 ( .A0(n2619), .A1(GFidata[62]), .Z(n2588));
Q_AN02 U2132 ( .A0(n2619), .A1(GFidata[63]), .Z(n2587));
Q_AN02 U2133 ( .A0(n2619), .A1(GFidata[64]), .Z(n2586));
Q_AN02 U2134 ( .A0(n2619), .A1(GFidata[65]), .Z(n2585));
Q_AN02 U2135 ( .A0(n2619), .A1(GFidata[66]), .Z(n2584));
Q_AN02 U2136 ( .A0(n2619), .A1(GFidata[67]), .Z(n2583));
Q_AN02 U2137 ( .A0(n2619), .A1(GFidata[68]), .Z(n2582));
Q_AN02 U2138 ( .A0(n2619), .A1(GFidata[69]), .Z(n2581));
Q_AN02 U2139 ( .A0(n2619), .A1(GFidata[70]), .Z(n2580));
Q_AN02 U2140 ( .A0(n2619), .A1(GFidata[71]), .Z(n2579));
Q_AN02 U2141 ( .A0(n2619), .A1(GFidata[72]), .Z(n2578));
Q_AN02 U2142 ( .A0(n2619), .A1(GFidata[73]), .Z(n2577));
Q_AN02 U2143 ( .A0(n2619), .A1(GFidata[74]), .Z(n2576));
Q_AN02 U2144 ( .A0(n2619), .A1(GFidata[75]), .Z(n2575));
Q_AN02 U2145 ( .A0(n2619), .A1(GFidata[76]), .Z(n2574));
Q_AN02 U2146 ( .A0(n2619), .A1(GFidata[77]), .Z(n2573));
Q_AN02 U2147 ( .A0(n2619), .A1(GFidata[78]), .Z(n2572));
Q_AN02 U2148 ( .A0(n2619), .A1(GFidata[79]), .Z(n2571));
Q_AN02 U2149 ( .A0(n2619), .A1(GFidata[80]), .Z(n2570));
Q_AN02 U2150 ( .A0(n2619), .A1(GFidata[81]), .Z(n2569));
Q_AN02 U2151 ( .A0(n2619), .A1(GFidata[82]), .Z(n2568));
Q_AN02 U2152 ( .A0(n2619), .A1(GFidata[83]), .Z(n2567));
Q_AN02 U2153 ( .A0(n2619), .A1(GFidata[84]), .Z(n2566));
Q_AN02 U2154 ( .A0(n2619), .A1(GFidata[85]), .Z(n2565));
Q_AN02 U2155 ( .A0(n2619), .A1(GFidata[86]), .Z(n2564));
Q_AN02 U2156 ( .A0(n2619), .A1(GFidata[87]), .Z(n2563));
Q_AN02 U2157 ( .A0(n2619), .A1(GFidata[88]), .Z(n2562));
Q_AN02 U2158 ( .A0(n2619), .A1(GFidata[89]), .Z(n2561));
Q_AN02 U2159 ( .A0(n2619), .A1(GFidata[90]), .Z(n2560));
Q_AN02 U2160 ( .A0(n2619), .A1(GFidata[91]), .Z(n2559));
Q_AN02 U2161 ( .A0(n2619), .A1(GFidata[92]), .Z(n2558));
Q_AN02 U2162 ( .A0(n2619), .A1(GFidata[93]), .Z(n2557));
Q_AN02 U2163 ( .A0(n2619), .A1(GFidata[94]), .Z(n2556));
Q_AN02 U2164 ( .A0(n2619), .A1(GFidata[95]), .Z(n2555));
Q_AN02 U2165 ( .A0(n2619), .A1(GFidata[96]), .Z(n2554));
Q_AN02 U2166 ( .A0(n2619), .A1(GFidata[97]), .Z(n2553));
Q_AN02 U2167 ( .A0(n2619), .A1(GFidata[98]), .Z(n2552));
Q_AN02 U2168 ( .A0(n2619), .A1(GFidata[99]), .Z(n2551));
Q_AN02 U2169 ( .A0(n2619), .A1(GFidata[100]), .Z(n2550));
Q_AN02 U2170 ( .A0(n2619), .A1(GFidata[101]), .Z(n2549));
Q_AN02 U2171 ( .A0(n2619), .A1(GFidata[102]), .Z(n2548));
Q_AN02 U2172 ( .A0(n2619), .A1(GFidata[103]), .Z(n2547));
Q_AN02 U2173 ( .A0(n2619), .A1(GFidata[104]), .Z(n2546));
Q_AN02 U2174 ( .A0(n2619), .A1(GFidata[105]), .Z(n2545));
Q_AN02 U2175 ( .A0(n2619), .A1(GFidata[106]), .Z(n2544));
Q_AN02 U2176 ( .A0(n2619), .A1(GFidata[107]), .Z(n2543));
Q_AN02 U2177 ( .A0(n2619), .A1(GFidata[108]), .Z(n2542));
Q_AN02 U2178 ( .A0(n2619), .A1(GFidata[109]), .Z(n2541));
Q_AN02 U2179 ( .A0(n2619), .A1(GFidata[110]), .Z(n2540));
Q_AN02 U2180 ( .A0(n2619), .A1(GFidata[111]), .Z(n2539));
Q_AN02 U2181 ( .A0(n2619), .A1(GFidata[112]), .Z(n2538));
Q_AN02 U2182 ( .A0(n2619), .A1(GFidata[113]), .Z(n2537));
Q_AN02 U2183 ( .A0(n2619), .A1(GFidata[114]), .Z(n2536));
Q_AN02 U2184 ( .A0(n2619), .A1(GFidata[115]), .Z(n2535));
Q_AN02 U2185 ( .A0(n2619), .A1(GFidata[116]), .Z(n2534));
Q_AN02 U2186 ( .A0(n2619), .A1(GFidata[117]), .Z(n2533));
Q_AN02 U2187 ( .A0(n2619), .A1(GFidata[118]), .Z(n2532));
Q_AN02 U2188 ( .A0(n2619), .A1(GFidata[119]), .Z(n2531));
Q_AN02 U2189 ( .A0(n2619), .A1(GFidata[120]), .Z(n2530));
Q_AN02 U2190 ( .A0(n2619), .A1(GFidata[121]), .Z(n2529));
Q_AN02 U2191 ( .A0(n2619), .A1(GFidata[122]), .Z(n2528));
Q_AN02 U2192 ( .A0(n2619), .A1(GFidata[123]), .Z(n2527));
Q_AN02 U2193 ( .A0(n2619), .A1(GFidata[124]), .Z(n2526));
Q_AN02 U2194 ( .A0(n2619), .A1(GFidata[125]), .Z(n2525));
Q_AN02 U2195 ( .A0(n2619), .A1(GFidata[126]), .Z(n2524));
Q_AN02 U2196 ( .A0(n2619), .A1(GFidata[127]), .Z(n2523));
Q_AN02 U2197 ( .A0(n2619), .A1(GFidata[128]), .Z(n2522));
Q_AN02 U2198 ( .A0(n2619), .A1(GFidata[129]), .Z(n2521));
Q_AN02 U2199 ( .A0(n2619), .A1(GFidata[130]), .Z(n2520));
Q_AN02 U2200 ( .A0(n2619), .A1(GFidata[131]), .Z(n2519));
Q_AN02 U2201 ( .A0(n2619), .A1(GFidata[132]), .Z(n2518));
Q_AN02 U2202 ( .A0(n2619), .A1(GFidata[133]), .Z(n2517));
Q_AN02 U2203 ( .A0(n2619), .A1(GFidata[134]), .Z(n2516));
Q_AN02 U2204 ( .A0(n2619), .A1(GFidata[135]), .Z(n2515));
Q_AN02 U2205 ( .A0(n2619), .A1(GFidata[136]), .Z(n2514));
Q_AN02 U2206 ( .A0(n2619), .A1(GFidata[137]), .Z(n2513));
Q_AN02 U2207 ( .A0(n2619), .A1(GFidata[138]), .Z(n2512));
Q_AN02 U2208 ( .A0(n2619), .A1(GFidata[139]), .Z(n2511));
Q_AN02 U2209 ( .A0(n2619), .A1(GFidata[140]), .Z(n2510));
Q_AN02 U2210 ( .A0(n2619), .A1(GFidata[141]), .Z(n2509));
Q_AN02 U2211 ( .A0(n2619), .A1(GFidata[142]), .Z(n2508));
Q_AN02 U2212 ( .A0(n2619), .A1(GFidata[143]), .Z(n2507));
Q_AN02 U2213 ( .A0(n2619), .A1(GFidata[144]), .Z(n2506));
Q_AN02 U2214 ( .A0(n2619), .A1(GFidata[145]), .Z(n2505));
Q_AN02 U2215 ( .A0(n2619), .A1(GFidata[146]), .Z(n2504));
Q_AN02 U2216 ( .A0(n2619), .A1(GFidata[147]), .Z(n2503));
Q_AN02 U2217 ( .A0(n2619), .A1(GFidata[148]), .Z(n2502));
Q_AN02 U2218 ( .A0(n2619), .A1(GFidata[149]), .Z(n2501));
Q_AN02 U2219 ( .A0(n2619), .A1(GFidata[150]), .Z(n2500));
Q_AN02 U2220 ( .A0(n2619), .A1(GFidata[151]), .Z(n2499));
Q_AN02 U2221 ( .A0(n2619), .A1(GFidata[152]), .Z(n2498));
Q_AN02 U2222 ( .A0(n2619), .A1(GFidata[153]), .Z(n2497));
Q_AN02 U2223 ( .A0(n2619), .A1(GFidata[154]), .Z(n2496));
Q_AN02 U2224 ( .A0(n2619), .A1(GFidata[155]), .Z(n2495));
Q_AN02 U2225 ( .A0(n2619), .A1(GFidata[156]), .Z(n2494));
Q_AN02 U2226 ( .A0(n2619), .A1(GFidata[157]), .Z(n2493));
Q_AN02 U2227 ( .A0(n2619), .A1(GFidata[158]), .Z(n2492));
Q_AN02 U2228 ( .A0(n2619), .A1(GFidata[159]), .Z(n2491));
Q_AN02 U2229 ( .A0(n2619), .A1(GFidata[160]), .Z(n2490));
Q_AN02 U2230 ( .A0(n2619), .A1(GFidata[161]), .Z(n2489));
Q_AN02 U2231 ( .A0(n2619), .A1(GFidata[162]), .Z(n2488));
Q_AN02 U2232 ( .A0(n2619), .A1(GFidata[163]), .Z(n2487));
Q_AN02 U2233 ( .A0(n2619), .A1(GFidata[164]), .Z(n2486));
Q_AN02 U2234 ( .A0(n2619), .A1(GFidata[165]), .Z(n2485));
Q_AN02 U2235 ( .A0(n2619), .A1(GFidata[166]), .Z(n2484));
Q_AN02 U2236 ( .A0(n2619), .A1(GFidata[167]), .Z(n2483));
Q_AN02 U2237 ( .A0(n2619), .A1(GFidata[168]), .Z(n2482));
Q_AN02 U2238 ( .A0(n2619), .A1(GFidata[169]), .Z(n2481));
Q_AN02 U2239 ( .A0(n2619), .A1(GFidata[170]), .Z(n2480));
Q_AN02 U2240 ( .A0(n2619), .A1(GFidata[171]), .Z(n2479));
Q_AN02 U2241 ( .A0(n2619), .A1(GFidata[172]), .Z(n2478));
Q_AN02 U2242 ( .A0(n2619), .A1(GFidata[173]), .Z(n2477));
Q_AN02 U2243 ( .A0(n2619), .A1(GFidata[174]), .Z(n2476));
Q_AN02 U2244 ( .A0(n2619), .A1(GFidata[175]), .Z(n2475));
Q_AN02 U2245 ( .A0(n2619), .A1(GFidata[176]), .Z(n2474));
Q_AN02 U2246 ( .A0(n2619), .A1(GFidata[177]), .Z(n2473));
Q_AN02 U2247 ( .A0(n2619), .A1(GFidata[178]), .Z(n2472));
Q_AN02 U2248 ( .A0(n2619), .A1(GFidata[179]), .Z(n2471));
Q_AN02 U2249 ( .A0(n2619), .A1(GFidata[180]), .Z(n2470));
Q_AN02 U2250 ( .A0(n2619), .A1(GFidata[181]), .Z(n2469));
Q_AN02 U2251 ( .A0(n2619), .A1(GFidata[182]), .Z(n2468));
Q_AN02 U2252 ( .A0(n2619), .A1(GFidata[183]), .Z(n2467));
Q_AN02 U2253 ( .A0(n2619), .A1(GFidata[184]), .Z(n2466));
Q_AN02 U2254 ( .A0(n2619), .A1(GFidata[185]), .Z(n2465));
Q_AN02 U2255 ( .A0(n2619), .A1(GFidata[186]), .Z(n2464));
Q_AN02 U2256 ( .A0(n2619), .A1(GFidata[187]), .Z(n2463));
Q_AN02 U2257 ( .A0(n2619), .A1(GFidata[188]), .Z(n2462));
Q_AN02 U2258 ( .A0(n2619), .A1(GFidata[189]), .Z(n2461));
Q_AN02 U2259 ( .A0(n2619), .A1(GFidata[190]), .Z(n2460));
Q_AN02 U2260 ( .A0(n2619), .A1(GFidata[191]), .Z(n2459));
Q_AN02 U2261 ( .A0(n2619), .A1(GFidata[192]), .Z(n2458));
Q_AN02 U2262 ( .A0(n2619), .A1(GFidata[193]), .Z(n2457));
Q_AN02 U2263 ( .A0(n2619), .A1(GFidata[194]), .Z(n2456));
Q_AN02 U2264 ( .A0(n2619), .A1(GFidata[195]), .Z(n2455));
Q_AN02 U2265 ( .A0(n2619), .A1(GFidata[196]), .Z(n2454));
Q_AN02 U2266 ( .A0(n2619), .A1(GFidata[197]), .Z(n2453));
Q_AN02 U2267 ( .A0(n2619), .A1(GFidata[198]), .Z(n2452));
Q_AN02 U2268 ( .A0(n2619), .A1(GFidata[199]), .Z(n2451));
Q_AN02 U2269 ( .A0(n2619), .A1(GFidata[200]), .Z(n2450));
Q_AN02 U2270 ( .A0(n2619), .A1(GFidata[201]), .Z(n2449));
Q_AN02 U2271 ( .A0(n2619), .A1(GFidata[202]), .Z(n2448));
Q_AN02 U2272 ( .A0(n2619), .A1(GFidata[203]), .Z(n2447));
Q_AN02 U2273 ( .A0(n2619), .A1(GFidata[204]), .Z(n2446));
Q_AN02 U2274 ( .A0(n2619), .A1(GFidata[205]), .Z(n2445));
Q_AN02 U2275 ( .A0(n2619), .A1(GFidata[206]), .Z(n2444));
Q_AN02 U2276 ( .A0(n2619), .A1(GFidata[207]), .Z(n2443));
Q_AN02 U2277 ( .A0(n2619), .A1(GFidata[208]), .Z(n2442));
Q_AN02 U2278 ( .A0(n2619), .A1(GFidata[209]), .Z(n2441));
Q_AN02 U2279 ( .A0(n2619), .A1(GFidata[210]), .Z(n2440));
Q_AN02 U2280 ( .A0(n2619), .A1(GFidata[211]), .Z(n2439));
Q_AN02 U2281 ( .A0(n2619), .A1(GFidata[212]), .Z(n2438));
Q_AN02 U2282 ( .A0(n2619), .A1(GFidata[213]), .Z(n2437));
Q_AN02 U2283 ( .A0(n2619), .A1(GFidata[214]), .Z(n2436));
Q_AN02 U2284 ( .A0(n2619), .A1(GFidata[215]), .Z(n2435));
Q_AN02 U2285 ( .A0(n2619), .A1(GFidata[216]), .Z(n2434));
Q_AN02 U2286 ( .A0(n2619), .A1(GFidata[217]), .Z(n2433));
Q_AN02 U2287 ( .A0(n2619), .A1(GFidata[218]), .Z(n2432));
Q_AN02 U2288 ( .A0(n2619), .A1(GFidata[219]), .Z(n2431));
Q_AN02 U2289 ( .A0(n2619), .A1(GFidata[220]), .Z(n2430));
Q_AN02 U2290 ( .A0(n2619), .A1(GFidata[221]), .Z(n2429));
Q_AN02 U2291 ( .A0(n2619), .A1(GFidata[222]), .Z(n2428));
Q_AN02 U2292 ( .A0(n2619), .A1(GFidata[223]), .Z(n2427));
Q_AN02 U2293 ( .A0(n2619), .A1(GFidata[224]), .Z(n2426));
Q_AN02 U2294 ( .A0(n2619), .A1(GFidata[225]), .Z(n2425));
Q_AN02 U2295 ( .A0(n2619), .A1(GFidata[226]), .Z(n2424));
Q_AN02 U2296 ( .A0(n2619), .A1(GFidata[227]), .Z(n2423));
Q_AN02 U2297 ( .A0(n2619), .A1(GFidata[228]), .Z(n2422));
Q_AN02 U2298 ( .A0(n2619), .A1(GFidata[229]), .Z(n2421));
Q_AN02 U2299 ( .A0(n2619), .A1(GFidata[230]), .Z(n2420));
Q_AN02 U2300 ( .A0(n2619), .A1(GFidata[231]), .Z(n2419));
Q_AN02 U2301 ( .A0(n2619), .A1(GFidata[232]), .Z(n2418));
Q_AN02 U2302 ( .A0(n2619), .A1(GFidata[233]), .Z(n2417));
Q_AN02 U2303 ( .A0(n2619), .A1(GFidata[234]), .Z(n2416));
Q_AN02 U2304 ( .A0(n2619), .A1(GFidata[235]), .Z(n2415));
Q_AN02 U2305 ( .A0(n2619), .A1(GFidata[236]), .Z(n2414));
Q_AN02 U2306 ( .A0(n2619), .A1(GFidata[237]), .Z(n2413));
Q_AN02 U2307 ( .A0(n2619), .A1(GFidata[238]), .Z(n2412));
Q_AN02 U2308 ( .A0(n2619), .A1(GFidata[239]), .Z(n2411));
Q_AN02 U2309 ( .A0(n2619), .A1(GFidata[240]), .Z(n2410));
Q_AN02 U2310 ( .A0(n2619), .A1(GFidata[241]), .Z(n2409));
Q_AN02 U2311 ( .A0(n2619), .A1(GFidata[242]), .Z(n2408));
Q_AN02 U2312 ( .A0(n2619), .A1(GFidata[243]), .Z(n2407));
Q_AN02 U2313 ( .A0(n2619), .A1(GFidata[244]), .Z(n2406));
Q_AN02 U2314 ( .A0(n2619), .A1(GFidata[245]), .Z(n2405));
Q_AN02 U2315 ( .A0(n2619), .A1(GFidata[246]), .Z(n2404));
Q_AN02 U2316 ( .A0(n2619), .A1(GFidata[247]), .Z(n2403));
Q_AN02 U2317 ( .A0(n2619), .A1(GFidata[248]), .Z(n2402));
Q_AN02 U2318 ( .A0(n2619), .A1(GFidata[249]), .Z(n2401));
Q_AN02 U2319 ( .A0(n2619), .A1(GFidata[250]), .Z(n2400));
Q_AN02 U2320 ( .A0(n2619), .A1(GFidata[251]), .Z(n2399));
Q_AN02 U2321 ( .A0(n2619), .A1(GFidata[252]), .Z(n2398));
Q_AN02 U2322 ( .A0(n2619), .A1(GFidata[253]), .Z(n2397));
Q_AN02 U2323 ( .A0(n2619), .A1(GFidata[254]), .Z(n2396));
Q_AN02 U2324 ( .A0(n2619), .A1(GFidata[255]), .Z(n2395));
Q_AN02 U2325 ( .A0(n2619), .A1(GFidata[256]), .Z(n2394));
Q_AN02 U2326 ( .A0(n2619), .A1(GFidata[257]), .Z(n2393));
Q_AN02 U2327 ( .A0(n2619), .A1(GFidata[258]), .Z(n2392));
Q_AN02 U2328 ( .A0(n2619), .A1(GFidata[259]), .Z(n2391));
Q_AN02 U2329 ( .A0(n2619), .A1(GFidata[260]), .Z(n2390));
Q_AN02 U2330 ( .A0(n2619), .A1(GFidata[261]), .Z(n2389));
Q_AN02 U2331 ( .A0(n2619), .A1(GFidata[262]), .Z(n2388));
Q_AN02 U2332 ( .A0(n2619), .A1(GFidata[263]), .Z(n2387));
Q_AN02 U2333 ( .A0(n2619), .A1(GFidata[264]), .Z(n2386));
Q_AN02 U2334 ( .A0(n2619), .A1(GFidata[265]), .Z(n2385));
Q_AN02 U2335 ( .A0(n2619), .A1(GFidata[266]), .Z(n2384));
Q_AN02 U2336 ( .A0(n2619), .A1(GFidata[267]), .Z(n2383));
Q_AN02 U2337 ( .A0(n2619), .A1(GFidata[268]), .Z(n2382));
Q_AN02 U2338 ( .A0(n2619), .A1(GFidata[269]), .Z(n2381));
Q_AN02 U2339 ( .A0(n2619), .A1(GFidata[270]), .Z(n2380));
Q_AN02 U2340 ( .A0(n2619), .A1(GFidata[271]), .Z(n2379));
Q_AN02 U2341 ( .A0(n2619), .A1(GFidata[272]), .Z(n2378));
Q_AN02 U2342 ( .A0(n2619), .A1(GFidata[273]), .Z(n2377));
Q_AN02 U2343 ( .A0(n2619), .A1(GFidata[274]), .Z(n2376));
Q_AN02 U2344 ( .A0(n2619), .A1(GFidata[275]), .Z(n2375));
Q_AN02 U2345 ( .A0(n2619), .A1(GFidata[276]), .Z(n2374));
Q_AN02 U2346 ( .A0(n2619), .A1(GFidata[277]), .Z(n2373));
Q_AN02 U2347 ( .A0(n2619), .A1(GFidata[278]), .Z(n2372));
Q_AN02 U2348 ( .A0(n2619), .A1(GFidata[279]), .Z(n2371));
Q_AN02 U2349 ( .A0(n2619), .A1(GFidata[280]), .Z(n2370));
Q_AN02 U2350 ( .A0(n2619), .A1(GFidata[281]), .Z(n2369));
Q_AN02 U2351 ( .A0(n2619), .A1(GFidata[282]), .Z(n2368));
Q_AN02 U2352 ( .A0(n2619), .A1(GFidata[283]), .Z(n2367));
Q_AN02 U2353 ( .A0(n2619), .A1(GFidata[284]), .Z(n2366));
Q_AN02 U2354 ( .A0(n2619), .A1(GFidata[285]), .Z(n2365));
Q_AN02 U2355 ( .A0(n2619), .A1(GFidata[286]), .Z(n2364));
Q_AN02 U2356 ( .A0(n2619), .A1(GFidata[287]), .Z(n2363));
Q_AN02 U2357 ( .A0(n2619), .A1(GFidata[288]), .Z(n2362));
Q_AN02 U2358 ( .A0(n2619), .A1(GFidata[289]), .Z(n2361));
Q_AN02 U2359 ( .A0(n2619), .A1(GFidata[290]), .Z(n2360));
Q_AN02 U2360 ( .A0(n2619), .A1(GFidata[291]), .Z(n2359));
Q_AN02 U2361 ( .A0(n2619), .A1(GFidata[292]), .Z(n2358));
Q_AN02 U2362 ( .A0(n2619), .A1(GFidata[293]), .Z(n2357));
Q_AN02 U2363 ( .A0(n2619), .A1(GFidata[294]), .Z(n2356));
Q_AN02 U2364 ( .A0(n2619), .A1(GFidata[295]), .Z(n2355));
Q_AN02 U2365 ( .A0(n2619), .A1(GFidata[296]), .Z(n2354));
Q_AN02 U2366 ( .A0(n2619), .A1(GFidata[297]), .Z(n2353));
Q_AN02 U2367 ( .A0(n2619), .A1(GFidata[298]), .Z(n2352));
Q_AN02 U2368 ( .A0(n2619), .A1(GFidata[299]), .Z(n2351));
Q_AN02 U2369 ( .A0(n2619), .A1(GFidata[300]), .Z(n2350));
Q_AN02 U2370 ( .A0(n2619), .A1(GFidata[301]), .Z(n2349));
Q_AN02 U2371 ( .A0(n2619), .A1(GFidata[302]), .Z(n2348));
Q_AN02 U2372 ( .A0(n2619), .A1(GFidata[303]), .Z(n2347));
Q_AN02 U2373 ( .A0(n2619), .A1(GFidata[304]), .Z(n2346));
Q_AN02 U2374 ( .A0(n2619), .A1(GFidata[305]), .Z(n2345));
Q_AN02 U2375 ( .A0(n2619), .A1(GFidata[306]), .Z(n2344));
Q_AN02 U2376 ( .A0(n2619), .A1(GFidata[307]), .Z(n2343));
Q_AN02 U2377 ( .A0(n2619), .A1(GFidata[308]), .Z(n2342));
Q_AN02 U2378 ( .A0(n2619), .A1(GFidata[309]), .Z(n2341));
Q_AN02 U2379 ( .A0(n2619), .A1(GFidata[310]), .Z(n2340));
Q_AN02 U2380 ( .A0(n2619), .A1(GFidata[311]), .Z(n2339));
Q_AN02 U2381 ( .A0(n2619), .A1(GFidata[312]), .Z(n2338));
Q_AN02 U2382 ( .A0(n2619), .A1(GFidata[313]), .Z(n2337));
Q_AN02 U2383 ( .A0(n2619), .A1(GFidata[314]), .Z(n2336));
Q_AN02 U2384 ( .A0(n2619), .A1(GFidata[315]), .Z(n2335));
Q_AN02 U2385 ( .A0(n2619), .A1(GFidata[316]), .Z(n2334));
Q_AN02 U2386 ( .A0(n2619), .A1(GFidata[317]), .Z(n2333));
Q_AN02 U2387 ( .A0(n2619), .A1(GFidata[318]), .Z(n2332));
Q_AN02 U2388 ( .A0(n2619), .A1(GFidata[319]), .Z(n2331));
Q_AN02 U2389 ( .A0(n2619), .A1(GFidata[320]), .Z(n2330));
Q_AN02 U2390 ( .A0(n2619), .A1(GFidata[321]), .Z(n2329));
Q_AN02 U2391 ( .A0(n2619), .A1(GFidata[322]), .Z(n2328));
Q_AN02 U2392 ( .A0(n2619), .A1(GFidata[323]), .Z(n2327));
Q_AN02 U2393 ( .A0(n2619), .A1(GFidata[324]), .Z(n2326));
Q_AN02 U2394 ( .A0(n2619), .A1(GFidata[325]), .Z(n2325));
Q_AN02 U2395 ( .A0(n2619), .A1(GFidata[326]), .Z(n2324));
Q_AN02 U2396 ( .A0(n2619), .A1(GFidata[327]), .Z(n2323));
Q_AN02 U2397 ( .A0(n2619), .A1(GFidata[328]), .Z(n2322));
Q_AN02 U2398 ( .A0(n2619), .A1(GFidata[329]), .Z(n2321));
Q_AN02 U2399 ( .A0(n2619), .A1(GFidata[330]), .Z(n2320));
Q_AN02 U2400 ( .A0(n2619), .A1(GFidata[331]), .Z(n2319));
Q_AN02 U2401 ( .A0(n2619), .A1(GFidata[332]), .Z(n2318));
Q_AN02 U2402 ( .A0(n2619), .A1(GFidata[333]), .Z(n2317));
Q_AN02 U2403 ( .A0(n2619), .A1(GFidata[334]), .Z(n2316));
Q_AN02 U2404 ( .A0(n2619), .A1(GFidata[335]), .Z(n2315));
Q_AN02 U2405 ( .A0(n2619), .A1(GFidata[336]), .Z(n2314));
Q_AN02 U2406 ( .A0(n2619), .A1(GFidata[337]), .Z(n2313));
Q_AN02 U2407 ( .A0(n2619), .A1(GFidata[338]), .Z(n2312));
Q_AN02 U2408 ( .A0(n2619), .A1(GFidata[339]), .Z(n2311));
Q_AN02 U2409 ( .A0(n2619), .A1(GFidata[340]), .Z(n2310));
Q_AN02 U2410 ( .A0(n2619), .A1(GFidata[341]), .Z(n2309));
Q_AN02 U2411 ( .A0(n2619), .A1(GFidata[342]), .Z(n2308));
Q_AN02 U2412 ( .A0(n2619), .A1(GFidata[343]), .Z(n2307));
Q_AN02 U2413 ( .A0(n2619), .A1(GFidata[344]), .Z(n2306));
Q_AN02 U2414 ( .A0(n2619), .A1(GFidata[345]), .Z(n2305));
Q_AN02 U2415 ( .A0(n2619), .A1(GFidata[346]), .Z(n2304));
Q_AN02 U2416 ( .A0(n2619), .A1(GFidata[347]), .Z(n2303));
Q_AN02 U2417 ( .A0(n2619), .A1(GFidata[348]), .Z(n2302));
Q_AN02 U2418 ( .A0(n2619), .A1(GFidata[349]), .Z(n2301));
Q_AN02 U2419 ( .A0(n2619), .A1(GFidata[350]), .Z(n2300));
Q_AN02 U2420 ( .A0(n2619), .A1(GFidata[351]), .Z(n2299));
Q_AN02 U2421 ( .A0(n2619), .A1(GFidata[352]), .Z(n2298));
Q_AN02 U2422 ( .A0(n2619), .A1(GFidata[353]), .Z(n2297));
Q_AN02 U2423 ( .A0(n2619), .A1(GFidata[354]), .Z(n2296));
Q_AN02 U2424 ( .A0(n2619), .A1(GFidata[355]), .Z(n2295));
Q_AN02 U2425 ( .A0(n2619), .A1(GFidata[356]), .Z(n2294));
Q_AN02 U2426 ( .A0(n2619), .A1(GFidata[357]), .Z(n2293));
Q_AN02 U2427 ( .A0(n2619), .A1(GFidata[358]), .Z(n2292));
Q_AN02 U2428 ( .A0(n2619), .A1(GFidata[359]), .Z(n2291));
Q_AN02 U2429 ( .A0(n2619), .A1(GFidata[360]), .Z(n2290));
Q_AN02 U2430 ( .A0(n2619), .A1(GFidata[361]), .Z(n2289));
Q_AN02 U2431 ( .A0(n2619), .A1(GFidata[362]), .Z(n2288));
Q_AN02 U2432 ( .A0(n2619), .A1(GFidata[363]), .Z(n2287));
Q_AN02 U2433 ( .A0(n2619), .A1(GFidata[364]), .Z(n2286));
Q_AN02 U2434 ( .A0(n2619), .A1(GFidata[365]), .Z(n2285));
Q_AN02 U2435 ( .A0(n2619), .A1(GFidata[366]), .Z(n2284));
Q_AN02 U2436 ( .A0(n2619), .A1(GFidata[367]), .Z(n2283));
Q_AN02 U2437 ( .A0(n2619), .A1(GFidata[368]), .Z(n2282));
Q_AN02 U2438 ( .A0(n2619), .A1(GFidata[369]), .Z(n2281));
Q_AN02 U2439 ( .A0(n2619), .A1(GFidata[370]), .Z(n2280));
Q_AN02 U2440 ( .A0(n2619), .A1(GFidata[371]), .Z(n2279));
Q_AN02 U2441 ( .A0(n2619), .A1(GFidata[372]), .Z(n2278));
Q_AN02 U2442 ( .A0(n2619), .A1(GFidata[373]), .Z(n2277));
Q_AN02 U2443 ( .A0(n2619), .A1(GFidata[374]), .Z(n2276));
Q_AN02 U2444 ( .A0(n2619), .A1(GFidata[375]), .Z(n2275));
Q_AN02 U2445 ( .A0(n2619), .A1(GFidata[376]), .Z(n2274));
Q_AN02 U2446 ( .A0(n2619), .A1(GFidata[377]), .Z(n2273));
Q_AN02 U2447 ( .A0(n2619), .A1(GFidata[378]), .Z(n2272));
Q_AN02 U2448 ( .A0(n2619), .A1(GFidata[379]), .Z(n2271));
Q_AN02 U2449 ( .A0(n2619), .A1(GFidata[380]), .Z(n2270));
Q_AN02 U2450 ( .A0(n2619), .A1(GFidata[381]), .Z(n2269));
Q_AN02 U2451 ( .A0(n2619), .A1(GFidata[382]), .Z(n2268));
Q_AN02 U2452 ( .A0(n2619), .A1(GFidata[383]), .Z(n2267));
Q_AN02 U2453 ( .A0(n2619), .A1(GFidata[384]), .Z(n2266));
Q_AN02 U2454 ( .A0(n2619), .A1(GFidata[385]), .Z(n2265));
Q_AN02 U2455 ( .A0(n2619), .A1(GFidata[386]), .Z(n2264));
Q_AN02 U2456 ( .A0(n2619), .A1(GFidata[387]), .Z(n2263));
Q_AN02 U2457 ( .A0(n2619), .A1(GFidata[388]), .Z(n2262));
Q_AN02 U2458 ( .A0(n2619), .A1(GFidata[389]), .Z(n2261));
Q_AN02 U2459 ( .A0(n2619), .A1(GFidata[390]), .Z(n2260));
Q_AN02 U2460 ( .A0(n2619), .A1(GFidata[391]), .Z(n2259));
Q_AN02 U2461 ( .A0(n2619), .A1(GFidata[392]), .Z(n2258));
Q_AN02 U2462 ( .A0(n2619), .A1(GFidata[393]), .Z(n2257));
Q_AN02 U2463 ( .A0(n2619), .A1(GFidata[394]), .Z(n2256));
Q_AN02 U2464 ( .A0(n2619), .A1(GFidata[395]), .Z(n2255));
Q_AN02 U2465 ( .A0(n2619), .A1(GFidata[396]), .Z(n2254));
Q_AN02 U2466 ( .A0(n2619), .A1(GFidata[397]), .Z(n2253));
Q_AN02 U2467 ( .A0(n2619), .A1(GFidata[398]), .Z(n2252));
Q_AN02 U2468 ( .A0(n2619), .A1(GFidata[399]), .Z(n2251));
Q_AN02 U2469 ( .A0(n2619), .A1(GFidata[400]), .Z(n2250));
Q_AN02 U2470 ( .A0(n2619), .A1(GFidata[401]), .Z(n2249));
Q_AN02 U2471 ( .A0(n2619), .A1(GFidata[402]), .Z(n2248));
Q_AN02 U2472 ( .A0(n2619), .A1(GFidata[403]), .Z(n2247));
Q_AN02 U2473 ( .A0(n2619), .A1(GFidata[404]), .Z(n2246));
Q_AN02 U2474 ( .A0(n2619), .A1(GFidata[405]), .Z(n2245));
Q_AN02 U2475 ( .A0(n2619), .A1(GFidata[406]), .Z(n2244));
Q_AN02 U2476 ( .A0(n2619), .A1(GFidata[407]), .Z(n2243));
Q_AN02 U2477 ( .A0(n2619), .A1(GFidata[408]), .Z(n2242));
Q_AN02 U2478 ( .A0(n2619), .A1(GFidata[409]), .Z(n2241));
Q_AN02 U2479 ( .A0(n2619), .A1(GFidata[410]), .Z(n2240));
Q_AN02 U2480 ( .A0(n2619), .A1(GFidata[411]), .Z(n2239));
Q_AN02 U2481 ( .A0(n2619), .A1(GFidata[412]), .Z(n2238));
Q_AN02 U2482 ( .A0(n2619), .A1(GFidata[413]), .Z(n2237));
Q_AN02 U2483 ( .A0(n2619), .A1(GFidata[414]), .Z(n2236));
Q_AN02 U2484 ( .A0(n2619), .A1(GFidata[415]), .Z(n2235));
Q_AN02 U2485 ( .A0(n2619), .A1(GFidata[416]), .Z(n2234));
Q_AN02 U2486 ( .A0(n2619), .A1(GFidata[417]), .Z(n2233));
Q_AN02 U2487 ( .A0(n2619), .A1(GFidata[418]), .Z(n2232));
Q_AN02 U2488 ( .A0(n2619), .A1(GFidata[419]), .Z(n2231));
Q_AN02 U2489 ( .A0(n2619), .A1(GFidata[420]), .Z(n2230));
Q_AN02 U2490 ( .A0(n2619), .A1(GFidata[421]), .Z(n2229));
Q_AN02 U2491 ( .A0(n2619), .A1(GFidata[422]), .Z(n2228));
Q_AN02 U2492 ( .A0(n2619), .A1(GFidata[423]), .Z(n2227));
Q_AN02 U2493 ( .A0(n2619), .A1(GFidata[424]), .Z(n2226));
Q_AN02 U2494 ( .A0(n2619), .A1(GFidata[425]), .Z(n2225));
Q_AN02 U2495 ( .A0(n2619), .A1(GFidata[426]), .Z(n2224));
Q_AN02 U2496 ( .A0(n2619), .A1(GFidata[427]), .Z(n2223));
Q_AN02 U2497 ( .A0(n2619), .A1(GFidata[428]), .Z(n2222));
Q_AN02 U2498 ( .A0(n2619), .A1(GFidata[429]), .Z(n2221));
Q_AN02 U2499 ( .A0(n2619), .A1(GFidata[430]), .Z(n2220));
Q_AN02 U2500 ( .A0(n2619), .A1(GFidata[431]), .Z(n2219));
Q_AN02 U2501 ( .A0(n2619), .A1(GFidata[432]), .Z(n2218));
Q_AN02 U2502 ( .A0(n2619), .A1(GFidata[433]), .Z(n2217));
Q_AN02 U2503 ( .A0(n2619), .A1(GFidata[434]), .Z(n2216));
Q_AN02 U2504 ( .A0(n2619), .A1(GFidata[435]), .Z(n2215));
Q_AN02 U2505 ( .A0(n2619), .A1(GFidata[436]), .Z(n2214));
Q_AN02 U2506 ( .A0(n2619), .A1(GFidata[437]), .Z(n2213));
Q_AN02 U2507 ( .A0(n2619), .A1(GFidata[438]), .Z(n2212));
Q_AN02 U2508 ( .A0(n2619), .A1(GFidata[439]), .Z(n2211));
Q_AN02 U2509 ( .A0(n2619), .A1(GFidata[440]), .Z(n2210));
Q_AN02 U2510 ( .A0(n2619), .A1(GFidata[441]), .Z(n2209));
Q_AN02 U2511 ( .A0(n2619), .A1(GFidata[442]), .Z(n2208));
Q_AN02 U2512 ( .A0(n2619), .A1(GFidata[443]), .Z(n2207));
Q_AN02 U2513 ( .A0(n2619), .A1(GFidata[444]), .Z(n2206));
Q_AN02 U2514 ( .A0(n2619), .A1(GFidata[445]), .Z(n2205));
Q_AN02 U2515 ( .A0(n2619), .A1(GFidata[446]), .Z(n2204));
Q_AN02 U2516 ( .A0(n2619), .A1(GFidata[447]), .Z(n2203));
Q_AN02 U2517 ( .A0(n2619), .A1(GFidata[448]), .Z(n2202));
Q_AN02 U2518 ( .A0(n2619), .A1(GFidata[449]), .Z(n2201));
Q_AN02 U2519 ( .A0(n2619), .A1(GFidata[450]), .Z(n2200));
Q_AN02 U2520 ( .A0(n2619), .A1(GFidata[451]), .Z(n2199));
Q_AN02 U2521 ( .A0(n2619), .A1(GFidata[452]), .Z(n2198));
Q_AN02 U2522 ( .A0(n2619), .A1(GFidata[453]), .Z(n2197));
Q_AN02 U2523 ( .A0(n2619), .A1(GFidata[454]), .Z(n2196));
Q_AN02 U2524 ( .A0(n2619), .A1(GFidata[455]), .Z(n2195));
Q_AN02 U2525 ( .A0(n2619), .A1(GFidata[456]), .Z(n2194));
Q_AN02 U2526 ( .A0(n2619), .A1(GFidata[457]), .Z(n2193));
Q_AN02 U2527 ( .A0(n2619), .A1(GFidata[458]), .Z(n2192));
Q_AN02 U2528 ( .A0(n2619), .A1(GFidata[459]), .Z(n2191));
Q_AN02 U2529 ( .A0(n2619), .A1(GFidata[460]), .Z(n2190));
Q_AN02 U2530 ( .A0(n2619), .A1(GFidata[461]), .Z(n2189));
Q_AN02 U2531 ( .A0(n2619), .A1(GFidata[462]), .Z(n2188));
Q_AN02 U2532 ( .A0(n2619), .A1(GFidata[463]), .Z(n2187));
Q_AN02 U2533 ( .A0(n2619), .A1(GFidata[464]), .Z(n2186));
Q_AN02 U2534 ( .A0(n2619), .A1(GFidata[465]), .Z(n2185));
Q_AN02 U2535 ( .A0(n2619), .A1(GFidata[466]), .Z(n2184));
Q_AN02 U2536 ( .A0(n2619), .A1(GFidata[467]), .Z(n2183));
Q_AN02 U2537 ( .A0(n2619), .A1(GFidata[468]), .Z(n2182));
Q_AN02 U2538 ( .A0(n2619), .A1(GFidata[469]), .Z(n2181));
Q_AN02 U2539 ( .A0(n2619), .A1(GFidata[470]), .Z(n2180));
Q_AN02 U2540 ( .A0(n2619), .A1(GFidata[471]), .Z(n2179));
Q_AN02 U2541 ( .A0(n2619), .A1(GFidata[472]), .Z(n2178));
Q_AN02 U2542 ( .A0(n2619), .A1(GFidata[473]), .Z(n2177));
Q_AN02 U2543 ( .A0(n2619), .A1(GFidata[474]), .Z(n2176));
Q_AN02 U2544 ( .A0(n2619), .A1(GFidata[475]), .Z(n2175));
Q_AN02 U2545 ( .A0(n2619), .A1(GFidata[476]), .Z(n2174));
Q_AN02 U2546 ( .A0(n2619), .A1(GFidata[477]), .Z(n2173));
Q_AN02 U2547 ( .A0(n2619), .A1(GFidata[478]), .Z(n2172));
Q_AN02 U2548 ( .A0(n2619), .A1(GFidata[479]), .Z(n2171));
Q_AN03 U2549 ( .A0(n2619), .A1(GFidata[480]), .A2(n786), .Z(n921));
Q_AN03 U2550 ( .A0(n2619), .A1(GFidata[481]), .A2(n786), .Z(n920));
Q_AN03 U2551 ( .A0(n2619), .A1(GFidata[482]), .A2(n786), .Z(n919));
Q_AN03 U2552 ( .A0(n2619), .A1(GFidata[483]), .A2(n786), .Z(n918));
Q_AN03 U2553 ( .A0(n2619), .A1(GFidata[484]), .A2(n786), .Z(n917));
Q_AN03 U2554 ( .A0(n2619), .A1(GFidata[485]), .A2(n786), .Z(n916));
Q_AN03 U2555 ( .A0(n2619), .A1(GFidata[486]), .A2(n786), .Z(n915));
Q_AN03 U2556 ( .A0(n2619), .A1(GFidata[487]), .A2(n786), .Z(n914));
Q_AN03 U2557 ( .A0(n2619), .A1(GFidata[488]), .A2(n786), .Z(n913));
Q_AN03 U2558 ( .A0(n2619), .A1(GFidata[489]), .A2(n786), .Z(n912));
Q_AN03 U2559 ( .A0(n2619), .A1(GFidata[490]), .A2(n786), .Z(n911));
Q_AN03 U2560 ( .A0(n2619), .A1(GFidata[491]), .A2(n786), .Z(n910));
Q_AN03 U2561 ( .A0(n2619), .A1(GFidata[492]), .A2(n786), .Z(n909));
Q_AN03 U2562 ( .A0(n2619), .A1(GFidata[493]), .A2(n786), .Z(n908));
Q_AN03 U2563 ( .A0(n2619), .A1(GFidata[494]), .A2(n786), .Z(n907));
Q_AN03 U2564 ( .A0(n2619), .A1(GFidata[495]), .A2(n786), .Z(n906));
Q_AN03 U2565 ( .A0(n2619), .A1(GFidata[496]), .A2(n786), .Z(n905));
Q_AN03 U2566 ( .A0(n2619), .A1(GFidata[497]), .A2(n786), .Z(n904));
Q_AN03 U2567 ( .A0(n2619), .A1(GFidata[498]), .A2(n786), .Z(n903));
Q_AN03 U2568 ( .A0(n2619), .A1(GFidata[499]), .A2(n786), .Z(n902));
Q_AN03 U2569 ( .A0(n2619), .A1(GFidata[500]), .A2(n786), .Z(n901));
Q_AN03 U2570 ( .A0(n2619), .A1(GFidata[501]), .A2(n786), .Z(n900));
Q_AN03 U2571 ( .A0(n2619), .A1(GFidata[502]), .A2(n786), .Z(n899));
Q_AN03 U2572 ( .A0(n2619), .A1(GFidata[503]), .A2(n786), .Z(n898));
Q_AN03 U2573 ( .A0(n2619), .A1(GFidata[504]), .A2(n786), .Z(n897));
Q_AN03 U2574 ( .A0(n2619), .A1(GFidata[505]), .A2(n786), .Z(n896));
Q_AN03 U2575 ( .A0(n2619), .A1(GFidata[506]), .A2(n786), .Z(n895));
Q_AN03 U2576 ( .A0(n2619), .A1(GFidata[507]), .A2(n786), .Z(n894));
Q_AN03 U2577 ( .A0(n2619), .A1(GFidata[508]), .A2(n786), .Z(n893));
Q_AN03 U2578 ( .A0(n2619), .A1(GFidata[509]), .A2(n786), .Z(n892));
Q_AN03 U2579 ( .A0(n2619), .A1(GFidata[510]), .A2(n786), .Z(n891));
Q_AN03 U2580 ( .A0(n2619), .A1(GFidata[511]), .A2(n786), .Z(n890));
Q_AD01HF U2581 ( .A0(n2160), .B0(n2161), .S(n2170), .CO(n2169));
Q_AD01HF U2582 ( .A0(n2169), .B0(n2159), .S(n2168), .CO(n2167));
Q_AD01HF U2583 ( .A0(n2167), .B0(n2158), .S(n2166), .CO(n2165));
Q_AD01HF U2584 ( .A0(n2165), .B0(n2157), .S(n2164), .CO(n2163));
Q_AN02 U2585 ( .A0(n787), .A1(GFlen[0]), .Z(n2161));
Q_AN02 U2586 ( .A0(n787), .A1(GFlen[1]), .Z(n2160));
Q_AN02 U2587 ( .A0(n787), .A1(GFlen[2]), .Z(n2159));
Q_AN02 U2588 ( .A0(n787), .A1(GFlen[3]), .Z(n2158));
Q_OR02 U2589 ( .A0(n783), .A1(GFlen[4]), .Z(n2157));
Q_AN02 U2590 ( .A0(n787), .A1(GFlen[5]), .Z(n2156));
Q_MX02 U2591 ( .S(n813), .A0(GFlen[0]), .A1(argLen[0]), .Z(n2155));
Q_MX02 U2592 ( .S(n813), .A0(GFlen[1]), .A1(argLen[1]), .Z(n2154));
Q_MX02 U2593 ( .S(n813), .A0(GFlen[2]), .A1(argLen[2]), .Z(n2153));
Q_MX02 U2594 ( .S(n813), .A0(GFlen[3]), .A1(argLen[3]), .Z(n2152));
Q_MX02 U2595 ( .S(n813), .A0(GFlen[4]), .A1(argLen[4]), .Z(n2151));
Q_MX02 U2596 ( .S(n813), .A0(GFlen[5]), .A1(argLen[5]), .Z(n2150));
Q_MX02 U2597 ( .S(n813), .A0(GFlen[6]), .A1(argLen[6]), .Z(n2149));
Q_MX02 U2598 ( .S(n813), .A0(GFlen[7]), .A1(argLen[7]), .Z(n2148));
Q_MX02 U2599 ( .S(n813), .A0(GFlen[8]), .A1(argLen[8]), .Z(n2147));
Q_MX02 U2600 ( .S(n813), .A0(GFlen[9]), .A1(argLen[9]), .Z(n2146));
Q_MX02 U2601 ( .S(n813), .A0(GFlen[10]), .A1(argLen[10]), .Z(n2145));
Q_MX02 U2602 ( .S(n813), .A0(GFlen[11]), .A1(argLen[11]), .Z(n2144));
Q_XNR2 U2603 ( .A0(wrtCnt[0]), .A1(n2155), .Z(n2143));
Q_OR02 U2604 ( .A0(wrtCnt[0]), .A1(n2155), .Z(n2142));
Q_AD01 U2605 ( .CI(n2142), .A0(wrtCnt[1]), .B0(n2154), .S(n2141), .CO(n2140));
Q_AD02 U2606 ( .CI(n2140), .A0(wrtCnt[2]), .A1(wrtCnt[3]), .B0(n2153), .B1(n2152), .S0(n2139), .S1(n2138), .CO(n2137));
Q_AD02 U2607 ( .CI(n2137), .A0(wrtCnt[4]), .A1(wrtCnt[5]), .B0(n2151), .B1(n2150), .S0(n2136), .S1(n2135), .CO(n2134));
Q_AD02 U2608 ( .CI(n2134), .A0(wrtCnt[6]), .A1(wrtCnt[7]), .B0(n2149), .B1(n2148), .S0(n2133), .S1(n2132), .CO(n2131));
Q_AD02 U2609 ( .CI(n2131), .A0(wrtCnt[8]), .A1(wrtCnt[9]), .B0(n2147), .B1(n2146), .S0(n2130), .S1(n2129), .CO(n2128));
Q_AD02 U2610 ( .CI(n2128), .A0(wrtCnt[10]), .A1(wrtCnt[11]), .B0(n2145), .B1(n2144), .S0(n2127), .S1(n2126), .CO(n2125));
Q_AD01HF U2611 ( .A0(wrtCnt[12]), .B0(n2125), .S(n2124), .CO(n2123));
Q_AD01HF U2612 ( .A0(wrtCnt[13]), .B0(n2123), .S(n2122), .CO(n2121));
Q_AD01HF U2613 ( .A0(wrtCnt[14]), .B0(n2121), .S(n2120), .CO(n2119));
Q_AD01HF U2614 ( .A0(wrtCnt[15]), .B0(n2119), .S(n2118), .CO(n2117));
Q_AD01HF U2615 ( .A0(wrtCnt[16]), .B0(n2117), .S(n2116), .CO(n2115));
Q_AD01HF U2616 ( .A0(wrtCnt[17]), .B0(n2115), .S(n2114), .CO(n2113));
Q_AD01HF U2617 ( .A0(wrtCnt[18]), .B0(n2113), .S(n2112), .CO(n2111));
Q_AD01HF U2618 ( .A0(wrtCnt[19]), .B0(n2111), .S(n2110), .CO(n2109));
Q_AD01HF U2619 ( .A0(wrtCnt[20]), .B0(n2109), .S(n2108), .CO(n2107));
Q_AD01HF U2620 ( .A0(wrtCnt[21]), .B0(n2107), .S(n2106), .CO(n2105));
Q_AD01HF U2621 ( .A0(wrtCnt[22]), .B0(n2105), .S(n2104), .CO(n2103));
Q_AD01HF U2622 ( .A0(wrtCnt[23]), .B0(n2103), .S(n2102), .CO(n2101));
Q_AD01HF U2623 ( .A0(wrtCnt[24]), .B0(n2101), .S(n2100), .CO(n2099));
Q_AD01HF U2624 ( .A0(wrtCnt[25]), .B0(n2099), .S(n2098), .CO(n2097));
Q_AD01HF U2625 ( .A0(wrtCnt[26]), .B0(n2097), .S(n2096), .CO(n2095));
Q_AD01HF U2626 ( .A0(wrtCnt[27]), .B0(n2095), .S(n2094), .CO(n2093));
Q_AD01HF U2627 ( .A0(wrtCnt[28]), .B0(n2093), .S(n2092), .CO(n2091));
Q_AD01HF U2628 ( .A0(wrtCnt[29]), .B0(n2091), .S(n2090), .CO(n2089));
Q_AD01HF U2629 ( .A0(wrtCnt[30]), .B0(n2089), .S(n2088), .CO(n2087));
Q_AD01HF U2630 ( .A0(wrtCnt[31]), .B0(n2087), .S(n2086), .CO(n2085));
Q_AD01HF U2631 ( .A0(wrtCnt[32]), .B0(n2085), .S(n2084), .CO(n2083));
Q_AD01HF U2632 ( .A0(wrtCnt[33]), .B0(n2083), .S(n2082), .CO(n2081));
Q_AD01HF U2633 ( .A0(wrtCnt[34]), .B0(n2081), .S(n2080), .CO(n2079));
Q_AD01HF U2634 ( .A0(wrtCnt[35]), .B0(n2079), .S(n2078), .CO(n2077));
Q_AD01HF U2635 ( .A0(wrtCnt[36]), .B0(n2077), .S(n2076), .CO(n2075));
Q_AD01HF U2636 ( .A0(wrtCnt[37]), .B0(n2075), .S(n2074), .CO(n2073));
Q_AD01HF U2637 ( .A0(wrtCnt[38]), .B0(n2073), .S(n2072), .CO(n2071));
Q_AD01HF U2638 ( .A0(wrtCnt[39]), .B0(n2071), .S(n2070), .CO(n2069));
Q_AD01HF U2639 ( .A0(wrtCnt[40]), .B0(n2069), .S(n2068), .CO(n2067));
Q_AD01HF U2640 ( .A0(wrtCnt[41]), .B0(n2067), .S(n2066), .CO(n2065));
Q_AD01HF U2641 ( .A0(wrtCnt[42]), .B0(n2065), .S(n2064), .CO(n2063));
Q_AD01HF U2642 ( .A0(wrtCnt[43]), .B0(n2063), .S(n2062), .CO(n2061));
Q_AD01HF U2643 ( .A0(wrtCnt[44]), .B0(n2061), .S(n2060), .CO(n2059));
Q_AD01HF U2644 ( .A0(wrtCnt[45]), .B0(n2059), .S(n2058), .CO(n2057));
Q_AD01HF U2645 ( .A0(wrtCnt[46]), .B0(n2057), .S(n2056), .CO(n2055));
Q_AD01HF U2646 ( .A0(wrtCnt[47]), .B0(n2055), .S(n2054), .CO(n2053));
Q_AD01HF U2647 ( .A0(wrtCnt[48]), .B0(n2053), .S(n2052), .CO(n2051));
Q_AD01HF U2648 ( .A0(wrtCnt[49]), .B0(n2051), .S(n2050), .CO(n2049));
Q_AD01HF U2649 ( .A0(wrtCnt[50]), .B0(n2049), .S(n2048), .CO(n2047));
Q_AD01HF U2650 ( .A0(wrtCnt[51]), .B0(n2047), .S(n2046), .CO(n2045));
Q_AD01HF U2651 ( .A0(wrtCnt[52]), .B0(n2045), .S(n2044), .CO(n2043));
Q_AD01HF U2652 ( .A0(wrtCnt[53]), .B0(n2043), .S(n2042), .CO(n2041));
Q_AD01HF U2653 ( .A0(wrtCnt[54]), .B0(n2041), .S(n2040), .CO(n2039));
Q_AD01HF U2654 ( .A0(wrtCnt[55]), .B0(n2039), .S(n2038), .CO(n2037));
Q_AD01HF U2655 ( .A0(wrtCnt[56]), .B0(n2037), .S(n2036), .CO(n2035));
Q_AD01HF U2656 ( .A0(wrtCnt[57]), .B0(n2035), .S(n2034), .CO(n2033));
Q_AD01HF U2657 ( .A0(wrtCnt[58]), .B0(n2033), .S(n2032), .CO(n2031));
Q_AD01HF U2658 ( .A0(wrtCnt[59]), .B0(n2031), .S(n2030), .CO(n2029));
Q_AD01HF U2659 ( .A0(wrtCnt[60]), .B0(n2029), .S(n2028), .CO(n2027));
Q_AD01HF U2660 ( .A0(wrtCnt[61]), .B0(n2027), .S(n2026), .CO(n2025));
Q_AD01HF U2661 ( .A0(wrtCnt[62]), .B0(n2025), .S(n2024), .CO(n2023));
Q_XOR2 U2662 ( .A0(wrtCnt[63]), .A1(n2023), .Z(n2022));
Q_NR02 U2663 ( .A0(n808), .A1(n2161), .Z(n2021));
Q_MX02 U2664 ( .S(n785), .A0(n2021), .A1(n2161), .Z(n2020));
Q_AN02 U2665 ( .A0(n786), .A1(n2170), .Z(n2019));
Q_MX02 U2666 ( .S(n785), .A0(n2019), .A1(n2160), .Z(n2018));
Q_AN02 U2667 ( .A0(n786), .A1(n2168), .Z(n2017));
Q_MX02 U2668 ( .S(n785), .A0(n2017), .A1(n2159), .Z(n2016));
Q_AN02 U2669 ( .A0(n786), .A1(n2166), .Z(n2015));
Q_MX02 U2670 ( .S(n785), .A0(n2015), .A1(n2158), .Z(n2014));
Q_AN02 U2671 ( .A0(n786), .A1(n2164), .Z(n2013));
Q_MX02 U2672 ( .S(n785), .A0(n2013), .A1(n2157), .Z(n2012));
Q_AN02 U2673 ( .A0(n786), .A1(n2162), .Z(n2011));
Q_MX02 U2674 ( .S(n785), .A0(n2011), .A1(n2156), .Z(n2010));
Q_AN02 U2675 ( .A0(n65), .A1(n2143), .Z(n2009));
Q_AN02 U2676 ( .A0(n65), .A1(n2141), .Z(n2008));
Q_AN02 U2677 ( .A0(n65), .A1(n2139), .Z(n2007));
Q_AN02 U2678 ( .A0(n65), .A1(n2138), .Z(n2006));
Q_AN02 U2679 ( .A0(n65), .A1(n2136), .Z(n2005));
Q_AN02 U2680 ( .A0(n65), .A1(n2135), .Z(n2004));
Q_AN02 U2681 ( .A0(n65), .A1(n2133), .Z(n2003));
Q_AN02 U2682 ( .A0(n65), .A1(n2132), .Z(n2002));
Q_AN02 U2683 ( .A0(n65), .A1(n2130), .Z(n2001));
Q_AN02 U2684 ( .A0(n65), .A1(n2129), .Z(n2000));
Q_AN02 U2685 ( .A0(n65), .A1(n2127), .Z(n1999));
Q_AN02 U2686 ( .A0(n65), .A1(n2126), .Z(n1998));
Q_AN02 U2687 ( .A0(n65), .A1(n2124), .Z(n1997));
Q_AN02 U2688 ( .A0(n65), .A1(n2122), .Z(n1996));
Q_AN02 U2689 ( .A0(n65), .A1(n2120), .Z(n1995));
Q_AN02 U2690 ( .A0(n65), .A1(n2118), .Z(n1994));
Q_AN02 U2691 ( .A0(n65), .A1(n2116), .Z(n1993));
Q_AN02 U2692 ( .A0(n65), .A1(n2114), .Z(n1992));
Q_AN02 U2693 ( .A0(n65), .A1(n2112), .Z(n1991));
Q_AN02 U2694 ( .A0(n65), .A1(n2110), .Z(n1990));
Q_AN02 U2695 ( .A0(n65), .A1(n2108), .Z(n1989));
Q_AN02 U2696 ( .A0(n65), .A1(n2106), .Z(n1988));
Q_AN02 U2697 ( .A0(n65), .A1(n2104), .Z(n1987));
Q_AN02 U2698 ( .A0(n65), .A1(n2102), .Z(n1986));
Q_AN02 U2699 ( .A0(n65), .A1(n2100), .Z(n1985));
Q_AN02 U2700 ( .A0(n65), .A1(n2098), .Z(n1984));
Q_AN02 U2701 ( .A0(n65), .A1(n2096), .Z(n1983));
Q_AN02 U2702 ( .A0(n65), .A1(n2094), .Z(n1982));
Q_AN02 U2703 ( .A0(n65), .A1(n2092), .Z(n1981));
Q_AN02 U2704 ( .A0(n65), .A1(n2090), .Z(n1980));
Q_AN02 U2705 ( .A0(n65), .A1(n2088), .Z(n1979));
Q_AN02 U2706 ( .A0(n65), .A1(n2086), .Z(n1978));
Q_AN02 U2707 ( .A0(n65), .A1(n2084), .Z(n1977));
Q_AN02 U2708 ( .A0(n65), .A1(n2082), .Z(n1976));
Q_AN02 U2709 ( .A0(n65), .A1(n2080), .Z(n1975));
Q_AN02 U2710 ( .A0(n65), .A1(n2078), .Z(n1974));
Q_AN02 U2711 ( .A0(n65), .A1(n2076), .Z(n1973));
Q_AN02 U2712 ( .A0(n65), .A1(n2074), .Z(n1972));
Q_AN02 U2713 ( .A0(n65), .A1(n2072), .Z(n1971));
Q_AN02 U2714 ( .A0(n65), .A1(n2070), .Z(n1970));
Q_AN02 U2715 ( .A0(n65), .A1(n2068), .Z(n1969));
Q_AN02 U2716 ( .A0(n65), .A1(n2066), .Z(n1968));
Q_AN02 U2717 ( .A0(n65), .A1(n2064), .Z(n1967));
Q_AN02 U2718 ( .A0(n65), .A1(n2062), .Z(n1966));
Q_AN02 U2719 ( .A0(n65), .A1(n2060), .Z(n1965));
Q_AN02 U2720 ( .A0(n65), .A1(n2058), .Z(n1964));
Q_AN02 U2721 ( .A0(n65), .A1(n2056), .Z(n1963));
Q_AN02 U2722 ( .A0(n65), .A1(n2054), .Z(n1962));
Q_AN02 U2723 ( .A0(n65), .A1(n2052), .Z(n1961));
Q_AN02 U2724 ( .A0(n65), .A1(n2050), .Z(n1960));
Q_AN02 U2725 ( .A0(n65), .A1(n2048), .Z(n1959));
Q_AN02 U2726 ( .A0(n65), .A1(n2046), .Z(n1958));
Q_AN02 U2727 ( .A0(n65), .A1(n2044), .Z(n1957));
Q_AN02 U2728 ( .A0(n65), .A1(n2042), .Z(n1956));
Q_AN02 U2729 ( .A0(n65), .A1(n2040), .Z(n1955));
Q_AN02 U2730 ( .A0(n65), .A1(n2038), .Z(n1954));
Q_AN02 U2731 ( .A0(n65), .A1(n2036), .Z(n1953));
Q_AN02 U2732 ( .A0(n65), .A1(n2034), .Z(n1952));
Q_AN02 U2733 ( .A0(n65), .A1(n2032), .Z(n1951));
Q_AN02 U2734 ( .A0(n65), .A1(n2030), .Z(n1950));
Q_AN02 U2735 ( .A0(n65), .A1(n2028), .Z(n1949));
Q_AN02 U2736 ( .A0(n65), .A1(n2026), .Z(n1948));
Q_AN02 U2737 ( .A0(n65), .A1(n2024), .Z(n1947));
Q_AN02 U2738 ( .A0(n65), .A1(n2022), .Z(n1946));
Q_AN02 U2739 ( .A0(n785), .A1(GFidata[0]), .Z(n1945));
Q_MX03 U2740 ( .S0(n788), .S1(n808), .A0(GFcbid[0]), .A1(timeStampPkt[0]), .A2(n1945), .Z(n1944));
Q_AN02 U2741 ( .A0(n785), .A1(GFidata[1]), .Z(n1943));
Q_MX03 U2742 ( .S0(n788), .S1(n808), .A0(GFcbid[1]), .A1(timeStampPkt[1]), .A2(n1943), .Z(n1942));
Q_AN02 U2743 ( .A0(n785), .A1(GFidata[2]), .Z(n1941));
Q_MX03 U2744 ( .S0(n788), .S1(n808), .A0(GFcbid[2]), .A1(timeStampPkt[2]), .A2(n1941), .Z(n1940));
Q_AN02 U2745 ( .A0(n785), .A1(GFidata[3]), .Z(n1939));
Q_MX03 U2746 ( .S0(n788), .S1(n808), .A0(GFcbid[3]), .A1(timeStampPkt[3]), .A2(n1939), .Z(n1938));
Q_AN02 U2747 ( .A0(n785), .A1(GFidata[4]), .Z(n1937));
Q_MX03 U2748 ( .S0(n788), .S1(n808), .A0(GFcbid[4]), .A1(timeStampPkt[4]), .A2(n1937), .Z(n1936));
Q_AN02 U2749 ( .A0(n785), .A1(GFidata[5]), .Z(n1935));
Q_MX03 U2750 ( .S0(n788), .S1(n808), .A0(GFcbid[5]), .A1(timeStampPkt[5]), .A2(n1935), .Z(n1934));
Q_AN02 U2751 ( .A0(n785), .A1(GFidata[6]), .Z(n1933));
Q_MX03 U2752 ( .S0(n788), .S1(n808), .A0(GFcbid[6]), .A1(timeStampPkt[6]), .A2(n1933), .Z(n1932));
Q_AN02 U2753 ( .A0(n785), .A1(GFidata[7]), .Z(n1931));
Q_MX03 U2754 ( .S0(n788), .S1(n808), .A0(GFcbid[7]), .A1(timeStampPkt[7]), .A2(n1931), .Z(n1930));
Q_AN02 U2755 ( .A0(n785), .A1(GFidata[8]), .Z(n1929));
Q_MX03 U2756 ( .S0(n788), .S1(n808), .A0(GFcbid[8]), .A1(timeStampPkt[8]), .A2(n1929), .Z(n1928));
Q_AN02 U2757 ( .A0(n785), .A1(GFidata[9]), .Z(n1927));
Q_MX03 U2758 ( .S0(n788), .S1(n808), .A0(GFcbid[9]), .A1(timeStampPkt[9]), .A2(n1927), .Z(n1926));
Q_AN02 U2759 ( .A0(n785), .A1(GFidata[10]), .Z(n1925));
Q_MX03 U2760 ( .S0(n788), .S1(n808), .A0(GFcbid[10]), .A1(timeStampPkt[10]), .A2(n1925), .Z(n1924));
Q_AN02 U2761 ( .A0(n785), .A1(GFidata[11]), .Z(n1923));
Q_MX03 U2762 ( .S0(n788), .S1(n808), .A0(GFcbid[11]), .A1(timeStampPkt[11]), .A2(n1923), .Z(n1922));
Q_AN02 U2763 ( .A0(n785), .A1(GFidata[12]), .Z(n1921));
Q_MX03 U2764 ( .S0(n788), .S1(n808), .A0(GFcbid[12]), .A1(timeStampPkt[12]), .A2(n1921), .Z(n1920));
Q_AN02 U2765 ( .A0(n785), .A1(GFidata[13]), .Z(n1919));
Q_MX03 U2766 ( .S0(n788), .S1(n808), .A0(GFcbid[13]), .A1(timeStampPkt[13]), .A2(n1919), .Z(n1918));
Q_AN02 U2767 ( .A0(n785), .A1(GFidata[14]), .Z(n1917));
Q_MX03 U2768 ( .S0(n788), .S1(n808), .A0(GFcbid[14]), .A1(timeStampPkt[14]), .A2(n1917), .Z(n1916));
Q_AN02 U2769 ( .A0(n785), .A1(GFidata[15]), .Z(n1915));
Q_MX03 U2770 ( .S0(n788), .S1(n808), .A0(GFcbid[15]), .A1(timeStampPkt[15]), .A2(n1915), .Z(n1914));
Q_AN02 U2771 ( .A0(n785), .A1(GFidata[16]), .Z(n1913));
Q_MX03 U2772 ( .S0(n788), .S1(n808), .A0(GFcbid[16]), .A1(timeStampPkt[16]), .A2(n1913), .Z(n1912));
Q_AN02 U2773 ( .A0(n785), .A1(GFidata[17]), .Z(n1911));
Q_MX03 U2774 ( .S0(n788), .S1(n808), .A0(GFcbid[17]), .A1(timeStampPkt[17]), .A2(n1911), .Z(n1910));
Q_AN02 U2775 ( .A0(n785), .A1(GFidata[18]), .Z(n1909));
Q_MX03 U2776 ( .S0(n788), .S1(n808), .A0(GFcbid[18]), .A1(timeStampPkt[18]), .A2(n1909), .Z(n1908));
Q_AN02 U2777 ( .A0(n785), .A1(GFidata[19]), .Z(n1907));
Q_MX03 U2778 ( .S0(n788), .S1(n808), .A0(GFcbid[19]), .A1(timeStampPkt[19]), .A2(n1907), .Z(n1906));
Q_AN02 U2779 ( .A0(n785), .A1(GFidata[20]), .Z(n1905));
Q_MX03 U2780 ( .S0(n788), .S1(n808), .A0(GFlen[0]), .A1(timeStampPkt[20]), .A2(n1905), .Z(n1904));
Q_AN02 U2781 ( .A0(n785), .A1(GFidata[21]), .Z(n1903));
Q_MX03 U2782 ( .S0(n788), .S1(n808), .A0(GFlen[1]), .A1(timeStampPkt[21]), .A2(n1903), .Z(n1902));
Q_AN02 U2783 ( .A0(n785), .A1(GFidata[22]), .Z(n1901));
Q_MX03 U2784 ( .S0(n788), .S1(n808), .A0(GFlen[2]), .A1(timeStampPkt[22]), .A2(n1901), .Z(n1900));
Q_AN02 U2785 ( .A0(n785), .A1(GFidata[23]), .Z(n1899));
Q_MX03 U2786 ( .S0(n788), .S1(n808), .A0(GFlen[3]), .A1(timeStampPkt[23]), .A2(n1899), .Z(n1898));
Q_AN02 U2787 ( .A0(n785), .A1(GFidata[24]), .Z(n1897));
Q_MX03 U2788 ( .S0(n788), .S1(n808), .A0(GFlen[4]), .A1(timeStampPkt[24]), .A2(n1897), .Z(n1896));
Q_AN02 U2789 ( .A0(n785), .A1(GFidata[25]), .Z(n1895));
Q_MX03 U2790 ( .S0(n788), .S1(n808), .A0(GFlen[5]), .A1(timeStampPkt[25]), .A2(n1895), .Z(n1894));
Q_AN02 U2791 ( .A0(n785), .A1(GFidata[26]), .Z(n1893));
Q_MX03 U2792 ( .S0(n788), .S1(n808), .A0(GFlen[6]), .A1(timeStampPkt[26]), .A2(n1893), .Z(n1892));
Q_AN02 U2793 ( .A0(n785), .A1(GFidata[27]), .Z(n1891));
Q_MX03 U2794 ( .S0(n788), .S1(n808), .A0(GFlen[7]), .A1(timeStampPkt[27]), .A2(n1891), .Z(n1890));
Q_AN02 U2795 ( .A0(n785), .A1(GFidata[28]), .Z(n1889));
Q_MX03 U2796 ( .S0(n788), .S1(n808), .A0(GFlen[8]), .A1(timeStampPkt[28]), .A2(n1889), .Z(n1888));
Q_AN02 U2797 ( .A0(n785), .A1(GFidata[29]), .Z(n1887));
Q_MX03 U2798 ( .S0(n788), .S1(n808), .A0(GFlen[9]), .A1(timeStampPkt[29]), .A2(n1887), .Z(n1886));
Q_AN02 U2799 ( .A0(n785), .A1(GFidata[30]), .Z(n1885));
Q_MX03 U2800 ( .S0(n788), .S1(n808), .A0(GFlen[10]), .A1(timeStampPkt[30]), .A2(n1885), .Z(n1884));
Q_AN02 U2801 ( .A0(n785), .A1(GFidata[31]), .Z(n1883));
Q_MX02 U2802 ( .S(n808), .A0(n2620), .A1(n1883), .Z(n1882));
Q_AN02 U2803 ( .A0(n785), .A1(GFidata[32]), .Z(n1881));
Q_MX03 U2804 ( .S0(n788), .S1(n808), .A0(GFidata[0]), .A1(timeStampPkt[32]), .A2(n1881), .Z(n1880));
Q_AN02 U2805 ( .A0(n785), .A1(GFidata[33]), .Z(n1879));
Q_MX03 U2806 ( .S0(n788), .S1(n808), .A0(GFidata[1]), .A1(timeStampPkt[33]), .A2(n1879), .Z(n1878));
Q_AN02 U2807 ( .A0(n785), .A1(GFidata[34]), .Z(n1877));
Q_MX03 U2808 ( .S0(n788), .S1(n808), .A0(GFidata[2]), .A1(timeStampPkt[34]), .A2(n1877), .Z(n1876));
Q_AN02 U2809 ( .A0(n785), .A1(GFidata[35]), .Z(n1875));
Q_MX03 U2810 ( .S0(n788), .S1(n808), .A0(GFidata[3]), .A1(timeStampPkt[35]), .A2(n1875), .Z(n1874));
Q_AN02 U2811 ( .A0(n785), .A1(GFidata[36]), .Z(n1873));
Q_MX03 U2812 ( .S0(n788), .S1(n808), .A0(GFidata[4]), .A1(timeStampPkt[36]), .A2(n1873), .Z(n1872));
Q_AN02 U2813 ( .A0(n785), .A1(GFidata[37]), .Z(n1871));
Q_MX03 U2814 ( .S0(n788), .S1(n808), .A0(GFidata[5]), .A1(timeStampPkt[37]), .A2(n1871), .Z(n1870));
Q_AN02 U2815 ( .A0(n785), .A1(GFidata[38]), .Z(n1869));
Q_MX03 U2816 ( .S0(n788), .S1(n808), .A0(GFidata[6]), .A1(timeStampPkt[38]), .A2(n1869), .Z(n1868));
Q_AN02 U2817 ( .A0(n785), .A1(GFidata[39]), .Z(n1867));
Q_MX03 U2818 ( .S0(n788), .S1(n808), .A0(GFidata[7]), .A1(timeStampPkt[39]), .A2(n1867), .Z(n1866));
Q_AN02 U2819 ( .A0(n785), .A1(GFidata[40]), .Z(n1865));
Q_MX03 U2820 ( .S0(n788), .S1(n808), .A0(GFidata[8]), .A1(timeStampPkt[40]), .A2(n1865), .Z(n1864));
Q_AN02 U2821 ( .A0(n785), .A1(GFidata[41]), .Z(n1863));
Q_MX03 U2822 ( .S0(n788), .S1(n808), .A0(GFidata[9]), .A1(timeStampPkt[41]), .A2(n1863), .Z(n1862));
Q_AN02 U2823 ( .A0(n785), .A1(GFidata[42]), .Z(n1861));
Q_MX03 U2824 ( .S0(n788), .S1(n808), .A0(GFidata[10]), .A1(timeStampPkt[42]), .A2(n1861), .Z(n1860));
Q_AN02 U2825 ( .A0(n785), .A1(GFidata[43]), .Z(n1859));
Q_MX03 U2826 ( .S0(n788), .S1(n808), .A0(GFidata[11]), .A1(timeStampPkt[43]), .A2(n1859), .Z(n1858));
Q_AN02 U2827 ( .A0(n785), .A1(GFidata[44]), .Z(n1857));
Q_MX03 U2828 ( .S0(n788), .S1(n808), .A0(GFidata[12]), .A1(timeStampPkt[44]), .A2(n1857), .Z(n1856));
Q_AN02 U2829 ( .A0(n785), .A1(GFidata[45]), .Z(n1855));
Q_MX03 U2830 ( .S0(n788), .S1(n808), .A0(GFidata[13]), .A1(timeStampPkt[45]), .A2(n1855), .Z(n1854));
Q_AN02 U2831 ( .A0(n785), .A1(GFidata[46]), .Z(n1853));
Q_MX03 U2832 ( .S0(n788), .S1(n808), .A0(GFidata[14]), .A1(timeStampPkt[46]), .A2(n1853), .Z(n1852));
Q_AN02 U2833 ( .A0(n785), .A1(GFidata[47]), .Z(n1851));
Q_MX03 U2834 ( .S0(n788), .S1(n808), .A0(GFidata[15]), .A1(timeStampPkt[47]), .A2(n1851), .Z(n1850));
Q_AN02 U2835 ( .A0(n785), .A1(GFidata[48]), .Z(n1849));
Q_MX03 U2836 ( .S0(n788), .S1(n808), .A0(GFidata[16]), .A1(timeStampPkt[48]), .A2(n1849), .Z(n1848));
Q_AN02 U2837 ( .A0(n785), .A1(GFidata[49]), .Z(n1847));
Q_MX03 U2838 ( .S0(n788), .S1(n808), .A0(GFidata[17]), .A1(timeStampPkt[49]), .A2(n1847), .Z(n1846));
Q_AN02 U2839 ( .A0(n785), .A1(GFidata[50]), .Z(n1845));
Q_MX03 U2840 ( .S0(n788), .S1(n808), .A0(GFidata[18]), .A1(timeStampPkt[50]), .A2(n1845), .Z(n1844));
Q_AN02 U2841 ( .A0(n785), .A1(GFidata[51]), .Z(n1843));
Q_MX03 U2842 ( .S0(n788), .S1(n808), .A0(GFidata[19]), .A1(timeStampPkt[51]), .A2(n1843), .Z(n1842));
Q_AN02 U2843 ( .A0(n785), .A1(GFidata[52]), .Z(n1841));
Q_MX03 U2844 ( .S0(n788), .S1(n808), .A0(GFidata[20]), .A1(timeStampPkt[52]), .A2(n1841), .Z(n1840));
Q_AN02 U2845 ( .A0(n785), .A1(GFidata[53]), .Z(n1839));
Q_MX03 U2846 ( .S0(n788), .S1(n808), .A0(GFidata[21]), .A1(timeStampPkt[53]), .A2(n1839), .Z(n1838));
Q_AN02 U2847 ( .A0(n785), .A1(GFidata[54]), .Z(n1837));
Q_MX03 U2848 ( .S0(n788), .S1(n808), .A0(GFidata[22]), .A1(timeStampPkt[54]), .A2(n1837), .Z(n1836));
Q_AN02 U2849 ( .A0(n785), .A1(GFidata[55]), .Z(n1835));
Q_MX03 U2850 ( .S0(n788), .S1(n808), .A0(GFidata[23]), .A1(timeStampPkt[55]), .A2(n1835), .Z(n1834));
Q_AN02 U2851 ( .A0(n785), .A1(GFidata[56]), .Z(n1833));
Q_MX03 U2852 ( .S0(n788), .S1(n808), .A0(GFidata[24]), .A1(timeStampPkt[56]), .A2(n1833), .Z(n1832));
Q_AN02 U2853 ( .A0(n785), .A1(GFidata[57]), .Z(n1831));
Q_MX03 U2854 ( .S0(n788), .S1(n808), .A0(GFidata[25]), .A1(timeStampPkt[57]), .A2(n1831), .Z(n1830));
Q_AN02 U2855 ( .A0(n785), .A1(GFidata[58]), .Z(n1829));
Q_MX03 U2856 ( .S0(n788), .S1(n808), .A0(GFidata[26]), .A1(timeStampPkt[58]), .A2(n1829), .Z(n1828));
Q_AN02 U2857 ( .A0(n785), .A1(GFidata[59]), .Z(n1827));
Q_MX03 U2858 ( .S0(n788), .S1(n808), .A0(GFidata[27]), .A1(timeStampPkt[59]), .A2(n1827), .Z(n1826));
Q_AN02 U2859 ( .A0(n785), .A1(GFidata[60]), .Z(n1825));
Q_MX03 U2860 ( .S0(n788), .S1(n808), .A0(GFidata[28]), .A1(timeStampPkt[60]), .A2(n1825), .Z(n1824));
Q_AN02 U2861 ( .A0(n785), .A1(GFidata[61]), .Z(n1823));
Q_MX03 U2862 ( .S0(n788), .S1(n808), .A0(GFidata[29]), .A1(timeStampPkt[61]), .A2(n1823), .Z(n1822));
Q_AN02 U2863 ( .A0(n785), .A1(GFidata[62]), .Z(n1821));
Q_MX03 U2864 ( .S0(n788), .S1(n808), .A0(GFidata[30]), .A1(timeStampPkt[62]), .A2(n1821), .Z(n1820));
Q_AN02 U2865 ( .A0(n785), .A1(GFidata[63]), .Z(n1819));
Q_MX03 U2866 ( .S0(n788), .S1(n808), .A0(GFidata[31]), .A1(timeStampPkt[63]), .A2(n1819), .Z(n1818));
Q_AN02 U2867 ( .A0(n785), .A1(GFidata[64]), .Z(n1817));
Q_MX02 U2868 ( .S(n808), .A0(n2618), .A1(n1817), .Z(n1816));
Q_AN02 U2869 ( .A0(n785), .A1(GFidata[65]), .Z(n1815));
Q_MX02 U2870 ( .S(n808), .A0(n2617), .A1(n1815), .Z(n1814));
Q_AN02 U2871 ( .A0(n785), .A1(GFidata[66]), .Z(n1813));
Q_MX02 U2872 ( .S(n808), .A0(n2616), .A1(n1813), .Z(n1812));
Q_AN02 U2873 ( .A0(n785), .A1(GFidata[67]), .Z(n1811));
Q_MX02 U2874 ( .S(n808), .A0(n2615), .A1(n1811), .Z(n1810));
Q_AN02 U2875 ( .A0(n785), .A1(GFidata[68]), .Z(n1809));
Q_MX02 U2876 ( .S(n808), .A0(n2614), .A1(n1809), .Z(n1808));
Q_AN02 U2877 ( .A0(n785), .A1(GFidata[69]), .Z(n1807));
Q_MX02 U2878 ( .S(n808), .A0(n2613), .A1(n1807), .Z(n1806));
Q_AN02 U2879 ( .A0(n785), .A1(GFidata[70]), .Z(n1805));
Q_MX02 U2880 ( .S(n808), .A0(n2612), .A1(n1805), .Z(n1804));
Q_AN02 U2881 ( .A0(n785), .A1(GFidata[71]), .Z(n1803));
Q_MX02 U2882 ( .S(n808), .A0(n2611), .A1(n1803), .Z(n1802));
Q_AN02 U2883 ( .A0(n785), .A1(GFidata[72]), .Z(n1801));
Q_MX02 U2884 ( .S(n808), .A0(n2610), .A1(n1801), .Z(n1800));
Q_AN02 U2885 ( .A0(n785), .A1(GFidata[73]), .Z(n1799));
Q_MX02 U2886 ( .S(n808), .A0(n2609), .A1(n1799), .Z(n1798));
Q_AN02 U2887 ( .A0(n785), .A1(GFidata[74]), .Z(n1797));
Q_MX02 U2888 ( .S(n808), .A0(n2608), .A1(n1797), .Z(n1796));
Q_AN02 U2889 ( .A0(n785), .A1(GFidata[75]), .Z(n1795));
Q_MX02 U2890 ( .S(n808), .A0(n2607), .A1(n1795), .Z(n1794));
Q_AN02 U2891 ( .A0(n785), .A1(GFidata[76]), .Z(n1793));
Q_MX02 U2892 ( .S(n808), .A0(n2606), .A1(n1793), .Z(n1792));
Q_AN02 U2893 ( .A0(n785), .A1(GFidata[77]), .Z(n1791));
Q_MX02 U2894 ( .S(n808), .A0(n2605), .A1(n1791), .Z(n1790));
Q_AN02 U2895 ( .A0(n785), .A1(GFidata[78]), .Z(n1789));
Q_MX02 U2896 ( .S(n808), .A0(n2604), .A1(n1789), .Z(n1788));
Q_AN02 U2897 ( .A0(n785), .A1(GFidata[79]), .Z(n1787));
Q_MX02 U2898 ( .S(n808), .A0(n2603), .A1(n1787), .Z(n1786));
Q_AN02 U2899 ( .A0(n785), .A1(GFidata[80]), .Z(n1785));
Q_MX02 U2900 ( .S(n808), .A0(n2602), .A1(n1785), .Z(n1784));
Q_AN02 U2901 ( .A0(n785), .A1(GFidata[81]), .Z(n1783));
Q_MX02 U2902 ( .S(n808), .A0(n2601), .A1(n1783), .Z(n1782));
Q_AN02 U2903 ( .A0(n785), .A1(GFidata[82]), .Z(n1781));
Q_MX02 U2904 ( .S(n808), .A0(n2600), .A1(n1781), .Z(n1780));
Q_AN02 U2905 ( .A0(n785), .A1(GFidata[83]), .Z(n1779));
Q_MX02 U2906 ( .S(n808), .A0(n2599), .A1(n1779), .Z(n1778));
Q_AN02 U2907 ( .A0(n785), .A1(GFidata[84]), .Z(n1777));
Q_MX02 U2908 ( .S(n808), .A0(n2598), .A1(n1777), .Z(n1776));
Q_AN02 U2909 ( .A0(n785), .A1(GFidata[85]), .Z(n1775));
Q_MX02 U2910 ( .S(n808), .A0(n2597), .A1(n1775), .Z(n1774));
Q_AN02 U2911 ( .A0(n785), .A1(GFidata[86]), .Z(n1773));
Q_MX02 U2912 ( .S(n808), .A0(n2596), .A1(n1773), .Z(n1772));
Q_AN02 U2913 ( .A0(n785), .A1(GFidata[87]), .Z(n1771));
Q_MX02 U2914 ( .S(n808), .A0(n2595), .A1(n1771), .Z(n1770));
Q_AN02 U2915 ( .A0(n785), .A1(GFidata[88]), .Z(n1769));
Q_MX02 U2916 ( .S(n808), .A0(n2594), .A1(n1769), .Z(n1768));
Q_AN02 U2917 ( .A0(n785), .A1(GFidata[89]), .Z(n1767));
Q_MX02 U2918 ( .S(n808), .A0(n2593), .A1(n1767), .Z(n1766));
Q_AN02 U2919 ( .A0(n785), .A1(GFidata[90]), .Z(n1765));
Q_MX02 U2920 ( .S(n808), .A0(n2592), .A1(n1765), .Z(n1764));
Q_AN02 U2921 ( .A0(n785), .A1(GFidata[91]), .Z(n1763));
Q_MX02 U2922 ( .S(n808), .A0(n2591), .A1(n1763), .Z(n1762));
Q_AN02 U2923 ( .A0(n785), .A1(GFidata[92]), .Z(n1761));
Q_MX02 U2924 ( .S(n808), .A0(n2590), .A1(n1761), .Z(n1760));
Q_AN02 U2925 ( .A0(n785), .A1(GFidata[93]), .Z(n1759));
Q_MX02 U2926 ( .S(n808), .A0(n2589), .A1(n1759), .Z(n1758));
Q_AN02 U2927 ( .A0(n785), .A1(GFidata[94]), .Z(n1757));
Q_MX02 U2928 ( .S(n808), .A0(n2588), .A1(n1757), .Z(n1756));
Q_AN02 U2929 ( .A0(n785), .A1(GFidata[95]), .Z(n1755));
Q_MX02 U2930 ( .S(n808), .A0(n2587), .A1(n1755), .Z(n1754));
Q_AN02 U2931 ( .A0(n785), .A1(GFidata[96]), .Z(n1753));
Q_MX02 U2932 ( .S(n808), .A0(n2586), .A1(n1753), .Z(n1752));
Q_AN02 U2933 ( .A0(n785), .A1(GFidata[97]), .Z(n1751));
Q_MX02 U2934 ( .S(n808), .A0(n2585), .A1(n1751), .Z(n1750));
Q_AN02 U2935 ( .A0(n785), .A1(GFidata[98]), .Z(n1749));
Q_MX02 U2936 ( .S(n808), .A0(n2584), .A1(n1749), .Z(n1748));
Q_AN02 U2937 ( .A0(n785), .A1(GFidata[99]), .Z(n1747));
Q_MX02 U2938 ( .S(n808), .A0(n2583), .A1(n1747), .Z(n1746));
Q_AN02 U2939 ( .A0(n785), .A1(GFidata[100]), .Z(n1745));
Q_MX02 U2940 ( .S(n808), .A0(n2582), .A1(n1745), .Z(n1744));
Q_AN02 U2941 ( .A0(n785), .A1(GFidata[101]), .Z(n1743));
Q_MX02 U2942 ( .S(n808), .A0(n2581), .A1(n1743), .Z(n1742));
Q_AN02 U2943 ( .A0(n785), .A1(GFidata[102]), .Z(n1741));
Q_MX02 U2944 ( .S(n808), .A0(n2580), .A1(n1741), .Z(n1740));
Q_AN02 U2945 ( .A0(n785), .A1(GFidata[103]), .Z(n1739));
Q_MX02 U2946 ( .S(n808), .A0(n2579), .A1(n1739), .Z(n1738));
Q_AN02 U2947 ( .A0(n785), .A1(GFidata[104]), .Z(n1737));
Q_MX02 U2948 ( .S(n808), .A0(n2578), .A1(n1737), .Z(n1736));
Q_AN02 U2949 ( .A0(n785), .A1(GFidata[105]), .Z(n1735));
Q_MX02 U2950 ( .S(n808), .A0(n2577), .A1(n1735), .Z(n1734));
Q_AN02 U2951 ( .A0(n785), .A1(GFidata[106]), .Z(n1733));
Q_MX02 U2952 ( .S(n808), .A0(n2576), .A1(n1733), .Z(n1732));
Q_AN02 U2953 ( .A0(n785), .A1(GFidata[107]), .Z(n1731));
Q_MX02 U2954 ( .S(n808), .A0(n2575), .A1(n1731), .Z(n1730));
Q_AN02 U2955 ( .A0(n785), .A1(GFidata[108]), .Z(n1729));
Q_MX02 U2956 ( .S(n808), .A0(n2574), .A1(n1729), .Z(n1728));
Q_AN02 U2957 ( .A0(n785), .A1(GFidata[109]), .Z(n1727));
Q_MX02 U2958 ( .S(n808), .A0(n2573), .A1(n1727), .Z(n1726));
Q_AN02 U2959 ( .A0(n785), .A1(GFidata[110]), .Z(n1725));
Q_MX02 U2960 ( .S(n808), .A0(n2572), .A1(n1725), .Z(n1724));
Q_AN02 U2961 ( .A0(n785), .A1(GFidata[111]), .Z(n1723));
Q_MX02 U2962 ( .S(n808), .A0(n2571), .A1(n1723), .Z(n1722));
Q_AN02 U2963 ( .A0(n785), .A1(GFidata[112]), .Z(n1721));
Q_MX02 U2964 ( .S(n808), .A0(n2570), .A1(n1721), .Z(n1720));
Q_AN02 U2965 ( .A0(n785), .A1(GFidata[113]), .Z(n1719));
Q_MX02 U2966 ( .S(n808), .A0(n2569), .A1(n1719), .Z(n1718));
Q_AN02 U2967 ( .A0(n785), .A1(GFidata[114]), .Z(n1717));
Q_MX02 U2968 ( .S(n808), .A0(n2568), .A1(n1717), .Z(n1716));
Q_AN02 U2969 ( .A0(n785), .A1(GFidata[115]), .Z(n1715));
Q_MX02 U2970 ( .S(n808), .A0(n2567), .A1(n1715), .Z(n1714));
Q_AN02 U2971 ( .A0(n785), .A1(GFidata[116]), .Z(n1713));
Q_MX02 U2972 ( .S(n808), .A0(n2566), .A1(n1713), .Z(n1712));
Q_AN02 U2973 ( .A0(n785), .A1(GFidata[117]), .Z(n1711));
Q_MX02 U2974 ( .S(n808), .A0(n2565), .A1(n1711), .Z(n1710));
Q_AN02 U2975 ( .A0(n785), .A1(GFidata[118]), .Z(n1709));
Q_MX02 U2976 ( .S(n808), .A0(n2564), .A1(n1709), .Z(n1708));
Q_AN02 U2977 ( .A0(n785), .A1(GFidata[119]), .Z(n1707));
Q_MX02 U2978 ( .S(n808), .A0(n2563), .A1(n1707), .Z(n1706));
Q_AN02 U2979 ( .A0(n785), .A1(GFidata[120]), .Z(n1705));
Q_MX02 U2980 ( .S(n808), .A0(n2562), .A1(n1705), .Z(n1704));
Q_AN02 U2981 ( .A0(n785), .A1(GFidata[121]), .Z(n1703));
Q_MX02 U2982 ( .S(n808), .A0(n2561), .A1(n1703), .Z(n1702));
Q_AN02 U2983 ( .A0(n785), .A1(GFidata[122]), .Z(n1701));
Q_MX02 U2984 ( .S(n808), .A0(n2560), .A1(n1701), .Z(n1700));
Q_AN02 U2985 ( .A0(n785), .A1(GFidata[123]), .Z(n1699));
Q_MX02 U2986 ( .S(n808), .A0(n2559), .A1(n1699), .Z(n1698));
Q_AN02 U2987 ( .A0(n785), .A1(GFidata[124]), .Z(n1697));
Q_MX02 U2988 ( .S(n808), .A0(n2558), .A1(n1697), .Z(n1696));
Q_AN02 U2989 ( .A0(n785), .A1(GFidata[125]), .Z(n1695));
Q_MX02 U2990 ( .S(n808), .A0(n2557), .A1(n1695), .Z(n1694));
Q_AN02 U2991 ( .A0(n785), .A1(GFidata[126]), .Z(n1693));
Q_MX02 U2992 ( .S(n808), .A0(n2556), .A1(n1693), .Z(n1692));
Q_AN02 U2993 ( .A0(n785), .A1(GFidata[127]), .Z(n1691));
Q_MX02 U2994 ( .S(n808), .A0(n2555), .A1(n1691), .Z(n1690));
Q_AN02 U2995 ( .A0(n785), .A1(GFidata[128]), .Z(n1689));
Q_MX02 U2996 ( .S(n808), .A0(n2554), .A1(n1689), .Z(n1688));
Q_AN02 U2997 ( .A0(n785), .A1(GFidata[129]), .Z(n1687));
Q_MX02 U2998 ( .S(n808), .A0(n2553), .A1(n1687), .Z(n1686));
Q_AN02 U2999 ( .A0(n785), .A1(GFidata[130]), .Z(n1685));
Q_MX02 U3000 ( .S(n808), .A0(n2552), .A1(n1685), .Z(n1684));
Q_AN02 U3001 ( .A0(n785), .A1(GFidata[131]), .Z(n1683));
Q_MX02 U3002 ( .S(n808), .A0(n2551), .A1(n1683), .Z(n1682));
Q_AN02 U3003 ( .A0(n785), .A1(GFidata[132]), .Z(n1681));
Q_MX02 U3004 ( .S(n808), .A0(n2550), .A1(n1681), .Z(n1680));
Q_AN02 U3005 ( .A0(n785), .A1(GFidata[133]), .Z(n1679));
Q_MX02 U3006 ( .S(n808), .A0(n2549), .A1(n1679), .Z(n1678));
Q_AN02 U3007 ( .A0(n785), .A1(GFidata[134]), .Z(n1677));
Q_MX02 U3008 ( .S(n808), .A0(n2548), .A1(n1677), .Z(n1676));
Q_AN02 U3009 ( .A0(n785), .A1(GFidata[135]), .Z(n1675));
Q_MX02 U3010 ( .S(n808), .A0(n2547), .A1(n1675), .Z(n1674));
Q_AN02 U3011 ( .A0(n785), .A1(GFidata[136]), .Z(n1673));
Q_MX02 U3012 ( .S(n808), .A0(n2546), .A1(n1673), .Z(n1672));
Q_AN02 U3013 ( .A0(n785), .A1(GFidata[137]), .Z(n1671));
Q_MX02 U3014 ( .S(n808), .A0(n2545), .A1(n1671), .Z(n1670));
Q_AN02 U3015 ( .A0(n785), .A1(GFidata[138]), .Z(n1669));
Q_MX02 U3016 ( .S(n808), .A0(n2544), .A1(n1669), .Z(n1668));
Q_AN02 U3017 ( .A0(n785), .A1(GFidata[139]), .Z(n1667));
Q_MX02 U3018 ( .S(n808), .A0(n2543), .A1(n1667), .Z(n1666));
Q_AN02 U3019 ( .A0(n785), .A1(GFidata[140]), .Z(n1665));
Q_MX02 U3020 ( .S(n808), .A0(n2542), .A1(n1665), .Z(n1664));
Q_AN02 U3021 ( .A0(n785), .A1(GFidata[141]), .Z(n1663));
Q_MX02 U3022 ( .S(n808), .A0(n2541), .A1(n1663), .Z(n1662));
Q_AN02 U3023 ( .A0(n785), .A1(GFidata[142]), .Z(n1661));
Q_MX02 U3024 ( .S(n808), .A0(n2540), .A1(n1661), .Z(n1660));
Q_AN02 U3025 ( .A0(n785), .A1(GFidata[143]), .Z(n1659));
Q_MX02 U3026 ( .S(n808), .A0(n2539), .A1(n1659), .Z(n1658));
Q_AN02 U3027 ( .A0(n785), .A1(GFidata[144]), .Z(n1657));
Q_MX02 U3028 ( .S(n808), .A0(n2538), .A1(n1657), .Z(n1656));
Q_AN02 U3029 ( .A0(n785), .A1(GFidata[145]), .Z(n1655));
Q_MX02 U3030 ( .S(n808), .A0(n2537), .A1(n1655), .Z(n1654));
Q_AN02 U3031 ( .A0(n785), .A1(GFidata[146]), .Z(n1653));
Q_MX02 U3032 ( .S(n808), .A0(n2536), .A1(n1653), .Z(n1652));
Q_AN02 U3033 ( .A0(n785), .A1(GFidata[147]), .Z(n1651));
Q_MX02 U3034 ( .S(n808), .A0(n2535), .A1(n1651), .Z(n1650));
Q_AN02 U3035 ( .A0(n785), .A1(GFidata[148]), .Z(n1649));
Q_MX02 U3036 ( .S(n808), .A0(n2534), .A1(n1649), .Z(n1648));
Q_AN02 U3037 ( .A0(n785), .A1(GFidata[149]), .Z(n1647));
Q_MX02 U3038 ( .S(n808), .A0(n2533), .A1(n1647), .Z(n1646));
Q_AN02 U3039 ( .A0(n785), .A1(GFidata[150]), .Z(n1645));
Q_MX02 U3040 ( .S(n808), .A0(n2532), .A1(n1645), .Z(n1644));
Q_AN02 U3041 ( .A0(n785), .A1(GFidata[151]), .Z(n1643));
Q_MX02 U3042 ( .S(n808), .A0(n2531), .A1(n1643), .Z(n1642));
Q_AN02 U3043 ( .A0(n785), .A1(GFidata[152]), .Z(n1641));
Q_MX02 U3044 ( .S(n808), .A0(n2530), .A1(n1641), .Z(n1640));
Q_AN02 U3045 ( .A0(n785), .A1(GFidata[153]), .Z(n1639));
Q_MX02 U3046 ( .S(n808), .A0(n2529), .A1(n1639), .Z(n1638));
Q_AN02 U3047 ( .A0(n785), .A1(GFidata[154]), .Z(n1637));
Q_MX02 U3048 ( .S(n808), .A0(n2528), .A1(n1637), .Z(n1636));
Q_AN02 U3049 ( .A0(n785), .A1(GFidata[155]), .Z(n1635));
Q_MX02 U3050 ( .S(n808), .A0(n2527), .A1(n1635), .Z(n1634));
Q_AN02 U3051 ( .A0(n785), .A1(GFidata[156]), .Z(n1633));
Q_MX02 U3052 ( .S(n808), .A0(n2526), .A1(n1633), .Z(n1632));
Q_AN02 U3053 ( .A0(n785), .A1(GFidata[157]), .Z(n1631));
Q_MX02 U3054 ( .S(n808), .A0(n2525), .A1(n1631), .Z(n1630));
Q_AN02 U3055 ( .A0(n785), .A1(GFidata[158]), .Z(n1629));
Q_MX02 U3056 ( .S(n808), .A0(n2524), .A1(n1629), .Z(n1628));
Q_AN02 U3057 ( .A0(n785), .A1(GFidata[159]), .Z(n1627));
Q_MX02 U3058 ( .S(n808), .A0(n2523), .A1(n1627), .Z(n1626));
Q_AN02 U3059 ( .A0(n785), .A1(GFidata[160]), .Z(n1625));
Q_MX02 U3060 ( .S(n808), .A0(n2522), .A1(n1625), .Z(n1624));
Q_AN02 U3061 ( .A0(n785), .A1(GFidata[161]), .Z(n1623));
Q_MX02 U3062 ( .S(n808), .A0(n2521), .A1(n1623), .Z(n1622));
Q_AN02 U3063 ( .A0(n785), .A1(GFidata[162]), .Z(n1621));
Q_MX02 U3064 ( .S(n808), .A0(n2520), .A1(n1621), .Z(n1620));
Q_AN02 U3065 ( .A0(n785), .A1(GFidata[163]), .Z(n1619));
Q_MX02 U3066 ( .S(n808), .A0(n2519), .A1(n1619), .Z(n1618));
Q_AN02 U3067 ( .A0(n785), .A1(GFidata[164]), .Z(n1617));
Q_MX02 U3068 ( .S(n808), .A0(n2518), .A1(n1617), .Z(n1616));
Q_AN02 U3069 ( .A0(n785), .A1(GFidata[165]), .Z(n1615));
Q_MX02 U3070 ( .S(n808), .A0(n2517), .A1(n1615), .Z(n1614));
Q_AN02 U3071 ( .A0(n785), .A1(GFidata[166]), .Z(n1613));
Q_MX02 U3072 ( .S(n808), .A0(n2516), .A1(n1613), .Z(n1612));
Q_AN02 U3073 ( .A0(n785), .A1(GFidata[167]), .Z(n1611));
Q_MX02 U3074 ( .S(n808), .A0(n2515), .A1(n1611), .Z(n1610));
Q_AN02 U3075 ( .A0(n785), .A1(GFidata[168]), .Z(n1609));
Q_MX02 U3076 ( .S(n808), .A0(n2514), .A1(n1609), .Z(n1608));
Q_AN02 U3077 ( .A0(n785), .A1(GFidata[169]), .Z(n1607));
Q_MX02 U3078 ( .S(n808), .A0(n2513), .A1(n1607), .Z(n1606));
Q_AN02 U3079 ( .A0(n785), .A1(GFidata[170]), .Z(n1605));
Q_MX02 U3080 ( .S(n808), .A0(n2512), .A1(n1605), .Z(n1604));
Q_AN02 U3081 ( .A0(n785), .A1(GFidata[171]), .Z(n1603));
Q_MX02 U3082 ( .S(n808), .A0(n2511), .A1(n1603), .Z(n1602));
Q_AN02 U3083 ( .A0(n785), .A1(GFidata[172]), .Z(n1601));
Q_MX02 U3084 ( .S(n808), .A0(n2510), .A1(n1601), .Z(n1600));
Q_AN02 U3085 ( .A0(n785), .A1(GFidata[173]), .Z(n1599));
Q_MX02 U3086 ( .S(n808), .A0(n2509), .A1(n1599), .Z(n1598));
Q_AN02 U3087 ( .A0(n785), .A1(GFidata[174]), .Z(n1597));
Q_MX02 U3088 ( .S(n808), .A0(n2508), .A1(n1597), .Z(n1596));
Q_AN02 U3089 ( .A0(n785), .A1(GFidata[175]), .Z(n1595));
Q_MX02 U3090 ( .S(n808), .A0(n2507), .A1(n1595), .Z(n1594));
Q_AN02 U3091 ( .A0(n785), .A1(GFidata[176]), .Z(n1593));
Q_MX02 U3092 ( .S(n808), .A0(n2506), .A1(n1593), .Z(n1592));
Q_AN02 U3093 ( .A0(n785), .A1(GFidata[177]), .Z(n1591));
Q_MX02 U3094 ( .S(n808), .A0(n2505), .A1(n1591), .Z(n1590));
Q_AN02 U3095 ( .A0(n785), .A1(GFidata[178]), .Z(n1589));
Q_MX02 U3096 ( .S(n808), .A0(n2504), .A1(n1589), .Z(n1588));
Q_AN02 U3097 ( .A0(n785), .A1(GFidata[179]), .Z(n1587));
Q_MX02 U3098 ( .S(n808), .A0(n2503), .A1(n1587), .Z(n1586));
Q_AN02 U3099 ( .A0(n785), .A1(GFidata[180]), .Z(n1585));
Q_MX02 U3100 ( .S(n808), .A0(n2502), .A1(n1585), .Z(n1584));
Q_AN02 U3101 ( .A0(n785), .A1(GFidata[181]), .Z(n1583));
Q_MX02 U3102 ( .S(n808), .A0(n2501), .A1(n1583), .Z(n1582));
Q_AN02 U3103 ( .A0(n785), .A1(GFidata[182]), .Z(n1581));
Q_MX02 U3104 ( .S(n808), .A0(n2500), .A1(n1581), .Z(n1580));
Q_AN02 U3105 ( .A0(n785), .A1(GFidata[183]), .Z(n1579));
Q_MX02 U3106 ( .S(n808), .A0(n2499), .A1(n1579), .Z(n1578));
Q_AN02 U3107 ( .A0(n785), .A1(GFidata[184]), .Z(n1577));
Q_MX02 U3108 ( .S(n808), .A0(n2498), .A1(n1577), .Z(n1576));
Q_AN02 U3109 ( .A0(n785), .A1(GFidata[185]), .Z(n1575));
Q_MX02 U3110 ( .S(n808), .A0(n2497), .A1(n1575), .Z(n1574));
Q_AN02 U3111 ( .A0(n785), .A1(GFidata[186]), .Z(n1573));
Q_MX02 U3112 ( .S(n808), .A0(n2496), .A1(n1573), .Z(n1572));
Q_AN02 U3113 ( .A0(n785), .A1(GFidata[187]), .Z(n1571));
Q_MX02 U3114 ( .S(n808), .A0(n2495), .A1(n1571), .Z(n1570));
Q_AN02 U3115 ( .A0(n785), .A1(GFidata[188]), .Z(n1569));
Q_MX02 U3116 ( .S(n808), .A0(n2494), .A1(n1569), .Z(n1568));
Q_AN02 U3117 ( .A0(n785), .A1(GFidata[189]), .Z(n1567));
Q_MX02 U3118 ( .S(n808), .A0(n2493), .A1(n1567), .Z(n1566));
Q_AN02 U3119 ( .A0(n785), .A1(GFidata[190]), .Z(n1565));
Q_MX02 U3120 ( .S(n808), .A0(n2492), .A1(n1565), .Z(n1564));
Q_AN02 U3121 ( .A0(n785), .A1(GFidata[191]), .Z(n1563));
Q_MX02 U3122 ( .S(n808), .A0(n2491), .A1(n1563), .Z(n1562));
Q_AN02 U3123 ( .A0(n785), .A1(GFidata[192]), .Z(n1561));
Q_MX02 U3124 ( .S(n808), .A0(n2490), .A1(n1561), .Z(n1560));
Q_AN02 U3125 ( .A0(n785), .A1(GFidata[193]), .Z(n1559));
Q_MX02 U3126 ( .S(n808), .A0(n2489), .A1(n1559), .Z(n1558));
Q_AN02 U3127 ( .A0(n785), .A1(GFidata[194]), .Z(n1557));
Q_MX02 U3128 ( .S(n808), .A0(n2488), .A1(n1557), .Z(n1556));
Q_AN02 U3129 ( .A0(n785), .A1(GFidata[195]), .Z(n1555));
Q_MX02 U3130 ( .S(n808), .A0(n2487), .A1(n1555), .Z(n1554));
Q_AN02 U3131 ( .A0(n785), .A1(GFidata[196]), .Z(n1553));
Q_MX02 U3132 ( .S(n808), .A0(n2486), .A1(n1553), .Z(n1552));
Q_AN02 U3133 ( .A0(n785), .A1(GFidata[197]), .Z(n1551));
Q_MX02 U3134 ( .S(n808), .A0(n2485), .A1(n1551), .Z(n1550));
Q_AN02 U3135 ( .A0(n785), .A1(GFidata[198]), .Z(n1549));
Q_MX02 U3136 ( .S(n808), .A0(n2484), .A1(n1549), .Z(n1548));
Q_AN02 U3137 ( .A0(n785), .A1(GFidata[199]), .Z(n1547));
Q_MX02 U3138 ( .S(n808), .A0(n2483), .A1(n1547), .Z(n1546));
Q_AN02 U3139 ( .A0(n785), .A1(GFidata[200]), .Z(n1545));
Q_MX02 U3140 ( .S(n808), .A0(n2482), .A1(n1545), .Z(n1544));
Q_AN02 U3141 ( .A0(n785), .A1(GFidata[201]), .Z(n1543));
Q_MX02 U3142 ( .S(n808), .A0(n2481), .A1(n1543), .Z(n1542));
Q_AN02 U3143 ( .A0(n785), .A1(GFidata[202]), .Z(n1541));
Q_MX02 U3144 ( .S(n808), .A0(n2480), .A1(n1541), .Z(n1540));
Q_AN02 U3145 ( .A0(n785), .A1(GFidata[203]), .Z(n1539));
Q_MX02 U3146 ( .S(n808), .A0(n2479), .A1(n1539), .Z(n1538));
Q_AN02 U3147 ( .A0(n785), .A1(GFidata[204]), .Z(n1537));
Q_MX02 U3148 ( .S(n808), .A0(n2478), .A1(n1537), .Z(n1536));
Q_AN02 U3149 ( .A0(n785), .A1(GFidata[205]), .Z(n1535));
Q_MX02 U3150 ( .S(n808), .A0(n2477), .A1(n1535), .Z(n1534));
Q_AN02 U3151 ( .A0(n785), .A1(GFidata[206]), .Z(n1533));
Q_MX02 U3152 ( .S(n808), .A0(n2476), .A1(n1533), .Z(n1532));
Q_AN02 U3153 ( .A0(n785), .A1(GFidata[207]), .Z(n1531));
Q_MX02 U3154 ( .S(n808), .A0(n2475), .A1(n1531), .Z(n1530));
Q_AN02 U3155 ( .A0(n785), .A1(GFidata[208]), .Z(n1529));
Q_MX02 U3156 ( .S(n808), .A0(n2474), .A1(n1529), .Z(n1528));
Q_AN02 U3157 ( .A0(n785), .A1(GFidata[209]), .Z(n1527));
Q_MX02 U3158 ( .S(n808), .A0(n2473), .A1(n1527), .Z(n1526));
Q_AN02 U3159 ( .A0(n785), .A1(GFidata[210]), .Z(n1525));
Q_MX02 U3160 ( .S(n808), .A0(n2472), .A1(n1525), .Z(n1524));
Q_AN02 U3161 ( .A0(n785), .A1(GFidata[211]), .Z(n1523));
Q_MX02 U3162 ( .S(n808), .A0(n2471), .A1(n1523), .Z(n1522));
Q_AN02 U3163 ( .A0(n785), .A1(GFidata[212]), .Z(n1521));
Q_MX02 U3164 ( .S(n808), .A0(n2470), .A1(n1521), .Z(n1520));
Q_AN02 U3165 ( .A0(n785), .A1(GFidata[213]), .Z(n1519));
Q_MX02 U3166 ( .S(n808), .A0(n2469), .A1(n1519), .Z(n1518));
Q_AN02 U3167 ( .A0(n785), .A1(GFidata[214]), .Z(n1517));
Q_MX02 U3168 ( .S(n808), .A0(n2468), .A1(n1517), .Z(n1516));
Q_AN02 U3169 ( .A0(n785), .A1(GFidata[215]), .Z(n1515));
Q_MX02 U3170 ( .S(n808), .A0(n2467), .A1(n1515), .Z(n1514));
Q_AN02 U3171 ( .A0(n785), .A1(GFidata[216]), .Z(n1513));
Q_MX02 U3172 ( .S(n808), .A0(n2466), .A1(n1513), .Z(n1512));
Q_AN02 U3173 ( .A0(n785), .A1(GFidata[217]), .Z(n1511));
Q_MX02 U3174 ( .S(n808), .A0(n2465), .A1(n1511), .Z(n1510));
Q_AN02 U3175 ( .A0(n785), .A1(GFidata[218]), .Z(n1509));
Q_MX02 U3176 ( .S(n808), .A0(n2464), .A1(n1509), .Z(n1508));
Q_AN02 U3177 ( .A0(n785), .A1(GFidata[219]), .Z(n1507));
Q_MX02 U3178 ( .S(n808), .A0(n2463), .A1(n1507), .Z(n1506));
Q_AN02 U3179 ( .A0(n785), .A1(GFidata[220]), .Z(n1505));
Q_MX02 U3180 ( .S(n808), .A0(n2462), .A1(n1505), .Z(n1504));
Q_AN02 U3181 ( .A0(n785), .A1(GFidata[221]), .Z(n1503));
Q_MX02 U3182 ( .S(n808), .A0(n2461), .A1(n1503), .Z(n1502));
Q_AN02 U3183 ( .A0(n785), .A1(GFidata[222]), .Z(n1501));
Q_MX02 U3184 ( .S(n808), .A0(n2460), .A1(n1501), .Z(n1500));
Q_AN02 U3185 ( .A0(n785), .A1(GFidata[223]), .Z(n1499));
Q_MX02 U3186 ( .S(n808), .A0(n2459), .A1(n1499), .Z(n1498));
Q_AN02 U3187 ( .A0(n785), .A1(GFidata[224]), .Z(n1497));
Q_MX02 U3188 ( .S(n808), .A0(n2458), .A1(n1497), .Z(n1496));
Q_AN02 U3189 ( .A0(n785), .A1(GFidata[225]), .Z(n1495));
Q_MX02 U3190 ( .S(n808), .A0(n2457), .A1(n1495), .Z(n1494));
Q_AN02 U3191 ( .A0(n785), .A1(GFidata[226]), .Z(n1493));
Q_MX02 U3192 ( .S(n808), .A0(n2456), .A1(n1493), .Z(n1492));
Q_AN02 U3193 ( .A0(n785), .A1(GFidata[227]), .Z(n1491));
Q_MX02 U3194 ( .S(n808), .A0(n2455), .A1(n1491), .Z(n1490));
Q_AN02 U3195 ( .A0(n785), .A1(GFidata[228]), .Z(n1489));
Q_MX02 U3196 ( .S(n808), .A0(n2454), .A1(n1489), .Z(n1488));
Q_AN02 U3197 ( .A0(n785), .A1(GFidata[229]), .Z(n1487));
Q_MX02 U3198 ( .S(n808), .A0(n2453), .A1(n1487), .Z(n1486));
Q_AN02 U3199 ( .A0(n785), .A1(GFidata[230]), .Z(n1485));
Q_MX02 U3200 ( .S(n808), .A0(n2452), .A1(n1485), .Z(n1484));
Q_AN02 U3201 ( .A0(n785), .A1(GFidata[231]), .Z(n1483));
Q_MX02 U3202 ( .S(n808), .A0(n2451), .A1(n1483), .Z(n1482));
Q_AN02 U3203 ( .A0(n785), .A1(GFidata[232]), .Z(n1481));
Q_MX02 U3204 ( .S(n808), .A0(n2450), .A1(n1481), .Z(n1480));
Q_AN02 U3205 ( .A0(n785), .A1(GFidata[233]), .Z(n1479));
Q_MX02 U3206 ( .S(n808), .A0(n2449), .A1(n1479), .Z(n1478));
Q_AN02 U3207 ( .A0(n785), .A1(GFidata[234]), .Z(n1477));
Q_MX02 U3208 ( .S(n808), .A0(n2448), .A1(n1477), .Z(n1476));
Q_AN02 U3209 ( .A0(n785), .A1(GFidata[235]), .Z(n1475));
Q_MX02 U3210 ( .S(n808), .A0(n2447), .A1(n1475), .Z(n1474));
Q_AN02 U3211 ( .A0(n785), .A1(GFidata[236]), .Z(n1473));
Q_MX02 U3212 ( .S(n808), .A0(n2446), .A1(n1473), .Z(n1472));
Q_AN02 U3213 ( .A0(n785), .A1(GFidata[237]), .Z(n1471));
Q_MX02 U3214 ( .S(n808), .A0(n2445), .A1(n1471), .Z(n1470));
Q_AN02 U3215 ( .A0(n785), .A1(GFidata[238]), .Z(n1469));
Q_MX02 U3216 ( .S(n808), .A0(n2444), .A1(n1469), .Z(n1468));
Q_AN02 U3217 ( .A0(n785), .A1(GFidata[239]), .Z(n1467));
Q_MX02 U3218 ( .S(n808), .A0(n2443), .A1(n1467), .Z(n1466));
Q_AN02 U3219 ( .A0(n785), .A1(GFidata[240]), .Z(n1465));
Q_MX02 U3220 ( .S(n808), .A0(n2442), .A1(n1465), .Z(n1464));
Q_AN02 U3221 ( .A0(n785), .A1(GFidata[241]), .Z(n1463));
Q_MX02 U3222 ( .S(n808), .A0(n2441), .A1(n1463), .Z(n1462));
Q_AN02 U3223 ( .A0(n785), .A1(GFidata[242]), .Z(n1461));
Q_MX02 U3224 ( .S(n808), .A0(n2440), .A1(n1461), .Z(n1460));
Q_AN02 U3225 ( .A0(n785), .A1(GFidata[243]), .Z(n1459));
Q_MX02 U3226 ( .S(n808), .A0(n2439), .A1(n1459), .Z(n1458));
Q_AN02 U3227 ( .A0(n785), .A1(GFidata[244]), .Z(n1457));
Q_MX02 U3228 ( .S(n808), .A0(n2438), .A1(n1457), .Z(n1456));
Q_AN02 U3229 ( .A0(n785), .A1(GFidata[245]), .Z(n1455));
Q_MX02 U3230 ( .S(n808), .A0(n2437), .A1(n1455), .Z(n1454));
Q_AN02 U3231 ( .A0(n785), .A1(GFidata[246]), .Z(n1453));
Q_MX02 U3232 ( .S(n808), .A0(n2436), .A1(n1453), .Z(n1452));
Q_AN02 U3233 ( .A0(n785), .A1(GFidata[247]), .Z(n1451));
Q_MX02 U3234 ( .S(n808), .A0(n2435), .A1(n1451), .Z(n1450));
Q_AN02 U3235 ( .A0(n785), .A1(GFidata[248]), .Z(n1449));
Q_MX02 U3236 ( .S(n808), .A0(n2434), .A1(n1449), .Z(n1448));
Q_AN02 U3237 ( .A0(n785), .A1(GFidata[249]), .Z(n1447));
Q_MX02 U3238 ( .S(n808), .A0(n2433), .A1(n1447), .Z(n1446));
Q_AN02 U3239 ( .A0(n785), .A1(GFidata[250]), .Z(n1445));
Q_MX02 U3240 ( .S(n808), .A0(n2432), .A1(n1445), .Z(n1444));
Q_AN02 U3241 ( .A0(n785), .A1(GFidata[251]), .Z(n1443));
Q_MX02 U3242 ( .S(n808), .A0(n2431), .A1(n1443), .Z(n1442));
Q_AN02 U3243 ( .A0(n785), .A1(GFidata[252]), .Z(n1441));
Q_MX02 U3244 ( .S(n808), .A0(n2430), .A1(n1441), .Z(n1440));
Q_AN02 U3245 ( .A0(n785), .A1(GFidata[253]), .Z(n1439));
Q_MX02 U3246 ( .S(n808), .A0(n2429), .A1(n1439), .Z(n1438));
Q_AN02 U3247 ( .A0(n785), .A1(GFidata[254]), .Z(n1437));
Q_MX02 U3248 ( .S(n808), .A0(n2428), .A1(n1437), .Z(n1436));
Q_AN02 U3249 ( .A0(n785), .A1(GFidata[255]), .Z(n1435));
Q_MX02 U3250 ( .S(n808), .A0(n2427), .A1(n1435), .Z(n1434));
Q_AN02 U3251 ( .A0(n785), .A1(GFidata[256]), .Z(n1433));
Q_MX02 U3252 ( .S(n808), .A0(n2426), .A1(n1433), .Z(n1432));
Q_AN02 U3253 ( .A0(n785), .A1(GFidata[257]), .Z(n1431));
Q_MX02 U3254 ( .S(n808), .A0(n2425), .A1(n1431), .Z(n1430));
Q_AN02 U3255 ( .A0(n785), .A1(GFidata[258]), .Z(n1429));
Q_MX02 U3256 ( .S(n808), .A0(n2424), .A1(n1429), .Z(n1428));
Q_AN02 U3257 ( .A0(n785), .A1(GFidata[259]), .Z(n1427));
Q_MX02 U3258 ( .S(n808), .A0(n2423), .A1(n1427), .Z(n1426));
Q_AN02 U3259 ( .A0(n785), .A1(GFidata[260]), .Z(n1425));
Q_MX02 U3260 ( .S(n808), .A0(n2422), .A1(n1425), .Z(n1424));
Q_AN02 U3261 ( .A0(n785), .A1(GFidata[261]), .Z(n1423));
Q_MX02 U3262 ( .S(n808), .A0(n2421), .A1(n1423), .Z(n1422));
Q_AN02 U3263 ( .A0(n785), .A1(GFidata[262]), .Z(n1421));
Q_MX02 U3264 ( .S(n808), .A0(n2420), .A1(n1421), .Z(n1420));
Q_AN02 U3265 ( .A0(n785), .A1(GFidata[263]), .Z(n1419));
Q_MX02 U3266 ( .S(n808), .A0(n2419), .A1(n1419), .Z(n1418));
Q_AN02 U3267 ( .A0(n785), .A1(GFidata[264]), .Z(n1417));
Q_MX02 U3268 ( .S(n808), .A0(n2418), .A1(n1417), .Z(n1416));
Q_AN02 U3269 ( .A0(n785), .A1(GFidata[265]), .Z(n1415));
Q_MX02 U3270 ( .S(n808), .A0(n2417), .A1(n1415), .Z(n1414));
Q_AN02 U3271 ( .A0(n785), .A1(GFidata[266]), .Z(n1413));
Q_MX02 U3272 ( .S(n808), .A0(n2416), .A1(n1413), .Z(n1412));
Q_AN02 U3273 ( .A0(n785), .A1(GFidata[267]), .Z(n1411));
Q_MX02 U3274 ( .S(n808), .A0(n2415), .A1(n1411), .Z(n1410));
Q_AN02 U3275 ( .A0(n785), .A1(GFidata[268]), .Z(n1409));
Q_MX02 U3276 ( .S(n808), .A0(n2414), .A1(n1409), .Z(n1408));
Q_AN02 U3277 ( .A0(n785), .A1(GFidata[269]), .Z(n1407));
Q_MX02 U3278 ( .S(n808), .A0(n2413), .A1(n1407), .Z(n1406));
Q_AN02 U3279 ( .A0(n785), .A1(GFidata[270]), .Z(n1405));
Q_MX02 U3280 ( .S(n808), .A0(n2412), .A1(n1405), .Z(n1404));
Q_AN02 U3281 ( .A0(n785), .A1(GFidata[271]), .Z(n1403));
Q_MX02 U3282 ( .S(n808), .A0(n2411), .A1(n1403), .Z(n1402));
Q_AN02 U3283 ( .A0(n785), .A1(GFidata[272]), .Z(n1401));
Q_MX02 U3284 ( .S(n808), .A0(n2410), .A1(n1401), .Z(n1400));
Q_AN02 U3285 ( .A0(n785), .A1(GFidata[273]), .Z(n1399));
Q_MX02 U3286 ( .S(n808), .A0(n2409), .A1(n1399), .Z(n1398));
Q_AN02 U3287 ( .A0(n785), .A1(GFidata[274]), .Z(n1397));
Q_MX02 U3288 ( .S(n808), .A0(n2408), .A1(n1397), .Z(n1396));
Q_AN02 U3289 ( .A0(n785), .A1(GFidata[275]), .Z(n1395));
Q_MX02 U3290 ( .S(n808), .A0(n2407), .A1(n1395), .Z(n1394));
Q_AN02 U3291 ( .A0(n785), .A1(GFidata[276]), .Z(n1393));
Q_MX02 U3292 ( .S(n808), .A0(n2406), .A1(n1393), .Z(n1392));
Q_AN02 U3293 ( .A0(n785), .A1(GFidata[277]), .Z(n1391));
Q_MX02 U3294 ( .S(n808), .A0(n2405), .A1(n1391), .Z(n1390));
Q_AN02 U3295 ( .A0(n785), .A1(GFidata[278]), .Z(n1389));
Q_MX02 U3296 ( .S(n808), .A0(n2404), .A1(n1389), .Z(n1388));
Q_AN02 U3297 ( .A0(n785), .A1(GFidata[279]), .Z(n1387));
Q_MX02 U3298 ( .S(n808), .A0(n2403), .A1(n1387), .Z(n1386));
Q_AN02 U3299 ( .A0(n785), .A1(GFidata[280]), .Z(n1385));
Q_MX02 U3300 ( .S(n808), .A0(n2402), .A1(n1385), .Z(n1384));
Q_AN02 U3301 ( .A0(n785), .A1(GFidata[281]), .Z(n1383));
Q_MX02 U3302 ( .S(n808), .A0(n2401), .A1(n1383), .Z(n1382));
Q_AN02 U3303 ( .A0(n785), .A1(GFidata[282]), .Z(n1381));
Q_MX02 U3304 ( .S(n808), .A0(n2400), .A1(n1381), .Z(n1380));
Q_AN02 U3305 ( .A0(n785), .A1(GFidata[283]), .Z(n1379));
Q_MX02 U3306 ( .S(n808), .A0(n2399), .A1(n1379), .Z(n1378));
Q_AN02 U3307 ( .A0(n785), .A1(GFidata[284]), .Z(n1377));
Q_MX02 U3308 ( .S(n808), .A0(n2398), .A1(n1377), .Z(n1376));
Q_AN02 U3309 ( .A0(n785), .A1(GFidata[285]), .Z(n1375));
Q_MX02 U3310 ( .S(n808), .A0(n2397), .A1(n1375), .Z(n1374));
Q_AN02 U3311 ( .A0(n785), .A1(GFidata[286]), .Z(n1373));
Q_MX02 U3312 ( .S(n808), .A0(n2396), .A1(n1373), .Z(n1372));
Q_AN02 U3313 ( .A0(n785), .A1(GFidata[287]), .Z(n1371));
Q_MX02 U3314 ( .S(n808), .A0(n2395), .A1(n1371), .Z(n1370));
Q_AN02 U3315 ( .A0(n785), .A1(GFidata[288]), .Z(n1369));
Q_MX02 U3316 ( .S(n808), .A0(n2394), .A1(n1369), .Z(n1368));
Q_AN02 U3317 ( .A0(n785), .A1(GFidata[289]), .Z(n1367));
Q_MX02 U3318 ( .S(n808), .A0(n2393), .A1(n1367), .Z(n1366));
Q_AN02 U3319 ( .A0(n785), .A1(GFidata[290]), .Z(n1365));
Q_MX02 U3320 ( .S(n808), .A0(n2392), .A1(n1365), .Z(n1364));
Q_AN02 U3321 ( .A0(n785), .A1(GFidata[291]), .Z(n1363));
Q_MX02 U3322 ( .S(n808), .A0(n2391), .A1(n1363), .Z(n1362));
Q_AN02 U3323 ( .A0(n785), .A1(GFidata[292]), .Z(n1361));
Q_MX02 U3324 ( .S(n808), .A0(n2390), .A1(n1361), .Z(n1360));
Q_AN02 U3325 ( .A0(n785), .A1(GFidata[293]), .Z(n1359));
Q_MX02 U3326 ( .S(n808), .A0(n2389), .A1(n1359), .Z(n1358));
Q_AN02 U3327 ( .A0(n785), .A1(GFidata[294]), .Z(n1357));
Q_MX02 U3328 ( .S(n808), .A0(n2388), .A1(n1357), .Z(n1356));
Q_AN02 U3329 ( .A0(n785), .A1(GFidata[295]), .Z(n1355));
Q_MX02 U3330 ( .S(n808), .A0(n2387), .A1(n1355), .Z(n1354));
Q_AN02 U3331 ( .A0(n785), .A1(GFidata[296]), .Z(n1353));
Q_MX02 U3332 ( .S(n808), .A0(n2386), .A1(n1353), .Z(n1352));
Q_AN02 U3333 ( .A0(n785), .A1(GFidata[297]), .Z(n1351));
Q_MX02 U3334 ( .S(n808), .A0(n2385), .A1(n1351), .Z(n1350));
Q_AN02 U3335 ( .A0(n785), .A1(GFidata[298]), .Z(n1349));
Q_MX02 U3336 ( .S(n808), .A0(n2384), .A1(n1349), .Z(n1348));
Q_AN02 U3337 ( .A0(n785), .A1(GFidata[299]), .Z(n1347));
Q_MX02 U3338 ( .S(n808), .A0(n2383), .A1(n1347), .Z(n1346));
Q_AN02 U3339 ( .A0(n785), .A1(GFidata[300]), .Z(n1345));
Q_MX02 U3340 ( .S(n808), .A0(n2382), .A1(n1345), .Z(n1344));
Q_AN02 U3341 ( .A0(n785), .A1(GFidata[301]), .Z(n1343));
Q_MX02 U3342 ( .S(n808), .A0(n2381), .A1(n1343), .Z(n1342));
Q_AN02 U3343 ( .A0(n785), .A1(GFidata[302]), .Z(n1341));
Q_MX02 U3344 ( .S(n808), .A0(n2380), .A1(n1341), .Z(n1340));
Q_AN02 U3345 ( .A0(n785), .A1(GFidata[303]), .Z(n1339));
Q_MX02 U3346 ( .S(n808), .A0(n2379), .A1(n1339), .Z(n1338));
Q_AN02 U3347 ( .A0(n785), .A1(GFidata[304]), .Z(n1337));
Q_MX02 U3348 ( .S(n808), .A0(n2378), .A1(n1337), .Z(n1336));
Q_AN02 U3349 ( .A0(n785), .A1(GFidata[305]), .Z(n1335));
Q_MX02 U3350 ( .S(n808), .A0(n2377), .A1(n1335), .Z(n1334));
Q_AN02 U3351 ( .A0(n785), .A1(GFidata[306]), .Z(n1333));
Q_MX02 U3352 ( .S(n808), .A0(n2376), .A1(n1333), .Z(n1332));
Q_AN02 U3353 ( .A0(n785), .A1(GFidata[307]), .Z(n1331));
Q_MX02 U3354 ( .S(n808), .A0(n2375), .A1(n1331), .Z(n1330));
Q_AN02 U3355 ( .A0(n785), .A1(GFidata[308]), .Z(n1329));
Q_MX02 U3356 ( .S(n808), .A0(n2374), .A1(n1329), .Z(n1328));
Q_AN02 U3357 ( .A0(n785), .A1(GFidata[309]), .Z(n1327));
Q_MX02 U3358 ( .S(n808), .A0(n2373), .A1(n1327), .Z(n1326));
Q_AN02 U3359 ( .A0(n785), .A1(GFidata[310]), .Z(n1325));
Q_MX02 U3360 ( .S(n808), .A0(n2372), .A1(n1325), .Z(n1324));
Q_AN02 U3361 ( .A0(n785), .A1(GFidata[311]), .Z(n1323));
Q_MX02 U3362 ( .S(n808), .A0(n2371), .A1(n1323), .Z(n1322));
Q_AN02 U3363 ( .A0(n785), .A1(GFidata[312]), .Z(n1321));
Q_MX02 U3364 ( .S(n808), .A0(n2370), .A1(n1321), .Z(n1320));
Q_AN02 U3365 ( .A0(n785), .A1(GFidata[313]), .Z(n1319));
Q_MX02 U3366 ( .S(n808), .A0(n2369), .A1(n1319), .Z(n1318));
Q_AN02 U3367 ( .A0(n785), .A1(GFidata[314]), .Z(n1317));
Q_MX02 U3368 ( .S(n808), .A0(n2368), .A1(n1317), .Z(n1316));
Q_AN02 U3369 ( .A0(n785), .A1(GFidata[315]), .Z(n1315));
Q_MX02 U3370 ( .S(n808), .A0(n2367), .A1(n1315), .Z(n1314));
Q_AN02 U3371 ( .A0(n785), .A1(GFidata[316]), .Z(n1313));
Q_MX02 U3372 ( .S(n808), .A0(n2366), .A1(n1313), .Z(n1312));
Q_AN02 U3373 ( .A0(n785), .A1(GFidata[317]), .Z(n1311));
Q_MX02 U3374 ( .S(n808), .A0(n2365), .A1(n1311), .Z(n1310));
Q_AN02 U3375 ( .A0(n785), .A1(GFidata[318]), .Z(n1309));
Q_MX02 U3376 ( .S(n808), .A0(n2364), .A1(n1309), .Z(n1308));
Q_AN02 U3377 ( .A0(n785), .A1(GFidata[319]), .Z(n1307));
Q_MX02 U3378 ( .S(n808), .A0(n2363), .A1(n1307), .Z(n1306));
Q_AN02 U3379 ( .A0(n785), .A1(GFidata[320]), .Z(n1305));
Q_MX02 U3380 ( .S(n808), .A0(n2362), .A1(n1305), .Z(n1304));
Q_AN02 U3381 ( .A0(n785), .A1(GFidata[321]), .Z(n1303));
Q_MX02 U3382 ( .S(n808), .A0(n2361), .A1(n1303), .Z(n1302));
Q_AN02 U3383 ( .A0(n785), .A1(GFidata[322]), .Z(n1301));
Q_MX02 U3384 ( .S(n808), .A0(n2360), .A1(n1301), .Z(n1300));
Q_AN02 U3385 ( .A0(n785), .A1(GFidata[323]), .Z(n1299));
Q_MX02 U3386 ( .S(n808), .A0(n2359), .A1(n1299), .Z(n1298));
Q_AN02 U3387 ( .A0(n785), .A1(GFidata[324]), .Z(n1297));
Q_MX02 U3388 ( .S(n808), .A0(n2358), .A1(n1297), .Z(n1296));
Q_AN02 U3389 ( .A0(n785), .A1(GFidata[325]), .Z(n1295));
Q_MX02 U3390 ( .S(n808), .A0(n2357), .A1(n1295), .Z(n1294));
Q_AN02 U3391 ( .A0(n785), .A1(GFidata[326]), .Z(n1293));
Q_MX02 U3392 ( .S(n808), .A0(n2356), .A1(n1293), .Z(n1292));
Q_AN02 U3393 ( .A0(n785), .A1(GFidata[327]), .Z(n1291));
Q_MX02 U3394 ( .S(n808), .A0(n2355), .A1(n1291), .Z(n1290));
Q_AN02 U3395 ( .A0(n785), .A1(GFidata[328]), .Z(n1289));
Q_MX02 U3396 ( .S(n808), .A0(n2354), .A1(n1289), .Z(n1288));
Q_AN02 U3397 ( .A0(n785), .A1(GFidata[329]), .Z(n1287));
Q_MX02 U3398 ( .S(n808), .A0(n2353), .A1(n1287), .Z(n1286));
Q_AN02 U3399 ( .A0(n785), .A1(GFidata[330]), .Z(n1285));
Q_MX02 U3400 ( .S(n808), .A0(n2352), .A1(n1285), .Z(n1284));
Q_AN02 U3401 ( .A0(n785), .A1(GFidata[331]), .Z(n1283));
Q_MX02 U3402 ( .S(n808), .A0(n2351), .A1(n1283), .Z(n1282));
Q_AN02 U3403 ( .A0(n785), .A1(GFidata[332]), .Z(n1281));
Q_MX02 U3404 ( .S(n808), .A0(n2350), .A1(n1281), .Z(n1280));
Q_AN02 U3405 ( .A0(n785), .A1(GFidata[333]), .Z(n1279));
Q_MX02 U3406 ( .S(n808), .A0(n2349), .A1(n1279), .Z(n1278));
Q_AN02 U3407 ( .A0(n785), .A1(GFidata[334]), .Z(n1277));
Q_MX02 U3408 ( .S(n808), .A0(n2348), .A1(n1277), .Z(n1276));
Q_AN02 U3409 ( .A0(n785), .A1(GFidata[335]), .Z(n1275));
Q_MX02 U3410 ( .S(n808), .A0(n2347), .A1(n1275), .Z(n1274));
Q_AN02 U3411 ( .A0(n785), .A1(GFidata[336]), .Z(n1273));
Q_MX02 U3412 ( .S(n808), .A0(n2346), .A1(n1273), .Z(n1272));
Q_AN02 U3413 ( .A0(n785), .A1(GFidata[337]), .Z(n1271));
Q_MX02 U3414 ( .S(n808), .A0(n2345), .A1(n1271), .Z(n1270));
Q_AN02 U3415 ( .A0(n785), .A1(GFidata[338]), .Z(n1269));
Q_MX02 U3416 ( .S(n808), .A0(n2344), .A1(n1269), .Z(n1268));
Q_AN02 U3417 ( .A0(n785), .A1(GFidata[339]), .Z(n1267));
Q_MX02 U3418 ( .S(n808), .A0(n2343), .A1(n1267), .Z(n1266));
Q_AN02 U3419 ( .A0(n785), .A1(GFidata[340]), .Z(n1265));
Q_MX02 U3420 ( .S(n808), .A0(n2342), .A1(n1265), .Z(n1264));
Q_AN02 U3421 ( .A0(n785), .A1(GFidata[341]), .Z(n1263));
Q_MX02 U3422 ( .S(n808), .A0(n2341), .A1(n1263), .Z(n1262));
Q_AN02 U3423 ( .A0(n785), .A1(GFidata[342]), .Z(n1261));
Q_MX02 U3424 ( .S(n808), .A0(n2340), .A1(n1261), .Z(n1260));
Q_AN02 U3425 ( .A0(n785), .A1(GFidata[343]), .Z(n1259));
Q_MX02 U3426 ( .S(n808), .A0(n2339), .A1(n1259), .Z(n1258));
Q_AN02 U3427 ( .A0(n785), .A1(GFidata[344]), .Z(n1257));
Q_MX02 U3428 ( .S(n808), .A0(n2338), .A1(n1257), .Z(n1256));
Q_AN02 U3429 ( .A0(n785), .A1(GFidata[345]), .Z(n1255));
Q_MX02 U3430 ( .S(n808), .A0(n2337), .A1(n1255), .Z(n1254));
Q_AN02 U3431 ( .A0(n785), .A1(GFidata[346]), .Z(n1253));
Q_MX02 U3432 ( .S(n808), .A0(n2336), .A1(n1253), .Z(n1252));
Q_AN02 U3433 ( .A0(n785), .A1(GFidata[347]), .Z(n1251));
Q_MX02 U3434 ( .S(n808), .A0(n2335), .A1(n1251), .Z(n1250));
Q_AN02 U3435 ( .A0(n785), .A1(GFidata[348]), .Z(n1249));
Q_MX02 U3436 ( .S(n808), .A0(n2334), .A1(n1249), .Z(n1248));
Q_AN02 U3437 ( .A0(n785), .A1(GFidata[349]), .Z(n1247));
Q_MX02 U3438 ( .S(n808), .A0(n2333), .A1(n1247), .Z(n1246));
Q_AN02 U3439 ( .A0(n785), .A1(GFidata[350]), .Z(n1245));
Q_MX02 U3440 ( .S(n808), .A0(n2332), .A1(n1245), .Z(n1244));
Q_AN02 U3441 ( .A0(n785), .A1(GFidata[351]), .Z(n1243));
Q_MX02 U3442 ( .S(n808), .A0(n2331), .A1(n1243), .Z(n1242));
Q_AN02 U3443 ( .A0(n785), .A1(GFidata[352]), .Z(n1241));
Q_MX02 U3444 ( .S(n808), .A0(n2330), .A1(n1241), .Z(n1240));
Q_AN02 U3445 ( .A0(n785), .A1(GFidata[353]), .Z(n1239));
Q_MX02 U3446 ( .S(n808), .A0(n2329), .A1(n1239), .Z(n1238));
Q_AN02 U3447 ( .A0(n785), .A1(GFidata[354]), .Z(n1237));
Q_MX02 U3448 ( .S(n808), .A0(n2328), .A1(n1237), .Z(n1236));
Q_AN02 U3449 ( .A0(n785), .A1(GFidata[355]), .Z(n1235));
Q_MX02 U3450 ( .S(n808), .A0(n2327), .A1(n1235), .Z(n1234));
Q_AN02 U3451 ( .A0(n785), .A1(GFidata[356]), .Z(n1233));
Q_MX02 U3452 ( .S(n808), .A0(n2326), .A1(n1233), .Z(n1232));
Q_AN02 U3453 ( .A0(n785), .A1(GFidata[357]), .Z(n1231));
Q_MX02 U3454 ( .S(n808), .A0(n2325), .A1(n1231), .Z(n1230));
Q_AN02 U3455 ( .A0(n785), .A1(GFidata[358]), .Z(n1229));
Q_MX02 U3456 ( .S(n808), .A0(n2324), .A1(n1229), .Z(n1228));
Q_AN02 U3457 ( .A0(n785), .A1(GFidata[359]), .Z(n1227));
Q_MX02 U3458 ( .S(n808), .A0(n2323), .A1(n1227), .Z(n1226));
Q_AN02 U3459 ( .A0(n785), .A1(GFidata[360]), .Z(n1225));
Q_MX02 U3460 ( .S(n808), .A0(n2322), .A1(n1225), .Z(n1224));
Q_AN02 U3461 ( .A0(n785), .A1(GFidata[361]), .Z(n1223));
Q_MX02 U3462 ( .S(n808), .A0(n2321), .A1(n1223), .Z(n1222));
Q_AN02 U3463 ( .A0(n785), .A1(GFidata[362]), .Z(n1221));
Q_MX02 U3464 ( .S(n808), .A0(n2320), .A1(n1221), .Z(n1220));
Q_AN02 U3465 ( .A0(n785), .A1(GFidata[363]), .Z(n1219));
Q_MX02 U3466 ( .S(n808), .A0(n2319), .A1(n1219), .Z(n1218));
Q_AN02 U3467 ( .A0(n785), .A1(GFidata[364]), .Z(n1217));
Q_MX02 U3468 ( .S(n808), .A0(n2318), .A1(n1217), .Z(n1216));
Q_AN02 U3469 ( .A0(n785), .A1(GFidata[365]), .Z(n1215));
Q_MX02 U3470 ( .S(n808), .A0(n2317), .A1(n1215), .Z(n1214));
Q_AN02 U3471 ( .A0(n785), .A1(GFidata[366]), .Z(n1213));
Q_MX02 U3472 ( .S(n808), .A0(n2316), .A1(n1213), .Z(n1212));
Q_AN02 U3473 ( .A0(n785), .A1(GFidata[367]), .Z(n1211));
Q_MX02 U3474 ( .S(n808), .A0(n2315), .A1(n1211), .Z(n1210));
Q_AN02 U3475 ( .A0(n785), .A1(GFidata[368]), .Z(n1209));
Q_MX02 U3476 ( .S(n808), .A0(n2314), .A1(n1209), .Z(n1208));
Q_AN02 U3477 ( .A0(n785), .A1(GFidata[369]), .Z(n1207));
Q_MX02 U3478 ( .S(n808), .A0(n2313), .A1(n1207), .Z(n1206));
Q_AN02 U3479 ( .A0(n785), .A1(GFidata[370]), .Z(n1205));
Q_MX02 U3480 ( .S(n808), .A0(n2312), .A1(n1205), .Z(n1204));
Q_AN02 U3481 ( .A0(n785), .A1(GFidata[371]), .Z(n1203));
Q_MX02 U3482 ( .S(n808), .A0(n2311), .A1(n1203), .Z(n1202));
Q_AN02 U3483 ( .A0(n785), .A1(GFidata[372]), .Z(n1201));
Q_MX02 U3484 ( .S(n808), .A0(n2310), .A1(n1201), .Z(n1200));
Q_AN02 U3485 ( .A0(n785), .A1(GFidata[373]), .Z(n1199));
Q_MX02 U3486 ( .S(n808), .A0(n2309), .A1(n1199), .Z(n1198));
Q_AN02 U3487 ( .A0(n785), .A1(GFidata[374]), .Z(n1197));
Q_MX02 U3488 ( .S(n808), .A0(n2308), .A1(n1197), .Z(n1196));
Q_AN02 U3489 ( .A0(n785), .A1(GFidata[375]), .Z(n1195));
Q_MX02 U3490 ( .S(n808), .A0(n2307), .A1(n1195), .Z(n1194));
Q_AN02 U3491 ( .A0(n785), .A1(GFidata[376]), .Z(n1193));
Q_MX02 U3492 ( .S(n808), .A0(n2306), .A1(n1193), .Z(n1192));
Q_AN02 U3493 ( .A0(n785), .A1(GFidata[377]), .Z(n1191));
Q_MX02 U3494 ( .S(n808), .A0(n2305), .A1(n1191), .Z(n1190));
Q_AN02 U3495 ( .A0(n785), .A1(GFidata[378]), .Z(n1189));
Q_MX02 U3496 ( .S(n808), .A0(n2304), .A1(n1189), .Z(n1188));
Q_AN02 U3497 ( .A0(n785), .A1(GFidata[379]), .Z(n1187));
Q_MX02 U3498 ( .S(n808), .A0(n2303), .A1(n1187), .Z(n1186));
Q_AN02 U3499 ( .A0(n785), .A1(GFidata[380]), .Z(n1185));
Q_MX02 U3500 ( .S(n808), .A0(n2302), .A1(n1185), .Z(n1184));
Q_AN02 U3501 ( .A0(n785), .A1(GFidata[381]), .Z(n1183));
Q_MX02 U3502 ( .S(n808), .A0(n2301), .A1(n1183), .Z(n1182));
Q_AN02 U3503 ( .A0(n785), .A1(GFidata[382]), .Z(n1181));
Q_MX02 U3504 ( .S(n808), .A0(n2300), .A1(n1181), .Z(n1180));
Q_AN02 U3505 ( .A0(n785), .A1(GFidata[383]), .Z(n1179));
Q_MX02 U3506 ( .S(n808), .A0(n2299), .A1(n1179), .Z(n1178));
Q_AN02 U3507 ( .A0(n785), .A1(GFidata[384]), .Z(n1177));
Q_MX02 U3508 ( .S(n808), .A0(n2298), .A1(n1177), .Z(n1176));
Q_AN02 U3509 ( .A0(n785), .A1(GFidata[385]), .Z(n1175));
Q_MX02 U3510 ( .S(n808), .A0(n2297), .A1(n1175), .Z(n1174));
Q_AN02 U3511 ( .A0(n785), .A1(GFidata[386]), .Z(n1173));
Q_MX02 U3512 ( .S(n808), .A0(n2296), .A1(n1173), .Z(n1172));
Q_AN02 U3513 ( .A0(n785), .A1(GFidata[387]), .Z(n1171));
Q_MX02 U3514 ( .S(n808), .A0(n2295), .A1(n1171), .Z(n1170));
Q_AN02 U3515 ( .A0(n785), .A1(GFidata[388]), .Z(n1169));
Q_MX02 U3516 ( .S(n808), .A0(n2294), .A1(n1169), .Z(n1168));
Q_AN02 U3517 ( .A0(n785), .A1(GFidata[389]), .Z(n1167));
Q_MX02 U3518 ( .S(n808), .A0(n2293), .A1(n1167), .Z(n1166));
Q_AN02 U3519 ( .A0(n785), .A1(GFidata[390]), .Z(n1165));
Q_MX02 U3520 ( .S(n808), .A0(n2292), .A1(n1165), .Z(n1164));
Q_AN02 U3521 ( .A0(n785), .A1(GFidata[391]), .Z(n1163));
Q_MX02 U3522 ( .S(n808), .A0(n2291), .A1(n1163), .Z(n1162));
Q_AN02 U3523 ( .A0(n785), .A1(GFidata[392]), .Z(n1161));
Q_MX02 U3524 ( .S(n808), .A0(n2290), .A1(n1161), .Z(n1160));
Q_AN02 U3525 ( .A0(n785), .A1(GFidata[393]), .Z(n1159));
Q_MX02 U3526 ( .S(n808), .A0(n2289), .A1(n1159), .Z(n1158));
Q_AN02 U3527 ( .A0(n785), .A1(GFidata[394]), .Z(n1157));
Q_MX02 U3528 ( .S(n808), .A0(n2288), .A1(n1157), .Z(n1156));
Q_AN02 U3529 ( .A0(n785), .A1(GFidata[395]), .Z(n1155));
Q_MX02 U3530 ( .S(n808), .A0(n2287), .A1(n1155), .Z(n1154));
Q_AN02 U3531 ( .A0(n785), .A1(GFidata[396]), .Z(n1153));
Q_MX02 U3532 ( .S(n808), .A0(n2286), .A1(n1153), .Z(n1152));
Q_AN02 U3533 ( .A0(n785), .A1(GFidata[397]), .Z(n1151));
Q_MX02 U3534 ( .S(n808), .A0(n2285), .A1(n1151), .Z(n1150));
Q_AN02 U3535 ( .A0(n785), .A1(GFidata[398]), .Z(n1149));
Q_MX02 U3536 ( .S(n808), .A0(n2284), .A1(n1149), .Z(n1148));
Q_AN02 U3537 ( .A0(n785), .A1(GFidata[399]), .Z(n1147));
Q_MX02 U3538 ( .S(n808), .A0(n2283), .A1(n1147), .Z(n1146));
Q_AN02 U3539 ( .A0(n785), .A1(GFidata[400]), .Z(n1145));
Q_MX02 U3540 ( .S(n808), .A0(n2282), .A1(n1145), .Z(n1144));
Q_AN02 U3541 ( .A0(n785), .A1(GFidata[401]), .Z(n1143));
Q_MX02 U3542 ( .S(n808), .A0(n2281), .A1(n1143), .Z(n1142));
Q_AN02 U3543 ( .A0(n785), .A1(GFidata[402]), .Z(n1141));
Q_MX02 U3544 ( .S(n808), .A0(n2280), .A1(n1141), .Z(n1140));
Q_AN02 U3545 ( .A0(n785), .A1(GFidata[403]), .Z(n1139));
Q_MX02 U3546 ( .S(n808), .A0(n2279), .A1(n1139), .Z(n1138));
Q_AN02 U3547 ( .A0(n785), .A1(GFidata[404]), .Z(n1137));
Q_MX02 U3548 ( .S(n808), .A0(n2278), .A1(n1137), .Z(n1136));
Q_AN02 U3549 ( .A0(n785), .A1(GFidata[405]), .Z(n1135));
Q_MX02 U3550 ( .S(n808), .A0(n2277), .A1(n1135), .Z(n1134));
Q_AN02 U3551 ( .A0(n785), .A1(GFidata[406]), .Z(n1133));
Q_MX02 U3552 ( .S(n808), .A0(n2276), .A1(n1133), .Z(n1132));
Q_AN02 U3553 ( .A0(n785), .A1(GFidata[407]), .Z(n1131));
Q_MX02 U3554 ( .S(n808), .A0(n2275), .A1(n1131), .Z(n1130));
Q_AN02 U3555 ( .A0(n785), .A1(GFidata[408]), .Z(n1129));
Q_MX02 U3556 ( .S(n808), .A0(n2274), .A1(n1129), .Z(n1128));
Q_AN02 U3557 ( .A0(n785), .A1(GFidata[409]), .Z(n1127));
Q_MX02 U3558 ( .S(n808), .A0(n2273), .A1(n1127), .Z(n1126));
Q_AN02 U3559 ( .A0(n785), .A1(GFidata[410]), .Z(n1125));
Q_MX02 U3560 ( .S(n808), .A0(n2272), .A1(n1125), .Z(n1124));
Q_AN02 U3561 ( .A0(n785), .A1(GFidata[411]), .Z(n1123));
Q_MX02 U3562 ( .S(n808), .A0(n2271), .A1(n1123), .Z(n1122));
Q_AN02 U3563 ( .A0(n785), .A1(GFidata[412]), .Z(n1121));
Q_MX02 U3564 ( .S(n808), .A0(n2270), .A1(n1121), .Z(n1120));
Q_AN02 U3565 ( .A0(n785), .A1(GFidata[413]), .Z(n1119));
Q_MX02 U3566 ( .S(n808), .A0(n2269), .A1(n1119), .Z(n1118));
Q_AN02 U3567 ( .A0(n785), .A1(GFidata[414]), .Z(n1117));
Q_MX02 U3568 ( .S(n808), .A0(n2268), .A1(n1117), .Z(n1116));
Q_AN02 U3569 ( .A0(n785), .A1(GFidata[415]), .Z(n1115));
Q_MX02 U3570 ( .S(n808), .A0(n2267), .A1(n1115), .Z(n1114));
Q_AN02 U3571 ( .A0(n785), .A1(GFidata[416]), .Z(n1113));
Q_MX02 U3572 ( .S(n808), .A0(n2266), .A1(n1113), .Z(n1112));
Q_AN02 U3573 ( .A0(n785), .A1(GFidata[417]), .Z(n1111));
Q_MX02 U3574 ( .S(n808), .A0(n2265), .A1(n1111), .Z(n1110));
Q_AN02 U3575 ( .A0(n785), .A1(GFidata[418]), .Z(n1109));
Q_MX02 U3576 ( .S(n808), .A0(n2264), .A1(n1109), .Z(n1108));
Q_AN02 U3577 ( .A0(n785), .A1(GFidata[419]), .Z(n1107));
Q_MX02 U3578 ( .S(n808), .A0(n2263), .A1(n1107), .Z(n1106));
Q_AN02 U3579 ( .A0(n785), .A1(GFidata[420]), .Z(n1105));
Q_MX02 U3580 ( .S(n808), .A0(n2262), .A1(n1105), .Z(n1104));
Q_AN02 U3581 ( .A0(n785), .A1(GFidata[421]), .Z(n1103));
Q_MX02 U3582 ( .S(n808), .A0(n2261), .A1(n1103), .Z(n1102));
Q_AN02 U3583 ( .A0(n785), .A1(GFidata[422]), .Z(n1101));
Q_MX02 U3584 ( .S(n808), .A0(n2260), .A1(n1101), .Z(n1100));
Q_AN02 U3585 ( .A0(n785), .A1(GFidata[423]), .Z(n1099));
Q_MX02 U3586 ( .S(n808), .A0(n2259), .A1(n1099), .Z(n1098));
Q_AN02 U3587 ( .A0(n785), .A1(GFidata[424]), .Z(n1097));
Q_MX02 U3588 ( .S(n808), .A0(n2258), .A1(n1097), .Z(n1096));
Q_AN02 U3589 ( .A0(n785), .A1(GFidata[425]), .Z(n1095));
Q_MX02 U3590 ( .S(n808), .A0(n2257), .A1(n1095), .Z(n1094));
Q_AN02 U3591 ( .A0(n785), .A1(GFidata[426]), .Z(n1093));
Q_MX02 U3592 ( .S(n808), .A0(n2256), .A1(n1093), .Z(n1092));
Q_AN02 U3593 ( .A0(n785), .A1(GFidata[427]), .Z(n1091));
Q_MX02 U3594 ( .S(n808), .A0(n2255), .A1(n1091), .Z(n1090));
Q_AN02 U3595 ( .A0(n785), .A1(GFidata[428]), .Z(n1089));
Q_MX02 U3596 ( .S(n808), .A0(n2254), .A1(n1089), .Z(n1088));
Q_AN02 U3597 ( .A0(n785), .A1(GFidata[429]), .Z(n1087));
Q_MX02 U3598 ( .S(n808), .A0(n2253), .A1(n1087), .Z(n1086));
Q_AN02 U3599 ( .A0(n785), .A1(GFidata[430]), .Z(n1085));
Q_MX02 U3600 ( .S(n808), .A0(n2252), .A1(n1085), .Z(n1084));
Q_AN02 U3601 ( .A0(n785), .A1(GFidata[431]), .Z(n1083));
Q_MX02 U3602 ( .S(n808), .A0(n2251), .A1(n1083), .Z(n1082));
Q_AN02 U3603 ( .A0(n785), .A1(GFidata[432]), .Z(n1081));
Q_MX02 U3604 ( .S(n808), .A0(n2250), .A1(n1081), .Z(n1080));
Q_AN02 U3605 ( .A0(n785), .A1(GFidata[433]), .Z(n1079));
Q_MX02 U3606 ( .S(n808), .A0(n2249), .A1(n1079), .Z(n1078));
Q_AN02 U3607 ( .A0(n785), .A1(GFidata[434]), .Z(n1077));
Q_MX02 U3608 ( .S(n808), .A0(n2248), .A1(n1077), .Z(n1076));
Q_AN02 U3609 ( .A0(n785), .A1(GFidata[435]), .Z(n1075));
Q_MX02 U3610 ( .S(n808), .A0(n2247), .A1(n1075), .Z(n1074));
Q_AN02 U3611 ( .A0(n785), .A1(GFidata[436]), .Z(n1073));
Q_MX02 U3612 ( .S(n808), .A0(n2246), .A1(n1073), .Z(n1072));
Q_AN02 U3613 ( .A0(n785), .A1(GFidata[437]), .Z(n1071));
Q_MX02 U3614 ( .S(n808), .A0(n2245), .A1(n1071), .Z(n1070));
Q_AN02 U3615 ( .A0(n785), .A1(GFidata[438]), .Z(n1069));
Q_MX02 U3616 ( .S(n808), .A0(n2244), .A1(n1069), .Z(n1068));
Q_AN02 U3617 ( .A0(n785), .A1(GFidata[439]), .Z(n1067));
Q_MX02 U3618 ( .S(n808), .A0(n2243), .A1(n1067), .Z(n1066));
Q_AN02 U3619 ( .A0(n785), .A1(GFidata[440]), .Z(n1065));
Q_MX02 U3620 ( .S(n808), .A0(n2242), .A1(n1065), .Z(n1064));
Q_AN02 U3621 ( .A0(n785), .A1(GFidata[441]), .Z(n1063));
Q_MX02 U3622 ( .S(n808), .A0(n2241), .A1(n1063), .Z(n1062));
Q_AN02 U3623 ( .A0(n785), .A1(GFidata[442]), .Z(n1061));
Q_MX02 U3624 ( .S(n808), .A0(n2240), .A1(n1061), .Z(n1060));
Q_AN02 U3625 ( .A0(n785), .A1(GFidata[443]), .Z(n1059));
Q_MX02 U3626 ( .S(n808), .A0(n2239), .A1(n1059), .Z(n1058));
Q_AN02 U3627 ( .A0(n785), .A1(GFidata[444]), .Z(n1057));
Q_MX02 U3628 ( .S(n808), .A0(n2238), .A1(n1057), .Z(n1056));
Q_AN02 U3629 ( .A0(n785), .A1(GFidata[445]), .Z(n1055));
Q_MX02 U3630 ( .S(n808), .A0(n2237), .A1(n1055), .Z(n1054));
Q_AN02 U3631 ( .A0(n785), .A1(GFidata[446]), .Z(n1053));
Q_MX02 U3632 ( .S(n808), .A0(n2236), .A1(n1053), .Z(n1052));
Q_AN02 U3633 ( .A0(n785), .A1(GFidata[447]), .Z(n1051));
Q_MX02 U3634 ( .S(n808), .A0(n2235), .A1(n1051), .Z(n1050));
Q_AN02 U3635 ( .A0(n785), .A1(GFidata[448]), .Z(n1049));
Q_MX02 U3636 ( .S(n808), .A0(n2234), .A1(n1049), .Z(n1048));
Q_AN02 U3637 ( .A0(n785), .A1(GFidata[449]), .Z(n1047));
Q_MX02 U3638 ( .S(n808), .A0(n2233), .A1(n1047), .Z(n1046));
Q_AN02 U3639 ( .A0(n785), .A1(GFidata[450]), .Z(n1045));
Q_MX02 U3640 ( .S(n808), .A0(n2232), .A1(n1045), .Z(n1044));
Q_AN02 U3641 ( .A0(n785), .A1(GFidata[451]), .Z(n1043));
Q_MX02 U3642 ( .S(n808), .A0(n2231), .A1(n1043), .Z(n1042));
Q_AN02 U3643 ( .A0(n785), .A1(GFidata[452]), .Z(n1041));
Q_MX02 U3644 ( .S(n808), .A0(n2230), .A1(n1041), .Z(n1040));
Q_AN02 U3645 ( .A0(n785), .A1(GFidata[453]), .Z(n1039));
Q_MX02 U3646 ( .S(n808), .A0(n2229), .A1(n1039), .Z(n1038));
Q_AN02 U3647 ( .A0(n785), .A1(GFidata[454]), .Z(n1037));
Q_MX02 U3648 ( .S(n808), .A0(n2228), .A1(n1037), .Z(n1036));
Q_AN02 U3649 ( .A0(n785), .A1(GFidata[455]), .Z(n1035));
Q_MX02 U3650 ( .S(n808), .A0(n2227), .A1(n1035), .Z(n1034));
Q_AN02 U3651 ( .A0(n785), .A1(GFidata[456]), .Z(n1033));
Q_MX02 U3652 ( .S(n808), .A0(n2226), .A1(n1033), .Z(n1032));
Q_AN02 U3653 ( .A0(n785), .A1(GFidata[457]), .Z(n1031));
Q_MX02 U3654 ( .S(n808), .A0(n2225), .A1(n1031), .Z(n1030));
Q_AN02 U3655 ( .A0(n785), .A1(GFidata[458]), .Z(n1029));
Q_MX02 U3656 ( .S(n808), .A0(n2224), .A1(n1029), .Z(n1028));
Q_AN02 U3657 ( .A0(n785), .A1(GFidata[459]), .Z(n1027));
Q_MX02 U3658 ( .S(n808), .A0(n2223), .A1(n1027), .Z(n1026));
Q_AN02 U3659 ( .A0(n785), .A1(GFidata[460]), .Z(n1025));
Q_MX02 U3660 ( .S(n808), .A0(n2222), .A1(n1025), .Z(n1024));
Q_AN02 U3661 ( .A0(n785), .A1(GFidata[461]), .Z(n1023));
Q_MX02 U3662 ( .S(n808), .A0(n2221), .A1(n1023), .Z(n1022));
Q_AN02 U3663 ( .A0(n785), .A1(GFidata[462]), .Z(n1021));
Q_MX02 U3664 ( .S(n808), .A0(n2220), .A1(n1021), .Z(n1020));
Q_AN02 U3665 ( .A0(n785), .A1(GFidata[463]), .Z(n1019));
Q_MX02 U3666 ( .S(n808), .A0(n2219), .A1(n1019), .Z(n1018));
Q_AN02 U3667 ( .A0(n785), .A1(GFidata[464]), .Z(n1017));
Q_MX02 U3668 ( .S(n808), .A0(n2218), .A1(n1017), .Z(n1016));
Q_AN02 U3669 ( .A0(n785), .A1(GFidata[465]), .Z(n1015));
Q_MX02 U3670 ( .S(n808), .A0(n2217), .A1(n1015), .Z(n1014));
Q_AN02 U3671 ( .A0(n785), .A1(GFidata[466]), .Z(n1013));
Q_MX02 U3672 ( .S(n808), .A0(n2216), .A1(n1013), .Z(n1012));
Q_AN02 U3673 ( .A0(n785), .A1(GFidata[467]), .Z(n1011));
Q_MX02 U3674 ( .S(n808), .A0(n2215), .A1(n1011), .Z(n1010));
Q_AN02 U3675 ( .A0(n785), .A1(GFidata[468]), .Z(n1009));
Q_MX02 U3676 ( .S(n808), .A0(n2214), .A1(n1009), .Z(n1008));
Q_AN02 U3677 ( .A0(n785), .A1(GFidata[469]), .Z(n1007));
Q_MX02 U3678 ( .S(n808), .A0(n2213), .A1(n1007), .Z(n1006));
Q_AN02 U3679 ( .A0(n785), .A1(GFidata[470]), .Z(n1005));
Q_MX02 U3680 ( .S(n808), .A0(n2212), .A1(n1005), .Z(n1004));
Q_AN02 U3681 ( .A0(n785), .A1(GFidata[471]), .Z(n1003));
Q_MX02 U3682 ( .S(n808), .A0(n2211), .A1(n1003), .Z(n1002));
Q_AN02 U3683 ( .A0(n785), .A1(GFidata[472]), .Z(n1001));
Q_MX02 U3684 ( .S(n808), .A0(n2210), .A1(n1001), .Z(n1000));
Q_AN02 U3685 ( .A0(n785), .A1(GFidata[473]), .Z(n999));
Q_MX02 U3686 ( .S(n808), .A0(n2209), .A1(n999), .Z(n998));
Q_AN02 U3687 ( .A0(n785), .A1(GFidata[474]), .Z(n997));
Q_MX02 U3688 ( .S(n808), .A0(n2208), .A1(n997), .Z(n996));
Q_AN02 U3689 ( .A0(n785), .A1(GFidata[475]), .Z(n995));
Q_MX02 U3690 ( .S(n808), .A0(n2207), .A1(n995), .Z(n994));
Q_AN02 U3691 ( .A0(n785), .A1(GFidata[476]), .Z(n993));
Q_MX02 U3692 ( .S(n808), .A0(n2206), .A1(n993), .Z(n992));
Q_AN02 U3693 ( .A0(n785), .A1(GFidata[477]), .Z(n991));
Q_MX02 U3694 ( .S(n808), .A0(n2205), .A1(n991), .Z(n990));
Q_AN02 U3695 ( .A0(n785), .A1(GFidata[478]), .Z(n989));
Q_MX02 U3696 ( .S(n808), .A0(n2204), .A1(n989), .Z(n988));
Q_AN02 U3697 ( .A0(n785), .A1(GFidata[479]), .Z(n987));
Q_MX02 U3698 ( .S(n808), .A0(n2203), .A1(n987), .Z(n986));
Q_AN02 U3699 ( .A0(n785), .A1(GFidata[480]), .Z(n985));
Q_MX02 U3700 ( .S(n808), .A0(n2202), .A1(n985), .Z(n984));
Q_AN02 U3701 ( .A0(n785), .A1(GFidata[481]), .Z(n983));
Q_MX02 U3702 ( .S(n808), .A0(n2201), .A1(n983), .Z(n982));
Q_AN02 U3703 ( .A0(n785), .A1(GFidata[482]), .Z(n981));
Q_MX02 U3704 ( .S(n808), .A0(n2200), .A1(n981), .Z(n980));
Q_AN02 U3705 ( .A0(n785), .A1(GFidata[483]), .Z(n979));
Q_MX02 U3706 ( .S(n808), .A0(n2199), .A1(n979), .Z(n978));
Q_AN02 U3707 ( .A0(n785), .A1(GFidata[484]), .Z(n977));
Q_MX02 U3708 ( .S(n808), .A0(n2198), .A1(n977), .Z(n976));
Q_AN02 U3709 ( .A0(n785), .A1(GFidata[485]), .Z(n975));
Q_MX02 U3710 ( .S(n808), .A0(n2197), .A1(n975), .Z(n974));
Q_AN02 U3711 ( .A0(n785), .A1(GFidata[486]), .Z(n973));
Q_MX02 U3712 ( .S(n808), .A0(n2196), .A1(n973), .Z(n972));
Q_AN02 U3713 ( .A0(n785), .A1(GFidata[487]), .Z(n971));
Q_MX02 U3714 ( .S(n808), .A0(n2195), .A1(n971), .Z(n970));
Q_AN02 U3715 ( .A0(n785), .A1(GFidata[488]), .Z(n969));
Q_MX02 U3716 ( .S(n808), .A0(n2194), .A1(n969), .Z(n968));
Q_AN02 U3717 ( .A0(n785), .A1(GFidata[489]), .Z(n967));
Q_MX02 U3718 ( .S(n808), .A0(n2193), .A1(n967), .Z(n966));
Q_AN02 U3719 ( .A0(n785), .A1(GFidata[490]), .Z(n965));
Q_MX02 U3720 ( .S(n808), .A0(n2192), .A1(n965), .Z(n964));
Q_AN02 U3721 ( .A0(n785), .A1(GFidata[491]), .Z(n963));
Q_MX02 U3722 ( .S(n808), .A0(n2191), .A1(n963), .Z(n962));
Q_AN02 U3723 ( .A0(n785), .A1(GFidata[492]), .Z(n961));
Q_MX02 U3724 ( .S(n808), .A0(n2190), .A1(n961), .Z(n960));
Q_AN02 U3725 ( .A0(n785), .A1(GFidata[493]), .Z(n959));
Q_MX02 U3726 ( .S(n808), .A0(n2189), .A1(n959), .Z(n958));
Q_AN02 U3727 ( .A0(n785), .A1(GFidata[494]), .Z(n957));
Q_MX02 U3728 ( .S(n808), .A0(n2188), .A1(n957), .Z(n956));
Q_AN02 U3729 ( .A0(n785), .A1(GFidata[495]), .Z(n955));
Q_MX02 U3730 ( .S(n808), .A0(n2187), .A1(n955), .Z(n954));
Q_AN02 U3731 ( .A0(n785), .A1(GFidata[496]), .Z(n953));
Q_MX02 U3732 ( .S(n808), .A0(n2186), .A1(n953), .Z(n952));
Q_AN02 U3733 ( .A0(n785), .A1(GFidata[497]), .Z(n951));
Q_MX02 U3734 ( .S(n808), .A0(n2185), .A1(n951), .Z(n950));
Q_AN02 U3735 ( .A0(n785), .A1(GFidata[498]), .Z(n949));
Q_MX02 U3736 ( .S(n808), .A0(n2184), .A1(n949), .Z(n948));
Q_AN02 U3737 ( .A0(n785), .A1(GFidata[499]), .Z(n947));
Q_MX02 U3738 ( .S(n808), .A0(n2183), .A1(n947), .Z(n946));
Q_AN02 U3739 ( .A0(n785), .A1(GFidata[500]), .Z(n945));
Q_MX02 U3740 ( .S(n808), .A0(n2182), .A1(n945), .Z(n944));
Q_AN02 U3741 ( .A0(n785), .A1(GFidata[501]), .Z(n943));
Q_MX02 U3742 ( .S(n808), .A0(n2181), .A1(n943), .Z(n942));
Q_AN02 U3743 ( .A0(n785), .A1(GFidata[502]), .Z(n941));
Q_MX02 U3744 ( .S(n808), .A0(n2180), .A1(n941), .Z(n940));
Q_AN02 U3745 ( .A0(n785), .A1(GFidata[503]), .Z(n939));
Q_MX02 U3746 ( .S(n808), .A0(n2179), .A1(n939), .Z(n938));
Q_AN02 U3747 ( .A0(n785), .A1(GFidata[504]), .Z(n937));
Q_MX02 U3748 ( .S(n808), .A0(n2178), .A1(n937), .Z(n936));
Q_AN02 U3749 ( .A0(n785), .A1(GFidata[505]), .Z(n935));
Q_MX02 U3750 ( .S(n808), .A0(n2177), .A1(n935), .Z(n934));
Q_AN02 U3751 ( .A0(n785), .A1(GFidata[506]), .Z(n933));
Q_MX02 U3752 ( .S(n808), .A0(n2176), .A1(n933), .Z(n932));
Q_AN02 U3753 ( .A0(n785), .A1(GFidata[507]), .Z(n931));
Q_MX02 U3754 ( .S(n808), .A0(n2175), .A1(n931), .Z(n930));
Q_AN02 U3755 ( .A0(n785), .A1(GFidata[508]), .Z(n929));
Q_MX02 U3756 ( .S(n808), .A0(n2174), .A1(n929), .Z(n928));
Q_AN02 U3757 ( .A0(n785), .A1(GFidata[509]), .Z(n927));
Q_MX02 U3758 ( .S(n808), .A0(n2173), .A1(n927), .Z(n926));
Q_AN02 U3759 ( .A0(n785), .A1(GFidata[510]), .Z(n925));
Q_MX02 U3760 ( .S(n808), .A0(n2172), .A1(n925), .Z(n924));
Q_AN02 U3761 ( .A0(n785), .A1(GFidata[511]), .Z(n923));
Q_MX02 U3762 ( .S(n808), .A0(n2171), .A1(n923), .Z(n922));
Q_FDP0UA U3763 ( .D(n890), .QTFCLK( ), .Q(xdata[543]));
Q_FDP0UA U3764 ( .D(n891), .QTFCLK( ), .Q(xdata[542]));
Q_FDP0UA U3765 ( .D(n892), .QTFCLK( ), .Q(xdata[541]));
Q_FDP0UA U3766 ( .D(n893), .QTFCLK( ), .Q(xdata[540]));
Q_FDP0UA U3767 ( .D(n894), .QTFCLK( ), .Q(xdata[539]));
Q_FDP0UA U3768 ( .D(n895), .QTFCLK( ), .Q(xdata[538]));
Q_FDP0UA U3769 ( .D(n896), .QTFCLK( ), .Q(xdata[537]));
Q_FDP0UA U3770 ( .D(n897), .QTFCLK( ), .Q(xdata[536]));
Q_FDP0UA U3771 ( .D(n898), .QTFCLK( ), .Q(xdata[535]));
Q_FDP0UA U3772 ( .D(n899), .QTFCLK( ), .Q(xdata[534]));
Q_FDP0UA U3773 ( .D(n900), .QTFCLK( ), .Q(xdata[533]));
Q_FDP0UA U3774 ( .D(n901), .QTFCLK( ), .Q(xdata[532]));
Q_FDP0UA U3775 ( .D(n902), .QTFCLK( ), .Q(xdata[531]));
Q_FDP0UA U3776 ( .D(n903), .QTFCLK( ), .Q(xdata[530]));
Q_FDP0UA U3777 ( .D(n904), .QTFCLK( ), .Q(xdata[529]));
Q_FDP0UA U3778 ( .D(n905), .QTFCLK( ), .Q(xdata[528]));
Q_FDP0UA U3779 ( .D(n906), .QTFCLK( ), .Q(xdata[527]));
Q_FDP0UA U3780 ( .D(n907), .QTFCLK( ), .Q(xdata[526]));
Q_FDP0UA U3781 ( .D(n908), .QTFCLK( ), .Q(xdata[525]));
Q_FDP0UA U3782 ( .D(n909), .QTFCLK( ), .Q(xdata[524]));
Q_FDP0UA U3783 ( .D(n910), .QTFCLK( ), .Q(xdata[523]));
Q_FDP0UA U3784 ( .D(n911), .QTFCLK( ), .Q(xdata[522]));
Q_FDP0UA U3785 ( .D(n912), .QTFCLK( ), .Q(xdata[521]));
Q_FDP0UA U3786 ( .D(n913), .QTFCLK( ), .Q(xdata[520]));
Q_FDP0UA U3787 ( .D(n914), .QTFCLK( ), .Q(xdata[519]));
Q_FDP0UA U3788 ( .D(n915), .QTFCLK( ), .Q(xdata[518]));
Q_FDP0UA U3789 ( .D(n916), .QTFCLK( ), .Q(xdata[517]));
Q_FDP0UA U3790 ( .D(n917), .QTFCLK( ), .Q(xdata[516]));
Q_FDP0UA U3791 ( .D(n918), .QTFCLK( ), .Q(xdata[515]));
Q_FDP0UA U3792 ( .D(n919), .QTFCLK( ), .Q(xdata[514]));
Q_FDP0UA U3793 ( .D(n920), .QTFCLK( ), .Q(xdata[513]));
Q_FDP0UA U3794 ( .D(n921), .QTFCLK( ), .Q(xdata[512]));
Q_FDP0UA U3795 ( .D(n922), .QTFCLK( ), .Q(xdata[511]));
Q_FDP0UA U3796 ( .D(n924), .QTFCLK( ), .Q(xdata[510]));
Q_FDP0UA U3797 ( .D(n926), .QTFCLK( ), .Q(xdata[509]));
Q_FDP0UA U3798 ( .D(n928), .QTFCLK( ), .Q(xdata[508]));
Q_FDP0UA U3799 ( .D(n930), .QTFCLK( ), .Q(xdata[507]));
Q_FDP0UA U3800 ( .D(n932), .QTFCLK( ), .Q(xdata[506]));
Q_FDP0UA U3801 ( .D(n934), .QTFCLK( ), .Q(xdata[505]));
Q_FDP0UA U3802 ( .D(n936), .QTFCLK( ), .Q(xdata[504]));
Q_FDP0UA U3803 ( .D(n938), .QTFCLK( ), .Q(xdata[503]));
Q_FDP0UA U3804 ( .D(n940), .QTFCLK( ), .Q(xdata[502]));
Q_FDP0UA U3805 ( .D(n942), .QTFCLK( ), .Q(xdata[501]));
Q_FDP0UA U3806 ( .D(n944), .QTFCLK( ), .Q(xdata[500]));
Q_FDP0UA U3807 ( .D(n946), .QTFCLK( ), .Q(xdata[499]));
Q_FDP0UA U3808 ( .D(n948), .QTFCLK( ), .Q(xdata[498]));
Q_FDP0UA U3809 ( .D(n950), .QTFCLK( ), .Q(xdata[497]));
Q_FDP0UA U3810 ( .D(n952), .QTFCLK( ), .Q(xdata[496]));
Q_FDP0UA U3811 ( .D(n954), .QTFCLK( ), .Q(xdata[495]));
Q_FDP0UA U3812 ( .D(n956), .QTFCLK( ), .Q(xdata[494]));
Q_FDP0UA U3813 ( .D(n958), .QTFCLK( ), .Q(xdata[493]));
Q_FDP0UA U3814 ( .D(n960), .QTFCLK( ), .Q(xdata[492]));
Q_FDP0UA U3815 ( .D(n962), .QTFCLK( ), .Q(xdata[491]));
Q_FDP0UA U3816 ( .D(n964), .QTFCLK( ), .Q(xdata[490]));
Q_FDP0UA U3817 ( .D(n966), .QTFCLK( ), .Q(xdata[489]));
Q_FDP0UA U3818 ( .D(n968), .QTFCLK( ), .Q(xdata[488]));
Q_FDP0UA U3819 ( .D(n970), .QTFCLK( ), .Q(xdata[487]));
Q_FDP0UA U3820 ( .D(n972), .QTFCLK( ), .Q(xdata[486]));
Q_FDP0UA U3821 ( .D(n974), .QTFCLK( ), .Q(xdata[485]));
Q_FDP0UA U3822 ( .D(n976), .QTFCLK( ), .Q(xdata[484]));
Q_FDP0UA U3823 ( .D(n978), .QTFCLK( ), .Q(xdata[483]));
Q_FDP0UA U3824 ( .D(n980), .QTFCLK( ), .Q(xdata[482]));
Q_FDP0UA U3825 ( .D(n982), .QTFCLK( ), .Q(xdata[481]));
Q_FDP0UA U3826 ( .D(n984), .QTFCLK( ), .Q(xdata[480]));
Q_FDP0UA U3827 ( .D(n986), .QTFCLK( ), .Q(xdata[479]));
Q_FDP0UA U3828 ( .D(n988), .QTFCLK( ), .Q(xdata[478]));
Q_FDP0UA U3829 ( .D(n990), .QTFCLK( ), .Q(xdata[477]));
Q_FDP0UA U3830 ( .D(n992), .QTFCLK( ), .Q(xdata[476]));
Q_FDP0UA U3831 ( .D(n994), .QTFCLK( ), .Q(xdata[475]));
Q_FDP0UA U3832 ( .D(n996), .QTFCLK( ), .Q(xdata[474]));
Q_FDP0UA U3833 ( .D(n998), .QTFCLK( ), .Q(xdata[473]));
Q_FDP0UA U3834 ( .D(n1000), .QTFCLK( ), .Q(xdata[472]));
Q_FDP0UA U3835 ( .D(n1002), .QTFCLK( ), .Q(xdata[471]));
Q_FDP0UA U3836 ( .D(n1004), .QTFCLK( ), .Q(xdata[470]));
Q_FDP0UA U3837 ( .D(n1006), .QTFCLK( ), .Q(xdata[469]));
Q_FDP0UA U3838 ( .D(n1008), .QTFCLK( ), .Q(xdata[468]));
Q_FDP0UA U3839 ( .D(n1010), .QTFCLK( ), .Q(xdata[467]));
Q_FDP0UA U3840 ( .D(n1012), .QTFCLK( ), .Q(xdata[466]));
Q_FDP0UA U3841 ( .D(n1014), .QTFCLK( ), .Q(xdata[465]));
Q_FDP0UA U3842 ( .D(n1016), .QTFCLK( ), .Q(xdata[464]));
Q_FDP0UA U3843 ( .D(n1018), .QTFCLK( ), .Q(xdata[463]));
Q_FDP0UA U3844 ( .D(n1020), .QTFCLK( ), .Q(xdata[462]));
Q_FDP0UA U3845 ( .D(n1022), .QTFCLK( ), .Q(xdata[461]));
Q_FDP0UA U3846 ( .D(n1024), .QTFCLK( ), .Q(xdata[460]));
Q_FDP0UA U3847 ( .D(n1026), .QTFCLK( ), .Q(xdata[459]));
Q_FDP0UA U3848 ( .D(n1028), .QTFCLK( ), .Q(xdata[458]));
Q_FDP0UA U3849 ( .D(n1030), .QTFCLK( ), .Q(xdata[457]));
Q_FDP0UA U3850 ( .D(n1032), .QTFCLK( ), .Q(xdata[456]));
Q_FDP0UA U3851 ( .D(n1034), .QTFCLK( ), .Q(xdata[455]));
Q_FDP0UA U3852 ( .D(n1036), .QTFCLK( ), .Q(xdata[454]));
Q_FDP0UA U3853 ( .D(n1038), .QTFCLK( ), .Q(xdata[453]));
Q_FDP0UA U3854 ( .D(n1040), .QTFCLK( ), .Q(xdata[452]));
Q_FDP0UA U3855 ( .D(n1042), .QTFCLK( ), .Q(xdata[451]));
Q_FDP0UA U3856 ( .D(n1044), .QTFCLK( ), .Q(xdata[450]));
Q_FDP0UA U3857 ( .D(n1046), .QTFCLK( ), .Q(xdata[449]));
Q_FDP0UA U3858 ( .D(n1048), .QTFCLK( ), .Q(xdata[448]));
Q_FDP0UA U3859 ( .D(n1050), .QTFCLK( ), .Q(xdata[447]));
Q_FDP0UA U3860 ( .D(n1052), .QTFCLK( ), .Q(xdata[446]));
Q_FDP0UA U3861 ( .D(n1054), .QTFCLK( ), .Q(xdata[445]));
Q_FDP0UA U3862 ( .D(n1056), .QTFCLK( ), .Q(xdata[444]));
Q_FDP0UA U3863 ( .D(n1058), .QTFCLK( ), .Q(xdata[443]));
Q_FDP0UA U3864 ( .D(n1060), .QTFCLK( ), .Q(xdata[442]));
Q_FDP0UA U3865 ( .D(n1062), .QTFCLK( ), .Q(xdata[441]));
Q_FDP0UA U3866 ( .D(n1064), .QTFCLK( ), .Q(xdata[440]));
Q_FDP0UA U3867 ( .D(n1066), .QTFCLK( ), .Q(xdata[439]));
Q_FDP0UA U3868 ( .D(n1068), .QTFCLK( ), .Q(xdata[438]));
Q_FDP0UA U3869 ( .D(n1070), .QTFCLK( ), .Q(xdata[437]));
Q_FDP0UA U3870 ( .D(n1072), .QTFCLK( ), .Q(xdata[436]));
Q_FDP0UA U3871 ( .D(n1074), .QTFCLK( ), .Q(xdata[435]));
Q_FDP0UA U3872 ( .D(n1076), .QTFCLK( ), .Q(xdata[434]));
Q_FDP0UA U3873 ( .D(n1078), .QTFCLK( ), .Q(xdata[433]));
Q_FDP0UA U3874 ( .D(n1080), .QTFCLK( ), .Q(xdata[432]));
Q_FDP0UA U3875 ( .D(n1082), .QTFCLK( ), .Q(xdata[431]));
Q_FDP0UA U3876 ( .D(n1084), .QTFCLK( ), .Q(xdata[430]));
Q_FDP0UA U3877 ( .D(n1086), .QTFCLK( ), .Q(xdata[429]));
Q_FDP0UA U3878 ( .D(n1088), .QTFCLK( ), .Q(xdata[428]));
Q_FDP0UA U3879 ( .D(n1090), .QTFCLK( ), .Q(xdata[427]));
Q_FDP0UA U3880 ( .D(n1092), .QTFCLK( ), .Q(xdata[426]));
Q_FDP0UA U3881 ( .D(n1094), .QTFCLK( ), .Q(xdata[425]));
Q_FDP0UA U3882 ( .D(n1096), .QTFCLK( ), .Q(xdata[424]));
Q_FDP0UA U3883 ( .D(n1098), .QTFCLK( ), .Q(xdata[423]));
Q_FDP0UA U3884 ( .D(n1100), .QTFCLK( ), .Q(xdata[422]));
Q_FDP0UA U3885 ( .D(n1102), .QTFCLK( ), .Q(xdata[421]));
Q_FDP0UA U3886 ( .D(n1104), .QTFCLK( ), .Q(xdata[420]));
Q_FDP0UA U3887 ( .D(n1106), .QTFCLK( ), .Q(xdata[419]));
Q_FDP0UA U3888 ( .D(n1108), .QTFCLK( ), .Q(xdata[418]));
Q_FDP0UA U3889 ( .D(n1110), .QTFCLK( ), .Q(xdata[417]));
Q_FDP0UA U3890 ( .D(n1112), .QTFCLK( ), .Q(xdata[416]));
Q_FDP0UA U3891 ( .D(n1114), .QTFCLK( ), .Q(xdata[415]));
Q_FDP0UA U3892 ( .D(n1116), .QTFCLK( ), .Q(xdata[414]));
Q_FDP0UA U3893 ( .D(n1118), .QTFCLK( ), .Q(xdata[413]));
Q_FDP0UA U3894 ( .D(n1120), .QTFCLK( ), .Q(xdata[412]));
Q_FDP0UA U3895 ( .D(n1122), .QTFCLK( ), .Q(xdata[411]));
Q_FDP0UA U3896 ( .D(n1124), .QTFCLK( ), .Q(xdata[410]));
Q_FDP0UA U3897 ( .D(n1126), .QTFCLK( ), .Q(xdata[409]));
Q_FDP0UA U3898 ( .D(n1128), .QTFCLK( ), .Q(xdata[408]));
Q_FDP0UA U3899 ( .D(n1130), .QTFCLK( ), .Q(xdata[407]));
Q_FDP0UA U3900 ( .D(n1132), .QTFCLK( ), .Q(xdata[406]));
Q_FDP0UA U3901 ( .D(n1134), .QTFCLK( ), .Q(xdata[405]));
Q_FDP0UA U3902 ( .D(n1136), .QTFCLK( ), .Q(xdata[404]));
Q_FDP0UA U3903 ( .D(n1138), .QTFCLK( ), .Q(xdata[403]));
Q_FDP0UA U3904 ( .D(n1140), .QTFCLK( ), .Q(xdata[402]));
Q_FDP0UA U3905 ( .D(n1142), .QTFCLK( ), .Q(xdata[401]));
Q_FDP0UA U3906 ( .D(n1144), .QTFCLK( ), .Q(xdata[400]));
Q_FDP0UA U3907 ( .D(n1146), .QTFCLK( ), .Q(xdata[399]));
Q_FDP0UA U3908 ( .D(n1148), .QTFCLK( ), .Q(xdata[398]));
Q_FDP0UA U3909 ( .D(n1150), .QTFCLK( ), .Q(xdata[397]));
Q_FDP0UA U3910 ( .D(n1152), .QTFCLK( ), .Q(xdata[396]));
Q_FDP0UA U3911 ( .D(n1154), .QTFCLK( ), .Q(xdata[395]));
Q_FDP0UA U3912 ( .D(n1156), .QTFCLK( ), .Q(xdata[394]));
Q_FDP0UA U3913 ( .D(n1158), .QTFCLK( ), .Q(xdata[393]));
Q_FDP0UA U3914 ( .D(n1160), .QTFCLK( ), .Q(xdata[392]));
Q_FDP0UA U3915 ( .D(n1162), .QTFCLK( ), .Q(xdata[391]));
Q_FDP0UA U3916 ( .D(n1164), .QTFCLK( ), .Q(xdata[390]));
Q_FDP0UA U3917 ( .D(n1166), .QTFCLK( ), .Q(xdata[389]));
Q_FDP0UA U3918 ( .D(n1168), .QTFCLK( ), .Q(xdata[388]));
Q_FDP0UA U3919 ( .D(n1170), .QTFCLK( ), .Q(xdata[387]));
Q_FDP0UA U3920 ( .D(n1172), .QTFCLK( ), .Q(xdata[386]));
Q_FDP0UA U3921 ( .D(n1174), .QTFCLK( ), .Q(xdata[385]));
Q_FDP0UA U3922 ( .D(n1176), .QTFCLK( ), .Q(xdata[384]));
Q_FDP0UA U3923 ( .D(n1178), .QTFCLK( ), .Q(xdata[383]));
Q_FDP0UA U3924 ( .D(n1180), .QTFCLK( ), .Q(xdata[382]));
Q_FDP0UA U3925 ( .D(n1182), .QTFCLK( ), .Q(xdata[381]));
Q_FDP0UA U3926 ( .D(n1184), .QTFCLK( ), .Q(xdata[380]));
Q_FDP0UA U3927 ( .D(n1186), .QTFCLK( ), .Q(xdata[379]));
Q_FDP0UA U3928 ( .D(n1188), .QTFCLK( ), .Q(xdata[378]));
Q_FDP0UA U3929 ( .D(n1190), .QTFCLK( ), .Q(xdata[377]));
Q_FDP0UA U3930 ( .D(n1192), .QTFCLK( ), .Q(xdata[376]));
Q_FDP0UA U3931 ( .D(n1194), .QTFCLK( ), .Q(xdata[375]));
Q_FDP0UA U3932 ( .D(n1196), .QTFCLK( ), .Q(xdata[374]));
Q_FDP0UA U3933 ( .D(n1198), .QTFCLK( ), .Q(xdata[373]));
Q_FDP0UA U3934 ( .D(n1200), .QTFCLK( ), .Q(xdata[372]));
Q_FDP0UA U3935 ( .D(n1202), .QTFCLK( ), .Q(xdata[371]));
Q_FDP0UA U3936 ( .D(n1204), .QTFCLK( ), .Q(xdata[370]));
Q_FDP0UA U3937 ( .D(n1206), .QTFCLK( ), .Q(xdata[369]));
Q_FDP0UA U3938 ( .D(n1208), .QTFCLK( ), .Q(xdata[368]));
Q_FDP0UA U3939 ( .D(n1210), .QTFCLK( ), .Q(xdata[367]));
Q_FDP0UA U3940 ( .D(n1212), .QTFCLK( ), .Q(xdata[366]));
Q_FDP0UA U3941 ( .D(n1214), .QTFCLK( ), .Q(xdata[365]));
Q_FDP0UA U3942 ( .D(n1216), .QTFCLK( ), .Q(xdata[364]));
Q_FDP0UA U3943 ( .D(n1218), .QTFCLK( ), .Q(xdata[363]));
Q_FDP0UA U3944 ( .D(n1220), .QTFCLK( ), .Q(xdata[362]));
Q_FDP0UA U3945 ( .D(n1222), .QTFCLK( ), .Q(xdata[361]));
Q_FDP0UA U3946 ( .D(n1224), .QTFCLK( ), .Q(xdata[360]));
Q_FDP0UA U3947 ( .D(n1226), .QTFCLK( ), .Q(xdata[359]));
Q_FDP0UA U3948 ( .D(n1228), .QTFCLK( ), .Q(xdata[358]));
Q_FDP0UA U3949 ( .D(n1230), .QTFCLK( ), .Q(xdata[357]));
Q_FDP0UA U3950 ( .D(n1232), .QTFCLK( ), .Q(xdata[356]));
Q_FDP0UA U3951 ( .D(n1234), .QTFCLK( ), .Q(xdata[355]));
Q_FDP0UA U3952 ( .D(n1236), .QTFCLK( ), .Q(xdata[354]));
Q_FDP0UA U3953 ( .D(n1238), .QTFCLK( ), .Q(xdata[353]));
Q_FDP0UA U3954 ( .D(n1240), .QTFCLK( ), .Q(xdata[352]));
Q_FDP0UA U3955 ( .D(n1242), .QTFCLK( ), .Q(xdata[351]));
Q_FDP0UA U3956 ( .D(n1244), .QTFCLK( ), .Q(xdata[350]));
Q_FDP0UA U3957 ( .D(n1246), .QTFCLK( ), .Q(xdata[349]));
Q_FDP0UA U3958 ( .D(n1248), .QTFCLK( ), .Q(xdata[348]));
Q_FDP0UA U3959 ( .D(n1250), .QTFCLK( ), .Q(xdata[347]));
Q_FDP0UA U3960 ( .D(n1252), .QTFCLK( ), .Q(xdata[346]));
Q_FDP0UA U3961 ( .D(n1254), .QTFCLK( ), .Q(xdata[345]));
Q_FDP0UA U3962 ( .D(n1256), .QTFCLK( ), .Q(xdata[344]));
Q_FDP0UA U3963 ( .D(n1258), .QTFCLK( ), .Q(xdata[343]));
Q_FDP0UA U3964 ( .D(n1260), .QTFCLK( ), .Q(xdata[342]));
Q_FDP0UA U3965 ( .D(n1262), .QTFCLK( ), .Q(xdata[341]));
Q_FDP0UA U3966 ( .D(n1264), .QTFCLK( ), .Q(xdata[340]));
Q_FDP0UA U3967 ( .D(n1266), .QTFCLK( ), .Q(xdata[339]));
Q_FDP0UA U3968 ( .D(n1268), .QTFCLK( ), .Q(xdata[338]));
Q_FDP0UA U3969 ( .D(n1270), .QTFCLK( ), .Q(xdata[337]));
Q_FDP0UA U3970 ( .D(n1272), .QTFCLK( ), .Q(xdata[336]));
Q_FDP0UA U3971 ( .D(n1274), .QTFCLK( ), .Q(xdata[335]));
Q_FDP0UA U3972 ( .D(n1276), .QTFCLK( ), .Q(xdata[334]));
Q_FDP0UA U3973 ( .D(n1278), .QTFCLK( ), .Q(xdata[333]));
Q_FDP0UA U3974 ( .D(n1280), .QTFCLK( ), .Q(xdata[332]));
Q_FDP0UA U3975 ( .D(n1282), .QTFCLK( ), .Q(xdata[331]));
Q_FDP0UA U3976 ( .D(n1284), .QTFCLK( ), .Q(xdata[330]));
Q_FDP0UA U3977 ( .D(n1286), .QTFCLK( ), .Q(xdata[329]));
Q_FDP0UA U3978 ( .D(n1288), .QTFCLK( ), .Q(xdata[328]));
Q_FDP0UA U3979 ( .D(n1290), .QTFCLK( ), .Q(xdata[327]));
Q_FDP0UA U3980 ( .D(n1292), .QTFCLK( ), .Q(xdata[326]));
Q_FDP0UA U3981 ( .D(n1294), .QTFCLK( ), .Q(xdata[325]));
Q_FDP0UA U3982 ( .D(n1296), .QTFCLK( ), .Q(xdata[324]));
Q_FDP0UA U3983 ( .D(n1298), .QTFCLK( ), .Q(xdata[323]));
Q_FDP0UA U3984 ( .D(n1300), .QTFCLK( ), .Q(xdata[322]));
Q_FDP0UA U3985 ( .D(n1302), .QTFCLK( ), .Q(xdata[321]));
Q_FDP0UA U3986 ( .D(n1304), .QTFCLK( ), .Q(xdata[320]));
Q_FDP0UA U3987 ( .D(n1306), .QTFCLK( ), .Q(xdata[319]));
Q_FDP0UA U3988 ( .D(n1308), .QTFCLK( ), .Q(xdata[318]));
Q_FDP0UA U3989 ( .D(n1310), .QTFCLK( ), .Q(xdata[317]));
Q_FDP0UA U3990 ( .D(n1312), .QTFCLK( ), .Q(xdata[316]));
Q_FDP0UA U3991 ( .D(n1314), .QTFCLK( ), .Q(xdata[315]));
Q_FDP0UA U3992 ( .D(n1316), .QTFCLK( ), .Q(xdata[314]));
Q_FDP0UA U3993 ( .D(n1318), .QTFCLK( ), .Q(xdata[313]));
Q_FDP0UA U3994 ( .D(n1320), .QTFCLK( ), .Q(xdata[312]));
Q_FDP0UA U3995 ( .D(n1322), .QTFCLK( ), .Q(xdata[311]));
Q_FDP0UA U3996 ( .D(n1324), .QTFCLK( ), .Q(xdata[310]));
Q_FDP0UA U3997 ( .D(n1326), .QTFCLK( ), .Q(xdata[309]));
Q_FDP0UA U3998 ( .D(n1328), .QTFCLK( ), .Q(xdata[308]));
Q_FDP0UA U3999 ( .D(n1330), .QTFCLK( ), .Q(xdata[307]));
Q_FDP0UA U4000 ( .D(n1332), .QTFCLK( ), .Q(xdata[306]));
Q_FDP0UA U4001 ( .D(n1334), .QTFCLK( ), .Q(xdata[305]));
Q_FDP0UA U4002 ( .D(n1336), .QTFCLK( ), .Q(xdata[304]));
Q_FDP0UA U4003 ( .D(n1338), .QTFCLK( ), .Q(xdata[303]));
Q_FDP0UA U4004 ( .D(n1340), .QTFCLK( ), .Q(xdata[302]));
Q_FDP0UA U4005 ( .D(n1342), .QTFCLK( ), .Q(xdata[301]));
Q_FDP0UA U4006 ( .D(n1344), .QTFCLK( ), .Q(xdata[300]));
Q_FDP0UA U4007 ( .D(n1346), .QTFCLK( ), .Q(xdata[299]));
Q_FDP0UA U4008 ( .D(n1348), .QTFCLK( ), .Q(xdata[298]));
Q_FDP0UA U4009 ( .D(n1350), .QTFCLK( ), .Q(xdata[297]));
Q_FDP0UA U4010 ( .D(n1352), .QTFCLK( ), .Q(xdata[296]));
Q_FDP0UA U4011 ( .D(n1354), .QTFCLK( ), .Q(xdata[295]));
Q_FDP0UA U4012 ( .D(n1356), .QTFCLK( ), .Q(xdata[294]));
Q_FDP0UA U4013 ( .D(n1358), .QTFCLK( ), .Q(xdata[293]));
Q_FDP0UA U4014 ( .D(n1360), .QTFCLK( ), .Q(xdata[292]));
Q_FDP0UA U4015 ( .D(n1362), .QTFCLK( ), .Q(xdata[291]));
Q_FDP0UA U4016 ( .D(n1364), .QTFCLK( ), .Q(xdata[290]));
Q_FDP0UA U4017 ( .D(n1366), .QTFCLK( ), .Q(xdata[289]));
Q_FDP0UA U4018 ( .D(n1368), .QTFCLK( ), .Q(xdata[288]));
Q_FDP0UA U4019 ( .D(n1370), .QTFCLK( ), .Q(xdata[287]));
Q_FDP0UA U4020 ( .D(n1372), .QTFCLK( ), .Q(xdata[286]));
Q_FDP0UA U4021 ( .D(n1374), .QTFCLK( ), .Q(xdata[285]));
Q_FDP0UA U4022 ( .D(n1376), .QTFCLK( ), .Q(xdata[284]));
Q_FDP0UA U4023 ( .D(n1378), .QTFCLK( ), .Q(xdata[283]));
Q_FDP0UA U4024 ( .D(n1380), .QTFCLK( ), .Q(xdata[282]));
Q_FDP0UA U4025 ( .D(n1382), .QTFCLK( ), .Q(xdata[281]));
Q_FDP0UA U4026 ( .D(n1384), .QTFCLK( ), .Q(xdata[280]));
Q_FDP0UA U4027 ( .D(n1386), .QTFCLK( ), .Q(xdata[279]));
Q_FDP0UA U4028 ( .D(n1388), .QTFCLK( ), .Q(xdata[278]));
Q_FDP0UA U4029 ( .D(n1390), .QTFCLK( ), .Q(xdata[277]));
Q_FDP0UA U4030 ( .D(n1392), .QTFCLK( ), .Q(xdata[276]));
Q_FDP0UA U4031 ( .D(n1394), .QTFCLK( ), .Q(xdata[275]));
Q_FDP0UA U4032 ( .D(n1396), .QTFCLK( ), .Q(xdata[274]));
Q_FDP0UA U4033 ( .D(n1398), .QTFCLK( ), .Q(xdata[273]));
Q_FDP0UA U4034 ( .D(n1400), .QTFCLK( ), .Q(xdata[272]));
Q_FDP0UA U4035 ( .D(n1402), .QTFCLK( ), .Q(xdata[271]));
Q_FDP0UA U4036 ( .D(n1404), .QTFCLK( ), .Q(xdata[270]));
Q_FDP0UA U4037 ( .D(n1406), .QTFCLK( ), .Q(xdata[269]));
Q_FDP0UA U4038 ( .D(n1408), .QTFCLK( ), .Q(xdata[268]));
Q_FDP0UA U4039 ( .D(n1410), .QTFCLK( ), .Q(xdata[267]));
Q_FDP0UA U4040 ( .D(n1412), .QTFCLK( ), .Q(xdata[266]));
Q_FDP0UA U4041 ( .D(n1414), .QTFCLK( ), .Q(xdata[265]));
Q_FDP0UA U4042 ( .D(n1416), .QTFCLK( ), .Q(xdata[264]));
Q_FDP0UA U4043 ( .D(n1418), .QTFCLK( ), .Q(xdata[263]));
Q_FDP0UA U4044 ( .D(n1420), .QTFCLK( ), .Q(xdata[262]));
Q_FDP0UA U4045 ( .D(n1422), .QTFCLK( ), .Q(xdata[261]));
Q_FDP0UA U4046 ( .D(n1424), .QTFCLK( ), .Q(xdata[260]));
Q_FDP0UA U4047 ( .D(n1426), .QTFCLK( ), .Q(xdata[259]));
Q_FDP0UA U4048 ( .D(n1428), .QTFCLK( ), .Q(xdata[258]));
Q_FDP0UA U4049 ( .D(n1430), .QTFCLK( ), .Q(xdata[257]));
Q_FDP0UA U4050 ( .D(n1432), .QTFCLK( ), .Q(xdata[256]));
Q_FDP0UA U4051 ( .D(n1434), .QTFCLK( ), .Q(xdata[255]));
Q_FDP0UA U4052 ( .D(n1436), .QTFCLK( ), .Q(xdata[254]));
Q_FDP0UA U4053 ( .D(n1438), .QTFCLK( ), .Q(xdata[253]));
Q_FDP0UA U4054 ( .D(n1440), .QTFCLK( ), .Q(xdata[252]));
Q_FDP0UA U4055 ( .D(n1442), .QTFCLK( ), .Q(xdata[251]));
Q_FDP0UA U4056 ( .D(n1444), .QTFCLK( ), .Q(xdata[250]));
Q_FDP0UA U4057 ( .D(n1446), .QTFCLK( ), .Q(xdata[249]));
Q_FDP0UA U4058 ( .D(n1448), .QTFCLK( ), .Q(xdata[248]));
Q_FDP0UA U4059 ( .D(n1450), .QTFCLK( ), .Q(xdata[247]));
Q_FDP0UA U4060 ( .D(n1452), .QTFCLK( ), .Q(xdata[246]));
Q_FDP0UA U4061 ( .D(n1454), .QTFCLK( ), .Q(xdata[245]));
Q_FDP0UA U4062 ( .D(n1456), .QTFCLK( ), .Q(xdata[244]));
Q_FDP0UA U4063 ( .D(n1458), .QTFCLK( ), .Q(xdata[243]));
Q_FDP0UA U4064 ( .D(n1460), .QTFCLK( ), .Q(xdata[242]));
Q_FDP0UA U4065 ( .D(n1462), .QTFCLK( ), .Q(xdata[241]));
Q_FDP0UA U4066 ( .D(n1464), .QTFCLK( ), .Q(xdata[240]));
Q_FDP0UA U4067 ( .D(n1466), .QTFCLK( ), .Q(xdata[239]));
Q_FDP0UA U4068 ( .D(n1468), .QTFCLK( ), .Q(xdata[238]));
Q_FDP0UA U4069 ( .D(n1470), .QTFCLK( ), .Q(xdata[237]));
Q_FDP0UA U4070 ( .D(n1472), .QTFCLK( ), .Q(xdata[236]));
Q_FDP0UA U4071 ( .D(n1474), .QTFCLK( ), .Q(xdata[235]));
Q_FDP0UA U4072 ( .D(n1476), .QTFCLK( ), .Q(xdata[234]));
Q_FDP0UA U4073 ( .D(n1478), .QTFCLK( ), .Q(xdata[233]));
Q_FDP0UA U4074 ( .D(n1480), .QTFCLK( ), .Q(xdata[232]));
Q_FDP0UA U4075 ( .D(n1482), .QTFCLK( ), .Q(xdata[231]));
Q_FDP0UA U4076 ( .D(n1484), .QTFCLK( ), .Q(xdata[230]));
Q_FDP0UA U4077 ( .D(n1486), .QTFCLK( ), .Q(xdata[229]));
Q_FDP0UA U4078 ( .D(n1488), .QTFCLK( ), .Q(xdata[228]));
Q_FDP0UA U4079 ( .D(n1490), .QTFCLK( ), .Q(xdata[227]));
Q_FDP0UA U4080 ( .D(n1492), .QTFCLK( ), .Q(xdata[226]));
Q_FDP0UA U4081 ( .D(n1494), .QTFCLK( ), .Q(xdata[225]));
Q_FDP0UA U4082 ( .D(n1496), .QTFCLK( ), .Q(xdata[224]));
Q_FDP0UA U4083 ( .D(n1498), .QTFCLK( ), .Q(xdata[223]));
Q_FDP0UA U4084 ( .D(n1500), .QTFCLK( ), .Q(xdata[222]));
Q_FDP0UA U4085 ( .D(n1502), .QTFCLK( ), .Q(xdata[221]));
Q_FDP0UA U4086 ( .D(n1504), .QTFCLK( ), .Q(xdata[220]));
Q_FDP0UA U4087 ( .D(n1506), .QTFCLK( ), .Q(xdata[219]));
Q_FDP0UA U4088 ( .D(n1508), .QTFCLK( ), .Q(xdata[218]));
Q_FDP0UA U4089 ( .D(n1510), .QTFCLK( ), .Q(xdata[217]));
Q_FDP0UA U4090 ( .D(n1512), .QTFCLK( ), .Q(xdata[216]));
Q_FDP0UA U4091 ( .D(n1514), .QTFCLK( ), .Q(xdata[215]));
Q_FDP0UA U4092 ( .D(n1516), .QTFCLK( ), .Q(xdata[214]));
Q_FDP0UA U4093 ( .D(n1518), .QTFCLK( ), .Q(xdata[213]));
Q_FDP0UA U4094 ( .D(n1520), .QTFCLK( ), .Q(xdata[212]));
Q_FDP0UA U4095 ( .D(n1522), .QTFCLK( ), .Q(xdata[211]));
Q_FDP0UA U4096 ( .D(n1524), .QTFCLK( ), .Q(xdata[210]));
Q_FDP0UA U4097 ( .D(n1526), .QTFCLK( ), .Q(xdata[209]));
Q_FDP0UA U4098 ( .D(n1528), .QTFCLK( ), .Q(xdata[208]));
Q_FDP0UA U4099 ( .D(n1530), .QTFCLK( ), .Q(xdata[207]));
Q_FDP0UA U4100 ( .D(n1532), .QTFCLK( ), .Q(xdata[206]));
Q_FDP0UA U4101 ( .D(n1534), .QTFCLK( ), .Q(xdata[205]));
Q_FDP0UA U4102 ( .D(n1536), .QTFCLK( ), .Q(xdata[204]));
Q_FDP0UA U4103 ( .D(n1538), .QTFCLK( ), .Q(xdata[203]));
Q_FDP0UA U4104 ( .D(n1540), .QTFCLK( ), .Q(xdata[202]));
Q_FDP0UA U4105 ( .D(n1542), .QTFCLK( ), .Q(xdata[201]));
Q_FDP0UA U4106 ( .D(n1544), .QTFCLK( ), .Q(xdata[200]));
Q_FDP0UA U4107 ( .D(n1546), .QTFCLK( ), .Q(xdata[199]));
Q_FDP0UA U4108 ( .D(n1548), .QTFCLK( ), .Q(xdata[198]));
Q_FDP0UA U4109 ( .D(n1550), .QTFCLK( ), .Q(xdata[197]));
Q_FDP0UA U4110 ( .D(n1552), .QTFCLK( ), .Q(xdata[196]));
Q_FDP0UA U4111 ( .D(n1554), .QTFCLK( ), .Q(xdata[195]));
Q_FDP0UA U4112 ( .D(n1556), .QTFCLK( ), .Q(xdata[194]));
Q_FDP0UA U4113 ( .D(n1558), .QTFCLK( ), .Q(xdata[193]));
Q_FDP0UA U4114 ( .D(n1560), .QTFCLK( ), .Q(xdata[192]));
Q_FDP0UA U4115 ( .D(n1562), .QTFCLK( ), .Q(xdata[191]));
Q_FDP0UA U4116 ( .D(n1564), .QTFCLK( ), .Q(xdata[190]));
Q_FDP0UA U4117 ( .D(n1566), .QTFCLK( ), .Q(xdata[189]));
Q_FDP0UA U4118 ( .D(n1568), .QTFCLK( ), .Q(xdata[188]));
Q_FDP0UA U4119 ( .D(n1570), .QTFCLK( ), .Q(xdata[187]));
Q_FDP0UA U4120 ( .D(n1572), .QTFCLK( ), .Q(xdata[186]));
Q_FDP0UA U4121 ( .D(n1574), .QTFCLK( ), .Q(xdata[185]));
Q_FDP0UA U4122 ( .D(n1576), .QTFCLK( ), .Q(xdata[184]));
Q_FDP0UA U4123 ( .D(n1578), .QTFCLK( ), .Q(xdata[183]));
Q_FDP0UA U4124 ( .D(n1580), .QTFCLK( ), .Q(xdata[182]));
Q_FDP0UA U4125 ( .D(n1582), .QTFCLK( ), .Q(xdata[181]));
Q_FDP0UA U4126 ( .D(n1584), .QTFCLK( ), .Q(xdata[180]));
Q_FDP0UA U4127 ( .D(n1586), .QTFCLK( ), .Q(xdata[179]));
Q_FDP0UA U4128 ( .D(n1588), .QTFCLK( ), .Q(xdata[178]));
Q_FDP0UA U4129 ( .D(n1590), .QTFCLK( ), .Q(xdata[177]));
Q_FDP0UA U4130 ( .D(n1592), .QTFCLK( ), .Q(xdata[176]));
Q_FDP0UA U4131 ( .D(n1594), .QTFCLK( ), .Q(xdata[175]));
Q_FDP0UA U4132 ( .D(n1596), .QTFCLK( ), .Q(xdata[174]));
Q_FDP0UA U4133 ( .D(n1598), .QTFCLK( ), .Q(xdata[173]));
Q_FDP0UA U4134 ( .D(n1600), .QTFCLK( ), .Q(xdata[172]));
Q_FDP0UA U4135 ( .D(n1602), .QTFCLK( ), .Q(xdata[171]));
Q_FDP0UA U4136 ( .D(n1604), .QTFCLK( ), .Q(xdata[170]));
Q_FDP0UA U4137 ( .D(n1606), .QTFCLK( ), .Q(xdata[169]));
Q_FDP0UA U4138 ( .D(n1608), .QTFCLK( ), .Q(xdata[168]));
Q_FDP0UA U4139 ( .D(n1610), .QTFCLK( ), .Q(xdata[167]));
Q_FDP0UA U4140 ( .D(n1612), .QTFCLK( ), .Q(xdata[166]));
Q_FDP0UA U4141 ( .D(n1614), .QTFCLK( ), .Q(xdata[165]));
Q_FDP0UA U4142 ( .D(n1616), .QTFCLK( ), .Q(xdata[164]));
Q_FDP0UA U4143 ( .D(n1618), .QTFCLK( ), .Q(xdata[163]));
Q_FDP0UA U4144 ( .D(n1620), .QTFCLK( ), .Q(xdata[162]));
Q_FDP0UA U4145 ( .D(n1622), .QTFCLK( ), .Q(xdata[161]));
Q_FDP0UA U4146 ( .D(n1624), .QTFCLK( ), .Q(xdata[160]));
Q_FDP0UA U4147 ( .D(n1626), .QTFCLK( ), .Q(xdata[159]));
Q_FDP0UA U4148 ( .D(n1628), .QTFCLK( ), .Q(xdata[158]));
Q_FDP0UA U4149 ( .D(n1630), .QTFCLK( ), .Q(xdata[157]));
Q_FDP0UA U4150 ( .D(n1632), .QTFCLK( ), .Q(xdata[156]));
Q_FDP0UA U4151 ( .D(n1634), .QTFCLK( ), .Q(xdata[155]));
Q_FDP0UA U4152 ( .D(n1636), .QTFCLK( ), .Q(xdata[154]));
Q_FDP0UA U4153 ( .D(n1638), .QTFCLK( ), .Q(xdata[153]));
Q_FDP0UA U4154 ( .D(n1640), .QTFCLK( ), .Q(xdata[152]));
Q_FDP0UA U4155 ( .D(n1642), .QTFCLK( ), .Q(xdata[151]));
Q_FDP0UA U4156 ( .D(n1644), .QTFCLK( ), .Q(xdata[150]));
Q_FDP0UA U4157 ( .D(n1646), .QTFCLK( ), .Q(xdata[149]));
Q_FDP0UA U4158 ( .D(n1648), .QTFCLK( ), .Q(xdata[148]));
Q_FDP0UA U4159 ( .D(n1650), .QTFCLK( ), .Q(xdata[147]));
Q_FDP0UA U4160 ( .D(n1652), .QTFCLK( ), .Q(xdata[146]));
Q_FDP0UA U4161 ( .D(n1654), .QTFCLK( ), .Q(xdata[145]));
Q_FDP0UA U4162 ( .D(n1656), .QTFCLK( ), .Q(xdata[144]));
Q_FDP0UA U4163 ( .D(n1658), .QTFCLK( ), .Q(xdata[143]));
Q_FDP0UA U4164 ( .D(n1660), .QTFCLK( ), .Q(xdata[142]));
Q_FDP0UA U4165 ( .D(n1662), .QTFCLK( ), .Q(xdata[141]));
Q_FDP0UA U4166 ( .D(n1664), .QTFCLK( ), .Q(xdata[140]));
Q_FDP0UA U4167 ( .D(n1666), .QTFCLK( ), .Q(xdata[139]));
Q_FDP0UA U4168 ( .D(n1668), .QTFCLK( ), .Q(xdata[138]));
Q_FDP0UA U4169 ( .D(n1670), .QTFCLK( ), .Q(xdata[137]));
Q_FDP0UA U4170 ( .D(n1672), .QTFCLK( ), .Q(xdata[136]));
Q_FDP0UA U4171 ( .D(n1674), .QTFCLK( ), .Q(xdata[135]));
Q_FDP0UA U4172 ( .D(n1676), .QTFCLK( ), .Q(xdata[134]));
Q_FDP0UA U4173 ( .D(n1678), .QTFCLK( ), .Q(xdata[133]));
Q_FDP0UA U4174 ( .D(n1680), .QTFCLK( ), .Q(xdata[132]));
Q_FDP0UA U4175 ( .D(n1682), .QTFCLK( ), .Q(xdata[131]));
Q_FDP0UA U4176 ( .D(n1684), .QTFCLK( ), .Q(xdata[130]));
Q_FDP0UA U4177 ( .D(n1686), .QTFCLK( ), .Q(xdata[129]));
Q_FDP0UA U4178 ( .D(n1688), .QTFCLK( ), .Q(xdata[128]));
Q_FDP0UA U4179 ( .D(n1690), .QTFCLK( ), .Q(xdata[127]));
Q_FDP0UA U4180 ( .D(n1692), .QTFCLK( ), .Q(xdata[126]));
Q_FDP0UA U4181 ( .D(n1694), .QTFCLK( ), .Q(xdata[125]));
Q_FDP0UA U4182 ( .D(n1696), .QTFCLK( ), .Q(xdata[124]));
Q_FDP0UA U4183 ( .D(n1698), .QTFCLK( ), .Q(xdata[123]));
Q_FDP0UA U4184 ( .D(n1700), .QTFCLK( ), .Q(xdata[122]));
Q_FDP0UA U4185 ( .D(n1702), .QTFCLK( ), .Q(xdata[121]));
Q_FDP0UA U4186 ( .D(n1704), .QTFCLK( ), .Q(xdata[120]));
Q_FDP0UA U4187 ( .D(n1706), .QTFCLK( ), .Q(xdata[119]));
Q_FDP0UA U4188 ( .D(n1708), .QTFCLK( ), .Q(xdata[118]));
Q_FDP0UA U4189 ( .D(n1710), .QTFCLK( ), .Q(xdata[117]));
Q_FDP0UA U4190 ( .D(n1712), .QTFCLK( ), .Q(xdata[116]));
Q_FDP0UA U4191 ( .D(n1714), .QTFCLK( ), .Q(xdata[115]));
Q_FDP0UA U4192 ( .D(n1716), .QTFCLK( ), .Q(xdata[114]));
Q_FDP0UA U4193 ( .D(n1718), .QTFCLK( ), .Q(xdata[113]));
Q_FDP0UA U4194 ( .D(n1720), .QTFCLK( ), .Q(xdata[112]));
Q_FDP0UA U4195 ( .D(n1722), .QTFCLK( ), .Q(xdata[111]));
Q_FDP0UA U4196 ( .D(n1724), .QTFCLK( ), .Q(xdata[110]));
Q_FDP0UA U4197 ( .D(n1726), .QTFCLK( ), .Q(xdata[109]));
Q_FDP0UA U4198 ( .D(n1728), .QTFCLK( ), .Q(xdata[108]));
Q_FDP0UA U4199 ( .D(n1730), .QTFCLK( ), .Q(xdata[107]));
Q_FDP0UA U4200 ( .D(n1732), .QTFCLK( ), .Q(xdata[106]));
Q_FDP0UA U4201 ( .D(n1734), .QTFCLK( ), .Q(xdata[105]));
Q_FDP0UA U4202 ( .D(n1736), .QTFCLK( ), .Q(xdata[104]));
Q_FDP0UA U4203 ( .D(n1738), .QTFCLK( ), .Q(xdata[103]));
Q_FDP0UA U4204 ( .D(n1740), .QTFCLK( ), .Q(xdata[102]));
Q_FDP0UA U4205 ( .D(n1742), .QTFCLK( ), .Q(xdata[101]));
Q_FDP0UA U4206 ( .D(n1744), .QTFCLK( ), .Q(xdata[100]));
Q_FDP0UA U4207 ( .D(n1746), .QTFCLK( ), .Q(xdata[99]));
Q_FDP0UA U4208 ( .D(n1748), .QTFCLK( ), .Q(xdata[98]));
Q_FDP0UA U4209 ( .D(n1750), .QTFCLK( ), .Q(xdata[97]));
Q_FDP0UA U4210 ( .D(n1752), .QTFCLK( ), .Q(xdata[96]));
Q_FDP0UA U4211 ( .D(n1754), .QTFCLK( ), .Q(xdata[95]));
Q_FDP0UA U4212 ( .D(n1756), .QTFCLK( ), .Q(xdata[94]));
Q_FDP0UA U4213 ( .D(n1758), .QTFCLK( ), .Q(xdata[93]));
Q_FDP0UA U4214 ( .D(n1760), .QTFCLK( ), .Q(xdata[92]));
Q_FDP0UA U4215 ( .D(n1762), .QTFCLK( ), .Q(xdata[91]));
Q_FDP0UA U4216 ( .D(n1764), .QTFCLK( ), .Q(xdata[90]));
Q_FDP0UA U4217 ( .D(n1766), .QTFCLK( ), .Q(xdata[89]));
Q_FDP0UA U4218 ( .D(n1768), .QTFCLK( ), .Q(xdata[88]));
Q_FDP0UA U4219 ( .D(n1770), .QTFCLK( ), .Q(xdata[87]));
Q_FDP0UA U4220 ( .D(n1772), .QTFCLK( ), .Q(xdata[86]));
Q_FDP0UA U4221 ( .D(n1774), .QTFCLK( ), .Q(xdata[85]));
Q_FDP0UA U4222 ( .D(n1776), .QTFCLK( ), .Q(xdata[84]));
Q_FDP0UA U4223 ( .D(n1778), .QTFCLK( ), .Q(xdata[83]));
Q_FDP0UA U4224 ( .D(n1780), .QTFCLK( ), .Q(xdata[82]));
Q_FDP0UA U4225 ( .D(n1782), .QTFCLK( ), .Q(xdata[81]));
Q_FDP0UA U4226 ( .D(n1784), .QTFCLK( ), .Q(xdata[80]));
Q_FDP0UA U4227 ( .D(n1786), .QTFCLK( ), .Q(xdata[79]));
Q_FDP0UA U4228 ( .D(n1788), .QTFCLK( ), .Q(xdata[78]));
Q_FDP0UA U4229 ( .D(n1790), .QTFCLK( ), .Q(xdata[77]));
Q_FDP0UA U4230 ( .D(n1792), .QTFCLK( ), .Q(xdata[76]));
Q_FDP0UA U4231 ( .D(n1794), .QTFCLK( ), .Q(xdata[75]));
Q_FDP0UA U4232 ( .D(n1796), .QTFCLK( ), .Q(xdata[74]));
Q_FDP0UA U4233 ( .D(n1798), .QTFCLK( ), .Q(xdata[73]));
Q_FDP0UA U4234 ( .D(n1800), .QTFCLK( ), .Q(xdata[72]));
Q_FDP0UA U4235 ( .D(n1802), .QTFCLK( ), .Q(xdata[71]));
Q_FDP0UA U4236 ( .D(n1804), .QTFCLK( ), .Q(xdata[70]));
Q_FDP0UA U4237 ( .D(n1806), .QTFCLK( ), .Q(xdata[69]));
Q_FDP0UA U4238 ( .D(n1808), .QTFCLK( ), .Q(xdata[68]));
Q_FDP0UA U4239 ( .D(n1810), .QTFCLK( ), .Q(xdata[67]));
Q_FDP0UA U4240 ( .D(n1812), .QTFCLK( ), .Q(xdata[66]));
Q_FDP0UA U4241 ( .D(n1814), .QTFCLK( ), .Q(xdata[65]));
Q_FDP0UA U4242 ( .D(n1816), .QTFCLK( ), .Q(xdata[64]));
Q_FDP0UA U4243 ( .D(n1818), .QTFCLK( ), .Q(xdata[63]));
Q_FDP0UA U4244 ( .D(n1820), .QTFCLK( ), .Q(xdata[62]));
Q_FDP0UA U4245 ( .D(n1822), .QTFCLK( ), .Q(xdata[61]));
Q_FDP0UA U4246 ( .D(n1824), .QTFCLK( ), .Q(xdata[60]));
Q_FDP0UA U4247 ( .D(n1826), .QTFCLK( ), .Q(xdata[59]));
Q_FDP0UA U4248 ( .D(n1828), .QTFCLK( ), .Q(xdata[58]));
Q_FDP0UA U4249 ( .D(n1830), .QTFCLK( ), .Q(xdata[57]));
Q_FDP0UA U4250 ( .D(n1832), .QTFCLK( ), .Q(xdata[56]));
Q_FDP0UA U4251 ( .D(n1834), .QTFCLK( ), .Q(xdata[55]));
Q_FDP0UA U4252 ( .D(n1836), .QTFCLK( ), .Q(xdata[54]));
Q_FDP0UA U4253 ( .D(n1838), .QTFCLK( ), .Q(xdata[53]));
Q_FDP0UA U4254 ( .D(n1840), .QTFCLK( ), .Q(xdata[52]));
Q_FDP0UA U4255 ( .D(n1842), .QTFCLK( ), .Q(xdata[51]));
Q_FDP0UA U4256 ( .D(n1844), .QTFCLK( ), .Q(xdata[50]));
Q_FDP0UA U4257 ( .D(n1846), .QTFCLK( ), .Q(xdata[49]));
Q_FDP0UA U4258 ( .D(n1848), .QTFCLK( ), .Q(xdata[48]));
Q_FDP0UA U4259 ( .D(n1850), .QTFCLK( ), .Q(xdata[47]));
Q_FDP0UA U4260 ( .D(n1852), .QTFCLK( ), .Q(xdata[46]));
Q_FDP0UA U4261 ( .D(n1854), .QTFCLK( ), .Q(xdata[45]));
Q_FDP0UA U4262 ( .D(n1856), .QTFCLK( ), .Q(xdata[44]));
Q_FDP0UA U4263 ( .D(n1858), .QTFCLK( ), .Q(xdata[43]));
Q_FDP0UA U4264 ( .D(n1860), .QTFCLK( ), .Q(xdata[42]));
Q_FDP0UA U4265 ( .D(n1862), .QTFCLK( ), .Q(xdata[41]));
Q_FDP0UA U4266 ( .D(n1864), .QTFCLK( ), .Q(xdata[40]));
Q_FDP0UA U4267 ( .D(n1866), .QTFCLK( ), .Q(xdata[39]));
Q_FDP0UA U4268 ( .D(n1868), .QTFCLK( ), .Q(xdata[38]));
Q_FDP0UA U4269 ( .D(n1870), .QTFCLK( ), .Q(xdata[37]));
Q_FDP0UA U4270 ( .D(n1872), .QTFCLK( ), .Q(xdata[36]));
Q_FDP0UA U4271 ( .D(n1874), .QTFCLK( ), .Q(xdata[35]));
Q_FDP0UA U4272 ( .D(n1876), .QTFCLK( ), .Q(xdata[34]));
Q_FDP0UA U4273 ( .D(n1878), .QTFCLK( ), .Q(xdata[33]));
Q_FDP0UA U4274 ( .D(n1880), .QTFCLK( ), .Q(xdata[32]));
Q_FDP0UA U4275 ( .D(n1882), .QTFCLK( ), .Q(xdata[31]));
Q_FDP0UA U4276 ( .D(n1884), .QTFCLK( ), .Q(xdata[30]));
Q_FDP0UA U4277 ( .D(n1886), .QTFCLK( ), .Q(xdata[29]));
Q_FDP0UA U4278 ( .D(n1888), .QTFCLK( ), .Q(xdata[28]));
Q_FDP0UA U4279 ( .D(n1890), .QTFCLK( ), .Q(xdata[27]));
Q_FDP0UA U4280 ( .D(n1892), .QTFCLK( ), .Q(xdata[26]));
Q_FDP0UA U4281 ( .D(n1894), .QTFCLK( ), .Q(xdata[25]));
Q_FDP0UA U4282 ( .D(n1896), .QTFCLK( ), .Q(xdata[24]));
Q_FDP0UA U4283 ( .D(n1898), .QTFCLK( ), .Q(xdata[23]));
Q_FDP0UA U4284 ( .D(n1900), .QTFCLK( ), .Q(xdata[22]));
Q_FDP0UA U4285 ( .D(n1902), .QTFCLK( ), .Q(xdata[21]));
Q_FDP0UA U4286 ( .D(n1904), .QTFCLK( ), .Q(xdata[20]));
Q_FDP0UA U4287 ( .D(n1906), .QTFCLK( ), .Q(xdata[19]));
Q_FDP0UA U4288 ( .D(n1908), .QTFCLK( ), .Q(xdata[18]));
Q_FDP0UA U4289 ( .D(n1910), .QTFCLK( ), .Q(xdata[17]));
Q_FDP0UA U4290 ( .D(n1912), .QTFCLK( ), .Q(xdata[16]));
Q_FDP0UA U4291 ( .D(n1914), .QTFCLK( ), .Q(xdata[15]));
Q_FDP0UA U4292 ( .D(n1916), .QTFCLK( ), .Q(xdata[14]));
Q_FDP0UA U4293 ( .D(n1918), .QTFCLK( ), .Q(xdata[13]));
Q_FDP0UA U4294 ( .D(n1920), .QTFCLK( ), .Q(xdata[12]));
Q_FDP0UA U4295 ( .D(n1922), .QTFCLK( ), .Q(xdata[11]));
Q_FDP0UA U4296 ( .D(n1924), .QTFCLK( ), .Q(xdata[10]));
Q_FDP0UA U4297 ( .D(n1926), .QTFCLK( ), .Q(xdata[9]));
Q_FDP0UA U4298 ( .D(n1928), .QTFCLK( ), .Q(xdata[8]));
Q_FDP0UA U4299 ( .D(n1930), .QTFCLK( ), .Q(xdata[7]));
Q_FDP0UA U4300 ( .D(n1932), .QTFCLK( ), .Q(xdata[6]));
Q_FDP0UA U4301 ( .D(n1934), .QTFCLK( ), .Q(xdata[5]));
Q_FDP0UA U4302 ( .D(n1936), .QTFCLK( ), .Q(xdata[4]));
Q_FDP0UA U4303 ( .D(n1938), .QTFCLK( ), .Q(xdata[3]));
Q_FDP0UA U4304 ( .D(n1940), .QTFCLK( ), .Q(xdata[2]));
Q_FDP0UA U4305 ( .D(n1942), .QTFCLK( ), .Q(xdata[1]));
Q_FDP0UA U4306 ( .D(n1944), .QTFCLK( ), .Q(xdata[0]));
Q_FDP0UA U4307 ( .D(n889), .QTFCLK( ), .Q(wrtCnt[63]));
Q_MX02 U4308 ( .S(n797), .A0(n1946), .A1(wrtCnt[63]), .Z(n889));
Q_FDP0UA U4309 ( .D(n888), .QTFCLK( ), .Q(wrtCnt[62]));
Q_MX02 U4310 ( .S(n797), .A0(n1947), .A1(wrtCnt[62]), .Z(n888));
Q_FDP0UA U4311 ( .D(n887), .QTFCLK( ), .Q(wrtCnt[61]));
Q_MX02 U4312 ( .S(n797), .A0(n1948), .A1(wrtCnt[61]), .Z(n887));
Q_FDP0UA U4313 ( .D(n886), .QTFCLK( ), .Q(wrtCnt[60]));
Q_MX02 U4314 ( .S(n797), .A0(n1949), .A1(wrtCnt[60]), .Z(n886));
Q_FDP0UA U4315 ( .D(n885), .QTFCLK( ), .Q(wrtCnt[59]));
Q_MX02 U4316 ( .S(n797), .A0(n1950), .A1(wrtCnt[59]), .Z(n885));
Q_FDP0UA U4317 ( .D(n884), .QTFCLK( ), .Q(wrtCnt[58]));
Q_MX02 U4318 ( .S(n797), .A0(n1951), .A1(wrtCnt[58]), .Z(n884));
Q_FDP0UA U4319 ( .D(n883), .QTFCLK( ), .Q(wrtCnt[57]));
Q_MX02 U4320 ( .S(n797), .A0(n1952), .A1(wrtCnt[57]), .Z(n883));
Q_FDP0UA U4321 ( .D(n882), .QTFCLK( ), .Q(wrtCnt[56]));
Q_MX02 U4322 ( .S(n797), .A0(n1953), .A1(wrtCnt[56]), .Z(n882));
Q_FDP0UA U4323 ( .D(n881), .QTFCLK( ), .Q(wrtCnt[55]));
Q_MX02 U4324 ( .S(n797), .A0(n1954), .A1(wrtCnt[55]), .Z(n881));
Q_FDP0UA U4325 ( .D(n880), .QTFCLK( ), .Q(wrtCnt[54]));
Q_MX02 U4326 ( .S(n797), .A0(n1955), .A1(wrtCnt[54]), .Z(n880));
Q_FDP0UA U4327 ( .D(n879), .QTFCLK( ), .Q(wrtCnt[53]));
Q_MX02 U4328 ( .S(n797), .A0(n1956), .A1(wrtCnt[53]), .Z(n879));
Q_FDP0UA U4329 ( .D(n878), .QTFCLK( ), .Q(wrtCnt[52]));
Q_MX02 U4330 ( .S(n797), .A0(n1957), .A1(wrtCnt[52]), .Z(n878));
Q_FDP0UA U4331 ( .D(n877), .QTFCLK( ), .Q(wrtCnt[51]));
Q_MX02 U4332 ( .S(n797), .A0(n1958), .A1(wrtCnt[51]), .Z(n877));
Q_FDP0UA U4333 ( .D(n876), .QTFCLK( ), .Q(wrtCnt[50]));
Q_MX02 U4334 ( .S(n797), .A0(n1959), .A1(wrtCnt[50]), .Z(n876));
Q_FDP0UA U4335 ( .D(n875), .QTFCLK( ), .Q(wrtCnt[49]));
Q_MX02 U4336 ( .S(n797), .A0(n1960), .A1(wrtCnt[49]), .Z(n875));
Q_FDP0UA U4337 ( .D(n874), .QTFCLK( ), .Q(wrtCnt[48]));
Q_MX02 U4338 ( .S(n797), .A0(n1961), .A1(wrtCnt[48]), .Z(n874));
Q_FDP0UA U4339 ( .D(n873), .QTFCLK( ), .Q(wrtCnt[47]));
Q_MX02 U4340 ( .S(n797), .A0(n1962), .A1(wrtCnt[47]), .Z(n873));
Q_FDP0UA U4341 ( .D(n872), .QTFCLK( ), .Q(wrtCnt[46]));
Q_MX02 U4342 ( .S(n797), .A0(n1963), .A1(wrtCnt[46]), .Z(n872));
Q_FDP0UA U4343 ( .D(n871), .QTFCLK( ), .Q(wrtCnt[45]));
Q_MX02 U4344 ( .S(n797), .A0(n1964), .A1(wrtCnt[45]), .Z(n871));
Q_FDP0UA U4345 ( .D(n870), .QTFCLK( ), .Q(wrtCnt[44]));
Q_MX02 U4346 ( .S(n797), .A0(n1965), .A1(wrtCnt[44]), .Z(n870));
Q_FDP0UA U4347 ( .D(n869), .QTFCLK( ), .Q(wrtCnt[43]));
Q_MX02 U4348 ( .S(n797), .A0(n1966), .A1(wrtCnt[43]), .Z(n869));
Q_FDP0UA U4349 ( .D(n868), .QTFCLK( ), .Q(wrtCnt[42]));
Q_MX02 U4350 ( .S(n797), .A0(n1967), .A1(wrtCnt[42]), .Z(n868));
Q_FDP0UA U4351 ( .D(n867), .QTFCLK( ), .Q(wrtCnt[41]));
Q_MX02 U4352 ( .S(n797), .A0(n1968), .A1(wrtCnt[41]), .Z(n867));
Q_FDP0UA U4353 ( .D(n866), .QTFCLK( ), .Q(wrtCnt[40]));
Q_MX02 U4354 ( .S(n797), .A0(n1969), .A1(wrtCnt[40]), .Z(n866));
Q_FDP0UA U4355 ( .D(n865), .QTFCLK( ), .Q(wrtCnt[39]));
Q_MX02 U4356 ( .S(n797), .A0(n1970), .A1(wrtCnt[39]), .Z(n865));
Q_FDP0UA U4357 ( .D(n864), .QTFCLK( ), .Q(wrtCnt[38]));
Q_MX02 U4358 ( .S(n797), .A0(n1971), .A1(wrtCnt[38]), .Z(n864));
Q_FDP0UA U4359 ( .D(n863), .QTFCLK( ), .Q(wrtCnt[37]));
Q_MX02 U4360 ( .S(n797), .A0(n1972), .A1(wrtCnt[37]), .Z(n863));
Q_FDP0UA U4361 ( .D(n862), .QTFCLK( ), .Q(wrtCnt[36]));
Q_MX02 U4362 ( .S(n797), .A0(n1973), .A1(wrtCnt[36]), .Z(n862));
Q_FDP0UA U4363 ( .D(n861), .QTFCLK( ), .Q(wrtCnt[35]));
Q_MX02 U4364 ( .S(n797), .A0(n1974), .A1(wrtCnt[35]), .Z(n861));
Q_FDP0UA U4365 ( .D(n860), .QTFCLK( ), .Q(wrtCnt[34]));
Q_MX02 U4366 ( .S(n797), .A0(n1975), .A1(wrtCnt[34]), .Z(n860));
Q_FDP0UA U4367 ( .D(n859), .QTFCLK( ), .Q(wrtCnt[33]));
Q_MX02 U4368 ( .S(n797), .A0(n1976), .A1(wrtCnt[33]), .Z(n859));
Q_FDP0UA U4369 ( .D(n858), .QTFCLK( ), .Q(wrtCnt[32]));
Q_MX02 U4370 ( .S(n797), .A0(n1977), .A1(wrtCnt[32]), .Z(n858));
Q_FDP0UA U4371 ( .D(n857), .QTFCLK( ), .Q(wrtCnt[31]));
Q_MX02 U4372 ( .S(n797), .A0(n1978), .A1(wrtCnt[31]), .Z(n857));
Q_FDP0UA U4373 ( .D(n856), .QTFCLK( ), .Q(wrtCnt[30]));
Q_MX02 U4374 ( .S(n797), .A0(n1979), .A1(wrtCnt[30]), .Z(n856));
Q_FDP0UA U4375 ( .D(n855), .QTFCLK( ), .Q(wrtCnt[29]));
Q_MX02 U4376 ( .S(n797), .A0(n1980), .A1(wrtCnt[29]), .Z(n855));
Q_FDP0UA U4377 ( .D(n854), .QTFCLK( ), .Q(wrtCnt[28]));
Q_MX02 U4378 ( .S(n797), .A0(n1981), .A1(wrtCnt[28]), .Z(n854));
Q_FDP0UA U4379 ( .D(n853), .QTFCLK( ), .Q(wrtCnt[27]));
Q_MX02 U4380 ( .S(n797), .A0(n1982), .A1(wrtCnt[27]), .Z(n853));
Q_FDP0UA U4381 ( .D(n852), .QTFCLK( ), .Q(wrtCnt[26]));
Q_MX02 U4382 ( .S(n797), .A0(n1983), .A1(wrtCnt[26]), .Z(n852));
Q_FDP0UA U4383 ( .D(n851), .QTFCLK( ), .Q(wrtCnt[25]));
Q_MX02 U4384 ( .S(n797), .A0(n1984), .A1(wrtCnt[25]), .Z(n851));
Q_FDP0UA U4385 ( .D(n850), .QTFCLK( ), .Q(wrtCnt[24]));
Q_MX02 U4386 ( .S(n797), .A0(n1985), .A1(wrtCnt[24]), .Z(n850));
Q_FDP0UA U4387 ( .D(n849), .QTFCLK( ), .Q(wrtCnt[23]));
Q_MX02 U4388 ( .S(n797), .A0(n1986), .A1(wrtCnt[23]), .Z(n849));
Q_FDP0UA U4389 ( .D(n848), .QTFCLK( ), .Q(wrtCnt[22]));
Q_MX02 U4390 ( .S(n797), .A0(n1987), .A1(wrtCnt[22]), .Z(n848));
Q_FDP0UA U4391 ( .D(n847), .QTFCLK( ), .Q(wrtCnt[21]));
Q_MX02 U4392 ( .S(n797), .A0(n1988), .A1(wrtCnt[21]), .Z(n847));
Q_FDP0UA U4393 ( .D(n846), .QTFCLK( ), .Q(wrtCnt[20]));
Q_MX02 U4394 ( .S(n797), .A0(n1989), .A1(wrtCnt[20]), .Z(n846));
Q_FDP0UA U4395 ( .D(n845), .QTFCLK( ), .Q(wrtCnt[19]));
Q_MX02 U4396 ( .S(n797), .A0(n1990), .A1(wrtCnt[19]), .Z(n845));
Q_FDP0UA U4397 ( .D(n844), .QTFCLK( ), .Q(wrtCnt[18]));
Q_MX02 U4398 ( .S(n797), .A0(n1991), .A1(wrtCnt[18]), .Z(n844));
Q_FDP0UA U4399 ( .D(n843), .QTFCLK( ), .Q(wrtCnt[17]));
Q_MX02 U4400 ( .S(n797), .A0(n1992), .A1(wrtCnt[17]), .Z(n843));
Q_FDP0UA U4401 ( .D(n842), .QTFCLK( ), .Q(wrtCnt[16]));
Q_MX02 U4402 ( .S(n797), .A0(n1993), .A1(wrtCnt[16]), .Z(n842));
Q_FDP0UA U4403 ( .D(n841), .QTFCLK( ), .Q(wrtCnt[15]));
Q_MX02 U4404 ( .S(n797), .A0(n1994), .A1(wrtCnt[15]), .Z(n841));
Q_FDP0UA U4405 ( .D(n840), .QTFCLK( ), .Q(wrtCnt[14]));
Q_MX02 U4406 ( .S(n797), .A0(n1995), .A1(wrtCnt[14]), .Z(n840));
Q_FDP0UA U4407 ( .D(n839), .QTFCLK( ), .Q(wrtCnt[13]));
Q_MX02 U4408 ( .S(n797), .A0(n1996), .A1(wrtCnt[13]), .Z(n839));
Q_FDP0UA U4409 ( .D(n838), .QTFCLK( ), .Q(wrtCnt[12]));
Q_MX02 U4410 ( .S(n797), .A0(n1997), .A1(wrtCnt[12]), .Z(n838));
Q_FDP0UA U4411 ( .D(n837), .QTFCLK( ), .Q(wrtCnt[11]));
Q_MX02 U4412 ( .S(n797), .A0(n1998), .A1(wrtCnt[11]), .Z(n837));
Q_FDP0UA U4413 ( .D(n836), .QTFCLK( ), .Q(wrtCnt[10]));
Q_MX02 U4414 ( .S(n797), .A0(n1999), .A1(wrtCnt[10]), .Z(n836));
Q_FDP0UA U4415 ( .D(n835), .QTFCLK( ), .Q(wrtCnt[9]));
Q_MX02 U4416 ( .S(n797), .A0(n2000), .A1(wrtCnt[9]), .Z(n835));
Q_FDP0UA U4417 ( .D(n834), .QTFCLK( ), .Q(wrtCnt[8]));
Q_MX02 U4418 ( .S(n797), .A0(n2001), .A1(wrtCnt[8]), .Z(n834));
Q_FDP0UA U4419 ( .D(n833), .QTFCLK( ), .Q(wrtCnt[7]));
Q_MX02 U4420 ( .S(n797), .A0(n2002), .A1(wrtCnt[7]), .Z(n833));
Q_FDP0UA U4421 ( .D(n832), .QTFCLK( ), .Q(wrtCnt[6]));
Q_MX02 U4422 ( .S(n797), .A0(n2003), .A1(wrtCnt[6]), .Z(n832));
Q_FDP0UA U4423 ( .D(n831), .QTFCLK( ), .Q(wrtCnt[5]));
Q_MX02 U4424 ( .S(n797), .A0(n2004), .A1(wrtCnt[5]), .Z(n831));
Q_FDP0UA U4425 ( .D(n830), .QTFCLK( ), .Q(wrtCnt[4]));
Q_MX02 U4426 ( .S(n797), .A0(n2005), .A1(wrtCnt[4]), .Z(n830));
Q_FDP0UA U4427 ( .D(n829), .QTFCLK( ), .Q(wrtCnt[3]));
Q_MX02 U4428 ( .S(n797), .A0(n2006), .A1(wrtCnt[3]), .Z(n829));
Q_FDP0UA U4429 ( .D(n828), .QTFCLK( ), .Q(wrtCnt[2]));
Q_MX02 U4430 ( .S(n797), .A0(n2007), .A1(wrtCnt[2]), .Z(n828));
Q_FDP0UA U4431 ( .D(n827), .QTFCLK( ), .Q(wrtCnt[1]));
Q_MX02 U4432 ( .S(n797), .A0(n2008), .A1(wrtCnt[1]), .Z(n827));
Q_FDP0UA U4433 ( .D(n826), .QTFCLK( ), .Q(wrtCnt[0]));
Q_MX02 U4434 ( .S(n797), .A0(n2009), .A1(wrtCnt[0]), .Z(n826));
Q_FDP0UA U4435 ( .D(n2010), .QTFCLK( ), .Q(writeLen[5]));
Q_FDP0UA U4436 ( .D(n2012), .QTFCLK( ), .Q(writeLen[4]));
Q_FDP0UA U4437 ( .D(n2014), .QTFCLK( ), .Q(writeLen[3]));
Q_FDP0UA U4438 ( .D(n2016), .QTFCLK( ), .Q(writeLen[2]));
Q_FDP0UA U4439 ( .D(n2018), .QTFCLK( ), .Q(writeLen[1]));
Q_FDP0UA U4440 ( .D(n2020), .QTFCLK( ), .Q(writeLen[0]));
Q_FDP0UA U4441 ( .D(n825), .QTFCLK( ), .Q(argLen[11]));
Q_MX02 U4442 ( .S(n807), .A0(n2144), .A1(argLen[11]), .Z(n825));
Q_FDP0UA U4443 ( .D(n824), .QTFCLK( ), .Q(argLen[10]));
Q_MX02 U4444 ( .S(n807), .A0(n2145), .A1(argLen[10]), .Z(n824));
Q_FDP0UA U4445 ( .D(n823), .QTFCLK( ), .Q(argLen[9]));
Q_MX02 U4446 ( .S(n807), .A0(n2146), .A1(argLen[9]), .Z(n823));
Q_FDP0UA U4447 ( .D(n822), .QTFCLK( ), .Q(argLen[8]));
Q_MX02 U4448 ( .S(n807), .A0(n2147), .A1(argLen[8]), .Z(n822));
Q_FDP0UA U4449 ( .D(n821), .QTFCLK( ), .Q(argLen[7]));
Q_MX02 U4450 ( .S(n807), .A0(n2148), .A1(argLen[7]), .Z(n821));
Q_FDP0UA U4451 ( .D(n820), .QTFCLK( ), .Q(argLen[6]));
Q_MX02 U4452 ( .S(n807), .A0(n2149), .A1(argLen[6]), .Z(n820));
Q_FDP0UA U4453 ( .D(n819), .QTFCLK( ), .Q(argLen[5]));
Q_MX02 U4454 ( .S(n807), .A0(n2150), .A1(argLen[5]), .Z(n819));
Q_FDP0UA U4455 ( .D(n818), .QTFCLK( ), .Q(argLen[4]));
Q_MX02 U4456 ( .S(n807), .A0(n2151), .A1(argLen[4]), .Z(n818));
Q_FDP0UA U4457 ( .D(n817), .QTFCLK( ), .Q(argLen[3]));
Q_MX02 U4458 ( .S(n807), .A0(n2152), .A1(argLen[3]), .Z(n817));
Q_FDP0UA U4459 ( .D(n816), .QTFCLK( ), .Q(argLen[2]));
Q_MX02 U4460 ( .S(n807), .A0(n2153), .A1(argLen[2]), .Z(n816));
Q_FDP0UA U4461 ( .D(n815), .QTFCLK( ), .Q(argLen[1]));
Q_MX02 U4462 ( .S(n807), .A0(n2154), .A1(argLen[1]), .Z(n815));
Q_FDP0UA U4463 ( .D(n814), .QTFCLK( ), .Q(argLen[0]));
Q_MX02 U4464 ( .S(n807), .A0(n2155), .A1(argLen[0]), .Z(n814));
Q_INV U4465 ( .A(n783), .Z(n787));
Q_AN02 U4466 ( .A0(n812), .A1(n811), .Z(n813));
Q_AN03 U4467 ( .A0(n809), .A1(GFcbid[0]), .A2(n810), .Z(n811));
Q_INV U4468 ( .A(n808), .Z(n786));
Q_OR02 U4469 ( .A0(n785), .A1(n807), .Z(n808));
Q_AN03 U4470 ( .A0(n810), .A1(n805), .A2(n806), .Z(n785));
Q_AN03 U4471 ( .A0(GFcbid[1]), .A1(GFcbid[0]), .A2(n809), .Z(n805));
Q_AN02 U4472 ( .A0(n804), .A1(n803), .Z(n806));
Q_AN03 U4473 ( .A0(n801), .A1(n800), .A2(n802), .Z(n804));
Q_AN02 U4474 ( .A0(n65), .A1(n784), .Z(n801));
Q_OR02 U4475 ( .A0(n799), .A1(n798), .Z(n807));
Q_INV U4476 ( .A(n801), .Z(n798));
Q_AN02 U4477 ( .A0(n65), .A1(n796), .Z(n797));
Q_INV U4478 ( .A(n784), .Z(n795));
Q_OR03 U4479 ( .A0(n795), .A1(n783), .A2(n799), .Z(n796));
Q_AN03 U4480 ( .A0(n810), .A1(n794), .A2(n812), .Z(n799));
Q_AN03 U4481 ( .A0(n793), .A1(GFcbid[0]), .A2(n809), .Z(n794));
Q_INV U4482 ( .A(GFcbid[1]), .Z(n793));
Q_AN02 U4483 ( .A0(GFcbid[3]), .A1(GFcbid[2]), .Z(n809));
Q_AN03 U4484 ( .A0(GFcbid[5]), .A1(GFcbid[4]), .A2(n792), .Z(n810));
Q_AN03 U4485 ( .A0(GFcbid[7]), .A1(GFcbid[6]), .A2(n791), .Z(n792));
Q_AN02 U4486 ( .A0(GFcbid[9]), .A1(GFcbid[8]), .Z(n791));
Q_AN03 U4487 ( .A0(GFcbid[11]), .A1(GFcbid[10]), .A2(n790), .Z(n803));
Q_AN03 U4488 ( .A0(GFcbid[13]), .A1(GFcbid[12]), .A2(n789), .Z(n790));
Q_AN02 U4489 ( .A0(GFcbid[15]), .A1(GFcbid[14]), .Z(n789));
Q_AN03 U4490 ( .A0(n800), .A1(n802), .A2(n803), .Z(n812));
Q_AN02 U4491 ( .A0(GFcbid[17]), .A1(GFcbid[16]), .Z(n802));
Q_AN02 U4492 ( .A0(GFcbid[19]), .A1(GFcbid[18]), .Z(n800));
Q_AN02 U4493 ( .A0(n65), .A1(ofifoDataN[0]), .Z(n782));
Q_AN02 U4494 ( .A0(n65), .A1(ofifoDataN[1]), .Z(n781));
Q_AN02 U4495 ( .A0(n65), .A1(ofifoDataN[2]), .Z(n780));
Q_AN02 U4496 ( .A0(n65), .A1(ofifoDataN[3]), .Z(n779));
Q_AN02 U4497 ( .A0(n65), .A1(ofifoDataN[4]), .Z(n778));
Q_AN02 U4498 ( .A0(n65), .A1(ofifoDataN[5]), .Z(n777));
Q_AN02 U4499 ( .A0(n65), .A1(ofifoDataN[6]), .Z(n776));
Q_AN02 U4500 ( .A0(n65), .A1(ofifoDataN[7]), .Z(n775));
Q_AN02 U4501 ( .A0(n65), .A1(ofifoDataN[8]), .Z(n774));
Q_AN02 U4502 ( .A0(n65), .A1(ofifoDataN[9]), .Z(n773));
Q_AN02 U4503 ( .A0(n65), .A1(ofifoDataN[10]), .Z(n772));
Q_AN02 U4504 ( .A0(n65), .A1(ofifoDataN[11]), .Z(n771));
Q_AN02 U4505 ( .A0(n65), .A1(ofifoDataN[12]), .Z(n770));
Q_AN02 U4506 ( .A0(n65), .A1(ofifoDataN[13]), .Z(n769));
Q_AN02 U4507 ( .A0(n65), .A1(ofifoDataN[14]), .Z(n768));
Q_AN02 U4508 ( .A0(n65), .A1(ofifoDataN[15]), .Z(n767));
Q_AN02 U4509 ( .A0(n65), .A1(ofifoDataN[16]), .Z(n766));
Q_AN02 U4510 ( .A0(n65), .A1(ofifoDataN[17]), .Z(n765));
Q_AN02 U4511 ( .A0(n65), .A1(ofifoDataN[18]), .Z(n764));
Q_AN02 U4512 ( .A0(n65), .A1(ofifoDataN[19]), .Z(n763));
Q_AN02 U4513 ( .A0(n65), .A1(ofifoDataN[20]), .Z(n762));
Q_AN02 U4514 ( .A0(n65), .A1(ofifoDataN[21]), .Z(n761));
Q_AN02 U4515 ( .A0(n65), .A1(ofifoDataN[22]), .Z(n760));
Q_AN02 U4516 ( .A0(n65), .A1(ofifoDataN[23]), .Z(n759));
Q_AN02 U4517 ( .A0(n65), .A1(ofifoDataN[24]), .Z(n758));
Q_AN02 U4518 ( .A0(n65), .A1(ofifoDataN[25]), .Z(n757));
Q_AN02 U4519 ( .A0(n65), .A1(ofifoDataN[26]), .Z(n756));
Q_AN02 U4520 ( .A0(n65), .A1(ofifoDataN[27]), .Z(n755));
Q_AN02 U4521 ( .A0(n65), .A1(ofifoDataN[28]), .Z(n754));
Q_AN02 U4522 ( .A0(n65), .A1(ofifoDataN[29]), .Z(n753));
Q_AN02 U4523 ( .A0(n65), .A1(ofifoDataN[30]), .Z(n752));
Q_AN02 U4524 ( .A0(n65), .A1(ofifoDataN[31]), .Z(n751));
Q_AN02 U4525 ( .A0(n65), .A1(ofifoDataN[32]), .Z(n750));
Q_AN02 U4526 ( .A0(n65), .A1(ofifoDataN[33]), .Z(n749));
Q_AN02 U4527 ( .A0(n65), .A1(ofifoDataN[34]), .Z(n748));
Q_AN02 U4528 ( .A0(n65), .A1(ofifoDataN[35]), .Z(n747));
Q_AN02 U4529 ( .A0(n65), .A1(ofifoDataN[36]), .Z(n746));
Q_AN02 U4530 ( .A0(n65), .A1(ofifoDataN[37]), .Z(n745));
Q_AN02 U4531 ( .A0(n65), .A1(ofifoDataN[38]), .Z(n744));
Q_AN02 U4532 ( .A0(n65), .A1(ofifoDataN[39]), .Z(n743));
Q_AN02 U4533 ( .A0(n65), .A1(ofifoDataN[40]), .Z(n742));
Q_AN02 U4534 ( .A0(n65), .A1(ofifoDataN[41]), .Z(n741));
Q_AN02 U4535 ( .A0(n65), .A1(ofifoDataN[42]), .Z(n740));
Q_AN02 U4536 ( .A0(n65), .A1(ofifoDataN[43]), .Z(n739));
Q_AN02 U4537 ( .A0(n65), .A1(ofifoDataN[44]), .Z(n738));
Q_AN02 U4538 ( .A0(n65), .A1(ofifoDataN[45]), .Z(n737));
Q_AN02 U4539 ( .A0(n65), .A1(ofifoDataN[46]), .Z(n736));
Q_AN02 U4540 ( .A0(n65), .A1(ofifoDataN[47]), .Z(n735));
Q_AN02 U4541 ( .A0(n65), .A1(ofifoDataN[48]), .Z(n734));
Q_AN02 U4542 ( .A0(n65), .A1(ofifoDataN[49]), .Z(n733));
Q_AN02 U4543 ( .A0(n65), .A1(ofifoDataN[50]), .Z(n732));
Q_AN02 U4544 ( .A0(n65), .A1(ofifoDataN[51]), .Z(n731));
Q_AN02 U4545 ( .A0(n65), .A1(ofifoDataN[52]), .Z(n730));
Q_AN02 U4546 ( .A0(n65), .A1(ofifoDataN[53]), .Z(n729));
Q_AN02 U4547 ( .A0(n65), .A1(ofifoDataN[54]), .Z(n728));
Q_AN02 U4548 ( .A0(n65), .A1(ofifoDataN[55]), .Z(n727));
Q_AN02 U4549 ( .A0(n65), .A1(ofifoDataN[56]), .Z(n726));
Q_AN02 U4550 ( .A0(n65), .A1(ofifoDataN[57]), .Z(n725));
Q_AN02 U4551 ( .A0(n65), .A1(ofifoDataN[58]), .Z(n724));
Q_AN02 U4552 ( .A0(n65), .A1(ofifoDataN[59]), .Z(n723));
Q_AN02 U4553 ( .A0(n65), .A1(ofifoDataN[60]), .Z(n722));
Q_AN02 U4554 ( .A0(n65), .A1(ofifoDataN[61]), .Z(n721));
Q_AN02 U4555 ( .A0(n65), .A1(ofifoDataN[62]), .Z(n720));
Q_AN02 U4556 ( .A0(n65), .A1(ofifoDataN[63]), .Z(n719));
Q_AN02 U4557 ( .A0(n65), .A1(ofifoDataN[64]), .Z(n718));
Q_AN02 U4558 ( .A0(n65), .A1(ofifoDataN[65]), .Z(n717));
Q_AN02 U4559 ( .A0(n65), .A1(ofifoDataN[66]), .Z(n716));
Q_AN02 U4560 ( .A0(n65), .A1(ofifoDataN[67]), .Z(n715));
Q_AN02 U4561 ( .A0(n65), .A1(ofifoDataN[68]), .Z(n714));
Q_AN02 U4562 ( .A0(n65), .A1(ofifoDataN[69]), .Z(n713));
Q_AN02 U4563 ( .A0(n65), .A1(ofifoDataN[70]), .Z(n712));
Q_AN02 U4564 ( .A0(n65), .A1(ofifoDataN[71]), .Z(n711));
Q_AN02 U4565 ( .A0(n65), .A1(ofifoDataN[72]), .Z(n710));
Q_AN02 U4566 ( .A0(n65), .A1(ofifoDataN[73]), .Z(n709));
Q_AN02 U4567 ( .A0(n65), .A1(ofifoDataN[74]), .Z(n708));
Q_AN02 U4568 ( .A0(n65), .A1(ofifoDataN[75]), .Z(n707));
Q_AN02 U4569 ( .A0(n65), .A1(ofifoDataN[76]), .Z(n706));
Q_AN02 U4570 ( .A0(n65), .A1(ofifoDataN[77]), .Z(n705));
Q_AN02 U4571 ( .A0(n65), .A1(ofifoDataN[78]), .Z(n704));
Q_AN02 U4572 ( .A0(n65), .A1(ofifoDataN[79]), .Z(n703));
Q_AN02 U4573 ( .A0(n65), .A1(ofifoDataN[80]), .Z(n702));
Q_AN02 U4574 ( .A0(n65), .A1(ofifoDataN[81]), .Z(n701));
Q_AN02 U4575 ( .A0(n65), .A1(ofifoDataN[82]), .Z(n700));
Q_AN02 U4576 ( .A0(n65), .A1(ofifoDataN[83]), .Z(n699));
Q_AN02 U4577 ( .A0(n65), .A1(ofifoDataN[84]), .Z(n698));
Q_AN02 U4578 ( .A0(n65), .A1(ofifoDataN[85]), .Z(n697));
Q_AN02 U4579 ( .A0(n65), .A1(ofifoDataN[86]), .Z(n696));
Q_AN02 U4580 ( .A0(n65), .A1(ofifoDataN[87]), .Z(n695));
Q_AN02 U4581 ( .A0(n65), .A1(ofifoDataN[88]), .Z(n694));
Q_AN02 U4582 ( .A0(n65), .A1(ofifoDataN[89]), .Z(n693));
Q_AN02 U4583 ( .A0(n65), .A1(ofifoDataN[90]), .Z(n692));
Q_AN02 U4584 ( .A0(n65), .A1(ofifoDataN[91]), .Z(n691));
Q_AN02 U4585 ( .A0(n65), .A1(ofifoDataN[92]), .Z(n690));
Q_AN02 U4586 ( .A0(n65), .A1(ofifoDataN[93]), .Z(n689));
Q_AN02 U4587 ( .A0(n65), .A1(ofifoDataN[94]), .Z(n688));
Q_AN02 U4588 ( .A0(n65), .A1(ofifoDataN[95]), .Z(n687));
Q_AN02 U4589 ( .A0(n65), .A1(ofifoDataN[96]), .Z(n686));
Q_AN02 U4590 ( .A0(n65), .A1(ofifoDataN[97]), .Z(n685));
Q_AN02 U4591 ( .A0(n65), .A1(ofifoDataN[98]), .Z(n684));
Q_AN02 U4592 ( .A0(n65), .A1(ofifoDataN[99]), .Z(n683));
Q_AN02 U4593 ( .A0(n65), .A1(ofifoDataN[100]), .Z(n682));
Q_AN02 U4594 ( .A0(n65), .A1(ofifoDataN[101]), .Z(n681));
Q_AN02 U4595 ( .A0(n65), .A1(ofifoDataN[102]), .Z(n680));
Q_AN02 U4596 ( .A0(n65), .A1(ofifoDataN[103]), .Z(n679));
Q_AN02 U4597 ( .A0(n65), .A1(ofifoDataN[104]), .Z(n678));
Q_AN02 U4598 ( .A0(n65), .A1(ofifoDataN[105]), .Z(n677));
Q_AN02 U4599 ( .A0(n65), .A1(ofifoDataN[106]), .Z(n676));
Q_AN02 U4600 ( .A0(n65), .A1(ofifoDataN[107]), .Z(n675));
Q_AN02 U4601 ( .A0(n65), .A1(ofifoDataN[108]), .Z(n674));
Q_AN02 U4602 ( .A0(n65), .A1(ofifoDataN[109]), .Z(n673));
Q_AN02 U4603 ( .A0(n65), .A1(ofifoDataN[110]), .Z(n672));
Q_AN02 U4604 ( .A0(n65), .A1(ofifoDataN[111]), .Z(n671));
Q_AN02 U4605 ( .A0(n65), .A1(ofifoDataN[112]), .Z(n670));
Q_AN02 U4606 ( .A0(n65), .A1(ofifoDataN[113]), .Z(n669));
Q_AN02 U4607 ( .A0(n65), .A1(ofifoDataN[114]), .Z(n668));
Q_AN02 U4608 ( .A0(n65), .A1(ofifoDataN[115]), .Z(n667));
Q_AN02 U4609 ( .A0(n65), .A1(ofifoDataN[116]), .Z(n666));
Q_AN02 U4610 ( .A0(n65), .A1(ofifoDataN[117]), .Z(n665));
Q_AN02 U4611 ( .A0(n65), .A1(ofifoDataN[118]), .Z(n664));
Q_AN02 U4612 ( .A0(n65), .A1(ofifoDataN[119]), .Z(n663));
Q_AN02 U4613 ( .A0(n65), .A1(ofifoDataN[120]), .Z(n662));
Q_AN02 U4614 ( .A0(n65), .A1(ofifoDataN[121]), .Z(n661));
Q_AN02 U4615 ( .A0(n65), .A1(ofifoDataN[122]), .Z(n660));
Q_AN02 U4616 ( .A0(n65), .A1(ofifoDataN[123]), .Z(n659));
Q_AN02 U4617 ( .A0(n65), .A1(ofifoDataN[124]), .Z(n658));
Q_AN02 U4618 ( .A0(n65), .A1(ofifoDataN[125]), .Z(n657));
Q_AN02 U4619 ( .A0(n65), .A1(ofifoDataN[126]), .Z(n656));
Q_AN02 U4620 ( .A0(n65), .A1(ofifoDataN[127]), .Z(n655));
Q_AN02 U4621 ( .A0(n65), .A1(ofifoDataN[128]), .Z(n654));
Q_AN02 U4622 ( .A0(n65), .A1(ofifoDataN[129]), .Z(n653));
Q_AN02 U4623 ( .A0(n65), .A1(ofifoDataN[130]), .Z(n652));
Q_AN02 U4624 ( .A0(n65), .A1(ofifoDataN[131]), .Z(n651));
Q_AN02 U4625 ( .A0(n65), .A1(ofifoDataN[132]), .Z(n650));
Q_AN02 U4626 ( .A0(n65), .A1(ofifoDataN[133]), .Z(n649));
Q_AN02 U4627 ( .A0(n65), .A1(ofifoDataN[134]), .Z(n648));
Q_AN02 U4628 ( .A0(n65), .A1(ofifoDataN[135]), .Z(n647));
Q_AN02 U4629 ( .A0(n65), .A1(ofifoDataN[136]), .Z(n646));
Q_AN02 U4630 ( .A0(n65), .A1(ofifoDataN[137]), .Z(n645));
Q_AN02 U4631 ( .A0(n65), .A1(ofifoDataN[138]), .Z(n644));
Q_AN02 U4632 ( .A0(n65), .A1(ofifoDataN[139]), .Z(n643));
Q_AN02 U4633 ( .A0(n65), .A1(ofifoDataN[140]), .Z(n642));
Q_AN02 U4634 ( .A0(n65), .A1(ofifoDataN[141]), .Z(n641));
Q_AN02 U4635 ( .A0(n65), .A1(ofifoDataN[142]), .Z(n640));
Q_AN02 U4636 ( .A0(n65), .A1(ofifoDataN[143]), .Z(n639));
Q_AN02 U4637 ( .A0(n65), .A1(ofifoDataN[144]), .Z(n638));
Q_AN02 U4638 ( .A0(n65), .A1(ofifoDataN[145]), .Z(n637));
Q_AN02 U4639 ( .A0(n65), .A1(ofifoDataN[146]), .Z(n636));
Q_AN02 U4640 ( .A0(n65), .A1(ofifoDataN[147]), .Z(n635));
Q_AN02 U4641 ( .A0(n65), .A1(ofifoDataN[148]), .Z(n634));
Q_AN02 U4642 ( .A0(n65), .A1(ofifoDataN[149]), .Z(n633));
Q_AN02 U4643 ( .A0(n65), .A1(ofifoDataN[150]), .Z(n632));
Q_AN02 U4644 ( .A0(n65), .A1(ofifoDataN[151]), .Z(n631));
Q_AN02 U4645 ( .A0(n65), .A1(ofifoDataN[152]), .Z(n630));
Q_AN02 U4646 ( .A0(n65), .A1(ofifoDataN[153]), .Z(n629));
Q_AN02 U4647 ( .A0(n65), .A1(ofifoDataN[154]), .Z(n628));
Q_AN02 U4648 ( .A0(n65), .A1(ofifoDataN[155]), .Z(n627));
Q_AN02 U4649 ( .A0(n65), .A1(ofifoDataN[156]), .Z(n626));
Q_AN02 U4650 ( .A0(n65), .A1(ofifoDataN[157]), .Z(n625));
Q_AN02 U4651 ( .A0(n65), .A1(ofifoDataN[158]), .Z(n624));
Q_AN02 U4652 ( .A0(n65), .A1(ofifoDataN[159]), .Z(n623));
Q_AN02 U4653 ( .A0(n65), .A1(ofifoDataN[160]), .Z(n622));
Q_AN02 U4654 ( .A0(n65), .A1(ofifoDataN[161]), .Z(n621));
Q_AN02 U4655 ( .A0(n65), .A1(ofifoDataN[162]), .Z(n620));
Q_AN02 U4656 ( .A0(n65), .A1(ofifoDataN[163]), .Z(n619));
Q_AN02 U4657 ( .A0(n65), .A1(ofifoDataN[164]), .Z(n618));
Q_AN02 U4658 ( .A0(n65), .A1(ofifoDataN[165]), .Z(n617));
Q_AN02 U4659 ( .A0(n65), .A1(ofifoDataN[166]), .Z(n616));
Q_AN02 U4660 ( .A0(n65), .A1(ofifoDataN[167]), .Z(n615));
Q_AN02 U4661 ( .A0(n65), .A1(ofifoDataN[168]), .Z(n614));
Q_AN02 U4662 ( .A0(n65), .A1(ofifoDataN[169]), .Z(n613));
Q_AN02 U4663 ( .A0(n65), .A1(ofifoDataN[170]), .Z(n612));
Q_AN02 U4664 ( .A0(n65), .A1(ofifoDataN[171]), .Z(n611));
Q_AN02 U4665 ( .A0(n65), .A1(ofifoDataN[172]), .Z(n610));
Q_AN02 U4666 ( .A0(n65), .A1(ofifoDataN[173]), .Z(n609));
Q_AN02 U4667 ( .A0(n65), .A1(ofifoDataN[174]), .Z(n608));
Q_AN02 U4668 ( .A0(n65), .A1(ofifoDataN[175]), .Z(n607));
Q_AN02 U4669 ( .A0(n65), .A1(ofifoDataN[176]), .Z(n606));
Q_AN02 U4670 ( .A0(n65), .A1(ofifoDataN[177]), .Z(n605));
Q_AN02 U4671 ( .A0(n65), .A1(ofifoDataN[178]), .Z(n604));
Q_AN02 U4672 ( .A0(n65), .A1(ofifoDataN[179]), .Z(n603));
Q_AN02 U4673 ( .A0(n65), .A1(ofifoDataN[180]), .Z(n602));
Q_AN02 U4674 ( .A0(n65), .A1(ofifoDataN[181]), .Z(n601));
Q_AN02 U4675 ( .A0(n65), .A1(ofifoDataN[182]), .Z(n600));
Q_AN02 U4676 ( .A0(n65), .A1(ofifoDataN[183]), .Z(n599));
Q_AN02 U4677 ( .A0(n65), .A1(ofifoDataN[184]), .Z(n598));
Q_AN02 U4678 ( .A0(n65), .A1(ofifoDataN[185]), .Z(n597));
Q_AN02 U4679 ( .A0(n65), .A1(ofifoDataN[186]), .Z(n596));
Q_AN02 U4680 ( .A0(n65), .A1(ofifoDataN[187]), .Z(n595));
Q_AN02 U4681 ( .A0(n65), .A1(ofifoDataN[188]), .Z(n594));
Q_AN02 U4682 ( .A0(n65), .A1(ofifoDataN[189]), .Z(n593));
Q_AN02 U4683 ( .A0(n65), .A1(ofifoDataN[190]), .Z(n592));
Q_AN02 U4684 ( .A0(n65), .A1(ofifoDataN[191]), .Z(n591));
Q_AN02 U4685 ( .A0(n65), .A1(ofifoDataN[192]), .Z(n590));
Q_AN02 U4686 ( .A0(n65), .A1(ofifoDataN[193]), .Z(n589));
Q_AN02 U4687 ( .A0(n65), .A1(ofifoDataN[194]), .Z(n588));
Q_AN02 U4688 ( .A0(n65), .A1(ofifoDataN[195]), .Z(n587));
Q_AN02 U4689 ( .A0(n65), .A1(ofifoDataN[196]), .Z(n586));
Q_AN02 U4690 ( .A0(n65), .A1(ofifoDataN[197]), .Z(n585));
Q_AN02 U4691 ( .A0(n65), .A1(ofifoDataN[198]), .Z(n584));
Q_AN02 U4692 ( .A0(n65), .A1(ofifoDataN[199]), .Z(n583));
Q_AN02 U4693 ( .A0(n65), .A1(ofifoDataN[200]), .Z(n582));
Q_AN02 U4694 ( .A0(n65), .A1(ofifoDataN[201]), .Z(n581));
Q_AN02 U4695 ( .A0(n65), .A1(ofifoDataN[202]), .Z(n580));
Q_AN02 U4696 ( .A0(n65), .A1(ofifoDataN[203]), .Z(n579));
Q_AN02 U4697 ( .A0(n65), .A1(ofifoDataN[204]), .Z(n578));
Q_AN02 U4698 ( .A0(n65), .A1(ofifoDataN[205]), .Z(n577));
Q_AN02 U4699 ( .A0(n65), .A1(ofifoDataN[206]), .Z(n576));
Q_AN02 U4700 ( .A0(n65), .A1(ofifoDataN[207]), .Z(n575));
Q_AN02 U4701 ( .A0(n65), .A1(ofifoDataN[208]), .Z(n574));
Q_AN02 U4702 ( .A0(n65), .A1(ofifoDataN[209]), .Z(n573));
Q_AN02 U4703 ( .A0(n65), .A1(ofifoDataN[210]), .Z(n572));
Q_AN02 U4704 ( .A0(n65), .A1(ofifoDataN[211]), .Z(n571));
Q_AN02 U4705 ( .A0(n65), .A1(ofifoDataN[212]), .Z(n570));
Q_AN02 U4706 ( .A0(n65), .A1(ofifoDataN[213]), .Z(n569));
Q_AN02 U4707 ( .A0(n65), .A1(ofifoDataN[214]), .Z(n568));
Q_AN02 U4708 ( .A0(n65), .A1(ofifoDataN[215]), .Z(n567));
Q_AN02 U4709 ( .A0(n65), .A1(ofifoDataN[216]), .Z(n566));
Q_AN02 U4710 ( .A0(n65), .A1(ofifoDataN[217]), .Z(n565));
Q_AN02 U4711 ( .A0(n65), .A1(ofifoDataN[218]), .Z(n564));
Q_AN02 U4712 ( .A0(n65), .A1(ofifoDataN[219]), .Z(n563));
Q_AN02 U4713 ( .A0(n65), .A1(ofifoDataN[220]), .Z(n562));
Q_AN02 U4714 ( .A0(n65), .A1(ofifoDataN[221]), .Z(n561));
Q_AN02 U4715 ( .A0(n65), .A1(ofifoDataN[222]), .Z(n560));
Q_AN02 U4716 ( .A0(n65), .A1(ofifoDataN[223]), .Z(n559));
Q_AN02 U4717 ( .A0(n65), .A1(ofifoDataN[224]), .Z(n558));
Q_AN02 U4718 ( .A0(n65), .A1(ofifoDataN[225]), .Z(n557));
Q_AN02 U4719 ( .A0(n65), .A1(ofifoDataN[226]), .Z(n556));
Q_AN02 U4720 ( .A0(n65), .A1(ofifoDataN[227]), .Z(n555));
Q_AN02 U4721 ( .A0(n65), .A1(ofifoDataN[228]), .Z(n554));
Q_AN02 U4722 ( .A0(n65), .A1(ofifoDataN[229]), .Z(n553));
Q_AN02 U4723 ( .A0(n65), .A1(ofifoDataN[230]), .Z(n552));
Q_AN02 U4724 ( .A0(n65), .A1(ofifoDataN[231]), .Z(n551));
Q_AN02 U4725 ( .A0(n65), .A1(ofifoDataN[232]), .Z(n550));
Q_AN02 U4726 ( .A0(n65), .A1(ofifoDataN[233]), .Z(n549));
Q_AN02 U4727 ( .A0(n65), .A1(ofifoDataN[234]), .Z(n548));
Q_AN02 U4728 ( .A0(n65), .A1(ofifoDataN[235]), .Z(n547));
Q_AN02 U4729 ( .A0(n65), .A1(ofifoDataN[236]), .Z(n546));
Q_AN02 U4730 ( .A0(n65), .A1(ofifoDataN[237]), .Z(n545));
Q_AN02 U4731 ( .A0(n65), .A1(ofifoDataN[238]), .Z(n544));
Q_AN02 U4732 ( .A0(n65), .A1(ofifoDataN[239]), .Z(n543));
Q_AN02 U4733 ( .A0(n65), .A1(ofifoDataN[240]), .Z(n542));
Q_AN02 U4734 ( .A0(n65), .A1(ofifoDataN[241]), .Z(n541));
Q_AN02 U4735 ( .A0(n65), .A1(ofifoDataN[242]), .Z(n540));
Q_AN02 U4736 ( .A0(n65), .A1(ofifoDataN[243]), .Z(n539));
Q_AN02 U4737 ( .A0(n65), .A1(ofifoDataN[244]), .Z(n538));
Q_AN02 U4738 ( .A0(n65), .A1(ofifoDataN[245]), .Z(n537));
Q_AN02 U4739 ( .A0(n65), .A1(ofifoDataN[246]), .Z(n536));
Q_AN02 U4740 ( .A0(n65), .A1(ofifoDataN[247]), .Z(n535));
Q_AN02 U4741 ( .A0(n65), .A1(ofifoDataN[248]), .Z(n534));
Q_AN02 U4742 ( .A0(n65), .A1(ofifoDataN[249]), .Z(n533));
Q_AN02 U4743 ( .A0(n65), .A1(ofifoDataN[250]), .Z(n532));
Q_AN02 U4744 ( .A0(n65), .A1(ofifoDataN[251]), .Z(n531));
Q_AN02 U4745 ( .A0(n65), .A1(ofifoDataN[252]), .Z(n530));
Q_AN02 U4746 ( .A0(n65), .A1(ofifoDataN[253]), .Z(n529));
Q_AN02 U4747 ( .A0(n65), .A1(ofifoDataN[254]), .Z(n528));
Q_AN02 U4748 ( .A0(n65), .A1(ofifoDataN[255]), .Z(n527));
Q_AN02 U4749 ( .A0(n65), .A1(ofifoDataN[256]), .Z(n526));
Q_AN02 U4750 ( .A0(n65), .A1(ofifoDataN[257]), .Z(n525));
Q_AN02 U4751 ( .A0(n65), .A1(ofifoDataN[258]), .Z(n524));
Q_AN02 U4752 ( .A0(n65), .A1(ofifoDataN[259]), .Z(n523));
Q_AN02 U4753 ( .A0(n65), .A1(ofifoDataN[260]), .Z(n522));
Q_AN02 U4754 ( .A0(n65), .A1(ofifoDataN[261]), .Z(n521));
Q_AN02 U4755 ( .A0(n65), .A1(ofifoDataN[262]), .Z(n520));
Q_AN02 U4756 ( .A0(n65), .A1(ofifoDataN[263]), .Z(n519));
Q_AN02 U4757 ( .A0(n65), .A1(ofifoDataN[264]), .Z(n518));
Q_AN02 U4758 ( .A0(n65), .A1(ofifoDataN[265]), .Z(n517));
Q_AN02 U4759 ( .A0(n65), .A1(ofifoDataN[266]), .Z(n516));
Q_AN02 U4760 ( .A0(n65), .A1(ofifoDataN[267]), .Z(n515));
Q_AN02 U4761 ( .A0(n65), .A1(ofifoDataN[268]), .Z(n514));
Q_AN02 U4762 ( .A0(n65), .A1(ofifoDataN[269]), .Z(n513));
Q_AN02 U4763 ( .A0(n65), .A1(ofifoDataN[270]), .Z(n512));
Q_AN02 U4764 ( .A0(n65), .A1(ofifoDataN[271]), .Z(n511));
Q_AN02 U4765 ( .A0(n65), .A1(ofifoDataN[272]), .Z(n510));
Q_AN02 U4766 ( .A0(n65), .A1(ofifoDataN[273]), .Z(n509));
Q_AN02 U4767 ( .A0(n65), .A1(ofifoDataN[274]), .Z(n508));
Q_AN02 U4768 ( .A0(n65), .A1(ofifoDataN[275]), .Z(n507));
Q_AN02 U4769 ( .A0(n65), .A1(ofifoDataN[276]), .Z(n506));
Q_AN02 U4770 ( .A0(n65), .A1(ofifoDataN[277]), .Z(n505));
Q_AN02 U4771 ( .A0(n65), .A1(ofifoDataN[278]), .Z(n504));
Q_AN02 U4772 ( .A0(n65), .A1(ofifoDataN[279]), .Z(n503));
Q_AN02 U4773 ( .A0(n65), .A1(ofifoDataN[280]), .Z(n502));
Q_AN02 U4774 ( .A0(n65), .A1(ofifoDataN[281]), .Z(n501));
Q_AN02 U4775 ( .A0(n65), .A1(ofifoDataN[282]), .Z(n500));
Q_AN02 U4776 ( .A0(n65), .A1(ofifoDataN[283]), .Z(n499));
Q_AN02 U4777 ( .A0(n65), .A1(ofifoDataN[284]), .Z(n498));
Q_AN02 U4778 ( .A0(n65), .A1(ofifoDataN[285]), .Z(n497));
Q_AN02 U4779 ( .A0(n65), .A1(ofifoDataN[286]), .Z(n496));
Q_AN02 U4780 ( .A0(n65), .A1(ofifoDataN[287]), .Z(n495));
Q_AN02 U4781 ( .A0(n65), .A1(ofifoDataN[288]), .Z(n494));
Q_AN02 U4782 ( .A0(n65), .A1(ofifoDataN[289]), .Z(n493));
Q_AN02 U4783 ( .A0(n65), .A1(ofifoDataN[290]), .Z(n492));
Q_AN02 U4784 ( .A0(n65), .A1(ofifoDataN[291]), .Z(n491));
Q_AN02 U4785 ( .A0(n65), .A1(ofifoDataN[292]), .Z(n490));
Q_AN02 U4786 ( .A0(n65), .A1(ofifoDataN[293]), .Z(n489));
Q_AN02 U4787 ( .A0(n65), .A1(ofifoDataN[294]), .Z(n488));
Q_AN02 U4788 ( .A0(n65), .A1(ofifoDataN[295]), .Z(n487));
Q_AN02 U4789 ( .A0(n65), .A1(ofifoDataN[296]), .Z(n486));
Q_AN02 U4790 ( .A0(n65), .A1(ofifoDataN[297]), .Z(n485));
Q_AN02 U4791 ( .A0(n65), .A1(ofifoDataN[298]), .Z(n484));
Q_AN02 U4792 ( .A0(n65), .A1(ofifoDataN[299]), .Z(n483));
Q_AN02 U4793 ( .A0(n65), .A1(ofifoDataN[300]), .Z(n482));
Q_AN02 U4794 ( .A0(n65), .A1(ofifoDataN[301]), .Z(n481));
Q_AN02 U4795 ( .A0(n65), .A1(ofifoDataN[302]), .Z(n480));
Q_AN02 U4796 ( .A0(n65), .A1(ofifoDataN[303]), .Z(n479));
Q_AN02 U4797 ( .A0(n65), .A1(ofifoDataN[304]), .Z(n478));
Q_AN02 U4798 ( .A0(n65), .A1(ofifoDataN[305]), .Z(n477));
Q_AN02 U4799 ( .A0(n65), .A1(ofifoDataN[306]), .Z(n476));
Q_AN02 U4800 ( .A0(n65), .A1(ofifoDataN[307]), .Z(n475));
Q_AN02 U4801 ( .A0(n65), .A1(ofifoDataN[308]), .Z(n474));
Q_AN02 U4802 ( .A0(n65), .A1(ofifoDataN[309]), .Z(n473));
Q_AN02 U4803 ( .A0(n65), .A1(ofifoDataN[310]), .Z(n472));
Q_AN02 U4804 ( .A0(n65), .A1(ofifoDataN[311]), .Z(n471));
Q_AN02 U4805 ( .A0(n65), .A1(ofifoDataN[312]), .Z(n470));
Q_AN02 U4806 ( .A0(n65), .A1(ofifoDataN[313]), .Z(n469));
Q_AN02 U4807 ( .A0(n65), .A1(ofifoDataN[314]), .Z(n468));
Q_AN02 U4808 ( .A0(n65), .A1(ofifoDataN[315]), .Z(n467));
Q_AN02 U4809 ( .A0(n65), .A1(ofifoDataN[316]), .Z(n466));
Q_AN02 U4810 ( .A0(n65), .A1(ofifoDataN[317]), .Z(n465));
Q_AN02 U4811 ( .A0(n65), .A1(ofifoDataN[318]), .Z(n464));
Q_AN02 U4812 ( .A0(n65), .A1(ofifoDataN[319]), .Z(n463));
Q_AN02 U4813 ( .A0(n65), .A1(ofifoDataN[320]), .Z(n462));
Q_AN02 U4814 ( .A0(n65), .A1(ofifoDataN[321]), .Z(n461));
Q_AN02 U4815 ( .A0(n65), .A1(ofifoDataN[322]), .Z(n460));
Q_AN02 U4816 ( .A0(n65), .A1(ofifoDataN[323]), .Z(n459));
Q_AN02 U4817 ( .A0(n65), .A1(ofifoDataN[324]), .Z(n458));
Q_AN02 U4818 ( .A0(n65), .A1(ofifoDataN[325]), .Z(n457));
Q_AN02 U4819 ( .A0(n65), .A1(ofifoDataN[326]), .Z(n456));
Q_AN02 U4820 ( .A0(n65), .A1(ofifoDataN[327]), .Z(n455));
Q_AN02 U4821 ( .A0(n65), .A1(ofifoDataN[328]), .Z(n454));
Q_AN02 U4822 ( .A0(n65), .A1(ofifoDataN[329]), .Z(n453));
Q_AN02 U4823 ( .A0(n65), .A1(ofifoDataN[330]), .Z(n452));
Q_AN02 U4824 ( .A0(n65), .A1(ofifoDataN[331]), .Z(n451));
Q_AN02 U4825 ( .A0(n65), .A1(ofifoDataN[332]), .Z(n450));
Q_AN02 U4826 ( .A0(n65), .A1(ofifoDataN[333]), .Z(n449));
Q_AN02 U4827 ( .A0(n65), .A1(ofifoDataN[334]), .Z(n448));
Q_AN02 U4828 ( .A0(n65), .A1(ofifoDataN[335]), .Z(n447));
Q_AN02 U4829 ( .A0(n65), .A1(ofifoDataN[336]), .Z(n446));
Q_AN02 U4830 ( .A0(n65), .A1(ofifoDataN[337]), .Z(n445));
Q_AN02 U4831 ( .A0(n65), .A1(ofifoDataN[338]), .Z(n444));
Q_AN02 U4832 ( .A0(n65), .A1(ofifoDataN[339]), .Z(n443));
Q_AN02 U4833 ( .A0(n65), .A1(ofifoDataN[340]), .Z(n442));
Q_AN02 U4834 ( .A0(n65), .A1(ofifoDataN[341]), .Z(n441));
Q_AN02 U4835 ( .A0(n65), .A1(ofifoDataN[342]), .Z(n440));
Q_AN02 U4836 ( .A0(n65), .A1(ofifoDataN[343]), .Z(n439));
Q_AN02 U4837 ( .A0(n65), .A1(ofifoDataN[344]), .Z(n438));
Q_AN02 U4838 ( .A0(n65), .A1(ofifoDataN[345]), .Z(n437));
Q_AN02 U4839 ( .A0(n65), .A1(ofifoDataN[346]), .Z(n436));
Q_AN02 U4840 ( .A0(n65), .A1(ofifoDataN[347]), .Z(n435));
Q_AN02 U4841 ( .A0(n65), .A1(ofifoDataN[348]), .Z(n434));
Q_AN02 U4842 ( .A0(n65), .A1(ofifoDataN[349]), .Z(n433));
Q_AN02 U4843 ( .A0(n65), .A1(ofifoDataN[350]), .Z(n432));
Q_AN02 U4844 ( .A0(n65), .A1(ofifoDataN[351]), .Z(n431));
Q_AN02 U4845 ( .A0(n65), .A1(ofifoDataN[352]), .Z(n430));
Q_AN02 U4846 ( .A0(n65), .A1(ofifoDataN[353]), .Z(n429));
Q_AN02 U4847 ( .A0(n65), .A1(ofifoDataN[354]), .Z(n428));
Q_AN02 U4848 ( .A0(n65), .A1(ofifoDataN[355]), .Z(n427));
Q_AN02 U4849 ( .A0(n65), .A1(ofifoDataN[356]), .Z(n426));
Q_AN02 U4850 ( .A0(n65), .A1(ofifoDataN[357]), .Z(n425));
Q_AN02 U4851 ( .A0(n65), .A1(ofifoDataN[358]), .Z(n424));
Q_AN02 U4852 ( .A0(n65), .A1(ofifoDataN[359]), .Z(n423));
Q_AN02 U4853 ( .A0(n65), .A1(ofifoDataN[360]), .Z(n422));
Q_AN02 U4854 ( .A0(n65), .A1(ofifoDataN[361]), .Z(n421));
Q_AN02 U4855 ( .A0(n65), .A1(ofifoDataN[362]), .Z(n420));
Q_AN02 U4856 ( .A0(n65), .A1(ofifoDataN[363]), .Z(n419));
Q_AN02 U4857 ( .A0(n65), .A1(ofifoDataN[364]), .Z(n418));
Q_AN02 U4858 ( .A0(n65), .A1(ofifoDataN[365]), .Z(n417));
Q_AN02 U4859 ( .A0(n65), .A1(ofifoDataN[366]), .Z(n416));
Q_AN02 U4860 ( .A0(n65), .A1(ofifoDataN[367]), .Z(n415));
Q_AN02 U4861 ( .A0(n65), .A1(ofifoDataN[368]), .Z(n414));
Q_AN02 U4862 ( .A0(n65), .A1(ofifoDataN[369]), .Z(n413));
Q_AN02 U4863 ( .A0(n65), .A1(ofifoDataN[370]), .Z(n412));
Q_AN02 U4864 ( .A0(n65), .A1(ofifoDataN[371]), .Z(n411));
Q_AN02 U4865 ( .A0(n65), .A1(ofifoDataN[372]), .Z(n410));
Q_AN02 U4866 ( .A0(n65), .A1(ofifoDataN[373]), .Z(n409));
Q_AN02 U4867 ( .A0(n65), .A1(ofifoDataN[374]), .Z(n408));
Q_AN02 U4868 ( .A0(n65), .A1(ofifoDataN[375]), .Z(n407));
Q_AN02 U4869 ( .A0(n65), .A1(ofifoDataN[376]), .Z(n406));
Q_AN02 U4870 ( .A0(n65), .A1(ofifoDataN[377]), .Z(n405));
Q_AN02 U4871 ( .A0(n65), .A1(ofifoDataN[378]), .Z(n404));
Q_AN02 U4872 ( .A0(n65), .A1(ofifoDataN[379]), .Z(n403));
Q_AN02 U4873 ( .A0(n65), .A1(ofifoDataN[380]), .Z(n402));
Q_AN02 U4874 ( .A0(n65), .A1(ofifoDataN[381]), .Z(n401));
Q_AN02 U4875 ( .A0(n65), .A1(ofifoDataN[382]), .Z(n400));
Q_AN02 U4876 ( .A0(n65), .A1(ofifoDataN[383]), .Z(n399));
Q_AN02 U4877 ( .A0(n65), .A1(ofifoDataN[384]), .Z(n398));
Q_AN02 U4878 ( .A0(n65), .A1(ofifoDataN[385]), .Z(n397));
Q_AN02 U4879 ( .A0(n65), .A1(ofifoDataN[386]), .Z(n396));
Q_AN02 U4880 ( .A0(n65), .A1(ofifoDataN[387]), .Z(n395));
Q_AN02 U4881 ( .A0(n65), .A1(ofifoDataN[388]), .Z(n394));
Q_AN02 U4882 ( .A0(n65), .A1(ofifoDataN[389]), .Z(n393));
Q_AN02 U4883 ( .A0(n65), .A1(ofifoDataN[390]), .Z(n392));
Q_AN02 U4884 ( .A0(n65), .A1(ofifoDataN[391]), .Z(n391));
Q_AN02 U4885 ( .A0(n65), .A1(ofifoDataN[392]), .Z(n390));
Q_AN02 U4886 ( .A0(n65), .A1(ofifoDataN[393]), .Z(n389));
Q_AN02 U4887 ( .A0(n65), .A1(ofifoDataN[394]), .Z(n388));
Q_AN02 U4888 ( .A0(n65), .A1(ofifoDataN[395]), .Z(n387));
Q_AN02 U4889 ( .A0(n65), .A1(ofifoDataN[396]), .Z(n386));
Q_AN02 U4890 ( .A0(n65), .A1(ofifoDataN[397]), .Z(n385));
Q_AN02 U4891 ( .A0(n65), .A1(ofifoDataN[398]), .Z(n384));
Q_AN02 U4892 ( .A0(n65), .A1(ofifoDataN[399]), .Z(n383));
Q_AN02 U4893 ( .A0(n65), .A1(ofifoDataN[400]), .Z(n382));
Q_AN02 U4894 ( .A0(n65), .A1(ofifoDataN[401]), .Z(n381));
Q_AN02 U4895 ( .A0(n65), .A1(ofifoDataN[402]), .Z(n380));
Q_AN02 U4896 ( .A0(n65), .A1(ofifoDataN[403]), .Z(n379));
Q_AN02 U4897 ( .A0(n65), .A1(ofifoDataN[404]), .Z(n378));
Q_AN02 U4898 ( .A0(n65), .A1(ofifoDataN[405]), .Z(n377));
Q_AN02 U4899 ( .A0(n65), .A1(ofifoDataN[406]), .Z(n376));
Q_AN02 U4900 ( .A0(n65), .A1(ofifoDataN[407]), .Z(n375));
Q_AN02 U4901 ( .A0(n65), .A1(ofifoDataN[408]), .Z(n374));
Q_AN02 U4902 ( .A0(n65), .A1(ofifoDataN[409]), .Z(n373));
Q_AN02 U4903 ( .A0(n65), .A1(ofifoDataN[410]), .Z(n372));
Q_AN02 U4904 ( .A0(n65), .A1(ofifoDataN[411]), .Z(n371));
Q_AN02 U4905 ( .A0(n65), .A1(ofifoDataN[412]), .Z(n370));
Q_AN02 U4906 ( .A0(n65), .A1(ofifoDataN[413]), .Z(n369));
Q_AN02 U4907 ( .A0(n65), .A1(ofifoDataN[414]), .Z(n368));
Q_AN02 U4908 ( .A0(n65), .A1(ofifoDataN[415]), .Z(n367));
Q_AN02 U4909 ( .A0(n65), .A1(ofifoDataN[416]), .Z(n366));
Q_AN02 U4910 ( .A0(n65), .A1(ofifoDataN[417]), .Z(n365));
Q_AN02 U4911 ( .A0(n65), .A1(ofifoDataN[418]), .Z(n364));
Q_AN02 U4912 ( .A0(n65), .A1(ofifoDataN[419]), .Z(n363));
Q_AN02 U4913 ( .A0(n65), .A1(ofifoDataN[420]), .Z(n362));
Q_AN02 U4914 ( .A0(n65), .A1(ofifoDataN[421]), .Z(n361));
Q_AN02 U4915 ( .A0(n65), .A1(ofifoDataN[422]), .Z(n360));
Q_AN02 U4916 ( .A0(n65), .A1(ofifoDataN[423]), .Z(n359));
Q_AN02 U4917 ( .A0(n65), .A1(ofifoDataN[424]), .Z(n358));
Q_AN02 U4918 ( .A0(n65), .A1(ofifoDataN[425]), .Z(n357));
Q_AN02 U4919 ( .A0(n65), .A1(ofifoDataN[426]), .Z(n356));
Q_AN02 U4920 ( .A0(n65), .A1(ofifoDataN[427]), .Z(n355));
Q_AN02 U4921 ( .A0(n65), .A1(ofifoDataN[428]), .Z(n354));
Q_AN02 U4922 ( .A0(n65), .A1(ofifoDataN[429]), .Z(n353));
Q_AN02 U4923 ( .A0(n65), .A1(ofifoDataN[430]), .Z(n352));
Q_AN02 U4924 ( .A0(n65), .A1(ofifoDataN[431]), .Z(n351));
Q_AN02 U4925 ( .A0(n65), .A1(ofifoDataN[432]), .Z(n350));
Q_AN02 U4926 ( .A0(n65), .A1(ofifoDataN[433]), .Z(n349));
Q_AN02 U4927 ( .A0(n65), .A1(ofifoDataN[434]), .Z(n348));
Q_AN02 U4928 ( .A0(n65), .A1(ofifoDataN[435]), .Z(n347));
Q_AN02 U4929 ( .A0(n65), .A1(ofifoDataN[436]), .Z(n346));
Q_AN02 U4930 ( .A0(n65), .A1(ofifoDataN[437]), .Z(n345));
Q_AN02 U4931 ( .A0(n65), .A1(ofifoDataN[438]), .Z(n344));
Q_AN02 U4932 ( .A0(n65), .A1(ofifoDataN[439]), .Z(n343));
Q_AN02 U4933 ( .A0(n65), .A1(ofifoDataN[440]), .Z(n342));
Q_AN02 U4934 ( .A0(n65), .A1(ofifoDataN[441]), .Z(n341));
Q_AN02 U4935 ( .A0(n65), .A1(ofifoDataN[442]), .Z(n340));
Q_AN02 U4936 ( .A0(n65), .A1(ofifoDataN[443]), .Z(n339));
Q_AN02 U4937 ( .A0(n65), .A1(ofifoDataN[444]), .Z(n338));
Q_AN02 U4938 ( .A0(n65), .A1(ofifoDataN[445]), .Z(n337));
Q_AN02 U4939 ( .A0(n65), .A1(ofifoDataN[446]), .Z(n336));
Q_AN02 U4940 ( .A0(n65), .A1(ofifoDataN[447]), .Z(n335));
Q_AN02 U4941 ( .A0(n65), .A1(ofifoDataN[448]), .Z(n334));
Q_AN02 U4942 ( .A0(n65), .A1(ofifoDataN[449]), .Z(n333));
Q_AN02 U4943 ( .A0(n65), .A1(ofifoDataN[450]), .Z(n332));
Q_AN02 U4944 ( .A0(n65), .A1(ofifoDataN[451]), .Z(n331));
Q_AN02 U4945 ( .A0(n65), .A1(ofifoDataN[452]), .Z(n330));
Q_AN02 U4946 ( .A0(n65), .A1(ofifoDataN[453]), .Z(n329));
Q_AN02 U4947 ( .A0(n65), .A1(ofifoDataN[454]), .Z(n328));
Q_AN02 U4948 ( .A0(n65), .A1(ofifoDataN[455]), .Z(n327));
Q_AN02 U4949 ( .A0(n65), .A1(ofifoDataN[456]), .Z(n326));
Q_AN02 U4950 ( .A0(n65), .A1(ofifoDataN[457]), .Z(n325));
Q_AN02 U4951 ( .A0(n65), .A1(ofifoDataN[458]), .Z(n324));
Q_AN02 U4952 ( .A0(n65), .A1(ofifoDataN[459]), .Z(n323));
Q_AN02 U4953 ( .A0(n65), .A1(ofifoDataN[460]), .Z(n322));
Q_AN02 U4954 ( .A0(n65), .A1(ofifoDataN[461]), .Z(n321));
Q_AN02 U4955 ( .A0(n65), .A1(ofifoDataN[462]), .Z(n320));
Q_AN02 U4956 ( .A0(n65), .A1(ofifoDataN[463]), .Z(n319));
Q_AN02 U4957 ( .A0(n65), .A1(ofifoDataN[464]), .Z(n318));
Q_AN02 U4958 ( .A0(n65), .A1(ofifoDataN[465]), .Z(n317));
Q_AN02 U4959 ( .A0(n65), .A1(ofifoDataN[466]), .Z(n316));
Q_AN02 U4960 ( .A0(n65), .A1(ofifoDataN[467]), .Z(n315));
Q_AN02 U4961 ( .A0(n65), .A1(ofifoDataN[468]), .Z(n314));
Q_AN02 U4962 ( .A0(n65), .A1(ofifoDataN[469]), .Z(n313));
Q_AN02 U4963 ( .A0(n65), .A1(ofifoDataN[470]), .Z(n312));
Q_AN02 U4964 ( .A0(n65), .A1(ofifoDataN[471]), .Z(n311));
Q_AN02 U4965 ( .A0(n65), .A1(ofifoDataN[472]), .Z(n310));
Q_AN02 U4966 ( .A0(n65), .A1(ofifoDataN[473]), .Z(n309));
Q_AN02 U4967 ( .A0(n65), .A1(ofifoDataN[474]), .Z(n308));
Q_AN02 U4968 ( .A0(n65), .A1(ofifoDataN[475]), .Z(n307));
Q_AN02 U4969 ( .A0(n65), .A1(ofifoDataN[476]), .Z(n306));
Q_AN02 U4970 ( .A0(n65), .A1(ofifoDataN[477]), .Z(n305));
Q_AN02 U4971 ( .A0(n65), .A1(ofifoDataN[478]), .Z(n304));
Q_AN02 U4972 ( .A0(n65), .A1(ofifoDataN[479]), .Z(n303));
Q_AN02 U4973 ( .A0(n65), .A1(ofifoDataN[480]), .Z(n302));
Q_AN02 U4974 ( .A0(n65), .A1(ofifoDataN[481]), .Z(n301));
Q_AN02 U4975 ( .A0(n65), .A1(ofifoDataN[482]), .Z(n300));
Q_AN02 U4976 ( .A0(n65), .A1(ofifoDataN[483]), .Z(n299));
Q_AN02 U4977 ( .A0(n65), .A1(ofifoDataN[484]), .Z(n298));
Q_AN02 U4978 ( .A0(n65), .A1(ofifoDataN[485]), .Z(n297));
Q_AN02 U4979 ( .A0(n65), .A1(ofifoDataN[486]), .Z(n296));
Q_AN02 U4980 ( .A0(n65), .A1(ofifoDataN[487]), .Z(n295));
Q_AN02 U4981 ( .A0(n65), .A1(ofifoDataN[488]), .Z(n294));
Q_AN02 U4982 ( .A0(n65), .A1(ofifoDataN[489]), .Z(n293));
Q_AN02 U4983 ( .A0(n65), .A1(ofifoDataN[490]), .Z(n292));
Q_AN02 U4984 ( .A0(n65), .A1(ofifoDataN[491]), .Z(n291));
Q_AN02 U4985 ( .A0(n65), .A1(ofifoDataN[492]), .Z(n290));
Q_AN02 U4986 ( .A0(n65), .A1(ofifoDataN[493]), .Z(n289));
Q_AN02 U4987 ( .A0(n65), .A1(ofifoDataN[494]), .Z(n288));
Q_AN02 U4988 ( .A0(n65), .A1(ofifoDataN[495]), .Z(n287));
Q_AN02 U4989 ( .A0(n65), .A1(ofifoDataN[496]), .Z(n286));
Q_AN02 U4990 ( .A0(n65), .A1(ofifoDataN[497]), .Z(n285));
Q_AN02 U4991 ( .A0(n65), .A1(ofifoDataN[498]), .Z(n284));
Q_AN02 U4992 ( .A0(n65), .A1(ofifoDataN[499]), .Z(n283));
Q_AN02 U4993 ( .A0(n65), .A1(ofifoDataN[500]), .Z(n282));
Q_AN02 U4994 ( .A0(n65), .A1(ofifoDataN[501]), .Z(n281));
Q_AN02 U4995 ( .A0(n65), .A1(ofifoDataN[502]), .Z(n280));
Q_AN02 U4996 ( .A0(n65), .A1(ofifoDataN[503]), .Z(n279));
Q_AN02 U4997 ( .A0(n65), .A1(ofifoDataN[504]), .Z(n278));
Q_AN02 U4998 ( .A0(n65), .A1(ofifoDataN[505]), .Z(n277));
Q_AN02 U4999 ( .A0(n65), .A1(ofifoDataN[506]), .Z(n276));
Q_AN02 U5000 ( .A0(n65), .A1(ofifoDataN[507]), .Z(n275));
Q_AN02 U5001 ( .A0(n65), .A1(ofifoDataN[508]), .Z(n274));
Q_AN02 U5002 ( .A0(n65), .A1(ofifoDataN[509]), .Z(n273));
Q_AN02 U5003 ( .A0(n65), .A1(ofifoDataN[510]), .Z(n272));
Q_AN02 U5004 ( .A0(n65), .A1(ofifoDataN[511]), .Z(n271));
Q_AN02 U5005 ( .A0(n65), .A1(ofifoDataN[512]), .Z(n270));
Q_AN02 U5006 ( .A0(n65), .A1(ofifoDataN[513]), .Z(n269));
Q_AN02 U5007 ( .A0(n65), .A1(ofifoDataN[514]), .Z(n268));
Q_AN02 U5008 ( .A0(n65), .A1(ofifoDataN[515]), .Z(n267));
Q_AN02 U5009 ( .A0(n65), .A1(ofifoDataN[516]), .Z(n266));
Q_AN02 U5010 ( .A0(n65), .A1(ofifoDataN[517]), .Z(n265));
Q_AN02 U5011 ( .A0(n65), .A1(ofifoDataN[518]), .Z(n264));
Q_AN02 U5012 ( .A0(n65), .A1(ofifoDataN[519]), .Z(n263));
Q_AN02 U5013 ( .A0(n65), .A1(ofifoDataN[520]), .Z(n262));
Q_AN02 U5014 ( .A0(n65), .A1(ofifoDataN[521]), .Z(n261));
Q_AN02 U5015 ( .A0(n65), .A1(ofifoDataN[522]), .Z(n260));
Q_AN02 U5016 ( .A0(n65), .A1(ofifoDataN[523]), .Z(n259));
Q_AN02 U5017 ( .A0(n65), .A1(ofifoDataN[524]), .Z(n258));
Q_AN02 U5018 ( .A0(n65), .A1(ofifoDataN[525]), .Z(n257));
Q_AN02 U5019 ( .A0(n65), .A1(ofifoDataN[526]), .Z(n256));
Q_AN02 U5020 ( .A0(n65), .A1(ofifoDataN[527]), .Z(n255));
Q_AN02 U5021 ( .A0(n65), .A1(ofifoDataN[528]), .Z(n254));
Q_AN02 U5022 ( .A0(n65), .A1(ofifoDataN[529]), .Z(n253));
Q_AN02 U5023 ( .A0(n65), .A1(ofifoDataN[530]), .Z(n252));
Q_AN02 U5024 ( .A0(n65), .A1(ofifoDataN[531]), .Z(n251));
Q_AN02 U5025 ( .A0(n65), .A1(ofifoDataN[532]), .Z(n250));
Q_AN02 U5026 ( .A0(n65), .A1(ofifoDataN[533]), .Z(n249));
Q_AN02 U5027 ( .A0(n65), .A1(ofifoDataN[534]), .Z(n248));
Q_AN02 U5028 ( .A0(n65), .A1(ofifoDataN[535]), .Z(n247));
Q_AN02 U5029 ( .A0(n65), .A1(ofifoDataN[536]), .Z(n246));
Q_AN02 U5030 ( .A0(n65), .A1(ofifoDataN[537]), .Z(n245));
Q_AN02 U5031 ( .A0(n65), .A1(ofifoDataN[538]), .Z(n244));
Q_AN02 U5032 ( .A0(n65), .A1(ofifoDataN[539]), .Z(n243));
Q_AN02 U5033 ( .A0(n65), .A1(ofifoDataN[540]), .Z(n242));
Q_AN02 U5034 ( .A0(n65), .A1(ofifoDataN[541]), .Z(n241));
Q_AN02 U5035 ( .A0(n65), .A1(ofifoDataN[542]), .Z(n240));
Q_AN02 U5036 ( .A0(n65), .A1(ofifoDataN[543]), .Z(n239));
Q_AN02 U5037 ( .A0(n65), .A1(ofifoDataN[544]), .Z(n238));
Q_AN02 U5038 ( .A0(n65), .A1(ofifoDataN[545]), .Z(n237));
Q_AN02 U5039 ( .A0(n65), .A1(ofifoDataN[546]), .Z(n236));
Q_AN02 U5040 ( .A0(n65), .A1(ofifoDataN[547]), .Z(n235));
Q_AN02 U5041 ( .A0(n65), .A1(ofifoDataN[548]), .Z(n234));
Q_AN02 U5042 ( .A0(n65), .A1(ofifoDataN[549]), .Z(n233));
Q_AN02 U5043 ( .A0(n65), .A1(ofifoDataN[550]), .Z(n232));
Q_AN02 U5044 ( .A0(n65), .A1(ofifoDataN[551]), .Z(n231));
Q_AN02 U5045 ( .A0(n65), .A1(ofifoDataN[552]), .Z(n230));
Q_AN02 U5046 ( .A0(n65), .A1(ofifoDataN[553]), .Z(n229));
Q_AN02 U5047 ( .A0(n65), .A1(ofifoDataN[554]), .Z(n228));
Q_AN02 U5048 ( .A0(n65), .A1(ofifoDataN[555]), .Z(n227));
Q_AN02 U5049 ( .A0(n65), .A1(ofifoDataN[556]), .Z(n226));
Q_AN02 U5050 ( .A0(n65), .A1(ofifoDataN[557]), .Z(n225));
Q_AN02 U5051 ( .A0(n65), .A1(ofifoDataN[558]), .Z(n224));
Q_AN02 U5052 ( .A0(n65), .A1(ofifoDataN[559]), .Z(n223));
Q_AN02 U5053 ( .A0(n65), .A1(ofifoDataN[560]), .Z(n222));
Q_AN02 U5054 ( .A0(n65), .A1(ofifoDataN[561]), .Z(n221));
Q_AN02 U5055 ( .A0(n65), .A1(ofifoDataN[562]), .Z(n220));
Q_AN02 U5056 ( .A0(n65), .A1(ofifoDataN[563]), .Z(n219));
Q_AN02 U5057 ( .A0(n65), .A1(ofifoDataN[564]), .Z(n218));
Q_AN02 U5058 ( .A0(n65), .A1(ofifoDataN[565]), .Z(n217));
Q_AN02 U5059 ( .A0(n65), .A1(ofifoDataN[566]), .Z(n216));
Q_AN02 U5060 ( .A0(n65), .A1(ofifoDataN[567]), .Z(n215));
Q_AN02 U5061 ( .A0(n65), .A1(ofifoDataN[568]), .Z(n214));
Q_AN02 U5062 ( .A0(n65), .A1(ofifoDataN[569]), .Z(n213));
Q_AN02 U5063 ( .A0(n65), .A1(ofifoDataN[570]), .Z(n212));
Q_AN02 U5064 ( .A0(n65), .A1(ofifoDataN[571]), .Z(n211));
Q_AN02 U5065 ( .A0(n65), .A1(ofifoDataN[572]), .Z(n210));
Q_AN02 U5066 ( .A0(n65), .A1(ofifoDataN[573]), .Z(n209));
Q_AN02 U5067 ( .A0(n65), .A1(ofifoDataN[574]), .Z(n208));
Q_AN02 U5068 ( .A0(n65), .A1(ofifoDataN[575]), .Z(n207));
Q_AN02 U5069 ( .A0(n65), .A1(ofifoWptrN[0]), .Z(n206));
Q_AN02 U5070 ( .A0(n65), .A1(ofifoWptrN[1]), .Z(n205));
Q_AN02 U5071 ( .A0(n65), .A1(ofifoWptrN[2]), .Z(n204));
Q_AN02 U5072 ( .A0(n65), .A1(ofifoWptrN[3]), .Z(n203));
Q_AN02 U5073 ( .A0(n65), .A1(ofifoWptrN[4]), .Z(n202));
Q_AN02 U5074 ( .A0(n65), .A1(ofifoWptrN[5]), .Z(n201));
Q_AN02 U5075 ( .A0(n65), .A1(ofifoWptrN[6]), .Z(n200));
Q_AN02 U5076 ( .A0(n65), .A1(ofifoWptrN[7]), .Z(n199));
Q_AN02 U5077 ( .A0(n65), .A1(ofifoWptrN[8]), .Z(n198));
Q_AN02 U5078 ( .A0(n65), .A1(ofifoWptrN[9]), .Z(n197));
Q_AN02 U5079 ( .A0(n65), .A1(ofifoWptrN[10]), .Z(n196));
Q_AN02 U5080 ( .A0(n65), .A1(ofifoWptrN[11]), .Z(n195));
Q_AN02 U5081 ( .A0(n65), .A1(ofifoWptrN[12]), .Z(n194));
Q_AN02 U5082 ( .A0(n65), .A1(ofifoWptrN[13]), .Z(n193));
Q_AN02 U5083 ( .A0(n65), .A1(ofifoWptrN[14]), .Z(n192));
Q_AN02 U5084 ( .A0(n65), .A1(ofifoWptrN[15]), .Z(n191));
Q_AN02 U5085 ( .A0(n65), .A1(ofifoWptrN[16]), .Z(n190));
Q_AN02 U5086 ( .A0(n65), .A1(oFillN[0]), .Z(n189));
Q_AN02 U5087 ( .A0(n65), .A1(oFillN[1]), .Z(n188));
Q_AN02 U5088 ( .A0(n65), .A1(oFillN[2]), .Z(n187));
Q_AN02 U5089 ( .A0(n65), .A1(oFillN[3]), .Z(n186));
Q_AN02 U5090 ( .A0(n65), .A1(oFillN[4]), .Z(n185));
Q_AN02 U5091 ( .A0(n65), .A1(ofifoAddr8N[4]), .Z(n184));
Q_AN02 U5092 ( .A0(n65), .A1(ofifoAddr8N[5]), .Z(n183));
Q_AN02 U5093 ( .A0(n65), .A1(ofifoAddr8N[6]), .Z(n182));
Q_AN02 U5094 ( .A0(n65), .A1(ofifoAddr8N[7]), .Z(n181));
Q_AN02 U5095 ( .A0(n65), .A1(ofifoAddr8N[8]), .Z(n180));
Q_AN02 U5096 ( .A0(n65), .A1(ofifoAddr8N[9]), .Z(n179));
Q_AN02 U5097 ( .A0(n65), .A1(ofifoAddr8N[10]), .Z(n178));
Q_AN02 U5098 ( .A0(n65), .A1(ofifoAddr8N[11]), .Z(n177));
Q_AN02 U5099 ( .A0(n65), .A1(ofifoAddr8N[12]), .Z(n176));
Q_AN02 U5100 ( .A0(n65), .A1(ofifoAddr8N[13]), .Z(n175));
Q_AN02 U5101 ( .A0(n65), .A1(ofifoAddr8N[14]), .Z(n174));
Q_AN02 U5102 ( .A0(n65), .A1(ofifoAddr8N[15]), .Z(n173));
Q_AN02 U5103 ( .A0(n65), .A1(ofifoAddr8N[16]), .Z(n172));
Q_OR02 U5104 ( .A0(xc_top.GFReset), .A1(ofifoAddr7N[2]), .Z(n171));
Q_AN02 U5105 ( .A0(n65), .A1(ofifoAddr7N[3]), .Z(n170));
Q_AN02 U5106 ( .A0(n65), .A1(ofifoAddr7N[4]), .Z(n169));
Q_AN02 U5107 ( .A0(n65), .A1(ofifoAddr7N[5]), .Z(n168));
Q_AN02 U5108 ( .A0(n65), .A1(ofifoAddr7N[6]), .Z(n167));
Q_AN02 U5109 ( .A0(n65), .A1(ofifoAddr7N[7]), .Z(n166));
Q_AN02 U5110 ( .A0(n65), .A1(ofifoAddr7N[8]), .Z(n165));
Q_AN02 U5111 ( .A0(n65), .A1(ofifoAddr7N[9]), .Z(n164));
Q_AN02 U5112 ( .A0(n65), .A1(ofifoAddr7N[10]), .Z(n163));
Q_AN02 U5113 ( .A0(n65), .A1(ofifoAddr7N[11]), .Z(n162));
Q_AN02 U5114 ( .A0(n65), .A1(ofifoAddr7N[12]), .Z(n161));
Q_AN02 U5115 ( .A0(n65), .A1(ofifoAddr7N[13]), .Z(n160));
Q_AN02 U5116 ( .A0(n65), .A1(ofifoAddr7N[14]), .Z(n159));
Q_AN02 U5117 ( .A0(n65), .A1(ofifoAddr7N[15]), .Z(n158));
Q_AN02 U5118 ( .A0(n65), .A1(ofifoAddr7N[16]), .Z(n157));
Q_AN02 U5119 ( .A0(n65), .A1(ofifoAddr6N[3]), .Z(n156));
Q_AN02 U5120 ( .A0(n65), .A1(ofifoAddr6N[4]), .Z(n155));
Q_AN02 U5121 ( .A0(n65), .A1(ofifoAddr6N[5]), .Z(n154));
Q_AN02 U5122 ( .A0(n65), .A1(ofifoAddr6N[6]), .Z(n153));
Q_AN02 U5123 ( .A0(n65), .A1(ofifoAddr6N[7]), .Z(n152));
Q_AN02 U5124 ( .A0(n65), .A1(ofifoAddr6N[8]), .Z(n151));
Q_AN02 U5125 ( .A0(n65), .A1(ofifoAddr6N[9]), .Z(n150));
Q_AN02 U5126 ( .A0(n65), .A1(ofifoAddr6N[10]), .Z(n149));
Q_AN02 U5127 ( .A0(n65), .A1(ofifoAddr6N[11]), .Z(n148));
Q_AN02 U5128 ( .A0(n65), .A1(ofifoAddr6N[12]), .Z(n147));
Q_AN02 U5129 ( .A0(n65), .A1(ofifoAddr6N[13]), .Z(n146));
Q_AN02 U5130 ( .A0(n65), .A1(ofifoAddr6N[14]), .Z(n145));
Q_AN02 U5131 ( .A0(n65), .A1(ofifoAddr6N[15]), .Z(n144));
Q_AN02 U5132 ( .A0(n65), .A1(ofifoAddr6N[16]), .Z(n143));
Q_AN02 U5133 ( .A0(n65), .A1(ofifoAddr5N[3]), .Z(n142));
Q_AN02 U5134 ( .A0(n65), .A1(ofifoAddr5N[4]), .Z(n141));
Q_AN02 U5135 ( .A0(n65), .A1(ofifoAddr5N[5]), .Z(n140));
Q_AN02 U5136 ( .A0(n65), .A1(ofifoAddr5N[6]), .Z(n139));
Q_AN02 U5137 ( .A0(n65), .A1(ofifoAddr5N[7]), .Z(n138));
Q_AN02 U5138 ( .A0(n65), .A1(ofifoAddr5N[8]), .Z(n137));
Q_AN02 U5139 ( .A0(n65), .A1(ofifoAddr5N[9]), .Z(n136));
Q_AN02 U5140 ( .A0(n65), .A1(ofifoAddr5N[10]), .Z(n135));
Q_AN02 U5141 ( .A0(n65), .A1(ofifoAddr5N[11]), .Z(n134));
Q_AN02 U5142 ( .A0(n65), .A1(ofifoAddr5N[12]), .Z(n133));
Q_AN02 U5143 ( .A0(n65), .A1(ofifoAddr5N[13]), .Z(n132));
Q_AN02 U5144 ( .A0(n65), .A1(ofifoAddr5N[14]), .Z(n131));
Q_AN02 U5145 ( .A0(n65), .A1(ofifoAddr5N[15]), .Z(n130));
Q_AN02 U5146 ( .A0(n65), .A1(ofifoAddr5N[16]), .Z(n129));
Q_AN02 U5147 ( .A0(n65), .A1(ofifoAddr4N[3]), .Z(n128));
Q_AN02 U5148 ( .A0(n65), .A1(ofifoAddr4N[4]), .Z(n127));
Q_AN02 U5149 ( .A0(n65), .A1(ofifoAddr4N[5]), .Z(n126));
Q_AN02 U5150 ( .A0(n65), .A1(ofifoAddr4N[6]), .Z(n125));
Q_AN02 U5151 ( .A0(n65), .A1(ofifoAddr4N[7]), .Z(n124));
Q_AN02 U5152 ( .A0(n65), .A1(ofifoAddr4N[8]), .Z(n123));
Q_AN02 U5153 ( .A0(n65), .A1(ofifoAddr4N[9]), .Z(n122));
Q_AN02 U5154 ( .A0(n65), .A1(ofifoAddr4N[10]), .Z(n121));
Q_AN02 U5155 ( .A0(n65), .A1(ofifoAddr4N[11]), .Z(n120));
Q_AN02 U5156 ( .A0(n65), .A1(ofifoAddr4N[12]), .Z(n119));
Q_AN02 U5157 ( .A0(n65), .A1(ofifoAddr4N[13]), .Z(n118));
Q_AN02 U5158 ( .A0(n65), .A1(ofifoAddr4N[14]), .Z(n117));
Q_AN02 U5159 ( .A0(n65), .A1(ofifoAddr4N[15]), .Z(n116));
Q_AN02 U5160 ( .A0(n65), .A1(ofifoAddr4N[16]), .Z(n115));
Q_OR02 U5161 ( .A0(xc_top.GFReset), .A1(ofifoAddr0N[0]), .Z(n114));
Q_NR02 U5162 ( .A0(xc_top.GFReset), .A1(ofifoAddr6N[2]), .Z(n113));
Q_AN02 U5163 ( .A0(n65), .A1(ofifoAddr2N[3]), .Z(n112));
Q_AN02 U5164 ( .A0(n65), .A1(ofifoAddr2N[4]), .Z(n111));
Q_AN02 U5165 ( .A0(n65), .A1(ofifoAddr2N[5]), .Z(n110));
Q_AN02 U5166 ( .A0(n65), .A1(ofifoAddr2N[6]), .Z(n109));
Q_AN02 U5167 ( .A0(n65), .A1(ofifoAddr2N[7]), .Z(n108));
Q_AN02 U5168 ( .A0(n65), .A1(ofifoAddr2N[8]), .Z(n107));
Q_AN02 U5169 ( .A0(n65), .A1(ofifoAddr2N[9]), .Z(n106));
Q_AN02 U5170 ( .A0(n65), .A1(ofifoAddr2N[10]), .Z(n105));
Q_AN02 U5171 ( .A0(n65), .A1(ofifoAddr2N[11]), .Z(n104));
Q_AN02 U5172 ( .A0(n65), .A1(ofifoAddr2N[12]), .Z(n103));
Q_AN02 U5173 ( .A0(n65), .A1(ofifoAddr2N[13]), .Z(n102));
Q_AN02 U5174 ( .A0(n65), .A1(ofifoAddr2N[14]), .Z(n101));
Q_AN02 U5175 ( .A0(n65), .A1(ofifoAddr2N[15]), .Z(n100));
Q_AN02 U5176 ( .A0(n65), .A1(ofifoAddr2N[16]), .Z(n99));
Q_NR02 U5177 ( .A0(xc_top.GFReset), .A1(ofifoAddr7N[1]), .Z(n98));
Q_NR02 U5178 ( .A0(xc_top.GFReset), .A1(ofifoAddr5N[2]), .Z(n97));
Q_AN02 U5179 ( .A0(n65), .A1(ofifoAddr1N[3]), .Z(n96));
Q_AN02 U5180 ( .A0(n65), .A1(ofifoAddr1N[4]), .Z(n95));
Q_AN02 U5181 ( .A0(n65), .A1(ofifoAddr1N[5]), .Z(n94));
Q_AN02 U5182 ( .A0(n65), .A1(ofifoAddr1N[6]), .Z(n93));
Q_AN02 U5183 ( .A0(n65), .A1(ofifoAddr1N[7]), .Z(n92));
Q_AN02 U5184 ( .A0(n65), .A1(ofifoAddr1N[8]), .Z(n91));
Q_AN02 U5185 ( .A0(n65), .A1(ofifoAddr1N[9]), .Z(n90));
Q_AN02 U5186 ( .A0(n65), .A1(ofifoAddr1N[10]), .Z(n89));
Q_AN02 U5187 ( .A0(n65), .A1(ofifoAddr1N[11]), .Z(n88));
Q_AN02 U5188 ( .A0(n65), .A1(ofifoAddr1N[12]), .Z(n87));
Q_AN02 U5189 ( .A0(n65), .A1(ofifoAddr1N[13]), .Z(n86));
Q_AN02 U5190 ( .A0(n65), .A1(ofifoAddr1N[14]), .Z(n85));
Q_AN02 U5191 ( .A0(n65), .A1(ofifoAddr1N[15]), .Z(n84));
Q_AN02 U5192 ( .A0(n65), .A1(ofifoAddr1N[16]), .Z(n83));
Q_AN02 U5193 ( .A0(n65), .A1(ofifoAddr0N[0]), .Z(n82));
Q_AN02 U5194 ( .A0(n65), .A1(ofifoAddr0N[1]), .Z(n81));
Q_AN02 U5195 ( .A0(n65), .A1(ofifoAddr0N[2]), .Z(n80));
Q_AN02 U5196 ( .A0(n65), .A1(ofifoAddr0N[3]), .Z(n79));
Q_AN02 U5197 ( .A0(n65), .A1(ofifoAddr0N[4]), .Z(n78));
Q_AN02 U5198 ( .A0(n65), .A1(ofifoAddr0N[5]), .Z(n77));
Q_AN02 U5199 ( .A0(n65), .A1(ofifoAddr0N[6]), .Z(n76));
Q_AN02 U5200 ( .A0(n65), .A1(ofifoAddr0N[7]), .Z(n75));
Q_AN02 U5201 ( .A0(n65), .A1(ofifoAddr0N[8]), .Z(n74));
Q_AN02 U5202 ( .A0(n65), .A1(ofifoAddr0N[9]), .Z(n73));
Q_AN02 U5203 ( .A0(n65), .A1(ofifoAddr0N[10]), .Z(n72));
Q_AN02 U5204 ( .A0(n65), .A1(ofifoAddr0N[11]), .Z(n71));
Q_AN02 U5205 ( .A0(n65), .A1(ofifoAddr0N[12]), .Z(n70));
Q_AN02 U5206 ( .A0(n65), .A1(ofifoAddr0N[13]), .Z(n69));
Q_AN02 U5207 ( .A0(n65), .A1(ofifoAddr0N[14]), .Z(n68));
Q_AN02 U5208 ( .A0(n65), .A1(ofifoAddr0N[15]), .Z(n67));
Q_AN02 U5209 ( .A0(n65), .A1(ofifoAddr0N[16]), .Z(n66));
Q_FDP0UA U5210 ( .D(n66), .QTFCLK( ), .Q(ofifoAddr0[16]));
Q_FDP0UA U5211 ( .D(n67), .QTFCLK( ), .Q(ofifoAddr0[15]));
Q_FDP0UA U5212 ( .D(n68), .QTFCLK( ), .Q(ofifoAddr0[14]));
Q_FDP0UA U5213 ( .D(n69), .QTFCLK( ), .Q(ofifoAddr0[13]));
Q_FDP0UA U5214 ( .D(n70), .QTFCLK( ), .Q(ofifoAddr0[12]));
Q_FDP0UA U5215 ( .D(n71), .QTFCLK( ), .Q(ofifoAddr0[11]));
Q_FDP0UA U5216 ( .D(n72), .QTFCLK( ), .Q(ofifoAddr0[10]));
Q_FDP0UA U5217 ( .D(n73), .QTFCLK( ), .Q(ofifoAddr0[9]));
Q_FDP0UA U5218 ( .D(n74), .QTFCLK( ), .Q(ofifoAddr0[8]));
Q_FDP0UA U5219 ( .D(n75), .QTFCLK( ), .Q(ofifoAddr0[7]));
Q_FDP0UA U5220 ( .D(n76), .QTFCLK( ), .Q(ofifoAddr0[6]));
Q_FDP0UA U5221 ( .D(n77), .QTFCLK( ), .Q(ofifoAddr0[5]));
Q_FDP0UA U5222 ( .D(n78), .QTFCLK( ), .Q(ofifoAddr0[4]));
Q_FDP0UA U5223 ( .D(n79), .QTFCLK( ), .Q(ofifoAddr0[3]));
Q_FDP0UA U5224 ( .D(n80), .QTFCLK( ), .Q(ofifoAddr0[2]));
Q_FDP0UA U5225 ( .D(n81), .QTFCLK( ), .Q(ofifoAddr0[1]));
Q_FDP0UA U5226 ( .D(n82), .QTFCLK( ), .Q(ofifoAddr0[0]));
Q_FDP0UA U5227 ( .D(n83), .QTFCLK( ), .Q(ofifoAddr1[16]));
Q_FDP0UA U5228 ( .D(n84), .QTFCLK( ), .Q(ofifoAddr1[15]));
Q_FDP0UA U5229 ( .D(n85), .QTFCLK( ), .Q(ofifoAddr1[14]));
Q_FDP0UA U5230 ( .D(n86), .QTFCLK( ), .Q(ofifoAddr1[13]));
Q_FDP0UA U5231 ( .D(n87), .QTFCLK( ), .Q(ofifoAddr1[12]));
Q_FDP0UA U5232 ( .D(n88), .QTFCLK( ), .Q(ofifoAddr1[11]));
Q_FDP0UA U5233 ( .D(n89), .QTFCLK( ), .Q(ofifoAddr1[10]));
Q_FDP0UA U5234 ( .D(n90), .QTFCLK( ), .Q(ofifoAddr1[9]));
Q_FDP0UA U5235 ( .D(n91), .QTFCLK( ), .Q(ofifoAddr1[8]));
Q_FDP0UA U5236 ( .D(n92), .QTFCLK( ), .Q(ofifoAddr1[7]));
Q_FDP0UA U5237 ( .D(n93), .QTFCLK( ), .Q(ofifoAddr1[6]));
Q_FDP0UA U5238 ( .D(n94), .QTFCLK( ), .Q(ofifoAddr1[5]));
Q_FDP0UA U5239 ( .D(n95), .QTFCLK( ), .Q(ofifoAddr1[4]));
Q_FDP0UA U5240 ( .D(n96), .QTFCLK( ), .Q(ofifoAddr1[3]));
Q_FDP0UA U5241 ( .D(n97), .QTFCLK( ), .Q(ofifoAddr1[2]));
Q_FDP0UA U5242 ( .D(n98), .QTFCLK( ), .Q(ofifoAddr1[1]));
Q_FDP0UA U5243 ( .D(n3341), .QTFCLK( ), .Q(ofifoAddr1[0]));
Q_FDP0UA U5244 ( .D(n99), .QTFCLK( ), .Q(ofifoAddr2[16]));
Q_FDP0UA U5245 ( .D(n100), .QTFCLK( ), .Q(ofifoAddr2[15]));
Q_FDP0UA U5246 ( .D(n101), .QTFCLK( ), .Q(ofifoAddr2[14]));
Q_FDP0UA U5247 ( .D(n102), .QTFCLK( ), .Q(ofifoAddr2[13]));
Q_FDP0UA U5248 ( .D(n103), .QTFCLK( ), .Q(ofifoAddr2[12]));
Q_FDP0UA U5249 ( .D(n104), .QTFCLK( ), .Q(ofifoAddr2[11]));
Q_FDP0UA U5250 ( .D(n105), .QTFCLK( ), .Q(ofifoAddr2[10]));
Q_FDP0UA U5251 ( .D(n106), .QTFCLK( ), .Q(ofifoAddr2[9]));
Q_FDP0UA U5252 ( .D(n107), .QTFCLK( ), .Q(ofifoAddr2[8]));
Q_FDP0UA U5253 ( .D(n108), .QTFCLK( ), .Q(ofifoAddr2[7]));
Q_FDP0UA U5254 ( .D(n109), .QTFCLK( ), .Q(ofifoAddr2[6]));
Q_FDP0UA U5255 ( .D(n110), .QTFCLK( ), .Q(ofifoAddr2[5]));
Q_FDP0UA U5256 ( .D(n111), .QTFCLK( ), .Q(ofifoAddr2[4]));
Q_FDP0UA U5257 ( .D(n112), .QTFCLK( ), .Q(ofifoAddr2[3]));
Q_FDP0UA U5258 ( .D(n113), .QTFCLK( ), .Q(ofifoAddr2[2]));
Q_FDP0UA U5259 ( .D(n3342), .QTFCLK( ), .Q(ofifoAddr2[1]));
Q_FDP0UA U5260 ( .D(n82), .QTFCLK( ), .Q(ofifoAddr2[0]));
Q_FDP0UA U5261 ( .D(n99), .QTFCLK( ), .Q(ofifoAddr3[16]));
Q_FDP0UA U5262 ( .D(n100), .QTFCLK( ), .Q(ofifoAddr3[15]));
Q_FDP0UA U5263 ( .D(n101), .QTFCLK( ), .Q(ofifoAddr3[14]));
Q_FDP0UA U5264 ( .D(n102), .QTFCLK( ), .Q(ofifoAddr3[13]));
Q_FDP0UA U5265 ( .D(n103), .QTFCLK( ), .Q(ofifoAddr3[12]));
Q_FDP0UA U5266 ( .D(n104), .QTFCLK( ), .Q(ofifoAddr3[11]));
Q_FDP0UA U5267 ( .D(n105), .QTFCLK( ), .Q(ofifoAddr3[10]));
Q_FDP0UA U5268 ( .D(n106), .QTFCLK( ), .Q(ofifoAddr3[9]));
Q_FDP0UA U5269 ( .D(n107), .QTFCLK( ), .Q(ofifoAddr3[8]));
Q_FDP0UA U5270 ( .D(n108), .QTFCLK( ), .Q(ofifoAddr3[7]));
Q_FDP0UA U5271 ( .D(n109), .QTFCLK( ), .Q(ofifoAddr3[6]));
Q_FDP0UA U5272 ( .D(n110), .QTFCLK( ), .Q(ofifoAddr3[5]));
Q_FDP0UA U5273 ( .D(n111), .QTFCLK( ), .Q(ofifoAddr3[4]));
Q_FDP0UA U5274 ( .D(n112), .QTFCLK( ), .Q(ofifoAddr3[3]));
Q_FDP0UA U5275 ( .D(n113), .QTFCLK( ), .Q(ofifoAddr3[2]));
Q_FDP0UA U5276 ( .D(n3342), .QTFCLK( ), .Q(ofifoAddr3[1]));
Q_FDP0UA U5277 ( .D(n114), .QTFCLK( ), .Q(ofifoAddr3[0]));
Q_FDP0UA U5278 ( .D(n115), .QTFCLK( ), .Q(ofifoAddr4[16]));
Q_FDP0UA U5279 ( .D(n116), .QTFCLK( ), .Q(ofifoAddr4[15]));
Q_FDP0UA U5280 ( .D(n117), .QTFCLK( ), .Q(ofifoAddr4[14]));
Q_FDP0UA U5281 ( .D(n118), .QTFCLK( ), .Q(ofifoAddr4[13]));
Q_FDP0UA U5282 ( .D(n119), .QTFCLK( ), .Q(ofifoAddr4[12]));
Q_FDP0UA U5283 ( .D(n120), .QTFCLK( ), .Q(ofifoAddr4[11]));
Q_FDP0UA U5284 ( .D(n121), .QTFCLK( ), .Q(ofifoAddr4[10]));
Q_FDP0UA U5285 ( .D(n122), .QTFCLK( ), .Q(ofifoAddr4[9]));
Q_FDP0UA U5286 ( .D(n123), .QTFCLK( ), .Q(ofifoAddr4[8]));
Q_FDP0UA U5287 ( .D(n124), .QTFCLK( ), .Q(ofifoAddr4[7]));
Q_FDP0UA U5288 ( .D(n125), .QTFCLK( ), .Q(ofifoAddr4[6]));
Q_FDP0UA U5289 ( .D(n126), .QTFCLK( ), .Q(ofifoAddr4[5]));
Q_FDP0UA U5290 ( .D(n127), .QTFCLK( ), .Q(ofifoAddr4[4]));
Q_FDP0UA U5291 ( .D(n128), .QTFCLK( ), .Q(ofifoAddr4[3]));
Q_FDP0UA U5292 ( .D(n3343), .QTFCLK( ), .Q(ofifoAddr4[2]));
Q_FDP0UA U5293 ( .D(n81), .QTFCLK( ), .Q(ofifoAddr4[1]));
Q_FDP0UA U5294 ( .D(n82), .QTFCLK( ), .Q(ofifoAddr4[0]));
Q_FDP0UA U5295 ( .D(n129), .QTFCLK( ), .Q(ofifoAddr5[16]));
Q_FDP0UA U5296 ( .D(n130), .QTFCLK( ), .Q(ofifoAddr5[15]));
Q_FDP0UA U5297 ( .D(n131), .QTFCLK( ), .Q(ofifoAddr5[14]));
Q_FDP0UA U5298 ( .D(n132), .QTFCLK( ), .Q(ofifoAddr5[13]));
Q_FDP0UA U5299 ( .D(n133), .QTFCLK( ), .Q(ofifoAddr5[12]));
Q_FDP0UA U5300 ( .D(n134), .QTFCLK( ), .Q(ofifoAddr5[11]));
Q_FDP0UA U5301 ( .D(n135), .QTFCLK( ), .Q(ofifoAddr5[10]));
Q_FDP0UA U5302 ( .D(n136), .QTFCLK( ), .Q(ofifoAddr5[9]));
Q_FDP0UA U5303 ( .D(n137), .QTFCLK( ), .Q(ofifoAddr5[8]));
Q_FDP0UA U5304 ( .D(n138), .QTFCLK( ), .Q(ofifoAddr5[7]));
Q_FDP0UA U5305 ( .D(n139), .QTFCLK( ), .Q(ofifoAddr5[6]));
Q_FDP0UA U5306 ( .D(n140), .QTFCLK( ), .Q(ofifoAddr5[5]));
Q_FDP0UA U5307 ( .D(n141), .QTFCLK( ), .Q(ofifoAddr5[4]));
Q_FDP0UA U5308 ( .D(n142), .QTFCLK( ), .Q(ofifoAddr5[3]));
Q_FDP0UA U5309 ( .D(n3347), .QTFCLK( ), .Q(ofifoAddr5[2]));
Q_FDP0UA U5310 ( .D(n98), .QTFCLK( ), .Q(ofifoAddr5[1]));
Q_FDP0UA U5311 ( .D(n3341), .QTFCLK( ), .Q(ofifoAddr5[0]));
Q_FDP0UA U5312 ( .D(n143), .QTFCLK( ), .Q(ofifoAddr6[16]));
Q_FDP0UA U5313 ( .D(n144), .QTFCLK( ), .Q(ofifoAddr6[15]));
Q_FDP0UA U5314 ( .D(n145), .QTFCLK( ), .Q(ofifoAddr6[14]));
Q_FDP0UA U5315 ( .D(n146), .QTFCLK( ), .Q(ofifoAddr6[13]));
Q_FDP0UA U5316 ( .D(n147), .QTFCLK( ), .Q(ofifoAddr6[12]));
Q_FDP0UA U5317 ( .D(n148), .QTFCLK( ), .Q(ofifoAddr6[11]));
Q_FDP0UA U5318 ( .D(n149), .QTFCLK( ), .Q(ofifoAddr6[10]));
Q_FDP0UA U5319 ( .D(n150), .QTFCLK( ), .Q(ofifoAddr6[9]));
Q_FDP0UA U5320 ( .D(n151), .QTFCLK( ), .Q(ofifoAddr6[8]));
Q_FDP0UA U5321 ( .D(n152), .QTFCLK( ), .Q(ofifoAddr6[7]));
Q_FDP0UA U5322 ( .D(n153), .QTFCLK( ), .Q(ofifoAddr6[6]));
Q_FDP0UA U5323 ( .D(n154), .QTFCLK( ), .Q(ofifoAddr6[5]));
Q_FDP0UA U5324 ( .D(n155), .QTFCLK( ), .Q(ofifoAddr6[4]));
Q_FDP0UA U5325 ( .D(n156), .QTFCLK( ), .Q(ofifoAddr6[3]));
Q_FDP0UA U5326 ( .D(n3346), .QTFCLK( ), .Q(ofifoAddr6[2]));
Q_FDP0UA U5327 ( .D(n3342), .QTFCLK( ), .Q(ofifoAddr6[1]));
Q_FDP0UA U5328 ( .D(n82), .QTFCLK( ), .Q(ofifoAddr6[0]));
Q_FDP0UA U5329 ( .D(n157), .QTFCLK( ), .Q(ofifoAddr7[16]));
Q_FDP0UA U5330 ( .D(n158), .QTFCLK( ), .Q(ofifoAddr7[15]));
Q_FDP0UA U5331 ( .D(n159), .QTFCLK( ), .Q(ofifoAddr7[14]));
Q_FDP0UA U5332 ( .D(n160), .QTFCLK( ), .Q(ofifoAddr7[13]));
Q_FDP0UA U5333 ( .D(n161), .QTFCLK( ), .Q(ofifoAddr7[12]));
Q_FDP0UA U5334 ( .D(n162), .QTFCLK( ), .Q(ofifoAddr7[11]));
Q_FDP0UA U5335 ( .D(n163), .QTFCLK( ), .Q(ofifoAddr7[10]));
Q_FDP0UA U5336 ( .D(n164), .QTFCLK( ), .Q(ofifoAddr7[9]));
Q_FDP0UA U5337 ( .D(n165), .QTFCLK( ), .Q(ofifoAddr7[8]));
Q_FDP0UA U5338 ( .D(n166), .QTFCLK( ), .Q(ofifoAddr7[7]));
Q_FDP0UA U5339 ( .D(n167), .QTFCLK( ), .Q(ofifoAddr7[6]));
Q_FDP0UA U5340 ( .D(n168), .QTFCLK( ), .Q(ofifoAddr7[5]));
Q_FDP0UA U5341 ( .D(n169), .QTFCLK( ), .Q(ofifoAddr7[4]));
Q_FDP0UA U5342 ( .D(n170), .QTFCLK( ), .Q(ofifoAddr7[3]));
Q_FDP0UA U5343 ( .D(n171), .QTFCLK( ), .Q(ofifoAddr7[2]));
Q_FDP0UA U5344 ( .D(n3345), .QTFCLK( ), .Q(ofifoAddr7[1]));
Q_FDP0UA U5345 ( .D(n3341), .QTFCLK( ), .Q(ofifoAddr7[0]));
Q_FDP0UA U5346 ( .D(n172), .QTFCLK( ), .Q(ofifoAddr8[16]));
Q_FDP0UA U5347 ( .D(n173), .QTFCLK( ), .Q(ofifoAddr8[15]));
Q_FDP0UA U5348 ( .D(n174), .QTFCLK( ), .Q(ofifoAddr8[14]));
Q_FDP0UA U5349 ( .D(n175), .QTFCLK( ), .Q(ofifoAddr8[13]));
Q_FDP0UA U5350 ( .D(n176), .QTFCLK( ), .Q(ofifoAddr8[12]));
Q_FDP0UA U5351 ( .D(n177), .QTFCLK( ), .Q(ofifoAddr8[11]));
Q_FDP0UA U5352 ( .D(n178), .QTFCLK( ), .Q(ofifoAddr8[10]));
Q_FDP0UA U5353 ( .D(n179), .QTFCLK( ), .Q(ofifoAddr8[9]));
Q_FDP0UA U5354 ( .D(n180), .QTFCLK( ), .Q(ofifoAddr8[8]));
Q_FDP0UA U5355 ( .D(n181), .QTFCLK( ), .Q(ofifoAddr8[7]));
Q_FDP0UA U5356 ( .D(n182), .QTFCLK( ), .Q(ofifoAddr8[6]));
Q_FDP0UA U5357 ( .D(n183), .QTFCLK( ), .Q(ofifoAddr8[5]));
Q_FDP0UA U5358 ( .D(n184), .QTFCLK( ), .Q(ofifoAddr8[4]));
Q_FDP0UA U5359 ( .D(n3344), .QTFCLK( ), .Q(ofifoAddr8[3]));
Q_FDP0UA U5360 ( .D(n80), .QTFCLK( ), .Q(ofifoAddr8[2]));
Q_FDP0UA U5361 ( .D(n81), .QTFCLK( ), .Q(ofifoAddr8[1]));
Q_FDP0UA U5362 ( .D(n82), .QTFCLK( ), .Q(ofifoAddr8[0]));
Q_FDP0UA U5363 ( .D(n185), .QTFCLK( ), .Q(oFill[4]));
Q_FDP0UA U5364 ( .D(n186), .QTFCLK( ), .Q(oFill[3]));
Q_FDP0UA U5365 ( .D(n187), .QTFCLK( ), .Q(oFill[2]));
Q_FDP0UA U5366 ( .D(n188), .QTFCLK( ), .Q(oFill[1]));
Q_FDP0UA U5367 ( .D(n189), .QTFCLK( ), .Q(oFill[0]));
Q_FDP0UA U5368 ( .D(n190), .QTFCLK( ), .Q(ofifoWptr[16]));
Q_FDP0UA U5369 ( .D(n191), .QTFCLK( ), .Q(ofifoWptr[15]));
Q_FDP0UA U5370 ( .D(n192), .QTFCLK( ), .Q(ofifoWptr[14]));
Q_FDP0UA U5371 ( .D(n193), .QTFCLK( ), .Q(ofifoWptr[13]));
Q_FDP0UA U5372 ( .D(n194), .QTFCLK( ), .Q(ofifoWptr[12]));
Q_FDP0UA U5373 ( .D(n195), .QTFCLK( ), .Q(ofifoWptr[11]));
Q_FDP0UA U5374 ( .D(n196), .QTFCLK( ), .Q(ofifoWptr[10]));
Q_FDP0UA U5375 ( .D(n197), .QTFCLK( ), .Q(ofifoWptr[9]));
Q_FDP0UA U5376 ( .D(n198), .QTFCLK( ), .Q(ofifoWptr[8]));
Q_FDP0UA U5377 ( .D(n199), .QTFCLK( ), .Q(ofifoWptr[7]));
Q_FDP0UA U5378 ( .D(n200), .QTFCLK( ), .Q(ofifoWptr[6]));
Q_FDP0UA U5379 ( .D(n201), .QTFCLK( ), .Q(ofifoWptr[5]));
Q_FDP0UA U5380 ( .D(n202), .QTFCLK( ), .Q(ofifoWptr[4]));
Q_FDP0UA U5381 ( .D(n203), .QTFCLK( ), .Q(ofifoWptr[3]));
Q_FDP0UA U5382 ( .D(n204), .QTFCLK( ), .Q(ofifoWptr[2]));
Q_FDP0UA U5383 ( .D(n205), .QTFCLK( ), .Q(ofifoWptr[1]));
Q_FDP0UA U5384 ( .D(n206), .QTFCLK( ), .Q(ofifoWptr[0]));
Q_INV U5385 ( .A(xc_top.GFReset), .Z(n65));
Q_FDP0UA U5386 ( .D(n782), .QTFCLK( ), .Q(ofifoData[0]));
Q_FDP0UA U5387 ( .D(n781), .QTFCLK( ), .Q(ofifoData[1]));
Q_FDP0UA U5388 ( .D(n780), .QTFCLK( ), .Q(ofifoData[2]));
Q_FDP0UA U5389 ( .D(n779), .QTFCLK( ), .Q(ofifoData[3]));
Q_FDP0UA U5390 ( .D(n778), .QTFCLK( ), .Q(ofifoData[4]));
Q_FDP0UA U5391 ( .D(n777), .QTFCLK( ), .Q(ofifoData[5]));
Q_FDP0UA U5392 ( .D(n776), .QTFCLK( ), .Q(ofifoData[6]));
Q_FDP0UA U5393 ( .D(n775), .QTFCLK( ), .Q(ofifoData[7]));
Q_FDP0UA U5394 ( .D(n774), .QTFCLK( ), .Q(ofifoData[8]));
Q_FDP0UA U5395 ( .D(n773), .QTFCLK( ), .Q(ofifoData[9]));
Q_FDP0UA U5396 ( .D(n772), .QTFCLK( ), .Q(ofifoData[10]));
Q_FDP0UA U5397 ( .D(n771), .QTFCLK( ), .Q(ofifoData[11]));
Q_FDP0UA U5398 ( .D(n770), .QTFCLK( ), .Q(ofifoData[12]));
Q_FDP0UA U5399 ( .D(n769), .QTFCLK( ), .Q(ofifoData[13]));
Q_FDP0UA U5400 ( .D(n768), .QTFCLK( ), .Q(ofifoData[14]));
Q_FDP0UA U5401 ( .D(n767), .QTFCLK( ), .Q(ofifoData[15]));
Q_FDP0UA U5402 ( .D(n766), .QTFCLK( ), .Q(ofifoData[16]));
Q_FDP0UA U5403 ( .D(n765), .QTFCLK( ), .Q(ofifoData[17]));
Q_FDP0UA U5404 ( .D(n764), .QTFCLK( ), .Q(ofifoData[18]));
Q_FDP0UA U5405 ( .D(n763), .QTFCLK( ), .Q(ofifoData[19]));
Q_FDP0UA U5406 ( .D(n762), .QTFCLK( ), .Q(ofifoData[20]));
Q_FDP0UA U5407 ( .D(n761), .QTFCLK( ), .Q(ofifoData[21]));
Q_FDP0UA U5408 ( .D(n760), .QTFCLK( ), .Q(ofifoData[22]));
Q_FDP0UA U5409 ( .D(n759), .QTFCLK( ), .Q(ofifoData[23]));
Q_FDP0UA U5410 ( .D(n758), .QTFCLK( ), .Q(ofifoData[24]));
Q_FDP0UA U5411 ( .D(n757), .QTFCLK( ), .Q(ofifoData[25]));
Q_FDP0UA U5412 ( .D(n756), .QTFCLK( ), .Q(ofifoData[26]));
Q_FDP0UA U5413 ( .D(n755), .QTFCLK( ), .Q(ofifoData[27]));
Q_FDP0UA U5414 ( .D(n754), .QTFCLK( ), .Q(ofifoData[28]));
Q_FDP0UA U5415 ( .D(n753), .QTFCLK( ), .Q(ofifoData[29]));
Q_FDP0UA U5416 ( .D(n752), .QTFCLK( ), .Q(ofifoData[30]));
Q_FDP0UA U5417 ( .D(n751), .QTFCLK( ), .Q(ofifoData[31]));
Q_FDP0UA U5418 ( .D(n750), .QTFCLK( ), .Q(ofifoData[32]));
Q_FDP0UA U5419 ( .D(n749), .QTFCLK( ), .Q(ofifoData[33]));
Q_FDP0UA U5420 ( .D(n748), .QTFCLK( ), .Q(ofifoData[34]));
Q_FDP0UA U5421 ( .D(n747), .QTFCLK( ), .Q(ofifoData[35]));
Q_FDP0UA U5422 ( .D(n746), .QTFCLK( ), .Q(ofifoData[36]));
Q_FDP0UA U5423 ( .D(n745), .QTFCLK( ), .Q(ofifoData[37]));
Q_FDP0UA U5424 ( .D(n744), .QTFCLK( ), .Q(ofifoData[38]));
Q_FDP0UA U5425 ( .D(n743), .QTFCLK( ), .Q(ofifoData[39]));
Q_FDP0UA U5426 ( .D(n742), .QTFCLK( ), .Q(ofifoData[40]));
Q_FDP0UA U5427 ( .D(n741), .QTFCLK( ), .Q(ofifoData[41]));
Q_FDP0UA U5428 ( .D(n740), .QTFCLK( ), .Q(ofifoData[42]));
Q_FDP0UA U5429 ( .D(n739), .QTFCLK( ), .Q(ofifoData[43]));
Q_FDP0UA U5430 ( .D(n738), .QTFCLK( ), .Q(ofifoData[44]));
Q_FDP0UA U5431 ( .D(n737), .QTFCLK( ), .Q(ofifoData[45]));
Q_FDP0UA U5432 ( .D(n736), .QTFCLK( ), .Q(ofifoData[46]));
Q_FDP0UA U5433 ( .D(n735), .QTFCLK( ), .Q(ofifoData[47]));
Q_FDP0UA U5434 ( .D(n734), .QTFCLK( ), .Q(ofifoData[48]));
Q_FDP0UA U5435 ( .D(n733), .QTFCLK( ), .Q(ofifoData[49]));
Q_FDP0UA U5436 ( .D(n732), .QTFCLK( ), .Q(ofifoData[50]));
Q_FDP0UA U5437 ( .D(n731), .QTFCLK( ), .Q(ofifoData[51]));
Q_FDP0UA U5438 ( .D(n730), .QTFCLK( ), .Q(ofifoData[52]));
Q_FDP0UA U5439 ( .D(n729), .QTFCLK( ), .Q(ofifoData[53]));
Q_FDP0UA U5440 ( .D(n728), .QTFCLK( ), .Q(ofifoData[54]));
Q_FDP0UA U5441 ( .D(n727), .QTFCLK( ), .Q(ofifoData[55]));
Q_FDP0UA U5442 ( .D(n726), .QTFCLK( ), .Q(ofifoData[56]));
Q_FDP0UA U5443 ( .D(n725), .QTFCLK( ), .Q(ofifoData[57]));
Q_FDP0UA U5444 ( .D(n724), .QTFCLK( ), .Q(ofifoData[58]));
Q_FDP0UA U5445 ( .D(n723), .QTFCLK( ), .Q(ofifoData[59]));
Q_FDP0UA U5446 ( .D(n722), .QTFCLK( ), .Q(ofifoData[60]));
Q_FDP0UA U5447 ( .D(n721), .QTFCLK( ), .Q(ofifoData[61]));
Q_FDP0UA U5448 ( .D(n720), .QTFCLK( ), .Q(ofifoData[62]));
Q_FDP0UA U5449 ( .D(n719), .QTFCLK( ), .Q(ofifoData[63]));
Q_FDP0UA U5450 ( .D(n718), .QTFCLK( ), .Q(ofifoData[64]));
Q_FDP0UA U5451 ( .D(n717), .QTFCLK( ), .Q(ofifoData[65]));
Q_FDP0UA U5452 ( .D(n716), .QTFCLK( ), .Q(ofifoData[66]));
Q_FDP0UA U5453 ( .D(n715), .QTFCLK( ), .Q(ofifoData[67]));
Q_FDP0UA U5454 ( .D(n714), .QTFCLK( ), .Q(ofifoData[68]));
Q_FDP0UA U5455 ( .D(n713), .QTFCLK( ), .Q(ofifoData[69]));
Q_FDP0UA U5456 ( .D(n712), .QTFCLK( ), .Q(ofifoData[70]));
Q_FDP0UA U5457 ( .D(n711), .QTFCLK( ), .Q(ofifoData[71]));
Q_FDP0UA U5458 ( .D(n710), .QTFCLK( ), .Q(ofifoData[72]));
Q_FDP0UA U5459 ( .D(n709), .QTFCLK( ), .Q(ofifoData[73]));
Q_FDP0UA U5460 ( .D(n708), .QTFCLK( ), .Q(ofifoData[74]));
Q_FDP0UA U5461 ( .D(n707), .QTFCLK( ), .Q(ofifoData[75]));
Q_FDP0UA U5462 ( .D(n706), .QTFCLK( ), .Q(ofifoData[76]));
Q_FDP0UA U5463 ( .D(n705), .QTFCLK( ), .Q(ofifoData[77]));
Q_FDP0UA U5464 ( .D(n704), .QTFCLK( ), .Q(ofifoData[78]));
Q_FDP0UA U5465 ( .D(n703), .QTFCLK( ), .Q(ofifoData[79]));
Q_FDP0UA U5466 ( .D(n702), .QTFCLK( ), .Q(ofifoData[80]));
Q_FDP0UA U5467 ( .D(n701), .QTFCLK( ), .Q(ofifoData[81]));
Q_FDP0UA U5468 ( .D(n700), .QTFCLK( ), .Q(ofifoData[82]));
Q_FDP0UA U5469 ( .D(n699), .QTFCLK( ), .Q(ofifoData[83]));
Q_FDP0UA U5470 ( .D(n698), .QTFCLK( ), .Q(ofifoData[84]));
Q_FDP0UA U5471 ( .D(n697), .QTFCLK( ), .Q(ofifoData[85]));
Q_FDP0UA U5472 ( .D(n696), .QTFCLK( ), .Q(ofifoData[86]));
Q_FDP0UA U5473 ( .D(n695), .QTFCLK( ), .Q(ofifoData[87]));
Q_FDP0UA U5474 ( .D(n694), .QTFCLK( ), .Q(ofifoData[88]));
Q_FDP0UA U5475 ( .D(n693), .QTFCLK( ), .Q(ofifoData[89]));
Q_FDP0UA U5476 ( .D(n692), .QTFCLK( ), .Q(ofifoData[90]));
Q_FDP0UA U5477 ( .D(n691), .QTFCLK( ), .Q(ofifoData[91]));
Q_FDP0UA U5478 ( .D(n690), .QTFCLK( ), .Q(ofifoData[92]));
Q_FDP0UA U5479 ( .D(n689), .QTFCLK( ), .Q(ofifoData[93]));
Q_FDP0UA U5480 ( .D(n688), .QTFCLK( ), .Q(ofifoData[94]));
Q_FDP0UA U5481 ( .D(n687), .QTFCLK( ), .Q(ofifoData[95]));
Q_FDP0UA U5482 ( .D(n686), .QTFCLK( ), .Q(ofifoData[96]));
Q_FDP0UA U5483 ( .D(n685), .QTFCLK( ), .Q(ofifoData[97]));
Q_FDP0UA U5484 ( .D(n684), .QTFCLK( ), .Q(ofifoData[98]));
Q_FDP0UA U5485 ( .D(n683), .QTFCLK( ), .Q(ofifoData[99]));
Q_FDP0UA U5486 ( .D(n682), .QTFCLK( ), .Q(ofifoData[100]));
Q_FDP0UA U5487 ( .D(n681), .QTFCLK( ), .Q(ofifoData[101]));
Q_FDP0UA U5488 ( .D(n680), .QTFCLK( ), .Q(ofifoData[102]));
Q_FDP0UA U5489 ( .D(n679), .QTFCLK( ), .Q(ofifoData[103]));
Q_FDP0UA U5490 ( .D(n678), .QTFCLK( ), .Q(ofifoData[104]));
Q_FDP0UA U5491 ( .D(n677), .QTFCLK( ), .Q(ofifoData[105]));
Q_FDP0UA U5492 ( .D(n676), .QTFCLK( ), .Q(ofifoData[106]));
Q_FDP0UA U5493 ( .D(n675), .QTFCLK( ), .Q(ofifoData[107]));
Q_FDP0UA U5494 ( .D(n674), .QTFCLK( ), .Q(ofifoData[108]));
Q_FDP0UA U5495 ( .D(n673), .QTFCLK( ), .Q(ofifoData[109]));
Q_FDP0UA U5496 ( .D(n672), .QTFCLK( ), .Q(ofifoData[110]));
Q_FDP0UA U5497 ( .D(n671), .QTFCLK( ), .Q(ofifoData[111]));
Q_FDP0UA U5498 ( .D(n670), .QTFCLK( ), .Q(ofifoData[112]));
Q_FDP0UA U5499 ( .D(n669), .QTFCLK( ), .Q(ofifoData[113]));
Q_FDP0UA U5500 ( .D(n668), .QTFCLK( ), .Q(ofifoData[114]));
Q_FDP0UA U5501 ( .D(n667), .QTFCLK( ), .Q(ofifoData[115]));
Q_FDP0UA U5502 ( .D(n666), .QTFCLK( ), .Q(ofifoData[116]));
Q_FDP0UA U5503 ( .D(n665), .QTFCLK( ), .Q(ofifoData[117]));
Q_FDP0UA U5504 ( .D(n664), .QTFCLK( ), .Q(ofifoData[118]));
Q_FDP0UA U5505 ( .D(n663), .QTFCLK( ), .Q(ofifoData[119]));
Q_FDP0UA U5506 ( .D(n662), .QTFCLK( ), .Q(ofifoData[120]));
Q_FDP0UA U5507 ( .D(n661), .QTFCLK( ), .Q(ofifoData[121]));
Q_FDP0UA U5508 ( .D(n660), .QTFCLK( ), .Q(ofifoData[122]));
Q_FDP0UA U5509 ( .D(n659), .QTFCLK( ), .Q(ofifoData[123]));
Q_FDP0UA U5510 ( .D(n658), .QTFCLK( ), .Q(ofifoData[124]));
Q_FDP0UA U5511 ( .D(n657), .QTFCLK( ), .Q(ofifoData[125]));
Q_FDP0UA U5512 ( .D(n656), .QTFCLK( ), .Q(ofifoData[126]));
Q_FDP0UA U5513 ( .D(n655), .QTFCLK( ), .Q(ofifoData[127]));
Q_FDP0UA U5514 ( .D(n654), .QTFCLK( ), .Q(ofifoData[128]));
Q_FDP0UA U5515 ( .D(n653), .QTFCLK( ), .Q(ofifoData[129]));
Q_FDP0UA U5516 ( .D(n652), .QTFCLK( ), .Q(ofifoData[130]));
Q_FDP0UA U5517 ( .D(n651), .QTFCLK( ), .Q(ofifoData[131]));
Q_FDP0UA U5518 ( .D(n650), .QTFCLK( ), .Q(ofifoData[132]));
Q_FDP0UA U5519 ( .D(n649), .QTFCLK( ), .Q(ofifoData[133]));
Q_FDP0UA U5520 ( .D(n648), .QTFCLK( ), .Q(ofifoData[134]));
Q_FDP0UA U5521 ( .D(n647), .QTFCLK( ), .Q(ofifoData[135]));
Q_FDP0UA U5522 ( .D(n646), .QTFCLK( ), .Q(ofifoData[136]));
Q_FDP0UA U5523 ( .D(n645), .QTFCLK( ), .Q(ofifoData[137]));
Q_FDP0UA U5524 ( .D(n644), .QTFCLK( ), .Q(ofifoData[138]));
Q_FDP0UA U5525 ( .D(n643), .QTFCLK( ), .Q(ofifoData[139]));
Q_FDP0UA U5526 ( .D(n642), .QTFCLK( ), .Q(ofifoData[140]));
Q_FDP0UA U5527 ( .D(n641), .QTFCLK( ), .Q(ofifoData[141]));
Q_FDP0UA U5528 ( .D(n640), .QTFCLK( ), .Q(ofifoData[142]));
Q_FDP0UA U5529 ( .D(n639), .QTFCLK( ), .Q(ofifoData[143]));
Q_FDP0UA U5530 ( .D(n638), .QTFCLK( ), .Q(ofifoData[144]));
Q_FDP0UA U5531 ( .D(n637), .QTFCLK( ), .Q(ofifoData[145]));
Q_FDP0UA U5532 ( .D(n636), .QTFCLK( ), .Q(ofifoData[146]));
Q_FDP0UA U5533 ( .D(n635), .QTFCLK( ), .Q(ofifoData[147]));
Q_FDP0UA U5534 ( .D(n634), .QTFCLK( ), .Q(ofifoData[148]));
Q_FDP0UA U5535 ( .D(n633), .QTFCLK( ), .Q(ofifoData[149]));
Q_FDP0UA U5536 ( .D(n632), .QTFCLK( ), .Q(ofifoData[150]));
Q_FDP0UA U5537 ( .D(n631), .QTFCLK( ), .Q(ofifoData[151]));
Q_FDP0UA U5538 ( .D(n630), .QTFCLK( ), .Q(ofifoData[152]));
Q_FDP0UA U5539 ( .D(n629), .QTFCLK( ), .Q(ofifoData[153]));
Q_FDP0UA U5540 ( .D(n628), .QTFCLK( ), .Q(ofifoData[154]));
Q_FDP0UA U5541 ( .D(n627), .QTFCLK( ), .Q(ofifoData[155]));
Q_FDP0UA U5542 ( .D(n626), .QTFCLK( ), .Q(ofifoData[156]));
Q_FDP0UA U5543 ( .D(n625), .QTFCLK( ), .Q(ofifoData[157]));
Q_FDP0UA U5544 ( .D(n624), .QTFCLK( ), .Q(ofifoData[158]));
Q_FDP0UA U5545 ( .D(n623), .QTFCLK( ), .Q(ofifoData[159]));
Q_FDP0UA U5546 ( .D(n622), .QTFCLK( ), .Q(ofifoData[160]));
Q_FDP0UA U5547 ( .D(n621), .QTFCLK( ), .Q(ofifoData[161]));
Q_FDP0UA U5548 ( .D(n620), .QTFCLK( ), .Q(ofifoData[162]));
Q_FDP0UA U5549 ( .D(n619), .QTFCLK( ), .Q(ofifoData[163]));
Q_FDP0UA U5550 ( .D(n618), .QTFCLK( ), .Q(ofifoData[164]));
Q_FDP0UA U5551 ( .D(n617), .QTFCLK( ), .Q(ofifoData[165]));
Q_FDP0UA U5552 ( .D(n616), .QTFCLK( ), .Q(ofifoData[166]));
Q_FDP0UA U5553 ( .D(n615), .QTFCLK( ), .Q(ofifoData[167]));
Q_FDP0UA U5554 ( .D(n614), .QTFCLK( ), .Q(ofifoData[168]));
Q_FDP0UA U5555 ( .D(n613), .QTFCLK( ), .Q(ofifoData[169]));
Q_FDP0UA U5556 ( .D(n612), .QTFCLK( ), .Q(ofifoData[170]));
Q_FDP0UA U5557 ( .D(n611), .QTFCLK( ), .Q(ofifoData[171]));
Q_FDP0UA U5558 ( .D(n610), .QTFCLK( ), .Q(ofifoData[172]));
Q_FDP0UA U5559 ( .D(n609), .QTFCLK( ), .Q(ofifoData[173]));
Q_FDP0UA U5560 ( .D(n608), .QTFCLK( ), .Q(ofifoData[174]));
Q_FDP0UA U5561 ( .D(n607), .QTFCLK( ), .Q(ofifoData[175]));
Q_FDP0UA U5562 ( .D(n606), .QTFCLK( ), .Q(ofifoData[176]));
Q_FDP0UA U5563 ( .D(n605), .QTFCLK( ), .Q(ofifoData[177]));
Q_FDP0UA U5564 ( .D(n604), .QTFCLK( ), .Q(ofifoData[178]));
Q_FDP0UA U5565 ( .D(n603), .QTFCLK( ), .Q(ofifoData[179]));
Q_FDP0UA U5566 ( .D(n602), .QTFCLK( ), .Q(ofifoData[180]));
Q_FDP0UA U5567 ( .D(n601), .QTFCLK( ), .Q(ofifoData[181]));
Q_FDP0UA U5568 ( .D(n600), .QTFCLK( ), .Q(ofifoData[182]));
Q_FDP0UA U5569 ( .D(n599), .QTFCLK( ), .Q(ofifoData[183]));
Q_FDP0UA U5570 ( .D(n598), .QTFCLK( ), .Q(ofifoData[184]));
Q_FDP0UA U5571 ( .D(n597), .QTFCLK( ), .Q(ofifoData[185]));
Q_FDP0UA U5572 ( .D(n596), .QTFCLK( ), .Q(ofifoData[186]));
Q_FDP0UA U5573 ( .D(n595), .QTFCLK( ), .Q(ofifoData[187]));
Q_FDP0UA U5574 ( .D(n594), .QTFCLK( ), .Q(ofifoData[188]));
Q_FDP0UA U5575 ( .D(n593), .QTFCLK( ), .Q(ofifoData[189]));
Q_FDP0UA U5576 ( .D(n592), .QTFCLK( ), .Q(ofifoData[190]));
Q_FDP0UA U5577 ( .D(n591), .QTFCLK( ), .Q(ofifoData[191]));
Q_FDP0UA U5578 ( .D(n590), .QTFCLK( ), .Q(ofifoData[192]));
Q_FDP0UA U5579 ( .D(n589), .QTFCLK( ), .Q(ofifoData[193]));
Q_FDP0UA U5580 ( .D(n588), .QTFCLK( ), .Q(ofifoData[194]));
Q_FDP0UA U5581 ( .D(n587), .QTFCLK( ), .Q(ofifoData[195]));
Q_FDP0UA U5582 ( .D(n586), .QTFCLK( ), .Q(ofifoData[196]));
Q_FDP0UA U5583 ( .D(n585), .QTFCLK( ), .Q(ofifoData[197]));
Q_FDP0UA U5584 ( .D(n584), .QTFCLK( ), .Q(ofifoData[198]));
Q_FDP0UA U5585 ( .D(n583), .QTFCLK( ), .Q(ofifoData[199]));
Q_FDP0UA U5586 ( .D(n582), .QTFCLK( ), .Q(ofifoData[200]));
Q_FDP0UA U5587 ( .D(n581), .QTFCLK( ), .Q(ofifoData[201]));
Q_FDP0UA U5588 ( .D(n580), .QTFCLK( ), .Q(ofifoData[202]));
Q_FDP0UA U5589 ( .D(n579), .QTFCLK( ), .Q(ofifoData[203]));
Q_FDP0UA U5590 ( .D(n578), .QTFCLK( ), .Q(ofifoData[204]));
Q_FDP0UA U5591 ( .D(n577), .QTFCLK( ), .Q(ofifoData[205]));
Q_FDP0UA U5592 ( .D(n576), .QTFCLK( ), .Q(ofifoData[206]));
Q_FDP0UA U5593 ( .D(n575), .QTFCLK( ), .Q(ofifoData[207]));
Q_FDP0UA U5594 ( .D(n574), .QTFCLK( ), .Q(ofifoData[208]));
Q_FDP0UA U5595 ( .D(n573), .QTFCLK( ), .Q(ofifoData[209]));
Q_FDP0UA U5596 ( .D(n572), .QTFCLK( ), .Q(ofifoData[210]));
Q_FDP0UA U5597 ( .D(n571), .QTFCLK( ), .Q(ofifoData[211]));
Q_FDP0UA U5598 ( .D(n570), .QTFCLK( ), .Q(ofifoData[212]));
Q_FDP0UA U5599 ( .D(n569), .QTFCLK( ), .Q(ofifoData[213]));
Q_FDP0UA U5600 ( .D(n568), .QTFCLK( ), .Q(ofifoData[214]));
Q_FDP0UA U5601 ( .D(n567), .QTFCLK( ), .Q(ofifoData[215]));
Q_FDP0UA U5602 ( .D(n566), .QTFCLK( ), .Q(ofifoData[216]));
Q_FDP0UA U5603 ( .D(n565), .QTFCLK( ), .Q(ofifoData[217]));
Q_FDP0UA U5604 ( .D(n564), .QTFCLK( ), .Q(ofifoData[218]));
Q_FDP0UA U5605 ( .D(n563), .QTFCLK( ), .Q(ofifoData[219]));
Q_FDP0UA U5606 ( .D(n562), .QTFCLK( ), .Q(ofifoData[220]));
Q_FDP0UA U5607 ( .D(n561), .QTFCLK( ), .Q(ofifoData[221]));
Q_FDP0UA U5608 ( .D(n560), .QTFCLK( ), .Q(ofifoData[222]));
Q_FDP0UA U5609 ( .D(n559), .QTFCLK( ), .Q(ofifoData[223]));
Q_FDP0UA U5610 ( .D(n558), .QTFCLK( ), .Q(ofifoData[224]));
Q_FDP0UA U5611 ( .D(n557), .QTFCLK( ), .Q(ofifoData[225]));
Q_FDP0UA U5612 ( .D(n556), .QTFCLK( ), .Q(ofifoData[226]));
Q_FDP0UA U5613 ( .D(n555), .QTFCLK( ), .Q(ofifoData[227]));
Q_FDP0UA U5614 ( .D(n554), .QTFCLK( ), .Q(ofifoData[228]));
Q_FDP0UA U5615 ( .D(n553), .QTFCLK( ), .Q(ofifoData[229]));
Q_FDP0UA U5616 ( .D(n552), .QTFCLK( ), .Q(ofifoData[230]));
Q_FDP0UA U5617 ( .D(n551), .QTFCLK( ), .Q(ofifoData[231]));
Q_FDP0UA U5618 ( .D(n550), .QTFCLK( ), .Q(ofifoData[232]));
Q_FDP0UA U5619 ( .D(n549), .QTFCLK( ), .Q(ofifoData[233]));
Q_FDP0UA U5620 ( .D(n548), .QTFCLK( ), .Q(ofifoData[234]));
Q_FDP0UA U5621 ( .D(n547), .QTFCLK( ), .Q(ofifoData[235]));
Q_FDP0UA U5622 ( .D(n546), .QTFCLK( ), .Q(ofifoData[236]));
Q_FDP0UA U5623 ( .D(n545), .QTFCLK( ), .Q(ofifoData[237]));
Q_FDP0UA U5624 ( .D(n544), .QTFCLK( ), .Q(ofifoData[238]));
Q_FDP0UA U5625 ( .D(n543), .QTFCLK( ), .Q(ofifoData[239]));
Q_FDP0UA U5626 ( .D(n542), .QTFCLK( ), .Q(ofifoData[240]));
Q_FDP0UA U5627 ( .D(n541), .QTFCLK( ), .Q(ofifoData[241]));
Q_FDP0UA U5628 ( .D(n540), .QTFCLK( ), .Q(ofifoData[242]));
Q_FDP0UA U5629 ( .D(n539), .QTFCLK( ), .Q(ofifoData[243]));
Q_FDP0UA U5630 ( .D(n538), .QTFCLK( ), .Q(ofifoData[244]));
Q_FDP0UA U5631 ( .D(n537), .QTFCLK( ), .Q(ofifoData[245]));
Q_FDP0UA U5632 ( .D(n536), .QTFCLK( ), .Q(ofifoData[246]));
Q_FDP0UA U5633 ( .D(n535), .QTFCLK( ), .Q(ofifoData[247]));
Q_FDP0UA U5634 ( .D(n534), .QTFCLK( ), .Q(ofifoData[248]));
Q_FDP0UA U5635 ( .D(n533), .QTFCLK( ), .Q(ofifoData[249]));
Q_FDP0UA U5636 ( .D(n532), .QTFCLK( ), .Q(ofifoData[250]));
Q_FDP0UA U5637 ( .D(n531), .QTFCLK( ), .Q(ofifoData[251]));
Q_FDP0UA U5638 ( .D(n530), .QTFCLK( ), .Q(ofifoData[252]));
Q_FDP0UA U5639 ( .D(n529), .QTFCLK( ), .Q(ofifoData[253]));
Q_FDP0UA U5640 ( .D(n528), .QTFCLK( ), .Q(ofifoData[254]));
Q_FDP0UA U5641 ( .D(n527), .QTFCLK( ), .Q(ofifoData[255]));
Q_FDP0UA U5642 ( .D(n526), .QTFCLK( ), .Q(ofifoData[256]));
Q_FDP0UA U5643 ( .D(n525), .QTFCLK( ), .Q(ofifoData[257]));
Q_FDP0UA U5644 ( .D(n524), .QTFCLK( ), .Q(ofifoData[258]));
Q_FDP0UA U5645 ( .D(n523), .QTFCLK( ), .Q(ofifoData[259]));
Q_FDP0UA U5646 ( .D(n522), .QTFCLK( ), .Q(ofifoData[260]));
Q_FDP0UA U5647 ( .D(n521), .QTFCLK( ), .Q(ofifoData[261]));
Q_FDP0UA U5648 ( .D(n520), .QTFCLK( ), .Q(ofifoData[262]));
Q_FDP0UA U5649 ( .D(n519), .QTFCLK( ), .Q(ofifoData[263]));
Q_FDP0UA U5650 ( .D(n518), .QTFCLK( ), .Q(ofifoData[264]));
Q_FDP0UA U5651 ( .D(n517), .QTFCLK( ), .Q(ofifoData[265]));
Q_FDP0UA U5652 ( .D(n516), .QTFCLK( ), .Q(ofifoData[266]));
Q_FDP0UA U5653 ( .D(n515), .QTFCLK( ), .Q(ofifoData[267]));
Q_FDP0UA U5654 ( .D(n514), .QTFCLK( ), .Q(ofifoData[268]));
Q_FDP0UA U5655 ( .D(n513), .QTFCLK( ), .Q(ofifoData[269]));
Q_FDP0UA U5656 ( .D(n512), .QTFCLK( ), .Q(ofifoData[270]));
Q_FDP0UA U5657 ( .D(n511), .QTFCLK( ), .Q(ofifoData[271]));
Q_FDP0UA U5658 ( .D(n510), .QTFCLK( ), .Q(ofifoData[272]));
Q_FDP0UA U5659 ( .D(n509), .QTFCLK( ), .Q(ofifoData[273]));
Q_FDP0UA U5660 ( .D(n508), .QTFCLK( ), .Q(ofifoData[274]));
Q_FDP0UA U5661 ( .D(n507), .QTFCLK( ), .Q(ofifoData[275]));
Q_FDP0UA U5662 ( .D(n506), .QTFCLK( ), .Q(ofifoData[276]));
Q_FDP0UA U5663 ( .D(n505), .QTFCLK( ), .Q(ofifoData[277]));
Q_FDP0UA U5664 ( .D(n504), .QTFCLK( ), .Q(ofifoData[278]));
Q_FDP0UA U5665 ( .D(n503), .QTFCLK( ), .Q(ofifoData[279]));
Q_FDP0UA U5666 ( .D(n502), .QTFCLK( ), .Q(ofifoData[280]));
Q_FDP0UA U5667 ( .D(n501), .QTFCLK( ), .Q(ofifoData[281]));
Q_FDP0UA U5668 ( .D(n500), .QTFCLK( ), .Q(ofifoData[282]));
Q_FDP0UA U5669 ( .D(n499), .QTFCLK( ), .Q(ofifoData[283]));
Q_FDP0UA U5670 ( .D(n498), .QTFCLK( ), .Q(ofifoData[284]));
Q_FDP0UA U5671 ( .D(n497), .QTFCLK( ), .Q(ofifoData[285]));
Q_FDP0UA U5672 ( .D(n496), .QTFCLK( ), .Q(ofifoData[286]));
Q_FDP0UA U5673 ( .D(n495), .QTFCLK( ), .Q(ofifoData[287]));
Q_FDP0UA U5674 ( .D(n494), .QTFCLK( ), .Q(ofifoData[288]));
Q_FDP0UA U5675 ( .D(n493), .QTFCLK( ), .Q(ofifoData[289]));
Q_FDP0UA U5676 ( .D(n492), .QTFCLK( ), .Q(ofifoData[290]));
Q_FDP0UA U5677 ( .D(n491), .QTFCLK( ), .Q(ofifoData[291]));
Q_FDP0UA U5678 ( .D(n490), .QTFCLK( ), .Q(ofifoData[292]));
Q_FDP0UA U5679 ( .D(n489), .QTFCLK( ), .Q(ofifoData[293]));
Q_FDP0UA U5680 ( .D(n488), .QTFCLK( ), .Q(ofifoData[294]));
Q_FDP0UA U5681 ( .D(n487), .QTFCLK( ), .Q(ofifoData[295]));
Q_FDP0UA U5682 ( .D(n486), .QTFCLK( ), .Q(ofifoData[296]));
Q_FDP0UA U5683 ( .D(n485), .QTFCLK( ), .Q(ofifoData[297]));
Q_FDP0UA U5684 ( .D(n484), .QTFCLK( ), .Q(ofifoData[298]));
Q_FDP0UA U5685 ( .D(n483), .QTFCLK( ), .Q(ofifoData[299]));
Q_FDP0UA U5686 ( .D(n482), .QTFCLK( ), .Q(ofifoData[300]));
Q_FDP0UA U5687 ( .D(n481), .QTFCLK( ), .Q(ofifoData[301]));
Q_FDP0UA U5688 ( .D(n480), .QTFCLK( ), .Q(ofifoData[302]));
Q_FDP0UA U5689 ( .D(n479), .QTFCLK( ), .Q(ofifoData[303]));
Q_FDP0UA U5690 ( .D(n478), .QTFCLK( ), .Q(ofifoData[304]));
Q_FDP0UA U5691 ( .D(n477), .QTFCLK( ), .Q(ofifoData[305]));
Q_FDP0UA U5692 ( .D(n476), .QTFCLK( ), .Q(ofifoData[306]));
Q_FDP0UA U5693 ( .D(n475), .QTFCLK( ), .Q(ofifoData[307]));
Q_FDP0UA U5694 ( .D(n474), .QTFCLK( ), .Q(ofifoData[308]));
Q_FDP0UA U5695 ( .D(n473), .QTFCLK( ), .Q(ofifoData[309]));
Q_FDP0UA U5696 ( .D(n472), .QTFCLK( ), .Q(ofifoData[310]));
Q_FDP0UA U5697 ( .D(n471), .QTFCLK( ), .Q(ofifoData[311]));
Q_FDP0UA U5698 ( .D(n470), .QTFCLK( ), .Q(ofifoData[312]));
Q_FDP0UA U5699 ( .D(n469), .QTFCLK( ), .Q(ofifoData[313]));
Q_FDP0UA U5700 ( .D(n468), .QTFCLK( ), .Q(ofifoData[314]));
Q_FDP0UA U5701 ( .D(n467), .QTFCLK( ), .Q(ofifoData[315]));
Q_FDP0UA U5702 ( .D(n466), .QTFCLK( ), .Q(ofifoData[316]));
Q_FDP0UA U5703 ( .D(n465), .QTFCLK( ), .Q(ofifoData[317]));
Q_FDP0UA U5704 ( .D(n464), .QTFCLK( ), .Q(ofifoData[318]));
Q_FDP0UA U5705 ( .D(n463), .QTFCLK( ), .Q(ofifoData[319]));
Q_FDP0UA U5706 ( .D(n462), .QTFCLK( ), .Q(ofifoData[320]));
Q_FDP0UA U5707 ( .D(n461), .QTFCLK( ), .Q(ofifoData[321]));
Q_FDP0UA U5708 ( .D(n460), .QTFCLK( ), .Q(ofifoData[322]));
Q_FDP0UA U5709 ( .D(n459), .QTFCLK( ), .Q(ofifoData[323]));
Q_FDP0UA U5710 ( .D(n458), .QTFCLK( ), .Q(ofifoData[324]));
Q_FDP0UA U5711 ( .D(n457), .QTFCLK( ), .Q(ofifoData[325]));
Q_FDP0UA U5712 ( .D(n456), .QTFCLK( ), .Q(ofifoData[326]));
Q_FDP0UA U5713 ( .D(n455), .QTFCLK( ), .Q(ofifoData[327]));
Q_FDP0UA U5714 ( .D(n454), .QTFCLK( ), .Q(ofifoData[328]));
Q_FDP0UA U5715 ( .D(n453), .QTFCLK( ), .Q(ofifoData[329]));
Q_FDP0UA U5716 ( .D(n452), .QTFCLK( ), .Q(ofifoData[330]));
Q_FDP0UA U5717 ( .D(n451), .QTFCLK( ), .Q(ofifoData[331]));
Q_FDP0UA U5718 ( .D(n450), .QTFCLK( ), .Q(ofifoData[332]));
Q_FDP0UA U5719 ( .D(n449), .QTFCLK( ), .Q(ofifoData[333]));
Q_FDP0UA U5720 ( .D(n448), .QTFCLK( ), .Q(ofifoData[334]));
Q_FDP0UA U5721 ( .D(n447), .QTFCLK( ), .Q(ofifoData[335]));
Q_FDP0UA U5722 ( .D(n446), .QTFCLK( ), .Q(ofifoData[336]));
Q_FDP0UA U5723 ( .D(n445), .QTFCLK( ), .Q(ofifoData[337]));
Q_FDP0UA U5724 ( .D(n444), .QTFCLK( ), .Q(ofifoData[338]));
Q_FDP0UA U5725 ( .D(n443), .QTFCLK( ), .Q(ofifoData[339]));
Q_FDP0UA U5726 ( .D(n442), .QTFCLK( ), .Q(ofifoData[340]));
Q_FDP0UA U5727 ( .D(n441), .QTFCLK( ), .Q(ofifoData[341]));
Q_FDP0UA U5728 ( .D(n440), .QTFCLK( ), .Q(ofifoData[342]));
Q_FDP0UA U5729 ( .D(n439), .QTFCLK( ), .Q(ofifoData[343]));
Q_FDP0UA U5730 ( .D(n438), .QTFCLK( ), .Q(ofifoData[344]));
Q_FDP0UA U5731 ( .D(n437), .QTFCLK( ), .Q(ofifoData[345]));
Q_FDP0UA U5732 ( .D(n436), .QTFCLK( ), .Q(ofifoData[346]));
Q_FDP0UA U5733 ( .D(n435), .QTFCLK( ), .Q(ofifoData[347]));
Q_FDP0UA U5734 ( .D(n434), .QTFCLK( ), .Q(ofifoData[348]));
Q_FDP0UA U5735 ( .D(n433), .QTFCLK( ), .Q(ofifoData[349]));
Q_FDP0UA U5736 ( .D(n432), .QTFCLK( ), .Q(ofifoData[350]));
Q_FDP0UA U5737 ( .D(n431), .QTFCLK( ), .Q(ofifoData[351]));
Q_FDP0UA U5738 ( .D(n430), .QTFCLK( ), .Q(ofifoData[352]));
Q_FDP0UA U5739 ( .D(n429), .QTFCLK( ), .Q(ofifoData[353]));
Q_FDP0UA U5740 ( .D(n428), .QTFCLK( ), .Q(ofifoData[354]));
Q_FDP0UA U5741 ( .D(n427), .QTFCLK( ), .Q(ofifoData[355]));
Q_FDP0UA U5742 ( .D(n426), .QTFCLK( ), .Q(ofifoData[356]));
Q_FDP0UA U5743 ( .D(n425), .QTFCLK( ), .Q(ofifoData[357]));
Q_FDP0UA U5744 ( .D(n424), .QTFCLK( ), .Q(ofifoData[358]));
Q_FDP0UA U5745 ( .D(n423), .QTFCLK( ), .Q(ofifoData[359]));
Q_FDP0UA U5746 ( .D(n422), .QTFCLK( ), .Q(ofifoData[360]));
Q_FDP0UA U5747 ( .D(n421), .QTFCLK( ), .Q(ofifoData[361]));
Q_FDP0UA U5748 ( .D(n420), .QTFCLK( ), .Q(ofifoData[362]));
Q_FDP0UA U5749 ( .D(n419), .QTFCLK( ), .Q(ofifoData[363]));
Q_FDP0UA U5750 ( .D(n418), .QTFCLK( ), .Q(ofifoData[364]));
Q_FDP0UA U5751 ( .D(n417), .QTFCLK( ), .Q(ofifoData[365]));
Q_FDP0UA U5752 ( .D(n416), .QTFCLK( ), .Q(ofifoData[366]));
Q_FDP0UA U5753 ( .D(n415), .QTFCLK( ), .Q(ofifoData[367]));
Q_FDP0UA U5754 ( .D(n414), .QTFCLK( ), .Q(ofifoData[368]));
Q_FDP0UA U5755 ( .D(n413), .QTFCLK( ), .Q(ofifoData[369]));
Q_FDP0UA U5756 ( .D(n412), .QTFCLK( ), .Q(ofifoData[370]));
Q_FDP0UA U5757 ( .D(n411), .QTFCLK( ), .Q(ofifoData[371]));
Q_FDP0UA U5758 ( .D(n410), .QTFCLK( ), .Q(ofifoData[372]));
Q_FDP0UA U5759 ( .D(n409), .QTFCLK( ), .Q(ofifoData[373]));
Q_FDP0UA U5760 ( .D(n408), .QTFCLK( ), .Q(ofifoData[374]));
Q_FDP0UA U5761 ( .D(n407), .QTFCLK( ), .Q(ofifoData[375]));
Q_FDP0UA U5762 ( .D(n406), .QTFCLK( ), .Q(ofifoData[376]));
Q_FDP0UA U5763 ( .D(n405), .QTFCLK( ), .Q(ofifoData[377]));
Q_FDP0UA U5764 ( .D(n404), .QTFCLK( ), .Q(ofifoData[378]));
Q_FDP0UA U5765 ( .D(n403), .QTFCLK( ), .Q(ofifoData[379]));
Q_FDP0UA U5766 ( .D(n402), .QTFCLK( ), .Q(ofifoData[380]));
Q_FDP0UA U5767 ( .D(n401), .QTFCLK( ), .Q(ofifoData[381]));
Q_FDP0UA U5768 ( .D(n400), .QTFCLK( ), .Q(ofifoData[382]));
Q_FDP0UA U5769 ( .D(n399), .QTFCLK( ), .Q(ofifoData[383]));
Q_FDP0UA U5770 ( .D(n398), .QTFCLK( ), .Q(ofifoData[384]));
Q_FDP0UA U5771 ( .D(n397), .QTFCLK( ), .Q(ofifoData[385]));
Q_FDP0UA U5772 ( .D(n396), .QTFCLK( ), .Q(ofifoData[386]));
Q_FDP0UA U5773 ( .D(n395), .QTFCLK( ), .Q(ofifoData[387]));
Q_FDP0UA U5774 ( .D(n394), .QTFCLK( ), .Q(ofifoData[388]));
Q_FDP0UA U5775 ( .D(n393), .QTFCLK( ), .Q(ofifoData[389]));
Q_FDP0UA U5776 ( .D(n392), .QTFCLK( ), .Q(ofifoData[390]));
Q_FDP0UA U5777 ( .D(n391), .QTFCLK( ), .Q(ofifoData[391]));
Q_FDP0UA U5778 ( .D(n390), .QTFCLK( ), .Q(ofifoData[392]));
Q_FDP0UA U5779 ( .D(n389), .QTFCLK( ), .Q(ofifoData[393]));
Q_FDP0UA U5780 ( .D(n388), .QTFCLK( ), .Q(ofifoData[394]));
Q_FDP0UA U5781 ( .D(n387), .QTFCLK( ), .Q(ofifoData[395]));
Q_FDP0UA U5782 ( .D(n386), .QTFCLK( ), .Q(ofifoData[396]));
Q_FDP0UA U5783 ( .D(n385), .QTFCLK( ), .Q(ofifoData[397]));
Q_FDP0UA U5784 ( .D(n384), .QTFCLK( ), .Q(ofifoData[398]));
Q_FDP0UA U5785 ( .D(n383), .QTFCLK( ), .Q(ofifoData[399]));
Q_FDP0UA U5786 ( .D(n382), .QTFCLK( ), .Q(ofifoData[400]));
Q_FDP0UA U5787 ( .D(n381), .QTFCLK( ), .Q(ofifoData[401]));
Q_FDP0UA U5788 ( .D(n380), .QTFCLK( ), .Q(ofifoData[402]));
Q_FDP0UA U5789 ( .D(n379), .QTFCLK( ), .Q(ofifoData[403]));
Q_FDP0UA U5790 ( .D(n378), .QTFCLK( ), .Q(ofifoData[404]));
Q_FDP0UA U5791 ( .D(n377), .QTFCLK( ), .Q(ofifoData[405]));
Q_FDP0UA U5792 ( .D(n376), .QTFCLK( ), .Q(ofifoData[406]));
Q_FDP0UA U5793 ( .D(n375), .QTFCLK( ), .Q(ofifoData[407]));
Q_FDP0UA U5794 ( .D(n374), .QTFCLK( ), .Q(ofifoData[408]));
Q_FDP0UA U5795 ( .D(n373), .QTFCLK( ), .Q(ofifoData[409]));
Q_FDP0UA U5796 ( .D(n372), .QTFCLK( ), .Q(ofifoData[410]));
Q_FDP0UA U5797 ( .D(n371), .QTFCLK( ), .Q(ofifoData[411]));
Q_FDP0UA U5798 ( .D(n370), .QTFCLK( ), .Q(ofifoData[412]));
Q_FDP0UA U5799 ( .D(n369), .QTFCLK( ), .Q(ofifoData[413]));
Q_FDP0UA U5800 ( .D(n368), .QTFCLK( ), .Q(ofifoData[414]));
Q_FDP0UA U5801 ( .D(n367), .QTFCLK( ), .Q(ofifoData[415]));
Q_FDP0UA U5802 ( .D(n366), .QTFCLK( ), .Q(ofifoData[416]));
Q_FDP0UA U5803 ( .D(n365), .QTFCLK( ), .Q(ofifoData[417]));
Q_FDP0UA U5804 ( .D(n364), .QTFCLK( ), .Q(ofifoData[418]));
Q_FDP0UA U5805 ( .D(n363), .QTFCLK( ), .Q(ofifoData[419]));
Q_FDP0UA U5806 ( .D(n362), .QTFCLK( ), .Q(ofifoData[420]));
Q_FDP0UA U5807 ( .D(n361), .QTFCLK( ), .Q(ofifoData[421]));
Q_FDP0UA U5808 ( .D(n360), .QTFCLK( ), .Q(ofifoData[422]));
Q_FDP0UA U5809 ( .D(n359), .QTFCLK( ), .Q(ofifoData[423]));
Q_FDP0UA U5810 ( .D(n358), .QTFCLK( ), .Q(ofifoData[424]));
Q_FDP0UA U5811 ( .D(n357), .QTFCLK( ), .Q(ofifoData[425]));
Q_FDP0UA U5812 ( .D(n356), .QTFCLK( ), .Q(ofifoData[426]));
Q_FDP0UA U5813 ( .D(n355), .QTFCLK( ), .Q(ofifoData[427]));
Q_FDP0UA U5814 ( .D(n354), .QTFCLK( ), .Q(ofifoData[428]));
Q_FDP0UA U5815 ( .D(n353), .QTFCLK( ), .Q(ofifoData[429]));
Q_FDP0UA U5816 ( .D(n352), .QTFCLK( ), .Q(ofifoData[430]));
Q_FDP0UA U5817 ( .D(n351), .QTFCLK( ), .Q(ofifoData[431]));
Q_FDP0UA U5818 ( .D(n350), .QTFCLK( ), .Q(ofifoData[432]));
Q_FDP0UA U5819 ( .D(n349), .QTFCLK( ), .Q(ofifoData[433]));
Q_FDP0UA U5820 ( .D(n348), .QTFCLK( ), .Q(ofifoData[434]));
Q_FDP0UA U5821 ( .D(n347), .QTFCLK( ), .Q(ofifoData[435]));
Q_FDP0UA U5822 ( .D(n346), .QTFCLK( ), .Q(ofifoData[436]));
Q_FDP0UA U5823 ( .D(n345), .QTFCLK( ), .Q(ofifoData[437]));
Q_FDP0UA U5824 ( .D(n344), .QTFCLK( ), .Q(ofifoData[438]));
Q_FDP0UA U5825 ( .D(n343), .QTFCLK( ), .Q(ofifoData[439]));
Q_FDP0UA U5826 ( .D(n342), .QTFCLK( ), .Q(ofifoData[440]));
Q_FDP0UA U5827 ( .D(n341), .QTFCLK( ), .Q(ofifoData[441]));
Q_FDP0UA U5828 ( .D(n340), .QTFCLK( ), .Q(ofifoData[442]));
Q_FDP0UA U5829 ( .D(n339), .QTFCLK( ), .Q(ofifoData[443]));
Q_FDP0UA U5830 ( .D(n338), .QTFCLK( ), .Q(ofifoData[444]));
Q_FDP0UA U5831 ( .D(n337), .QTFCLK( ), .Q(ofifoData[445]));
Q_FDP0UA U5832 ( .D(n336), .QTFCLK( ), .Q(ofifoData[446]));
Q_FDP0UA U5833 ( .D(n335), .QTFCLK( ), .Q(ofifoData[447]));
Q_FDP0UA U5834 ( .D(n334), .QTFCLK( ), .Q(ofifoData[448]));
Q_FDP0UA U5835 ( .D(n333), .QTFCLK( ), .Q(ofifoData[449]));
Q_FDP0UA U5836 ( .D(n332), .QTFCLK( ), .Q(ofifoData[450]));
Q_FDP0UA U5837 ( .D(n331), .QTFCLK( ), .Q(ofifoData[451]));
Q_FDP0UA U5838 ( .D(n330), .QTFCLK( ), .Q(ofifoData[452]));
Q_FDP0UA U5839 ( .D(n329), .QTFCLK( ), .Q(ofifoData[453]));
Q_FDP0UA U5840 ( .D(n328), .QTFCLK( ), .Q(ofifoData[454]));
Q_FDP0UA U5841 ( .D(n327), .QTFCLK( ), .Q(ofifoData[455]));
Q_FDP0UA U5842 ( .D(n326), .QTFCLK( ), .Q(ofifoData[456]));
Q_FDP0UA U5843 ( .D(n325), .QTFCLK( ), .Q(ofifoData[457]));
Q_FDP0UA U5844 ( .D(n324), .QTFCLK( ), .Q(ofifoData[458]));
Q_FDP0UA U5845 ( .D(n323), .QTFCLK( ), .Q(ofifoData[459]));
Q_FDP0UA U5846 ( .D(n322), .QTFCLK( ), .Q(ofifoData[460]));
Q_FDP0UA U5847 ( .D(n321), .QTFCLK( ), .Q(ofifoData[461]));
Q_FDP0UA U5848 ( .D(n320), .QTFCLK( ), .Q(ofifoData[462]));
Q_FDP0UA U5849 ( .D(n319), .QTFCLK( ), .Q(ofifoData[463]));
Q_FDP0UA U5850 ( .D(n318), .QTFCLK( ), .Q(ofifoData[464]));
Q_FDP0UA U5851 ( .D(n317), .QTFCLK( ), .Q(ofifoData[465]));
Q_FDP0UA U5852 ( .D(n316), .QTFCLK( ), .Q(ofifoData[466]));
Q_FDP0UA U5853 ( .D(n315), .QTFCLK( ), .Q(ofifoData[467]));
Q_FDP0UA U5854 ( .D(n314), .QTFCLK( ), .Q(ofifoData[468]));
Q_FDP0UA U5855 ( .D(n313), .QTFCLK( ), .Q(ofifoData[469]));
Q_FDP0UA U5856 ( .D(n312), .QTFCLK( ), .Q(ofifoData[470]));
Q_FDP0UA U5857 ( .D(n311), .QTFCLK( ), .Q(ofifoData[471]));
Q_FDP0UA U5858 ( .D(n310), .QTFCLK( ), .Q(ofifoData[472]));
Q_FDP0UA U5859 ( .D(n309), .QTFCLK( ), .Q(ofifoData[473]));
Q_FDP0UA U5860 ( .D(n308), .QTFCLK( ), .Q(ofifoData[474]));
Q_FDP0UA U5861 ( .D(n307), .QTFCLK( ), .Q(ofifoData[475]));
Q_FDP0UA U5862 ( .D(n306), .QTFCLK( ), .Q(ofifoData[476]));
Q_FDP0UA U5863 ( .D(n305), .QTFCLK( ), .Q(ofifoData[477]));
Q_FDP0UA U5864 ( .D(n304), .QTFCLK( ), .Q(ofifoData[478]));
Q_FDP0UA U5865 ( .D(n303), .QTFCLK( ), .Q(ofifoData[479]));
Q_FDP0UA U5866 ( .D(n302), .QTFCLK( ), .Q(ofifoData[480]));
Q_FDP0UA U5867 ( .D(n301), .QTFCLK( ), .Q(ofifoData[481]));
Q_FDP0UA U5868 ( .D(n300), .QTFCLK( ), .Q(ofifoData[482]));
Q_FDP0UA U5869 ( .D(n299), .QTFCLK( ), .Q(ofifoData[483]));
Q_FDP0UA U5870 ( .D(n298), .QTFCLK( ), .Q(ofifoData[484]));
Q_FDP0UA U5871 ( .D(n297), .QTFCLK( ), .Q(ofifoData[485]));
Q_FDP0UA U5872 ( .D(n296), .QTFCLK( ), .Q(ofifoData[486]));
Q_FDP0UA U5873 ( .D(n295), .QTFCLK( ), .Q(ofifoData[487]));
Q_FDP0UA U5874 ( .D(n294), .QTFCLK( ), .Q(ofifoData[488]));
Q_FDP0UA U5875 ( .D(n293), .QTFCLK( ), .Q(ofifoData[489]));
Q_FDP0UA U5876 ( .D(n292), .QTFCLK( ), .Q(ofifoData[490]));
Q_FDP0UA U5877 ( .D(n291), .QTFCLK( ), .Q(ofifoData[491]));
Q_FDP0UA U5878 ( .D(n290), .QTFCLK( ), .Q(ofifoData[492]));
Q_FDP0UA U5879 ( .D(n289), .QTFCLK( ), .Q(ofifoData[493]));
Q_FDP0UA U5880 ( .D(n288), .QTFCLK( ), .Q(ofifoData[494]));
Q_FDP0UA U5881 ( .D(n287), .QTFCLK( ), .Q(ofifoData[495]));
Q_FDP0UA U5882 ( .D(n286), .QTFCLK( ), .Q(ofifoData[496]));
Q_FDP0UA U5883 ( .D(n285), .QTFCLK( ), .Q(ofifoData[497]));
Q_FDP0UA U5884 ( .D(n284), .QTFCLK( ), .Q(ofifoData[498]));
Q_FDP0UA U5885 ( .D(n283), .QTFCLK( ), .Q(ofifoData[499]));
Q_FDP0UA U5886 ( .D(n282), .QTFCLK( ), .Q(ofifoData[500]));
Q_FDP0UA U5887 ( .D(n281), .QTFCLK( ), .Q(ofifoData[501]));
Q_FDP0UA U5888 ( .D(n280), .QTFCLK( ), .Q(ofifoData[502]));
Q_FDP0UA U5889 ( .D(n279), .QTFCLK( ), .Q(ofifoData[503]));
Q_FDP0UA U5890 ( .D(n278), .QTFCLK( ), .Q(ofifoData[504]));
Q_FDP0UA U5891 ( .D(n277), .QTFCLK( ), .Q(ofifoData[505]));
Q_FDP0UA U5892 ( .D(n276), .QTFCLK( ), .Q(ofifoData[506]));
Q_FDP0UA U5893 ( .D(n275), .QTFCLK( ), .Q(ofifoData[507]));
Q_FDP0UA U5894 ( .D(n274), .QTFCLK( ), .Q(ofifoData[508]));
Q_FDP0UA U5895 ( .D(n273), .QTFCLK( ), .Q(ofifoData[509]));
Q_FDP0UA U5896 ( .D(n272), .QTFCLK( ), .Q(ofifoData[510]));
Q_FDP0UA U5897 ( .D(n271), .QTFCLK( ), .Q(ofifoData[511]));
Q_FDP0UA U5898 ( .D(n270), .QTFCLK( ), .Q(ofifoData[512]));
Q_FDP0UA U5899 ( .D(n269), .QTFCLK( ), .Q(ofifoData[513]));
Q_FDP0UA U5900 ( .D(n268), .QTFCLK( ), .Q(ofifoData[514]));
Q_FDP0UA U5901 ( .D(n267), .QTFCLK( ), .Q(ofifoData[515]));
Q_FDP0UA U5902 ( .D(n266), .QTFCLK( ), .Q(ofifoData[516]));
Q_FDP0UA U5903 ( .D(n265), .QTFCLK( ), .Q(ofifoData[517]));
Q_FDP0UA U5904 ( .D(n264), .QTFCLK( ), .Q(ofifoData[518]));
Q_FDP0UA U5905 ( .D(n263), .QTFCLK( ), .Q(ofifoData[519]));
Q_FDP0UA U5906 ( .D(n262), .QTFCLK( ), .Q(ofifoData[520]));
Q_FDP0UA U5907 ( .D(n261), .QTFCLK( ), .Q(ofifoData[521]));
Q_FDP0UA U5908 ( .D(n260), .QTFCLK( ), .Q(ofifoData[522]));
Q_FDP0UA U5909 ( .D(n259), .QTFCLK( ), .Q(ofifoData[523]));
Q_FDP0UA U5910 ( .D(n258), .QTFCLK( ), .Q(ofifoData[524]));
Q_FDP0UA U5911 ( .D(n257), .QTFCLK( ), .Q(ofifoData[525]));
Q_FDP0UA U5912 ( .D(n256), .QTFCLK( ), .Q(ofifoData[526]));
Q_FDP0UA U5913 ( .D(n255), .QTFCLK( ), .Q(ofifoData[527]));
Q_FDP0UA U5914 ( .D(n254), .QTFCLK( ), .Q(ofifoData[528]));
Q_FDP0UA U5915 ( .D(n253), .QTFCLK( ), .Q(ofifoData[529]));
Q_FDP0UA U5916 ( .D(n252), .QTFCLK( ), .Q(ofifoData[530]));
Q_FDP0UA U5917 ( .D(n251), .QTFCLK( ), .Q(ofifoData[531]));
Q_FDP0UA U5918 ( .D(n250), .QTFCLK( ), .Q(ofifoData[532]));
Q_FDP0UA U5919 ( .D(n249), .QTFCLK( ), .Q(ofifoData[533]));
Q_FDP0UA U5920 ( .D(n248), .QTFCLK( ), .Q(ofifoData[534]));
Q_FDP0UA U5921 ( .D(n247), .QTFCLK( ), .Q(ofifoData[535]));
Q_FDP0UA U5922 ( .D(n246), .QTFCLK( ), .Q(ofifoData[536]));
Q_FDP0UA U5923 ( .D(n245), .QTFCLK( ), .Q(ofifoData[537]));
Q_FDP0UA U5924 ( .D(n244), .QTFCLK( ), .Q(ofifoData[538]));
Q_FDP0UA U5925 ( .D(n243), .QTFCLK( ), .Q(ofifoData[539]));
Q_FDP0UA U5926 ( .D(n242), .QTFCLK( ), .Q(ofifoData[540]));
Q_FDP0UA U5927 ( .D(n241), .QTFCLK( ), .Q(ofifoData[541]));
Q_FDP0UA U5928 ( .D(n240), .QTFCLK( ), .Q(ofifoData[542]));
Q_FDP0UA U5929 ( .D(n239), .QTFCLK( ), .Q(ofifoData[543]));
Q_FDP0UA U5930 ( .D(n238), .QTFCLK( ), .Q(ofifoData[544]));
Q_FDP0UA U5931 ( .D(n237), .QTFCLK( ), .Q(ofifoData[545]));
Q_FDP0UA U5932 ( .D(n236), .QTFCLK( ), .Q(ofifoData[546]));
Q_FDP0UA U5933 ( .D(n235), .QTFCLK( ), .Q(ofifoData[547]));
Q_FDP0UA U5934 ( .D(n234), .QTFCLK( ), .Q(ofifoData[548]));
Q_FDP0UA U5935 ( .D(n233), .QTFCLK( ), .Q(ofifoData[549]));
Q_FDP0UA U5936 ( .D(n232), .QTFCLK( ), .Q(ofifoData[550]));
Q_FDP0UA U5937 ( .D(n231), .QTFCLK( ), .Q(ofifoData[551]));
Q_FDP0UA U5938 ( .D(n230), .QTFCLK( ), .Q(ofifoData[552]));
Q_FDP0UA U5939 ( .D(n229), .QTFCLK( ), .Q(ofifoData[553]));
Q_FDP0UA U5940 ( .D(n228), .QTFCLK( ), .Q(ofifoData[554]));
Q_FDP0UA U5941 ( .D(n227), .QTFCLK( ), .Q(ofifoData[555]));
Q_FDP0UA U5942 ( .D(n226), .QTFCLK( ), .Q(ofifoData[556]));
Q_FDP0UA U5943 ( .D(n225), .QTFCLK( ), .Q(ofifoData[557]));
Q_FDP0UA U5944 ( .D(n224), .QTFCLK( ), .Q(ofifoData[558]));
Q_FDP0UA U5945 ( .D(n223), .QTFCLK( ), .Q(ofifoData[559]));
Q_FDP0UA U5946 ( .D(n222), .QTFCLK( ), .Q(ofifoData[560]));
Q_FDP0UA U5947 ( .D(n221), .QTFCLK( ), .Q(ofifoData[561]));
Q_FDP0UA U5948 ( .D(n220), .QTFCLK( ), .Q(ofifoData[562]));
Q_FDP0UA U5949 ( .D(n219), .QTFCLK( ), .Q(ofifoData[563]));
Q_FDP0UA U5950 ( .D(n218), .QTFCLK( ), .Q(ofifoData[564]));
Q_FDP0UA U5951 ( .D(n217), .QTFCLK( ), .Q(ofifoData[565]));
Q_FDP0UA U5952 ( .D(n216), .QTFCLK( ), .Q(ofifoData[566]));
Q_FDP0UA U5953 ( .D(n215), .QTFCLK( ), .Q(ofifoData[567]));
Q_FDP0UA U5954 ( .D(n214), .QTFCLK( ), .Q(ofifoData[568]));
Q_FDP0UA U5955 ( .D(n213), .QTFCLK( ), .Q(ofifoData[569]));
Q_FDP0UA U5956 ( .D(n212), .QTFCLK( ), .Q(ofifoData[570]));
Q_FDP0UA U5957 ( .D(n211), .QTFCLK( ), .Q(ofifoData[571]));
Q_FDP0UA U5958 ( .D(n210), .QTFCLK( ), .Q(ofifoData[572]));
Q_FDP0UA U5959 ( .D(n209), .QTFCLK( ), .Q(ofifoData[573]));
Q_FDP0UA U5960 ( .D(n208), .QTFCLK( ), .Q(ofifoData[574]));
Q_FDP0UA U5961 ( .D(n207), .QTFCLK( ), .Q(ofifoData[575]));
Q_MX08 U5962 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[0]), .A1(ofifoData[64]), .A2(ofifoData[128]), .A3(ofifoData[192]), .A4(ofifoData[256]), .A5(ofifoData[320]), .A6(ofifoData[384]), .A7(ofifoData[448]), .Z(n64));
Q_MX02 U5963 ( .S(oFill[4]), .A0(n64), .A1(ofifoData[512]), .Z(n63));
Q_MX08 U5964 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[1]), .A1(ofifoData[65]), .A2(ofifoData[129]), .A3(ofifoData[193]), .A4(ofifoData[257]), .A5(ofifoData[321]), .A6(ofifoData[385]), .A7(ofifoData[449]), .Z(n62));
Q_MX02 U5965 ( .S(oFill[4]), .A0(n62), .A1(ofifoData[513]), .Z(n61));
Q_MX08 U5966 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[2]), .A1(ofifoData[66]), .A2(ofifoData[130]), .A3(ofifoData[194]), .A4(ofifoData[258]), .A5(ofifoData[322]), .A6(ofifoData[386]), .A7(ofifoData[450]), .Z(n60));
Q_MX02 U5967 ( .S(oFill[4]), .A0(n60), .A1(ofifoData[514]), .Z(n59));
Q_MX08 U5968 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[3]), .A1(ofifoData[67]), .A2(ofifoData[131]), .A3(ofifoData[195]), .A4(ofifoData[259]), .A5(ofifoData[323]), .A6(ofifoData[387]), .A7(ofifoData[451]), .Z(n58));
Q_MX02 U5969 ( .S(oFill[4]), .A0(n58), .A1(ofifoData[515]), .Z(n57));
Q_MX08 U5970 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[4]), .A1(ofifoData[68]), .A2(ofifoData[132]), .A3(ofifoData[196]), .A4(ofifoData[260]), .A5(ofifoData[324]), .A6(ofifoData[388]), .A7(ofifoData[452]), .Z(n56));
Q_MX02 U5971 ( .S(oFill[4]), .A0(n56), .A1(ofifoData[516]), .Z(n55));
Q_MX08 U5972 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[5]), .A1(ofifoData[69]), .A2(ofifoData[133]), .A3(ofifoData[197]), .A4(ofifoData[261]), .A5(ofifoData[325]), .A6(ofifoData[389]), .A7(ofifoData[453]), .Z(n54));
Q_MX02 U5973 ( .S(oFill[4]), .A0(n54), .A1(ofifoData[517]), .Z(n53));
Q_MX08 U5974 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[6]), .A1(ofifoData[70]), .A2(ofifoData[134]), .A3(ofifoData[198]), .A4(ofifoData[262]), .A5(ofifoData[326]), .A6(ofifoData[390]), .A7(ofifoData[454]), .Z(n52));
Q_MX02 U5975 ( .S(oFill[4]), .A0(n52), .A1(ofifoData[518]), .Z(n51));
Q_MX08 U5976 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[7]), .A1(ofifoData[71]), .A2(ofifoData[135]), .A3(ofifoData[199]), .A4(ofifoData[263]), .A5(ofifoData[327]), .A6(ofifoData[391]), .A7(ofifoData[455]), .Z(n50));
Q_MX02 U5977 ( .S(oFill[4]), .A0(n50), .A1(ofifoData[519]), .Z(n49));
Q_MX08 U5978 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[8]), .A1(ofifoData[72]), .A2(ofifoData[136]), .A3(ofifoData[200]), .A4(ofifoData[264]), .A5(ofifoData[328]), .A6(ofifoData[392]), .A7(ofifoData[456]), .Z(n48));
Q_MX02 U5979 ( .S(oFill[4]), .A0(n48), .A1(ofifoData[520]), .Z(n47));
Q_MX08 U5980 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[9]), .A1(ofifoData[73]), .A2(ofifoData[137]), .A3(ofifoData[201]), .A4(ofifoData[265]), .A5(ofifoData[329]), .A6(ofifoData[393]), .A7(ofifoData[457]), .Z(n46));
Q_MX02 U5981 ( .S(oFill[4]), .A0(n46), .A1(ofifoData[521]), .Z(n45));
Q_MX08 U5982 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[10]), .A1(ofifoData[74]), .A2(ofifoData[138]), .A3(ofifoData[202]), .A4(ofifoData[266]), .A5(ofifoData[330]), .A6(ofifoData[394]), .A7(ofifoData[458]), .Z(n44));
Q_MX02 U5983 ( .S(oFill[4]), .A0(n44), .A1(ofifoData[522]), .Z(n43));
Q_MX08 U5984 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[11]), .A1(ofifoData[75]), .A2(ofifoData[139]), .A3(ofifoData[203]), .A4(ofifoData[267]), .A5(ofifoData[331]), .A6(ofifoData[395]), .A7(ofifoData[459]), .Z(n42));
Q_MX02 U5985 ( .S(oFill[4]), .A0(n42), .A1(ofifoData[523]), .Z(n41));
Q_MX08 U5986 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[12]), .A1(ofifoData[76]), .A2(ofifoData[140]), .A3(ofifoData[204]), .A4(ofifoData[268]), .A5(ofifoData[332]), .A6(ofifoData[396]), .A7(ofifoData[460]), .Z(n40));
Q_MX02 U5987 ( .S(oFill[4]), .A0(n40), .A1(ofifoData[524]), .Z(n39));
Q_MX08 U5988 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[13]), .A1(ofifoData[77]), .A2(ofifoData[141]), .A3(ofifoData[205]), .A4(ofifoData[269]), .A5(ofifoData[333]), .A6(ofifoData[397]), .A7(ofifoData[461]), .Z(n38));
Q_MX02 U5989 ( .S(oFill[4]), .A0(n38), .A1(ofifoData[525]), .Z(n37));
Q_MX08 U5990 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[14]), .A1(ofifoData[78]), .A2(ofifoData[142]), .A3(ofifoData[206]), .A4(ofifoData[270]), .A5(ofifoData[334]), .A6(ofifoData[398]), .A7(ofifoData[462]), .Z(n36));
Q_MX02 U5991 ( .S(oFill[4]), .A0(n36), .A1(ofifoData[526]), .Z(n35));
Q_MX08 U5992 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[15]), .A1(ofifoData[79]), .A2(ofifoData[143]), .A3(ofifoData[207]), .A4(ofifoData[271]), .A5(ofifoData[335]), .A6(ofifoData[399]), .A7(ofifoData[463]), .Z(n34));
Q_MX02 U5993 ( .S(oFill[4]), .A0(n34), .A1(ofifoData[527]), .Z(n33));
Q_MX08 U5994 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[16]), .A1(ofifoData[80]), .A2(ofifoData[144]), .A3(ofifoData[208]), .A4(ofifoData[272]), .A5(ofifoData[336]), .A6(ofifoData[400]), .A7(ofifoData[464]), .Z(n32));
Q_MX02 U5995 ( .S(oFill[4]), .A0(n32), .A1(ofifoData[528]), .Z(n31));
Q_MX08 U5996 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[17]), .A1(ofifoData[81]), .A2(ofifoData[145]), .A3(ofifoData[209]), .A4(ofifoData[273]), .A5(ofifoData[337]), .A6(ofifoData[401]), .A7(ofifoData[465]), .Z(n30));
Q_MX02 U5997 ( .S(oFill[4]), .A0(n30), .A1(ofifoData[529]), .Z(n29));
Q_MX08 U5998 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[18]), .A1(ofifoData[82]), .A2(ofifoData[146]), .A3(ofifoData[210]), .A4(ofifoData[274]), .A5(ofifoData[338]), .A6(ofifoData[402]), .A7(ofifoData[466]), .Z(n28));
Q_MX02 U5999 ( .S(oFill[4]), .A0(n28), .A1(ofifoData[530]), .Z(n27));
Q_MX08 U6000 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[19]), .A1(ofifoData[83]), .A2(ofifoData[147]), .A3(ofifoData[211]), .A4(ofifoData[275]), .A5(ofifoData[339]), .A6(ofifoData[403]), .A7(ofifoData[467]), .Z(n26));
Q_MX02 U6001 ( .S(oFill[4]), .A0(n26), .A1(ofifoData[531]), .Z(n25));
Q_MX08 U6002 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[20]), .A1(ofifoData[84]), .A2(ofifoData[148]), .A3(ofifoData[212]), .A4(ofifoData[276]), .A5(ofifoData[340]), .A6(ofifoData[404]), .A7(ofifoData[468]), .Z(n24));
Q_MX02 U6003 ( .S(oFill[4]), .A0(n24), .A1(ofifoData[532]), .Z(n23));
Q_MX08 U6004 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[21]), .A1(ofifoData[85]), .A2(ofifoData[149]), .A3(ofifoData[213]), .A4(ofifoData[277]), .A5(ofifoData[341]), .A6(ofifoData[405]), .A7(ofifoData[469]), .Z(n22));
Q_MX02 U6005 ( .S(oFill[4]), .A0(n22), .A1(ofifoData[533]), .Z(n21));
Q_MX08 U6006 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[22]), .A1(ofifoData[86]), .A2(ofifoData[150]), .A3(ofifoData[214]), .A4(ofifoData[278]), .A5(ofifoData[342]), .A6(ofifoData[406]), .A7(ofifoData[470]), .Z(n20));
Q_MX02 U6007 ( .S(oFill[4]), .A0(n20), .A1(ofifoData[534]), .Z(n19));
Q_MX08 U6008 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[23]), .A1(ofifoData[87]), .A2(ofifoData[151]), .A3(ofifoData[215]), .A4(ofifoData[279]), .A5(ofifoData[343]), .A6(ofifoData[407]), .A7(ofifoData[471]), .Z(n18));
Q_MX02 U6009 ( .S(oFill[4]), .A0(n18), .A1(ofifoData[535]), .Z(n17));
Q_MX08 U6010 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[24]), .A1(ofifoData[88]), .A2(ofifoData[152]), .A3(ofifoData[216]), .A4(ofifoData[280]), .A5(ofifoData[344]), .A6(ofifoData[408]), .A7(ofifoData[472]), .Z(n16));
Q_MX02 U6011 ( .S(oFill[4]), .A0(n16), .A1(ofifoData[536]), .Z(n15));
Q_MX08 U6012 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[25]), .A1(ofifoData[89]), .A2(ofifoData[153]), .A3(ofifoData[217]), .A4(ofifoData[281]), .A5(ofifoData[345]), .A6(ofifoData[409]), .A7(ofifoData[473]), .Z(n14));
Q_MX02 U6013 ( .S(oFill[4]), .A0(n14), .A1(ofifoData[537]), .Z(n13));
Q_MX08 U6014 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[26]), .A1(ofifoData[90]), .A2(ofifoData[154]), .A3(ofifoData[218]), .A4(ofifoData[282]), .A5(ofifoData[346]), .A6(ofifoData[410]), .A7(ofifoData[474]), .Z(n12));
Q_MX02 U6015 ( .S(oFill[4]), .A0(n12), .A1(ofifoData[538]), .Z(n11));
Q_MX08 U6016 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[27]), .A1(ofifoData[91]), .A2(ofifoData[155]), .A3(ofifoData[219]), .A4(ofifoData[283]), .A5(ofifoData[347]), .A6(ofifoData[411]), .A7(ofifoData[475]), .Z(n10));
Q_MX02 U6017 ( .S(oFill[4]), .A0(n10), .A1(ofifoData[539]), .Z(n9));
Q_MX08 U6018 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[28]), .A1(ofifoData[92]), .A2(ofifoData[156]), .A3(ofifoData[220]), .A4(ofifoData[284]), .A5(ofifoData[348]), .A6(ofifoData[412]), .A7(ofifoData[476]), .Z(n8));
Q_MX02 U6019 ( .S(oFill[4]), .A0(n8), .A1(ofifoData[540]), .Z(n7));
Q_MX08 U6020 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[29]), .A1(ofifoData[93]), .A2(ofifoData[157]), .A3(ofifoData[221]), .A4(ofifoData[285]), .A5(ofifoData[349]), .A6(ofifoData[413]), .A7(ofifoData[477]), .Z(n6));
Q_MX02 U6021 ( .S(oFill[4]), .A0(n6), .A1(ofifoData[541]), .Z(n5));
Q_MX08 U6022 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[30]), .A1(ofifoData[94]), .A2(ofifoData[158]), .A3(ofifoData[222]), .A4(ofifoData[286]), .A5(ofifoData[350]), .A6(ofifoData[414]), .A7(ofifoData[478]), .Z(n4));
Q_MX02 U6023 ( .S(oFill[4]), .A0(n4), .A1(ofifoData[542]), .Z(n3));
Q_MX08 U6024 ( .S0(oFill[1]), .S1(oFill[2]), .S2(oFill[3]), .A0(ofifoData[31]), .A1(ofifoData[95]), .A2(ofifoData[159]), .A3(ofifoData[223]), .A4(ofifoData[287]), .A5(ofifoData[351]), .A6(ofifoData[415]), .A7(ofifoData[479]), .Z(n2));
Q_MX02 U6025 ( .S(oFill[4]), .A0(n2), .A1(ofifoData[543]), .Z(n1));
Q_XOR2 U6026 ( .A0(n2163), .A1(n2156), .Z(n2162));
Q_OR02 U6027 ( .A0(n788), .A1(GFlen[11]), .Z(n2620));
Q_XOR2 U6028 ( .A0(writeLen[4]), .A1(n3202), .Z(oFillN[4]));
Q_AN02 U6029 ( .A0(ofifoAddr0N[1]), .A1(ofifoAddr0N[0]), .Z(n3261));
Q_AN02 U6030 ( .A0(ofifoAddr0N[2]), .A1(n3232), .Z(n3288));
Q_AN02 U6031 ( .A0(ofifoAddr0N[2]), .A1(ofifoAddr0N[1]), .Z(n3302));
Q_AN02 U6032 ( .A0(ofifoAddr0N[2]), .A1(n3261), .Z(n3316));
`ifdef CBV

reg [63:0] ixc_gfm_ctl [0:0];
always @(n3317 or wrtCntD[63] or wrtCntD[62] or wrtCntD[61] or wrtCntD[60]
 or wrtCntD[59] or wrtCntD[58] or wrtCntD[57] or wrtCntD[56] or wrtCntD[55] or wrtCntD[54] or wrtCntD[53] or wrtCntD[52]
 or wrtCntD[51] or wrtCntD[50] or wrtCntD[49] or wrtCntD[48] or wrtCntD[47] or wrtCntD[46] or wrtCntD[45] or wrtCntD[44]
 or wrtCntD[43] or wrtCntD[42] or wrtCntD[41] or wrtCntD[40] or wrtCntD[39] or wrtCntD[38] or wrtCntD[37] or wrtCntD[36]
 or wrtCntD[35] or wrtCntD[34] or wrtCntD[33] or wrtCntD[32] or wrtCntD[31] or wrtCntD[30] or wrtCntD[29] or wrtCntD[28]
 or wrtCntD[27] or wrtCntD[26] or wrtCntD[25] or wrtCntD[24] or wrtCntD[23] or wrtCntD[22] or wrtCntD[21] or wrtCntD[20]
 or wrtCntD[19] or wrtCntD[18] or wrtCntD[17] or wrtCntD[16] or wrtCntD[15] or wrtCntD[14] or wrtCntD[13] or wrtCntD[12]
 or wrtCntD[11] or wrtCntD[10] or wrtCntD[9] or wrtCntD[8] or wrtCntD[7] or wrtCntD[6] or wrtCntD[5] or wrtCntD[4]
 or wrtCntD[3] or wrtCntD[2] or wrtCntD[1] or wrtCntD[0] or n3318)
#0 begin
if (n3318)
ixc_gfm_ctl[{n3317}] =
{wrtCntD[63], wrtCntD[62], wrtCntD[61], wrtCntD[60], wrtCntD[59],
 wrtCntD[58], wrtCntD[57], wrtCntD[56], wrtCntD[55], wrtCntD[54], wrtCntD[53], wrtCntD[52], wrtCntD[51],
 wrtCntD[50], wrtCntD[49], wrtCntD[48], wrtCntD[47], wrtCntD[46], wrtCntD[45], wrtCntD[44], wrtCntD[43],
 wrtCntD[42], wrtCntD[41], wrtCntD[40], wrtCntD[39], wrtCntD[38], wrtCntD[37], wrtCntD[36], wrtCntD[35],
 wrtCntD[34], wrtCntD[33], wrtCntD[32], wrtCntD[31], wrtCntD[30], wrtCntD[29], wrtCntD[28], wrtCntD[27],
 wrtCntD[26], wrtCntD[25], wrtCntD[24], wrtCntD[23], wrtCntD[22], wrtCntD[21], wrtCntD[20], wrtCntD[19],
 wrtCntD[18], wrtCntD[17], wrtCntD[16], wrtCntD[15], wrtCntD[14], wrtCntD[13], wrtCntD[12], wrtCntD[11],
 wrtCntD[10], wrtCntD[9], wrtCntD[8], wrtCntD[7], wrtCntD[6], wrtCntD[5], wrtCntD[4], wrtCntD[3],
 wrtCntD[2], wrtCntD[1], wrtCntD[0]};
end
`else

MPW2X64 ixc_gfm_ctl ( .A0(n3317), .DI63(wrtCntD[63]), .DI62(wrtCntD[62]), .DI61(wrtCntD[61]), .DI60(wrtCntD[60]), .DI59(wrtCntD[59]),
 .DI58(wrtCntD[58]), .DI57(wrtCntD[57]), .DI56(wrtCntD[56]), .DI55(wrtCntD[55]), .DI54(wrtCntD[54]), .DI53(wrtCntD[53]), .DI52(wrtCntD[52]), .DI51(wrtCntD[51]),
 .DI50(wrtCntD[50]), .DI49(wrtCntD[49]), .DI48(wrtCntD[48]), .DI47(wrtCntD[47]), .DI46(wrtCntD[46]), .DI45(wrtCntD[45]), .DI44(wrtCntD[44]), .DI43(wrtCntD[43]),
 .DI42(wrtCntD[42]), .DI41(wrtCntD[41]), .DI40(wrtCntD[40]), .DI39(wrtCntD[39]), .DI38(wrtCntD[38]), .DI37(wrtCntD[37]), .DI36(wrtCntD[36]), .DI35(wrtCntD[35]),
 .DI34(wrtCntD[34]), .DI33(wrtCntD[33]), .DI32(wrtCntD[32]), .DI31(wrtCntD[31]), .DI30(wrtCntD[30]), .DI29(wrtCntD[29]), .DI28(wrtCntD[28]), .DI27(wrtCntD[27]),
 .DI26(wrtCntD[26]), .DI25(wrtCntD[25]), .DI24(wrtCntD[24]), .DI23(wrtCntD[23]), .DI22(wrtCntD[22]), .DI21(wrtCntD[21]), .DI20(wrtCntD[20]), .DI19(wrtCntD[19]),
 .DI18(wrtCntD[18]), .DI17(wrtCntD[17]), .DI16(wrtCntD[16]), .DI15(wrtCntD[15]), .DI14(wrtCntD[14]), .DI13(wrtCntD[13]), .DI12(wrtCntD[12]), .DI11(wrtCntD[11]),
 .DI10(wrtCntD[10]), .DI9(wrtCntD[9]), .DI8(wrtCntD[8]), .DI7(wrtCntD[7]), .DI6(wrtCntD[6]), .DI5(wrtCntD[5]), .DI4(wrtCntD[4]), .DI3(wrtCntD[3]),
 .DI2(wrtCntD[2]), .DI1(wrtCntD[1]), .DI0(wrtCntD[0]), .WE(n3318), .SYNC_IN(n3317), .SYNC_OUT( ));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ctl" HDL_MEMORY_DECL "1 63 0 0 0"
`endif
`ifdef CBV

reg [63:0] ixc_gfm_ofifo [0:131071];
always @(ofifoAddr0N[16] or ofifoAddr0N[15] or ofifoAddr0N[14] or ofifoAddr0N[13] or ofifoAddr0N[12]
 or ofifoAddr0N[11] or ofifoAddr0N[10] or ofifoAddr0N[9] or ofifoAddr0N[8] or ofifoAddr0N[7] or ofifoAddr0N[6] or ofifoAddr0N[5] or ofifoAddr0N[4]
 or ofifoAddr0N[3] or ofifoAddr0N[2] or ofifoAddr0N[1] or ofifoAddr0N[0] or ofifoDataN[63] or ofifoDataN[62] or ofifoDataN[61] or ofifoDataN[60]
 or ofifoDataN[59] or ofifoDataN[58] or ofifoDataN[57] or ofifoDataN[56] or ofifoDataN[55] or ofifoDataN[54] or ofifoDataN[53] or ofifoDataN[52]
 or ofifoDataN[51] or ofifoDataN[50] or ofifoDataN[49] or ofifoDataN[48] or ofifoDataN[47] or ofifoDataN[46] or ofifoDataN[45] or ofifoDataN[44]
 or ofifoDataN[43] or ofifoDataN[42] or ofifoDataN[41] or ofifoDataN[40] or ofifoDataN[39] or ofifoDataN[38] or ofifoDataN[37] or ofifoDataN[36]
 or ofifoDataN[35] or ofifoDataN[34] or ofifoDataN[33] or ofifoDataN[32] or ofifoDataN[31] or ofifoDataN[30] or ofifoDataN[29] or ofifoDataN[28]
 or ofifoDataN[27] or ofifoDataN[26] or ofifoDataN[25] or ofifoDataN[24] or ofifoDataN[23] or ofifoDataN[22] or ofifoDataN[21] or ofifoDataN[20]
 or ofifoDataN[19] or ofifoDataN[18] or ofifoDataN[17] or ofifoDataN[16] or ofifoDataN[15] or ofifoDataN[14] or ofifoDataN[13] or ofifoDataN[12]
 or ofifoDataN[11] or ofifoDataN[10] or ofifoDataN[9] or ofifoDataN[8] or ofifoDataN[7] or ofifoDataN[6] or ofifoDataN[5] or ofifoDataN[4]
 or ofifoDataN[3] or ofifoDataN[2] or ofifoDataN[1] or ofifoDataN[0] or n3318 or ofifoAddr1N[16] or ofifoAddr1N[15] or ofifoAddr1N[14]
 or ofifoAddr1N[13] or ofifoAddr1N[12] or ofifoAddr1N[11] or ofifoAddr1N[10] or ofifoAddr1N[9] or ofifoAddr1N[8] or ofifoAddr1N[7] or ofifoAddr1N[6]
 or ofifoAddr1N[5] or ofifoAddr1N[4] or ofifoAddr1N[3] or ofifoAddr1N[2] or ofifoAddr1N[1] or ofifoAddr7N[0] or ofifoDataN[127] or ofifoDataN[126]
 or ofifoDataN[125] or ofifoDataN[124] or ofifoDataN[123] or ofifoDataN[122] or ofifoDataN[121] or ofifoDataN[120] or ofifoDataN[119] or ofifoDataN[118]
 or ofifoDataN[117] or ofifoDataN[116] or ofifoDataN[115] or ofifoDataN[114] or ofifoDataN[113] or ofifoDataN[112] or ofifoDataN[111] or ofifoDataN[110]
 or ofifoDataN[109] or ofifoDataN[108] or ofifoDataN[107] or ofifoDataN[106] or ofifoDataN[105] or ofifoDataN[104] or ofifoDataN[103] or ofifoDataN[102]
 or ofifoDataN[101] or ofifoDataN[100] or ofifoDataN[99] or ofifoDataN[98] or ofifoDataN[97] or ofifoDataN[96] or ofifoDataN[95] or ofifoDataN[94]
 or ofifoDataN[93] or ofifoDataN[92] or ofifoDataN[91] or ofifoDataN[90] or ofifoDataN[89] or ofifoDataN[88] or ofifoDataN[87] or ofifoDataN[86]
 or ofifoDataN[85] or ofifoDataN[84] or ofifoDataN[83] or ofifoDataN[82] or ofifoDataN[81] or ofifoDataN[80] or ofifoDataN[79] or ofifoDataN[78]
 or ofifoDataN[77] or ofifoDataN[76] or ofifoDataN[75] or ofifoDataN[74] or ofifoDataN[73] or ofifoDataN[72] or ofifoDataN[71] or ofifoDataN[70]
 or ofifoDataN[69] or ofifoDataN[68] or ofifoDataN[67] or ofifoDataN[66] or ofifoDataN[65] or ofifoDataN[64] or ofifoAddr2N[16] or ofifoAddr2N[15]
 or ofifoAddr2N[14] or ofifoAddr2N[13] or ofifoAddr2N[12] or ofifoAddr2N[11] or ofifoAddr2N[10] or ofifoAddr2N[9] or ofifoAddr2N[8] or ofifoAddr2N[7]
 or ofifoAddr2N[6] or ofifoAddr2N[5] or ofifoAddr2N[4] or ofifoAddr2N[3] or ofifoAddr2N[2] or ofifoAddr6N[1] or ofifoDataN[191] or ofifoDataN[190]
 or ofifoDataN[189] or ofifoDataN[188] or ofifoDataN[187] or ofifoDataN[186] or ofifoDataN[185] or ofifoDataN[184] or ofifoDataN[183] or ofifoDataN[182]
 or ofifoDataN[181] or ofifoDataN[180] or ofifoDataN[179] or ofifoDataN[178] or ofifoDataN[177] or ofifoDataN[176] or ofifoDataN[175] or ofifoDataN[174]
 or ofifoDataN[173] or ofifoDataN[172] or ofifoDataN[171] or ofifoDataN[170] or ofifoDataN[169] or ofifoDataN[168] or ofifoDataN[167] or ofifoDataN[166]
 or ofifoDataN[165] or ofifoDataN[164] or ofifoDataN[163] or ofifoDataN[162] or ofifoDataN[161] or ofifoDataN[160] or ofifoDataN[159] or ofifoDataN[158]
 or ofifoDataN[157] or ofifoDataN[156] or ofifoDataN[155] or ofifoDataN[154] or ofifoDataN[153] or ofifoDataN[152] or ofifoDataN[151] or ofifoDataN[150]
 or ofifoDataN[149] or ofifoDataN[148] or ofifoDataN[147] or ofifoDataN[146] or ofifoDataN[145] or ofifoDataN[144] or ofifoDataN[143] or ofifoDataN[142]
 or ofifoDataN[141] or ofifoDataN[140] or ofifoDataN[139] or ofifoDataN[138] or ofifoDataN[137] or ofifoDataN[136] or ofifoDataN[135] or ofifoDataN[134]
 or ofifoDataN[133] or ofifoDataN[132] or ofifoDataN[131] or ofifoDataN[130] or ofifoDataN[129] or ofifoDataN[128] or ofifoAddr3N[16] or ofifoAddr3N[15]
 or ofifoAddr3N[14] or ofifoAddr3N[13] or ofifoAddr3N[12] or ofifoAddr3N[11] or ofifoAddr3N[10] or ofifoAddr3N[9] or ofifoAddr3N[8] or ofifoAddr3N[7]
 or ofifoAddr3N[6] or ofifoAddr3N[5] or ofifoAddr3N[4] or ofifoAddr3N[3] or ofifoAddr3N[2] or ofifoAddr7N[1] or ofifoDataN[255] or ofifoDataN[254]
 or ofifoDataN[253] or ofifoDataN[252] or ofifoDataN[251] or ofifoDataN[250] or ofifoDataN[249] or ofifoDataN[248] or ofifoDataN[247] or ofifoDataN[246]
 or ofifoDataN[245] or ofifoDataN[244] or ofifoDataN[243] or ofifoDataN[242] or ofifoDataN[241] or ofifoDataN[240] or ofifoDataN[239] or ofifoDataN[238]
 or ofifoDataN[237] or ofifoDataN[236] or ofifoDataN[235] or ofifoDataN[234] or ofifoDataN[233] or ofifoDataN[232] or ofifoDataN[231] or ofifoDataN[230]
 or ofifoDataN[229] or ofifoDataN[228] or ofifoDataN[227] or ofifoDataN[226] or ofifoDataN[225] or ofifoDataN[224] or ofifoDataN[223] or ofifoDataN[222]
 or ofifoDataN[221] or ofifoDataN[220] or ofifoDataN[219] or ofifoDataN[218] or ofifoDataN[217] or ofifoDataN[216] or ofifoDataN[215] or ofifoDataN[214]
 or ofifoDataN[213] or ofifoDataN[212] or ofifoDataN[211] or ofifoDataN[210] or ofifoDataN[209] or ofifoDataN[208] or ofifoDataN[207] or ofifoDataN[206]
 or ofifoDataN[205] or ofifoDataN[204] or ofifoDataN[203] or ofifoDataN[202] or ofifoDataN[201] or ofifoDataN[200] or ofifoDataN[199] or ofifoDataN[198]
 or ofifoDataN[197] or ofifoDataN[196] or ofifoDataN[195] or ofifoDataN[194] or ofifoDataN[193] or ofifoDataN[192] or ofifoAddr4N[16] or ofifoAddr4N[15]
 or ofifoAddr4N[14] or ofifoAddr4N[13] or ofifoAddr4N[12] or ofifoAddr4N[11] or ofifoAddr4N[10] or ofifoAddr4N[9] or ofifoAddr4N[8] or ofifoAddr4N[7]
 or ofifoAddr4N[6] or ofifoAddr4N[5] or ofifoAddr4N[4] or ofifoAddr4N[3] or ofifoAddr4N[2] or ofifoDataN[319] or ofifoDataN[318] or ofifoDataN[317]
 or ofifoDataN[316] or ofifoDataN[315] or ofifoDataN[314] or ofifoDataN[313] or ofifoDataN[312] or ofifoDataN[311] or ofifoDataN[310] or ofifoDataN[309]
 or ofifoDataN[308] or ofifoDataN[307] or ofifoDataN[306] or ofifoDataN[305] or ofifoDataN[304] or ofifoDataN[303] or ofifoDataN[302] or ofifoDataN[301]
 or ofifoDataN[300] or ofifoDataN[299] or ofifoDataN[298] or ofifoDataN[297] or ofifoDataN[296] or ofifoDataN[295] or ofifoDataN[294] or ofifoDataN[293]
 or ofifoDataN[292] or ofifoDataN[291] or ofifoDataN[290] or ofifoDataN[289] or ofifoDataN[288] or ofifoDataN[287] or ofifoDataN[286] or ofifoDataN[285]
 or ofifoDataN[284] or ofifoDataN[283] or ofifoDataN[282] or ofifoDataN[281] or ofifoDataN[280] or ofifoDataN[279] or ofifoDataN[278] or ofifoDataN[277]
 or ofifoDataN[276] or ofifoDataN[275] or ofifoDataN[274] or ofifoDataN[273] or ofifoDataN[272] or ofifoDataN[271] or ofifoDataN[270] or ofifoDataN[269]
 or ofifoDataN[268] or ofifoDataN[267] or ofifoDataN[266] or ofifoDataN[265] or ofifoDataN[264] or ofifoDataN[263] or ofifoDataN[262] or ofifoDataN[261]
 or ofifoDataN[260] or ofifoDataN[259] or ofifoDataN[258] or ofifoDataN[257] or ofifoDataN[256] or ofifoAddr5N[16] or ofifoAddr5N[15] or ofifoAddr5N[14]
 or ofifoAddr5N[13] or ofifoAddr5N[12] or ofifoAddr5N[11] or ofifoAddr5N[10] or ofifoAddr5N[9] or ofifoAddr5N[8] or ofifoAddr5N[7] or ofifoAddr5N[6]
 or ofifoAddr5N[5] or ofifoAddr5N[4] or ofifoAddr5N[3] or ofifoAddr5N[2] or ofifoDataN[383] or ofifoDataN[382] or ofifoDataN[381] or ofifoDataN[380]
 or ofifoDataN[379] or ofifoDataN[378] or ofifoDataN[377] or ofifoDataN[376] or ofifoDataN[375] or ofifoDataN[374] or ofifoDataN[373] or ofifoDataN[372]
 or ofifoDataN[371] or ofifoDataN[370] or ofifoDataN[369] or ofifoDataN[368] or ofifoDataN[367] or ofifoDataN[366] or ofifoDataN[365] or ofifoDataN[364]
 or ofifoDataN[363] or ofifoDataN[362] or ofifoDataN[361] or ofifoDataN[360] or ofifoDataN[359] or ofifoDataN[358] or ofifoDataN[357] or ofifoDataN[356]
 or ofifoDataN[355] or ofifoDataN[354] or ofifoDataN[353] or ofifoDataN[352] or ofifoDataN[351] or ofifoDataN[350] or ofifoDataN[349] or ofifoDataN[348]
 or ofifoDataN[347] or ofifoDataN[346] or ofifoDataN[345] or ofifoDataN[344] or ofifoDataN[343] or ofifoDataN[342] or ofifoDataN[341] or ofifoDataN[340]
 or ofifoDataN[339] or ofifoDataN[338] or ofifoDataN[337] or ofifoDataN[336] or ofifoDataN[335] or ofifoDataN[334] or ofifoDataN[333] or ofifoDataN[332]
 or ofifoDataN[331] or ofifoDataN[330] or ofifoDataN[329] or ofifoDataN[328] or ofifoDataN[327] or ofifoDataN[326] or ofifoDataN[325] or ofifoDataN[324]
 or ofifoDataN[323] or ofifoDataN[322] or ofifoDataN[321] or ofifoDataN[320] or ofifoAddr6N[16] or ofifoAddr6N[15] or ofifoAddr6N[14] or ofifoAddr6N[13]
 or ofifoAddr6N[12] or ofifoAddr6N[11] or ofifoAddr6N[10] or ofifoAddr6N[9] or ofifoAddr6N[8] or ofifoAddr6N[7] or ofifoAddr6N[6] or ofifoAddr6N[5]
 or ofifoAddr6N[4] or ofifoAddr6N[3] or ofifoAddr6N[2] or ofifoDataN[447] or ofifoDataN[446] or ofifoDataN[445] or ofifoDataN[444] or ofifoDataN[443]
 or ofifoDataN[442] or ofifoDataN[441] or ofifoDataN[440] or ofifoDataN[439] or ofifoDataN[438] or ofifoDataN[437] or ofifoDataN[436] or ofifoDataN[435]
 or ofifoDataN[434] or ofifoDataN[433] or ofifoDataN[432] or ofifoDataN[431] or ofifoDataN[430] or ofifoDataN[429] or ofifoDataN[428] or ofifoDataN[427]
 or ofifoDataN[426] or ofifoDataN[425] or ofifoDataN[424] or ofifoDataN[423] or ofifoDataN[422] or ofifoDataN[421] or ofifoDataN[420] or ofifoDataN[419]
 or ofifoDataN[418] or ofifoDataN[417] or ofifoDataN[416] or ofifoDataN[415] or ofifoDataN[414] or ofifoDataN[413] or ofifoDataN[412] or ofifoDataN[411]
 or ofifoDataN[410] or ofifoDataN[409] or ofifoDataN[408] or ofifoDataN[407] or ofifoDataN[406] or ofifoDataN[405] or ofifoDataN[404] or ofifoDataN[403]
 or ofifoDataN[402] or ofifoDataN[401] or ofifoDataN[400] or ofifoDataN[399] or ofifoDataN[398] or ofifoDataN[397] or ofifoDataN[396] or ofifoDataN[395]
 or ofifoDataN[394] or ofifoDataN[393] or ofifoDataN[392] or ofifoDataN[391] or ofifoDataN[390] or ofifoDataN[389] or ofifoDataN[388] or ofifoDataN[387]
 or ofifoDataN[386] or ofifoDataN[385] or ofifoDataN[384] or ofifoAddr7N[16] or ofifoAddr7N[15] or ofifoAddr7N[14] or ofifoAddr7N[13] or ofifoAddr7N[12]
 or ofifoAddr7N[11] or ofifoAddr7N[10] or ofifoAddr7N[9] or ofifoAddr7N[8] or ofifoAddr7N[7] or ofifoAddr7N[6] or ofifoAddr7N[5] or ofifoAddr7N[4]
 or ofifoAddr7N[3] or ofifoAddr7N[2] or ofifoDataN[511] or ofifoDataN[510] or ofifoDataN[509] or ofifoDataN[508] or ofifoDataN[507] or ofifoDataN[506]
 or ofifoDataN[505] or ofifoDataN[504] or ofifoDataN[503] or ofifoDataN[502] or ofifoDataN[501] or ofifoDataN[500] or ofifoDataN[499] or ofifoDataN[498]
 or ofifoDataN[497] or ofifoDataN[496] or ofifoDataN[495] or ofifoDataN[494] or ofifoDataN[493] or ofifoDataN[492] or ofifoDataN[491] or ofifoDataN[490]
 or ofifoDataN[489] or ofifoDataN[488] or ofifoDataN[487] or ofifoDataN[486] or ofifoDataN[485] or ofifoDataN[484] or ofifoDataN[483] or ofifoDataN[482]
 or ofifoDataN[481] or ofifoDataN[480] or ofifoDataN[479] or ofifoDataN[478] or ofifoDataN[477] or ofifoDataN[476] or ofifoDataN[475] or ofifoDataN[474]
 or ofifoDataN[473] or ofifoDataN[472] or ofifoDataN[471] or ofifoDataN[470] or ofifoDataN[469] or ofifoDataN[468] or ofifoDataN[467] or ofifoDataN[466]
 or ofifoDataN[465] or ofifoDataN[464] or ofifoDataN[463] or ofifoDataN[462] or ofifoDataN[461] or ofifoDataN[460] or ofifoDataN[459] or ofifoDataN[458]
 or ofifoDataN[457] or ofifoDataN[456] or ofifoDataN[455] or ofifoDataN[454] or ofifoDataN[453] or ofifoDataN[452] or ofifoDataN[451] or ofifoDataN[450]
 or ofifoDataN[449] or ofifoDataN[448] or ofifoAddr8N[16] or ofifoAddr8N[15] or ofifoAddr8N[14] or ofifoAddr8N[13] or ofifoAddr8N[12] or ofifoAddr8N[11]
 or ofifoAddr8N[10] or ofifoAddr8N[9] or ofifoAddr8N[8] or ofifoAddr8N[7] or ofifoAddr8N[6] or ofifoAddr8N[5] or ofifoAddr8N[4] or ofifoAddr8N[3]
 or ofifoDataN[575] or ofifoDataN[574] or ofifoDataN[573] or ofifoDataN[572] or ofifoDataN[571] or ofifoDataN[570] or ofifoDataN[569] or ofifoDataN[568]
 or ofifoDataN[567] or ofifoDataN[566] or ofifoDataN[565] or ofifoDataN[564] or ofifoDataN[563] or ofifoDataN[562] or ofifoDataN[561] or ofifoDataN[560]
 or ofifoDataN[559] or ofifoDataN[558] or ofifoDataN[557] or ofifoDataN[556] or ofifoDataN[555] or ofifoDataN[554] or ofifoDataN[553] or ofifoDataN[552]
 or ofifoDataN[551] or ofifoDataN[550] or ofifoDataN[549] or ofifoDataN[548] or ofifoDataN[547] or ofifoDataN[546] or ofifoDataN[545] or ofifoDataN[544]
 or ofifoDataN[543] or ofifoDataN[542] or ofifoDataN[541] or ofifoDataN[540] or ofifoDataN[539] or ofifoDataN[538] or ofifoDataN[537] or ofifoDataN[536]
 or ofifoDataN[535] or ofifoDataN[534] or ofifoDataN[533] or ofifoDataN[532] or ofifoDataN[531] or ofifoDataN[530] or ofifoDataN[529] or ofifoDataN[528]
 or ofifoDataN[527] or ofifoDataN[526] or ofifoDataN[525] or ofifoDataN[524] or ofifoDataN[523] or ofifoDataN[522] or ofifoDataN[521] or ofifoDataN[520]
 or ofifoDataN[519] or ofifoDataN[518] or ofifoDataN[517] or ofifoDataN[516] or ofifoDataN[515] or ofifoDataN[514] or ofifoDataN[513] or ofifoDataN[512])
#0 begin
if (n3318)
ixc_gfm_ofifo[{ofifoAddr0N[16], ofifoAddr0N[15], ofifoAddr0N[14], ofifoAddr0N[13], ofifoAddr0N[12],
 ofifoAddr0N[11], ofifoAddr0N[10], ofifoAddr0N[9], ofifoAddr0N[8], ofifoAddr0N[7], ofifoAddr0N[6], ofifoAddr0N[5], ofifoAddr0N[4],
 ofifoAddr0N[3], ofifoAddr0N[2], ofifoAddr0N[1], ofifoAddr0N[0]}] =
{ofifoDataN[63], ofifoDataN[62], ofifoDataN[61], ofifoDataN[60], ofifoDataN[59],
 ofifoDataN[58], ofifoDataN[57], ofifoDataN[56], ofifoDataN[55], ofifoDataN[54], ofifoDataN[53], ofifoDataN[52], ofifoDataN[51],
 ofifoDataN[50], ofifoDataN[49], ofifoDataN[48], ofifoDataN[47], ofifoDataN[46], ofifoDataN[45], ofifoDataN[44], ofifoDataN[43],
 ofifoDataN[42], ofifoDataN[41], ofifoDataN[40], ofifoDataN[39], ofifoDataN[38], ofifoDataN[37], ofifoDataN[36], ofifoDataN[35],
 ofifoDataN[34], ofifoDataN[33], ofifoDataN[32], ofifoDataN[31], ofifoDataN[30], ofifoDataN[29], ofifoDataN[28], ofifoDataN[27],
 ofifoDataN[26], ofifoDataN[25], ofifoDataN[24], ofifoDataN[23], ofifoDataN[22], ofifoDataN[21], ofifoDataN[20], ofifoDataN[19],
 ofifoDataN[18], ofifoDataN[17], ofifoDataN[16], ofifoDataN[15], ofifoDataN[14], ofifoDataN[13], ofifoDataN[12], ofifoDataN[11],
 ofifoDataN[10], ofifoDataN[9], ofifoDataN[8], ofifoDataN[7], ofifoDataN[6], ofifoDataN[5], ofifoDataN[4], ofifoDataN[3],
 ofifoDataN[2], ofifoDataN[1], ofifoDataN[0]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr1N[16], ofifoAddr1N[15], ofifoAddr1N[14], ofifoAddr1N[13], ofifoAddr1N[12],
 ofifoAddr1N[11], ofifoAddr1N[10], ofifoAddr1N[9], ofifoAddr1N[8], ofifoAddr1N[7], ofifoAddr1N[6], ofifoAddr1N[5], ofifoAddr1N[4],
 ofifoAddr1N[3], ofifoAddr1N[2], ofifoAddr1N[1], ofifoAddr7N[0]}] =
{ofifoDataN[127], ofifoDataN[126], ofifoDataN[125], ofifoDataN[124], ofifoDataN[123],
 ofifoDataN[122], ofifoDataN[121], ofifoDataN[120], ofifoDataN[119], ofifoDataN[118], ofifoDataN[117], ofifoDataN[116], ofifoDataN[115],
 ofifoDataN[114], ofifoDataN[113], ofifoDataN[112], ofifoDataN[111], ofifoDataN[110], ofifoDataN[109], ofifoDataN[108], ofifoDataN[107],
 ofifoDataN[106], ofifoDataN[105], ofifoDataN[104], ofifoDataN[103], ofifoDataN[102], ofifoDataN[101], ofifoDataN[100], ofifoDataN[99],
 ofifoDataN[98], ofifoDataN[97], ofifoDataN[96], ofifoDataN[95], ofifoDataN[94], ofifoDataN[93], ofifoDataN[92], ofifoDataN[91],
 ofifoDataN[90], ofifoDataN[89], ofifoDataN[88], ofifoDataN[87], ofifoDataN[86], ofifoDataN[85], ofifoDataN[84], ofifoDataN[83],
 ofifoDataN[82], ofifoDataN[81], ofifoDataN[80], ofifoDataN[79], ofifoDataN[78], ofifoDataN[77], ofifoDataN[76], ofifoDataN[75],
 ofifoDataN[74], ofifoDataN[73], ofifoDataN[72], ofifoDataN[71], ofifoDataN[70], ofifoDataN[69], ofifoDataN[68], ofifoDataN[67],
 ofifoDataN[66], ofifoDataN[65], ofifoDataN[64]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr2N[16], ofifoAddr2N[15], ofifoAddr2N[14], ofifoAddr2N[13], ofifoAddr2N[12],
 ofifoAddr2N[11], ofifoAddr2N[10], ofifoAddr2N[9], ofifoAddr2N[8], ofifoAddr2N[7], ofifoAddr2N[6], ofifoAddr2N[5], ofifoAddr2N[4],
 ofifoAddr2N[3], ofifoAddr2N[2], ofifoAddr6N[1], ofifoAddr0N[0]}] =
{ofifoDataN[191], ofifoDataN[190], ofifoDataN[189], ofifoDataN[188], ofifoDataN[187],
 ofifoDataN[186], ofifoDataN[185], ofifoDataN[184], ofifoDataN[183], ofifoDataN[182], ofifoDataN[181], ofifoDataN[180], ofifoDataN[179],
 ofifoDataN[178], ofifoDataN[177], ofifoDataN[176], ofifoDataN[175], ofifoDataN[174], ofifoDataN[173], ofifoDataN[172], ofifoDataN[171],
 ofifoDataN[170], ofifoDataN[169], ofifoDataN[168], ofifoDataN[167], ofifoDataN[166], ofifoDataN[165], ofifoDataN[164], ofifoDataN[163],
 ofifoDataN[162], ofifoDataN[161], ofifoDataN[160], ofifoDataN[159], ofifoDataN[158], ofifoDataN[157], ofifoDataN[156], ofifoDataN[155],
 ofifoDataN[154], ofifoDataN[153], ofifoDataN[152], ofifoDataN[151], ofifoDataN[150], ofifoDataN[149], ofifoDataN[148], ofifoDataN[147],
 ofifoDataN[146], ofifoDataN[145], ofifoDataN[144], ofifoDataN[143], ofifoDataN[142], ofifoDataN[141], ofifoDataN[140], ofifoDataN[139],
 ofifoDataN[138], ofifoDataN[137], ofifoDataN[136], ofifoDataN[135], ofifoDataN[134], ofifoDataN[133], ofifoDataN[132], ofifoDataN[131],
 ofifoDataN[130], ofifoDataN[129], ofifoDataN[128]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr3N[16], ofifoAddr3N[15], ofifoAddr3N[14], ofifoAddr3N[13], ofifoAddr3N[12],
 ofifoAddr3N[11], ofifoAddr3N[10], ofifoAddr3N[9], ofifoAddr3N[8], ofifoAddr3N[7], ofifoAddr3N[6], ofifoAddr3N[5], ofifoAddr3N[4],
 ofifoAddr3N[3], ofifoAddr3N[2], ofifoAddr7N[1], ofifoAddr7N[0]}] =
{ofifoDataN[255], ofifoDataN[254], ofifoDataN[253], ofifoDataN[252], ofifoDataN[251],
 ofifoDataN[250], ofifoDataN[249], ofifoDataN[248], ofifoDataN[247], ofifoDataN[246], ofifoDataN[245], ofifoDataN[244], ofifoDataN[243],
 ofifoDataN[242], ofifoDataN[241], ofifoDataN[240], ofifoDataN[239], ofifoDataN[238], ofifoDataN[237], ofifoDataN[236], ofifoDataN[235],
 ofifoDataN[234], ofifoDataN[233], ofifoDataN[232], ofifoDataN[231], ofifoDataN[230], ofifoDataN[229], ofifoDataN[228], ofifoDataN[227],
 ofifoDataN[226], ofifoDataN[225], ofifoDataN[224], ofifoDataN[223], ofifoDataN[222], ofifoDataN[221], ofifoDataN[220], ofifoDataN[219],
 ofifoDataN[218], ofifoDataN[217], ofifoDataN[216], ofifoDataN[215], ofifoDataN[214], ofifoDataN[213], ofifoDataN[212], ofifoDataN[211],
 ofifoDataN[210], ofifoDataN[209], ofifoDataN[208], ofifoDataN[207], ofifoDataN[206], ofifoDataN[205], ofifoDataN[204], ofifoDataN[203],
 ofifoDataN[202], ofifoDataN[201], ofifoDataN[200], ofifoDataN[199], ofifoDataN[198], ofifoDataN[197], ofifoDataN[196], ofifoDataN[195],
 ofifoDataN[194], ofifoDataN[193], ofifoDataN[192]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr4N[16], ofifoAddr4N[15], ofifoAddr4N[14], ofifoAddr4N[13], ofifoAddr4N[12],
 ofifoAddr4N[11], ofifoAddr4N[10], ofifoAddr4N[9], ofifoAddr4N[8], ofifoAddr4N[7], ofifoAddr4N[6], ofifoAddr4N[5], ofifoAddr4N[4],
 ofifoAddr4N[3], ofifoAddr4N[2], ofifoAddr0N[1], ofifoAddr0N[0]}] =
{ofifoDataN[319], ofifoDataN[318], ofifoDataN[317], ofifoDataN[316], ofifoDataN[315],
 ofifoDataN[314], ofifoDataN[313], ofifoDataN[312], ofifoDataN[311], ofifoDataN[310], ofifoDataN[309], ofifoDataN[308], ofifoDataN[307],
 ofifoDataN[306], ofifoDataN[305], ofifoDataN[304], ofifoDataN[303], ofifoDataN[302], ofifoDataN[301], ofifoDataN[300], ofifoDataN[299],
 ofifoDataN[298], ofifoDataN[297], ofifoDataN[296], ofifoDataN[295], ofifoDataN[294], ofifoDataN[293], ofifoDataN[292], ofifoDataN[291],
 ofifoDataN[290], ofifoDataN[289], ofifoDataN[288], ofifoDataN[287], ofifoDataN[286], ofifoDataN[285], ofifoDataN[284], ofifoDataN[283],
 ofifoDataN[282], ofifoDataN[281], ofifoDataN[280], ofifoDataN[279], ofifoDataN[278], ofifoDataN[277], ofifoDataN[276], ofifoDataN[275],
 ofifoDataN[274], ofifoDataN[273], ofifoDataN[272], ofifoDataN[271], ofifoDataN[270], ofifoDataN[269], ofifoDataN[268], ofifoDataN[267],
 ofifoDataN[266], ofifoDataN[265], ofifoDataN[264], ofifoDataN[263], ofifoDataN[262], ofifoDataN[261], ofifoDataN[260], ofifoDataN[259],
 ofifoDataN[258], ofifoDataN[257], ofifoDataN[256]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr5N[16], ofifoAddr5N[15], ofifoAddr5N[14], ofifoAddr5N[13], ofifoAddr5N[12],
 ofifoAddr5N[11], ofifoAddr5N[10], ofifoAddr5N[9], ofifoAddr5N[8], ofifoAddr5N[7], ofifoAddr5N[6], ofifoAddr5N[5], ofifoAddr5N[4],
 ofifoAddr5N[3], ofifoAddr5N[2], ofifoAddr1N[1], ofifoAddr7N[0]}] =
{ofifoDataN[383], ofifoDataN[382], ofifoDataN[381], ofifoDataN[380], ofifoDataN[379],
 ofifoDataN[378], ofifoDataN[377], ofifoDataN[376], ofifoDataN[375], ofifoDataN[374], ofifoDataN[373], ofifoDataN[372], ofifoDataN[371],
 ofifoDataN[370], ofifoDataN[369], ofifoDataN[368], ofifoDataN[367], ofifoDataN[366], ofifoDataN[365], ofifoDataN[364], ofifoDataN[363],
 ofifoDataN[362], ofifoDataN[361], ofifoDataN[360], ofifoDataN[359], ofifoDataN[358], ofifoDataN[357], ofifoDataN[356], ofifoDataN[355],
 ofifoDataN[354], ofifoDataN[353], ofifoDataN[352], ofifoDataN[351], ofifoDataN[350], ofifoDataN[349], ofifoDataN[348], ofifoDataN[347],
 ofifoDataN[346], ofifoDataN[345], ofifoDataN[344], ofifoDataN[343], ofifoDataN[342], ofifoDataN[341], ofifoDataN[340], ofifoDataN[339],
 ofifoDataN[338], ofifoDataN[337], ofifoDataN[336], ofifoDataN[335], ofifoDataN[334], ofifoDataN[333], ofifoDataN[332], ofifoDataN[331],
 ofifoDataN[330], ofifoDataN[329], ofifoDataN[328], ofifoDataN[327], ofifoDataN[326], ofifoDataN[325], ofifoDataN[324], ofifoDataN[323],
 ofifoDataN[322], ofifoDataN[321], ofifoDataN[320]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr6N[16], ofifoAddr6N[15], ofifoAddr6N[14], ofifoAddr6N[13], ofifoAddr6N[12],
 ofifoAddr6N[11], ofifoAddr6N[10], ofifoAddr6N[9], ofifoAddr6N[8], ofifoAddr6N[7], ofifoAddr6N[6], ofifoAddr6N[5], ofifoAddr6N[4],
 ofifoAddr6N[3], ofifoAddr6N[2], ofifoAddr6N[1], ofifoAddr0N[0]}] =
{ofifoDataN[447], ofifoDataN[446], ofifoDataN[445], ofifoDataN[444], ofifoDataN[443],
 ofifoDataN[442], ofifoDataN[441], ofifoDataN[440], ofifoDataN[439], ofifoDataN[438], ofifoDataN[437], ofifoDataN[436], ofifoDataN[435],
 ofifoDataN[434], ofifoDataN[433], ofifoDataN[432], ofifoDataN[431], ofifoDataN[430], ofifoDataN[429], ofifoDataN[428], ofifoDataN[427],
 ofifoDataN[426], ofifoDataN[425], ofifoDataN[424], ofifoDataN[423], ofifoDataN[422], ofifoDataN[421], ofifoDataN[420], ofifoDataN[419],
 ofifoDataN[418], ofifoDataN[417], ofifoDataN[416], ofifoDataN[415], ofifoDataN[414], ofifoDataN[413], ofifoDataN[412], ofifoDataN[411],
 ofifoDataN[410], ofifoDataN[409], ofifoDataN[408], ofifoDataN[407], ofifoDataN[406], ofifoDataN[405], ofifoDataN[404], ofifoDataN[403],
 ofifoDataN[402], ofifoDataN[401], ofifoDataN[400], ofifoDataN[399], ofifoDataN[398], ofifoDataN[397], ofifoDataN[396], ofifoDataN[395],
 ofifoDataN[394], ofifoDataN[393], ofifoDataN[392], ofifoDataN[391], ofifoDataN[390], ofifoDataN[389], ofifoDataN[388], ofifoDataN[387],
 ofifoDataN[386], ofifoDataN[385], ofifoDataN[384]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr7N[16], ofifoAddr7N[15], ofifoAddr7N[14], ofifoAddr7N[13], ofifoAddr7N[12],
 ofifoAddr7N[11], ofifoAddr7N[10], ofifoAddr7N[9], ofifoAddr7N[8], ofifoAddr7N[7], ofifoAddr7N[6], ofifoAddr7N[5], ofifoAddr7N[4],
 ofifoAddr7N[3], ofifoAddr7N[2], ofifoAddr7N[1], ofifoAddr7N[0]}] =
{ofifoDataN[511], ofifoDataN[510], ofifoDataN[509], ofifoDataN[508], ofifoDataN[507],
 ofifoDataN[506], ofifoDataN[505], ofifoDataN[504], ofifoDataN[503], ofifoDataN[502], ofifoDataN[501], ofifoDataN[500], ofifoDataN[499],
 ofifoDataN[498], ofifoDataN[497], ofifoDataN[496], ofifoDataN[495], ofifoDataN[494], ofifoDataN[493], ofifoDataN[492], ofifoDataN[491],
 ofifoDataN[490], ofifoDataN[489], ofifoDataN[488], ofifoDataN[487], ofifoDataN[486], ofifoDataN[485], ofifoDataN[484], ofifoDataN[483],
 ofifoDataN[482], ofifoDataN[481], ofifoDataN[480], ofifoDataN[479], ofifoDataN[478], ofifoDataN[477], ofifoDataN[476], ofifoDataN[475],
 ofifoDataN[474], ofifoDataN[473], ofifoDataN[472], ofifoDataN[471], ofifoDataN[470], ofifoDataN[469], ofifoDataN[468], ofifoDataN[467],
 ofifoDataN[466], ofifoDataN[465], ofifoDataN[464], ofifoDataN[463], ofifoDataN[462], ofifoDataN[461], ofifoDataN[460], ofifoDataN[459],
 ofifoDataN[458], ofifoDataN[457], ofifoDataN[456], ofifoDataN[455], ofifoDataN[454], ofifoDataN[453], ofifoDataN[452], ofifoDataN[451],
 ofifoDataN[450], ofifoDataN[449], ofifoDataN[448]};
if (n3318)
ixc_gfm_ofifo[{ofifoAddr8N[16], ofifoAddr8N[15], ofifoAddr8N[14], ofifoAddr8N[13], ofifoAddr8N[12],
 ofifoAddr8N[11], ofifoAddr8N[10], ofifoAddr8N[9], ofifoAddr8N[8], ofifoAddr8N[7], ofifoAddr8N[6], ofifoAddr8N[5], ofifoAddr8N[4],
 ofifoAddr8N[3], ofifoAddr0N[2], ofifoAddr0N[1], ofifoAddr0N[0]}] =
{ofifoDataN[575], ofifoDataN[574], ofifoDataN[573], ofifoDataN[572], ofifoDataN[571],
 ofifoDataN[570], ofifoDataN[569], ofifoDataN[568], ofifoDataN[567], ofifoDataN[566], ofifoDataN[565], ofifoDataN[564], ofifoDataN[563],
 ofifoDataN[562], ofifoDataN[561], ofifoDataN[560], ofifoDataN[559], ofifoDataN[558], ofifoDataN[557], ofifoDataN[556], ofifoDataN[555],
 ofifoDataN[554], ofifoDataN[553], ofifoDataN[552], ofifoDataN[551], ofifoDataN[550], ofifoDataN[549], ofifoDataN[548], ofifoDataN[547],
 ofifoDataN[546], ofifoDataN[545], ofifoDataN[544], ofifoDataN[543], ofifoDataN[542], ofifoDataN[541], ofifoDataN[540], ofifoDataN[539],
 ofifoDataN[538], ofifoDataN[537], ofifoDataN[536], ofifoDataN[535], ofifoDataN[534], ofifoDataN[533], ofifoDataN[532], ofifoDataN[531],
 ofifoDataN[530], ofifoDataN[529], ofifoDataN[528], ofifoDataN[527], ofifoDataN[526], ofifoDataN[525], ofifoDataN[524], ofifoDataN[523],
 ofifoDataN[522], ofifoDataN[521], ofifoDataN[520], ofifoDataN[519], ofifoDataN[518], ofifoDataN[517], ofifoDataN[516], ofifoDataN[515],
 ofifoDataN[514], ofifoDataN[513], ofifoDataN[512]};
end
`else

MPW128KX64 ixc_gfm_ofifo ( .A16(ofifoAddr0N[16]), .A15(ofifoAddr0N[15]), .A14(ofifoAddr0N[14]), .A13(ofifoAddr0N[13]), .A12(ofifoAddr0N[12]), .A11(ofifoAddr0N[11]),
 .A10(ofifoAddr0N[10]), .A9(ofifoAddr0N[9]), .A8(ofifoAddr0N[8]), .A7(ofifoAddr0N[7]), .A6(ofifoAddr0N[6]), .A5(ofifoAddr0N[5]), .A4(ofifoAddr0N[4]), .A3(ofifoAddr0N[3]),
 .A2(ofifoAddr0N[2]), .A1(ofifoAddr0N[1]), .A0(ofifoAddr0N[0]), .DI63(ofifoDataN[63]), .DI62(ofifoDataN[62]), .DI61(ofifoDataN[61]), .DI60(ofifoDataN[60]), .DI59(ofifoDataN[59]),
 .DI58(ofifoDataN[58]), .DI57(ofifoDataN[57]), .DI56(ofifoDataN[56]), .DI55(ofifoDataN[55]), .DI54(ofifoDataN[54]), .DI53(ofifoDataN[53]), .DI52(ofifoDataN[52]), .DI51(ofifoDataN[51]),
 .DI50(ofifoDataN[50]), .DI49(ofifoDataN[49]), .DI48(ofifoDataN[48]), .DI47(ofifoDataN[47]), .DI46(ofifoDataN[46]), .DI45(ofifoDataN[45]), .DI44(ofifoDataN[44]), .DI43(ofifoDataN[43]),
 .DI42(ofifoDataN[42]), .DI41(ofifoDataN[41]), .DI40(ofifoDataN[40]), .DI39(ofifoDataN[39]), .DI38(ofifoDataN[38]), .DI37(ofifoDataN[37]), .DI36(ofifoDataN[36]), .DI35(ofifoDataN[35]),
 .DI34(ofifoDataN[34]), .DI33(ofifoDataN[33]), .DI32(ofifoDataN[32]), .DI31(ofifoDataN[31]), .DI30(ofifoDataN[30]), .DI29(ofifoDataN[29]), .DI28(ofifoDataN[28]), .DI27(ofifoDataN[27]),
 .DI26(ofifoDataN[26]), .DI25(ofifoDataN[25]), .DI24(ofifoDataN[24]), .DI23(ofifoDataN[23]), .DI22(ofifoDataN[22]), .DI21(ofifoDataN[21]), .DI20(ofifoDataN[20]), .DI19(ofifoDataN[19]),
 .DI18(ofifoDataN[18]), .DI17(ofifoDataN[17]), .DI16(ofifoDataN[16]), .DI15(ofifoDataN[15]), .DI14(ofifoDataN[14]), .DI13(ofifoDataN[13]), .DI12(ofifoDataN[12]), .DI11(ofifoDataN[11]),
 .DI10(ofifoDataN[10]), .DI9(ofifoDataN[9]), .DI8(ofifoDataN[8]), .DI7(ofifoDataN[7]), .DI6(ofifoDataN[6]), .DI5(ofifoDataN[5]), .DI4(ofifoDataN[4]), .DI3(ofifoDataN[3]),
 .DI2(ofifoDataN[2]), .DI1(ofifoDataN[1]), .DI0(ofifoDataN[0]), .WE(n3318), .SYNC_IN(n3317), .SYNC_OUT(n4790));
// pragma CVASTRPROP INSTANCE "ixc_gfm_ofifo" HDL_MEMORY_DECL "1 63 0 0 131071"
MPW128KX64 U6035 ( .A16(ofifoAddr1N[16]), .A15(ofifoAddr1N[15]), .A14(ofifoAddr1N[14]), .A13(ofifoAddr1N[13]), .A12(ofifoAddr1N[12]), .A11(ofifoAddr1N[11]),
 .A10(ofifoAddr1N[10]), .A9(ofifoAddr1N[9]), .A8(ofifoAddr1N[8]), .A7(ofifoAddr1N[7]), .A6(ofifoAddr1N[6]), .A5(ofifoAddr1N[5]), .A4(ofifoAddr1N[4]), .A3(ofifoAddr1N[3]),
 .A2(ofifoAddr1N[2]), .A1(ofifoAddr1N[1]), .A0(ofifoAddr7N[0]), .DI63(ofifoDataN[127]), .DI62(ofifoDataN[126]), .DI61(ofifoDataN[125]), .DI60(ofifoDataN[124]), .DI59(ofifoDataN[123]),
 .DI58(ofifoDataN[122]), .DI57(ofifoDataN[121]), .DI56(ofifoDataN[120]), .DI55(ofifoDataN[119]), .DI54(ofifoDataN[118]), .DI53(ofifoDataN[117]), .DI52(ofifoDataN[116]), .DI51(ofifoDataN[115]),
 .DI50(ofifoDataN[114]), .DI49(ofifoDataN[113]), .DI48(ofifoDataN[112]), .DI47(ofifoDataN[111]), .DI46(ofifoDataN[110]), .DI45(ofifoDataN[109]), .DI44(ofifoDataN[108]), .DI43(ofifoDataN[107]),
 .DI42(ofifoDataN[106]), .DI41(ofifoDataN[105]), .DI40(ofifoDataN[104]), .DI39(ofifoDataN[103]), .DI38(ofifoDataN[102]), .DI37(ofifoDataN[101]), .DI36(ofifoDataN[100]), .DI35(ofifoDataN[99]),
 .DI34(ofifoDataN[98]), .DI33(ofifoDataN[97]), .DI32(ofifoDataN[96]), .DI31(ofifoDataN[95]), .DI30(ofifoDataN[94]), .DI29(ofifoDataN[93]), .DI28(ofifoDataN[92]), .DI27(ofifoDataN[91]),
 .DI26(ofifoDataN[90]), .DI25(ofifoDataN[89]), .DI24(ofifoDataN[88]), .DI23(ofifoDataN[87]), .DI22(ofifoDataN[86]), .DI21(ofifoDataN[85]), .DI20(ofifoDataN[84]), .DI19(ofifoDataN[83]),
 .DI18(ofifoDataN[82]), .DI17(ofifoDataN[81]), .DI16(ofifoDataN[80]), .DI15(ofifoDataN[79]), .DI14(ofifoDataN[78]), .DI13(ofifoDataN[77]), .DI12(ofifoDataN[76]), .DI11(ofifoDataN[75]),
 .DI10(ofifoDataN[74]), .DI9(ofifoDataN[73]), .DI8(ofifoDataN[72]), .DI7(ofifoDataN[71]), .DI6(ofifoDataN[70]), .DI5(ofifoDataN[69]), .DI4(ofifoDataN[68]), .DI3(ofifoDataN[67]),
 .DI2(ofifoDataN[66]), .DI1(ofifoDataN[65]), .DI0(ofifoDataN[64]), .WE(n3318), .SYNC_IN(n4790), .SYNC_OUT(n4791));
MPW128KX64 U6036 ( .A16(ofifoAddr2N[16]), .A15(ofifoAddr2N[15]), .A14(ofifoAddr2N[14]), .A13(ofifoAddr2N[13]), .A12(ofifoAddr2N[12]), .A11(ofifoAddr2N[11]),
 .A10(ofifoAddr2N[10]), .A9(ofifoAddr2N[9]), .A8(ofifoAddr2N[8]), .A7(ofifoAddr2N[7]), .A6(ofifoAddr2N[6]), .A5(ofifoAddr2N[5]), .A4(ofifoAddr2N[4]), .A3(ofifoAddr2N[3]),
 .A2(ofifoAddr2N[2]), .A1(ofifoAddr6N[1]), .A0(ofifoAddr0N[0]), .DI63(ofifoDataN[191]), .DI62(ofifoDataN[190]), .DI61(ofifoDataN[189]), .DI60(ofifoDataN[188]), .DI59(ofifoDataN[187]),
 .DI58(ofifoDataN[186]), .DI57(ofifoDataN[185]), .DI56(ofifoDataN[184]), .DI55(ofifoDataN[183]), .DI54(ofifoDataN[182]), .DI53(ofifoDataN[181]), .DI52(ofifoDataN[180]), .DI51(ofifoDataN[179]),
 .DI50(ofifoDataN[178]), .DI49(ofifoDataN[177]), .DI48(ofifoDataN[176]), .DI47(ofifoDataN[175]), .DI46(ofifoDataN[174]), .DI45(ofifoDataN[173]), .DI44(ofifoDataN[172]), .DI43(ofifoDataN[171]),
 .DI42(ofifoDataN[170]), .DI41(ofifoDataN[169]), .DI40(ofifoDataN[168]), .DI39(ofifoDataN[167]), .DI38(ofifoDataN[166]), .DI37(ofifoDataN[165]), .DI36(ofifoDataN[164]), .DI35(ofifoDataN[163]),
 .DI34(ofifoDataN[162]), .DI33(ofifoDataN[161]), .DI32(ofifoDataN[160]), .DI31(ofifoDataN[159]), .DI30(ofifoDataN[158]), .DI29(ofifoDataN[157]), .DI28(ofifoDataN[156]), .DI27(ofifoDataN[155]),
 .DI26(ofifoDataN[154]), .DI25(ofifoDataN[153]), .DI24(ofifoDataN[152]), .DI23(ofifoDataN[151]), .DI22(ofifoDataN[150]), .DI21(ofifoDataN[149]), .DI20(ofifoDataN[148]), .DI19(ofifoDataN[147]),
 .DI18(ofifoDataN[146]), .DI17(ofifoDataN[145]), .DI16(ofifoDataN[144]), .DI15(ofifoDataN[143]), .DI14(ofifoDataN[142]), .DI13(ofifoDataN[141]), .DI12(ofifoDataN[140]), .DI11(ofifoDataN[139]),
 .DI10(ofifoDataN[138]), .DI9(ofifoDataN[137]), .DI8(ofifoDataN[136]), .DI7(ofifoDataN[135]), .DI6(ofifoDataN[134]), .DI5(ofifoDataN[133]), .DI4(ofifoDataN[132]), .DI3(ofifoDataN[131]),
 .DI2(ofifoDataN[130]), .DI1(ofifoDataN[129]), .DI0(ofifoDataN[128]), .WE(n3318), .SYNC_IN(n4791), .SYNC_OUT(n4792));
MPW128KX64 U6037 ( .A16(ofifoAddr3N[16]), .A15(ofifoAddr3N[15]), .A14(ofifoAddr3N[14]), .A13(ofifoAddr3N[13]), .A12(ofifoAddr3N[12]), .A11(ofifoAddr3N[11]),
 .A10(ofifoAddr3N[10]), .A9(ofifoAddr3N[9]), .A8(ofifoAddr3N[8]), .A7(ofifoAddr3N[7]), .A6(ofifoAddr3N[6]), .A5(ofifoAddr3N[5]), .A4(ofifoAddr3N[4]), .A3(ofifoAddr3N[3]),
 .A2(ofifoAddr3N[2]), .A1(ofifoAddr7N[1]), .A0(ofifoAddr7N[0]), .DI63(ofifoDataN[255]), .DI62(ofifoDataN[254]), .DI61(ofifoDataN[253]), .DI60(ofifoDataN[252]), .DI59(ofifoDataN[251]),
 .DI58(ofifoDataN[250]), .DI57(ofifoDataN[249]), .DI56(ofifoDataN[248]), .DI55(ofifoDataN[247]), .DI54(ofifoDataN[246]), .DI53(ofifoDataN[245]), .DI52(ofifoDataN[244]), .DI51(ofifoDataN[243]),
 .DI50(ofifoDataN[242]), .DI49(ofifoDataN[241]), .DI48(ofifoDataN[240]), .DI47(ofifoDataN[239]), .DI46(ofifoDataN[238]), .DI45(ofifoDataN[237]), .DI44(ofifoDataN[236]), .DI43(ofifoDataN[235]),
 .DI42(ofifoDataN[234]), .DI41(ofifoDataN[233]), .DI40(ofifoDataN[232]), .DI39(ofifoDataN[231]), .DI38(ofifoDataN[230]), .DI37(ofifoDataN[229]), .DI36(ofifoDataN[228]), .DI35(ofifoDataN[227]),
 .DI34(ofifoDataN[226]), .DI33(ofifoDataN[225]), .DI32(ofifoDataN[224]), .DI31(ofifoDataN[223]), .DI30(ofifoDataN[222]), .DI29(ofifoDataN[221]), .DI28(ofifoDataN[220]), .DI27(ofifoDataN[219]),
 .DI26(ofifoDataN[218]), .DI25(ofifoDataN[217]), .DI24(ofifoDataN[216]), .DI23(ofifoDataN[215]), .DI22(ofifoDataN[214]), .DI21(ofifoDataN[213]), .DI20(ofifoDataN[212]), .DI19(ofifoDataN[211]),
 .DI18(ofifoDataN[210]), .DI17(ofifoDataN[209]), .DI16(ofifoDataN[208]), .DI15(ofifoDataN[207]), .DI14(ofifoDataN[206]), .DI13(ofifoDataN[205]), .DI12(ofifoDataN[204]), .DI11(ofifoDataN[203]),
 .DI10(ofifoDataN[202]), .DI9(ofifoDataN[201]), .DI8(ofifoDataN[200]), .DI7(ofifoDataN[199]), .DI6(ofifoDataN[198]), .DI5(ofifoDataN[197]), .DI4(ofifoDataN[196]), .DI3(ofifoDataN[195]),
 .DI2(ofifoDataN[194]), .DI1(ofifoDataN[193]), .DI0(ofifoDataN[192]), .WE(n3318), .SYNC_IN(n4792), .SYNC_OUT(n4793));
MPW128KX64 U6038 ( .A16(ofifoAddr4N[16]), .A15(ofifoAddr4N[15]), .A14(ofifoAddr4N[14]), .A13(ofifoAddr4N[13]), .A12(ofifoAddr4N[12]), .A11(ofifoAddr4N[11]),
 .A10(ofifoAddr4N[10]), .A9(ofifoAddr4N[9]), .A8(ofifoAddr4N[8]), .A7(ofifoAddr4N[7]), .A6(ofifoAddr4N[6]), .A5(ofifoAddr4N[5]), .A4(ofifoAddr4N[4]), .A3(ofifoAddr4N[3]),
 .A2(ofifoAddr4N[2]), .A1(ofifoAddr0N[1]), .A0(ofifoAddr0N[0]), .DI63(ofifoDataN[319]), .DI62(ofifoDataN[318]), .DI61(ofifoDataN[317]), .DI60(ofifoDataN[316]), .DI59(ofifoDataN[315]),
 .DI58(ofifoDataN[314]), .DI57(ofifoDataN[313]), .DI56(ofifoDataN[312]), .DI55(ofifoDataN[311]), .DI54(ofifoDataN[310]), .DI53(ofifoDataN[309]), .DI52(ofifoDataN[308]), .DI51(ofifoDataN[307]),
 .DI50(ofifoDataN[306]), .DI49(ofifoDataN[305]), .DI48(ofifoDataN[304]), .DI47(ofifoDataN[303]), .DI46(ofifoDataN[302]), .DI45(ofifoDataN[301]), .DI44(ofifoDataN[300]), .DI43(ofifoDataN[299]),
 .DI42(ofifoDataN[298]), .DI41(ofifoDataN[297]), .DI40(ofifoDataN[296]), .DI39(ofifoDataN[295]), .DI38(ofifoDataN[294]), .DI37(ofifoDataN[293]), .DI36(ofifoDataN[292]), .DI35(ofifoDataN[291]),
 .DI34(ofifoDataN[290]), .DI33(ofifoDataN[289]), .DI32(ofifoDataN[288]), .DI31(ofifoDataN[287]), .DI30(ofifoDataN[286]), .DI29(ofifoDataN[285]), .DI28(ofifoDataN[284]), .DI27(ofifoDataN[283]),
 .DI26(ofifoDataN[282]), .DI25(ofifoDataN[281]), .DI24(ofifoDataN[280]), .DI23(ofifoDataN[279]), .DI22(ofifoDataN[278]), .DI21(ofifoDataN[277]), .DI20(ofifoDataN[276]), .DI19(ofifoDataN[275]),
 .DI18(ofifoDataN[274]), .DI17(ofifoDataN[273]), .DI16(ofifoDataN[272]), .DI15(ofifoDataN[271]), .DI14(ofifoDataN[270]), .DI13(ofifoDataN[269]), .DI12(ofifoDataN[268]), .DI11(ofifoDataN[267]),
 .DI10(ofifoDataN[266]), .DI9(ofifoDataN[265]), .DI8(ofifoDataN[264]), .DI7(ofifoDataN[263]), .DI6(ofifoDataN[262]), .DI5(ofifoDataN[261]), .DI4(ofifoDataN[260]), .DI3(ofifoDataN[259]),
 .DI2(ofifoDataN[258]), .DI1(ofifoDataN[257]), .DI0(ofifoDataN[256]), .WE(n3318), .SYNC_IN(n4793), .SYNC_OUT(n4794));
MPW128KX64 U6039 ( .A16(ofifoAddr5N[16]), .A15(ofifoAddr5N[15]), .A14(ofifoAddr5N[14]), .A13(ofifoAddr5N[13]), .A12(ofifoAddr5N[12]), .A11(ofifoAddr5N[11]),
 .A10(ofifoAddr5N[10]), .A9(ofifoAddr5N[9]), .A8(ofifoAddr5N[8]), .A7(ofifoAddr5N[7]), .A6(ofifoAddr5N[6]), .A5(ofifoAddr5N[5]), .A4(ofifoAddr5N[4]), .A3(ofifoAddr5N[3]),
 .A2(ofifoAddr5N[2]), .A1(ofifoAddr1N[1]), .A0(ofifoAddr7N[0]), .DI63(ofifoDataN[383]), .DI62(ofifoDataN[382]), .DI61(ofifoDataN[381]), .DI60(ofifoDataN[380]), .DI59(ofifoDataN[379]),
 .DI58(ofifoDataN[378]), .DI57(ofifoDataN[377]), .DI56(ofifoDataN[376]), .DI55(ofifoDataN[375]), .DI54(ofifoDataN[374]), .DI53(ofifoDataN[373]), .DI52(ofifoDataN[372]), .DI51(ofifoDataN[371]),
 .DI50(ofifoDataN[370]), .DI49(ofifoDataN[369]), .DI48(ofifoDataN[368]), .DI47(ofifoDataN[367]), .DI46(ofifoDataN[366]), .DI45(ofifoDataN[365]), .DI44(ofifoDataN[364]), .DI43(ofifoDataN[363]),
 .DI42(ofifoDataN[362]), .DI41(ofifoDataN[361]), .DI40(ofifoDataN[360]), .DI39(ofifoDataN[359]), .DI38(ofifoDataN[358]), .DI37(ofifoDataN[357]), .DI36(ofifoDataN[356]), .DI35(ofifoDataN[355]),
 .DI34(ofifoDataN[354]), .DI33(ofifoDataN[353]), .DI32(ofifoDataN[352]), .DI31(ofifoDataN[351]), .DI30(ofifoDataN[350]), .DI29(ofifoDataN[349]), .DI28(ofifoDataN[348]), .DI27(ofifoDataN[347]),
 .DI26(ofifoDataN[346]), .DI25(ofifoDataN[345]), .DI24(ofifoDataN[344]), .DI23(ofifoDataN[343]), .DI22(ofifoDataN[342]), .DI21(ofifoDataN[341]), .DI20(ofifoDataN[340]), .DI19(ofifoDataN[339]),
 .DI18(ofifoDataN[338]), .DI17(ofifoDataN[337]), .DI16(ofifoDataN[336]), .DI15(ofifoDataN[335]), .DI14(ofifoDataN[334]), .DI13(ofifoDataN[333]), .DI12(ofifoDataN[332]), .DI11(ofifoDataN[331]),
 .DI10(ofifoDataN[330]), .DI9(ofifoDataN[329]), .DI8(ofifoDataN[328]), .DI7(ofifoDataN[327]), .DI6(ofifoDataN[326]), .DI5(ofifoDataN[325]), .DI4(ofifoDataN[324]), .DI3(ofifoDataN[323]),
 .DI2(ofifoDataN[322]), .DI1(ofifoDataN[321]), .DI0(ofifoDataN[320]), .WE(n3318), .SYNC_IN(n4794), .SYNC_OUT(n4795));
MPW128KX64 U6040 ( .A16(ofifoAddr6N[16]), .A15(ofifoAddr6N[15]), .A14(ofifoAddr6N[14]), .A13(ofifoAddr6N[13]), .A12(ofifoAddr6N[12]), .A11(ofifoAddr6N[11]),
 .A10(ofifoAddr6N[10]), .A9(ofifoAddr6N[9]), .A8(ofifoAddr6N[8]), .A7(ofifoAddr6N[7]), .A6(ofifoAddr6N[6]), .A5(ofifoAddr6N[5]), .A4(ofifoAddr6N[4]), .A3(ofifoAddr6N[3]),
 .A2(ofifoAddr6N[2]), .A1(ofifoAddr6N[1]), .A0(ofifoAddr0N[0]), .DI63(ofifoDataN[447]), .DI62(ofifoDataN[446]), .DI61(ofifoDataN[445]), .DI60(ofifoDataN[444]), .DI59(ofifoDataN[443]),
 .DI58(ofifoDataN[442]), .DI57(ofifoDataN[441]), .DI56(ofifoDataN[440]), .DI55(ofifoDataN[439]), .DI54(ofifoDataN[438]), .DI53(ofifoDataN[437]), .DI52(ofifoDataN[436]), .DI51(ofifoDataN[435]),
 .DI50(ofifoDataN[434]), .DI49(ofifoDataN[433]), .DI48(ofifoDataN[432]), .DI47(ofifoDataN[431]), .DI46(ofifoDataN[430]), .DI45(ofifoDataN[429]), .DI44(ofifoDataN[428]), .DI43(ofifoDataN[427]),
 .DI42(ofifoDataN[426]), .DI41(ofifoDataN[425]), .DI40(ofifoDataN[424]), .DI39(ofifoDataN[423]), .DI38(ofifoDataN[422]), .DI37(ofifoDataN[421]), .DI36(ofifoDataN[420]), .DI35(ofifoDataN[419]),
 .DI34(ofifoDataN[418]), .DI33(ofifoDataN[417]), .DI32(ofifoDataN[416]), .DI31(ofifoDataN[415]), .DI30(ofifoDataN[414]), .DI29(ofifoDataN[413]), .DI28(ofifoDataN[412]), .DI27(ofifoDataN[411]),
 .DI26(ofifoDataN[410]), .DI25(ofifoDataN[409]), .DI24(ofifoDataN[408]), .DI23(ofifoDataN[407]), .DI22(ofifoDataN[406]), .DI21(ofifoDataN[405]), .DI20(ofifoDataN[404]), .DI19(ofifoDataN[403]),
 .DI18(ofifoDataN[402]), .DI17(ofifoDataN[401]), .DI16(ofifoDataN[400]), .DI15(ofifoDataN[399]), .DI14(ofifoDataN[398]), .DI13(ofifoDataN[397]), .DI12(ofifoDataN[396]), .DI11(ofifoDataN[395]),
 .DI10(ofifoDataN[394]), .DI9(ofifoDataN[393]), .DI8(ofifoDataN[392]), .DI7(ofifoDataN[391]), .DI6(ofifoDataN[390]), .DI5(ofifoDataN[389]), .DI4(ofifoDataN[388]), .DI3(ofifoDataN[387]),
 .DI2(ofifoDataN[386]), .DI1(ofifoDataN[385]), .DI0(ofifoDataN[384]), .WE(n3318), .SYNC_IN(n4795), .SYNC_OUT(n4796));
MPW128KX64 U6041 ( .A16(ofifoAddr7N[16]), .A15(ofifoAddr7N[15]), .A14(ofifoAddr7N[14]), .A13(ofifoAddr7N[13]), .A12(ofifoAddr7N[12]), .A11(ofifoAddr7N[11]),
 .A10(ofifoAddr7N[10]), .A9(ofifoAddr7N[9]), .A8(ofifoAddr7N[8]), .A7(ofifoAddr7N[7]), .A6(ofifoAddr7N[6]), .A5(ofifoAddr7N[5]), .A4(ofifoAddr7N[4]), .A3(ofifoAddr7N[3]),
 .A2(ofifoAddr7N[2]), .A1(ofifoAddr7N[1]), .A0(ofifoAddr7N[0]), .DI63(ofifoDataN[511]), .DI62(ofifoDataN[510]), .DI61(ofifoDataN[509]), .DI60(ofifoDataN[508]), .DI59(ofifoDataN[507]),
 .DI58(ofifoDataN[506]), .DI57(ofifoDataN[505]), .DI56(ofifoDataN[504]), .DI55(ofifoDataN[503]), .DI54(ofifoDataN[502]), .DI53(ofifoDataN[501]), .DI52(ofifoDataN[500]), .DI51(ofifoDataN[499]),
 .DI50(ofifoDataN[498]), .DI49(ofifoDataN[497]), .DI48(ofifoDataN[496]), .DI47(ofifoDataN[495]), .DI46(ofifoDataN[494]), .DI45(ofifoDataN[493]), .DI44(ofifoDataN[492]), .DI43(ofifoDataN[491]),
 .DI42(ofifoDataN[490]), .DI41(ofifoDataN[489]), .DI40(ofifoDataN[488]), .DI39(ofifoDataN[487]), .DI38(ofifoDataN[486]), .DI37(ofifoDataN[485]), .DI36(ofifoDataN[484]), .DI35(ofifoDataN[483]),
 .DI34(ofifoDataN[482]), .DI33(ofifoDataN[481]), .DI32(ofifoDataN[480]), .DI31(ofifoDataN[479]), .DI30(ofifoDataN[478]), .DI29(ofifoDataN[477]), .DI28(ofifoDataN[476]), .DI27(ofifoDataN[475]),
 .DI26(ofifoDataN[474]), .DI25(ofifoDataN[473]), .DI24(ofifoDataN[472]), .DI23(ofifoDataN[471]), .DI22(ofifoDataN[470]), .DI21(ofifoDataN[469]), .DI20(ofifoDataN[468]), .DI19(ofifoDataN[467]),
 .DI18(ofifoDataN[466]), .DI17(ofifoDataN[465]), .DI16(ofifoDataN[464]), .DI15(ofifoDataN[463]), .DI14(ofifoDataN[462]), .DI13(ofifoDataN[461]), .DI12(ofifoDataN[460]), .DI11(ofifoDataN[459]),
 .DI10(ofifoDataN[458]), .DI9(ofifoDataN[457]), .DI8(ofifoDataN[456]), .DI7(ofifoDataN[455]), .DI6(ofifoDataN[454]), .DI5(ofifoDataN[453]), .DI4(ofifoDataN[452]), .DI3(ofifoDataN[451]),
 .DI2(ofifoDataN[450]), .DI1(ofifoDataN[449]), .DI0(ofifoDataN[448]), .WE(n3318), .SYNC_IN(n4796), .SYNC_OUT(n4797));
MPW128KX64 U6042 ( .A16(ofifoAddr8N[16]), .A15(ofifoAddr8N[15]), .A14(ofifoAddr8N[14]), .A13(ofifoAddr8N[13]), .A12(ofifoAddr8N[12]), .A11(ofifoAddr8N[11]),
 .A10(ofifoAddr8N[10]), .A9(ofifoAddr8N[9]), .A8(ofifoAddr8N[8]), .A7(ofifoAddr8N[7]), .A6(ofifoAddr8N[6]), .A5(ofifoAddr8N[5]), .A4(ofifoAddr8N[4]), .A3(ofifoAddr8N[3]),
 .A2(ofifoAddr0N[2]), .A1(ofifoAddr0N[1]), .A0(ofifoAddr0N[0]), .DI63(ofifoDataN[575]), .DI62(ofifoDataN[574]), .DI61(ofifoDataN[573]), .DI60(ofifoDataN[572]), .DI59(ofifoDataN[571]),
 .DI58(ofifoDataN[570]), .DI57(ofifoDataN[569]), .DI56(ofifoDataN[568]), .DI55(ofifoDataN[567]), .DI54(ofifoDataN[566]), .DI53(ofifoDataN[565]), .DI52(ofifoDataN[564]), .DI51(ofifoDataN[563]),
 .DI50(ofifoDataN[562]), .DI49(ofifoDataN[561]), .DI48(ofifoDataN[560]), .DI47(ofifoDataN[559]), .DI46(ofifoDataN[558]), .DI45(ofifoDataN[557]), .DI44(ofifoDataN[556]), .DI43(ofifoDataN[555]),
 .DI42(ofifoDataN[554]), .DI41(ofifoDataN[553]), .DI40(ofifoDataN[552]), .DI39(ofifoDataN[551]), .DI38(ofifoDataN[550]), .DI37(ofifoDataN[549]), .DI36(ofifoDataN[548]), .DI35(ofifoDataN[547]),
 .DI34(ofifoDataN[546]), .DI33(ofifoDataN[545]), .DI32(ofifoDataN[544]), .DI31(ofifoDataN[543]), .DI30(ofifoDataN[542]), .DI29(ofifoDataN[541]), .DI28(ofifoDataN[540]), .DI27(ofifoDataN[539]),
 .DI26(ofifoDataN[538]), .DI25(ofifoDataN[537]), .DI24(ofifoDataN[536]), .DI23(ofifoDataN[535]), .DI22(ofifoDataN[534]), .DI21(ofifoDataN[533]), .DI20(ofifoDataN[532]), .DI19(ofifoDataN[531]),
 .DI18(ofifoDataN[530]), .DI17(ofifoDataN[529]), .DI16(ofifoDataN[528]), .DI15(ofifoDataN[527]), .DI14(ofifoDataN[526]), .DI13(ofifoDataN[525]), .DI12(ofifoDataN[524]), .DI11(ofifoDataN[523]),
 .DI10(ofifoDataN[522]), .DI9(ofifoDataN[521]), .DI8(ofifoDataN[520]), .DI7(ofifoDataN[519]), .DI6(ofifoDataN[518]), .DI5(ofifoDataN[517]), .DI4(ofifoDataN[516]), .DI3(ofifoDataN[515]),
 .DI2(ofifoDataN[514]), .DI1(ofifoDataN[513]), .DI0(ofifoDataN[512]), .WE(n3318), .SYNC_IN(n4797), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "ixc_gfm_ofifo 1 63 0 0 131071"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m2 "ixc_gfm_ctl 1 63 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "2"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
`ifdef CBV
`else
`ifdef MPW2X64_MPR2X64
`else
module MPW2X64( A0, DI63, DI62, DI61, DI60, DI59, DI58,
 DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42,
 DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34,
 DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26,
 DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18,
 DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2,
 DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A0, DI63, DI62, DI61, DI60, DI59, DI58, DI57,
 DI56, DI55, DI54, DI53, DI52, DI51, DI50, DI49, DI48, DI47,
 DI46, DI45, DI44, DI43, DI42, DI41, DI40, DI39, DI38, DI37,
 DI36, DI35, DI34, DI33, DI32, DI31, DI30, DI29, DI28, DI27,
 DI26, DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18, DI17,
 DI16, DI15, DI14, DI13, DI12, DI11, DI10, DI9, DI8, DI7,
 DI6, DI5, DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR2X64_
`else
module MPR2X64( A0, SYNC_IN, DO63, DO62, DO61, DO60, DO59,
 DO58, DO57, DO56, DO55, DO54, DO53, DO52, DO51,
 DO50, DO49, DO48, DO47, DO46, DO45, DO44, DO43,
 DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35,
 DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27,
 DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19,
 DO18, DO17, DO16, DO15, DO14, DO13, DO12, DO11,
 DO10, DO9, DO8, DO7, DO6, DO5, DO4, DO3,
 DO2, DO1, DO0, SYNC_OUT);
input  A0, SYNC_IN;
output  DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56,
 DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26,
 DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16,
 DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR2X64_
`endif
`define MPW2X64_MPR2X64
`endif
`ifdef MPW128KX64_MPR128KX64
`else
module MPW128KX64( A16, A15, A14, A13, A12, A11, A10,
 A9, A8, A7, A6, A5, A4, A3, A2,
 A1, A0, DI63, DI62, DI61, DI60, DI59, DI58,
 DI57, DI56, DI55, DI54, DI53, DI52, DI51, DI50,
 DI49, DI48, DI47, DI46, DI45, DI44, DI43, DI42,
 DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34,
 DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26,
 DI25, DI24, DI23, DI22, DI21, DI20, DI19, DI18,
 DI17, DI16, DI15, DI14, DI13, DI12, DI11, DI10,
 DI9, DI8, DI7, DI6, DI5, DI4, DI3, DI2,
 DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A16, A15, A14, A13, A12, A11, A10, A9,
 A8, A7, A6, A5, A4, A3, A2, A1, A0, DI63,
 DI62, DI61, DI60, DI59, DI58, DI57, DI56, DI55, DI54, DI53,
 DI52, DI51, DI50, DI49, DI48, DI47, DI46, DI45, DI44, DI43,
 DI42, DI41, DI40, DI39, DI38, DI37, DI36, DI35, DI34, DI33,
 DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24, DI23,
 DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5, DI4, DI3,
 DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR128KX64_
`else
module MPR128KX64( A16, A15, A14, A13, A12, A11, A10,
 A9, A8, A7, A6, A5, A4, A3, A2,
 A1, A0, SYNC_IN, DO63, DO62, DO61, DO60, DO59,
 DO58, DO57, DO56, DO55, DO54, DO53, DO52, DO51,
 DO50, DO49, DO48, DO47, DO46, DO45, DO44, DO43,
 DO42, DO41, DO40, DO39, DO38, DO37, DO36, DO35,
 DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27,
 DO26, DO25, DO24, DO23, DO22, DO21, DO20, DO19,
 DO18, DO17, DO16, DO15, DO14, DO13, DO12, DO11,
 DO10, DO9, DO8, DO7, DO6, DO5, DO4, DO3,
 DO2, DO1, DO0, SYNC_OUT);
input  A16, A15, A14, A13, A12, A11, A10, A9,
 A8, A7, A6, A5, A4, A3, A2, A1, A0, SYNC_IN;
output  DO63, DO62, DO61, DO60, DO59, DO58, DO57, DO56,
 DO55, DO54, DO53, DO52, DO51, DO50, DO49, DO48, DO47, DO46,
 DO45, DO44, DO43, DO42, DO41, DO40, DO39, DO38, DO37, DO36,
 DO35, DO34, DO33, DO32, DO31, DO30, DO29, DO28, DO27, DO26,
 DO25, DO24, DO23, DO22, DO21, DO20, DO19, DO18, DO17, DO16,
 DO15, DO14, DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT;
endmodule
`define _MPR128KX64_
`endif
`define MPW128KX64_MPR128KX64
`endif
`endif
