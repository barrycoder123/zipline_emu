
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_regs ( clk, i_reset_, i_sw_init, i_addr, i_wr_strb, i_wr_data, 
	i_rd_strb, o_rd_data, o_ack, o_err_ack, o_spare_config, 
	o_cceip0_out_ia_wdata_part0, o_cceip0_out_ia_wdata_part1, 
	o_cceip0_out_ia_wdata_part2, o_cceip0_out_ia_config, 
	o_cceip0_out_im_config, o_cceip0_out_im_read_done, 
	o_cceip1_out_ia_wdata_part0, o_cceip1_out_ia_wdata_part1, 
	o_cceip1_out_ia_wdata_part2, o_cceip1_out_ia_config, 
	o_cceip1_out_im_config, o_cceip1_out_im_read_done, 
	o_cceip2_out_ia_wdata_part0, o_cceip2_out_ia_wdata_part1, 
	o_cceip2_out_ia_wdata_part2, o_cceip2_out_ia_config, 
	o_cceip2_out_im_config, o_cceip2_out_im_read_done, 
	o_cceip3_out_ia_wdata_part0, o_cceip3_out_ia_wdata_part1, 
	o_cceip3_out_ia_wdata_part2, o_cceip3_out_ia_config, 
	o_cceip3_out_im_config, o_cceip3_out_im_read_done, 
	o_cddip0_out_ia_wdata_part0, o_cddip0_out_ia_wdata_part1, 
	o_cddip0_out_ia_wdata_part2, o_cddip0_out_ia_config, 
	o_cddip0_out_im_config, o_cddip0_out_im_read_done, 
	o_cddip1_out_ia_wdata_part0, o_cddip1_out_ia_wdata_part1, 
	o_cddip1_out_ia_wdata_part2, o_cddip1_out_ia_config, 
	o_cddip1_out_im_config, o_cddip1_out_im_read_done, 
	o_cddip2_out_ia_wdata_part0, o_cddip2_out_ia_wdata_part1, 
	o_cddip2_out_ia_wdata_part2, o_cddip2_out_ia_config, 
	o_cddip2_out_im_config, o_cddip2_out_im_read_done, 
	o_cddip3_out_ia_wdata_part0, o_cddip3_out_ia_wdata_part1, 
	o_cddip3_out_ia_wdata_part2, o_cddip3_out_ia_config, 
	o_cddip3_out_im_config, o_cddip3_out_im_read_done, 
	o_ckv_ia_wdata_part0, o_ckv_ia_wdata_part1, o_ckv_ia_config, 
	o_kim_ia_wdata_part0, o_kim_ia_wdata_part1, o_kim_ia_config, 
	o_label0_config, o_label0_data7, o_label0_data6, o_label0_data5, 
	o_label0_data4, o_label0_data3, o_label0_data2, o_label0_data1, 
	o_label0_data0, o_label1_config, o_label1_data7, o_label1_data6, 
	o_label1_data5, o_label1_data4, o_label1_data3, o_label1_data2, 
	o_label1_data1, o_label1_data0, o_label2_config, o_label2_data7, 
	o_label2_data6, o_label2_data5, o_label2_data4, o_label2_data3, 
	o_label2_data2, o_label2_data1, o_label2_data0, o_label3_config, 
	o_label3_data7, o_label3_data6, o_label3_data5, o_label3_data4, 
	o_label3_data3, o_label3_data2, o_label3_data1, o_label3_data0, 
	o_label4_config, o_label4_data7, o_label4_data6, o_label4_data5, 
	o_label4_data4, o_label4_data3, o_label4_data2, o_label4_data1, 
	o_label4_data0, o_label5_config, o_label5_data7, o_label5_data6, 
	o_label5_data5, o_label5_data4, o_label5_data3, o_label5_data2, 
	o_label5_data1, o_label5_data0, o_label6_config, o_label6_data7, 
	o_label6_data6, o_label6_data5, o_label6_data4, o_label6_data3, 
	o_label6_data2, o_label6_data1, o_label6_data0, o_label7_config, 
	o_label7_data7, o_label7_data6, o_label7_data5, o_label7_data4, 
	o_label7_data3, o_label7_data2, o_label7_data1, o_label7_data0, 
	o_kdf_drbg_ctrl, o_kdf_drbg_seed_0_state_key_31_0, 
	o_kdf_drbg_seed_0_state_key_63_32, o_kdf_drbg_seed_0_state_key_95_64, 
	o_kdf_drbg_seed_0_state_key_127_96, 
	o_kdf_drbg_seed_0_state_key_159_128, 
	o_kdf_drbg_seed_0_state_key_191_160, 
	o_kdf_drbg_seed_0_state_key_223_192, 
	o_kdf_drbg_seed_0_state_key_255_224, 
	o_kdf_drbg_seed_0_state_value_31_0, 
	o_kdf_drbg_seed_0_state_value_63_32, 
	o_kdf_drbg_seed_0_state_value_95_64, 
	o_kdf_drbg_seed_0_state_value_127_96, 
	o_kdf_drbg_seed_0_reseed_interval_0, 
	o_kdf_drbg_seed_0_reseed_interval_1, 
	o_kdf_drbg_seed_1_state_key_31_0, o_kdf_drbg_seed_1_state_key_63_32, 
	o_kdf_drbg_seed_1_state_key_95_64, 
	o_kdf_drbg_seed_1_state_key_127_96, 
	o_kdf_drbg_seed_1_state_key_159_128, 
	o_kdf_drbg_seed_1_state_key_191_160, 
	o_kdf_drbg_seed_1_state_key_223_192, 
	o_kdf_drbg_seed_1_state_key_255_224, 
	o_kdf_drbg_seed_1_state_value_31_0, 
	o_kdf_drbg_seed_1_state_value_63_32, 
	o_kdf_drbg_seed_1_state_value_95_64, 
	o_kdf_drbg_seed_1_state_value_127_96, 
	o_kdf_drbg_seed_1_reseed_interval_0, 
	o_kdf_drbg_seed_1_reseed_interval_1, o_interrupt_status, 
	o_interrupt_mask, o_engine_sticky_status, o_bimc_monitor_mask, 
	o_bimc_ecc_uncorrectable_error_cnt, o_bimc_ecc_correctable_error_cnt, 
	o_bimc_parity_error_cnt, o_bimc_global_config, o_bimc_eccpar_debug, 
	o_bimc_cmd2, o_bimc_cmd1, o_bimc_cmd0, o_bimc_rxcmd2, o_bimc_rxrsp2, 
	o_bimc_pollrsp2, o_bimc_dbgcmd2, o_im_consumed, o_tready_override, 
	o_regs_sa_ctrl, o_sa_snapshot_ia_wdata_part0, 
	o_sa_snapshot_ia_wdata_part1, o_sa_snapshot_ia_config, 
	o_sa_count_ia_wdata_part0, o_sa_count_ia_wdata_part1, 
	o_sa_count_ia_config, o_cceip_encrypt_kop_fifo_override, 
	o_cceip_validate_kop_fifo_override, 
	o_cddip_decrypt_kop_fifo_override, o_sa_global_ctrl, 
	o_sa_ctrl_ia_wdata_part0, o_sa_ctrl_ia_config, 
	o_kdf_test_key_size_config, i_blkid_revid_config, i_revision_config, 
	i_spare_config, i_cceip0_out_ia_capability, i_cceip0_out_ia_status, 
	i_cceip0_out_ia_rdata_part0, i_cceip0_out_ia_rdata_part1, 
	i_cceip0_out_ia_rdata_part2, i_cceip0_out_im_status, 
	i_cceip0_out_im_read_done, i_cceip1_out_ia_capability, 
	i_cceip1_out_ia_status, i_cceip1_out_ia_rdata_part0, 
	i_cceip1_out_ia_rdata_part1, i_cceip1_out_ia_rdata_part2, 
	i_cceip1_out_im_status, i_cceip1_out_im_read_done, 
	i_cceip2_out_ia_capability, i_cceip2_out_ia_status, 
	i_cceip2_out_ia_rdata_part0, i_cceip2_out_ia_rdata_part1, 
	i_cceip2_out_ia_rdata_part2, i_cceip2_out_im_status, 
	i_cceip2_out_im_read_done, i_cceip3_out_ia_capability, 
	i_cceip3_out_ia_status, i_cceip3_out_ia_rdata_part0, 
	i_cceip3_out_ia_rdata_part1, i_cceip3_out_ia_rdata_part2, 
	i_cceip3_out_im_status, i_cceip3_out_im_read_done, 
	i_cddip0_out_ia_capability, i_cddip0_out_ia_status, 
	i_cddip0_out_ia_rdata_part0, i_cddip0_out_ia_rdata_part1, 
	i_cddip0_out_ia_rdata_part2, i_cddip0_out_im_status, 
	i_cddip0_out_im_read_done, i_cddip1_out_ia_capability, 
	i_cddip1_out_ia_status, i_cddip1_out_ia_rdata_part0, 
	i_cddip1_out_ia_rdata_part1, i_cddip1_out_ia_rdata_part2, 
	i_cddip1_out_im_status, i_cddip1_out_im_read_done, 
	i_cddip2_out_ia_capability, i_cddip2_out_ia_status, 
	i_cddip2_out_ia_rdata_part0, i_cddip2_out_ia_rdata_part1, 
	i_cddip2_out_ia_rdata_part2, i_cddip2_out_im_status, 
	i_cddip2_out_im_read_done, i_cddip3_out_ia_capability, 
	i_cddip3_out_ia_status, i_cddip3_out_ia_rdata_part0, 
	i_cddip3_out_ia_rdata_part1, i_cddip3_out_ia_rdata_part2, 
	i_cddip3_out_im_status, i_cddip3_out_im_read_done, 
	i_ckv_ia_capability, i_ckv_ia_status, i_ckv_ia_rdata_part0, 
	i_ckv_ia_rdata_part1, i_kim_ia_capability, i_kim_ia_status, 
	i_kim_ia_rdata_part0, i_kim_ia_rdata_part1, i_kdf_drbg_ctrl, 
	i_interrupt_status, i_engine_sticky_status, i_bimc_monitor, 
	i_bimc_ecc_uncorrectable_error_cnt, i_bimc_ecc_correctable_error_cnt, 
	i_bimc_parity_error_cnt, i_bimc_global_config, i_bimc_memid, 
	i_bimc_eccpar_debug, i_bimc_cmd2, i_bimc_rxcmd2, i_bimc_rxcmd1, 
	i_bimc_rxcmd0, i_bimc_rxrsp2, i_bimc_rxrsp1, i_bimc_rxrsp0, 
	i_bimc_pollrsp2, i_bimc_pollrsp1, i_bimc_pollrsp0, i_bimc_dbgcmd2, 
	i_bimc_dbgcmd1, i_bimc_dbgcmd0, i_im_available, i_im_consumed, 
	i_tready_override, i_regs_sa_ctrl, i_sa_snapshot_ia_capability, 
	i_sa_snapshot_ia_status, i_sa_snapshot_ia_rdata_part0, 
	i_sa_snapshot_ia_rdata_part1, i_sa_count_ia_capability, 
	i_sa_count_ia_status, i_sa_count_ia_rdata_part0, 
	i_sa_count_ia_rdata_part1, i_idle_components, i_sa_global_ctrl, 
	i_sa_ctrl_ia_capability, i_sa_ctrl_ia_status, 
	i_sa_ctrl_ia_rdata_part0, o_reg_written, o_reg_read, o_reg_wr_data, 
	o_reg_addr);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input i_reset_;
input i_sw_init;
input [10:0] i_addr;
input i_wr_strb;
input [31:0] i_wr_data;
input i_rd_strb;
output [31:0] o_rd_data;
output o_ack;
output o_err_ack;
output [31:0] o_spare_config;
output [31:0] o_cceip0_out_ia_wdata_part0;
output [31:0] o_cceip0_out_ia_wdata_part1;
output [31:0] o_cceip0_out_ia_wdata_part2;
output [12:0] o_cceip0_out_ia_config;
output [11:0] o_cceip0_out_im_config;
output [1:0] o_cceip0_out_im_read_done;
output [31:0] o_cceip1_out_ia_wdata_part0;
output [31:0] o_cceip1_out_ia_wdata_part1;
output [31:0] o_cceip1_out_ia_wdata_part2;
output [12:0] o_cceip1_out_ia_config;
output [11:0] o_cceip1_out_im_config;
output [1:0] o_cceip1_out_im_read_done;
output [31:0] o_cceip2_out_ia_wdata_part0;
output [31:0] o_cceip2_out_ia_wdata_part1;
output [31:0] o_cceip2_out_ia_wdata_part2;
output [12:0] o_cceip2_out_ia_config;
output [11:0] o_cceip2_out_im_config;
output [1:0] o_cceip2_out_im_read_done;
output [31:0] o_cceip3_out_ia_wdata_part0;
output [31:0] o_cceip3_out_ia_wdata_part1;
output [31:0] o_cceip3_out_ia_wdata_part2;
output [12:0] o_cceip3_out_ia_config;
output [11:0] o_cceip3_out_im_config;
output [1:0] o_cceip3_out_im_read_done;
output [31:0] o_cddip0_out_ia_wdata_part0;
output [31:0] o_cddip0_out_ia_wdata_part1;
output [31:0] o_cddip0_out_ia_wdata_part2;
output [12:0] o_cddip0_out_ia_config;
output [11:0] o_cddip0_out_im_config;
output [1:0] o_cddip0_out_im_read_done;
output [31:0] o_cddip1_out_ia_wdata_part0;
output [31:0] o_cddip1_out_ia_wdata_part1;
output [31:0] o_cddip1_out_ia_wdata_part2;
output [12:0] o_cddip1_out_ia_config;
output [11:0] o_cddip1_out_im_config;
output [1:0] o_cddip1_out_im_read_done;
output [31:0] o_cddip2_out_ia_wdata_part0;
output [31:0] o_cddip2_out_ia_wdata_part1;
output [31:0] o_cddip2_out_ia_wdata_part2;
output [12:0] o_cddip2_out_ia_config;
output [11:0] o_cddip2_out_im_config;
output [1:0] o_cddip2_out_im_read_done;
output [31:0] o_cddip3_out_ia_wdata_part0;
output [31:0] o_cddip3_out_ia_wdata_part1;
output [31:0] o_cddip3_out_ia_wdata_part2;
output [12:0] o_cddip3_out_ia_config;
output [11:0] o_cddip3_out_im_config;
output [1:0] o_cddip3_out_im_read_done;
output [31:0] o_ckv_ia_wdata_part0;
output [31:0] o_ckv_ia_wdata_part1;
output [18:0] o_ckv_ia_config;
output [20:0] o_kim_ia_wdata_part0;
output [16:0] o_kim_ia_wdata_part1;
output [17:0] o_kim_ia_config;
output [15:0] o_label0_config;
output [31:0] o_label0_data7;
output [31:0] o_label0_data6;
output [31:0] o_label0_data5;
output [31:0] o_label0_data4;
output [31:0] o_label0_data3;
output [31:0] o_label0_data2;
output [31:0] o_label0_data1;
output [31:0] o_label0_data0;
output [15:0] o_label1_config;
output [31:0] o_label1_data7;
output [31:0] o_label1_data6;
output [31:0] o_label1_data5;
output [31:0] o_label1_data4;
output [31:0] o_label1_data3;
output [31:0] o_label1_data2;
output [31:0] o_label1_data1;
output [31:0] o_label1_data0;
output [15:0] o_label2_config;
output [31:0] o_label2_data7;
output [31:0] o_label2_data6;
output [31:0] o_label2_data5;
output [31:0] o_label2_data4;
output [31:0] o_label2_data3;
output [31:0] o_label2_data2;
output [31:0] o_label2_data1;
output [31:0] o_label2_data0;
output [15:0] o_label3_config;
output [31:0] o_label3_data7;
output [31:0] o_label3_data6;
output [31:0] o_label3_data5;
output [31:0] o_label3_data4;
output [31:0] o_label3_data3;
output [31:0] o_label3_data2;
output [31:0] o_label3_data1;
output [31:0] o_label3_data0;
output [15:0] o_label4_config;
output [31:0] o_label4_data7;
output [31:0] o_label4_data6;
output [31:0] o_label4_data5;
output [31:0] o_label4_data4;
output [31:0] o_label4_data3;
output [31:0] o_label4_data2;
output [31:0] o_label4_data1;
output [31:0] o_label4_data0;
output [15:0] o_label5_config;
output [31:0] o_label5_data7;
output [31:0] o_label5_data6;
output [31:0] o_label5_data5;
output [31:0] o_label5_data4;
output [31:0] o_label5_data3;
output [31:0] o_label5_data2;
output [31:0] o_label5_data1;
output [31:0] o_label5_data0;
output [15:0] o_label6_config;
output [31:0] o_label6_data7;
output [31:0] o_label6_data6;
output [31:0] o_label6_data5;
output [31:0] o_label6_data4;
output [31:0] o_label6_data3;
output [31:0] o_label6_data2;
output [31:0] o_label6_data1;
output [31:0] o_label6_data0;
output [15:0] o_label7_config;
output [31:0] o_label7_data7;
output [31:0] o_label7_data6;
output [31:0] o_label7_data5;
output [31:0] o_label7_data4;
output [31:0] o_label7_data3;
output [31:0] o_label7_data2;
output [31:0] o_label7_data1;
output [31:0] o_label7_data0;
output [1:0] o_kdf_drbg_ctrl;
output [31:0] o_kdf_drbg_seed_0_state_key_31_0;
output [31:0] o_kdf_drbg_seed_0_state_key_63_32;
output [31:0] o_kdf_drbg_seed_0_state_key_95_64;
output [31:0] o_kdf_drbg_seed_0_state_key_127_96;
output [31:0] o_kdf_drbg_seed_0_state_key_159_128;
output [31:0] o_kdf_drbg_seed_0_state_key_191_160;
output [31:0] o_kdf_drbg_seed_0_state_key_223_192;
output [31:0] o_kdf_drbg_seed_0_state_key_255_224;
output [31:0] o_kdf_drbg_seed_0_state_value_31_0;
output [31:0] o_kdf_drbg_seed_0_state_value_63_32;
output [31:0] o_kdf_drbg_seed_0_state_value_95_64;
output [31:0] o_kdf_drbg_seed_0_state_value_127_96;
output [31:0] o_kdf_drbg_seed_0_reseed_interval_0;
output [15:0] o_kdf_drbg_seed_0_reseed_interval_1;
output [31:0] o_kdf_drbg_seed_1_state_key_31_0;
output [31:0] o_kdf_drbg_seed_1_state_key_63_32;
output [31:0] o_kdf_drbg_seed_1_state_key_95_64;
output [31:0] o_kdf_drbg_seed_1_state_key_127_96;
output [31:0] o_kdf_drbg_seed_1_state_key_159_128;
output [31:0] o_kdf_drbg_seed_1_state_key_191_160;
output [31:0] o_kdf_drbg_seed_1_state_key_223_192;
output [31:0] o_kdf_drbg_seed_1_state_key_255_224;
output [31:0] o_kdf_drbg_seed_1_state_value_31_0;
output [31:0] o_kdf_drbg_seed_1_state_value_63_32;
output [31:0] o_kdf_drbg_seed_1_state_value_95_64;
output [31:0] o_kdf_drbg_seed_1_state_value_127_96;
output [31:0] o_kdf_drbg_seed_1_reseed_interval_0;
output [15:0] o_kdf_drbg_seed_1_reseed_interval_1;
output [4:0] o_interrupt_status;
output [4:0] o_interrupt_mask;
output [7:0] o_engine_sticky_status;
output [6:0] o_bimc_monitor_mask;
output [31:0] o_bimc_ecc_uncorrectable_error_cnt;
output [31:0] o_bimc_ecc_correctable_error_cnt;
output [31:0] o_bimc_parity_error_cnt;
output [31:0] o_bimc_global_config;
output [28:0] o_bimc_eccpar_debug;
output [10:0] o_bimc_cmd2;
output [31:0] o_bimc_cmd1;
output [31:0] o_bimc_cmd0;
output [9:0] o_bimc_rxcmd2;
output [9:0] o_bimc_rxrsp2;
output [9:0] o_bimc_pollrsp2;
output [9:0] o_bimc_dbgcmd2;
output [15:0] o_im_consumed;
output [8:0] o_tready_override;
output [31:0] o_regs_sa_ctrl;
output [31:0] o_sa_snapshot_ia_wdata_part0;
output [31:0] o_sa_snapshot_ia_wdata_part1;
output [8:0] o_sa_snapshot_ia_config;
output [31:0] o_sa_count_ia_wdata_part0;
output [31:0] o_sa_count_ia_wdata_part1;
output [8:0] o_sa_count_ia_config;
output [6:0] o_cceip_encrypt_kop_fifo_override;
output [6:0] o_cceip_validate_kop_fifo_override;
output [6:0] o_cddip_decrypt_kop_fifo_override;
output [31:0] o_sa_global_ctrl;
output [31:0] o_sa_ctrl_ia_wdata_part0;
output [8:0] o_sa_ctrl_ia_config;
output [31:0] o_kdf_test_key_size_config;
input [31:0] i_blkid_revid_config;
input [7:0] i_revision_config;
input [31:0] i_spare_config;
input [19:0] i_cceip0_out_ia_capability;
input [16:0] i_cceip0_out_ia_status;
input [31:0] i_cceip0_out_ia_rdata_part0;
input [31:0] i_cceip0_out_ia_rdata_part1;
input [31:0] i_cceip0_out_ia_rdata_part2;
input [11:0] i_cceip0_out_im_status;
input [1:0] i_cceip0_out_im_read_done;
input [19:0] i_cceip1_out_ia_capability;
input [16:0] i_cceip1_out_ia_status;
input [31:0] i_cceip1_out_ia_rdata_part0;
input [31:0] i_cceip1_out_ia_rdata_part1;
input [31:0] i_cceip1_out_ia_rdata_part2;
input [11:0] i_cceip1_out_im_status;
input [1:0] i_cceip1_out_im_read_done;
input [19:0] i_cceip2_out_ia_capability;
input [16:0] i_cceip2_out_ia_status;
input [31:0] i_cceip2_out_ia_rdata_part0;
input [31:0] i_cceip2_out_ia_rdata_part1;
input [31:0] i_cceip2_out_ia_rdata_part2;
input [11:0] i_cceip2_out_im_status;
input [1:0] i_cceip2_out_im_read_done;
input [19:0] i_cceip3_out_ia_capability;
input [16:0] i_cceip3_out_ia_status;
input [31:0] i_cceip3_out_ia_rdata_part0;
input [31:0] i_cceip3_out_ia_rdata_part1;
input [31:0] i_cceip3_out_ia_rdata_part2;
input [11:0] i_cceip3_out_im_status;
input [1:0] i_cceip3_out_im_read_done;
input [19:0] i_cddip0_out_ia_capability;
input [16:0] i_cddip0_out_ia_status;
input [31:0] i_cddip0_out_ia_rdata_part0;
input [31:0] i_cddip0_out_ia_rdata_part1;
input [31:0] i_cddip0_out_ia_rdata_part2;
input [11:0] i_cddip0_out_im_status;
input [1:0] i_cddip0_out_im_read_done;
input [19:0] i_cddip1_out_ia_capability;
input [16:0] i_cddip1_out_ia_status;
input [31:0] i_cddip1_out_ia_rdata_part0;
input [31:0] i_cddip1_out_ia_rdata_part1;
input [31:0] i_cddip1_out_ia_rdata_part2;
input [11:0] i_cddip1_out_im_status;
input [1:0] i_cddip1_out_im_read_done;
input [19:0] i_cddip2_out_ia_capability;
input [16:0] i_cddip2_out_ia_status;
input [31:0] i_cddip2_out_ia_rdata_part0;
input [31:0] i_cddip2_out_ia_rdata_part1;
input [31:0] i_cddip2_out_ia_rdata_part2;
input [11:0] i_cddip2_out_im_status;
input [1:0] i_cddip2_out_im_read_done;
input [19:0] i_cddip3_out_ia_capability;
input [16:0] i_cddip3_out_ia_status;
input [31:0] i_cddip3_out_ia_rdata_part0;
input [31:0] i_cddip3_out_ia_rdata_part1;
input [31:0] i_cddip3_out_ia_rdata_part2;
input [11:0] i_cddip3_out_im_status;
input [1:0] i_cddip3_out_im_read_done;
input [19:0] i_ckv_ia_capability;
input [22:0] i_ckv_ia_status;
input [31:0] i_ckv_ia_rdata_part0;
input [31:0] i_ckv_ia_rdata_part1;
input [19:0] i_kim_ia_capability;
input [21:0] i_kim_ia_status;
input [20:0] i_kim_ia_rdata_part0;
input [16:0] i_kim_ia_rdata_part1;
input [1:0] i_kdf_drbg_ctrl;
input [4:0] i_interrupt_status;
input [7:0] i_engine_sticky_status;
input [6:0] i_bimc_monitor;
input [31:0] i_bimc_ecc_uncorrectable_error_cnt;
input [31:0] i_bimc_ecc_correctable_error_cnt;
input [31:0] i_bimc_parity_error_cnt;
input [31:0] i_bimc_global_config;
input [11:0] i_bimc_memid;
input [28:0] i_bimc_eccpar_debug;
input [10:0] i_bimc_cmd2;
input [9:0] i_bimc_rxcmd2;
input [31:0] i_bimc_rxcmd1;
input [31:0] i_bimc_rxcmd0;
input [9:0] i_bimc_rxrsp2;
input [31:0] i_bimc_rxrsp1;
input [31:0] i_bimc_rxrsp0;
input [9:0] i_bimc_pollrsp2;
input [31:0] i_bimc_pollrsp1;
input [31:0] i_bimc_pollrsp0;
input [9:0] i_bimc_dbgcmd2;
input [31:0] i_bimc_dbgcmd1;
input [31:0] i_bimc_dbgcmd0;
input [15:0] i_im_available;
input [15:0] i_im_consumed;
input [8:0] i_tready_override;
input [31:0] i_regs_sa_ctrl;
input [19:0] i_sa_snapshot_ia_capability;
input [12:0] i_sa_snapshot_ia_status;
input [31:0] i_sa_snapshot_ia_rdata_part0;
input [31:0] i_sa_snapshot_ia_rdata_part1;
input [19:0] i_sa_count_ia_capability;
input [12:0] i_sa_count_ia_status;
input [31:0] i_sa_count_ia_rdata_part0;
input [31:0] i_sa_count_ia_rdata_part1;
input [31:0] i_idle_components;
input [31:0] i_sa_global_ctrl;
input [19:0] i_sa_ctrl_ia_capability;
input [12:0] i_sa_ctrl_ia_status;
input [31:0] i_sa_ctrl_ia_rdata_part0;
output o_reg_written;
output o_reg_read;
output [31:0] o_reg_wr_data;
output [10:0] o_reg_addr;
wire [10:0] ws_read_addr;
wire [10:0] ws_addr;
wire n_wr_strobe;
wire n_rd_strobe;
wire w_32b_aligned;
wire w_valid_rd_addr;
wire w_valid_wr_addr;
wire w_valid_addr;
wire w_do_write;
wire w_do_read;
wire [2:0] w_next_state;
wire w_next_ack;
wire w_next_err_ack;
wire [31:0] r32_formatted_reg_data;
wire w_load_spare_config;
wire w_load_cceip0_out_ia_wdata_part0;
wire w_load_cceip0_out_ia_wdata_part1;
wire w_load_cceip0_out_ia_wdata_part2;
wire w_load_cceip0_out_ia_config;
wire w_load_cceip0_out_im_config;
wire w_load_cceip0_out_im_read_done;
wire w_load_cceip1_out_ia_wdata_part0;
wire w_load_cceip1_out_ia_wdata_part1;
wire w_load_cceip1_out_ia_wdata_part2;
wire w_load_cceip1_out_ia_config;
wire w_load_cceip1_out_im_config;
wire w_load_cceip1_out_im_read_done;
wire w_load_cceip2_out_ia_wdata_part0;
wire w_load_cceip2_out_ia_wdata_part1;
wire w_load_cceip2_out_ia_wdata_part2;
wire w_load_cceip2_out_ia_config;
wire w_load_cceip2_out_im_config;
wire w_load_cceip2_out_im_read_done;
wire w_load_cceip3_out_ia_wdata_part0;
wire w_load_cceip3_out_ia_wdata_part1;
wire w_load_cceip3_out_ia_wdata_part2;
wire w_load_cceip3_out_ia_config;
wire w_load_cceip3_out_im_config;
wire w_load_cceip3_out_im_read_done;
wire w_load_cddip0_out_ia_wdata_part0;
wire w_load_cddip0_out_ia_wdata_part1;
wire w_load_cddip0_out_ia_wdata_part2;
wire w_load_cddip0_out_ia_config;
wire w_load_cddip0_out_im_config;
wire w_load_cddip0_out_im_read_done;
wire w_load_cddip1_out_ia_wdata_part0;
wire w_load_cddip1_out_ia_wdata_part1;
wire w_load_cddip1_out_ia_wdata_part2;
wire w_load_cddip1_out_ia_config;
wire w_load_cddip1_out_im_config;
wire w_load_cddip1_out_im_read_done;
wire w_load_cddip2_out_ia_wdata_part0;
wire w_load_cddip2_out_ia_wdata_part1;
wire w_load_cddip2_out_ia_wdata_part2;
wire w_load_cddip2_out_ia_config;
wire w_load_cddip2_out_im_config;
wire w_load_cddip2_out_im_read_done;
wire w_load_cddip3_out_ia_wdata_part0;
wire w_load_cddip3_out_ia_wdata_part1;
wire w_load_cddip3_out_ia_wdata_part2;
wire w_load_cddip3_out_ia_config;
wire w_load_cddip3_out_im_config;
wire w_load_cddip3_out_im_read_done;
wire w_load_ckv_ia_wdata_part0;
wire w_load_ckv_ia_wdata_part1;
wire w_load_ckv_ia_config;
wire w_load_kim_ia_wdata_part0;
wire w_load_kim_ia_wdata_part1;
wire w_load_kim_ia_config;
wire w_load_label0_config;
wire w_load_label0_data7;
wire w_load_label0_data6;
wire w_load_label0_data5;
wire w_load_label0_data4;
wire w_load_label0_data3;
wire w_load_label0_data2;
wire w_load_label0_data1;
wire w_load_label0_data0;
wire w_load_label1_config;
wire w_load_label1_data7;
wire w_load_label1_data6;
wire w_load_label1_data5;
wire w_load_label1_data4;
wire w_load_label1_data3;
wire w_load_label1_data2;
wire w_load_label1_data1;
wire w_load_label1_data0;
wire w_load_label2_config;
wire w_load_label2_data7;
wire w_load_label2_data6;
wire w_load_label2_data5;
wire w_load_label2_data4;
wire w_load_label2_data3;
wire w_load_label2_data2;
wire w_load_label2_data1;
wire w_load_label2_data0;
wire w_load_label3_config;
wire w_load_label3_data7;
wire w_load_label3_data6;
wire w_load_label3_data5;
wire w_load_label3_data4;
wire w_load_label3_data3;
wire w_load_label3_data2;
wire w_load_label3_data1;
wire w_load_label3_data0;
wire w_load_label4_config;
wire w_load_label4_data7;
wire w_load_label4_data6;
wire w_load_label4_data5;
wire w_load_label4_data4;
wire w_load_label4_data3;
wire w_load_label4_data2;
wire w_load_label4_data1;
wire w_load_label4_data0;
wire w_load_label5_config;
wire w_load_label5_data7;
wire w_load_label5_data6;
wire w_load_label5_data5;
wire w_load_label5_data4;
wire w_load_label5_data3;
wire w_load_label5_data2;
wire w_load_label5_data1;
wire w_load_label5_data0;
wire w_load_label6_config;
wire w_load_label6_data7;
wire w_load_label6_data6;
wire w_load_label6_data5;
wire w_load_label6_data4;
wire w_load_label6_data3;
wire w_load_label6_data2;
wire w_load_label6_data1;
wire w_load_label6_data0;
wire w_load_label7_config;
wire w_load_label7_data7;
wire w_load_label7_data6;
wire w_load_label7_data5;
wire w_load_label7_data4;
wire w_load_label7_data3;
wire w_load_label7_data2;
wire w_load_label7_data1;
wire w_load_label7_data0;
wire w_load_kdf_drbg_ctrl;
wire w_load_kdf_drbg_seed_0_state_key_31_0;
wire w_load_kdf_drbg_seed_0_state_key_63_32;
wire w_load_kdf_drbg_seed_0_state_key_95_64;
wire w_load_kdf_drbg_seed_0_state_key_127_96;
wire w_load_kdf_drbg_seed_0_state_key_159_128;
wire w_load_kdf_drbg_seed_0_state_key_191_160;
wire w_load_kdf_drbg_seed_0_state_key_223_192;
wire w_load_kdf_drbg_seed_0_state_key_255_224;
wire w_load_kdf_drbg_seed_0_state_value_31_0;
wire w_load_kdf_drbg_seed_0_state_value_63_32;
wire w_load_kdf_drbg_seed_0_state_value_95_64;
wire w_load_kdf_drbg_seed_0_state_value_127_96;
wire w_load_kdf_drbg_seed_0_reseed_interval_0;
wire w_load_kdf_drbg_seed_0_reseed_interval_1;
wire w_load_kdf_drbg_seed_1_state_key_31_0;
wire w_load_kdf_drbg_seed_1_state_key_63_32;
wire w_load_kdf_drbg_seed_1_state_key_95_64;
wire w_load_kdf_drbg_seed_1_state_key_127_96;
wire w_load_kdf_drbg_seed_1_state_key_159_128;
wire w_load_kdf_drbg_seed_1_state_key_191_160;
wire w_load_kdf_drbg_seed_1_state_key_223_192;
wire w_load_kdf_drbg_seed_1_state_key_255_224;
wire w_load_kdf_drbg_seed_1_state_value_31_0;
wire w_load_kdf_drbg_seed_1_state_value_63_32;
wire w_load_kdf_drbg_seed_1_state_value_95_64;
wire w_load_kdf_drbg_seed_1_state_value_127_96;
wire w_load_kdf_drbg_seed_1_reseed_interval_0;
wire w_load_kdf_drbg_seed_1_reseed_interval_1;
wire w_load_interrupt_status;
wire w_load_interrupt_mask;
wire w_load_engine_sticky_status;
wire w_load_bimc_monitor_mask;
wire w_load_bimc_ecc_uncorrectable_error_cnt;
wire w_load_bimc_ecc_correctable_error_cnt;
wire w_load_bimc_parity_error_cnt;
wire w_load_bimc_global_config;
wire w_load_bimc_eccpar_debug;
wire w_load_bimc_cmd2;
wire w_load_bimc_cmd1;
wire w_load_bimc_cmd0;
wire w_load_bimc_rxcmd2;
wire w_load_bimc_rxrsp2;
wire w_load_bimc_pollrsp2;
wire w_load_bimc_dbgcmd2;
wire w_load_im_consumed;
wire w_load_tready_override;
wire w_load_regs_sa_ctrl;
wire w_load_sa_snapshot_ia_wdata_part0;
wire w_load_sa_snapshot_ia_wdata_part1;
wire w_load_sa_snapshot_ia_config;
wire w_load_sa_count_ia_wdata_part0;
wire w_load_sa_count_ia_wdata_part1;
wire w_load_sa_count_ia_config;
wire w_load_cceip_encrypt_kop_fifo_override;
wire w_load_cceip_validate_kop_fifo_override;
wire w_load_cddip_decrypt_kop_fifo_override;
wire w_load_sa_global_ctrl;
wire w_load_sa_ctrl_ia_wdata_part0;
wire w_load_sa_ctrl_ia_config;
wire w_load_kdf_test_key_size_config;
wire _zy_simnet_o_reg_written_0_w$;
wire _zy_simnet_o_reg_read_1_w$;
wire [0:10] _zy_simnet_o_reg_addr_2_w$;
wire [0:31] _zy_simnet_f32_data_3_w$;
wire n_write;
wire [2:0] f_state;
wire f_prev_do_read;
wire f_ack;
wire f_err_ack;
wire [31:0] r32_mux_0_data;
wire [31:0] f32_mux_0_data;
wire [31:0] r32_mux_1_data;
wire [31:0] f32_mux_1_data;
wire [31:0] r32_mux_2_data;
wire [31:0] f32_mux_2_data;
wire [31:0] r32_mux_3_data;
wire [31:0] f32_mux_3_data;
wire [31:0] r32_mux_4_data;
wire [31:0] f32_mux_4_data;
wire [31:0] r32_mux_5_data;
wire [31:0] f32_mux_5_data;
wire [31:0] r32_mux_6_data;
wire [31:0] f32_mux_6_data;
wire [31:0] r32_mux_7_data;
wire [31:0] f32_mux_7_data;
wire [31:0] r32_mux_8_data;
wire [31:0] f32_mux_8_data;
wire [31:0] f32_data;
supply0 n4920;
Q_BUF U0 ( .A(w_next_ack), .Z(w_do_read));
Q_BUF U1 ( .A(w_valid_addr), .Z(w_valid_rd_addr));
Q_BUF U2 ( .A(w_valid_wr_addr), .Z(w_valid_addr));
cr_kme_regs_flops u_cr_kme_regs_flops ( .clk( clk), .i_reset_( i_reset_), 
	.i_sw_init( i_sw_init), .o_spare_config( o_spare_config[31:0]), 
	.o_cceip0_out_ia_wdata_part0( o_cceip0_out_ia_wdata_part0[31:0]), 
	.o_cceip0_out_ia_wdata_part1( o_cceip0_out_ia_wdata_part1[31:0]), 
	.o_cceip0_out_ia_wdata_part2( o_cceip0_out_ia_wdata_part2[31:0]), 
	.o_cceip0_out_ia_config( o_cceip0_out_ia_config[12:0]), 
	.o_cceip0_out_im_config( o_cceip0_out_im_config[11:0]), 
	.o_cceip0_out_im_read_done( o_cceip0_out_im_read_done[1:0]), 
	.o_cceip1_out_ia_wdata_part0( o_cceip1_out_ia_wdata_part0[31:0]), 
	.o_cceip1_out_ia_wdata_part1( o_cceip1_out_ia_wdata_part1[31:0]), 
	.o_cceip1_out_ia_wdata_part2( o_cceip1_out_ia_wdata_part2[31:0]), 
	.o_cceip1_out_ia_config( o_cceip1_out_ia_config[12:0]), 
	.o_cceip1_out_im_config( o_cceip1_out_im_config[11:0]), 
	.o_cceip1_out_im_read_done( o_cceip1_out_im_read_done[1:0]), 
	.o_cceip2_out_ia_wdata_part0( o_cceip2_out_ia_wdata_part0[31:0]), 
	.o_cceip2_out_ia_wdata_part1( o_cceip2_out_ia_wdata_part1[31:0]), 
	.o_cceip2_out_ia_wdata_part2( o_cceip2_out_ia_wdata_part2[31:0]), 
	.o_cceip2_out_ia_config( o_cceip2_out_ia_config[12:0]), 
	.o_cceip2_out_im_config( o_cceip2_out_im_config[11:0]), 
	.o_cceip2_out_im_read_done( o_cceip2_out_im_read_done[1:0]), 
	.o_cceip3_out_ia_wdata_part0( o_cceip3_out_ia_wdata_part0[31:0]), 
	.o_cceip3_out_ia_wdata_part1( o_cceip3_out_ia_wdata_part1[31:0]), 
	.o_cceip3_out_ia_wdata_part2( o_cceip3_out_ia_wdata_part2[31:0]), 
	.o_cceip3_out_ia_config( o_cceip3_out_ia_config[12:0]), 
	.o_cceip3_out_im_config( o_cceip3_out_im_config[11:0]), 
	.o_cceip3_out_im_read_done( o_cceip3_out_im_read_done[1:0]), 
	.o_cddip0_out_ia_wdata_part0( o_cddip0_out_ia_wdata_part0[31:0]), 
	.o_cddip0_out_ia_wdata_part1( o_cddip0_out_ia_wdata_part1[31:0]), 
	.o_cddip0_out_ia_wdata_part2( o_cddip0_out_ia_wdata_part2[31:0]), 
	.o_cddip0_out_ia_config( o_cddip0_out_ia_config[12:0]), 
	.o_cddip0_out_im_config( o_cddip0_out_im_config[11:0]), 
	.o_cddip0_out_im_read_done( o_cddip0_out_im_read_done[1:0]), 
	.o_cddip1_out_ia_wdata_part0( o_cddip1_out_ia_wdata_part0[31:0]), 
	.o_cddip1_out_ia_wdata_part1( o_cddip1_out_ia_wdata_part1[31:0]), 
	.o_cddip1_out_ia_wdata_part2( o_cddip1_out_ia_wdata_part2[31:0]), 
	.o_cddip1_out_ia_config( o_cddip1_out_ia_config[12:0]), 
	.o_cddip1_out_im_config( o_cddip1_out_im_config[11:0]), 
	.o_cddip1_out_im_read_done( o_cddip1_out_im_read_done[1:0]), 
	.o_cddip2_out_ia_wdata_part0( o_cddip2_out_ia_wdata_part0[31:0]), 
	.o_cddip2_out_ia_wdata_part1( o_cddip2_out_ia_wdata_part1[31:0]), 
	.o_cddip2_out_ia_wdata_part2( o_cddip2_out_ia_wdata_part2[31:0]), 
	.o_cddip2_out_ia_config( o_cddip2_out_ia_config[12:0]), 
	.o_cddip2_out_im_config( o_cddip2_out_im_config[11:0]), 
	.o_cddip2_out_im_read_done( o_cddip2_out_im_read_done[1:0]), 
	.o_cddip3_out_ia_wdata_part0( o_cddip3_out_ia_wdata_part0[31:0]), 
	.o_cddip3_out_ia_wdata_part1( o_cddip3_out_ia_wdata_part1[31:0]), 
	.o_cddip3_out_ia_wdata_part2( o_cddip3_out_ia_wdata_part2[31:0]), 
	.o_cddip3_out_ia_config( o_cddip3_out_ia_config[12:0]), 
	.o_cddip3_out_im_config( o_cddip3_out_im_config[11:0]), 
	.o_cddip3_out_im_read_done( o_cddip3_out_im_read_done[1:0]), 
	.o_ckv_ia_wdata_part0( o_ckv_ia_wdata_part0[31:0]), 
	.o_ckv_ia_wdata_part1( o_ckv_ia_wdata_part1[31:0]), 
	.o_ckv_ia_config( o_ckv_ia_config[18:0]), .o_kim_ia_wdata_part0( 
	o_kim_ia_wdata_part0[20:0]), .o_kim_ia_wdata_part1( 
	o_kim_ia_wdata_part1[16:0]), .o_kim_ia_config( 
	o_kim_ia_config[17:0]), .o_label0_config( o_label0_config[15:0]), 
	.o_label0_data7( o_label0_data7[31:0]), .o_label0_data6( 
	o_label0_data6[31:0]), .o_label0_data5( o_label0_data5[31:0]), 
	.o_label0_data4( o_label0_data4[31:0]), .o_label0_data3( 
	o_label0_data3[31:0]), .o_label0_data2( o_label0_data2[31:0]), 
	.o_label0_data1( o_label0_data1[31:0]), .o_label0_data0( 
	o_label0_data0[31:0]), .o_label1_config( o_label1_config[15:0]), 
	.o_label1_data7( o_label1_data7[31:0]), .o_label1_data6( 
	o_label1_data6[31:0]), .o_label1_data5( o_label1_data5[31:0]), 
	.o_label1_data4( o_label1_data4[31:0]), .o_label1_data3( 
	o_label1_data3[31:0]), .o_label1_data2( o_label1_data2[31:0]), 
	.o_label1_data1( o_label1_data1[31:0]), .o_label1_data0( 
	o_label1_data0[31:0]), .o_label2_config( o_label2_config[15:0]), 
	.o_label2_data7( o_label2_data7[31:0]), .o_label2_data6( 
	o_label2_data6[31:0]), .o_label2_data5( o_label2_data5[31:0]), 
	.o_label2_data4( o_label2_data4[31:0]), .o_label2_data3( 
	o_label2_data3[31:0]), .o_label2_data2( o_label2_data2[31:0]), 
	.o_label2_data1( o_label2_data1[31:0]), .o_label2_data0( 
	o_label2_data0[31:0]), .o_label3_config( o_label3_config[15:0]), 
	.o_label3_data7( o_label3_data7[31:0]), .o_label3_data6( 
	o_label3_data6[31:0]), .o_label3_data5( o_label3_data5[31:0]), 
	.o_label3_data4( o_label3_data4[31:0]), .o_label3_data3( 
	o_label3_data3[31:0]), .o_label3_data2( o_label3_data2[31:0]), 
	.o_label3_data1( o_label3_data1[31:0]), .o_label3_data0( 
	o_label3_data0[31:0]), .o_label4_config( o_label4_config[15:0]), 
	.o_label4_data7( o_label4_data7[31:0]), .o_label4_data6( 
	o_label4_data6[31:0]), .o_label4_data5( o_label4_data5[31:0]), 
	.o_label4_data4( o_label4_data4[31:0]), .o_label4_data3( 
	o_label4_data3[31:0]), .o_label4_data2( o_label4_data2[31:0]), 
	.o_label4_data1( o_label4_data1[31:0]), .o_label4_data0( 
	o_label4_data0[31:0]), .o_label5_config( o_label5_config[15:0]), 
	.o_label5_data7( o_label5_data7[31:0]), .o_label5_data6( 
	o_label5_data6[31:0]), .o_label5_data5( o_label5_data5[31:0]), 
	.o_label5_data4( o_label5_data4[31:0]), .o_label5_data3( 
	o_label5_data3[31:0]), .o_label5_data2( o_label5_data2[31:0]), 
	.o_label5_data1( o_label5_data1[31:0]), .o_label5_data0( 
	o_label5_data0[31:0]), .o_label6_config( o_label6_config[15:0]), 
	.o_label6_data7( o_label6_data7[31:0]), .o_label6_data6( 
	o_label6_data6[31:0]), .o_label6_data5( o_label6_data5[31:0]), 
	.o_label6_data4( o_label6_data4[31:0]), .o_label6_data3( 
	o_label6_data3[31:0]), .o_label6_data2( o_label6_data2[31:0]), 
	.o_label6_data1( o_label6_data1[31:0]), .o_label6_data0( 
	o_label6_data0[31:0]), .o_label7_config( o_label7_config[15:0]), 
	.o_label7_data7( o_label7_data7[31:0]), .o_label7_data6( 
	o_label7_data6[31:0]), .o_label7_data5( o_label7_data5[31:0]), 
	.o_label7_data4( o_label7_data4[31:0]), .o_label7_data3( 
	o_label7_data3[31:0]), .o_label7_data2( o_label7_data2[31:0]), 
	.o_label7_data1( o_label7_data1[31:0]), .o_label7_data0( 
	o_label7_data0[31:0]), .o_kdf_drbg_ctrl( o_kdf_drbg_ctrl[1:0]), 
	.o_kdf_drbg_seed_0_state_key_31_0( 
	o_kdf_drbg_seed_0_state_key_31_0[31:0]), 
	.o_kdf_drbg_seed_0_state_key_63_32( 
	o_kdf_drbg_seed_0_state_key_63_32[31:0]), 
	.o_kdf_drbg_seed_0_state_key_95_64( 
	o_kdf_drbg_seed_0_state_key_95_64[31:0]), 
	.o_kdf_drbg_seed_0_state_key_127_96( 
	o_kdf_drbg_seed_0_state_key_127_96[31:0]), 
	.o_kdf_drbg_seed_0_state_key_159_128( 
	o_kdf_drbg_seed_0_state_key_159_128[31:0]), 
	.o_kdf_drbg_seed_0_state_key_191_160( 
	o_kdf_drbg_seed_0_state_key_191_160[31:0]), 
	.o_kdf_drbg_seed_0_state_key_223_192( 
	o_kdf_drbg_seed_0_state_key_223_192[31:0]), 
	.o_kdf_drbg_seed_0_state_key_255_224( 
	o_kdf_drbg_seed_0_state_key_255_224[31:0]), 
	.o_kdf_drbg_seed_0_state_value_31_0( 
	o_kdf_drbg_seed_0_state_value_31_0[31:0]), 
	.o_kdf_drbg_seed_0_state_value_63_32( 
	o_kdf_drbg_seed_0_state_value_63_32[31:0]), 
	.o_kdf_drbg_seed_0_state_value_95_64( 
	o_kdf_drbg_seed_0_state_value_95_64[31:0]), 
	.o_kdf_drbg_seed_0_state_value_127_96( 
	o_kdf_drbg_seed_0_state_value_127_96[31:0]), 
	.o_kdf_drbg_seed_0_reseed_interval_0( 
	o_kdf_drbg_seed_0_reseed_interval_0[31:0]), 
	.o_kdf_drbg_seed_0_reseed_interval_1( 
	o_kdf_drbg_seed_0_reseed_interval_1[15:0]), 
	.o_kdf_drbg_seed_1_state_key_31_0( 
	o_kdf_drbg_seed_1_state_key_31_0[31:0]), 
	.o_kdf_drbg_seed_1_state_key_63_32( 
	o_kdf_drbg_seed_1_state_key_63_32[31:0]), 
	.o_kdf_drbg_seed_1_state_key_95_64( 
	o_kdf_drbg_seed_1_state_key_95_64[31:0]), 
	.o_kdf_drbg_seed_1_state_key_127_96( 
	o_kdf_drbg_seed_1_state_key_127_96[31:0]), 
	.o_kdf_drbg_seed_1_state_key_159_128( 
	o_kdf_drbg_seed_1_state_key_159_128[31:0]), 
	.o_kdf_drbg_seed_1_state_key_191_160( 
	o_kdf_drbg_seed_1_state_key_191_160[31:0]), 
	.o_kdf_drbg_seed_1_state_key_223_192( 
	o_kdf_drbg_seed_1_state_key_223_192[31:0]), 
	.o_kdf_drbg_seed_1_state_key_255_224( 
	o_kdf_drbg_seed_1_state_key_255_224[31:0]), 
	.o_kdf_drbg_seed_1_state_value_31_0( 
	o_kdf_drbg_seed_1_state_value_31_0[31:0]), 
	.o_kdf_drbg_seed_1_state_value_63_32( 
	o_kdf_drbg_seed_1_state_value_63_32[31:0]), 
	.o_kdf_drbg_seed_1_state_value_95_64( 
	o_kdf_drbg_seed_1_state_value_95_64[31:0]), 
	.o_kdf_drbg_seed_1_state_value_127_96( 
	o_kdf_drbg_seed_1_state_value_127_96[31:0]), 
	.o_kdf_drbg_seed_1_reseed_interval_0( 
	o_kdf_drbg_seed_1_reseed_interval_0[31:0]), 
	.o_kdf_drbg_seed_1_reseed_interval_1( 
	o_kdf_drbg_seed_1_reseed_interval_1[15:0]), .o_interrupt_status( 
	o_interrupt_status[4:0]), .o_interrupt_mask( o_interrupt_mask[4:0]), 
	.o_engine_sticky_status( o_engine_sticky_status[7:0]), 
	.o_bimc_monitor_mask( o_bimc_monitor_mask[6:0]), 
	.o_bimc_ecc_uncorrectable_error_cnt( 
	o_bimc_ecc_uncorrectable_error_cnt[31:0]), 
	.o_bimc_ecc_correctable_error_cnt( 
	o_bimc_ecc_correctable_error_cnt[31:0]), .o_bimc_parity_error_cnt( 
	o_bimc_parity_error_cnt[31:0]), .o_bimc_global_config( 
	o_bimc_global_config[31:0]), .o_bimc_eccpar_debug( 
	o_bimc_eccpar_debug[28:0]), .o_bimc_cmd2( o_bimc_cmd2[10:0]), 
	.o_bimc_cmd1( o_bimc_cmd1[31:0]), .o_bimc_cmd0( 
	o_bimc_cmd0[31:0]), .o_bimc_rxcmd2( o_bimc_rxcmd2[9:0]), 
	.o_bimc_rxrsp2( o_bimc_rxrsp2[9:0]), .o_bimc_pollrsp2( 
	o_bimc_pollrsp2[9:0]), .o_bimc_dbgcmd2( o_bimc_dbgcmd2[9:0]), 
	.o_im_consumed( o_im_consumed[15:0]), .o_tready_override( 
	o_tready_override[8:0]), .o_regs_sa_ctrl( o_regs_sa_ctrl[31:0]), 
	.o_sa_snapshot_ia_wdata_part0( o_sa_snapshot_ia_wdata_part0[31:0]), 
	.o_sa_snapshot_ia_wdata_part1( o_sa_snapshot_ia_wdata_part1[31:0]), 
	.o_sa_snapshot_ia_config( o_sa_snapshot_ia_config[8:0]), 
	.o_sa_count_ia_wdata_part0( o_sa_count_ia_wdata_part0[31:0]), 
	.o_sa_count_ia_wdata_part1( o_sa_count_ia_wdata_part1[31:0]), 
	.o_sa_count_ia_config( o_sa_count_ia_config[8:0]), 
	.o_cceip_encrypt_kop_fifo_override( 
	o_cceip_encrypt_kop_fifo_override[6:0]), 
	.o_cceip_validate_kop_fifo_override( 
	o_cceip_validate_kop_fifo_override[6:0]), 
	.o_cddip_decrypt_kop_fifo_override( 
	o_cddip_decrypt_kop_fifo_override[6:0]), .o_sa_global_ctrl( 
	o_sa_global_ctrl[31:0]), .o_sa_ctrl_ia_wdata_part0( 
	o_sa_ctrl_ia_wdata_part0[31:0]), .o_sa_ctrl_ia_config( 
	o_sa_ctrl_ia_config[8:0]), .o_kdf_test_key_size_config( 
	o_kdf_test_key_size_config[31:0]), .w_load_spare_config( 
	w_load_spare_config), .w_load_cceip0_out_ia_wdata_part0( 
	w_load_cceip0_out_ia_wdata_part0), 
	.w_load_cceip0_out_ia_wdata_part1( w_load_cceip0_out_ia_wdata_part1), 
	.w_load_cceip0_out_ia_wdata_part2( w_load_cceip0_out_ia_wdata_part2), 
	.w_load_cceip0_out_ia_config( w_load_cceip0_out_ia_config), 
	.w_load_cceip0_out_im_config( w_load_cceip0_out_im_config), 
	.w_load_cceip0_out_im_read_done( w_load_cceip0_out_im_read_done), 
	.w_load_cceip1_out_ia_wdata_part0( w_load_cceip1_out_ia_wdata_part0), 
	.w_load_cceip1_out_ia_wdata_part1( w_load_cceip1_out_ia_wdata_part1), 
	.w_load_cceip1_out_ia_wdata_part2( w_load_cceip1_out_ia_wdata_part2), 
	.w_load_cceip1_out_ia_config( w_load_cceip1_out_ia_config), 
	.w_load_cceip1_out_im_config( w_load_cceip1_out_im_config), 
	.w_load_cceip1_out_im_read_done( w_load_cceip1_out_im_read_done), 
	.w_load_cceip2_out_ia_wdata_part0( w_load_cceip2_out_ia_wdata_part0), 
	.w_load_cceip2_out_ia_wdata_part1( w_load_cceip2_out_ia_wdata_part1), 
	.w_load_cceip2_out_ia_wdata_part2( w_load_cceip2_out_ia_wdata_part2), 
	.w_load_cceip2_out_ia_config( w_load_cceip2_out_ia_config), 
	.w_load_cceip2_out_im_config( w_load_cceip2_out_im_config), 
	.w_load_cceip2_out_im_read_done( w_load_cceip2_out_im_read_done), 
	.w_load_cceip3_out_ia_wdata_part0( w_load_cceip3_out_ia_wdata_part0), 
	.w_load_cceip3_out_ia_wdata_part1( w_load_cceip3_out_ia_wdata_part1), 
	.w_load_cceip3_out_ia_wdata_part2( w_load_cceip3_out_ia_wdata_part2), 
	.w_load_cceip3_out_ia_config( w_load_cceip3_out_ia_config), 
	.w_load_cceip3_out_im_config( w_load_cceip3_out_im_config), 
	.w_load_cceip3_out_im_read_done( w_load_cceip3_out_im_read_done), 
	.w_load_cddip0_out_ia_wdata_part0( w_load_cddip0_out_ia_wdata_part0), 
	.w_load_cddip0_out_ia_wdata_part1( w_load_cddip0_out_ia_wdata_part1), 
	.w_load_cddip0_out_ia_wdata_part2( w_load_cddip0_out_ia_wdata_part2), 
	.w_load_cddip0_out_ia_config( w_load_cddip0_out_ia_config), 
	.w_load_cddip0_out_im_config( w_load_cddip0_out_im_config), 
	.w_load_cddip0_out_im_read_done( w_load_cddip0_out_im_read_done), 
	.w_load_cddip1_out_ia_wdata_part0( w_load_cddip1_out_ia_wdata_part0), 
	.w_load_cddip1_out_ia_wdata_part1( w_load_cddip1_out_ia_wdata_part1), 
	.w_load_cddip1_out_ia_wdata_part2( w_load_cddip1_out_ia_wdata_part2), 
	.w_load_cddip1_out_ia_config( w_load_cddip1_out_ia_config), 
	.w_load_cddip1_out_im_config( w_load_cddip1_out_im_config), 
	.w_load_cddip1_out_im_read_done( w_load_cddip1_out_im_read_done), 
	.w_load_cddip2_out_ia_wdata_part0( w_load_cddip2_out_ia_wdata_part0), 
	.w_load_cddip2_out_ia_wdata_part1( w_load_cddip2_out_ia_wdata_part1), 
	.w_load_cddip2_out_ia_wdata_part2( w_load_cddip2_out_ia_wdata_part2), 
	.w_load_cddip2_out_ia_config( w_load_cddip2_out_ia_config), 
	.w_load_cddip2_out_im_config( w_load_cddip2_out_im_config), 
	.w_load_cddip2_out_im_read_done( w_load_cddip2_out_im_read_done), 
	.w_load_cddip3_out_ia_wdata_part0( w_load_cddip3_out_ia_wdata_part0), 
	.w_load_cddip3_out_ia_wdata_part1( w_load_cddip3_out_ia_wdata_part1), 
	.w_load_cddip3_out_ia_wdata_part2( w_load_cddip3_out_ia_wdata_part2), 
	.w_load_cddip3_out_ia_config( w_load_cddip3_out_ia_config), 
	.w_load_cddip3_out_im_config( w_load_cddip3_out_im_config), 
	.w_load_cddip3_out_im_read_done( w_load_cddip3_out_im_read_done), 
	.w_load_ckv_ia_wdata_part0( w_load_ckv_ia_wdata_part0), 
	.w_load_ckv_ia_wdata_part1( w_load_ckv_ia_wdata_part1), 
	.w_load_ckv_ia_config( w_load_ckv_ia_config), 
	.w_load_kim_ia_wdata_part0( w_load_kim_ia_wdata_part0), 
	.w_load_kim_ia_wdata_part1( w_load_kim_ia_wdata_part1), 
	.w_load_kim_ia_config( w_load_kim_ia_config), 
	.w_load_label0_config( w_load_label0_config), .w_load_label0_data7( 
	w_load_label0_data7), .w_load_label0_data6( w_load_label0_data6), 
	.w_load_label0_data5( w_load_label0_data5), .w_load_label0_data4( 
	w_load_label0_data4), .w_load_label0_data3( w_load_label0_data3), 
	.w_load_label0_data2( w_load_label0_data2), .w_load_label0_data1( 
	w_load_label0_data1), .w_load_label0_data0( w_load_label0_data0), 
	.w_load_label1_config( w_load_label1_config), .w_load_label1_data7( 
	w_load_label1_data7), .w_load_label1_data6( w_load_label1_data6), 
	.w_load_label1_data5( w_load_label1_data5), .w_load_label1_data4( 
	w_load_label1_data4), .w_load_label1_data3( w_load_label1_data3), 
	.w_load_label1_data2( w_load_label1_data2), .w_load_label1_data1( 
	w_load_label1_data1), .w_load_label1_data0( w_load_label1_data0), 
	.w_load_label2_config( w_load_label2_config), .w_load_label2_data7( 
	w_load_label2_data7), .w_load_label2_data6( w_load_label2_data6), 
	.w_load_label2_data5( w_load_label2_data5), .w_load_label2_data4( 
	w_load_label2_data4), .w_load_label2_data3( w_load_label2_data3), 
	.w_load_label2_data2( w_load_label2_data2), .w_load_label2_data1( 
	w_load_label2_data1), .w_load_label2_data0( w_load_label2_data0), 
	.w_load_label3_config( w_load_label3_config), .w_load_label3_data7( 
	w_load_label3_data7), .w_load_label3_data6( w_load_label3_data6), 
	.w_load_label3_data5( w_load_label3_data5), .w_load_label3_data4( 
	w_load_label3_data4), .w_load_label3_data3( w_load_label3_data3), 
	.w_load_label3_data2( w_load_label3_data2), .w_load_label3_data1( 
	w_load_label3_data1), .w_load_label3_data0( w_load_label3_data0), 
	.w_load_label4_config( w_load_label4_config), .w_load_label4_data7( 
	w_load_label4_data7), .w_load_label4_data6( w_load_label4_data6), 
	.w_load_label4_data5( w_load_label4_data5), .w_load_label4_data4( 
	w_load_label4_data4), .w_load_label4_data3( w_load_label4_data3), 
	.w_load_label4_data2( w_load_label4_data2), .w_load_label4_data1( 
	w_load_label4_data1), .w_load_label4_data0( w_load_label4_data0), 
	.w_load_label5_config( w_load_label5_config), .w_load_label5_data7( 
	w_load_label5_data7), .w_load_label5_data6( w_load_label5_data6), 
	.w_load_label5_data5( w_load_label5_data5), .w_load_label5_data4( 
	w_load_label5_data4), .w_load_label5_data3( w_load_label5_data3), 
	.w_load_label5_data2( w_load_label5_data2), .w_load_label5_data1( 
	w_load_label5_data1), .w_load_label5_data0( w_load_label5_data0), 
	.w_load_label6_config( w_load_label6_config), .w_load_label6_data7( 
	w_load_label6_data7), .w_load_label6_data6( w_load_label6_data6), 
	.w_load_label6_data5( w_load_label6_data5), .w_load_label6_data4( 
	w_load_label6_data4), .w_load_label6_data3( w_load_label6_data3), 
	.w_load_label6_data2( w_load_label6_data2), .w_load_label6_data1( 
	w_load_label6_data1), .w_load_label6_data0( w_load_label6_data0), 
	.w_load_label7_config( w_load_label7_config), .w_load_label7_data7( 
	w_load_label7_data7), .w_load_label7_data6( w_load_label7_data6), 
	.w_load_label7_data5( w_load_label7_data5), .w_load_label7_data4( 
	w_load_label7_data4), .w_load_label7_data3( w_load_label7_data3), 
	.w_load_label7_data2( w_load_label7_data2), .w_load_label7_data1( 
	w_load_label7_data1), .w_load_label7_data0( w_load_label7_data0), 
	.w_load_kdf_drbg_ctrl( w_load_kdf_drbg_ctrl), 
	.w_load_kdf_drbg_seed_0_state_key_31_0( 
	w_load_kdf_drbg_seed_0_state_key_31_0), 
	.w_load_kdf_drbg_seed_0_state_key_63_32( 
	w_load_kdf_drbg_seed_0_state_key_63_32), 
	.w_load_kdf_drbg_seed_0_state_key_95_64( 
	w_load_kdf_drbg_seed_0_state_key_95_64), 
	.w_load_kdf_drbg_seed_0_state_key_127_96( 
	w_load_kdf_drbg_seed_0_state_key_127_96), 
	.w_load_kdf_drbg_seed_0_state_key_159_128( 
	w_load_kdf_drbg_seed_0_state_key_159_128), 
	.w_load_kdf_drbg_seed_0_state_key_191_160( 
	w_load_kdf_drbg_seed_0_state_key_191_160), 
	.w_load_kdf_drbg_seed_0_state_key_223_192( 
	w_load_kdf_drbg_seed_0_state_key_223_192), 
	.w_load_kdf_drbg_seed_0_state_key_255_224( 
	w_load_kdf_drbg_seed_0_state_key_255_224), 
	.w_load_kdf_drbg_seed_0_state_value_31_0( 
	w_load_kdf_drbg_seed_0_state_value_31_0), 
	.w_load_kdf_drbg_seed_0_state_value_63_32( 
	w_load_kdf_drbg_seed_0_state_value_63_32), 
	.w_load_kdf_drbg_seed_0_state_value_95_64( 
	w_load_kdf_drbg_seed_0_state_value_95_64), 
	.w_load_kdf_drbg_seed_0_state_value_127_96( 
	w_load_kdf_drbg_seed_0_state_value_127_96), 
	.w_load_kdf_drbg_seed_0_reseed_interval_0( 
	w_load_kdf_drbg_seed_0_reseed_interval_0), 
	.w_load_kdf_drbg_seed_0_reseed_interval_1( 
	w_load_kdf_drbg_seed_0_reseed_interval_1), 
	.w_load_kdf_drbg_seed_1_state_key_31_0( 
	w_load_kdf_drbg_seed_1_state_key_31_0), 
	.w_load_kdf_drbg_seed_1_state_key_63_32( 
	w_load_kdf_drbg_seed_1_state_key_63_32), 
	.w_load_kdf_drbg_seed_1_state_key_95_64( 
	w_load_kdf_drbg_seed_1_state_key_95_64), 
	.w_load_kdf_drbg_seed_1_state_key_127_96( 
	w_load_kdf_drbg_seed_1_state_key_127_96), 
	.w_load_kdf_drbg_seed_1_state_key_159_128( 
	w_load_kdf_drbg_seed_1_state_key_159_128), 
	.w_load_kdf_drbg_seed_1_state_key_191_160( 
	w_load_kdf_drbg_seed_1_state_key_191_160), 
	.w_load_kdf_drbg_seed_1_state_key_223_192( 
	w_load_kdf_drbg_seed_1_state_key_223_192), 
	.w_load_kdf_drbg_seed_1_state_key_255_224( 
	w_load_kdf_drbg_seed_1_state_key_255_224), 
	.w_load_kdf_drbg_seed_1_state_value_31_0( 
	w_load_kdf_drbg_seed_1_state_value_31_0), 
	.w_load_kdf_drbg_seed_1_state_value_63_32( 
	w_load_kdf_drbg_seed_1_state_value_63_32), 
	.w_load_kdf_drbg_seed_1_state_value_95_64( 
	w_load_kdf_drbg_seed_1_state_value_95_64), 
	.w_load_kdf_drbg_seed_1_state_value_127_96( 
	w_load_kdf_drbg_seed_1_state_value_127_96), 
	.w_load_kdf_drbg_seed_1_reseed_interval_0( 
	w_load_kdf_drbg_seed_1_reseed_interval_0), 
	.w_load_kdf_drbg_seed_1_reseed_interval_1( 
	w_load_kdf_drbg_seed_1_reseed_interval_1), .w_load_interrupt_status( 
	w_load_interrupt_status), .w_load_interrupt_mask( 
	w_load_interrupt_mask), .w_load_engine_sticky_status( 
	w_load_engine_sticky_status), .w_load_bimc_monitor_mask( 
	w_load_bimc_monitor_mask), .w_load_bimc_ecc_uncorrectable_error_cnt( 
	w_load_bimc_ecc_uncorrectable_error_cnt), 
	.w_load_bimc_ecc_correctable_error_cnt( 
	w_load_bimc_ecc_correctable_error_cnt), 
	.w_load_bimc_parity_error_cnt( w_load_bimc_parity_error_cnt), 
	.w_load_bimc_global_config( w_load_bimc_global_config), 
	.w_load_bimc_eccpar_debug( w_load_bimc_eccpar_debug), 
	.w_load_bimc_cmd2( w_load_bimc_cmd2), .w_load_bimc_cmd1( 
	w_load_bimc_cmd1), .w_load_bimc_cmd0( w_load_bimc_cmd0), 
	.w_load_bimc_rxcmd2( w_load_bimc_rxcmd2), .w_load_bimc_rxrsp2( 
	w_load_bimc_rxrsp2), .w_load_bimc_pollrsp2( w_load_bimc_pollrsp2), 
	.w_load_bimc_dbgcmd2( w_load_bimc_dbgcmd2), .w_load_im_consumed( 
	w_load_im_consumed), .w_load_tready_override( 
	w_load_tready_override), .w_load_regs_sa_ctrl( w_load_regs_sa_ctrl), 
	.w_load_sa_snapshot_ia_wdata_part0( 
	w_load_sa_snapshot_ia_wdata_part0), 
	.w_load_sa_snapshot_ia_wdata_part1( 
	w_load_sa_snapshot_ia_wdata_part1), .w_load_sa_snapshot_ia_config( 
	w_load_sa_snapshot_ia_config), .w_load_sa_count_ia_wdata_part0( 
	w_load_sa_count_ia_wdata_part0), .w_load_sa_count_ia_wdata_part1( 
	w_load_sa_count_ia_wdata_part1), .w_load_sa_count_ia_config( 
	w_load_sa_count_ia_config), .w_load_cceip_encrypt_kop_fifo_override( 
	w_load_cceip_encrypt_kop_fifo_override), 
	.w_load_cceip_validate_kop_fifo_override( 
	w_load_cceip_validate_kop_fifo_override), 
	.w_load_cddip_decrypt_kop_fifo_override( 
	w_load_cddip_decrypt_kop_fifo_override), .w_load_sa_global_ctrl( 
	w_load_sa_global_ctrl), .w_load_sa_ctrl_ia_wdata_part0( 
	w_load_sa_ctrl_ia_wdata_part0), .w_load_sa_ctrl_ia_config( 
	w_load_sa_ctrl_ia_config), .w_load_kdf_test_key_size_config( 
	w_load_kdf_test_key_size_config), .f32_data( 
	_zy_simnet_f32_data_3_w$[0:31]));
ixc_assign_32 _zz_strnp_8 ( _zy_simnet_f32_data_3_w$[0:31], f32_data[31:0]);
ixc_assign_11 _zz_strnp_7 ( _zy_simnet_o_reg_addr_2_w$[0:10], 
	o_reg_addr[10:0]);
ixc_assign _zz_strnp_6 ( _zy_simnet_o_reg_read_1_w$, o_reg_read);
ixc_assign _zz_strnp_5 ( _zy_simnet_o_reg_written_0_w$, o_reg_written);
Q_NR02 U8 ( .A0(n122), .A1(n434), .Z(w_load_kdf_test_key_size_config));
Q_OR03 U9 ( .A0(n238), .A1(n230), .A2(n421), .Z(n434));
Q_NR02 U10 ( .A0(n122), .A1(n433), .Z(w_load_sa_ctrl_ia_config));
Q_OR03 U11 ( .A0(n238), .A1(n226), .A2(n421), .Z(n433));
Q_NR02 U12 ( .A0(n122), .A1(n432), .Z(w_load_sa_ctrl_ia_wdata_part0));
Q_OR03 U13 ( .A0(n238), .A1(n235), .A2(n421), .Z(n432));
Q_NR02 U14 ( .A0(n122), .A1(n431), .Z(w_load_sa_global_ctrl));
Q_OR03 U15 ( .A0(n238), .A1(n239), .A2(n421), .Z(n431));
Q_NR02 U16 ( .A0(n122), .A1(n430), .Z(w_load_cddip_decrypt_kop_fifo_override));
Q_OR03 U17 ( .A0(n238), .A1(n233), .A2(n421), .Z(n430));
Q_NR02 U18 ( .A0(n122), .A1(n429), .Z(w_load_cceip_validate_kop_fifo_override));
Q_OR03 U19 ( .A0(n232), .A1(n230), .A2(n421), .Z(n429));
Q_NR02 U20 ( .A0(n122), .A1(n428), .Z(w_load_cceip_encrypt_kop_fifo_override));
Q_OR03 U21 ( .A0(n232), .A1(n228), .A2(n421), .Z(n428));
Q_NR02 U22 ( .A0(n122), .A1(n427), .Z(w_load_sa_count_ia_config));
Q_OR03 U23 ( .A0(n232), .A1(n223), .A2(n421), .Z(n427));
Q_NR02 U24 ( .A0(n122), .A1(n426), .Z(w_load_sa_count_ia_wdata_part1));
Q_OR03 U25 ( .A0(n232), .A1(n239), .A2(n421), .Z(n426));
Q_NR02 U26 ( .A0(n122), .A1(n425), .Z(w_load_sa_count_ia_wdata_part0));
Q_OR03 U27 ( .A0(n232), .A1(n233), .A2(n421), .Z(n425));
Q_NR02 U28 ( .A0(n122), .A1(n424), .Z(w_load_sa_snapshot_ia_config));
Q_OR03 U29 ( .A0(n222), .A1(n242), .A2(n421), .Z(n424));
Q_NR02 U30 ( .A0(n122), .A1(n423), .Z(w_load_sa_snapshot_ia_wdata_part1));
Q_OR03 U31 ( .A0(n222), .A1(n223), .A2(n421), .Z(n423));
Q_NR02 U32 ( .A0(n122), .A1(n422), .Z(w_load_sa_snapshot_ia_wdata_part0));
Q_OR03 U33 ( .A0(n222), .A1(n239), .A2(n421), .Z(n422));
Q_OR03 U34 ( .A0(ws_addr[1]), .A1(ws_addr[0]), .A2(n420), .Z(n421));
Q_OR03 U35 ( .A0(n7), .A1(ws_addr[9]), .A2(ws_addr[8]), .Z(n420));
Q_AN02 U36 ( .A0(w_do_write), .A1(n419), .Z(w_load_regs_sa_ctrl));
Q_NR03 U37 ( .A0(n266), .A1(n228), .A2(n370), .Z(n419));
Q_AN02 U38 ( .A0(w_do_write), .A1(n418), .Z(w_load_tready_override));
Q_NR03 U39 ( .A0(n266), .A1(n226), .A2(n370), .Z(n418));
Q_AN02 U40 ( .A0(w_do_write), .A1(n417), .Z(w_load_im_consumed));
Q_NR03 U41 ( .A0(n266), .A1(n235), .A2(n370), .Z(n417));
Q_AN02 U42 ( .A0(w_do_write), .A1(n416), .Z(w_load_bimc_dbgcmd2));
Q_NR03 U43 ( .A0(n260), .A1(n230), .A2(n370), .Z(n416));
Q_NR02 U44 ( .A0(n122), .A1(n415), .Z(w_load_bimc_pollrsp2));
Q_OR03 U45 ( .A0(n260), .A1(n235), .A2(n370), .Z(n415));
Q_NR02 U46 ( .A0(n122), .A1(n414), .Z(w_load_bimc_rxrsp2));
Q_OR03 U47 ( .A0(n260), .A1(n239), .A2(n370), .Z(n414));
Q_AN02 U48 ( .A0(w_do_write), .A1(n413), .Z(w_load_bimc_rxcmd2));
Q_NR03 U49 ( .A0(n255), .A1(n228), .A2(n370), .Z(n413));
Q_AN02 U50 ( .A0(w_do_write), .A1(n412), .Z(w_load_bimc_cmd0));
Q_NR03 U51 ( .A0(n255), .A1(n226), .A2(n370), .Z(n412));
Q_NR02 U52 ( .A0(n122), .A1(n411), .Z(w_load_bimc_cmd1));
Q_OR03 U53 ( .A0(n255), .A1(n235), .A2(n370), .Z(n411));
Q_AN02 U54 ( .A0(w_do_write), .A1(n410), .Z(w_load_bimc_cmd2));
Q_NR03 U55 ( .A0(n255), .A1(n242), .A2(n370), .Z(n410));
Q_NR02 U56 ( .A0(n122), .A1(n409), .Z(w_load_bimc_eccpar_debug));
Q_OR03 U57 ( .A0(n255), .A1(n223), .A2(n370), .Z(n409));
Q_NR02 U58 ( .A0(n122), .A1(n408), .Z(w_load_bimc_global_config));
Q_OR03 U59 ( .A0(n255), .A1(n233), .A2(n370), .Z(n408));
Q_AN02 U60 ( .A0(w_do_write), .A1(n407), .Z(w_load_bimc_parity_error_cnt));
Q_NR03 U61 ( .A0(n251), .A1(n230), .A2(n370), .Z(n407));
Q_NR02 U62 ( .A0(n122), .A1(n406), .Z(w_load_bimc_ecc_correctable_error_cnt));
Q_OR03 U63 ( .A0(n251), .A1(n228), .A2(n370), .Z(n406));
Q_NR02 U64 ( .A0(n122), .A1(n405), .Z(w_load_bimc_ecc_uncorrectable_error_cnt));
Q_OR03 U65 ( .A0(n251), .A1(n226), .A2(n370), .Z(n405));
Q_NR02 U66 ( .A0(n122), .A1(n404), .Z(w_load_bimc_monitor_mask));
Q_OR03 U67 ( .A0(n251), .A1(n235), .A2(n370), .Z(n404));
Q_NR02 U68 ( .A0(n122), .A1(n403), .Z(w_load_engine_sticky_status));
Q_OR03 U69 ( .A0(n251), .A1(n239), .A2(n370), .Z(n403));
Q_NR02 U70 ( .A0(n122), .A1(n402), .Z(w_load_interrupt_mask));
Q_OR03 U71 ( .A0(n251), .A1(n233), .A2(n370), .Z(n402));
Q_AN02 U72 ( .A0(w_do_write), .A1(n401), .Z(w_load_interrupt_status));
Q_NR03 U73 ( .A0(n245), .A1(n230), .A2(n370), .Z(n401));
Q_AN02 U74 ( .A0(w_do_write), .A1(n400), .Z(w_load_kdf_drbg_seed_1_reseed_interval_1));
Q_NR03 U75 ( .A0(n245), .A1(n228), .A2(n370), .Z(n400));
Q_AN02 U76 ( .A0(w_do_write), .A1(n399), .Z(w_load_kdf_drbg_seed_1_reseed_interval_0));
Q_NR03 U77 ( .A0(n245), .A1(n226), .A2(n370), .Z(n399));
Q_NR02 U78 ( .A0(n122), .A1(n398), .Z(w_load_kdf_drbg_seed_1_state_value_127_96));
Q_OR03 U79 ( .A0(n245), .A1(n235), .A2(n370), .Z(n398));
Q_AN02 U80 ( .A0(w_do_write), .A1(n397), .Z(w_load_kdf_drbg_seed_1_state_value_95_64));
Q_NR03 U81 ( .A0(n245), .A1(n242), .A2(n370), .Z(n397));
Q_NR02 U82 ( .A0(n122), .A1(n396), .Z(w_load_kdf_drbg_seed_1_state_value_63_32));
Q_OR03 U83 ( .A0(n245), .A1(n223), .A2(n370), .Z(n396));
Q_NR02 U84 ( .A0(n122), .A1(n395), .Z(w_load_kdf_drbg_seed_1_state_value_31_0));
Q_OR03 U85 ( .A0(n245), .A1(n239), .A2(n370), .Z(n395));
Q_NR02 U86 ( .A0(n122), .A1(n394), .Z(w_load_kdf_drbg_seed_1_state_key_255_224));
Q_OR03 U87 ( .A0(n245), .A1(n233), .A2(n370), .Z(n394));
Q_AN02 U88 ( .A0(w_do_write), .A1(n393), .Z(w_load_kdf_drbg_seed_1_state_key_223_192));
Q_NR03 U89 ( .A0(n238), .A1(n230), .A2(n370), .Z(n393));
Q_NR02 U90 ( .A0(n122), .A1(n392), .Z(w_load_kdf_drbg_seed_1_state_key_191_160));
Q_OR03 U91 ( .A0(n238), .A1(n228), .A2(n370), .Z(n392));
Q_NR02 U92 ( .A0(n122), .A1(n391), .Z(w_load_kdf_drbg_seed_1_state_key_159_128));
Q_OR03 U93 ( .A0(n238), .A1(n226), .A2(n370), .Z(n391));
Q_NR02 U94 ( .A0(n122), .A1(n390), .Z(w_load_kdf_drbg_seed_1_state_key_127_96));
Q_OR03 U95 ( .A0(n238), .A1(n235), .A2(n370), .Z(n390));
Q_NR02 U96 ( .A0(n122), .A1(n389), .Z(w_load_kdf_drbg_seed_1_state_key_95_64));
Q_OR03 U97 ( .A0(n238), .A1(n242), .A2(n370), .Z(n389));
Q_NR02 U98 ( .A0(n122), .A1(n388), .Z(w_load_kdf_drbg_seed_1_state_key_63_32));
Q_OR03 U99 ( .A0(n238), .A1(n223), .A2(n370), .Z(n388));
Q_NR02 U100 ( .A0(n122), .A1(n387), .Z(w_load_kdf_drbg_seed_1_state_key_31_0));
Q_OR03 U101 ( .A0(n238), .A1(n239), .A2(n370), .Z(n387));
Q_NR02 U102 ( .A0(n122), .A1(n386), .Z(w_load_kdf_drbg_seed_0_reseed_interval_1));
Q_OR03 U103 ( .A0(n238), .A1(n233), .A2(n370), .Z(n386));
Q_AN02 U104 ( .A0(w_do_write), .A1(n385), .Z(w_load_kdf_drbg_seed_0_reseed_interval_0));
Q_NR03 U105 ( .A0(n232), .A1(n230), .A2(n370), .Z(n385));
Q_NR02 U106 ( .A0(n122), .A1(n384), .Z(w_load_kdf_drbg_seed_0_state_value_127_96));
Q_OR03 U107 ( .A0(n232), .A1(n228), .A2(n370), .Z(n384));
Q_NR02 U108 ( .A0(n122), .A1(n383), .Z(w_load_kdf_drbg_seed_0_state_value_95_64));
Q_OR03 U109 ( .A0(n232), .A1(n226), .A2(n370), .Z(n383));
Q_NR02 U110 ( .A0(n122), .A1(n382), .Z(w_load_kdf_drbg_seed_0_state_value_63_32));
Q_OR03 U111 ( .A0(n232), .A1(n235), .A2(n370), .Z(n382));
Q_NR02 U112 ( .A0(n122), .A1(n381), .Z(w_load_kdf_drbg_seed_0_state_value_31_0));
Q_OR03 U113 ( .A0(n232), .A1(n242), .A2(n370), .Z(n381));
Q_NR02 U114 ( .A0(n122), .A1(n380), .Z(w_load_kdf_drbg_seed_0_state_key_255_224));
Q_OR03 U115 ( .A0(n232), .A1(n223), .A2(n370), .Z(n380));
Q_NR02 U116 ( .A0(n122), .A1(n379), .Z(w_load_kdf_drbg_seed_0_state_key_223_192));
Q_OR03 U117 ( .A0(n232), .A1(n239), .A2(n370), .Z(n379));
Q_NR02 U118 ( .A0(n122), .A1(n378), .Z(w_load_kdf_drbg_seed_0_state_key_191_160));
Q_OR03 U119 ( .A0(n232), .A1(n233), .A2(n370), .Z(n378));
Q_NR02 U120 ( .A0(n122), .A1(n377), .Z(w_load_kdf_drbg_seed_0_state_key_159_128));
Q_OR03 U121 ( .A0(n222), .A1(n230), .A2(n370), .Z(n377));
Q_NR02 U122 ( .A0(n122), .A1(n376), .Z(w_load_kdf_drbg_seed_0_state_key_127_96));
Q_OR03 U123 ( .A0(n222), .A1(n228), .A2(n370), .Z(n376));
Q_NR02 U124 ( .A0(n122), .A1(n375), .Z(w_load_kdf_drbg_seed_0_state_key_95_64));
Q_OR03 U125 ( .A0(n222), .A1(n226), .A2(n370), .Z(n375));
Q_NR02 U126 ( .A0(n122), .A1(n374), .Z(w_load_kdf_drbg_seed_0_state_key_63_32));
Q_OR03 U127 ( .A0(n222), .A1(n235), .A2(n370), .Z(n374));
Q_NR02 U128 ( .A0(n122), .A1(n373), .Z(w_load_kdf_drbg_seed_0_state_key_31_0));
Q_OR03 U129 ( .A0(n222), .A1(n242), .A2(n370), .Z(n373));
Q_NR02 U130 ( .A0(n122), .A1(n372), .Z(w_load_kdf_drbg_ctrl));
Q_OR03 U131 ( .A0(n222), .A1(n223), .A2(n370), .Z(n372));
Q_NR02 U132 ( .A0(n122), .A1(n371), .Z(w_load_label7_data0));
Q_OR03 U133 ( .A0(n222), .A1(n233), .A2(n370), .Z(n371));
Q_OR03 U134 ( .A0(ws_addr[1]), .A1(ws_addr[0]), .A2(n369), .Z(n370));
Q_OR03 U135 ( .A0(ws_addr[10]), .A1(n8), .A2(n9), .Z(n369));
Q_AN02 U136 ( .A0(w_do_write), .A1(n368), .Z(w_load_label7_data1));
Q_NR03 U137 ( .A0(n266), .A1(n230), .A2(n310), .Z(n368));
Q_AN02 U138 ( .A0(w_do_write), .A1(n367), .Z(w_load_label7_data2));
Q_NR03 U139 ( .A0(n266), .A1(n228), .A2(n310), .Z(n367));
Q_AN02 U140 ( .A0(w_do_write), .A1(n366), .Z(w_load_label7_data3));
Q_NR03 U141 ( .A0(n266), .A1(n226), .A2(n310), .Z(n366));
Q_NR02 U142 ( .A0(n122), .A1(n365), .Z(w_load_label7_data4));
Q_OR03 U143 ( .A0(n266), .A1(n235), .A2(n310), .Z(n365));
Q_AN02 U144 ( .A0(w_do_write), .A1(n364), .Z(w_load_label7_data5));
Q_NR03 U145 ( .A0(n266), .A1(n242), .A2(n310), .Z(n364));
Q_NR02 U146 ( .A0(n122), .A1(n363), .Z(w_load_label7_data6));
Q_OR03 U147 ( .A0(n266), .A1(n223), .A2(n310), .Z(n363));
Q_NR02 U148 ( .A0(n122), .A1(n362), .Z(w_load_label7_data7));
Q_OR03 U149 ( .A0(n266), .A1(n239), .A2(n310), .Z(n362));
Q_NR02 U150 ( .A0(n122), .A1(n361), .Z(w_load_label7_config));
Q_OR03 U151 ( .A0(n266), .A1(n233), .A2(n310), .Z(n361));
Q_NR02 U152 ( .A0(n122), .A1(n360), .Z(w_load_label6_data0));
Q_OR03 U153 ( .A0(n260), .A1(n228), .A2(n310), .Z(n360));
Q_NR02 U154 ( .A0(n122), .A1(n359), .Z(w_load_label6_data1));
Q_OR03 U155 ( .A0(n260), .A1(n226), .A2(n310), .Z(n359));
Q_NR02 U156 ( .A0(n122), .A1(n358), .Z(w_load_label6_data2));
Q_OR03 U157 ( .A0(n260), .A1(n235), .A2(n310), .Z(n358));
Q_NR02 U158 ( .A0(n122), .A1(n357), .Z(w_load_label6_data3));
Q_OR03 U159 ( .A0(n260), .A1(n242), .A2(n310), .Z(n357));
Q_NR02 U160 ( .A0(n122), .A1(n356), .Z(w_load_label6_data4));
Q_OR03 U161 ( .A0(n260), .A1(n223), .A2(n310), .Z(n356));
Q_NR02 U162 ( .A0(n122), .A1(n355), .Z(w_load_label6_data5));
Q_OR03 U163 ( .A0(n260), .A1(n239), .A2(n310), .Z(n355));
Q_NR02 U164 ( .A0(n122), .A1(n354), .Z(w_load_label6_data6));
Q_OR03 U165 ( .A0(n260), .A1(n233), .A2(n310), .Z(n354));
Q_AN02 U166 ( .A0(w_do_write), .A1(n353), .Z(w_load_label6_data7));
Q_NR03 U167 ( .A0(n255), .A1(n230), .A2(n310), .Z(n353));
Q_NR02 U168 ( .A0(n122), .A1(n352), .Z(w_load_label6_config));
Q_OR03 U169 ( .A0(n255), .A1(n228), .A2(n310), .Z(n352));
Q_NR02 U170 ( .A0(n122), .A1(n351), .Z(w_load_label5_data0));
Q_OR03 U171 ( .A0(n255), .A1(n235), .A2(n310), .Z(n351));
Q_NR02 U172 ( .A0(n122), .A1(n350), .Z(w_load_label5_data1));
Q_OR03 U173 ( .A0(n255), .A1(n242), .A2(n310), .Z(n350));
Q_NR02 U174 ( .A0(n122), .A1(n349), .Z(w_load_label5_data2));
Q_OR03 U175 ( .A0(n255), .A1(n223), .A2(n310), .Z(n349));
Q_NR02 U176 ( .A0(n122), .A1(n348), .Z(w_load_label5_data3));
Q_OR03 U177 ( .A0(n255), .A1(n239), .A2(n310), .Z(n348));
Q_NR02 U178 ( .A0(n122), .A1(n347), .Z(w_load_label5_data4));
Q_OR03 U179 ( .A0(n255), .A1(n233), .A2(n310), .Z(n347));
Q_NR02 U180 ( .A0(n122), .A1(n346), .Z(w_load_label5_data5));
Q_OR03 U181 ( .A0(n251), .A1(n230), .A2(n310), .Z(n346));
Q_NR02 U182 ( .A0(n122), .A1(n345), .Z(w_load_label5_data6));
Q_OR03 U183 ( .A0(n251), .A1(n228), .A2(n310), .Z(n345));
Q_NR02 U184 ( .A0(n122), .A1(n344), .Z(w_load_label5_data7));
Q_OR03 U185 ( .A0(n251), .A1(n226), .A2(n310), .Z(n344));
Q_NR02 U186 ( .A0(n122), .A1(n343), .Z(w_load_label5_config));
Q_OR03 U187 ( .A0(n251), .A1(n235), .A2(n310), .Z(n343));
Q_NR02 U188 ( .A0(n122), .A1(n342), .Z(w_load_label4_data0));
Q_OR03 U189 ( .A0(n251), .A1(n223), .A2(n310), .Z(n342));
Q_NR02 U190 ( .A0(n122), .A1(n341), .Z(w_load_label4_data1));
Q_OR03 U191 ( .A0(n251), .A1(n239), .A2(n310), .Z(n341));
Q_NR02 U192 ( .A0(n122), .A1(n340), .Z(w_load_label4_data2));
Q_OR03 U193 ( .A0(n251), .A1(n233), .A2(n310), .Z(n340));
Q_AN02 U194 ( .A0(w_do_write), .A1(n339), .Z(w_load_label4_data3));
Q_NR03 U195 ( .A0(n245), .A1(n230), .A2(n310), .Z(n339));
Q_NR02 U196 ( .A0(n122), .A1(n338), .Z(w_load_label4_data4));
Q_OR03 U197 ( .A0(n245), .A1(n228), .A2(n310), .Z(n338));
Q_NR02 U198 ( .A0(n122), .A1(n337), .Z(w_load_label4_data5));
Q_OR03 U199 ( .A0(n245), .A1(n226), .A2(n310), .Z(n337));
Q_NR02 U200 ( .A0(n122), .A1(n336), .Z(w_load_label4_data6));
Q_OR03 U201 ( .A0(n245), .A1(n235), .A2(n310), .Z(n336));
Q_NR02 U202 ( .A0(n122), .A1(n335), .Z(w_load_label4_data7));
Q_OR03 U203 ( .A0(n245), .A1(n242), .A2(n310), .Z(n335));
Q_NR02 U204 ( .A0(n122), .A1(n334), .Z(w_load_label4_config));
Q_OR03 U205 ( .A0(n245), .A1(n223), .A2(n310), .Z(n334));
Q_NR02 U206 ( .A0(n122), .A1(n333), .Z(w_load_label3_data0));
Q_OR03 U207 ( .A0(n245), .A1(n233), .A2(n310), .Z(n333));
Q_NR02 U208 ( .A0(n122), .A1(n332), .Z(w_load_label3_data1));
Q_OR03 U209 ( .A0(n238), .A1(n230), .A2(n310), .Z(n332));
Q_NR02 U210 ( .A0(n122), .A1(n331), .Z(w_load_label3_data2));
Q_OR03 U211 ( .A0(n238), .A1(n228), .A2(n310), .Z(n331));
Q_NR02 U212 ( .A0(n122), .A1(n330), .Z(w_load_label3_data3));
Q_OR03 U213 ( .A0(n238), .A1(n226), .A2(n310), .Z(n330));
Q_NR02 U214 ( .A0(n122), .A1(n329), .Z(w_load_label3_data4));
Q_OR03 U215 ( .A0(n238), .A1(n235), .A2(n310), .Z(n329));
Q_NR02 U216 ( .A0(n122), .A1(n328), .Z(w_load_label3_data5));
Q_OR03 U217 ( .A0(n238), .A1(n242), .A2(n310), .Z(n328));
Q_NR02 U218 ( .A0(n122), .A1(n327), .Z(w_load_label3_data6));
Q_OR03 U219 ( .A0(n238), .A1(n223), .A2(n310), .Z(n327));
Q_NR02 U220 ( .A0(n122), .A1(n326), .Z(w_load_label3_data7));
Q_OR03 U221 ( .A0(n238), .A1(n239), .A2(n310), .Z(n326));
Q_NR02 U222 ( .A0(n122), .A1(n325), .Z(w_load_label3_config));
Q_OR03 U223 ( .A0(n238), .A1(n233), .A2(n310), .Z(n325));
Q_NR02 U224 ( .A0(n122), .A1(n324), .Z(w_load_label2_data0));
Q_OR03 U225 ( .A0(n232), .A1(n228), .A2(n310), .Z(n324));
Q_NR02 U226 ( .A0(n122), .A1(n323), .Z(w_load_label2_data1));
Q_OR03 U227 ( .A0(n232), .A1(n226), .A2(n310), .Z(n323));
Q_NR02 U228 ( .A0(n122), .A1(n322), .Z(w_load_label2_data2));
Q_OR03 U229 ( .A0(n232), .A1(n235), .A2(n310), .Z(n322));
Q_NR02 U230 ( .A0(n122), .A1(n321), .Z(w_load_label2_data3));
Q_OR03 U231 ( .A0(n232), .A1(n242), .A2(n310), .Z(n321));
Q_NR02 U232 ( .A0(n122), .A1(n320), .Z(w_load_label2_data4));
Q_OR03 U233 ( .A0(n232), .A1(n223), .A2(n310), .Z(n320));
Q_NR02 U234 ( .A0(n122), .A1(n319), .Z(w_load_label2_data5));
Q_OR03 U235 ( .A0(n232), .A1(n239), .A2(n310), .Z(n319));
Q_NR02 U236 ( .A0(n122), .A1(n318), .Z(w_load_label2_data6));
Q_OR03 U237 ( .A0(n232), .A1(n233), .A2(n310), .Z(n318));
Q_NR02 U238 ( .A0(n122), .A1(n317), .Z(w_load_label2_data7));
Q_OR03 U239 ( .A0(n222), .A1(n230), .A2(n310), .Z(n317));
Q_NR02 U240 ( .A0(n122), .A1(n316), .Z(w_load_label2_config));
Q_OR03 U241 ( .A0(n222), .A1(n228), .A2(n310), .Z(n316));
Q_NR02 U242 ( .A0(n122), .A1(n315), .Z(w_load_label1_data0));
Q_OR03 U243 ( .A0(n222), .A1(n235), .A2(n310), .Z(n315));
Q_NR02 U244 ( .A0(n122), .A1(n314), .Z(w_load_label1_data1));
Q_OR03 U245 ( .A0(n222), .A1(n242), .A2(n310), .Z(n314));
Q_NR02 U246 ( .A0(n122), .A1(n313), .Z(w_load_label1_data2));
Q_OR03 U247 ( .A0(n222), .A1(n223), .A2(n310), .Z(n313));
Q_NR02 U248 ( .A0(n122), .A1(n312), .Z(w_load_label1_data3));
Q_OR03 U249 ( .A0(n222), .A1(n239), .A2(n310), .Z(n312));
Q_NR02 U250 ( .A0(n122), .A1(n311), .Z(w_load_label1_data4));
Q_OR03 U251 ( .A0(n222), .A1(n233), .A2(n310), .Z(n311));
Q_OR03 U252 ( .A0(ws_addr[1]), .A1(ws_addr[0]), .A2(n309), .Z(n310));
Q_OR03 U253 ( .A0(ws_addr[10]), .A1(n8), .A2(ws_addr[8]), .Z(n309));
Q_AN02 U254 ( .A0(w_do_write), .A1(n308), .Z(w_load_label1_data5));
Q_NR03 U255 ( .A0(n266), .A1(n230), .A2(n271), .Z(n308));
Q_AN02 U256 ( .A0(w_do_write), .A1(n307), .Z(w_load_label1_data6));
Q_NR03 U257 ( .A0(n266), .A1(n228), .A2(n271), .Z(n307));
Q_AN02 U258 ( .A0(w_do_write), .A1(n306), .Z(w_load_label1_data7));
Q_NR03 U259 ( .A0(n266), .A1(n226), .A2(n271), .Z(n306));
Q_NR02 U260 ( .A0(n122), .A1(n305), .Z(w_load_label1_config));
Q_OR03 U261 ( .A0(n266), .A1(n235), .A2(n271), .Z(n305));
Q_NR02 U262 ( .A0(n122), .A1(n304), .Z(w_load_label0_data0));
Q_OR03 U263 ( .A0(n266), .A1(n223), .A2(n271), .Z(n304));
Q_NR02 U264 ( .A0(n122), .A1(n303), .Z(w_load_label0_data1));
Q_OR03 U265 ( .A0(n266), .A1(n239), .A2(n271), .Z(n303));
Q_NR02 U266 ( .A0(n122), .A1(n302), .Z(w_load_label0_data2));
Q_OR03 U267 ( .A0(n266), .A1(n233), .A2(n271), .Z(n302));
Q_AN02 U268 ( .A0(w_do_write), .A1(n301), .Z(w_load_label0_data3));
Q_NR03 U269 ( .A0(n260), .A1(n230), .A2(n271), .Z(n301));
Q_NR02 U270 ( .A0(n122), .A1(n300), .Z(w_load_label0_data4));
Q_OR03 U271 ( .A0(n260), .A1(n228), .A2(n271), .Z(n300));
Q_NR02 U272 ( .A0(n122), .A1(n299), .Z(w_load_label0_data5));
Q_OR03 U273 ( .A0(n260), .A1(n226), .A2(n271), .Z(n299));
Q_NR02 U274 ( .A0(n122), .A1(n298), .Z(w_load_label0_data6));
Q_OR03 U275 ( .A0(n260), .A1(n235), .A2(n271), .Z(n298));
Q_NR02 U276 ( .A0(n122), .A1(n297), .Z(w_load_label0_data7));
Q_OR03 U277 ( .A0(n260), .A1(n242), .A2(n271), .Z(n297));
Q_NR02 U278 ( .A0(n122), .A1(n296), .Z(w_load_label0_config));
Q_OR03 U279 ( .A0(n260), .A1(n223), .A2(n271), .Z(n296));
Q_NR02 U280 ( .A0(n122), .A1(n295), .Z(w_load_kim_ia_config));
Q_OR03 U281 ( .A0(n255), .A1(n228), .A2(n271), .Z(n295));
Q_NR02 U282 ( .A0(n122), .A1(n294), .Z(w_load_kim_ia_wdata_part1));
Q_OR03 U283 ( .A0(n255), .A1(n226), .A2(n271), .Z(n294));
Q_NR02 U284 ( .A0(n122), .A1(n293), .Z(w_load_kim_ia_wdata_part0));
Q_OR03 U285 ( .A0(n255), .A1(n235), .A2(n271), .Z(n293));
Q_NR02 U286 ( .A0(n122), .A1(n292), .Z(w_load_ckv_ia_config));
Q_OR03 U287 ( .A0(n251), .A1(n230), .A2(n271), .Z(n292));
Q_NR02 U288 ( .A0(n122), .A1(n291), .Z(w_load_ckv_ia_wdata_part1));
Q_OR03 U289 ( .A0(n251), .A1(n228), .A2(n271), .Z(n291));
Q_NR02 U290 ( .A0(n122), .A1(n290), .Z(w_load_ckv_ia_wdata_part0));
Q_OR03 U291 ( .A0(n251), .A1(n226), .A2(n271), .Z(n290));
Q_NR02 U292 ( .A0(n122), .A1(n289), .Z(w_load_cddip3_out_im_read_done));
Q_OR03 U293 ( .A0(n251), .A1(n223), .A2(n271), .Z(n289));
Q_NR02 U294 ( .A0(n122), .A1(n288), .Z(w_load_cddip3_out_im_config));
Q_OR03 U295 ( .A0(n251), .A1(n233), .A2(n271), .Z(n288));
Q_NR02 U296 ( .A0(n122), .A1(n287), .Z(w_load_cddip3_out_ia_config));
Q_OR03 U297 ( .A0(n245), .A1(n235), .A2(n271), .Z(n287));
Q_NR02 U298 ( .A0(n122), .A1(n286), .Z(w_load_cddip3_out_ia_wdata_part2));
Q_OR03 U299 ( .A0(n245), .A1(n242), .A2(n271), .Z(n286));
Q_NR02 U300 ( .A0(n122), .A1(n285), .Z(w_load_cddip3_out_ia_wdata_part1));
Q_OR03 U301 ( .A0(n245), .A1(n223), .A2(n271), .Z(n285));
Q_NR02 U302 ( .A0(n122), .A1(n284), .Z(w_load_cddip3_out_ia_wdata_part0));
Q_OR03 U303 ( .A0(n245), .A1(n239), .A2(n271), .Z(n284));
Q_NR02 U304 ( .A0(n122), .A1(n283), .Z(w_load_cddip2_out_im_read_done));
Q_OR03 U305 ( .A0(n238), .A1(n228), .A2(n271), .Z(n283));
Q_NR02 U306 ( .A0(n122), .A1(n282), .Z(w_load_cddip2_out_im_config));
Q_OR03 U307 ( .A0(n238), .A1(n235), .A2(n271), .Z(n282));
Q_NR02 U308 ( .A0(n122), .A1(n281), .Z(w_load_cddip2_out_ia_config));
Q_OR03 U309 ( .A0(n238), .A1(n233), .A2(n271), .Z(n281));
Q_NR02 U310 ( .A0(n122), .A1(n280), .Z(w_load_cddip2_out_ia_wdata_part2));
Q_OR03 U311 ( .A0(n232), .A1(n230), .A2(n271), .Z(n280));
Q_NR02 U312 ( .A0(n122), .A1(n279), .Z(w_load_cddip2_out_ia_wdata_part1));
Q_OR03 U313 ( .A0(n232), .A1(n228), .A2(n271), .Z(n279));
Q_NR02 U314 ( .A0(n122), .A1(n278), .Z(w_load_cddip2_out_ia_wdata_part0));
Q_OR03 U315 ( .A0(n232), .A1(n226), .A2(n271), .Z(n278));
Q_NR02 U316 ( .A0(n122), .A1(n277), .Z(w_load_cddip1_out_im_read_done));
Q_OR03 U317 ( .A0(n232), .A1(n223), .A2(n271), .Z(n277));
Q_NR02 U318 ( .A0(n122), .A1(n276), .Z(w_load_cddip1_out_im_config));
Q_OR03 U319 ( .A0(n232), .A1(n233), .A2(n271), .Z(n276));
Q_NR02 U320 ( .A0(n122), .A1(n275), .Z(w_load_cddip1_out_ia_config));
Q_OR03 U321 ( .A0(n222), .A1(n235), .A2(n271), .Z(n275));
Q_NR02 U322 ( .A0(n122), .A1(n274), .Z(w_load_cddip1_out_ia_wdata_part2));
Q_OR03 U323 ( .A0(n222), .A1(n242), .A2(n271), .Z(n274));
Q_NR02 U324 ( .A0(n122), .A1(n273), .Z(w_load_cddip1_out_ia_wdata_part1));
Q_OR03 U325 ( .A0(n222), .A1(n223), .A2(n271), .Z(n273));
Q_NR02 U326 ( .A0(n122), .A1(n272), .Z(w_load_cddip1_out_ia_wdata_part0));
Q_OR03 U327 ( .A0(n222), .A1(n239), .A2(n271), .Z(n272));
Q_OR03 U328 ( .A0(ws_addr[1]), .A1(ws_addr[0]), .A2(n270), .Z(n271));
Q_OR03 U329 ( .A0(ws_addr[10]), .A1(ws_addr[9]), .A2(n9), .Z(n270));
Q_NR02 U330 ( .A0(n122), .A1(n269), .Z(w_load_cddip0_out_im_read_done));
Q_OR03 U331 ( .A0(n266), .A1(n228), .A2(n224), .Z(n269));
Q_NR02 U332 ( .A0(n122), .A1(n268), .Z(w_load_cddip0_out_im_config));
Q_OR03 U333 ( .A0(n266), .A1(n235), .A2(n224), .Z(n268));
Q_NR02 U334 ( .A0(n122), .A1(n267), .Z(w_load_cddip0_out_ia_config));
Q_OR03 U335 ( .A0(n266), .A1(n233), .A2(n224), .Z(n267));
Q_ND03 U336 ( .A0(ws_addr[7]), .A1(ws_addr[6]), .A2(ws_addr[5]), .Z(n266));
Q_NR02 U337 ( .A0(n122), .A1(n265), .Z(w_load_cddip0_out_ia_wdata_part2));
Q_OR03 U338 ( .A0(n260), .A1(n230), .A2(n224), .Z(n265));
Q_NR02 U339 ( .A0(n122), .A1(n264), .Z(w_load_cddip0_out_ia_wdata_part1));
Q_OR03 U340 ( .A0(n260), .A1(n228), .A2(n224), .Z(n264));
Q_NR02 U341 ( .A0(n122), .A1(n263), .Z(w_load_cddip0_out_ia_wdata_part0));
Q_OR03 U342 ( .A0(n260), .A1(n226), .A2(n224), .Z(n263));
Q_NR02 U343 ( .A0(n122), .A1(n262), .Z(w_load_cceip3_out_im_read_done));
Q_OR03 U344 ( .A0(n260), .A1(n223), .A2(n224), .Z(n262));
Q_NR02 U345 ( .A0(n122), .A1(n261), .Z(w_load_cceip3_out_im_config));
Q_OR03 U346 ( .A0(n260), .A1(n233), .A2(n224), .Z(n261));
Q_OR03 U347 ( .A0(n10), .A1(n13), .A2(ws_addr[5]), .Z(n260));
Q_NR02 U348 ( .A0(n122), .A1(n259), .Z(w_load_cceip3_out_ia_config));
Q_OR03 U349 ( .A0(n255), .A1(n235), .A2(n224), .Z(n259));
Q_NR02 U350 ( .A0(n122), .A1(n258), .Z(w_load_cceip3_out_ia_wdata_part2));
Q_OR03 U351 ( .A0(n255), .A1(n242), .A2(n224), .Z(n258));
Q_NR02 U352 ( .A0(n122), .A1(n257), .Z(w_load_cceip3_out_ia_wdata_part1));
Q_OR03 U353 ( .A0(n255), .A1(n223), .A2(n224), .Z(n257));
Q_NR02 U354 ( .A0(n122), .A1(n256), .Z(w_load_cceip3_out_ia_wdata_part0));
Q_OR03 U355 ( .A0(n255), .A1(n239), .A2(n224), .Z(n256));
Q_OR03 U356 ( .A0(n10), .A1(ws_addr[6]), .A2(n14), .Z(n255));
Q_NR02 U357 ( .A0(n122), .A1(n254), .Z(w_load_cceip2_out_im_read_done));
Q_OR03 U358 ( .A0(n251), .A1(n228), .A2(n224), .Z(n254));
Q_NR02 U359 ( .A0(n122), .A1(n253), .Z(w_load_cceip2_out_im_config));
Q_OR03 U360 ( .A0(n251), .A1(n235), .A2(n224), .Z(n253));
Q_NR02 U361 ( .A0(n122), .A1(n252), .Z(w_load_cceip2_out_ia_config));
Q_OR03 U362 ( .A0(n251), .A1(n233), .A2(n224), .Z(n252));
Q_OR03 U363 ( .A0(n10), .A1(ws_addr[6]), .A2(ws_addr[5]), .Z(n251));
Q_NR02 U364 ( .A0(n122), .A1(n250), .Z(w_load_cceip2_out_ia_wdata_part2));
Q_OR03 U365 ( .A0(n245), .A1(n230), .A2(n224), .Z(n250));
Q_NR02 U366 ( .A0(n122), .A1(n249), .Z(w_load_cceip2_out_ia_wdata_part1));
Q_OR03 U367 ( .A0(n245), .A1(n228), .A2(n224), .Z(n249));
Q_NR02 U368 ( .A0(n122), .A1(n248), .Z(w_load_cceip2_out_ia_wdata_part0));
Q_OR03 U369 ( .A0(n245), .A1(n226), .A2(n224), .Z(n248));
Q_NR02 U370 ( .A0(n122), .A1(n247), .Z(w_load_cceip1_out_im_read_done));
Q_OR03 U371 ( .A0(n245), .A1(n223), .A2(n224), .Z(n247));
Q_NR02 U372 ( .A0(n122), .A1(n246), .Z(w_load_cceip1_out_im_config));
Q_OR03 U373 ( .A0(n245), .A1(n233), .A2(n224), .Z(n246));
Q_OR03 U374 ( .A0(ws_addr[7]), .A1(n13), .A2(n14), .Z(n245));
Q_NR02 U375 ( .A0(n122), .A1(n244), .Z(w_load_cceip1_out_ia_config));
Q_OR03 U376 ( .A0(n238), .A1(n235), .A2(n224), .Z(n244));
Q_NR02 U377 ( .A0(n122), .A1(n243), .Z(w_load_cceip1_out_ia_wdata_part2));
Q_OR03 U378 ( .A0(n238), .A1(n242), .A2(n224), .Z(n243));
Q_OR03 U379 ( .A0(ws_addr[4]), .A1(n16), .A2(n19), .Z(n242));
Q_NR02 U380 ( .A0(n122), .A1(n241), .Z(w_load_cceip1_out_ia_wdata_part1));
Q_OR03 U381 ( .A0(n238), .A1(n223), .A2(n224), .Z(n241));
Q_NR02 U382 ( .A0(n122), .A1(n240), .Z(w_load_cceip1_out_ia_wdata_part0));
Q_OR03 U383 ( .A0(n238), .A1(n239), .A2(n224), .Z(n240));
Q_OR03 U384 ( .A0(ws_addr[4]), .A1(ws_addr[3]), .A2(n19), .Z(n239));
Q_OR03 U385 ( .A0(ws_addr[7]), .A1(n13), .A2(ws_addr[5]), .Z(n238));
Q_NR02 U386 ( .A0(n122), .A1(n237), .Z(w_load_cceip0_out_im_read_done));
Q_OR03 U387 ( .A0(n232), .A1(n228), .A2(n224), .Z(n237));
Q_NR02 U388 ( .A0(n122), .A1(n236), .Z(w_load_cceip0_out_im_config));
Q_OR03 U389 ( .A0(n232), .A1(n235), .A2(n224), .Z(n236));
Q_OR03 U390 ( .A0(n15), .A1(ws_addr[3]), .A2(ws_addr[2]), .Z(n235));
Q_NR02 U391 ( .A0(n122), .A1(n234), .Z(w_load_cceip0_out_ia_config));
Q_OR03 U392 ( .A0(n232), .A1(n233), .A2(n224), .Z(n234));
Q_OR03 U393 ( .A0(ws_addr[4]), .A1(ws_addr[3]), .A2(ws_addr[2]), .Z(n233));
Q_OR03 U394 ( .A0(ws_addr[7]), .A1(ws_addr[6]), .A2(n14), .Z(n232));
Q_NR02 U395 ( .A0(n122), .A1(n231), .Z(w_load_cceip0_out_ia_wdata_part2));
Q_OR03 U396 ( .A0(n222), .A1(n230), .A2(n224), .Z(n231));
Q_ND03 U397 ( .A0(ws_addr[4]), .A1(ws_addr[3]), .A2(ws_addr[2]), .Z(n230));
Q_NR02 U398 ( .A0(n122), .A1(n229), .Z(w_load_cceip0_out_ia_wdata_part1));
Q_OR03 U399 ( .A0(n222), .A1(n228), .A2(n224), .Z(n229));
Q_OR03 U400 ( .A0(n15), .A1(n16), .A2(ws_addr[2]), .Z(n228));
Q_NR02 U401 ( .A0(n122), .A1(n227), .Z(w_load_cceip0_out_ia_wdata_part0));
Q_OR03 U402 ( .A0(n222), .A1(n226), .A2(n224), .Z(n227));
Q_OR03 U403 ( .A0(n15), .A1(ws_addr[3]), .A2(n19), .Z(n226));
Q_NR02 U404 ( .A0(n122), .A1(n225), .Z(w_load_spare_config));
Q_OR03 U405 ( .A0(n222), .A1(n223), .A2(n224), .Z(n225));
Q_OR03 U406 ( .A0(ws_addr[1]), .A1(ws_addr[0]), .A2(n221), .Z(n224));
Q_OR03 U407 ( .A0(ws_addr[4]), .A1(n16), .A2(ws_addr[2]), .Z(n223));
Q_OR03 U408 ( .A0(ws_addr[7]), .A1(ws_addr[6]), .A2(ws_addr[5]), .Z(n222));
Q_OR03 U409 ( .A0(ws_addr[10]), .A1(ws_addr[9]), .A2(ws_addr[8]), .Z(n221));
ixc_assign_32 _zz_strnp_4 ( o_reg_wr_data[31:0], f32_data[31:0]);
Q_OR03 U411 ( .A0(n218), .A1(n219), .A2(n220), .Z(r32_formatted_reg_data[31]));
Q_OR03 U412 ( .A0(f32_mux_2_data[31]), .A1(f32_mux_1_data[31]), .A2(f32_mux_0_data[31]), .Z(n220));
Q_OR03 U413 ( .A0(f32_mux_5_data[31]), .A1(f32_mux_4_data[31]), .A2(f32_mux_3_data[31]), .Z(n219));
Q_OR03 U414 ( .A0(f32_mux_8_data[31]), .A1(f32_mux_7_data[31]), .A2(f32_mux_6_data[31]), .Z(n218));
Q_OR03 U415 ( .A0(n215), .A1(n216), .A2(n217), .Z(r32_formatted_reg_data[30]));
Q_OR03 U416 ( .A0(f32_mux_2_data[30]), .A1(f32_mux_1_data[30]), .A2(f32_mux_0_data[30]), .Z(n217));
Q_OR03 U417 ( .A0(f32_mux_5_data[30]), .A1(f32_mux_4_data[30]), .A2(f32_mux_3_data[30]), .Z(n216));
Q_OR03 U418 ( .A0(f32_mux_8_data[30]), .A1(f32_mux_7_data[30]), .A2(f32_mux_6_data[30]), .Z(n215));
Q_OR03 U419 ( .A0(n212), .A1(n213), .A2(n214), .Z(r32_formatted_reg_data[29]));
Q_OR03 U420 ( .A0(f32_mux_2_data[29]), .A1(f32_mux_1_data[29]), .A2(f32_mux_0_data[29]), .Z(n214));
Q_OR03 U421 ( .A0(f32_mux_5_data[29]), .A1(f32_mux_4_data[29]), .A2(f32_mux_3_data[29]), .Z(n213));
Q_OR03 U422 ( .A0(f32_mux_8_data[29]), .A1(f32_mux_7_data[29]), .A2(f32_mux_6_data[29]), .Z(n212));
Q_OR03 U423 ( .A0(n209), .A1(n210), .A2(n211), .Z(r32_formatted_reg_data[28]));
Q_OR03 U424 ( .A0(f32_mux_2_data[28]), .A1(f32_mux_1_data[28]), .A2(f32_mux_0_data[28]), .Z(n211));
Q_OR03 U425 ( .A0(f32_mux_5_data[28]), .A1(f32_mux_4_data[28]), .A2(f32_mux_3_data[28]), .Z(n210));
Q_OR03 U426 ( .A0(f32_mux_8_data[28]), .A1(f32_mux_7_data[28]), .A2(f32_mux_6_data[28]), .Z(n209));
Q_OR03 U427 ( .A0(n206), .A1(n207), .A2(n208), .Z(r32_formatted_reg_data[27]));
Q_OR03 U428 ( .A0(f32_mux_2_data[27]), .A1(f32_mux_1_data[27]), .A2(f32_mux_0_data[27]), .Z(n208));
Q_OR03 U429 ( .A0(f32_mux_5_data[27]), .A1(f32_mux_4_data[27]), .A2(f32_mux_3_data[27]), .Z(n207));
Q_OR03 U430 ( .A0(f32_mux_8_data[27]), .A1(f32_mux_7_data[27]), .A2(f32_mux_6_data[27]), .Z(n206));
Q_OR03 U431 ( .A0(n203), .A1(n204), .A2(n205), .Z(r32_formatted_reg_data[26]));
Q_OR03 U432 ( .A0(f32_mux_2_data[26]), .A1(f32_mux_1_data[26]), .A2(f32_mux_0_data[26]), .Z(n205));
Q_OR03 U433 ( .A0(f32_mux_5_data[26]), .A1(f32_mux_4_data[26]), .A2(f32_mux_3_data[26]), .Z(n204));
Q_OR03 U434 ( .A0(f32_mux_8_data[26]), .A1(f32_mux_7_data[26]), .A2(f32_mux_6_data[26]), .Z(n203));
Q_OR03 U435 ( .A0(n200), .A1(n201), .A2(n202), .Z(r32_formatted_reg_data[25]));
Q_OR03 U436 ( .A0(f32_mux_2_data[25]), .A1(f32_mux_1_data[25]), .A2(f32_mux_0_data[25]), .Z(n202));
Q_OR03 U437 ( .A0(f32_mux_5_data[25]), .A1(f32_mux_4_data[25]), .A2(f32_mux_3_data[25]), .Z(n201));
Q_OR03 U438 ( .A0(f32_mux_8_data[25]), .A1(f32_mux_7_data[25]), .A2(f32_mux_6_data[25]), .Z(n200));
Q_OR03 U439 ( .A0(n197), .A1(n198), .A2(n199), .Z(r32_formatted_reg_data[24]));
Q_OR03 U440 ( .A0(f32_mux_2_data[24]), .A1(f32_mux_1_data[24]), .A2(f32_mux_0_data[24]), .Z(n199));
Q_OR03 U441 ( .A0(f32_mux_5_data[24]), .A1(f32_mux_4_data[24]), .A2(f32_mux_3_data[24]), .Z(n198));
Q_OR03 U442 ( .A0(f32_mux_8_data[24]), .A1(f32_mux_7_data[24]), .A2(f32_mux_6_data[24]), .Z(n197));
Q_OR03 U443 ( .A0(n194), .A1(n195), .A2(n196), .Z(r32_formatted_reg_data[23]));
Q_OR03 U444 ( .A0(f32_mux_2_data[23]), .A1(f32_mux_1_data[23]), .A2(f32_mux_0_data[23]), .Z(n196));
Q_OR03 U445 ( .A0(f32_mux_5_data[23]), .A1(f32_mux_4_data[23]), .A2(f32_mux_3_data[23]), .Z(n195));
Q_OR03 U446 ( .A0(f32_mux_8_data[23]), .A1(f32_mux_7_data[23]), .A2(f32_mux_6_data[23]), .Z(n194));
Q_OR03 U447 ( .A0(n191), .A1(n192), .A2(n193), .Z(r32_formatted_reg_data[22]));
Q_OR03 U448 ( .A0(f32_mux_2_data[22]), .A1(f32_mux_1_data[22]), .A2(f32_mux_0_data[22]), .Z(n193));
Q_OR03 U449 ( .A0(f32_mux_5_data[22]), .A1(f32_mux_4_data[22]), .A2(f32_mux_3_data[22]), .Z(n192));
Q_OR03 U450 ( .A0(f32_mux_8_data[22]), .A1(f32_mux_7_data[22]), .A2(f32_mux_6_data[22]), .Z(n191));
Q_OR03 U451 ( .A0(n188), .A1(n189), .A2(n190), .Z(r32_formatted_reg_data[21]));
Q_OR03 U452 ( .A0(f32_mux_2_data[21]), .A1(f32_mux_1_data[21]), .A2(f32_mux_0_data[21]), .Z(n190));
Q_OR03 U453 ( .A0(f32_mux_5_data[21]), .A1(f32_mux_4_data[21]), .A2(f32_mux_3_data[21]), .Z(n189));
Q_OR03 U454 ( .A0(f32_mux_8_data[21]), .A1(f32_mux_7_data[21]), .A2(f32_mux_6_data[21]), .Z(n188));
Q_OR03 U455 ( .A0(n185), .A1(n186), .A2(n187), .Z(r32_formatted_reg_data[20]));
Q_OR03 U456 ( .A0(f32_mux_2_data[20]), .A1(f32_mux_1_data[20]), .A2(f32_mux_0_data[20]), .Z(n187));
Q_OR03 U457 ( .A0(f32_mux_5_data[20]), .A1(f32_mux_4_data[20]), .A2(f32_mux_3_data[20]), .Z(n186));
Q_OR03 U458 ( .A0(f32_mux_8_data[20]), .A1(f32_mux_7_data[20]), .A2(f32_mux_6_data[20]), .Z(n185));
Q_OR03 U459 ( .A0(n182), .A1(n183), .A2(n184), .Z(r32_formatted_reg_data[19]));
Q_OR03 U460 ( .A0(f32_mux_2_data[19]), .A1(f32_mux_1_data[19]), .A2(f32_mux_0_data[19]), .Z(n184));
Q_OR03 U461 ( .A0(f32_mux_5_data[19]), .A1(f32_mux_4_data[19]), .A2(f32_mux_3_data[19]), .Z(n183));
Q_OR03 U462 ( .A0(f32_mux_8_data[19]), .A1(f32_mux_7_data[19]), .A2(f32_mux_6_data[19]), .Z(n182));
Q_OR03 U463 ( .A0(n179), .A1(n180), .A2(n181), .Z(r32_formatted_reg_data[18]));
Q_OR03 U464 ( .A0(f32_mux_2_data[18]), .A1(f32_mux_1_data[18]), .A2(f32_mux_0_data[18]), .Z(n181));
Q_OR03 U465 ( .A0(f32_mux_5_data[18]), .A1(f32_mux_4_data[18]), .A2(f32_mux_3_data[18]), .Z(n180));
Q_OR03 U466 ( .A0(f32_mux_8_data[18]), .A1(f32_mux_7_data[18]), .A2(f32_mux_6_data[18]), .Z(n179));
Q_OR03 U467 ( .A0(n176), .A1(n177), .A2(n178), .Z(r32_formatted_reg_data[17]));
Q_OR03 U468 ( .A0(f32_mux_2_data[17]), .A1(f32_mux_1_data[17]), .A2(f32_mux_0_data[17]), .Z(n178));
Q_OR03 U469 ( .A0(f32_mux_5_data[17]), .A1(f32_mux_4_data[17]), .A2(f32_mux_3_data[17]), .Z(n177));
Q_OR03 U470 ( .A0(f32_mux_8_data[17]), .A1(f32_mux_7_data[17]), .A2(f32_mux_6_data[17]), .Z(n176));
Q_OR03 U471 ( .A0(n173), .A1(n174), .A2(n175), .Z(r32_formatted_reg_data[16]));
Q_OR03 U472 ( .A0(f32_mux_2_data[16]), .A1(f32_mux_1_data[16]), .A2(f32_mux_0_data[16]), .Z(n175));
Q_OR03 U473 ( .A0(f32_mux_5_data[16]), .A1(f32_mux_4_data[16]), .A2(f32_mux_3_data[16]), .Z(n174));
Q_OR03 U474 ( .A0(f32_mux_8_data[16]), .A1(f32_mux_7_data[16]), .A2(f32_mux_6_data[16]), .Z(n173));
Q_OR03 U475 ( .A0(n170), .A1(n171), .A2(n172), .Z(r32_formatted_reg_data[15]));
Q_OR03 U476 ( .A0(f32_mux_2_data[15]), .A1(f32_mux_1_data[15]), .A2(f32_mux_0_data[15]), .Z(n172));
Q_OR03 U477 ( .A0(f32_mux_5_data[15]), .A1(f32_mux_4_data[15]), .A2(f32_mux_3_data[15]), .Z(n171));
Q_OR03 U478 ( .A0(f32_mux_8_data[15]), .A1(f32_mux_7_data[15]), .A2(f32_mux_6_data[15]), .Z(n170));
Q_OR03 U479 ( .A0(n167), .A1(n168), .A2(n169), .Z(r32_formatted_reg_data[14]));
Q_OR03 U480 ( .A0(f32_mux_2_data[14]), .A1(f32_mux_1_data[14]), .A2(f32_mux_0_data[14]), .Z(n169));
Q_OR03 U481 ( .A0(f32_mux_5_data[14]), .A1(f32_mux_4_data[14]), .A2(f32_mux_3_data[14]), .Z(n168));
Q_OR03 U482 ( .A0(f32_mux_8_data[14]), .A1(f32_mux_7_data[14]), .A2(f32_mux_6_data[14]), .Z(n167));
Q_OR03 U483 ( .A0(n164), .A1(n165), .A2(n166), .Z(r32_formatted_reg_data[13]));
Q_OR03 U484 ( .A0(f32_mux_2_data[13]), .A1(f32_mux_1_data[13]), .A2(f32_mux_0_data[13]), .Z(n166));
Q_OR03 U485 ( .A0(f32_mux_5_data[13]), .A1(f32_mux_4_data[13]), .A2(f32_mux_3_data[13]), .Z(n165));
Q_OR03 U486 ( .A0(f32_mux_8_data[13]), .A1(f32_mux_7_data[13]), .A2(f32_mux_6_data[13]), .Z(n164));
Q_OR03 U487 ( .A0(n161), .A1(n162), .A2(n163), .Z(r32_formatted_reg_data[12]));
Q_OR03 U488 ( .A0(f32_mux_2_data[12]), .A1(f32_mux_1_data[12]), .A2(f32_mux_0_data[12]), .Z(n163));
Q_OR03 U489 ( .A0(f32_mux_5_data[12]), .A1(f32_mux_4_data[12]), .A2(f32_mux_3_data[12]), .Z(n162));
Q_OR03 U490 ( .A0(f32_mux_8_data[12]), .A1(f32_mux_7_data[12]), .A2(f32_mux_6_data[12]), .Z(n161));
Q_OR03 U491 ( .A0(n158), .A1(n159), .A2(n160), .Z(r32_formatted_reg_data[11]));
Q_OR03 U492 ( .A0(f32_mux_2_data[11]), .A1(f32_mux_1_data[11]), .A2(f32_mux_0_data[11]), .Z(n160));
Q_OR03 U493 ( .A0(f32_mux_5_data[11]), .A1(f32_mux_4_data[11]), .A2(f32_mux_3_data[11]), .Z(n159));
Q_OR03 U494 ( .A0(f32_mux_8_data[11]), .A1(f32_mux_7_data[11]), .A2(f32_mux_6_data[11]), .Z(n158));
Q_OR03 U495 ( .A0(n155), .A1(n156), .A2(n157), .Z(r32_formatted_reg_data[10]));
Q_OR03 U496 ( .A0(f32_mux_2_data[10]), .A1(f32_mux_1_data[10]), .A2(f32_mux_0_data[10]), .Z(n157));
Q_OR03 U497 ( .A0(f32_mux_5_data[10]), .A1(f32_mux_4_data[10]), .A2(f32_mux_3_data[10]), .Z(n156));
Q_OR03 U498 ( .A0(f32_mux_8_data[10]), .A1(f32_mux_7_data[10]), .A2(f32_mux_6_data[10]), .Z(n155));
Q_OR03 U499 ( .A0(n152), .A1(n153), .A2(n154), .Z(r32_formatted_reg_data[9]));
Q_OR03 U500 ( .A0(f32_mux_2_data[9]), .A1(f32_mux_1_data[9]), .A2(f32_mux_0_data[9]), .Z(n154));
Q_OR03 U501 ( .A0(f32_mux_5_data[9]), .A1(f32_mux_4_data[9]), .A2(f32_mux_3_data[9]), .Z(n153));
Q_OR03 U502 ( .A0(f32_mux_8_data[9]), .A1(f32_mux_7_data[9]), .A2(f32_mux_6_data[9]), .Z(n152));
Q_OR03 U503 ( .A0(n149), .A1(n150), .A2(n151), .Z(r32_formatted_reg_data[8]));
Q_OR03 U504 ( .A0(f32_mux_2_data[8]), .A1(f32_mux_1_data[8]), .A2(f32_mux_0_data[8]), .Z(n151));
Q_OR03 U505 ( .A0(f32_mux_5_data[8]), .A1(f32_mux_4_data[8]), .A2(f32_mux_3_data[8]), .Z(n150));
Q_OR03 U506 ( .A0(f32_mux_8_data[8]), .A1(f32_mux_7_data[8]), .A2(f32_mux_6_data[8]), .Z(n149));
Q_OR03 U507 ( .A0(n146), .A1(n147), .A2(n148), .Z(r32_formatted_reg_data[7]));
Q_OR03 U508 ( .A0(f32_mux_2_data[7]), .A1(f32_mux_1_data[7]), .A2(f32_mux_0_data[7]), .Z(n148));
Q_OR03 U509 ( .A0(f32_mux_5_data[7]), .A1(f32_mux_4_data[7]), .A2(f32_mux_3_data[7]), .Z(n147));
Q_OR03 U510 ( .A0(f32_mux_8_data[7]), .A1(f32_mux_7_data[7]), .A2(f32_mux_6_data[7]), .Z(n146));
Q_OR03 U511 ( .A0(n143), .A1(n144), .A2(n145), .Z(r32_formatted_reg_data[6]));
Q_OR03 U512 ( .A0(f32_mux_2_data[6]), .A1(f32_mux_1_data[6]), .A2(f32_mux_0_data[6]), .Z(n145));
Q_OR03 U513 ( .A0(f32_mux_5_data[6]), .A1(f32_mux_4_data[6]), .A2(f32_mux_3_data[6]), .Z(n144));
Q_OR03 U514 ( .A0(f32_mux_8_data[6]), .A1(f32_mux_7_data[6]), .A2(f32_mux_6_data[6]), .Z(n143));
Q_OR03 U515 ( .A0(n140), .A1(n141), .A2(n142), .Z(r32_formatted_reg_data[5]));
Q_OR03 U516 ( .A0(f32_mux_2_data[5]), .A1(f32_mux_1_data[5]), .A2(f32_mux_0_data[5]), .Z(n142));
Q_OR03 U517 ( .A0(f32_mux_5_data[5]), .A1(f32_mux_4_data[5]), .A2(f32_mux_3_data[5]), .Z(n141));
Q_OR03 U518 ( .A0(f32_mux_8_data[5]), .A1(f32_mux_7_data[5]), .A2(f32_mux_6_data[5]), .Z(n140));
Q_OR03 U519 ( .A0(n137), .A1(n138), .A2(n139), .Z(r32_formatted_reg_data[4]));
Q_OR03 U520 ( .A0(f32_mux_2_data[4]), .A1(f32_mux_1_data[4]), .A2(f32_mux_0_data[4]), .Z(n139));
Q_OR03 U521 ( .A0(f32_mux_5_data[4]), .A1(f32_mux_4_data[4]), .A2(f32_mux_3_data[4]), .Z(n138));
Q_OR03 U522 ( .A0(f32_mux_8_data[4]), .A1(f32_mux_7_data[4]), .A2(f32_mux_6_data[4]), .Z(n137));
Q_OR03 U523 ( .A0(n134), .A1(n135), .A2(n136), .Z(r32_formatted_reg_data[3]));
Q_OR03 U524 ( .A0(f32_mux_2_data[3]), .A1(f32_mux_1_data[3]), .A2(f32_mux_0_data[3]), .Z(n136));
Q_OR03 U525 ( .A0(f32_mux_5_data[3]), .A1(f32_mux_4_data[3]), .A2(f32_mux_3_data[3]), .Z(n135));
Q_OR03 U526 ( .A0(f32_mux_8_data[3]), .A1(f32_mux_7_data[3]), .A2(f32_mux_6_data[3]), .Z(n134));
Q_OR03 U527 ( .A0(n131), .A1(n132), .A2(n133), .Z(r32_formatted_reg_data[2]));
Q_OR03 U528 ( .A0(f32_mux_2_data[2]), .A1(f32_mux_1_data[2]), .A2(f32_mux_0_data[2]), .Z(n133));
Q_OR03 U529 ( .A0(f32_mux_5_data[2]), .A1(f32_mux_4_data[2]), .A2(f32_mux_3_data[2]), .Z(n132));
Q_OR03 U530 ( .A0(f32_mux_8_data[2]), .A1(f32_mux_7_data[2]), .A2(f32_mux_6_data[2]), .Z(n131));
Q_OR03 U531 ( .A0(n128), .A1(n129), .A2(n130), .Z(r32_formatted_reg_data[1]));
Q_OR03 U532 ( .A0(f32_mux_2_data[1]), .A1(f32_mux_1_data[1]), .A2(f32_mux_0_data[1]), .Z(n130));
Q_OR03 U533 ( .A0(f32_mux_5_data[1]), .A1(f32_mux_4_data[1]), .A2(f32_mux_3_data[1]), .Z(n129));
Q_OR03 U534 ( .A0(f32_mux_8_data[1]), .A1(f32_mux_7_data[1]), .A2(f32_mux_6_data[1]), .Z(n128));
Q_OR03 U535 ( .A0(n125), .A1(n126), .A2(n127), .Z(r32_formatted_reg_data[0]));
Q_OR03 U536 ( .A0(f32_mux_2_data[0]), .A1(f32_mux_1_data[0]), .A2(f32_mux_0_data[0]), .Z(n127));
Q_OR03 U537 ( .A0(f32_mux_5_data[0]), .A1(f32_mux_4_data[0]), .A2(f32_mux_3_data[0]), .Z(n126));
Q_OR03 U538 ( .A0(f32_mux_8_data[0]), .A1(f32_mux_7_data[0]), .A2(f32_mux_6_data[0]), .Z(n125));
Q_OR02 U539 ( .A0(f_err_ack), .A1(n124), .Z(o_err_ack));
Q_NR02 U540 ( .A0(n122), .A1(w_valid_rd_addr), .Z(n124));
Q_INV U541 ( .A(w_valid_rd_addr), .Z(n123));
Q_OR02 U542 ( .A0(f_ack), .A1(w_do_write), .Z(o_ack));
Q_INV U543 ( .A(n122), .Z(w_do_write));
Q_OR03 U544 ( .A0(n435), .A1(f_state[1]), .A2(f_state[2]), .Z(n122));
Q_AN02 U545 ( .A0(w_do_read), .A1(n123), .Z(w_next_err_ack));
Q_AN03 U546 ( .A0(f_state[0]), .A1(n121), .A2(f_state[2]), .Z(w_next_ack));
Q_OR02 U547 ( .A0(n119), .A1(n120), .Z(w_valid_wr_addr));
Q_OR03 U548 ( .A0(n116), .A1(n117), .A2(n118), .Z(n120));
Q_OR03 U549 ( .A0(n67), .A1(n95), .A2(n115), .Z(n119));
Q_OR03 U550 ( .A0(n37), .A1(n43), .A2(n55), .Z(n118));
Q_OR03 U551 ( .A0(n31), .A1(n6), .A2(n25), .Z(n117));
Q_OR03 U552 ( .A0(n81), .A1(n74), .A2(n48), .Z(n116));
Q_NR03 U553 ( .A0(n1), .A1(n105), .A2(n114), .Z(n115));
Q_OR03 U554 ( .A0(n107), .A1(n113), .A2(n112), .Z(n114));
Q_AN02 U555 ( .A0(ws_addr[10]), .A1(n109), .Z(n113));
Q_AN03 U556 ( .A0(ws_addr[10]), .A1(n110), .A2(n111), .Z(n112));
Q_OA21 U557 ( .A0(ws_addr[1]), .A1(ws_addr[0]), .B0(ws_addr[2]), .Z(n111));
Q_AN02 U558 ( .A0(n108), .A1(ws_addr[3]), .Z(n110));
Q_AN02 U559 ( .A0(ws_addr[6]), .A1(ws_addr[5]), .Z(n109));
Q_AN02 U560 ( .A0(ws_addr[6]), .A1(ws_addr[4]), .Z(n108));
Q_AO21 U561 ( .A0(ws_addr[10]), .A1(ws_addr[9]), .B0(n106), .Z(n107));
Q_OA21 U562 ( .A0(ws_addr[8]), .A1(ws_addr[7]), .B0(ws_addr[10]), .Z(n106));
Q_OR03 U563 ( .A0(n99), .A1(n104), .A2(n103), .Z(n105));
Q_AN02 U564 ( .A0(n7), .A1(n101), .Z(n104));
Q_AN02 U565 ( .A0(n102), .A1(n19), .Z(n103));
Q_NR02 U566 ( .A0(ws_addr[10]), .A1(ws_addr[4]), .Z(n102));
Q_OR02 U567 ( .A0(n4922), .A1(n100), .Z(n101));
Q_NR02 U568 ( .A0(ws_addr[4]), .A1(ws_addr[3]), .Z(n100));
Q_NR02 U569 ( .A0(ws_addr[10]), .A1(ws_addr[9]), .Z(n98));
Q_OR03 U570 ( .A0(n97), .A1(n96), .A2(n98), .Z(n99));
Q_NR02 U571 ( .A0(ws_addr[10]), .A1(ws_addr[8]), .Z(n97));
Q_NR02 U572 ( .A0(ws_addr[10]), .A1(ws_addr[7]), .Z(n96));
Q_NR03 U573 ( .A0(n1), .A1(n87), .A2(n94), .Z(n95));
Q_OR03 U574 ( .A0(ws_addr[10]), .A1(n93), .A2(n92), .Z(n94));
Q_AN02 U575 ( .A0(n88), .A1(n91), .Z(n93));
Q_AN03 U576 ( .A0(n88), .A1(n109), .A2(n111), .Z(n92));
Q_OR02 U577 ( .A0(n90), .A1(n89), .Z(n91));
Q_AN02 U578 ( .A0(n109), .A1(ws_addr[4]), .Z(n90));
Q_AN02 U579 ( .A0(n109), .A1(ws_addr[3]), .Z(n89));
Q_AN02 U580 ( .A0(n77), .A1(ws_addr[7]), .Z(n88));
Q_OR03 U581 ( .A0(n99), .A1(n86), .A2(n85), .Z(n87));
Q_AN02 U582 ( .A0(n7), .A1(n84), .Z(n86));
Q_AN03 U583 ( .A0(n7), .A1(n83), .A2(n19), .Z(n85));
Q_AN02 U584 ( .A0(n83), .A1(n16), .Z(n84));
Q_AN02 U585 ( .A0(n82), .A1(n15), .Z(n83));
Q_NR02 U586 ( .A0(ws_addr[6]), .A1(ws_addr[5]), .Z(n82));
Q_NR03 U587 ( .A0(n1), .A1(n76), .A2(n80), .Z(n81));
Q_OR03 U588 ( .A0(ws_addr[10]), .A1(n79), .A2(n78), .Z(n80));
Q_AN02 U589 ( .A0(n88), .A1(n70), .Z(n79));
Q_AN02 U590 ( .A0(n88), .A1(n111), .Z(n78));
Q_AN02 U591 ( .A0(ws_addr[9]), .A1(ws_addr[8]), .Z(n77));
Q_AN02 U592 ( .A0(n96), .A1(n84), .Z(n75));
Q_OR03 U593 ( .A0(n98), .A1(n97), .A2(n75), .Z(n76));
Q_NR03 U594 ( .A0(n1), .A1(n68), .A2(n73), .Z(n74));
Q_OR03 U595 ( .A0(n69), .A1(n72), .A2(n71), .Z(n73));
Q_AN02 U596 ( .A0(n77), .A1(n70), .Z(n72));
Q_AN02 U597 ( .A0(n77), .A1(n63), .Z(n71));
Q_ND02 U598 ( .A0(n82), .A1(n100), .Z(n70));
Q_OR02 U599 ( .A0(ws_addr[10]), .A1(n88), .Z(n69));
Q_AO21 U600 ( .A0(n97), .A1(n4922), .B0(n57), .Z(n68));
Q_NR03 U601 ( .A0(n1), .A1(n60), .A2(n66), .Z(n67));
Q_OR03 U602 ( .A0(n61), .A1(n65), .A2(n64), .Z(n66));
Q_AN02 U603 ( .A0(n62), .A1(n109), .Z(n65));
Q_AN03 U604 ( .A0(n62), .A1(n110), .A2(n63), .Z(n64));
Q_OR03 U605 ( .A0(ws_addr[2]), .A1(ws_addr[1]), .A2(ws_addr[0]), .Z(n63));
Q_AN02 U606 ( .A0(ws_addr[9]), .A1(ws_addr[7]), .Z(n62));
Q_OR02 U607 ( .A0(ws_addr[10]), .A1(n77), .Z(n61));
Q_AO21 U608 ( .A0(n97), .A1(n59), .B0(n57), .Z(n60));
Q_AO21 U609 ( .A0(n13), .A1(n58), .B0(n82), .Z(n59));
Q_ND02 U610 ( .A0(ws_addr[4]), .A1(ws_addr[3]), .Z(n58));
Q_OR02 U611 ( .A0(n98), .A1(n56), .Z(n57));
Q_AN02 U612 ( .A0(n97), .A1(n10), .Z(n56));
Q_NR03 U613 ( .A0(n1), .A1(n49), .A2(n54), .Z(n55));
Q_OR03 U614 ( .A0(n61), .A1(n53), .A2(n52), .Z(n54));
Q_AN03 U615 ( .A0(n62), .A1(n50), .A2(n63), .Z(n52));
Q_OA21 U616 ( .A0(ws_addr[6]), .A1(n51), .B0(n62), .Z(n53));
Q_AN02 U617 ( .A0(n50), .A1(ws_addr[3]), .Z(n51));
Q_AN02 U618 ( .A0(ws_addr[5]), .A1(ws_addr[4]), .Z(n50));
Q_AO21 U619 ( .A0(n97), .A1(n83), .B0(n57), .Z(n49));
Q_NR03 U620 ( .A0(n1), .A1(n44), .A2(n47), .Z(n48));
Q_OR03 U621 ( .A0(n61), .A1(n46), .A2(n45), .Z(n47));
Q_AN02 U622 ( .A0(n62), .A1(n4925), .Z(n46));
Q_AN03 U623 ( .A0(n62), .A1(ws_addr[3]), .A2(n63), .Z(n45));
Q_AO21 U624 ( .A0(n56), .A1(n101), .B0(n98), .Z(n44));
Q_NR03 U625 ( .A0(n1), .A1(n38), .A2(n42), .Z(n43));
Q_OR03 U626 ( .A0(n39), .A1(n41), .A2(n40), .Z(n42));
Q_AN02 U627 ( .A0(ws_addr[9]), .A1(n91), .Z(n41));
Q_AN03 U628 ( .A0(ws_addr[9]), .A1(n109), .A2(n63), .Z(n40));
Q_OR03 U629 ( .A0(n77), .A1(n62), .A2(ws_addr[10]), .Z(n39));
Q_AO21 U630 ( .A0(n56), .A1(n13), .B0(n98), .Z(n38));
Q_NR03 U631 ( .A0(n1), .A1(n33), .A2(n36), .Z(n37));
Q_OR03 U632 ( .A0(n39), .A1(n35), .A2(n34), .Z(n36));
Q_AN02 U633 ( .A0(ws_addr[9]), .A1(ws_addr[6]), .Z(n35));
Q_AN03 U634 ( .A0(ws_addr[9]), .A1(n51), .A2(n63), .Z(n34));
Q_AO21 U635 ( .A0(n56), .A1(n32), .B0(n98), .Z(n33));
Q_AO21 U636 ( .A0(n82), .A1(n16), .B0(n83), .Z(n32));
Q_NR03 U637 ( .A0(n1), .A1(n26), .A2(n30), .Z(n31));
Q_OR03 U638 ( .A0(n39), .A1(n29), .A2(n28), .Z(n30));
Q_AN02 U639 ( .A0(ws_addr[9]), .A1(n27), .Z(n29));
Q_AN03 U640 ( .A0(ws_addr[9]), .A1(ws_addr[4]), .A2(n63), .Z(n28));
Q_AO21 U641 ( .A0(ws_addr[4]), .A1(ws_addr[3]), .B0(n4923), .Z(n27));
Q_AO21 U642 ( .A0(n98), .A1(n4924), .B0(n12), .Z(n26));
Q_NR03 U643 ( .A0(n1), .A1(n20), .A2(n24), .Z(n25));
Q_OR03 U644 ( .A0(n4921), .A1(n23), .A2(n22), .Z(n24));
Q_AN02 U645 ( .A0(n21), .A1(n90), .Z(n23));
Q_AN03 U646 ( .A0(n21), .A1(n89), .A2(n63), .Z(n22));
Q_AN02 U647 ( .A0(ws_addr[8]), .A1(ws_addr[7]), .Z(n21));
Q_AO21 U648 ( .A0(n98), .A1(n18), .B0(n12), .Z(n20));
Q_INV U649 ( .A(ws_addr[2]), .Z(n19));
Q_AO21 U650 ( .A0(n17), .A1(n16), .B0(n13), .Z(n18));
Q_NR02 U651 ( .A0(ws_addr[5]), .A1(ws_addr[4]), .Z(n17));
Q_INV U652 ( .A(ws_addr[3]), .Z(n16));
Q_INV U653 ( .A(ws_addr[4]), .Z(n15));
Q_INV U654 ( .A(ws_addr[5]), .Z(n14));
Q_INV U655 ( .A(ws_addr[6]), .Z(n13));
Q_AN02 U656 ( .A0(n98), .A1(n11), .Z(n12));
Q_ND02 U657 ( .A0(ws_addr[8]), .A1(ws_addr[7]), .Z(n11));
Q_INV U658 ( .A(ws_addr[7]), .Z(n10));
Q_INV U659 ( .A(ws_addr[8]), .Z(n9));
Q_INV U660 ( .A(ws_addr[9]), .Z(n8));
Q_INV U661 ( .A(ws_addr[10]), .Z(n7));
Q_NR02 U662 ( .A0(n1), .A1(n5), .Z(n6));
Q_OR03 U663 ( .A0(n4921), .A1(n4), .A2(n3), .Z(n5));
Q_AN03 U664 ( .A0(n21), .A1(ws_addr[6]), .A2(n63), .Z(n3));
Q_OA21 U665 ( .A0(n109), .A1(n2), .B0(n21), .Z(n4));
Q_AO21 U666 ( .A0(ws_addr[6]), .A1(ws_addr[3]), .B0(n108), .Z(n2));
Q_INV U667 ( .A(n1), .Z(w_32b_aligned));
Q_OR02 U668 ( .A0(o_reg_addr[0]), .A1(o_reg_addr[1]), .Z(n1));
ixc_assign _zz_strnp_3 ( n_rd_strobe, i_rd_strb);
ixc_assign _zz_strnp_2 ( n_wr_strobe, i_wr_strb);
ixc_assign_11 _zz_strnp_1 ( ws_addr[10:0], o_reg_addr[10:0]);
ixc_assign_11 _zz_strnp_0 ( ws_read_addr[10:0], o_reg_addr[10:0]);
Q_OR02 U673 ( .A0(f_state[1]), .A1(n435), .Z(n441));
Q_OA21 U674 ( .A0(n436), .A1(n441), .B0(n437), .Z(n438));
Q_INV U675 ( .A(n_rd_strobe), .Z(n437));
Q_OR02 U676 ( .A0(n_wr_strobe), .A1(n438), .Z(n439));
Q_INV U677 ( .A(n439), .Z(w_next_state[2]));
Q_OR02 U678 ( .A0(n443), .A1(n441), .Z(n440));
Q_INV U679 ( .A(n440), .Z(w_next_state[1]));
Q_INV U680 ( .A(n441), .Z(n442));
Q_OR02 U681 ( .A0(n_wr_strobe), .A1(n_rd_strobe), .Z(n443));
Q_OR02 U682 ( .A0(n443), .A1(n442), .Z(w_next_state[0]));
Q_AN02 U683 ( .A0(n445), .A1(r32_formatted_reg_data[0]), .Z(o_rd_data[0]));
Q_AN02 U684 ( .A0(n445), .A1(r32_formatted_reg_data[1]), .Z(o_rd_data[1]));
Q_AN02 U685 ( .A0(n445), .A1(r32_formatted_reg_data[2]), .Z(o_rd_data[2]));
Q_AN02 U686 ( .A0(n445), .A1(r32_formatted_reg_data[3]), .Z(o_rd_data[3]));
Q_AN02 U687 ( .A0(n445), .A1(r32_formatted_reg_data[4]), .Z(o_rd_data[4]));
Q_AN02 U688 ( .A0(n445), .A1(r32_formatted_reg_data[5]), .Z(o_rd_data[5]));
Q_AN02 U689 ( .A0(n445), .A1(r32_formatted_reg_data[6]), .Z(o_rd_data[6]));
Q_AN02 U690 ( .A0(n445), .A1(r32_formatted_reg_data[7]), .Z(o_rd_data[7]));
Q_AN02 U691 ( .A0(n445), .A1(r32_formatted_reg_data[8]), .Z(o_rd_data[8]));
Q_AN02 U692 ( .A0(n445), .A1(r32_formatted_reg_data[9]), .Z(o_rd_data[9]));
Q_AN02 U693 ( .A0(n445), .A1(r32_formatted_reg_data[10]), .Z(o_rd_data[10]));
Q_AN02 U694 ( .A0(n445), .A1(r32_formatted_reg_data[11]), .Z(o_rd_data[11]));
Q_AN02 U695 ( .A0(n445), .A1(r32_formatted_reg_data[12]), .Z(o_rd_data[12]));
Q_AN02 U696 ( .A0(n445), .A1(r32_formatted_reg_data[13]), .Z(o_rd_data[13]));
Q_AN02 U697 ( .A0(n445), .A1(r32_formatted_reg_data[14]), .Z(o_rd_data[14]));
Q_AN02 U698 ( .A0(n445), .A1(r32_formatted_reg_data[15]), .Z(o_rd_data[15]));
Q_AN02 U699 ( .A0(n445), .A1(r32_formatted_reg_data[16]), .Z(o_rd_data[16]));
Q_AN02 U700 ( .A0(n445), .A1(r32_formatted_reg_data[17]), .Z(o_rd_data[17]));
Q_AN02 U701 ( .A0(n445), .A1(r32_formatted_reg_data[18]), .Z(o_rd_data[18]));
Q_AN02 U702 ( .A0(n445), .A1(r32_formatted_reg_data[19]), .Z(o_rd_data[19]));
Q_AN02 U703 ( .A0(n445), .A1(r32_formatted_reg_data[20]), .Z(o_rd_data[20]));
Q_AN02 U704 ( .A0(n445), .A1(r32_formatted_reg_data[21]), .Z(o_rd_data[21]));
Q_AN02 U705 ( .A0(n445), .A1(r32_formatted_reg_data[22]), .Z(o_rd_data[22]));
Q_AN02 U706 ( .A0(n445), .A1(r32_formatted_reg_data[23]), .Z(o_rd_data[23]));
Q_AN02 U707 ( .A0(n445), .A1(r32_formatted_reg_data[24]), .Z(o_rd_data[24]));
Q_AN02 U708 ( .A0(n445), .A1(r32_formatted_reg_data[25]), .Z(o_rd_data[25]));
Q_AN02 U709 ( .A0(n445), .A1(r32_formatted_reg_data[26]), .Z(o_rd_data[26]));
Q_AN02 U710 ( .A0(n445), .A1(r32_formatted_reg_data[27]), .Z(o_rd_data[27]));
Q_AN02 U711 ( .A0(n445), .A1(r32_formatted_reg_data[28]), .Z(o_rd_data[28]));
Q_AN02 U712 ( .A0(n445), .A1(r32_formatted_reg_data[29]), .Z(o_rd_data[29]));
Q_AN02 U713 ( .A0(n445), .A1(r32_formatted_reg_data[30]), .Z(o_rd_data[30]));
Q_AN02 U714 ( .A0(n445), .A1(r32_formatted_reg_data[31]), .Z(o_rd_data[31]));
Q_AN02 U715 ( .A0(o_ack), .A1(n444), .Z(n445));
Q_AN02 U716 ( .A0(n446), .A1(i_wr_strb), .Z(n451));
Q_ND02 U717 ( .A0(n448), .A1(n449), .Z(n447));
Q_INV U718 ( .A(o_ack), .Z(n449));
Q_NR02 U719 ( .A0(i_sw_init), .A1(i_wr_strb), .Z(n448));
Q_INV U720 ( .A(i_wr_strb), .Z(n450));
Q_INV U721 ( .A(i_sw_init), .Z(n446));
Q_MX02 U722 ( .S(n4313), .A0(i_im_consumed[0]), .A1(i_im_available[0]), .Z(n452));
Q_MX04 U723 ( .S0(n4313), .S1(n4314), .A0(i_sa_snapshot_ia_status[0]), .A1(i_sa_snapshot_ia_capability[0]), .A2(i_regs_sa_ctrl[0]), .A3(i_tready_override[0]), .Z(n453));
Q_MX02 U724 ( .S(n4315), .A0(n453), .A1(n452), .Z(n454));
Q_MX08 U725 ( .S0(n4313), .S1(n4314), .S2(n4315), .A0(o_sa_count_ia_wdata_part0[0]), .A1(i_sa_count_ia_status[0]), .A2(i_sa_count_ia_capability[0]), .A3(i_sa_snapshot_ia_rdata_part1[0]), .A4(i_sa_snapshot_ia_rdata_part0[0]), .A5(o_sa_snapshot_ia_config[0]), .A6(o_sa_snapshot_ia_wdata_part1[0]), .A7(o_sa_snapshot_ia_wdata_part0[0]), .Z(n455));
Q_MX02 U726 ( .S(n4316), .A0(n455), .A1(n454), .Z(n456));
Q_MX04 U727 ( .S0(n4313), .S1(n4314), .A0(i_sa_count_ia_rdata_part1[0]), .A1(i_sa_count_ia_rdata_part0[0]), .A2(o_sa_count_ia_config[0]), .A3(o_sa_count_ia_wdata_part1[0]), .Z(n457));
Q_MX04 U728 ( .S0(n4313), .S1(n4314), .A0(o_cddip_decrypt_kop_fifo_override[0]), .A1(o_cceip_validate_kop_fifo_override[0]), .A2(o_cceip_encrypt_kop_fifo_override[0]), .A3(i_idle_components[0]), .Z(n458));
Q_MX04 U729 ( .S0(n4313), .S1(n4314), .A0(o_sa_ctrl_ia_wdata_part0[0]), .A1(i_sa_ctrl_ia_status[0]), .A2(i_sa_ctrl_ia_capability[0]), .A3(i_sa_global_ctrl[0]), .Z(n459));
Q_MX02 U730 ( .S(n4313), .A0(i_sa_ctrl_ia_rdata_part0[0]), .A1(o_sa_ctrl_ia_config[0]), .Z(n460));
Q_AN02 U731 ( .A0(n4313), .A1(o_kdf_test_key_size_config[0]), .Z(n461));
Q_MX02 U732 ( .S(n4314), .A0(n461), .A1(n460), .Z(n462));
Q_MX04 U733 ( .S0(n4315), .S1(n4316), .A0(n462), .A1(n459), .A2(n458), .A3(n457), .Z(n463));
Q_MX02 U734 ( .S(n4317), .A0(n463), .A1(n456), .Z(r32_mux_8_data[0]));
Q_MX02 U735 ( .S(n4313), .A0(i_im_consumed[1]), .A1(i_im_available[1]), .Z(n464));
Q_MX04 U736 ( .S0(n4313), .S1(n4314), .A0(i_sa_snapshot_ia_status[1]), .A1(i_sa_snapshot_ia_capability[1]), .A2(i_regs_sa_ctrl[1]), .A3(i_tready_override[1]), .Z(n465));
Q_MX02 U737 ( .S(n4315), .A0(n465), .A1(n464), .Z(n466));
Q_MX08 U738 ( .S0(n4313), .S1(n4314), .S2(n4315), .A0(o_sa_count_ia_wdata_part0[1]), .A1(i_sa_count_ia_status[1]), .A2(i_sa_count_ia_capability[1]), .A3(i_sa_snapshot_ia_rdata_part1[1]), .A4(i_sa_snapshot_ia_rdata_part0[1]), .A5(o_sa_snapshot_ia_config[1]), .A6(o_sa_snapshot_ia_wdata_part1[1]), .A7(o_sa_snapshot_ia_wdata_part0[1]), .Z(n467));
Q_MX02 U739 ( .S(n4316), .A0(n467), .A1(n466), .Z(n468));
Q_MX04 U740 ( .S0(n4313), .S1(n4314), .A0(i_sa_count_ia_rdata_part1[1]), .A1(i_sa_count_ia_rdata_part0[1]), .A2(o_sa_count_ia_config[1]), .A3(o_sa_count_ia_wdata_part1[1]), .Z(n469));
Q_MX04 U741 ( .S0(n4313), .S1(n4314), .A0(o_cddip_decrypt_kop_fifo_override[1]), .A1(o_cceip_validate_kop_fifo_override[1]), .A2(o_cceip_encrypt_kop_fifo_override[1]), .A3(i_idle_components[1]), .Z(n470));
Q_MX04 U742 ( .S0(n4313), .S1(n4314), .A0(o_sa_ctrl_ia_wdata_part0[1]), .A1(i_sa_ctrl_ia_status[1]), .A2(i_sa_ctrl_ia_capability[1]), .A3(i_sa_global_ctrl[1]), .Z(n471));
Q_MX02 U743 ( .S(n4313), .A0(i_sa_ctrl_ia_rdata_part0[1]), .A1(o_sa_ctrl_ia_config[1]), .Z(n472));
Q_AN02 U744 ( .A0(n4313), .A1(o_kdf_test_key_size_config[1]), .Z(n473));
Q_MX02 U745 ( .S(n4314), .A0(n473), .A1(n472), .Z(n474));
Q_MX04 U746 ( .S0(n4315), .S1(n4316), .A0(n474), .A1(n471), .A2(n470), .A3(n469), .Z(n475));
Q_MX02 U747 ( .S(n4317), .A0(n475), .A1(n468), .Z(r32_mux_8_data[1]));
Q_MX02 U748 ( .S(n4313), .A0(i_im_consumed[2]), .A1(i_im_available[2]), .Z(n476));
Q_MX04 U749 ( .S0(n4313), .S1(n4314), .A0(i_sa_snapshot_ia_status[2]), .A1(i_sa_snapshot_ia_capability[2]), .A2(i_regs_sa_ctrl[2]), .A3(i_tready_override[2]), .Z(n477));
Q_MX02 U750 ( .S(n4315), .A0(n477), .A1(n476), .Z(n478));
Q_MX08 U751 ( .S0(n4313), .S1(n4314), .S2(n4315), .A0(o_sa_count_ia_wdata_part0[2]), .A1(i_sa_count_ia_status[2]), .A2(i_sa_count_ia_capability[2]), .A3(i_sa_snapshot_ia_rdata_part1[2]), .A4(i_sa_snapshot_ia_rdata_part0[2]), .A5(o_sa_snapshot_ia_config[2]), .A6(o_sa_snapshot_ia_wdata_part1[2]), .A7(o_sa_snapshot_ia_wdata_part0[2]), .Z(n479));
Q_MX02 U752 ( .S(n4316), .A0(n479), .A1(n478), .Z(n480));
Q_MX04 U753 ( .S0(n4313), .S1(n4314), .A0(i_sa_count_ia_rdata_part1[2]), .A1(i_sa_count_ia_rdata_part0[2]), .A2(o_sa_count_ia_config[2]), .A3(o_sa_count_ia_wdata_part1[2]), .Z(n481));
Q_MX04 U754 ( .S0(n4313), .S1(n4314), .A0(o_cddip_decrypt_kop_fifo_override[2]), .A1(o_cceip_validate_kop_fifo_override[2]), .A2(o_cceip_encrypt_kop_fifo_override[2]), .A3(i_idle_components[2]), .Z(n482));
Q_MX04 U755 ( .S0(n4313), .S1(n4314), .A0(o_sa_ctrl_ia_wdata_part0[2]), .A1(i_sa_ctrl_ia_status[2]), .A2(i_sa_ctrl_ia_capability[2]), .A3(i_sa_global_ctrl[2]), .Z(n483));
Q_MX02 U756 ( .S(n4313), .A0(i_sa_ctrl_ia_rdata_part0[2]), .A1(o_sa_ctrl_ia_config[2]), .Z(n484));
Q_AN02 U757 ( .A0(n4313), .A1(o_kdf_test_key_size_config[2]), .Z(n485));
Q_MX02 U758 ( .S(n4314), .A0(n485), .A1(n484), .Z(n486));
Q_MX04 U759 ( .S0(n4315), .S1(n4316), .A0(n486), .A1(n483), .A2(n482), .A3(n481), .Z(n487));
Q_MX02 U760 ( .S(n4317), .A0(n487), .A1(n480), .Z(r32_mux_8_data[2]));
Q_MX02 U761 ( .S(n4313), .A0(i_im_consumed[3]), .A1(i_im_available[3]), .Z(n488));
Q_MX04 U762 ( .S0(n4313), .S1(n4314), .A0(i_sa_snapshot_ia_status[3]), .A1(i_sa_snapshot_ia_capability[3]), .A2(i_regs_sa_ctrl[3]), .A3(i_tready_override[3]), .Z(n489));
Q_MX02 U763 ( .S(n4315), .A0(n489), .A1(n488), .Z(n490));
Q_MX08 U764 ( .S0(n4313), .S1(n4314), .S2(n4315), .A0(o_sa_count_ia_wdata_part0[3]), .A1(i_sa_count_ia_status[3]), .A2(i_sa_count_ia_capability[3]), .A3(i_sa_snapshot_ia_rdata_part1[3]), .A4(i_sa_snapshot_ia_rdata_part0[3]), .A5(o_sa_snapshot_ia_config[3]), .A6(o_sa_snapshot_ia_wdata_part1[3]), .A7(o_sa_snapshot_ia_wdata_part0[3]), .Z(n491));
Q_MX02 U765 ( .S(n4316), .A0(n491), .A1(n490), .Z(n492));
Q_MX04 U766 ( .S0(n4313), .S1(n4314), .A0(i_sa_count_ia_rdata_part1[3]), .A1(i_sa_count_ia_rdata_part0[3]), .A2(o_sa_count_ia_config[3]), .A3(o_sa_count_ia_wdata_part1[3]), .Z(n493));
Q_MX04 U767 ( .S0(n4313), .S1(n4314), .A0(o_cddip_decrypt_kop_fifo_override[3]), .A1(o_cceip_validate_kop_fifo_override[3]), .A2(o_cceip_encrypt_kop_fifo_override[3]), .A3(i_idle_components[3]), .Z(n494));
Q_MX04 U768 ( .S0(n4313), .S1(n4314), .A0(o_sa_ctrl_ia_wdata_part0[3]), .A1(i_sa_ctrl_ia_status[3]), .A2(i_sa_ctrl_ia_capability[3]), .A3(i_sa_global_ctrl[3]), .Z(n495));
Q_MX02 U769 ( .S(n4313), .A0(i_sa_ctrl_ia_rdata_part0[3]), .A1(o_sa_ctrl_ia_config[3]), .Z(n496));
Q_AN02 U770 ( .A0(n4313), .A1(o_kdf_test_key_size_config[3]), .Z(n497));
Q_MX02 U771 ( .S(n4314), .A0(n497), .A1(n496), .Z(n498));
Q_MX04 U772 ( .S0(n4315), .S1(n4316), .A0(n498), .A1(n495), .A2(n494), .A3(n493), .Z(n499));
Q_MX02 U773 ( .S(n4317), .A0(n499), .A1(n492), .Z(r32_mux_8_data[3]));
Q_MX02 U774 ( .S(n4313), .A0(i_im_consumed[4]), .A1(i_im_available[4]), .Z(n500));
Q_MX04 U775 ( .S0(n4313), .S1(n4314), .A0(i_sa_snapshot_ia_status[4]), .A1(i_sa_snapshot_ia_capability[4]), .A2(i_regs_sa_ctrl[4]), .A3(i_tready_override[4]), .Z(n501));
Q_MX02 U776 ( .S(n4315), .A0(n501), .A1(n500), .Z(n502));
Q_MX08 U777 ( .S0(n4313), .S1(n4314), .S2(n4315), .A0(o_sa_count_ia_wdata_part0[4]), .A1(i_sa_count_ia_status[4]), .A2(i_sa_count_ia_capability[4]), .A3(i_sa_snapshot_ia_rdata_part1[4]), .A4(i_sa_snapshot_ia_rdata_part0[4]), .A5(o_sa_snapshot_ia_config[4]), .A6(o_sa_snapshot_ia_wdata_part1[4]), .A7(o_sa_snapshot_ia_wdata_part0[4]), .Z(n503));
Q_MX02 U778 ( .S(n4316), .A0(n503), .A1(n502), .Z(n504));
Q_MX04 U779 ( .S0(n4313), .S1(n4314), .A0(i_sa_count_ia_rdata_part1[4]), .A1(i_sa_count_ia_rdata_part0[4]), .A2(o_sa_count_ia_config[4]), .A3(o_sa_count_ia_wdata_part1[4]), .Z(n505));
Q_MX04 U780 ( .S0(n4313), .S1(n4314), .A0(o_cddip_decrypt_kop_fifo_override[4]), .A1(o_cceip_validate_kop_fifo_override[4]), .A2(o_cceip_encrypt_kop_fifo_override[4]), .A3(i_idle_components[4]), .Z(n506));
Q_MX04 U781 ( .S0(n4313), .S1(n4314), .A0(o_sa_ctrl_ia_wdata_part0[4]), .A1(i_sa_ctrl_ia_status[4]), .A2(i_sa_ctrl_ia_capability[4]), .A3(i_sa_global_ctrl[4]), .Z(n507));
Q_MX02 U782 ( .S(n4313), .A0(i_sa_ctrl_ia_rdata_part0[4]), .A1(o_sa_ctrl_ia_config[4]), .Z(n508));
Q_AN02 U783 ( .A0(n4313), .A1(o_kdf_test_key_size_config[4]), .Z(n509));
Q_MX02 U784 ( .S(n4314), .A0(n509), .A1(n508), .Z(n510));
Q_MX04 U785 ( .S0(n4315), .S1(n4316), .A0(n510), .A1(n507), .A2(n506), .A3(n505), .Z(n511));
Q_MX02 U786 ( .S(n4317), .A0(n511), .A1(n504), .Z(r32_mux_8_data[4]));
Q_MX08 U787 ( .S0(n4318), .S1(n4319), .S2(n4320), .A0(i_sa_snapshot_ia_rdata_part0[5]), .A1(o_sa_snapshot_ia_wdata_part1[5]), .A2(o_sa_snapshot_ia_wdata_part0[5]), .A3(i_sa_snapshot_ia_capability[5]), .A4(i_regs_sa_ctrl[5]), .A5(i_tready_override[5]), .A6(i_im_consumed[5]), .A7(i_im_available[5]), .Z(n512));
Q_MX04 U788 ( .S0(n4318), .S1(n4319), .A0(o_sa_count_ia_wdata_part1[5]), .A1(o_sa_count_ia_wdata_part0[5]), .A2(i_sa_count_ia_capability[5]), .A3(i_sa_snapshot_ia_rdata_part1[5]), .Z(n513));
Q_MX04 U789 ( .S0(n4318), .S1(n4319), .A0(o_cceip_encrypt_kop_fifo_override[5]), .A1(i_idle_components[5]), .A2(i_sa_count_ia_rdata_part1[5]), .A3(i_sa_count_ia_rdata_part0[5]), .Z(n514));
Q_MX04 U790 ( .S0(n4318), .S1(n4319), .A0(i_sa_ctrl_ia_capability[5]), .A1(i_sa_global_ctrl[5]), .A2(o_cddip_decrypt_kop_fifo_override[5]), .A3(o_cceip_validate_kop_fifo_override[5]), .Z(n515));
Q_MX02 U791 ( .S(n4318), .A0(i_sa_ctrl_ia_rdata_part0[5]), .A1(o_sa_ctrl_ia_wdata_part0[5]), .Z(n516));
Q_AN02 U792 ( .A0(n4318), .A1(o_kdf_test_key_size_config[5]), .Z(n517));
Q_MX02 U793 ( .S(n4319), .A0(n517), .A1(n516), .Z(n518));
Q_MX04 U794 ( .S0(n4320), .S1(n4321), .A0(n518), .A1(n515), .A2(n514), .A3(n513), .Z(n519));
Q_MX02 U795 ( .S(n4322), .A0(n519), .A1(n512), .Z(r32_mux_8_data[5]));
Q_MX08 U796 ( .S0(n4318), .S1(n4319), .S2(n4320), .A0(i_sa_snapshot_ia_rdata_part0[6]), .A1(o_sa_snapshot_ia_wdata_part1[6]), .A2(o_sa_snapshot_ia_wdata_part0[6]), .A3(i_sa_snapshot_ia_capability[6]), .A4(i_regs_sa_ctrl[6]), .A5(i_tready_override[6]), .A6(i_im_consumed[6]), .A7(i_im_available[6]), .Z(n520));
Q_MX04 U797 ( .S0(n4318), .S1(n4319), .A0(o_sa_count_ia_wdata_part1[6]), .A1(o_sa_count_ia_wdata_part0[6]), .A2(i_sa_count_ia_capability[6]), .A3(i_sa_snapshot_ia_rdata_part1[6]), .Z(n521));
Q_MX04 U798 ( .S0(n4318), .S1(n4319), .A0(o_cceip_encrypt_kop_fifo_override[6]), .A1(i_idle_components[6]), .A2(i_sa_count_ia_rdata_part1[6]), .A3(i_sa_count_ia_rdata_part0[6]), .Z(n522));
Q_MX04 U799 ( .S0(n4318), .S1(n4319), .A0(i_sa_ctrl_ia_capability[6]), .A1(i_sa_global_ctrl[6]), .A2(o_cddip_decrypt_kop_fifo_override[6]), .A3(o_cceip_validate_kop_fifo_override[6]), .Z(n523));
Q_MX02 U800 ( .S(n4318), .A0(i_sa_ctrl_ia_rdata_part0[6]), .A1(o_sa_ctrl_ia_wdata_part0[6]), .Z(n524));
Q_AN02 U801 ( .A0(n4318), .A1(o_kdf_test_key_size_config[6]), .Z(n525));
Q_MX02 U802 ( .S(n4319), .A0(n525), .A1(n524), .Z(n526));
Q_MX04 U803 ( .S0(n4320), .S1(n4321), .A0(n526), .A1(n523), .A2(n522), .A3(n521), .Z(n527));
Q_MX02 U804 ( .S(n4322), .A0(n527), .A1(n520), .Z(r32_mux_8_data[6]));
Q_MX04 U805 ( .S0(n4323), .S1(n4324), .A0(i_sa_snapshot_ia_capability[7]), .A1(i_regs_sa_ctrl[7]), .A2(i_tready_override[7]), .A3(i_im_consumed[7]), .Z(n528));
Q_MX02 U806 ( .S(n4325), .A0(n528), .A1(i_im_available[7]), .Z(n529));
Q_MX04 U807 ( .S0(n4323), .S1(n4324), .A0(i_sa_snapshot_ia_rdata_part1[7]), .A1(i_sa_snapshot_ia_rdata_part0[7]), .A2(o_sa_snapshot_ia_wdata_part1[7]), .A3(o_sa_snapshot_ia_wdata_part0[7]), .Z(n530));
Q_MX04 U808 ( .S0(n4323), .S1(n4324), .A0(i_sa_count_ia_rdata_part0[7]), .A1(o_sa_count_ia_wdata_part1[7]), .A2(o_sa_count_ia_wdata_part0[7]), .A3(i_sa_count_ia_capability[7]), .Z(n531));
Q_MX04 U809 ( .S0(n4323), .S1(n4324), .A0(i_sa_ctrl_ia_capability[7]), .A1(i_sa_global_ctrl[7]), .A2(i_idle_components[7]), .A3(i_sa_count_ia_rdata_part1[7]), .Z(n532));
Q_MX02 U810 ( .S(n4323), .A0(i_sa_ctrl_ia_rdata_part0[7]), .A1(o_sa_ctrl_ia_wdata_part0[7]), .Z(n533));
Q_AN02 U811 ( .A0(n4323), .A1(o_kdf_test_key_size_config[7]), .Z(n534));
Q_MX02 U812 ( .S(n4324), .A0(n534), .A1(n533), .Z(n535));
Q_MX04 U813 ( .S0(n4325), .S1(n4326), .A0(n535), .A1(n532), .A2(n531), .A3(n530), .Z(n536));
Q_MX02 U814 ( .S(n4327), .A0(n536), .A1(n529), .Z(r32_mux_8_data[7]));
Q_MX04 U815 ( .S0(n4323), .S1(n4324), .A0(i_sa_snapshot_ia_capability[8]), .A1(i_regs_sa_ctrl[8]), .A2(i_tready_override[8]), .A3(i_im_consumed[8]), .Z(n537));
Q_MX02 U816 ( .S(n4325), .A0(n537), .A1(i_im_available[8]), .Z(n538));
Q_MX04 U817 ( .S0(n4323), .S1(n4324), .A0(i_sa_snapshot_ia_rdata_part1[8]), .A1(i_sa_snapshot_ia_rdata_part0[8]), .A2(o_sa_snapshot_ia_wdata_part1[8]), .A3(o_sa_snapshot_ia_wdata_part0[8]), .Z(n539));
Q_MX04 U818 ( .S0(n4323), .S1(n4324), .A0(i_sa_count_ia_rdata_part0[8]), .A1(o_sa_count_ia_wdata_part1[8]), .A2(o_sa_count_ia_wdata_part0[8]), .A3(i_sa_count_ia_capability[8]), .Z(n540));
Q_MX04 U819 ( .S0(n4323), .S1(n4324), .A0(i_sa_ctrl_ia_capability[8]), .A1(i_sa_global_ctrl[8]), .A2(i_idle_components[8]), .A3(i_sa_count_ia_rdata_part1[8]), .Z(n541));
Q_MX02 U820 ( .S(n4323), .A0(i_sa_ctrl_ia_rdata_part0[8]), .A1(o_sa_ctrl_ia_wdata_part0[8]), .Z(n542));
Q_AN02 U821 ( .A0(n4323), .A1(o_kdf_test_key_size_config[8]), .Z(n543));
Q_MX02 U822 ( .S(n4324), .A0(n543), .A1(n542), .Z(n544));
Q_MX04 U823 ( .S0(n4325), .S1(n4326), .A0(n544), .A1(n541), .A2(n540), .A3(n539), .Z(n545));
Q_MX02 U824 ( .S(n4327), .A0(n545), .A1(n538), .Z(r32_mux_8_data[8]));
Q_MX04 U825 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[9]), .A1(i_regs_sa_ctrl[9]), .A2(i_im_consumed[9]), .A3(i_im_available[9]), .Z(n546));
Q_MX04 U826 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[9]), .A1(i_sa_snapshot_ia_rdata_part0[9]), .A2(o_sa_snapshot_ia_wdata_part1[9]), .A3(o_sa_snapshot_ia_wdata_part0[9]), .Z(n547));
Q_MX04 U827 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[9]), .A1(o_sa_count_ia_wdata_part1[9]), .A2(o_sa_count_ia_wdata_part0[9]), .A3(i_sa_count_ia_capability[9]), .Z(n548));
Q_MX04 U828 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[9]), .A1(i_sa_global_ctrl[9]), .A2(i_idle_components[9]), .A3(i_sa_count_ia_rdata_part1[9]), .Z(n549));
Q_MX02 U829 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[9]), .A1(o_sa_ctrl_ia_wdata_part0[9]), .Z(n550));
Q_AN02 U830 ( .A0(n4328), .A1(o_kdf_test_key_size_config[9]), .Z(n551));
Q_MX02 U831 ( .S(n4329), .A0(n551), .A1(n550), .Z(n552));
Q_MX04 U832 ( .S0(n4330), .S1(n4326), .A0(n552), .A1(n549), .A2(n548), .A3(n547), .Z(n553));
Q_MX02 U833 ( .S(n4331), .A0(n553), .A1(n546), .Z(r32_mux_8_data[9]));
Q_MX04 U834 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[10]), .A1(i_regs_sa_ctrl[10]), .A2(i_im_consumed[10]), .A3(i_im_available[10]), .Z(n554));
Q_MX04 U835 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[10]), .A1(i_sa_snapshot_ia_rdata_part0[10]), .A2(o_sa_snapshot_ia_wdata_part1[10]), .A3(o_sa_snapshot_ia_wdata_part0[10]), .Z(n555));
Q_MX04 U836 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[10]), .A1(o_sa_count_ia_wdata_part1[10]), .A2(o_sa_count_ia_wdata_part0[10]), .A3(i_sa_count_ia_capability[10]), .Z(n556));
Q_MX04 U837 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[10]), .A1(i_sa_global_ctrl[10]), .A2(i_idle_components[10]), .A3(i_sa_count_ia_rdata_part1[10]), .Z(n557));
Q_MX02 U838 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[10]), .A1(o_sa_ctrl_ia_wdata_part0[10]), .Z(n558));
Q_AN02 U839 ( .A0(n4328), .A1(o_kdf_test_key_size_config[10]), .Z(n559));
Q_MX02 U840 ( .S(n4329), .A0(n559), .A1(n558), .Z(n560));
Q_MX04 U841 ( .S0(n4330), .S1(n4326), .A0(n560), .A1(n557), .A2(n556), .A3(n555), .Z(n561));
Q_MX02 U842 ( .S(n4331), .A0(n561), .A1(n554), .Z(r32_mux_8_data[10]));
Q_MX04 U843 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[11]), .A1(i_regs_sa_ctrl[11]), .A2(i_im_consumed[11]), .A3(i_im_available[11]), .Z(n562));
Q_MX04 U844 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[11]), .A1(i_sa_snapshot_ia_rdata_part0[11]), .A2(o_sa_snapshot_ia_wdata_part1[11]), .A3(o_sa_snapshot_ia_wdata_part0[11]), .Z(n563));
Q_MX04 U845 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[11]), .A1(o_sa_count_ia_wdata_part1[11]), .A2(o_sa_count_ia_wdata_part0[11]), .A3(i_sa_count_ia_capability[11]), .Z(n564));
Q_MX04 U846 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[11]), .A1(i_sa_global_ctrl[11]), .A2(i_idle_components[11]), .A3(i_sa_count_ia_rdata_part1[11]), .Z(n565));
Q_MX02 U847 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[11]), .A1(o_sa_ctrl_ia_wdata_part0[11]), .Z(n566));
Q_AN02 U848 ( .A0(n4328), .A1(o_kdf_test_key_size_config[11]), .Z(n567));
Q_MX02 U849 ( .S(n4329), .A0(n567), .A1(n566), .Z(n568));
Q_MX04 U850 ( .S0(n4330), .S1(n4326), .A0(n568), .A1(n565), .A2(n564), .A3(n563), .Z(n569));
Q_MX02 U851 ( .S(n4331), .A0(n569), .A1(n562), .Z(r32_mux_8_data[11]));
Q_MX04 U852 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[12]), .A1(i_regs_sa_ctrl[12]), .A2(i_im_consumed[12]), .A3(i_im_available[12]), .Z(n570));
Q_MX04 U853 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[12]), .A1(i_sa_snapshot_ia_rdata_part0[12]), .A2(o_sa_snapshot_ia_wdata_part1[12]), .A3(o_sa_snapshot_ia_wdata_part0[12]), .Z(n571));
Q_MX04 U854 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[12]), .A1(o_sa_count_ia_wdata_part1[12]), .A2(o_sa_count_ia_wdata_part0[12]), .A3(i_sa_count_ia_capability[12]), .Z(n572));
Q_MX04 U855 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[12]), .A1(i_sa_global_ctrl[12]), .A2(i_idle_components[12]), .A3(i_sa_count_ia_rdata_part1[12]), .Z(n573));
Q_MX02 U856 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[12]), .A1(o_sa_ctrl_ia_wdata_part0[12]), .Z(n574));
Q_AN02 U857 ( .A0(n4328), .A1(o_kdf_test_key_size_config[12]), .Z(n575));
Q_MX02 U858 ( .S(n4329), .A0(n575), .A1(n574), .Z(n576));
Q_MX04 U859 ( .S0(n4330), .S1(n4326), .A0(n576), .A1(n573), .A2(n572), .A3(n571), .Z(n577));
Q_MX02 U860 ( .S(n4331), .A0(n577), .A1(n570), .Z(r32_mux_8_data[12]));
Q_MX04 U861 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[13]), .A1(i_regs_sa_ctrl[13]), .A2(i_im_consumed[13]), .A3(i_im_available[13]), .Z(n578));
Q_MX04 U862 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[13]), .A1(i_sa_snapshot_ia_rdata_part0[13]), .A2(o_sa_snapshot_ia_wdata_part1[13]), .A3(o_sa_snapshot_ia_wdata_part0[13]), .Z(n579));
Q_MX04 U863 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[13]), .A1(o_sa_count_ia_wdata_part1[13]), .A2(o_sa_count_ia_wdata_part0[13]), .A3(i_sa_count_ia_capability[13]), .Z(n580));
Q_MX04 U864 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[13]), .A1(i_sa_global_ctrl[13]), .A2(i_idle_components[13]), .A3(i_sa_count_ia_rdata_part1[13]), .Z(n581));
Q_MX02 U865 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[13]), .A1(o_sa_ctrl_ia_wdata_part0[13]), .Z(n582));
Q_AN02 U866 ( .A0(n4328), .A1(o_kdf_test_key_size_config[13]), .Z(n583));
Q_MX02 U867 ( .S(n4329), .A0(n583), .A1(n582), .Z(n584));
Q_MX04 U868 ( .S0(n4330), .S1(n4326), .A0(n584), .A1(n581), .A2(n580), .A3(n579), .Z(n585));
Q_MX02 U869 ( .S(n4331), .A0(n585), .A1(n578), .Z(r32_mux_8_data[13]));
Q_MX04 U870 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[14]), .A1(i_regs_sa_ctrl[14]), .A2(i_im_consumed[14]), .A3(i_im_available[14]), .Z(n586));
Q_MX04 U871 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[14]), .A1(i_sa_snapshot_ia_rdata_part0[14]), .A2(o_sa_snapshot_ia_wdata_part1[14]), .A3(o_sa_snapshot_ia_wdata_part0[14]), .Z(n587));
Q_MX04 U872 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[14]), .A1(o_sa_count_ia_wdata_part1[14]), .A2(o_sa_count_ia_wdata_part0[14]), .A3(i_sa_count_ia_capability[14]), .Z(n588));
Q_MX04 U873 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[14]), .A1(i_sa_global_ctrl[14]), .A2(i_idle_components[14]), .A3(i_sa_count_ia_rdata_part1[14]), .Z(n589));
Q_MX02 U874 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[14]), .A1(o_sa_ctrl_ia_wdata_part0[14]), .Z(n590));
Q_AN02 U875 ( .A0(n4328), .A1(o_kdf_test_key_size_config[14]), .Z(n591));
Q_MX02 U876 ( .S(n4329), .A0(n591), .A1(n590), .Z(n592));
Q_MX04 U877 ( .S0(n4330), .S1(n4326), .A0(n592), .A1(n589), .A2(n588), .A3(n587), .Z(n593));
Q_MX02 U878 ( .S(n4331), .A0(n593), .A1(n586), .Z(r32_mux_8_data[14]));
Q_MX04 U879 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_capability[15]), .A1(i_regs_sa_ctrl[15]), .A2(i_im_consumed[15]), .A3(i_im_available[15]), .Z(n594));
Q_MX04 U880 ( .S0(n4328), .S1(n4329), .A0(i_sa_snapshot_ia_rdata_part1[15]), .A1(i_sa_snapshot_ia_rdata_part0[15]), .A2(o_sa_snapshot_ia_wdata_part1[15]), .A3(o_sa_snapshot_ia_wdata_part0[15]), .Z(n595));
Q_MX04 U881 ( .S0(n4328), .S1(n4329), .A0(i_sa_count_ia_rdata_part0[15]), .A1(o_sa_count_ia_wdata_part1[15]), .A2(o_sa_count_ia_wdata_part0[15]), .A3(i_sa_count_ia_capability[15]), .Z(n596));
Q_MX04 U882 ( .S0(n4328), .S1(n4329), .A0(i_sa_ctrl_ia_capability[15]), .A1(i_sa_global_ctrl[15]), .A2(i_idle_components[15]), .A3(i_sa_count_ia_rdata_part1[15]), .Z(n597));
Q_MX02 U883 ( .S(n4328), .A0(i_sa_ctrl_ia_rdata_part0[15]), .A1(o_sa_ctrl_ia_wdata_part0[15]), .Z(n598));
Q_AN02 U884 ( .A0(n4328), .A1(o_kdf_test_key_size_config[15]), .Z(n599));
Q_MX02 U885 ( .S(n4329), .A0(n599), .A1(n598), .Z(n600));
Q_MX04 U886 ( .S0(n4330), .S1(n4326), .A0(n600), .A1(n597), .A2(n596), .A3(n595), .Z(n601));
Q_MX02 U887 ( .S(n4331), .A0(n601), .A1(n594), .Z(r32_mux_8_data[15]));
Q_MX03 U888 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[16]), .A1(o_sa_snapshot_ia_wdata_part0[16]), .A2(i_regs_sa_ctrl[16]), .Z(n602));
Q_MX04 U889 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[16]), .A1(o_sa_count_ia_wdata_part0[16]), .A2(i_sa_snapshot_ia_rdata_part1[16]), .A3(i_sa_snapshot_ia_rdata_part0[16]), .Z(n603));
Q_MX02 U890 ( .S(n4334), .A0(n603), .A1(n602), .Z(n604));
Q_MX04 U891 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[16]), .A1(i_idle_components[16]), .A2(i_sa_count_ia_rdata_part1[16]), .A3(i_sa_count_ia_rdata_part0[16]), .Z(n605));
Q_MX02 U892 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[16]), .A1(o_sa_ctrl_ia_wdata_part0[16]), .Z(n606));
Q_AN02 U893 ( .A0(n4332), .A1(o_kdf_test_key_size_config[16]), .Z(n607));
Q_MX03 U894 ( .S0(n4333), .S1(n4334), .A0(n607), .A1(n606), .A2(n605), .Z(n608));
Q_MX02 U895 ( .S(n4335), .A0(n608), .A1(n604), .Z(r32_mux_8_data[16]));
Q_MX03 U896 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[17]), .A1(o_sa_snapshot_ia_wdata_part0[17]), .A2(i_regs_sa_ctrl[17]), .Z(n609));
Q_MX04 U897 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[17]), .A1(o_sa_count_ia_wdata_part0[17]), .A2(i_sa_snapshot_ia_rdata_part1[17]), .A3(i_sa_snapshot_ia_rdata_part0[17]), .Z(n610));
Q_MX02 U898 ( .S(n4334), .A0(n610), .A1(n609), .Z(n611));
Q_MX04 U899 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[17]), .A1(i_idle_components[17]), .A2(i_sa_count_ia_rdata_part1[17]), .A3(i_sa_count_ia_rdata_part0[17]), .Z(n612));
Q_MX02 U900 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[17]), .A1(o_sa_ctrl_ia_wdata_part0[17]), .Z(n613));
Q_AN02 U901 ( .A0(n4332), .A1(o_kdf_test_key_size_config[17]), .Z(n614));
Q_MX03 U902 ( .S0(n4333), .S1(n4334), .A0(n614), .A1(n613), .A2(n612), .Z(n615));
Q_MX02 U903 ( .S(n4335), .A0(n615), .A1(n611), .Z(r32_mux_8_data[17]));
Q_MX03 U904 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[18]), .A1(o_sa_snapshot_ia_wdata_part0[18]), .A2(i_regs_sa_ctrl[18]), .Z(n616));
Q_MX04 U905 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[18]), .A1(o_sa_count_ia_wdata_part0[18]), .A2(i_sa_snapshot_ia_rdata_part1[18]), .A3(i_sa_snapshot_ia_rdata_part0[18]), .Z(n617));
Q_MX02 U906 ( .S(n4334), .A0(n617), .A1(n616), .Z(n618));
Q_MX04 U907 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[18]), .A1(i_idle_components[18]), .A2(i_sa_count_ia_rdata_part1[18]), .A3(i_sa_count_ia_rdata_part0[18]), .Z(n619));
Q_MX02 U908 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[18]), .A1(o_sa_ctrl_ia_wdata_part0[18]), .Z(n620));
Q_AN02 U909 ( .A0(n4332), .A1(o_kdf_test_key_size_config[18]), .Z(n621));
Q_MX03 U910 ( .S0(n4333), .S1(n4334), .A0(n621), .A1(n620), .A2(n619), .Z(n622));
Q_MX02 U911 ( .S(n4335), .A0(n622), .A1(n618), .Z(r32_mux_8_data[18]));
Q_MX03 U912 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[19]), .A1(o_sa_snapshot_ia_wdata_part0[19]), .A2(i_regs_sa_ctrl[19]), .Z(n623));
Q_MX04 U913 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[19]), .A1(o_sa_count_ia_wdata_part0[19]), .A2(i_sa_snapshot_ia_rdata_part1[19]), .A3(i_sa_snapshot_ia_rdata_part0[19]), .Z(n624));
Q_MX02 U914 ( .S(n4334), .A0(n624), .A1(n623), .Z(n625));
Q_MX04 U915 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[19]), .A1(i_idle_components[19]), .A2(i_sa_count_ia_rdata_part1[19]), .A3(i_sa_count_ia_rdata_part0[19]), .Z(n626));
Q_MX02 U916 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[19]), .A1(o_sa_ctrl_ia_wdata_part0[19]), .Z(n627));
Q_AN02 U917 ( .A0(n4332), .A1(o_kdf_test_key_size_config[19]), .Z(n628));
Q_MX03 U918 ( .S0(n4333), .S1(n4334), .A0(n628), .A1(n627), .A2(n626), .Z(n629));
Q_MX02 U919 ( .S(n4335), .A0(n629), .A1(n625), .Z(r32_mux_8_data[19]));
Q_MX03 U920 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[20]), .A1(o_sa_snapshot_ia_wdata_part0[20]), .A2(i_regs_sa_ctrl[20]), .Z(n630));
Q_MX04 U921 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[20]), .A1(o_sa_count_ia_wdata_part0[20]), .A2(i_sa_snapshot_ia_rdata_part1[20]), .A3(i_sa_snapshot_ia_rdata_part0[20]), .Z(n631));
Q_MX02 U922 ( .S(n4334), .A0(n631), .A1(n630), .Z(n632));
Q_MX04 U923 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[20]), .A1(i_idle_components[20]), .A2(i_sa_count_ia_rdata_part1[20]), .A3(i_sa_count_ia_rdata_part0[20]), .Z(n633));
Q_MX02 U924 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[20]), .A1(o_sa_ctrl_ia_wdata_part0[20]), .Z(n634));
Q_AN02 U925 ( .A0(n4332), .A1(o_kdf_test_key_size_config[20]), .Z(n635));
Q_MX03 U926 ( .S0(n4333), .S1(n4334), .A0(n635), .A1(n634), .A2(n633), .Z(n636));
Q_MX02 U927 ( .S(n4335), .A0(n636), .A1(n632), .Z(r32_mux_8_data[20]));
Q_MX03 U928 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[21]), .A1(o_sa_snapshot_ia_wdata_part0[21]), .A2(i_regs_sa_ctrl[21]), .Z(n637));
Q_MX04 U929 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[21]), .A1(o_sa_count_ia_wdata_part0[21]), .A2(i_sa_snapshot_ia_rdata_part1[21]), .A3(i_sa_snapshot_ia_rdata_part0[21]), .Z(n638));
Q_MX02 U930 ( .S(n4334), .A0(n638), .A1(n637), .Z(n639));
Q_MX04 U931 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[21]), .A1(i_idle_components[21]), .A2(i_sa_count_ia_rdata_part1[21]), .A3(i_sa_count_ia_rdata_part0[21]), .Z(n640));
Q_MX02 U932 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[21]), .A1(o_sa_ctrl_ia_wdata_part0[21]), .Z(n641));
Q_AN02 U933 ( .A0(n4332), .A1(o_kdf_test_key_size_config[21]), .Z(n642));
Q_MX03 U934 ( .S0(n4333), .S1(n4334), .A0(n642), .A1(n641), .A2(n640), .Z(n643));
Q_MX02 U935 ( .S(n4335), .A0(n643), .A1(n639), .Z(r32_mux_8_data[21]));
Q_MX03 U936 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[22]), .A1(o_sa_snapshot_ia_wdata_part0[22]), .A2(i_regs_sa_ctrl[22]), .Z(n644));
Q_MX04 U937 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[22]), .A1(o_sa_count_ia_wdata_part0[22]), .A2(i_sa_snapshot_ia_rdata_part1[22]), .A3(i_sa_snapshot_ia_rdata_part0[22]), .Z(n645));
Q_MX02 U938 ( .S(n4334), .A0(n645), .A1(n644), .Z(n646));
Q_MX04 U939 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[22]), .A1(i_idle_components[22]), .A2(i_sa_count_ia_rdata_part1[22]), .A3(i_sa_count_ia_rdata_part0[22]), .Z(n647));
Q_MX02 U940 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[22]), .A1(o_sa_ctrl_ia_wdata_part0[22]), .Z(n648));
Q_AN02 U941 ( .A0(n4332), .A1(o_kdf_test_key_size_config[22]), .Z(n649));
Q_MX03 U942 ( .S0(n4333), .S1(n4334), .A0(n649), .A1(n648), .A2(n647), .Z(n650));
Q_MX02 U943 ( .S(n4335), .A0(n650), .A1(n646), .Z(r32_mux_8_data[22]));
Q_MX03 U944 ( .S0(n4332), .S1(n4333), .A0(o_sa_snapshot_ia_wdata_part1[23]), .A1(o_sa_snapshot_ia_wdata_part0[23]), .A2(i_regs_sa_ctrl[23]), .Z(n651));
Q_MX04 U945 ( .S0(n4332), .S1(n4333), .A0(o_sa_count_ia_wdata_part1[23]), .A1(o_sa_count_ia_wdata_part0[23]), .A2(i_sa_snapshot_ia_rdata_part1[23]), .A3(i_sa_snapshot_ia_rdata_part0[23]), .Z(n652));
Q_MX02 U946 ( .S(n4334), .A0(n652), .A1(n651), .Z(n653));
Q_MX04 U947 ( .S0(n4332), .S1(n4333), .A0(i_sa_global_ctrl[23]), .A1(i_idle_components[23]), .A2(i_sa_count_ia_rdata_part1[23]), .A3(i_sa_count_ia_rdata_part0[23]), .Z(n654));
Q_MX02 U948 ( .S(n4332), .A0(i_sa_ctrl_ia_rdata_part0[23]), .A1(o_sa_ctrl_ia_wdata_part0[23]), .Z(n655));
Q_AN02 U949 ( .A0(n4332), .A1(o_kdf_test_key_size_config[23]), .Z(n656));
Q_MX03 U950 ( .S0(n4333), .S1(n4334), .A0(n656), .A1(n655), .A2(n654), .Z(n657));
Q_MX02 U951 ( .S(n4335), .A0(n657), .A1(n653), .Z(r32_mux_8_data[23]));
Q_MX02 U952 ( .S(n4336), .A0(i_sa_snapshot_ia_status[5]), .A1(i_regs_sa_ctrl[24]), .Z(n658));
Q_MX04 U953 ( .S0(n4336), .S1(n4337), .A0(i_sa_snapshot_ia_rdata_part1[24]), .A1(i_sa_snapshot_ia_rdata_part0[24]), .A2(o_sa_snapshot_ia_wdata_part1[24]), .A3(o_sa_snapshot_ia_wdata_part0[24]), .Z(n659));
Q_MX04 U954 ( .S0(n4336), .S1(n4337), .A0(i_sa_count_ia_rdata_part0[24]), .A1(o_sa_count_ia_wdata_part1[24]), .A2(o_sa_count_ia_wdata_part0[24]), .A3(i_sa_count_ia_status[5]), .Z(n660));
Q_MX04 U955 ( .S0(n4336), .S1(n4337), .A0(i_sa_ctrl_ia_status[5]), .A1(i_sa_global_ctrl[24]), .A2(i_idle_components[24]), .A3(i_sa_count_ia_rdata_part1[24]), .Z(n661));
Q_MX02 U956 ( .S(n4336), .A0(i_sa_ctrl_ia_rdata_part0[24]), .A1(o_sa_ctrl_ia_wdata_part0[24]), .Z(n662));
Q_AN02 U957 ( .A0(n4336), .A1(o_kdf_test_key_size_config[24]), .Z(n663));
Q_MX02 U958 ( .S(n4337), .A0(n663), .A1(n662), .Z(n664));
Q_MX04 U959 ( .S0(n4338), .S1(n4339), .A0(n664), .A1(n661), .A2(n660), .A3(n659), .Z(n665));
Q_MX02 U960 ( .S(n4340), .A0(n665), .A1(n658), .Z(r32_mux_8_data[24]));
Q_MX02 U961 ( .S(n4336), .A0(i_sa_snapshot_ia_status[6]), .A1(i_regs_sa_ctrl[25]), .Z(n666));
Q_MX04 U962 ( .S0(n4336), .S1(n4337), .A0(i_sa_snapshot_ia_rdata_part1[25]), .A1(i_sa_snapshot_ia_rdata_part0[25]), .A2(o_sa_snapshot_ia_wdata_part1[25]), .A3(o_sa_snapshot_ia_wdata_part0[25]), .Z(n667));
Q_MX04 U963 ( .S0(n4336), .S1(n4337), .A0(i_sa_count_ia_rdata_part0[25]), .A1(o_sa_count_ia_wdata_part1[25]), .A2(o_sa_count_ia_wdata_part0[25]), .A3(i_sa_count_ia_status[6]), .Z(n668));
Q_MX04 U964 ( .S0(n4336), .S1(n4337), .A0(i_sa_ctrl_ia_status[6]), .A1(i_sa_global_ctrl[25]), .A2(i_idle_components[25]), .A3(i_sa_count_ia_rdata_part1[25]), .Z(n669));
Q_MX02 U965 ( .S(n4336), .A0(i_sa_ctrl_ia_rdata_part0[25]), .A1(o_sa_ctrl_ia_wdata_part0[25]), .Z(n670));
Q_AN02 U966 ( .A0(n4336), .A1(o_kdf_test_key_size_config[25]), .Z(n671));
Q_MX02 U967 ( .S(n4337), .A0(n671), .A1(n670), .Z(n672));
Q_MX04 U968 ( .S0(n4338), .S1(n4339), .A0(n672), .A1(n669), .A2(n668), .A3(n667), .Z(n673));
Q_MX02 U969 ( .S(n4340), .A0(n673), .A1(n666), .Z(r32_mux_8_data[25]));
Q_MX02 U970 ( .S(n4336), .A0(i_sa_snapshot_ia_status[7]), .A1(i_regs_sa_ctrl[26]), .Z(n674));
Q_MX04 U971 ( .S0(n4336), .S1(n4337), .A0(i_sa_snapshot_ia_rdata_part1[26]), .A1(i_sa_snapshot_ia_rdata_part0[26]), .A2(o_sa_snapshot_ia_wdata_part1[26]), .A3(o_sa_snapshot_ia_wdata_part0[26]), .Z(n675));
Q_MX04 U972 ( .S0(n4336), .S1(n4337), .A0(i_sa_count_ia_rdata_part0[26]), .A1(o_sa_count_ia_wdata_part1[26]), .A2(o_sa_count_ia_wdata_part0[26]), .A3(i_sa_count_ia_status[7]), .Z(n676));
Q_MX04 U973 ( .S0(n4336), .S1(n4337), .A0(i_sa_ctrl_ia_status[7]), .A1(i_sa_global_ctrl[26]), .A2(i_idle_components[26]), .A3(i_sa_count_ia_rdata_part1[26]), .Z(n677));
Q_MX02 U974 ( .S(n4336), .A0(i_sa_ctrl_ia_rdata_part0[26]), .A1(o_sa_ctrl_ia_wdata_part0[26]), .Z(n678));
Q_AN02 U975 ( .A0(n4336), .A1(o_kdf_test_key_size_config[26]), .Z(n679));
Q_MX02 U976 ( .S(n4337), .A0(n679), .A1(n678), .Z(n680));
Q_MX04 U977 ( .S0(n4338), .S1(n4339), .A0(n680), .A1(n677), .A2(n676), .A3(n675), .Z(n681));
Q_MX02 U978 ( .S(n4340), .A0(n681), .A1(n674), .Z(r32_mux_8_data[26]));
Q_MX02 U979 ( .S(n4336), .A0(i_sa_snapshot_ia_status[8]), .A1(i_regs_sa_ctrl[27]), .Z(n682));
Q_MX04 U980 ( .S0(n4336), .S1(n4337), .A0(i_sa_snapshot_ia_rdata_part1[27]), .A1(i_sa_snapshot_ia_rdata_part0[27]), .A2(o_sa_snapshot_ia_wdata_part1[27]), .A3(o_sa_snapshot_ia_wdata_part0[27]), .Z(n683));
Q_MX04 U981 ( .S0(n4336), .S1(n4337), .A0(i_sa_count_ia_rdata_part0[27]), .A1(o_sa_count_ia_wdata_part1[27]), .A2(o_sa_count_ia_wdata_part0[27]), .A3(i_sa_count_ia_status[8]), .Z(n684));
Q_MX04 U982 ( .S0(n4336), .S1(n4337), .A0(i_sa_ctrl_ia_status[8]), .A1(i_sa_global_ctrl[27]), .A2(i_idle_components[27]), .A3(i_sa_count_ia_rdata_part1[27]), .Z(n685));
Q_MX02 U983 ( .S(n4336), .A0(i_sa_ctrl_ia_rdata_part0[27]), .A1(o_sa_ctrl_ia_wdata_part0[27]), .Z(n686));
Q_AN02 U984 ( .A0(n4336), .A1(o_kdf_test_key_size_config[27]), .Z(n687));
Q_MX02 U985 ( .S(n4337), .A0(n687), .A1(n686), .Z(n688));
Q_MX04 U986 ( .S0(n4338), .S1(n4339), .A0(n688), .A1(n685), .A2(n684), .A3(n683), .Z(n689));
Q_MX02 U987 ( .S(n4340), .A0(n689), .A1(n682), .Z(r32_mux_8_data[27]));
Q_MX08 U988 ( .S0(n4341), .S1(n4342), .S2(n4343), .A0(i_sa_snapshot_ia_rdata_part1[28]), .A1(i_sa_snapshot_ia_rdata_part0[28]), .A2(o_sa_snapshot_ia_config[5]), .A3(o_sa_snapshot_ia_wdata_part1[28]), .A4(o_sa_snapshot_ia_wdata_part0[28]), .A5(i_sa_snapshot_ia_status[9]), .A6(i_sa_snapshot_ia_capability[16]), .A7(i_regs_sa_ctrl[28]), .Z(n690));
Q_MX04 U989 ( .S0(n4341), .S1(n4342), .A0(o_sa_count_ia_wdata_part1[28]), .A1(o_sa_count_ia_wdata_part0[28]), .A2(i_sa_count_ia_status[9]), .A3(i_sa_count_ia_capability[16]), .Z(n691));
Q_MX04 U990 ( .S0(n4341), .S1(n4342), .A0(i_idle_components[28]), .A1(i_sa_count_ia_rdata_part1[28]), .A2(i_sa_count_ia_rdata_part0[28]), .A3(o_sa_count_ia_config[5]), .Z(n692));
Q_MX04 U991 ( .S0(n4341), .S1(n4342), .A0(o_sa_ctrl_ia_wdata_part0[28]), .A1(i_sa_ctrl_ia_status[9]), .A2(i_sa_ctrl_ia_capability[16]), .A3(i_sa_global_ctrl[28]), .Z(n693));
Q_MX02 U992 ( .S(n4341), .A0(i_sa_ctrl_ia_rdata_part0[28]), .A1(o_sa_ctrl_ia_config[5]), .Z(n694));
Q_AN02 U993 ( .A0(n4341), .A1(o_kdf_test_key_size_config[28]), .Z(n695));
Q_MX02 U994 ( .S(n4342), .A0(n695), .A1(n694), .Z(n696));
Q_MX04 U995 ( .S0(n4343), .S1(n4344), .A0(n696), .A1(n693), .A2(n692), .A3(n691), .Z(n697));
Q_MX02 U996 ( .S(n4345), .A0(n697), .A1(n690), .Z(r32_mux_8_data[28]));
Q_MX08 U997 ( .S0(n4341), .S1(n4342), .S2(n4343), .A0(i_sa_snapshot_ia_rdata_part1[29]), .A1(i_sa_snapshot_ia_rdata_part0[29]), .A2(o_sa_snapshot_ia_config[6]), .A3(o_sa_snapshot_ia_wdata_part1[29]), .A4(o_sa_snapshot_ia_wdata_part0[29]), .A5(i_sa_snapshot_ia_status[10]), .A6(i_sa_snapshot_ia_capability[17]), .A7(i_regs_sa_ctrl[29]), .Z(n698));
Q_MX04 U998 ( .S0(n4341), .S1(n4342), .A0(o_sa_count_ia_wdata_part1[29]), .A1(o_sa_count_ia_wdata_part0[29]), .A2(i_sa_count_ia_status[10]), .A3(i_sa_count_ia_capability[17]), .Z(n699));
Q_MX04 U999 ( .S0(n4341), .S1(n4342), .A0(i_idle_components[29]), .A1(i_sa_count_ia_rdata_part1[29]), .A2(i_sa_count_ia_rdata_part0[29]), .A3(o_sa_count_ia_config[6]), .Z(n700));
Q_MX04 U1000 ( .S0(n4341), .S1(n4342), .A0(o_sa_ctrl_ia_wdata_part0[29]), .A1(i_sa_ctrl_ia_status[10]), .A2(i_sa_ctrl_ia_capability[17]), .A3(i_sa_global_ctrl[29]), .Z(n701));
Q_MX02 U1001 ( .S(n4341), .A0(i_sa_ctrl_ia_rdata_part0[29]), .A1(o_sa_ctrl_ia_config[6]), .Z(n702));
Q_AN02 U1002 ( .A0(n4341), .A1(o_kdf_test_key_size_config[29]), .Z(n703));
Q_MX02 U1003 ( .S(n4342), .A0(n703), .A1(n702), .Z(n704));
Q_MX04 U1004 ( .S0(n4343), .S1(n4344), .A0(n704), .A1(n701), .A2(n700), .A3(n699), .Z(n705));
Q_MX02 U1005 ( .S(n4345), .A0(n705), .A1(n698), .Z(r32_mux_8_data[29]));
Q_MX08 U1006 ( .S0(n4341), .S1(n4342), .S2(n4343), .A0(i_sa_snapshot_ia_rdata_part1[30]), .A1(i_sa_snapshot_ia_rdata_part0[30]), .A2(o_sa_snapshot_ia_config[7]), .A3(o_sa_snapshot_ia_wdata_part1[30]), .A4(o_sa_snapshot_ia_wdata_part0[30]), .A5(i_sa_snapshot_ia_status[11]), .A6(i_sa_snapshot_ia_capability[18]), .A7(i_regs_sa_ctrl[30]), .Z(n706));
Q_MX04 U1007 ( .S0(n4341), .S1(n4342), .A0(o_sa_count_ia_wdata_part1[30]), .A1(o_sa_count_ia_wdata_part0[30]), .A2(i_sa_count_ia_status[11]), .A3(i_sa_count_ia_capability[18]), .Z(n707));
Q_MX04 U1008 ( .S0(n4341), .S1(n4342), .A0(i_idle_components[30]), .A1(i_sa_count_ia_rdata_part1[30]), .A2(i_sa_count_ia_rdata_part0[30]), .A3(o_sa_count_ia_config[7]), .Z(n708));
Q_MX04 U1009 ( .S0(n4341), .S1(n4342), .A0(o_sa_ctrl_ia_wdata_part0[30]), .A1(i_sa_ctrl_ia_status[11]), .A2(i_sa_ctrl_ia_capability[18]), .A3(i_sa_global_ctrl[30]), .Z(n709));
Q_MX02 U1010 ( .S(n4341), .A0(i_sa_ctrl_ia_rdata_part0[30]), .A1(o_sa_ctrl_ia_config[7]), .Z(n710));
Q_AN02 U1011 ( .A0(n4341), .A1(o_kdf_test_key_size_config[30]), .Z(n711));
Q_MX02 U1012 ( .S(n4342), .A0(n711), .A1(n710), .Z(n712));
Q_MX04 U1013 ( .S0(n4343), .S1(n4344), .A0(n712), .A1(n709), .A2(n708), .A3(n707), .Z(n713));
Q_MX02 U1014 ( .S(n4345), .A0(n713), .A1(n706), .Z(r32_mux_8_data[30]));
Q_MX08 U1015 ( .S0(n4341), .S1(n4342), .S2(n4343), .A0(i_sa_snapshot_ia_rdata_part1[31]), .A1(i_sa_snapshot_ia_rdata_part0[31]), .A2(o_sa_snapshot_ia_config[8]), .A3(o_sa_snapshot_ia_wdata_part1[31]), .A4(o_sa_snapshot_ia_wdata_part0[31]), .A5(i_sa_snapshot_ia_status[12]), .A6(i_sa_snapshot_ia_capability[19]), .A7(i_regs_sa_ctrl[31]), .Z(n714));
Q_MX04 U1016 ( .S0(n4341), .S1(n4342), .A0(o_sa_count_ia_wdata_part1[31]), .A1(o_sa_count_ia_wdata_part0[31]), .A2(i_sa_count_ia_status[12]), .A3(i_sa_count_ia_capability[19]), .Z(n715));
Q_MX04 U1017 ( .S0(n4341), .S1(n4342), .A0(i_idle_components[31]), .A1(i_sa_count_ia_rdata_part1[31]), .A2(i_sa_count_ia_rdata_part0[31]), .A3(o_sa_count_ia_config[8]), .Z(n716));
Q_MX04 U1018 ( .S0(n4341), .S1(n4342), .A0(o_sa_ctrl_ia_wdata_part0[31]), .A1(i_sa_ctrl_ia_status[12]), .A2(i_sa_ctrl_ia_capability[19]), .A3(i_sa_global_ctrl[31]), .Z(n717));
Q_MX02 U1019 ( .S(n4341), .A0(i_sa_ctrl_ia_rdata_part0[31]), .A1(o_sa_ctrl_ia_config[8]), .Z(n718));
Q_AN02 U1020 ( .A0(n4341), .A1(o_kdf_test_key_size_config[31]), .Z(n719));
Q_MX02 U1021 ( .S(n4342), .A0(n719), .A1(n718), .Z(n720));
Q_MX04 U1022 ( .S0(n4343), .S1(n4344), .A0(n720), .A1(n717), .A2(n716), .A3(n715), .Z(n721));
Q_MX02 U1023 ( .S(n4345), .A0(n721), .A1(n714), .Z(r32_mux_8_data[31]));
Q_MX03 U1024 ( .S0(n4346), .S1(n4347), .A0(o_kdf_drbg_seed_1_reseed_interval_0[0]), .A1(o_kdf_drbg_seed_1_state_value_127_96[0]), .A2(o_kdf_drbg_seed_1_state_value_95_64[0]), .Z(n722));
Q_MX04 U1025 ( .S0(n4346), .S1(n4347), .A0(i_engine_sticky_status[0]), .A1(o_interrupt_mask[0]), .A2(i_interrupt_status[0]), .A3(o_kdf_drbg_seed_1_reseed_interval_1[0]), .Z(n723));
Q_MX02 U1026 ( .S(n4348), .A0(n723), .A1(n722), .Z(n724));
Q_MX08 U1027 ( .S0(n4346), .S1(n4347), .S2(n4348), .A0(i_bimc_eccpar_debug[0]), .A1(i_bimc_memid[0]), .A2(i_bimc_global_config[0]), .A3(i_bimc_parity_error_cnt[0]), .A4(i_bimc_ecc_correctable_error_cnt[0]), .A5(i_bimc_ecc_uncorrectable_error_cnt[0]), .A6(o_bimc_monitor_mask[0]), .A7(i_bimc_monitor[0]), .Z(n725));
Q_MX02 U1028 ( .S(n4349), .A0(n725), .A1(n724), .Z(n726));
Q_MX04 U1029 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxcmd2[0]), .A1(o_bimc_cmd0[0]), .A2(o_bimc_cmd1[0]), .A3(i_bimc_cmd2[0]), .Z(n727));
Q_MX04 U1030 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxrsp1[0]), .A1(i_bimc_rxrsp2[0]), .A2(i_bimc_rxcmd0[0]), .A3(i_bimc_rxcmd1[0]), .Z(n728));
Q_MX04 U1031 ( .S0(n4346), .S1(n4347), .A0(i_bimc_pollrsp0[0]), .A1(i_bimc_pollrsp1[0]), .A2(i_bimc_pollrsp2[0]), .A3(i_bimc_rxrsp0[0]), .Z(n729));
Q_MX02 U1032 ( .S(n4346), .A0(i_bimc_dbgcmd1[0]), .A1(i_bimc_dbgcmd2[0]), .Z(n730));
Q_AN02 U1033 ( .A0(n4346), .A1(i_bimc_dbgcmd0[0]), .Z(n731));
Q_MX02 U1034 ( .S(n4347), .A0(n731), .A1(n730), .Z(n732));
Q_MX04 U1035 ( .S0(n4348), .S1(n4349), .A0(n732), .A1(n729), .A2(n728), .A3(n727), .Z(n733));
Q_MX02 U1036 ( .S(n4350), .A0(n733), .A1(n726), .Z(r32_mux_7_data[0]));
Q_MX03 U1037 ( .S0(n4346), .S1(n4347), .A0(o_kdf_drbg_seed_1_reseed_interval_0[1]), .A1(o_kdf_drbg_seed_1_state_value_127_96[1]), .A2(o_kdf_drbg_seed_1_state_value_95_64[1]), .Z(n734));
Q_MX04 U1038 ( .S0(n4346), .S1(n4347), .A0(i_engine_sticky_status[1]), .A1(o_interrupt_mask[1]), .A2(i_interrupt_status[1]), .A3(o_kdf_drbg_seed_1_reseed_interval_1[1]), .Z(n735));
Q_MX02 U1039 ( .S(n4348), .A0(n735), .A1(n734), .Z(n736));
Q_MX08 U1040 ( .S0(n4346), .S1(n4347), .S2(n4348), .A0(i_bimc_eccpar_debug[1]), .A1(i_bimc_memid[1]), .A2(i_bimc_global_config[1]), .A3(i_bimc_parity_error_cnt[1]), .A4(i_bimc_ecc_correctable_error_cnt[1]), .A5(i_bimc_ecc_uncorrectable_error_cnt[1]), .A6(o_bimc_monitor_mask[1]), .A7(i_bimc_monitor[1]), .Z(n737));
Q_MX02 U1041 ( .S(n4349), .A0(n737), .A1(n736), .Z(n738));
Q_MX04 U1042 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxcmd2[1]), .A1(o_bimc_cmd0[1]), .A2(o_bimc_cmd1[1]), .A3(i_bimc_cmd2[1]), .Z(n739));
Q_MX04 U1043 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxrsp1[1]), .A1(i_bimc_rxrsp2[1]), .A2(i_bimc_rxcmd0[1]), .A3(i_bimc_rxcmd1[1]), .Z(n740));
Q_MX04 U1044 ( .S0(n4346), .S1(n4347), .A0(i_bimc_pollrsp0[1]), .A1(i_bimc_pollrsp1[1]), .A2(i_bimc_pollrsp2[1]), .A3(i_bimc_rxrsp0[1]), .Z(n741));
Q_MX02 U1045 ( .S(n4346), .A0(i_bimc_dbgcmd1[1]), .A1(i_bimc_dbgcmd2[1]), .Z(n742));
Q_AN02 U1046 ( .A0(n4346), .A1(i_bimc_dbgcmd0[1]), .Z(n743));
Q_MX02 U1047 ( .S(n4347), .A0(n743), .A1(n742), .Z(n744));
Q_MX04 U1048 ( .S0(n4348), .S1(n4349), .A0(n744), .A1(n741), .A2(n740), .A3(n739), .Z(n745));
Q_MX02 U1049 ( .S(n4350), .A0(n745), .A1(n738), .Z(r32_mux_7_data[1]));
Q_MX03 U1050 ( .S0(n4346), .S1(n4347), .A0(o_kdf_drbg_seed_1_reseed_interval_0[2]), .A1(o_kdf_drbg_seed_1_state_value_127_96[2]), .A2(o_kdf_drbg_seed_1_state_value_95_64[2]), .Z(n746));
Q_MX04 U1051 ( .S0(n4346), .S1(n4347), .A0(i_engine_sticky_status[2]), .A1(o_interrupt_mask[2]), .A2(i_interrupt_status[2]), .A3(o_kdf_drbg_seed_1_reseed_interval_1[2]), .Z(n747));
Q_MX02 U1052 ( .S(n4348), .A0(n747), .A1(n746), .Z(n748));
Q_MX08 U1053 ( .S0(n4346), .S1(n4347), .S2(n4348), .A0(i_bimc_eccpar_debug[2]), .A1(i_bimc_memid[2]), .A2(i_bimc_global_config[2]), .A3(i_bimc_parity_error_cnt[2]), .A4(i_bimc_ecc_correctable_error_cnt[2]), .A5(i_bimc_ecc_uncorrectable_error_cnt[2]), .A6(o_bimc_monitor_mask[2]), .A7(i_bimc_monitor[2]), .Z(n749));
Q_MX02 U1054 ( .S(n4349), .A0(n749), .A1(n748), .Z(n750));
Q_MX04 U1055 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxcmd2[2]), .A1(o_bimc_cmd0[2]), .A2(o_bimc_cmd1[2]), .A3(i_bimc_cmd2[2]), .Z(n751));
Q_MX04 U1056 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxrsp1[2]), .A1(i_bimc_rxrsp2[2]), .A2(i_bimc_rxcmd0[2]), .A3(i_bimc_rxcmd1[2]), .Z(n752));
Q_MX04 U1057 ( .S0(n4346), .S1(n4347), .A0(i_bimc_pollrsp0[2]), .A1(i_bimc_pollrsp1[2]), .A2(i_bimc_pollrsp2[2]), .A3(i_bimc_rxrsp0[2]), .Z(n753));
Q_MX02 U1058 ( .S(n4346), .A0(i_bimc_dbgcmd1[2]), .A1(i_bimc_dbgcmd2[2]), .Z(n754));
Q_AN02 U1059 ( .A0(n4346), .A1(i_bimc_dbgcmd0[2]), .Z(n755));
Q_MX02 U1060 ( .S(n4347), .A0(n755), .A1(n754), .Z(n756));
Q_MX04 U1061 ( .S0(n4348), .S1(n4349), .A0(n756), .A1(n753), .A2(n752), .A3(n751), .Z(n757));
Q_MX02 U1062 ( .S(n4350), .A0(n757), .A1(n750), .Z(r32_mux_7_data[2]));
Q_MX03 U1063 ( .S0(n4346), .S1(n4347), .A0(o_kdf_drbg_seed_1_reseed_interval_0[3]), .A1(o_kdf_drbg_seed_1_state_value_127_96[3]), .A2(o_kdf_drbg_seed_1_state_value_95_64[3]), .Z(n758));
Q_MX04 U1064 ( .S0(n4346), .S1(n4347), .A0(i_engine_sticky_status[3]), .A1(o_interrupt_mask[3]), .A2(i_interrupt_status[3]), .A3(o_kdf_drbg_seed_1_reseed_interval_1[3]), .Z(n759));
Q_MX02 U1065 ( .S(n4348), .A0(n759), .A1(n758), .Z(n760));
Q_MX08 U1066 ( .S0(n4346), .S1(n4347), .S2(n4348), .A0(i_bimc_eccpar_debug[3]), .A1(i_bimc_memid[3]), .A2(i_bimc_global_config[3]), .A3(i_bimc_parity_error_cnt[3]), .A4(i_bimc_ecc_correctable_error_cnt[3]), .A5(i_bimc_ecc_uncorrectable_error_cnt[3]), .A6(o_bimc_monitor_mask[3]), .A7(i_bimc_monitor[3]), .Z(n761));
Q_MX02 U1067 ( .S(n4349), .A0(n761), .A1(n760), .Z(n762));
Q_MX04 U1068 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxcmd2[3]), .A1(o_bimc_cmd0[3]), .A2(o_bimc_cmd1[3]), .A3(i_bimc_cmd2[3]), .Z(n763));
Q_MX04 U1069 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxrsp1[3]), .A1(i_bimc_rxrsp2[3]), .A2(i_bimc_rxcmd0[3]), .A3(i_bimc_rxcmd1[3]), .Z(n764));
Q_MX04 U1070 ( .S0(n4346), .S1(n4347), .A0(i_bimc_pollrsp0[3]), .A1(i_bimc_pollrsp1[3]), .A2(i_bimc_pollrsp2[3]), .A3(i_bimc_rxrsp0[3]), .Z(n765));
Q_MX02 U1071 ( .S(n4346), .A0(i_bimc_dbgcmd1[3]), .A1(i_bimc_dbgcmd2[3]), .Z(n766));
Q_AN02 U1072 ( .A0(n4346), .A1(i_bimc_dbgcmd0[3]), .Z(n767));
Q_MX02 U1073 ( .S(n4347), .A0(n767), .A1(n766), .Z(n768));
Q_MX04 U1074 ( .S0(n4348), .S1(n4349), .A0(n768), .A1(n765), .A2(n764), .A3(n763), .Z(n769));
Q_MX02 U1075 ( .S(n4350), .A0(n769), .A1(n762), .Z(r32_mux_7_data[3]));
Q_MX03 U1076 ( .S0(n4346), .S1(n4347), .A0(o_kdf_drbg_seed_1_reseed_interval_0[4]), .A1(o_kdf_drbg_seed_1_state_value_127_96[4]), .A2(o_kdf_drbg_seed_1_state_value_95_64[4]), .Z(n770));
Q_MX04 U1077 ( .S0(n4346), .S1(n4347), .A0(i_engine_sticky_status[4]), .A1(o_interrupt_mask[4]), .A2(i_interrupt_status[4]), .A3(o_kdf_drbg_seed_1_reseed_interval_1[4]), .Z(n771));
Q_MX02 U1078 ( .S(n4348), .A0(n771), .A1(n770), .Z(n772));
Q_MX08 U1079 ( .S0(n4346), .S1(n4347), .S2(n4348), .A0(i_bimc_eccpar_debug[4]), .A1(i_bimc_memid[4]), .A2(i_bimc_global_config[4]), .A3(i_bimc_parity_error_cnt[4]), .A4(i_bimc_ecc_correctable_error_cnt[4]), .A5(i_bimc_ecc_uncorrectable_error_cnt[4]), .A6(o_bimc_monitor_mask[4]), .A7(i_bimc_monitor[4]), .Z(n773));
Q_MX02 U1080 ( .S(n4349), .A0(n773), .A1(n772), .Z(n774));
Q_MX04 U1081 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxcmd2[4]), .A1(o_bimc_cmd0[4]), .A2(o_bimc_cmd1[4]), .A3(i_bimc_cmd2[4]), .Z(n775));
Q_MX04 U1082 ( .S0(n4346), .S1(n4347), .A0(i_bimc_rxrsp1[4]), .A1(i_bimc_rxrsp2[4]), .A2(i_bimc_rxcmd0[4]), .A3(i_bimc_rxcmd1[4]), .Z(n776));
Q_MX04 U1083 ( .S0(n4346), .S1(n4347), .A0(i_bimc_pollrsp0[4]), .A1(i_bimc_pollrsp1[4]), .A2(i_bimc_pollrsp2[4]), .A3(i_bimc_rxrsp0[4]), .Z(n777));
Q_MX02 U1084 ( .S(n4346), .A0(i_bimc_dbgcmd1[4]), .A1(i_bimc_dbgcmd2[4]), .Z(n778));
Q_AN02 U1085 ( .A0(n4346), .A1(i_bimc_dbgcmd0[4]), .Z(n779));
Q_MX02 U1086 ( .S(n4347), .A0(n779), .A1(n778), .Z(n780));
Q_MX04 U1087 ( .S0(n4348), .S1(n4349), .A0(n780), .A1(n777), .A2(n776), .A3(n775), .Z(n781));
Q_MX02 U1088 ( .S(n4350), .A0(n781), .A1(n774), .Z(r32_mux_7_data[4]));
Q_MX04 U1089 ( .S0(n4351), .S1(n4352), .A0(i_engine_sticky_status[5]), .A1(o_kdf_drbg_seed_1_reseed_interval_1[5]), .A2(o_kdf_drbg_seed_1_reseed_interval_0[5]), .A3(o_kdf_drbg_seed_1_state_value_127_96[5]), .Z(n782));
Q_MX02 U1090 ( .S(n4353), .A0(n782), .A1(o_kdf_drbg_seed_1_state_value_95_64[5]), .Z(n783));
Q_MX08 U1091 ( .S0(n4351), .S1(n4352), .S2(n4353), .A0(i_bimc_eccpar_debug[5]), .A1(i_bimc_memid[5]), .A2(i_bimc_global_config[5]), .A3(i_bimc_parity_error_cnt[5]), .A4(i_bimc_ecc_correctable_error_cnt[5]), .A5(i_bimc_ecc_uncorrectable_error_cnt[5]), .A6(o_bimc_monitor_mask[5]), .A7(i_bimc_monitor[5]), .Z(n784));
Q_MX02 U1092 ( .S(n4354), .A0(n784), .A1(n783), .Z(n785));
Q_MX04 U1093 ( .S0(n4351), .S1(n4352), .A0(i_bimc_rxcmd2[5]), .A1(o_bimc_cmd0[5]), .A2(o_bimc_cmd1[5]), .A3(i_bimc_cmd2[5]), .Z(n786));
Q_MX04 U1094 ( .S0(n4351), .S1(n4352), .A0(i_bimc_rxrsp1[5]), .A1(i_bimc_rxrsp2[5]), .A2(i_bimc_rxcmd0[5]), .A3(i_bimc_rxcmd1[5]), .Z(n787));
Q_MX04 U1095 ( .S0(n4351), .S1(n4352), .A0(i_bimc_pollrsp0[5]), .A1(i_bimc_pollrsp1[5]), .A2(i_bimc_pollrsp2[5]), .A3(i_bimc_rxrsp0[5]), .Z(n788));
Q_MX02 U1096 ( .S(n4351), .A0(i_bimc_dbgcmd1[5]), .A1(i_bimc_dbgcmd2[5]), .Z(n789));
Q_AN02 U1097 ( .A0(n4351), .A1(i_bimc_dbgcmd0[5]), .Z(n790));
Q_MX02 U1098 ( .S(n4352), .A0(n790), .A1(n789), .Z(n791));
Q_MX04 U1099 ( .S0(n4353), .S1(n4354), .A0(n791), .A1(n788), .A2(n787), .A3(n786), .Z(n792));
Q_MX02 U1100 ( .S(n4355), .A0(n792), .A1(n785), .Z(r32_mux_7_data[5]));
Q_MX04 U1101 ( .S0(n4351), .S1(n4352), .A0(i_engine_sticky_status[6]), .A1(o_kdf_drbg_seed_1_reseed_interval_1[6]), .A2(o_kdf_drbg_seed_1_reseed_interval_0[6]), .A3(o_kdf_drbg_seed_1_state_value_127_96[6]), .Z(n793));
Q_MX02 U1102 ( .S(n4353), .A0(n793), .A1(o_kdf_drbg_seed_1_state_value_95_64[6]), .Z(n794));
Q_MX08 U1103 ( .S0(n4351), .S1(n4352), .S2(n4353), .A0(i_bimc_eccpar_debug[6]), .A1(i_bimc_memid[6]), .A2(i_bimc_global_config[6]), .A3(i_bimc_parity_error_cnt[6]), .A4(i_bimc_ecc_correctable_error_cnt[6]), .A5(i_bimc_ecc_uncorrectable_error_cnt[6]), .A6(o_bimc_monitor_mask[6]), .A7(i_bimc_monitor[6]), .Z(n795));
Q_MX02 U1104 ( .S(n4354), .A0(n795), .A1(n794), .Z(n796));
Q_MX04 U1105 ( .S0(n4351), .S1(n4352), .A0(i_bimc_rxcmd2[6]), .A1(o_bimc_cmd0[6]), .A2(o_bimc_cmd1[6]), .A3(i_bimc_cmd2[6]), .Z(n797));
Q_MX04 U1106 ( .S0(n4351), .S1(n4352), .A0(i_bimc_rxrsp1[6]), .A1(i_bimc_rxrsp2[6]), .A2(i_bimc_rxcmd0[6]), .A3(i_bimc_rxcmd1[6]), .Z(n798));
Q_MX04 U1107 ( .S0(n4351), .S1(n4352), .A0(i_bimc_pollrsp0[6]), .A1(i_bimc_pollrsp1[6]), .A2(i_bimc_pollrsp2[6]), .A3(i_bimc_rxrsp0[6]), .Z(n799));
Q_MX02 U1108 ( .S(n4351), .A0(i_bimc_dbgcmd1[6]), .A1(i_bimc_dbgcmd2[6]), .Z(n800));
Q_AN02 U1109 ( .A0(n4351), .A1(i_bimc_dbgcmd0[6]), .Z(n801));
Q_MX02 U1110 ( .S(n4352), .A0(n801), .A1(n800), .Z(n802));
Q_MX04 U1111 ( .S0(n4353), .S1(n4354), .A0(n802), .A1(n799), .A2(n798), .A3(n797), .Z(n803));
Q_MX02 U1112 ( .S(n4355), .A0(n803), .A1(n796), .Z(r32_mux_7_data[6]));
Q_MX03 U1113 ( .S0(n4356), .S1(n4357), .A0(o_kdf_drbg_seed_1_reseed_interval_0[7]), .A1(o_kdf_drbg_seed_1_state_value_127_96[7]), .A2(o_kdf_drbg_seed_1_state_value_95_64[7]), .Z(n804));
Q_MX08 U1114 ( .S0(n4356), .S1(n4357), .S2(n4358), .A0(i_bimc_eccpar_debug[7]), .A1(i_bimc_memid[7]), .A2(i_bimc_global_config[7]), .A3(i_bimc_parity_error_cnt[7]), .A4(i_bimc_ecc_correctable_error_cnt[7]), .A5(i_bimc_ecc_uncorrectable_error_cnt[7]), .A6(i_engine_sticky_status[7]), .A7(o_kdf_drbg_seed_1_reseed_interval_1[7]), .Z(n805));
Q_MX02 U1115 ( .S(n4359), .A0(n805), .A1(n804), .Z(n806));
Q_MX04 U1116 ( .S0(n4356), .S1(n4357), .A0(i_bimc_rxcmd2[7]), .A1(o_bimc_cmd0[7]), .A2(o_bimc_cmd1[7]), .A3(i_bimc_cmd2[7]), .Z(n807));
Q_MX04 U1117 ( .S0(n4356), .S1(n4357), .A0(i_bimc_rxrsp1[7]), .A1(i_bimc_rxrsp2[7]), .A2(i_bimc_rxcmd0[7]), .A3(i_bimc_rxcmd1[7]), .Z(n808));
Q_MX04 U1118 ( .S0(n4356), .S1(n4357), .A0(i_bimc_pollrsp0[7]), .A1(i_bimc_pollrsp1[7]), .A2(i_bimc_pollrsp2[7]), .A3(i_bimc_rxrsp0[7]), .Z(n809));
Q_MX02 U1119 ( .S(n4356), .A0(i_bimc_dbgcmd1[7]), .A1(i_bimc_dbgcmd2[7]), .Z(n810));
Q_AN02 U1120 ( .A0(n4356), .A1(i_bimc_dbgcmd0[7]), .Z(n811));
Q_MX02 U1121 ( .S(n4357), .A0(n811), .A1(n810), .Z(n812));
Q_MX04 U1122 ( .S0(n4358), .S1(n4359), .A0(n812), .A1(n809), .A2(n808), .A3(n807), .Z(n813));
Q_MX02 U1123 ( .S(n4360), .A0(n813), .A1(n806), .Z(r32_mux_7_data[7]));
Q_MX02 U1124 ( .S(n4361), .A0(o_kdf_drbg_seed_1_state_value_127_96[8]), .A1(o_kdf_drbg_seed_1_state_value_95_64[8]), .Z(n814));
Q_MX08 U1125 ( .S0(n4361), .S1(n4362), .S2(n4363), .A0(i_bimc_eccpar_debug[8]), .A1(i_bimc_memid[8]), .A2(i_bimc_global_config[8]), .A3(i_bimc_parity_error_cnt[8]), .A4(i_bimc_ecc_correctable_error_cnt[8]), .A5(i_bimc_ecc_uncorrectable_error_cnt[8]), .A6(o_kdf_drbg_seed_1_reseed_interval_1[8]), .A7(o_kdf_drbg_seed_1_reseed_interval_0[8]), .Z(n815));
Q_MX02 U1126 ( .S(n4364), .A0(n815), .A1(n814), .Z(n816));
Q_MX04 U1127 ( .S0(n4361), .S1(n4362), .A0(i_bimc_rxcmd2[8]), .A1(o_bimc_cmd0[8]), .A2(o_bimc_cmd1[8]), .A3(i_bimc_cmd2[8]), .Z(n817));
Q_MX04 U1128 ( .S0(n4361), .S1(n4362), .A0(i_bimc_rxrsp1[8]), .A1(i_bimc_rxrsp2[8]), .A2(i_bimc_rxcmd0[8]), .A3(i_bimc_rxcmd1[8]), .Z(n818));
Q_MX04 U1129 ( .S0(n4361), .S1(n4362), .A0(i_bimc_pollrsp0[8]), .A1(i_bimc_pollrsp1[8]), .A2(i_bimc_pollrsp2[8]), .A3(i_bimc_rxrsp0[8]), .Z(n819));
Q_MX02 U1130 ( .S(n4361), .A0(i_bimc_dbgcmd1[8]), .A1(i_bimc_dbgcmd2[8]), .Z(n820));
Q_AN02 U1131 ( .A0(n4361), .A1(i_bimc_dbgcmd0[8]), .Z(n821));
Q_MX02 U1132 ( .S(n4362), .A0(n821), .A1(n820), .Z(n822));
Q_MX04 U1133 ( .S0(n4363), .S1(n4364), .A0(n822), .A1(n819), .A2(n818), .A3(n817), .Z(n823));
Q_MX02 U1134 ( .S(n4365), .A0(n823), .A1(n816), .Z(r32_mux_7_data[8]));
Q_MX02 U1135 ( .S(n4361), .A0(o_kdf_drbg_seed_1_state_value_127_96[9]), .A1(o_kdf_drbg_seed_1_state_value_95_64[9]), .Z(n824));
Q_MX08 U1136 ( .S0(n4361), .S1(n4362), .S2(n4363), .A0(i_bimc_eccpar_debug[9]), .A1(i_bimc_memid[9]), .A2(i_bimc_global_config[9]), .A3(i_bimc_parity_error_cnt[9]), .A4(i_bimc_ecc_correctable_error_cnt[9]), .A5(i_bimc_ecc_uncorrectable_error_cnt[9]), .A6(o_kdf_drbg_seed_1_reseed_interval_1[9]), .A7(o_kdf_drbg_seed_1_reseed_interval_0[9]), .Z(n825));
Q_MX02 U1137 ( .S(n4364), .A0(n825), .A1(n824), .Z(n826));
Q_MX04 U1138 ( .S0(n4361), .S1(n4362), .A0(i_bimc_rxcmd2[9]), .A1(o_bimc_cmd0[9]), .A2(o_bimc_cmd1[9]), .A3(i_bimc_cmd2[9]), .Z(n827));
Q_MX04 U1139 ( .S0(n4361), .S1(n4362), .A0(i_bimc_rxrsp1[9]), .A1(i_bimc_rxrsp2[9]), .A2(i_bimc_rxcmd0[9]), .A3(i_bimc_rxcmd1[9]), .Z(n828));
Q_MX04 U1140 ( .S0(n4361), .S1(n4362), .A0(i_bimc_pollrsp0[9]), .A1(i_bimc_pollrsp1[9]), .A2(i_bimc_pollrsp2[9]), .A3(i_bimc_rxrsp0[9]), .Z(n829));
Q_MX02 U1141 ( .S(n4361), .A0(i_bimc_dbgcmd1[9]), .A1(i_bimc_dbgcmd2[9]), .Z(n830));
Q_AN02 U1142 ( .A0(n4361), .A1(i_bimc_dbgcmd0[9]), .Z(n831));
Q_MX02 U1143 ( .S(n4362), .A0(n831), .A1(n830), .Z(n832));
Q_MX04 U1144 ( .S0(n4363), .S1(n4364), .A0(n832), .A1(n829), .A2(n828), .A3(n827), .Z(n833));
Q_MX02 U1145 ( .S(n4365), .A0(n833), .A1(n826), .Z(r32_mux_7_data[9]));
Q_MX02 U1146 ( .S(n4366), .A0(o_kdf_drbg_seed_1_state_value_127_96[10]), .A1(o_kdf_drbg_seed_1_state_value_95_64[10]), .Z(n834));
Q_MX04 U1147 ( .S0(n4366), .S1(n4367), .A0(i_bimc_ecc_correctable_error_cnt[10]), .A1(i_bimc_ecc_uncorrectable_error_cnt[10]), .A2(o_kdf_drbg_seed_1_reseed_interval_1[10]), .A3(o_kdf_drbg_seed_1_reseed_interval_0[10]), .Z(n835));
Q_MX02 U1148 ( .S(n4368), .A0(n835), .A1(n834), .Z(n836));
Q_MX04 U1149 ( .S0(n4366), .S1(n4367), .A0(i_bimc_eccpar_debug[10]), .A1(i_bimc_memid[10]), .A2(i_bimc_global_config[10]), .A3(i_bimc_parity_error_cnt[10]), .Z(n837));
Q_MX04 U1150 ( .S0(n4366), .S1(n4367), .A0(i_bimc_rxcmd1[10]), .A1(o_bimc_cmd0[10]), .A2(o_bimc_cmd1[10]), .A3(i_bimc_cmd2[10]), .Z(n838));
Q_MX04 U1151 ( .S0(n4366), .S1(n4367), .A0(i_bimc_pollrsp1[10]), .A1(i_bimc_rxrsp0[10]), .A2(i_bimc_rxrsp1[10]), .A3(i_bimc_rxcmd0[10]), .Z(n839));
Q_MX02 U1152 ( .S(n4366), .A0(i_bimc_dbgcmd1[10]), .A1(i_bimc_pollrsp0[10]), .Z(n840));
Q_AN02 U1153 ( .A0(n4366), .A1(i_bimc_dbgcmd0[10]), .Z(n841));
Q_MX02 U1154 ( .S(n4367), .A0(n841), .A1(n840), .Z(n842));
Q_MX04 U1155 ( .S0(n4368), .S1(n4369), .A0(n842), .A1(n839), .A2(n838), .A3(n837), .Z(n843));
Q_MX02 U1156 ( .S(n4370), .A0(n843), .A1(n836), .Z(r32_mux_7_data[10]));
Q_MX04 U1157 ( .S0(n4371), .S1(n4372), .A0(i_bimc_ecc_uncorrectable_error_cnt[11]), .A1(o_kdf_drbg_seed_1_reseed_interval_1[11]), .A2(o_kdf_drbg_seed_1_reseed_interval_0[11]), .A3(o_kdf_drbg_seed_1_state_value_127_96[11]), .Z(n844));
Q_MX02 U1158 ( .S(n4373), .A0(n844), .A1(o_kdf_drbg_seed_1_state_value_95_64[11]), .Z(n845));
Q_MX04 U1159 ( .S0(n4371), .S1(n4372), .A0(i_bimc_memid[11]), .A1(i_bimc_global_config[11]), .A2(i_bimc_parity_error_cnt[11]), .A3(i_bimc_ecc_correctable_error_cnt[11]), .Z(n846));
Q_MX04 U1160 ( .S0(n4371), .S1(n4372), .A0(i_bimc_rxcmd1[11]), .A1(o_bimc_cmd0[11]), .A2(o_bimc_cmd1[11]), .A3(i_bimc_eccpar_debug[11]), .Z(n847));
Q_MX04 U1161 ( .S0(n4371), .S1(n4372), .A0(i_bimc_pollrsp1[11]), .A1(i_bimc_rxrsp0[11]), .A2(i_bimc_rxrsp1[11]), .A3(i_bimc_rxcmd0[11]), .Z(n848));
Q_MX02 U1162 ( .S(n4371), .A0(i_bimc_dbgcmd1[11]), .A1(i_bimc_pollrsp0[11]), .Z(n849));
Q_AN02 U1163 ( .A0(n4371), .A1(i_bimc_dbgcmd0[11]), .Z(n850));
Q_MX02 U1164 ( .S(n4372), .A0(n850), .A1(n849), .Z(n851));
Q_MX04 U1165 ( .S0(n4373), .S1(n4374), .A0(n851), .A1(n848), .A2(n847), .A3(n846), .Z(n852));
Q_MX02 U1166 ( .S(n4375), .A0(n852), .A1(n845), .Z(r32_mux_7_data[11]));
Q_MX04 U1167 ( .S0(n4376), .S1(n4377), .A0(o_kdf_drbg_seed_1_reseed_interval_1[12]), .A1(o_kdf_drbg_seed_1_reseed_interval_0[12]), .A2(o_kdf_drbg_seed_1_state_value_127_96[12]), .A3(o_kdf_drbg_seed_1_state_value_95_64[12]), .Z(n853));
Q_MX04 U1168 ( .S0(n4376), .S1(n4377), .A0(i_bimc_global_config[12]), .A1(i_bimc_parity_error_cnt[12]), .A2(i_bimc_ecc_correctable_error_cnt[12]), .A3(i_bimc_ecc_uncorrectable_error_cnt[12]), .Z(n854));
Q_MX04 U1169 ( .S0(n4376), .S1(n4377), .A0(i_bimc_rxcmd1[12]), .A1(o_bimc_cmd0[12]), .A2(o_bimc_cmd1[12]), .A3(i_bimc_eccpar_debug[12]), .Z(n855));
Q_MX04 U1170 ( .S0(n4376), .S1(n4377), .A0(i_bimc_pollrsp1[12]), .A1(i_bimc_rxrsp0[12]), .A2(i_bimc_rxrsp1[12]), .A3(i_bimc_rxcmd0[12]), .Z(n856));
Q_MX02 U1171 ( .S(n4376), .A0(i_bimc_dbgcmd1[12]), .A1(i_bimc_pollrsp0[12]), .Z(n857));
Q_AN02 U1172 ( .A0(n4376), .A1(i_bimc_dbgcmd0[12]), .Z(n858));
Q_MX02 U1173 ( .S(n4377), .A0(n858), .A1(n857), .Z(n859));
Q_MX04 U1174 ( .S0(n4378), .S1(n4379), .A0(n859), .A1(n856), .A2(n855), .A3(n854), .Z(n860));
Q_MX02 U1175 ( .S(n4380), .A0(n860), .A1(n853), .Z(r32_mux_7_data[12]));
Q_MX04 U1176 ( .S0(n4376), .S1(n4377), .A0(o_kdf_drbg_seed_1_reseed_interval_1[13]), .A1(o_kdf_drbg_seed_1_reseed_interval_0[13]), .A2(o_kdf_drbg_seed_1_state_value_127_96[13]), .A3(o_kdf_drbg_seed_1_state_value_95_64[13]), .Z(n861));
Q_MX04 U1177 ( .S0(n4376), .S1(n4377), .A0(i_bimc_global_config[13]), .A1(i_bimc_parity_error_cnt[13]), .A2(i_bimc_ecc_correctable_error_cnt[13]), .A3(i_bimc_ecc_uncorrectable_error_cnt[13]), .Z(n862));
Q_MX04 U1178 ( .S0(n4376), .S1(n4377), .A0(i_bimc_rxcmd1[13]), .A1(o_bimc_cmd0[13]), .A2(o_bimc_cmd1[13]), .A3(i_bimc_eccpar_debug[13]), .Z(n863));
Q_MX04 U1179 ( .S0(n4376), .S1(n4377), .A0(i_bimc_pollrsp1[13]), .A1(i_bimc_rxrsp0[13]), .A2(i_bimc_rxrsp1[13]), .A3(i_bimc_rxcmd0[13]), .Z(n864));
Q_MX02 U1180 ( .S(n4376), .A0(i_bimc_dbgcmd1[13]), .A1(i_bimc_pollrsp0[13]), .Z(n865));
Q_AN02 U1181 ( .A0(n4376), .A1(i_bimc_dbgcmd0[13]), .Z(n866));
Q_MX02 U1182 ( .S(n4377), .A0(n866), .A1(n865), .Z(n867));
Q_MX04 U1183 ( .S0(n4378), .S1(n4379), .A0(n867), .A1(n864), .A2(n863), .A3(n862), .Z(n868));
Q_MX02 U1184 ( .S(n4380), .A0(n868), .A1(n861), .Z(r32_mux_7_data[13]));
Q_MX04 U1185 ( .S0(n4376), .S1(n4377), .A0(o_kdf_drbg_seed_1_reseed_interval_1[14]), .A1(o_kdf_drbg_seed_1_reseed_interval_0[14]), .A2(o_kdf_drbg_seed_1_state_value_127_96[14]), .A3(o_kdf_drbg_seed_1_state_value_95_64[14]), .Z(n869));
Q_MX04 U1186 ( .S0(n4376), .S1(n4377), .A0(i_bimc_global_config[14]), .A1(i_bimc_parity_error_cnt[14]), .A2(i_bimc_ecc_correctable_error_cnt[14]), .A3(i_bimc_ecc_uncorrectable_error_cnt[14]), .Z(n870));
Q_MX04 U1187 ( .S0(n4376), .S1(n4377), .A0(i_bimc_rxcmd1[14]), .A1(o_bimc_cmd0[14]), .A2(o_bimc_cmd1[14]), .A3(i_bimc_eccpar_debug[14]), .Z(n871));
Q_MX04 U1188 ( .S0(n4376), .S1(n4377), .A0(i_bimc_pollrsp1[14]), .A1(i_bimc_rxrsp0[14]), .A2(i_bimc_rxrsp1[14]), .A3(i_bimc_rxcmd0[14]), .Z(n872));
Q_MX02 U1189 ( .S(n4376), .A0(i_bimc_dbgcmd1[14]), .A1(i_bimc_pollrsp0[14]), .Z(n873));
Q_AN02 U1190 ( .A0(n4376), .A1(i_bimc_dbgcmd0[14]), .Z(n874));
Q_MX02 U1191 ( .S(n4377), .A0(n874), .A1(n873), .Z(n875));
Q_MX04 U1192 ( .S0(n4378), .S1(n4379), .A0(n875), .A1(n872), .A2(n871), .A3(n870), .Z(n876));
Q_MX02 U1193 ( .S(n4380), .A0(n876), .A1(n869), .Z(r32_mux_7_data[14]));
Q_MX04 U1194 ( .S0(n4376), .S1(n4377), .A0(o_kdf_drbg_seed_1_reseed_interval_1[15]), .A1(o_kdf_drbg_seed_1_reseed_interval_0[15]), .A2(o_kdf_drbg_seed_1_state_value_127_96[15]), .A3(o_kdf_drbg_seed_1_state_value_95_64[15]), .Z(n877));
Q_MX04 U1195 ( .S0(n4376), .S1(n4377), .A0(i_bimc_global_config[15]), .A1(i_bimc_parity_error_cnt[15]), .A2(i_bimc_ecc_correctable_error_cnt[15]), .A3(i_bimc_ecc_uncorrectable_error_cnt[15]), .Z(n878));
Q_MX04 U1196 ( .S0(n4376), .S1(n4377), .A0(i_bimc_rxcmd1[15]), .A1(o_bimc_cmd0[15]), .A2(o_bimc_cmd1[15]), .A3(i_bimc_eccpar_debug[15]), .Z(n879));
Q_MX04 U1197 ( .S0(n4376), .S1(n4377), .A0(i_bimc_pollrsp1[15]), .A1(i_bimc_rxrsp0[15]), .A2(i_bimc_rxrsp1[15]), .A3(i_bimc_rxcmd0[15]), .Z(n880));
Q_MX02 U1198 ( .S(n4376), .A0(i_bimc_dbgcmd1[15]), .A1(i_bimc_pollrsp0[15]), .Z(n881));
Q_AN02 U1199 ( .A0(n4376), .A1(i_bimc_dbgcmd0[15]), .Z(n882));
Q_MX02 U1200 ( .S(n4377), .A0(n882), .A1(n881), .Z(n883));
Q_MX04 U1201 ( .S0(n4378), .S1(n4379), .A0(n883), .A1(n880), .A2(n879), .A3(n878), .Z(n884));
Q_MX02 U1202 ( .S(n4380), .A0(n884), .A1(n877), .Z(r32_mux_7_data[15]));
Q_MX03 U1203 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[16]), .A1(o_kdf_drbg_seed_1_state_value_127_96[16]), .A2(o_kdf_drbg_seed_1_state_value_95_64[16]), .Z(n885));
Q_MX04 U1204 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[16]), .A1(i_bimc_parity_error_cnt[16]), .A2(i_bimc_ecc_correctable_error_cnt[16]), .A3(i_bimc_ecc_uncorrectable_error_cnt[16]), .Z(n886));
Q_MX04 U1205 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[16]), .A1(o_bimc_cmd0[16]), .A2(o_bimc_cmd1[16]), .A3(i_bimc_eccpar_debug[16]), .Z(n887));
Q_MX04 U1206 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[16]), .A1(i_bimc_rxrsp0[16]), .A2(i_bimc_rxrsp1[16]), .A3(i_bimc_rxcmd0[16]), .Z(n888));
Q_MX02 U1207 ( .S(n4381), .A0(i_bimc_dbgcmd1[16]), .A1(i_bimc_pollrsp0[16]), .Z(n889));
Q_AN02 U1208 ( .A0(n4381), .A1(i_bimc_dbgcmd0[16]), .Z(n890));
Q_MX02 U1209 ( .S(n4382), .A0(n890), .A1(n889), .Z(n891));
Q_MX04 U1210 ( .S0(n4378), .S1(n4379), .A0(n891), .A1(n888), .A2(n887), .A3(n886), .Z(n892));
Q_MX02 U1211 ( .S(n4383), .A0(n892), .A1(n885), .Z(r32_mux_7_data[16]));
Q_MX03 U1212 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[17]), .A1(o_kdf_drbg_seed_1_state_value_127_96[17]), .A2(o_kdf_drbg_seed_1_state_value_95_64[17]), .Z(n893));
Q_MX04 U1213 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[17]), .A1(i_bimc_parity_error_cnt[17]), .A2(i_bimc_ecc_correctable_error_cnt[17]), .A3(i_bimc_ecc_uncorrectable_error_cnt[17]), .Z(n894));
Q_MX04 U1214 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[17]), .A1(o_bimc_cmd0[17]), .A2(o_bimc_cmd1[17]), .A3(i_bimc_eccpar_debug[17]), .Z(n895));
Q_MX04 U1215 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[17]), .A1(i_bimc_rxrsp0[17]), .A2(i_bimc_rxrsp1[17]), .A3(i_bimc_rxcmd0[17]), .Z(n896));
Q_MX02 U1216 ( .S(n4381), .A0(i_bimc_dbgcmd1[17]), .A1(i_bimc_pollrsp0[17]), .Z(n897));
Q_AN02 U1217 ( .A0(n4381), .A1(i_bimc_dbgcmd0[17]), .Z(n898));
Q_MX02 U1218 ( .S(n4382), .A0(n898), .A1(n897), .Z(n899));
Q_MX04 U1219 ( .S0(n4378), .S1(n4379), .A0(n899), .A1(n896), .A2(n895), .A3(n894), .Z(n900));
Q_MX02 U1220 ( .S(n4383), .A0(n900), .A1(n893), .Z(r32_mux_7_data[17]));
Q_MX03 U1221 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[18]), .A1(o_kdf_drbg_seed_1_state_value_127_96[18]), .A2(o_kdf_drbg_seed_1_state_value_95_64[18]), .Z(n901));
Q_MX04 U1222 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[18]), .A1(i_bimc_parity_error_cnt[18]), .A2(i_bimc_ecc_correctable_error_cnt[18]), .A3(i_bimc_ecc_uncorrectable_error_cnt[18]), .Z(n902));
Q_MX04 U1223 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[18]), .A1(o_bimc_cmd0[18]), .A2(o_bimc_cmd1[18]), .A3(i_bimc_eccpar_debug[18]), .Z(n903));
Q_MX04 U1224 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[18]), .A1(i_bimc_rxrsp0[18]), .A2(i_bimc_rxrsp1[18]), .A3(i_bimc_rxcmd0[18]), .Z(n904));
Q_MX02 U1225 ( .S(n4381), .A0(i_bimc_dbgcmd1[18]), .A1(i_bimc_pollrsp0[18]), .Z(n905));
Q_AN02 U1226 ( .A0(n4381), .A1(i_bimc_dbgcmd0[18]), .Z(n906));
Q_MX02 U1227 ( .S(n4382), .A0(n906), .A1(n905), .Z(n907));
Q_MX04 U1228 ( .S0(n4378), .S1(n4379), .A0(n907), .A1(n904), .A2(n903), .A3(n902), .Z(n908));
Q_MX02 U1229 ( .S(n4383), .A0(n908), .A1(n901), .Z(r32_mux_7_data[18]));
Q_MX03 U1230 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[19]), .A1(o_kdf_drbg_seed_1_state_value_127_96[19]), .A2(o_kdf_drbg_seed_1_state_value_95_64[19]), .Z(n909));
Q_MX04 U1231 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[19]), .A1(i_bimc_parity_error_cnt[19]), .A2(i_bimc_ecc_correctable_error_cnt[19]), .A3(i_bimc_ecc_uncorrectable_error_cnt[19]), .Z(n910));
Q_MX04 U1232 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[19]), .A1(o_bimc_cmd0[19]), .A2(o_bimc_cmd1[19]), .A3(i_bimc_eccpar_debug[19]), .Z(n911));
Q_MX04 U1233 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[19]), .A1(i_bimc_rxrsp0[19]), .A2(i_bimc_rxrsp1[19]), .A3(i_bimc_rxcmd0[19]), .Z(n912));
Q_MX02 U1234 ( .S(n4381), .A0(i_bimc_dbgcmd1[19]), .A1(i_bimc_pollrsp0[19]), .Z(n913));
Q_AN02 U1235 ( .A0(n4381), .A1(i_bimc_dbgcmd0[19]), .Z(n914));
Q_MX02 U1236 ( .S(n4382), .A0(n914), .A1(n913), .Z(n915));
Q_MX04 U1237 ( .S0(n4378), .S1(n4379), .A0(n915), .A1(n912), .A2(n911), .A3(n910), .Z(n916));
Q_MX02 U1238 ( .S(n4383), .A0(n916), .A1(n909), .Z(r32_mux_7_data[19]));
Q_MX03 U1239 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[20]), .A1(o_kdf_drbg_seed_1_state_value_127_96[20]), .A2(o_kdf_drbg_seed_1_state_value_95_64[20]), .Z(n917));
Q_MX04 U1240 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[20]), .A1(i_bimc_parity_error_cnt[20]), .A2(i_bimc_ecc_correctable_error_cnt[20]), .A3(i_bimc_ecc_uncorrectable_error_cnt[20]), .Z(n918));
Q_MX04 U1241 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[20]), .A1(o_bimc_cmd0[20]), .A2(o_bimc_cmd1[20]), .A3(i_bimc_eccpar_debug[20]), .Z(n919));
Q_MX04 U1242 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[20]), .A1(i_bimc_rxrsp0[20]), .A2(i_bimc_rxrsp1[20]), .A3(i_bimc_rxcmd0[20]), .Z(n920));
Q_MX02 U1243 ( .S(n4381), .A0(i_bimc_dbgcmd1[20]), .A1(i_bimc_pollrsp0[20]), .Z(n921));
Q_AN02 U1244 ( .A0(n4381), .A1(i_bimc_dbgcmd0[20]), .Z(n922));
Q_MX02 U1245 ( .S(n4382), .A0(n922), .A1(n921), .Z(n923));
Q_MX04 U1246 ( .S0(n4378), .S1(n4379), .A0(n923), .A1(n920), .A2(n919), .A3(n918), .Z(n924));
Q_MX02 U1247 ( .S(n4383), .A0(n924), .A1(n917), .Z(r32_mux_7_data[20]));
Q_MX03 U1248 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[21]), .A1(o_kdf_drbg_seed_1_state_value_127_96[21]), .A2(o_kdf_drbg_seed_1_state_value_95_64[21]), .Z(n925));
Q_MX04 U1249 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[21]), .A1(i_bimc_parity_error_cnt[21]), .A2(i_bimc_ecc_correctable_error_cnt[21]), .A3(i_bimc_ecc_uncorrectable_error_cnt[21]), .Z(n926));
Q_MX04 U1250 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[21]), .A1(o_bimc_cmd0[21]), .A2(o_bimc_cmd1[21]), .A3(i_bimc_eccpar_debug[21]), .Z(n927));
Q_MX04 U1251 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[21]), .A1(i_bimc_rxrsp0[21]), .A2(i_bimc_rxrsp1[21]), .A3(i_bimc_rxcmd0[21]), .Z(n928));
Q_MX02 U1252 ( .S(n4381), .A0(i_bimc_dbgcmd1[21]), .A1(i_bimc_pollrsp0[21]), .Z(n929));
Q_AN02 U1253 ( .A0(n4381), .A1(i_bimc_dbgcmd0[21]), .Z(n930));
Q_MX02 U1254 ( .S(n4382), .A0(n930), .A1(n929), .Z(n931));
Q_MX04 U1255 ( .S0(n4378), .S1(n4379), .A0(n931), .A1(n928), .A2(n927), .A3(n926), .Z(n932));
Q_MX02 U1256 ( .S(n4383), .A0(n932), .A1(n925), .Z(r32_mux_7_data[21]));
Q_MX03 U1257 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[22]), .A1(o_kdf_drbg_seed_1_state_value_127_96[22]), .A2(o_kdf_drbg_seed_1_state_value_95_64[22]), .Z(n933));
Q_MX04 U1258 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[22]), .A1(i_bimc_parity_error_cnt[22]), .A2(i_bimc_ecc_correctable_error_cnt[22]), .A3(i_bimc_ecc_uncorrectable_error_cnt[22]), .Z(n934));
Q_MX04 U1259 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[22]), .A1(o_bimc_cmd0[22]), .A2(o_bimc_cmd1[22]), .A3(i_bimc_eccpar_debug[22]), .Z(n935));
Q_MX04 U1260 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[22]), .A1(i_bimc_rxrsp0[22]), .A2(i_bimc_rxrsp1[22]), .A3(i_bimc_rxcmd0[22]), .Z(n936));
Q_MX02 U1261 ( .S(n4381), .A0(i_bimc_dbgcmd1[22]), .A1(i_bimc_pollrsp0[22]), .Z(n937));
Q_AN02 U1262 ( .A0(n4381), .A1(i_bimc_dbgcmd0[22]), .Z(n938));
Q_MX02 U1263 ( .S(n4382), .A0(n938), .A1(n937), .Z(n939));
Q_MX04 U1264 ( .S0(n4378), .S1(n4379), .A0(n939), .A1(n936), .A2(n935), .A3(n934), .Z(n940));
Q_MX02 U1265 ( .S(n4383), .A0(n940), .A1(n933), .Z(r32_mux_7_data[22]));
Q_MX03 U1266 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[23]), .A1(o_kdf_drbg_seed_1_state_value_127_96[23]), .A2(o_kdf_drbg_seed_1_state_value_95_64[23]), .Z(n941));
Q_MX04 U1267 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[23]), .A1(i_bimc_parity_error_cnt[23]), .A2(i_bimc_ecc_correctable_error_cnt[23]), .A3(i_bimc_ecc_uncorrectable_error_cnt[23]), .Z(n942));
Q_MX04 U1268 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[23]), .A1(o_bimc_cmd0[23]), .A2(o_bimc_cmd1[23]), .A3(i_bimc_eccpar_debug[23]), .Z(n943));
Q_MX04 U1269 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[23]), .A1(i_bimc_rxrsp0[23]), .A2(i_bimc_rxrsp1[23]), .A3(i_bimc_rxcmd0[23]), .Z(n944));
Q_MX02 U1270 ( .S(n4381), .A0(i_bimc_dbgcmd1[23]), .A1(i_bimc_pollrsp0[23]), .Z(n945));
Q_AN02 U1271 ( .A0(n4381), .A1(i_bimc_dbgcmd0[23]), .Z(n946));
Q_MX02 U1272 ( .S(n4382), .A0(n946), .A1(n945), .Z(n947));
Q_MX04 U1273 ( .S0(n4378), .S1(n4379), .A0(n947), .A1(n944), .A2(n943), .A3(n942), .Z(n948));
Q_MX02 U1274 ( .S(n4383), .A0(n948), .A1(n941), .Z(r32_mux_7_data[23]));
Q_MX03 U1275 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[24]), .A1(o_kdf_drbg_seed_1_state_value_127_96[24]), .A2(o_kdf_drbg_seed_1_state_value_95_64[24]), .Z(n949));
Q_MX04 U1276 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[24]), .A1(i_bimc_parity_error_cnt[24]), .A2(i_bimc_ecc_correctable_error_cnt[24]), .A3(i_bimc_ecc_uncorrectable_error_cnt[24]), .Z(n950));
Q_MX04 U1277 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[24]), .A1(o_bimc_cmd0[24]), .A2(o_bimc_cmd1[24]), .A3(i_bimc_eccpar_debug[24]), .Z(n951));
Q_MX04 U1278 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[24]), .A1(i_bimc_rxrsp0[24]), .A2(i_bimc_rxrsp1[24]), .A3(i_bimc_rxcmd0[24]), .Z(n952));
Q_MX02 U1279 ( .S(n4381), .A0(i_bimc_dbgcmd1[24]), .A1(i_bimc_pollrsp0[24]), .Z(n953));
Q_AN02 U1280 ( .A0(n4381), .A1(i_bimc_dbgcmd0[24]), .Z(n954));
Q_MX02 U1281 ( .S(n4382), .A0(n954), .A1(n953), .Z(n955));
Q_MX04 U1282 ( .S0(n4378), .S1(n4379), .A0(n955), .A1(n952), .A2(n951), .A3(n950), .Z(n956));
Q_MX02 U1283 ( .S(n4383), .A0(n956), .A1(n949), .Z(r32_mux_7_data[24]));
Q_MX03 U1284 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[25]), .A1(o_kdf_drbg_seed_1_state_value_127_96[25]), .A2(o_kdf_drbg_seed_1_state_value_95_64[25]), .Z(n957));
Q_MX04 U1285 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[25]), .A1(i_bimc_parity_error_cnt[25]), .A2(i_bimc_ecc_correctable_error_cnt[25]), .A3(i_bimc_ecc_uncorrectable_error_cnt[25]), .Z(n958));
Q_MX04 U1286 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[25]), .A1(o_bimc_cmd0[25]), .A2(o_bimc_cmd1[25]), .A3(i_bimc_eccpar_debug[25]), .Z(n959));
Q_MX04 U1287 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[25]), .A1(i_bimc_rxrsp0[25]), .A2(i_bimc_rxrsp1[25]), .A3(i_bimc_rxcmd0[25]), .Z(n960));
Q_MX02 U1288 ( .S(n4381), .A0(i_bimc_dbgcmd1[25]), .A1(i_bimc_pollrsp0[25]), .Z(n961));
Q_AN02 U1289 ( .A0(n4381), .A1(i_bimc_dbgcmd0[25]), .Z(n962));
Q_MX02 U1290 ( .S(n4382), .A0(n962), .A1(n961), .Z(n963));
Q_MX04 U1291 ( .S0(n4378), .S1(n4379), .A0(n963), .A1(n960), .A2(n959), .A3(n958), .Z(n964));
Q_MX02 U1292 ( .S(n4383), .A0(n964), .A1(n957), .Z(r32_mux_7_data[25]));
Q_MX03 U1293 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[26]), .A1(o_kdf_drbg_seed_1_state_value_127_96[26]), .A2(o_kdf_drbg_seed_1_state_value_95_64[26]), .Z(n965));
Q_MX04 U1294 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[26]), .A1(i_bimc_parity_error_cnt[26]), .A2(i_bimc_ecc_correctable_error_cnt[26]), .A3(i_bimc_ecc_uncorrectable_error_cnt[26]), .Z(n966));
Q_MX04 U1295 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[26]), .A1(o_bimc_cmd0[26]), .A2(o_bimc_cmd1[26]), .A3(i_bimc_eccpar_debug[26]), .Z(n967));
Q_MX04 U1296 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[26]), .A1(i_bimc_rxrsp0[26]), .A2(i_bimc_rxrsp1[26]), .A3(i_bimc_rxcmd0[26]), .Z(n968));
Q_MX02 U1297 ( .S(n4381), .A0(i_bimc_dbgcmd1[26]), .A1(i_bimc_pollrsp0[26]), .Z(n969));
Q_AN02 U1298 ( .A0(n4381), .A1(i_bimc_dbgcmd0[26]), .Z(n970));
Q_MX02 U1299 ( .S(n4382), .A0(n970), .A1(n969), .Z(n971));
Q_MX04 U1300 ( .S0(n4378), .S1(n4379), .A0(n971), .A1(n968), .A2(n967), .A3(n966), .Z(n972));
Q_MX02 U1301 ( .S(n4383), .A0(n972), .A1(n965), .Z(r32_mux_7_data[26]));
Q_MX03 U1302 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[27]), .A1(o_kdf_drbg_seed_1_state_value_127_96[27]), .A2(o_kdf_drbg_seed_1_state_value_95_64[27]), .Z(n973));
Q_MX04 U1303 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[27]), .A1(i_bimc_parity_error_cnt[27]), .A2(i_bimc_ecc_correctable_error_cnt[27]), .A3(i_bimc_ecc_uncorrectable_error_cnt[27]), .Z(n974));
Q_MX04 U1304 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[27]), .A1(o_bimc_cmd0[27]), .A2(o_bimc_cmd1[27]), .A3(i_bimc_eccpar_debug[27]), .Z(n975));
Q_MX04 U1305 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[27]), .A1(i_bimc_rxrsp0[27]), .A2(i_bimc_rxrsp1[27]), .A3(i_bimc_rxcmd0[27]), .Z(n976));
Q_MX02 U1306 ( .S(n4381), .A0(i_bimc_dbgcmd1[27]), .A1(i_bimc_pollrsp0[27]), .Z(n977));
Q_AN02 U1307 ( .A0(n4381), .A1(i_bimc_dbgcmd0[27]), .Z(n978));
Q_MX02 U1308 ( .S(n4382), .A0(n978), .A1(n977), .Z(n979));
Q_MX04 U1309 ( .S0(n4378), .S1(n4379), .A0(n979), .A1(n976), .A2(n975), .A3(n974), .Z(n980));
Q_MX02 U1310 ( .S(n4383), .A0(n980), .A1(n973), .Z(r32_mux_7_data[27]));
Q_MX03 U1311 ( .S0(n4381), .S1(n4382), .A0(o_kdf_drbg_seed_1_reseed_interval_0[28]), .A1(o_kdf_drbg_seed_1_state_value_127_96[28]), .A2(o_kdf_drbg_seed_1_state_value_95_64[28]), .Z(n981));
Q_MX04 U1312 ( .S0(n4381), .S1(n4382), .A0(i_bimc_global_config[28]), .A1(i_bimc_parity_error_cnt[28]), .A2(i_bimc_ecc_correctable_error_cnt[28]), .A3(i_bimc_ecc_uncorrectable_error_cnt[28]), .Z(n982));
Q_MX04 U1313 ( .S0(n4381), .S1(n4382), .A0(i_bimc_rxcmd1[28]), .A1(o_bimc_cmd0[28]), .A2(o_bimc_cmd1[28]), .A3(i_bimc_eccpar_debug[28]), .Z(n983));
Q_MX04 U1314 ( .S0(n4381), .S1(n4382), .A0(i_bimc_pollrsp1[28]), .A1(i_bimc_rxrsp0[28]), .A2(i_bimc_rxrsp1[28]), .A3(i_bimc_rxcmd0[28]), .Z(n984));
Q_MX02 U1315 ( .S(n4381), .A0(i_bimc_dbgcmd1[28]), .A1(i_bimc_pollrsp0[28]), .Z(n985));
Q_AN02 U1316 ( .A0(n4381), .A1(i_bimc_dbgcmd0[28]), .Z(n986));
Q_MX02 U1317 ( .S(n4382), .A0(n986), .A1(n985), .Z(n987));
Q_MX04 U1318 ( .S0(n4378), .S1(n4379), .A0(n987), .A1(n984), .A2(n983), .A3(n982), .Z(n988));
Q_MX02 U1319 ( .S(n4383), .A0(n988), .A1(n981), .Z(r32_mux_7_data[28]));
Q_MX02 U1320 ( .S(n4384), .A0(o_kdf_drbg_seed_1_state_value_127_96[29]), .A1(o_kdf_drbg_seed_1_state_value_95_64[29]), .Z(n989));
Q_MX04 U1321 ( .S0(n4384), .S1(n4385), .A0(i_bimc_parity_error_cnt[29]), .A1(i_bimc_ecc_correctable_error_cnt[29]), .A2(i_bimc_ecc_uncorrectable_error_cnt[29]), .A3(o_kdf_drbg_seed_1_reseed_interval_0[29]), .Z(n990));
Q_MX04 U1322 ( .S0(n4384), .S1(n4385), .A0(i_bimc_rxcmd1[29]), .A1(o_bimc_cmd0[29]), .A2(o_bimc_cmd1[29]), .A3(i_bimc_global_config[29]), .Z(n991));
Q_MX04 U1323 ( .S0(n4384), .S1(n4385), .A0(i_bimc_pollrsp1[29]), .A1(i_bimc_rxrsp0[29]), .A2(i_bimc_rxrsp1[29]), .A3(i_bimc_rxcmd0[29]), .Z(n992));
Q_MX02 U1324 ( .S(n4384), .A0(i_bimc_dbgcmd1[29]), .A1(i_bimc_pollrsp0[29]), .Z(n993));
Q_AN02 U1325 ( .A0(n4384), .A1(i_bimc_dbgcmd0[29]), .Z(n994));
Q_MX02 U1326 ( .S(n4385), .A0(n994), .A1(n993), .Z(n995));
Q_MX04 U1327 ( .S0(n4386), .S1(n4387), .A0(n995), .A1(n992), .A2(n991), .A3(n990), .Z(n996));
Q_MX02 U1328 ( .S(n4388), .A0(n996), .A1(n989), .Z(r32_mux_7_data[29]));
Q_MX02 U1329 ( .S(n4384), .A0(o_kdf_drbg_seed_1_state_value_127_96[30]), .A1(o_kdf_drbg_seed_1_state_value_95_64[30]), .Z(n997));
Q_MX04 U1330 ( .S0(n4384), .S1(n4385), .A0(i_bimc_parity_error_cnt[30]), .A1(i_bimc_ecc_correctable_error_cnt[30]), .A2(i_bimc_ecc_uncorrectable_error_cnt[30]), .A3(o_kdf_drbg_seed_1_reseed_interval_0[30]), .Z(n998));
Q_MX04 U1331 ( .S0(n4384), .S1(n4385), .A0(i_bimc_rxcmd1[30]), .A1(o_bimc_cmd0[30]), .A2(o_bimc_cmd1[30]), .A3(i_bimc_global_config[30]), .Z(n999));
Q_MX04 U1332 ( .S0(n4384), .S1(n4385), .A0(i_bimc_pollrsp1[30]), .A1(i_bimc_rxrsp0[30]), .A2(i_bimc_rxrsp1[30]), .A3(i_bimc_rxcmd0[30]), .Z(n1000));
Q_MX02 U1333 ( .S(n4384), .A0(i_bimc_dbgcmd1[30]), .A1(i_bimc_pollrsp0[30]), .Z(n1001));
Q_AN02 U1334 ( .A0(n4384), .A1(i_bimc_dbgcmd0[30]), .Z(n1002));
Q_MX02 U1335 ( .S(n4385), .A0(n1002), .A1(n1001), .Z(n1003));
Q_MX04 U1336 ( .S0(n4386), .S1(n4387), .A0(n1003), .A1(n1000), .A2(n999), .A3(n998), .Z(n1004));
Q_MX02 U1337 ( .S(n4388), .A0(n1004), .A1(n997), .Z(r32_mux_7_data[30]));
Q_MX02 U1338 ( .S(n4384), .A0(o_kdf_drbg_seed_1_state_value_127_96[31]), .A1(o_kdf_drbg_seed_1_state_value_95_64[31]), .Z(n1005));
Q_MX04 U1339 ( .S0(n4384), .S1(n4385), .A0(i_bimc_parity_error_cnt[31]), .A1(i_bimc_ecc_correctable_error_cnt[31]), .A2(i_bimc_ecc_uncorrectable_error_cnt[31]), .A3(o_kdf_drbg_seed_1_reseed_interval_0[31]), .Z(n1006));
Q_MX04 U1340 ( .S0(n4384), .S1(n4385), .A0(i_bimc_rxcmd1[31]), .A1(o_bimc_cmd0[31]), .A2(o_bimc_cmd1[31]), .A3(i_bimc_global_config[31]), .Z(n1007));
Q_MX04 U1341 ( .S0(n4384), .S1(n4385), .A0(i_bimc_pollrsp1[31]), .A1(i_bimc_rxrsp0[31]), .A2(i_bimc_rxrsp1[31]), .A3(i_bimc_rxcmd0[31]), .Z(n1008));
Q_MX02 U1342 ( .S(n4384), .A0(i_bimc_dbgcmd1[31]), .A1(i_bimc_pollrsp0[31]), .Z(n1009));
Q_AN02 U1343 ( .A0(n4384), .A1(i_bimc_dbgcmd0[31]), .Z(n1010));
Q_MX02 U1344 ( .S(n4385), .A0(n1010), .A1(n1009), .Z(n1011));
Q_MX04 U1345 ( .S0(n4386), .S1(n4387), .A0(n1011), .A1(n1008), .A2(n1007), .A3(n1006), .Z(n1012));
Q_MX02 U1346 ( .S(n4388), .A0(n1012), .A1(n1005), .Z(r32_mux_7_data[31]));
Q_MX03 U1347 ( .S0(n4389), .S1(n4390), .A0(o_label7_data2[0]), .A1(o_label7_data3[0]), .A2(o_label7_data4[0]), .Z(n1013));
Q_MX04 U1348 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_0_state_key_31_0[0]), .A1(i_kdf_drbg_ctrl[0]), .A2(o_label7_data0[0]), .A3(o_label7_data1[0]), .Z(n1014));
Q_MX02 U1349 ( .S(n4391), .A0(n1014), .A1(n1013), .Z(n1015));
Q_MX08 U1350 ( .S0(n4389), .S1(n4390), .S2(n4391), .A0(o_kdf_drbg_seed_0_state_value_31_0[0]), .A1(o_kdf_drbg_seed_0_state_key_255_224[0]), .A2(o_kdf_drbg_seed_0_state_key_223_192[0]), .A3(o_kdf_drbg_seed_0_state_key_191_160[0]), .A4(o_kdf_drbg_seed_0_state_key_159_128[0]), .A5(o_kdf_drbg_seed_0_state_key_127_96[0]), .A6(o_kdf_drbg_seed_0_state_key_95_64[0]), .A7(o_kdf_drbg_seed_0_state_key_63_32[0]), .Z(n1016));
Q_MX02 U1351 ( .S(n4392), .A0(n1016), .A1(n1015), .Z(n1017));
Q_MX04 U1352 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_0_reseed_interval_0[0]), .A1(o_kdf_drbg_seed_0_state_value_127_96[0]), .A2(o_kdf_drbg_seed_0_state_value_95_64[0]), .A3(o_kdf_drbg_seed_0_state_value_63_32[0]), .Z(n1018));
Q_MX04 U1353 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_1_state_key_95_64[0]), .A1(o_kdf_drbg_seed_1_state_key_63_32[0]), .A2(o_kdf_drbg_seed_1_state_key_31_0[0]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[0]), .Z(n1019));
Q_MX04 U1354 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_1_state_key_223_192[0]), .A1(o_kdf_drbg_seed_1_state_key_191_160[0]), .A2(o_kdf_drbg_seed_1_state_key_159_128[0]), .A3(o_kdf_drbg_seed_1_state_key_127_96[0]), .Z(n1020));
Q_MX02 U1355 ( .S(n4389), .A0(o_kdf_drbg_seed_1_state_value_31_0[0]), .A1(o_kdf_drbg_seed_1_state_key_255_224[0]), .Z(n1021));
Q_AN02 U1356 ( .A0(n4389), .A1(o_kdf_drbg_seed_1_state_value_63_32[0]), .Z(n1022));
Q_MX02 U1357 ( .S(n4390), .A0(n1022), .A1(n1021), .Z(n1023));
Q_MX04 U1358 ( .S0(n4391), .S1(n4392), .A0(n1023), .A1(n1020), .A2(n1019), .A3(n1018), .Z(n1024));
Q_MX02 U1359 ( .S(n4393), .A0(n1024), .A1(n1017), .Z(r32_mux_6_data[0]));
Q_MX03 U1360 ( .S0(n4389), .S1(n4390), .A0(o_label7_data2[1]), .A1(o_label7_data3[1]), .A2(o_label7_data4[1]), .Z(n1025));
Q_MX04 U1361 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_0_state_key_31_0[1]), .A1(i_kdf_drbg_ctrl[1]), .A2(o_label7_data0[1]), .A3(o_label7_data1[1]), .Z(n1026));
Q_MX02 U1362 ( .S(n4391), .A0(n1026), .A1(n1025), .Z(n1027));
Q_MX08 U1363 ( .S0(n4389), .S1(n4390), .S2(n4391), .A0(o_kdf_drbg_seed_0_state_value_31_0[1]), .A1(o_kdf_drbg_seed_0_state_key_255_224[1]), .A2(o_kdf_drbg_seed_0_state_key_223_192[1]), .A3(o_kdf_drbg_seed_0_state_key_191_160[1]), .A4(o_kdf_drbg_seed_0_state_key_159_128[1]), .A5(o_kdf_drbg_seed_0_state_key_127_96[1]), .A6(o_kdf_drbg_seed_0_state_key_95_64[1]), .A7(o_kdf_drbg_seed_0_state_key_63_32[1]), .Z(n1028));
Q_MX02 U1364 ( .S(n4392), .A0(n1028), .A1(n1027), .Z(n1029));
Q_MX04 U1365 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_0_reseed_interval_0[1]), .A1(o_kdf_drbg_seed_0_state_value_127_96[1]), .A2(o_kdf_drbg_seed_0_state_value_95_64[1]), .A3(o_kdf_drbg_seed_0_state_value_63_32[1]), .Z(n1030));
Q_MX04 U1366 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_1_state_key_95_64[1]), .A1(o_kdf_drbg_seed_1_state_key_63_32[1]), .A2(o_kdf_drbg_seed_1_state_key_31_0[1]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[1]), .Z(n1031));
Q_MX04 U1367 ( .S0(n4389), .S1(n4390), .A0(o_kdf_drbg_seed_1_state_key_223_192[1]), .A1(o_kdf_drbg_seed_1_state_key_191_160[1]), .A2(o_kdf_drbg_seed_1_state_key_159_128[1]), .A3(o_kdf_drbg_seed_1_state_key_127_96[1]), .Z(n1032));
Q_MX02 U1368 ( .S(n4389), .A0(o_kdf_drbg_seed_1_state_value_31_0[1]), .A1(o_kdf_drbg_seed_1_state_key_255_224[1]), .Z(n1033));
Q_AN02 U1369 ( .A0(n4389), .A1(o_kdf_drbg_seed_1_state_value_63_32[1]), .Z(n1034));
Q_MX02 U1370 ( .S(n4390), .A0(n1034), .A1(n1033), .Z(n1035));
Q_MX04 U1371 ( .S0(n4391), .S1(n4392), .A0(n1035), .A1(n1032), .A2(n1031), .A3(n1030), .Z(n1036));
Q_MX02 U1372 ( .S(n4393), .A0(n1036), .A1(n1029), .Z(r32_mux_6_data[1]));
Q_MX02 U1373 ( .S(n4394), .A0(o_label7_data3[2]), .A1(o_label7_data4[2]), .Z(n1037));
Q_MX04 U1374 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[2]), .A1(o_label7_data0[2]), .A2(o_label7_data1[2]), .A3(o_label7_data2[2]), .Z(n1038));
Q_MX02 U1375 ( .S(n4396), .A0(n1038), .A1(n1037), .Z(n1039));
Q_MX08 U1376 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[2]), .A1(o_kdf_drbg_seed_0_state_key_255_224[2]), .A2(o_kdf_drbg_seed_0_state_key_223_192[2]), .A3(o_kdf_drbg_seed_0_state_key_191_160[2]), .A4(o_kdf_drbg_seed_0_state_key_159_128[2]), .A5(o_kdf_drbg_seed_0_state_key_127_96[2]), .A6(o_kdf_drbg_seed_0_state_key_95_64[2]), .A7(o_kdf_drbg_seed_0_state_key_63_32[2]), .Z(n1040));
Q_MX02 U1377 ( .S(n4397), .A0(n1040), .A1(n1039), .Z(n1041));
Q_MX04 U1378 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[2]), .A1(o_kdf_drbg_seed_0_state_value_127_96[2]), .A2(o_kdf_drbg_seed_0_state_value_95_64[2]), .A3(o_kdf_drbg_seed_0_state_value_63_32[2]), .Z(n1042));
Q_MX04 U1379 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[2]), .A1(o_kdf_drbg_seed_1_state_key_63_32[2]), .A2(o_kdf_drbg_seed_1_state_key_31_0[2]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[2]), .Z(n1043));
Q_MX04 U1380 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[2]), .A1(o_kdf_drbg_seed_1_state_key_191_160[2]), .A2(o_kdf_drbg_seed_1_state_key_159_128[2]), .A3(o_kdf_drbg_seed_1_state_key_127_96[2]), .Z(n1044));
Q_MX02 U1381 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[2]), .A1(o_kdf_drbg_seed_1_state_key_255_224[2]), .Z(n1045));
Q_AN02 U1382 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[2]), .Z(n1046));
Q_MX02 U1383 ( .S(n4395), .A0(n1046), .A1(n1045), .Z(n1047));
Q_MX04 U1384 ( .S0(n4396), .S1(n4397), .A0(n1047), .A1(n1044), .A2(n1043), .A3(n1042), .Z(n1048));
Q_MX02 U1385 ( .S(n4398), .A0(n1048), .A1(n1041), .Z(r32_mux_6_data[2]));
Q_MX02 U1386 ( .S(n4394), .A0(o_label7_data3[3]), .A1(o_label7_data4[3]), .Z(n1049));
Q_MX04 U1387 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[3]), .A1(o_label7_data0[3]), .A2(o_label7_data1[3]), .A3(o_label7_data2[3]), .Z(n1050));
Q_MX02 U1388 ( .S(n4396), .A0(n1050), .A1(n1049), .Z(n1051));
Q_MX08 U1389 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[3]), .A1(o_kdf_drbg_seed_0_state_key_255_224[3]), .A2(o_kdf_drbg_seed_0_state_key_223_192[3]), .A3(o_kdf_drbg_seed_0_state_key_191_160[3]), .A4(o_kdf_drbg_seed_0_state_key_159_128[3]), .A5(o_kdf_drbg_seed_0_state_key_127_96[3]), .A6(o_kdf_drbg_seed_0_state_key_95_64[3]), .A7(o_kdf_drbg_seed_0_state_key_63_32[3]), .Z(n1052));
Q_MX02 U1390 ( .S(n4397), .A0(n1052), .A1(n1051), .Z(n1053));
Q_MX04 U1391 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[3]), .A1(o_kdf_drbg_seed_0_state_value_127_96[3]), .A2(o_kdf_drbg_seed_0_state_value_95_64[3]), .A3(o_kdf_drbg_seed_0_state_value_63_32[3]), .Z(n1054));
Q_MX04 U1392 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[3]), .A1(o_kdf_drbg_seed_1_state_key_63_32[3]), .A2(o_kdf_drbg_seed_1_state_key_31_0[3]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[3]), .Z(n1055));
Q_MX04 U1393 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[3]), .A1(o_kdf_drbg_seed_1_state_key_191_160[3]), .A2(o_kdf_drbg_seed_1_state_key_159_128[3]), .A3(o_kdf_drbg_seed_1_state_key_127_96[3]), .Z(n1056));
Q_MX02 U1394 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[3]), .A1(o_kdf_drbg_seed_1_state_key_255_224[3]), .Z(n1057));
Q_AN02 U1395 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[3]), .Z(n1058));
Q_MX02 U1396 ( .S(n4395), .A0(n1058), .A1(n1057), .Z(n1059));
Q_MX04 U1397 ( .S0(n4396), .S1(n4397), .A0(n1059), .A1(n1056), .A2(n1055), .A3(n1054), .Z(n1060));
Q_MX02 U1398 ( .S(n4398), .A0(n1060), .A1(n1053), .Z(r32_mux_6_data[3]));
Q_MX02 U1399 ( .S(n4394), .A0(o_label7_data3[4]), .A1(o_label7_data4[4]), .Z(n1061));
Q_MX04 U1400 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[4]), .A1(o_label7_data0[4]), .A2(o_label7_data1[4]), .A3(o_label7_data2[4]), .Z(n1062));
Q_MX02 U1401 ( .S(n4396), .A0(n1062), .A1(n1061), .Z(n1063));
Q_MX08 U1402 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[4]), .A1(o_kdf_drbg_seed_0_state_key_255_224[4]), .A2(o_kdf_drbg_seed_0_state_key_223_192[4]), .A3(o_kdf_drbg_seed_0_state_key_191_160[4]), .A4(o_kdf_drbg_seed_0_state_key_159_128[4]), .A5(o_kdf_drbg_seed_0_state_key_127_96[4]), .A6(o_kdf_drbg_seed_0_state_key_95_64[4]), .A7(o_kdf_drbg_seed_0_state_key_63_32[4]), .Z(n1064));
Q_MX02 U1403 ( .S(n4397), .A0(n1064), .A1(n1063), .Z(n1065));
Q_MX04 U1404 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[4]), .A1(o_kdf_drbg_seed_0_state_value_127_96[4]), .A2(o_kdf_drbg_seed_0_state_value_95_64[4]), .A3(o_kdf_drbg_seed_0_state_value_63_32[4]), .Z(n1066));
Q_MX04 U1405 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[4]), .A1(o_kdf_drbg_seed_1_state_key_63_32[4]), .A2(o_kdf_drbg_seed_1_state_key_31_0[4]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[4]), .Z(n1067));
Q_MX04 U1406 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[4]), .A1(o_kdf_drbg_seed_1_state_key_191_160[4]), .A2(o_kdf_drbg_seed_1_state_key_159_128[4]), .A3(o_kdf_drbg_seed_1_state_key_127_96[4]), .Z(n1068));
Q_MX02 U1407 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[4]), .A1(o_kdf_drbg_seed_1_state_key_255_224[4]), .Z(n1069));
Q_AN02 U1408 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[4]), .Z(n1070));
Q_MX02 U1409 ( .S(n4395), .A0(n1070), .A1(n1069), .Z(n1071));
Q_MX04 U1410 ( .S0(n4396), .S1(n4397), .A0(n1071), .A1(n1068), .A2(n1067), .A3(n1066), .Z(n1072));
Q_MX02 U1411 ( .S(n4398), .A0(n1072), .A1(n1065), .Z(r32_mux_6_data[4]));
Q_MX02 U1412 ( .S(n4394), .A0(o_label7_data3[5]), .A1(o_label7_data4[5]), .Z(n1073));
Q_MX04 U1413 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[5]), .A1(o_label7_data0[5]), .A2(o_label7_data1[5]), .A3(o_label7_data2[5]), .Z(n1074));
Q_MX02 U1414 ( .S(n4396), .A0(n1074), .A1(n1073), .Z(n1075));
Q_MX08 U1415 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[5]), .A1(o_kdf_drbg_seed_0_state_key_255_224[5]), .A2(o_kdf_drbg_seed_0_state_key_223_192[5]), .A3(o_kdf_drbg_seed_0_state_key_191_160[5]), .A4(o_kdf_drbg_seed_0_state_key_159_128[5]), .A5(o_kdf_drbg_seed_0_state_key_127_96[5]), .A6(o_kdf_drbg_seed_0_state_key_95_64[5]), .A7(o_kdf_drbg_seed_0_state_key_63_32[5]), .Z(n1076));
Q_MX02 U1416 ( .S(n4397), .A0(n1076), .A1(n1075), .Z(n1077));
Q_MX04 U1417 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[5]), .A1(o_kdf_drbg_seed_0_state_value_127_96[5]), .A2(o_kdf_drbg_seed_0_state_value_95_64[5]), .A3(o_kdf_drbg_seed_0_state_value_63_32[5]), .Z(n1078));
Q_MX04 U1418 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[5]), .A1(o_kdf_drbg_seed_1_state_key_63_32[5]), .A2(o_kdf_drbg_seed_1_state_key_31_0[5]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[5]), .Z(n1079));
Q_MX04 U1419 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[5]), .A1(o_kdf_drbg_seed_1_state_key_191_160[5]), .A2(o_kdf_drbg_seed_1_state_key_159_128[5]), .A3(o_kdf_drbg_seed_1_state_key_127_96[5]), .Z(n1080));
Q_MX02 U1420 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[5]), .A1(o_kdf_drbg_seed_1_state_key_255_224[5]), .Z(n1081));
Q_AN02 U1421 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[5]), .Z(n1082));
Q_MX02 U1422 ( .S(n4395), .A0(n1082), .A1(n1081), .Z(n1083));
Q_MX04 U1423 ( .S0(n4396), .S1(n4397), .A0(n1083), .A1(n1080), .A2(n1079), .A3(n1078), .Z(n1084));
Q_MX02 U1424 ( .S(n4398), .A0(n1084), .A1(n1077), .Z(r32_mux_6_data[5]));
Q_MX02 U1425 ( .S(n4394), .A0(o_label7_data3[6]), .A1(o_label7_data4[6]), .Z(n1085));
Q_MX04 U1426 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[6]), .A1(o_label7_data0[6]), .A2(o_label7_data1[6]), .A3(o_label7_data2[6]), .Z(n1086));
Q_MX02 U1427 ( .S(n4396), .A0(n1086), .A1(n1085), .Z(n1087));
Q_MX08 U1428 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[6]), .A1(o_kdf_drbg_seed_0_state_key_255_224[6]), .A2(o_kdf_drbg_seed_0_state_key_223_192[6]), .A3(o_kdf_drbg_seed_0_state_key_191_160[6]), .A4(o_kdf_drbg_seed_0_state_key_159_128[6]), .A5(o_kdf_drbg_seed_0_state_key_127_96[6]), .A6(o_kdf_drbg_seed_0_state_key_95_64[6]), .A7(o_kdf_drbg_seed_0_state_key_63_32[6]), .Z(n1088));
Q_MX02 U1429 ( .S(n4397), .A0(n1088), .A1(n1087), .Z(n1089));
Q_MX04 U1430 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[6]), .A1(o_kdf_drbg_seed_0_state_value_127_96[6]), .A2(o_kdf_drbg_seed_0_state_value_95_64[6]), .A3(o_kdf_drbg_seed_0_state_value_63_32[6]), .Z(n1090));
Q_MX04 U1431 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[6]), .A1(o_kdf_drbg_seed_1_state_key_63_32[6]), .A2(o_kdf_drbg_seed_1_state_key_31_0[6]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[6]), .Z(n1091));
Q_MX04 U1432 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[6]), .A1(o_kdf_drbg_seed_1_state_key_191_160[6]), .A2(o_kdf_drbg_seed_1_state_key_159_128[6]), .A3(o_kdf_drbg_seed_1_state_key_127_96[6]), .Z(n1092));
Q_MX02 U1433 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[6]), .A1(o_kdf_drbg_seed_1_state_key_255_224[6]), .Z(n1093));
Q_AN02 U1434 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[6]), .Z(n1094));
Q_MX02 U1435 ( .S(n4395), .A0(n1094), .A1(n1093), .Z(n1095));
Q_MX04 U1436 ( .S0(n4396), .S1(n4397), .A0(n1095), .A1(n1092), .A2(n1091), .A3(n1090), .Z(n1096));
Q_MX02 U1437 ( .S(n4398), .A0(n1096), .A1(n1089), .Z(r32_mux_6_data[6]));
Q_MX02 U1438 ( .S(n4394), .A0(o_label7_data3[7]), .A1(o_label7_data4[7]), .Z(n1097));
Q_MX04 U1439 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[7]), .A1(o_label7_data0[7]), .A2(o_label7_data1[7]), .A3(o_label7_data2[7]), .Z(n1098));
Q_MX02 U1440 ( .S(n4396), .A0(n1098), .A1(n1097), .Z(n1099));
Q_MX08 U1441 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[7]), .A1(o_kdf_drbg_seed_0_state_key_255_224[7]), .A2(o_kdf_drbg_seed_0_state_key_223_192[7]), .A3(o_kdf_drbg_seed_0_state_key_191_160[7]), .A4(o_kdf_drbg_seed_0_state_key_159_128[7]), .A5(o_kdf_drbg_seed_0_state_key_127_96[7]), .A6(o_kdf_drbg_seed_0_state_key_95_64[7]), .A7(o_kdf_drbg_seed_0_state_key_63_32[7]), .Z(n1100));
Q_MX02 U1442 ( .S(n4397), .A0(n1100), .A1(n1099), .Z(n1101));
Q_MX04 U1443 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[7]), .A1(o_kdf_drbg_seed_0_state_value_127_96[7]), .A2(o_kdf_drbg_seed_0_state_value_95_64[7]), .A3(o_kdf_drbg_seed_0_state_value_63_32[7]), .Z(n1102));
Q_MX04 U1444 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[7]), .A1(o_kdf_drbg_seed_1_state_key_63_32[7]), .A2(o_kdf_drbg_seed_1_state_key_31_0[7]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[7]), .Z(n1103));
Q_MX04 U1445 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[7]), .A1(o_kdf_drbg_seed_1_state_key_191_160[7]), .A2(o_kdf_drbg_seed_1_state_key_159_128[7]), .A3(o_kdf_drbg_seed_1_state_key_127_96[7]), .Z(n1104));
Q_MX02 U1446 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[7]), .A1(o_kdf_drbg_seed_1_state_key_255_224[7]), .Z(n1105));
Q_AN02 U1447 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[7]), .Z(n1106));
Q_MX02 U1448 ( .S(n4395), .A0(n1106), .A1(n1105), .Z(n1107));
Q_MX04 U1449 ( .S0(n4396), .S1(n4397), .A0(n1107), .A1(n1104), .A2(n1103), .A3(n1102), .Z(n1108));
Q_MX02 U1450 ( .S(n4398), .A0(n1108), .A1(n1101), .Z(r32_mux_6_data[7]));
Q_MX02 U1451 ( .S(n4394), .A0(o_label7_data3[8]), .A1(o_label7_data4[8]), .Z(n1109));
Q_MX04 U1452 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[8]), .A1(o_label7_data0[8]), .A2(o_label7_data1[8]), .A3(o_label7_data2[8]), .Z(n1110));
Q_MX02 U1453 ( .S(n4396), .A0(n1110), .A1(n1109), .Z(n1111));
Q_MX08 U1454 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[8]), .A1(o_kdf_drbg_seed_0_state_key_255_224[8]), .A2(o_kdf_drbg_seed_0_state_key_223_192[8]), .A3(o_kdf_drbg_seed_0_state_key_191_160[8]), .A4(o_kdf_drbg_seed_0_state_key_159_128[8]), .A5(o_kdf_drbg_seed_0_state_key_127_96[8]), .A6(o_kdf_drbg_seed_0_state_key_95_64[8]), .A7(o_kdf_drbg_seed_0_state_key_63_32[8]), .Z(n1112));
Q_MX02 U1455 ( .S(n4397), .A0(n1112), .A1(n1111), .Z(n1113));
Q_MX04 U1456 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[8]), .A1(o_kdf_drbg_seed_0_state_value_127_96[8]), .A2(o_kdf_drbg_seed_0_state_value_95_64[8]), .A3(o_kdf_drbg_seed_0_state_value_63_32[8]), .Z(n1114));
Q_MX04 U1457 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[8]), .A1(o_kdf_drbg_seed_1_state_key_63_32[8]), .A2(o_kdf_drbg_seed_1_state_key_31_0[8]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[8]), .Z(n1115));
Q_MX04 U1458 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[8]), .A1(o_kdf_drbg_seed_1_state_key_191_160[8]), .A2(o_kdf_drbg_seed_1_state_key_159_128[8]), .A3(o_kdf_drbg_seed_1_state_key_127_96[8]), .Z(n1116));
Q_MX02 U1459 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[8]), .A1(o_kdf_drbg_seed_1_state_key_255_224[8]), .Z(n1117));
Q_AN02 U1460 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[8]), .Z(n1118));
Q_MX02 U1461 ( .S(n4395), .A0(n1118), .A1(n1117), .Z(n1119));
Q_MX04 U1462 ( .S0(n4396), .S1(n4397), .A0(n1119), .A1(n1116), .A2(n1115), .A3(n1114), .Z(n1120));
Q_MX02 U1463 ( .S(n4398), .A0(n1120), .A1(n1113), .Z(r32_mux_6_data[8]));
Q_MX02 U1464 ( .S(n4394), .A0(o_label7_data3[9]), .A1(o_label7_data4[9]), .Z(n1121));
Q_MX04 U1465 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[9]), .A1(o_label7_data0[9]), .A2(o_label7_data1[9]), .A3(o_label7_data2[9]), .Z(n1122));
Q_MX02 U1466 ( .S(n4396), .A0(n1122), .A1(n1121), .Z(n1123));
Q_MX08 U1467 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[9]), .A1(o_kdf_drbg_seed_0_state_key_255_224[9]), .A2(o_kdf_drbg_seed_0_state_key_223_192[9]), .A3(o_kdf_drbg_seed_0_state_key_191_160[9]), .A4(o_kdf_drbg_seed_0_state_key_159_128[9]), .A5(o_kdf_drbg_seed_0_state_key_127_96[9]), .A6(o_kdf_drbg_seed_0_state_key_95_64[9]), .A7(o_kdf_drbg_seed_0_state_key_63_32[9]), .Z(n1124));
Q_MX02 U1468 ( .S(n4397), .A0(n1124), .A1(n1123), .Z(n1125));
Q_MX04 U1469 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[9]), .A1(o_kdf_drbg_seed_0_state_value_127_96[9]), .A2(o_kdf_drbg_seed_0_state_value_95_64[9]), .A3(o_kdf_drbg_seed_0_state_value_63_32[9]), .Z(n1126));
Q_MX04 U1470 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[9]), .A1(o_kdf_drbg_seed_1_state_key_63_32[9]), .A2(o_kdf_drbg_seed_1_state_key_31_0[9]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[9]), .Z(n1127));
Q_MX04 U1471 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[9]), .A1(o_kdf_drbg_seed_1_state_key_191_160[9]), .A2(o_kdf_drbg_seed_1_state_key_159_128[9]), .A3(o_kdf_drbg_seed_1_state_key_127_96[9]), .Z(n1128));
Q_MX02 U1472 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[9]), .A1(o_kdf_drbg_seed_1_state_key_255_224[9]), .Z(n1129));
Q_AN02 U1473 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[9]), .Z(n1130));
Q_MX02 U1474 ( .S(n4395), .A0(n1130), .A1(n1129), .Z(n1131));
Q_MX04 U1475 ( .S0(n4396), .S1(n4397), .A0(n1131), .A1(n1128), .A2(n1127), .A3(n1126), .Z(n1132));
Q_MX02 U1476 ( .S(n4398), .A0(n1132), .A1(n1125), .Z(r32_mux_6_data[9]));
Q_MX02 U1477 ( .S(n4394), .A0(o_label7_data3[10]), .A1(o_label7_data4[10]), .Z(n1133));
Q_MX04 U1478 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[10]), .A1(o_label7_data0[10]), .A2(o_label7_data1[10]), .A3(o_label7_data2[10]), .Z(n1134));
Q_MX02 U1479 ( .S(n4396), .A0(n1134), .A1(n1133), .Z(n1135));
Q_MX08 U1480 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[10]), .A1(o_kdf_drbg_seed_0_state_key_255_224[10]), .A2(o_kdf_drbg_seed_0_state_key_223_192[10]), .A3(o_kdf_drbg_seed_0_state_key_191_160[10]), .A4(o_kdf_drbg_seed_0_state_key_159_128[10]), .A5(o_kdf_drbg_seed_0_state_key_127_96[10]), .A6(o_kdf_drbg_seed_0_state_key_95_64[10]), .A7(o_kdf_drbg_seed_0_state_key_63_32[10]), .Z(n1136));
Q_MX02 U1481 ( .S(n4397), .A0(n1136), .A1(n1135), .Z(n1137));
Q_MX04 U1482 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[10]), .A1(o_kdf_drbg_seed_0_state_value_127_96[10]), .A2(o_kdf_drbg_seed_0_state_value_95_64[10]), .A3(o_kdf_drbg_seed_0_state_value_63_32[10]), .Z(n1138));
Q_MX04 U1483 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[10]), .A1(o_kdf_drbg_seed_1_state_key_63_32[10]), .A2(o_kdf_drbg_seed_1_state_key_31_0[10]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[10]), .Z(n1139));
Q_MX04 U1484 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[10]), .A1(o_kdf_drbg_seed_1_state_key_191_160[10]), .A2(o_kdf_drbg_seed_1_state_key_159_128[10]), .A3(o_kdf_drbg_seed_1_state_key_127_96[10]), .Z(n1140));
Q_MX02 U1485 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[10]), .A1(o_kdf_drbg_seed_1_state_key_255_224[10]), .Z(n1141));
Q_AN02 U1486 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[10]), .Z(n1142));
Q_MX02 U1487 ( .S(n4395), .A0(n1142), .A1(n1141), .Z(n1143));
Q_MX04 U1488 ( .S0(n4396), .S1(n4397), .A0(n1143), .A1(n1140), .A2(n1139), .A3(n1138), .Z(n1144));
Q_MX02 U1489 ( .S(n4398), .A0(n1144), .A1(n1137), .Z(r32_mux_6_data[10]));
Q_MX02 U1490 ( .S(n4394), .A0(o_label7_data3[11]), .A1(o_label7_data4[11]), .Z(n1145));
Q_MX04 U1491 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[11]), .A1(o_label7_data0[11]), .A2(o_label7_data1[11]), .A3(o_label7_data2[11]), .Z(n1146));
Q_MX02 U1492 ( .S(n4396), .A0(n1146), .A1(n1145), .Z(n1147));
Q_MX08 U1493 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[11]), .A1(o_kdf_drbg_seed_0_state_key_255_224[11]), .A2(o_kdf_drbg_seed_0_state_key_223_192[11]), .A3(o_kdf_drbg_seed_0_state_key_191_160[11]), .A4(o_kdf_drbg_seed_0_state_key_159_128[11]), .A5(o_kdf_drbg_seed_0_state_key_127_96[11]), .A6(o_kdf_drbg_seed_0_state_key_95_64[11]), .A7(o_kdf_drbg_seed_0_state_key_63_32[11]), .Z(n1148));
Q_MX02 U1494 ( .S(n4397), .A0(n1148), .A1(n1147), .Z(n1149));
Q_MX04 U1495 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[11]), .A1(o_kdf_drbg_seed_0_state_value_127_96[11]), .A2(o_kdf_drbg_seed_0_state_value_95_64[11]), .A3(o_kdf_drbg_seed_0_state_value_63_32[11]), .Z(n1150));
Q_MX04 U1496 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[11]), .A1(o_kdf_drbg_seed_1_state_key_63_32[11]), .A2(o_kdf_drbg_seed_1_state_key_31_0[11]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[11]), .Z(n1151));
Q_MX04 U1497 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[11]), .A1(o_kdf_drbg_seed_1_state_key_191_160[11]), .A2(o_kdf_drbg_seed_1_state_key_159_128[11]), .A3(o_kdf_drbg_seed_1_state_key_127_96[11]), .Z(n1152));
Q_MX02 U1498 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[11]), .A1(o_kdf_drbg_seed_1_state_key_255_224[11]), .Z(n1153));
Q_AN02 U1499 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[11]), .Z(n1154));
Q_MX02 U1500 ( .S(n4395), .A0(n1154), .A1(n1153), .Z(n1155));
Q_MX04 U1501 ( .S0(n4396), .S1(n4397), .A0(n1155), .A1(n1152), .A2(n1151), .A3(n1150), .Z(n1156));
Q_MX02 U1502 ( .S(n4398), .A0(n1156), .A1(n1149), .Z(r32_mux_6_data[11]));
Q_MX02 U1503 ( .S(n4394), .A0(o_label7_data3[12]), .A1(o_label7_data4[12]), .Z(n1157));
Q_MX04 U1504 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[12]), .A1(o_label7_data0[12]), .A2(o_label7_data1[12]), .A3(o_label7_data2[12]), .Z(n1158));
Q_MX02 U1505 ( .S(n4396), .A0(n1158), .A1(n1157), .Z(n1159));
Q_MX08 U1506 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[12]), .A1(o_kdf_drbg_seed_0_state_key_255_224[12]), .A2(o_kdf_drbg_seed_0_state_key_223_192[12]), .A3(o_kdf_drbg_seed_0_state_key_191_160[12]), .A4(o_kdf_drbg_seed_0_state_key_159_128[12]), .A5(o_kdf_drbg_seed_0_state_key_127_96[12]), .A6(o_kdf_drbg_seed_0_state_key_95_64[12]), .A7(o_kdf_drbg_seed_0_state_key_63_32[12]), .Z(n1160));
Q_MX02 U1507 ( .S(n4397), .A0(n1160), .A1(n1159), .Z(n1161));
Q_MX04 U1508 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[12]), .A1(o_kdf_drbg_seed_0_state_value_127_96[12]), .A2(o_kdf_drbg_seed_0_state_value_95_64[12]), .A3(o_kdf_drbg_seed_0_state_value_63_32[12]), .Z(n1162));
Q_MX04 U1509 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[12]), .A1(o_kdf_drbg_seed_1_state_key_63_32[12]), .A2(o_kdf_drbg_seed_1_state_key_31_0[12]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[12]), .Z(n1163));
Q_MX04 U1510 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[12]), .A1(o_kdf_drbg_seed_1_state_key_191_160[12]), .A2(o_kdf_drbg_seed_1_state_key_159_128[12]), .A3(o_kdf_drbg_seed_1_state_key_127_96[12]), .Z(n1164));
Q_MX02 U1511 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[12]), .A1(o_kdf_drbg_seed_1_state_key_255_224[12]), .Z(n1165));
Q_AN02 U1512 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[12]), .Z(n1166));
Q_MX02 U1513 ( .S(n4395), .A0(n1166), .A1(n1165), .Z(n1167));
Q_MX04 U1514 ( .S0(n4396), .S1(n4397), .A0(n1167), .A1(n1164), .A2(n1163), .A3(n1162), .Z(n1168));
Q_MX02 U1515 ( .S(n4398), .A0(n1168), .A1(n1161), .Z(r32_mux_6_data[12]));
Q_MX02 U1516 ( .S(n4394), .A0(o_label7_data3[13]), .A1(o_label7_data4[13]), .Z(n1169));
Q_MX04 U1517 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[13]), .A1(o_label7_data0[13]), .A2(o_label7_data1[13]), .A3(o_label7_data2[13]), .Z(n1170));
Q_MX02 U1518 ( .S(n4396), .A0(n1170), .A1(n1169), .Z(n1171));
Q_MX08 U1519 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[13]), .A1(o_kdf_drbg_seed_0_state_key_255_224[13]), .A2(o_kdf_drbg_seed_0_state_key_223_192[13]), .A3(o_kdf_drbg_seed_0_state_key_191_160[13]), .A4(o_kdf_drbg_seed_0_state_key_159_128[13]), .A5(o_kdf_drbg_seed_0_state_key_127_96[13]), .A6(o_kdf_drbg_seed_0_state_key_95_64[13]), .A7(o_kdf_drbg_seed_0_state_key_63_32[13]), .Z(n1172));
Q_MX02 U1520 ( .S(n4397), .A0(n1172), .A1(n1171), .Z(n1173));
Q_MX04 U1521 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[13]), .A1(o_kdf_drbg_seed_0_state_value_127_96[13]), .A2(o_kdf_drbg_seed_0_state_value_95_64[13]), .A3(o_kdf_drbg_seed_0_state_value_63_32[13]), .Z(n1174));
Q_MX04 U1522 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[13]), .A1(o_kdf_drbg_seed_1_state_key_63_32[13]), .A2(o_kdf_drbg_seed_1_state_key_31_0[13]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[13]), .Z(n1175));
Q_MX04 U1523 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[13]), .A1(o_kdf_drbg_seed_1_state_key_191_160[13]), .A2(o_kdf_drbg_seed_1_state_key_159_128[13]), .A3(o_kdf_drbg_seed_1_state_key_127_96[13]), .Z(n1176));
Q_MX02 U1524 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[13]), .A1(o_kdf_drbg_seed_1_state_key_255_224[13]), .Z(n1177));
Q_AN02 U1525 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[13]), .Z(n1178));
Q_MX02 U1526 ( .S(n4395), .A0(n1178), .A1(n1177), .Z(n1179));
Q_MX04 U1527 ( .S0(n4396), .S1(n4397), .A0(n1179), .A1(n1176), .A2(n1175), .A3(n1174), .Z(n1180));
Q_MX02 U1528 ( .S(n4398), .A0(n1180), .A1(n1173), .Z(r32_mux_6_data[13]));
Q_MX02 U1529 ( .S(n4394), .A0(o_label7_data3[14]), .A1(o_label7_data4[14]), .Z(n1181));
Q_MX04 U1530 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[14]), .A1(o_label7_data0[14]), .A2(o_label7_data1[14]), .A3(o_label7_data2[14]), .Z(n1182));
Q_MX02 U1531 ( .S(n4396), .A0(n1182), .A1(n1181), .Z(n1183));
Q_MX08 U1532 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[14]), .A1(o_kdf_drbg_seed_0_state_key_255_224[14]), .A2(o_kdf_drbg_seed_0_state_key_223_192[14]), .A3(o_kdf_drbg_seed_0_state_key_191_160[14]), .A4(o_kdf_drbg_seed_0_state_key_159_128[14]), .A5(o_kdf_drbg_seed_0_state_key_127_96[14]), .A6(o_kdf_drbg_seed_0_state_key_95_64[14]), .A7(o_kdf_drbg_seed_0_state_key_63_32[14]), .Z(n1184));
Q_MX02 U1533 ( .S(n4397), .A0(n1184), .A1(n1183), .Z(n1185));
Q_MX04 U1534 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[14]), .A1(o_kdf_drbg_seed_0_state_value_127_96[14]), .A2(o_kdf_drbg_seed_0_state_value_95_64[14]), .A3(o_kdf_drbg_seed_0_state_value_63_32[14]), .Z(n1186));
Q_MX04 U1535 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[14]), .A1(o_kdf_drbg_seed_1_state_key_63_32[14]), .A2(o_kdf_drbg_seed_1_state_key_31_0[14]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[14]), .Z(n1187));
Q_MX04 U1536 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[14]), .A1(o_kdf_drbg_seed_1_state_key_191_160[14]), .A2(o_kdf_drbg_seed_1_state_key_159_128[14]), .A3(o_kdf_drbg_seed_1_state_key_127_96[14]), .Z(n1188));
Q_MX02 U1537 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[14]), .A1(o_kdf_drbg_seed_1_state_key_255_224[14]), .Z(n1189));
Q_AN02 U1538 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[14]), .Z(n1190));
Q_MX02 U1539 ( .S(n4395), .A0(n1190), .A1(n1189), .Z(n1191));
Q_MX04 U1540 ( .S0(n4396), .S1(n4397), .A0(n1191), .A1(n1188), .A2(n1187), .A3(n1186), .Z(n1192));
Q_MX02 U1541 ( .S(n4398), .A0(n1192), .A1(n1185), .Z(r32_mux_6_data[14]));
Q_MX02 U1542 ( .S(n4394), .A0(o_label7_data3[15]), .A1(o_label7_data4[15]), .Z(n1193));
Q_MX04 U1543 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_state_key_31_0[15]), .A1(o_label7_data0[15]), .A2(o_label7_data1[15]), .A3(o_label7_data2[15]), .Z(n1194));
Q_MX02 U1544 ( .S(n4396), .A0(n1194), .A1(n1193), .Z(n1195));
Q_MX08 U1545 ( .S0(n4394), .S1(n4395), .S2(n4396), .A0(o_kdf_drbg_seed_0_state_value_31_0[15]), .A1(o_kdf_drbg_seed_0_state_key_255_224[15]), .A2(o_kdf_drbg_seed_0_state_key_223_192[15]), .A3(o_kdf_drbg_seed_0_state_key_191_160[15]), .A4(o_kdf_drbg_seed_0_state_key_159_128[15]), .A5(o_kdf_drbg_seed_0_state_key_127_96[15]), .A6(o_kdf_drbg_seed_0_state_key_95_64[15]), .A7(o_kdf_drbg_seed_0_state_key_63_32[15]), .Z(n1196));
Q_MX02 U1546 ( .S(n4397), .A0(n1196), .A1(n1195), .Z(n1197));
Q_MX04 U1547 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_0_reseed_interval_0[15]), .A1(o_kdf_drbg_seed_0_state_value_127_96[15]), .A2(o_kdf_drbg_seed_0_state_value_95_64[15]), .A3(o_kdf_drbg_seed_0_state_value_63_32[15]), .Z(n1198));
Q_MX04 U1548 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_95_64[15]), .A1(o_kdf_drbg_seed_1_state_key_63_32[15]), .A2(o_kdf_drbg_seed_1_state_key_31_0[15]), .A3(o_kdf_drbg_seed_0_reseed_interval_1[15]), .Z(n1199));
Q_MX04 U1549 ( .S0(n4394), .S1(n4395), .A0(o_kdf_drbg_seed_1_state_key_223_192[15]), .A1(o_kdf_drbg_seed_1_state_key_191_160[15]), .A2(o_kdf_drbg_seed_1_state_key_159_128[15]), .A3(o_kdf_drbg_seed_1_state_key_127_96[15]), .Z(n1200));
Q_MX02 U1550 ( .S(n4394), .A0(o_kdf_drbg_seed_1_state_value_31_0[15]), .A1(o_kdf_drbg_seed_1_state_key_255_224[15]), .Z(n1201));
Q_AN02 U1551 ( .A0(n4394), .A1(o_kdf_drbg_seed_1_state_value_63_32[15]), .Z(n1202));
Q_MX02 U1552 ( .S(n4395), .A0(n1202), .A1(n1201), .Z(n1203));
Q_MX04 U1553 ( .S0(n4396), .S1(n4397), .A0(n1203), .A1(n1200), .A2(n1199), .A3(n1198), .Z(n1204));
Q_MX02 U1554 ( .S(n4398), .A0(n1204), .A1(n1197), .Z(r32_mux_6_data[15]));
Q_MX04 U1555 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[16]), .A1(o_label7_data1[16]), .A2(o_label7_data2[16]), .A3(o_label7_data3[16]), .Z(n1205));
Q_MX02 U1556 ( .S(n4401), .A0(n1205), .A1(o_label7_data4[16]), .Z(n1206));
Q_MX08 U1557 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[16]), .A1(o_kdf_drbg_seed_0_state_key_223_192[16]), .A2(o_kdf_drbg_seed_0_state_key_191_160[16]), .A3(o_kdf_drbg_seed_0_state_key_159_128[16]), .A4(o_kdf_drbg_seed_0_state_key_127_96[16]), .A5(o_kdf_drbg_seed_0_state_key_95_64[16]), .A6(o_kdf_drbg_seed_0_state_key_63_32[16]), .A7(o_kdf_drbg_seed_0_state_key_31_0[16]), .Z(n1207));
Q_MX02 U1558 ( .S(n4402), .A0(n1207), .A1(n1206), .Z(n1208));
Q_MX04 U1559 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[16]), .A1(o_kdf_drbg_seed_0_state_value_95_64[16]), .A2(o_kdf_drbg_seed_0_state_value_63_32[16]), .A3(o_kdf_drbg_seed_0_state_value_31_0[16]), .Z(n1209));
Q_MX04 U1560 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[16]), .A1(o_kdf_drbg_seed_1_state_key_63_32[16]), .A2(o_kdf_drbg_seed_1_state_key_31_0[16]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[16]), .Z(n1210));
Q_MX04 U1561 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[16]), .A1(o_kdf_drbg_seed_1_state_key_191_160[16]), .A2(o_kdf_drbg_seed_1_state_key_159_128[16]), .A3(o_kdf_drbg_seed_1_state_key_127_96[16]), .Z(n1211));
Q_MX02 U1562 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[16]), .A1(o_kdf_drbg_seed_1_state_key_255_224[16]), .Z(n1212));
Q_AN02 U1563 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[16]), .Z(n1213));
Q_MX02 U1564 ( .S(n4400), .A0(n1213), .A1(n1212), .Z(n1214));
Q_MX04 U1565 ( .S0(n4401), .S1(n4402), .A0(n1214), .A1(n1211), .A2(n1210), .A3(n1209), .Z(n1215));
Q_MX02 U1566 ( .S(n4403), .A0(n1215), .A1(n1208), .Z(r32_mux_6_data[16]));
Q_MX04 U1567 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[17]), .A1(o_label7_data1[17]), .A2(o_label7_data2[17]), .A3(o_label7_data3[17]), .Z(n1216));
Q_MX02 U1568 ( .S(n4401), .A0(n1216), .A1(o_label7_data4[17]), .Z(n1217));
Q_MX08 U1569 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[17]), .A1(o_kdf_drbg_seed_0_state_key_223_192[17]), .A2(o_kdf_drbg_seed_0_state_key_191_160[17]), .A3(o_kdf_drbg_seed_0_state_key_159_128[17]), .A4(o_kdf_drbg_seed_0_state_key_127_96[17]), .A5(o_kdf_drbg_seed_0_state_key_95_64[17]), .A6(o_kdf_drbg_seed_0_state_key_63_32[17]), .A7(o_kdf_drbg_seed_0_state_key_31_0[17]), .Z(n1218));
Q_MX02 U1570 ( .S(n4402), .A0(n1218), .A1(n1217), .Z(n1219));
Q_MX04 U1571 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[17]), .A1(o_kdf_drbg_seed_0_state_value_95_64[17]), .A2(o_kdf_drbg_seed_0_state_value_63_32[17]), .A3(o_kdf_drbg_seed_0_state_value_31_0[17]), .Z(n1220));
Q_MX04 U1572 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[17]), .A1(o_kdf_drbg_seed_1_state_key_63_32[17]), .A2(o_kdf_drbg_seed_1_state_key_31_0[17]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[17]), .Z(n1221));
Q_MX04 U1573 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[17]), .A1(o_kdf_drbg_seed_1_state_key_191_160[17]), .A2(o_kdf_drbg_seed_1_state_key_159_128[17]), .A3(o_kdf_drbg_seed_1_state_key_127_96[17]), .Z(n1222));
Q_MX02 U1574 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[17]), .A1(o_kdf_drbg_seed_1_state_key_255_224[17]), .Z(n1223));
Q_AN02 U1575 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[17]), .Z(n1224));
Q_MX02 U1576 ( .S(n4400), .A0(n1224), .A1(n1223), .Z(n1225));
Q_MX04 U1577 ( .S0(n4401), .S1(n4402), .A0(n1225), .A1(n1222), .A2(n1221), .A3(n1220), .Z(n1226));
Q_MX02 U1578 ( .S(n4403), .A0(n1226), .A1(n1219), .Z(r32_mux_6_data[17]));
Q_MX04 U1579 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[18]), .A1(o_label7_data1[18]), .A2(o_label7_data2[18]), .A3(o_label7_data3[18]), .Z(n1227));
Q_MX02 U1580 ( .S(n4401), .A0(n1227), .A1(o_label7_data4[18]), .Z(n1228));
Q_MX08 U1581 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[18]), .A1(o_kdf_drbg_seed_0_state_key_223_192[18]), .A2(o_kdf_drbg_seed_0_state_key_191_160[18]), .A3(o_kdf_drbg_seed_0_state_key_159_128[18]), .A4(o_kdf_drbg_seed_0_state_key_127_96[18]), .A5(o_kdf_drbg_seed_0_state_key_95_64[18]), .A6(o_kdf_drbg_seed_0_state_key_63_32[18]), .A7(o_kdf_drbg_seed_0_state_key_31_0[18]), .Z(n1229));
Q_MX02 U1582 ( .S(n4402), .A0(n1229), .A1(n1228), .Z(n1230));
Q_MX04 U1583 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[18]), .A1(o_kdf_drbg_seed_0_state_value_95_64[18]), .A2(o_kdf_drbg_seed_0_state_value_63_32[18]), .A3(o_kdf_drbg_seed_0_state_value_31_0[18]), .Z(n1231));
Q_MX04 U1584 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[18]), .A1(o_kdf_drbg_seed_1_state_key_63_32[18]), .A2(o_kdf_drbg_seed_1_state_key_31_0[18]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[18]), .Z(n1232));
Q_MX04 U1585 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[18]), .A1(o_kdf_drbg_seed_1_state_key_191_160[18]), .A2(o_kdf_drbg_seed_1_state_key_159_128[18]), .A3(o_kdf_drbg_seed_1_state_key_127_96[18]), .Z(n1233));
Q_MX02 U1586 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[18]), .A1(o_kdf_drbg_seed_1_state_key_255_224[18]), .Z(n1234));
Q_AN02 U1587 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[18]), .Z(n1235));
Q_MX02 U1588 ( .S(n4400), .A0(n1235), .A1(n1234), .Z(n1236));
Q_MX04 U1589 ( .S0(n4401), .S1(n4402), .A0(n1236), .A1(n1233), .A2(n1232), .A3(n1231), .Z(n1237));
Q_MX02 U1590 ( .S(n4403), .A0(n1237), .A1(n1230), .Z(r32_mux_6_data[18]));
Q_MX04 U1591 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[19]), .A1(o_label7_data1[19]), .A2(o_label7_data2[19]), .A3(o_label7_data3[19]), .Z(n1238));
Q_MX02 U1592 ( .S(n4401), .A0(n1238), .A1(o_label7_data4[19]), .Z(n1239));
Q_MX08 U1593 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[19]), .A1(o_kdf_drbg_seed_0_state_key_223_192[19]), .A2(o_kdf_drbg_seed_0_state_key_191_160[19]), .A3(o_kdf_drbg_seed_0_state_key_159_128[19]), .A4(o_kdf_drbg_seed_0_state_key_127_96[19]), .A5(o_kdf_drbg_seed_0_state_key_95_64[19]), .A6(o_kdf_drbg_seed_0_state_key_63_32[19]), .A7(o_kdf_drbg_seed_0_state_key_31_0[19]), .Z(n1240));
Q_MX02 U1594 ( .S(n4402), .A0(n1240), .A1(n1239), .Z(n1241));
Q_MX04 U1595 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[19]), .A1(o_kdf_drbg_seed_0_state_value_95_64[19]), .A2(o_kdf_drbg_seed_0_state_value_63_32[19]), .A3(o_kdf_drbg_seed_0_state_value_31_0[19]), .Z(n1242));
Q_MX04 U1596 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[19]), .A1(o_kdf_drbg_seed_1_state_key_63_32[19]), .A2(o_kdf_drbg_seed_1_state_key_31_0[19]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[19]), .Z(n1243));
Q_MX04 U1597 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[19]), .A1(o_kdf_drbg_seed_1_state_key_191_160[19]), .A2(o_kdf_drbg_seed_1_state_key_159_128[19]), .A3(o_kdf_drbg_seed_1_state_key_127_96[19]), .Z(n1244));
Q_MX02 U1598 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[19]), .A1(o_kdf_drbg_seed_1_state_key_255_224[19]), .Z(n1245));
Q_AN02 U1599 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[19]), .Z(n1246));
Q_MX02 U1600 ( .S(n4400), .A0(n1246), .A1(n1245), .Z(n1247));
Q_MX04 U1601 ( .S0(n4401), .S1(n4402), .A0(n1247), .A1(n1244), .A2(n1243), .A3(n1242), .Z(n1248));
Q_MX02 U1602 ( .S(n4403), .A0(n1248), .A1(n1241), .Z(r32_mux_6_data[19]));
Q_MX04 U1603 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[20]), .A1(o_label7_data1[20]), .A2(o_label7_data2[20]), .A3(o_label7_data3[20]), .Z(n1249));
Q_MX02 U1604 ( .S(n4401), .A0(n1249), .A1(o_label7_data4[20]), .Z(n1250));
Q_MX08 U1605 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[20]), .A1(o_kdf_drbg_seed_0_state_key_223_192[20]), .A2(o_kdf_drbg_seed_0_state_key_191_160[20]), .A3(o_kdf_drbg_seed_0_state_key_159_128[20]), .A4(o_kdf_drbg_seed_0_state_key_127_96[20]), .A5(o_kdf_drbg_seed_0_state_key_95_64[20]), .A6(o_kdf_drbg_seed_0_state_key_63_32[20]), .A7(o_kdf_drbg_seed_0_state_key_31_0[20]), .Z(n1251));
Q_MX02 U1606 ( .S(n4402), .A0(n1251), .A1(n1250), .Z(n1252));
Q_MX04 U1607 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[20]), .A1(o_kdf_drbg_seed_0_state_value_95_64[20]), .A2(o_kdf_drbg_seed_0_state_value_63_32[20]), .A3(o_kdf_drbg_seed_0_state_value_31_0[20]), .Z(n1253));
Q_MX04 U1608 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[20]), .A1(o_kdf_drbg_seed_1_state_key_63_32[20]), .A2(o_kdf_drbg_seed_1_state_key_31_0[20]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[20]), .Z(n1254));
Q_MX04 U1609 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[20]), .A1(o_kdf_drbg_seed_1_state_key_191_160[20]), .A2(o_kdf_drbg_seed_1_state_key_159_128[20]), .A3(o_kdf_drbg_seed_1_state_key_127_96[20]), .Z(n1255));
Q_MX02 U1610 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[20]), .A1(o_kdf_drbg_seed_1_state_key_255_224[20]), .Z(n1256));
Q_AN02 U1611 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[20]), .Z(n1257));
Q_MX02 U1612 ( .S(n4400), .A0(n1257), .A1(n1256), .Z(n1258));
Q_MX04 U1613 ( .S0(n4401), .S1(n4402), .A0(n1258), .A1(n1255), .A2(n1254), .A3(n1253), .Z(n1259));
Q_MX02 U1614 ( .S(n4403), .A0(n1259), .A1(n1252), .Z(r32_mux_6_data[20]));
Q_MX04 U1615 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[21]), .A1(o_label7_data1[21]), .A2(o_label7_data2[21]), .A3(o_label7_data3[21]), .Z(n1260));
Q_MX02 U1616 ( .S(n4401), .A0(n1260), .A1(o_label7_data4[21]), .Z(n1261));
Q_MX08 U1617 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[21]), .A1(o_kdf_drbg_seed_0_state_key_223_192[21]), .A2(o_kdf_drbg_seed_0_state_key_191_160[21]), .A3(o_kdf_drbg_seed_0_state_key_159_128[21]), .A4(o_kdf_drbg_seed_0_state_key_127_96[21]), .A5(o_kdf_drbg_seed_0_state_key_95_64[21]), .A6(o_kdf_drbg_seed_0_state_key_63_32[21]), .A7(o_kdf_drbg_seed_0_state_key_31_0[21]), .Z(n1262));
Q_MX02 U1618 ( .S(n4402), .A0(n1262), .A1(n1261), .Z(n1263));
Q_MX04 U1619 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[21]), .A1(o_kdf_drbg_seed_0_state_value_95_64[21]), .A2(o_kdf_drbg_seed_0_state_value_63_32[21]), .A3(o_kdf_drbg_seed_0_state_value_31_0[21]), .Z(n1264));
Q_MX04 U1620 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[21]), .A1(o_kdf_drbg_seed_1_state_key_63_32[21]), .A2(o_kdf_drbg_seed_1_state_key_31_0[21]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[21]), .Z(n1265));
Q_MX04 U1621 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[21]), .A1(o_kdf_drbg_seed_1_state_key_191_160[21]), .A2(o_kdf_drbg_seed_1_state_key_159_128[21]), .A3(o_kdf_drbg_seed_1_state_key_127_96[21]), .Z(n1266));
Q_MX02 U1622 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[21]), .A1(o_kdf_drbg_seed_1_state_key_255_224[21]), .Z(n1267));
Q_AN02 U1623 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[21]), .Z(n1268));
Q_MX02 U1624 ( .S(n4400), .A0(n1268), .A1(n1267), .Z(n1269));
Q_MX04 U1625 ( .S0(n4401), .S1(n4402), .A0(n1269), .A1(n1266), .A2(n1265), .A3(n1264), .Z(n1270));
Q_MX02 U1626 ( .S(n4403), .A0(n1270), .A1(n1263), .Z(r32_mux_6_data[21]));
Q_MX04 U1627 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[22]), .A1(o_label7_data1[22]), .A2(o_label7_data2[22]), .A3(o_label7_data3[22]), .Z(n1271));
Q_MX02 U1628 ( .S(n4401), .A0(n1271), .A1(o_label7_data4[22]), .Z(n1272));
Q_MX08 U1629 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[22]), .A1(o_kdf_drbg_seed_0_state_key_223_192[22]), .A2(o_kdf_drbg_seed_0_state_key_191_160[22]), .A3(o_kdf_drbg_seed_0_state_key_159_128[22]), .A4(o_kdf_drbg_seed_0_state_key_127_96[22]), .A5(o_kdf_drbg_seed_0_state_key_95_64[22]), .A6(o_kdf_drbg_seed_0_state_key_63_32[22]), .A7(o_kdf_drbg_seed_0_state_key_31_0[22]), .Z(n1273));
Q_MX02 U1630 ( .S(n4402), .A0(n1273), .A1(n1272), .Z(n1274));
Q_MX04 U1631 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[22]), .A1(o_kdf_drbg_seed_0_state_value_95_64[22]), .A2(o_kdf_drbg_seed_0_state_value_63_32[22]), .A3(o_kdf_drbg_seed_0_state_value_31_0[22]), .Z(n1275));
Q_MX04 U1632 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[22]), .A1(o_kdf_drbg_seed_1_state_key_63_32[22]), .A2(o_kdf_drbg_seed_1_state_key_31_0[22]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[22]), .Z(n1276));
Q_MX04 U1633 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[22]), .A1(o_kdf_drbg_seed_1_state_key_191_160[22]), .A2(o_kdf_drbg_seed_1_state_key_159_128[22]), .A3(o_kdf_drbg_seed_1_state_key_127_96[22]), .Z(n1277));
Q_MX02 U1634 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[22]), .A1(o_kdf_drbg_seed_1_state_key_255_224[22]), .Z(n1278));
Q_AN02 U1635 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[22]), .Z(n1279));
Q_MX02 U1636 ( .S(n4400), .A0(n1279), .A1(n1278), .Z(n1280));
Q_MX04 U1637 ( .S0(n4401), .S1(n4402), .A0(n1280), .A1(n1277), .A2(n1276), .A3(n1275), .Z(n1281));
Q_MX02 U1638 ( .S(n4403), .A0(n1281), .A1(n1274), .Z(r32_mux_6_data[22]));
Q_MX04 U1639 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[23]), .A1(o_label7_data1[23]), .A2(o_label7_data2[23]), .A3(o_label7_data3[23]), .Z(n1282));
Q_MX02 U1640 ( .S(n4401), .A0(n1282), .A1(o_label7_data4[23]), .Z(n1283));
Q_MX08 U1641 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[23]), .A1(o_kdf_drbg_seed_0_state_key_223_192[23]), .A2(o_kdf_drbg_seed_0_state_key_191_160[23]), .A3(o_kdf_drbg_seed_0_state_key_159_128[23]), .A4(o_kdf_drbg_seed_0_state_key_127_96[23]), .A5(o_kdf_drbg_seed_0_state_key_95_64[23]), .A6(o_kdf_drbg_seed_0_state_key_63_32[23]), .A7(o_kdf_drbg_seed_0_state_key_31_0[23]), .Z(n1284));
Q_MX02 U1642 ( .S(n4402), .A0(n1284), .A1(n1283), .Z(n1285));
Q_MX04 U1643 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[23]), .A1(o_kdf_drbg_seed_0_state_value_95_64[23]), .A2(o_kdf_drbg_seed_0_state_value_63_32[23]), .A3(o_kdf_drbg_seed_0_state_value_31_0[23]), .Z(n1286));
Q_MX04 U1644 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[23]), .A1(o_kdf_drbg_seed_1_state_key_63_32[23]), .A2(o_kdf_drbg_seed_1_state_key_31_0[23]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[23]), .Z(n1287));
Q_MX04 U1645 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[23]), .A1(o_kdf_drbg_seed_1_state_key_191_160[23]), .A2(o_kdf_drbg_seed_1_state_key_159_128[23]), .A3(o_kdf_drbg_seed_1_state_key_127_96[23]), .Z(n1288));
Q_MX02 U1646 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[23]), .A1(o_kdf_drbg_seed_1_state_key_255_224[23]), .Z(n1289));
Q_AN02 U1647 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[23]), .Z(n1290));
Q_MX02 U1648 ( .S(n4400), .A0(n1290), .A1(n1289), .Z(n1291));
Q_MX04 U1649 ( .S0(n4401), .S1(n4402), .A0(n1291), .A1(n1288), .A2(n1287), .A3(n1286), .Z(n1292));
Q_MX02 U1650 ( .S(n4403), .A0(n1292), .A1(n1285), .Z(r32_mux_6_data[23]));
Q_MX04 U1651 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[24]), .A1(o_label7_data1[24]), .A2(o_label7_data2[24]), .A3(o_label7_data3[24]), .Z(n1293));
Q_MX02 U1652 ( .S(n4401), .A0(n1293), .A1(o_label7_data4[24]), .Z(n1294));
Q_MX08 U1653 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[24]), .A1(o_kdf_drbg_seed_0_state_key_223_192[24]), .A2(o_kdf_drbg_seed_0_state_key_191_160[24]), .A3(o_kdf_drbg_seed_0_state_key_159_128[24]), .A4(o_kdf_drbg_seed_0_state_key_127_96[24]), .A5(o_kdf_drbg_seed_0_state_key_95_64[24]), .A6(o_kdf_drbg_seed_0_state_key_63_32[24]), .A7(o_kdf_drbg_seed_0_state_key_31_0[24]), .Z(n1295));
Q_MX02 U1654 ( .S(n4402), .A0(n1295), .A1(n1294), .Z(n1296));
Q_MX04 U1655 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[24]), .A1(o_kdf_drbg_seed_0_state_value_95_64[24]), .A2(o_kdf_drbg_seed_0_state_value_63_32[24]), .A3(o_kdf_drbg_seed_0_state_value_31_0[24]), .Z(n1297));
Q_MX04 U1656 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[24]), .A1(o_kdf_drbg_seed_1_state_key_63_32[24]), .A2(o_kdf_drbg_seed_1_state_key_31_0[24]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[24]), .Z(n1298));
Q_MX04 U1657 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[24]), .A1(o_kdf_drbg_seed_1_state_key_191_160[24]), .A2(o_kdf_drbg_seed_1_state_key_159_128[24]), .A3(o_kdf_drbg_seed_1_state_key_127_96[24]), .Z(n1299));
Q_MX02 U1658 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[24]), .A1(o_kdf_drbg_seed_1_state_key_255_224[24]), .Z(n1300));
Q_AN02 U1659 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[24]), .Z(n1301));
Q_MX02 U1660 ( .S(n4400), .A0(n1301), .A1(n1300), .Z(n1302));
Q_MX04 U1661 ( .S0(n4401), .S1(n4402), .A0(n1302), .A1(n1299), .A2(n1298), .A3(n1297), .Z(n1303));
Q_MX02 U1662 ( .S(n4403), .A0(n1303), .A1(n1296), .Z(r32_mux_6_data[24]));
Q_MX04 U1663 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[25]), .A1(o_label7_data1[25]), .A2(o_label7_data2[25]), .A3(o_label7_data3[25]), .Z(n1304));
Q_MX02 U1664 ( .S(n4401), .A0(n1304), .A1(o_label7_data4[25]), .Z(n1305));
Q_MX08 U1665 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[25]), .A1(o_kdf_drbg_seed_0_state_key_223_192[25]), .A2(o_kdf_drbg_seed_0_state_key_191_160[25]), .A3(o_kdf_drbg_seed_0_state_key_159_128[25]), .A4(o_kdf_drbg_seed_0_state_key_127_96[25]), .A5(o_kdf_drbg_seed_0_state_key_95_64[25]), .A6(o_kdf_drbg_seed_0_state_key_63_32[25]), .A7(o_kdf_drbg_seed_0_state_key_31_0[25]), .Z(n1306));
Q_MX02 U1666 ( .S(n4402), .A0(n1306), .A1(n1305), .Z(n1307));
Q_MX04 U1667 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[25]), .A1(o_kdf_drbg_seed_0_state_value_95_64[25]), .A2(o_kdf_drbg_seed_0_state_value_63_32[25]), .A3(o_kdf_drbg_seed_0_state_value_31_0[25]), .Z(n1308));
Q_MX04 U1668 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[25]), .A1(o_kdf_drbg_seed_1_state_key_63_32[25]), .A2(o_kdf_drbg_seed_1_state_key_31_0[25]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[25]), .Z(n1309));
Q_MX04 U1669 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[25]), .A1(o_kdf_drbg_seed_1_state_key_191_160[25]), .A2(o_kdf_drbg_seed_1_state_key_159_128[25]), .A3(o_kdf_drbg_seed_1_state_key_127_96[25]), .Z(n1310));
Q_MX02 U1670 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[25]), .A1(o_kdf_drbg_seed_1_state_key_255_224[25]), .Z(n1311));
Q_AN02 U1671 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[25]), .Z(n1312));
Q_MX02 U1672 ( .S(n4400), .A0(n1312), .A1(n1311), .Z(n1313));
Q_MX04 U1673 ( .S0(n4401), .S1(n4402), .A0(n1313), .A1(n1310), .A2(n1309), .A3(n1308), .Z(n1314));
Q_MX02 U1674 ( .S(n4403), .A0(n1314), .A1(n1307), .Z(r32_mux_6_data[25]));
Q_MX04 U1675 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[26]), .A1(o_label7_data1[26]), .A2(o_label7_data2[26]), .A3(o_label7_data3[26]), .Z(n1315));
Q_MX02 U1676 ( .S(n4401), .A0(n1315), .A1(o_label7_data4[26]), .Z(n1316));
Q_MX08 U1677 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[26]), .A1(o_kdf_drbg_seed_0_state_key_223_192[26]), .A2(o_kdf_drbg_seed_0_state_key_191_160[26]), .A3(o_kdf_drbg_seed_0_state_key_159_128[26]), .A4(o_kdf_drbg_seed_0_state_key_127_96[26]), .A5(o_kdf_drbg_seed_0_state_key_95_64[26]), .A6(o_kdf_drbg_seed_0_state_key_63_32[26]), .A7(o_kdf_drbg_seed_0_state_key_31_0[26]), .Z(n1317));
Q_MX02 U1678 ( .S(n4402), .A0(n1317), .A1(n1316), .Z(n1318));
Q_MX04 U1679 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[26]), .A1(o_kdf_drbg_seed_0_state_value_95_64[26]), .A2(o_kdf_drbg_seed_0_state_value_63_32[26]), .A3(o_kdf_drbg_seed_0_state_value_31_0[26]), .Z(n1319));
Q_MX04 U1680 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[26]), .A1(o_kdf_drbg_seed_1_state_key_63_32[26]), .A2(o_kdf_drbg_seed_1_state_key_31_0[26]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[26]), .Z(n1320));
Q_MX04 U1681 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[26]), .A1(o_kdf_drbg_seed_1_state_key_191_160[26]), .A2(o_kdf_drbg_seed_1_state_key_159_128[26]), .A3(o_kdf_drbg_seed_1_state_key_127_96[26]), .Z(n1321));
Q_MX02 U1682 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[26]), .A1(o_kdf_drbg_seed_1_state_key_255_224[26]), .Z(n1322));
Q_AN02 U1683 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[26]), .Z(n1323));
Q_MX02 U1684 ( .S(n4400), .A0(n1323), .A1(n1322), .Z(n1324));
Q_MX04 U1685 ( .S0(n4401), .S1(n4402), .A0(n1324), .A1(n1321), .A2(n1320), .A3(n1319), .Z(n1325));
Q_MX02 U1686 ( .S(n4403), .A0(n1325), .A1(n1318), .Z(r32_mux_6_data[26]));
Q_MX04 U1687 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[27]), .A1(o_label7_data1[27]), .A2(o_label7_data2[27]), .A3(o_label7_data3[27]), .Z(n1326));
Q_MX02 U1688 ( .S(n4401), .A0(n1326), .A1(o_label7_data4[27]), .Z(n1327));
Q_MX08 U1689 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[27]), .A1(o_kdf_drbg_seed_0_state_key_223_192[27]), .A2(o_kdf_drbg_seed_0_state_key_191_160[27]), .A3(o_kdf_drbg_seed_0_state_key_159_128[27]), .A4(o_kdf_drbg_seed_0_state_key_127_96[27]), .A5(o_kdf_drbg_seed_0_state_key_95_64[27]), .A6(o_kdf_drbg_seed_0_state_key_63_32[27]), .A7(o_kdf_drbg_seed_0_state_key_31_0[27]), .Z(n1328));
Q_MX02 U1690 ( .S(n4402), .A0(n1328), .A1(n1327), .Z(n1329));
Q_MX04 U1691 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[27]), .A1(o_kdf_drbg_seed_0_state_value_95_64[27]), .A2(o_kdf_drbg_seed_0_state_value_63_32[27]), .A3(o_kdf_drbg_seed_0_state_value_31_0[27]), .Z(n1330));
Q_MX04 U1692 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[27]), .A1(o_kdf_drbg_seed_1_state_key_63_32[27]), .A2(o_kdf_drbg_seed_1_state_key_31_0[27]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[27]), .Z(n1331));
Q_MX04 U1693 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[27]), .A1(o_kdf_drbg_seed_1_state_key_191_160[27]), .A2(o_kdf_drbg_seed_1_state_key_159_128[27]), .A3(o_kdf_drbg_seed_1_state_key_127_96[27]), .Z(n1332));
Q_MX02 U1694 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[27]), .A1(o_kdf_drbg_seed_1_state_key_255_224[27]), .Z(n1333));
Q_AN02 U1695 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[27]), .Z(n1334));
Q_MX02 U1696 ( .S(n4400), .A0(n1334), .A1(n1333), .Z(n1335));
Q_MX04 U1697 ( .S0(n4401), .S1(n4402), .A0(n1335), .A1(n1332), .A2(n1331), .A3(n1330), .Z(n1336));
Q_MX02 U1698 ( .S(n4403), .A0(n1336), .A1(n1329), .Z(r32_mux_6_data[27]));
Q_MX04 U1699 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[28]), .A1(o_label7_data1[28]), .A2(o_label7_data2[28]), .A3(o_label7_data3[28]), .Z(n1337));
Q_MX02 U1700 ( .S(n4401), .A0(n1337), .A1(o_label7_data4[28]), .Z(n1338));
Q_MX08 U1701 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[28]), .A1(o_kdf_drbg_seed_0_state_key_223_192[28]), .A2(o_kdf_drbg_seed_0_state_key_191_160[28]), .A3(o_kdf_drbg_seed_0_state_key_159_128[28]), .A4(o_kdf_drbg_seed_0_state_key_127_96[28]), .A5(o_kdf_drbg_seed_0_state_key_95_64[28]), .A6(o_kdf_drbg_seed_0_state_key_63_32[28]), .A7(o_kdf_drbg_seed_0_state_key_31_0[28]), .Z(n1339));
Q_MX02 U1702 ( .S(n4402), .A0(n1339), .A1(n1338), .Z(n1340));
Q_MX04 U1703 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[28]), .A1(o_kdf_drbg_seed_0_state_value_95_64[28]), .A2(o_kdf_drbg_seed_0_state_value_63_32[28]), .A3(o_kdf_drbg_seed_0_state_value_31_0[28]), .Z(n1341));
Q_MX04 U1704 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[28]), .A1(o_kdf_drbg_seed_1_state_key_63_32[28]), .A2(o_kdf_drbg_seed_1_state_key_31_0[28]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[28]), .Z(n1342));
Q_MX04 U1705 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[28]), .A1(o_kdf_drbg_seed_1_state_key_191_160[28]), .A2(o_kdf_drbg_seed_1_state_key_159_128[28]), .A3(o_kdf_drbg_seed_1_state_key_127_96[28]), .Z(n1343));
Q_MX02 U1706 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[28]), .A1(o_kdf_drbg_seed_1_state_key_255_224[28]), .Z(n1344));
Q_AN02 U1707 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[28]), .Z(n1345));
Q_MX02 U1708 ( .S(n4400), .A0(n1345), .A1(n1344), .Z(n1346));
Q_MX04 U1709 ( .S0(n4401), .S1(n4402), .A0(n1346), .A1(n1343), .A2(n1342), .A3(n1341), .Z(n1347));
Q_MX02 U1710 ( .S(n4403), .A0(n1347), .A1(n1340), .Z(r32_mux_6_data[28]));
Q_MX04 U1711 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[29]), .A1(o_label7_data1[29]), .A2(o_label7_data2[29]), .A3(o_label7_data3[29]), .Z(n1348));
Q_MX02 U1712 ( .S(n4401), .A0(n1348), .A1(o_label7_data4[29]), .Z(n1349));
Q_MX08 U1713 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[29]), .A1(o_kdf_drbg_seed_0_state_key_223_192[29]), .A2(o_kdf_drbg_seed_0_state_key_191_160[29]), .A3(o_kdf_drbg_seed_0_state_key_159_128[29]), .A4(o_kdf_drbg_seed_0_state_key_127_96[29]), .A5(o_kdf_drbg_seed_0_state_key_95_64[29]), .A6(o_kdf_drbg_seed_0_state_key_63_32[29]), .A7(o_kdf_drbg_seed_0_state_key_31_0[29]), .Z(n1350));
Q_MX02 U1714 ( .S(n4402), .A0(n1350), .A1(n1349), .Z(n1351));
Q_MX04 U1715 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[29]), .A1(o_kdf_drbg_seed_0_state_value_95_64[29]), .A2(o_kdf_drbg_seed_0_state_value_63_32[29]), .A3(o_kdf_drbg_seed_0_state_value_31_0[29]), .Z(n1352));
Q_MX04 U1716 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[29]), .A1(o_kdf_drbg_seed_1_state_key_63_32[29]), .A2(o_kdf_drbg_seed_1_state_key_31_0[29]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[29]), .Z(n1353));
Q_MX04 U1717 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[29]), .A1(o_kdf_drbg_seed_1_state_key_191_160[29]), .A2(o_kdf_drbg_seed_1_state_key_159_128[29]), .A3(o_kdf_drbg_seed_1_state_key_127_96[29]), .Z(n1354));
Q_MX02 U1718 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[29]), .A1(o_kdf_drbg_seed_1_state_key_255_224[29]), .Z(n1355));
Q_AN02 U1719 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[29]), .Z(n1356));
Q_MX02 U1720 ( .S(n4400), .A0(n1356), .A1(n1355), .Z(n1357));
Q_MX04 U1721 ( .S0(n4401), .S1(n4402), .A0(n1357), .A1(n1354), .A2(n1353), .A3(n1352), .Z(n1358));
Q_MX02 U1722 ( .S(n4403), .A0(n1358), .A1(n1351), .Z(r32_mux_6_data[29]));
Q_MX04 U1723 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[30]), .A1(o_label7_data1[30]), .A2(o_label7_data2[30]), .A3(o_label7_data3[30]), .Z(n1359));
Q_MX02 U1724 ( .S(n4401), .A0(n1359), .A1(o_label7_data4[30]), .Z(n1360));
Q_MX08 U1725 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[30]), .A1(o_kdf_drbg_seed_0_state_key_223_192[30]), .A2(o_kdf_drbg_seed_0_state_key_191_160[30]), .A3(o_kdf_drbg_seed_0_state_key_159_128[30]), .A4(o_kdf_drbg_seed_0_state_key_127_96[30]), .A5(o_kdf_drbg_seed_0_state_key_95_64[30]), .A6(o_kdf_drbg_seed_0_state_key_63_32[30]), .A7(o_kdf_drbg_seed_0_state_key_31_0[30]), .Z(n1361));
Q_MX02 U1726 ( .S(n4402), .A0(n1361), .A1(n1360), .Z(n1362));
Q_MX04 U1727 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[30]), .A1(o_kdf_drbg_seed_0_state_value_95_64[30]), .A2(o_kdf_drbg_seed_0_state_value_63_32[30]), .A3(o_kdf_drbg_seed_0_state_value_31_0[30]), .Z(n1363));
Q_MX04 U1728 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[30]), .A1(o_kdf_drbg_seed_1_state_key_63_32[30]), .A2(o_kdf_drbg_seed_1_state_key_31_0[30]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[30]), .Z(n1364));
Q_MX04 U1729 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[30]), .A1(o_kdf_drbg_seed_1_state_key_191_160[30]), .A2(o_kdf_drbg_seed_1_state_key_159_128[30]), .A3(o_kdf_drbg_seed_1_state_key_127_96[30]), .Z(n1365));
Q_MX02 U1730 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[30]), .A1(o_kdf_drbg_seed_1_state_key_255_224[30]), .Z(n1366));
Q_AN02 U1731 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[30]), .Z(n1367));
Q_MX02 U1732 ( .S(n4400), .A0(n1367), .A1(n1366), .Z(n1368));
Q_MX04 U1733 ( .S0(n4401), .S1(n4402), .A0(n1368), .A1(n1365), .A2(n1364), .A3(n1363), .Z(n1369));
Q_MX02 U1734 ( .S(n4403), .A0(n1369), .A1(n1362), .Z(r32_mux_6_data[30]));
Q_MX04 U1735 ( .S0(n4399), .S1(n4400), .A0(o_label7_data0[31]), .A1(o_label7_data1[31]), .A2(o_label7_data2[31]), .A3(o_label7_data3[31]), .Z(n1370));
Q_MX02 U1736 ( .S(n4401), .A0(n1370), .A1(o_label7_data4[31]), .Z(n1371));
Q_MX08 U1737 ( .S0(n4399), .S1(n4400), .S2(n4401), .A0(o_kdf_drbg_seed_0_state_key_255_224[31]), .A1(o_kdf_drbg_seed_0_state_key_223_192[31]), .A2(o_kdf_drbg_seed_0_state_key_191_160[31]), .A3(o_kdf_drbg_seed_0_state_key_159_128[31]), .A4(o_kdf_drbg_seed_0_state_key_127_96[31]), .A5(o_kdf_drbg_seed_0_state_key_95_64[31]), .A6(o_kdf_drbg_seed_0_state_key_63_32[31]), .A7(o_kdf_drbg_seed_0_state_key_31_0[31]), .Z(n1372));
Q_MX02 U1738 ( .S(n4402), .A0(n1372), .A1(n1371), .Z(n1373));
Q_MX04 U1739 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_0_state_value_127_96[31]), .A1(o_kdf_drbg_seed_0_state_value_95_64[31]), .A2(o_kdf_drbg_seed_0_state_value_63_32[31]), .A3(o_kdf_drbg_seed_0_state_value_31_0[31]), .Z(n1374));
Q_MX04 U1740 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_95_64[31]), .A1(o_kdf_drbg_seed_1_state_key_63_32[31]), .A2(o_kdf_drbg_seed_1_state_key_31_0[31]), .A3(o_kdf_drbg_seed_0_reseed_interval_0[31]), .Z(n1375));
Q_MX04 U1741 ( .S0(n4399), .S1(n4400), .A0(o_kdf_drbg_seed_1_state_key_223_192[31]), .A1(o_kdf_drbg_seed_1_state_key_191_160[31]), .A2(o_kdf_drbg_seed_1_state_key_159_128[31]), .A3(o_kdf_drbg_seed_1_state_key_127_96[31]), .Z(n1376));
Q_MX02 U1742 ( .S(n4399), .A0(o_kdf_drbg_seed_1_state_value_31_0[31]), .A1(o_kdf_drbg_seed_1_state_key_255_224[31]), .Z(n1377));
Q_AN02 U1743 ( .A0(n4399), .A1(o_kdf_drbg_seed_1_state_value_63_32[31]), .Z(n1378));
Q_MX02 U1744 ( .S(n4400), .A0(n1378), .A1(n1377), .Z(n1379));
Q_MX04 U1745 ( .S0(n4401), .S1(n4402), .A0(n1379), .A1(n1376), .A2(n1375), .A3(n1374), .Z(n1380));
Q_MX02 U1746 ( .S(n4403), .A0(n1380), .A1(n1373), .Z(r32_mux_6_data[31]));
Q_MX03 U1747 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[0]), .A1(o_label4_data6[0]), .A2(o_label4_data7[0]), .Z(n1381));
Q_MX04 U1748 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[0]), .A1(o_label4_data2[0]), .A2(o_label4_data3[0]), .A3(o_label4_data4[0]), .Z(n1382));
Q_MX02 U1749 ( .S(n4406), .A0(n1382), .A1(n1381), .Z(n1383));
Q_MX08 U1750 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[0]), .A1(o_label5_data3[0]), .A2(o_label5_data4[0]), .A3(o_label5_data5[0]), .A4(o_label5_data6[0]), .A5(o_label5_data7[0]), .A6(o_label5_config[0]), .A7(o_label4_data0[0]), .Z(n1384));
Q_MX02 U1751 ( .S(n4407), .A0(n1384), .A1(n1383), .Z(n1385));
Q_MX04 U1752 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[0]), .A1(o_label6_config[0]), .A2(o_label5_data0[0]), .A3(o_label5_data1[0]), .Z(n1386));
Q_MX04 U1753 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[0]), .A1(o_label6_data4[0]), .A2(o_label6_data5[0]), .A3(o_label6_data6[0]), .Z(n1387));
Q_MX04 U1754 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[0]), .A1(o_label6_data0[0]), .A2(o_label6_data1[0]), .A3(o_label6_data2[0]), .Z(n1388));
Q_MX02 U1755 ( .S(n4404), .A0(o_label7_data6[0]), .A1(o_label7_data7[0]), .Z(n1389));
Q_AN02 U1756 ( .A0(n4404), .A1(o_label7_data5[0]), .Z(n1390));
Q_MX02 U1757 ( .S(n4405), .A0(n1390), .A1(n1389), .Z(n1391));
Q_MX04 U1758 ( .S0(n4406), .S1(n4407), .A0(n1391), .A1(n1388), .A2(n1387), .A3(n1386), .Z(n1392));
Q_MX02 U1759 ( .S(n4408), .A0(n1392), .A1(n1385), .Z(r32_mux_5_data[0]));
Q_MX03 U1760 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[1]), .A1(o_label4_data6[1]), .A2(o_label4_data7[1]), .Z(n1393));
Q_MX04 U1761 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[1]), .A1(o_label4_data2[1]), .A2(o_label4_data3[1]), .A3(o_label4_data4[1]), .Z(n1394));
Q_MX02 U1762 ( .S(n4406), .A0(n1394), .A1(n1393), .Z(n1395));
Q_MX08 U1763 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[1]), .A1(o_label5_data3[1]), .A2(o_label5_data4[1]), .A3(o_label5_data5[1]), .A4(o_label5_data6[1]), .A5(o_label5_data7[1]), .A6(o_label5_config[1]), .A7(o_label4_data0[1]), .Z(n1396));
Q_MX02 U1764 ( .S(n4407), .A0(n1396), .A1(n1395), .Z(n1397));
Q_MX04 U1765 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[1]), .A1(o_label6_config[1]), .A2(o_label5_data0[1]), .A3(o_label5_data1[1]), .Z(n1398));
Q_MX04 U1766 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[1]), .A1(o_label6_data4[1]), .A2(o_label6_data5[1]), .A3(o_label6_data6[1]), .Z(n1399));
Q_MX04 U1767 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[1]), .A1(o_label6_data0[1]), .A2(o_label6_data1[1]), .A3(o_label6_data2[1]), .Z(n1400));
Q_MX02 U1768 ( .S(n4404), .A0(o_label7_data6[1]), .A1(o_label7_data7[1]), .Z(n1401));
Q_AN02 U1769 ( .A0(n4404), .A1(o_label7_data5[1]), .Z(n1402));
Q_MX02 U1770 ( .S(n4405), .A0(n1402), .A1(n1401), .Z(n1403));
Q_MX04 U1771 ( .S0(n4406), .S1(n4407), .A0(n1403), .A1(n1400), .A2(n1399), .A3(n1398), .Z(n1404));
Q_MX02 U1772 ( .S(n4408), .A0(n1404), .A1(n1397), .Z(r32_mux_5_data[1]));
Q_MX03 U1773 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[2]), .A1(o_label4_data6[2]), .A2(o_label4_data7[2]), .Z(n1405));
Q_MX04 U1774 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[2]), .A1(o_label4_data2[2]), .A2(o_label4_data3[2]), .A3(o_label4_data4[2]), .Z(n1406));
Q_MX02 U1775 ( .S(n4406), .A0(n1406), .A1(n1405), .Z(n1407));
Q_MX08 U1776 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[2]), .A1(o_label5_data3[2]), .A2(o_label5_data4[2]), .A3(o_label5_data5[2]), .A4(o_label5_data6[2]), .A5(o_label5_data7[2]), .A6(o_label5_config[2]), .A7(o_label4_data0[2]), .Z(n1408));
Q_MX02 U1777 ( .S(n4407), .A0(n1408), .A1(n1407), .Z(n1409));
Q_MX04 U1778 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[2]), .A1(o_label6_config[2]), .A2(o_label5_data0[2]), .A3(o_label5_data1[2]), .Z(n1410));
Q_MX04 U1779 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[2]), .A1(o_label6_data4[2]), .A2(o_label6_data5[2]), .A3(o_label6_data6[2]), .Z(n1411));
Q_MX04 U1780 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[2]), .A1(o_label6_data0[2]), .A2(o_label6_data1[2]), .A3(o_label6_data2[2]), .Z(n1412));
Q_MX02 U1781 ( .S(n4404), .A0(o_label7_data6[2]), .A1(o_label7_data7[2]), .Z(n1413));
Q_AN02 U1782 ( .A0(n4404), .A1(o_label7_data5[2]), .Z(n1414));
Q_MX02 U1783 ( .S(n4405), .A0(n1414), .A1(n1413), .Z(n1415));
Q_MX04 U1784 ( .S0(n4406), .S1(n4407), .A0(n1415), .A1(n1412), .A2(n1411), .A3(n1410), .Z(n1416));
Q_MX02 U1785 ( .S(n4408), .A0(n1416), .A1(n1409), .Z(r32_mux_5_data[2]));
Q_MX03 U1786 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[3]), .A1(o_label4_data6[3]), .A2(o_label4_data7[3]), .Z(n1417));
Q_MX04 U1787 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[3]), .A1(o_label4_data2[3]), .A2(o_label4_data3[3]), .A3(o_label4_data4[3]), .Z(n1418));
Q_MX02 U1788 ( .S(n4406), .A0(n1418), .A1(n1417), .Z(n1419));
Q_MX08 U1789 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[3]), .A1(o_label5_data3[3]), .A2(o_label5_data4[3]), .A3(o_label5_data5[3]), .A4(o_label5_data6[3]), .A5(o_label5_data7[3]), .A6(o_label5_config[3]), .A7(o_label4_data0[3]), .Z(n1420));
Q_MX02 U1790 ( .S(n4407), .A0(n1420), .A1(n1419), .Z(n1421));
Q_MX04 U1791 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[3]), .A1(o_label6_config[3]), .A2(o_label5_data0[3]), .A3(o_label5_data1[3]), .Z(n1422));
Q_MX04 U1792 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[3]), .A1(o_label6_data4[3]), .A2(o_label6_data5[3]), .A3(o_label6_data6[3]), .Z(n1423));
Q_MX04 U1793 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[3]), .A1(o_label6_data0[3]), .A2(o_label6_data1[3]), .A3(o_label6_data2[3]), .Z(n1424));
Q_MX02 U1794 ( .S(n4404), .A0(o_label7_data6[3]), .A1(o_label7_data7[3]), .Z(n1425));
Q_AN02 U1795 ( .A0(n4404), .A1(o_label7_data5[3]), .Z(n1426));
Q_MX02 U1796 ( .S(n4405), .A0(n1426), .A1(n1425), .Z(n1427));
Q_MX04 U1797 ( .S0(n4406), .S1(n4407), .A0(n1427), .A1(n1424), .A2(n1423), .A3(n1422), .Z(n1428));
Q_MX02 U1798 ( .S(n4408), .A0(n1428), .A1(n1421), .Z(r32_mux_5_data[3]));
Q_MX03 U1799 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[4]), .A1(o_label4_data6[4]), .A2(o_label4_data7[4]), .Z(n1429));
Q_MX04 U1800 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[4]), .A1(o_label4_data2[4]), .A2(o_label4_data3[4]), .A3(o_label4_data4[4]), .Z(n1430));
Q_MX02 U1801 ( .S(n4406), .A0(n1430), .A1(n1429), .Z(n1431));
Q_MX08 U1802 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[4]), .A1(o_label5_data3[4]), .A2(o_label5_data4[4]), .A3(o_label5_data5[4]), .A4(o_label5_data6[4]), .A5(o_label5_data7[4]), .A6(o_label5_config[4]), .A7(o_label4_data0[4]), .Z(n1432));
Q_MX02 U1803 ( .S(n4407), .A0(n1432), .A1(n1431), .Z(n1433));
Q_MX04 U1804 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[4]), .A1(o_label6_config[4]), .A2(o_label5_data0[4]), .A3(o_label5_data1[4]), .Z(n1434));
Q_MX04 U1805 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[4]), .A1(o_label6_data4[4]), .A2(o_label6_data5[4]), .A3(o_label6_data6[4]), .Z(n1435));
Q_MX04 U1806 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[4]), .A1(o_label6_data0[4]), .A2(o_label6_data1[4]), .A3(o_label6_data2[4]), .Z(n1436));
Q_MX02 U1807 ( .S(n4404), .A0(o_label7_data6[4]), .A1(o_label7_data7[4]), .Z(n1437));
Q_AN02 U1808 ( .A0(n4404), .A1(o_label7_data5[4]), .Z(n1438));
Q_MX02 U1809 ( .S(n4405), .A0(n1438), .A1(n1437), .Z(n1439));
Q_MX04 U1810 ( .S0(n4406), .S1(n4407), .A0(n1439), .A1(n1436), .A2(n1435), .A3(n1434), .Z(n1440));
Q_MX02 U1811 ( .S(n4408), .A0(n1440), .A1(n1433), .Z(r32_mux_5_data[4]));
Q_MX03 U1812 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[5]), .A1(o_label4_data6[5]), .A2(o_label4_data7[5]), .Z(n1441));
Q_MX04 U1813 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[5]), .A1(o_label4_data2[5]), .A2(o_label4_data3[5]), .A3(o_label4_data4[5]), .Z(n1442));
Q_MX02 U1814 ( .S(n4406), .A0(n1442), .A1(n1441), .Z(n1443));
Q_MX08 U1815 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[5]), .A1(o_label5_data3[5]), .A2(o_label5_data4[5]), .A3(o_label5_data5[5]), .A4(o_label5_data6[5]), .A5(o_label5_data7[5]), .A6(o_label5_config[5]), .A7(o_label4_data0[5]), .Z(n1444));
Q_MX02 U1816 ( .S(n4407), .A0(n1444), .A1(n1443), .Z(n1445));
Q_MX04 U1817 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[5]), .A1(o_label6_config[5]), .A2(o_label5_data0[5]), .A3(o_label5_data1[5]), .Z(n1446));
Q_MX04 U1818 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[5]), .A1(o_label6_data4[5]), .A2(o_label6_data5[5]), .A3(o_label6_data6[5]), .Z(n1447));
Q_MX04 U1819 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[5]), .A1(o_label6_data0[5]), .A2(o_label6_data1[5]), .A3(o_label6_data2[5]), .Z(n1448));
Q_MX02 U1820 ( .S(n4404), .A0(o_label7_data6[5]), .A1(o_label7_data7[5]), .Z(n1449));
Q_AN02 U1821 ( .A0(n4404), .A1(o_label7_data5[5]), .Z(n1450));
Q_MX02 U1822 ( .S(n4405), .A0(n1450), .A1(n1449), .Z(n1451));
Q_MX04 U1823 ( .S0(n4406), .S1(n4407), .A0(n1451), .A1(n1448), .A2(n1447), .A3(n1446), .Z(n1452));
Q_MX02 U1824 ( .S(n4408), .A0(n1452), .A1(n1445), .Z(r32_mux_5_data[5]));
Q_MX03 U1825 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[6]), .A1(o_label4_data6[6]), .A2(o_label4_data7[6]), .Z(n1453));
Q_MX04 U1826 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[6]), .A1(o_label4_data2[6]), .A2(o_label4_data3[6]), .A3(o_label4_data4[6]), .Z(n1454));
Q_MX02 U1827 ( .S(n4406), .A0(n1454), .A1(n1453), .Z(n1455));
Q_MX08 U1828 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[6]), .A1(o_label5_data3[6]), .A2(o_label5_data4[6]), .A3(o_label5_data5[6]), .A4(o_label5_data6[6]), .A5(o_label5_data7[6]), .A6(o_label5_config[6]), .A7(o_label4_data0[6]), .Z(n1456));
Q_MX02 U1829 ( .S(n4407), .A0(n1456), .A1(n1455), .Z(n1457));
Q_MX04 U1830 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[6]), .A1(o_label6_config[6]), .A2(o_label5_data0[6]), .A3(o_label5_data1[6]), .Z(n1458));
Q_MX04 U1831 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[6]), .A1(o_label6_data4[6]), .A2(o_label6_data5[6]), .A3(o_label6_data6[6]), .Z(n1459));
Q_MX04 U1832 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[6]), .A1(o_label6_data0[6]), .A2(o_label6_data1[6]), .A3(o_label6_data2[6]), .Z(n1460));
Q_MX02 U1833 ( .S(n4404), .A0(o_label7_data6[6]), .A1(o_label7_data7[6]), .Z(n1461));
Q_AN02 U1834 ( .A0(n4404), .A1(o_label7_data5[6]), .Z(n1462));
Q_MX02 U1835 ( .S(n4405), .A0(n1462), .A1(n1461), .Z(n1463));
Q_MX04 U1836 ( .S0(n4406), .S1(n4407), .A0(n1463), .A1(n1460), .A2(n1459), .A3(n1458), .Z(n1464));
Q_MX02 U1837 ( .S(n4408), .A0(n1464), .A1(n1457), .Z(r32_mux_5_data[6]));
Q_MX03 U1838 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[7]), .A1(o_label4_data6[7]), .A2(o_label4_data7[7]), .Z(n1465));
Q_MX04 U1839 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[7]), .A1(o_label4_data2[7]), .A2(o_label4_data3[7]), .A3(o_label4_data4[7]), .Z(n1466));
Q_MX02 U1840 ( .S(n4406), .A0(n1466), .A1(n1465), .Z(n1467));
Q_MX08 U1841 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[7]), .A1(o_label5_data3[7]), .A2(o_label5_data4[7]), .A3(o_label5_data5[7]), .A4(o_label5_data6[7]), .A5(o_label5_data7[7]), .A6(o_label5_config[7]), .A7(o_label4_data0[7]), .Z(n1468));
Q_MX02 U1842 ( .S(n4407), .A0(n1468), .A1(n1467), .Z(n1469));
Q_MX04 U1843 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[7]), .A1(o_label6_config[7]), .A2(o_label5_data0[7]), .A3(o_label5_data1[7]), .Z(n1470));
Q_MX04 U1844 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[7]), .A1(o_label6_data4[7]), .A2(o_label6_data5[7]), .A3(o_label6_data6[7]), .Z(n1471));
Q_MX04 U1845 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[7]), .A1(o_label6_data0[7]), .A2(o_label6_data1[7]), .A3(o_label6_data2[7]), .Z(n1472));
Q_MX02 U1846 ( .S(n4404), .A0(o_label7_data6[7]), .A1(o_label7_data7[7]), .Z(n1473));
Q_AN02 U1847 ( .A0(n4404), .A1(o_label7_data5[7]), .Z(n1474));
Q_MX02 U1848 ( .S(n4405), .A0(n1474), .A1(n1473), .Z(n1475));
Q_MX04 U1849 ( .S0(n4406), .S1(n4407), .A0(n1475), .A1(n1472), .A2(n1471), .A3(n1470), .Z(n1476));
Q_MX02 U1850 ( .S(n4408), .A0(n1476), .A1(n1469), .Z(r32_mux_5_data[7]));
Q_MX03 U1851 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[8]), .A1(o_label4_data6[8]), .A2(o_label4_data7[8]), .Z(n1477));
Q_MX04 U1852 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[8]), .A1(o_label4_data2[8]), .A2(o_label4_data3[8]), .A3(o_label4_data4[8]), .Z(n1478));
Q_MX02 U1853 ( .S(n4406), .A0(n1478), .A1(n1477), .Z(n1479));
Q_MX08 U1854 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[8]), .A1(o_label5_data3[8]), .A2(o_label5_data4[8]), .A3(o_label5_data5[8]), .A4(o_label5_data6[8]), .A5(o_label5_data7[8]), .A6(o_label5_config[8]), .A7(o_label4_data0[8]), .Z(n1480));
Q_MX02 U1855 ( .S(n4407), .A0(n1480), .A1(n1479), .Z(n1481));
Q_MX04 U1856 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[8]), .A1(o_label6_config[8]), .A2(o_label5_data0[8]), .A3(o_label5_data1[8]), .Z(n1482));
Q_MX04 U1857 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[8]), .A1(o_label6_data4[8]), .A2(o_label6_data5[8]), .A3(o_label6_data6[8]), .Z(n1483));
Q_MX04 U1858 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[8]), .A1(o_label6_data0[8]), .A2(o_label6_data1[8]), .A3(o_label6_data2[8]), .Z(n1484));
Q_MX02 U1859 ( .S(n4404), .A0(o_label7_data6[8]), .A1(o_label7_data7[8]), .Z(n1485));
Q_AN02 U1860 ( .A0(n4404), .A1(o_label7_data5[8]), .Z(n1486));
Q_MX02 U1861 ( .S(n4405), .A0(n1486), .A1(n1485), .Z(n1487));
Q_MX04 U1862 ( .S0(n4406), .S1(n4407), .A0(n1487), .A1(n1484), .A2(n1483), .A3(n1482), .Z(n1488));
Q_MX02 U1863 ( .S(n4408), .A0(n1488), .A1(n1481), .Z(r32_mux_5_data[8]));
Q_MX04 U1864 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[9]), .A1(o_label4_data5[9]), .A2(o_label4_data6[9]), .A3(o_label4_data7[9]), .Z(n1489));
Q_MX08 U1865 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[9]), .A1(o_label5_data5[9]), .A2(o_label5_data6[9]), .A3(o_label5_data7[9]), .A4(o_label4_data0[9]), .A5(o_label4_data1[9]), .A6(o_label4_data2[9]), .A7(o_label4_data3[9]), .Z(n1490));
Q_MX02 U1866 ( .S(n4412), .A0(n1490), .A1(n1489), .Z(n1491));
Q_MX04 U1867 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[9]), .A1(o_label5_data1[9]), .A2(o_label5_data2[9]), .A3(o_label5_data3[9]), .Z(n1492));
Q_MX04 U1868 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[9]), .A1(o_label6_data5[9]), .A2(o_label6_data6[9]), .A3(o_label6_data7[9]), .Z(n1493));
Q_MX04 U1869 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[9]), .A1(o_label6_data1[9]), .A2(o_label6_data2[9]), .A3(o_label6_data3[9]), .Z(n1494));
Q_MX02 U1870 ( .S(n4409), .A0(o_label7_data6[9]), .A1(o_label7_data7[9]), .Z(n1495));
Q_AN02 U1871 ( .A0(n4409), .A1(o_label7_data5[9]), .Z(n1496));
Q_MX02 U1872 ( .S(n4410), .A0(n1496), .A1(n1495), .Z(n1497));
Q_MX04 U1873 ( .S0(n4411), .S1(n4412), .A0(n1497), .A1(n1494), .A2(n1493), .A3(n1492), .Z(n1498));
Q_MX02 U1874 ( .S(n4413), .A0(n1498), .A1(n1491), .Z(r32_mux_5_data[9]));
Q_MX04 U1875 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[10]), .A1(o_label4_data5[10]), .A2(o_label4_data6[10]), .A3(o_label4_data7[10]), .Z(n1499));
Q_MX08 U1876 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[10]), .A1(o_label5_data5[10]), .A2(o_label5_data6[10]), .A3(o_label5_data7[10]), .A4(o_label4_data0[10]), .A5(o_label4_data1[10]), .A6(o_label4_data2[10]), .A7(o_label4_data3[10]), .Z(n1500));
Q_MX02 U1877 ( .S(n4412), .A0(n1500), .A1(n1499), .Z(n1501));
Q_MX04 U1878 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[10]), .A1(o_label5_data1[10]), .A2(o_label5_data2[10]), .A3(o_label5_data3[10]), .Z(n1502));
Q_MX04 U1879 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[10]), .A1(o_label6_data5[10]), .A2(o_label6_data6[10]), .A3(o_label6_data7[10]), .Z(n1503));
Q_MX04 U1880 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[10]), .A1(o_label6_data1[10]), .A2(o_label6_data2[10]), .A3(o_label6_data3[10]), .Z(n1504));
Q_MX02 U1881 ( .S(n4409), .A0(o_label7_data6[10]), .A1(o_label7_data7[10]), .Z(n1505));
Q_AN02 U1882 ( .A0(n4409), .A1(o_label7_data5[10]), .Z(n1506));
Q_MX02 U1883 ( .S(n4410), .A0(n1506), .A1(n1505), .Z(n1507));
Q_MX04 U1884 ( .S0(n4411), .S1(n4412), .A0(n1507), .A1(n1504), .A2(n1503), .A3(n1502), .Z(n1508));
Q_MX02 U1885 ( .S(n4413), .A0(n1508), .A1(n1501), .Z(r32_mux_5_data[10]));
Q_MX04 U1886 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[11]), .A1(o_label4_data5[11]), .A2(o_label4_data6[11]), .A3(o_label4_data7[11]), .Z(n1509));
Q_MX08 U1887 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[11]), .A1(o_label5_data5[11]), .A2(o_label5_data6[11]), .A3(o_label5_data7[11]), .A4(o_label4_data0[11]), .A5(o_label4_data1[11]), .A6(o_label4_data2[11]), .A7(o_label4_data3[11]), .Z(n1510));
Q_MX02 U1888 ( .S(n4412), .A0(n1510), .A1(n1509), .Z(n1511));
Q_MX04 U1889 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[11]), .A1(o_label5_data1[11]), .A2(o_label5_data2[11]), .A3(o_label5_data3[11]), .Z(n1512));
Q_MX04 U1890 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[11]), .A1(o_label6_data5[11]), .A2(o_label6_data6[11]), .A3(o_label6_data7[11]), .Z(n1513));
Q_MX04 U1891 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[11]), .A1(o_label6_data1[11]), .A2(o_label6_data2[11]), .A3(o_label6_data3[11]), .Z(n1514));
Q_MX02 U1892 ( .S(n4409), .A0(o_label7_data6[11]), .A1(o_label7_data7[11]), .Z(n1515));
Q_AN02 U1893 ( .A0(n4409), .A1(o_label7_data5[11]), .Z(n1516));
Q_MX02 U1894 ( .S(n4410), .A0(n1516), .A1(n1515), .Z(n1517));
Q_MX04 U1895 ( .S0(n4411), .S1(n4412), .A0(n1517), .A1(n1514), .A2(n1513), .A3(n1512), .Z(n1518));
Q_MX02 U1896 ( .S(n4413), .A0(n1518), .A1(n1511), .Z(r32_mux_5_data[11]));
Q_MX04 U1897 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[12]), .A1(o_label4_data5[12]), .A2(o_label4_data6[12]), .A3(o_label4_data7[12]), .Z(n1519));
Q_MX08 U1898 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[12]), .A1(o_label5_data5[12]), .A2(o_label5_data6[12]), .A3(o_label5_data7[12]), .A4(o_label4_data0[12]), .A5(o_label4_data1[12]), .A6(o_label4_data2[12]), .A7(o_label4_data3[12]), .Z(n1520));
Q_MX02 U1899 ( .S(n4412), .A0(n1520), .A1(n1519), .Z(n1521));
Q_MX04 U1900 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[12]), .A1(o_label5_data1[12]), .A2(o_label5_data2[12]), .A3(o_label5_data3[12]), .Z(n1522));
Q_MX04 U1901 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[12]), .A1(o_label6_data5[12]), .A2(o_label6_data6[12]), .A3(o_label6_data7[12]), .Z(n1523));
Q_MX04 U1902 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[12]), .A1(o_label6_data1[12]), .A2(o_label6_data2[12]), .A3(o_label6_data3[12]), .Z(n1524));
Q_MX02 U1903 ( .S(n4409), .A0(o_label7_data6[12]), .A1(o_label7_data7[12]), .Z(n1525));
Q_AN02 U1904 ( .A0(n4409), .A1(o_label7_data5[12]), .Z(n1526));
Q_MX02 U1905 ( .S(n4410), .A0(n1526), .A1(n1525), .Z(n1527));
Q_MX04 U1906 ( .S0(n4411), .S1(n4412), .A0(n1527), .A1(n1524), .A2(n1523), .A3(n1522), .Z(n1528));
Q_MX02 U1907 ( .S(n4413), .A0(n1528), .A1(n1521), .Z(r32_mux_5_data[12]));
Q_MX04 U1908 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[13]), .A1(o_label4_data5[13]), .A2(o_label4_data6[13]), .A3(o_label4_data7[13]), .Z(n1529));
Q_MX08 U1909 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[13]), .A1(o_label5_data5[13]), .A2(o_label5_data6[13]), .A3(o_label5_data7[13]), .A4(o_label4_data0[13]), .A5(o_label4_data1[13]), .A6(o_label4_data2[13]), .A7(o_label4_data3[13]), .Z(n1530));
Q_MX02 U1910 ( .S(n4412), .A0(n1530), .A1(n1529), .Z(n1531));
Q_MX04 U1911 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[13]), .A1(o_label5_data1[13]), .A2(o_label5_data2[13]), .A3(o_label5_data3[13]), .Z(n1532));
Q_MX04 U1912 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[13]), .A1(o_label6_data5[13]), .A2(o_label6_data6[13]), .A3(o_label6_data7[13]), .Z(n1533));
Q_MX04 U1913 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[13]), .A1(o_label6_data1[13]), .A2(o_label6_data2[13]), .A3(o_label6_data3[13]), .Z(n1534));
Q_MX02 U1914 ( .S(n4409), .A0(o_label7_data6[13]), .A1(o_label7_data7[13]), .Z(n1535));
Q_AN02 U1915 ( .A0(n4409), .A1(o_label7_data5[13]), .Z(n1536));
Q_MX02 U1916 ( .S(n4410), .A0(n1536), .A1(n1535), .Z(n1537));
Q_MX04 U1917 ( .S0(n4411), .S1(n4412), .A0(n1537), .A1(n1534), .A2(n1533), .A3(n1532), .Z(n1538));
Q_MX02 U1918 ( .S(n4413), .A0(n1538), .A1(n1531), .Z(r32_mux_5_data[13]));
Q_MX04 U1919 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[14]), .A1(o_label4_data5[14]), .A2(o_label4_data6[14]), .A3(o_label4_data7[14]), .Z(n1539));
Q_MX08 U1920 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[14]), .A1(o_label5_data5[14]), .A2(o_label5_data6[14]), .A3(o_label5_data7[14]), .A4(o_label4_data0[14]), .A5(o_label4_data1[14]), .A6(o_label4_data2[14]), .A7(o_label4_data3[14]), .Z(n1540));
Q_MX02 U1921 ( .S(n4412), .A0(n1540), .A1(n1539), .Z(n1541));
Q_MX04 U1922 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[14]), .A1(o_label5_data1[14]), .A2(o_label5_data2[14]), .A3(o_label5_data3[14]), .Z(n1542));
Q_MX04 U1923 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[14]), .A1(o_label6_data5[14]), .A2(o_label6_data6[14]), .A3(o_label6_data7[14]), .Z(n1543));
Q_MX04 U1924 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[14]), .A1(o_label6_data1[14]), .A2(o_label6_data2[14]), .A3(o_label6_data3[14]), .Z(n1544));
Q_MX02 U1925 ( .S(n4409), .A0(o_label7_data6[14]), .A1(o_label7_data7[14]), .Z(n1545));
Q_AN02 U1926 ( .A0(n4409), .A1(o_label7_data5[14]), .Z(n1546));
Q_MX02 U1927 ( .S(n4410), .A0(n1546), .A1(n1545), .Z(n1547));
Q_MX04 U1928 ( .S0(n4411), .S1(n4412), .A0(n1547), .A1(n1544), .A2(n1543), .A3(n1542), .Z(n1548));
Q_MX02 U1929 ( .S(n4413), .A0(n1548), .A1(n1541), .Z(r32_mux_5_data[14]));
Q_MX04 U1930 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[15]), .A1(o_label4_data5[15]), .A2(o_label4_data6[15]), .A3(o_label4_data7[15]), .Z(n1549));
Q_MX08 U1931 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[15]), .A1(o_label5_data5[15]), .A2(o_label5_data6[15]), .A3(o_label5_data7[15]), .A4(o_label4_data0[15]), .A5(o_label4_data1[15]), .A6(o_label4_data2[15]), .A7(o_label4_data3[15]), .Z(n1550));
Q_MX02 U1932 ( .S(n4412), .A0(n1550), .A1(n1549), .Z(n1551));
Q_MX04 U1933 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[15]), .A1(o_label5_data1[15]), .A2(o_label5_data2[15]), .A3(o_label5_data3[15]), .Z(n1552));
Q_MX04 U1934 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[15]), .A1(o_label6_data5[15]), .A2(o_label6_data6[15]), .A3(o_label6_data7[15]), .Z(n1553));
Q_MX04 U1935 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[15]), .A1(o_label6_data1[15]), .A2(o_label6_data2[15]), .A3(o_label6_data3[15]), .Z(n1554));
Q_MX02 U1936 ( .S(n4409), .A0(o_label7_data6[15]), .A1(o_label7_data7[15]), .Z(n1555));
Q_AN02 U1937 ( .A0(n4409), .A1(o_label7_data5[15]), .Z(n1556));
Q_MX02 U1938 ( .S(n4410), .A0(n1556), .A1(n1555), .Z(n1557));
Q_MX04 U1939 ( .S0(n4411), .S1(n4412), .A0(n1557), .A1(n1554), .A2(n1553), .A3(n1552), .Z(n1558));
Q_MX02 U1940 ( .S(n4413), .A0(n1558), .A1(n1551), .Z(r32_mux_5_data[15]));
Q_MX04 U1941 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[16]), .A1(o_label4_data5[16]), .A2(o_label4_data6[16]), .A3(o_label4_data7[16]), .Z(n1559));
Q_MX08 U1942 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[16]), .A1(o_label5_data5[16]), .A2(o_label5_data6[16]), .A3(o_label5_data7[16]), .A4(o_label4_data0[16]), .A5(o_label4_data1[16]), .A6(o_label4_data2[16]), .A7(o_label4_data3[16]), .Z(n1560));
Q_MX02 U1943 ( .S(n4412), .A0(n1560), .A1(n1559), .Z(n1561));
Q_MX04 U1944 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[16]), .A1(o_label5_data1[16]), .A2(o_label5_data2[16]), .A3(o_label5_data3[16]), .Z(n1562));
Q_MX04 U1945 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[16]), .A1(o_label6_data5[16]), .A2(o_label6_data6[16]), .A3(o_label6_data7[16]), .Z(n1563));
Q_MX04 U1946 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[16]), .A1(o_label6_data1[16]), .A2(o_label6_data2[16]), .A3(o_label6_data3[16]), .Z(n1564));
Q_MX02 U1947 ( .S(n4409), .A0(o_label7_data6[16]), .A1(o_label7_data7[16]), .Z(n1565));
Q_AN02 U1948 ( .A0(n4409), .A1(o_label7_data5[16]), .Z(n1566));
Q_MX02 U1949 ( .S(n4410), .A0(n1566), .A1(n1565), .Z(n1567));
Q_MX04 U1950 ( .S0(n4411), .S1(n4412), .A0(n1567), .A1(n1564), .A2(n1563), .A3(n1562), .Z(n1568));
Q_MX02 U1951 ( .S(n4413), .A0(n1568), .A1(n1561), .Z(r32_mux_5_data[16]));
Q_MX04 U1952 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[17]), .A1(o_label4_data5[17]), .A2(o_label4_data6[17]), .A3(o_label4_data7[17]), .Z(n1569));
Q_MX08 U1953 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[17]), .A1(o_label5_data5[17]), .A2(o_label5_data6[17]), .A3(o_label5_data7[17]), .A4(o_label4_data0[17]), .A5(o_label4_data1[17]), .A6(o_label4_data2[17]), .A7(o_label4_data3[17]), .Z(n1570));
Q_MX02 U1954 ( .S(n4412), .A0(n1570), .A1(n1569), .Z(n1571));
Q_MX04 U1955 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[17]), .A1(o_label5_data1[17]), .A2(o_label5_data2[17]), .A3(o_label5_data3[17]), .Z(n1572));
Q_MX04 U1956 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[17]), .A1(o_label6_data5[17]), .A2(o_label6_data6[17]), .A3(o_label6_data7[17]), .Z(n1573));
Q_MX04 U1957 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[17]), .A1(o_label6_data1[17]), .A2(o_label6_data2[17]), .A3(o_label6_data3[17]), .Z(n1574));
Q_MX02 U1958 ( .S(n4409), .A0(o_label7_data6[17]), .A1(o_label7_data7[17]), .Z(n1575));
Q_AN02 U1959 ( .A0(n4409), .A1(o_label7_data5[17]), .Z(n1576));
Q_MX02 U1960 ( .S(n4410), .A0(n1576), .A1(n1575), .Z(n1577));
Q_MX04 U1961 ( .S0(n4411), .S1(n4412), .A0(n1577), .A1(n1574), .A2(n1573), .A3(n1572), .Z(n1578));
Q_MX02 U1962 ( .S(n4413), .A0(n1578), .A1(n1571), .Z(r32_mux_5_data[17]));
Q_MX04 U1963 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[18]), .A1(o_label4_data5[18]), .A2(o_label4_data6[18]), .A3(o_label4_data7[18]), .Z(n1579));
Q_MX08 U1964 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[18]), .A1(o_label5_data5[18]), .A2(o_label5_data6[18]), .A3(o_label5_data7[18]), .A4(o_label4_data0[18]), .A5(o_label4_data1[18]), .A6(o_label4_data2[18]), .A7(o_label4_data3[18]), .Z(n1580));
Q_MX02 U1965 ( .S(n4412), .A0(n1580), .A1(n1579), .Z(n1581));
Q_MX04 U1966 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[18]), .A1(o_label5_data1[18]), .A2(o_label5_data2[18]), .A3(o_label5_data3[18]), .Z(n1582));
Q_MX04 U1967 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[18]), .A1(o_label6_data5[18]), .A2(o_label6_data6[18]), .A3(o_label6_data7[18]), .Z(n1583));
Q_MX04 U1968 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[18]), .A1(o_label6_data1[18]), .A2(o_label6_data2[18]), .A3(o_label6_data3[18]), .Z(n1584));
Q_MX02 U1969 ( .S(n4409), .A0(o_label7_data6[18]), .A1(o_label7_data7[18]), .Z(n1585));
Q_AN02 U1970 ( .A0(n4409), .A1(o_label7_data5[18]), .Z(n1586));
Q_MX02 U1971 ( .S(n4410), .A0(n1586), .A1(n1585), .Z(n1587));
Q_MX04 U1972 ( .S0(n4411), .S1(n4412), .A0(n1587), .A1(n1584), .A2(n1583), .A3(n1582), .Z(n1588));
Q_MX02 U1973 ( .S(n4413), .A0(n1588), .A1(n1581), .Z(r32_mux_5_data[18]));
Q_MX04 U1974 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[19]), .A1(o_label4_data5[19]), .A2(o_label4_data6[19]), .A3(o_label4_data7[19]), .Z(n1589));
Q_MX08 U1975 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[19]), .A1(o_label5_data5[19]), .A2(o_label5_data6[19]), .A3(o_label5_data7[19]), .A4(o_label4_data0[19]), .A5(o_label4_data1[19]), .A6(o_label4_data2[19]), .A7(o_label4_data3[19]), .Z(n1590));
Q_MX02 U1976 ( .S(n4412), .A0(n1590), .A1(n1589), .Z(n1591));
Q_MX04 U1977 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[19]), .A1(o_label5_data1[19]), .A2(o_label5_data2[19]), .A3(o_label5_data3[19]), .Z(n1592));
Q_MX04 U1978 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[19]), .A1(o_label6_data5[19]), .A2(o_label6_data6[19]), .A3(o_label6_data7[19]), .Z(n1593));
Q_MX04 U1979 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[19]), .A1(o_label6_data1[19]), .A2(o_label6_data2[19]), .A3(o_label6_data3[19]), .Z(n1594));
Q_MX02 U1980 ( .S(n4409), .A0(o_label7_data6[19]), .A1(o_label7_data7[19]), .Z(n1595));
Q_AN02 U1981 ( .A0(n4409), .A1(o_label7_data5[19]), .Z(n1596));
Q_MX02 U1982 ( .S(n4410), .A0(n1596), .A1(n1595), .Z(n1597));
Q_MX04 U1983 ( .S0(n4411), .S1(n4412), .A0(n1597), .A1(n1594), .A2(n1593), .A3(n1592), .Z(n1598));
Q_MX02 U1984 ( .S(n4413), .A0(n1598), .A1(n1591), .Z(r32_mux_5_data[19]));
Q_MX04 U1985 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[20]), .A1(o_label4_data5[20]), .A2(o_label4_data6[20]), .A3(o_label4_data7[20]), .Z(n1599));
Q_MX08 U1986 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[20]), .A1(o_label5_data5[20]), .A2(o_label5_data6[20]), .A3(o_label5_data7[20]), .A4(o_label4_data0[20]), .A5(o_label4_data1[20]), .A6(o_label4_data2[20]), .A7(o_label4_data3[20]), .Z(n1600));
Q_MX02 U1987 ( .S(n4412), .A0(n1600), .A1(n1599), .Z(n1601));
Q_MX04 U1988 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[20]), .A1(o_label5_data1[20]), .A2(o_label5_data2[20]), .A3(o_label5_data3[20]), .Z(n1602));
Q_MX04 U1989 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[20]), .A1(o_label6_data5[20]), .A2(o_label6_data6[20]), .A3(o_label6_data7[20]), .Z(n1603));
Q_MX04 U1990 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[20]), .A1(o_label6_data1[20]), .A2(o_label6_data2[20]), .A3(o_label6_data3[20]), .Z(n1604));
Q_MX02 U1991 ( .S(n4409), .A0(o_label7_data6[20]), .A1(o_label7_data7[20]), .Z(n1605));
Q_AN02 U1992 ( .A0(n4409), .A1(o_label7_data5[20]), .Z(n1606));
Q_MX02 U1993 ( .S(n4410), .A0(n1606), .A1(n1605), .Z(n1607));
Q_MX04 U1994 ( .S0(n4411), .S1(n4412), .A0(n1607), .A1(n1604), .A2(n1603), .A3(n1602), .Z(n1608));
Q_MX02 U1995 ( .S(n4413), .A0(n1608), .A1(n1601), .Z(r32_mux_5_data[20]));
Q_MX04 U1996 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[21]), .A1(o_label4_data5[21]), .A2(o_label4_data6[21]), .A3(o_label4_data7[21]), .Z(n1609));
Q_MX08 U1997 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[21]), .A1(o_label5_data5[21]), .A2(o_label5_data6[21]), .A3(o_label5_data7[21]), .A4(o_label4_data0[21]), .A5(o_label4_data1[21]), .A6(o_label4_data2[21]), .A7(o_label4_data3[21]), .Z(n1610));
Q_MX02 U1998 ( .S(n4412), .A0(n1610), .A1(n1609), .Z(n1611));
Q_MX04 U1999 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[21]), .A1(o_label5_data1[21]), .A2(o_label5_data2[21]), .A3(o_label5_data3[21]), .Z(n1612));
Q_MX04 U2000 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[21]), .A1(o_label6_data5[21]), .A2(o_label6_data6[21]), .A3(o_label6_data7[21]), .Z(n1613));
Q_MX04 U2001 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[21]), .A1(o_label6_data1[21]), .A2(o_label6_data2[21]), .A3(o_label6_data3[21]), .Z(n1614));
Q_MX02 U2002 ( .S(n4409), .A0(o_label7_data6[21]), .A1(o_label7_data7[21]), .Z(n1615));
Q_AN02 U2003 ( .A0(n4409), .A1(o_label7_data5[21]), .Z(n1616));
Q_MX02 U2004 ( .S(n4410), .A0(n1616), .A1(n1615), .Z(n1617));
Q_MX04 U2005 ( .S0(n4411), .S1(n4412), .A0(n1617), .A1(n1614), .A2(n1613), .A3(n1612), .Z(n1618));
Q_MX02 U2006 ( .S(n4413), .A0(n1618), .A1(n1611), .Z(r32_mux_5_data[21]));
Q_MX04 U2007 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[22]), .A1(o_label4_data5[22]), .A2(o_label4_data6[22]), .A3(o_label4_data7[22]), .Z(n1619));
Q_MX08 U2008 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[22]), .A1(o_label5_data5[22]), .A2(o_label5_data6[22]), .A3(o_label5_data7[22]), .A4(o_label4_data0[22]), .A5(o_label4_data1[22]), .A6(o_label4_data2[22]), .A7(o_label4_data3[22]), .Z(n1620));
Q_MX02 U2009 ( .S(n4412), .A0(n1620), .A1(n1619), .Z(n1621));
Q_MX04 U2010 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[22]), .A1(o_label5_data1[22]), .A2(o_label5_data2[22]), .A3(o_label5_data3[22]), .Z(n1622));
Q_MX04 U2011 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[22]), .A1(o_label6_data5[22]), .A2(o_label6_data6[22]), .A3(o_label6_data7[22]), .Z(n1623));
Q_MX04 U2012 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[22]), .A1(o_label6_data1[22]), .A2(o_label6_data2[22]), .A3(o_label6_data3[22]), .Z(n1624));
Q_MX02 U2013 ( .S(n4409), .A0(o_label7_data6[22]), .A1(o_label7_data7[22]), .Z(n1625));
Q_AN02 U2014 ( .A0(n4409), .A1(o_label7_data5[22]), .Z(n1626));
Q_MX02 U2015 ( .S(n4410), .A0(n1626), .A1(n1625), .Z(n1627));
Q_MX04 U2016 ( .S0(n4411), .S1(n4412), .A0(n1627), .A1(n1624), .A2(n1623), .A3(n1622), .Z(n1628));
Q_MX02 U2017 ( .S(n4413), .A0(n1628), .A1(n1621), .Z(r32_mux_5_data[22]));
Q_MX04 U2018 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[23]), .A1(o_label4_data5[23]), .A2(o_label4_data6[23]), .A3(o_label4_data7[23]), .Z(n1629));
Q_MX08 U2019 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[23]), .A1(o_label5_data5[23]), .A2(o_label5_data6[23]), .A3(o_label5_data7[23]), .A4(o_label4_data0[23]), .A5(o_label4_data1[23]), .A6(o_label4_data2[23]), .A7(o_label4_data3[23]), .Z(n1630));
Q_MX02 U2020 ( .S(n4412), .A0(n1630), .A1(n1629), .Z(n1631));
Q_MX04 U2021 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[23]), .A1(o_label5_data1[23]), .A2(o_label5_data2[23]), .A3(o_label5_data3[23]), .Z(n1632));
Q_MX04 U2022 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[23]), .A1(o_label6_data5[23]), .A2(o_label6_data6[23]), .A3(o_label6_data7[23]), .Z(n1633));
Q_MX04 U2023 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[23]), .A1(o_label6_data1[23]), .A2(o_label6_data2[23]), .A3(o_label6_data3[23]), .Z(n1634));
Q_MX02 U2024 ( .S(n4409), .A0(o_label7_data6[23]), .A1(o_label7_data7[23]), .Z(n1635));
Q_AN02 U2025 ( .A0(n4409), .A1(o_label7_data5[23]), .Z(n1636));
Q_MX02 U2026 ( .S(n4410), .A0(n1636), .A1(n1635), .Z(n1637));
Q_MX04 U2027 ( .S0(n4411), .S1(n4412), .A0(n1637), .A1(n1634), .A2(n1633), .A3(n1632), .Z(n1638));
Q_MX02 U2028 ( .S(n4413), .A0(n1638), .A1(n1631), .Z(r32_mux_5_data[23]));
Q_MX04 U2029 ( .S0(n4409), .S1(n4410), .A0(o_label4_data4[24]), .A1(o_label4_data5[24]), .A2(o_label4_data6[24]), .A3(o_label4_data7[24]), .Z(n1639));
Q_MX08 U2030 ( .S0(n4409), .S1(n4410), .S2(n4411), .A0(o_label5_data4[24]), .A1(o_label5_data5[24]), .A2(o_label5_data6[24]), .A3(o_label5_data7[24]), .A4(o_label4_data0[24]), .A5(o_label4_data1[24]), .A6(o_label4_data2[24]), .A7(o_label4_data3[24]), .Z(n1640));
Q_MX02 U2031 ( .S(n4412), .A0(n1640), .A1(n1639), .Z(n1641));
Q_MX04 U2032 ( .S0(n4409), .S1(n4410), .A0(o_label5_data0[24]), .A1(o_label5_data1[24]), .A2(o_label5_data2[24]), .A3(o_label5_data3[24]), .Z(n1642));
Q_MX04 U2033 ( .S0(n4409), .S1(n4410), .A0(o_label6_data4[24]), .A1(o_label6_data5[24]), .A2(o_label6_data6[24]), .A3(o_label6_data7[24]), .Z(n1643));
Q_MX04 U2034 ( .S0(n4409), .S1(n4410), .A0(o_label6_data0[24]), .A1(o_label6_data1[24]), .A2(o_label6_data2[24]), .A3(o_label6_data3[24]), .Z(n1644));
Q_MX02 U2035 ( .S(n4409), .A0(o_label7_data6[24]), .A1(o_label7_data7[24]), .Z(n1645));
Q_AN02 U2036 ( .A0(n4409), .A1(o_label7_data5[24]), .Z(n1646));
Q_MX02 U2037 ( .S(n4410), .A0(n1646), .A1(n1645), .Z(n1647));
Q_MX04 U2038 ( .S0(n4411), .S1(n4412), .A0(n1647), .A1(n1644), .A2(n1643), .A3(n1642), .Z(n1648));
Q_MX02 U2039 ( .S(n4413), .A0(n1648), .A1(n1641), .Z(r32_mux_5_data[24]));
Q_MX03 U2040 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[25]), .A1(o_label4_data6[25]), .A2(o_label4_data7[25]), .Z(n1649));
Q_MX04 U2041 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[25]), .A1(o_label4_data2[25]), .A2(o_label4_data3[25]), .A3(o_label4_data4[25]), .Z(n1650));
Q_MX02 U2042 ( .S(n4406), .A0(n1650), .A1(n1649), .Z(n1651));
Q_MX08 U2043 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[25]), .A1(o_label5_data3[25]), .A2(o_label5_data4[25]), .A3(o_label5_data5[25]), .A4(o_label5_data6[25]), .A5(o_label5_data7[25]), .A6(o_label5_config[9]), .A7(o_label4_data0[25]), .Z(n1652));
Q_MX02 U2044 ( .S(n4407), .A0(n1652), .A1(n1651), .Z(n1653));
Q_MX04 U2045 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[25]), .A1(o_label6_config[9]), .A2(o_label5_data0[25]), .A3(o_label5_data1[25]), .Z(n1654));
Q_MX04 U2046 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[25]), .A1(o_label6_data4[25]), .A2(o_label6_data5[25]), .A3(o_label6_data6[25]), .Z(n1655));
Q_MX04 U2047 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[9]), .A1(o_label6_data0[25]), .A2(o_label6_data1[25]), .A3(o_label6_data2[25]), .Z(n1656));
Q_MX02 U2048 ( .S(n4404), .A0(o_label7_data6[25]), .A1(o_label7_data7[25]), .Z(n1657));
Q_AN02 U2049 ( .A0(n4404), .A1(o_label7_data5[25]), .Z(n1658));
Q_MX02 U2050 ( .S(n4405), .A0(n1658), .A1(n1657), .Z(n1659));
Q_MX04 U2051 ( .S0(n4406), .S1(n4407), .A0(n1659), .A1(n1656), .A2(n1655), .A3(n1654), .Z(n1660));
Q_MX02 U2052 ( .S(n4408), .A0(n1660), .A1(n1653), .Z(r32_mux_5_data[25]));
Q_MX03 U2053 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[26]), .A1(o_label4_data6[26]), .A2(o_label4_data7[26]), .Z(n1661));
Q_MX04 U2054 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[26]), .A1(o_label4_data2[26]), .A2(o_label4_data3[26]), .A3(o_label4_data4[26]), .Z(n1662));
Q_MX02 U2055 ( .S(n4406), .A0(n1662), .A1(n1661), .Z(n1663));
Q_MX08 U2056 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[26]), .A1(o_label5_data3[26]), .A2(o_label5_data4[26]), .A3(o_label5_data5[26]), .A4(o_label5_data6[26]), .A5(o_label5_data7[26]), .A6(o_label5_config[10]), .A7(o_label4_data0[26]), .Z(n1664));
Q_MX02 U2057 ( .S(n4407), .A0(n1664), .A1(n1663), .Z(n1665));
Q_MX04 U2058 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[26]), .A1(o_label6_config[10]), .A2(o_label5_data0[26]), .A3(o_label5_data1[26]), .Z(n1666));
Q_MX04 U2059 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[26]), .A1(o_label6_data4[26]), .A2(o_label6_data5[26]), .A3(o_label6_data6[26]), .Z(n1667));
Q_MX04 U2060 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[10]), .A1(o_label6_data0[26]), .A2(o_label6_data1[26]), .A3(o_label6_data2[26]), .Z(n1668));
Q_MX02 U2061 ( .S(n4404), .A0(o_label7_data6[26]), .A1(o_label7_data7[26]), .Z(n1669));
Q_AN02 U2062 ( .A0(n4404), .A1(o_label7_data5[26]), .Z(n1670));
Q_MX02 U2063 ( .S(n4405), .A0(n1670), .A1(n1669), .Z(n1671));
Q_MX04 U2064 ( .S0(n4406), .S1(n4407), .A0(n1671), .A1(n1668), .A2(n1667), .A3(n1666), .Z(n1672));
Q_MX02 U2065 ( .S(n4408), .A0(n1672), .A1(n1665), .Z(r32_mux_5_data[26]));
Q_MX03 U2066 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[27]), .A1(o_label4_data6[27]), .A2(o_label4_data7[27]), .Z(n1673));
Q_MX04 U2067 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[27]), .A1(o_label4_data2[27]), .A2(o_label4_data3[27]), .A3(o_label4_data4[27]), .Z(n1674));
Q_MX02 U2068 ( .S(n4406), .A0(n1674), .A1(n1673), .Z(n1675));
Q_MX08 U2069 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[27]), .A1(o_label5_data3[27]), .A2(o_label5_data4[27]), .A3(o_label5_data5[27]), .A4(o_label5_data6[27]), .A5(o_label5_data7[27]), .A6(o_label5_config[11]), .A7(o_label4_data0[27]), .Z(n1676));
Q_MX02 U2070 ( .S(n4407), .A0(n1676), .A1(n1675), .Z(n1677));
Q_MX04 U2071 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[27]), .A1(o_label6_config[11]), .A2(o_label5_data0[27]), .A3(o_label5_data1[27]), .Z(n1678));
Q_MX04 U2072 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[27]), .A1(o_label6_data4[27]), .A2(o_label6_data5[27]), .A3(o_label6_data6[27]), .Z(n1679));
Q_MX04 U2073 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[11]), .A1(o_label6_data0[27]), .A2(o_label6_data1[27]), .A3(o_label6_data2[27]), .Z(n1680));
Q_MX02 U2074 ( .S(n4404), .A0(o_label7_data6[27]), .A1(o_label7_data7[27]), .Z(n1681));
Q_AN02 U2075 ( .A0(n4404), .A1(o_label7_data5[27]), .Z(n1682));
Q_MX02 U2076 ( .S(n4405), .A0(n1682), .A1(n1681), .Z(n1683));
Q_MX04 U2077 ( .S0(n4406), .S1(n4407), .A0(n1683), .A1(n1680), .A2(n1679), .A3(n1678), .Z(n1684));
Q_MX02 U2078 ( .S(n4408), .A0(n1684), .A1(n1677), .Z(r32_mux_5_data[27]));
Q_MX03 U2079 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[28]), .A1(o_label4_data6[28]), .A2(o_label4_data7[28]), .Z(n1685));
Q_MX04 U2080 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[28]), .A1(o_label4_data2[28]), .A2(o_label4_data3[28]), .A3(o_label4_data4[28]), .Z(n1686));
Q_MX02 U2081 ( .S(n4406), .A0(n1686), .A1(n1685), .Z(n1687));
Q_MX08 U2082 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[28]), .A1(o_label5_data3[28]), .A2(o_label5_data4[28]), .A3(o_label5_data5[28]), .A4(o_label5_data6[28]), .A5(o_label5_data7[28]), .A6(o_label5_config[12]), .A7(o_label4_data0[28]), .Z(n1688));
Q_MX02 U2083 ( .S(n4407), .A0(n1688), .A1(n1687), .Z(n1689));
Q_MX04 U2084 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[28]), .A1(o_label6_config[12]), .A2(o_label5_data0[28]), .A3(o_label5_data1[28]), .Z(n1690));
Q_MX04 U2085 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[28]), .A1(o_label6_data4[28]), .A2(o_label6_data5[28]), .A3(o_label6_data6[28]), .Z(n1691));
Q_MX04 U2086 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[12]), .A1(o_label6_data0[28]), .A2(o_label6_data1[28]), .A3(o_label6_data2[28]), .Z(n1692));
Q_MX02 U2087 ( .S(n4404), .A0(o_label7_data6[28]), .A1(o_label7_data7[28]), .Z(n1693));
Q_AN02 U2088 ( .A0(n4404), .A1(o_label7_data5[28]), .Z(n1694));
Q_MX02 U2089 ( .S(n4405), .A0(n1694), .A1(n1693), .Z(n1695));
Q_MX04 U2090 ( .S0(n4406), .S1(n4407), .A0(n1695), .A1(n1692), .A2(n1691), .A3(n1690), .Z(n1696));
Q_MX02 U2091 ( .S(n4408), .A0(n1696), .A1(n1689), .Z(r32_mux_5_data[28]));
Q_MX03 U2092 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[29]), .A1(o_label4_data6[29]), .A2(o_label4_data7[29]), .Z(n1697));
Q_MX04 U2093 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[29]), .A1(o_label4_data2[29]), .A2(o_label4_data3[29]), .A3(o_label4_data4[29]), .Z(n1698));
Q_MX02 U2094 ( .S(n4406), .A0(n1698), .A1(n1697), .Z(n1699));
Q_MX08 U2095 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[29]), .A1(o_label5_data3[29]), .A2(o_label5_data4[29]), .A3(o_label5_data5[29]), .A4(o_label5_data6[29]), .A5(o_label5_data7[29]), .A6(o_label5_config[13]), .A7(o_label4_data0[29]), .Z(n1700));
Q_MX02 U2096 ( .S(n4407), .A0(n1700), .A1(n1699), .Z(n1701));
Q_MX04 U2097 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[29]), .A1(o_label6_config[13]), .A2(o_label5_data0[29]), .A3(o_label5_data1[29]), .Z(n1702));
Q_MX04 U2098 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[29]), .A1(o_label6_data4[29]), .A2(o_label6_data5[29]), .A3(o_label6_data6[29]), .Z(n1703));
Q_MX04 U2099 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[13]), .A1(o_label6_data0[29]), .A2(o_label6_data1[29]), .A3(o_label6_data2[29]), .Z(n1704));
Q_MX02 U2100 ( .S(n4404), .A0(o_label7_data6[29]), .A1(o_label7_data7[29]), .Z(n1705));
Q_AN02 U2101 ( .A0(n4404), .A1(o_label7_data5[29]), .Z(n1706));
Q_MX02 U2102 ( .S(n4405), .A0(n1706), .A1(n1705), .Z(n1707));
Q_MX04 U2103 ( .S0(n4406), .S1(n4407), .A0(n1707), .A1(n1704), .A2(n1703), .A3(n1702), .Z(n1708));
Q_MX02 U2104 ( .S(n4408), .A0(n1708), .A1(n1701), .Z(r32_mux_5_data[29]));
Q_MX03 U2105 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[30]), .A1(o_label4_data6[30]), .A2(o_label4_data7[30]), .Z(n1709));
Q_MX04 U2106 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[30]), .A1(o_label4_data2[30]), .A2(o_label4_data3[30]), .A3(o_label4_data4[30]), .Z(n1710));
Q_MX02 U2107 ( .S(n4406), .A0(n1710), .A1(n1709), .Z(n1711));
Q_MX08 U2108 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[30]), .A1(o_label5_data3[30]), .A2(o_label5_data4[30]), .A3(o_label5_data5[30]), .A4(o_label5_data6[30]), .A5(o_label5_data7[30]), .A6(o_label5_config[14]), .A7(o_label4_data0[30]), .Z(n1712));
Q_MX02 U2109 ( .S(n4407), .A0(n1712), .A1(n1711), .Z(n1713));
Q_MX04 U2110 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[30]), .A1(o_label6_config[14]), .A2(o_label5_data0[30]), .A3(o_label5_data1[30]), .Z(n1714));
Q_MX04 U2111 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[30]), .A1(o_label6_data4[30]), .A2(o_label6_data5[30]), .A3(o_label6_data6[30]), .Z(n1715));
Q_MX04 U2112 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[14]), .A1(o_label6_data0[30]), .A2(o_label6_data1[30]), .A3(o_label6_data2[30]), .Z(n1716));
Q_MX02 U2113 ( .S(n4404), .A0(o_label7_data6[30]), .A1(o_label7_data7[30]), .Z(n1717));
Q_AN02 U2114 ( .A0(n4404), .A1(o_label7_data5[30]), .Z(n1718));
Q_MX02 U2115 ( .S(n4405), .A0(n1718), .A1(n1717), .Z(n1719));
Q_MX04 U2116 ( .S0(n4406), .S1(n4407), .A0(n1719), .A1(n1716), .A2(n1715), .A3(n1714), .Z(n1720));
Q_MX02 U2117 ( .S(n4408), .A0(n1720), .A1(n1713), .Z(r32_mux_5_data[30]));
Q_MX03 U2118 ( .S0(n4404), .S1(n4405), .A0(o_label4_data5[31]), .A1(o_label4_data6[31]), .A2(o_label4_data7[31]), .Z(n1721));
Q_MX04 U2119 ( .S0(n4404), .S1(n4405), .A0(o_label4_data1[31]), .A1(o_label4_data2[31]), .A2(o_label4_data3[31]), .A3(o_label4_data4[31]), .Z(n1722));
Q_MX02 U2120 ( .S(n4406), .A0(n1722), .A1(n1721), .Z(n1723));
Q_MX08 U2121 ( .S0(n4404), .S1(n4405), .S2(n4406), .A0(o_label5_data2[31]), .A1(o_label5_data3[31]), .A2(o_label5_data4[31]), .A3(o_label5_data5[31]), .A4(o_label5_data6[31]), .A5(o_label5_data7[31]), .A6(o_label5_config[15]), .A7(o_label4_data0[31]), .Z(n1724));
Q_MX02 U2122 ( .S(n4407), .A0(n1724), .A1(n1723), .Z(n1725));
Q_MX04 U2123 ( .S0(n4404), .S1(n4405), .A0(o_label6_data7[31]), .A1(o_label6_config[15]), .A2(o_label5_data0[31]), .A3(o_label5_data1[31]), .Z(n1726));
Q_MX04 U2124 ( .S0(n4404), .S1(n4405), .A0(o_label6_data3[31]), .A1(o_label6_data4[31]), .A2(o_label6_data5[31]), .A3(o_label6_data6[31]), .Z(n1727));
Q_MX04 U2125 ( .S0(n4404), .S1(n4405), .A0(o_label7_config[15]), .A1(o_label6_data0[31]), .A2(o_label6_data1[31]), .A3(o_label6_data2[31]), .Z(n1728));
Q_MX02 U2126 ( .S(n4404), .A0(o_label7_data6[31]), .A1(o_label7_data7[31]), .Z(n1729));
Q_AN02 U2127 ( .A0(n4404), .A1(o_label7_data5[31]), .Z(n1730));
Q_MX02 U2128 ( .S(n4405), .A0(n1730), .A1(n1729), .Z(n1731));
Q_MX04 U2129 ( .S0(n4406), .S1(n4407), .A0(n1731), .A1(n1728), .A2(n1727), .A3(n1726), .Z(n1732));
Q_MX02 U2130 ( .S(n4408), .A0(n1732), .A1(n1725), .Z(r32_mux_5_data[31]));
Q_MX03 U2131 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[0]), .A1(o_label0_data0[0]), .A2(o_label0_data1[0]), .Z(n1733));
Q_MX04 U2132 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[0]), .A1(o_label1_data5[0]), .A2(o_label1_data6[0]), .A3(o_label1_data7[0]), .Z(n1734));
Q_MX02 U2133 ( .S(n4416), .A0(n1734), .A1(n1733), .Z(n1735));
Q_MX08 U2134 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[0]), .A1(o_label2_data6[0]), .A2(o_label2_data7[0]), .A3(o_label2_config[0]), .A4(o_label1_data0[0]), .A5(o_label1_data1[0]), .A6(o_label1_data2[0]), .A7(o_label1_data3[0]), .Z(n1736));
Q_MX02 U2135 ( .S(n4417), .A0(n1736), .A1(n1735), .Z(n1737));
Q_MX04 U2136 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[0]), .A1(o_label2_data2[0]), .A2(o_label2_data3[0]), .A3(o_label2_data4[0]), .Z(n1738));
Q_MX04 U2137 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[0]), .A1(o_label3_data7[0]), .A2(o_label3_config[0]), .A3(o_label2_data0[0]), .Z(n1739));
Q_MX04 U2138 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[0]), .A1(o_label3_data3[0]), .A2(o_label3_data4[0]), .A3(o_label3_data5[0]), .Z(n1740));
Q_MX02 U2139 ( .S(n4414), .A0(o_label3_data0[0]), .A1(o_label3_data1[0]), .Z(n1741));
Q_AN02 U2140 ( .A0(n4414), .A1(o_label4_config[0]), .Z(n1742));
Q_MX02 U2141 ( .S(n4415), .A0(n1742), .A1(n1741), .Z(n1743));
Q_MX04 U2142 ( .S0(n4416), .S1(n4417), .A0(n1743), .A1(n1740), .A2(n1739), .A3(n1738), .Z(n1744));
Q_MX02 U2143 ( .S(n4418), .A0(n1744), .A1(n1737), .Z(r32_mux_4_data[0]));
Q_MX03 U2144 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[1]), .A1(o_label0_data0[1]), .A2(o_label0_data1[1]), .Z(n1745));
Q_MX04 U2145 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[1]), .A1(o_label1_data5[1]), .A2(o_label1_data6[1]), .A3(o_label1_data7[1]), .Z(n1746));
Q_MX02 U2146 ( .S(n4416), .A0(n1746), .A1(n1745), .Z(n1747));
Q_MX08 U2147 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[1]), .A1(o_label2_data6[1]), .A2(o_label2_data7[1]), .A3(o_label2_config[1]), .A4(o_label1_data0[1]), .A5(o_label1_data1[1]), .A6(o_label1_data2[1]), .A7(o_label1_data3[1]), .Z(n1748));
Q_MX02 U2148 ( .S(n4417), .A0(n1748), .A1(n1747), .Z(n1749));
Q_MX04 U2149 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[1]), .A1(o_label2_data2[1]), .A2(o_label2_data3[1]), .A3(o_label2_data4[1]), .Z(n1750));
Q_MX04 U2150 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[1]), .A1(o_label3_data7[1]), .A2(o_label3_config[1]), .A3(o_label2_data0[1]), .Z(n1751));
Q_MX04 U2151 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[1]), .A1(o_label3_data3[1]), .A2(o_label3_data4[1]), .A3(o_label3_data5[1]), .Z(n1752));
Q_MX02 U2152 ( .S(n4414), .A0(o_label3_data0[1]), .A1(o_label3_data1[1]), .Z(n1753));
Q_AN02 U2153 ( .A0(n4414), .A1(o_label4_config[1]), .Z(n1754));
Q_MX02 U2154 ( .S(n4415), .A0(n1754), .A1(n1753), .Z(n1755));
Q_MX04 U2155 ( .S0(n4416), .S1(n4417), .A0(n1755), .A1(n1752), .A2(n1751), .A3(n1750), .Z(n1756));
Q_MX02 U2156 ( .S(n4418), .A0(n1756), .A1(n1749), .Z(r32_mux_4_data[1]));
Q_MX03 U2157 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[2]), .A1(o_label0_data0[2]), .A2(o_label0_data1[2]), .Z(n1757));
Q_MX04 U2158 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[2]), .A1(o_label1_data5[2]), .A2(o_label1_data6[2]), .A3(o_label1_data7[2]), .Z(n1758));
Q_MX02 U2159 ( .S(n4416), .A0(n1758), .A1(n1757), .Z(n1759));
Q_MX08 U2160 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[2]), .A1(o_label2_data6[2]), .A2(o_label2_data7[2]), .A3(o_label2_config[2]), .A4(o_label1_data0[2]), .A5(o_label1_data1[2]), .A6(o_label1_data2[2]), .A7(o_label1_data3[2]), .Z(n1760));
Q_MX02 U2161 ( .S(n4417), .A0(n1760), .A1(n1759), .Z(n1761));
Q_MX04 U2162 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[2]), .A1(o_label2_data2[2]), .A2(o_label2_data3[2]), .A3(o_label2_data4[2]), .Z(n1762));
Q_MX04 U2163 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[2]), .A1(o_label3_data7[2]), .A2(o_label3_config[2]), .A3(o_label2_data0[2]), .Z(n1763));
Q_MX04 U2164 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[2]), .A1(o_label3_data3[2]), .A2(o_label3_data4[2]), .A3(o_label3_data5[2]), .Z(n1764));
Q_MX02 U2165 ( .S(n4414), .A0(o_label3_data0[2]), .A1(o_label3_data1[2]), .Z(n1765));
Q_AN02 U2166 ( .A0(n4414), .A1(o_label4_config[2]), .Z(n1766));
Q_MX02 U2167 ( .S(n4415), .A0(n1766), .A1(n1765), .Z(n1767));
Q_MX04 U2168 ( .S0(n4416), .S1(n4417), .A0(n1767), .A1(n1764), .A2(n1763), .A3(n1762), .Z(n1768));
Q_MX02 U2169 ( .S(n4418), .A0(n1768), .A1(n1761), .Z(r32_mux_4_data[2]));
Q_MX03 U2170 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[3]), .A1(o_label0_data0[3]), .A2(o_label0_data1[3]), .Z(n1769));
Q_MX04 U2171 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[3]), .A1(o_label1_data5[3]), .A2(o_label1_data6[3]), .A3(o_label1_data7[3]), .Z(n1770));
Q_MX02 U2172 ( .S(n4416), .A0(n1770), .A1(n1769), .Z(n1771));
Q_MX08 U2173 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[3]), .A1(o_label2_data6[3]), .A2(o_label2_data7[3]), .A3(o_label2_config[3]), .A4(o_label1_data0[3]), .A5(o_label1_data1[3]), .A6(o_label1_data2[3]), .A7(o_label1_data3[3]), .Z(n1772));
Q_MX02 U2174 ( .S(n4417), .A0(n1772), .A1(n1771), .Z(n1773));
Q_MX04 U2175 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[3]), .A1(o_label2_data2[3]), .A2(o_label2_data3[3]), .A3(o_label2_data4[3]), .Z(n1774));
Q_MX04 U2176 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[3]), .A1(o_label3_data7[3]), .A2(o_label3_config[3]), .A3(o_label2_data0[3]), .Z(n1775));
Q_MX04 U2177 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[3]), .A1(o_label3_data3[3]), .A2(o_label3_data4[3]), .A3(o_label3_data5[3]), .Z(n1776));
Q_MX02 U2178 ( .S(n4414), .A0(o_label3_data0[3]), .A1(o_label3_data1[3]), .Z(n1777));
Q_AN02 U2179 ( .A0(n4414), .A1(o_label4_config[3]), .Z(n1778));
Q_MX02 U2180 ( .S(n4415), .A0(n1778), .A1(n1777), .Z(n1779));
Q_MX04 U2181 ( .S0(n4416), .S1(n4417), .A0(n1779), .A1(n1776), .A2(n1775), .A3(n1774), .Z(n1780));
Q_MX02 U2182 ( .S(n4418), .A0(n1780), .A1(n1773), .Z(r32_mux_4_data[3]));
Q_MX03 U2183 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[4]), .A1(o_label0_data0[4]), .A2(o_label0_data1[4]), .Z(n1781));
Q_MX04 U2184 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[4]), .A1(o_label1_data5[4]), .A2(o_label1_data6[4]), .A3(o_label1_data7[4]), .Z(n1782));
Q_MX02 U2185 ( .S(n4416), .A0(n1782), .A1(n1781), .Z(n1783));
Q_MX08 U2186 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[4]), .A1(o_label2_data6[4]), .A2(o_label2_data7[4]), .A3(o_label2_config[4]), .A4(o_label1_data0[4]), .A5(o_label1_data1[4]), .A6(o_label1_data2[4]), .A7(o_label1_data3[4]), .Z(n1784));
Q_MX02 U2187 ( .S(n4417), .A0(n1784), .A1(n1783), .Z(n1785));
Q_MX04 U2188 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[4]), .A1(o_label2_data2[4]), .A2(o_label2_data3[4]), .A3(o_label2_data4[4]), .Z(n1786));
Q_MX04 U2189 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[4]), .A1(o_label3_data7[4]), .A2(o_label3_config[4]), .A3(o_label2_data0[4]), .Z(n1787));
Q_MX04 U2190 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[4]), .A1(o_label3_data3[4]), .A2(o_label3_data4[4]), .A3(o_label3_data5[4]), .Z(n1788));
Q_MX02 U2191 ( .S(n4414), .A0(o_label3_data0[4]), .A1(o_label3_data1[4]), .Z(n1789));
Q_AN02 U2192 ( .A0(n4414), .A1(o_label4_config[4]), .Z(n1790));
Q_MX02 U2193 ( .S(n4415), .A0(n1790), .A1(n1789), .Z(n1791));
Q_MX04 U2194 ( .S0(n4416), .S1(n4417), .A0(n1791), .A1(n1788), .A2(n1787), .A3(n1786), .Z(n1792));
Q_MX02 U2195 ( .S(n4418), .A0(n1792), .A1(n1785), .Z(r32_mux_4_data[4]));
Q_MX03 U2196 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[5]), .A1(o_label0_data0[5]), .A2(o_label0_data1[5]), .Z(n1793));
Q_MX04 U2197 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[5]), .A1(o_label1_data5[5]), .A2(o_label1_data6[5]), .A3(o_label1_data7[5]), .Z(n1794));
Q_MX02 U2198 ( .S(n4416), .A0(n1794), .A1(n1793), .Z(n1795));
Q_MX08 U2199 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[5]), .A1(o_label2_data6[5]), .A2(o_label2_data7[5]), .A3(o_label2_config[5]), .A4(o_label1_data0[5]), .A5(o_label1_data1[5]), .A6(o_label1_data2[5]), .A7(o_label1_data3[5]), .Z(n1796));
Q_MX02 U2200 ( .S(n4417), .A0(n1796), .A1(n1795), .Z(n1797));
Q_MX04 U2201 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[5]), .A1(o_label2_data2[5]), .A2(o_label2_data3[5]), .A3(o_label2_data4[5]), .Z(n1798));
Q_MX04 U2202 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[5]), .A1(o_label3_data7[5]), .A2(o_label3_config[5]), .A3(o_label2_data0[5]), .Z(n1799));
Q_MX04 U2203 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[5]), .A1(o_label3_data3[5]), .A2(o_label3_data4[5]), .A3(o_label3_data5[5]), .Z(n1800));
Q_MX02 U2204 ( .S(n4414), .A0(o_label3_data0[5]), .A1(o_label3_data1[5]), .Z(n1801));
Q_AN02 U2205 ( .A0(n4414), .A1(o_label4_config[5]), .Z(n1802));
Q_MX02 U2206 ( .S(n4415), .A0(n1802), .A1(n1801), .Z(n1803));
Q_MX04 U2207 ( .S0(n4416), .S1(n4417), .A0(n1803), .A1(n1800), .A2(n1799), .A3(n1798), .Z(n1804));
Q_MX02 U2208 ( .S(n4418), .A0(n1804), .A1(n1797), .Z(r32_mux_4_data[5]));
Q_MX03 U2209 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[6]), .A1(o_label0_data0[6]), .A2(o_label0_data1[6]), .Z(n1805));
Q_MX04 U2210 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[6]), .A1(o_label1_data5[6]), .A2(o_label1_data6[6]), .A3(o_label1_data7[6]), .Z(n1806));
Q_MX02 U2211 ( .S(n4416), .A0(n1806), .A1(n1805), .Z(n1807));
Q_MX08 U2212 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[6]), .A1(o_label2_data6[6]), .A2(o_label2_data7[6]), .A3(o_label2_config[6]), .A4(o_label1_data0[6]), .A5(o_label1_data1[6]), .A6(o_label1_data2[6]), .A7(o_label1_data3[6]), .Z(n1808));
Q_MX02 U2213 ( .S(n4417), .A0(n1808), .A1(n1807), .Z(n1809));
Q_MX04 U2214 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[6]), .A1(o_label2_data2[6]), .A2(o_label2_data3[6]), .A3(o_label2_data4[6]), .Z(n1810));
Q_MX04 U2215 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[6]), .A1(o_label3_data7[6]), .A2(o_label3_config[6]), .A3(o_label2_data0[6]), .Z(n1811));
Q_MX04 U2216 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[6]), .A1(o_label3_data3[6]), .A2(o_label3_data4[6]), .A3(o_label3_data5[6]), .Z(n1812));
Q_MX02 U2217 ( .S(n4414), .A0(o_label3_data0[6]), .A1(o_label3_data1[6]), .Z(n1813));
Q_AN02 U2218 ( .A0(n4414), .A1(o_label4_config[6]), .Z(n1814));
Q_MX02 U2219 ( .S(n4415), .A0(n1814), .A1(n1813), .Z(n1815));
Q_MX04 U2220 ( .S0(n4416), .S1(n4417), .A0(n1815), .A1(n1812), .A2(n1811), .A3(n1810), .Z(n1816));
Q_MX02 U2221 ( .S(n4418), .A0(n1816), .A1(n1809), .Z(r32_mux_4_data[6]));
Q_MX03 U2222 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[7]), .A1(o_label0_data0[7]), .A2(o_label0_data1[7]), .Z(n1817));
Q_MX04 U2223 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[7]), .A1(o_label1_data5[7]), .A2(o_label1_data6[7]), .A3(o_label1_data7[7]), .Z(n1818));
Q_MX02 U2224 ( .S(n4416), .A0(n1818), .A1(n1817), .Z(n1819));
Q_MX08 U2225 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[7]), .A1(o_label2_data6[7]), .A2(o_label2_data7[7]), .A3(o_label2_config[7]), .A4(o_label1_data0[7]), .A5(o_label1_data1[7]), .A6(o_label1_data2[7]), .A7(o_label1_data3[7]), .Z(n1820));
Q_MX02 U2226 ( .S(n4417), .A0(n1820), .A1(n1819), .Z(n1821));
Q_MX04 U2227 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[7]), .A1(o_label2_data2[7]), .A2(o_label2_data3[7]), .A3(o_label2_data4[7]), .Z(n1822));
Q_MX04 U2228 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[7]), .A1(o_label3_data7[7]), .A2(o_label3_config[7]), .A3(o_label2_data0[7]), .Z(n1823));
Q_MX04 U2229 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[7]), .A1(o_label3_data3[7]), .A2(o_label3_data4[7]), .A3(o_label3_data5[7]), .Z(n1824));
Q_MX02 U2230 ( .S(n4414), .A0(o_label3_data0[7]), .A1(o_label3_data1[7]), .Z(n1825));
Q_AN02 U2231 ( .A0(n4414), .A1(o_label4_config[7]), .Z(n1826));
Q_MX02 U2232 ( .S(n4415), .A0(n1826), .A1(n1825), .Z(n1827));
Q_MX04 U2233 ( .S0(n4416), .S1(n4417), .A0(n1827), .A1(n1824), .A2(n1823), .A3(n1822), .Z(n1828));
Q_MX02 U2234 ( .S(n4418), .A0(n1828), .A1(n1821), .Z(r32_mux_4_data[7]));
Q_MX03 U2235 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[8]), .A1(o_label0_data0[8]), .A2(o_label0_data1[8]), .Z(n1829));
Q_MX04 U2236 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[8]), .A1(o_label1_data5[8]), .A2(o_label1_data6[8]), .A3(o_label1_data7[8]), .Z(n1830));
Q_MX02 U2237 ( .S(n4416), .A0(n1830), .A1(n1829), .Z(n1831));
Q_MX08 U2238 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[8]), .A1(o_label2_data6[8]), .A2(o_label2_data7[8]), .A3(o_label2_config[8]), .A4(o_label1_data0[8]), .A5(o_label1_data1[8]), .A6(o_label1_data2[8]), .A7(o_label1_data3[8]), .Z(n1832));
Q_MX02 U2239 ( .S(n4417), .A0(n1832), .A1(n1831), .Z(n1833));
Q_MX04 U2240 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[8]), .A1(o_label2_data2[8]), .A2(o_label2_data3[8]), .A3(o_label2_data4[8]), .Z(n1834));
Q_MX04 U2241 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[8]), .A1(o_label3_data7[8]), .A2(o_label3_config[8]), .A3(o_label2_data0[8]), .Z(n1835));
Q_MX04 U2242 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[8]), .A1(o_label3_data3[8]), .A2(o_label3_data4[8]), .A3(o_label3_data5[8]), .Z(n1836));
Q_MX02 U2243 ( .S(n4414), .A0(o_label3_data0[8]), .A1(o_label3_data1[8]), .Z(n1837));
Q_AN02 U2244 ( .A0(n4414), .A1(o_label4_config[8]), .Z(n1838));
Q_MX02 U2245 ( .S(n4415), .A0(n1838), .A1(n1837), .Z(n1839));
Q_MX04 U2246 ( .S0(n4416), .S1(n4417), .A0(n1839), .A1(n1836), .A2(n1835), .A3(n1834), .Z(n1840));
Q_MX02 U2247 ( .S(n4418), .A0(n1840), .A1(n1833), .Z(r32_mux_4_data[8]));
Q_MX03 U2248 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[9]), .A1(o_label0_data0[9]), .A2(o_label0_data1[9]), .Z(n1841));
Q_MX08 U2249 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[9]), .A1(o_label1_data0[9]), .A2(o_label1_data1[9]), .A3(o_label1_data2[9]), .A4(o_label1_data3[9]), .A5(o_label1_data4[9]), .A6(o_label1_data5[9]), .A7(o_label1_data6[9]), .Z(n1842));
Q_MX02 U2250 ( .S(n4422), .A0(n1842), .A1(n1841), .Z(n1843));
Q_MX04 U2251 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[9]), .A1(o_label2_data4[9]), .A2(o_label2_data5[9]), .A3(o_label2_data6[9]), .Z(n1844));
Q_MX04 U2252 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[9]), .A1(o_label2_data0[9]), .A2(o_label2_data1[9]), .A3(o_label2_data2[9]), .Z(n1845));
Q_MX04 U2253 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[9]), .A1(o_label3_data4[9]), .A2(o_label3_data5[9]), .A3(o_label3_data6[9]), .Z(n1846));
Q_MX02 U2254 ( .S(n4419), .A0(o_label3_data1[9]), .A1(o_label3_data2[9]), .Z(n1847));
Q_AN02 U2255 ( .A0(n4419), .A1(o_label3_data0[9]), .Z(n1848));
Q_MX02 U2256 ( .S(n4420), .A0(n1848), .A1(n1847), .Z(n1849));
Q_MX04 U2257 ( .S0(n4421), .S1(n4422), .A0(n1849), .A1(n1846), .A2(n1845), .A3(n1844), .Z(n1850));
Q_MX02 U2258 ( .S(n4423), .A0(n1850), .A1(n1843), .Z(r32_mux_4_data[9]));
Q_MX03 U2259 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[10]), .A1(o_label0_data0[10]), .A2(o_label0_data1[10]), .Z(n1851));
Q_MX08 U2260 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[10]), .A1(o_label1_data0[10]), .A2(o_label1_data1[10]), .A3(o_label1_data2[10]), .A4(o_label1_data3[10]), .A5(o_label1_data4[10]), .A6(o_label1_data5[10]), .A7(o_label1_data6[10]), .Z(n1852));
Q_MX02 U2261 ( .S(n4422), .A0(n1852), .A1(n1851), .Z(n1853));
Q_MX04 U2262 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[10]), .A1(o_label2_data4[10]), .A2(o_label2_data5[10]), .A3(o_label2_data6[10]), .Z(n1854));
Q_MX04 U2263 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[10]), .A1(o_label2_data0[10]), .A2(o_label2_data1[10]), .A3(o_label2_data2[10]), .Z(n1855));
Q_MX04 U2264 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[10]), .A1(o_label3_data4[10]), .A2(o_label3_data5[10]), .A3(o_label3_data6[10]), .Z(n1856));
Q_MX02 U2265 ( .S(n4419), .A0(o_label3_data1[10]), .A1(o_label3_data2[10]), .Z(n1857));
Q_AN02 U2266 ( .A0(n4419), .A1(o_label3_data0[10]), .Z(n1858));
Q_MX02 U2267 ( .S(n4420), .A0(n1858), .A1(n1857), .Z(n1859));
Q_MX04 U2268 ( .S0(n4421), .S1(n4422), .A0(n1859), .A1(n1856), .A2(n1855), .A3(n1854), .Z(n1860));
Q_MX02 U2269 ( .S(n4423), .A0(n1860), .A1(n1853), .Z(r32_mux_4_data[10]));
Q_MX03 U2270 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[11]), .A1(o_label0_data0[11]), .A2(o_label0_data1[11]), .Z(n1861));
Q_MX08 U2271 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[11]), .A1(o_label1_data0[11]), .A2(o_label1_data1[11]), .A3(o_label1_data2[11]), .A4(o_label1_data3[11]), .A5(o_label1_data4[11]), .A6(o_label1_data5[11]), .A7(o_label1_data6[11]), .Z(n1862));
Q_MX02 U2272 ( .S(n4422), .A0(n1862), .A1(n1861), .Z(n1863));
Q_MX04 U2273 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[11]), .A1(o_label2_data4[11]), .A2(o_label2_data5[11]), .A3(o_label2_data6[11]), .Z(n1864));
Q_MX04 U2274 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[11]), .A1(o_label2_data0[11]), .A2(o_label2_data1[11]), .A3(o_label2_data2[11]), .Z(n1865));
Q_MX04 U2275 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[11]), .A1(o_label3_data4[11]), .A2(o_label3_data5[11]), .A3(o_label3_data6[11]), .Z(n1866));
Q_MX02 U2276 ( .S(n4419), .A0(o_label3_data1[11]), .A1(o_label3_data2[11]), .Z(n1867));
Q_AN02 U2277 ( .A0(n4419), .A1(o_label3_data0[11]), .Z(n1868));
Q_MX02 U2278 ( .S(n4420), .A0(n1868), .A1(n1867), .Z(n1869));
Q_MX04 U2279 ( .S0(n4421), .S1(n4422), .A0(n1869), .A1(n1866), .A2(n1865), .A3(n1864), .Z(n1870));
Q_MX02 U2280 ( .S(n4423), .A0(n1870), .A1(n1863), .Z(r32_mux_4_data[11]));
Q_MX03 U2281 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[12]), .A1(o_label0_data0[12]), .A2(o_label0_data1[12]), .Z(n1871));
Q_MX08 U2282 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[12]), .A1(o_label1_data0[12]), .A2(o_label1_data1[12]), .A3(o_label1_data2[12]), .A4(o_label1_data3[12]), .A5(o_label1_data4[12]), .A6(o_label1_data5[12]), .A7(o_label1_data6[12]), .Z(n1872));
Q_MX02 U2283 ( .S(n4422), .A0(n1872), .A1(n1871), .Z(n1873));
Q_MX04 U2284 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[12]), .A1(o_label2_data4[12]), .A2(o_label2_data5[12]), .A3(o_label2_data6[12]), .Z(n1874));
Q_MX04 U2285 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[12]), .A1(o_label2_data0[12]), .A2(o_label2_data1[12]), .A3(o_label2_data2[12]), .Z(n1875));
Q_MX04 U2286 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[12]), .A1(o_label3_data4[12]), .A2(o_label3_data5[12]), .A3(o_label3_data6[12]), .Z(n1876));
Q_MX02 U2287 ( .S(n4419), .A0(o_label3_data1[12]), .A1(o_label3_data2[12]), .Z(n1877));
Q_AN02 U2288 ( .A0(n4419), .A1(o_label3_data0[12]), .Z(n1878));
Q_MX02 U2289 ( .S(n4420), .A0(n1878), .A1(n1877), .Z(n1879));
Q_MX04 U2290 ( .S0(n4421), .S1(n4422), .A0(n1879), .A1(n1876), .A2(n1875), .A3(n1874), .Z(n1880));
Q_MX02 U2291 ( .S(n4423), .A0(n1880), .A1(n1873), .Z(r32_mux_4_data[12]));
Q_MX03 U2292 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[13]), .A1(o_label0_data0[13]), .A2(o_label0_data1[13]), .Z(n1881));
Q_MX08 U2293 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[13]), .A1(o_label1_data0[13]), .A2(o_label1_data1[13]), .A3(o_label1_data2[13]), .A4(o_label1_data3[13]), .A5(o_label1_data4[13]), .A6(o_label1_data5[13]), .A7(o_label1_data6[13]), .Z(n1882));
Q_MX02 U2294 ( .S(n4422), .A0(n1882), .A1(n1881), .Z(n1883));
Q_MX04 U2295 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[13]), .A1(o_label2_data4[13]), .A2(o_label2_data5[13]), .A3(o_label2_data6[13]), .Z(n1884));
Q_MX04 U2296 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[13]), .A1(o_label2_data0[13]), .A2(o_label2_data1[13]), .A3(o_label2_data2[13]), .Z(n1885));
Q_MX04 U2297 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[13]), .A1(o_label3_data4[13]), .A2(o_label3_data5[13]), .A3(o_label3_data6[13]), .Z(n1886));
Q_MX02 U2298 ( .S(n4419), .A0(o_label3_data1[13]), .A1(o_label3_data2[13]), .Z(n1887));
Q_AN02 U2299 ( .A0(n4419), .A1(o_label3_data0[13]), .Z(n1888));
Q_MX02 U2300 ( .S(n4420), .A0(n1888), .A1(n1887), .Z(n1889));
Q_MX04 U2301 ( .S0(n4421), .S1(n4422), .A0(n1889), .A1(n1886), .A2(n1885), .A3(n1884), .Z(n1890));
Q_MX02 U2302 ( .S(n4423), .A0(n1890), .A1(n1883), .Z(r32_mux_4_data[13]));
Q_MX03 U2303 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[14]), .A1(o_label0_data0[14]), .A2(o_label0_data1[14]), .Z(n1891));
Q_MX08 U2304 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[14]), .A1(o_label1_data0[14]), .A2(o_label1_data1[14]), .A3(o_label1_data2[14]), .A4(o_label1_data3[14]), .A5(o_label1_data4[14]), .A6(o_label1_data5[14]), .A7(o_label1_data6[14]), .Z(n1892));
Q_MX02 U2305 ( .S(n4422), .A0(n1892), .A1(n1891), .Z(n1893));
Q_MX04 U2306 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[14]), .A1(o_label2_data4[14]), .A2(o_label2_data5[14]), .A3(o_label2_data6[14]), .Z(n1894));
Q_MX04 U2307 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[14]), .A1(o_label2_data0[14]), .A2(o_label2_data1[14]), .A3(o_label2_data2[14]), .Z(n1895));
Q_MX04 U2308 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[14]), .A1(o_label3_data4[14]), .A2(o_label3_data5[14]), .A3(o_label3_data6[14]), .Z(n1896));
Q_MX02 U2309 ( .S(n4419), .A0(o_label3_data1[14]), .A1(o_label3_data2[14]), .Z(n1897));
Q_AN02 U2310 ( .A0(n4419), .A1(o_label3_data0[14]), .Z(n1898));
Q_MX02 U2311 ( .S(n4420), .A0(n1898), .A1(n1897), .Z(n1899));
Q_MX04 U2312 ( .S0(n4421), .S1(n4422), .A0(n1899), .A1(n1896), .A2(n1895), .A3(n1894), .Z(n1900));
Q_MX02 U2313 ( .S(n4423), .A0(n1900), .A1(n1893), .Z(r32_mux_4_data[14]));
Q_MX03 U2314 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[15]), .A1(o_label0_data0[15]), .A2(o_label0_data1[15]), .Z(n1901));
Q_MX08 U2315 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[15]), .A1(o_label1_data0[15]), .A2(o_label1_data1[15]), .A3(o_label1_data2[15]), .A4(o_label1_data3[15]), .A5(o_label1_data4[15]), .A6(o_label1_data5[15]), .A7(o_label1_data6[15]), .Z(n1902));
Q_MX02 U2316 ( .S(n4422), .A0(n1902), .A1(n1901), .Z(n1903));
Q_MX04 U2317 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[15]), .A1(o_label2_data4[15]), .A2(o_label2_data5[15]), .A3(o_label2_data6[15]), .Z(n1904));
Q_MX04 U2318 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[15]), .A1(o_label2_data0[15]), .A2(o_label2_data1[15]), .A3(o_label2_data2[15]), .Z(n1905));
Q_MX04 U2319 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[15]), .A1(o_label3_data4[15]), .A2(o_label3_data5[15]), .A3(o_label3_data6[15]), .Z(n1906));
Q_MX02 U2320 ( .S(n4419), .A0(o_label3_data1[15]), .A1(o_label3_data2[15]), .Z(n1907));
Q_AN02 U2321 ( .A0(n4419), .A1(o_label3_data0[15]), .Z(n1908));
Q_MX02 U2322 ( .S(n4420), .A0(n1908), .A1(n1907), .Z(n1909));
Q_MX04 U2323 ( .S0(n4421), .S1(n4422), .A0(n1909), .A1(n1906), .A2(n1905), .A3(n1904), .Z(n1910));
Q_MX02 U2324 ( .S(n4423), .A0(n1910), .A1(n1903), .Z(r32_mux_4_data[15]));
Q_MX03 U2325 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[16]), .A1(o_label0_data0[16]), .A2(o_label0_data1[16]), .Z(n1911));
Q_MX08 U2326 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[16]), .A1(o_label1_data0[16]), .A2(o_label1_data1[16]), .A3(o_label1_data2[16]), .A4(o_label1_data3[16]), .A5(o_label1_data4[16]), .A6(o_label1_data5[16]), .A7(o_label1_data6[16]), .Z(n1912));
Q_MX02 U2327 ( .S(n4422), .A0(n1912), .A1(n1911), .Z(n1913));
Q_MX04 U2328 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[16]), .A1(o_label2_data4[16]), .A2(o_label2_data5[16]), .A3(o_label2_data6[16]), .Z(n1914));
Q_MX04 U2329 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[16]), .A1(o_label2_data0[16]), .A2(o_label2_data1[16]), .A3(o_label2_data2[16]), .Z(n1915));
Q_MX04 U2330 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[16]), .A1(o_label3_data4[16]), .A2(o_label3_data5[16]), .A3(o_label3_data6[16]), .Z(n1916));
Q_MX02 U2331 ( .S(n4419), .A0(o_label3_data1[16]), .A1(o_label3_data2[16]), .Z(n1917));
Q_AN02 U2332 ( .A0(n4419), .A1(o_label3_data0[16]), .Z(n1918));
Q_MX02 U2333 ( .S(n4420), .A0(n1918), .A1(n1917), .Z(n1919));
Q_MX04 U2334 ( .S0(n4421), .S1(n4422), .A0(n1919), .A1(n1916), .A2(n1915), .A3(n1914), .Z(n1920));
Q_MX02 U2335 ( .S(n4423), .A0(n1920), .A1(n1913), .Z(r32_mux_4_data[16]));
Q_MX03 U2336 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[17]), .A1(o_label0_data0[17]), .A2(o_label0_data1[17]), .Z(n1921));
Q_MX08 U2337 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[17]), .A1(o_label1_data0[17]), .A2(o_label1_data1[17]), .A3(o_label1_data2[17]), .A4(o_label1_data3[17]), .A5(o_label1_data4[17]), .A6(o_label1_data5[17]), .A7(o_label1_data6[17]), .Z(n1922));
Q_MX02 U2338 ( .S(n4422), .A0(n1922), .A1(n1921), .Z(n1923));
Q_MX04 U2339 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[17]), .A1(o_label2_data4[17]), .A2(o_label2_data5[17]), .A3(o_label2_data6[17]), .Z(n1924));
Q_MX04 U2340 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[17]), .A1(o_label2_data0[17]), .A2(o_label2_data1[17]), .A3(o_label2_data2[17]), .Z(n1925));
Q_MX04 U2341 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[17]), .A1(o_label3_data4[17]), .A2(o_label3_data5[17]), .A3(o_label3_data6[17]), .Z(n1926));
Q_MX02 U2342 ( .S(n4419), .A0(o_label3_data1[17]), .A1(o_label3_data2[17]), .Z(n1927));
Q_AN02 U2343 ( .A0(n4419), .A1(o_label3_data0[17]), .Z(n1928));
Q_MX02 U2344 ( .S(n4420), .A0(n1928), .A1(n1927), .Z(n1929));
Q_MX04 U2345 ( .S0(n4421), .S1(n4422), .A0(n1929), .A1(n1926), .A2(n1925), .A3(n1924), .Z(n1930));
Q_MX02 U2346 ( .S(n4423), .A0(n1930), .A1(n1923), .Z(r32_mux_4_data[17]));
Q_MX03 U2347 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[18]), .A1(o_label0_data0[18]), .A2(o_label0_data1[18]), .Z(n1931));
Q_MX08 U2348 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[18]), .A1(o_label1_data0[18]), .A2(o_label1_data1[18]), .A3(o_label1_data2[18]), .A4(o_label1_data3[18]), .A5(o_label1_data4[18]), .A6(o_label1_data5[18]), .A7(o_label1_data6[18]), .Z(n1932));
Q_MX02 U2349 ( .S(n4422), .A0(n1932), .A1(n1931), .Z(n1933));
Q_MX04 U2350 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[18]), .A1(o_label2_data4[18]), .A2(o_label2_data5[18]), .A3(o_label2_data6[18]), .Z(n1934));
Q_MX04 U2351 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[18]), .A1(o_label2_data0[18]), .A2(o_label2_data1[18]), .A3(o_label2_data2[18]), .Z(n1935));
Q_MX04 U2352 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[18]), .A1(o_label3_data4[18]), .A2(o_label3_data5[18]), .A3(o_label3_data6[18]), .Z(n1936));
Q_MX02 U2353 ( .S(n4419), .A0(o_label3_data1[18]), .A1(o_label3_data2[18]), .Z(n1937));
Q_AN02 U2354 ( .A0(n4419), .A1(o_label3_data0[18]), .Z(n1938));
Q_MX02 U2355 ( .S(n4420), .A0(n1938), .A1(n1937), .Z(n1939));
Q_MX04 U2356 ( .S0(n4421), .S1(n4422), .A0(n1939), .A1(n1936), .A2(n1935), .A3(n1934), .Z(n1940));
Q_MX02 U2357 ( .S(n4423), .A0(n1940), .A1(n1933), .Z(r32_mux_4_data[18]));
Q_MX03 U2358 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[19]), .A1(o_label0_data0[19]), .A2(o_label0_data1[19]), .Z(n1941));
Q_MX08 U2359 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[19]), .A1(o_label1_data0[19]), .A2(o_label1_data1[19]), .A3(o_label1_data2[19]), .A4(o_label1_data3[19]), .A5(o_label1_data4[19]), .A6(o_label1_data5[19]), .A7(o_label1_data6[19]), .Z(n1942));
Q_MX02 U2360 ( .S(n4422), .A0(n1942), .A1(n1941), .Z(n1943));
Q_MX04 U2361 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[19]), .A1(o_label2_data4[19]), .A2(o_label2_data5[19]), .A3(o_label2_data6[19]), .Z(n1944));
Q_MX04 U2362 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[19]), .A1(o_label2_data0[19]), .A2(o_label2_data1[19]), .A3(o_label2_data2[19]), .Z(n1945));
Q_MX04 U2363 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[19]), .A1(o_label3_data4[19]), .A2(o_label3_data5[19]), .A3(o_label3_data6[19]), .Z(n1946));
Q_MX02 U2364 ( .S(n4419), .A0(o_label3_data1[19]), .A1(o_label3_data2[19]), .Z(n1947));
Q_AN02 U2365 ( .A0(n4419), .A1(o_label3_data0[19]), .Z(n1948));
Q_MX02 U2366 ( .S(n4420), .A0(n1948), .A1(n1947), .Z(n1949));
Q_MX04 U2367 ( .S0(n4421), .S1(n4422), .A0(n1949), .A1(n1946), .A2(n1945), .A3(n1944), .Z(n1950));
Q_MX02 U2368 ( .S(n4423), .A0(n1950), .A1(n1943), .Z(r32_mux_4_data[19]));
Q_MX03 U2369 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[20]), .A1(o_label0_data0[20]), .A2(o_label0_data1[20]), .Z(n1951));
Q_MX08 U2370 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[20]), .A1(o_label1_data0[20]), .A2(o_label1_data1[20]), .A3(o_label1_data2[20]), .A4(o_label1_data3[20]), .A5(o_label1_data4[20]), .A6(o_label1_data5[20]), .A7(o_label1_data6[20]), .Z(n1952));
Q_MX02 U2371 ( .S(n4422), .A0(n1952), .A1(n1951), .Z(n1953));
Q_MX04 U2372 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[20]), .A1(o_label2_data4[20]), .A2(o_label2_data5[20]), .A3(o_label2_data6[20]), .Z(n1954));
Q_MX04 U2373 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[20]), .A1(o_label2_data0[20]), .A2(o_label2_data1[20]), .A3(o_label2_data2[20]), .Z(n1955));
Q_MX04 U2374 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[20]), .A1(o_label3_data4[20]), .A2(o_label3_data5[20]), .A3(o_label3_data6[20]), .Z(n1956));
Q_MX02 U2375 ( .S(n4419), .A0(o_label3_data1[20]), .A1(o_label3_data2[20]), .Z(n1957));
Q_AN02 U2376 ( .A0(n4419), .A1(o_label3_data0[20]), .Z(n1958));
Q_MX02 U2377 ( .S(n4420), .A0(n1958), .A1(n1957), .Z(n1959));
Q_MX04 U2378 ( .S0(n4421), .S1(n4422), .A0(n1959), .A1(n1956), .A2(n1955), .A3(n1954), .Z(n1960));
Q_MX02 U2379 ( .S(n4423), .A0(n1960), .A1(n1953), .Z(r32_mux_4_data[20]));
Q_MX03 U2380 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[21]), .A1(o_label0_data0[21]), .A2(o_label0_data1[21]), .Z(n1961));
Q_MX08 U2381 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[21]), .A1(o_label1_data0[21]), .A2(o_label1_data1[21]), .A3(o_label1_data2[21]), .A4(o_label1_data3[21]), .A5(o_label1_data4[21]), .A6(o_label1_data5[21]), .A7(o_label1_data6[21]), .Z(n1962));
Q_MX02 U2382 ( .S(n4422), .A0(n1962), .A1(n1961), .Z(n1963));
Q_MX04 U2383 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[21]), .A1(o_label2_data4[21]), .A2(o_label2_data5[21]), .A3(o_label2_data6[21]), .Z(n1964));
Q_MX04 U2384 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[21]), .A1(o_label2_data0[21]), .A2(o_label2_data1[21]), .A3(o_label2_data2[21]), .Z(n1965));
Q_MX04 U2385 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[21]), .A1(o_label3_data4[21]), .A2(o_label3_data5[21]), .A3(o_label3_data6[21]), .Z(n1966));
Q_MX02 U2386 ( .S(n4419), .A0(o_label3_data1[21]), .A1(o_label3_data2[21]), .Z(n1967));
Q_AN02 U2387 ( .A0(n4419), .A1(o_label3_data0[21]), .Z(n1968));
Q_MX02 U2388 ( .S(n4420), .A0(n1968), .A1(n1967), .Z(n1969));
Q_MX04 U2389 ( .S0(n4421), .S1(n4422), .A0(n1969), .A1(n1966), .A2(n1965), .A3(n1964), .Z(n1970));
Q_MX02 U2390 ( .S(n4423), .A0(n1970), .A1(n1963), .Z(r32_mux_4_data[21]));
Q_MX03 U2391 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[22]), .A1(o_label0_data0[22]), .A2(o_label0_data1[22]), .Z(n1971));
Q_MX08 U2392 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[22]), .A1(o_label1_data0[22]), .A2(o_label1_data1[22]), .A3(o_label1_data2[22]), .A4(o_label1_data3[22]), .A5(o_label1_data4[22]), .A6(o_label1_data5[22]), .A7(o_label1_data6[22]), .Z(n1972));
Q_MX02 U2393 ( .S(n4422), .A0(n1972), .A1(n1971), .Z(n1973));
Q_MX04 U2394 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[22]), .A1(o_label2_data4[22]), .A2(o_label2_data5[22]), .A3(o_label2_data6[22]), .Z(n1974));
Q_MX04 U2395 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[22]), .A1(o_label2_data0[22]), .A2(o_label2_data1[22]), .A3(o_label2_data2[22]), .Z(n1975));
Q_MX04 U2396 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[22]), .A1(o_label3_data4[22]), .A2(o_label3_data5[22]), .A3(o_label3_data6[22]), .Z(n1976));
Q_MX02 U2397 ( .S(n4419), .A0(o_label3_data1[22]), .A1(o_label3_data2[22]), .Z(n1977));
Q_AN02 U2398 ( .A0(n4419), .A1(o_label3_data0[22]), .Z(n1978));
Q_MX02 U2399 ( .S(n4420), .A0(n1978), .A1(n1977), .Z(n1979));
Q_MX04 U2400 ( .S0(n4421), .S1(n4422), .A0(n1979), .A1(n1976), .A2(n1975), .A3(n1974), .Z(n1980));
Q_MX02 U2401 ( .S(n4423), .A0(n1980), .A1(n1973), .Z(r32_mux_4_data[22]));
Q_MX03 U2402 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[23]), .A1(o_label0_data0[23]), .A2(o_label0_data1[23]), .Z(n1981));
Q_MX08 U2403 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[23]), .A1(o_label1_data0[23]), .A2(o_label1_data1[23]), .A3(o_label1_data2[23]), .A4(o_label1_data3[23]), .A5(o_label1_data4[23]), .A6(o_label1_data5[23]), .A7(o_label1_data6[23]), .Z(n1982));
Q_MX02 U2404 ( .S(n4422), .A0(n1982), .A1(n1981), .Z(n1983));
Q_MX04 U2405 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[23]), .A1(o_label2_data4[23]), .A2(o_label2_data5[23]), .A3(o_label2_data6[23]), .Z(n1984));
Q_MX04 U2406 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[23]), .A1(o_label2_data0[23]), .A2(o_label2_data1[23]), .A3(o_label2_data2[23]), .Z(n1985));
Q_MX04 U2407 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[23]), .A1(o_label3_data4[23]), .A2(o_label3_data5[23]), .A3(o_label3_data6[23]), .Z(n1986));
Q_MX02 U2408 ( .S(n4419), .A0(o_label3_data1[23]), .A1(o_label3_data2[23]), .Z(n1987));
Q_AN02 U2409 ( .A0(n4419), .A1(o_label3_data0[23]), .Z(n1988));
Q_MX02 U2410 ( .S(n4420), .A0(n1988), .A1(n1987), .Z(n1989));
Q_MX04 U2411 ( .S0(n4421), .S1(n4422), .A0(n1989), .A1(n1986), .A2(n1985), .A3(n1984), .Z(n1990));
Q_MX02 U2412 ( .S(n4423), .A0(n1990), .A1(n1983), .Z(r32_mux_4_data[23]));
Q_MX03 U2413 ( .S0(n4419), .S1(n4420), .A0(o_label1_data7[24]), .A1(o_label0_data0[24]), .A2(o_label0_data1[24]), .Z(n1991));
Q_MX08 U2414 ( .S0(n4419), .S1(n4420), .S2(n4421), .A0(o_label2_data7[24]), .A1(o_label1_data0[24]), .A2(o_label1_data1[24]), .A3(o_label1_data2[24]), .A4(o_label1_data3[24]), .A5(o_label1_data4[24]), .A6(o_label1_data5[24]), .A7(o_label1_data6[24]), .Z(n1992));
Q_MX02 U2415 ( .S(n4422), .A0(n1992), .A1(n1991), .Z(n1993));
Q_MX04 U2416 ( .S0(n4419), .S1(n4420), .A0(o_label2_data3[24]), .A1(o_label2_data4[24]), .A2(o_label2_data5[24]), .A3(o_label2_data6[24]), .Z(n1994));
Q_MX04 U2417 ( .S0(n4419), .S1(n4420), .A0(o_label3_data7[24]), .A1(o_label2_data0[24]), .A2(o_label2_data1[24]), .A3(o_label2_data2[24]), .Z(n1995));
Q_MX04 U2418 ( .S0(n4419), .S1(n4420), .A0(o_label3_data3[24]), .A1(o_label3_data4[24]), .A2(o_label3_data5[24]), .A3(o_label3_data6[24]), .Z(n1996));
Q_MX02 U2419 ( .S(n4419), .A0(o_label3_data1[24]), .A1(o_label3_data2[24]), .Z(n1997));
Q_AN02 U2420 ( .A0(n4419), .A1(o_label3_data0[24]), .Z(n1998));
Q_MX02 U2421 ( .S(n4420), .A0(n1998), .A1(n1997), .Z(n1999));
Q_MX04 U2422 ( .S0(n4421), .S1(n4422), .A0(n1999), .A1(n1996), .A2(n1995), .A3(n1994), .Z(n2000));
Q_MX02 U2423 ( .S(n4423), .A0(n2000), .A1(n1993), .Z(r32_mux_4_data[24]));
Q_MX03 U2424 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[9]), .A1(o_label0_data0[25]), .A2(o_label0_data1[25]), .Z(n2001));
Q_MX04 U2425 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[25]), .A1(o_label1_data5[25]), .A2(o_label1_data6[25]), .A3(o_label1_data7[25]), .Z(n2002));
Q_MX02 U2426 ( .S(n4416), .A0(n2002), .A1(n2001), .Z(n2003));
Q_MX08 U2427 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[25]), .A1(o_label2_data6[25]), .A2(o_label2_data7[25]), .A3(o_label2_config[9]), .A4(o_label1_data0[25]), .A5(o_label1_data1[25]), .A6(o_label1_data2[25]), .A7(o_label1_data3[25]), .Z(n2004));
Q_MX02 U2428 ( .S(n4417), .A0(n2004), .A1(n2003), .Z(n2005));
Q_MX04 U2429 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[25]), .A1(o_label2_data2[25]), .A2(o_label2_data3[25]), .A3(o_label2_data4[25]), .Z(n2006));
Q_MX04 U2430 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[25]), .A1(o_label3_data7[25]), .A2(o_label3_config[9]), .A3(o_label2_data0[25]), .Z(n2007));
Q_MX04 U2431 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[25]), .A1(o_label3_data3[25]), .A2(o_label3_data4[25]), .A3(o_label3_data5[25]), .Z(n2008));
Q_MX02 U2432 ( .S(n4414), .A0(o_label3_data0[25]), .A1(o_label3_data1[25]), .Z(n2009));
Q_AN02 U2433 ( .A0(n4414), .A1(o_label4_config[9]), .Z(n2010));
Q_MX02 U2434 ( .S(n4415), .A0(n2010), .A1(n2009), .Z(n2011));
Q_MX04 U2435 ( .S0(n4416), .S1(n4417), .A0(n2011), .A1(n2008), .A2(n2007), .A3(n2006), .Z(n2012));
Q_MX02 U2436 ( .S(n4418), .A0(n2012), .A1(n2005), .Z(r32_mux_4_data[25]));
Q_MX03 U2437 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[10]), .A1(o_label0_data0[26]), .A2(o_label0_data1[26]), .Z(n2013));
Q_MX04 U2438 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[26]), .A1(o_label1_data5[26]), .A2(o_label1_data6[26]), .A3(o_label1_data7[26]), .Z(n2014));
Q_MX02 U2439 ( .S(n4416), .A0(n2014), .A1(n2013), .Z(n2015));
Q_MX08 U2440 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[26]), .A1(o_label2_data6[26]), .A2(o_label2_data7[26]), .A3(o_label2_config[10]), .A4(o_label1_data0[26]), .A5(o_label1_data1[26]), .A6(o_label1_data2[26]), .A7(o_label1_data3[26]), .Z(n2016));
Q_MX02 U2441 ( .S(n4417), .A0(n2016), .A1(n2015), .Z(n2017));
Q_MX04 U2442 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[26]), .A1(o_label2_data2[26]), .A2(o_label2_data3[26]), .A3(o_label2_data4[26]), .Z(n2018));
Q_MX04 U2443 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[26]), .A1(o_label3_data7[26]), .A2(o_label3_config[10]), .A3(o_label2_data0[26]), .Z(n2019));
Q_MX04 U2444 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[26]), .A1(o_label3_data3[26]), .A2(o_label3_data4[26]), .A3(o_label3_data5[26]), .Z(n2020));
Q_MX02 U2445 ( .S(n4414), .A0(o_label3_data0[26]), .A1(o_label3_data1[26]), .Z(n2021));
Q_AN02 U2446 ( .A0(n4414), .A1(o_label4_config[10]), .Z(n2022));
Q_MX02 U2447 ( .S(n4415), .A0(n2022), .A1(n2021), .Z(n2023));
Q_MX04 U2448 ( .S0(n4416), .S1(n4417), .A0(n2023), .A1(n2020), .A2(n2019), .A3(n2018), .Z(n2024));
Q_MX02 U2449 ( .S(n4418), .A0(n2024), .A1(n2017), .Z(r32_mux_4_data[26]));
Q_MX03 U2450 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[11]), .A1(o_label0_data0[27]), .A2(o_label0_data1[27]), .Z(n2025));
Q_MX04 U2451 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[27]), .A1(o_label1_data5[27]), .A2(o_label1_data6[27]), .A3(o_label1_data7[27]), .Z(n2026));
Q_MX02 U2452 ( .S(n4416), .A0(n2026), .A1(n2025), .Z(n2027));
Q_MX08 U2453 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[27]), .A1(o_label2_data6[27]), .A2(o_label2_data7[27]), .A3(o_label2_config[11]), .A4(o_label1_data0[27]), .A5(o_label1_data1[27]), .A6(o_label1_data2[27]), .A7(o_label1_data3[27]), .Z(n2028));
Q_MX02 U2454 ( .S(n4417), .A0(n2028), .A1(n2027), .Z(n2029));
Q_MX04 U2455 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[27]), .A1(o_label2_data2[27]), .A2(o_label2_data3[27]), .A3(o_label2_data4[27]), .Z(n2030));
Q_MX04 U2456 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[27]), .A1(o_label3_data7[27]), .A2(o_label3_config[11]), .A3(o_label2_data0[27]), .Z(n2031));
Q_MX04 U2457 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[27]), .A1(o_label3_data3[27]), .A2(o_label3_data4[27]), .A3(o_label3_data5[27]), .Z(n2032));
Q_MX02 U2458 ( .S(n4414), .A0(o_label3_data0[27]), .A1(o_label3_data1[27]), .Z(n2033));
Q_AN02 U2459 ( .A0(n4414), .A1(o_label4_config[11]), .Z(n2034));
Q_MX02 U2460 ( .S(n4415), .A0(n2034), .A1(n2033), .Z(n2035));
Q_MX04 U2461 ( .S0(n4416), .S1(n4417), .A0(n2035), .A1(n2032), .A2(n2031), .A3(n2030), .Z(n2036));
Q_MX02 U2462 ( .S(n4418), .A0(n2036), .A1(n2029), .Z(r32_mux_4_data[27]));
Q_MX03 U2463 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[12]), .A1(o_label0_data0[28]), .A2(o_label0_data1[28]), .Z(n2037));
Q_MX04 U2464 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[28]), .A1(o_label1_data5[28]), .A2(o_label1_data6[28]), .A3(o_label1_data7[28]), .Z(n2038));
Q_MX02 U2465 ( .S(n4416), .A0(n2038), .A1(n2037), .Z(n2039));
Q_MX08 U2466 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[28]), .A1(o_label2_data6[28]), .A2(o_label2_data7[28]), .A3(o_label2_config[12]), .A4(o_label1_data0[28]), .A5(o_label1_data1[28]), .A6(o_label1_data2[28]), .A7(o_label1_data3[28]), .Z(n2040));
Q_MX02 U2467 ( .S(n4417), .A0(n2040), .A1(n2039), .Z(n2041));
Q_MX04 U2468 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[28]), .A1(o_label2_data2[28]), .A2(o_label2_data3[28]), .A3(o_label2_data4[28]), .Z(n2042));
Q_MX04 U2469 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[28]), .A1(o_label3_data7[28]), .A2(o_label3_config[12]), .A3(o_label2_data0[28]), .Z(n2043));
Q_MX04 U2470 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[28]), .A1(o_label3_data3[28]), .A2(o_label3_data4[28]), .A3(o_label3_data5[28]), .Z(n2044));
Q_MX02 U2471 ( .S(n4414), .A0(o_label3_data0[28]), .A1(o_label3_data1[28]), .Z(n2045));
Q_AN02 U2472 ( .A0(n4414), .A1(o_label4_config[12]), .Z(n2046));
Q_MX02 U2473 ( .S(n4415), .A0(n2046), .A1(n2045), .Z(n2047));
Q_MX04 U2474 ( .S0(n4416), .S1(n4417), .A0(n2047), .A1(n2044), .A2(n2043), .A3(n2042), .Z(n2048));
Q_MX02 U2475 ( .S(n4418), .A0(n2048), .A1(n2041), .Z(r32_mux_4_data[28]));
Q_MX03 U2476 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[13]), .A1(o_label0_data0[29]), .A2(o_label0_data1[29]), .Z(n2049));
Q_MX04 U2477 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[29]), .A1(o_label1_data5[29]), .A2(o_label1_data6[29]), .A3(o_label1_data7[29]), .Z(n2050));
Q_MX02 U2478 ( .S(n4416), .A0(n2050), .A1(n2049), .Z(n2051));
Q_MX08 U2479 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[29]), .A1(o_label2_data6[29]), .A2(o_label2_data7[29]), .A3(o_label2_config[13]), .A4(o_label1_data0[29]), .A5(o_label1_data1[29]), .A6(o_label1_data2[29]), .A7(o_label1_data3[29]), .Z(n2052));
Q_MX02 U2480 ( .S(n4417), .A0(n2052), .A1(n2051), .Z(n2053));
Q_MX04 U2481 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[29]), .A1(o_label2_data2[29]), .A2(o_label2_data3[29]), .A3(o_label2_data4[29]), .Z(n2054));
Q_MX04 U2482 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[29]), .A1(o_label3_data7[29]), .A2(o_label3_config[13]), .A3(o_label2_data0[29]), .Z(n2055));
Q_MX04 U2483 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[29]), .A1(o_label3_data3[29]), .A2(o_label3_data4[29]), .A3(o_label3_data5[29]), .Z(n2056));
Q_MX02 U2484 ( .S(n4414), .A0(o_label3_data0[29]), .A1(o_label3_data1[29]), .Z(n2057));
Q_AN02 U2485 ( .A0(n4414), .A1(o_label4_config[13]), .Z(n2058));
Q_MX02 U2486 ( .S(n4415), .A0(n2058), .A1(n2057), .Z(n2059));
Q_MX04 U2487 ( .S0(n4416), .S1(n4417), .A0(n2059), .A1(n2056), .A2(n2055), .A3(n2054), .Z(n2060));
Q_MX02 U2488 ( .S(n4418), .A0(n2060), .A1(n2053), .Z(r32_mux_4_data[29]));
Q_MX03 U2489 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[14]), .A1(o_label0_data0[30]), .A2(o_label0_data1[30]), .Z(n2061));
Q_MX04 U2490 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[30]), .A1(o_label1_data5[30]), .A2(o_label1_data6[30]), .A3(o_label1_data7[30]), .Z(n2062));
Q_MX02 U2491 ( .S(n4416), .A0(n2062), .A1(n2061), .Z(n2063));
Q_MX08 U2492 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[30]), .A1(o_label2_data6[30]), .A2(o_label2_data7[30]), .A3(o_label2_config[14]), .A4(o_label1_data0[30]), .A5(o_label1_data1[30]), .A6(o_label1_data2[30]), .A7(o_label1_data3[30]), .Z(n2064));
Q_MX02 U2493 ( .S(n4417), .A0(n2064), .A1(n2063), .Z(n2065));
Q_MX04 U2494 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[30]), .A1(o_label2_data2[30]), .A2(o_label2_data3[30]), .A3(o_label2_data4[30]), .Z(n2066));
Q_MX04 U2495 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[30]), .A1(o_label3_data7[30]), .A2(o_label3_config[14]), .A3(o_label2_data0[30]), .Z(n2067));
Q_MX04 U2496 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[30]), .A1(o_label3_data3[30]), .A2(o_label3_data4[30]), .A3(o_label3_data5[30]), .Z(n2068));
Q_MX02 U2497 ( .S(n4414), .A0(o_label3_data0[30]), .A1(o_label3_data1[30]), .Z(n2069));
Q_AN02 U2498 ( .A0(n4414), .A1(o_label4_config[14]), .Z(n2070));
Q_MX02 U2499 ( .S(n4415), .A0(n2070), .A1(n2069), .Z(n2071));
Q_MX04 U2500 ( .S0(n4416), .S1(n4417), .A0(n2071), .A1(n2068), .A2(n2067), .A3(n2066), .Z(n2072));
Q_MX02 U2501 ( .S(n4418), .A0(n2072), .A1(n2065), .Z(r32_mux_4_data[30]));
Q_MX03 U2502 ( .S0(n4414), .S1(n4415), .A0(o_label1_config[15]), .A1(o_label0_data0[31]), .A2(o_label0_data1[31]), .Z(n2073));
Q_MX04 U2503 ( .S0(n4414), .S1(n4415), .A0(o_label1_data4[31]), .A1(o_label1_data5[31]), .A2(o_label1_data6[31]), .A3(o_label1_data7[31]), .Z(n2074));
Q_MX02 U2504 ( .S(n4416), .A0(n2074), .A1(n2073), .Z(n2075));
Q_MX08 U2505 ( .S0(n4414), .S1(n4415), .S2(n4416), .A0(o_label2_data5[31]), .A1(o_label2_data6[31]), .A2(o_label2_data7[31]), .A3(o_label2_config[15]), .A4(o_label1_data0[31]), .A5(o_label1_data1[31]), .A6(o_label1_data2[31]), .A7(o_label1_data3[31]), .Z(n2076));
Q_MX02 U2506 ( .S(n4417), .A0(n2076), .A1(n2075), .Z(n2077));
Q_MX04 U2507 ( .S0(n4414), .S1(n4415), .A0(o_label2_data1[31]), .A1(o_label2_data2[31]), .A2(o_label2_data3[31]), .A3(o_label2_data4[31]), .Z(n2078));
Q_MX04 U2508 ( .S0(n4414), .S1(n4415), .A0(o_label3_data6[31]), .A1(o_label3_data7[31]), .A2(o_label3_config[15]), .A3(o_label2_data0[31]), .Z(n2079));
Q_MX04 U2509 ( .S0(n4414), .S1(n4415), .A0(o_label3_data2[31]), .A1(o_label3_data3[31]), .A2(o_label3_data4[31]), .A3(o_label3_data5[31]), .Z(n2080));
Q_MX02 U2510 ( .S(n4414), .A0(o_label3_data0[31]), .A1(o_label3_data1[31]), .Z(n2081));
Q_AN02 U2511 ( .A0(n4414), .A1(o_label4_config[15]), .Z(n2082));
Q_MX02 U2512 ( .S(n4415), .A0(n2082), .A1(n2081), .Z(n2083));
Q_MX04 U2513 ( .S0(n4416), .S1(n4417), .A0(n2083), .A1(n2080), .A2(n2079), .A3(n2078), .Z(n2084));
Q_MX02 U2514 ( .S(n4418), .A0(n2084), .A1(n2077), .Z(r32_mux_4_data[31]));
Q_MX02 U2515 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[0]), .A1(o_cddip3_out_ia_wdata_part1[0]), .Z(n2085));
Q_MX04 U2516 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[0]), .A1(i_cddip3_out_ia_rdata_part1[0]), .A2(i_cddip3_out_ia_rdata_part0[0]), .A3(o_cddip3_out_ia_config[0]), .Z(n2086));
Q_MX02 U2517 ( .S(n4426), .A0(n2086), .A1(n2085), .Z(n2087));
Q_MX08 U2518 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[0]), .A1(o_ckv_ia_config[0]), .A2(o_ckv_ia_wdata_part1[0]), .A3(o_ckv_ia_wdata_part0[0]), .A4(i_ckv_ia_status[0]), .A5(i_ckv_ia_capability[0]), .A6(i_cddip3_out_im_status[0]), .A7(o_cddip3_out_im_config[0]), .Z(n2088));
Q_MX02 U2519 ( .S(n4427), .A0(n2088), .A1(n2087), .Z(n2089));
Q_MX04 U2520 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[0]), .A1(i_kim_ia_status[0]), .A2(i_kim_ia_capability[0]), .A3(i_ckv_ia_rdata_part1[0]), .Z(n2090));
Q_MX04 U2521 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[0]), .A1(i_kim_ia_rdata_part0[0]), .A2(o_kim_ia_config[0]), .A3(o_kim_ia_wdata_part1[0]), .Z(n2091));
Q_MX04 U2522 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[0]), .A1(o_label0_data6[0]), .A2(o_label0_data7[0]), .A3(o_label0_config[0]), .Z(n2092));
Q_MX02 U2523 ( .S(n4424), .A0(o_label0_data3[0]), .A1(o_label0_data4[0]), .Z(n2093));
Q_AN02 U2524 ( .A0(n4424), .A1(o_label0_data2[0]), .Z(n2094));
Q_MX02 U2525 ( .S(n4425), .A0(n2094), .A1(n2093), .Z(n2095));
Q_MX04 U2526 ( .S0(n4426), .S1(n4427), .A0(n2095), .A1(n2092), .A2(n2091), .A3(n2090), .Z(n2096));
Q_MX02 U2527 ( .S(n4428), .A0(n2096), .A1(n2089), .Z(r32_mux_3_data[0]));
Q_MX02 U2528 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[1]), .A1(o_cddip3_out_ia_wdata_part1[1]), .Z(n2097));
Q_MX04 U2529 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[1]), .A1(i_cddip3_out_ia_rdata_part1[1]), .A2(i_cddip3_out_ia_rdata_part0[1]), .A3(o_cddip3_out_ia_config[1]), .Z(n2098));
Q_MX02 U2530 ( .S(n4426), .A0(n2098), .A1(n2097), .Z(n2099));
Q_MX08 U2531 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[1]), .A1(o_ckv_ia_config[1]), .A2(o_ckv_ia_wdata_part1[1]), .A3(o_ckv_ia_wdata_part0[1]), .A4(i_ckv_ia_status[1]), .A5(i_ckv_ia_capability[1]), .A6(i_cddip3_out_im_status[1]), .A7(o_cddip3_out_im_config[1]), .Z(n2100));
Q_MX02 U2532 ( .S(n4427), .A0(n2100), .A1(n2099), .Z(n2101));
Q_MX04 U2533 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[1]), .A1(i_kim_ia_status[1]), .A2(i_kim_ia_capability[1]), .A3(i_ckv_ia_rdata_part1[1]), .Z(n2102));
Q_MX04 U2534 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[1]), .A1(i_kim_ia_rdata_part0[1]), .A2(o_kim_ia_config[1]), .A3(o_kim_ia_wdata_part1[1]), .Z(n2103));
Q_MX04 U2535 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[1]), .A1(o_label0_data6[1]), .A2(o_label0_data7[1]), .A3(o_label0_config[1]), .Z(n2104));
Q_MX02 U2536 ( .S(n4424), .A0(o_label0_data3[1]), .A1(o_label0_data4[1]), .Z(n2105));
Q_AN02 U2537 ( .A0(n4424), .A1(o_label0_data2[1]), .Z(n2106));
Q_MX02 U2538 ( .S(n4425), .A0(n2106), .A1(n2105), .Z(n2107));
Q_MX04 U2539 ( .S0(n4426), .S1(n4427), .A0(n2107), .A1(n2104), .A2(n2103), .A3(n2102), .Z(n2108));
Q_MX02 U2540 ( .S(n4428), .A0(n2108), .A1(n2101), .Z(r32_mux_3_data[1]));
Q_MX02 U2541 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[2]), .A1(o_cddip3_out_ia_wdata_part1[2]), .Z(n2109));
Q_MX04 U2542 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[2]), .A1(i_cddip3_out_ia_rdata_part1[2]), .A2(i_cddip3_out_ia_rdata_part0[2]), .A3(o_cddip3_out_ia_config[2]), .Z(n2110));
Q_MX02 U2543 ( .S(n4426), .A0(n2110), .A1(n2109), .Z(n2111));
Q_MX08 U2544 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[2]), .A1(o_ckv_ia_config[2]), .A2(o_ckv_ia_wdata_part1[2]), .A3(o_ckv_ia_wdata_part0[2]), .A4(i_ckv_ia_status[2]), .A5(i_ckv_ia_capability[2]), .A6(i_cddip3_out_im_status[2]), .A7(o_cddip3_out_im_config[2]), .Z(n2112));
Q_MX02 U2545 ( .S(n4427), .A0(n2112), .A1(n2111), .Z(n2113));
Q_MX04 U2546 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[2]), .A1(i_kim_ia_status[2]), .A2(i_kim_ia_capability[2]), .A3(i_ckv_ia_rdata_part1[2]), .Z(n2114));
Q_MX04 U2547 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[2]), .A1(i_kim_ia_rdata_part0[2]), .A2(o_kim_ia_config[2]), .A3(o_kim_ia_wdata_part1[2]), .Z(n2115));
Q_MX04 U2548 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[2]), .A1(o_label0_data6[2]), .A2(o_label0_data7[2]), .A3(o_label0_config[2]), .Z(n2116));
Q_MX02 U2549 ( .S(n4424), .A0(o_label0_data3[2]), .A1(o_label0_data4[2]), .Z(n2117));
Q_AN02 U2550 ( .A0(n4424), .A1(o_label0_data2[2]), .Z(n2118));
Q_MX02 U2551 ( .S(n4425), .A0(n2118), .A1(n2117), .Z(n2119));
Q_MX04 U2552 ( .S0(n4426), .S1(n4427), .A0(n2119), .A1(n2116), .A2(n2115), .A3(n2114), .Z(n2120));
Q_MX02 U2553 ( .S(n4428), .A0(n2120), .A1(n2113), .Z(r32_mux_3_data[2]));
Q_MX02 U2554 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[3]), .A1(o_cddip3_out_ia_wdata_part1[3]), .Z(n2121));
Q_MX04 U2555 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[3]), .A1(i_cddip3_out_ia_rdata_part1[3]), .A2(i_cddip3_out_ia_rdata_part0[3]), .A3(o_cddip3_out_ia_config[3]), .Z(n2122));
Q_MX02 U2556 ( .S(n4426), .A0(n2122), .A1(n2121), .Z(n2123));
Q_MX08 U2557 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[3]), .A1(o_ckv_ia_config[3]), .A2(o_ckv_ia_wdata_part1[3]), .A3(o_ckv_ia_wdata_part0[3]), .A4(i_ckv_ia_status[3]), .A5(i_ckv_ia_capability[3]), .A6(i_cddip3_out_im_status[3]), .A7(o_cddip3_out_im_config[3]), .Z(n2124));
Q_MX02 U2558 ( .S(n4427), .A0(n2124), .A1(n2123), .Z(n2125));
Q_MX04 U2559 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[3]), .A1(i_kim_ia_status[3]), .A2(i_kim_ia_capability[3]), .A3(i_ckv_ia_rdata_part1[3]), .Z(n2126));
Q_MX04 U2560 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[3]), .A1(i_kim_ia_rdata_part0[3]), .A2(o_kim_ia_config[3]), .A3(o_kim_ia_wdata_part1[3]), .Z(n2127));
Q_MX04 U2561 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[3]), .A1(o_label0_data6[3]), .A2(o_label0_data7[3]), .A3(o_label0_config[3]), .Z(n2128));
Q_MX02 U2562 ( .S(n4424), .A0(o_label0_data3[3]), .A1(o_label0_data4[3]), .Z(n2129));
Q_AN02 U2563 ( .A0(n4424), .A1(o_label0_data2[3]), .Z(n2130));
Q_MX02 U2564 ( .S(n4425), .A0(n2130), .A1(n2129), .Z(n2131));
Q_MX04 U2565 ( .S0(n4426), .S1(n4427), .A0(n2131), .A1(n2128), .A2(n2127), .A3(n2126), .Z(n2132));
Q_MX02 U2566 ( .S(n4428), .A0(n2132), .A1(n2125), .Z(r32_mux_3_data[3]));
Q_MX02 U2567 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[4]), .A1(o_cddip3_out_ia_wdata_part1[4]), .Z(n2133));
Q_MX04 U2568 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[4]), .A1(i_cddip3_out_ia_rdata_part1[4]), .A2(i_cddip3_out_ia_rdata_part0[4]), .A3(o_cddip3_out_ia_config[4]), .Z(n2134));
Q_MX02 U2569 ( .S(n4426), .A0(n2134), .A1(n2133), .Z(n2135));
Q_MX08 U2570 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[4]), .A1(o_ckv_ia_config[4]), .A2(o_ckv_ia_wdata_part1[4]), .A3(o_ckv_ia_wdata_part0[4]), .A4(i_ckv_ia_status[4]), .A5(i_ckv_ia_capability[4]), .A6(i_cddip3_out_im_status[4]), .A7(o_cddip3_out_im_config[4]), .Z(n2136));
Q_MX02 U2571 ( .S(n4427), .A0(n2136), .A1(n2135), .Z(n2137));
Q_MX04 U2572 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[4]), .A1(i_kim_ia_status[4]), .A2(i_kim_ia_capability[4]), .A3(i_ckv_ia_rdata_part1[4]), .Z(n2138));
Q_MX04 U2573 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[4]), .A1(i_kim_ia_rdata_part0[4]), .A2(o_kim_ia_config[4]), .A3(o_kim_ia_wdata_part1[4]), .Z(n2139));
Q_MX04 U2574 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[4]), .A1(o_label0_data6[4]), .A2(o_label0_data7[4]), .A3(o_label0_config[4]), .Z(n2140));
Q_MX02 U2575 ( .S(n4424), .A0(o_label0_data3[4]), .A1(o_label0_data4[4]), .Z(n2141));
Q_AN02 U2576 ( .A0(n4424), .A1(o_label0_data2[4]), .Z(n2142));
Q_MX02 U2577 ( .S(n4425), .A0(n2142), .A1(n2141), .Z(n2143));
Q_MX04 U2578 ( .S0(n4426), .S1(n4427), .A0(n2143), .A1(n2140), .A2(n2139), .A3(n2138), .Z(n2144));
Q_MX02 U2579 ( .S(n4428), .A0(n2144), .A1(n2137), .Z(r32_mux_3_data[4]));
Q_MX02 U2580 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[5]), .A1(o_cddip3_out_ia_wdata_part1[5]), .Z(n2145));
Q_MX04 U2581 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[5]), .A1(i_cddip3_out_ia_rdata_part1[5]), .A2(i_cddip3_out_ia_rdata_part0[5]), .A3(o_cddip3_out_ia_config[5]), .Z(n2146));
Q_MX02 U2582 ( .S(n4426), .A0(n2146), .A1(n2145), .Z(n2147));
Q_MX08 U2583 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[5]), .A1(o_ckv_ia_config[5]), .A2(o_ckv_ia_wdata_part1[5]), .A3(o_ckv_ia_wdata_part0[5]), .A4(i_ckv_ia_status[5]), .A5(i_ckv_ia_capability[5]), .A6(i_cddip3_out_im_status[5]), .A7(o_cddip3_out_im_config[5]), .Z(n2148));
Q_MX02 U2584 ( .S(n4427), .A0(n2148), .A1(n2147), .Z(n2149));
Q_MX04 U2585 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[5]), .A1(i_kim_ia_status[5]), .A2(i_kim_ia_capability[5]), .A3(i_ckv_ia_rdata_part1[5]), .Z(n2150));
Q_MX04 U2586 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[5]), .A1(i_kim_ia_rdata_part0[5]), .A2(o_kim_ia_config[5]), .A3(o_kim_ia_wdata_part1[5]), .Z(n2151));
Q_MX04 U2587 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[5]), .A1(o_label0_data6[5]), .A2(o_label0_data7[5]), .A3(o_label0_config[5]), .Z(n2152));
Q_MX02 U2588 ( .S(n4424), .A0(o_label0_data3[5]), .A1(o_label0_data4[5]), .Z(n2153));
Q_AN02 U2589 ( .A0(n4424), .A1(o_label0_data2[5]), .Z(n2154));
Q_MX02 U2590 ( .S(n4425), .A0(n2154), .A1(n2153), .Z(n2155));
Q_MX04 U2591 ( .S0(n4426), .S1(n4427), .A0(n2155), .A1(n2152), .A2(n2151), .A3(n2150), .Z(n2156));
Q_MX02 U2592 ( .S(n4428), .A0(n2156), .A1(n2149), .Z(r32_mux_3_data[5]));
Q_MX02 U2593 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[6]), .A1(o_cddip3_out_ia_wdata_part1[6]), .Z(n2157));
Q_MX04 U2594 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[6]), .A1(i_cddip3_out_ia_rdata_part1[6]), .A2(i_cddip3_out_ia_rdata_part0[6]), .A3(o_cddip3_out_ia_config[6]), .Z(n2158));
Q_MX02 U2595 ( .S(n4426), .A0(n2158), .A1(n2157), .Z(n2159));
Q_MX08 U2596 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[6]), .A1(o_ckv_ia_config[6]), .A2(o_ckv_ia_wdata_part1[6]), .A3(o_ckv_ia_wdata_part0[6]), .A4(i_ckv_ia_status[6]), .A5(i_ckv_ia_capability[6]), .A6(i_cddip3_out_im_status[6]), .A7(o_cddip3_out_im_config[6]), .Z(n2160));
Q_MX02 U2597 ( .S(n4427), .A0(n2160), .A1(n2159), .Z(n2161));
Q_MX04 U2598 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[6]), .A1(i_kim_ia_status[6]), .A2(i_kim_ia_capability[6]), .A3(i_ckv_ia_rdata_part1[6]), .Z(n2162));
Q_MX04 U2599 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[6]), .A1(i_kim_ia_rdata_part0[6]), .A2(o_kim_ia_config[6]), .A3(o_kim_ia_wdata_part1[6]), .Z(n2163));
Q_MX04 U2600 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[6]), .A1(o_label0_data6[6]), .A2(o_label0_data7[6]), .A3(o_label0_config[6]), .Z(n2164));
Q_MX02 U2601 ( .S(n4424), .A0(o_label0_data3[6]), .A1(o_label0_data4[6]), .Z(n2165));
Q_AN02 U2602 ( .A0(n4424), .A1(o_label0_data2[6]), .Z(n2166));
Q_MX02 U2603 ( .S(n4425), .A0(n2166), .A1(n2165), .Z(n2167));
Q_MX04 U2604 ( .S0(n4426), .S1(n4427), .A0(n2167), .A1(n2164), .A2(n2163), .A3(n2162), .Z(n2168));
Q_MX02 U2605 ( .S(n4428), .A0(n2168), .A1(n2161), .Z(r32_mux_3_data[6]));
Q_MX02 U2606 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[7]), .A1(o_cddip3_out_ia_wdata_part1[7]), .Z(n2169));
Q_MX04 U2607 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[7]), .A1(i_cddip3_out_ia_rdata_part1[7]), .A2(i_cddip3_out_ia_rdata_part0[7]), .A3(o_cddip3_out_ia_config[7]), .Z(n2170));
Q_MX02 U2608 ( .S(n4426), .A0(n2170), .A1(n2169), .Z(n2171));
Q_MX08 U2609 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[7]), .A1(o_ckv_ia_config[7]), .A2(o_ckv_ia_wdata_part1[7]), .A3(o_ckv_ia_wdata_part0[7]), .A4(i_ckv_ia_status[7]), .A5(i_ckv_ia_capability[7]), .A6(i_cddip3_out_im_status[7]), .A7(o_cddip3_out_im_config[7]), .Z(n2172));
Q_MX02 U2610 ( .S(n4427), .A0(n2172), .A1(n2171), .Z(n2173));
Q_MX04 U2611 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[7]), .A1(i_kim_ia_status[7]), .A2(i_kim_ia_capability[7]), .A3(i_ckv_ia_rdata_part1[7]), .Z(n2174));
Q_MX04 U2612 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[7]), .A1(i_kim_ia_rdata_part0[7]), .A2(o_kim_ia_config[7]), .A3(o_kim_ia_wdata_part1[7]), .Z(n2175));
Q_MX04 U2613 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[7]), .A1(o_label0_data6[7]), .A2(o_label0_data7[7]), .A3(o_label0_config[7]), .Z(n2176));
Q_MX02 U2614 ( .S(n4424), .A0(o_label0_data3[7]), .A1(o_label0_data4[7]), .Z(n2177));
Q_AN02 U2615 ( .A0(n4424), .A1(o_label0_data2[7]), .Z(n2178));
Q_MX02 U2616 ( .S(n4425), .A0(n2178), .A1(n2177), .Z(n2179));
Q_MX04 U2617 ( .S0(n4426), .S1(n4427), .A0(n2179), .A1(n2176), .A2(n2175), .A3(n2174), .Z(n2180));
Q_MX02 U2618 ( .S(n4428), .A0(n2180), .A1(n2173), .Z(r32_mux_3_data[7]));
Q_MX02 U2619 ( .S(n4424), .A0(o_cddip3_out_ia_wdata_part2[8]), .A1(o_cddip3_out_ia_wdata_part1[8]), .Z(n2181));
Q_MX04 U2620 ( .S0(n4424), .S1(n4425), .A0(i_cddip3_out_ia_rdata_part2[8]), .A1(i_cddip3_out_ia_rdata_part1[8]), .A2(i_cddip3_out_ia_rdata_part0[8]), .A3(o_cddip3_out_ia_config[8]), .Z(n2182));
Q_MX02 U2621 ( .S(n4426), .A0(n2182), .A1(n2181), .Z(n2183));
Q_MX08 U2622 ( .S0(n4424), .S1(n4425), .S2(n4426), .A0(i_ckv_ia_rdata_part0[8]), .A1(o_ckv_ia_config[8]), .A2(o_ckv_ia_wdata_part1[8]), .A3(o_ckv_ia_wdata_part0[8]), .A4(i_ckv_ia_status[8]), .A5(i_ckv_ia_capability[8]), .A6(i_cddip3_out_im_status[8]), .A7(o_cddip3_out_im_config[8]), .Z(n2184));
Q_MX02 U2623 ( .S(n4427), .A0(n2184), .A1(n2183), .Z(n2185));
Q_MX04 U2624 ( .S0(n4424), .S1(n4425), .A0(o_kim_ia_wdata_part0[8]), .A1(i_kim_ia_status[8]), .A2(i_kim_ia_capability[8]), .A3(i_ckv_ia_rdata_part1[8]), .Z(n2186));
Q_MX04 U2625 ( .S0(n4424), .S1(n4425), .A0(i_kim_ia_rdata_part1[8]), .A1(i_kim_ia_rdata_part0[8]), .A2(o_kim_ia_config[8]), .A3(o_kim_ia_wdata_part1[8]), .Z(n2187));
Q_MX04 U2626 ( .S0(n4424), .S1(n4425), .A0(o_label0_data5[8]), .A1(o_label0_data6[8]), .A2(o_label0_data7[8]), .A3(o_label0_config[8]), .Z(n2188));
Q_MX02 U2627 ( .S(n4424), .A0(o_label0_data3[8]), .A1(o_label0_data4[8]), .Z(n2189));
Q_AN02 U2628 ( .A0(n4424), .A1(o_label0_data2[8]), .Z(n2190));
Q_MX02 U2629 ( .S(n4425), .A0(n2190), .A1(n2189), .Z(n2191));
Q_MX04 U2630 ( .S0(n4426), .S1(n4427), .A0(n2191), .A1(n2188), .A2(n2187), .A3(n2186), .Z(n2192));
Q_MX02 U2631 ( .S(n4428), .A0(n2192), .A1(n2185), .Z(r32_mux_3_data[8]));
Q_MX03 U2632 ( .S0(n4429), .S1(n4430), .A0(i_cddip3_out_ia_rdata_part0[9]), .A1(o_cddip3_out_ia_wdata_part2[9]), .A2(o_cddip3_out_ia_wdata_part1[9]), .Z(n2193));
Q_MX08 U2633 ( .S0(n4429), .S1(n4430), .S2(n4431), .A0(o_ckv_ia_config[9]), .A1(o_ckv_ia_wdata_part1[9]), .A2(o_ckv_ia_wdata_part0[9]), .A3(i_ckv_ia_status[9]), .A4(i_ckv_ia_capability[9]), .A5(o_cddip3_out_im_config[9]), .A6(i_cddip3_out_ia_rdata_part2[9]), .A7(i_cddip3_out_ia_rdata_part1[9]), .Z(n2194));
Q_MX02 U2634 ( .S(n4432), .A0(n2194), .A1(n2193), .Z(n2195));
Q_MX04 U2635 ( .S0(n4429), .S1(n4430), .A0(i_kim_ia_status[9]), .A1(i_kim_ia_capability[9]), .A2(i_ckv_ia_rdata_part1[9]), .A3(i_ckv_ia_rdata_part0[9]), .Z(n2196));
Q_MX04 U2636 ( .S0(n4429), .S1(n4430), .A0(i_kim_ia_rdata_part0[9]), .A1(o_kim_ia_config[9]), .A2(o_kim_ia_wdata_part1[9]), .A3(o_kim_ia_wdata_part0[9]), .Z(n2197));
Q_MX04 U2637 ( .S0(n4429), .S1(n4430), .A0(o_label0_data5[9]), .A1(o_label0_data6[9]), .A2(o_label0_data7[9]), .A3(i_kim_ia_rdata_part1[9]), .Z(n2198));
Q_MX02 U2638 ( .S(n4429), .A0(o_label0_data3[9]), .A1(o_label0_data4[9]), .Z(n2199));
Q_AN02 U2639 ( .A0(n4429), .A1(o_label0_data2[9]), .Z(n2200));
Q_MX02 U2640 ( .S(n4430), .A0(n2200), .A1(n2199), .Z(n2201));
Q_MX04 U2641 ( .S0(n4431), .S1(n4432), .A0(n2201), .A1(n2198), .A2(n2197), .A3(n2196), .Z(n2202));
Q_MX02 U2642 ( .S(n4433), .A0(n2202), .A1(n2195), .Z(r32_mux_3_data[9]));
Q_MX02 U2643 ( .S(n4434), .A0(o_cddip3_out_ia_wdata_part2[10]), .A1(o_cddip3_out_ia_wdata_part1[10]), .Z(n2203));
Q_MX08 U2644 ( .S0(n4434), .S1(n4435), .S2(n4436), .A0(o_ckv_ia_config[10]), .A1(o_ckv_ia_wdata_part1[10]), .A2(o_ckv_ia_wdata_part0[10]), .A3(i_ckv_ia_status[10]), .A4(i_ckv_ia_capability[10]), .A5(i_cddip3_out_ia_rdata_part2[10]), .A6(i_cddip3_out_ia_rdata_part1[10]), .A7(i_cddip3_out_ia_rdata_part0[10]), .Z(n2204));
Q_MX02 U2645 ( .S(n4437), .A0(n2204), .A1(n2203), .Z(n2205));
Q_MX04 U2646 ( .S0(n4434), .S1(n4435), .A0(i_kim_ia_status[10]), .A1(i_kim_ia_capability[10]), .A2(i_ckv_ia_rdata_part1[10]), .A3(i_ckv_ia_rdata_part0[10]), .Z(n2206));
Q_MX04 U2647 ( .S0(n4434), .S1(n4435), .A0(i_kim_ia_rdata_part0[10]), .A1(o_kim_ia_config[10]), .A2(o_kim_ia_wdata_part1[10]), .A3(o_kim_ia_wdata_part0[10]), .Z(n2207));
Q_MX04 U2648 ( .S0(n4434), .S1(n4435), .A0(o_label0_data5[10]), .A1(o_label0_data6[10]), .A2(o_label0_data7[10]), .A3(i_kim_ia_rdata_part1[10]), .Z(n2208));
Q_MX02 U2649 ( .S(n4434), .A0(o_label0_data3[10]), .A1(o_label0_data4[10]), .Z(n2209));
Q_AN02 U2650 ( .A0(n4434), .A1(o_label0_data2[10]), .Z(n2210));
Q_MX02 U2651 ( .S(n4435), .A0(n2210), .A1(n2209), .Z(n2211));
Q_MX04 U2652 ( .S0(n4436), .S1(n4437), .A0(n2211), .A1(n2208), .A2(n2207), .A3(n2206), .Z(n2212));
Q_MX02 U2653 ( .S(n4438), .A0(n2212), .A1(n2205), .Z(r32_mux_3_data[10]));
Q_MX02 U2654 ( .S(n4434), .A0(o_cddip3_out_ia_wdata_part2[11]), .A1(o_cddip3_out_ia_wdata_part1[11]), .Z(n2213));
Q_MX08 U2655 ( .S0(n4434), .S1(n4435), .S2(n4436), .A0(o_ckv_ia_config[11]), .A1(o_ckv_ia_wdata_part1[11]), .A2(o_ckv_ia_wdata_part0[11]), .A3(i_ckv_ia_status[11]), .A4(i_ckv_ia_capability[11]), .A5(i_cddip3_out_ia_rdata_part2[11]), .A6(i_cddip3_out_ia_rdata_part1[11]), .A7(i_cddip3_out_ia_rdata_part0[11]), .Z(n2214));
Q_MX02 U2656 ( .S(n4437), .A0(n2214), .A1(n2213), .Z(n2215));
Q_MX04 U2657 ( .S0(n4434), .S1(n4435), .A0(i_kim_ia_status[11]), .A1(i_kim_ia_capability[11]), .A2(i_ckv_ia_rdata_part1[11]), .A3(i_ckv_ia_rdata_part0[11]), .Z(n2216));
Q_MX04 U2658 ( .S0(n4434), .S1(n4435), .A0(i_kim_ia_rdata_part0[11]), .A1(o_kim_ia_config[11]), .A2(o_kim_ia_wdata_part1[11]), .A3(o_kim_ia_wdata_part0[11]), .Z(n2217));
Q_MX04 U2659 ( .S0(n4434), .S1(n4435), .A0(o_label0_data5[11]), .A1(o_label0_data6[11]), .A2(o_label0_data7[11]), .A3(i_kim_ia_rdata_part1[11]), .Z(n2218));
Q_MX02 U2660 ( .S(n4434), .A0(o_label0_data3[11]), .A1(o_label0_data4[11]), .Z(n2219));
Q_AN02 U2661 ( .A0(n4434), .A1(o_label0_data2[11]), .Z(n2220));
Q_MX02 U2662 ( .S(n4435), .A0(n2220), .A1(n2219), .Z(n2221));
Q_MX04 U2663 ( .S0(n4436), .S1(n4437), .A0(n2221), .A1(n2218), .A2(n2217), .A3(n2216), .Z(n2222));
Q_MX02 U2664 ( .S(n4438), .A0(n2222), .A1(n2215), .Z(r32_mux_3_data[11]));
Q_MX02 U2665 ( .S(n4434), .A0(o_cddip3_out_ia_wdata_part2[12]), .A1(o_cddip3_out_ia_wdata_part1[12]), .Z(n2223));
Q_MX08 U2666 ( .S0(n4434), .S1(n4435), .S2(n4436), .A0(o_ckv_ia_config[12]), .A1(o_ckv_ia_wdata_part1[12]), .A2(o_ckv_ia_wdata_part0[12]), .A3(i_ckv_ia_status[12]), .A4(i_ckv_ia_capability[12]), .A5(i_cddip3_out_ia_rdata_part2[12]), .A6(i_cddip3_out_ia_rdata_part1[12]), .A7(i_cddip3_out_ia_rdata_part0[12]), .Z(n2224));
Q_MX02 U2667 ( .S(n4437), .A0(n2224), .A1(n2223), .Z(n2225));
Q_MX04 U2668 ( .S0(n4434), .S1(n4435), .A0(i_kim_ia_status[12]), .A1(i_kim_ia_capability[12]), .A2(i_ckv_ia_rdata_part1[12]), .A3(i_ckv_ia_rdata_part0[12]), .Z(n2226));
Q_MX04 U2669 ( .S0(n4434), .S1(n4435), .A0(i_kim_ia_rdata_part0[12]), .A1(o_kim_ia_config[12]), .A2(o_kim_ia_wdata_part1[12]), .A3(o_kim_ia_wdata_part0[12]), .Z(n2227));
Q_MX04 U2670 ( .S0(n4434), .S1(n4435), .A0(o_label0_data5[12]), .A1(o_label0_data6[12]), .A2(o_label0_data7[12]), .A3(i_kim_ia_rdata_part1[12]), .Z(n2228));
Q_MX02 U2671 ( .S(n4434), .A0(o_label0_data3[12]), .A1(o_label0_data4[12]), .Z(n2229));
Q_AN02 U2672 ( .A0(n4434), .A1(o_label0_data2[12]), .Z(n2230));
Q_MX02 U2673 ( .S(n4435), .A0(n2230), .A1(n2229), .Z(n2231));
Q_MX04 U2674 ( .S0(n4436), .S1(n4437), .A0(n2231), .A1(n2228), .A2(n2227), .A3(n2226), .Z(n2232));
Q_MX02 U2675 ( .S(n4438), .A0(n2232), .A1(n2225), .Z(r32_mux_3_data[12]));
Q_MX08 U2676 ( .S0(n4439), .S1(n4440), .S2(n4441), .A0(o_ckv_ia_wdata_part0[13]), .A1(i_ckv_ia_status[13]), .A2(i_ckv_ia_capability[13]), .A3(i_cddip3_out_ia_rdata_part2[13]), .A4(i_cddip3_out_ia_rdata_part1[13]), .A5(i_cddip3_out_ia_rdata_part0[13]), .A6(o_cddip3_out_ia_wdata_part2[13]), .A7(o_cddip3_out_ia_wdata_part1[13]), .Z(n2233));
Q_MX04 U2677 ( .S0(n4439), .S1(n4440), .A0(i_ckv_ia_rdata_part1[13]), .A1(i_ckv_ia_rdata_part0[13]), .A2(o_ckv_ia_config[13]), .A3(o_ckv_ia_wdata_part1[13]), .Z(n2234));
Q_MX04 U2678 ( .S0(n4439), .S1(n4440), .A0(o_kim_ia_config[13]), .A1(o_kim_ia_wdata_part0[13]), .A2(i_kim_ia_status[13]), .A3(i_kim_ia_capability[13]), .Z(n2235));
Q_MX04 U2679 ( .S0(n4439), .S1(n4440), .A0(o_label0_data5[13]), .A1(o_label0_data6[13]), .A2(o_label0_data7[13]), .A3(i_kim_ia_rdata_part0[13]), .Z(n2236));
Q_MX02 U2680 ( .S(n4439), .A0(o_label0_data3[13]), .A1(o_label0_data4[13]), .Z(n2237));
Q_AN02 U2681 ( .A0(n4439), .A1(o_label0_data2[13]), .Z(n2238));
Q_MX02 U2682 ( .S(n4440), .A0(n2238), .A1(n2237), .Z(n2239));
Q_MX04 U2683 ( .S0(n4441), .S1(n4442), .A0(n2239), .A1(n2236), .A2(n2235), .A3(n2234), .Z(n2240));
Q_MX02 U2684 ( .S(n4443), .A0(n2240), .A1(n2233), .Z(r32_mux_3_data[13]));
Q_MX02 U2685 ( .S(n4444), .A0(o_cddip3_out_ia_wdata_part2[14]), .A1(o_cddip3_out_ia_wdata_part1[14]), .Z(n2241));
Q_MX04 U2686 ( .S0(n4444), .S1(n4445), .A0(i_ckv_ia_capability[14]), .A1(i_cddip3_out_ia_rdata_part2[14]), .A2(i_cddip3_out_ia_rdata_part1[14]), .A3(i_cddip3_out_ia_rdata_part0[14]), .Z(n2242));
Q_MX02 U2687 ( .S(n4446), .A0(n2242), .A1(n2241), .Z(n2243));
Q_MX04 U2688 ( .S0(n4444), .S1(n4445), .A0(o_ckv_ia_config[14]), .A1(o_ckv_ia_wdata_part1[14]), .A2(o_ckv_ia_wdata_part0[14]), .A3(i_ckv_ia_status[14]), .Z(n2244));
Q_MX04 U2689 ( .S0(n4444), .S1(n4445), .A0(o_kim_ia_wdata_part0[14]), .A1(i_kim_ia_capability[14]), .A2(i_ckv_ia_rdata_part1[14]), .A3(i_ckv_ia_rdata_part0[14]), .Z(n2245));
Q_MX04 U2690 ( .S0(n4444), .S1(n4445), .A0(o_label0_data5[14]), .A1(o_label0_data6[14]), .A2(o_label0_data7[14]), .A3(i_kim_ia_rdata_part0[14]), .Z(n2246));
Q_MX02 U2691 ( .S(n4444), .A0(o_label0_data3[14]), .A1(o_label0_data4[14]), .Z(n2247));
Q_AN02 U2692 ( .A0(n4444), .A1(o_label0_data2[14]), .Z(n2248));
Q_MX02 U2693 ( .S(n4445), .A0(n2248), .A1(n2247), .Z(n2249));
Q_MX04 U2694 ( .S0(n4446), .S1(n4447), .A0(n2249), .A1(n2246), .A2(n2245), .A3(n2244), .Z(n2250));
Q_MX02 U2695 ( .S(n4448), .A0(n2250), .A1(n2243), .Z(r32_mux_3_data[14]));
Q_MX02 U2696 ( .S(n4449), .A0(o_cddip3_out_ia_wdata_part2[15]), .A1(o_cddip3_out_ia_wdata_part1[15]), .Z(n2251));
Q_MX04 U2697 ( .S0(n4449), .S1(n4450), .A0(i_ckv_ia_capability[15]), .A1(i_cddip3_out_ia_rdata_part2[15]), .A2(i_cddip3_out_ia_rdata_part1[15]), .A3(i_cddip3_out_ia_rdata_part0[15]), .Z(n2252));
Q_MX04 U2698 ( .S0(n4449), .S1(n4450), .A0(i_ckv_ia_rdata_part1[15]), .A1(i_ckv_ia_rdata_part0[15]), .A2(o_ckv_ia_wdata_part1[15]), .A3(o_ckv_ia_wdata_part0[15]), .Z(n2253));
Q_MX04 U2699 ( .S0(n4449), .S1(n4450), .A0(o_label0_data5[15]), .A1(o_label0_data6[15]), .A2(o_label0_data7[15]), .A3(i_kim_ia_capability[15]), .Z(n2254));
Q_MX02 U2700 ( .S(n4449), .A0(o_label0_data3[15]), .A1(o_label0_data4[15]), .Z(n2255));
Q_AN02 U2701 ( .A0(n4449), .A1(o_label0_data2[15]), .Z(n2256));
Q_MX02 U2702 ( .S(n4450), .A0(n2256), .A1(n2255), .Z(n2257));
Q_MX04 U2703 ( .S0(n4451), .S1(n4452), .A0(n2257), .A1(n2254), .A2(n2253), .A3(n2252), .Z(n2258));
Q_MX02 U2704 ( .S(n4453), .A0(n2258), .A1(n2251), .Z(r32_mux_3_data[15]));
Q_MX04 U2705 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[16]), .A1(i_cddip3_out_ia_rdata_part0[16]), .A2(o_cddip3_out_ia_wdata_part2[16]), .A3(o_cddip3_out_ia_wdata_part1[16]), .Z(n2259));
Q_MX04 U2706 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[16]), .A1(o_ckv_ia_wdata_part1[16]), .A2(o_ckv_ia_wdata_part0[16]), .A3(i_cddip3_out_ia_rdata_part2[16]), .Z(n2260));
Q_MX04 U2707 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[16]), .A1(o_label0_data6[16]), .A2(o_label0_data7[16]), .A3(i_ckv_ia_rdata_part1[16]), .Z(n2261));
Q_MX02 U2708 ( .S(n4454), .A0(o_label0_data3[16]), .A1(o_label0_data4[16]), .Z(n2262));
Q_AN02 U2709 ( .A0(n4454), .A1(o_label0_data2[16]), .Z(n2263));
Q_MX02 U2710 ( .S(n4455), .A0(n2263), .A1(n2262), .Z(n2264));
Q_MX04 U2711 ( .S0(n4456), .S1(n4457), .A0(n2264), .A1(n2261), .A2(n2260), .A3(n2259), .Z(r32_mux_3_data[16]));
Q_MX04 U2712 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[17]), .A1(i_cddip3_out_ia_rdata_part0[17]), .A2(o_cddip3_out_ia_wdata_part2[17]), .A3(o_cddip3_out_ia_wdata_part1[17]), .Z(n2265));
Q_MX04 U2713 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[17]), .A1(o_ckv_ia_wdata_part1[17]), .A2(o_ckv_ia_wdata_part0[17]), .A3(i_cddip3_out_ia_rdata_part2[17]), .Z(n2266));
Q_MX04 U2714 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[17]), .A1(o_label0_data6[17]), .A2(o_label0_data7[17]), .A3(i_ckv_ia_rdata_part1[17]), .Z(n2267));
Q_MX02 U2715 ( .S(n4454), .A0(o_label0_data3[17]), .A1(o_label0_data4[17]), .Z(n2268));
Q_AN02 U2716 ( .A0(n4454), .A1(o_label0_data2[17]), .Z(n2269));
Q_MX02 U2717 ( .S(n4455), .A0(n2269), .A1(n2268), .Z(n2270));
Q_MX04 U2718 ( .S0(n4456), .S1(n4457), .A0(n2270), .A1(n2267), .A2(n2266), .A3(n2265), .Z(r32_mux_3_data[17]));
Q_MX04 U2719 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[18]), .A1(i_cddip3_out_ia_rdata_part0[18]), .A2(o_cddip3_out_ia_wdata_part2[18]), .A3(o_cddip3_out_ia_wdata_part1[18]), .Z(n2271));
Q_MX04 U2720 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[18]), .A1(o_ckv_ia_wdata_part1[18]), .A2(o_ckv_ia_wdata_part0[18]), .A3(i_cddip3_out_ia_rdata_part2[18]), .Z(n2272));
Q_MX04 U2721 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[18]), .A1(o_label0_data6[18]), .A2(o_label0_data7[18]), .A3(i_ckv_ia_rdata_part1[18]), .Z(n2273));
Q_MX02 U2722 ( .S(n4454), .A0(o_label0_data3[18]), .A1(o_label0_data4[18]), .Z(n2274));
Q_AN02 U2723 ( .A0(n4454), .A1(o_label0_data2[18]), .Z(n2275));
Q_MX02 U2724 ( .S(n4455), .A0(n2275), .A1(n2274), .Z(n2276));
Q_MX04 U2725 ( .S0(n4456), .S1(n4457), .A0(n2276), .A1(n2273), .A2(n2272), .A3(n2271), .Z(r32_mux_3_data[18]));
Q_MX04 U2726 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[19]), .A1(i_cddip3_out_ia_rdata_part0[19]), .A2(o_cddip3_out_ia_wdata_part2[19]), .A3(o_cddip3_out_ia_wdata_part1[19]), .Z(n2277));
Q_MX04 U2727 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[19]), .A1(o_ckv_ia_wdata_part1[19]), .A2(o_ckv_ia_wdata_part0[19]), .A3(i_cddip3_out_ia_rdata_part2[19]), .Z(n2278));
Q_MX04 U2728 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[19]), .A1(o_label0_data6[19]), .A2(o_label0_data7[19]), .A3(i_ckv_ia_rdata_part1[19]), .Z(n2279));
Q_MX02 U2729 ( .S(n4454), .A0(o_label0_data3[19]), .A1(o_label0_data4[19]), .Z(n2280));
Q_AN02 U2730 ( .A0(n4454), .A1(o_label0_data2[19]), .Z(n2281));
Q_MX02 U2731 ( .S(n4455), .A0(n2281), .A1(n2280), .Z(n2282));
Q_MX04 U2732 ( .S0(n4456), .S1(n4457), .A0(n2282), .A1(n2279), .A2(n2278), .A3(n2277), .Z(r32_mux_3_data[19]));
Q_MX04 U2733 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[20]), .A1(i_cddip3_out_ia_rdata_part0[20]), .A2(o_cddip3_out_ia_wdata_part2[20]), .A3(o_cddip3_out_ia_wdata_part1[20]), .Z(n2283));
Q_MX04 U2734 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[20]), .A1(o_ckv_ia_wdata_part1[20]), .A2(o_ckv_ia_wdata_part0[20]), .A3(i_cddip3_out_ia_rdata_part2[20]), .Z(n2284));
Q_MX04 U2735 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[20]), .A1(o_label0_data6[20]), .A2(o_label0_data7[20]), .A3(i_ckv_ia_rdata_part1[20]), .Z(n2285));
Q_MX02 U2736 ( .S(n4454), .A0(o_label0_data3[20]), .A1(o_label0_data4[20]), .Z(n2286));
Q_AN02 U2737 ( .A0(n4454), .A1(o_label0_data2[20]), .Z(n2287));
Q_MX02 U2738 ( .S(n4455), .A0(n2287), .A1(n2286), .Z(n2288));
Q_MX04 U2739 ( .S0(n4456), .S1(n4457), .A0(n2288), .A1(n2285), .A2(n2284), .A3(n2283), .Z(r32_mux_3_data[20]));
Q_MX04 U2740 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[21]), .A1(i_cddip3_out_ia_rdata_part0[21]), .A2(o_cddip3_out_ia_wdata_part2[21]), .A3(o_cddip3_out_ia_wdata_part1[21]), .Z(n2289));
Q_MX04 U2741 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[21]), .A1(o_ckv_ia_wdata_part1[21]), .A2(o_ckv_ia_wdata_part0[21]), .A3(i_cddip3_out_ia_rdata_part2[21]), .Z(n2290));
Q_MX04 U2742 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[21]), .A1(o_label0_data6[21]), .A2(o_label0_data7[21]), .A3(i_ckv_ia_rdata_part1[21]), .Z(n2291));
Q_MX02 U2743 ( .S(n4454), .A0(o_label0_data3[21]), .A1(o_label0_data4[21]), .Z(n2292));
Q_AN02 U2744 ( .A0(n4454), .A1(o_label0_data2[21]), .Z(n2293));
Q_MX02 U2745 ( .S(n4455), .A0(n2293), .A1(n2292), .Z(n2294));
Q_MX04 U2746 ( .S0(n4456), .S1(n4457), .A0(n2294), .A1(n2291), .A2(n2290), .A3(n2289), .Z(r32_mux_3_data[21]));
Q_MX04 U2747 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[22]), .A1(i_cddip3_out_ia_rdata_part0[22]), .A2(o_cddip3_out_ia_wdata_part2[22]), .A3(o_cddip3_out_ia_wdata_part1[22]), .Z(n2295));
Q_MX04 U2748 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[22]), .A1(o_ckv_ia_wdata_part1[22]), .A2(o_ckv_ia_wdata_part0[22]), .A3(i_cddip3_out_ia_rdata_part2[22]), .Z(n2296));
Q_MX04 U2749 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[22]), .A1(o_label0_data6[22]), .A2(o_label0_data7[22]), .A3(i_ckv_ia_rdata_part1[22]), .Z(n2297));
Q_MX02 U2750 ( .S(n4454), .A0(o_label0_data3[22]), .A1(o_label0_data4[22]), .Z(n2298));
Q_AN02 U2751 ( .A0(n4454), .A1(o_label0_data2[22]), .Z(n2299));
Q_MX02 U2752 ( .S(n4455), .A0(n2299), .A1(n2298), .Z(n2300));
Q_MX04 U2753 ( .S0(n4456), .S1(n4457), .A0(n2300), .A1(n2297), .A2(n2296), .A3(n2295), .Z(r32_mux_3_data[22]));
Q_MX04 U2754 ( .S0(n4454), .S1(n4455), .A0(i_cddip3_out_ia_rdata_part1[23]), .A1(i_cddip3_out_ia_rdata_part0[23]), .A2(o_cddip3_out_ia_wdata_part2[23]), .A3(o_cddip3_out_ia_wdata_part1[23]), .Z(n2301));
Q_MX04 U2755 ( .S0(n4454), .S1(n4455), .A0(i_ckv_ia_rdata_part0[23]), .A1(o_ckv_ia_wdata_part1[23]), .A2(o_ckv_ia_wdata_part0[23]), .A3(i_cddip3_out_ia_rdata_part2[23]), .Z(n2302));
Q_MX04 U2756 ( .S0(n4454), .S1(n4455), .A0(o_label0_data5[23]), .A1(o_label0_data6[23]), .A2(o_label0_data7[23]), .A3(i_ckv_ia_rdata_part1[23]), .Z(n2303));
Q_MX02 U2757 ( .S(n4454), .A0(o_label0_data3[23]), .A1(o_label0_data4[23]), .Z(n2304));
Q_AN02 U2758 ( .A0(n4454), .A1(o_label0_data2[23]), .Z(n2305));
Q_MX02 U2759 ( .S(n4455), .A0(n2305), .A1(n2304), .Z(n2306));
Q_MX04 U2760 ( .S0(n4456), .S1(n4457), .A0(n2306), .A1(n2303), .A2(n2302), .A3(n2301), .Z(r32_mux_3_data[23]));
Q_MX02 U2761 ( .S(n4458), .A0(o_cddip3_out_ia_wdata_part2[24]), .A1(o_cddip3_out_ia_wdata_part1[24]), .Z(n2307));
Q_MX04 U2762 ( .S0(n4458), .S1(n4459), .A0(i_ckv_ia_status[15]), .A1(i_cddip3_out_ia_rdata_part2[24]), .A2(i_cddip3_out_ia_rdata_part1[24]), .A3(i_cddip3_out_ia_rdata_part0[24]), .Z(n2308));
Q_MX04 U2763 ( .S0(n4458), .S1(n4459), .A0(i_ckv_ia_rdata_part1[24]), .A1(i_ckv_ia_rdata_part0[24]), .A2(o_ckv_ia_wdata_part1[24]), .A3(o_ckv_ia_wdata_part0[24]), .Z(n2309));
Q_MX04 U2764 ( .S0(n4458), .S1(n4459), .A0(o_label0_data5[24]), .A1(o_label0_data6[24]), .A2(o_label0_data7[24]), .A3(i_kim_ia_status[14]), .Z(n2310));
Q_MX02 U2765 ( .S(n4458), .A0(o_label0_data3[24]), .A1(o_label0_data4[24]), .Z(n2311));
Q_AN02 U2766 ( .A0(n4458), .A1(o_label0_data2[24]), .Z(n2312));
Q_MX02 U2767 ( .S(n4459), .A0(n2312), .A1(n2311), .Z(n2313));
Q_MX04 U2768 ( .S0(n4460), .S1(n4461), .A0(n2313), .A1(n2310), .A2(n2309), .A3(n2308), .Z(n2314));
Q_MX02 U2769 ( .S(n4453), .A0(n2314), .A1(n2307), .Z(r32_mux_3_data[24]));
Q_MX03 U2770 ( .S0(n4462), .S1(n4463), .A0(i_cddip3_out_ia_rdata_part0[25]), .A1(o_cddip3_out_ia_wdata_part2[25]), .A2(o_cddip3_out_ia_wdata_part1[25]), .Z(n2315));
Q_MX04 U2771 ( .S0(n4462), .S1(n4463), .A0(o_ckv_ia_wdata_part0[25]), .A1(i_ckv_ia_status[16]), .A2(i_cddip3_out_ia_rdata_part2[25]), .A3(i_cddip3_out_ia_rdata_part1[25]), .Z(n2316));
Q_MX04 U2772 ( .S0(n4462), .S1(n4463), .A0(i_kim_ia_status[15]), .A1(i_ckv_ia_rdata_part1[25]), .A2(i_ckv_ia_rdata_part0[25]), .A3(o_ckv_ia_wdata_part1[25]), .Z(n2317));
Q_MX04 U2773 ( .S0(n4462), .S1(n4463), .A0(o_label0_data5[25]), .A1(o_label0_data6[25]), .A2(o_label0_data7[25]), .A3(o_label0_config[9]), .Z(n2318));
Q_MX02 U2774 ( .S(n4462), .A0(o_label0_data3[25]), .A1(o_label0_data4[25]), .Z(n2319));
Q_AN02 U2775 ( .A0(n4462), .A1(o_label0_data2[25]), .Z(n2320));
Q_MX02 U2776 ( .S(n4463), .A0(n2320), .A1(n2319), .Z(n2321));
Q_MX04 U2777 ( .S0(n4464), .S1(n4465), .A0(n2321), .A1(n2318), .A2(n2317), .A3(n2316), .Z(n2322));
Q_MX02 U2778 ( .S(n4466), .A0(n2322), .A1(n2315), .Z(r32_mux_3_data[25]));
Q_MX04 U2779 ( .S0(n4467), .S1(n4468), .A0(i_cddip3_out_ia_rdata_part2[26]), .A1(i_cddip3_out_ia_rdata_part1[26]), .A2(i_cddip3_out_ia_rdata_part0[26]), .A3(o_cddip3_out_ia_wdata_part2[26]), .Z(n2323));
Q_MX02 U2780 ( .S(n4469), .A0(n2323), .A1(o_cddip3_out_ia_wdata_part1[26]), .Z(n2324));
Q_MX04 U2781 ( .S0(n4467), .S1(n4468), .A0(i_ckv_ia_rdata_part0[26]), .A1(o_ckv_ia_wdata_part1[26]), .A2(o_ckv_ia_wdata_part0[26]), .A3(i_ckv_ia_status[17]), .Z(n2325));
Q_MX04 U2782 ( .S0(n4467), .S1(n4468), .A0(i_kim_ia_rdata_part0[15]), .A1(o_kim_ia_wdata_part0[15]), .A2(i_kim_ia_status[16]), .A3(i_ckv_ia_rdata_part1[26]), .Z(n2326));
Q_MX04 U2783 ( .S0(n4467), .S1(n4468), .A0(o_label0_data5[26]), .A1(o_label0_data6[26]), .A2(o_label0_data7[26]), .A3(o_label0_config[10]), .Z(n2327));
Q_MX02 U2784 ( .S(n4467), .A0(o_label0_data3[26]), .A1(o_label0_data4[26]), .Z(n2328));
Q_AN02 U2785 ( .A0(n4467), .A1(o_label0_data2[26]), .Z(n2329));
Q_MX02 U2786 ( .S(n4468), .A0(n2329), .A1(n2328), .Z(n2330));
Q_MX04 U2787 ( .S0(n4469), .S1(n4470), .A0(n2330), .A1(n2327), .A2(n2326), .A3(n2325), .Z(n2331));
Q_MX02 U2788 ( .S(n4471), .A0(n2331), .A1(n2324), .Z(r32_mux_3_data[26]));
Q_MX04 U2789 ( .S0(n4467), .S1(n4468), .A0(i_cddip3_out_ia_rdata_part2[27]), .A1(i_cddip3_out_ia_rdata_part1[27]), .A2(i_cddip3_out_ia_rdata_part0[27]), .A3(o_cddip3_out_ia_wdata_part2[27]), .Z(n2332));
Q_MX02 U2790 ( .S(n4469), .A0(n2332), .A1(o_cddip3_out_ia_wdata_part1[27]), .Z(n2333));
Q_MX04 U2791 ( .S0(n4467), .S1(n4468), .A0(i_ckv_ia_rdata_part0[27]), .A1(o_ckv_ia_wdata_part1[27]), .A2(o_ckv_ia_wdata_part0[27]), .A3(i_ckv_ia_status[18]), .Z(n2334));
Q_MX04 U2792 ( .S0(n4467), .S1(n4468), .A0(i_kim_ia_rdata_part0[16]), .A1(o_kim_ia_wdata_part0[16]), .A2(i_kim_ia_status[17]), .A3(i_ckv_ia_rdata_part1[27]), .Z(n2335));
Q_MX04 U2793 ( .S0(n4467), .S1(n4468), .A0(o_label0_data5[27]), .A1(o_label0_data6[27]), .A2(o_label0_data7[27]), .A3(o_label0_config[11]), .Z(n2336));
Q_MX02 U2794 ( .S(n4467), .A0(o_label0_data3[27]), .A1(o_label0_data4[27]), .Z(n2337));
Q_AN02 U2795 ( .A0(n4467), .A1(o_label0_data2[27]), .Z(n2338));
Q_MX02 U2796 ( .S(n4468), .A0(n2338), .A1(n2337), .Z(n2339));
Q_MX04 U2797 ( .S0(n4469), .S1(n4470), .A0(n2339), .A1(n2336), .A2(n2335), .A3(n2334), .Z(n2340));
Q_MX02 U2798 ( .S(n4471), .A0(n2340), .A1(n2333), .Z(r32_mux_3_data[27]));
Q_MX04 U2799 ( .S0(n4472), .S1(n4473), .A0(i_cddip3_out_ia_rdata_part0[28]), .A1(o_cddip3_out_ia_config[9]), .A2(o_cddip3_out_ia_wdata_part2[28]), .A3(o_cddip3_out_ia_wdata_part1[28]), .Z(n2341));
Q_MX08 U2800 ( .S0(n4472), .S1(n4473), .S2(n4474), .A0(i_ckv_ia_rdata_part0[28]), .A1(o_ckv_ia_config[15]), .A2(o_ckv_ia_wdata_part1[28]), .A3(o_ckv_ia_wdata_part0[28]), .A4(i_ckv_ia_status[19]), .A5(i_ckv_ia_capability[16]), .A6(i_cddip3_out_ia_rdata_part2[28]), .A7(i_cddip3_out_ia_rdata_part1[28]), .Z(n2342));
Q_MX02 U2801 ( .S(n4475), .A0(n2342), .A1(n2341), .Z(n2343));
Q_MX04 U2802 ( .S0(n4472), .S1(n4473), .A0(o_kim_ia_wdata_part0[17]), .A1(i_kim_ia_status[18]), .A2(i_kim_ia_capability[16]), .A3(i_ckv_ia_rdata_part1[28]), .Z(n2344));
Q_MX04 U2803 ( .S0(n4472), .S1(n4473), .A0(i_kim_ia_rdata_part1[13]), .A1(i_kim_ia_rdata_part0[17]), .A2(o_kim_ia_config[14]), .A3(o_kim_ia_wdata_part1[13]), .Z(n2345));
Q_MX04 U2804 ( .S0(n4472), .S1(n4473), .A0(o_label0_data5[28]), .A1(o_label0_data6[28]), .A2(o_label0_data7[28]), .A3(o_label0_config[12]), .Z(n2346));
Q_MX02 U2805 ( .S(n4472), .A0(o_label0_data3[28]), .A1(o_label0_data4[28]), .Z(n2347));
Q_AN02 U2806 ( .A0(n4472), .A1(o_label0_data2[28]), .Z(n2348));
Q_MX02 U2807 ( .S(n4473), .A0(n2348), .A1(n2347), .Z(n2349));
Q_MX04 U2808 ( .S0(n4474), .S1(n4475), .A0(n2349), .A1(n2346), .A2(n2345), .A3(n2344), .Z(n2350));
Q_MX02 U2809 ( .S(n4476), .A0(n2350), .A1(n2343), .Z(r32_mux_3_data[28]));
Q_MX04 U2810 ( .S0(n4477), .S1(n4478), .A0(i_cddip3_out_ia_rdata_part1[29]), .A1(i_cddip3_out_ia_rdata_part0[29]), .A2(o_cddip3_out_ia_config[10]), .A3(o_cddip3_out_ia_wdata_part2[29]), .Z(n2351));
Q_MX02 U2811 ( .S(n4479), .A0(n2351), .A1(o_cddip3_out_ia_wdata_part1[29]), .Z(n2352));
Q_MX08 U2812 ( .S0(n4477), .S1(n4478), .S2(n4479), .A0(i_ckv_ia_rdata_part0[29]), .A1(o_ckv_ia_config[16]), .A2(o_ckv_ia_wdata_part1[29]), .A3(o_ckv_ia_wdata_part0[29]), .A4(i_ckv_ia_status[20]), .A5(i_ckv_ia_capability[17]), .A6(i_cddip3_out_im_status[9]), .A7(i_cddip3_out_ia_rdata_part2[29]), .Z(n2353));
Q_MX02 U2813 ( .S(n4480), .A0(n2353), .A1(n2352), .Z(n2354));
Q_MX04 U2814 ( .S0(n4477), .S1(n4478), .A0(o_kim_ia_wdata_part0[18]), .A1(i_kim_ia_status[19]), .A2(i_kim_ia_capability[17]), .A3(i_ckv_ia_rdata_part1[29]), .Z(n2355));
Q_MX04 U2815 ( .S0(n4477), .S1(n4478), .A0(i_kim_ia_rdata_part1[14]), .A1(i_kim_ia_rdata_part0[18]), .A2(o_kim_ia_config[15]), .A3(o_kim_ia_wdata_part1[14]), .Z(n2356));
Q_MX04 U2816 ( .S0(n4477), .S1(n4478), .A0(o_label0_data5[29]), .A1(o_label0_data6[29]), .A2(o_label0_data7[29]), .A3(o_label0_config[13]), .Z(n2357));
Q_MX02 U2817 ( .S(n4477), .A0(o_label0_data3[29]), .A1(o_label0_data4[29]), .Z(n2358));
Q_AN02 U2818 ( .A0(n4477), .A1(o_label0_data2[29]), .Z(n2359));
Q_MX02 U2819 ( .S(n4478), .A0(n2359), .A1(n2358), .Z(n2360));
Q_MX04 U2820 ( .S0(n4479), .S1(n4480), .A0(n2360), .A1(n2357), .A2(n2356), .A3(n2355), .Z(n2361));
Q_MX02 U2821 ( .S(n4481), .A0(n2361), .A1(n2354), .Z(r32_mux_3_data[29]));
Q_MX03 U2822 ( .S0(n4482), .S1(n4483), .A0(o_cddip3_out_ia_config[11]), .A1(o_cddip3_out_ia_wdata_part2[30]), .A2(o_cddip3_out_ia_wdata_part1[30]), .Z(n2362));
Q_MX04 U2823 ( .S0(n4482), .S1(n4483), .A0(o_cddip3_out_im_config[10]), .A1(i_cddip3_out_ia_rdata_part2[30]), .A2(i_cddip3_out_ia_rdata_part1[30]), .A3(i_cddip3_out_ia_rdata_part0[30]), .Z(n2363));
Q_MX02 U2824 ( .S(n4484), .A0(n2363), .A1(n2362), .Z(n2364));
Q_MX08 U2825 ( .S0(n4482), .S1(n4483), .S2(n4484), .A0(i_ckv_ia_rdata_part0[30]), .A1(o_ckv_ia_config[17]), .A2(o_ckv_ia_wdata_part1[30]), .A3(o_ckv_ia_wdata_part0[30]), .A4(i_ckv_ia_status[21]), .A5(i_ckv_ia_capability[18]), .A6(i_cddip3_out_im_read_done[0]), .A7(i_cddip3_out_im_status[10]), .Z(n2365));
Q_MX02 U2826 ( .S(n4485), .A0(n2365), .A1(n2364), .Z(n2366));
Q_MX04 U2827 ( .S0(n4482), .S1(n4483), .A0(o_kim_ia_wdata_part0[19]), .A1(i_kim_ia_status[20]), .A2(i_kim_ia_capability[18]), .A3(i_ckv_ia_rdata_part1[30]), .Z(n2367));
Q_MX04 U2828 ( .S0(n4482), .S1(n4483), .A0(i_kim_ia_rdata_part1[15]), .A1(i_kim_ia_rdata_part0[19]), .A2(o_kim_ia_config[16]), .A3(o_kim_ia_wdata_part1[15]), .Z(n2368));
Q_MX04 U2829 ( .S0(n4482), .S1(n4483), .A0(o_label0_data5[30]), .A1(o_label0_data6[30]), .A2(o_label0_data7[30]), .A3(o_label0_config[14]), .Z(n2369));
Q_MX02 U2830 ( .S(n4482), .A0(o_label0_data3[30]), .A1(o_label0_data4[30]), .Z(n2370));
Q_AN02 U2831 ( .A0(n4482), .A1(o_label0_data2[30]), .Z(n2371));
Q_MX02 U2832 ( .S(n4483), .A0(n2371), .A1(n2370), .Z(n2372));
Q_MX04 U2833 ( .S0(n4484), .S1(n4485), .A0(n2372), .A1(n2369), .A2(n2368), .A3(n2367), .Z(n2373));
Q_MX02 U2834 ( .S(n4486), .A0(n2373), .A1(n2366), .Z(r32_mux_3_data[30]));
Q_MX03 U2835 ( .S0(n4482), .S1(n4483), .A0(o_cddip3_out_ia_config[12]), .A1(o_cddip3_out_ia_wdata_part2[31]), .A2(o_cddip3_out_ia_wdata_part1[31]), .Z(n2374));
Q_MX04 U2836 ( .S0(n4482), .S1(n4483), .A0(o_cddip3_out_im_config[11]), .A1(i_cddip3_out_ia_rdata_part2[31]), .A2(i_cddip3_out_ia_rdata_part1[31]), .A3(i_cddip3_out_ia_rdata_part0[31]), .Z(n2375));
Q_MX02 U2837 ( .S(n4484), .A0(n2375), .A1(n2374), .Z(n2376));
Q_MX08 U2838 ( .S0(n4482), .S1(n4483), .S2(n4484), .A0(i_ckv_ia_rdata_part0[31]), .A1(o_ckv_ia_config[18]), .A2(o_ckv_ia_wdata_part1[31]), .A3(o_ckv_ia_wdata_part0[31]), .A4(i_ckv_ia_status[22]), .A5(i_ckv_ia_capability[19]), .A6(i_cddip3_out_im_read_done[1]), .A7(i_cddip3_out_im_status[11]), .Z(n2377));
Q_MX02 U2839 ( .S(n4485), .A0(n2377), .A1(n2376), .Z(n2378));
Q_MX04 U2840 ( .S0(n4482), .S1(n4483), .A0(o_kim_ia_wdata_part0[20]), .A1(i_kim_ia_status[21]), .A2(i_kim_ia_capability[19]), .A3(i_ckv_ia_rdata_part1[31]), .Z(n2379));
Q_MX04 U2841 ( .S0(n4482), .S1(n4483), .A0(i_kim_ia_rdata_part1[16]), .A1(i_kim_ia_rdata_part0[20]), .A2(o_kim_ia_config[17]), .A3(o_kim_ia_wdata_part1[16]), .Z(n2380));
Q_MX04 U2842 ( .S0(n4482), .S1(n4483), .A0(o_label0_data5[31]), .A1(o_label0_data6[31]), .A2(o_label0_data7[31]), .A3(o_label0_config[15]), .Z(n2381));
Q_MX02 U2843 ( .S(n4482), .A0(o_label0_data3[31]), .A1(o_label0_data4[31]), .Z(n2382));
Q_AN02 U2844 ( .A0(n4482), .A1(o_label0_data2[31]), .Z(n2383));
Q_MX02 U2845 ( .S(n4483), .A0(n2383), .A1(n2382), .Z(n2384));
Q_MX04 U2846 ( .S0(n4484), .S1(n4485), .A0(n2384), .A1(n2381), .A2(n2380), .A3(n2379), .Z(n2385));
Q_MX02 U2847 ( .S(n4486), .A0(n2385), .A1(n2378), .Z(r32_mux_3_data[31]));
Q_MX04 U2848 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[0]), .A1(i_cddip1_out_ia_capability[0]), .A2(i_cddip0_out_im_status[0]), .A3(o_cddip0_out_im_config[0]), .Z(n2386));
Q_MX08 U2849 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[0]), .A1(i_cddip1_out_ia_rdata_part2[0]), .A2(i_cddip1_out_ia_rdata_part1[0]), .A3(i_cddip1_out_ia_rdata_part0[0]), .A4(o_cddip1_out_ia_config[0]), .A5(o_cddip1_out_ia_wdata_part2[0]), .A6(o_cddip1_out_ia_wdata_part1[0]), .A7(o_cddip1_out_ia_wdata_part0[0]), .Z(n2387));
Q_MX02 U2850 ( .S(n4490), .A0(n2387), .A1(n2386), .Z(n2388));
Q_MX04 U2851 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[0]), .A1(i_cddip2_out_ia_status[0]), .A2(i_cddip2_out_ia_capability[0]), .A3(i_cddip1_out_im_status[0]), .Z(n2389));
Q_MX04 U2852 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[0]), .A1(o_cddip2_out_ia_config[0]), .A2(o_cddip2_out_ia_wdata_part2[0]), .A3(o_cddip2_out_ia_wdata_part1[0]), .Z(n2390));
Q_MX04 U2853 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[0]), .A1(o_cddip2_out_im_config[0]), .A2(i_cddip2_out_ia_rdata_part2[0]), .A3(i_cddip2_out_ia_rdata_part1[0]), .Z(n2391));
Q_MX02 U2854 ( .S(n4487), .A0(i_cddip3_out_ia_status[0]), .A1(i_cddip3_out_ia_capability[0]), .Z(n2392));
Q_AN02 U2855 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[0]), .Z(n2393));
Q_MX02 U2856 ( .S(n4488), .A0(n2393), .A1(n2392), .Z(n2394));
Q_MX04 U2857 ( .S0(n4489), .S1(n4490), .A0(n2394), .A1(n2391), .A2(n2390), .A3(n2389), .Z(n2395));
Q_MX02 U2858 ( .S(n4491), .A0(n2395), .A1(n2388), .Z(r32_mux_2_data[0]));
Q_MX04 U2859 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[1]), .A1(i_cddip1_out_ia_capability[1]), .A2(i_cddip0_out_im_status[1]), .A3(o_cddip0_out_im_config[1]), .Z(n2396));
Q_MX08 U2860 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[1]), .A1(i_cddip1_out_ia_rdata_part2[1]), .A2(i_cddip1_out_ia_rdata_part1[1]), .A3(i_cddip1_out_ia_rdata_part0[1]), .A4(o_cddip1_out_ia_config[1]), .A5(o_cddip1_out_ia_wdata_part2[1]), .A6(o_cddip1_out_ia_wdata_part1[1]), .A7(o_cddip1_out_ia_wdata_part0[1]), .Z(n2397));
Q_MX02 U2861 ( .S(n4490), .A0(n2397), .A1(n2396), .Z(n2398));
Q_MX04 U2862 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[1]), .A1(i_cddip2_out_ia_status[1]), .A2(i_cddip2_out_ia_capability[1]), .A3(i_cddip1_out_im_status[1]), .Z(n2399));
Q_MX04 U2863 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[1]), .A1(o_cddip2_out_ia_config[1]), .A2(o_cddip2_out_ia_wdata_part2[1]), .A3(o_cddip2_out_ia_wdata_part1[1]), .Z(n2400));
Q_MX04 U2864 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[1]), .A1(o_cddip2_out_im_config[1]), .A2(i_cddip2_out_ia_rdata_part2[1]), .A3(i_cddip2_out_ia_rdata_part1[1]), .Z(n2401));
Q_MX02 U2865 ( .S(n4487), .A0(i_cddip3_out_ia_status[1]), .A1(i_cddip3_out_ia_capability[1]), .Z(n2402));
Q_AN02 U2866 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[1]), .Z(n2403));
Q_MX02 U2867 ( .S(n4488), .A0(n2403), .A1(n2402), .Z(n2404));
Q_MX04 U2868 ( .S0(n4489), .S1(n4490), .A0(n2404), .A1(n2401), .A2(n2400), .A3(n2399), .Z(n2405));
Q_MX02 U2869 ( .S(n4491), .A0(n2405), .A1(n2398), .Z(r32_mux_2_data[1]));
Q_MX04 U2870 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[2]), .A1(i_cddip1_out_ia_capability[2]), .A2(i_cddip0_out_im_status[2]), .A3(o_cddip0_out_im_config[2]), .Z(n2406));
Q_MX08 U2871 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[2]), .A1(i_cddip1_out_ia_rdata_part2[2]), .A2(i_cddip1_out_ia_rdata_part1[2]), .A3(i_cddip1_out_ia_rdata_part0[2]), .A4(o_cddip1_out_ia_config[2]), .A5(o_cddip1_out_ia_wdata_part2[2]), .A6(o_cddip1_out_ia_wdata_part1[2]), .A7(o_cddip1_out_ia_wdata_part0[2]), .Z(n2407));
Q_MX02 U2872 ( .S(n4490), .A0(n2407), .A1(n2406), .Z(n2408));
Q_MX04 U2873 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[2]), .A1(i_cddip2_out_ia_status[2]), .A2(i_cddip2_out_ia_capability[2]), .A3(i_cddip1_out_im_status[2]), .Z(n2409));
Q_MX04 U2874 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[2]), .A1(o_cddip2_out_ia_config[2]), .A2(o_cddip2_out_ia_wdata_part2[2]), .A3(o_cddip2_out_ia_wdata_part1[2]), .Z(n2410));
Q_MX04 U2875 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[2]), .A1(o_cddip2_out_im_config[2]), .A2(i_cddip2_out_ia_rdata_part2[2]), .A3(i_cddip2_out_ia_rdata_part1[2]), .Z(n2411));
Q_MX02 U2876 ( .S(n4487), .A0(i_cddip3_out_ia_status[2]), .A1(i_cddip3_out_ia_capability[2]), .Z(n2412));
Q_AN02 U2877 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[2]), .Z(n2413));
Q_MX02 U2878 ( .S(n4488), .A0(n2413), .A1(n2412), .Z(n2414));
Q_MX04 U2879 ( .S0(n4489), .S1(n4490), .A0(n2414), .A1(n2411), .A2(n2410), .A3(n2409), .Z(n2415));
Q_MX02 U2880 ( .S(n4491), .A0(n2415), .A1(n2408), .Z(r32_mux_2_data[2]));
Q_MX04 U2881 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[3]), .A1(i_cddip1_out_ia_capability[3]), .A2(i_cddip0_out_im_status[3]), .A3(o_cddip0_out_im_config[3]), .Z(n2416));
Q_MX08 U2882 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[3]), .A1(i_cddip1_out_ia_rdata_part2[3]), .A2(i_cddip1_out_ia_rdata_part1[3]), .A3(i_cddip1_out_ia_rdata_part0[3]), .A4(o_cddip1_out_ia_config[3]), .A5(o_cddip1_out_ia_wdata_part2[3]), .A6(o_cddip1_out_ia_wdata_part1[3]), .A7(o_cddip1_out_ia_wdata_part0[3]), .Z(n2417));
Q_MX02 U2883 ( .S(n4490), .A0(n2417), .A1(n2416), .Z(n2418));
Q_MX04 U2884 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[3]), .A1(i_cddip2_out_ia_status[3]), .A2(i_cddip2_out_ia_capability[3]), .A3(i_cddip1_out_im_status[3]), .Z(n2419));
Q_MX04 U2885 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[3]), .A1(o_cddip2_out_ia_config[3]), .A2(o_cddip2_out_ia_wdata_part2[3]), .A3(o_cddip2_out_ia_wdata_part1[3]), .Z(n2420));
Q_MX04 U2886 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[3]), .A1(o_cddip2_out_im_config[3]), .A2(i_cddip2_out_ia_rdata_part2[3]), .A3(i_cddip2_out_ia_rdata_part1[3]), .Z(n2421));
Q_MX02 U2887 ( .S(n4487), .A0(i_cddip3_out_ia_status[3]), .A1(i_cddip3_out_ia_capability[3]), .Z(n2422));
Q_AN02 U2888 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[3]), .Z(n2423));
Q_MX02 U2889 ( .S(n4488), .A0(n2423), .A1(n2422), .Z(n2424));
Q_MX04 U2890 ( .S0(n4489), .S1(n4490), .A0(n2424), .A1(n2421), .A2(n2420), .A3(n2419), .Z(n2425));
Q_MX02 U2891 ( .S(n4491), .A0(n2425), .A1(n2418), .Z(r32_mux_2_data[3]));
Q_MX04 U2892 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[4]), .A1(i_cddip1_out_ia_capability[4]), .A2(i_cddip0_out_im_status[4]), .A3(o_cddip0_out_im_config[4]), .Z(n2426));
Q_MX08 U2893 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[4]), .A1(i_cddip1_out_ia_rdata_part2[4]), .A2(i_cddip1_out_ia_rdata_part1[4]), .A3(i_cddip1_out_ia_rdata_part0[4]), .A4(o_cddip1_out_ia_config[4]), .A5(o_cddip1_out_ia_wdata_part2[4]), .A6(o_cddip1_out_ia_wdata_part1[4]), .A7(o_cddip1_out_ia_wdata_part0[4]), .Z(n2427));
Q_MX02 U2894 ( .S(n4490), .A0(n2427), .A1(n2426), .Z(n2428));
Q_MX04 U2895 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[4]), .A1(i_cddip2_out_ia_status[4]), .A2(i_cddip2_out_ia_capability[4]), .A3(i_cddip1_out_im_status[4]), .Z(n2429));
Q_MX04 U2896 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[4]), .A1(o_cddip2_out_ia_config[4]), .A2(o_cddip2_out_ia_wdata_part2[4]), .A3(o_cddip2_out_ia_wdata_part1[4]), .Z(n2430));
Q_MX04 U2897 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[4]), .A1(o_cddip2_out_im_config[4]), .A2(i_cddip2_out_ia_rdata_part2[4]), .A3(i_cddip2_out_ia_rdata_part1[4]), .Z(n2431));
Q_MX02 U2898 ( .S(n4487), .A0(i_cddip3_out_ia_status[4]), .A1(i_cddip3_out_ia_capability[4]), .Z(n2432));
Q_AN02 U2899 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[4]), .Z(n2433));
Q_MX02 U2900 ( .S(n4488), .A0(n2433), .A1(n2432), .Z(n2434));
Q_MX04 U2901 ( .S0(n4489), .S1(n4490), .A0(n2434), .A1(n2431), .A2(n2430), .A3(n2429), .Z(n2435));
Q_MX02 U2902 ( .S(n4491), .A0(n2435), .A1(n2428), .Z(r32_mux_2_data[4]));
Q_MX04 U2903 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[5]), .A1(i_cddip1_out_ia_capability[5]), .A2(i_cddip0_out_im_status[5]), .A3(o_cddip0_out_im_config[5]), .Z(n2436));
Q_MX08 U2904 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[5]), .A1(i_cddip1_out_ia_rdata_part2[5]), .A2(i_cddip1_out_ia_rdata_part1[5]), .A3(i_cddip1_out_ia_rdata_part0[5]), .A4(o_cddip1_out_ia_config[5]), .A5(o_cddip1_out_ia_wdata_part2[5]), .A6(o_cddip1_out_ia_wdata_part1[5]), .A7(o_cddip1_out_ia_wdata_part0[5]), .Z(n2437));
Q_MX02 U2905 ( .S(n4490), .A0(n2437), .A1(n2436), .Z(n2438));
Q_MX04 U2906 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[5]), .A1(i_cddip2_out_ia_status[5]), .A2(i_cddip2_out_ia_capability[5]), .A3(i_cddip1_out_im_status[5]), .Z(n2439));
Q_MX04 U2907 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[5]), .A1(o_cddip2_out_ia_config[5]), .A2(o_cddip2_out_ia_wdata_part2[5]), .A3(o_cddip2_out_ia_wdata_part1[5]), .Z(n2440));
Q_MX04 U2908 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[5]), .A1(o_cddip2_out_im_config[5]), .A2(i_cddip2_out_ia_rdata_part2[5]), .A3(i_cddip2_out_ia_rdata_part1[5]), .Z(n2441));
Q_MX02 U2909 ( .S(n4487), .A0(i_cddip3_out_ia_status[5]), .A1(i_cddip3_out_ia_capability[5]), .Z(n2442));
Q_AN02 U2910 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[5]), .Z(n2443));
Q_MX02 U2911 ( .S(n4488), .A0(n2443), .A1(n2442), .Z(n2444));
Q_MX04 U2912 ( .S0(n4489), .S1(n4490), .A0(n2444), .A1(n2441), .A2(n2440), .A3(n2439), .Z(n2445));
Q_MX02 U2913 ( .S(n4491), .A0(n2445), .A1(n2438), .Z(r32_mux_2_data[5]));
Q_MX04 U2914 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[6]), .A1(i_cddip1_out_ia_capability[6]), .A2(i_cddip0_out_im_status[6]), .A3(o_cddip0_out_im_config[6]), .Z(n2446));
Q_MX08 U2915 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[6]), .A1(i_cddip1_out_ia_rdata_part2[6]), .A2(i_cddip1_out_ia_rdata_part1[6]), .A3(i_cddip1_out_ia_rdata_part0[6]), .A4(o_cddip1_out_ia_config[6]), .A5(o_cddip1_out_ia_wdata_part2[6]), .A6(o_cddip1_out_ia_wdata_part1[6]), .A7(o_cddip1_out_ia_wdata_part0[6]), .Z(n2447));
Q_MX02 U2916 ( .S(n4490), .A0(n2447), .A1(n2446), .Z(n2448));
Q_MX04 U2917 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[6]), .A1(i_cddip2_out_ia_status[6]), .A2(i_cddip2_out_ia_capability[6]), .A3(i_cddip1_out_im_status[6]), .Z(n2449));
Q_MX04 U2918 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[6]), .A1(o_cddip2_out_ia_config[6]), .A2(o_cddip2_out_ia_wdata_part2[6]), .A3(o_cddip2_out_ia_wdata_part1[6]), .Z(n2450));
Q_MX04 U2919 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[6]), .A1(o_cddip2_out_im_config[6]), .A2(i_cddip2_out_ia_rdata_part2[6]), .A3(i_cddip2_out_ia_rdata_part1[6]), .Z(n2451));
Q_MX02 U2920 ( .S(n4487), .A0(i_cddip3_out_ia_status[6]), .A1(i_cddip3_out_ia_capability[6]), .Z(n2452));
Q_AN02 U2921 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[6]), .Z(n2453));
Q_MX02 U2922 ( .S(n4488), .A0(n2453), .A1(n2452), .Z(n2454));
Q_MX04 U2923 ( .S0(n4489), .S1(n4490), .A0(n2454), .A1(n2451), .A2(n2450), .A3(n2449), .Z(n2455));
Q_MX02 U2924 ( .S(n4491), .A0(n2455), .A1(n2448), .Z(r32_mux_2_data[6]));
Q_MX04 U2925 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[7]), .A1(i_cddip1_out_ia_capability[7]), .A2(i_cddip0_out_im_status[7]), .A3(o_cddip0_out_im_config[7]), .Z(n2456));
Q_MX08 U2926 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[7]), .A1(i_cddip1_out_ia_rdata_part2[7]), .A2(i_cddip1_out_ia_rdata_part1[7]), .A3(i_cddip1_out_ia_rdata_part0[7]), .A4(o_cddip1_out_ia_config[7]), .A5(o_cddip1_out_ia_wdata_part2[7]), .A6(o_cddip1_out_ia_wdata_part1[7]), .A7(o_cddip1_out_ia_wdata_part0[7]), .Z(n2457));
Q_MX02 U2927 ( .S(n4490), .A0(n2457), .A1(n2456), .Z(n2458));
Q_MX04 U2928 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[7]), .A1(i_cddip2_out_ia_status[7]), .A2(i_cddip2_out_ia_capability[7]), .A3(i_cddip1_out_im_status[7]), .Z(n2459));
Q_MX04 U2929 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[7]), .A1(o_cddip2_out_ia_config[7]), .A2(o_cddip2_out_ia_wdata_part2[7]), .A3(o_cddip2_out_ia_wdata_part1[7]), .Z(n2460));
Q_MX04 U2930 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[7]), .A1(o_cddip2_out_im_config[7]), .A2(i_cddip2_out_ia_rdata_part2[7]), .A3(i_cddip2_out_ia_rdata_part1[7]), .Z(n2461));
Q_MX02 U2931 ( .S(n4487), .A0(i_cddip3_out_ia_status[7]), .A1(i_cddip3_out_ia_capability[7]), .Z(n2462));
Q_AN02 U2932 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[7]), .Z(n2463));
Q_MX02 U2933 ( .S(n4488), .A0(n2463), .A1(n2462), .Z(n2464));
Q_MX04 U2934 ( .S0(n4489), .S1(n4490), .A0(n2464), .A1(n2461), .A2(n2460), .A3(n2459), .Z(n2465));
Q_MX02 U2935 ( .S(n4491), .A0(n2465), .A1(n2458), .Z(r32_mux_2_data[7]));
Q_MX04 U2936 ( .S0(n4487), .S1(n4488), .A0(i_cddip1_out_ia_status[8]), .A1(i_cddip1_out_ia_capability[8]), .A2(i_cddip0_out_im_status[8]), .A3(o_cddip0_out_im_config[8]), .Z(n2466));
Q_MX08 U2937 ( .S0(n4487), .S1(n4488), .S2(n4489), .A0(o_cddip1_out_im_config[8]), .A1(i_cddip1_out_ia_rdata_part2[8]), .A2(i_cddip1_out_ia_rdata_part1[8]), .A3(i_cddip1_out_ia_rdata_part0[8]), .A4(o_cddip1_out_ia_config[8]), .A5(o_cddip1_out_ia_wdata_part2[8]), .A6(o_cddip1_out_ia_wdata_part1[8]), .A7(o_cddip1_out_ia_wdata_part0[8]), .Z(n2467));
Q_MX02 U2938 ( .S(n4490), .A0(n2467), .A1(n2466), .Z(n2468));
Q_MX04 U2939 ( .S0(n4487), .S1(n4488), .A0(o_cddip2_out_ia_wdata_part0[8]), .A1(i_cddip2_out_ia_status[8]), .A2(i_cddip2_out_ia_capability[8]), .A3(i_cddip1_out_im_status[8]), .Z(n2469));
Q_MX04 U2940 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_ia_rdata_part0[8]), .A1(o_cddip2_out_ia_config[8]), .A2(o_cddip2_out_ia_wdata_part2[8]), .A3(o_cddip2_out_ia_wdata_part1[8]), .Z(n2470));
Q_MX04 U2941 ( .S0(n4487), .S1(n4488), .A0(i_cddip2_out_im_status[8]), .A1(o_cddip2_out_im_config[8]), .A2(i_cddip2_out_ia_rdata_part2[8]), .A3(i_cddip2_out_ia_rdata_part1[8]), .Z(n2471));
Q_MX02 U2942 ( .S(n4487), .A0(i_cddip3_out_ia_status[8]), .A1(i_cddip3_out_ia_capability[8]), .Z(n2472));
Q_AN02 U2943 ( .A0(n4487), .A1(o_cddip3_out_ia_wdata_part0[8]), .Z(n2473));
Q_MX02 U2944 ( .S(n4488), .A0(n2473), .A1(n2472), .Z(n2474));
Q_MX04 U2945 ( .S0(n4489), .S1(n4490), .A0(n2474), .A1(n2471), .A2(n2470), .A3(n2469), .Z(n2475));
Q_MX02 U2946 ( .S(n4491), .A0(n2475), .A1(n2468), .Z(r32_mux_2_data[8]));
Q_MX04 U2947 ( .S0(n4492), .S1(n4493), .A0(o_cddip1_out_ia_wdata_part1[9]), .A1(o_cddip1_out_ia_wdata_part0[9]), .A2(i_cddip1_out_ia_capability[9]), .A3(o_cddip0_out_im_config[9]), .Z(n2476));
Q_MX04 U2948 ( .S0(n4492), .S1(n4493), .A0(i_cddip1_out_ia_rdata_part2[9]), .A1(i_cddip1_out_ia_rdata_part1[9]), .A2(i_cddip1_out_ia_rdata_part0[9]), .A3(o_cddip1_out_ia_wdata_part2[9]), .Z(n2477));
Q_MX04 U2949 ( .S0(n4492), .S1(n4493), .A0(o_cddip2_out_ia_wdata_part1[9]), .A1(o_cddip2_out_ia_wdata_part0[9]), .A2(i_cddip2_out_ia_capability[9]), .A3(o_cddip1_out_im_config[9]), .Z(n2478));
Q_MX04 U2950 ( .S0(n4492), .S1(n4493), .A0(i_cddip2_out_ia_rdata_part2[9]), .A1(i_cddip2_out_ia_rdata_part1[9]), .A2(i_cddip2_out_ia_rdata_part0[9]), .A3(o_cddip2_out_ia_wdata_part2[9]), .Z(n2479));
Q_MX02 U2951 ( .S(n4492), .A0(i_cddip3_out_ia_capability[9]), .A1(o_cddip2_out_im_config[9]), .Z(n2480));
Q_AN02 U2952 ( .A0(n4492), .A1(o_cddip3_out_ia_wdata_part0[9]), .Z(n2481));
Q_MX02 U2953 ( .S(n4493), .A0(n2481), .A1(n2480), .Z(n2482));
Q_MX04 U2954 ( .S0(n4494), .S1(n4495), .A0(n2482), .A1(n2479), .A2(n2478), .A3(n2477), .Z(n2483));
Q_MX02 U2955 ( .S(n4496), .A0(n2483), .A1(n2476), .Z(r32_mux_2_data[9]));
Q_MX04 U2956 ( .S0(n4497), .S1(n4498), .A0(i_cddip1_out_ia_rdata_part0[10]), .A1(o_cddip1_out_ia_wdata_part2[10]), .A2(o_cddip1_out_ia_wdata_part1[10]), .A3(o_cddip1_out_ia_wdata_part0[10]), .Z(n2484));
Q_MX04 U2957 ( .S0(n4497), .S1(n4498), .A0(o_cddip2_out_ia_wdata_part0[10]), .A1(i_cddip2_out_ia_capability[10]), .A2(i_cddip1_out_ia_rdata_part2[10]), .A3(i_cddip1_out_ia_rdata_part1[10]), .Z(n2485));
Q_MX04 U2958 ( .S0(n4497), .S1(n4498), .A0(i_cddip2_out_ia_rdata_part1[10]), .A1(i_cddip2_out_ia_rdata_part0[10]), .A2(o_cddip2_out_ia_wdata_part2[10]), .A3(o_cddip2_out_ia_wdata_part1[10]), .Z(n2486));
Q_MX02 U2959 ( .S(n4497), .A0(i_cddip3_out_ia_capability[10]), .A1(i_cddip2_out_ia_rdata_part2[10]), .Z(n2487));
Q_AN02 U2960 ( .A0(n4497), .A1(o_cddip3_out_ia_wdata_part0[10]), .Z(n2488));
Q_MX02 U2961 ( .S(n4498), .A0(n2488), .A1(n2487), .Z(n2489));
Q_MX04 U2962 ( .S0(n4499), .S1(n4500), .A0(n2489), .A1(n2486), .A2(n2485), .A3(n2484), .Z(n2490));
Q_MX02 U2963 ( .S(n4501), .A0(n2490), .A1(i_cddip1_out_ia_capability[10]), .Z(r32_mux_2_data[10]));
Q_MX04 U2964 ( .S0(n4497), .S1(n4498), .A0(i_cddip1_out_ia_rdata_part0[11]), .A1(o_cddip1_out_ia_wdata_part2[11]), .A2(o_cddip1_out_ia_wdata_part1[11]), .A3(o_cddip1_out_ia_wdata_part0[11]), .Z(n2491));
Q_MX04 U2965 ( .S0(n4497), .S1(n4498), .A0(o_cddip2_out_ia_wdata_part0[11]), .A1(i_cddip2_out_ia_capability[11]), .A2(i_cddip1_out_ia_rdata_part2[11]), .A3(i_cddip1_out_ia_rdata_part1[11]), .Z(n2492));
Q_MX04 U2966 ( .S0(n4497), .S1(n4498), .A0(i_cddip2_out_ia_rdata_part1[11]), .A1(i_cddip2_out_ia_rdata_part0[11]), .A2(o_cddip2_out_ia_wdata_part2[11]), .A3(o_cddip2_out_ia_wdata_part1[11]), .Z(n2493));
Q_MX02 U2967 ( .S(n4497), .A0(i_cddip3_out_ia_capability[11]), .A1(i_cddip2_out_ia_rdata_part2[11]), .Z(n2494));
Q_AN02 U2968 ( .A0(n4497), .A1(o_cddip3_out_ia_wdata_part0[11]), .Z(n2495));
Q_MX02 U2969 ( .S(n4498), .A0(n2495), .A1(n2494), .Z(n2496));
Q_MX04 U2970 ( .S0(n4499), .S1(n4500), .A0(n2496), .A1(n2493), .A2(n2492), .A3(n2491), .Z(n2497));
Q_MX02 U2971 ( .S(n4501), .A0(n2497), .A1(i_cddip1_out_ia_capability[11]), .Z(r32_mux_2_data[11]));
Q_MX04 U2972 ( .S0(n4497), .S1(n4498), .A0(i_cddip1_out_ia_rdata_part0[12]), .A1(o_cddip1_out_ia_wdata_part2[12]), .A2(o_cddip1_out_ia_wdata_part1[12]), .A3(o_cddip1_out_ia_wdata_part0[12]), .Z(n2498));
Q_MX04 U2973 ( .S0(n4497), .S1(n4498), .A0(o_cddip2_out_ia_wdata_part0[12]), .A1(i_cddip2_out_ia_capability[12]), .A2(i_cddip1_out_ia_rdata_part2[12]), .A3(i_cddip1_out_ia_rdata_part1[12]), .Z(n2499));
Q_MX04 U2974 ( .S0(n4497), .S1(n4498), .A0(i_cddip2_out_ia_rdata_part1[12]), .A1(i_cddip2_out_ia_rdata_part0[12]), .A2(o_cddip2_out_ia_wdata_part2[12]), .A3(o_cddip2_out_ia_wdata_part1[12]), .Z(n2500));
Q_MX02 U2975 ( .S(n4497), .A0(i_cddip3_out_ia_capability[12]), .A1(i_cddip2_out_ia_rdata_part2[12]), .Z(n2501));
Q_AN02 U2976 ( .A0(n4497), .A1(o_cddip3_out_ia_wdata_part0[12]), .Z(n2502));
Q_MX02 U2977 ( .S(n4498), .A0(n2502), .A1(n2501), .Z(n2503));
Q_MX04 U2978 ( .S0(n4499), .S1(n4500), .A0(n2503), .A1(n2500), .A2(n2499), .A3(n2498), .Z(n2504));
Q_MX02 U2979 ( .S(n4501), .A0(n2504), .A1(i_cddip1_out_ia_capability[12]), .Z(r32_mux_2_data[12]));
Q_MX04 U2980 ( .S0(n4497), .S1(n4498), .A0(i_cddip1_out_ia_rdata_part0[13]), .A1(o_cddip1_out_ia_wdata_part2[13]), .A2(o_cddip1_out_ia_wdata_part1[13]), .A3(o_cddip1_out_ia_wdata_part0[13]), .Z(n2505));
Q_MX04 U2981 ( .S0(n4497), .S1(n4498), .A0(o_cddip2_out_ia_wdata_part0[13]), .A1(i_cddip2_out_ia_capability[13]), .A2(i_cddip1_out_ia_rdata_part2[13]), .A3(i_cddip1_out_ia_rdata_part1[13]), .Z(n2506));
Q_MX04 U2982 ( .S0(n4497), .S1(n4498), .A0(i_cddip2_out_ia_rdata_part1[13]), .A1(i_cddip2_out_ia_rdata_part0[13]), .A2(o_cddip2_out_ia_wdata_part2[13]), .A3(o_cddip2_out_ia_wdata_part1[13]), .Z(n2507));
Q_MX02 U2983 ( .S(n4497), .A0(i_cddip3_out_ia_capability[13]), .A1(i_cddip2_out_ia_rdata_part2[13]), .Z(n2508));
Q_AN02 U2984 ( .A0(n4497), .A1(o_cddip3_out_ia_wdata_part0[13]), .Z(n2509));
Q_MX02 U2985 ( .S(n4498), .A0(n2509), .A1(n2508), .Z(n2510));
Q_MX04 U2986 ( .S0(n4499), .S1(n4500), .A0(n2510), .A1(n2507), .A2(n2506), .A3(n2505), .Z(n2511));
Q_MX02 U2987 ( .S(n4501), .A0(n2511), .A1(i_cddip1_out_ia_capability[13]), .Z(r32_mux_2_data[13]));
Q_MX04 U2988 ( .S0(n4497), .S1(n4498), .A0(i_cddip1_out_ia_rdata_part0[14]), .A1(o_cddip1_out_ia_wdata_part2[14]), .A2(o_cddip1_out_ia_wdata_part1[14]), .A3(o_cddip1_out_ia_wdata_part0[14]), .Z(n2512));
Q_MX04 U2989 ( .S0(n4497), .S1(n4498), .A0(o_cddip2_out_ia_wdata_part0[14]), .A1(i_cddip2_out_ia_capability[14]), .A2(i_cddip1_out_ia_rdata_part2[14]), .A3(i_cddip1_out_ia_rdata_part1[14]), .Z(n2513));
Q_MX04 U2990 ( .S0(n4497), .S1(n4498), .A0(i_cddip2_out_ia_rdata_part1[14]), .A1(i_cddip2_out_ia_rdata_part0[14]), .A2(o_cddip2_out_ia_wdata_part2[14]), .A3(o_cddip2_out_ia_wdata_part1[14]), .Z(n2514));
Q_MX02 U2991 ( .S(n4497), .A0(i_cddip3_out_ia_capability[14]), .A1(i_cddip2_out_ia_rdata_part2[14]), .Z(n2515));
Q_AN02 U2992 ( .A0(n4497), .A1(o_cddip3_out_ia_wdata_part0[14]), .Z(n2516));
Q_MX02 U2993 ( .S(n4498), .A0(n2516), .A1(n2515), .Z(n2517));
Q_MX04 U2994 ( .S0(n4499), .S1(n4500), .A0(n2517), .A1(n2514), .A2(n2513), .A3(n2512), .Z(n2518));
Q_MX02 U2995 ( .S(n4501), .A0(n2518), .A1(i_cddip1_out_ia_capability[14]), .Z(r32_mux_2_data[14]));
Q_MX04 U2996 ( .S0(n4497), .S1(n4498), .A0(i_cddip1_out_ia_rdata_part0[15]), .A1(o_cddip1_out_ia_wdata_part2[15]), .A2(o_cddip1_out_ia_wdata_part1[15]), .A3(o_cddip1_out_ia_wdata_part0[15]), .Z(n2519));
Q_MX04 U2997 ( .S0(n4497), .S1(n4498), .A0(o_cddip2_out_ia_wdata_part0[15]), .A1(i_cddip2_out_ia_capability[15]), .A2(i_cddip1_out_ia_rdata_part2[15]), .A3(i_cddip1_out_ia_rdata_part1[15]), .Z(n2520));
Q_MX04 U2998 ( .S0(n4497), .S1(n4498), .A0(i_cddip2_out_ia_rdata_part1[15]), .A1(i_cddip2_out_ia_rdata_part0[15]), .A2(o_cddip2_out_ia_wdata_part2[15]), .A3(o_cddip2_out_ia_wdata_part1[15]), .Z(n2521));
Q_MX02 U2999 ( .S(n4497), .A0(i_cddip3_out_ia_capability[15]), .A1(i_cddip2_out_ia_rdata_part2[15]), .Z(n2522));
Q_AN02 U3000 ( .A0(n4497), .A1(o_cddip3_out_ia_wdata_part0[15]), .Z(n2523));
Q_MX02 U3001 ( .S(n4498), .A0(n2523), .A1(n2522), .Z(n2524));
Q_MX04 U3002 ( .S0(n4499), .S1(n4500), .A0(n2524), .A1(n2521), .A2(n2520), .A3(n2519), .Z(n2525));
Q_MX02 U3003 ( .S(n4501), .A0(n2525), .A1(i_cddip1_out_ia_capability[15]), .Z(r32_mux_2_data[15]));
Q_MX02 U3004 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[16]), .A1(o_cddip1_out_ia_wdata_part0[16]), .Z(n2526));
Q_MX04 U3005 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[16]), .A1(i_cddip1_out_ia_rdata_part1[16]), .A2(i_cddip1_out_ia_rdata_part0[16]), .A3(o_cddip1_out_ia_wdata_part2[16]), .Z(n2527));
Q_MX02 U3006 ( .S(n4504), .A0(n2527), .A1(n2526), .Z(n2528));
Q_MX04 U3007 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[16]), .A1(o_cddip2_out_ia_wdata_part2[16]), .A2(o_cddip2_out_ia_wdata_part1[16]), .A3(o_cddip2_out_ia_wdata_part0[16]), .Z(n2529));
Q_MX02 U3008 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[16]), .A1(i_cddip2_out_ia_rdata_part1[16]), .Z(n2530));
Q_AN02 U3009 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[16]), .Z(n2531));
Q_MX03 U3010 ( .S0(n4503), .S1(n4504), .A0(n2531), .A1(n2530), .A2(n2529), .Z(n2532));
Q_MX02 U3011 ( .S(n4505), .A0(n2532), .A1(n2528), .Z(r32_mux_2_data[16]));
Q_MX02 U3012 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[17]), .A1(o_cddip1_out_ia_wdata_part0[17]), .Z(n2533));
Q_MX04 U3013 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[17]), .A1(i_cddip1_out_ia_rdata_part1[17]), .A2(i_cddip1_out_ia_rdata_part0[17]), .A3(o_cddip1_out_ia_wdata_part2[17]), .Z(n2534));
Q_MX02 U3014 ( .S(n4504), .A0(n2534), .A1(n2533), .Z(n2535));
Q_MX04 U3015 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[17]), .A1(o_cddip2_out_ia_wdata_part2[17]), .A2(o_cddip2_out_ia_wdata_part1[17]), .A3(o_cddip2_out_ia_wdata_part0[17]), .Z(n2536));
Q_MX02 U3016 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[17]), .A1(i_cddip2_out_ia_rdata_part1[17]), .Z(n2537));
Q_AN02 U3017 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[17]), .Z(n2538));
Q_MX03 U3018 ( .S0(n4503), .S1(n4504), .A0(n2538), .A1(n2537), .A2(n2536), .Z(n2539));
Q_MX02 U3019 ( .S(n4505), .A0(n2539), .A1(n2535), .Z(r32_mux_2_data[17]));
Q_MX02 U3020 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[18]), .A1(o_cddip1_out_ia_wdata_part0[18]), .Z(n2540));
Q_MX04 U3021 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[18]), .A1(i_cddip1_out_ia_rdata_part1[18]), .A2(i_cddip1_out_ia_rdata_part0[18]), .A3(o_cddip1_out_ia_wdata_part2[18]), .Z(n2541));
Q_MX02 U3022 ( .S(n4504), .A0(n2541), .A1(n2540), .Z(n2542));
Q_MX04 U3023 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[18]), .A1(o_cddip2_out_ia_wdata_part2[18]), .A2(o_cddip2_out_ia_wdata_part1[18]), .A3(o_cddip2_out_ia_wdata_part0[18]), .Z(n2543));
Q_MX02 U3024 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[18]), .A1(i_cddip2_out_ia_rdata_part1[18]), .Z(n2544));
Q_AN02 U3025 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[18]), .Z(n2545));
Q_MX03 U3026 ( .S0(n4503), .S1(n4504), .A0(n2545), .A1(n2544), .A2(n2543), .Z(n2546));
Q_MX02 U3027 ( .S(n4505), .A0(n2546), .A1(n2542), .Z(r32_mux_2_data[18]));
Q_MX02 U3028 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[19]), .A1(o_cddip1_out_ia_wdata_part0[19]), .Z(n2547));
Q_MX04 U3029 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[19]), .A1(i_cddip1_out_ia_rdata_part1[19]), .A2(i_cddip1_out_ia_rdata_part0[19]), .A3(o_cddip1_out_ia_wdata_part2[19]), .Z(n2548));
Q_MX02 U3030 ( .S(n4504), .A0(n2548), .A1(n2547), .Z(n2549));
Q_MX04 U3031 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[19]), .A1(o_cddip2_out_ia_wdata_part2[19]), .A2(o_cddip2_out_ia_wdata_part1[19]), .A3(o_cddip2_out_ia_wdata_part0[19]), .Z(n2550));
Q_MX02 U3032 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[19]), .A1(i_cddip2_out_ia_rdata_part1[19]), .Z(n2551));
Q_AN02 U3033 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[19]), .Z(n2552));
Q_MX03 U3034 ( .S0(n4503), .S1(n4504), .A0(n2552), .A1(n2551), .A2(n2550), .Z(n2553));
Q_MX02 U3035 ( .S(n4505), .A0(n2553), .A1(n2549), .Z(r32_mux_2_data[19]));
Q_MX02 U3036 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[20]), .A1(o_cddip1_out_ia_wdata_part0[20]), .Z(n2554));
Q_MX04 U3037 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[20]), .A1(i_cddip1_out_ia_rdata_part1[20]), .A2(i_cddip1_out_ia_rdata_part0[20]), .A3(o_cddip1_out_ia_wdata_part2[20]), .Z(n2555));
Q_MX02 U3038 ( .S(n4504), .A0(n2555), .A1(n2554), .Z(n2556));
Q_MX04 U3039 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[20]), .A1(o_cddip2_out_ia_wdata_part2[20]), .A2(o_cddip2_out_ia_wdata_part1[20]), .A3(o_cddip2_out_ia_wdata_part0[20]), .Z(n2557));
Q_MX02 U3040 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[20]), .A1(i_cddip2_out_ia_rdata_part1[20]), .Z(n2558));
Q_AN02 U3041 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[20]), .Z(n2559));
Q_MX03 U3042 ( .S0(n4503), .S1(n4504), .A0(n2559), .A1(n2558), .A2(n2557), .Z(n2560));
Q_MX02 U3043 ( .S(n4505), .A0(n2560), .A1(n2556), .Z(r32_mux_2_data[20]));
Q_MX02 U3044 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[21]), .A1(o_cddip1_out_ia_wdata_part0[21]), .Z(n2561));
Q_MX04 U3045 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[21]), .A1(i_cddip1_out_ia_rdata_part1[21]), .A2(i_cddip1_out_ia_rdata_part0[21]), .A3(o_cddip1_out_ia_wdata_part2[21]), .Z(n2562));
Q_MX02 U3046 ( .S(n4504), .A0(n2562), .A1(n2561), .Z(n2563));
Q_MX04 U3047 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[21]), .A1(o_cddip2_out_ia_wdata_part2[21]), .A2(o_cddip2_out_ia_wdata_part1[21]), .A3(o_cddip2_out_ia_wdata_part0[21]), .Z(n2564));
Q_MX02 U3048 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[21]), .A1(i_cddip2_out_ia_rdata_part1[21]), .Z(n2565));
Q_AN02 U3049 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[21]), .Z(n2566));
Q_MX03 U3050 ( .S0(n4503), .S1(n4504), .A0(n2566), .A1(n2565), .A2(n2564), .Z(n2567));
Q_MX02 U3051 ( .S(n4505), .A0(n2567), .A1(n2563), .Z(r32_mux_2_data[21]));
Q_MX02 U3052 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[22]), .A1(o_cddip1_out_ia_wdata_part0[22]), .Z(n2568));
Q_MX04 U3053 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[22]), .A1(i_cddip1_out_ia_rdata_part1[22]), .A2(i_cddip1_out_ia_rdata_part0[22]), .A3(o_cddip1_out_ia_wdata_part2[22]), .Z(n2569));
Q_MX02 U3054 ( .S(n4504), .A0(n2569), .A1(n2568), .Z(n2570));
Q_MX04 U3055 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[22]), .A1(o_cddip2_out_ia_wdata_part2[22]), .A2(o_cddip2_out_ia_wdata_part1[22]), .A3(o_cddip2_out_ia_wdata_part0[22]), .Z(n2571));
Q_MX02 U3056 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[22]), .A1(i_cddip2_out_ia_rdata_part1[22]), .Z(n2572));
Q_AN02 U3057 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[22]), .Z(n2573));
Q_MX03 U3058 ( .S0(n4503), .S1(n4504), .A0(n2573), .A1(n2572), .A2(n2571), .Z(n2574));
Q_MX02 U3059 ( .S(n4505), .A0(n2574), .A1(n2570), .Z(r32_mux_2_data[22]));
Q_MX02 U3060 ( .S(n4502), .A0(o_cddip1_out_ia_wdata_part1[23]), .A1(o_cddip1_out_ia_wdata_part0[23]), .Z(n2575));
Q_MX04 U3061 ( .S0(n4502), .S1(n4503), .A0(i_cddip1_out_ia_rdata_part2[23]), .A1(i_cddip1_out_ia_rdata_part1[23]), .A2(i_cddip1_out_ia_rdata_part0[23]), .A3(o_cddip1_out_ia_wdata_part2[23]), .Z(n2576));
Q_MX02 U3062 ( .S(n4504), .A0(n2576), .A1(n2575), .Z(n2577));
Q_MX04 U3063 ( .S0(n4502), .S1(n4503), .A0(i_cddip2_out_ia_rdata_part0[23]), .A1(o_cddip2_out_ia_wdata_part2[23]), .A2(o_cddip2_out_ia_wdata_part1[23]), .A3(o_cddip2_out_ia_wdata_part0[23]), .Z(n2578));
Q_MX02 U3064 ( .S(n4502), .A0(i_cddip2_out_ia_rdata_part2[23]), .A1(i_cddip2_out_ia_rdata_part1[23]), .Z(n2579));
Q_AN02 U3065 ( .A0(n4502), .A1(o_cddip3_out_ia_wdata_part0[23]), .Z(n2580));
Q_MX03 U3066 ( .S0(n4503), .S1(n4504), .A0(n2580), .A1(n2579), .A2(n2578), .Z(n2581));
Q_MX02 U3067 ( .S(n4505), .A0(n2581), .A1(n2577), .Z(r32_mux_2_data[23]));
Q_MX04 U3068 ( .S0(n4506), .S1(n4507), .A0(i_cddip1_out_ia_rdata_part0[24]), .A1(o_cddip1_out_ia_wdata_part2[24]), .A2(o_cddip1_out_ia_wdata_part1[24]), .A3(o_cddip1_out_ia_wdata_part0[24]), .Z(n2582));
Q_MX04 U3069 ( .S0(n4506), .S1(n4507), .A0(o_cddip2_out_ia_wdata_part0[24]), .A1(i_cddip2_out_ia_status[9]), .A2(i_cddip1_out_ia_rdata_part2[24]), .A3(i_cddip1_out_ia_rdata_part1[24]), .Z(n2583));
Q_MX04 U3070 ( .S0(n4506), .S1(n4507), .A0(i_cddip2_out_ia_rdata_part1[24]), .A1(i_cddip2_out_ia_rdata_part0[24]), .A2(o_cddip2_out_ia_wdata_part2[24]), .A3(o_cddip2_out_ia_wdata_part1[24]), .Z(n2584));
Q_MX02 U3071 ( .S(n4506), .A0(i_cddip3_out_ia_status[9]), .A1(i_cddip2_out_ia_rdata_part2[24]), .Z(n2585));
Q_AN02 U3072 ( .A0(n4506), .A1(o_cddip3_out_ia_wdata_part0[24]), .Z(n2586));
Q_MX02 U3073 ( .S(n4507), .A0(n2586), .A1(n2585), .Z(n2587));
Q_MX04 U3074 ( .S0(n4499), .S1(n4508), .A0(n2587), .A1(n2584), .A2(n2583), .A3(n2582), .Z(n2588));
Q_MX02 U3075 ( .S(n4509), .A0(n2588), .A1(i_cddip1_out_ia_status[9]), .Z(r32_mux_2_data[24]));
Q_MX04 U3076 ( .S0(n4506), .S1(n4507), .A0(i_cddip1_out_ia_rdata_part0[25]), .A1(o_cddip1_out_ia_wdata_part2[25]), .A2(o_cddip1_out_ia_wdata_part1[25]), .A3(o_cddip1_out_ia_wdata_part0[25]), .Z(n2589));
Q_MX04 U3077 ( .S0(n4506), .S1(n4507), .A0(o_cddip2_out_ia_wdata_part0[25]), .A1(i_cddip2_out_ia_status[10]), .A2(i_cddip1_out_ia_rdata_part2[25]), .A3(i_cddip1_out_ia_rdata_part1[25]), .Z(n2590));
Q_MX04 U3078 ( .S0(n4506), .S1(n4507), .A0(i_cddip2_out_ia_rdata_part1[25]), .A1(i_cddip2_out_ia_rdata_part0[25]), .A2(o_cddip2_out_ia_wdata_part2[25]), .A3(o_cddip2_out_ia_wdata_part1[25]), .Z(n2591));
Q_MX02 U3079 ( .S(n4506), .A0(i_cddip3_out_ia_status[10]), .A1(i_cddip2_out_ia_rdata_part2[25]), .Z(n2592));
Q_AN02 U3080 ( .A0(n4506), .A1(o_cddip3_out_ia_wdata_part0[25]), .Z(n2593));
Q_MX02 U3081 ( .S(n4507), .A0(n2593), .A1(n2592), .Z(n2594));
Q_MX04 U3082 ( .S0(n4499), .S1(n4508), .A0(n2594), .A1(n2591), .A2(n2590), .A3(n2589), .Z(n2595));
Q_MX02 U3083 ( .S(n4509), .A0(n2595), .A1(i_cddip1_out_ia_status[10]), .Z(r32_mux_2_data[25]));
Q_MX04 U3084 ( .S0(n4506), .S1(n4507), .A0(i_cddip1_out_ia_rdata_part0[26]), .A1(o_cddip1_out_ia_wdata_part2[26]), .A2(o_cddip1_out_ia_wdata_part1[26]), .A3(o_cddip1_out_ia_wdata_part0[26]), .Z(n2596));
Q_MX04 U3085 ( .S0(n4506), .S1(n4507), .A0(o_cddip2_out_ia_wdata_part0[26]), .A1(i_cddip2_out_ia_status[11]), .A2(i_cddip1_out_ia_rdata_part2[26]), .A3(i_cddip1_out_ia_rdata_part1[26]), .Z(n2597));
Q_MX04 U3086 ( .S0(n4506), .S1(n4507), .A0(i_cddip2_out_ia_rdata_part1[26]), .A1(i_cddip2_out_ia_rdata_part0[26]), .A2(o_cddip2_out_ia_wdata_part2[26]), .A3(o_cddip2_out_ia_wdata_part1[26]), .Z(n2598));
Q_MX02 U3087 ( .S(n4506), .A0(i_cddip3_out_ia_status[11]), .A1(i_cddip2_out_ia_rdata_part2[26]), .Z(n2599));
Q_AN02 U3088 ( .A0(n4506), .A1(o_cddip3_out_ia_wdata_part0[26]), .Z(n2600));
Q_MX02 U3089 ( .S(n4507), .A0(n2600), .A1(n2599), .Z(n2601));
Q_MX04 U3090 ( .S0(n4499), .S1(n4508), .A0(n2601), .A1(n2598), .A2(n2597), .A3(n2596), .Z(n2602));
Q_MX02 U3091 ( .S(n4509), .A0(n2602), .A1(i_cddip1_out_ia_status[11]), .Z(r32_mux_2_data[26]));
Q_MX04 U3092 ( .S0(n4506), .S1(n4507), .A0(i_cddip1_out_ia_rdata_part0[27]), .A1(o_cddip1_out_ia_wdata_part2[27]), .A2(o_cddip1_out_ia_wdata_part1[27]), .A3(o_cddip1_out_ia_wdata_part0[27]), .Z(n2603));
Q_MX04 U3093 ( .S0(n4506), .S1(n4507), .A0(o_cddip2_out_ia_wdata_part0[27]), .A1(i_cddip2_out_ia_status[12]), .A2(i_cddip1_out_ia_rdata_part2[27]), .A3(i_cddip1_out_ia_rdata_part1[27]), .Z(n2604));
Q_MX04 U3094 ( .S0(n4506), .S1(n4507), .A0(i_cddip2_out_ia_rdata_part1[27]), .A1(i_cddip2_out_ia_rdata_part0[27]), .A2(o_cddip2_out_ia_wdata_part2[27]), .A3(o_cddip2_out_ia_wdata_part1[27]), .Z(n2605));
Q_MX02 U3095 ( .S(n4506), .A0(i_cddip3_out_ia_status[12]), .A1(i_cddip2_out_ia_rdata_part2[27]), .Z(n2606));
Q_AN02 U3096 ( .A0(n4506), .A1(o_cddip3_out_ia_wdata_part0[27]), .Z(n2607));
Q_MX02 U3097 ( .S(n4507), .A0(n2607), .A1(n2606), .Z(n2608));
Q_MX04 U3098 ( .S0(n4499), .S1(n4508), .A0(n2608), .A1(n2605), .A2(n2604), .A3(n2603), .Z(n2609));
Q_MX02 U3099 ( .S(n4509), .A0(n2609), .A1(i_cddip1_out_ia_status[12]), .Z(r32_mux_2_data[27]));
Q_MX02 U3100 ( .S(n4510), .A0(i_cddip1_out_ia_status[13]), .A1(i_cddip1_out_ia_capability[16]), .Z(n2610));
Q_MX04 U3101 ( .S0(n4510), .S1(n4511), .A0(o_cddip1_out_ia_config[9]), .A1(o_cddip1_out_ia_wdata_part2[28]), .A2(o_cddip1_out_ia_wdata_part1[28]), .A3(o_cddip1_out_ia_wdata_part0[28]), .Z(n2611));
Q_MX02 U3102 ( .S(n4512), .A0(n2611), .A1(n2610), .Z(n2612));
Q_MX04 U3103 ( .S0(n4510), .S1(n4511), .A0(i_cddip2_out_ia_capability[16]), .A1(i_cddip1_out_ia_rdata_part2[28]), .A2(i_cddip1_out_ia_rdata_part1[28]), .A3(i_cddip1_out_ia_rdata_part0[28]), .Z(n2613));
Q_MX04 U3104 ( .S0(n4510), .S1(n4511), .A0(o_cddip2_out_ia_wdata_part2[28]), .A1(o_cddip2_out_ia_wdata_part1[28]), .A2(o_cddip2_out_ia_wdata_part0[28]), .A3(i_cddip2_out_ia_status[13]), .Z(n2614));
Q_MX04 U3105 ( .S0(n4510), .S1(n4511), .A0(i_cddip2_out_ia_rdata_part2[28]), .A1(i_cddip2_out_ia_rdata_part1[28]), .A2(i_cddip2_out_ia_rdata_part0[28]), .A3(o_cddip2_out_ia_config[9]), .Z(n2615));
Q_MX02 U3106 ( .S(n4510), .A0(i_cddip3_out_ia_status[13]), .A1(i_cddip3_out_ia_capability[16]), .Z(n2616));
Q_AN02 U3107 ( .A0(n4510), .A1(o_cddip3_out_ia_wdata_part0[28]), .Z(n2617));
Q_MX02 U3108 ( .S(n4511), .A0(n2617), .A1(n2616), .Z(n2618));
Q_MX04 U3109 ( .S0(n4512), .S1(n4513), .A0(n2618), .A1(n2615), .A2(n2614), .A3(n2613), .Z(n2619));
Q_MX02 U3110 ( .S(n4514), .A0(n2619), .A1(n2612), .Z(r32_mux_2_data[28]));
Q_MX08 U3111 ( .S0(n4515), .S1(n4516), .S2(n4517), .A0(i_cddip1_out_ia_rdata_part1[29]), .A1(i_cddip1_out_ia_rdata_part0[29]), .A2(o_cddip1_out_ia_config[10]), .A3(o_cddip1_out_ia_wdata_part2[29]), .A4(o_cddip1_out_ia_wdata_part1[29]), .A5(o_cddip1_out_ia_wdata_part0[29]), .A6(i_cddip1_out_ia_status[14]), .A7(i_cddip1_out_ia_capability[17]), .Z(n2620));
Q_MX02 U3112 ( .S(n4518), .A0(n2620), .A1(i_cddip0_out_im_status[9]), .Z(n2621));
Q_MX04 U3113 ( .S0(n4515), .S1(n4516), .A0(i_cddip2_out_ia_status[14]), .A1(i_cddip2_out_ia_capability[17]), .A2(i_cddip1_out_im_status[9]), .A3(i_cddip1_out_ia_rdata_part2[29]), .Z(n2622));
Q_MX04 U3114 ( .S0(n4515), .S1(n4516), .A0(o_cddip2_out_ia_config[10]), .A1(o_cddip2_out_ia_wdata_part2[29]), .A2(o_cddip2_out_ia_wdata_part1[29]), .A3(o_cddip2_out_ia_wdata_part0[29]), .Z(n2623));
Q_MX04 U3115 ( .S0(n4515), .S1(n4516), .A0(i_cddip2_out_im_status[9]), .A1(i_cddip2_out_ia_rdata_part2[29]), .A2(i_cddip2_out_ia_rdata_part1[29]), .A3(i_cddip2_out_ia_rdata_part0[29]), .Z(n2624));
Q_MX02 U3116 ( .S(n4515), .A0(i_cddip3_out_ia_status[14]), .A1(i_cddip3_out_ia_capability[17]), .Z(n2625));
Q_AN02 U3117 ( .A0(n4515), .A1(o_cddip3_out_ia_wdata_part0[29]), .Z(n2626));
Q_MX02 U3118 ( .S(n4516), .A0(n2626), .A1(n2625), .Z(n2627));
Q_MX04 U3119 ( .S0(n4517), .S1(n4518), .A0(n2627), .A1(n2624), .A2(n2623), .A3(n2622), .Z(n2628));
Q_MX02 U3120 ( .S(n4519), .A0(n2628), .A1(n2621), .Z(r32_mux_2_data[29]));
Q_MX03 U3121 ( .S0(n4520), .S1(n4521), .A0(i_cddip0_out_im_read_done[0]), .A1(i_cddip0_out_im_status[10]), .A2(o_cddip0_out_im_config[10]), .Z(n2629));
Q_MX04 U3122 ( .S0(n4520), .S1(n4521), .A0(o_cddip1_out_ia_wdata_part1[30]), .A1(o_cddip1_out_ia_wdata_part0[30]), .A2(i_cddip1_out_ia_status[15]), .A3(i_cddip1_out_ia_capability[18]), .Z(n2630));
Q_MX02 U3123 ( .S(n4522), .A0(n2630), .A1(n2629), .Z(n2631));
Q_MX08 U3124 ( .S0(n4520), .S1(n4521), .S2(n4522), .A0(i_cddip1_out_im_read_done[0]), .A1(i_cddip1_out_im_status[10]), .A2(o_cddip1_out_im_config[10]), .A3(i_cddip1_out_ia_rdata_part2[30]), .A4(i_cddip1_out_ia_rdata_part1[30]), .A5(i_cddip1_out_ia_rdata_part0[30]), .A6(o_cddip1_out_ia_config[11]), .A7(o_cddip1_out_ia_wdata_part2[30]), .Z(n2632));
Q_MX02 U3125 ( .S(n4523), .A0(n2632), .A1(n2631), .Z(n2633));
Q_MX04 U3126 ( .S0(n4520), .S1(n4521), .A0(o_cddip2_out_ia_wdata_part1[30]), .A1(o_cddip2_out_ia_wdata_part0[30]), .A2(i_cddip2_out_ia_status[15]), .A3(i_cddip2_out_ia_capability[18]), .Z(n2634));
Q_MX04 U3127 ( .S0(n4520), .S1(n4521), .A0(i_cddip2_out_ia_rdata_part1[30]), .A1(i_cddip2_out_ia_rdata_part0[30]), .A2(o_cddip2_out_ia_config[11]), .A3(o_cddip2_out_ia_wdata_part2[30]), .Z(n2635));
Q_MX04 U3128 ( .S0(n4520), .S1(n4521), .A0(i_cddip2_out_im_read_done[0]), .A1(i_cddip2_out_im_status[10]), .A2(o_cddip2_out_im_config[10]), .A3(i_cddip2_out_ia_rdata_part2[30]), .Z(n2636));
Q_MX02 U3129 ( .S(n4520), .A0(i_cddip3_out_ia_status[15]), .A1(i_cddip3_out_ia_capability[18]), .Z(n2637));
Q_AN02 U3130 ( .A0(n4520), .A1(o_cddip3_out_ia_wdata_part0[30]), .Z(n2638));
Q_MX02 U3131 ( .S(n4521), .A0(n2638), .A1(n2637), .Z(n2639));
Q_MX04 U3132 ( .S0(n4522), .S1(n4523), .A0(n2639), .A1(n2636), .A2(n2635), .A3(n2634), .Z(n2640));
Q_MX02 U3133 ( .S(n4524), .A0(n2640), .A1(n2633), .Z(r32_mux_2_data[30]));
Q_MX03 U3134 ( .S0(n4520), .S1(n4521), .A0(i_cddip0_out_im_read_done[1]), .A1(i_cddip0_out_im_status[11]), .A2(o_cddip0_out_im_config[11]), .Z(n2641));
Q_MX04 U3135 ( .S0(n4520), .S1(n4521), .A0(o_cddip1_out_ia_wdata_part1[31]), .A1(o_cddip1_out_ia_wdata_part0[31]), .A2(i_cddip1_out_ia_status[16]), .A3(i_cddip1_out_ia_capability[19]), .Z(n2642));
Q_MX02 U3136 ( .S(n4522), .A0(n2642), .A1(n2641), .Z(n2643));
Q_MX08 U3137 ( .S0(n4520), .S1(n4521), .S2(n4522), .A0(i_cddip1_out_im_read_done[1]), .A1(i_cddip1_out_im_status[11]), .A2(o_cddip1_out_im_config[11]), .A3(i_cddip1_out_ia_rdata_part2[31]), .A4(i_cddip1_out_ia_rdata_part1[31]), .A5(i_cddip1_out_ia_rdata_part0[31]), .A6(o_cddip1_out_ia_config[12]), .A7(o_cddip1_out_ia_wdata_part2[31]), .Z(n2644));
Q_MX02 U3138 ( .S(n4523), .A0(n2644), .A1(n2643), .Z(n2645));
Q_MX04 U3139 ( .S0(n4520), .S1(n4521), .A0(o_cddip2_out_ia_wdata_part1[31]), .A1(o_cddip2_out_ia_wdata_part0[31]), .A2(i_cddip2_out_ia_status[16]), .A3(i_cddip2_out_ia_capability[19]), .Z(n2646));
Q_MX04 U3140 ( .S0(n4520), .S1(n4521), .A0(i_cddip2_out_ia_rdata_part1[31]), .A1(i_cddip2_out_ia_rdata_part0[31]), .A2(o_cddip2_out_ia_config[12]), .A3(o_cddip2_out_ia_wdata_part2[31]), .Z(n2647));
Q_MX04 U3141 ( .S0(n4520), .S1(n4521), .A0(i_cddip2_out_im_read_done[1]), .A1(i_cddip2_out_im_status[11]), .A2(o_cddip2_out_im_config[11]), .A3(i_cddip2_out_ia_rdata_part2[31]), .Z(n2648));
Q_MX02 U3142 ( .S(n4520), .A0(i_cddip3_out_ia_status[16]), .A1(i_cddip3_out_ia_capability[19]), .Z(n2649));
Q_AN02 U3143 ( .A0(n4520), .A1(o_cddip3_out_ia_wdata_part0[31]), .Z(n2650));
Q_MX02 U3144 ( .S(n4521), .A0(n2650), .A1(n2649), .Z(n2651));
Q_MX04 U3145 ( .S0(n4522), .S1(n4523), .A0(n2651), .A1(n2648), .A2(n2647), .A3(n2646), .Z(n2652));
Q_MX02 U3146 ( .S(n4524), .A0(n2652), .A1(n2645), .Z(r32_mux_2_data[31]));
Q_MX04 U3147 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[0]), .A1(i_cceip2_out_ia_rdata_part0[0]), .A2(o_cceip2_out_ia_config[0]), .A3(o_cceip2_out_ia_wdata_part2[0]), .Z(n2653));
Q_MX02 U3148 ( .S(n4527), .A0(n2653), .A1(o_cceip2_out_ia_wdata_part1[0]), .Z(n2654));
Q_MX08 U3149 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[0]), .A1(o_cceip3_out_ia_wdata_part1[0]), .A2(o_cceip3_out_ia_wdata_part0[0]), .A3(i_cceip3_out_ia_status[0]), .A4(i_cceip3_out_ia_capability[0]), .A5(i_cceip2_out_im_status[0]), .A6(o_cceip2_out_im_config[0]), .A7(i_cceip2_out_ia_rdata_part2[0]), .Z(n2655));
Q_MX02 U3150 ( .S(n4528), .A0(n2655), .A1(n2654), .Z(n2656));
Q_MX04 U3151 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[0]), .A1(i_cceip3_out_ia_rdata_part1[0]), .A2(i_cceip3_out_ia_rdata_part0[0]), .A3(o_cceip3_out_ia_config[0]), .Z(n2657));
Q_MX04 U3152 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[0]), .A1(i_cddip0_out_ia_capability[0]), .A2(i_cceip3_out_im_status[0]), .A3(o_cceip3_out_im_config[0]), .Z(n2658));
Q_MX04 U3153 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[0]), .A1(o_cddip0_out_ia_wdata_part2[0]), .A2(o_cddip0_out_ia_wdata_part1[0]), .A3(o_cddip0_out_ia_wdata_part0[0]), .Z(n2659));
Q_MX02 U3154 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[0]), .A1(i_cddip0_out_ia_rdata_part0[0]), .Z(n2660));
Q_AN02 U3155 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[0]), .Z(n2661));
Q_MX02 U3156 ( .S(n4526), .A0(n2661), .A1(n2660), .Z(n2662));
Q_MX04 U3157 ( .S0(n4527), .S1(n4528), .A0(n2662), .A1(n2659), .A2(n2658), .A3(n2657), .Z(n2663));
Q_MX02 U3158 ( .S(n4529), .A0(n2663), .A1(n2656), .Z(r32_mux_1_data[0]));
Q_MX04 U3159 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[1]), .A1(i_cceip2_out_ia_rdata_part0[1]), .A2(o_cceip2_out_ia_config[1]), .A3(o_cceip2_out_ia_wdata_part2[1]), .Z(n2664));
Q_MX02 U3160 ( .S(n4527), .A0(n2664), .A1(o_cceip2_out_ia_wdata_part1[1]), .Z(n2665));
Q_MX08 U3161 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[1]), .A1(o_cceip3_out_ia_wdata_part1[1]), .A2(o_cceip3_out_ia_wdata_part0[1]), .A3(i_cceip3_out_ia_status[1]), .A4(i_cceip3_out_ia_capability[1]), .A5(i_cceip2_out_im_status[1]), .A6(o_cceip2_out_im_config[1]), .A7(i_cceip2_out_ia_rdata_part2[1]), .Z(n2666));
Q_MX02 U3162 ( .S(n4528), .A0(n2666), .A1(n2665), .Z(n2667));
Q_MX04 U3163 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[1]), .A1(i_cceip3_out_ia_rdata_part1[1]), .A2(i_cceip3_out_ia_rdata_part0[1]), .A3(o_cceip3_out_ia_config[1]), .Z(n2668));
Q_MX04 U3164 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[1]), .A1(i_cddip0_out_ia_capability[1]), .A2(i_cceip3_out_im_status[1]), .A3(o_cceip3_out_im_config[1]), .Z(n2669));
Q_MX04 U3165 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[1]), .A1(o_cddip0_out_ia_wdata_part2[1]), .A2(o_cddip0_out_ia_wdata_part1[1]), .A3(o_cddip0_out_ia_wdata_part0[1]), .Z(n2670));
Q_MX02 U3166 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[1]), .A1(i_cddip0_out_ia_rdata_part0[1]), .Z(n2671));
Q_AN02 U3167 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[1]), .Z(n2672));
Q_MX02 U3168 ( .S(n4526), .A0(n2672), .A1(n2671), .Z(n2673));
Q_MX04 U3169 ( .S0(n4527), .S1(n4528), .A0(n2673), .A1(n2670), .A2(n2669), .A3(n2668), .Z(n2674));
Q_MX02 U3170 ( .S(n4529), .A0(n2674), .A1(n2667), .Z(r32_mux_1_data[1]));
Q_MX04 U3171 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[2]), .A1(i_cceip2_out_ia_rdata_part0[2]), .A2(o_cceip2_out_ia_config[2]), .A3(o_cceip2_out_ia_wdata_part2[2]), .Z(n2675));
Q_MX02 U3172 ( .S(n4527), .A0(n2675), .A1(o_cceip2_out_ia_wdata_part1[2]), .Z(n2676));
Q_MX08 U3173 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[2]), .A1(o_cceip3_out_ia_wdata_part1[2]), .A2(o_cceip3_out_ia_wdata_part0[2]), .A3(i_cceip3_out_ia_status[2]), .A4(i_cceip3_out_ia_capability[2]), .A5(i_cceip2_out_im_status[2]), .A6(o_cceip2_out_im_config[2]), .A7(i_cceip2_out_ia_rdata_part2[2]), .Z(n2677));
Q_MX02 U3174 ( .S(n4528), .A0(n2677), .A1(n2676), .Z(n2678));
Q_MX04 U3175 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[2]), .A1(i_cceip3_out_ia_rdata_part1[2]), .A2(i_cceip3_out_ia_rdata_part0[2]), .A3(o_cceip3_out_ia_config[2]), .Z(n2679));
Q_MX04 U3176 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[2]), .A1(i_cddip0_out_ia_capability[2]), .A2(i_cceip3_out_im_status[2]), .A3(o_cceip3_out_im_config[2]), .Z(n2680));
Q_MX04 U3177 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[2]), .A1(o_cddip0_out_ia_wdata_part2[2]), .A2(o_cddip0_out_ia_wdata_part1[2]), .A3(o_cddip0_out_ia_wdata_part0[2]), .Z(n2681));
Q_MX02 U3178 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[2]), .A1(i_cddip0_out_ia_rdata_part0[2]), .Z(n2682));
Q_AN02 U3179 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[2]), .Z(n2683));
Q_MX02 U3180 ( .S(n4526), .A0(n2683), .A1(n2682), .Z(n2684));
Q_MX04 U3181 ( .S0(n4527), .S1(n4528), .A0(n2684), .A1(n2681), .A2(n2680), .A3(n2679), .Z(n2685));
Q_MX02 U3182 ( .S(n4529), .A0(n2685), .A1(n2678), .Z(r32_mux_1_data[2]));
Q_MX04 U3183 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[3]), .A1(i_cceip2_out_ia_rdata_part0[3]), .A2(o_cceip2_out_ia_config[3]), .A3(o_cceip2_out_ia_wdata_part2[3]), .Z(n2686));
Q_MX02 U3184 ( .S(n4527), .A0(n2686), .A1(o_cceip2_out_ia_wdata_part1[3]), .Z(n2687));
Q_MX08 U3185 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[3]), .A1(o_cceip3_out_ia_wdata_part1[3]), .A2(o_cceip3_out_ia_wdata_part0[3]), .A3(i_cceip3_out_ia_status[3]), .A4(i_cceip3_out_ia_capability[3]), .A5(i_cceip2_out_im_status[3]), .A6(o_cceip2_out_im_config[3]), .A7(i_cceip2_out_ia_rdata_part2[3]), .Z(n2688));
Q_MX02 U3186 ( .S(n4528), .A0(n2688), .A1(n2687), .Z(n2689));
Q_MX04 U3187 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[3]), .A1(i_cceip3_out_ia_rdata_part1[3]), .A2(i_cceip3_out_ia_rdata_part0[3]), .A3(o_cceip3_out_ia_config[3]), .Z(n2690));
Q_MX04 U3188 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[3]), .A1(i_cddip0_out_ia_capability[3]), .A2(i_cceip3_out_im_status[3]), .A3(o_cceip3_out_im_config[3]), .Z(n2691));
Q_MX04 U3189 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[3]), .A1(o_cddip0_out_ia_wdata_part2[3]), .A2(o_cddip0_out_ia_wdata_part1[3]), .A3(o_cddip0_out_ia_wdata_part0[3]), .Z(n2692));
Q_MX02 U3190 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[3]), .A1(i_cddip0_out_ia_rdata_part0[3]), .Z(n2693));
Q_AN02 U3191 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[3]), .Z(n2694));
Q_MX02 U3192 ( .S(n4526), .A0(n2694), .A1(n2693), .Z(n2695));
Q_MX04 U3193 ( .S0(n4527), .S1(n4528), .A0(n2695), .A1(n2692), .A2(n2691), .A3(n2690), .Z(n2696));
Q_MX02 U3194 ( .S(n4529), .A0(n2696), .A1(n2689), .Z(r32_mux_1_data[3]));
Q_MX04 U3195 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[4]), .A1(i_cceip2_out_ia_rdata_part0[4]), .A2(o_cceip2_out_ia_config[4]), .A3(o_cceip2_out_ia_wdata_part2[4]), .Z(n2697));
Q_MX02 U3196 ( .S(n4527), .A0(n2697), .A1(o_cceip2_out_ia_wdata_part1[4]), .Z(n2698));
Q_MX08 U3197 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[4]), .A1(o_cceip3_out_ia_wdata_part1[4]), .A2(o_cceip3_out_ia_wdata_part0[4]), .A3(i_cceip3_out_ia_status[4]), .A4(i_cceip3_out_ia_capability[4]), .A5(i_cceip2_out_im_status[4]), .A6(o_cceip2_out_im_config[4]), .A7(i_cceip2_out_ia_rdata_part2[4]), .Z(n2699));
Q_MX02 U3198 ( .S(n4528), .A0(n2699), .A1(n2698), .Z(n2700));
Q_MX04 U3199 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[4]), .A1(i_cceip3_out_ia_rdata_part1[4]), .A2(i_cceip3_out_ia_rdata_part0[4]), .A3(o_cceip3_out_ia_config[4]), .Z(n2701));
Q_MX04 U3200 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[4]), .A1(i_cddip0_out_ia_capability[4]), .A2(i_cceip3_out_im_status[4]), .A3(o_cceip3_out_im_config[4]), .Z(n2702));
Q_MX04 U3201 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[4]), .A1(o_cddip0_out_ia_wdata_part2[4]), .A2(o_cddip0_out_ia_wdata_part1[4]), .A3(o_cddip0_out_ia_wdata_part0[4]), .Z(n2703));
Q_MX02 U3202 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[4]), .A1(i_cddip0_out_ia_rdata_part0[4]), .Z(n2704));
Q_AN02 U3203 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[4]), .Z(n2705));
Q_MX02 U3204 ( .S(n4526), .A0(n2705), .A1(n2704), .Z(n2706));
Q_MX04 U3205 ( .S0(n4527), .S1(n4528), .A0(n2706), .A1(n2703), .A2(n2702), .A3(n2701), .Z(n2707));
Q_MX02 U3206 ( .S(n4529), .A0(n2707), .A1(n2700), .Z(r32_mux_1_data[4]));
Q_MX04 U3207 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[5]), .A1(i_cceip2_out_ia_rdata_part0[5]), .A2(o_cceip2_out_ia_config[5]), .A3(o_cceip2_out_ia_wdata_part2[5]), .Z(n2708));
Q_MX02 U3208 ( .S(n4527), .A0(n2708), .A1(o_cceip2_out_ia_wdata_part1[5]), .Z(n2709));
Q_MX08 U3209 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[5]), .A1(o_cceip3_out_ia_wdata_part1[5]), .A2(o_cceip3_out_ia_wdata_part0[5]), .A3(i_cceip3_out_ia_status[5]), .A4(i_cceip3_out_ia_capability[5]), .A5(i_cceip2_out_im_status[5]), .A6(o_cceip2_out_im_config[5]), .A7(i_cceip2_out_ia_rdata_part2[5]), .Z(n2710));
Q_MX02 U3210 ( .S(n4528), .A0(n2710), .A1(n2709), .Z(n2711));
Q_MX04 U3211 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[5]), .A1(i_cceip3_out_ia_rdata_part1[5]), .A2(i_cceip3_out_ia_rdata_part0[5]), .A3(o_cceip3_out_ia_config[5]), .Z(n2712));
Q_MX04 U3212 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[5]), .A1(i_cddip0_out_ia_capability[5]), .A2(i_cceip3_out_im_status[5]), .A3(o_cceip3_out_im_config[5]), .Z(n2713));
Q_MX04 U3213 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[5]), .A1(o_cddip0_out_ia_wdata_part2[5]), .A2(o_cddip0_out_ia_wdata_part1[5]), .A3(o_cddip0_out_ia_wdata_part0[5]), .Z(n2714));
Q_MX02 U3214 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[5]), .A1(i_cddip0_out_ia_rdata_part0[5]), .Z(n2715));
Q_AN02 U3215 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[5]), .Z(n2716));
Q_MX02 U3216 ( .S(n4526), .A0(n2716), .A1(n2715), .Z(n2717));
Q_MX04 U3217 ( .S0(n4527), .S1(n4528), .A0(n2717), .A1(n2714), .A2(n2713), .A3(n2712), .Z(n2718));
Q_MX02 U3218 ( .S(n4529), .A0(n2718), .A1(n2711), .Z(r32_mux_1_data[5]));
Q_MX04 U3219 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[6]), .A1(i_cceip2_out_ia_rdata_part0[6]), .A2(o_cceip2_out_ia_config[6]), .A3(o_cceip2_out_ia_wdata_part2[6]), .Z(n2719));
Q_MX02 U3220 ( .S(n4527), .A0(n2719), .A1(o_cceip2_out_ia_wdata_part1[6]), .Z(n2720));
Q_MX08 U3221 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[6]), .A1(o_cceip3_out_ia_wdata_part1[6]), .A2(o_cceip3_out_ia_wdata_part0[6]), .A3(i_cceip3_out_ia_status[6]), .A4(i_cceip3_out_ia_capability[6]), .A5(i_cceip2_out_im_status[6]), .A6(o_cceip2_out_im_config[6]), .A7(i_cceip2_out_ia_rdata_part2[6]), .Z(n2721));
Q_MX02 U3222 ( .S(n4528), .A0(n2721), .A1(n2720), .Z(n2722));
Q_MX04 U3223 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[6]), .A1(i_cceip3_out_ia_rdata_part1[6]), .A2(i_cceip3_out_ia_rdata_part0[6]), .A3(o_cceip3_out_ia_config[6]), .Z(n2723));
Q_MX04 U3224 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[6]), .A1(i_cddip0_out_ia_capability[6]), .A2(i_cceip3_out_im_status[6]), .A3(o_cceip3_out_im_config[6]), .Z(n2724));
Q_MX04 U3225 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[6]), .A1(o_cddip0_out_ia_wdata_part2[6]), .A2(o_cddip0_out_ia_wdata_part1[6]), .A3(o_cddip0_out_ia_wdata_part0[6]), .Z(n2725));
Q_MX02 U3226 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[6]), .A1(i_cddip0_out_ia_rdata_part0[6]), .Z(n2726));
Q_AN02 U3227 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[6]), .Z(n2727));
Q_MX02 U3228 ( .S(n4526), .A0(n2727), .A1(n2726), .Z(n2728));
Q_MX04 U3229 ( .S0(n4527), .S1(n4528), .A0(n2728), .A1(n2725), .A2(n2724), .A3(n2723), .Z(n2729));
Q_MX02 U3230 ( .S(n4529), .A0(n2729), .A1(n2722), .Z(r32_mux_1_data[6]));
Q_MX04 U3231 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[7]), .A1(i_cceip2_out_ia_rdata_part0[7]), .A2(o_cceip2_out_ia_config[7]), .A3(o_cceip2_out_ia_wdata_part2[7]), .Z(n2730));
Q_MX02 U3232 ( .S(n4527), .A0(n2730), .A1(o_cceip2_out_ia_wdata_part1[7]), .Z(n2731));
Q_MX08 U3233 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[7]), .A1(o_cceip3_out_ia_wdata_part1[7]), .A2(o_cceip3_out_ia_wdata_part0[7]), .A3(i_cceip3_out_ia_status[7]), .A4(i_cceip3_out_ia_capability[7]), .A5(i_cceip2_out_im_status[7]), .A6(o_cceip2_out_im_config[7]), .A7(i_cceip2_out_ia_rdata_part2[7]), .Z(n2732));
Q_MX02 U3234 ( .S(n4528), .A0(n2732), .A1(n2731), .Z(n2733));
Q_MX04 U3235 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[7]), .A1(i_cceip3_out_ia_rdata_part1[7]), .A2(i_cceip3_out_ia_rdata_part0[7]), .A3(o_cceip3_out_ia_config[7]), .Z(n2734));
Q_MX04 U3236 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[7]), .A1(i_cddip0_out_ia_capability[7]), .A2(i_cceip3_out_im_status[7]), .A3(o_cceip3_out_im_config[7]), .Z(n2735));
Q_MX04 U3237 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[7]), .A1(o_cddip0_out_ia_wdata_part2[7]), .A2(o_cddip0_out_ia_wdata_part1[7]), .A3(o_cddip0_out_ia_wdata_part0[7]), .Z(n2736));
Q_MX02 U3238 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[7]), .A1(i_cddip0_out_ia_rdata_part0[7]), .Z(n2737));
Q_AN02 U3239 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[7]), .Z(n2738));
Q_MX02 U3240 ( .S(n4526), .A0(n2738), .A1(n2737), .Z(n2739));
Q_MX04 U3241 ( .S0(n4527), .S1(n4528), .A0(n2739), .A1(n2736), .A2(n2735), .A3(n2734), .Z(n2740));
Q_MX02 U3242 ( .S(n4529), .A0(n2740), .A1(n2733), .Z(r32_mux_1_data[7]));
Q_MX04 U3243 ( .S0(n4525), .S1(n4526), .A0(i_cceip2_out_ia_rdata_part1[8]), .A1(i_cceip2_out_ia_rdata_part0[8]), .A2(o_cceip2_out_ia_config[8]), .A3(o_cceip2_out_ia_wdata_part2[8]), .Z(n2741));
Q_MX02 U3244 ( .S(n4527), .A0(n2741), .A1(o_cceip2_out_ia_wdata_part1[8]), .Z(n2742));
Q_MX08 U3245 ( .S0(n4525), .S1(n4526), .S2(n4527), .A0(o_cceip3_out_ia_wdata_part2[8]), .A1(o_cceip3_out_ia_wdata_part1[8]), .A2(o_cceip3_out_ia_wdata_part0[8]), .A3(i_cceip3_out_ia_status[8]), .A4(i_cceip3_out_ia_capability[8]), .A5(i_cceip2_out_im_status[8]), .A6(o_cceip2_out_im_config[8]), .A7(i_cceip2_out_ia_rdata_part2[8]), .Z(n2743));
Q_MX02 U3246 ( .S(n4528), .A0(n2743), .A1(n2742), .Z(n2744));
Q_MX04 U3247 ( .S0(n4525), .S1(n4526), .A0(i_cceip3_out_ia_rdata_part2[8]), .A1(i_cceip3_out_ia_rdata_part1[8]), .A2(i_cceip3_out_ia_rdata_part0[8]), .A3(o_cceip3_out_ia_config[8]), .Z(n2745));
Q_MX04 U3248 ( .S0(n4525), .S1(n4526), .A0(i_cddip0_out_ia_status[8]), .A1(i_cddip0_out_ia_capability[8]), .A2(i_cceip3_out_im_status[8]), .A3(o_cceip3_out_im_config[8]), .Z(n2746));
Q_MX04 U3249 ( .S0(n4525), .S1(n4526), .A0(o_cddip0_out_ia_config[8]), .A1(o_cddip0_out_ia_wdata_part2[8]), .A2(o_cddip0_out_ia_wdata_part1[8]), .A3(o_cddip0_out_ia_wdata_part0[8]), .Z(n2747));
Q_MX02 U3250 ( .S(n4525), .A0(i_cddip0_out_ia_rdata_part1[8]), .A1(i_cddip0_out_ia_rdata_part0[8]), .Z(n2748));
Q_AN02 U3251 ( .A0(n4525), .A1(i_cddip0_out_ia_rdata_part2[8]), .Z(n2749));
Q_MX02 U3252 ( .S(n4526), .A0(n2749), .A1(n2748), .Z(n2750));
Q_MX04 U3253 ( .S0(n4527), .S1(n4528), .A0(n2750), .A1(n2747), .A2(n2746), .A3(n2745), .Z(n2751));
Q_MX02 U3254 ( .S(n4529), .A0(n2751), .A1(n2744), .Z(r32_mux_1_data[8]));
Q_MX02 U3255 ( .S(n4530), .A0(o_cceip2_out_ia_wdata_part2[9]), .A1(o_cceip2_out_ia_wdata_part1[9]), .Z(n2752));
Q_MX04 U3256 ( .S0(n4530), .S1(n4531), .A0(o_cceip2_out_im_config[9]), .A1(i_cceip2_out_ia_rdata_part2[9]), .A2(i_cceip2_out_ia_rdata_part1[9]), .A3(i_cceip2_out_ia_rdata_part0[9]), .Z(n2753));
Q_MX02 U3257 ( .S(n4532), .A0(n2753), .A1(n2752), .Z(n2754));
Q_MX04 U3258 ( .S0(n4530), .S1(n4531), .A0(o_cceip3_out_ia_wdata_part2[9]), .A1(o_cceip3_out_ia_wdata_part1[9]), .A2(o_cceip3_out_ia_wdata_part0[9]), .A3(i_cceip3_out_ia_capability[9]), .Z(n2755));
Q_MX04 U3259 ( .S0(n4530), .S1(n4531), .A0(o_cceip3_out_im_config[9]), .A1(i_cceip3_out_ia_rdata_part2[9]), .A2(i_cceip3_out_ia_rdata_part1[9]), .A3(i_cceip3_out_ia_rdata_part0[9]), .Z(n2756));
Q_MX04 U3260 ( .S0(n4530), .S1(n4531), .A0(o_cddip0_out_ia_wdata_part2[9]), .A1(o_cddip0_out_ia_wdata_part1[9]), .A2(o_cddip0_out_ia_wdata_part0[9]), .A3(i_cddip0_out_ia_capability[9]), .Z(n2757));
Q_MX02 U3261 ( .S(n4530), .A0(i_cddip0_out_ia_rdata_part1[9]), .A1(i_cddip0_out_ia_rdata_part0[9]), .Z(n2758));
Q_AN02 U3262 ( .A0(n4530), .A1(i_cddip0_out_ia_rdata_part2[9]), .Z(n2759));
Q_MX02 U3263 ( .S(n4531), .A0(n2759), .A1(n2758), .Z(n2760));
Q_MX04 U3264 ( .S0(n4532), .S1(n4533), .A0(n2760), .A1(n2757), .A2(n2756), .A3(n2755), .Z(n2761));
Q_MX02 U3265 ( .S(n4534), .A0(n2761), .A1(n2754), .Z(r32_mux_1_data[9]));
Q_MX04 U3266 ( .S0(n4535), .S1(n4536), .A0(i_cceip2_out_ia_rdata_part1[10]), .A1(i_cceip2_out_ia_rdata_part0[10]), .A2(o_cceip2_out_ia_wdata_part2[10]), .A3(o_cceip2_out_ia_wdata_part1[10]), .Z(n2762));
Q_MX04 U3267 ( .S0(n4535), .S1(n4536), .A0(o_cceip3_out_ia_wdata_part1[10]), .A1(o_cceip3_out_ia_wdata_part0[10]), .A2(i_cceip3_out_ia_capability[10]), .A3(i_cceip2_out_ia_rdata_part2[10]), .Z(n2763));
Q_MX04 U3268 ( .S0(n4535), .S1(n4536), .A0(i_cceip3_out_ia_rdata_part2[10]), .A1(i_cceip3_out_ia_rdata_part1[10]), .A2(i_cceip3_out_ia_rdata_part0[10]), .A3(o_cceip3_out_ia_wdata_part2[10]), .Z(n2764));
Q_MX04 U3269 ( .S0(n4535), .S1(n4536), .A0(o_cddip0_out_ia_wdata_part2[10]), .A1(o_cddip0_out_ia_wdata_part1[10]), .A2(o_cddip0_out_ia_wdata_part0[10]), .A3(i_cddip0_out_ia_capability[10]), .Z(n2765));
Q_MX02 U3270 ( .S(n4535), .A0(i_cddip0_out_ia_rdata_part1[10]), .A1(i_cddip0_out_ia_rdata_part0[10]), .Z(n2766));
Q_AN02 U3271 ( .A0(n4535), .A1(i_cddip0_out_ia_rdata_part2[10]), .Z(n2767));
Q_MX02 U3272 ( .S(n4536), .A0(n2767), .A1(n2766), .Z(n2768));
Q_MX04 U3273 ( .S0(n4537), .S1(n4538), .A0(n2768), .A1(n2765), .A2(n2764), .A3(n2763), .Z(n2769));
Q_MX02 U3274 ( .S(n4539), .A0(n2769), .A1(n2762), .Z(r32_mux_1_data[10]));
Q_MX04 U3275 ( .S0(n4535), .S1(n4536), .A0(i_cceip2_out_ia_rdata_part1[11]), .A1(i_cceip2_out_ia_rdata_part0[11]), .A2(o_cceip2_out_ia_wdata_part2[11]), .A3(o_cceip2_out_ia_wdata_part1[11]), .Z(n2770));
Q_MX04 U3276 ( .S0(n4535), .S1(n4536), .A0(o_cceip3_out_ia_wdata_part1[11]), .A1(o_cceip3_out_ia_wdata_part0[11]), .A2(i_cceip3_out_ia_capability[11]), .A3(i_cceip2_out_ia_rdata_part2[11]), .Z(n2771));
Q_MX04 U3277 ( .S0(n4535), .S1(n4536), .A0(i_cceip3_out_ia_rdata_part2[11]), .A1(i_cceip3_out_ia_rdata_part1[11]), .A2(i_cceip3_out_ia_rdata_part0[11]), .A3(o_cceip3_out_ia_wdata_part2[11]), .Z(n2772));
Q_MX04 U3278 ( .S0(n4535), .S1(n4536), .A0(o_cddip0_out_ia_wdata_part2[11]), .A1(o_cddip0_out_ia_wdata_part1[11]), .A2(o_cddip0_out_ia_wdata_part0[11]), .A3(i_cddip0_out_ia_capability[11]), .Z(n2773));
Q_MX02 U3279 ( .S(n4535), .A0(i_cddip0_out_ia_rdata_part1[11]), .A1(i_cddip0_out_ia_rdata_part0[11]), .Z(n2774));
Q_AN02 U3280 ( .A0(n4535), .A1(i_cddip0_out_ia_rdata_part2[11]), .Z(n2775));
Q_MX02 U3281 ( .S(n4536), .A0(n2775), .A1(n2774), .Z(n2776));
Q_MX04 U3282 ( .S0(n4537), .S1(n4538), .A0(n2776), .A1(n2773), .A2(n2772), .A3(n2771), .Z(n2777));
Q_MX02 U3283 ( .S(n4539), .A0(n2777), .A1(n2770), .Z(r32_mux_1_data[11]));
Q_MX04 U3284 ( .S0(n4535), .S1(n4536), .A0(i_cceip2_out_ia_rdata_part1[12]), .A1(i_cceip2_out_ia_rdata_part0[12]), .A2(o_cceip2_out_ia_wdata_part2[12]), .A3(o_cceip2_out_ia_wdata_part1[12]), .Z(n2778));
Q_MX04 U3285 ( .S0(n4535), .S1(n4536), .A0(o_cceip3_out_ia_wdata_part1[12]), .A1(o_cceip3_out_ia_wdata_part0[12]), .A2(i_cceip3_out_ia_capability[12]), .A3(i_cceip2_out_ia_rdata_part2[12]), .Z(n2779));
Q_MX04 U3286 ( .S0(n4535), .S1(n4536), .A0(i_cceip3_out_ia_rdata_part2[12]), .A1(i_cceip3_out_ia_rdata_part1[12]), .A2(i_cceip3_out_ia_rdata_part0[12]), .A3(o_cceip3_out_ia_wdata_part2[12]), .Z(n2780));
Q_MX04 U3287 ( .S0(n4535), .S1(n4536), .A0(o_cddip0_out_ia_wdata_part2[12]), .A1(o_cddip0_out_ia_wdata_part1[12]), .A2(o_cddip0_out_ia_wdata_part0[12]), .A3(i_cddip0_out_ia_capability[12]), .Z(n2781));
Q_MX02 U3288 ( .S(n4535), .A0(i_cddip0_out_ia_rdata_part1[12]), .A1(i_cddip0_out_ia_rdata_part0[12]), .Z(n2782));
Q_AN02 U3289 ( .A0(n4535), .A1(i_cddip0_out_ia_rdata_part2[12]), .Z(n2783));
Q_MX02 U3290 ( .S(n4536), .A0(n2783), .A1(n2782), .Z(n2784));
Q_MX04 U3291 ( .S0(n4537), .S1(n4538), .A0(n2784), .A1(n2781), .A2(n2780), .A3(n2779), .Z(n2785));
Q_MX02 U3292 ( .S(n4539), .A0(n2785), .A1(n2778), .Z(r32_mux_1_data[12]));
Q_MX04 U3293 ( .S0(n4535), .S1(n4536), .A0(i_cceip2_out_ia_rdata_part1[13]), .A1(i_cceip2_out_ia_rdata_part0[13]), .A2(o_cceip2_out_ia_wdata_part2[13]), .A3(o_cceip2_out_ia_wdata_part1[13]), .Z(n2786));
Q_MX04 U3294 ( .S0(n4535), .S1(n4536), .A0(o_cceip3_out_ia_wdata_part1[13]), .A1(o_cceip3_out_ia_wdata_part0[13]), .A2(i_cceip3_out_ia_capability[13]), .A3(i_cceip2_out_ia_rdata_part2[13]), .Z(n2787));
Q_MX04 U3295 ( .S0(n4535), .S1(n4536), .A0(i_cceip3_out_ia_rdata_part2[13]), .A1(i_cceip3_out_ia_rdata_part1[13]), .A2(i_cceip3_out_ia_rdata_part0[13]), .A3(o_cceip3_out_ia_wdata_part2[13]), .Z(n2788));
Q_MX04 U3296 ( .S0(n4535), .S1(n4536), .A0(o_cddip0_out_ia_wdata_part2[13]), .A1(o_cddip0_out_ia_wdata_part1[13]), .A2(o_cddip0_out_ia_wdata_part0[13]), .A3(i_cddip0_out_ia_capability[13]), .Z(n2789));
Q_MX02 U3297 ( .S(n4535), .A0(i_cddip0_out_ia_rdata_part1[13]), .A1(i_cddip0_out_ia_rdata_part0[13]), .Z(n2790));
Q_AN02 U3298 ( .A0(n4535), .A1(i_cddip0_out_ia_rdata_part2[13]), .Z(n2791));
Q_MX02 U3299 ( .S(n4536), .A0(n2791), .A1(n2790), .Z(n2792));
Q_MX04 U3300 ( .S0(n4537), .S1(n4538), .A0(n2792), .A1(n2789), .A2(n2788), .A3(n2787), .Z(n2793));
Q_MX02 U3301 ( .S(n4539), .A0(n2793), .A1(n2786), .Z(r32_mux_1_data[13]));
Q_MX04 U3302 ( .S0(n4535), .S1(n4536), .A0(i_cceip2_out_ia_rdata_part1[14]), .A1(i_cceip2_out_ia_rdata_part0[14]), .A2(o_cceip2_out_ia_wdata_part2[14]), .A3(o_cceip2_out_ia_wdata_part1[14]), .Z(n2794));
Q_MX04 U3303 ( .S0(n4535), .S1(n4536), .A0(o_cceip3_out_ia_wdata_part1[14]), .A1(o_cceip3_out_ia_wdata_part0[14]), .A2(i_cceip3_out_ia_capability[14]), .A3(i_cceip2_out_ia_rdata_part2[14]), .Z(n2795));
Q_MX04 U3304 ( .S0(n4535), .S1(n4536), .A0(i_cceip3_out_ia_rdata_part2[14]), .A1(i_cceip3_out_ia_rdata_part1[14]), .A2(i_cceip3_out_ia_rdata_part0[14]), .A3(o_cceip3_out_ia_wdata_part2[14]), .Z(n2796));
Q_MX04 U3305 ( .S0(n4535), .S1(n4536), .A0(o_cddip0_out_ia_wdata_part2[14]), .A1(o_cddip0_out_ia_wdata_part1[14]), .A2(o_cddip0_out_ia_wdata_part0[14]), .A3(i_cddip0_out_ia_capability[14]), .Z(n2797));
Q_MX02 U3306 ( .S(n4535), .A0(i_cddip0_out_ia_rdata_part1[14]), .A1(i_cddip0_out_ia_rdata_part0[14]), .Z(n2798));
Q_AN02 U3307 ( .A0(n4535), .A1(i_cddip0_out_ia_rdata_part2[14]), .Z(n2799));
Q_MX02 U3308 ( .S(n4536), .A0(n2799), .A1(n2798), .Z(n2800));
Q_MX04 U3309 ( .S0(n4537), .S1(n4538), .A0(n2800), .A1(n2797), .A2(n2796), .A3(n2795), .Z(n2801));
Q_MX02 U3310 ( .S(n4539), .A0(n2801), .A1(n2794), .Z(r32_mux_1_data[14]));
Q_MX04 U3311 ( .S0(n4535), .S1(n4536), .A0(i_cceip2_out_ia_rdata_part1[15]), .A1(i_cceip2_out_ia_rdata_part0[15]), .A2(o_cceip2_out_ia_wdata_part2[15]), .A3(o_cceip2_out_ia_wdata_part1[15]), .Z(n2802));
Q_MX04 U3312 ( .S0(n4535), .S1(n4536), .A0(o_cceip3_out_ia_wdata_part1[15]), .A1(o_cceip3_out_ia_wdata_part0[15]), .A2(i_cceip3_out_ia_capability[15]), .A3(i_cceip2_out_ia_rdata_part2[15]), .Z(n2803));
Q_MX04 U3313 ( .S0(n4535), .S1(n4536), .A0(i_cceip3_out_ia_rdata_part2[15]), .A1(i_cceip3_out_ia_rdata_part1[15]), .A2(i_cceip3_out_ia_rdata_part0[15]), .A3(o_cceip3_out_ia_wdata_part2[15]), .Z(n2804));
Q_MX04 U3314 ( .S0(n4535), .S1(n4536), .A0(o_cddip0_out_ia_wdata_part2[15]), .A1(o_cddip0_out_ia_wdata_part1[15]), .A2(o_cddip0_out_ia_wdata_part0[15]), .A3(i_cddip0_out_ia_capability[15]), .Z(n2805));
Q_MX02 U3315 ( .S(n4535), .A0(i_cddip0_out_ia_rdata_part1[15]), .A1(i_cddip0_out_ia_rdata_part0[15]), .Z(n2806));
Q_AN02 U3316 ( .A0(n4535), .A1(i_cddip0_out_ia_rdata_part2[15]), .Z(n2807));
Q_MX02 U3317 ( .S(n4536), .A0(n2807), .A1(n2806), .Z(n2808));
Q_MX04 U3318 ( .S0(n4537), .S1(n4538), .A0(n2808), .A1(n2805), .A2(n2804), .A3(n2803), .Z(n2809));
Q_MX02 U3319 ( .S(n4539), .A0(n2809), .A1(n2802), .Z(r32_mux_1_data[15]));
Q_MX02 U3320 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[16]), .A1(o_cceip2_out_ia_wdata_part1[16]), .Z(n2810));
Q_MX04 U3321 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[16]), .A1(i_cceip2_out_ia_rdata_part2[16]), .A2(i_cceip2_out_ia_rdata_part1[16]), .A3(i_cceip2_out_ia_rdata_part0[16]), .Z(n2811));
Q_MX04 U3322 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[16]), .A1(i_cceip3_out_ia_rdata_part0[16]), .A2(o_cceip3_out_ia_wdata_part2[16]), .A3(o_cceip3_out_ia_wdata_part1[16]), .Z(n2812));
Q_MX04 U3323 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[16]), .A1(o_cddip0_out_ia_wdata_part1[16]), .A2(o_cddip0_out_ia_wdata_part0[16]), .A3(i_cceip3_out_ia_rdata_part2[16]), .Z(n2813));
Q_MX02 U3324 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[16]), .A1(i_cddip0_out_ia_rdata_part0[16]), .Z(n2814));
Q_AN02 U3325 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[16]), .Z(n2815));
Q_MX02 U3326 ( .S(n4541), .A0(n2815), .A1(n2814), .Z(n2816));
Q_MX04 U3327 ( .S0(n4542), .S1(n4543), .A0(n2816), .A1(n2813), .A2(n2812), .A3(n2811), .Z(n2817));
Q_MX02 U3328 ( .S(n4544), .A0(n2817), .A1(n2810), .Z(r32_mux_1_data[16]));
Q_MX02 U3329 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[17]), .A1(o_cceip2_out_ia_wdata_part1[17]), .Z(n2818));
Q_MX04 U3330 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[17]), .A1(i_cceip2_out_ia_rdata_part2[17]), .A2(i_cceip2_out_ia_rdata_part1[17]), .A3(i_cceip2_out_ia_rdata_part0[17]), .Z(n2819));
Q_MX04 U3331 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[17]), .A1(i_cceip3_out_ia_rdata_part0[17]), .A2(o_cceip3_out_ia_wdata_part2[17]), .A3(o_cceip3_out_ia_wdata_part1[17]), .Z(n2820));
Q_MX04 U3332 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[17]), .A1(o_cddip0_out_ia_wdata_part1[17]), .A2(o_cddip0_out_ia_wdata_part0[17]), .A3(i_cceip3_out_ia_rdata_part2[17]), .Z(n2821));
Q_MX02 U3333 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[17]), .A1(i_cddip0_out_ia_rdata_part0[17]), .Z(n2822));
Q_AN02 U3334 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[17]), .Z(n2823));
Q_MX02 U3335 ( .S(n4541), .A0(n2823), .A1(n2822), .Z(n2824));
Q_MX04 U3336 ( .S0(n4542), .S1(n4543), .A0(n2824), .A1(n2821), .A2(n2820), .A3(n2819), .Z(n2825));
Q_MX02 U3337 ( .S(n4544), .A0(n2825), .A1(n2818), .Z(r32_mux_1_data[17]));
Q_MX02 U3338 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[18]), .A1(o_cceip2_out_ia_wdata_part1[18]), .Z(n2826));
Q_MX04 U3339 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[18]), .A1(i_cceip2_out_ia_rdata_part2[18]), .A2(i_cceip2_out_ia_rdata_part1[18]), .A3(i_cceip2_out_ia_rdata_part0[18]), .Z(n2827));
Q_MX04 U3340 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[18]), .A1(i_cceip3_out_ia_rdata_part0[18]), .A2(o_cceip3_out_ia_wdata_part2[18]), .A3(o_cceip3_out_ia_wdata_part1[18]), .Z(n2828));
Q_MX04 U3341 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[18]), .A1(o_cddip0_out_ia_wdata_part1[18]), .A2(o_cddip0_out_ia_wdata_part0[18]), .A3(i_cceip3_out_ia_rdata_part2[18]), .Z(n2829));
Q_MX02 U3342 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[18]), .A1(i_cddip0_out_ia_rdata_part0[18]), .Z(n2830));
Q_AN02 U3343 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[18]), .Z(n2831));
Q_MX02 U3344 ( .S(n4541), .A0(n2831), .A1(n2830), .Z(n2832));
Q_MX04 U3345 ( .S0(n4542), .S1(n4543), .A0(n2832), .A1(n2829), .A2(n2828), .A3(n2827), .Z(n2833));
Q_MX02 U3346 ( .S(n4544), .A0(n2833), .A1(n2826), .Z(r32_mux_1_data[18]));
Q_MX02 U3347 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[19]), .A1(o_cceip2_out_ia_wdata_part1[19]), .Z(n2834));
Q_MX04 U3348 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[19]), .A1(i_cceip2_out_ia_rdata_part2[19]), .A2(i_cceip2_out_ia_rdata_part1[19]), .A3(i_cceip2_out_ia_rdata_part0[19]), .Z(n2835));
Q_MX04 U3349 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[19]), .A1(i_cceip3_out_ia_rdata_part0[19]), .A2(o_cceip3_out_ia_wdata_part2[19]), .A3(o_cceip3_out_ia_wdata_part1[19]), .Z(n2836));
Q_MX04 U3350 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[19]), .A1(o_cddip0_out_ia_wdata_part1[19]), .A2(o_cddip0_out_ia_wdata_part0[19]), .A3(i_cceip3_out_ia_rdata_part2[19]), .Z(n2837));
Q_MX02 U3351 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[19]), .A1(i_cddip0_out_ia_rdata_part0[19]), .Z(n2838));
Q_AN02 U3352 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[19]), .Z(n2839));
Q_MX02 U3353 ( .S(n4541), .A0(n2839), .A1(n2838), .Z(n2840));
Q_MX04 U3354 ( .S0(n4542), .S1(n4543), .A0(n2840), .A1(n2837), .A2(n2836), .A3(n2835), .Z(n2841));
Q_MX02 U3355 ( .S(n4544), .A0(n2841), .A1(n2834), .Z(r32_mux_1_data[19]));
Q_MX02 U3356 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[20]), .A1(o_cceip2_out_ia_wdata_part1[20]), .Z(n2842));
Q_MX04 U3357 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[20]), .A1(i_cceip2_out_ia_rdata_part2[20]), .A2(i_cceip2_out_ia_rdata_part1[20]), .A3(i_cceip2_out_ia_rdata_part0[20]), .Z(n2843));
Q_MX04 U3358 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[20]), .A1(i_cceip3_out_ia_rdata_part0[20]), .A2(o_cceip3_out_ia_wdata_part2[20]), .A3(o_cceip3_out_ia_wdata_part1[20]), .Z(n2844));
Q_MX04 U3359 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[20]), .A1(o_cddip0_out_ia_wdata_part1[20]), .A2(o_cddip0_out_ia_wdata_part0[20]), .A3(i_cceip3_out_ia_rdata_part2[20]), .Z(n2845));
Q_MX02 U3360 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[20]), .A1(i_cddip0_out_ia_rdata_part0[20]), .Z(n2846));
Q_AN02 U3361 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[20]), .Z(n2847));
Q_MX02 U3362 ( .S(n4541), .A0(n2847), .A1(n2846), .Z(n2848));
Q_MX04 U3363 ( .S0(n4542), .S1(n4543), .A0(n2848), .A1(n2845), .A2(n2844), .A3(n2843), .Z(n2849));
Q_MX02 U3364 ( .S(n4544), .A0(n2849), .A1(n2842), .Z(r32_mux_1_data[20]));
Q_MX02 U3365 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[21]), .A1(o_cceip2_out_ia_wdata_part1[21]), .Z(n2850));
Q_MX04 U3366 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[21]), .A1(i_cceip2_out_ia_rdata_part2[21]), .A2(i_cceip2_out_ia_rdata_part1[21]), .A3(i_cceip2_out_ia_rdata_part0[21]), .Z(n2851));
Q_MX04 U3367 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[21]), .A1(i_cceip3_out_ia_rdata_part0[21]), .A2(o_cceip3_out_ia_wdata_part2[21]), .A3(o_cceip3_out_ia_wdata_part1[21]), .Z(n2852));
Q_MX04 U3368 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[21]), .A1(o_cddip0_out_ia_wdata_part1[21]), .A2(o_cddip0_out_ia_wdata_part0[21]), .A3(i_cceip3_out_ia_rdata_part2[21]), .Z(n2853));
Q_MX02 U3369 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[21]), .A1(i_cddip0_out_ia_rdata_part0[21]), .Z(n2854));
Q_AN02 U3370 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[21]), .Z(n2855));
Q_MX02 U3371 ( .S(n4541), .A0(n2855), .A1(n2854), .Z(n2856));
Q_MX04 U3372 ( .S0(n4542), .S1(n4543), .A0(n2856), .A1(n2853), .A2(n2852), .A3(n2851), .Z(n2857));
Q_MX02 U3373 ( .S(n4544), .A0(n2857), .A1(n2850), .Z(r32_mux_1_data[21]));
Q_MX02 U3374 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[22]), .A1(o_cceip2_out_ia_wdata_part1[22]), .Z(n2858));
Q_MX04 U3375 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[22]), .A1(i_cceip2_out_ia_rdata_part2[22]), .A2(i_cceip2_out_ia_rdata_part1[22]), .A3(i_cceip2_out_ia_rdata_part0[22]), .Z(n2859));
Q_MX04 U3376 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[22]), .A1(i_cceip3_out_ia_rdata_part0[22]), .A2(o_cceip3_out_ia_wdata_part2[22]), .A3(o_cceip3_out_ia_wdata_part1[22]), .Z(n2860));
Q_MX04 U3377 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[22]), .A1(o_cddip0_out_ia_wdata_part1[22]), .A2(o_cddip0_out_ia_wdata_part0[22]), .A3(i_cceip3_out_ia_rdata_part2[22]), .Z(n2861));
Q_MX02 U3378 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[22]), .A1(i_cddip0_out_ia_rdata_part0[22]), .Z(n2862));
Q_AN02 U3379 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[22]), .Z(n2863));
Q_MX02 U3380 ( .S(n4541), .A0(n2863), .A1(n2862), .Z(n2864));
Q_MX04 U3381 ( .S0(n4542), .S1(n4543), .A0(n2864), .A1(n2861), .A2(n2860), .A3(n2859), .Z(n2865));
Q_MX02 U3382 ( .S(n4544), .A0(n2865), .A1(n2858), .Z(r32_mux_1_data[22]));
Q_MX02 U3383 ( .S(n4540), .A0(o_cceip2_out_ia_wdata_part2[23]), .A1(o_cceip2_out_ia_wdata_part1[23]), .Z(n2866));
Q_MX04 U3384 ( .S0(n4540), .S1(n4541), .A0(o_cceip3_out_ia_wdata_part0[23]), .A1(i_cceip2_out_ia_rdata_part2[23]), .A2(i_cceip2_out_ia_rdata_part1[23]), .A3(i_cceip2_out_ia_rdata_part0[23]), .Z(n2867));
Q_MX04 U3385 ( .S0(n4540), .S1(n4541), .A0(i_cceip3_out_ia_rdata_part1[23]), .A1(i_cceip3_out_ia_rdata_part0[23]), .A2(o_cceip3_out_ia_wdata_part2[23]), .A3(o_cceip3_out_ia_wdata_part1[23]), .Z(n2868));
Q_MX04 U3386 ( .S0(n4540), .S1(n4541), .A0(o_cddip0_out_ia_wdata_part2[23]), .A1(o_cddip0_out_ia_wdata_part1[23]), .A2(o_cddip0_out_ia_wdata_part0[23]), .A3(i_cceip3_out_ia_rdata_part2[23]), .Z(n2869));
Q_MX02 U3387 ( .S(n4540), .A0(i_cddip0_out_ia_rdata_part1[23]), .A1(i_cddip0_out_ia_rdata_part0[23]), .Z(n2870));
Q_AN02 U3388 ( .A0(n4540), .A1(i_cddip0_out_ia_rdata_part2[23]), .Z(n2871));
Q_MX02 U3389 ( .S(n4541), .A0(n2871), .A1(n2870), .Z(n2872));
Q_MX04 U3390 ( .S0(n4542), .S1(n4543), .A0(n2872), .A1(n2869), .A2(n2868), .A3(n2867), .Z(n2873));
Q_MX02 U3391 ( .S(n4544), .A0(n2873), .A1(n2866), .Z(r32_mux_1_data[23]));
Q_MX04 U3392 ( .S0(n4545), .S1(n4546), .A0(i_cceip2_out_ia_rdata_part1[24]), .A1(i_cceip2_out_ia_rdata_part0[24]), .A2(o_cceip2_out_ia_wdata_part2[24]), .A3(o_cceip2_out_ia_wdata_part1[24]), .Z(n2874));
Q_MX04 U3393 ( .S0(n4545), .S1(n4546), .A0(o_cceip3_out_ia_wdata_part1[24]), .A1(o_cceip3_out_ia_wdata_part0[24]), .A2(i_cceip3_out_ia_status[9]), .A3(i_cceip2_out_ia_rdata_part2[24]), .Z(n2875));
Q_MX04 U3394 ( .S0(n4545), .S1(n4546), .A0(i_cceip3_out_ia_rdata_part2[24]), .A1(i_cceip3_out_ia_rdata_part1[24]), .A2(i_cceip3_out_ia_rdata_part0[24]), .A3(o_cceip3_out_ia_wdata_part2[24]), .Z(n2876));
Q_MX04 U3395 ( .S0(n4545), .S1(n4546), .A0(o_cddip0_out_ia_wdata_part2[24]), .A1(o_cddip0_out_ia_wdata_part1[24]), .A2(o_cddip0_out_ia_wdata_part0[24]), .A3(i_cddip0_out_ia_status[9]), .Z(n2877));
Q_MX02 U3396 ( .S(n4545), .A0(i_cddip0_out_ia_rdata_part1[24]), .A1(i_cddip0_out_ia_rdata_part0[24]), .Z(n2878));
Q_AN02 U3397 ( .A0(n4545), .A1(i_cddip0_out_ia_rdata_part2[24]), .Z(n2879));
Q_MX02 U3398 ( .S(n4546), .A0(n2879), .A1(n2878), .Z(n2880));
Q_MX04 U3399 ( .S0(n4547), .S1(n4548), .A0(n2880), .A1(n2877), .A2(n2876), .A3(n2875), .Z(n2881));
Q_MX02 U3400 ( .S(n4539), .A0(n2881), .A1(n2874), .Z(r32_mux_1_data[24]));
Q_MX04 U3401 ( .S0(n4545), .S1(n4546), .A0(i_cceip2_out_ia_rdata_part1[25]), .A1(i_cceip2_out_ia_rdata_part0[25]), .A2(o_cceip2_out_ia_wdata_part2[25]), .A3(o_cceip2_out_ia_wdata_part1[25]), .Z(n2882));
Q_MX04 U3402 ( .S0(n4545), .S1(n4546), .A0(o_cceip3_out_ia_wdata_part1[25]), .A1(o_cceip3_out_ia_wdata_part0[25]), .A2(i_cceip3_out_ia_status[10]), .A3(i_cceip2_out_ia_rdata_part2[25]), .Z(n2883));
Q_MX04 U3403 ( .S0(n4545), .S1(n4546), .A0(i_cceip3_out_ia_rdata_part2[25]), .A1(i_cceip3_out_ia_rdata_part1[25]), .A2(i_cceip3_out_ia_rdata_part0[25]), .A3(o_cceip3_out_ia_wdata_part2[25]), .Z(n2884));
Q_MX04 U3404 ( .S0(n4545), .S1(n4546), .A0(o_cddip0_out_ia_wdata_part2[25]), .A1(o_cddip0_out_ia_wdata_part1[25]), .A2(o_cddip0_out_ia_wdata_part0[25]), .A3(i_cddip0_out_ia_status[10]), .Z(n2885));
Q_MX02 U3405 ( .S(n4545), .A0(i_cddip0_out_ia_rdata_part1[25]), .A1(i_cddip0_out_ia_rdata_part0[25]), .Z(n2886));
Q_AN02 U3406 ( .A0(n4545), .A1(i_cddip0_out_ia_rdata_part2[25]), .Z(n2887));
Q_MX02 U3407 ( .S(n4546), .A0(n2887), .A1(n2886), .Z(n2888));
Q_MX04 U3408 ( .S0(n4547), .S1(n4548), .A0(n2888), .A1(n2885), .A2(n2884), .A3(n2883), .Z(n2889));
Q_MX02 U3409 ( .S(n4539), .A0(n2889), .A1(n2882), .Z(r32_mux_1_data[25]));
Q_MX04 U3410 ( .S0(n4545), .S1(n4546), .A0(i_cceip2_out_ia_rdata_part1[26]), .A1(i_cceip2_out_ia_rdata_part0[26]), .A2(o_cceip2_out_ia_wdata_part2[26]), .A3(o_cceip2_out_ia_wdata_part1[26]), .Z(n2890));
Q_MX04 U3411 ( .S0(n4545), .S1(n4546), .A0(o_cceip3_out_ia_wdata_part1[26]), .A1(o_cceip3_out_ia_wdata_part0[26]), .A2(i_cceip3_out_ia_status[11]), .A3(i_cceip2_out_ia_rdata_part2[26]), .Z(n2891));
Q_MX04 U3412 ( .S0(n4545), .S1(n4546), .A0(i_cceip3_out_ia_rdata_part2[26]), .A1(i_cceip3_out_ia_rdata_part1[26]), .A2(i_cceip3_out_ia_rdata_part0[26]), .A3(o_cceip3_out_ia_wdata_part2[26]), .Z(n2892));
Q_MX04 U3413 ( .S0(n4545), .S1(n4546), .A0(o_cddip0_out_ia_wdata_part2[26]), .A1(o_cddip0_out_ia_wdata_part1[26]), .A2(o_cddip0_out_ia_wdata_part0[26]), .A3(i_cddip0_out_ia_status[11]), .Z(n2893));
Q_MX02 U3414 ( .S(n4545), .A0(i_cddip0_out_ia_rdata_part1[26]), .A1(i_cddip0_out_ia_rdata_part0[26]), .Z(n2894));
Q_AN02 U3415 ( .A0(n4545), .A1(i_cddip0_out_ia_rdata_part2[26]), .Z(n2895));
Q_MX02 U3416 ( .S(n4546), .A0(n2895), .A1(n2894), .Z(n2896));
Q_MX04 U3417 ( .S0(n4547), .S1(n4548), .A0(n2896), .A1(n2893), .A2(n2892), .A3(n2891), .Z(n2897));
Q_MX02 U3418 ( .S(n4539), .A0(n2897), .A1(n2890), .Z(r32_mux_1_data[26]));
Q_MX04 U3419 ( .S0(n4545), .S1(n4546), .A0(i_cceip2_out_ia_rdata_part1[27]), .A1(i_cceip2_out_ia_rdata_part0[27]), .A2(o_cceip2_out_ia_wdata_part2[27]), .A3(o_cceip2_out_ia_wdata_part1[27]), .Z(n2898));
Q_MX04 U3420 ( .S0(n4545), .S1(n4546), .A0(o_cceip3_out_ia_wdata_part1[27]), .A1(o_cceip3_out_ia_wdata_part0[27]), .A2(i_cceip3_out_ia_status[12]), .A3(i_cceip2_out_ia_rdata_part2[27]), .Z(n2899));
Q_MX04 U3421 ( .S0(n4545), .S1(n4546), .A0(i_cceip3_out_ia_rdata_part2[27]), .A1(i_cceip3_out_ia_rdata_part1[27]), .A2(i_cceip3_out_ia_rdata_part0[27]), .A3(o_cceip3_out_ia_wdata_part2[27]), .Z(n2900));
Q_MX04 U3422 ( .S0(n4545), .S1(n4546), .A0(o_cddip0_out_ia_wdata_part2[27]), .A1(o_cddip0_out_ia_wdata_part1[27]), .A2(o_cddip0_out_ia_wdata_part0[27]), .A3(i_cddip0_out_ia_status[12]), .Z(n2901));
Q_MX02 U3423 ( .S(n4545), .A0(i_cddip0_out_ia_rdata_part1[27]), .A1(i_cddip0_out_ia_rdata_part0[27]), .Z(n2902));
Q_AN02 U3424 ( .A0(n4545), .A1(i_cddip0_out_ia_rdata_part2[27]), .Z(n2903));
Q_MX02 U3425 ( .S(n4546), .A0(n2903), .A1(n2902), .Z(n2904));
Q_MX04 U3426 ( .S0(n4547), .S1(n4548), .A0(n2904), .A1(n2901), .A2(n2900), .A3(n2899), .Z(n2905));
Q_MX02 U3427 ( .S(n4539), .A0(n2905), .A1(n2898), .Z(r32_mux_1_data[27]));
Q_MX08 U3428 ( .S0(n4549), .S1(n4550), .S2(n4551), .A0(o_cceip3_out_ia_wdata_part0[28]), .A1(i_cceip3_out_ia_status[13]), .A2(i_cceip3_out_ia_capability[16]), .A3(i_cceip2_out_ia_rdata_part2[28]), .A4(i_cceip2_out_ia_rdata_part1[28]), .A5(i_cceip2_out_ia_rdata_part0[28]), .A6(o_cceip2_out_ia_config[9]), .A7(o_cceip2_out_ia_wdata_part2[28]), .Z(n2906));
Q_MX02 U3429 ( .S(n4552), .A0(n2906), .A1(o_cceip2_out_ia_wdata_part1[28]), .Z(n2907));
Q_MX04 U3430 ( .S0(n4549), .S1(n4550), .A0(i_cceip3_out_ia_rdata_part0[28]), .A1(o_cceip3_out_ia_config[9]), .A2(o_cceip3_out_ia_wdata_part2[28]), .A3(o_cceip3_out_ia_wdata_part1[28]), .Z(n2908));
Q_MX04 U3431 ( .S0(n4549), .S1(n4550), .A0(i_cddip0_out_ia_status[13]), .A1(i_cddip0_out_ia_capability[16]), .A2(i_cceip3_out_ia_rdata_part2[28]), .A3(i_cceip3_out_ia_rdata_part1[28]), .Z(n2909));
Q_MX04 U3432 ( .S0(n4549), .S1(n4550), .A0(o_cddip0_out_ia_config[9]), .A1(o_cddip0_out_ia_wdata_part2[28]), .A2(o_cddip0_out_ia_wdata_part1[28]), .A3(o_cddip0_out_ia_wdata_part0[28]), .Z(n2910));
Q_MX02 U3433 ( .S(n4549), .A0(i_cddip0_out_ia_rdata_part1[28]), .A1(i_cddip0_out_ia_rdata_part0[28]), .Z(n2911));
Q_AN02 U3434 ( .A0(n4549), .A1(i_cddip0_out_ia_rdata_part2[28]), .Z(n2912));
Q_MX02 U3435 ( .S(n4550), .A0(n2912), .A1(n2911), .Z(n2913));
Q_MX04 U3436 ( .S0(n4551), .S1(n4552), .A0(n2913), .A1(n2910), .A2(n2909), .A3(n2908), .Z(n2914));
Q_MX02 U3437 ( .S(n4553), .A0(n2914), .A1(n2907), .Z(r32_mux_1_data[28]));
Q_MX03 U3438 ( .S0(n4554), .S1(n4555), .A0(o_cceip2_out_ia_config[10]), .A1(o_cceip2_out_ia_wdata_part2[29]), .A2(o_cceip2_out_ia_wdata_part1[29]), .Z(n2915));
Q_MX08 U3439 ( .S0(n4554), .S1(n4555), .S2(n4556), .A0(o_cceip3_out_ia_wdata_part1[29]), .A1(o_cceip3_out_ia_wdata_part0[29]), .A2(i_cceip3_out_ia_status[14]), .A3(i_cceip3_out_ia_capability[17]), .A4(i_cceip2_out_im_status[9]), .A5(i_cceip2_out_ia_rdata_part2[29]), .A6(i_cceip2_out_ia_rdata_part1[29]), .A7(i_cceip2_out_ia_rdata_part0[29]), .Z(n2916));
Q_MX02 U3440 ( .S(n4557), .A0(n2916), .A1(n2915), .Z(n2917));
Q_MX04 U3441 ( .S0(n4554), .S1(n4555), .A0(i_cceip3_out_ia_rdata_part1[29]), .A1(i_cceip3_out_ia_rdata_part0[29]), .A2(o_cceip3_out_ia_config[10]), .A3(o_cceip3_out_ia_wdata_part2[29]), .Z(n2918));
Q_MX04 U3442 ( .S0(n4554), .S1(n4555), .A0(i_cddip0_out_ia_status[14]), .A1(i_cddip0_out_ia_capability[17]), .A2(i_cceip3_out_im_status[9]), .A3(i_cceip3_out_ia_rdata_part2[29]), .Z(n2919));
Q_MX04 U3443 ( .S0(n4554), .S1(n4555), .A0(o_cddip0_out_ia_config[10]), .A1(o_cddip0_out_ia_wdata_part2[29]), .A2(o_cddip0_out_ia_wdata_part1[29]), .A3(o_cddip0_out_ia_wdata_part0[29]), .Z(n2920));
Q_MX02 U3444 ( .S(n4554), .A0(i_cddip0_out_ia_rdata_part1[29]), .A1(i_cddip0_out_ia_rdata_part0[29]), .Z(n2921));
Q_AN02 U3445 ( .A0(n4554), .A1(i_cddip0_out_ia_rdata_part2[29]), .Z(n2922));
Q_MX02 U3446 ( .S(n4555), .A0(n2922), .A1(n2921), .Z(n2923));
Q_MX04 U3447 ( .S0(n4556), .S1(n4557), .A0(n2923), .A1(n2920), .A2(n2919), .A3(n2918), .Z(n2924));
Q_MX02 U3448 ( .S(n4558), .A0(n2924), .A1(n2917), .Z(r32_mux_1_data[29]));
Q_MX03 U3449 ( .S0(n4559), .S1(n4560), .A0(o_cceip2_out_ia_config[11]), .A1(o_cceip2_out_ia_wdata_part2[30]), .A2(o_cceip2_out_ia_wdata_part1[30]), .Z(n2925));
Q_MX04 U3450 ( .S0(n4559), .S1(n4560), .A0(o_cceip2_out_im_config[10]), .A1(i_cceip2_out_ia_rdata_part2[30]), .A2(i_cceip2_out_ia_rdata_part1[30]), .A3(i_cceip2_out_ia_rdata_part0[30]), .Z(n2926));
Q_MX02 U3451 ( .S(n4561), .A0(n2926), .A1(n2925), .Z(n2927));
Q_MX08 U3452 ( .S0(n4559), .S1(n4560), .S2(n4561), .A0(o_cceip3_out_ia_config[11]), .A1(o_cceip3_out_ia_wdata_part2[30]), .A2(o_cceip3_out_ia_wdata_part1[30]), .A3(o_cceip3_out_ia_wdata_part0[30]), .A4(i_cceip3_out_ia_status[15]), .A5(i_cceip3_out_ia_capability[18]), .A6(i_cceip2_out_im_read_done[0]), .A7(i_cceip2_out_im_status[10]), .Z(n2928));
Q_MX02 U3453 ( .S(n4562), .A0(n2928), .A1(n2927), .Z(n2929));
Q_MX04 U3454 ( .S0(n4559), .S1(n4560), .A0(o_cceip3_out_im_config[10]), .A1(i_cceip3_out_ia_rdata_part2[30]), .A2(i_cceip3_out_ia_rdata_part1[30]), .A3(i_cceip3_out_ia_rdata_part0[30]), .Z(n2930));
Q_MX04 U3455 ( .S0(n4559), .S1(n4560), .A0(i_cddip0_out_ia_status[15]), .A1(i_cddip0_out_ia_capability[18]), .A2(i_cceip3_out_im_read_done[0]), .A3(i_cceip3_out_im_status[10]), .Z(n2931));
Q_MX04 U3456 ( .S0(n4559), .S1(n4560), .A0(o_cddip0_out_ia_config[11]), .A1(o_cddip0_out_ia_wdata_part2[30]), .A2(o_cddip0_out_ia_wdata_part1[30]), .A3(o_cddip0_out_ia_wdata_part0[30]), .Z(n2932));
Q_MX02 U3457 ( .S(n4559), .A0(i_cddip0_out_ia_rdata_part1[30]), .A1(i_cddip0_out_ia_rdata_part0[30]), .Z(n2933));
Q_AN02 U3458 ( .A0(n4559), .A1(i_cddip0_out_ia_rdata_part2[30]), .Z(n2934));
Q_MX02 U3459 ( .S(n4560), .A0(n2934), .A1(n2933), .Z(n2935));
Q_MX04 U3460 ( .S0(n4561), .S1(n4562), .A0(n2935), .A1(n2932), .A2(n2931), .A3(n2930), .Z(n2936));
Q_MX02 U3461 ( .S(n4563), .A0(n2936), .A1(n2929), .Z(r32_mux_1_data[30]));
Q_MX03 U3462 ( .S0(n4559), .S1(n4560), .A0(o_cceip2_out_ia_config[12]), .A1(o_cceip2_out_ia_wdata_part2[31]), .A2(o_cceip2_out_ia_wdata_part1[31]), .Z(n2937));
Q_MX04 U3463 ( .S0(n4559), .S1(n4560), .A0(o_cceip2_out_im_config[11]), .A1(i_cceip2_out_ia_rdata_part2[31]), .A2(i_cceip2_out_ia_rdata_part1[31]), .A3(i_cceip2_out_ia_rdata_part0[31]), .Z(n2938));
Q_MX02 U3464 ( .S(n4561), .A0(n2938), .A1(n2937), .Z(n2939));
Q_MX08 U3465 ( .S0(n4559), .S1(n4560), .S2(n4561), .A0(o_cceip3_out_ia_config[12]), .A1(o_cceip3_out_ia_wdata_part2[31]), .A2(o_cceip3_out_ia_wdata_part1[31]), .A3(o_cceip3_out_ia_wdata_part0[31]), .A4(i_cceip3_out_ia_status[16]), .A5(i_cceip3_out_ia_capability[19]), .A6(i_cceip2_out_im_read_done[1]), .A7(i_cceip2_out_im_status[11]), .Z(n2940));
Q_MX02 U3466 ( .S(n4562), .A0(n2940), .A1(n2939), .Z(n2941));
Q_MX04 U3467 ( .S0(n4559), .S1(n4560), .A0(o_cceip3_out_im_config[11]), .A1(i_cceip3_out_ia_rdata_part2[31]), .A2(i_cceip3_out_ia_rdata_part1[31]), .A3(i_cceip3_out_ia_rdata_part0[31]), .Z(n2942));
Q_MX04 U3468 ( .S0(n4559), .S1(n4560), .A0(i_cddip0_out_ia_status[16]), .A1(i_cddip0_out_ia_capability[19]), .A2(i_cceip3_out_im_read_done[1]), .A3(i_cceip3_out_im_status[11]), .Z(n2943));
Q_MX04 U3469 ( .S0(n4559), .S1(n4560), .A0(o_cddip0_out_ia_config[12]), .A1(o_cddip0_out_ia_wdata_part2[31]), .A2(o_cddip0_out_ia_wdata_part1[31]), .A3(o_cddip0_out_ia_wdata_part0[31]), .Z(n2944));
Q_MX02 U3470 ( .S(n4559), .A0(i_cddip0_out_ia_rdata_part1[31]), .A1(i_cddip0_out_ia_rdata_part0[31]), .Z(n2945));
Q_AN02 U3471 ( .A0(n4559), .A1(i_cddip0_out_ia_rdata_part2[31]), .Z(n2946));
Q_MX02 U3472 ( .S(n4560), .A0(n2946), .A1(n2945), .Z(n2947));
Q_MX04 U3473 ( .S0(n4561), .S1(n4562), .A0(n2947), .A1(n2944), .A2(n2943), .A3(n2942), .Z(n2948));
Q_MX02 U3474 ( .S(n4563), .A0(n2948), .A1(n2941), .Z(r32_mux_1_data[31]));
Q_MX04 U3475 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[0]), .A1(i_cceip0_out_ia_capability[0]), .A2(i_spare_config[0]), .A3(i_revision_config[0]), .Z(n2949));
Q_MX02 U3476 ( .S(n4566), .A0(n2949), .A1(i_blkid_revid_config[0]), .Z(n2950));
Q_MX08 U3477 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[0]), .A1(i_cceip0_out_ia_rdata_part2[0]), .A2(i_cceip0_out_ia_rdata_part1[0]), .A3(i_cceip0_out_ia_rdata_part0[0]), .A4(o_cceip0_out_ia_config[0]), .A5(o_cceip0_out_ia_wdata_part2[0]), .A6(o_cceip0_out_ia_wdata_part1[0]), .A7(o_cceip0_out_ia_wdata_part0[0]), .Z(n2951));
Q_MX02 U3478 ( .S(n4567), .A0(n2951), .A1(n2950), .Z(n2952));
Q_MX04 U3479 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[0]), .A1(i_cceip1_out_ia_status[0]), .A2(i_cceip1_out_ia_capability[0]), .A3(i_cceip0_out_im_status[0]), .Z(n2953));
Q_MX04 U3480 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[0]), .A1(o_cceip1_out_ia_config[0]), .A2(o_cceip1_out_ia_wdata_part2[0]), .A3(o_cceip1_out_ia_wdata_part1[0]), .Z(n2954));
Q_MX04 U3481 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[0]), .A1(o_cceip1_out_im_config[0]), .A2(i_cceip1_out_ia_rdata_part2[0]), .A3(i_cceip1_out_ia_rdata_part1[0]), .Z(n2955));
Q_MX02 U3482 ( .S(n4564), .A0(i_cceip2_out_ia_status[0]), .A1(i_cceip2_out_ia_capability[0]), .Z(n2956));
Q_AN02 U3483 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[0]), .Z(n2957));
Q_MX02 U3484 ( .S(n4565), .A0(n2957), .A1(n2956), .Z(n2958));
Q_MX04 U3485 ( .S0(n4566), .S1(n4567), .A0(n2958), .A1(n2955), .A2(n2954), .A3(n2953), .Z(n2959));
Q_MX02 U3486 ( .S(n4568), .A0(n2959), .A1(n2952), .Z(r32_mux_0_data[0]));
Q_MX04 U3487 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[1]), .A1(i_cceip0_out_ia_capability[1]), .A2(i_spare_config[1]), .A3(i_revision_config[1]), .Z(n2960));
Q_MX02 U3488 ( .S(n4566), .A0(n2960), .A1(i_blkid_revid_config[1]), .Z(n2961));
Q_MX08 U3489 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[1]), .A1(i_cceip0_out_ia_rdata_part2[1]), .A2(i_cceip0_out_ia_rdata_part1[1]), .A3(i_cceip0_out_ia_rdata_part0[1]), .A4(o_cceip0_out_ia_config[1]), .A5(o_cceip0_out_ia_wdata_part2[1]), .A6(o_cceip0_out_ia_wdata_part1[1]), .A7(o_cceip0_out_ia_wdata_part0[1]), .Z(n2962));
Q_MX02 U3490 ( .S(n4567), .A0(n2962), .A1(n2961), .Z(n2963));
Q_MX04 U3491 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[1]), .A1(i_cceip1_out_ia_status[1]), .A2(i_cceip1_out_ia_capability[1]), .A3(i_cceip0_out_im_status[1]), .Z(n2964));
Q_MX04 U3492 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[1]), .A1(o_cceip1_out_ia_config[1]), .A2(o_cceip1_out_ia_wdata_part2[1]), .A3(o_cceip1_out_ia_wdata_part1[1]), .Z(n2965));
Q_MX04 U3493 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[1]), .A1(o_cceip1_out_im_config[1]), .A2(i_cceip1_out_ia_rdata_part2[1]), .A3(i_cceip1_out_ia_rdata_part1[1]), .Z(n2966));
Q_MX02 U3494 ( .S(n4564), .A0(i_cceip2_out_ia_status[1]), .A1(i_cceip2_out_ia_capability[1]), .Z(n2967));
Q_AN02 U3495 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[1]), .Z(n2968));
Q_MX02 U3496 ( .S(n4565), .A0(n2968), .A1(n2967), .Z(n2969));
Q_MX04 U3497 ( .S0(n4566), .S1(n4567), .A0(n2969), .A1(n2966), .A2(n2965), .A3(n2964), .Z(n2970));
Q_MX02 U3498 ( .S(n4568), .A0(n2970), .A1(n2963), .Z(r32_mux_0_data[1]));
Q_MX04 U3499 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[2]), .A1(i_cceip0_out_ia_capability[2]), .A2(i_spare_config[2]), .A3(i_revision_config[2]), .Z(n2971));
Q_MX02 U3500 ( .S(n4566), .A0(n2971), .A1(i_blkid_revid_config[2]), .Z(n2972));
Q_MX08 U3501 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[2]), .A1(i_cceip0_out_ia_rdata_part2[2]), .A2(i_cceip0_out_ia_rdata_part1[2]), .A3(i_cceip0_out_ia_rdata_part0[2]), .A4(o_cceip0_out_ia_config[2]), .A5(o_cceip0_out_ia_wdata_part2[2]), .A6(o_cceip0_out_ia_wdata_part1[2]), .A7(o_cceip0_out_ia_wdata_part0[2]), .Z(n2973));
Q_MX02 U3502 ( .S(n4567), .A0(n2973), .A1(n2972), .Z(n2974));
Q_MX04 U3503 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[2]), .A1(i_cceip1_out_ia_status[2]), .A2(i_cceip1_out_ia_capability[2]), .A3(i_cceip0_out_im_status[2]), .Z(n2975));
Q_MX04 U3504 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[2]), .A1(o_cceip1_out_ia_config[2]), .A2(o_cceip1_out_ia_wdata_part2[2]), .A3(o_cceip1_out_ia_wdata_part1[2]), .Z(n2976));
Q_MX04 U3505 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[2]), .A1(o_cceip1_out_im_config[2]), .A2(i_cceip1_out_ia_rdata_part2[2]), .A3(i_cceip1_out_ia_rdata_part1[2]), .Z(n2977));
Q_MX02 U3506 ( .S(n4564), .A0(i_cceip2_out_ia_status[2]), .A1(i_cceip2_out_ia_capability[2]), .Z(n2978));
Q_AN02 U3507 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[2]), .Z(n2979));
Q_MX02 U3508 ( .S(n4565), .A0(n2979), .A1(n2978), .Z(n2980));
Q_MX04 U3509 ( .S0(n4566), .S1(n4567), .A0(n2980), .A1(n2977), .A2(n2976), .A3(n2975), .Z(n2981));
Q_MX02 U3510 ( .S(n4568), .A0(n2981), .A1(n2974), .Z(r32_mux_0_data[2]));
Q_MX04 U3511 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[3]), .A1(i_cceip0_out_ia_capability[3]), .A2(i_spare_config[3]), .A3(i_revision_config[3]), .Z(n2982));
Q_MX02 U3512 ( .S(n4566), .A0(n2982), .A1(i_blkid_revid_config[3]), .Z(n2983));
Q_MX08 U3513 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[3]), .A1(i_cceip0_out_ia_rdata_part2[3]), .A2(i_cceip0_out_ia_rdata_part1[3]), .A3(i_cceip0_out_ia_rdata_part0[3]), .A4(o_cceip0_out_ia_config[3]), .A5(o_cceip0_out_ia_wdata_part2[3]), .A6(o_cceip0_out_ia_wdata_part1[3]), .A7(o_cceip0_out_ia_wdata_part0[3]), .Z(n2984));
Q_MX02 U3514 ( .S(n4567), .A0(n2984), .A1(n2983), .Z(n2985));
Q_MX04 U3515 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[3]), .A1(i_cceip1_out_ia_status[3]), .A2(i_cceip1_out_ia_capability[3]), .A3(i_cceip0_out_im_status[3]), .Z(n2986));
Q_MX04 U3516 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[3]), .A1(o_cceip1_out_ia_config[3]), .A2(o_cceip1_out_ia_wdata_part2[3]), .A3(o_cceip1_out_ia_wdata_part1[3]), .Z(n2987));
Q_MX04 U3517 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[3]), .A1(o_cceip1_out_im_config[3]), .A2(i_cceip1_out_ia_rdata_part2[3]), .A3(i_cceip1_out_ia_rdata_part1[3]), .Z(n2988));
Q_MX02 U3518 ( .S(n4564), .A0(i_cceip2_out_ia_status[3]), .A1(i_cceip2_out_ia_capability[3]), .Z(n2989));
Q_AN02 U3519 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[3]), .Z(n2990));
Q_MX02 U3520 ( .S(n4565), .A0(n2990), .A1(n2989), .Z(n2991));
Q_MX04 U3521 ( .S0(n4566), .S1(n4567), .A0(n2991), .A1(n2988), .A2(n2987), .A3(n2986), .Z(n2992));
Q_MX02 U3522 ( .S(n4568), .A0(n2992), .A1(n2985), .Z(r32_mux_0_data[3]));
Q_MX04 U3523 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[4]), .A1(i_cceip0_out_ia_capability[4]), .A2(i_spare_config[4]), .A3(i_revision_config[4]), .Z(n2993));
Q_MX02 U3524 ( .S(n4566), .A0(n2993), .A1(i_blkid_revid_config[4]), .Z(n2994));
Q_MX08 U3525 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[4]), .A1(i_cceip0_out_ia_rdata_part2[4]), .A2(i_cceip0_out_ia_rdata_part1[4]), .A3(i_cceip0_out_ia_rdata_part0[4]), .A4(o_cceip0_out_ia_config[4]), .A5(o_cceip0_out_ia_wdata_part2[4]), .A6(o_cceip0_out_ia_wdata_part1[4]), .A7(o_cceip0_out_ia_wdata_part0[4]), .Z(n2995));
Q_MX02 U3526 ( .S(n4567), .A0(n2995), .A1(n2994), .Z(n2996));
Q_MX04 U3527 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[4]), .A1(i_cceip1_out_ia_status[4]), .A2(i_cceip1_out_ia_capability[4]), .A3(i_cceip0_out_im_status[4]), .Z(n2997));
Q_MX04 U3528 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[4]), .A1(o_cceip1_out_ia_config[4]), .A2(o_cceip1_out_ia_wdata_part2[4]), .A3(o_cceip1_out_ia_wdata_part1[4]), .Z(n2998));
Q_MX04 U3529 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[4]), .A1(o_cceip1_out_im_config[4]), .A2(i_cceip1_out_ia_rdata_part2[4]), .A3(i_cceip1_out_ia_rdata_part1[4]), .Z(n2999));
Q_MX02 U3530 ( .S(n4564), .A0(i_cceip2_out_ia_status[4]), .A1(i_cceip2_out_ia_capability[4]), .Z(n3000));
Q_AN02 U3531 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[4]), .Z(n3001));
Q_MX02 U3532 ( .S(n4565), .A0(n3001), .A1(n3000), .Z(n3002));
Q_MX04 U3533 ( .S0(n4566), .S1(n4567), .A0(n3002), .A1(n2999), .A2(n2998), .A3(n2997), .Z(n3003));
Q_MX02 U3534 ( .S(n4568), .A0(n3003), .A1(n2996), .Z(r32_mux_0_data[4]));
Q_MX04 U3535 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[5]), .A1(i_cceip0_out_ia_capability[5]), .A2(i_spare_config[5]), .A3(i_revision_config[5]), .Z(n3004));
Q_MX02 U3536 ( .S(n4566), .A0(n3004), .A1(i_blkid_revid_config[5]), .Z(n3005));
Q_MX08 U3537 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[5]), .A1(i_cceip0_out_ia_rdata_part2[5]), .A2(i_cceip0_out_ia_rdata_part1[5]), .A3(i_cceip0_out_ia_rdata_part0[5]), .A4(o_cceip0_out_ia_config[5]), .A5(o_cceip0_out_ia_wdata_part2[5]), .A6(o_cceip0_out_ia_wdata_part1[5]), .A7(o_cceip0_out_ia_wdata_part0[5]), .Z(n3006));
Q_MX02 U3538 ( .S(n4567), .A0(n3006), .A1(n3005), .Z(n3007));
Q_MX04 U3539 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[5]), .A1(i_cceip1_out_ia_status[5]), .A2(i_cceip1_out_ia_capability[5]), .A3(i_cceip0_out_im_status[5]), .Z(n3008));
Q_MX04 U3540 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[5]), .A1(o_cceip1_out_ia_config[5]), .A2(o_cceip1_out_ia_wdata_part2[5]), .A3(o_cceip1_out_ia_wdata_part1[5]), .Z(n3009));
Q_MX04 U3541 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[5]), .A1(o_cceip1_out_im_config[5]), .A2(i_cceip1_out_ia_rdata_part2[5]), .A3(i_cceip1_out_ia_rdata_part1[5]), .Z(n3010));
Q_MX02 U3542 ( .S(n4564), .A0(i_cceip2_out_ia_status[5]), .A1(i_cceip2_out_ia_capability[5]), .Z(n3011));
Q_AN02 U3543 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[5]), .Z(n3012));
Q_MX02 U3544 ( .S(n4565), .A0(n3012), .A1(n3011), .Z(n3013));
Q_MX04 U3545 ( .S0(n4566), .S1(n4567), .A0(n3013), .A1(n3010), .A2(n3009), .A3(n3008), .Z(n3014));
Q_MX02 U3546 ( .S(n4568), .A0(n3014), .A1(n3007), .Z(r32_mux_0_data[5]));
Q_MX04 U3547 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[6]), .A1(i_cceip0_out_ia_capability[6]), .A2(i_spare_config[6]), .A3(i_revision_config[6]), .Z(n3015));
Q_MX02 U3548 ( .S(n4566), .A0(n3015), .A1(i_blkid_revid_config[6]), .Z(n3016));
Q_MX08 U3549 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[6]), .A1(i_cceip0_out_ia_rdata_part2[6]), .A2(i_cceip0_out_ia_rdata_part1[6]), .A3(i_cceip0_out_ia_rdata_part0[6]), .A4(o_cceip0_out_ia_config[6]), .A5(o_cceip0_out_ia_wdata_part2[6]), .A6(o_cceip0_out_ia_wdata_part1[6]), .A7(o_cceip0_out_ia_wdata_part0[6]), .Z(n3017));
Q_MX02 U3550 ( .S(n4567), .A0(n3017), .A1(n3016), .Z(n3018));
Q_MX04 U3551 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[6]), .A1(i_cceip1_out_ia_status[6]), .A2(i_cceip1_out_ia_capability[6]), .A3(i_cceip0_out_im_status[6]), .Z(n3019));
Q_MX04 U3552 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[6]), .A1(o_cceip1_out_ia_config[6]), .A2(o_cceip1_out_ia_wdata_part2[6]), .A3(o_cceip1_out_ia_wdata_part1[6]), .Z(n3020));
Q_MX04 U3553 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[6]), .A1(o_cceip1_out_im_config[6]), .A2(i_cceip1_out_ia_rdata_part2[6]), .A3(i_cceip1_out_ia_rdata_part1[6]), .Z(n3021));
Q_MX02 U3554 ( .S(n4564), .A0(i_cceip2_out_ia_status[6]), .A1(i_cceip2_out_ia_capability[6]), .Z(n3022));
Q_AN02 U3555 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[6]), .Z(n3023));
Q_MX02 U3556 ( .S(n4565), .A0(n3023), .A1(n3022), .Z(n3024));
Q_MX04 U3557 ( .S0(n4566), .S1(n4567), .A0(n3024), .A1(n3021), .A2(n3020), .A3(n3019), .Z(n3025));
Q_MX02 U3558 ( .S(n4568), .A0(n3025), .A1(n3018), .Z(r32_mux_0_data[6]));
Q_MX04 U3559 ( .S0(n4564), .S1(n4565), .A0(i_cceip0_out_ia_status[7]), .A1(i_cceip0_out_ia_capability[7]), .A2(i_spare_config[7]), .A3(i_revision_config[7]), .Z(n3026));
Q_MX02 U3560 ( .S(n4566), .A0(n3026), .A1(i_blkid_revid_config[7]), .Z(n3027));
Q_MX08 U3561 ( .S0(n4564), .S1(n4565), .S2(n4566), .A0(o_cceip0_out_im_config[7]), .A1(i_cceip0_out_ia_rdata_part2[7]), .A2(i_cceip0_out_ia_rdata_part1[7]), .A3(i_cceip0_out_ia_rdata_part0[7]), .A4(o_cceip0_out_ia_config[7]), .A5(o_cceip0_out_ia_wdata_part2[7]), .A6(o_cceip0_out_ia_wdata_part1[7]), .A7(o_cceip0_out_ia_wdata_part0[7]), .Z(n3028));
Q_MX02 U3562 ( .S(n4567), .A0(n3028), .A1(n3027), .Z(n3029));
Q_MX04 U3563 ( .S0(n4564), .S1(n4565), .A0(o_cceip1_out_ia_wdata_part0[7]), .A1(i_cceip1_out_ia_status[7]), .A2(i_cceip1_out_ia_capability[7]), .A3(i_cceip0_out_im_status[7]), .Z(n3030));
Q_MX04 U3564 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_ia_rdata_part0[7]), .A1(o_cceip1_out_ia_config[7]), .A2(o_cceip1_out_ia_wdata_part2[7]), .A3(o_cceip1_out_ia_wdata_part1[7]), .Z(n3031));
Q_MX04 U3565 ( .S0(n4564), .S1(n4565), .A0(i_cceip1_out_im_status[7]), .A1(o_cceip1_out_im_config[7]), .A2(i_cceip1_out_ia_rdata_part2[7]), .A3(i_cceip1_out_ia_rdata_part1[7]), .Z(n3032));
Q_MX02 U3566 ( .S(n4564), .A0(i_cceip2_out_ia_status[7]), .A1(i_cceip2_out_ia_capability[7]), .Z(n3033));
Q_AN02 U3567 ( .A0(n4564), .A1(o_cceip2_out_ia_wdata_part0[7]), .Z(n3034));
Q_MX02 U3568 ( .S(n4565), .A0(n3034), .A1(n3033), .Z(n3035));
Q_MX04 U3569 ( .S0(n4566), .S1(n4567), .A0(n3035), .A1(n3032), .A2(n3031), .A3(n3030), .Z(n3036));
Q_MX02 U3570 ( .S(n4568), .A0(n3036), .A1(n3029), .Z(r32_mux_0_data[7]));
Q_MX04 U3571 ( .S0(n4569), .S1(n4570), .A0(i_cceip0_out_ia_status[8]), .A1(i_cceip0_out_ia_capability[8]), .A2(i_spare_config[8]), .A3(i_blkid_revid_config[8]), .Z(n3037));
Q_MX08 U3572 ( .S0(n4569), .S1(n4570), .S2(n4571), .A0(o_cceip0_out_im_config[8]), .A1(i_cceip0_out_ia_rdata_part2[8]), .A2(i_cceip0_out_ia_rdata_part1[8]), .A3(i_cceip0_out_ia_rdata_part0[8]), .A4(o_cceip0_out_ia_config[8]), .A5(o_cceip0_out_ia_wdata_part2[8]), .A6(o_cceip0_out_ia_wdata_part1[8]), .A7(o_cceip0_out_ia_wdata_part0[8]), .Z(n3038));
Q_MX02 U3573 ( .S(n4572), .A0(n3038), .A1(n3037), .Z(n3039));
Q_MX04 U3574 ( .S0(n4569), .S1(n4570), .A0(o_cceip1_out_ia_wdata_part0[8]), .A1(i_cceip1_out_ia_status[8]), .A2(i_cceip1_out_ia_capability[8]), .A3(i_cceip0_out_im_status[8]), .Z(n3040));
Q_MX04 U3575 ( .S0(n4569), .S1(n4570), .A0(i_cceip1_out_ia_rdata_part0[8]), .A1(o_cceip1_out_ia_config[8]), .A2(o_cceip1_out_ia_wdata_part2[8]), .A3(o_cceip1_out_ia_wdata_part1[8]), .Z(n3041));
Q_MX04 U3576 ( .S0(n4569), .S1(n4570), .A0(i_cceip1_out_im_status[8]), .A1(o_cceip1_out_im_config[8]), .A2(i_cceip1_out_ia_rdata_part2[8]), .A3(i_cceip1_out_ia_rdata_part1[8]), .Z(n3042));
Q_MX02 U3577 ( .S(n4569), .A0(i_cceip2_out_ia_status[8]), .A1(i_cceip2_out_ia_capability[8]), .Z(n3043));
Q_AN02 U3578 ( .A0(n4569), .A1(o_cceip2_out_ia_wdata_part0[8]), .Z(n3044));
Q_MX02 U3579 ( .S(n4570), .A0(n3044), .A1(n3043), .Z(n3045));
Q_MX04 U3580 ( .S0(n4571), .S1(n4572), .A0(n3045), .A1(n3042), .A2(n3041), .A3(n3040), .Z(n3046));
Q_MX02 U3581 ( .S(n4573), .A0(n3046), .A1(n3039), .Z(r32_mux_0_data[8]));
Q_MX04 U3582 ( .S0(n4574), .S1(n4575), .A0(o_cceip0_out_ia_wdata_part1[9]), .A1(o_cceip0_out_ia_wdata_part0[9]), .A2(i_cceip0_out_ia_capability[9]), .A3(i_spare_config[9]), .Z(n3047));
Q_MX02 U3583 ( .S(n4576), .A0(n3047), .A1(i_blkid_revid_config[9]), .Z(n3048));
Q_MX04 U3584 ( .S0(n4574), .S1(n4575), .A0(i_cceip0_out_ia_rdata_part2[9]), .A1(i_cceip0_out_ia_rdata_part1[9]), .A2(i_cceip0_out_ia_rdata_part0[9]), .A3(o_cceip0_out_ia_wdata_part2[9]), .Z(n3049));
Q_MX04 U3585 ( .S0(n4574), .S1(n4575), .A0(o_cceip1_out_ia_wdata_part1[9]), .A1(o_cceip1_out_ia_wdata_part0[9]), .A2(i_cceip1_out_ia_capability[9]), .A3(o_cceip0_out_im_config[9]), .Z(n3050));
Q_MX04 U3586 ( .S0(n4574), .S1(n4575), .A0(i_cceip1_out_ia_rdata_part2[9]), .A1(i_cceip1_out_ia_rdata_part1[9]), .A2(i_cceip1_out_ia_rdata_part0[9]), .A3(o_cceip1_out_ia_wdata_part2[9]), .Z(n3051));
Q_MX02 U3587 ( .S(n4574), .A0(i_cceip2_out_ia_capability[9]), .A1(o_cceip1_out_im_config[9]), .Z(n3052));
Q_AN02 U3588 ( .A0(n4574), .A1(o_cceip2_out_ia_wdata_part0[9]), .Z(n3053));
Q_MX02 U3589 ( .S(n4575), .A0(n3053), .A1(n3052), .Z(n3054));
Q_MX04 U3590 ( .S0(n4576), .S1(n4577), .A0(n3054), .A1(n3051), .A2(n3050), .A3(n3049), .Z(n3055));
Q_MX02 U3591 ( .S(n4578), .A0(n3055), .A1(n3048), .Z(r32_mux_0_data[9]));
Q_MX03 U3592 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_capability[10]), .A1(i_spare_config[10]), .A2(i_blkid_revid_config[10]), .Z(n3056));
Q_MX04 U3593 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_rdata_part0[10]), .A1(o_cceip0_out_ia_wdata_part2[10]), .A2(o_cceip0_out_ia_wdata_part1[10]), .A3(o_cceip0_out_ia_wdata_part0[10]), .Z(n3057));
Q_MX04 U3594 ( .S0(n4579), .S1(n4580), .A0(o_cceip1_out_ia_wdata_part0[10]), .A1(i_cceip1_out_ia_capability[10]), .A2(i_cceip0_out_ia_rdata_part2[10]), .A3(i_cceip0_out_ia_rdata_part1[10]), .Z(n3058));
Q_MX04 U3595 ( .S0(n4579), .S1(n4580), .A0(i_cceip1_out_ia_rdata_part1[10]), .A1(i_cceip1_out_ia_rdata_part0[10]), .A2(o_cceip1_out_ia_wdata_part2[10]), .A3(o_cceip1_out_ia_wdata_part1[10]), .Z(n3059));
Q_MX02 U3596 ( .S(n4579), .A0(i_cceip2_out_ia_capability[10]), .A1(i_cceip1_out_ia_rdata_part2[10]), .Z(n3060));
Q_AN02 U3597 ( .A0(n4579), .A1(o_cceip2_out_ia_wdata_part0[10]), .Z(n3061));
Q_MX02 U3598 ( .S(n4580), .A0(n3061), .A1(n3060), .Z(n3062));
Q_MX04 U3599 ( .S0(n4581), .S1(n4582), .A0(n3062), .A1(n3059), .A2(n3058), .A3(n3057), .Z(n3063));
Q_MX02 U3600 ( .S(n4583), .A0(n3063), .A1(n3056), .Z(r32_mux_0_data[10]));
Q_MX03 U3601 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_capability[11]), .A1(i_spare_config[11]), .A2(i_blkid_revid_config[11]), .Z(n3064));
Q_MX04 U3602 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_rdata_part0[11]), .A1(o_cceip0_out_ia_wdata_part2[11]), .A2(o_cceip0_out_ia_wdata_part1[11]), .A3(o_cceip0_out_ia_wdata_part0[11]), .Z(n3065));
Q_MX04 U3603 ( .S0(n4579), .S1(n4580), .A0(o_cceip1_out_ia_wdata_part0[11]), .A1(i_cceip1_out_ia_capability[11]), .A2(i_cceip0_out_ia_rdata_part2[11]), .A3(i_cceip0_out_ia_rdata_part1[11]), .Z(n3066));
Q_MX04 U3604 ( .S0(n4579), .S1(n4580), .A0(i_cceip1_out_ia_rdata_part1[11]), .A1(i_cceip1_out_ia_rdata_part0[11]), .A2(o_cceip1_out_ia_wdata_part2[11]), .A3(o_cceip1_out_ia_wdata_part1[11]), .Z(n3067));
Q_MX02 U3605 ( .S(n4579), .A0(i_cceip2_out_ia_capability[11]), .A1(i_cceip1_out_ia_rdata_part2[11]), .Z(n3068));
Q_AN02 U3606 ( .A0(n4579), .A1(o_cceip2_out_ia_wdata_part0[11]), .Z(n3069));
Q_MX02 U3607 ( .S(n4580), .A0(n3069), .A1(n3068), .Z(n3070));
Q_MX04 U3608 ( .S0(n4581), .S1(n4582), .A0(n3070), .A1(n3067), .A2(n3066), .A3(n3065), .Z(n3071));
Q_MX02 U3609 ( .S(n4583), .A0(n3071), .A1(n3064), .Z(r32_mux_0_data[11]));
Q_MX03 U3610 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_capability[12]), .A1(i_spare_config[12]), .A2(i_blkid_revid_config[12]), .Z(n3072));
Q_MX04 U3611 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_rdata_part0[12]), .A1(o_cceip0_out_ia_wdata_part2[12]), .A2(o_cceip0_out_ia_wdata_part1[12]), .A3(o_cceip0_out_ia_wdata_part0[12]), .Z(n3073));
Q_MX04 U3612 ( .S0(n4579), .S1(n4580), .A0(o_cceip1_out_ia_wdata_part0[12]), .A1(i_cceip1_out_ia_capability[12]), .A2(i_cceip0_out_ia_rdata_part2[12]), .A3(i_cceip0_out_ia_rdata_part1[12]), .Z(n3074));
Q_MX04 U3613 ( .S0(n4579), .S1(n4580), .A0(i_cceip1_out_ia_rdata_part1[12]), .A1(i_cceip1_out_ia_rdata_part0[12]), .A2(o_cceip1_out_ia_wdata_part2[12]), .A3(o_cceip1_out_ia_wdata_part1[12]), .Z(n3075));
Q_MX02 U3614 ( .S(n4579), .A0(i_cceip2_out_ia_capability[12]), .A1(i_cceip1_out_ia_rdata_part2[12]), .Z(n3076));
Q_AN02 U3615 ( .A0(n4579), .A1(o_cceip2_out_ia_wdata_part0[12]), .Z(n3077));
Q_MX02 U3616 ( .S(n4580), .A0(n3077), .A1(n3076), .Z(n3078));
Q_MX04 U3617 ( .S0(n4581), .S1(n4582), .A0(n3078), .A1(n3075), .A2(n3074), .A3(n3073), .Z(n3079));
Q_MX02 U3618 ( .S(n4583), .A0(n3079), .A1(n3072), .Z(r32_mux_0_data[12]));
Q_MX03 U3619 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_capability[13]), .A1(i_spare_config[13]), .A2(i_blkid_revid_config[13]), .Z(n3080));
Q_MX04 U3620 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_rdata_part0[13]), .A1(o_cceip0_out_ia_wdata_part2[13]), .A2(o_cceip0_out_ia_wdata_part1[13]), .A3(o_cceip0_out_ia_wdata_part0[13]), .Z(n3081));
Q_MX04 U3621 ( .S0(n4579), .S1(n4580), .A0(o_cceip1_out_ia_wdata_part0[13]), .A1(i_cceip1_out_ia_capability[13]), .A2(i_cceip0_out_ia_rdata_part2[13]), .A3(i_cceip0_out_ia_rdata_part1[13]), .Z(n3082));
Q_MX04 U3622 ( .S0(n4579), .S1(n4580), .A0(i_cceip1_out_ia_rdata_part1[13]), .A1(i_cceip1_out_ia_rdata_part0[13]), .A2(o_cceip1_out_ia_wdata_part2[13]), .A3(o_cceip1_out_ia_wdata_part1[13]), .Z(n3083));
Q_MX02 U3623 ( .S(n4579), .A0(i_cceip2_out_ia_capability[13]), .A1(i_cceip1_out_ia_rdata_part2[13]), .Z(n3084));
Q_AN02 U3624 ( .A0(n4579), .A1(o_cceip2_out_ia_wdata_part0[13]), .Z(n3085));
Q_MX02 U3625 ( .S(n4580), .A0(n3085), .A1(n3084), .Z(n3086));
Q_MX04 U3626 ( .S0(n4581), .S1(n4582), .A0(n3086), .A1(n3083), .A2(n3082), .A3(n3081), .Z(n3087));
Q_MX02 U3627 ( .S(n4583), .A0(n3087), .A1(n3080), .Z(r32_mux_0_data[13]));
Q_MX03 U3628 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_capability[14]), .A1(i_spare_config[14]), .A2(i_blkid_revid_config[14]), .Z(n3088));
Q_MX04 U3629 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_rdata_part0[14]), .A1(o_cceip0_out_ia_wdata_part2[14]), .A2(o_cceip0_out_ia_wdata_part1[14]), .A3(o_cceip0_out_ia_wdata_part0[14]), .Z(n3089));
Q_MX04 U3630 ( .S0(n4579), .S1(n4580), .A0(o_cceip1_out_ia_wdata_part0[14]), .A1(i_cceip1_out_ia_capability[14]), .A2(i_cceip0_out_ia_rdata_part2[14]), .A3(i_cceip0_out_ia_rdata_part1[14]), .Z(n3090));
Q_MX04 U3631 ( .S0(n4579), .S1(n4580), .A0(i_cceip1_out_ia_rdata_part1[14]), .A1(i_cceip1_out_ia_rdata_part0[14]), .A2(o_cceip1_out_ia_wdata_part2[14]), .A3(o_cceip1_out_ia_wdata_part1[14]), .Z(n3091));
Q_MX02 U3632 ( .S(n4579), .A0(i_cceip2_out_ia_capability[14]), .A1(i_cceip1_out_ia_rdata_part2[14]), .Z(n3092));
Q_AN02 U3633 ( .A0(n4579), .A1(o_cceip2_out_ia_wdata_part0[14]), .Z(n3093));
Q_MX02 U3634 ( .S(n4580), .A0(n3093), .A1(n3092), .Z(n3094));
Q_MX04 U3635 ( .S0(n4581), .S1(n4582), .A0(n3094), .A1(n3091), .A2(n3090), .A3(n3089), .Z(n3095));
Q_MX02 U3636 ( .S(n4583), .A0(n3095), .A1(n3088), .Z(r32_mux_0_data[14]));
Q_MX03 U3637 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_capability[15]), .A1(i_spare_config[15]), .A2(i_blkid_revid_config[15]), .Z(n3096));
Q_MX04 U3638 ( .S0(n4579), .S1(n4580), .A0(i_cceip0_out_ia_rdata_part0[15]), .A1(o_cceip0_out_ia_wdata_part2[15]), .A2(o_cceip0_out_ia_wdata_part1[15]), .A3(o_cceip0_out_ia_wdata_part0[15]), .Z(n3097));
Q_MX04 U3639 ( .S0(n4579), .S1(n4580), .A0(o_cceip1_out_ia_wdata_part0[15]), .A1(i_cceip1_out_ia_capability[15]), .A2(i_cceip0_out_ia_rdata_part2[15]), .A3(i_cceip0_out_ia_rdata_part1[15]), .Z(n3098));
Q_MX04 U3640 ( .S0(n4579), .S1(n4580), .A0(i_cceip1_out_ia_rdata_part1[15]), .A1(i_cceip1_out_ia_rdata_part0[15]), .A2(o_cceip1_out_ia_wdata_part2[15]), .A3(o_cceip1_out_ia_wdata_part1[15]), .Z(n3099));
Q_MX02 U3641 ( .S(n4579), .A0(i_cceip2_out_ia_capability[15]), .A1(i_cceip1_out_ia_rdata_part2[15]), .Z(n3100));
Q_AN02 U3642 ( .A0(n4579), .A1(o_cceip2_out_ia_wdata_part0[15]), .Z(n3101));
Q_MX02 U3643 ( .S(n4580), .A0(n3101), .A1(n3100), .Z(n3102));
Q_MX04 U3644 ( .S0(n4581), .S1(n4582), .A0(n3102), .A1(n3099), .A2(n3098), .A3(n3097), .Z(n3103));
Q_MX02 U3645 ( .S(n4583), .A0(n3103), .A1(n3096), .Z(r32_mux_0_data[15]));
Q_MX04 U3646 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[16]), .A1(o_cceip0_out_ia_wdata_part0[16]), .A2(i_spare_config[16]), .A3(i_blkid_revid_config[16]), .Z(n3104));
Q_MX04 U3647 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[16]), .A1(i_cceip0_out_ia_rdata_part1[16]), .A2(i_cceip0_out_ia_rdata_part0[16]), .A3(o_cceip0_out_ia_wdata_part2[16]), .Z(n3105));
Q_MX04 U3648 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[16]), .A1(o_cceip1_out_ia_wdata_part2[16]), .A2(o_cceip1_out_ia_wdata_part1[16]), .A3(o_cceip1_out_ia_wdata_part0[16]), .Z(n3106));
Q_MX02 U3649 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[16]), .A1(i_cceip1_out_ia_rdata_part1[16]), .Z(n3107));
Q_AN02 U3650 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[16]), .Z(n3108));
Q_MX02 U3651 ( .S(n4585), .A0(n3108), .A1(n3107), .Z(n3109));
Q_MX04 U3652 ( .S0(n4586), .S1(n4587), .A0(n3109), .A1(n3106), .A2(n3105), .A3(n3104), .Z(r32_mux_0_data[16]));
Q_MX04 U3653 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[17]), .A1(o_cceip0_out_ia_wdata_part0[17]), .A2(i_spare_config[17]), .A3(i_blkid_revid_config[17]), .Z(n3110));
Q_MX04 U3654 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[17]), .A1(i_cceip0_out_ia_rdata_part1[17]), .A2(i_cceip0_out_ia_rdata_part0[17]), .A3(o_cceip0_out_ia_wdata_part2[17]), .Z(n3111));
Q_MX04 U3655 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[17]), .A1(o_cceip1_out_ia_wdata_part2[17]), .A2(o_cceip1_out_ia_wdata_part1[17]), .A3(o_cceip1_out_ia_wdata_part0[17]), .Z(n3112));
Q_MX02 U3656 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[17]), .A1(i_cceip1_out_ia_rdata_part1[17]), .Z(n3113));
Q_AN02 U3657 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[17]), .Z(n3114));
Q_MX02 U3658 ( .S(n4585), .A0(n3114), .A1(n3113), .Z(n3115));
Q_MX04 U3659 ( .S0(n4586), .S1(n4587), .A0(n3115), .A1(n3112), .A2(n3111), .A3(n3110), .Z(r32_mux_0_data[17]));
Q_MX04 U3660 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[18]), .A1(o_cceip0_out_ia_wdata_part0[18]), .A2(i_spare_config[18]), .A3(i_blkid_revid_config[18]), .Z(n3116));
Q_MX04 U3661 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[18]), .A1(i_cceip0_out_ia_rdata_part1[18]), .A2(i_cceip0_out_ia_rdata_part0[18]), .A3(o_cceip0_out_ia_wdata_part2[18]), .Z(n3117));
Q_MX04 U3662 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[18]), .A1(o_cceip1_out_ia_wdata_part2[18]), .A2(o_cceip1_out_ia_wdata_part1[18]), .A3(o_cceip1_out_ia_wdata_part0[18]), .Z(n3118));
Q_MX02 U3663 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[18]), .A1(i_cceip1_out_ia_rdata_part1[18]), .Z(n3119));
Q_AN02 U3664 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[18]), .Z(n3120));
Q_MX02 U3665 ( .S(n4585), .A0(n3120), .A1(n3119), .Z(n3121));
Q_MX04 U3666 ( .S0(n4586), .S1(n4587), .A0(n3121), .A1(n3118), .A2(n3117), .A3(n3116), .Z(r32_mux_0_data[18]));
Q_MX04 U3667 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[19]), .A1(o_cceip0_out_ia_wdata_part0[19]), .A2(i_spare_config[19]), .A3(i_blkid_revid_config[19]), .Z(n3122));
Q_MX04 U3668 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[19]), .A1(i_cceip0_out_ia_rdata_part1[19]), .A2(i_cceip0_out_ia_rdata_part0[19]), .A3(o_cceip0_out_ia_wdata_part2[19]), .Z(n3123));
Q_MX04 U3669 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[19]), .A1(o_cceip1_out_ia_wdata_part2[19]), .A2(o_cceip1_out_ia_wdata_part1[19]), .A3(o_cceip1_out_ia_wdata_part0[19]), .Z(n3124));
Q_MX02 U3670 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[19]), .A1(i_cceip1_out_ia_rdata_part1[19]), .Z(n3125));
Q_AN02 U3671 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[19]), .Z(n3126));
Q_MX02 U3672 ( .S(n4585), .A0(n3126), .A1(n3125), .Z(n3127));
Q_MX04 U3673 ( .S0(n4586), .S1(n4587), .A0(n3127), .A1(n3124), .A2(n3123), .A3(n3122), .Z(r32_mux_0_data[19]));
Q_MX04 U3674 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[20]), .A1(o_cceip0_out_ia_wdata_part0[20]), .A2(i_spare_config[20]), .A3(i_blkid_revid_config[20]), .Z(n3128));
Q_MX04 U3675 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[20]), .A1(i_cceip0_out_ia_rdata_part1[20]), .A2(i_cceip0_out_ia_rdata_part0[20]), .A3(o_cceip0_out_ia_wdata_part2[20]), .Z(n3129));
Q_MX04 U3676 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[20]), .A1(o_cceip1_out_ia_wdata_part2[20]), .A2(o_cceip1_out_ia_wdata_part1[20]), .A3(o_cceip1_out_ia_wdata_part0[20]), .Z(n3130));
Q_MX02 U3677 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[20]), .A1(i_cceip1_out_ia_rdata_part1[20]), .Z(n3131));
Q_AN02 U3678 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[20]), .Z(n3132));
Q_MX02 U3679 ( .S(n4585), .A0(n3132), .A1(n3131), .Z(n3133));
Q_MX04 U3680 ( .S0(n4586), .S1(n4587), .A0(n3133), .A1(n3130), .A2(n3129), .A3(n3128), .Z(r32_mux_0_data[20]));
Q_MX04 U3681 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[21]), .A1(o_cceip0_out_ia_wdata_part0[21]), .A2(i_spare_config[21]), .A3(i_blkid_revid_config[21]), .Z(n3134));
Q_MX04 U3682 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[21]), .A1(i_cceip0_out_ia_rdata_part1[21]), .A2(i_cceip0_out_ia_rdata_part0[21]), .A3(o_cceip0_out_ia_wdata_part2[21]), .Z(n3135));
Q_MX04 U3683 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[21]), .A1(o_cceip1_out_ia_wdata_part2[21]), .A2(o_cceip1_out_ia_wdata_part1[21]), .A3(o_cceip1_out_ia_wdata_part0[21]), .Z(n3136));
Q_MX02 U3684 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[21]), .A1(i_cceip1_out_ia_rdata_part1[21]), .Z(n3137));
Q_AN02 U3685 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[21]), .Z(n3138));
Q_MX02 U3686 ( .S(n4585), .A0(n3138), .A1(n3137), .Z(n3139));
Q_MX04 U3687 ( .S0(n4586), .S1(n4587), .A0(n3139), .A1(n3136), .A2(n3135), .A3(n3134), .Z(r32_mux_0_data[21]));
Q_MX04 U3688 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[22]), .A1(o_cceip0_out_ia_wdata_part0[22]), .A2(i_spare_config[22]), .A3(i_blkid_revid_config[22]), .Z(n3140));
Q_MX04 U3689 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[22]), .A1(i_cceip0_out_ia_rdata_part1[22]), .A2(i_cceip0_out_ia_rdata_part0[22]), .A3(o_cceip0_out_ia_wdata_part2[22]), .Z(n3141));
Q_MX04 U3690 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[22]), .A1(o_cceip1_out_ia_wdata_part2[22]), .A2(o_cceip1_out_ia_wdata_part1[22]), .A3(o_cceip1_out_ia_wdata_part0[22]), .Z(n3142));
Q_MX02 U3691 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[22]), .A1(i_cceip1_out_ia_rdata_part1[22]), .Z(n3143));
Q_AN02 U3692 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[22]), .Z(n3144));
Q_MX02 U3693 ( .S(n4585), .A0(n3144), .A1(n3143), .Z(n3145));
Q_MX04 U3694 ( .S0(n4586), .S1(n4587), .A0(n3145), .A1(n3142), .A2(n3141), .A3(n3140), .Z(r32_mux_0_data[22]));
Q_MX04 U3695 ( .S0(n4584), .S1(n4585), .A0(o_cceip0_out_ia_wdata_part1[23]), .A1(o_cceip0_out_ia_wdata_part0[23]), .A2(i_spare_config[23]), .A3(i_blkid_revid_config[23]), .Z(n3146));
Q_MX04 U3696 ( .S0(n4584), .S1(n4585), .A0(i_cceip0_out_ia_rdata_part2[23]), .A1(i_cceip0_out_ia_rdata_part1[23]), .A2(i_cceip0_out_ia_rdata_part0[23]), .A3(o_cceip0_out_ia_wdata_part2[23]), .Z(n3147));
Q_MX04 U3697 ( .S0(n4584), .S1(n4585), .A0(i_cceip1_out_ia_rdata_part0[23]), .A1(o_cceip1_out_ia_wdata_part2[23]), .A2(o_cceip1_out_ia_wdata_part1[23]), .A3(o_cceip1_out_ia_wdata_part0[23]), .Z(n3148));
Q_MX02 U3698 ( .S(n4584), .A0(i_cceip1_out_ia_rdata_part2[23]), .A1(i_cceip1_out_ia_rdata_part1[23]), .Z(n3149));
Q_AN02 U3699 ( .A0(n4584), .A1(o_cceip2_out_ia_wdata_part0[23]), .Z(n3150));
Q_MX02 U3700 ( .S(n4585), .A0(n3150), .A1(n3149), .Z(n3151));
Q_MX04 U3701 ( .S0(n4586), .S1(n4587), .A0(n3151), .A1(n3148), .A2(n3147), .A3(n3146), .Z(r32_mux_0_data[23]));
Q_MX03 U3702 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_status[9]), .A1(i_spare_config[24]), .A2(i_blkid_revid_config[24]), .Z(n3152));
Q_MX04 U3703 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_rdata_part0[24]), .A1(o_cceip0_out_ia_wdata_part2[24]), .A2(o_cceip0_out_ia_wdata_part1[24]), .A3(o_cceip0_out_ia_wdata_part0[24]), .Z(n3153));
Q_MX04 U3704 ( .S0(n4588), .S1(n4589), .A0(o_cceip1_out_ia_wdata_part0[24]), .A1(i_cceip1_out_ia_status[9]), .A2(i_cceip0_out_ia_rdata_part2[24]), .A3(i_cceip0_out_ia_rdata_part1[24]), .Z(n3154));
Q_MX04 U3705 ( .S0(n4588), .S1(n4589), .A0(i_cceip1_out_ia_rdata_part1[24]), .A1(i_cceip1_out_ia_rdata_part0[24]), .A2(o_cceip1_out_ia_wdata_part2[24]), .A3(o_cceip1_out_ia_wdata_part1[24]), .Z(n3155));
Q_MX02 U3706 ( .S(n4588), .A0(i_cceip2_out_ia_status[9]), .A1(i_cceip1_out_ia_rdata_part2[24]), .Z(n3156));
Q_AN02 U3707 ( .A0(n4588), .A1(o_cceip2_out_ia_wdata_part0[24]), .Z(n3157));
Q_MX02 U3708 ( .S(n4589), .A0(n3157), .A1(n3156), .Z(n3158));
Q_MX04 U3709 ( .S0(n4581), .S1(n4590), .A0(n3158), .A1(n3155), .A2(n3154), .A3(n3153), .Z(n3159));
Q_MX02 U3710 ( .S(n4591), .A0(n3159), .A1(n3152), .Z(r32_mux_0_data[24]));
Q_MX03 U3711 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_status[10]), .A1(i_spare_config[25]), .A2(i_blkid_revid_config[25]), .Z(n3160));
Q_MX04 U3712 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_rdata_part0[25]), .A1(o_cceip0_out_ia_wdata_part2[25]), .A2(o_cceip0_out_ia_wdata_part1[25]), .A3(o_cceip0_out_ia_wdata_part0[25]), .Z(n3161));
Q_MX04 U3713 ( .S0(n4588), .S1(n4589), .A0(o_cceip1_out_ia_wdata_part0[25]), .A1(i_cceip1_out_ia_status[10]), .A2(i_cceip0_out_ia_rdata_part2[25]), .A3(i_cceip0_out_ia_rdata_part1[25]), .Z(n3162));
Q_MX04 U3714 ( .S0(n4588), .S1(n4589), .A0(i_cceip1_out_ia_rdata_part1[25]), .A1(i_cceip1_out_ia_rdata_part0[25]), .A2(o_cceip1_out_ia_wdata_part2[25]), .A3(o_cceip1_out_ia_wdata_part1[25]), .Z(n3163));
Q_MX02 U3715 ( .S(n4588), .A0(i_cceip2_out_ia_status[10]), .A1(i_cceip1_out_ia_rdata_part2[25]), .Z(n3164));
Q_AN02 U3716 ( .A0(n4588), .A1(o_cceip2_out_ia_wdata_part0[25]), .Z(n3165));
Q_MX02 U3717 ( .S(n4589), .A0(n3165), .A1(n3164), .Z(n3166));
Q_MX04 U3718 ( .S0(n4581), .S1(n4590), .A0(n3166), .A1(n3163), .A2(n3162), .A3(n3161), .Z(n3167));
Q_MX02 U3719 ( .S(n4591), .A0(n3167), .A1(n3160), .Z(r32_mux_0_data[25]));
Q_MX03 U3720 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_status[11]), .A1(i_spare_config[26]), .A2(i_blkid_revid_config[26]), .Z(n3168));
Q_MX04 U3721 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_rdata_part0[26]), .A1(o_cceip0_out_ia_wdata_part2[26]), .A2(o_cceip0_out_ia_wdata_part1[26]), .A3(o_cceip0_out_ia_wdata_part0[26]), .Z(n3169));
Q_MX04 U3722 ( .S0(n4588), .S1(n4589), .A0(o_cceip1_out_ia_wdata_part0[26]), .A1(i_cceip1_out_ia_status[11]), .A2(i_cceip0_out_ia_rdata_part2[26]), .A3(i_cceip0_out_ia_rdata_part1[26]), .Z(n3170));
Q_MX04 U3723 ( .S0(n4588), .S1(n4589), .A0(i_cceip1_out_ia_rdata_part1[26]), .A1(i_cceip1_out_ia_rdata_part0[26]), .A2(o_cceip1_out_ia_wdata_part2[26]), .A3(o_cceip1_out_ia_wdata_part1[26]), .Z(n3171));
Q_MX02 U3724 ( .S(n4588), .A0(i_cceip2_out_ia_status[11]), .A1(i_cceip1_out_ia_rdata_part2[26]), .Z(n3172));
Q_AN02 U3725 ( .A0(n4588), .A1(o_cceip2_out_ia_wdata_part0[26]), .Z(n3173));
Q_MX02 U3726 ( .S(n4589), .A0(n3173), .A1(n3172), .Z(n3174));
Q_MX04 U3727 ( .S0(n4581), .S1(n4590), .A0(n3174), .A1(n3171), .A2(n3170), .A3(n3169), .Z(n3175));
Q_MX02 U3728 ( .S(n4591), .A0(n3175), .A1(n3168), .Z(r32_mux_0_data[26]));
Q_MX03 U3729 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_status[12]), .A1(i_spare_config[27]), .A2(i_blkid_revid_config[27]), .Z(n3176));
Q_MX04 U3730 ( .S0(n4588), .S1(n4589), .A0(i_cceip0_out_ia_rdata_part0[27]), .A1(o_cceip0_out_ia_wdata_part2[27]), .A2(o_cceip0_out_ia_wdata_part1[27]), .A3(o_cceip0_out_ia_wdata_part0[27]), .Z(n3177));
Q_MX04 U3731 ( .S0(n4588), .S1(n4589), .A0(o_cceip1_out_ia_wdata_part0[27]), .A1(i_cceip1_out_ia_status[12]), .A2(i_cceip0_out_ia_rdata_part2[27]), .A3(i_cceip0_out_ia_rdata_part1[27]), .Z(n3178));
Q_MX04 U3732 ( .S0(n4588), .S1(n4589), .A0(i_cceip1_out_ia_rdata_part1[27]), .A1(i_cceip1_out_ia_rdata_part0[27]), .A2(o_cceip1_out_ia_wdata_part2[27]), .A3(o_cceip1_out_ia_wdata_part1[27]), .Z(n3179));
Q_MX02 U3733 ( .S(n4588), .A0(i_cceip2_out_ia_status[12]), .A1(i_cceip1_out_ia_rdata_part2[27]), .Z(n3180));
Q_AN02 U3734 ( .A0(n4588), .A1(o_cceip2_out_ia_wdata_part0[27]), .Z(n3181));
Q_MX02 U3735 ( .S(n4589), .A0(n3181), .A1(n3180), .Z(n3182));
Q_MX04 U3736 ( .S0(n4581), .S1(n4590), .A0(n3182), .A1(n3179), .A2(n3178), .A3(n3177), .Z(n3183));
Q_MX02 U3737 ( .S(n4591), .A0(n3183), .A1(n3176), .Z(r32_mux_0_data[27]));
Q_MX08 U3738 ( .S0(n4592), .S1(n4593), .S2(n4594), .A0(o_cceip0_out_ia_config[9]), .A1(o_cceip0_out_ia_wdata_part2[28]), .A2(o_cceip0_out_ia_wdata_part1[28]), .A3(o_cceip0_out_ia_wdata_part0[28]), .A4(i_cceip0_out_ia_status[13]), .A5(i_cceip0_out_ia_capability[16]), .A6(i_spare_config[28]), .A7(i_blkid_revid_config[28]), .Z(n3184));
Q_MX04 U3739 ( .S0(n4592), .S1(n4593), .A0(i_cceip1_out_ia_capability[16]), .A1(i_cceip0_out_ia_rdata_part2[28]), .A2(i_cceip0_out_ia_rdata_part1[28]), .A3(i_cceip0_out_ia_rdata_part0[28]), .Z(n3185));
Q_MX04 U3740 ( .S0(n4592), .S1(n4593), .A0(o_cceip1_out_ia_wdata_part2[28]), .A1(o_cceip1_out_ia_wdata_part1[28]), .A2(o_cceip1_out_ia_wdata_part0[28]), .A3(i_cceip1_out_ia_status[13]), .Z(n3186));
Q_MX04 U3741 ( .S0(n4592), .S1(n4593), .A0(i_cceip1_out_ia_rdata_part2[28]), .A1(i_cceip1_out_ia_rdata_part1[28]), .A2(i_cceip1_out_ia_rdata_part0[28]), .A3(o_cceip1_out_ia_config[9]), .Z(n3187));
Q_MX02 U3742 ( .S(n4592), .A0(i_cceip2_out_ia_status[13]), .A1(i_cceip2_out_ia_capability[16]), .Z(n3188));
Q_AN02 U3743 ( .A0(n4592), .A1(o_cceip2_out_ia_wdata_part0[28]), .Z(n3189));
Q_MX02 U3744 ( .S(n4593), .A0(n3189), .A1(n3188), .Z(n3190));
Q_MX04 U3745 ( .S0(n4594), .S1(n4595), .A0(n3190), .A1(n3187), .A2(n3186), .A3(n3185), .Z(n3191));
Q_MX02 U3746 ( .S(n4596), .A0(n3191), .A1(n3184), .Z(r32_mux_0_data[28]));
Q_MX02 U3747 ( .S(n4597), .A0(i_spare_config[29]), .A1(i_blkid_revid_config[29]), .Z(n3192));
Q_MX08 U3748 ( .S0(n4597), .S1(n4598), .S2(n4599), .A0(i_cceip0_out_ia_rdata_part1[29]), .A1(i_cceip0_out_ia_rdata_part0[29]), .A2(o_cceip0_out_ia_config[10]), .A3(o_cceip0_out_ia_wdata_part2[29]), .A4(o_cceip0_out_ia_wdata_part1[29]), .A5(o_cceip0_out_ia_wdata_part0[29]), .A6(i_cceip0_out_ia_status[14]), .A7(i_cceip0_out_ia_capability[17]), .Z(n3193));
Q_MX02 U3749 ( .S(n4600), .A0(n3193), .A1(n3192), .Z(n3194));
Q_MX04 U3750 ( .S0(n4597), .S1(n4598), .A0(i_cceip1_out_ia_status[14]), .A1(i_cceip1_out_ia_capability[17]), .A2(i_cceip0_out_im_status[9]), .A3(i_cceip0_out_ia_rdata_part2[29]), .Z(n3195));
Q_MX04 U3751 ( .S0(n4597), .S1(n4598), .A0(o_cceip1_out_ia_config[10]), .A1(o_cceip1_out_ia_wdata_part2[29]), .A2(o_cceip1_out_ia_wdata_part1[29]), .A3(o_cceip1_out_ia_wdata_part0[29]), .Z(n3196));
Q_MX04 U3752 ( .S0(n4597), .S1(n4598), .A0(i_cceip1_out_im_status[9]), .A1(i_cceip1_out_ia_rdata_part2[29]), .A2(i_cceip1_out_ia_rdata_part1[29]), .A3(i_cceip1_out_ia_rdata_part0[29]), .Z(n3197));
Q_MX02 U3753 ( .S(n4597), .A0(i_cceip2_out_ia_status[14]), .A1(i_cceip2_out_ia_capability[17]), .Z(n3198));
Q_AN02 U3754 ( .A0(n4597), .A1(o_cceip2_out_ia_wdata_part0[29]), .Z(n3199));
Q_MX02 U3755 ( .S(n4598), .A0(n3199), .A1(n3198), .Z(n3200));
Q_MX04 U3756 ( .S0(n4599), .S1(n4600), .A0(n3200), .A1(n3197), .A2(n3196), .A3(n3195), .Z(n3201));
Q_MX02 U3757 ( .S(n4601), .A0(n3201), .A1(n3194), .Z(r32_mux_0_data[29]));
Q_MX02 U3758 ( .S(n4602), .A0(i_spare_config[30]), .A1(i_blkid_revid_config[30]), .Z(n3202));
Q_MX04 U3759 ( .S0(n4602), .S1(n4603), .A0(o_cceip0_out_ia_wdata_part1[30]), .A1(o_cceip0_out_ia_wdata_part0[30]), .A2(i_cceip0_out_ia_status[15]), .A3(i_cceip0_out_ia_capability[18]), .Z(n3203));
Q_MX02 U3760 ( .S(n4604), .A0(n3203), .A1(n3202), .Z(n3204));
Q_MX08 U3761 ( .S0(n4602), .S1(n4603), .S2(n4604), .A0(i_cceip0_out_im_read_done[0]), .A1(i_cceip0_out_im_status[10]), .A2(o_cceip0_out_im_config[10]), .A3(i_cceip0_out_ia_rdata_part2[30]), .A4(i_cceip0_out_ia_rdata_part1[30]), .A5(i_cceip0_out_ia_rdata_part0[30]), .A6(o_cceip0_out_ia_config[11]), .A7(o_cceip0_out_ia_wdata_part2[30]), .Z(n3205));
Q_MX02 U3762 ( .S(n4605), .A0(n3205), .A1(n3204), .Z(n3206));
Q_MX04 U3763 ( .S0(n4602), .S1(n4603), .A0(o_cceip1_out_ia_wdata_part1[30]), .A1(o_cceip1_out_ia_wdata_part0[30]), .A2(i_cceip1_out_ia_status[15]), .A3(i_cceip1_out_ia_capability[18]), .Z(n3207));
Q_MX04 U3764 ( .S0(n4602), .S1(n4603), .A0(i_cceip1_out_ia_rdata_part1[30]), .A1(i_cceip1_out_ia_rdata_part0[30]), .A2(o_cceip1_out_ia_config[11]), .A3(o_cceip1_out_ia_wdata_part2[30]), .Z(n3208));
Q_MX04 U3765 ( .S0(n4602), .S1(n4603), .A0(i_cceip1_out_im_read_done[0]), .A1(i_cceip1_out_im_status[10]), .A2(o_cceip1_out_im_config[10]), .A3(i_cceip1_out_ia_rdata_part2[30]), .Z(n3209));
Q_MX02 U3766 ( .S(n4602), .A0(i_cceip2_out_ia_status[15]), .A1(i_cceip2_out_ia_capability[18]), .Z(n3210));
Q_AN02 U3767 ( .A0(n4602), .A1(o_cceip2_out_ia_wdata_part0[30]), .Z(n3211));
Q_MX02 U3768 ( .S(n4603), .A0(n3211), .A1(n3210), .Z(n3212));
Q_MX04 U3769 ( .S0(n4604), .S1(n4605), .A0(n3212), .A1(n3209), .A2(n3208), .A3(n3207), .Z(n3213));
Q_MX02 U3770 ( .S(n4606), .A0(n3213), .A1(n3206), .Z(r32_mux_0_data[30]));
Q_MX02 U3771 ( .S(n4602), .A0(i_spare_config[31]), .A1(i_blkid_revid_config[31]), .Z(n3214));
Q_MX04 U3772 ( .S0(n4602), .S1(n4603), .A0(o_cceip0_out_ia_wdata_part1[31]), .A1(o_cceip0_out_ia_wdata_part0[31]), .A2(i_cceip0_out_ia_status[16]), .A3(i_cceip0_out_ia_capability[19]), .Z(n3215));
Q_MX02 U3773 ( .S(n4604), .A0(n3215), .A1(n3214), .Z(n3216));
Q_MX08 U3774 ( .S0(n4602), .S1(n4603), .S2(n4604), .A0(i_cceip0_out_im_read_done[1]), .A1(i_cceip0_out_im_status[11]), .A2(o_cceip0_out_im_config[11]), .A3(i_cceip0_out_ia_rdata_part2[31]), .A4(i_cceip0_out_ia_rdata_part1[31]), .A5(i_cceip0_out_ia_rdata_part0[31]), .A6(o_cceip0_out_ia_config[12]), .A7(o_cceip0_out_ia_wdata_part2[31]), .Z(n3217));
Q_MX02 U3775 ( .S(n4605), .A0(n3217), .A1(n3216), .Z(n3218));
Q_MX04 U3776 ( .S0(n4602), .S1(n4603), .A0(o_cceip1_out_ia_wdata_part1[31]), .A1(o_cceip1_out_ia_wdata_part0[31]), .A2(i_cceip1_out_ia_status[16]), .A3(i_cceip1_out_ia_capability[19]), .Z(n3219));
Q_MX04 U3777 ( .S0(n4602), .S1(n4603), .A0(i_cceip1_out_ia_rdata_part1[31]), .A1(i_cceip1_out_ia_rdata_part0[31]), .A2(o_cceip1_out_ia_config[12]), .A3(o_cceip1_out_ia_wdata_part2[31]), .Z(n3220));
Q_MX04 U3778 ( .S0(n4602), .S1(n4603), .A0(i_cceip1_out_im_read_done[1]), .A1(i_cceip1_out_im_status[11]), .A2(o_cceip1_out_im_config[11]), .A3(i_cceip1_out_ia_rdata_part2[31]), .Z(n3221));
Q_MX02 U3779 ( .S(n4602), .A0(i_cceip2_out_ia_status[16]), .A1(i_cceip2_out_ia_capability[19]), .Z(n3222));
Q_AN02 U3780 ( .A0(n4602), .A1(o_cceip2_out_ia_wdata_part0[31]), .Z(n3223));
Q_MX02 U3781 ( .S(n4603), .A0(n3223), .A1(n3222), .Z(n3224));
Q_MX04 U3782 ( .S0(n4604), .S1(n4605), .A0(n3224), .A1(n3221), .A2(n3220), .A3(n3219), .Z(n3225));
Q_MX02 U3783 ( .S(n4606), .A0(n3225), .A1(n3218), .Z(r32_mux_0_data[31]));
Q_OA21 U3784 ( .A0(n3227), .A1(n3228), .B0(n3226), .Z(n4313));
Q_AO21 U3785 ( .A0(n3229), .A1(n3230), .B0(n3231), .Z(n3227));
Q_AN02 U3786 ( .A0(n3232), .A1(n3233), .Z(n3228));
Q_OA21 U3787 ( .A0(n3235), .A1(n3236), .B0(n3234), .Z(n4314));
Q_AO21 U3788 ( .A0(n3238), .A1(n3231), .B0(n3237), .Z(n3235));
Q_OA21 U3789 ( .A0(n3239), .A1(n3240), .B0(n3230), .Z(n3237));
Q_OA21 U3790 ( .A0(n3241), .A1(n3242), .B0(n3234), .Z(n4315));
Q_AO21 U3791 ( .A0(n3244), .A1(n3231), .B0(n3243), .Z(n3242));
Q_OA21 U3792 ( .A0(n3245), .A1(n3246), .B0(n3230), .Z(n3241));
Q_OA21 U3793 ( .A0(n3247), .A1(n3248), .B0(n3234), .Z(n4316));
Q_AN02 U3794 ( .A0(n3249), .A1(n3230), .Z(n3247));
Q_OA21 U3795 ( .A0(n3250), .A1(n3248), .B0(n3234), .Z(n4317));
Q_AN02 U3796 ( .A0(n3251), .A1(n3252), .Z(n3250));
Q_OR03 U3797 ( .A0(n3253), .A1(n3236), .A2(n3243), .Z(n3248));
Q_AN02 U3798 ( .A0(n3233), .A1(n3255), .Z(n3254));
Q_AO21 U3799 ( .A0(n3231), .A1(n3256), .B0(n3254), .Z(n3253));
Q_OA21 U3800 ( .A0(n3257), .A1(n3258), .B0(n3234), .Z(n4318));
Q_AN03 U3801 ( .A0(n3232), .A1(ws_read_addr[2]), .A2(n3233), .Z(n3259));
Q_AO21 U3802 ( .A0(n3260), .A1(n3252), .B0(n3259), .Z(n3258));
Q_OR02 U3803 ( .A0(n3261), .A1(n3262), .Z(n3260));
Q_OA21 U3804 ( .A0(n3263), .A1(n3264), .B0(n3230), .Z(n3257));
Q_OA21 U3805 ( .A0(n3265), .A1(n3266), .B0(n3234), .Z(n4319));
Q_AN02 U3806 ( .A0(n3238), .A1(n3268), .Z(n3269));
Q_OR03 U3807 ( .A0(n3269), .A1(n3243), .A2(n3267), .Z(n3266));
Q_OA21 U3808 ( .A0(n3270), .A1(n3271), .B0(n3230), .Z(n3265));
Q_OA21 U3809 ( .A0(n3272), .A1(n3273), .B0(n3234), .Z(n4320));
Q_AN02 U3810 ( .A0(n3274), .A1(n3230), .Z(n3272));
Q_AN02 U3811 ( .A0(n3276), .A1(n3233), .Z(n3275));
Q_AO21 U3812 ( .A0(n3277), .A1(n3252), .B0(n3275), .Z(n3273));
Q_OA21 U3813 ( .A0(n3279), .A1(n3277), .B0(n3278), .Z(n4321));
Q_OR02 U3814 ( .A0(n3280), .A1(n3281), .Z(n3277));
Q_OA21 U3815 ( .A0(n3267), .A1(n3282), .B0(n3234), .Z(n4322));
Q_AO21 U3816 ( .A0(n3231), .A1(n3283), .B0(n3243), .Z(n3286));
Q_AN02 U3817 ( .A0(n3284), .A1(n3285), .Z(n3283));
Q_OR02 U3818 ( .A0(n3236), .A1(n3286), .Z(n3282));
Q_AN02 U3819 ( .A0(n3238), .A1(n3287), .Z(n3236));
Q_AN02 U3820 ( .A0(n3288), .A1(ws_read_addr[2]), .Z(n3267));
Q_OA21 U3821 ( .A0(n3289), .A1(n3290), .B0(n3234), .Z(n4323));
Q_AO21 U3822 ( .A0(n3233), .A1(n3292), .B0(n3291), .Z(n3290));
Q_OA21 U3823 ( .A0(n3293), .A1(n3294), .B0(n3234), .Z(n4324));
Q_AO21 U3824 ( .A0(n3233), .A1(n3296), .B0(n3295), .Z(n3294));
Q_OA21 U3825 ( .A0(n3297), .A1(n3298), .B0(n3234), .Z(n4325));
Q_AO21 U3826 ( .A0(n3299), .A1(n3230), .B0(n3300), .Z(n3298));
Q_AN02 U3827 ( .A0(n3233), .A1(n3301), .Z(n3300));
Q_AN02 U3828 ( .A0(n3302), .A1(n3231), .Z(n3297));
Q_AN02 U3829 ( .A0(n3303), .A1(n3304), .Z(n4327));
Q_INV U3830 ( .A(n3305), .Z(n3304));
Q_OA21 U3831 ( .A0(n3289), .A1(n3306), .B0(n3234), .Z(n4328));
Q_AO21 U3832 ( .A0(n3233), .A1(n3307), .B0(n3291), .Z(n3306));
Q_AN02 U3833 ( .A0(n3308), .A1(ws_read_addr[3]), .Z(n3307));
Q_OA21 U3834 ( .A0(n3292), .A1(n3309), .B0(n3231), .Z(n3291));
Q_OA21 U3835 ( .A0(n3293), .A1(n3310), .B0(n3234), .Z(n4329));
Q_AN03 U3836 ( .A0(n3230), .A1(ws_read_addr[4]), .A2(n3311), .Z(n3295));
Q_OR02 U3837 ( .A0(n3295), .A1(n3243), .Z(n3310));
Q_AN02 U3838 ( .A0(n3312), .A1(n3233), .Z(n3243));
Q_OA21 U3839 ( .A0(n3313), .A1(n3314), .B0(n3252), .Z(n3293));
Q_OA21 U3840 ( .A0(n3299), .A1(n3316), .B0(n3315), .Z(n4330));
Q_OR02 U3841 ( .A0(n3317), .A1(n3318), .Z(n3299));
Q_OA21 U3842 ( .A0(n3319), .A1(n3320), .B0(n3278), .Z(n4326));
Q_OR02 U3843 ( .A0(n3321), .A1(n3314), .Z(n3320));
Q_AN02 U3844 ( .A0(n3303), .A1(n3322), .Z(n4331));
Q_AN02 U3845 ( .A0(n3233), .A1(n3234), .Z(n3303));
Q_OA21 U3846 ( .A0(n3323), .A1(n3324), .B0(n3315), .Z(n4332));
Q_NR02 U3847 ( .A0(ws_read_addr[6]), .A1(ws_read_addr[3]), .Z(n3325));
Q_OA21 U3848 ( .A0(n3328), .A1(n3329), .B0(n3325), .Z(n3324));
Q_AN02 U3849 ( .A0(n3330), .A1(n3285), .Z(n3328));
Q_AO21 U3850 ( .A0(n3284), .A1(n3332), .B0(n3331), .Z(n3323));
Q_OA21 U3851 ( .A0(n3333), .A1(n3334), .B0(n3234), .Z(n4333));
Q_OA21 U3852 ( .A0(n3335), .A1(n3336), .B0(ws_read_addr[4]), .Z(n3334));
Q_AN02 U3853 ( .A0(n3233), .A1(n3337), .Z(n3336));
Q_AN02 U3854 ( .A0(n3231), .A1(n3327), .Z(n3335));
Q_OA21 U3855 ( .A0(n3270), .A1(n3338), .B0(n3230), .Z(n3333));
Q_OA21 U3856 ( .A0(n3339), .A1(n3340), .B0(n3234), .Z(n4334));
Q_OA21 U3857 ( .A0(n3341), .A1(n3338), .B0(n3230), .Z(n3339));
Q_AN02 U3858 ( .A0(n3342), .A1(n3343), .Z(n3341));
Q_OA21 U3859 ( .A0(n3344), .A1(n3340), .B0(n3234), .Z(n4335));
Q_AN02 U3860 ( .A0(n3252), .A1(n3345), .Z(n3344));
Q_AN02 U3861 ( .A0(n3330), .A1(n3327), .Z(n3345));
Q_AO21 U3862 ( .A0(n3238), .A1(n3347), .B0(n3346), .Z(n3340));
Q_OA21 U3863 ( .A0(n3289), .A1(n3348), .B0(n3234), .Z(n4336));
Q_AO21 U3864 ( .A0(n3350), .A1(n3268), .B0(n3349), .Z(n3348));
Q_AN02 U3865 ( .A0(n3233), .A1(n3351), .Z(n3346));
Q_AO21 U3866 ( .A0(n3231), .A1(n3309), .B0(n3346), .Z(n3349));
Q_OA21 U3867 ( .A0(n3263), .A1(n3352), .B0(n3230), .Z(n3289));
Q_AN02 U3868 ( .A0(n3308), .A1(n3353), .Z(n3352));
Q_AN02 U3869 ( .A0(n3354), .A1(n3355), .Z(n3263));
Q_INV U3870 ( .A(n3356), .Z(n3354));
Q_OA21 U3871 ( .A0(n3357), .A1(n3358), .B0(n3315), .Z(n4337));
Q_AN02 U3872 ( .A0(n3311), .A1(ws_read_addr[4]), .Z(n3357));
Q_OA21 U3873 ( .A0(n3359), .A1(n3314), .B0(n3326), .Z(n3358));
Q_AO21 U3874 ( .A0(n3355), .A1(n3285), .B0(n3353), .Z(n3311));
Q_AN02 U3875 ( .A0(n3230), .A1(n3234), .Z(n3315));
Q_OA21 U3876 ( .A0(n3360), .A1(n3316), .B0(n3315), .Z(n4338));
Q_AN02 U3877 ( .A0(n3302), .A1(n3361), .Z(n3316));
Q_INV U3878 ( .A(n3362), .Z(n3302));
Q_OR02 U3879 ( .A0(n3363), .A1(n3318), .Z(n3360));
Q_OA21 U3880 ( .A0(n3359), .A1(n3364), .B0(n3278), .Z(n4339));
Q_OR02 U3881 ( .A0(n3321), .A1(n3365), .Z(n3366));
Q_OR02 U3882 ( .A0(n3366), .A1(n3314), .Z(n3364));
Q_AN02 U3883 ( .A0(n3367), .A1(n3288), .Z(n4340));
Q_OA21 U3884 ( .A0(n3368), .A1(n3369), .B0(n3234), .Z(n4341));
Q_OA21 U3885 ( .A0(n3370), .A1(n3371), .B0(n3285), .Z(n3369));
Q_AN02 U3886 ( .A0(n3372), .A1(n3252), .Z(n3370));
Q_OA21 U3887 ( .A0(n3373), .A1(n3374), .B0(n3230), .Z(n3368));
Q_AO21 U3888 ( .A0(n3232), .A1(n3375), .B0(n3376), .Z(n3374));
Q_AN02 U3889 ( .A0(n3377), .A1(n3378), .Z(n3376));
Q_AN02 U3890 ( .A0(n3379), .A1(n3327), .Z(n3373));
Q_OA21 U3891 ( .A0(n3380), .A1(n3381), .B0(n3234), .Z(n4342));
Q_OA21 U3892 ( .A0(n3268), .A1(n3382), .B0(ws_read_addr[3]), .Z(n3381));
Q_AN02 U3893 ( .A0(n3231), .A1(ws_read_addr[4]), .Z(n3268));
Q_OR02 U3894 ( .A0(n3347), .A1(n3287), .Z(n3382));
Q_AN02 U3895 ( .A0(n3233), .A1(ws_read_addr[4]), .Z(n3287));
Q_OA21 U3896 ( .A0(n3383), .A1(n3384), .B0(n3230), .Z(n3380));
Q_AN02 U3897 ( .A0(n3385), .A1(n3386), .Z(n3384));
Q_AN02 U3898 ( .A0(n3238), .A1(n3387), .Z(n3383));
Q_OA21 U3899 ( .A0(n3388), .A1(n3288), .B0(n3234), .Z(n4343));
Q_AN03 U3900 ( .A0(n3230), .A1(n3355), .A2(n3244), .Z(n3389));
Q_AO21 U3901 ( .A0(n3390), .A1(n3252), .B0(n3389), .Z(n3388));
Q_AO21 U3902 ( .A0(n3231), .A1(n3392), .B0(n3391), .Z(n3288));
Q_AN02 U3903 ( .A0(n3278), .A1(n3393), .Z(n4344));
Q_AN02 U3904 ( .A0(n3252), .A1(n3234), .Z(n3278));
Q_AN02 U3905 ( .A0(n3230), .A1(n3326), .Z(n3252));
Q_OA21 U3906 ( .A0(n3394), .A1(n3371), .B0(n3234), .Z(n4345));
Q_AN02 U3907 ( .A0(n3231), .A1(n3296), .Z(n3394));
Q_OR02 U3908 ( .A0(n3347), .A1(n3391), .Z(n3371));
Q_AN02 U3909 ( .A0(n3233), .A1(n3395), .Z(n3391));
Q_AN02 U3910 ( .A0(n3396), .A1(n3397), .Z(n3233));
Q_AN02 U3911 ( .A0(n3231), .A1(n3386), .Z(n3347));
Q_AN02 U3912 ( .A0(n3230), .A1(n3361), .Z(n3231));
Q_AN03 U3913 ( .A0(ws_read_addr[10]), .A1(n3399), .A2(n3398), .Z(n3230));
Q_OA21 U3914 ( .A0(n3401), .A1(n3402), .B0(n3400), .Z(n4346));
Q_AN02 U3915 ( .A0(n3403), .A1(n3404), .Z(n3401));
Q_OR02 U3916 ( .A0(n3405), .A1(n3406), .Z(n3402));
Q_OA21 U3917 ( .A0(n3407), .A1(n3408), .B0(n3400), .Z(n4347));
Q_AN02 U3918 ( .A0(n3409), .A1(ws_read_addr[7]), .Z(n3407));
Q_AO21 U3919 ( .A0(n3411), .A1(n3412), .B0(n3410), .Z(n3408));
Q_OA21 U3920 ( .A0(n3413), .A1(n3414), .B0(n3400), .Z(n4348));
Q_AN02 U3921 ( .A0(n3415), .A1(ws_read_addr[7]), .Z(n3413));
Q_AO21 U3922 ( .A0(n3276), .A1(n3417), .B0(n3416), .Z(n3414));
Q_OA21 U3923 ( .A0(n3418), .A1(n3419), .B0(n3400), .Z(n4349));
Q_AN02 U3924 ( .A0(n3420), .A1(ws_read_addr[7]), .Z(n3418));
Q_OA21 U3925 ( .A0(n3421), .A1(n3419), .B0(n3400), .Z(n4350));
Q_AN02 U3926 ( .A0(n3422), .A1(n3412), .Z(n3421));
Q_OA21 U3927 ( .A0(n3423), .A1(n3424), .B0(n3400), .Z(n4351));
Q_AO21 U3928 ( .A0(n3330), .A1(n3426), .B0(n3427), .Z(n3425));
Q_AN02 U3929 ( .A0(n3428), .A1(n3429), .Z(n3427));
Q_AO21 U3930 ( .A0(n3430), .A1(ws_read_addr[3]), .B0(n3425), .Z(n3424));
Q_AN02 U3931 ( .A0(n3428), .A1(n3292), .Z(n3431));
Q_AO21 U3932 ( .A0(n3417), .A1(n3432), .B0(n3431), .Z(n3430));
Q_OA21 U3933 ( .A0(n3433), .A1(n3434), .B0(n3400), .Z(n4352));
Q_OR03 U3934 ( .A0(n3436), .A1(n3437), .A2(n3435), .Z(n3434));
Q_OA21 U3935 ( .A0(n3438), .A1(n3439), .B0(n3400), .Z(n4353));
Q_AO21 U3936 ( .A0(n3441), .A1(n3412), .B0(n3440), .Z(n3439));
Q_OR02 U3937 ( .A0(n3436), .A1(n3442), .Z(n3440));
Q_OA21 U3938 ( .A0(n3443), .A1(n3444), .B0(n3400), .Z(n4354));
Q_OR03 U3939 ( .A0(n3446), .A1(n3416), .A2(n3445), .Z(n3444));
Q_OA21 U3940 ( .A0(n3447), .A1(n3448), .B0(n3400), .Z(n4355));
Q_AN02 U3941 ( .A0(n3449), .A1(n3412), .Z(n3447));
Q_OR03 U3942 ( .A0(n3436), .A1(n3446), .A2(n3416), .Z(n3448));
Q_OA21 U3943 ( .A0(n3423), .A1(n3450), .B0(n3400), .Z(n4356));
Q_AN02 U3944 ( .A0(n3451), .A1(n3404), .Z(n3423));
Q_AN02 U3945 ( .A0(ws_read_addr[7]), .A1(ws_read_addr[2]), .Z(n3404));
Q_AO21 U3946 ( .A0(n3453), .A1(n3426), .B0(n3452), .Z(n3450));
Q_OA21 U3947 ( .A0(n3454), .A1(n3455), .B0(ws_read_addr[4]), .Z(n3452));
Q_AN02 U3948 ( .A0(n3428), .A1(n3456), .Z(n3455));
Q_OA21 U3949 ( .A0(n3433), .A1(n3457), .B0(n3400), .Z(n4357));
Q_OR03 U3950 ( .A0(n3446), .A1(n3442), .A2(n3435), .Z(n3457));
Q_OA21 U3951 ( .A0(n3438), .A1(n3458), .B0(n3400), .Z(n4358));
Q_OR02 U3952 ( .A0(n3445), .A1(n3459), .Z(n3458));
Q_OA21 U3953 ( .A0(n3443), .A1(n3460), .B0(n3400), .Z(n4359));
Q_OA21 U3954 ( .A0(n3461), .A1(n3462), .B0(ws_read_addr[5]), .Z(n3460));
Q_AN02 U3955 ( .A0(n3463), .A1(n3464), .Z(n3462));
Q_OA21 U3956 ( .A0(n3465), .A1(n3466), .B0(n3400), .Z(n4360));
Q_OR02 U3957 ( .A0(n3459), .A1(n3416), .Z(n3466));
Q_OR02 U3958 ( .A0(n3467), .A1(n3446), .Z(n3459));
Q_AN03 U3959 ( .A0(n3469), .A1(n3226), .A2(n3468), .Z(n4361));
Q_AO21 U3960 ( .A0(n3451), .A1(ws_read_addr[7]), .B0(n3470), .Z(n3468));
Q_OR02 U3961 ( .A0(n3472), .A1(n3473), .Z(n3471));
Q_AO21 U3962 ( .A0(n3474), .A1(n3296), .B0(n3471), .Z(n3470));
Q_OR02 U3963 ( .A0(n3475), .A1(n3476), .Z(n3451));
Q_OA21 U3964 ( .A0(n3433), .A1(n3477), .B0(n3400), .Z(n4362));
Q_OR02 U3965 ( .A0(n3435), .A1(n3478), .Z(n3477));
Q_OA21 U3966 ( .A0(n3479), .A1(n3480), .B0(ws_read_addr[7]), .Z(n3433));
Q_OA21 U3967 ( .A0(n3438), .A1(n3481), .B0(n3400), .Z(n4363));
Q_OR02 U3968 ( .A0(n3445), .A1(n3482), .Z(n3481));
Q_OA21 U3969 ( .A0(n3483), .A1(n3484), .B0(ws_read_addr[7]), .Z(n3438));
Q_OA21 U3970 ( .A0(n3443), .A1(n3485), .B0(n3400), .Z(n4364));
Q_OA21 U3971 ( .A0(n3461), .A1(n3486), .B0(ws_read_addr[5]), .Z(n3485));
Q_AN02 U3972 ( .A0(n3312), .A1(n3464), .Z(n3486));
Q_AN02 U3973 ( .A0(n3312), .A1(n3412), .Z(n3461));
Q_OA21 U3974 ( .A0(n3274), .A1(n3484), .B0(ws_read_addr[7]), .Z(n3443));
Q_OA21 U3975 ( .A0(n3465), .A1(n3487), .B0(n3400), .Z(n4365));
Q_OA21 U3976 ( .A0(n3488), .A1(n3489), .B0(n3400), .Z(n4366));
Q_OA21 U3977 ( .A0(n3490), .A1(n3491), .B0(ws_read_addr[2]), .Z(n3489));
Q_AN02 U3978 ( .A0(n3284), .A1(n3428), .Z(n3491));
Q_AN02 U3979 ( .A0(n3372), .A1(n3412), .Z(n3490));
Q_OA21 U3980 ( .A0(n3492), .A1(n3493), .B0(ws_read_addr[7]), .Z(n3488));
Q_AO21 U3981 ( .A0(n3377), .A1(n3301), .B0(n3494), .Z(n3493));
Q_OA21 U3982 ( .A0(n3495), .A1(n3496), .B0(n3400), .Z(n4367));
Q_AO21 U3983 ( .A0(n3359), .A1(n3412), .B0(n3478), .Z(n3496));
Q_OA21 U3984 ( .A0(n3497), .A1(n3338), .B0(ws_read_addr[7]), .Z(n3495));
Q_OR02 U3985 ( .A0(n3498), .A1(n3499), .Z(n3497));
Q_OA21 U3986 ( .A0(n3465), .A1(n3500), .B0(n3400), .Z(n4368));
Q_OR02 U3987 ( .A0(n3501), .A1(n3502), .Z(n3500));
Q_OA21 U3988 ( .A0(n3504), .A1(n3505), .B0(n3503), .Z(n4369));
Q_OA21 U3989 ( .A0(n3506), .A1(n3312), .B0(ws_read_addr[5]), .Z(n3504));
Q_AN02 U3990 ( .A0(n3400), .A1(n3487), .Z(n4370));
Q_AO21 U3991 ( .A0(n3276), .A1(n3428), .B0(n3467), .Z(n3487));
Q_OA21 U3992 ( .A0(n3507), .A1(n3508), .B0(n3400), .Z(n4371));
Q_OA21 U3993 ( .A0(n3472), .A1(n3509), .B0(n3285), .Z(n3508));
Q_OA21 U3994 ( .A0(n3510), .A1(n3511), .B0(n3400), .Z(n4372));
Q_OR02 U3995 ( .A0(n3512), .A1(n3437), .Z(n3511));
Q_OA21 U3996 ( .A0(n3513), .A1(n3514), .B0(n3412), .Z(n3510));
Q_OA21 U3997 ( .A0(n3501), .A1(n3515), .B0(n3400), .Z(n4373));
Q_OR02 U3998 ( .A0(n3516), .A1(n3442), .Z(n3515));
Q_OA21 U3999 ( .A0(n3517), .A1(n3518), .B0(n3503), .Z(n4374));
Q_OR02 U4000 ( .A0(n3519), .A1(n3514), .Z(n3518));
Q_OA21 U4001 ( .A0(n3520), .A1(n3416), .B0(n3400), .Z(n4375));
Q_AN02 U4002 ( .A0(n3454), .A1(ws_read_addr[4]), .Z(n3520));
Q_AN02 U4003 ( .A0(n3428), .A1(n3337), .Z(n3521));
Q_AO21 U4004 ( .A0(n3417), .A1(n3343), .B0(n3521), .Z(n3454));
Q_OA21 U4005 ( .A0(n3507), .A1(n3522), .B0(n3400), .Z(n4376));
Q_AO21 U4006 ( .A0(n3524), .A1(n3412), .B0(n3523), .Z(n3522));
Q_AO21 U4007 ( .A0(n3526), .A1(n3527), .B0(n3525), .Z(n3524));
Q_OA21 U4008 ( .A0(n3528), .A1(n3529), .B0(n3400), .Z(n4377));
Q_OR02 U4009 ( .A0(n3512), .A1(n3502), .Z(n3529));
Q_AN02 U4010 ( .A0(n3530), .A1(n3412), .Z(n3528));
Q_OR02 U4011 ( .A0(n3513), .A1(n3281), .Z(n3530));
Q_AN02 U4012 ( .A0(n3531), .A1(n3276), .Z(n4380));
Q_OA21 U4013 ( .A0(n3507), .A1(n3532), .B0(n3400), .Z(n4381));
Q_AO21 U4014 ( .A0(n3534), .A1(n3535), .B0(n3533), .Z(n3532));
Q_OA21 U4015 ( .A0(n3536), .A1(n3537), .B0(n3296), .Z(n3533));
Q_AN02 U4016 ( .A0(n3417), .A1(ws_read_addr[2]), .Z(n3536));
Q_OA21 U4017 ( .A0(n3512), .A1(n3538), .B0(n3400), .Z(n4382));
Q_AN02 U4018 ( .A0(n3284), .A1(n3539), .Z(n3540));
Q_OR03 U4019 ( .A0(n3540), .A1(n3442), .A2(n3467), .Z(n3538));
Q_AN03 U4020 ( .A0(n3396), .A1(n3234), .A2(n3541), .Z(n4378));
Q_AN02 U4021 ( .A0(n3543), .A1(n3326), .Z(n3542));
Q_AO21 U4022 ( .A0(n3544), .A1(n3355), .B0(n3542), .Z(n3541));
Q_AN02 U4023 ( .A0(n3396), .A1(n3545), .Z(n3503));
Q_AN02 U4024 ( .A0(n3326), .A1(n3234), .Z(n3545));
Q_AN02 U4025 ( .A0(n3546), .A1(n3547), .Z(n3396));
Q_OA21 U4026 ( .A0(n3519), .A1(n3548), .B0(n3503), .Z(n4379));
Q_OR02 U4027 ( .A0(n3530), .A1(n3359), .Z(n3548));
Q_AN02 U4028 ( .A0(n3531), .A1(n3463), .Z(n4383));
Q_OA21 U4029 ( .A0(n3507), .A1(n3549), .B0(n3400), .Z(n4384));
Q_OR02 U4030 ( .A0(n3550), .A1(n3523), .Z(n3549));
Q_OA21 U4031 ( .A0(n3492), .A1(n3494), .B0(ws_read_addr[7]), .Z(n3507));
Q_AN02 U4032 ( .A0(n3551), .A1(n3327), .Z(n3494));
Q_OA21 U4033 ( .A0(n3552), .A1(n3553), .B0(ws_read_addr[6]), .Z(n3492));
Q_OA21 U4034 ( .A0(n3512), .A1(n3554), .B0(n3400), .Z(n4385));
Q_AN02 U4035 ( .A0(n3556), .A1(n3285), .Z(n3555));
Q_OA21 U4036 ( .A0(n3539), .A1(n3557), .B0(n3327), .Z(n3554));
Q_AN02 U4037 ( .A0(n3474), .A1(n3506), .Z(n3557));
Q_OA21 U4038 ( .A0(n3390), .A1(n3558), .B0(n3555), .Z(n3512));
Q_OA21 U4039 ( .A0(n3501), .A1(n3559), .B0(n3400), .Z(n4386));
Q_AN02 U4040 ( .A0(n3544), .A1(n3560), .Z(n3501));
Q_OA21 U4041 ( .A0(n3561), .A1(n3562), .B0(ws_read_addr[4]), .Z(n3559));
Q_AN02 U4042 ( .A0(n3474), .A1(n3343), .Z(n3562));
Q_AN02 U4043 ( .A0(n3417), .A1(ws_read_addr[3]), .Z(n3561));
Q_OR02 U4044 ( .A0(n3563), .A1(n3564), .Z(n3544));
Q_AN02 U4045 ( .A0(n3469), .A1(n3234), .Z(n3400));
Q_AN02 U4046 ( .A0(n3546), .A1(ws_read_addr[8]), .Z(n3469));
Q_OA21 U4047 ( .A0(n3565), .A1(n3566), .B0(n3400), .Z(n4387));
Q_AN02 U4048 ( .A0(n3567), .A1(n3506), .Z(n3565));
Q_AN02 U4049 ( .A0(n3474), .A1(n3527), .Z(n3568));
Q_AO21 U4050 ( .A0(n3569), .A1(n3412), .B0(n3568), .Z(n3566));
Q_OR02 U4051 ( .A0(n3417), .A1(n3428), .Z(n3474));
Q_OR02 U4052 ( .A0(n3570), .A1(n3514), .Z(n3569));
Q_AN02 U4053 ( .A0(n3531), .A1(n3312), .Z(n4388));
Q_AN02 U4054 ( .A0(n3397), .A1(n3234), .Z(n3571));
Q_AN03 U4055 ( .A0(n3546), .A1(n3572), .A2(n3571), .Z(n3531));
Q_OA21 U4056 ( .A0(n3574), .A1(n3575), .B0(n3573), .Z(n4389));
Q_AN03 U4057 ( .A0(n3572), .A1(n3285), .A2(n3576), .Z(n3577));
Q_AN02 U4058 ( .A0(n3578), .A1(n3328), .Z(n3579));
Q_OR03 U4059 ( .A0(n3579), .A1(n3580), .A2(n3577), .Z(n3575));
Q_OA21 U4060 ( .A0(n3581), .A1(n3582), .B0(ws_read_addr[3]), .Z(n3574));
Q_AN02 U4061 ( .A0(n3583), .A1(n3506), .Z(n3582));
Q_AN02 U4062 ( .A0(n3584), .A1(n3564), .Z(n3581));
Q_OA21 U4063 ( .A0(n3585), .A1(n3586), .B0(n3573), .Z(n4390));
Q_OR02 U4064 ( .A0(n3587), .A1(n3588), .Z(n3585));
Q_OA21 U4065 ( .A0(n3590), .A1(n3591), .B0(n3589), .Z(n4391));
Q_AN02 U4066 ( .A0(n3592), .A1(n3583), .Z(n3591));
Q_OA21 U4067 ( .A0(n3593), .A1(n3594), .B0(n3573), .Z(n4392));
Q_OA21 U4068 ( .A0(n3595), .A1(n3594), .B0(n3573), .Z(n4393));
Q_OR03 U4069 ( .A0(n3597), .A1(n3598), .A2(n3596), .Z(n3594));
Q_AN02 U4070 ( .A0(n3584), .A1(n3599), .Z(n3597));
Q_AN03 U4071 ( .A0(n3546), .A1(n3367), .A2(n3600), .Z(n4394));
Q_AN02 U4072 ( .A0(n3576), .A1(n3572), .Z(n3602));
Q_OR03 U4073 ( .A0(n3602), .A1(n3595), .A2(n3601), .Z(n3600));
Q_OA21 U4074 ( .A0(n3587), .A1(n3603), .B0(n3573), .Z(n4395));
Q_AN03 U4075 ( .A0(n3572), .A1(n3327), .A2(n3576), .Z(n3587));
Q_OR02 U4076 ( .A0(n3588), .A1(n3604), .Z(n3603));
Q_AN02 U4077 ( .A0(n3578), .A1(n3345), .Z(n3588));
Q_AN03 U4078 ( .A0(n3546), .A1(ws_read_addr[4]), .A2(n3234), .Z(n3589));
Q_OA21 U4079 ( .A0(n3590), .A1(n3605), .B0(n3589), .Z(n4396));
Q_AO21 U4080 ( .A0(n3229), .A1(n3572), .B0(n3584), .Z(n3590));
Q_AN02 U4081 ( .A0(n3583), .A1(n3327), .Z(n3605));
Q_OA21 U4082 ( .A0(n3593), .A1(n3606), .B0(n3573), .Z(n4397));
Q_AN02 U4083 ( .A0(n3342), .A1(n3572), .Z(n3593));
Q_OA21 U4084 ( .A0(n3595), .A1(n3606), .B0(n3573), .Z(n4398));
Q_OR02 U4085 ( .A0(n3604), .A1(n3608), .Z(n3607));
Q_AO21 U4086 ( .A0(n3350), .A1(n3609), .B0(n3607), .Z(n3606));
Q_OA21 U4087 ( .A0(n3610), .A1(n3611), .B0(n3573), .Z(n4399));
Q_OA21 U4088 ( .A0(n3612), .A1(n3613), .B0(ws_read_addr[2]), .Z(n3611));
Q_AN02 U4089 ( .A0(n3330), .A1(n3578), .Z(n3595));
Q_OR02 U4090 ( .A0(n3595), .A1(n3608), .Z(n3613));
Q_OA21 U4091 ( .A0(n3609), .A1(n3614), .B0(ws_read_addr[3]), .Z(n3612));
Q_OA21 U4092 ( .A0(n3615), .A1(n3616), .B0(n3572), .Z(n3610));
Q_AO21 U4093 ( .A0(n3330), .A1(n3617), .B0(n3618), .Z(n3616));
Q_AN02 U4094 ( .A0(n3377), .A1(n3527), .Z(n3618));
Q_OA21 U4095 ( .A0(n3619), .A1(n3620), .B0(n3573), .Z(n4400));
Q_AN02 U4096 ( .A0(n3622), .A1(n3578), .Z(n3619));
Q_OR03 U4097 ( .A0(n3623), .A1(n3624), .A2(n3621), .Z(n3620));
Q_AN02 U4098 ( .A0(n3238), .A1(n3614), .Z(n3624));
Q_OA21 U4099 ( .A0(n3625), .A1(n3626), .B0(n3572), .Z(n3621));
Q_AN03 U4100 ( .A0(ws_read_addr[6]), .A1(n3327), .A2(n3330), .Z(n3625));
Q_OA21 U4101 ( .A0(n3627), .A1(n3628), .B0(n3573), .Z(n4401));
Q_AN02 U4102 ( .A0(n3572), .A1(ws_read_addr[4]), .Z(n3629));
Q_OR03 U4103 ( .A0(n3630), .A1(n3631), .A2(n3623), .Z(n3628));
Q_AN02 U4104 ( .A0(n3441), .A1(n3578), .Z(n3627));
Q_OA21 U4105 ( .A0(n3355), .A1(n3240), .B0(n3629), .Z(n3630));
Q_OA21 U4106 ( .A0(n3632), .A1(n3633), .B0(n3573), .Z(n4402));
Q_AO21 U4107 ( .A0(n3312), .A1(n3635), .B0(n3634), .Z(n3633));
Q_OR02 U4108 ( .A0(n3596), .A1(n3598), .Z(n3634));
Q_OA21 U4109 ( .A0(n3636), .A1(n3484), .B0(n3572), .Z(n3632));
Q_AN02 U4110 ( .A0(n3546), .A1(n3234), .Z(n3573));
Q_OA21 U4111 ( .A0(n3637), .A1(n3638), .B0(n3573), .Z(n4403));
Q_AN02 U4112 ( .A0(n3449), .A1(n3578), .Z(n3637));
Q_OR02 U4113 ( .A0(n3639), .A1(n3598), .Z(n3638));
Q_OR02 U4114 ( .A0(n3640), .A1(n3543), .Z(n3449));
Q_AN03 U4115 ( .A0(n3642), .A1(n3226), .A2(n3641), .Z(n4409));
Q_AO21 U4116 ( .A0(n3644), .A1(ws_read_addr[7]), .B0(n3643), .Z(n3641));
Q_AO21 U4117 ( .A0(n3646), .A1(n3412), .B0(n3645), .Z(n3643));
Q_AO21 U4118 ( .A0(n3648), .A1(ws_read_addr[6]), .B0(n3647), .Z(n3644));
Q_OR02 U4119 ( .A0(n3649), .A1(n3650), .Z(n3647));
Q_OR02 U4120 ( .A0(n3651), .A1(n3652), .Z(n3648));
Q_OA21 U4121 ( .A0(n3654), .A1(n3655), .B0(n3653), .Z(n4410));
Q_OR03 U4122 ( .A0(n3657), .A1(n3502), .A2(n3656), .Z(n3655));
Q_OA21 U4123 ( .A0(n3658), .A1(n3480), .B0(ws_read_addr[7]), .Z(n3654));
Q_AN02 U4124 ( .A0(n3659), .A1(ws_read_addr[6]), .Z(n3658));
Q_OA21 U4125 ( .A0(n3660), .A1(n3661), .B0(n3653), .Z(n4411));
Q_OR02 U4126 ( .A0(n3662), .A1(n3657), .Z(n3661));
Q_OA21 U4127 ( .A0(n3483), .A1(n3338), .B0(ws_read_addr[7]), .Z(n3660));
Q_OA21 U4128 ( .A0(n3663), .A1(n3664), .B0(n3653), .Z(n4412));
Q_OA21 U4129 ( .A0(n3662), .A1(n3665), .B0(ws_read_addr[5]), .Z(n3664));
Q_AN02 U4130 ( .A0(n3276), .A1(n3464), .Z(n3665));
Q_OA21 U4131 ( .A0(n3274), .A1(n3338), .B0(ws_read_addr[7]), .Z(n3663));
Q_OA21 U4132 ( .A0(n3666), .A1(n3667), .B0(n3653), .Z(n4413));
Q_OR02 U4133 ( .A0(n3668), .A1(n3502), .Z(n3667));
Q_OA21 U4134 ( .A0(n3359), .A1(n3669), .B0(n3412), .Z(n3666));
Q_OA21 U4135 ( .A0(n3670), .A1(n3671), .B0(n3653), .Z(n4404));
Q_AO21 U4136 ( .A0(n3672), .A1(n3412), .B0(n3406), .Z(n3671));
Q_OA21 U4137 ( .A0(n3673), .A1(n3437), .B0(n3285), .Z(n3406));
Q_OR02 U4138 ( .A0(n3674), .A1(n3675), .Z(n3672));
Q_OA21 U4139 ( .A0(n3676), .A1(n3677), .B0(ws_read_addr[7]), .Z(n3670));
Q_AN02 U4140 ( .A0(n3678), .A1(ws_read_addr[6]), .Z(n3676));
Q_AO21 U4141 ( .A0(n3308), .A1(n3679), .B0(n3499), .Z(n3677));
Q_OA21 U4142 ( .A0(n3680), .A1(n3681), .B0(n3653), .Z(n4405));
Q_AN02 U4143 ( .A0(n3682), .A1(n3683), .Z(n3410));
Q_AO21 U4144 ( .A0(n3684), .A1(n3412), .B0(n3410), .Z(n3681));
Q_INV U4145 ( .A(n3564), .Z(n3682));
Q_OR02 U4146 ( .A0(n3359), .A1(n3685), .Z(n3684));
Q_OA21 U4147 ( .A0(n3686), .A1(n3687), .B0(ws_read_addr[7]), .Z(n3680));
Q_AN02 U4148 ( .A0(n3688), .A1(ws_read_addr[6]), .Z(n3686));
Q_OR02 U4149 ( .A0(n3689), .A1(n3338), .Z(n3687));
Q_OA21 U4150 ( .A0(n3690), .A1(n3691), .B0(n3653), .Z(n4406));
Q_AO21 U4151 ( .A0(n3692), .A1(n3417), .B0(n3416), .Z(n3691));
Q_OA21 U4152 ( .A0(n3693), .A1(n3694), .B0(ws_read_addr[7]), .Z(n3690));
Q_AN02 U4153 ( .A0(n3319), .A1(ws_read_addr[6]), .Z(n3693));
Q_OA21 U4154 ( .A0(n3695), .A1(n3419), .B0(n3653), .Z(n4407));
Q_OA21 U4155 ( .A0(n3696), .A1(n3694), .B0(ws_read_addr[7]), .Z(n3695));
Q_AN02 U4156 ( .A0(n3322), .A1(n3377), .Z(n3694));
Q_OR02 U4157 ( .A0(n3395), .A1(n3312), .Z(n3322));
Q_AN02 U4158 ( .A0(n3642), .A1(n3234), .Z(n3653));
Q_AN02 U4159 ( .A0(n3546), .A1(n3697), .Z(n3642));
Q_AN02 U4160 ( .A0(n3698), .A1(ws_read_addr[9]), .Z(n3546));
Q_OA21 U4161 ( .A0(n3699), .A1(n3419), .B0(n3653), .Z(n4408));
Q_OR02 U4162 ( .A0(n3673), .A1(n3416), .Z(n3419));
Q_AN02 U4163 ( .A0(n3463), .A1(n3428), .Z(n3416));
Q_OR02 U4164 ( .A0(n3296), .A1(n3301), .Z(n3463));
Q_OA21 U4165 ( .A0(n3505), .A1(n3700), .B0(n3412), .Z(n3699));
Q_AN02 U4166 ( .A0(n3692), .A1(n3526), .Z(n3700));
Q_OR02 U4167 ( .A0(n3761), .A1(n3283), .Z(n3692));
Q_AN03 U4168 ( .A0(n3698), .A1(n3367), .A2(n3701), .Z(n4419));
Q_AO21 U4169 ( .A0(n3703), .A1(n3704), .B0(n3702), .Z(n3701));
Q_OR03 U4170 ( .A0(n3707), .A1(n3708), .A2(n3705), .Z(n3702));
Q_AN02 U4171 ( .A0(n3709), .A1(n3599), .Z(n3708));
Q_OA21 U4172 ( .A0(n3345), .A1(n3710), .B0(n3706), .Z(n3707));
Q_OR02 U4173 ( .A0(n3475), .A1(n3711), .Z(n3703));
Q_OA21 U4174 ( .A0(n3713), .A1(n3714), .B0(n3712), .Z(n4420));
Q_AO21 U4175 ( .A0(n3706), .A1(n3716), .B0(n3715), .Z(n3714));
Q_AN02 U4176 ( .A0(n3717), .A1(n3386), .Z(n3716));
Q_OA21 U4177 ( .A0(n3395), .A1(n3309), .B0(n3709), .Z(n3715));
Q_OA21 U4178 ( .A0(n3718), .A1(n3318), .B0(n3704), .Z(n3713));
Q_OA21 U4179 ( .A0(n3719), .A1(n3705), .B0(n3712), .Z(n4421));
Q_OA21 U4180 ( .A0(n3720), .A1(n3721), .B0(n3704), .Z(n3719));
Q_AN02 U4181 ( .A0(n3377), .A1(n3392), .Z(n3721));
Q_OR02 U4182 ( .A0(n3722), .A1(n3650), .Z(n3720));
Q_OA21 U4183 ( .A0(n3723), .A1(n3724), .B0(n3712), .Z(n4422));
Q_OA21 U4184 ( .A0(n3725), .A1(n3726), .B0(ws_read_addr[5]), .Z(n3724));
Q_AN03 U4185 ( .A0(n3728), .A1(ws_read_addr[6]), .A2(n3727), .Z(n3726));
Q_AN02 U4186 ( .A0(n3706), .A1(n3392), .Z(n3725));
Q_OA21 U4187 ( .A0(n3729), .A1(n3730), .B0(n3704), .Z(n3723));
Q_OR02 U4188 ( .A0(n3318), .A1(n3650), .Z(n3730));
Q_OA21 U4189 ( .A0(n3731), .A1(n3732), .B0(n3712), .Z(n4423));
Q_AN02 U4190 ( .A0(n3733), .A1(n3734), .Z(n3731));
Q_AO21 U4191 ( .A0(n3727), .A1(n3709), .B0(n3705), .Z(n3732));
Q_OR02 U4192 ( .A0(n3735), .A1(n3309), .Z(n3727));
Q_AN02 U4193 ( .A0(n3709), .A1(n3395), .Z(n3736));
Q_AO21 U4194 ( .A0(n3734), .A1(n3392), .B0(n3736), .Z(n3705));
Q_OA21 U4195 ( .A0(n3737), .A1(n3738), .B0(n3712), .Z(n4414));
Q_AN02 U4196 ( .A0(n3740), .A1(n3709), .Z(n3739));
Q_AO21 U4197 ( .A0(n3741), .A1(n3706), .B0(n3739), .Z(n3738));
Q_OR02 U4198 ( .A0(n3313), .A1(n3329), .Z(n3741));
Q_OA21 U4199 ( .A0(n3742), .A1(n3743), .B0(n3704), .Z(n3737));
Q_AO21 U4200 ( .A0(n3284), .A1(n3744), .B0(n3729), .Z(n3743));
Q_OA21 U4201 ( .A0(n3525), .A1(n3745), .B0(ws_read_addr[6]), .Z(n3742));
Q_OA21 U4202 ( .A0(n3746), .A1(n3747), .B0(n3712), .Z(n4415));
Q_AO21 U4203 ( .A0(n3749), .A1(n3734), .B0(n3748), .Z(n3747));
Q_OA21 U4204 ( .A0(n3761), .A1(n3309), .B0(n3709), .Z(n3748));
Q_OA21 U4205 ( .A0(n3479), .A1(n3750), .B0(n3704), .Z(n3746));
Q_OR02 U4206 ( .A0(n3751), .A1(n3650), .Z(n3750));
Q_OA21 U4207 ( .A0(n3752), .A1(n3753), .B0(n3712), .Z(n4416));
Q_AO21 U4208 ( .A0(n3244), .A1(n3734), .B0(n3754), .Z(n3753));
Q_OA21 U4209 ( .A0(n3483), .A1(n3755), .B0(n3704), .Z(n3752));
Q_OA21 U4210 ( .A0(n3756), .A1(n3757), .B0(n3712), .Z(n4417));
Q_OA21 U4211 ( .A0(n3758), .A1(n3751), .B0(n3704), .Z(n3756));
Q_OR02 U4212 ( .A0(n3317), .A1(n3755), .Z(n3758));
Q_AN02 U4213 ( .A0(n3649), .A1(n3285), .Z(n3751));
Q_AN02 U4214 ( .A0(n3698), .A1(n3234), .Z(n3712));
Q_OA21 U4215 ( .A0(n3759), .A1(n3757), .B0(n3712), .Z(n4418));
Q_AN02 U4216 ( .A0(n3704), .A1(n3326), .Z(n3706));
Q_OA21 U4217 ( .A0(n3283), .A1(n3309), .B0(n3709), .Z(n3754));
Q_AO21 U4218 ( .A0(n3709), .A1(n3761), .B0(n3754), .Z(n3760));
Q_AN02 U4219 ( .A0(n3238), .A1(ws_read_addr[4]), .Z(n3761));
Q_OR03 U4220 ( .A0(n3762), .A1(n3763), .A2(n3760), .Z(n3757));
Q_AN02 U4221 ( .A0(n3709), .A1(n3255), .Z(n3763));
Q_AN02 U4222 ( .A0(n3728), .A1(n3397), .Z(n3709));
Q_AN02 U4223 ( .A0(n3399), .A1(n3547), .Z(n3728));
Q_AN02 U4224 ( .A0(n3734), .A1(n3256), .Z(n3762));
Q_AN02 U4225 ( .A0(n3704), .A1(n3361), .Z(n3734));
Q_AN02 U4226 ( .A0(ws_read_addr[9]), .A1(n3398), .Z(n3704));
Q_OA21 U4227 ( .A0(n3390), .A1(n3764), .B0(n3706), .Z(n3759));
Q_OA21 U4228 ( .A0(n3766), .A1(n3767), .B0(n3765), .Z(n4424));
Q_AO21 U4229 ( .A0(n3769), .A1(n3417), .B0(n3768), .Z(n3767));
Q_OR02 U4230 ( .A0(n3506), .A1(n3770), .Z(n3769));
Q_OA21 U4231 ( .A0(n3771), .A1(n3772), .B0(n3765), .Z(n4425));
Q_OR02 U4232 ( .A0(n3773), .A1(n3437), .Z(n3772));
Q_AN02 U4233 ( .A0(n3428), .A1(n3296), .Z(n3437));
Q_AN02 U4234 ( .A0(n3774), .A1(n3417), .Z(n3771));
Q_INV U4235 ( .A(n3733), .Z(n3774));
Q_OA21 U4236 ( .A0(n3775), .A1(n3776), .B0(n3765), .Z(n4426));
Q_AO21 U4237 ( .A0(n3777), .A1(n3417), .B0(n3473), .Z(n3776));
Q_OA21 U4238 ( .A0(n3778), .A1(n3645), .B0(n3765), .Z(n4427));
Q_OA21 U4239 ( .A0(n3779), .A1(n3645), .B0(n3765), .Z(n4428));
Q_OA21 U4240 ( .A0(n3543), .A1(n3780), .B0(n3412), .Z(n3779));
Q_AN02 U4241 ( .A0(n3777), .A1(n3526), .Z(n3780));
Q_OA21 U4242 ( .A0(n3781), .A1(n3782), .B0(n3765), .Z(n4429));
Q_OR02 U4243 ( .A0(n3784), .A1(n3442), .Z(n3783));
Q_AN02 U4244 ( .A0(n3428), .A1(n3301), .Z(n3442));
Q_AO21 U4245 ( .A0(n3673), .A1(n3285), .B0(n3783), .Z(n3782));
Q_OA21 U4246 ( .A0(n3785), .A1(n3786), .B0(n3765), .Z(n4430));
Q_OR02 U4247 ( .A0(n3787), .A1(n3788), .Z(n3786));
Q_OA21 U4248 ( .A0(n3789), .A1(n3790), .B0(n3765), .Z(n4431));
Q_OR02 U4249 ( .A0(n3791), .A1(n3792), .Z(n3790));
Q_OA21 U4250 ( .A0(n3794), .A1(n3795), .B0(n3793), .Z(n4432));
Q_AN02 U4251 ( .A0(n3797), .A1(n3464), .Z(n3795));
Q_AO21 U4252 ( .A0(n3412), .A1(n3392), .B0(n3796), .Z(n3794));
Q_OA21 U4253 ( .A0(n3798), .A1(n3799), .B0(n3765), .Z(n4433));
Q_AO21 U4254 ( .A0(n3797), .A1(n3428), .B0(n3792), .Z(n3799));
Q_AO21 U4255 ( .A0(n3350), .A1(n3801), .B0(n3800), .Z(n3792));
Q_OA21 U4256 ( .A0(n3781), .A1(n3802), .B0(n3765), .Z(n4434));
Q_OA21 U4257 ( .A0(n3804), .A1(n3711), .B0(n3803), .Z(n3781));
Q_AN02 U4258 ( .A0(n3232), .A1(n3377), .Z(n3711));
Q_AN02 U4259 ( .A0(n3646), .A1(ws_read_addr[6]), .Z(n3804));
Q_OR02 U4260 ( .A0(n3390), .A1(n3805), .Z(n3646));
Q_OA21 U4261 ( .A0(n3785), .A1(n3806), .B0(n3765), .Z(n4435));
Q_OR02 U4262 ( .A0(n3787), .A1(n3478), .Z(n3806));
Q_AN02 U4263 ( .A0(n3330), .A1(n3807), .Z(n3787));
Q_OA21 U4264 ( .A0(n3808), .A1(n3318), .B0(ws_read_addr[7]), .Z(n3785));
Q_AN02 U4265 ( .A0(n3362), .A1(n3355), .Z(n3808));
Q_OR02 U4266 ( .A0(n3395), .A1(n3770), .Z(n3362));
Q_OA21 U4267 ( .A0(n3789), .A1(n3809), .B0(n3765), .Z(n4436));
Q_OR02 U4268 ( .A0(n3791), .A1(n3810), .Z(n3809));
Q_OA21 U4269 ( .A0(n3811), .A1(n3650), .B0(ws_read_addr[7]), .Z(n3789));
Q_AN02 U4270 ( .A0(n3377), .A1(n3599), .Z(n3650));
Q_AN02 U4271 ( .A0(n3812), .A1(n3355), .Z(n3811));
Q_INV U4272 ( .A(n3749), .Z(n3812));
Q_NR02 U4273 ( .A0(n3238), .A1(ws_read_addr[4]), .Z(n3770));
Q_AN03 U4274 ( .A0(ws_read_addr[5]), .A1(n3234), .A2(n3813), .Z(n3793));
Q_OA21 U4275 ( .A0(n3796), .A1(n3814), .B0(n3793), .Z(n4437));
Q_AN02 U4276 ( .A0(n3232), .A1(n3412), .Z(n3796));
Q_OA21 U4277 ( .A0(n3807), .A1(n3815), .B0(n3386), .Z(n3814));
Q_AN02 U4278 ( .A0(n3464), .A1(ws_read_addr[3]), .Z(n3815));
Q_AN02 U4279 ( .A0(n3412), .A1(n3327), .Z(n3807));
Q_OA21 U4280 ( .A0(n3798), .A1(n3816), .B0(n3765), .Z(n4438));
Q_OA21 U4281 ( .A0(n3817), .A1(n3802), .B0(n3765), .Z(n4439));
Q_AO21 U4282 ( .A0(n3740), .A1(n3428), .B0(n3784), .Z(n3802));
Q_AN02 U4283 ( .A0(n3372), .A1(n3818), .Z(n3784));
Q_OR02 U4284 ( .A0(n3506), .A1(n3378), .Z(n3740));
Q_OA21 U4285 ( .A0(n3819), .A1(n3820), .B0(ws_read_addr[7]), .Z(n3817));
Q_OA21 U4286 ( .A0(n3821), .A1(n3378), .B0(n3377), .Z(n3820));
Q_AN03 U4287 ( .A0(n3813), .A1(n3823), .A2(n3822), .Z(n4440));
Q_AN02 U4288 ( .A0(ws_read_addr[3]), .A1(n3234), .Z(n3823));
Q_AO21 U4289 ( .A0(n3825), .A1(ws_read_addr[7]), .B0(n3824), .Z(n3822));
Q_AO21 U4290 ( .A0(n3428), .A1(n3386), .B0(n3798), .Z(n3826));
Q_AO21 U4291 ( .A0(n3827), .A1(ws_read_addr[2]), .B0(n3826), .Z(n3824));
Q_OR02 U4292 ( .A0(n3387), .A1(n3829), .Z(n3828));
Q_AO21 U4293 ( .A0(n3342), .A1(ws_read_addr[2]), .B0(n3828), .Z(n3825));
Q_OA21 U4294 ( .A0(n3830), .A1(n3831), .B0(n3765), .Z(n4441));
Q_OR02 U4295 ( .A0(n3516), .A1(n3832), .Z(n3831));
Q_AN02 U4296 ( .A0(n3390), .A1(n3412), .Z(n3516));
Q_OA21 U4297 ( .A0(n3834), .A1(n3390), .B0(n3833), .Z(n4442));
Q_OA21 U4298 ( .A0(n3292), .A1(n3599), .B0(ws_read_addr[5]), .Z(n3834));
Q_OA21 U4299 ( .A0(n3835), .A1(n3816), .B0(n3765), .Z(n4443));
Q_AN02 U4300 ( .A0(n3417), .A1(n3296), .Z(n3835));
Q_OA21 U4301 ( .A0(n3836), .A1(n3837), .B0(n3765), .Z(n4444));
Q_AO21 U4302 ( .A0(n3839), .A1(ws_read_addr[4]), .B0(n3838), .Z(n3837));
Q_OR02 U4303 ( .A0(n3840), .A1(n3841), .Z(n3839));
Q_OA21 U4304 ( .A0(n3819), .A1(n3842), .B0(ws_read_addr[7]), .Z(n3836));
Q_OA21 U4305 ( .A0(n3843), .A1(n3256), .B0(n3377), .Z(n3842));
Q_AN02 U4306 ( .A0(n3844), .A1(ws_read_addr[3]), .Z(n3843));
Q_OA21 U4307 ( .A0(n3845), .A1(n3846), .B0(n3765), .Z(n4445));
Q_OA21 U4308 ( .A0(n3847), .A1(n3848), .B0(ws_read_addr[4]), .Z(n3846));
Q_OA21 U4309 ( .A0(n3849), .A1(n3850), .B0(ws_read_addr[7]), .Z(n3845));
Q_OR02 U4310 ( .A0(n3851), .A1(n3721), .Z(n3850));
Q_OA21 U4311 ( .A0(n3830), .A1(n3852), .B0(n3765), .Z(n4446));
Q_OR02 U4312 ( .A0(n3798), .A1(n3473), .Z(n3852));
Q_OA21 U4313 ( .A0(n3853), .A1(n3849), .B0(ws_read_addr[7]), .Z(n3830));
Q_AN02 U4314 ( .A0(n3342), .A1(n3854), .Z(n3849));
Q_OA21 U4315 ( .A0(n3517), .A1(n3855), .B0(n3833), .Z(n4447));
Q_AN02 U4316 ( .A0(n3856), .A1(ws_read_addr[5]), .Z(n3517));
Q_INV U4317 ( .A(n3857), .Z(n3856));
Q_AN02 U4318 ( .A0(n3765), .A1(n3816), .Z(n4448));
Q_OR02 U4319 ( .A0(n3858), .A1(n3832), .Z(n3816));
Q_OA21 U4320 ( .A0(n3859), .A1(n3860), .B0(n3765), .Z(n4449));
Q_OA21 U4321 ( .A0(n3861), .A1(n3829), .B0(n3803), .Z(n3859));
Q_OA21 U4322 ( .A0(n3862), .A1(n3482), .B0(n3765), .Z(n4450));
Q_OA21 U4323 ( .A0(n3387), .A1(n3864), .B0(n3863), .Z(n3862));
Q_AN02 U4324 ( .A0(n3865), .A1(n3386), .Z(n3864));
Q_OA21 U4325 ( .A0(n3866), .A1(n3810), .B0(n3765), .Z(n4451));
Q_OR02 U4326 ( .A0(n3858), .A1(n3478), .Z(n3810));
Q_OA21 U4327 ( .A0(n3853), .A1(n3867), .B0(ws_read_addr[7]), .Z(n3866));
Q_AN02 U4328 ( .A0(n3865), .A1(n3599), .Z(n3867));
Q_OR02 U4329 ( .A0(n3375), .A1(n3744), .Z(n3865));
Q_AN02 U4330 ( .A0(n3377), .A1(n3285), .Z(n3744));
Q_OA21 U4331 ( .A0(n3791), .A1(n3868), .B0(n3765), .Z(n4452));
Q_OR03 U4332 ( .A0(n3467), .A1(n3478), .A2(n3858), .Z(n3868));
Q_AN02 U4333 ( .A0(n3827), .A1(n3854), .Z(n3858));
Q_AN02 U4334 ( .A0(n3238), .A1(n3798), .Z(n3467));
Q_AN02 U4335 ( .A0(n3417), .A1(ws_read_addr[4]), .Z(n3798));
Q_OR02 U4336 ( .A0(n3801), .A1(n3509), .Z(n3827));
Q_OA21 U4337 ( .A0(n3869), .A1(n3870), .B0(n3765), .Z(n4454));
Q_AO21 U4338 ( .A0(n3871), .A1(n3395), .B0(n3838), .Z(n3870));
Q_OR02 U4339 ( .A0(n3840), .A1(n3872), .Z(n3871));
Q_AN02 U4340 ( .A0(n3417), .A1(n3285), .Z(n3840));
Q_OA21 U4341 ( .A0(n3498), .A1(n3873), .B0(ws_read_addr[7]), .Z(n3869));
Q_AN02 U4342 ( .A0(n3390), .A1(n3617), .Z(n3498));
Q_OA21 U4343 ( .A0(n3270), .A1(n3874), .B0(n3327), .Z(n3873));
Q_AN02 U4344 ( .A0(n3377), .A1(n3432), .Z(n3874));
Q_AN02 U4345 ( .A0(n3355), .A1(n3292), .Z(n3270));
Q_OA21 U4346 ( .A0(n3875), .A1(n3876), .B0(n3765), .Z(n4455));
Q_OR02 U4347 ( .A0(n3877), .A1(n3473), .Z(n3876));
Q_AN02 U4348 ( .A0(n3428), .A1(n3599), .Z(n3473));
Q_OA21 U4349 ( .A0(n3851), .A1(n3878), .B0(ws_read_addr[7]), .Z(n3875));
Q_AN02 U4350 ( .A0(n3355), .A1(n3395), .Z(n3851));
Q_OA21 U4351 ( .A0(n3879), .A1(n3832), .B0(n3765), .Z(n4456));
Q_OA21 U4352 ( .A0(n3853), .A1(n3878), .B0(ws_read_addr[7]), .Z(n3879));
Q_OA21 U4353 ( .A0(n3718), .A1(n3353), .B0(n3432), .Z(n3878));
Q_AN02 U4354 ( .A0(n3377), .A1(n3327), .Z(n3353));
Q_OA21 U4355 ( .A0(n3880), .A1(n3877), .B0(n3765), .Z(n4457));
Q_AN02 U4356 ( .A0(n3881), .A1(n3428), .Z(n3832));
Q_OR02 U4357 ( .A0(n3550), .A1(n3832), .Z(n3880));
Q_OA21 U4358 ( .A0(n3882), .A1(n3860), .B0(n3765), .Z(n4458));
Q_OR02 U4359 ( .A0(n3877), .A1(n3838), .Z(n3860));
Q_AN02 U4360 ( .A0(n3735), .A1(n3428), .Z(n3838));
Q_AN02 U4361 ( .A0(n3883), .A1(n3506), .Z(n3877));
Q_OA21 U4362 ( .A0(n3819), .A1(n3884), .B0(ws_read_addr[7]), .Z(n3882));
Q_AN02 U4363 ( .A0(n3350), .A1(n3829), .Z(n3884));
Q_AN02 U4364 ( .A0(n3377), .A1(n3386), .Z(n3829));
Q_OA21 U4365 ( .A0(n3885), .A1(n3482), .B0(n3765), .Z(n4459));
Q_AN02 U4366 ( .A0(n3886), .A1(ws_read_addr[4]), .Z(n3482));
Q_AN02 U4367 ( .A0(ws_read_addr[7]), .A1(ws_read_addr[3]), .Z(n3863));
Q_OR02 U4368 ( .A0(n3887), .A1(n3848), .Z(n3886));
Q_OA21 U4369 ( .A0(n3387), .A1(n3888), .B0(n3863), .Z(n3885));
Q_AN02 U4370 ( .A0(n3229), .A1(n3432), .Z(n3888));
Q_OA21 U4371 ( .A0(n3889), .A1(n3890), .B0(n3765), .Z(n4460));
Q_OA21 U4372 ( .A0(n3891), .A1(n3848), .B0(ws_read_addr[4]), .Z(n3890));
Q_OA21 U4373 ( .A0(n3853), .A1(n3892), .B0(ws_read_addr[7]), .Z(n3889));
Q_AN02 U4374 ( .A0(n3229), .A1(n3301), .Z(n3892));
Q_AN02 U4375 ( .A0(n3355), .A1(n3296), .Z(n3853));
Q_OR02 U4376 ( .A0(n3355), .A1(n3377), .Z(n3229));
Q_OA21 U4377 ( .A0(n3791), .A1(n3893), .B0(n3765), .Z(n4461));
Q_OA21 U4378 ( .A0(n3886), .A1(n3891), .B0(ws_read_addr[4]), .Z(n3893));
Q_AN02 U4379 ( .A0(n3238), .A1(n3428), .Z(n3848));
Q_AN02 U4380 ( .A0(n3428), .A1(n3854), .Z(n3841));
Q_AO21 U4381 ( .A0(n3417), .A1(n3456), .B0(n3841), .Z(n3891));
Q_AN03 U4382 ( .A0(n3599), .A1(n3234), .A2(n3894), .Z(n4453));
Q_OA21 U4383 ( .A0(n3895), .A1(n3896), .B0(n3765), .Z(n4462));
Q_AO21 U4384 ( .A0(n3417), .A1(n3292), .B0(n3897), .Z(n3896));
Q_OA21 U4385 ( .A0(n3819), .A1(n3898), .B0(ws_read_addr[7]), .Z(n3895));
Q_AN02 U4386 ( .A0(n3372), .A1(n3617), .Z(n3819));
Q_OA21 U4387 ( .A0(n3899), .A1(n3900), .B0(n3386), .Z(n3898));
Q_AN02 U4388 ( .A0(n3377), .A1(n3343), .Z(n3900));
Q_AN02 U4389 ( .A0(n3355), .A1(n3337), .Z(n3899));
Q_OA21 U4390 ( .A0(n3901), .A1(n3902), .B0(n3765), .Z(n4463));
Q_OR02 U4391 ( .A0(n3550), .A1(n3788), .Z(n3902));
Q_AN02 U4392 ( .A0(n3903), .A1(n3683), .Z(n3788));
Q_AN02 U4393 ( .A0(n3390), .A1(n3818), .Z(n3550));
Q_AN02 U4394 ( .A0(n3412), .A1(n3285), .Z(n3818));
Q_INV U4395 ( .A(n3432), .Z(n3903));
Q_OA21 U4396 ( .A0(n3904), .A1(n3905), .B0(n3765), .Z(n4464));
Q_AN02 U4397 ( .A0(n3883), .A1(ws_read_addr[4]), .Z(n3905));
Q_OR02 U4398 ( .A0(n3847), .A1(n3683), .Z(n3883));
Q_AN02 U4399 ( .A0(n3417), .A1(n3327), .Z(n3847));
Q_OA21 U4400 ( .A0(n3906), .A1(n3907), .B0(n3765), .Z(n4465));
Q_AO21 U4401 ( .A0(n3567), .A1(n3432), .B0(n3800), .Z(n3907));
Q_AN02 U4402 ( .A0(n3908), .A1(n3797), .Z(n4466));
Q_OA21 U4403 ( .A0(n3909), .A1(n3910), .B0(n3765), .Z(n4467));
Q_AN02 U4404 ( .A0(ws_read_addr[7]), .A1(n3285), .Z(n3803));
Q_AN02 U4405 ( .A0(n3308), .A1(n3683), .Z(n3897));
Q_AO21 U4406 ( .A0(n3911), .A1(n3412), .B0(n3897), .Z(n3910));
Q_AO21 U4407 ( .A0(n3526), .A1(n3429), .B0(n3552), .Z(n3911));
Q_AO21 U4408 ( .A0(ws_read_addr[5]), .A1(n3309), .B0(n3912), .Z(n3552));
Q_OA21 U4409 ( .A0(n3861), .A1(n3913), .B0(n3803), .Z(n3909));
Q_AN02 U4410 ( .A0(n3372), .A1(ws_read_addr[6]), .Z(n3861));
Q_OR02 U4411 ( .A0(n3914), .A1(n3318), .Z(n3913));
Q_OR02 U4412 ( .A0(n3390), .A1(n3365), .Z(n3372));
Q_OA21 U4413 ( .A0(n3901), .A1(n3915), .B0(n3765), .Z(n4468));
Q_AN02 U4414 ( .A0(n3560), .A1(ws_read_addr[3]), .Z(n3901));
Q_AN02 U4415 ( .A0(n3284), .A1(n3872), .Z(n3523));
Q_AN02 U4416 ( .A0(n3428), .A1(ws_read_addr[2]), .Z(n3872));
Q_AO21 U4417 ( .A0(n3366), .A1(n3412), .B0(n3523), .Z(n3915));
Q_OA21 U4418 ( .A0(n3906), .A1(n3916), .B0(n3765), .Z(n4469));
Q_AN02 U4419 ( .A0(n3284), .A1(n3560), .Z(n3904));
Q_OR02 U4420 ( .A0(n3904), .A1(n3917), .Z(n3916));
Q_AN02 U4421 ( .A0(n3319), .A1(n3412), .Z(n3906));
Q_OR02 U4422 ( .A0(n3313), .A1(n3365), .Z(n3319));
Q_AN03 U4423 ( .A0(n3918), .A1(n3547), .A2(n3545), .Z(n3833));
Q_AN02 U4424 ( .A0(ws_read_addr[8]), .A1(ws_read_addr[7]), .Z(n3547));
Q_OA21 U4425 ( .A0(n3919), .A1(n3313), .B0(n3833), .Z(n4470));
Q_OR02 U4426 ( .A0(n3920), .A1(n3366), .Z(n3919));
Q_AN02 U4427 ( .A0(n3894), .A1(n3234), .Z(n3908));
Q_AN02 U4428 ( .A0(n3921), .A1(n3397), .Z(n3894));
Q_OA21 U4429 ( .A0(n3395), .A1(n3797), .B0(n3908), .Z(n4471));
Q_OR02 U4430 ( .A0(n3563), .A1(n3378), .Z(n3797));
Q_OA21 U4431 ( .A0(n3922), .A1(n3923), .B0(n3765), .Z(n4472));
Q_OR02 U4432 ( .A0(n3405), .A1(n3768), .Z(n3923));
Q_AN02 U4433 ( .A0(n3232), .A1(n3537), .Z(n3768));
Q_AN02 U4434 ( .A0(n3428), .A1(n3285), .Z(n3537));
Q_AN02 U4435 ( .A0(n3924), .A1(n3426), .Z(n3405));
Q_OA21 U4436 ( .A0(n3656), .A1(n3925), .B0(n3765), .Z(n4473));
Q_OR02 U4437 ( .A0(n3926), .A1(n3683), .Z(n3925));
Q_AN02 U4438 ( .A0(n3428), .A1(ws_read_addr[3]), .Z(n3683));
Q_OA21 U4439 ( .A0(n3927), .A1(n3928), .B0(n3765), .Z(n4474));
Q_OR02 U4440 ( .A0(n3929), .A1(n3800), .Z(n3928));
Q_OA21 U4441 ( .A0(n3930), .A1(n3931), .B0(n3765), .Z(n4475));
Q_OA21 U4442 ( .A0(n3662), .A1(n3932), .B0(ws_read_addr[5]), .Z(n3931));
Q_AN02 U4443 ( .A0(n3284), .A1(n3464), .Z(n3932));
Q_OA21 U4444 ( .A0(n3933), .A1(n3645), .B0(n3765), .Z(n4476));
Q_OA21 U4445 ( .A0(n3922), .A1(n3934), .B0(n3765), .Z(n4477));
Q_OA21 U4446 ( .A0(n3935), .A1(n3645), .B0(ws_read_addr[2]), .Z(n3934));
Q_AN02 U4447 ( .A0(n3924), .A1(n3412), .Z(n3935));
Q_OA21 U4448 ( .A0(n3936), .A1(n3264), .B0(ws_read_addr[7]), .Z(n3922));
Q_AN02 U4449 ( .A0(n3232), .A1(n3332), .Z(n3264));
Q_OA21 U4450 ( .A0(n3937), .A1(n3938), .B0(n3765), .Z(n4478));
Q_OR02 U4451 ( .A0(n3926), .A1(n3939), .Z(n3937));
Q_OR02 U4452 ( .A0(n3656), .A1(n3502), .Z(n3938));
Q_AN02 U4453 ( .A0(n3312), .A1(n3428), .Z(n3502));
Q_OA21 U4454 ( .A0(n3718), .A1(n3484), .B0(ws_read_addr[7]), .Z(n3926));
Q_OA21 U4455 ( .A0(n3929), .A1(n3940), .B0(n3765), .Z(n4479));
Q_AN02 U4456 ( .A0(n3659), .A1(n3412), .Z(n3927));
Q_OR03 U4457 ( .A0(n3939), .A1(n3917), .A2(n3927), .Z(n3940));
Q_AN02 U4458 ( .A0(n3428), .A1(n3378), .Z(n3917));
Q_OR02 U4459 ( .A0(n3640), .A1(n3941), .Z(n3659));
Q_OA21 U4460 ( .A0(n3722), .A1(n3338), .B0(ws_read_addr[7]), .Z(n3929));
Q_OA21 U4461 ( .A0(n3930), .A1(n3942), .B0(n3765), .Z(n4480));
Q_OA21 U4462 ( .A0(n3662), .A1(n3943), .B0(ws_read_addr[5]), .Z(n3942));
Q_AN03 U4463 ( .A0(n3412), .A1(n3386), .A2(n3238), .Z(n3662));
Q_OA21 U4464 ( .A0(n3761), .A1(n3944), .B0(n3464), .Z(n3943));
Q_OA21 U4465 ( .A0(n3945), .A1(n3338), .B0(ws_read_addr[7]), .Z(n3930));
Q_OA21 U4466 ( .A0(n3933), .A1(n3946), .B0(n3765), .Z(n4481));
Q_AN02 U4467 ( .A0(n3947), .A1(n3412), .Z(n3933));
Q_OR03 U4468 ( .A0(n3478), .A1(n3948), .A2(n3939), .Z(n3946));
Q_AN02 U4469 ( .A0(n3673), .A1(ws_read_addr[2]), .Z(n3939));
Q_AO21 U4470 ( .A0(n3417), .A1(n3392), .B0(n3800), .Z(n3673));
Q_OA21 U4471 ( .A0(n3766), .A1(n3949), .B0(n3765), .Z(n4482));
Q_OA21 U4472 ( .A0(n3417), .A1(n3645), .B0(ws_read_addr[2]), .Z(n3949));
Q_AN02 U4473 ( .A0(n3232), .A1(n3428), .Z(n3645));
Q_OA21 U4474 ( .A0(n3936), .A1(n3332), .B0(ws_read_addr[7]), .Z(n3766));
Q_AN02 U4475 ( .A0(n3377), .A1(ws_read_addr[2]), .Z(n3332));
Q_AN02 U4476 ( .A0(n3924), .A1(n3617), .Z(n3936));
Q_AN02 U4477 ( .A0(ws_read_addr[6]), .A1(n3285), .Z(n3617));
Q_OA21 U4478 ( .A0(n3950), .A1(n3951), .B0(n3765), .Z(n4483));
Q_OR02 U4479 ( .A0(n3773), .A1(n3887), .Z(n3950));
Q_AN02 U4480 ( .A0(n3238), .A1(n3417), .Z(n3887));
Q_OA21 U4481 ( .A0(n3761), .A1(n3378), .B0(n3428), .Z(n3951));
Q_OA21 U4482 ( .A0(n3718), .A1(n3240), .B0(ws_read_addr[7]), .Z(n3773));
Q_AN02 U4483 ( .A0(n3238), .A1(n3377), .Z(n3240));
Q_OA21 U4484 ( .A0(n3775), .A1(n3952), .B0(n3765), .Z(n4484));
Q_OR02 U4485 ( .A0(n3953), .A1(n3948), .Z(n3952));
Q_OA21 U4486 ( .A0(n3722), .A1(n3246), .B0(ws_read_addr[7]), .Z(n3775));
Q_OA21 U4487 ( .A0(n3778), .A1(n3954), .B0(n3765), .Z(n4485));
Q_AN02 U4488 ( .A0(n3249), .A1(ws_read_addr[7]), .Z(n3778));
Q_OR02 U4489 ( .A0(n3945), .A1(n3246), .Z(n3249));
Q_AN02 U4490 ( .A0(n3244), .A1(n3377), .Z(n3246));
Q_AN02 U4491 ( .A0(n3813), .A1(n3234), .Z(n3765));
Q_AN02 U4492 ( .A0(n3918), .A1(ws_read_addr[8]), .Z(n3813));
Q_OA21 U4493 ( .A0(n3955), .A1(n3954), .B0(n3765), .Z(n4486));
Q_AN02 U4494 ( .A0(n3251), .A1(n3412), .Z(n3955));
Q_OR02 U4495 ( .A0(n3668), .A1(n3948), .Z(n3954));
Q_AN02 U4496 ( .A0(n3944), .A1(n3428), .Z(n3948));
Q_OR02 U4497 ( .A0(n3312), .A1(n3378), .Z(n3944));
Q_OR02 U4498 ( .A0(n3657), .A1(n3478), .Z(n3668));
Q_AN02 U4499 ( .A0(n3238), .A1(n3509), .Z(n3478));
Q_AN02 U4500 ( .A0(n3428), .A1(ws_read_addr[4]), .Z(n3509));
Q_OR02 U4501 ( .A0(n3543), .A1(n3764), .Z(n3251));
Q_AN02 U4502 ( .A0(n3244), .A1(n3526), .Z(n3764));
Q_OA21 U4503 ( .A0(n3957), .A1(n3958), .B0(n3956), .Z(n4487));
Q_AO21 U4504 ( .A0(n3924), .A1(n3960), .B0(n3631), .Z(n3959));
Q_AO21 U4505 ( .A0(n3961), .A1(ws_read_addr[2]), .B0(n3959), .Z(n3958));
Q_OA21 U4506 ( .A0(n3962), .A1(n3963), .B0(n3572), .Z(n3957));
Q_OA21 U4507 ( .A0(n3674), .A1(n3685), .B0(ws_read_addr[6]), .Z(n3962));
Q_AN02 U4508 ( .A0(n3284), .A1(n3964), .Z(n3685));
Q_OA21 U4509 ( .A0(n3965), .A1(n3966), .B0(n3956), .Z(n4488));
Q_AO21 U4510 ( .A0(n3968), .A1(n3578), .B0(n3967), .Z(n3966));
Q_OR02 U4511 ( .A0(n3969), .A1(n3608), .Z(n3967));
Q_OR02 U4512 ( .A0(n3321), .A1(n3281), .Z(n3968));
Q_OA21 U4513 ( .A0(n3970), .A1(n3971), .B0(n3572), .Z(n3965));
Q_OA21 U4514 ( .A0(n3359), .A1(n3710), .B0(ws_read_addr[6]), .Z(n3970));
Q_OA21 U4515 ( .A0(n3973), .A1(n3974), .B0(n3972), .Z(n4489));
Q_OA21 U4516 ( .A0(n3320), .A1(n3941), .B0(n3326), .Z(n3974));
Q_OR02 U4517 ( .A0(n3722), .A1(n3318), .Z(n3973));
Q_OA21 U4518 ( .A0(n3975), .A1(n3976), .B0(n3956), .Z(n4490));
Q_AN02 U4519 ( .A0(n3476), .A1(n3572), .Z(n3975));
Q_AN02 U4520 ( .A0(n3635), .A1(n3432), .Z(n3977));
Q_AN02 U4521 ( .A0(n3572), .A1(n3377), .Z(n3635));
Q_OR03 U4522 ( .A0(n3977), .A1(n3608), .A2(n3596), .Z(n3976));
Q_OA21 U4523 ( .A0(n3978), .A1(n3979), .B0(n3956), .Z(n4491));
Q_AN02 U4524 ( .A0(n3947), .A1(n3578), .Z(n3978));
Q_OR02 U4525 ( .A0(n3980), .A1(n3608), .Z(n3979));
Q_OR02 U4526 ( .A0(n3359), .A1(n3981), .Z(n3947));
Q_OA21 U4527 ( .A0(n3982), .A1(n3983), .B0(n3956), .Z(n4492));
Q_AO21 U4528 ( .A0(n3985), .A1(n3578), .B0(n3984), .Z(n3983));
Q_OA21 U4529 ( .A0(n3986), .A1(n3987), .B0(n3327), .Z(n3984));
Q_AN02 U4530 ( .A0(n3583), .A1(n3292), .Z(n3987));
Q_AN02 U4531 ( .A0(n3584), .A1(n3432), .Z(n3986));
Q_OR02 U4532 ( .A0(n3313), .A1(n3553), .Z(n3985));
Q_AN02 U4533 ( .A0(n3526), .A1(n3301), .Z(n3553));
Q_OA21 U4534 ( .A0(n3988), .A1(n3989), .B0(n3572), .Z(n3982));
Q_OA21 U4535 ( .A0(n3990), .A1(n3262), .B0(ws_read_addr[6]), .Z(n3988));
Q_AN02 U4536 ( .A0(n3678), .A1(n3327), .Z(n3990));
Q_OA21 U4537 ( .A0(n3991), .A1(n3992), .B0(n3956), .Z(n4493));
Q_AO21 U4538 ( .A0(n3994), .A1(n3578), .B0(n3993), .Z(n3992));
Q_OA21 U4539 ( .A0(n3331), .A1(n3626), .B0(n3572), .Z(n3991));
Q_AN02 U4540 ( .A0(n3350), .A1(n3387), .Z(n3331));
Q_OA21 U4541 ( .A0(n3636), .A1(n3995), .B0(n3972), .Z(n4494));
Q_AN02 U4542 ( .A0(n3857), .A1(n3361), .Z(n3995));
Q_OR02 U4543 ( .A0(n3914), .A1(n3626), .Z(n3636));
Q_OA21 U4544 ( .A0(n3997), .A1(n3998), .B0(n3996), .Z(n4495));
Q_OR02 U4545 ( .A0(n3999), .A1(n4000), .Z(n3997));
Q_OR02 U4546 ( .A0(n3514), .A1(n3745), .Z(n3998));
Q_OA21 U4547 ( .A0(n3969), .A1(n3993), .B0(n3956), .Z(n4496));
Q_AN02 U4548 ( .A0(n3350), .A1(n3614), .Z(n3993));
Q_OA21 U4549 ( .A0(n4001), .A1(n4002), .B0(n3972), .Z(n4497));
Q_OA21 U4550 ( .A0(n4003), .A1(n3329), .B0(n3326), .Z(n4002));
Q_AN02 U4551 ( .A0(n3678), .A1(ws_read_addr[3]), .Z(n4003));
Q_AO21 U4552 ( .A0(n3526), .A1(n3292), .B0(n3321), .Z(n3678));
Q_OA21 U4553 ( .A0(n4004), .A1(n4005), .B0(n3972), .Z(n4498));
Q_OA21 U4554 ( .A0(n3375), .A1(n4006), .B0(ws_read_addr[3]), .Z(n4004));
Q_OA21 U4555 ( .A0(n4007), .A1(n4008), .B0(n3996), .Z(n4500));
Q_OR02 U4556 ( .A0(n4009), .A1(n3514), .Z(n4007));
Q_AN02 U4557 ( .A0(n3395), .A1(n3226), .Z(n4010));
Q_AN03 U4558 ( .A0(n4011), .A1(n3397), .A2(n4010), .Z(n4501));
Q_OA21 U4559 ( .A0(n4012), .A1(n4013), .B0(n3972), .Z(n4502));
Q_OA21 U4560 ( .A0(n3307), .A1(n3309), .B0(n3361), .Z(n4013));
Q_INV U4561 ( .A(n3844), .Z(n3308));
Q_AO21 U4562 ( .A0(n4014), .A1(n4015), .B0(n3989), .Z(n4012));
Q_OA21 U4563 ( .A0(n4016), .A1(n3484), .B0(n3972), .Z(n4503));
Q_AN03 U4564 ( .A0(n3361), .A1(ws_read_addr[2]), .A2(n3284), .Z(n4017));
Q_OR02 U4565 ( .A0(n3914), .A1(n4017), .Z(n4016));
Q_AN02 U4566 ( .A0(n3355), .A1(n3599), .Z(n3914));
Q_OA21 U4567 ( .A0(n3626), .A1(n4018), .B0(n3972), .Z(n4504));
Q_AN03 U4568 ( .A0(n3361), .A1(n3386), .A2(n3238), .Z(n4019));
Q_OR02 U4569 ( .A0(n3484), .A1(n4019), .Z(n4018));
Q_AN03 U4570 ( .A0(n3234), .A1(n4021), .A2(n4020), .Z(n4505));
Q_OA21 U4571 ( .A0(n4001), .A1(n4022), .B0(n3972), .Z(n4506));
Q_OA21 U4572 ( .A0(n4023), .A1(n3329), .B0(n3326), .Z(n4022));
Q_AN02 U4573 ( .A0(n3717), .A1(n3292), .Z(n4023));
Q_AO21 U4574 ( .A0(n3717), .A1(n4024), .B0(n3729), .Z(n4001));
Q_AN02 U4575 ( .A0(ws_read_addr[6]), .A1(n3432), .Z(n4024));
Q_AO21 U4576 ( .A0(n3355), .A1(n3309), .B0(n4025), .Z(n3729));
Q_OA21 U4577 ( .A0(n4026), .A1(n4005), .B0(n3972), .Z(n4507));
Q_AN02 U4578 ( .A0(n3749), .A1(n3361), .Z(n4005));
Q_AO21 U4579 ( .A0(n4027), .A1(n4015), .B0(n3971), .Z(n4026));
Q_AN02 U4580 ( .A0(ws_read_addr[6]), .A1(n3386), .Z(n4015));
Q_OA21 U4581 ( .A0(n4028), .A1(n4029), .B0(n3972), .Z(n4499));
Q_AN02 U4582 ( .A0(n4030), .A1(n3361), .Z(n4029));
Q_OR02 U4583 ( .A0(n3317), .A1(n3971), .Z(n4028));
Q_OA21 U4584 ( .A0(n4031), .A1(n4008), .B0(n3996), .Z(n4508));
Q_AN02 U4585 ( .A0(n3717), .A1(ws_read_addr[4]), .Z(n4031));
Q_AN03 U4586 ( .A0(n3392), .A1(n3367), .A2(n4020), .Z(n4509));
Q_AN02 U4587 ( .A0(n3921), .A1(n3361), .Z(n4020));
Q_OA21 U4588 ( .A0(n4032), .A1(n4033), .B0(n3956), .Z(n4510));
Q_OA21 U4589 ( .A0(n4034), .A1(n3961), .B0(ws_read_addr[2]), .Z(n4033));
Q_AN02 U4590 ( .A0(n3232), .A1(n3584), .Z(n4034));
Q_INV U4591 ( .A(n3392), .Z(n3232));
Q_OA21 U4592 ( .A0(n4035), .A1(n3963), .B0(n3572), .Z(n4032));
Q_AN02 U4593 ( .A0(n3476), .A1(n3285), .Z(n3963));
Q_OA21 U4594 ( .A0(n3674), .A1(n3262), .B0(ws_read_addr[6]), .Z(n4035));
Q_AN02 U4595 ( .A0(n3526), .A1(n3378), .Z(n3262));
Q_AN02 U4596 ( .A0(n3921), .A1(n3234), .Z(n3972));
Q_OA21 U4597 ( .A0(n4036), .A1(n4037), .B0(n3972), .Z(n4511));
Q_AO21 U4598 ( .A0(n3238), .A1(n3361), .B0(n4038), .Z(n4037));
Q_AN02 U4599 ( .A0(n3342), .A1(n3327), .Z(n4038));
Q_OA21 U4600 ( .A0(n4039), .A1(n4040), .B0(n3956), .Z(n4512));
Q_AO21 U4601 ( .A0(n4041), .A1(n3386), .B0(n3596), .Z(n4040));
Q_AN02 U4602 ( .A0(n4042), .A1(n3578), .Z(n4039));
Q_AN02 U4603 ( .A0(n3921), .A1(n3545), .Z(n3996));
Q_AN02 U4604 ( .A0(n3918), .A1(n3572), .Z(n3921));
Q_OA21 U4605 ( .A0(n4043), .A1(n4042), .B0(n3996), .Z(n4513));
Q_AO21 U4606 ( .A0(n3330), .A1(n3854), .B0(n3281), .Z(n4042));
Q_OA21 U4607 ( .A0(n3623), .A1(n3980), .B0(n3956), .Z(n4514));
Q_OA21 U4608 ( .A0(n4045), .A1(n4046), .B0(n4044), .Z(n4515));
Q_AO21 U4609 ( .A0(n4048), .A1(n3578), .B0(n4047), .Z(n4046));
Q_OR02 U4610 ( .A0(n3609), .A1(n3604), .Z(n4047));
Q_AO21 U4611 ( .A0(n3330), .A1(ws_read_addr[3]), .B0(n3365), .Z(n4048));
Q_OA21 U4612 ( .A0(n4049), .A1(n3476), .B0(n3572), .Z(n4045));
Q_OR02 U4613 ( .A0(n3649), .A1(n3318), .Z(n3476));
Q_OA21 U4614 ( .A0(n3390), .A1(n3710), .B0(ws_read_addr[6]), .Z(n4049));
Q_OA21 U4615 ( .A0(n4050), .A1(n4051), .B0(n3956), .Z(n4516));
Q_AO21 U4616 ( .A0(n3390), .A1(n3960), .B0(n3639), .Z(n4051));
Q_AN02 U4617 ( .A0(n3578), .A1(ws_read_addr[2]), .Z(n3960));
Q_OR02 U4618 ( .A0(n3623), .A1(n3596), .Z(n3639));
Q_AN02 U4619 ( .A0(n3312), .A1(n3584), .Z(n3623));
Q_OA21 U4620 ( .A0(n4036), .A1(n4052), .B0(n3572), .Z(n4050));
Q_AN02 U4621 ( .A0(n3359), .A1(ws_read_addr[6]), .Z(n4036));
Q_OA21 U4622 ( .A0(n4053), .A1(n4054), .B0(n3956), .Z(n4517));
Q_AO21 U4623 ( .A0(n4030), .A1(n4041), .B0(n3980), .Z(n4054));
Q_AN02 U4624 ( .A0(n3572), .A1(n3355), .Z(n4041));
Q_OA21 U4625 ( .A0(n4053), .A1(n4055), .B0(n3956), .Z(n4518));
Q_AO21 U4626 ( .A0(n3945), .A1(n3572), .B0(n3580), .Z(n4055));
Q_OA21 U4627 ( .A0(n4056), .A1(n3674), .B0(n3578), .Z(n4053));
Q_OA21 U4628 ( .A0(n4057), .A1(n4058), .B0(n3956), .Z(n4519));
Q_AO21 U4629 ( .A0(n3584), .A1(n3761), .B0(n3580), .Z(n4059));
Q_AN02 U4630 ( .A0(n3244), .A1(n3584), .Z(n4057));
Q_OR02 U4631 ( .A0(n3596), .A1(n4059), .Z(n4058));
Q_AN02 U4632 ( .A0(n3583), .A1(n3527), .Z(n3580));
Q_AN02 U4633 ( .A0(n3918), .A1(n3226), .Z(n4044));
Q_OA21 U4634 ( .A0(n4060), .A1(n4061), .B0(n4044), .Z(n4520));
Q_AN02 U4635 ( .A0(n3403), .A1(n3572), .Z(n4060));
Q_AO21 U4636 ( .A0(n3924), .A1(n3578), .B0(n3601), .Z(n4061));
Q_OR02 U4637 ( .A0(n3961), .A1(n3608), .Z(n3601));
Q_AN02 U4638 ( .A0(n3583), .A1(n3296), .Z(n3608));
Q_AN02 U4639 ( .A0(n3583), .A1(n3395), .Z(n3604));
Q_AO21 U4640 ( .A0(n3584), .A1(n3392), .B0(n3604), .Z(n3961));
Q_AN02 U4641 ( .A0(n3924), .A1(ws_read_addr[6]), .Z(n3475));
Q_OR03 U4642 ( .A0(n3649), .A1(n3755), .A2(n3475), .Z(n3403));
Q_AN02 U4643 ( .A0(n3284), .A1(n3377), .Z(n3755));
Q_OR02 U4644 ( .A0(n3390), .A1(n3652), .Z(n3924));
Q_AN02 U4645 ( .A0(n3284), .A1(n3526), .Z(n3652));
Q_OA21 U4646 ( .A0(n4062), .A1(n4063), .B0(n3956), .Z(n4521));
Q_AN02 U4647 ( .A0(n3409), .A1(n3572), .Z(n4062));
Q_AO21 U4648 ( .A0(n3411), .A1(n3578), .B0(n3586), .Z(n4063));
Q_OR02 U4649 ( .A0(n3596), .A1(n3631), .Z(n3586));
Q_AN02 U4650 ( .A0(n3583), .A1(n3429), .Z(n3631));
Q_OR02 U4651 ( .A0(n3479), .A1(n3271), .Z(n3409));
Q_AN02 U4652 ( .A0(n3411), .A1(ws_read_addr[6]), .Z(n3479));
Q_OR02 U4653 ( .A0(n3480), .A1(n3338), .Z(n3271));
Q_AN02 U4654 ( .A0(n3312), .A1(n3377), .Z(n3338));
Q_OR02 U4655 ( .A0(n3359), .A1(n3941), .Z(n3411));
Q_OA21 U4656 ( .A0(n4064), .A1(n4065), .B0(n3956), .Z(n4522));
Q_AN02 U4657 ( .A0(n3415), .A1(n3572), .Z(n4064));
Q_AO21 U4658 ( .A0(n3276), .A1(n3584), .B0(n3598), .Z(n4065));
Q_OR02 U4659 ( .A0(n3483), .A1(n4066), .Z(n3415));
Q_OA21 U4660 ( .A0(n4067), .A1(n4068), .B0(n3956), .Z(n4523));
Q_AN02 U4661 ( .A0(n3420), .A1(n3572), .Z(n4067));
Q_OR02 U4662 ( .A0(n3274), .A1(n4066), .Z(n3420));
Q_AN02 U4663 ( .A0(n3276), .A1(n3377), .Z(n4066));
Q_AN02 U4664 ( .A0(n3918), .A1(n3234), .Z(n3956));
Q_OA21 U4665 ( .A0(n4069), .A1(n4068), .B0(n3956), .Z(n4524));
Q_AN02 U4666 ( .A0(n3422), .A1(n3578), .Z(n4069));
Q_AN02 U4667 ( .A0(n3572), .A1(n3326), .Z(n3578));
Q_OR02 U4668 ( .A0(n3980), .A1(n3598), .Z(n4068));
Q_AN02 U4669 ( .A0(n3592), .A1(n3614), .Z(n3598));
Q_AN02 U4670 ( .A0(n3583), .A1(ws_read_addr[4]), .Z(n3614));
Q_OR02 U4671 ( .A0(n3969), .A1(n3596), .Z(n3980));
Q_AN02 U4672 ( .A0(n3238), .A1(n3609), .Z(n3969));
Q_AN02 U4673 ( .A0(n3584), .A1(n3386), .Z(n3609));
Q_AN02 U4674 ( .A0(n3583), .A1(n3255), .Z(n4070));
Q_AN02 U4675 ( .A0(n4071), .A1(n3397), .Z(n3583));
Q_AO21 U4676 ( .A0(n3584), .A1(n3256), .B0(n4070), .Z(n3596));
Q_AN02 U4677 ( .A0(n3572), .A1(n3361), .Z(n3584));
Q_AN02 U4678 ( .A0(ws_read_addr[8]), .A1(n4072), .Z(n3572));
Q_OR02 U4679 ( .A0(n3505), .A1(n3981), .Z(n3422));
Q_OA21 U4680 ( .A0(n4074), .A1(n4075), .B0(n4073), .Z(n4525));
Q_OR02 U4681 ( .A0(n4076), .A1(n4077), .Z(n4075));
Q_OA21 U4682 ( .A0(n3513), .A1(n3261), .B0(n3412), .Z(n4074));
Q_AN02 U4683 ( .A0(n3534), .A1(n3327), .Z(n3261));
Q_OA21 U4684 ( .A0(n4078), .A1(n4079), .B0(ws_read_addr[7]), .Z(n4076));
Q_AN02 U4685 ( .A0(n3330), .A1(n4080), .Z(n4078));
Q_AO21 U4686 ( .A0(n3350), .A1(n3696), .B0(n4025), .Z(n4079));
Q_OA21 U4687 ( .A0(n4081), .A1(n4082), .B0(n4073), .Z(n4526));
Q_AO21 U4688 ( .A0(n3567), .A1(n3327), .B0(n4083), .Z(n4082));
Q_OR02 U4689 ( .A0(n3436), .A1(n3657), .Z(n4083));
Q_OA21 U4690 ( .A0(n4084), .A1(n4085), .B0(n3556), .Z(n4081));
Q_OA21 U4691 ( .A0(n4086), .A1(n4087), .B0(n4073), .Z(n4527));
Q_AN02 U4692 ( .A0(n3412), .A1(ws_read_addr[4]), .Z(n4088));
Q_OR03 U4693 ( .A0(n4089), .A1(n4090), .A2(n3436), .Z(n4087));
Q_OA21 U4694 ( .A0(n4091), .A1(n4092), .B0(n4088), .Z(n4089));
Q_OA21 U4695 ( .A0(n4093), .A1(n3971), .B0(ws_read_addr[7]), .Z(n4086));
Q_OA21 U4696 ( .A0(n4094), .A1(n4095), .B0(n4073), .Z(n4528));
Q_AN02 U4697 ( .A0(n3567), .A1(n3296), .Z(n4097));
Q_OR03 U4698 ( .A0(n4097), .A1(n4098), .A2(n4096), .Z(n4095));
Q_OA21 U4699 ( .A0(n4099), .A1(n3971), .B0(ws_read_addr[7]), .Z(n4094));
Q_AN02 U4700 ( .A0(n3777), .A1(n3355), .Z(n4099));
Q_OR02 U4701 ( .A0(n3312), .A1(n3392), .Z(n3777));
Q_OA21 U4702 ( .A0(n4100), .A1(n4101), .B0(n4073), .Z(n4529));
Q_OA21 U4703 ( .A0(n4102), .A1(n4103), .B0(n3412), .Z(n4100));
Q_OR02 U4704 ( .A0(n3280), .A1(n4104), .Z(n4103));
Q_OA21 U4705 ( .A0(n4105), .A1(n4106), .B0(n4073), .Z(n4530));
Q_AO21 U4706 ( .A0(n4107), .A1(n3535), .B0(n3446), .Z(n4106));
Q_AN02 U4707 ( .A0(n3412), .A1(ws_read_addr[3]), .Z(n3535));
Q_OR02 U4708 ( .A0(n3534), .A1(n3329), .Z(n4107));
Q_OA21 U4709 ( .A0(n4108), .A1(n4109), .B0(ws_read_addr[7]), .Z(n4105));
Q_AN02 U4710 ( .A0(n4110), .A1(ws_read_addr[2]), .Z(n4109));
Q_OA21 U4711 ( .A0(n4112), .A1(n4113), .B0(n4111), .Z(n4531));
Q_OA21 U4712 ( .A0(n3674), .A1(n3314), .B0(n3326), .Z(n4113));
Q_OR03 U4713 ( .A0(n4115), .A1(n3484), .A2(n4114), .Z(n4112));
Q_OA21 U4714 ( .A0(n4116), .A1(n4117), .B0(n4073), .Z(n4532));
Q_AO21 U4715 ( .A0(n3857), .A1(n3560), .B0(n3800), .Z(n4117));
Q_AN02 U4716 ( .A0(ws_read_addr[7]), .A1(n3355), .Z(n3560));
Q_AN02 U4717 ( .A0(n4118), .A1(n3412), .Z(n4116));
Q_OA21 U4718 ( .A0(n3945), .A1(n4119), .B0(n4111), .Z(n4533));
Q_AN02 U4719 ( .A0(n4118), .A1(n3326), .Z(n4119));
Q_OA21 U4720 ( .A0(n3436), .A1(n4120), .B0(n4073), .Z(n4534));
Q_AN02 U4721 ( .A0(n3312), .A1(n3417), .Z(n3436));
Q_OA21 U4722 ( .A0(n4121), .A1(n4122), .B0(n4073), .Z(n4535));
Q_OA21 U4723 ( .A0(n4108), .A1(n4123), .B0(ws_read_addr[7]), .Z(n4121));
Q_AN02 U4724 ( .A0(n3379), .A1(ws_read_addr[3]), .Z(n4123));
Q_AO21 U4725 ( .A0(n3377), .A1(n3292), .B0(n3363), .Z(n3379));
Q_AN02 U4726 ( .A0(n3355), .A1(n3432), .Z(n3363));
Q_OA21 U4727 ( .A0(n4124), .A1(n4125), .B0(n4073), .Z(n4536));
Q_OR02 U4728 ( .A0(n4126), .A1(n3800), .Z(n4125));
Q_AN02 U4729 ( .A0(n3412), .A1(ws_read_addr[2]), .Z(n3426));
Q_OA21 U4730 ( .A0(n4127), .A1(n4128), .B0(n3426), .Z(n4124));
Q_OA21 U4731 ( .A0(n3640), .A1(n3745), .B0(n3556), .Z(n4126));
Q_OA21 U4732 ( .A0(n4129), .A1(n4130), .B0(n4111), .Z(n4537));
Q_OA21 U4733 ( .A0(n3640), .A1(n4131), .B0(n3326), .Z(n4130));
Q_OA21 U4734 ( .A0(n4133), .A1(n4134), .B0(n4073), .Z(n4540));
Q_AO21 U4735 ( .A0(n4135), .A1(n4136), .B0(n3446), .Z(n4134));
Q_AN02 U4736 ( .A0(n3412), .A1(n3599), .Z(n4136));
Q_OR02 U4737 ( .A0(n4137), .A1(n4092), .Z(n4135));
Q_OA21 U4738 ( .A0(n4108), .A1(n3989), .B0(ws_read_addr[7]), .Z(n4133));
Q_OA21 U4739 ( .A0(n4138), .A1(n4139), .B0(n4111), .Z(n4541));
Q_OA21 U4740 ( .A0(n4141), .A1(n3669), .B0(n4140), .Z(n4139));
Q_AO21 U4741 ( .A0(n4142), .A1(n3506), .B0(n4114), .Z(n4138));
Q_OA21 U4742 ( .A0(n4143), .A1(n4144), .B0(n4111), .Z(n4542));
Q_OA21 U4743 ( .A0(n4145), .A1(n3669), .B0(n4140), .Z(n4144));
Q_OA21 U4744 ( .A0(n3718), .A1(n4146), .B0(ws_read_addr[4]), .Z(n4143));
Q_AN02 U4745 ( .A0(n4142), .A1(ws_read_addr[2]), .Z(n4146));
Q_AN02 U4746 ( .A0(n3355), .A1(ws_read_addr[3]), .Z(n3718));
Q_OA21 U4747 ( .A0(n3999), .A1(n4147), .B0(n4132), .Z(n4543));
Q_NR02 U4748 ( .A0(n3456), .A1(ws_read_addr[4]), .Z(n4147));
Q_AN02 U4749 ( .A0(n3238), .A1(n4043), .Z(n3999));
Q_INV U4750 ( .A(n3456), .Z(n4021));
Q_OA21 U4751 ( .A0(n4141), .A1(n4145), .B0(n4132), .Z(n4538));
Q_AN02 U4752 ( .A0(n3717), .A1(ws_read_addr[2]), .Z(n4145));
Q_INV U4753 ( .A(n4148), .Z(n4141));
Q_AN02 U4754 ( .A0(n3395), .A1(n3234), .Z(n4150));
Q_AN03 U4755 ( .A0(n3397), .A1(n4150), .A2(n4149), .Z(n4544));
Q_OA21 U4756 ( .A0(n4151), .A1(n4122), .B0(n4073), .Z(n4545));
Q_AO21 U4757 ( .A0(n4152), .A1(n4153), .B0(n3446), .Z(n4122));
Q_AN02 U4758 ( .A0(n3412), .A1(n3432), .Z(n4153));
Q_AO21 U4759 ( .A0(n3417), .A1(n3309), .B0(n4090), .Z(n3446));
Q_AN02 U4760 ( .A0(n3392), .A1(ws_read_addr[2]), .Z(n3309));
Q_INV U4761 ( .A(n3805), .Z(n4152));
Q_OA21 U4762 ( .A0(n4108), .A1(n4154), .B0(ws_read_addr[7]), .Z(n4151));
Q_AN02 U4763 ( .A0(n4142), .A1(n3292), .Z(n4154));
Q_AN02 U4764 ( .A0(ws_read_addr[4]), .A1(n3285), .Z(n3292));
Q_AO21 U4765 ( .A0(n3355), .A1(n3327), .B0(n3679), .Z(n4142));
Q_OA21 U4766 ( .A0(n3321), .A1(n3912), .B0(ws_read_addr[6]), .Z(n4108));
Q_AN02 U4767 ( .A0(ws_read_addr[5]), .A1(n3432), .Z(n3321));
Q_OA21 U4768 ( .A0(n4155), .A1(n4156), .B0(n4073), .Z(n4546));
Q_AO21 U4769 ( .A0(n3688), .A1(n3556), .B0(n3800), .Z(n4156));
Q_OA21 U4770 ( .A0(n4009), .A1(n4157), .B0(n3412), .Z(n4155));
Q_OR02 U4771 ( .A0(n3640), .A1(n3365), .Z(n3688));
Q_AN02 U4772 ( .A0(n3526), .A1(n3296), .Z(n3365));
Q_OA21 U4773 ( .A0(n3387), .A1(n4158), .B0(n4111), .Z(n4547));
Q_NR02 U4774 ( .A0(ws_read_addr[6]), .A1(ws_read_addr[4]), .Z(n4140));
Q_OA21 U4775 ( .A0(n4159), .A1(n4027), .B0(n4140), .Z(n4158));
Q_AN02 U4776 ( .A0(n3238), .A1(ws_read_addr[5]), .Z(n4159));
Q_AN02 U4777 ( .A0(n4011), .A1(n3545), .Z(n4132));
Q_OA21 U4778 ( .A0(n4160), .A1(n4161), .B0(n4132), .Z(n4548));
Q_INV U4779 ( .A(n4162), .Z(n4163));
Q_OR02 U4780 ( .A0(n4163), .A1(n4157), .Z(n4161));
Q_AN02 U4781 ( .A0(n4027), .A1(n3386), .Z(n4157));
Q_AN02 U4782 ( .A0(n4030), .A1(ws_read_addr[5]), .Z(n4160));
Q_AN02 U4783 ( .A0(n4073), .A1(n4120), .Z(n4539));
Q_OR02 U4784 ( .A0(n4098), .A1(n3800), .Z(n4120));
Q_OA21 U4785 ( .A0(n4164), .A1(n4165), .B0(n4073), .Z(n4549));
Q_AN02 U4786 ( .A0(n4166), .A1(ws_read_addr[2]), .Z(n4077));
Q_AO21 U4787 ( .A0(n4167), .A1(n3539), .B0(n4077), .Z(n4165));
Q_AN02 U4788 ( .A0(n3567), .A1(n3285), .Z(n3539));
Q_OA21 U4789 ( .A0(n4168), .A1(n4169), .B0(ws_read_addr[7]), .Z(n4164));
Q_AN02 U4790 ( .A0(n3453), .A1(n4080), .Z(n4168));
Q_AN02 U4791 ( .A0(ws_read_addr[6]), .A1(ws_read_addr[2]), .Z(n4080));
Q_OR02 U4792 ( .A0(n4115), .A1(n4025), .Z(n4169));
Q_AN02 U4793 ( .A0(n3377), .A1(n3351), .Z(n4025));
Q_AN02 U4794 ( .A0(n3284), .A1(n3375), .Z(n4115));
Q_AN02 U4795 ( .A0(n3355), .A1(ws_read_addr[2]), .Z(n3375));
Q_OA21 U4796 ( .A0(n4170), .A1(n4171), .B0(n4073), .Z(n4550));
Q_AN02 U4797 ( .A0(n3567), .A1(n3599), .Z(n4172));
Q_OR03 U4798 ( .A0(n4172), .A1(n4173), .A2(n3657), .Z(n4171));
Q_AN02 U4799 ( .A0(n3417), .A1(n3854), .Z(n4173));
Q_OA21 U4800 ( .A0(n4114), .A1(n4174), .B0(ws_read_addr[7]), .Z(n4170));
Q_AN02 U4801 ( .A0(n3385), .A1(ws_read_addr[4]), .Z(n4174));
Q_AN03 U4802 ( .A0(n3397), .A1(n3386), .A2(n3238), .Z(n4114));
Q_OR02 U4803 ( .A0(n3239), .A1(n3679), .Z(n3385));
Q_AN02 U4804 ( .A0(n3377), .A1(ws_read_addr[3]), .Z(n3679));
Q_AN02 U4805 ( .A0(n3238), .A1(n3355), .Z(n3239));
Q_OA21 U4806 ( .A0(n4175), .A1(n4176), .B0(n4073), .Z(n4551));
Q_AN02 U4807 ( .A0(n3543), .A1(n3556), .Z(n4175));
Q_AN02 U4808 ( .A0(ws_read_addr[7]), .A1(ws_read_addr[6]), .Z(n3556));
Q_AO21 U4809 ( .A0(n3284), .A1(n3567), .B0(n4177), .Z(n4176));
Q_OR02 U4810 ( .A0(n4098), .A1(n3657), .Z(n4177));
Q_OA21 U4811 ( .A0(n4178), .A1(n4179), .B0(n4073), .Z(n4552));
Q_OA21 U4812 ( .A0(n4180), .A1(n4181), .B0(ws_read_addr[5]), .Z(n4179));
Q_AN02 U4813 ( .A0(n3464), .A1(n3351), .Z(n4181));
Q_AN02 U4814 ( .A0(n4072), .A1(ws_read_addr[6]), .Z(n3464));
Q_AN02 U4815 ( .A0(n3284), .A1(n3412), .Z(n4180));
Q_OA21 U4816 ( .A0(n4182), .A1(n3971), .B0(ws_read_addr[7]), .Z(n4178));
Q_OA21 U4817 ( .A0(n3791), .A1(n4183), .B0(n4073), .Z(n4553));
Q_AN02 U4818 ( .A0(n3567), .A1(n3392), .Z(n3791));
Q_AO21 U4819 ( .A0(n4184), .A1(n3417), .B0(n4096), .Z(n4183));
Q_OA21 U4820 ( .A0(n4186), .A1(n4187), .B0(n4185), .Z(n4554));
Q_OR02 U4821 ( .A0(n3472), .A1(n4166), .Z(n4187));
Q_AN02 U4822 ( .A0(n3453), .A1(n3412), .Z(n3472));
Q_OA21 U4823 ( .A0(n4188), .A1(n4110), .B0(ws_read_addr[7]), .Z(n4186));
Q_AN02 U4824 ( .A0(n3377), .A1(n3296), .Z(n3318));
Q_AO21 U4825 ( .A0(n3342), .A1(ws_read_addr[3]), .B0(n3318), .Z(n4110));
Q_OA21 U4826 ( .A0(n4189), .A1(n4190), .B0(n4073), .Z(n4555));
Q_OR02 U4827 ( .A0(n3435), .A1(n4191), .Z(n4190));
Q_AN02 U4828 ( .A0(n3622), .A1(n3412), .Z(n3435));
Q_OA21 U4829 ( .A0(n4192), .A1(n3626), .B0(ws_read_addr[7]), .Z(n4189));
Q_AN02 U4830 ( .A0(n4011), .A1(n3234), .Z(n4111));
Q_AN02 U4831 ( .A0(n3918), .A1(n4071), .Z(n4011));
Q_AN02 U4832 ( .A0(n3697), .A1(ws_read_addr[7]), .Z(n4071));
Q_OA21 U4833 ( .A0(n4193), .A1(n4194), .B0(n4111), .Z(n4556));
Q_OA21 U4834 ( .A0(n4056), .A1(n4008), .B0(n3326), .Z(n4194));
Q_AN02 U4835 ( .A0(n4030), .A1(n3526), .Z(n4008));
Q_OR02 U4836 ( .A0(n4093), .A1(n3484), .Z(n4193));
Q_OA21 U4837 ( .A0(n4195), .A1(n4196), .B0(n4073), .Z(n4557));
Q_OR02 U4838 ( .A0(n3445), .A1(n4096), .Z(n4196));
Q_AN02 U4839 ( .A0(n3312), .A1(n3567), .Z(n3445));
Q_AN02 U4840 ( .A0(ws_read_addr[7]), .A1(n3377), .Z(n3567));
Q_OA21 U4841 ( .A0(n4197), .A1(n3484), .B0(ws_read_addr[7]), .Z(n4195));
Q_OR02 U4842 ( .A0(n4182), .A1(n3626), .Z(n4197));
Q_OA21 U4843 ( .A0(n3465), .A1(n4198), .B0(n4073), .Z(n4558));
Q_AN02 U4844 ( .A0(n3505), .A1(n3412), .Z(n3465));
Q_AO21 U4845 ( .A0(n4030), .A1(n3417), .B0(n4096), .Z(n4198));
Q_AN02 U4846 ( .A0(n4199), .A1(n3226), .Z(n4185));
Q_AN03 U4847 ( .A0(ws_read_addr[2]), .A1(n4201), .A2(n4200), .Z(n3226));
Q_OA21 U4848 ( .A0(n4202), .A1(n4203), .B0(n4185), .Z(n4559));
Q_AN02 U4849 ( .A0(n3576), .A1(ws_read_addr[7]), .Z(n4202));
Q_AO21 U4850 ( .A0(n3330), .A1(n3412), .B0(n4166), .Z(n4203));
Q_OR02 U4851 ( .A0(n3801), .A1(n3800), .Z(n4166));
Q_AN02 U4852 ( .A0(n3428), .A1(n3395), .Z(n3800));
Q_OR02 U4853 ( .A0(n4188), .A1(n3342), .Z(n3576));
Q_AN02 U4854 ( .A0(n3330), .A1(ws_read_addr[6]), .Z(n4188));
Q_OR02 U4855 ( .A0(n3696), .A1(n4006), .Z(n3342));
Q_OA21 U4856 ( .A0(n4204), .A1(n4205), .B0(n4073), .Z(n4560));
Q_OR02 U4857 ( .A0(n3656), .A1(n4191), .Z(n4205));
Q_AN02 U4858 ( .A0(n4084), .A1(n3412), .Z(n3656));
Q_OR02 U4859 ( .A0(n4098), .A1(n4090), .Z(n4191));
Q_AN02 U4860 ( .A0(n3238), .A1(n3801), .Z(n4098));
Q_AN02 U4861 ( .A0(n3417), .A1(n3386), .Z(n3801));
Q_OA21 U4862 ( .A0(n4192), .A1(n4052), .B0(ws_read_addr[7]), .Z(n4204));
Q_AN02 U4863 ( .A0(n4084), .A1(ws_read_addr[6]), .Z(n4192));
Q_OR02 U4864 ( .A0(n3317), .A1(n3484), .Z(n4052));
Q_OR02 U4865 ( .A0(n3640), .A1(n3281), .Z(n4084));
Q_OA21 U4866 ( .A0(n4206), .A1(n4207), .B0(n4073), .Z(n4561));
Q_AO21 U4867 ( .A0(n3543), .A1(n3412), .B0(n4096), .Z(n4207));
Q_OA21 U4868 ( .A0(n4093), .A1(n3945), .B0(ws_read_addr[7]), .Z(n4206));
Q_AN02 U4869 ( .A0(n3543), .A1(ws_read_addr[6]), .Z(n4093));
Q_OA21 U4870 ( .A0(n4208), .A1(n4101), .B0(n4073), .Z(n4562));
Q_OA21 U4871 ( .A0(n3245), .A1(n3945), .B0(ws_read_addr[7]), .Z(n4208));
Q_OR02 U4872 ( .A0(n3480), .A1(n3484), .Z(n3945));
Q_AN02 U4873 ( .A0(n3238), .A1(n4006), .Z(n3484));
Q_AN02 U4874 ( .A0(n3377), .A1(ws_read_addr[4]), .Z(n4006));
Q_AN02 U4875 ( .A0(n4199), .A1(n3234), .Z(n4073));
Q_AN02 U4876 ( .A0(n3918), .A1(n3697), .Z(n4199));
Q_OA21 U4877 ( .A0(n4209), .A1(n4101), .B0(n4073), .Z(n4563));
Q_AN02 U4878 ( .A0(ws_read_addr[7]), .A1(n3326), .Z(n3412));
Q_OR02 U4879 ( .A0(n3953), .A1(n4096), .Z(n4101));
Q_AN02 U4880 ( .A0(n3244), .A1(n3417), .Z(n3953));
Q_OR02 U4881 ( .A0(n3657), .A1(n4090), .Z(n4096));
Q_AN02 U4882 ( .A0(n3428), .A1(n3351), .Z(n4090));
Q_AN02 U4883 ( .A0(n3428), .A1(n3255), .Z(n4210));
Q_AN02 U4884 ( .A0(n4072), .A1(n3397), .Z(n3428));
Q_AN02 U4885 ( .A0(ws_read_addr[6]), .A1(ws_read_addr[5]), .Z(n3397));
Q_AO21 U4886 ( .A0(n3417), .A1(n3256), .B0(n4210), .Z(n3657));
Q_AN02 U4887 ( .A0(ws_read_addr[7]), .A1(n3361), .Z(n3417));
Q_OA21 U4888 ( .A0(n4211), .A1(n3543), .B0(n3412), .Z(n4209));
Q_AN02 U4889 ( .A0(n3244), .A1(ws_read_addr[5]), .Z(n4211));
Q_OR02 U4890 ( .A0(n3359), .A1(n3281), .Z(n3543));
Q_OA21 U4891 ( .A0(n4213), .A1(n4214), .B0(n4212), .Z(n4564));
Q_AN03 U4892 ( .A0(n3326), .A1(ws_read_addr[2]), .A2(n4162), .Z(n4214));
Q_OR02 U4893 ( .A0(n3393), .A1(n4215), .Z(n4162));
Q_NR02 U4894 ( .A0(n3395), .A1(ws_read_addr[5]), .Z(n4215));
Q_OA21 U4895 ( .A0(n4216), .A1(n4217), .B0(n4212), .Z(n4565));
Q_OA21 U4896 ( .A0(n4218), .A1(n3669), .B0(n3326), .Z(n4217));
Q_AN02 U4897 ( .A0(n3238), .A1(n3526), .Z(n3669));
Q_OA21 U4898 ( .A0(n4219), .A1(n4220), .B0(n4212), .Z(n4566));
Q_OA21 U4899 ( .A0(n4221), .A1(n4222), .B0(n3326), .Z(n4220));
Q_OA21 U4900 ( .A0(n4223), .A1(n4224), .B0(n4212), .Z(n4567));
Q_OA21 U4901 ( .A0(n3519), .A1(n4225), .B0(n3326), .Z(n4224));
Q_OA21 U4902 ( .A0(n3312), .A1(n3305), .B0(n3526), .Z(n4225));
Q_OA21 U4903 ( .A0(n4227), .A1(n4228), .B0(n4226), .Z(n4568));
Q_NR02 U4904 ( .A0(n3255), .A1(ws_read_addr[5]), .Z(n4228));
Q_NR02 U4905 ( .A0(n3854), .A1(ws_read_addr[4]), .Z(n3305));
Q_INV U4906 ( .A(n3854), .Z(n3592));
Q_OA21 U4907 ( .A0(n4213), .A1(n4229), .B0(n4212), .Z(n4569));
Q_OA21 U4908 ( .A0(n4230), .A1(n3313), .B0(ws_read_addr[6]), .Z(n4213));
Q_OR02 U4909 ( .A0(n4009), .A1(n4231), .Z(n4230));
Q_AN02 U4910 ( .A0(n3390), .A1(n3285), .Z(n3313));
Q_OA21 U4911 ( .A0(n4216), .A1(n4232), .B0(n4212), .Z(n4570));
Q_OA21 U4912 ( .A0(n4218), .A1(n4233), .B0(n3326), .Z(n4232));
Q_OA21 U4913 ( .A0(n3506), .A1(n4234), .B0(ws_read_addr[5]), .Z(n4218));
Q_OA21 U4914 ( .A0(n4056), .A1(n4235), .B0(ws_read_addr[6]), .Z(n4216));
Q_OR02 U4915 ( .A0(n3514), .A1(n3710), .Z(n4235));
Q_OA21 U4916 ( .A0(n4219), .A1(n4236), .B0(n4212), .Z(n4571));
Q_OA21 U4917 ( .A0(n4221), .A1(n3281), .B0(n3326), .Z(n4236));
Q_OR02 U4918 ( .A0(n3519), .A1(n3359), .Z(n4221));
Q_OA21 U4919 ( .A0(n3390), .A1(n4085), .B0(ws_read_addr[6]), .Z(n4219));
Q_AN02 U4920 ( .A0(n3526), .A1(n3392), .Z(n4085));
Q_OA21 U4921 ( .A0(n4223), .A1(n4237), .B0(n4212), .Z(n4572));
Q_AN02 U4922 ( .A0(n4167), .A1(n3355), .Z(n4223));
Q_OA21 U4923 ( .A0(n3519), .A1(n4238), .B0(n3326), .Z(n4237));
Q_AN02 U4924 ( .A0(ws_read_addr[5]), .A1(n3506), .Z(n3519));
Q_OA21 U4925 ( .A0(n4227), .A1(n4239), .B0(n4226), .Z(n4573));
Q_OR02 U4926 ( .A0(n4056), .A1(n3505), .Z(n4227));
Q_AN02 U4927 ( .A0(n4212), .A1(n4240), .Z(n4574));
Q_MX02 U4928 ( .S(ws_read_addr[6]), .A0(n4241), .A1(n4242), .Z(n4240));
Q_OR03 U4929 ( .A0(n3513), .A1(n4243), .A2(n3675), .Z(n4241));
Q_AN02 U4930 ( .A0(n3284), .A1(n4137), .Z(n3513));
Q_AN02 U4931 ( .A0(ws_read_addr[5]), .A1(n3285), .Z(n4137));
Q_OR03 U4932 ( .A0(n4244), .A1(n3912), .A2(n3329), .Z(n4242));
Q_AN02 U4933 ( .A0(n3844), .A1(n4091), .Z(n4244));
Q_AN02 U4934 ( .A0(n4212), .A1(n4245), .Z(n4575));
Q_MX02 U4935 ( .S(ws_read_addr[6]), .A0(n4246), .A1(n3994), .Z(n4245));
Q_OR03 U4936 ( .A0(n3920), .A1(n3710), .A2(n3674), .Z(n4246));
Q_AN02 U4937 ( .A0(n3350), .A1(n4043), .Z(n3920));
Q_AN02 U4938 ( .A0(ws_read_addr[5]), .A1(ws_read_addr[4]), .Z(n4043));
Q_OR02 U4939 ( .A0(n4000), .A1(n3745), .Z(n3994));
Q_AN02 U4940 ( .A0(n3284), .A1(n4092), .Z(n3745));
Q_AN02 U4941 ( .A0(n3526), .A1(ws_read_addr[2]), .Z(n4092));
Q_AN02 U4942 ( .A0(n3350), .A1(n3651), .Z(n4000));
Q_OA21 U4943 ( .A0(n4129), .A1(n4247), .B0(n4212), .Z(n4576));
Q_AN02 U4944 ( .A0(n3857), .A1(n3355), .Z(n4129));
Q_OA21 U4945 ( .A0(n4118), .A1(n4248), .B0(n3326), .Z(n4247));
Q_AN02 U4946 ( .A0(n3526), .A1(n3256), .Z(n4248));
Q_OR02 U4947 ( .A0(n3395), .A1(n3563), .Z(n3857));
Q_OA21 U4948 ( .A0(n3317), .A1(n4249), .B0(n4212), .Z(n4577));
Q_OA21 U4949 ( .A0(n4250), .A1(n3674), .B0(n3326), .Z(n4249));
Q_AN02 U4950 ( .A0(n3733), .A1(ws_read_addr[5]), .Z(n4250));
Q_OR02 U4951 ( .A0(n3821), .A1(n3599), .Z(n3733));
Q_AN02 U4952 ( .A0(n3350), .A1(ws_read_addr[4]), .Z(n3821));
Q_INV U4953 ( .A(n3238), .Z(n3350));
Q_AN03 U4954 ( .A0(n4251), .A1(n3234), .A2(n3356), .Z(n4578));
Q_OR02 U4955 ( .A0(n3761), .A1(n4252), .Z(n3356));
Q_NR02 U4956 ( .A0(n3343), .A1(ws_read_addr[4]), .Z(n4252));
Q_OA21 U4957 ( .A0(n4253), .A1(n4254), .B0(n4212), .Z(n4579));
Q_AN02 U4958 ( .A0(n3551), .A1(ws_read_addr[3]), .Z(n3615));
Q_AO21 U4959 ( .A0(n4148), .A1(n4255), .B0(n3615), .Z(n4253));
Q_AN02 U4960 ( .A0(ws_read_addr[6]), .A1(n3506), .Z(n4255));
Q_OR02 U4961 ( .A0(n3499), .A1(n3989), .Z(n3551));
Q_AN02 U4962 ( .A0(n3377), .A1(n3506), .Z(n3989));
Q_AN02 U4963 ( .A0(n3355), .A1(n3564), .Z(n3499));
Q_OA21 U4964 ( .A0(n4256), .A1(n4257), .B0(n4212), .Z(n4580));
Q_AN02 U4965 ( .A0(ws_read_addr[6]), .A1(ws_read_addr[3]), .Z(n4258));
Q_OA21 U4966 ( .A0(n4259), .A1(n3558), .B0(n4258), .Z(n4256));
Q_AN02 U4967 ( .A0(n3330), .A1(ws_read_addr[2]), .Z(n4259));
Q_OR02 U4968 ( .A0(n3651), .A1(n3855), .Z(n3330));
Q_OA21 U4969 ( .A0(n3626), .A1(n4260), .B0(n4212), .Z(n4582));
Q_AN02 U4970 ( .A0(n3649), .A1(ws_read_addr[2]), .Z(n3626));
Q_AN03 U4971 ( .A0(n4252), .A1(n3234), .A2(n4251), .Z(n4583));
Q_AN02 U4972 ( .A0(n4212), .A1(n4261), .Z(n4584));
Q_MX02 U4973 ( .S(ws_read_addr[6]), .A0(n4262), .A1(n4263), .Z(n4261));
Q_AO21 U4974 ( .A0(n3844), .A1(n3805), .B0(n3525), .Z(n4262));
Q_OR02 U4975 ( .A0(n3506), .A1(n3564), .Z(n3844));
Q_AN02 U4976 ( .A0(n3526), .A1(n3432), .Z(n3329));
Q_AN02 U4977 ( .A0(n3386), .A1(ws_read_addr[2]), .Z(n3432));
Q_AO21 U4978 ( .A0(n4014), .A1(ws_read_addr[4]), .B0(n3329), .Z(n4263));
Q_MX02 U4979 ( .S(ws_read_addr[5]), .A0(n3337), .A1(n3343), .Z(n4014));
Q_OA21 U4980 ( .A0(n4264), .A1(n4265), .B0(n4212), .Z(n4585));
Q_AN02 U4981 ( .A0(n3749), .A1(n3355), .Z(n4264));
Q_OA21 U4982 ( .A0(n3674), .A1(n4266), .B0(n3326), .Z(n4265));
Q_OR02 U4983 ( .A0(n3395), .A1(n4234), .Z(n3749));
Q_AN03 U4984 ( .A0(n4149), .A1(n4268), .A2(n4267), .Z(n4586));
Q_AN02 U4985 ( .A0(n3526), .A1(n3234), .Z(n4268));
Q_MX02 U4986 ( .S(ws_read_addr[6]), .A0(n4269), .A1(n4030), .Z(n4267));
Q_OR02 U4987 ( .A0(n3563), .A1(n4234), .Z(n4030));
Q_OA21 U4988 ( .A0(n4118), .A1(n4233), .B0(n4226), .Z(n4587));
Q_OA21 U4989 ( .A0(n4270), .A1(n4254), .B0(n4212), .Z(n4588));
Q_OA21 U4990 ( .A0(n3525), .A1(n3675), .B0(n3326), .Z(n4254));
Q_AN02 U4991 ( .A0(n3735), .A1(n3526), .Z(n3675));
Q_AN02 U4992 ( .A0(n3534), .A1(ws_read_addr[3]), .Z(n3525));
Q_OR02 U4993 ( .A0(n3527), .A1(n3378), .Z(n3735));
Q_AN02 U4994 ( .A0(n3599), .A1(n3285), .Z(n3378));
Q_AN02 U4995 ( .A0(n3296), .A1(ws_read_addr[2]), .Z(n3527));
Q_AN02 U4996 ( .A0(n3526), .A1(n3506), .Z(n4104));
Q_AO21 U4997 ( .A0(ws_read_addr[5]), .A1(n3564), .B0(n4104), .Z(n3534));
Q_OA21 U4998 ( .A0(n4271), .A1(n4266), .B0(ws_read_addr[6]), .Z(n4270));
Q_AN02 U4999 ( .A0(n4148), .A1(n3506), .Z(n4271));
Q_AN02 U5000 ( .A0(ws_read_addr[4]), .A1(ws_read_addr[2]), .Z(n3506));
Q_OR02 U5001 ( .A0(n3717), .A1(n3805), .Z(n4148));
Q_OR02 U5002 ( .A0(n4091), .A1(n4128), .Z(n3717));
Q_AN02 U5003 ( .A0(n3526), .A1(ws_read_addr[3]), .Z(n4128));
Q_AN02 U5004 ( .A0(ws_read_addr[5]), .A1(n3327), .Z(n4091));
Q_OA21 U5005 ( .A0(n4272), .A1(n4257), .B0(n4212), .Z(n4589));
Q_OA21 U5006 ( .A0(n4102), .A1(n4222), .B0(n3326), .Z(n4257));
Q_OA21 U5007 ( .A0(n3761), .A1(n3256), .B0(n3526), .Z(n4222));
Q_OA21 U5008 ( .A0(n4273), .A1(n3710), .B0(ws_read_addr[6]), .Z(n4272));
Q_AN02 U5009 ( .A0(n3526), .A1(n3599), .Z(n3710));
Q_AN02 U5010 ( .A0(n4027), .A1(ws_read_addr[4]), .Z(n4273));
Q_OR02 U5011 ( .A0(n3570), .A1(n4131), .Z(n4027));
Q_AN02 U5012 ( .A0(n3526), .A1(n3854), .Z(n4131));
Q_AN02 U5013 ( .A0(ws_read_addr[5]), .A1(n3456), .Z(n3570));
Q_NR02 U5014 ( .A0(ws_read_addr[3]), .A1(ws_read_addr[2]), .Z(n3456));
Q_OA21 U5015 ( .A0(n4274), .A1(n4275), .B0(n4212), .Z(n4581));
Q_AN02 U5016 ( .A0(n4276), .A1(n3326), .Z(n4275));
Q_AN02 U5017 ( .A0(n3881), .A1(n3355), .Z(n4274));
Q_OR02 U5018 ( .A0(n3761), .A1(n3599), .Z(n3881));
Q_OA21 U5019 ( .A0(n3689), .A1(n4260), .B0(n4212), .Z(n4590));
Q_OA21 U5020 ( .A0(n4118), .A1(n3281), .B0(n3326), .Z(n4260));
Q_OR02 U5021 ( .A0(n4102), .A1(n3674), .Z(n4118));
Q_AN02 U5022 ( .A0(ws_read_addr[5]), .A1(n3599), .Z(n4102));
Q_AN03 U5023 ( .A0(n3367), .A1(n4167), .A2(n4251), .Z(n4591));
Q_AN02 U5024 ( .A0(n4277), .A1(n4200), .Z(n3367));
Q_NR02 U5025 ( .A0(ws_read_addr[2]), .A1(ws_read_addr[1]), .Z(n4277));
Q_AN02 U5026 ( .A0(n4149), .A1(n3361), .Z(n4251));
Q_OA21 U5027 ( .A0(n4278), .A1(n4279), .B0(n4212), .Z(n4592));
Q_OA21 U5028 ( .A0(n4280), .A1(n4231), .B0(ws_read_addr[6]), .Z(n4278));
Q_AN02 U5029 ( .A0(n4167), .A1(n3964), .Z(n4231));
Q_NR02 U5030 ( .A0(ws_read_addr[5]), .A1(ws_read_addr[2]), .Z(n3964));
Q_INV U5031 ( .A(n3395), .Z(n4167));
Q_OR02 U5032 ( .A0(n4009), .A1(n3912), .Z(n4280));
Q_AN02 U5033 ( .A0(n3526), .A1(n3351), .Z(n3912));
Q_AN02 U5034 ( .A0(n3395), .A1(n3285), .Z(n3351));
Q_AN02 U5035 ( .A0(n4212), .A1(n4281), .Z(n4593));
Q_MX02 U5036 ( .S(ws_read_addr[6]), .A0(n4282), .A1(n4283), .Z(n4281));
Q_OR02 U5037 ( .A0(n3640), .A1(n4233), .Z(n4282));
Q_AN02 U5038 ( .A0(n4269), .A1(n3526), .Z(n4233));
Q_OR02 U5039 ( .A0(n3761), .A1(n3564), .Z(n4269));
Q_OR02 U5040 ( .A0(n4056), .A1(n3805), .Z(n4283));
Q_NR02 U5041 ( .A0(ws_read_addr[5]), .A1(ws_read_addr[3]), .Z(n3805));
Q_OA21 U5042 ( .A0(n3387), .A1(n4284), .B0(n4212), .Z(n4594));
Q_AN02 U5043 ( .A0(n3355), .A1(ws_read_addr[4]), .Z(n3387));
Q_OA21 U5044 ( .A0(n4285), .A1(n4238), .B0(n3326), .Z(n4284));
Q_AN02 U5045 ( .A0(n4184), .A1(ws_read_addr[5]), .Z(n4285));
Q_OA21 U5046 ( .A0(n3312), .A1(n3564), .B0(n3526), .Z(n4238));
Q_OA21 U5047 ( .A0(n3696), .A1(n4286), .B0(n4212), .Z(n4595));
Q_AN02 U5048 ( .A0(n4184), .A1(n3377), .Z(n4286));
Q_OR02 U5049 ( .A0(n3854), .A1(n4234), .Z(n4184));
Q_AN02 U5050 ( .A0(ws_read_addr[3]), .A1(ws_read_addr[2]), .Z(n3854));
Q_OA21 U5051 ( .A0(n3359), .A1(n4239), .B0(n4226), .Z(n4596));
Q_OA21 U5052 ( .A0(n4287), .A1(n4279), .B0(n4212), .Z(n4597));
Q_OA21 U5053 ( .A0(n4288), .A1(n4289), .B0(n3326), .Z(n4279));
Q_AN02 U5054 ( .A0(n3453), .A1(ws_read_addr[2]), .Z(n4288));
Q_OR02 U5055 ( .A0(n3651), .A1(n3514), .Z(n3453));
Q_OA21 U5056 ( .A0(n4290), .A1(n4291), .B0(ws_read_addr[2]), .Z(n4287));
Q_OR02 U5057 ( .A0(n3696), .A1(n3971), .Z(n4291));
Q_OA21 U5058 ( .A0(n4127), .A1(n3855), .B0(ws_read_addr[6]), .Z(n4290));
Q_AN02 U5059 ( .A0(n4212), .A1(n4292), .Z(n4598));
Q_MX02 U5060 ( .S(ws_read_addr[6]), .A0(n4293), .A1(n4294), .Z(n4292));
Q_OR03 U5061 ( .A0(n4009), .A1(n3941), .A2(n3359), .Z(n4293));
Q_OR02 U5062 ( .A0(n3441), .A1(n3314), .Z(n4294));
Q_AN02 U5063 ( .A0(n3238), .A1(n3558), .Z(n3314));
Q_NR02 U5064 ( .A0(ws_read_addr[5]), .A1(ws_read_addr[4]), .Z(n3558));
Q_OR02 U5065 ( .A0(n4056), .A1(n3281), .Z(n3441));
Q_OA21 U5066 ( .A0(n4295), .A1(n4296), .B0(n4212), .Z(n4599));
Q_OA21 U5067 ( .A0(n4009), .A1(n3981), .B0(n3326), .Z(n4296));
Q_AN02 U5068 ( .A0(n3276), .A1(n3526), .Z(n3981));
Q_AO21 U5069 ( .A0(n4276), .A1(ws_read_addr[6]), .B0(n3480), .Z(n4295));
Q_OR02 U5070 ( .A0(n3674), .A1(n3281), .Z(n4276));
Q_AN02 U5071 ( .A0(n3238), .A1(n3855), .Z(n3281));
Q_AN02 U5072 ( .A0(n3526), .A1(ws_read_addr[4]), .Z(n3855));
Q_AN02 U5073 ( .A0(n3390), .A1(ws_read_addr[2]), .Z(n3674));
Q_OA21 U5074 ( .A0(n3245), .A1(n4297), .B0(n4212), .Z(n4600));
Q_OA21 U5075 ( .A0(n4009), .A1(n4266), .B0(n3326), .Z(n4298));
Q_AN03 U5076 ( .A0(ws_read_addr[5]), .A1(ws_read_addr[2]), .A2(n3284), .Z(n4009));
Q_OR02 U5077 ( .A0(n3480), .A1(n4298), .Z(n4297));
Q_AN02 U5078 ( .A0(n3244), .A1(n3355), .Z(n3245));
Q_OR02 U5079 ( .A0(n3312), .A1(n4234), .Z(n3244));
Q_AN02 U5080 ( .A0(n3238), .A1(n3386), .Z(n4234));
Q_OA21 U5081 ( .A0(n3505), .A1(n4239), .B0(n4226), .Z(n4601));
Q_OA21 U5082 ( .A0(n4299), .A1(n4229), .B0(n4212), .Z(n4602));
Q_OA21 U5083 ( .A0(n4300), .A1(n4289), .B0(n3326), .Z(n4229));
Q_AN02 U5084 ( .A0(n3393), .A1(ws_read_addr[2]), .Z(n4300));
Q_OA21 U5085 ( .A0(n3563), .A1(n3256), .B0(n3526), .Z(n4289));
Q_AN02 U5086 ( .A0(n3284), .A1(ws_read_addr[2]), .Z(n3563));
Q_OA21 U5087 ( .A0(n4301), .A1(n4302), .B0(ws_read_addr[2]), .Z(n4299));
Q_AN02 U5088 ( .A0(n3393), .A1(ws_read_addr[6]), .Z(n4301));
Q_OR02 U5089 ( .A0(n3722), .A1(n3649), .Z(n4302));
Q_AN02 U5090 ( .A0(n3284), .A1(n3355), .Z(n3722));
Q_OR02 U5091 ( .A0(n3689), .A1(n3971), .Z(n3649));
Q_AN02 U5092 ( .A0(n3377), .A1(n3395), .Z(n3971));
Q_AN02 U5093 ( .A0(n3355), .A1(n3392), .Z(n3689));
Q_OR02 U5094 ( .A0(n4127), .A1(n3390), .Z(n3393));
Q_AN02 U5095 ( .A0(n3284), .A1(ws_read_addr[5]), .Z(n4127));
Q_OR02 U5096 ( .A0(n3280), .A1(n3514), .Z(n3390));
Q_AN02 U5097 ( .A0(n3526), .A1(n3395), .Z(n3514));
Q_AN02 U5098 ( .A0(ws_read_addr[5]), .A1(n3392), .Z(n3280));
Q_OR02 U5099 ( .A0(n3296), .A1(n3599), .Z(n3284));
Q_OA21 U5100 ( .A0(n4303), .A1(n4304), .B0(n4212), .Z(n4603));
Q_OA21 U5101 ( .A0(n3622), .A1(n3941), .B0(n3326), .Z(n4304));
Q_AN02 U5102 ( .A0(n3312), .A1(n3526), .Z(n3941));
Q_AO21 U5103 ( .A0(n3622), .A1(ws_read_addr[6]), .B0(n4305), .Z(n4303));
Q_OR02 U5104 ( .A0(n4182), .A1(n3480), .Z(n4305));
Q_AN02 U5105 ( .A0(n3312), .A1(n3355), .Z(n4182));
Q_OR02 U5106 ( .A0(n4056), .A1(n3359), .Z(n3622));
Q_AN02 U5107 ( .A0(n3312), .A1(ws_read_addr[5]), .Z(n4056));
Q_OA21 U5108 ( .A0(n4306), .A1(n4307), .B0(n4212), .Z(n4604));
Q_OA21 U5109 ( .A0(n3505), .A1(n4266), .B0(n3326), .Z(n4307));
Q_AN02 U5110 ( .A0(n3526), .A1(n3564), .Z(n4266));
Q_AO21 U5111 ( .A0(n3505), .A1(ws_read_addr[6]), .B0(n3274), .Z(n4306));
Q_AN02 U5112 ( .A0(n4149), .A1(n3234), .Z(n4212));
Q_OA21 U5113 ( .A0(n4308), .A1(n4309), .B0(n4212), .Z(n4605));
Q_AN02 U5114 ( .A0(n4310), .A1(n3361), .Z(n4309));
Q_NR02 U5115 ( .A0(ws_read_addr[6]), .A1(ws_read_addr[5]), .Z(n3361));
Q_OR02 U5116 ( .A0(n3483), .A1(n3274), .Z(n4308));
Q_AN02 U5117 ( .A0(n3276), .A1(n3355), .Z(n3483));
Q_OR02 U5118 ( .A0(n3317), .A1(n3480), .Z(n3274));
Q_AN02 U5119 ( .A0(n3238), .A1(n3696), .Z(n3317));
Q_AN02 U5120 ( .A0(n3355), .A1(n3386), .Z(n3696));
Q_AN02 U5121 ( .A0(n3377), .A1(n3255), .Z(n4311));
Q_AN02 U5122 ( .A0(n3326), .A1(ws_read_addr[5]), .Z(n3377));
Q_AO21 U5123 ( .A0(n3355), .A1(n3256), .B0(n4311), .Z(n3480));
Q_AN02 U5124 ( .A0(ws_read_addr[6]), .A1(n3526), .Z(n3355));
Q_AN02 U5125 ( .A0(n4149), .A1(n3545), .Z(n4226));
Q_NR02 U5126 ( .A0(ws_read_addr[1]), .A1(ws_read_addr[0]), .Z(n3234));
Q_INV U5127 ( .A(ws_read_addr[0]), .Z(n4200));
Q_INV U5128 ( .A(ws_read_addr[1]), .Z(n4201));
Q_INV U5129 ( .A(ws_read_addr[6]), .Z(n3326));
Q_AN02 U5130 ( .A0(n3918), .A1(n3398), .Z(n4149));
Q_NR02 U5131 ( .A0(ws_read_addr[8]), .A1(ws_read_addr[7]), .Z(n3398));
Q_INV U5132 ( .A(ws_read_addr[7]), .Z(n4072));
Q_INV U5133 ( .A(ws_read_addr[8]), .Z(n3697));
Q_NR02 U5134 ( .A0(ws_read_addr[10]), .A1(ws_read_addr[9]), .Z(n3918));
Q_INV U5135 ( .A(ws_read_addr[9]), .Z(n3399));
Q_INV U5136 ( .A(ws_read_addr[10]), .Z(n3698));
Q_OA21 U5137 ( .A0(n4312), .A1(n4239), .B0(n4226), .Z(n4606));
Q_AN02 U5138 ( .A0(n4310), .A1(n3526), .Z(n4239));
Q_OR02 U5139 ( .A0(n3276), .A1(n3564), .Z(n4310));
Q_NR02 U5140 ( .A0(ws_read_addr[4]), .A1(ws_read_addr[2]), .Z(n3564));
Q_OR02 U5141 ( .A0(n3279), .A1(n3505), .Z(n4312));
Q_AN02 U5142 ( .A0(n3276), .A1(ws_read_addr[5]), .Z(n3279));
Q_OR02 U5143 ( .A0(n3640), .A1(n3359), .Z(n3505));
Q_AN02 U5144 ( .A0(n3238), .A1(n3651), .Z(n3640));
Q_AN02 U5145 ( .A0(ws_read_addr[5]), .A1(n3386), .Z(n3651));
Q_AN02 U5146 ( .A0(n3526), .A1(n3255), .Z(n4243));
Q_AN02 U5147 ( .A0(n3395), .A1(ws_read_addr[2]), .Z(n3255));
Q_AN02 U5148 ( .A0(ws_read_addr[4]), .A1(ws_read_addr[3]), .Z(n3395));
Q_INV U5149 ( .A(ws_read_addr[5]), .Z(n3526));
Q_AO21 U5150 ( .A0(ws_read_addr[5]), .A1(n3256), .B0(n4243), .Z(n3359));
Q_AN02 U5151 ( .A0(n3392), .A1(n3285), .Z(n3256));
Q_NR02 U5152 ( .A0(ws_read_addr[4]), .A1(ws_read_addr[3]), .Z(n3392));
Q_OR02 U5153 ( .A0(n3761), .A1(n3312), .Z(n3276));
Q_OR02 U5154 ( .A0(n3429), .A1(n3301), .Z(n3312));
Q_AN02 U5155 ( .A0(n3599), .A1(ws_read_addr[2]), .Z(n3301));
Q_AN02 U5156 ( .A0(n3386), .A1(ws_read_addr[3]), .Z(n3599));
Q_INV U5157 ( .A(ws_read_addr[4]), .Z(n3386));
Q_AN02 U5158 ( .A0(n3296), .A1(n3285), .Z(n3429));
Q_AN02 U5159 ( .A0(ws_read_addr[4]), .A1(n3327), .Z(n3296));
Q_OR02 U5160 ( .A0(n3337), .A1(n3343), .Z(n3238));
Q_AN02 U5161 ( .A0(n3327), .A1(ws_read_addr[2]), .Z(n3343));
Q_INV U5162 ( .A(ws_read_addr[3]), .Z(n3327));
Q_AN02 U5163 ( .A0(ws_read_addr[3]), .A1(n3285), .Z(n3337));
Q_INV U5164 ( .A(ws_read_addr[2]), .Z(n3285));
Q_INV U5165 ( .A(i_rd_strb), .Z(n4607));
Q_AN03 U5166 ( .A0(w_do_read), .A1(n450), .A2(n4607), .Z(n4608));
Q_AN03 U5167 ( .A0(w_do_write), .A1(w_32b_aligned), .A2(w_valid_rd_addr), .Z(n4609));
Q_AN03 U5168 ( .A0(w_do_read), .A1(w_32b_aligned), .A2(w_valid_rd_addr), .Z(n4610));
Q_AN02 U5169 ( .A0(n446), .A1(r32_mux_8_data[0]), .Z(n4611));
Q_AN02 U5170 ( .A0(n446), .A1(r32_mux_8_data[1]), .Z(n4612));
Q_AN02 U5171 ( .A0(n446), .A1(r32_mux_8_data[2]), .Z(n4613));
Q_AN02 U5172 ( .A0(n446), .A1(r32_mux_8_data[3]), .Z(n4614));
Q_AN02 U5173 ( .A0(n446), .A1(r32_mux_8_data[4]), .Z(n4615));
Q_AN02 U5174 ( .A0(n446), .A1(r32_mux_8_data[5]), .Z(n4616));
Q_AN02 U5175 ( .A0(n446), .A1(r32_mux_8_data[6]), .Z(n4617));
Q_AN02 U5176 ( .A0(n446), .A1(r32_mux_8_data[7]), .Z(n4618));
Q_AN02 U5177 ( .A0(n446), .A1(r32_mux_8_data[8]), .Z(n4619));
Q_AN02 U5178 ( .A0(n446), .A1(r32_mux_8_data[9]), .Z(n4620));
Q_AN02 U5179 ( .A0(n446), .A1(r32_mux_8_data[10]), .Z(n4621));
Q_AN02 U5180 ( .A0(n446), .A1(r32_mux_8_data[11]), .Z(n4622));
Q_AN02 U5181 ( .A0(n446), .A1(r32_mux_8_data[12]), .Z(n4623));
Q_AN02 U5182 ( .A0(n446), .A1(r32_mux_8_data[13]), .Z(n4624));
Q_AN02 U5183 ( .A0(n446), .A1(r32_mux_8_data[14]), .Z(n4625));
Q_AN02 U5184 ( .A0(n446), .A1(r32_mux_8_data[15]), .Z(n4626));
Q_AN02 U5185 ( .A0(n446), .A1(r32_mux_8_data[16]), .Z(n4627));
Q_AN02 U5186 ( .A0(n446), .A1(r32_mux_8_data[17]), .Z(n4628));
Q_AN02 U5187 ( .A0(n446), .A1(r32_mux_8_data[18]), .Z(n4629));
Q_AN02 U5188 ( .A0(n446), .A1(r32_mux_8_data[19]), .Z(n4630));
Q_AN02 U5189 ( .A0(n446), .A1(r32_mux_8_data[20]), .Z(n4631));
Q_AN02 U5190 ( .A0(n446), .A1(r32_mux_8_data[21]), .Z(n4632));
Q_AN02 U5191 ( .A0(n446), .A1(r32_mux_8_data[22]), .Z(n4633));
Q_AN02 U5192 ( .A0(n446), .A1(r32_mux_8_data[23]), .Z(n4634));
Q_AN02 U5193 ( .A0(n446), .A1(r32_mux_8_data[24]), .Z(n4635));
Q_AN02 U5194 ( .A0(n446), .A1(r32_mux_8_data[25]), .Z(n4636));
Q_AN02 U5195 ( .A0(n446), .A1(r32_mux_8_data[26]), .Z(n4637));
Q_AN02 U5196 ( .A0(n446), .A1(r32_mux_8_data[27]), .Z(n4638));
Q_AN02 U5197 ( .A0(n446), .A1(r32_mux_8_data[28]), .Z(n4639));
Q_AN02 U5198 ( .A0(n446), .A1(r32_mux_8_data[29]), .Z(n4640));
Q_AN02 U5199 ( .A0(n446), .A1(r32_mux_8_data[30]), .Z(n4641));
Q_AN02 U5200 ( .A0(n446), .A1(r32_mux_8_data[31]), .Z(n4642));
Q_AN02 U5201 ( .A0(n446), .A1(r32_mux_7_data[0]), .Z(n4643));
Q_AN02 U5202 ( .A0(n446), .A1(r32_mux_7_data[1]), .Z(n4644));
Q_AN02 U5203 ( .A0(n446), .A1(r32_mux_7_data[2]), .Z(n4645));
Q_AN02 U5204 ( .A0(n446), .A1(r32_mux_7_data[3]), .Z(n4646));
Q_AN02 U5205 ( .A0(n446), .A1(r32_mux_7_data[4]), .Z(n4647));
Q_AN02 U5206 ( .A0(n446), .A1(r32_mux_7_data[5]), .Z(n4648));
Q_AN02 U5207 ( .A0(n446), .A1(r32_mux_7_data[6]), .Z(n4649));
Q_AN02 U5208 ( .A0(n446), .A1(r32_mux_7_data[7]), .Z(n4650));
Q_AN02 U5209 ( .A0(n446), .A1(r32_mux_7_data[8]), .Z(n4651));
Q_AN02 U5210 ( .A0(n446), .A1(r32_mux_7_data[9]), .Z(n4652));
Q_AN02 U5211 ( .A0(n446), .A1(r32_mux_7_data[10]), .Z(n4653));
Q_AN02 U5212 ( .A0(n446), .A1(r32_mux_7_data[11]), .Z(n4654));
Q_AN02 U5213 ( .A0(n446), .A1(r32_mux_7_data[12]), .Z(n4655));
Q_AN02 U5214 ( .A0(n446), .A1(r32_mux_7_data[13]), .Z(n4656));
Q_AN02 U5215 ( .A0(n446), .A1(r32_mux_7_data[14]), .Z(n4657));
Q_AN02 U5216 ( .A0(n446), .A1(r32_mux_7_data[15]), .Z(n4658));
Q_AN02 U5217 ( .A0(n446), .A1(r32_mux_7_data[16]), .Z(n4659));
Q_AN02 U5218 ( .A0(n446), .A1(r32_mux_7_data[17]), .Z(n4660));
Q_AN02 U5219 ( .A0(n446), .A1(r32_mux_7_data[18]), .Z(n4661));
Q_AN02 U5220 ( .A0(n446), .A1(r32_mux_7_data[19]), .Z(n4662));
Q_AN02 U5221 ( .A0(n446), .A1(r32_mux_7_data[20]), .Z(n4663));
Q_AN02 U5222 ( .A0(n446), .A1(r32_mux_7_data[21]), .Z(n4664));
Q_AN02 U5223 ( .A0(n446), .A1(r32_mux_7_data[22]), .Z(n4665));
Q_AN02 U5224 ( .A0(n446), .A1(r32_mux_7_data[23]), .Z(n4666));
Q_AN02 U5225 ( .A0(n446), .A1(r32_mux_7_data[24]), .Z(n4667));
Q_AN02 U5226 ( .A0(n446), .A1(r32_mux_7_data[25]), .Z(n4668));
Q_AN02 U5227 ( .A0(n446), .A1(r32_mux_7_data[26]), .Z(n4669));
Q_AN02 U5228 ( .A0(n446), .A1(r32_mux_7_data[27]), .Z(n4670));
Q_AN02 U5229 ( .A0(n446), .A1(r32_mux_7_data[28]), .Z(n4671));
Q_AN02 U5230 ( .A0(n446), .A1(r32_mux_7_data[29]), .Z(n4672));
Q_AN02 U5231 ( .A0(n446), .A1(r32_mux_7_data[30]), .Z(n4673));
Q_AN02 U5232 ( .A0(n446), .A1(r32_mux_7_data[31]), .Z(n4674));
Q_AN02 U5233 ( .A0(n446), .A1(r32_mux_6_data[0]), .Z(n4675));
Q_AN02 U5234 ( .A0(n446), .A1(r32_mux_6_data[1]), .Z(n4676));
Q_AN02 U5235 ( .A0(n446), .A1(r32_mux_6_data[2]), .Z(n4677));
Q_AN02 U5236 ( .A0(n446), .A1(r32_mux_6_data[3]), .Z(n4678));
Q_AN02 U5237 ( .A0(n446), .A1(r32_mux_6_data[4]), .Z(n4679));
Q_AN02 U5238 ( .A0(n446), .A1(r32_mux_6_data[5]), .Z(n4680));
Q_AN02 U5239 ( .A0(n446), .A1(r32_mux_6_data[6]), .Z(n4681));
Q_AN02 U5240 ( .A0(n446), .A1(r32_mux_6_data[7]), .Z(n4682));
Q_AN02 U5241 ( .A0(n446), .A1(r32_mux_6_data[8]), .Z(n4683));
Q_AN02 U5242 ( .A0(n446), .A1(r32_mux_6_data[9]), .Z(n4684));
Q_AN02 U5243 ( .A0(n446), .A1(r32_mux_6_data[10]), .Z(n4685));
Q_AN02 U5244 ( .A0(n446), .A1(r32_mux_6_data[11]), .Z(n4686));
Q_AN02 U5245 ( .A0(n446), .A1(r32_mux_6_data[12]), .Z(n4687));
Q_AN02 U5246 ( .A0(n446), .A1(r32_mux_6_data[13]), .Z(n4688));
Q_AN02 U5247 ( .A0(n446), .A1(r32_mux_6_data[14]), .Z(n4689));
Q_AN02 U5248 ( .A0(n446), .A1(r32_mux_6_data[15]), .Z(n4690));
Q_AN02 U5249 ( .A0(n446), .A1(r32_mux_6_data[16]), .Z(n4691));
Q_AN02 U5250 ( .A0(n446), .A1(r32_mux_6_data[17]), .Z(n4692));
Q_AN02 U5251 ( .A0(n446), .A1(r32_mux_6_data[18]), .Z(n4693));
Q_AN02 U5252 ( .A0(n446), .A1(r32_mux_6_data[19]), .Z(n4694));
Q_AN02 U5253 ( .A0(n446), .A1(r32_mux_6_data[20]), .Z(n4695));
Q_AN02 U5254 ( .A0(n446), .A1(r32_mux_6_data[21]), .Z(n4696));
Q_AN02 U5255 ( .A0(n446), .A1(r32_mux_6_data[22]), .Z(n4697));
Q_AN02 U5256 ( .A0(n446), .A1(r32_mux_6_data[23]), .Z(n4698));
Q_AN02 U5257 ( .A0(n446), .A1(r32_mux_6_data[24]), .Z(n4699));
Q_AN02 U5258 ( .A0(n446), .A1(r32_mux_6_data[25]), .Z(n4700));
Q_AN02 U5259 ( .A0(n446), .A1(r32_mux_6_data[26]), .Z(n4701));
Q_AN02 U5260 ( .A0(n446), .A1(r32_mux_6_data[27]), .Z(n4702));
Q_AN02 U5261 ( .A0(n446), .A1(r32_mux_6_data[28]), .Z(n4703));
Q_AN02 U5262 ( .A0(n446), .A1(r32_mux_6_data[29]), .Z(n4704));
Q_AN02 U5263 ( .A0(n446), .A1(r32_mux_6_data[30]), .Z(n4705));
Q_AN02 U5264 ( .A0(n446), .A1(r32_mux_6_data[31]), .Z(n4706));
Q_AN02 U5265 ( .A0(n446), .A1(r32_mux_5_data[0]), .Z(n4707));
Q_AN02 U5266 ( .A0(n446), .A1(r32_mux_5_data[1]), .Z(n4708));
Q_AN02 U5267 ( .A0(n446), .A1(r32_mux_5_data[2]), .Z(n4709));
Q_AN02 U5268 ( .A0(n446), .A1(r32_mux_5_data[3]), .Z(n4710));
Q_AN02 U5269 ( .A0(n446), .A1(r32_mux_5_data[4]), .Z(n4711));
Q_AN02 U5270 ( .A0(n446), .A1(r32_mux_5_data[5]), .Z(n4712));
Q_AN02 U5271 ( .A0(n446), .A1(r32_mux_5_data[6]), .Z(n4713));
Q_AN02 U5272 ( .A0(n446), .A1(r32_mux_5_data[7]), .Z(n4714));
Q_AN02 U5273 ( .A0(n446), .A1(r32_mux_5_data[8]), .Z(n4715));
Q_AN02 U5274 ( .A0(n446), .A1(r32_mux_5_data[9]), .Z(n4716));
Q_AN02 U5275 ( .A0(n446), .A1(r32_mux_5_data[10]), .Z(n4717));
Q_AN02 U5276 ( .A0(n446), .A1(r32_mux_5_data[11]), .Z(n4718));
Q_AN02 U5277 ( .A0(n446), .A1(r32_mux_5_data[12]), .Z(n4719));
Q_AN02 U5278 ( .A0(n446), .A1(r32_mux_5_data[13]), .Z(n4720));
Q_AN02 U5279 ( .A0(n446), .A1(r32_mux_5_data[14]), .Z(n4721));
Q_AN02 U5280 ( .A0(n446), .A1(r32_mux_5_data[15]), .Z(n4722));
Q_AN02 U5281 ( .A0(n446), .A1(r32_mux_5_data[16]), .Z(n4723));
Q_AN02 U5282 ( .A0(n446), .A1(r32_mux_5_data[17]), .Z(n4724));
Q_AN02 U5283 ( .A0(n446), .A1(r32_mux_5_data[18]), .Z(n4725));
Q_AN02 U5284 ( .A0(n446), .A1(r32_mux_5_data[19]), .Z(n4726));
Q_AN02 U5285 ( .A0(n446), .A1(r32_mux_5_data[20]), .Z(n4727));
Q_AN02 U5286 ( .A0(n446), .A1(r32_mux_5_data[21]), .Z(n4728));
Q_AN02 U5287 ( .A0(n446), .A1(r32_mux_5_data[22]), .Z(n4729));
Q_AN02 U5288 ( .A0(n446), .A1(r32_mux_5_data[23]), .Z(n4730));
Q_AN02 U5289 ( .A0(n446), .A1(r32_mux_5_data[24]), .Z(n4731));
Q_AN02 U5290 ( .A0(n446), .A1(r32_mux_5_data[25]), .Z(n4732));
Q_AN02 U5291 ( .A0(n446), .A1(r32_mux_5_data[26]), .Z(n4733));
Q_AN02 U5292 ( .A0(n446), .A1(r32_mux_5_data[27]), .Z(n4734));
Q_AN02 U5293 ( .A0(n446), .A1(r32_mux_5_data[28]), .Z(n4735));
Q_AN02 U5294 ( .A0(n446), .A1(r32_mux_5_data[29]), .Z(n4736));
Q_AN02 U5295 ( .A0(n446), .A1(r32_mux_5_data[30]), .Z(n4737));
Q_AN02 U5296 ( .A0(n446), .A1(r32_mux_5_data[31]), .Z(n4738));
Q_AN02 U5297 ( .A0(n446), .A1(r32_mux_4_data[0]), .Z(n4739));
Q_AN02 U5298 ( .A0(n446), .A1(r32_mux_4_data[1]), .Z(n4740));
Q_AN02 U5299 ( .A0(n446), .A1(r32_mux_4_data[2]), .Z(n4741));
Q_AN02 U5300 ( .A0(n446), .A1(r32_mux_4_data[3]), .Z(n4742));
Q_AN02 U5301 ( .A0(n446), .A1(r32_mux_4_data[4]), .Z(n4743));
Q_AN02 U5302 ( .A0(n446), .A1(r32_mux_4_data[5]), .Z(n4744));
Q_AN02 U5303 ( .A0(n446), .A1(r32_mux_4_data[6]), .Z(n4745));
Q_AN02 U5304 ( .A0(n446), .A1(r32_mux_4_data[7]), .Z(n4746));
Q_AN02 U5305 ( .A0(n446), .A1(r32_mux_4_data[8]), .Z(n4747));
Q_AN02 U5306 ( .A0(n446), .A1(r32_mux_4_data[9]), .Z(n4748));
Q_AN02 U5307 ( .A0(n446), .A1(r32_mux_4_data[10]), .Z(n4749));
Q_AN02 U5308 ( .A0(n446), .A1(r32_mux_4_data[11]), .Z(n4750));
Q_AN02 U5309 ( .A0(n446), .A1(r32_mux_4_data[12]), .Z(n4751));
Q_AN02 U5310 ( .A0(n446), .A1(r32_mux_4_data[13]), .Z(n4752));
Q_AN02 U5311 ( .A0(n446), .A1(r32_mux_4_data[14]), .Z(n4753));
Q_AN02 U5312 ( .A0(n446), .A1(r32_mux_4_data[15]), .Z(n4754));
Q_AN02 U5313 ( .A0(n446), .A1(r32_mux_4_data[16]), .Z(n4755));
Q_AN02 U5314 ( .A0(n446), .A1(r32_mux_4_data[17]), .Z(n4756));
Q_AN02 U5315 ( .A0(n446), .A1(r32_mux_4_data[18]), .Z(n4757));
Q_AN02 U5316 ( .A0(n446), .A1(r32_mux_4_data[19]), .Z(n4758));
Q_AN02 U5317 ( .A0(n446), .A1(r32_mux_4_data[20]), .Z(n4759));
Q_AN02 U5318 ( .A0(n446), .A1(r32_mux_4_data[21]), .Z(n4760));
Q_AN02 U5319 ( .A0(n446), .A1(r32_mux_4_data[22]), .Z(n4761));
Q_AN02 U5320 ( .A0(n446), .A1(r32_mux_4_data[23]), .Z(n4762));
Q_AN02 U5321 ( .A0(n446), .A1(r32_mux_4_data[24]), .Z(n4763));
Q_AN02 U5322 ( .A0(n446), .A1(r32_mux_4_data[25]), .Z(n4764));
Q_AN02 U5323 ( .A0(n446), .A1(r32_mux_4_data[26]), .Z(n4765));
Q_AN02 U5324 ( .A0(n446), .A1(r32_mux_4_data[27]), .Z(n4766));
Q_AN02 U5325 ( .A0(n446), .A1(r32_mux_4_data[28]), .Z(n4767));
Q_AN02 U5326 ( .A0(n446), .A1(r32_mux_4_data[29]), .Z(n4768));
Q_AN02 U5327 ( .A0(n446), .A1(r32_mux_4_data[30]), .Z(n4769));
Q_AN02 U5328 ( .A0(n446), .A1(r32_mux_4_data[31]), .Z(n4770));
Q_AN02 U5329 ( .A0(n446), .A1(r32_mux_3_data[0]), .Z(n4771));
Q_AN02 U5330 ( .A0(n446), .A1(r32_mux_3_data[1]), .Z(n4772));
Q_AN02 U5331 ( .A0(n446), .A1(r32_mux_3_data[2]), .Z(n4773));
Q_AN02 U5332 ( .A0(n446), .A1(r32_mux_3_data[3]), .Z(n4774));
Q_AN02 U5333 ( .A0(n446), .A1(r32_mux_3_data[4]), .Z(n4775));
Q_AN02 U5334 ( .A0(n446), .A1(r32_mux_3_data[5]), .Z(n4776));
Q_AN02 U5335 ( .A0(n446), .A1(r32_mux_3_data[6]), .Z(n4777));
Q_AN02 U5336 ( .A0(n446), .A1(r32_mux_3_data[7]), .Z(n4778));
Q_AN02 U5337 ( .A0(n446), .A1(r32_mux_3_data[8]), .Z(n4779));
Q_AN02 U5338 ( .A0(n446), .A1(r32_mux_3_data[9]), .Z(n4780));
Q_AN02 U5339 ( .A0(n446), .A1(r32_mux_3_data[10]), .Z(n4781));
Q_AN02 U5340 ( .A0(n446), .A1(r32_mux_3_data[11]), .Z(n4782));
Q_AN02 U5341 ( .A0(n446), .A1(r32_mux_3_data[12]), .Z(n4783));
Q_AN02 U5342 ( .A0(n446), .A1(r32_mux_3_data[13]), .Z(n4784));
Q_AN02 U5343 ( .A0(n446), .A1(r32_mux_3_data[14]), .Z(n4785));
Q_AN02 U5344 ( .A0(n446), .A1(r32_mux_3_data[15]), .Z(n4786));
Q_AN02 U5345 ( .A0(n446), .A1(r32_mux_3_data[16]), .Z(n4787));
Q_AN02 U5346 ( .A0(n446), .A1(r32_mux_3_data[17]), .Z(n4788));
Q_AN02 U5347 ( .A0(n446), .A1(r32_mux_3_data[18]), .Z(n4789));
Q_AN02 U5348 ( .A0(n446), .A1(r32_mux_3_data[19]), .Z(n4790));
Q_AN02 U5349 ( .A0(n446), .A1(r32_mux_3_data[20]), .Z(n4791));
Q_AN02 U5350 ( .A0(n446), .A1(r32_mux_3_data[21]), .Z(n4792));
Q_AN02 U5351 ( .A0(n446), .A1(r32_mux_3_data[22]), .Z(n4793));
Q_AN02 U5352 ( .A0(n446), .A1(r32_mux_3_data[23]), .Z(n4794));
Q_AN02 U5353 ( .A0(n446), .A1(r32_mux_3_data[24]), .Z(n4795));
Q_AN02 U5354 ( .A0(n446), .A1(r32_mux_3_data[25]), .Z(n4796));
Q_AN02 U5355 ( .A0(n446), .A1(r32_mux_3_data[26]), .Z(n4797));
Q_AN02 U5356 ( .A0(n446), .A1(r32_mux_3_data[27]), .Z(n4798));
Q_AN02 U5357 ( .A0(n446), .A1(r32_mux_3_data[28]), .Z(n4799));
Q_AN02 U5358 ( .A0(n446), .A1(r32_mux_3_data[29]), .Z(n4800));
Q_AN02 U5359 ( .A0(n446), .A1(r32_mux_3_data[30]), .Z(n4801));
Q_AN02 U5360 ( .A0(n446), .A1(r32_mux_3_data[31]), .Z(n4802));
Q_AN02 U5361 ( .A0(n446), .A1(r32_mux_2_data[0]), .Z(n4803));
Q_AN02 U5362 ( .A0(n446), .A1(r32_mux_2_data[1]), .Z(n4804));
Q_AN02 U5363 ( .A0(n446), .A1(r32_mux_2_data[2]), .Z(n4805));
Q_AN02 U5364 ( .A0(n446), .A1(r32_mux_2_data[3]), .Z(n4806));
Q_AN02 U5365 ( .A0(n446), .A1(r32_mux_2_data[4]), .Z(n4807));
Q_AN02 U5366 ( .A0(n446), .A1(r32_mux_2_data[5]), .Z(n4808));
Q_AN02 U5367 ( .A0(n446), .A1(r32_mux_2_data[6]), .Z(n4809));
Q_AN02 U5368 ( .A0(n446), .A1(r32_mux_2_data[7]), .Z(n4810));
Q_AN02 U5369 ( .A0(n446), .A1(r32_mux_2_data[8]), .Z(n4811));
Q_AN02 U5370 ( .A0(n446), .A1(r32_mux_2_data[9]), .Z(n4812));
Q_AN02 U5371 ( .A0(n446), .A1(r32_mux_2_data[10]), .Z(n4813));
Q_AN02 U5372 ( .A0(n446), .A1(r32_mux_2_data[11]), .Z(n4814));
Q_AN02 U5373 ( .A0(n446), .A1(r32_mux_2_data[12]), .Z(n4815));
Q_AN02 U5374 ( .A0(n446), .A1(r32_mux_2_data[13]), .Z(n4816));
Q_AN02 U5375 ( .A0(n446), .A1(r32_mux_2_data[14]), .Z(n4817));
Q_AN02 U5376 ( .A0(n446), .A1(r32_mux_2_data[15]), .Z(n4818));
Q_AN02 U5377 ( .A0(n446), .A1(r32_mux_2_data[16]), .Z(n4819));
Q_AN02 U5378 ( .A0(n446), .A1(r32_mux_2_data[17]), .Z(n4820));
Q_AN02 U5379 ( .A0(n446), .A1(r32_mux_2_data[18]), .Z(n4821));
Q_AN02 U5380 ( .A0(n446), .A1(r32_mux_2_data[19]), .Z(n4822));
Q_AN02 U5381 ( .A0(n446), .A1(r32_mux_2_data[20]), .Z(n4823));
Q_AN02 U5382 ( .A0(n446), .A1(r32_mux_2_data[21]), .Z(n4824));
Q_AN02 U5383 ( .A0(n446), .A1(r32_mux_2_data[22]), .Z(n4825));
Q_AN02 U5384 ( .A0(n446), .A1(r32_mux_2_data[23]), .Z(n4826));
Q_AN02 U5385 ( .A0(n446), .A1(r32_mux_2_data[24]), .Z(n4827));
Q_AN02 U5386 ( .A0(n446), .A1(r32_mux_2_data[25]), .Z(n4828));
Q_AN02 U5387 ( .A0(n446), .A1(r32_mux_2_data[26]), .Z(n4829));
Q_AN02 U5388 ( .A0(n446), .A1(r32_mux_2_data[27]), .Z(n4830));
Q_AN02 U5389 ( .A0(n446), .A1(r32_mux_2_data[28]), .Z(n4831));
Q_AN02 U5390 ( .A0(n446), .A1(r32_mux_2_data[29]), .Z(n4832));
Q_AN02 U5391 ( .A0(n446), .A1(r32_mux_2_data[30]), .Z(n4833));
Q_AN02 U5392 ( .A0(n446), .A1(r32_mux_2_data[31]), .Z(n4834));
Q_AN02 U5393 ( .A0(n446), .A1(r32_mux_1_data[0]), .Z(n4835));
Q_AN02 U5394 ( .A0(n446), .A1(r32_mux_1_data[1]), .Z(n4836));
Q_AN02 U5395 ( .A0(n446), .A1(r32_mux_1_data[2]), .Z(n4837));
Q_AN02 U5396 ( .A0(n446), .A1(r32_mux_1_data[3]), .Z(n4838));
Q_AN02 U5397 ( .A0(n446), .A1(r32_mux_1_data[4]), .Z(n4839));
Q_AN02 U5398 ( .A0(n446), .A1(r32_mux_1_data[5]), .Z(n4840));
Q_AN02 U5399 ( .A0(n446), .A1(r32_mux_1_data[6]), .Z(n4841));
Q_AN02 U5400 ( .A0(n446), .A1(r32_mux_1_data[7]), .Z(n4842));
Q_AN02 U5401 ( .A0(n446), .A1(r32_mux_1_data[8]), .Z(n4843));
Q_AN02 U5402 ( .A0(n446), .A1(r32_mux_1_data[9]), .Z(n4844));
Q_AN02 U5403 ( .A0(n446), .A1(r32_mux_1_data[10]), .Z(n4845));
Q_AN02 U5404 ( .A0(n446), .A1(r32_mux_1_data[11]), .Z(n4846));
Q_AN02 U5405 ( .A0(n446), .A1(r32_mux_1_data[12]), .Z(n4847));
Q_AN02 U5406 ( .A0(n446), .A1(r32_mux_1_data[13]), .Z(n4848));
Q_AN02 U5407 ( .A0(n446), .A1(r32_mux_1_data[14]), .Z(n4849));
Q_AN02 U5408 ( .A0(n446), .A1(r32_mux_1_data[15]), .Z(n4850));
Q_AN02 U5409 ( .A0(n446), .A1(r32_mux_1_data[16]), .Z(n4851));
Q_AN02 U5410 ( .A0(n446), .A1(r32_mux_1_data[17]), .Z(n4852));
Q_AN02 U5411 ( .A0(n446), .A1(r32_mux_1_data[18]), .Z(n4853));
Q_AN02 U5412 ( .A0(n446), .A1(r32_mux_1_data[19]), .Z(n4854));
Q_AN02 U5413 ( .A0(n446), .A1(r32_mux_1_data[20]), .Z(n4855));
Q_AN02 U5414 ( .A0(n446), .A1(r32_mux_1_data[21]), .Z(n4856));
Q_AN02 U5415 ( .A0(n446), .A1(r32_mux_1_data[22]), .Z(n4857));
Q_AN02 U5416 ( .A0(n446), .A1(r32_mux_1_data[23]), .Z(n4858));
Q_AN02 U5417 ( .A0(n446), .A1(r32_mux_1_data[24]), .Z(n4859));
Q_AN02 U5418 ( .A0(n446), .A1(r32_mux_1_data[25]), .Z(n4860));
Q_AN02 U5419 ( .A0(n446), .A1(r32_mux_1_data[26]), .Z(n4861));
Q_AN02 U5420 ( .A0(n446), .A1(r32_mux_1_data[27]), .Z(n4862));
Q_AN02 U5421 ( .A0(n446), .A1(r32_mux_1_data[28]), .Z(n4863));
Q_AN02 U5422 ( .A0(n446), .A1(r32_mux_1_data[29]), .Z(n4864));
Q_AN02 U5423 ( .A0(n446), .A1(r32_mux_1_data[30]), .Z(n4865));
Q_AN02 U5424 ( .A0(n446), .A1(r32_mux_1_data[31]), .Z(n4866));
Q_AN02 U5425 ( .A0(n446), .A1(r32_mux_0_data[0]), .Z(n4867));
Q_AN02 U5426 ( .A0(n446), .A1(r32_mux_0_data[1]), .Z(n4868));
Q_AN02 U5427 ( .A0(n446), .A1(r32_mux_0_data[2]), .Z(n4869));
Q_AN02 U5428 ( .A0(n446), .A1(r32_mux_0_data[3]), .Z(n4870));
Q_AN02 U5429 ( .A0(n446), .A1(r32_mux_0_data[4]), .Z(n4871));
Q_AN02 U5430 ( .A0(n446), .A1(r32_mux_0_data[5]), .Z(n4872));
Q_AN02 U5431 ( .A0(n446), .A1(r32_mux_0_data[6]), .Z(n4873));
Q_AN02 U5432 ( .A0(n446), .A1(r32_mux_0_data[7]), .Z(n4874));
Q_AN02 U5433 ( .A0(n446), .A1(r32_mux_0_data[8]), .Z(n4875));
Q_AN02 U5434 ( .A0(n446), .A1(r32_mux_0_data[9]), .Z(n4876));
Q_AN02 U5435 ( .A0(n446), .A1(r32_mux_0_data[10]), .Z(n4877));
Q_AN02 U5436 ( .A0(n446), .A1(r32_mux_0_data[11]), .Z(n4878));
Q_AN02 U5437 ( .A0(n446), .A1(r32_mux_0_data[12]), .Z(n4879));
Q_AN02 U5438 ( .A0(n446), .A1(r32_mux_0_data[13]), .Z(n4880));
Q_AN02 U5439 ( .A0(n446), .A1(r32_mux_0_data[14]), .Z(n4881));
Q_AN02 U5440 ( .A0(n446), .A1(r32_mux_0_data[15]), .Z(n4882));
Q_AN02 U5441 ( .A0(n446), .A1(r32_mux_0_data[16]), .Z(n4883));
Q_AN02 U5442 ( .A0(n446), .A1(r32_mux_0_data[17]), .Z(n4884));
Q_AN02 U5443 ( .A0(n446), .A1(r32_mux_0_data[18]), .Z(n4885));
Q_AN02 U5444 ( .A0(n446), .A1(r32_mux_0_data[19]), .Z(n4886));
Q_AN02 U5445 ( .A0(n446), .A1(r32_mux_0_data[20]), .Z(n4887));
Q_AN02 U5446 ( .A0(n446), .A1(r32_mux_0_data[21]), .Z(n4888));
Q_AN02 U5447 ( .A0(n446), .A1(r32_mux_0_data[22]), .Z(n4889));
Q_AN02 U5448 ( .A0(n446), .A1(r32_mux_0_data[23]), .Z(n4890));
Q_AN02 U5449 ( .A0(n446), .A1(r32_mux_0_data[24]), .Z(n4891));
Q_AN02 U5450 ( .A0(n446), .A1(r32_mux_0_data[25]), .Z(n4892));
Q_AN02 U5451 ( .A0(n446), .A1(r32_mux_0_data[26]), .Z(n4893));
Q_AN02 U5452 ( .A0(n446), .A1(r32_mux_0_data[27]), .Z(n4894));
Q_AN02 U5453 ( .A0(n446), .A1(r32_mux_0_data[28]), .Z(n4895));
Q_AN02 U5454 ( .A0(n446), .A1(r32_mux_0_data[29]), .Z(n4896));
Q_AN02 U5455 ( .A0(n446), .A1(r32_mux_0_data[30]), .Z(n4897));
Q_AN02 U5456 ( .A0(n446), .A1(r32_mux_0_data[31]), .Z(n4898));
Q_AN02 U5457 ( .A0(n446), .A1(w_next_err_ack), .Z(n4899));
Q_AN02 U5458 ( .A0(n446), .A1(n4608), .Z(n4900));
Q_AN02 U5459 ( .A0(n446), .A1(w_do_read), .Z(n4901));
Q_AN02 U5460 ( .A0(n446), .A1(w_next_state[0]), .Z(n4902));
Q_NR02 U5461 ( .A0(i_sw_init), .A1(n440), .Z(n4903));
Q_NR02 U5462 ( .A0(i_sw_init), .A1(n439), .Z(n4904));
Q_AN02 U5463 ( .A0(n446), .A1(i_addr[0]), .Z(n4905));
Q_AN02 U5464 ( .A0(n446), .A1(i_addr[1]), .Z(n4906));
Q_AN02 U5465 ( .A0(n446), .A1(i_addr[2]), .Z(n4907));
Q_AN02 U5466 ( .A0(n446), .A1(i_addr[3]), .Z(n4908));
Q_AN02 U5467 ( .A0(n446), .A1(i_addr[4]), .Z(n4909));
Q_AN02 U5468 ( .A0(n446), .A1(i_addr[5]), .Z(n4910));
Q_AN02 U5469 ( .A0(n446), .A1(i_addr[6]), .Z(n4911));
Q_AN02 U5470 ( .A0(n446), .A1(i_addr[7]), .Z(n4912));
Q_AN02 U5471 ( .A0(n446), .A1(i_addr[8]), .Z(n4913));
Q_AN02 U5472 ( .A0(n446), .A1(i_addr[9]), .Z(n4914));
Q_AN02 U5473 ( .A0(n446), .A1(i_addr[10]), .Z(n4915));
Q_AN02 U5474 ( .A0(n446), .A1(n4610), .Z(n4916));
Q_AN02 U5475 ( .A0(n446), .A1(n4609), .Z(n4917));
Q_FDP1 o_reg_written_REG  ( .CK(clk), .R(i_reset_), .D(n4917), .Q(o_reg_written), .QN( ));
Q_FDP1 o_reg_read_REG  ( .CK(clk), .R(i_reset_), .D(n4916), .Q(o_reg_read), .QN( ));
Q_FDP1 \f_state_REG[2] ( .CK(clk), .R(i_reset_), .D(n4904), .Q(f_state[2]), .QN(n436));
Q_FDP1 \f_state_REG[1] ( .CK(clk), .R(i_reset_), .D(n4903), .Q(f_state[1]), .QN(n121));
Q_FDP1 \f_state_REG[0] ( .CK(clk), .R(i_reset_), .D(n4902), .Q(f_state[0]), .QN(n435));
Q_FDP1 f_prev_do_read_REG  ( .CK(clk), .R(i_reset_), .D(n4901), .Q(f_prev_do_read), .QN( ));
Q_FDP1 f_ack_REG  ( .CK(clk), .R(i_reset_), .D(n4900), .Q(f_ack), .QN( ));
Q_FDP1 f_err_ack_REG  ( .CK(clk), .R(i_reset_), .D(n4899), .Q(f_err_ack), .QN( ));
Q_ND02 U5484 ( .A0(n448), .A1(n4607), .Z(n4918));
Q_OR02 U5485 ( .A0(i_sw_init), .A1(w_do_read), .Z(n4919));
Q_INV U5486 ( .A(n98), .Z(n4921));
Q_INV U5487 ( .A(n109), .Z(n4922));
Q_INV U5488 ( .A(n82), .Z(n4923));
Q_INV U5489 ( .A(n90), .Z(n4924));
Q_INV U5490 ( .A(n83), .Z(n4925));
Q_FDP4EP \f32_data_REG[31] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[31]), .Q(f32_data[31]));
Q_FDP4EP \f32_data_REG[30] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[30]), .Q(f32_data[30]));
Q_FDP4EP \f32_data_REG[29] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[29]), .Q(f32_data[29]));
Q_FDP4EP \f32_data_REG[28] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[28]), .Q(f32_data[28]));
Q_FDP4EP \f32_data_REG[27] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[27]), .Q(f32_data[27]));
Q_FDP4EP \f32_data_REG[26] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[26]), .Q(f32_data[26]));
Q_FDP4EP \f32_data_REG[25] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[25]), .Q(f32_data[25]));
Q_FDP4EP \f32_data_REG[24] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[24]), .Q(f32_data[24]));
Q_FDP4EP \f32_data_REG[23] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[23]), .Q(f32_data[23]));
Q_FDP4EP \f32_data_REG[22] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[22]), .Q(f32_data[22]));
Q_FDP4EP \f32_data_REG[21] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[21]), .Q(f32_data[21]));
Q_FDP4EP \f32_data_REG[20] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[20]), .Q(f32_data[20]));
Q_FDP4EP \f32_data_REG[19] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[19]), .Q(f32_data[19]));
Q_FDP4EP \f32_data_REG[18] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[18]), .Q(f32_data[18]));
Q_FDP4EP \f32_data_REG[17] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[17]), .Q(f32_data[17]));
Q_FDP4EP \f32_data_REG[16] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[16]), .Q(f32_data[16]));
Q_FDP4EP \f32_data_REG[15] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[15]), .Q(f32_data[15]));
Q_FDP4EP \f32_data_REG[14] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[14]), .Q(f32_data[14]));
Q_FDP4EP \f32_data_REG[13] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[13]), .Q(f32_data[13]));
Q_FDP4EP \f32_data_REG[12] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[12]), .Q(f32_data[12]));
Q_FDP4EP \f32_data_REG[11] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[11]), .Q(f32_data[11]));
Q_FDP4EP \f32_data_REG[10] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[10]), .Q(f32_data[10]));
Q_FDP4EP \f32_data_REG[9] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[9]), .Q(f32_data[9]));
Q_FDP4EP \f32_data_REG[8] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[8]), .Q(f32_data[8]));
Q_FDP4EP \f32_data_REG[7] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[7]), .Q(f32_data[7]));
Q_FDP4EP \f32_data_REG[6] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[6]), .Q(f32_data[6]));
Q_FDP4EP \f32_data_REG[5] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[5]), .Q(f32_data[5]));
Q_FDP4EP \f32_data_REG[4] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[4]), .Q(f32_data[4]));
Q_FDP4EP \f32_data_REG[3] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[3]), .Q(f32_data[3]));
Q_FDP4EP \f32_data_REG[2] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[2]), .Q(f32_data[2]));
Q_FDP4EP \f32_data_REG[1] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[1]), .Q(f32_data[1]));
Q_FDP4EP \f32_data_REG[0] ( .CK(clk), .CE(i_wr_strb), .R(n4920), .D(i_wr_data[0]), .Q(f32_data[0]));
Q_FDP4EP \f32_mux_8_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4611), .Q(f32_mux_8_data[0]));
Q_INV U5524 ( .A(i_reset_), .Z(n4926));
Q_FDP4EP \f32_mux_8_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4612), .Q(f32_mux_8_data[1]));
Q_FDP4EP \f32_mux_8_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4613), .Q(f32_mux_8_data[2]));
Q_FDP4EP \f32_mux_8_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4614), .Q(f32_mux_8_data[3]));
Q_FDP4EP \f32_mux_8_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4615), .Q(f32_mux_8_data[4]));
Q_FDP4EP \f32_mux_8_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4616), .Q(f32_mux_8_data[5]));
Q_FDP4EP \f32_mux_8_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4617), .Q(f32_mux_8_data[6]));
Q_FDP4EP \f32_mux_8_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4618), .Q(f32_mux_8_data[7]));
Q_FDP4EP \f32_mux_8_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4619), .Q(f32_mux_8_data[8]));
Q_FDP4EP \f32_mux_8_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4620), .Q(f32_mux_8_data[9]));
Q_FDP4EP \f32_mux_8_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4621), .Q(f32_mux_8_data[10]));
Q_FDP4EP \f32_mux_8_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4622), .Q(f32_mux_8_data[11]));
Q_FDP4EP \f32_mux_8_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4623), .Q(f32_mux_8_data[12]));
Q_FDP4EP \f32_mux_8_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4624), .Q(f32_mux_8_data[13]));
Q_FDP4EP \f32_mux_8_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4625), .Q(f32_mux_8_data[14]));
Q_FDP4EP \f32_mux_8_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4626), .Q(f32_mux_8_data[15]));
Q_FDP4EP \f32_mux_8_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4627), .Q(f32_mux_8_data[16]));
Q_FDP4EP \f32_mux_8_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4628), .Q(f32_mux_8_data[17]));
Q_FDP4EP \f32_mux_8_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4629), .Q(f32_mux_8_data[18]));
Q_FDP4EP \f32_mux_8_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4630), .Q(f32_mux_8_data[19]));
Q_FDP4EP \f32_mux_8_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4631), .Q(f32_mux_8_data[20]));
Q_FDP4EP \f32_mux_8_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4632), .Q(f32_mux_8_data[21]));
Q_FDP4EP \f32_mux_8_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4633), .Q(f32_mux_8_data[22]));
Q_FDP4EP \f32_mux_8_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4634), .Q(f32_mux_8_data[23]));
Q_FDP4EP \f32_mux_8_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4635), .Q(f32_mux_8_data[24]));
Q_FDP4EP \f32_mux_8_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4636), .Q(f32_mux_8_data[25]));
Q_FDP4EP \f32_mux_8_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4637), .Q(f32_mux_8_data[26]));
Q_FDP4EP \f32_mux_8_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4638), .Q(f32_mux_8_data[27]));
Q_FDP4EP \f32_mux_8_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4639), .Q(f32_mux_8_data[28]));
Q_FDP4EP \f32_mux_8_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4640), .Q(f32_mux_8_data[29]));
Q_FDP4EP \f32_mux_8_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4641), .Q(f32_mux_8_data[30]));
Q_FDP4EP \f32_mux_8_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4642), .Q(f32_mux_8_data[31]));
Q_FDP4EP \f32_mux_7_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4643), .Q(f32_mux_7_data[0]));
Q_FDP4EP \f32_mux_7_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4644), .Q(f32_mux_7_data[1]));
Q_FDP4EP \f32_mux_7_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4645), .Q(f32_mux_7_data[2]));
Q_FDP4EP \f32_mux_7_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4646), .Q(f32_mux_7_data[3]));
Q_FDP4EP \f32_mux_7_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4647), .Q(f32_mux_7_data[4]));
Q_FDP4EP \f32_mux_7_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4648), .Q(f32_mux_7_data[5]));
Q_FDP4EP \f32_mux_7_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4649), .Q(f32_mux_7_data[6]));
Q_FDP4EP \f32_mux_7_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4650), .Q(f32_mux_7_data[7]));
Q_FDP4EP \f32_mux_7_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4651), .Q(f32_mux_7_data[8]));
Q_FDP4EP \f32_mux_7_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4652), .Q(f32_mux_7_data[9]));
Q_FDP4EP \f32_mux_7_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4653), .Q(f32_mux_7_data[10]));
Q_FDP4EP \f32_mux_7_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4654), .Q(f32_mux_7_data[11]));
Q_FDP4EP \f32_mux_7_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4655), .Q(f32_mux_7_data[12]));
Q_FDP4EP \f32_mux_7_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4656), .Q(f32_mux_7_data[13]));
Q_FDP4EP \f32_mux_7_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4657), .Q(f32_mux_7_data[14]));
Q_FDP4EP \f32_mux_7_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4658), .Q(f32_mux_7_data[15]));
Q_FDP4EP \f32_mux_7_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4659), .Q(f32_mux_7_data[16]));
Q_FDP4EP \f32_mux_7_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4660), .Q(f32_mux_7_data[17]));
Q_FDP4EP \f32_mux_7_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4661), .Q(f32_mux_7_data[18]));
Q_FDP4EP \f32_mux_7_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4662), .Q(f32_mux_7_data[19]));
Q_FDP4EP \f32_mux_7_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4663), .Q(f32_mux_7_data[20]));
Q_FDP4EP \f32_mux_7_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4664), .Q(f32_mux_7_data[21]));
Q_FDP4EP \f32_mux_7_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4665), .Q(f32_mux_7_data[22]));
Q_FDP4EP \f32_mux_7_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4666), .Q(f32_mux_7_data[23]));
Q_FDP4EP \f32_mux_7_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4667), .Q(f32_mux_7_data[24]));
Q_FDP4EP \f32_mux_7_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4668), .Q(f32_mux_7_data[25]));
Q_FDP4EP \f32_mux_7_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4669), .Q(f32_mux_7_data[26]));
Q_FDP4EP \f32_mux_7_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4670), .Q(f32_mux_7_data[27]));
Q_FDP4EP \f32_mux_7_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4671), .Q(f32_mux_7_data[28]));
Q_FDP4EP \f32_mux_7_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4672), .Q(f32_mux_7_data[29]));
Q_FDP4EP \f32_mux_7_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4673), .Q(f32_mux_7_data[30]));
Q_FDP4EP \f32_mux_7_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4674), .Q(f32_mux_7_data[31]));
Q_FDP4EP \f32_mux_6_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4675), .Q(f32_mux_6_data[0]));
Q_FDP4EP \f32_mux_6_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4676), .Q(f32_mux_6_data[1]));
Q_FDP4EP \f32_mux_6_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4677), .Q(f32_mux_6_data[2]));
Q_FDP4EP \f32_mux_6_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4678), .Q(f32_mux_6_data[3]));
Q_FDP4EP \f32_mux_6_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4679), .Q(f32_mux_6_data[4]));
Q_FDP4EP \f32_mux_6_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4680), .Q(f32_mux_6_data[5]));
Q_FDP4EP \f32_mux_6_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4681), .Q(f32_mux_6_data[6]));
Q_FDP4EP \f32_mux_6_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4682), .Q(f32_mux_6_data[7]));
Q_FDP4EP \f32_mux_6_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4683), .Q(f32_mux_6_data[8]));
Q_FDP4EP \f32_mux_6_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4684), .Q(f32_mux_6_data[9]));
Q_FDP4EP \f32_mux_6_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4685), .Q(f32_mux_6_data[10]));
Q_FDP4EP \f32_mux_6_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4686), .Q(f32_mux_6_data[11]));
Q_FDP4EP \f32_mux_6_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4687), .Q(f32_mux_6_data[12]));
Q_FDP4EP \f32_mux_6_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4688), .Q(f32_mux_6_data[13]));
Q_FDP4EP \f32_mux_6_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4689), .Q(f32_mux_6_data[14]));
Q_FDP4EP \f32_mux_6_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4690), .Q(f32_mux_6_data[15]));
Q_FDP4EP \f32_mux_6_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4691), .Q(f32_mux_6_data[16]));
Q_FDP4EP \f32_mux_6_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4692), .Q(f32_mux_6_data[17]));
Q_FDP4EP \f32_mux_6_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4693), .Q(f32_mux_6_data[18]));
Q_FDP4EP \f32_mux_6_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4694), .Q(f32_mux_6_data[19]));
Q_FDP4EP \f32_mux_6_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4695), .Q(f32_mux_6_data[20]));
Q_FDP4EP \f32_mux_6_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4696), .Q(f32_mux_6_data[21]));
Q_FDP4EP \f32_mux_6_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4697), .Q(f32_mux_6_data[22]));
Q_FDP4EP \f32_mux_6_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4698), .Q(f32_mux_6_data[23]));
Q_FDP4EP \f32_mux_6_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4699), .Q(f32_mux_6_data[24]));
Q_FDP4EP \f32_mux_6_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4700), .Q(f32_mux_6_data[25]));
Q_FDP4EP \f32_mux_6_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4701), .Q(f32_mux_6_data[26]));
Q_FDP4EP \f32_mux_6_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4702), .Q(f32_mux_6_data[27]));
Q_FDP4EP \f32_mux_6_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4703), .Q(f32_mux_6_data[28]));
Q_FDP4EP \f32_mux_6_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4704), .Q(f32_mux_6_data[29]));
Q_FDP4EP \f32_mux_6_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4705), .Q(f32_mux_6_data[30]));
Q_FDP4EP \f32_mux_6_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4706), .Q(f32_mux_6_data[31]));
Q_FDP4EP \f32_mux_5_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4707), .Q(f32_mux_5_data[0]));
Q_FDP4EP \f32_mux_5_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4708), .Q(f32_mux_5_data[1]));
Q_FDP4EP \f32_mux_5_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4709), .Q(f32_mux_5_data[2]));
Q_FDP4EP \f32_mux_5_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4710), .Q(f32_mux_5_data[3]));
Q_FDP4EP \f32_mux_5_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4711), .Q(f32_mux_5_data[4]));
Q_FDP4EP \f32_mux_5_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4712), .Q(f32_mux_5_data[5]));
Q_FDP4EP \f32_mux_5_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4713), .Q(f32_mux_5_data[6]));
Q_FDP4EP \f32_mux_5_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4714), .Q(f32_mux_5_data[7]));
Q_FDP4EP \f32_mux_5_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4715), .Q(f32_mux_5_data[8]));
Q_FDP4EP \f32_mux_5_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4716), .Q(f32_mux_5_data[9]));
Q_FDP4EP \f32_mux_5_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4717), .Q(f32_mux_5_data[10]));
Q_FDP4EP \f32_mux_5_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4718), .Q(f32_mux_5_data[11]));
Q_FDP4EP \f32_mux_5_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4719), .Q(f32_mux_5_data[12]));
Q_FDP4EP \f32_mux_5_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4720), .Q(f32_mux_5_data[13]));
Q_FDP4EP \f32_mux_5_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4721), .Q(f32_mux_5_data[14]));
Q_FDP4EP \f32_mux_5_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4722), .Q(f32_mux_5_data[15]));
Q_FDP4EP \f32_mux_5_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4723), .Q(f32_mux_5_data[16]));
Q_FDP4EP \f32_mux_5_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4724), .Q(f32_mux_5_data[17]));
Q_FDP4EP \f32_mux_5_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4725), .Q(f32_mux_5_data[18]));
Q_FDP4EP \f32_mux_5_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4726), .Q(f32_mux_5_data[19]));
Q_FDP4EP \f32_mux_5_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4727), .Q(f32_mux_5_data[20]));
Q_FDP4EP \f32_mux_5_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4728), .Q(f32_mux_5_data[21]));
Q_FDP4EP \f32_mux_5_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4729), .Q(f32_mux_5_data[22]));
Q_FDP4EP \f32_mux_5_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4730), .Q(f32_mux_5_data[23]));
Q_FDP4EP \f32_mux_5_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4731), .Q(f32_mux_5_data[24]));
Q_FDP4EP \f32_mux_5_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4732), .Q(f32_mux_5_data[25]));
Q_FDP4EP \f32_mux_5_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4733), .Q(f32_mux_5_data[26]));
Q_FDP4EP \f32_mux_5_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4734), .Q(f32_mux_5_data[27]));
Q_FDP4EP \f32_mux_5_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4735), .Q(f32_mux_5_data[28]));
Q_FDP4EP \f32_mux_5_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4736), .Q(f32_mux_5_data[29]));
Q_FDP4EP \f32_mux_5_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4737), .Q(f32_mux_5_data[30]));
Q_FDP4EP \f32_mux_5_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4738), .Q(f32_mux_5_data[31]));
Q_FDP4EP \f32_mux_4_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4739), .Q(f32_mux_4_data[0]));
Q_FDP4EP \f32_mux_4_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4740), .Q(f32_mux_4_data[1]));
Q_FDP4EP \f32_mux_4_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4741), .Q(f32_mux_4_data[2]));
Q_FDP4EP \f32_mux_4_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4742), .Q(f32_mux_4_data[3]));
Q_FDP4EP \f32_mux_4_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4743), .Q(f32_mux_4_data[4]));
Q_FDP4EP \f32_mux_4_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4744), .Q(f32_mux_4_data[5]));
Q_FDP4EP \f32_mux_4_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4745), .Q(f32_mux_4_data[6]));
Q_FDP4EP \f32_mux_4_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4746), .Q(f32_mux_4_data[7]));
Q_FDP4EP \f32_mux_4_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4747), .Q(f32_mux_4_data[8]));
Q_FDP4EP \f32_mux_4_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4748), .Q(f32_mux_4_data[9]));
Q_FDP4EP \f32_mux_4_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4749), .Q(f32_mux_4_data[10]));
Q_FDP4EP \f32_mux_4_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4750), .Q(f32_mux_4_data[11]));
Q_FDP4EP \f32_mux_4_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4751), .Q(f32_mux_4_data[12]));
Q_FDP4EP \f32_mux_4_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4752), .Q(f32_mux_4_data[13]));
Q_FDP4EP \f32_mux_4_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4753), .Q(f32_mux_4_data[14]));
Q_FDP4EP \f32_mux_4_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4754), .Q(f32_mux_4_data[15]));
Q_FDP4EP \f32_mux_4_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4755), .Q(f32_mux_4_data[16]));
Q_FDP4EP \f32_mux_4_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4756), .Q(f32_mux_4_data[17]));
Q_FDP4EP \f32_mux_4_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4757), .Q(f32_mux_4_data[18]));
Q_FDP4EP \f32_mux_4_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4758), .Q(f32_mux_4_data[19]));
Q_FDP4EP \f32_mux_4_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4759), .Q(f32_mux_4_data[20]));
Q_FDP4EP \f32_mux_4_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4760), .Q(f32_mux_4_data[21]));
Q_FDP4EP \f32_mux_4_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4761), .Q(f32_mux_4_data[22]));
Q_FDP4EP \f32_mux_4_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4762), .Q(f32_mux_4_data[23]));
Q_FDP4EP \f32_mux_4_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4763), .Q(f32_mux_4_data[24]));
Q_FDP4EP \f32_mux_4_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4764), .Q(f32_mux_4_data[25]));
Q_FDP4EP \f32_mux_4_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4765), .Q(f32_mux_4_data[26]));
Q_FDP4EP \f32_mux_4_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4766), .Q(f32_mux_4_data[27]));
Q_FDP4EP \f32_mux_4_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4767), .Q(f32_mux_4_data[28]));
Q_FDP4EP \f32_mux_4_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4768), .Q(f32_mux_4_data[29]));
Q_FDP4EP \f32_mux_4_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4769), .Q(f32_mux_4_data[30]));
Q_FDP4EP \f32_mux_4_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4770), .Q(f32_mux_4_data[31]));
Q_FDP4EP \f32_mux_3_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4771), .Q(f32_mux_3_data[0]));
Q_FDP4EP \f32_mux_3_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4772), .Q(f32_mux_3_data[1]));
Q_FDP4EP \f32_mux_3_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4773), .Q(f32_mux_3_data[2]));
Q_FDP4EP \f32_mux_3_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4774), .Q(f32_mux_3_data[3]));
Q_FDP4EP \f32_mux_3_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4775), .Q(f32_mux_3_data[4]));
Q_FDP4EP \f32_mux_3_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4776), .Q(f32_mux_3_data[5]));
Q_FDP4EP \f32_mux_3_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4777), .Q(f32_mux_3_data[6]));
Q_FDP4EP \f32_mux_3_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4778), .Q(f32_mux_3_data[7]));
Q_FDP4EP \f32_mux_3_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4779), .Q(f32_mux_3_data[8]));
Q_FDP4EP \f32_mux_3_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4780), .Q(f32_mux_3_data[9]));
Q_FDP4EP \f32_mux_3_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4781), .Q(f32_mux_3_data[10]));
Q_FDP4EP \f32_mux_3_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4782), .Q(f32_mux_3_data[11]));
Q_FDP4EP \f32_mux_3_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4783), .Q(f32_mux_3_data[12]));
Q_FDP4EP \f32_mux_3_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4784), .Q(f32_mux_3_data[13]));
Q_FDP4EP \f32_mux_3_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4785), .Q(f32_mux_3_data[14]));
Q_FDP4EP \f32_mux_3_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4786), .Q(f32_mux_3_data[15]));
Q_FDP4EP \f32_mux_3_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4787), .Q(f32_mux_3_data[16]));
Q_FDP4EP \f32_mux_3_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4788), .Q(f32_mux_3_data[17]));
Q_FDP4EP \f32_mux_3_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4789), .Q(f32_mux_3_data[18]));
Q_FDP4EP \f32_mux_3_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4790), .Q(f32_mux_3_data[19]));
Q_FDP4EP \f32_mux_3_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4791), .Q(f32_mux_3_data[20]));
Q_FDP4EP \f32_mux_3_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4792), .Q(f32_mux_3_data[21]));
Q_FDP4EP \f32_mux_3_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4793), .Q(f32_mux_3_data[22]));
Q_FDP4EP \f32_mux_3_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4794), .Q(f32_mux_3_data[23]));
Q_FDP4EP \f32_mux_3_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4795), .Q(f32_mux_3_data[24]));
Q_FDP4EP \f32_mux_3_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4796), .Q(f32_mux_3_data[25]));
Q_FDP4EP \f32_mux_3_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4797), .Q(f32_mux_3_data[26]));
Q_FDP4EP \f32_mux_3_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4798), .Q(f32_mux_3_data[27]));
Q_FDP4EP \f32_mux_3_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4799), .Q(f32_mux_3_data[28]));
Q_FDP4EP \f32_mux_3_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4800), .Q(f32_mux_3_data[29]));
Q_FDP4EP \f32_mux_3_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4801), .Q(f32_mux_3_data[30]));
Q_FDP4EP \f32_mux_3_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4802), .Q(f32_mux_3_data[31]));
Q_FDP4EP \f32_mux_2_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4803), .Q(f32_mux_2_data[0]));
Q_FDP4EP \f32_mux_2_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4804), .Q(f32_mux_2_data[1]));
Q_FDP4EP \f32_mux_2_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4805), .Q(f32_mux_2_data[2]));
Q_FDP4EP \f32_mux_2_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4806), .Q(f32_mux_2_data[3]));
Q_FDP4EP \f32_mux_2_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4807), .Q(f32_mux_2_data[4]));
Q_FDP4EP \f32_mux_2_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4808), .Q(f32_mux_2_data[5]));
Q_FDP4EP \f32_mux_2_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4809), .Q(f32_mux_2_data[6]));
Q_FDP4EP \f32_mux_2_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4810), .Q(f32_mux_2_data[7]));
Q_FDP4EP \f32_mux_2_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4811), .Q(f32_mux_2_data[8]));
Q_FDP4EP \f32_mux_2_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4812), .Q(f32_mux_2_data[9]));
Q_FDP4EP \f32_mux_2_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4813), .Q(f32_mux_2_data[10]));
Q_FDP4EP \f32_mux_2_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4814), .Q(f32_mux_2_data[11]));
Q_FDP4EP \f32_mux_2_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4815), .Q(f32_mux_2_data[12]));
Q_FDP4EP \f32_mux_2_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4816), .Q(f32_mux_2_data[13]));
Q_FDP4EP \f32_mux_2_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4817), .Q(f32_mux_2_data[14]));
Q_FDP4EP \f32_mux_2_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4818), .Q(f32_mux_2_data[15]));
Q_FDP4EP \f32_mux_2_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4819), .Q(f32_mux_2_data[16]));
Q_FDP4EP \f32_mux_2_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4820), .Q(f32_mux_2_data[17]));
Q_FDP4EP \f32_mux_2_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4821), .Q(f32_mux_2_data[18]));
Q_FDP4EP \f32_mux_2_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4822), .Q(f32_mux_2_data[19]));
Q_FDP4EP \f32_mux_2_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4823), .Q(f32_mux_2_data[20]));
Q_FDP4EP \f32_mux_2_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4824), .Q(f32_mux_2_data[21]));
Q_FDP4EP \f32_mux_2_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4825), .Q(f32_mux_2_data[22]));
Q_FDP4EP \f32_mux_2_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4826), .Q(f32_mux_2_data[23]));
Q_FDP4EP \f32_mux_2_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4827), .Q(f32_mux_2_data[24]));
Q_FDP4EP \f32_mux_2_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4828), .Q(f32_mux_2_data[25]));
Q_FDP4EP \f32_mux_2_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4829), .Q(f32_mux_2_data[26]));
Q_FDP4EP \f32_mux_2_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4830), .Q(f32_mux_2_data[27]));
Q_FDP4EP \f32_mux_2_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4831), .Q(f32_mux_2_data[28]));
Q_FDP4EP \f32_mux_2_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4832), .Q(f32_mux_2_data[29]));
Q_FDP4EP \f32_mux_2_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4833), .Q(f32_mux_2_data[30]));
Q_FDP4EP \f32_mux_2_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4834), .Q(f32_mux_2_data[31]));
Q_FDP4EP \f32_mux_1_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4835), .Q(f32_mux_1_data[0]));
Q_FDP4EP \f32_mux_1_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4836), .Q(f32_mux_1_data[1]));
Q_FDP4EP \f32_mux_1_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4837), .Q(f32_mux_1_data[2]));
Q_FDP4EP \f32_mux_1_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4838), .Q(f32_mux_1_data[3]));
Q_FDP4EP \f32_mux_1_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4839), .Q(f32_mux_1_data[4]));
Q_FDP4EP \f32_mux_1_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4840), .Q(f32_mux_1_data[5]));
Q_FDP4EP \f32_mux_1_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4841), .Q(f32_mux_1_data[6]));
Q_FDP4EP \f32_mux_1_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4842), .Q(f32_mux_1_data[7]));
Q_FDP4EP \f32_mux_1_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4843), .Q(f32_mux_1_data[8]));
Q_FDP4EP \f32_mux_1_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4844), .Q(f32_mux_1_data[9]));
Q_FDP4EP \f32_mux_1_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4845), .Q(f32_mux_1_data[10]));
Q_FDP4EP \f32_mux_1_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4846), .Q(f32_mux_1_data[11]));
Q_FDP4EP \f32_mux_1_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4847), .Q(f32_mux_1_data[12]));
Q_FDP4EP \f32_mux_1_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4848), .Q(f32_mux_1_data[13]));
Q_FDP4EP \f32_mux_1_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4849), .Q(f32_mux_1_data[14]));
Q_FDP4EP \f32_mux_1_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4850), .Q(f32_mux_1_data[15]));
Q_FDP4EP \f32_mux_1_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4851), .Q(f32_mux_1_data[16]));
Q_FDP4EP \f32_mux_1_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4852), .Q(f32_mux_1_data[17]));
Q_FDP4EP \f32_mux_1_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4853), .Q(f32_mux_1_data[18]));
Q_FDP4EP \f32_mux_1_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4854), .Q(f32_mux_1_data[19]));
Q_FDP4EP \f32_mux_1_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4855), .Q(f32_mux_1_data[20]));
Q_FDP4EP \f32_mux_1_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4856), .Q(f32_mux_1_data[21]));
Q_FDP4EP \f32_mux_1_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4857), .Q(f32_mux_1_data[22]));
Q_FDP4EP \f32_mux_1_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4858), .Q(f32_mux_1_data[23]));
Q_FDP4EP \f32_mux_1_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4859), .Q(f32_mux_1_data[24]));
Q_FDP4EP \f32_mux_1_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4860), .Q(f32_mux_1_data[25]));
Q_FDP4EP \f32_mux_1_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4861), .Q(f32_mux_1_data[26]));
Q_FDP4EP \f32_mux_1_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4862), .Q(f32_mux_1_data[27]));
Q_FDP4EP \f32_mux_1_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4863), .Q(f32_mux_1_data[28]));
Q_FDP4EP \f32_mux_1_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4864), .Q(f32_mux_1_data[29]));
Q_FDP4EP \f32_mux_1_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4865), .Q(f32_mux_1_data[30]));
Q_FDP4EP \f32_mux_1_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4866), .Q(f32_mux_1_data[31]));
Q_FDP4EP \f32_mux_0_data_REG[0] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4867), .Q(f32_mux_0_data[0]));
Q_FDP4EP \f32_mux_0_data_REG[1] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4868), .Q(f32_mux_0_data[1]));
Q_FDP4EP \f32_mux_0_data_REG[2] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4869), .Q(f32_mux_0_data[2]));
Q_FDP4EP \f32_mux_0_data_REG[3] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4870), .Q(f32_mux_0_data[3]));
Q_FDP4EP \f32_mux_0_data_REG[4] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4871), .Q(f32_mux_0_data[4]));
Q_FDP4EP \f32_mux_0_data_REG[5] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4872), .Q(f32_mux_0_data[5]));
Q_FDP4EP \f32_mux_0_data_REG[6] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4873), .Q(f32_mux_0_data[6]));
Q_FDP4EP \f32_mux_0_data_REG[7] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4874), .Q(f32_mux_0_data[7]));
Q_FDP4EP \f32_mux_0_data_REG[8] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4875), .Q(f32_mux_0_data[8]));
Q_FDP4EP \f32_mux_0_data_REG[9] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4876), .Q(f32_mux_0_data[9]));
Q_FDP4EP \f32_mux_0_data_REG[10] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4877), .Q(f32_mux_0_data[10]));
Q_FDP4EP \f32_mux_0_data_REG[11] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4878), .Q(f32_mux_0_data[11]));
Q_FDP4EP \f32_mux_0_data_REG[12] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4879), .Q(f32_mux_0_data[12]));
Q_FDP4EP \f32_mux_0_data_REG[13] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4880), .Q(f32_mux_0_data[13]));
Q_FDP4EP \f32_mux_0_data_REG[14] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4881), .Q(f32_mux_0_data[14]));
Q_FDP4EP \f32_mux_0_data_REG[15] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4882), .Q(f32_mux_0_data[15]));
Q_FDP4EP \f32_mux_0_data_REG[16] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4883), .Q(f32_mux_0_data[16]));
Q_FDP4EP \f32_mux_0_data_REG[17] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4884), .Q(f32_mux_0_data[17]));
Q_FDP4EP \f32_mux_0_data_REG[18] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4885), .Q(f32_mux_0_data[18]));
Q_FDP4EP \f32_mux_0_data_REG[19] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4886), .Q(f32_mux_0_data[19]));
Q_FDP4EP \f32_mux_0_data_REG[20] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4887), .Q(f32_mux_0_data[20]));
Q_FDP4EP \f32_mux_0_data_REG[21] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4888), .Q(f32_mux_0_data[21]));
Q_FDP4EP \f32_mux_0_data_REG[22] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4889), .Q(f32_mux_0_data[22]));
Q_FDP4EP \f32_mux_0_data_REG[23] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4890), .Q(f32_mux_0_data[23]));
Q_FDP4EP \f32_mux_0_data_REG[24] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4891), .Q(f32_mux_0_data[24]));
Q_FDP4EP \f32_mux_0_data_REG[25] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4892), .Q(f32_mux_0_data[25]));
Q_FDP4EP \f32_mux_0_data_REG[26] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4893), .Q(f32_mux_0_data[26]));
Q_FDP4EP \f32_mux_0_data_REG[27] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4894), .Q(f32_mux_0_data[27]));
Q_FDP4EP \f32_mux_0_data_REG[28] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4895), .Q(f32_mux_0_data[28]));
Q_FDP4EP \f32_mux_0_data_REG[29] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4896), .Q(f32_mux_0_data[29]));
Q_FDP4EP \f32_mux_0_data_REG[30] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4897), .Q(f32_mux_0_data[30]));
Q_FDP4EP \f32_mux_0_data_REG[31] ( .CK(clk), .CE(n4919), .R(n4926), .D(n4898), .Q(f32_mux_0_data[31]));
Q_FDP4EP \o_reg_addr_REG[0] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4905), .Q(o_reg_addr[0]));
Q_FDP4EP \o_reg_addr_REG[1] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4906), .Q(o_reg_addr[1]));
Q_FDP4EP \o_reg_addr_REG[2] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4907), .Q(o_reg_addr[2]));
Q_FDP4EP \o_reg_addr_REG[3] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4908), .Q(o_reg_addr[3]));
Q_FDP4EP \o_reg_addr_REG[4] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4909), .Q(o_reg_addr[4]));
Q_FDP4EP \o_reg_addr_REG[5] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4910), .Q(o_reg_addr[5]));
Q_FDP4EP \o_reg_addr_REG[6] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4911), .Q(o_reg_addr[6]));
Q_FDP4EP \o_reg_addr_REG[7] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4912), .Q(o_reg_addr[7]));
Q_FDP4EP \o_reg_addr_REG[8] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4913), .Q(o_reg_addr[8]));
Q_FDP4EP \o_reg_addr_REG[9] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4914), .Q(o_reg_addr[9]));
Q_FDP4EP \o_reg_addr_REG[10] ( .CK(clk), .CE(n4918), .R(n4926), .D(n4915), .Q(o_reg_addr[10]));
Q_FDP4EP n_write_REG  ( .CK(clk), .CE(n447), .R(n4926), .D(n451), .Q(n_write));
Q_INV U5824 ( .A(n_write), .Z(n444));
endmodule
