
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_kme_aes_256_drng ( seed_expired, drng_valid, drng_256_out, 
	drng_fifo_overflow, drng_fifo_underflow, drng_idle, start, seed, 
	seed_life, drng_ack, clk, rst_n);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output seed_expired;
output drng_valid;
output [127:0] drng_256_out;
output drng_fifo_overflow;
output drng_fifo_underflow;
output drng_idle;
input start;
input [383:0] seed;
input [47:0] seed_life;
input drng_ack;
input clk;
input rst_n;
wire CiphInStall;
wire KeyInStall;
wire fifo_in_stall;
wire [127:0] fifo_out;
wire _zy_simnet_seed_expired_0_w$;
wire _zy_simnet_drng_idle_1_w$;
wire [0:127] _zy_simnet_AesCiphOutR_2_w$;
wire _zy_simnet_AesCiphOutVldR_3_w$;
wire _zy_simnet_cio_4;
wire _zy_simnet_cio_5;
wire _zy_simnet_cio_6;
wire [0:127] _zy_simnet_CiphIn_7_w$;
wire _zy_simnet_CiphInVldR_8_w$;
wire _zy_simnet_CiphInLastR_9_w$;
wire _zy_simnet_cio_10;
wire [0:255] _zy_simnet_KeyIn_11_w$;
wire _zy_simnet_KeyInVld_12_w$;
wire _zy_simnet_cio_13;
wire [0:127] _zy_simnet_fifo_in_14_w$;
wire _zy_simnet_fifo_in_valid_15_w$;
wire _zy_simnet_cio_16;
wire [1:0] cur_state;
wire [1:0] nxt_state;
wire [127:0] CiphIn;
wire CiphInVldR;
wire CiphInLastR;
wire KeyInVld;
wire [255:0] KeyIn;
wire [127:0] AesCiphOutR;
wire AesCiphOutVldR;
wire fifo_in_valid;
wire [127:0] fifo_in;
wire [47:0] reseed_counter;
wire [47:0] reseed_counter_limit;
wire [255:0] internal_state_key;
wire [127:0] internal_state_value;
wire [2:0] in_count;
wire [2:0] out_count;
supply1 n1;
supply0 n2;
Q_BUF U0 ( .A(n2), .Z(_zy_simnet_cio_16));
Q_BUF U1 ( .A(n2), .Z(_zy_simnet_cio_13));
Q_BUF U2 ( .A(n1), .Z(_zy_simnet_cio_10));
Q_BUF U3 ( .A(n1), .Z(_zy_simnet_cio_6));
Q_BUF U4 ( .A(n2), .Z(_zy_simnet_cio_5));
Q_BUF U5 ( .A(n2), .Z(_zy_simnet_cio_4));
Q_XOR2 U6 ( .A0(out_count[1]), .A1(out_count[0]), .Z(n1150));
cr_kme_fifo_xcm59 rnd_fifo ( .fifo_in_stall( fifo_in_stall), .fifo_out( 
	fifo_out[127:0]), .fifo_out_valid( drng_valid), .fifo_overflow( 
	drng_fifo_overflow), .fifo_underflow( drng_fifo_underflow), .clk( 
	clk), .rst_n( rst_n), .fifo_in( _zy_simnet_fifo_in_14_w$[0:127]), 
	.fifo_in_valid( _zy_simnet_fifo_in_valid_15_w$), .fifo_out_ack( 
	drng_ack), .fifo_in_stall_override( _zy_simnet_cio_16));
AesSecIStub AesSecIStub ( .AesCiphOutR( _zy_simnet_AesCiphOutR_2_w$[0:127]), 
	.AesCiphOutVldR( _zy_simnet_AesCiphOutVldR_3_w$), .KeyInitStall( 
	KeyInStall), .CiphInStall( CiphInStall), .Aes128( _zy_simnet_cio_4), 
	.Aes192( _zy_simnet_cio_5), .Aes256( _zy_simnet_cio_6), .CiphIn( 
	_zy_simnet_CiphIn_7_w$[0:127]), .CiphInVldR( _zy_simnet_CiphInVldR_8_w$), 
	.CiphInLastR( _zy_simnet_CiphInLastR_9_w$), .EncryptEn( 
	_zy_simnet_cio_10), .KeyIn( _zy_simnet_KeyIn_11_w$[0:255]), 
	.KeyInitVldR( _zy_simnet_KeyInVld_12_w$), .AesCiphOutStall( 
	_zy_simnet_cio_13), .clk( clk), .rst_n( rst_n));
ixc_assign _zz_strnp_11 ( _zy_simnet_fifo_in_valid_15_w$, fifo_in_valid);
ixc_assign_128 _zz_strnp_10 ( _zy_simnet_fifo_in_14_w$[0:127], fifo_in[127:0]);
ixc_assign _zz_strnp_9 ( _zy_simnet_KeyInVld_12_w$, KeyInVld);
ixc_assign_256 _zz_strnp_8 ( _zy_simnet_KeyIn_11_w$[0:255], KeyIn[255:0]);
ixc_assign _zz_strnp_7 ( _zy_simnet_CiphInLastR_9_w$, CiphInLastR);
ixc_assign _zz_strnp_6 ( _zy_simnet_CiphInVldR_8_w$, CiphInVldR);
ixc_assign_128 _zz_strnp_5 ( _zy_simnet_CiphIn_7_w$[0:127], CiphIn[127:0]);
ixc_assign _zz_strnp_4 ( AesCiphOutVldR, _zy_simnet_AesCiphOutVldR_3_w$);
ixc_assign_128 _zz_strnp_3 ( AesCiphOutR[127:0], 
	_zy_simnet_AesCiphOutR_2_w$[0:127]);
ixc_assign _zz_strnp_2 ( _zy_simnet_drng_idle_1_w$, drng_idle);
ixc_assign _zz_strnp_1 ( _zy_simnet_seed_expired_0_w$, seed_expired);
ixc_assign_128 _zz_strnp_0 ( drng_256_out[127:0], fifo_out[127:0]);
Q_FDP1 \cur_state_REG[0] ( .CK(clk), .R(rst_n), .D(nxt_state[0]), .Q(cur_state[0]), .QN(n80));
Q_FDP1 \cur_state_REG[1] ( .CK(clk), .R(rst_n), .D(nxt_state[1]), .Q(cur_state[1]), .QN(n79));
Q_OR03 U23 ( .A0(out_count[0]), .A1(out_count[1]), .A2(n3), .Z(n4));
Q_INV U24 ( .A(n4), .Z(n85));
Q_XNR2 U25 ( .A0(reseed_counter_limit[0]), .A1(reseed_counter[0]), .Z(n5));
Q_XNR2 U26 ( .A0(reseed_counter_limit[1]), .A1(reseed_counter[1]), .Z(n6));
Q_XNR2 U27 ( .A0(reseed_counter_limit[2]), .A1(reseed_counter[2]), .Z(n7));
Q_XNR2 U28 ( .A0(reseed_counter_limit[3]), .A1(reseed_counter[3]), .Z(n8));
Q_XNR2 U29 ( .A0(reseed_counter_limit[4]), .A1(reseed_counter[4]), .Z(n9));
Q_XNR2 U30 ( .A0(reseed_counter_limit[5]), .A1(reseed_counter[5]), .Z(n10));
Q_XNR2 U31 ( .A0(reseed_counter_limit[6]), .A1(reseed_counter[6]), .Z(n11));
Q_XNR2 U32 ( .A0(reseed_counter_limit[7]), .A1(reseed_counter[7]), .Z(n12));
Q_XNR2 U33 ( .A0(reseed_counter_limit[8]), .A1(reseed_counter[8]), .Z(n13));
Q_XNR2 U34 ( .A0(reseed_counter_limit[9]), .A1(reseed_counter[9]), .Z(n14));
Q_XNR2 U35 ( .A0(reseed_counter_limit[10]), .A1(reseed_counter[10]), .Z(n15));
Q_XNR2 U36 ( .A0(reseed_counter_limit[11]), .A1(reseed_counter[11]), .Z(n16));
Q_XNR2 U37 ( .A0(reseed_counter_limit[12]), .A1(reseed_counter[12]), .Z(n17));
Q_XNR2 U38 ( .A0(reseed_counter_limit[13]), .A1(reseed_counter[13]), .Z(n18));
Q_XNR2 U39 ( .A0(reseed_counter_limit[14]), .A1(reseed_counter[14]), .Z(n19));
Q_XNR2 U40 ( .A0(reseed_counter_limit[15]), .A1(reseed_counter[15]), .Z(n20));
Q_XNR2 U41 ( .A0(reseed_counter_limit[16]), .A1(reseed_counter[16]), .Z(n21));
Q_XNR2 U42 ( .A0(reseed_counter_limit[17]), .A1(reseed_counter[17]), .Z(n22));
Q_XNR2 U43 ( .A0(reseed_counter_limit[18]), .A1(reseed_counter[18]), .Z(n23));
Q_XNR2 U44 ( .A0(reseed_counter_limit[19]), .A1(reseed_counter[19]), .Z(n24));
Q_XNR2 U45 ( .A0(reseed_counter_limit[20]), .A1(reseed_counter[20]), .Z(n25));
Q_XNR2 U46 ( .A0(reseed_counter_limit[21]), .A1(reseed_counter[21]), .Z(n26));
Q_XNR2 U47 ( .A0(reseed_counter_limit[22]), .A1(reseed_counter[22]), .Z(n27));
Q_XNR2 U48 ( .A0(reseed_counter_limit[23]), .A1(reseed_counter[23]), .Z(n28));
Q_XNR2 U49 ( .A0(reseed_counter_limit[24]), .A1(reseed_counter[24]), .Z(n29));
Q_XNR2 U50 ( .A0(reseed_counter_limit[25]), .A1(reseed_counter[25]), .Z(n30));
Q_XNR2 U51 ( .A0(reseed_counter_limit[26]), .A1(reseed_counter[26]), .Z(n31));
Q_XNR2 U52 ( .A0(reseed_counter_limit[27]), .A1(reseed_counter[27]), .Z(n32));
Q_XNR2 U53 ( .A0(reseed_counter_limit[28]), .A1(reseed_counter[28]), .Z(n33));
Q_XNR2 U54 ( .A0(reseed_counter_limit[29]), .A1(reseed_counter[29]), .Z(n34));
Q_XNR2 U55 ( .A0(reseed_counter_limit[30]), .A1(reseed_counter[30]), .Z(n35));
Q_XNR2 U56 ( .A0(reseed_counter_limit[31]), .A1(reseed_counter[31]), .Z(n36));
Q_XNR2 U57 ( .A0(reseed_counter_limit[32]), .A1(reseed_counter[32]), .Z(n37));
Q_XNR2 U58 ( .A0(reseed_counter_limit[33]), .A1(reseed_counter[33]), .Z(n38));
Q_XNR2 U59 ( .A0(reseed_counter_limit[34]), .A1(reseed_counter[34]), .Z(n39));
Q_XNR2 U60 ( .A0(reseed_counter_limit[35]), .A1(reseed_counter[35]), .Z(n40));
Q_XNR2 U61 ( .A0(reseed_counter_limit[36]), .A1(reseed_counter[36]), .Z(n41));
Q_XNR2 U62 ( .A0(reseed_counter_limit[37]), .A1(reseed_counter[37]), .Z(n42));
Q_XNR2 U63 ( .A0(reseed_counter_limit[38]), .A1(reseed_counter[38]), .Z(n43));
Q_XNR2 U64 ( .A0(reseed_counter_limit[39]), .A1(reseed_counter[39]), .Z(n44));
Q_XNR2 U65 ( .A0(reseed_counter_limit[40]), .A1(reseed_counter[40]), .Z(n45));
Q_XNR2 U66 ( .A0(reseed_counter_limit[41]), .A1(reseed_counter[41]), .Z(n46));
Q_XNR2 U67 ( .A0(reseed_counter_limit[42]), .A1(reseed_counter[42]), .Z(n47));
Q_XNR2 U68 ( .A0(reseed_counter_limit[43]), .A1(reseed_counter[43]), .Z(n48));
Q_XNR2 U69 ( .A0(reseed_counter_limit[44]), .A1(reseed_counter[44]), .Z(n49));
Q_XNR2 U70 ( .A0(reseed_counter_limit[45]), .A1(reseed_counter[45]), .Z(n50));
Q_XNR2 U71 ( .A0(reseed_counter_limit[46]), .A1(reseed_counter[46]), .Z(n51));
Q_XNR2 U72 ( .A0(reseed_counter_limit[47]), .A1(reseed_counter[47]), .Z(n52));
Q_AN03 U73 ( .A0(n52), .A1(n51), .A2(n50), .Z(n53));
Q_AN03 U74 ( .A0(n49), .A1(n48), .A2(n47), .Z(n54));
Q_AN03 U75 ( .A0(n46), .A1(n45), .A2(n44), .Z(n55));
Q_AN03 U76 ( .A0(n43), .A1(n42), .A2(n41), .Z(n56));
Q_AN03 U77 ( .A0(n40), .A1(n39), .A2(n38), .Z(n57));
Q_AN03 U78 ( .A0(n37), .A1(n36), .A2(n35), .Z(n58));
Q_AN03 U79 ( .A0(n34), .A1(n33), .A2(n32), .Z(n59));
Q_AN03 U80 ( .A0(n31), .A1(n30), .A2(n29), .Z(n60));
Q_AN03 U81 ( .A0(n28), .A1(n27), .A2(n26), .Z(n61));
Q_AN03 U82 ( .A0(n25), .A1(n24), .A2(n23), .Z(n62));
Q_AN03 U83 ( .A0(n22), .A1(n21), .A2(n20), .Z(n63));
Q_AN03 U84 ( .A0(n19), .A1(n18), .A2(n17), .Z(n64));
Q_AN03 U85 ( .A0(n16), .A1(n15), .A2(n14), .Z(n65));
Q_AN03 U86 ( .A0(n13), .A1(n12), .A2(n11), .Z(n66));
Q_AN03 U87 ( .A0(n10), .A1(n9), .A2(n8), .Z(n67));
Q_AN03 U88 ( .A0(n7), .A1(n6), .A2(n5), .Z(n68));
Q_AN03 U89 ( .A0(n53), .A1(n54), .A2(n55), .Z(n69));
Q_AN03 U90 ( .A0(n56), .A1(n57), .A2(n58), .Z(n70));
Q_AN03 U91 ( .A0(n59), .A1(n60), .A2(n61), .Z(n71));
Q_AN03 U92 ( .A0(n62), .A1(n63), .A2(n64), .Z(n72));
Q_AN03 U93 ( .A0(n65), .A1(n66), .A2(n67), .Z(n73));
Q_AN03 U94 ( .A0(n68), .A1(n69), .A2(n70), .Z(n74));
Q_AN03 U95 ( .A0(n71), .A1(n72), .A2(n73), .Z(n75));
Q_AO21 U96 ( .A0(n74), .A1(n75), .B0(n4), .Z(n81));
Q_XOR2 U97 ( .A0(n76), .A1(n84), .Z(nxt_state[0]));
Q_INV U98 ( .A(n84), .Z(nxt_state[1]));
Q_MX02 U99 ( .S(cur_state[1]), .A0(n77), .A1(n78), .Z(n76));
Q_NR02 U100 ( .A0(cur_state[0]), .A1(start), .Z(n77));
Q_MX02 U101 ( .S(cur_state[0]), .A0(CiphInLastR), .A1(n81), .Z(n78));
Q_MX02 U102 ( .S(cur_state[1]), .A0(n82), .A1(n83), .Z(n84));
Q_OR02 U103 ( .A0(n80), .A1(KeyInStall), .Z(n82));
Q_AN02 U104 ( .A0(cur_state[0]), .A1(n85), .Z(n83));
Q_NR02 U105 ( .A0(nxt_state[0]), .A1(nxt_state[1]), .Z(seed_expired));
Q_OR03 U106 ( .A0(in_count[0]), .A1(in_count[1]), .A2(n86), .Z(n87));
Q_INV U107 ( .A(n87), .Z(n88));
Q_AD01HF U108 ( .A0(internal_state_value[0]), .B0(in_count[0]), .S(n89), .CO(n90));
Q_AD02 U109 ( .CI(n90), .A0(internal_state_value[1]), .A1(internal_state_value[2]), .B0(in_count[1]), .B1(in_count[2]), .S0(n91), .S1(n92), .CO(n93));
Q_AD01HF U110 ( .A0(internal_state_value[3]), .B0(n93), .S(n94), .CO(n95));
Q_AD01HF U111 ( .A0(internal_state_value[4]), .B0(n95), .S(n96), .CO(n97));
Q_AD01HF U112 ( .A0(internal_state_value[5]), .B0(n97), .S(n98), .CO(n99));
Q_AD01HF U113 ( .A0(internal_state_value[6]), .B0(n99), .S(n100), .CO(n101));
Q_AD01HF U114 ( .A0(internal_state_value[7]), .B0(n101), .S(n102), .CO(n103));
Q_AD01HF U115 ( .A0(internal_state_value[8]), .B0(n103), .S(n104), .CO(n105));
Q_AD01HF U116 ( .A0(internal_state_value[9]), .B0(n105), .S(n106), .CO(n107));
Q_AD01HF U117 ( .A0(internal_state_value[10]), .B0(n107), .S(n108), .CO(n109));
Q_AD01HF U118 ( .A0(internal_state_value[11]), .B0(n109), .S(n110), .CO(n111));
Q_AD01HF U119 ( .A0(internal_state_value[12]), .B0(n111), .S(n112), .CO(n113));
Q_AD01HF U120 ( .A0(internal_state_value[13]), .B0(n113), .S(n114), .CO(n115));
Q_AD01HF U121 ( .A0(internal_state_value[14]), .B0(n115), .S(n116), .CO(n117));
Q_AD01HF U122 ( .A0(internal_state_value[15]), .B0(n117), .S(n118), .CO(n119));
Q_AD01HF U123 ( .A0(internal_state_value[16]), .B0(n119), .S(n120), .CO(n121));
Q_AD01HF U124 ( .A0(internal_state_value[17]), .B0(n121), .S(n122), .CO(n123));
Q_AD01HF U125 ( .A0(internal_state_value[18]), .B0(n123), .S(n124), .CO(n125));
Q_AD01HF U126 ( .A0(internal_state_value[19]), .B0(n125), .S(n126), .CO(n127));
Q_AD01HF U127 ( .A0(internal_state_value[20]), .B0(n127), .S(n128), .CO(n129));
Q_AD01HF U128 ( .A0(internal_state_value[21]), .B0(n129), .S(n130), .CO(n131));
Q_AD01HF U129 ( .A0(internal_state_value[22]), .B0(n131), .S(n132), .CO(n133));
Q_AD01HF U130 ( .A0(internal_state_value[23]), .B0(n133), .S(n134), .CO(n135));
Q_AD01HF U131 ( .A0(internal_state_value[24]), .B0(n135), .S(n136), .CO(n137));
Q_AD01HF U132 ( .A0(internal_state_value[25]), .B0(n137), .S(n138), .CO(n139));
Q_AD01HF U133 ( .A0(internal_state_value[26]), .B0(n139), .S(n140), .CO(n141));
Q_AD01HF U134 ( .A0(internal_state_value[27]), .B0(n141), .S(n142), .CO(n143));
Q_AD01HF U135 ( .A0(internal_state_value[28]), .B0(n143), .S(n144), .CO(n145));
Q_AD01HF U136 ( .A0(internal_state_value[29]), .B0(n145), .S(n146), .CO(n147));
Q_AD01HF U137 ( .A0(internal_state_value[30]), .B0(n147), .S(n148), .CO(n149));
Q_AD01HF U138 ( .A0(internal_state_value[31]), .B0(n149), .S(n150), .CO(n151));
Q_AD01HF U139 ( .A0(internal_state_value[32]), .B0(n151), .S(n152), .CO(n153));
Q_AD01HF U140 ( .A0(internal_state_value[33]), .B0(n153), .S(n154), .CO(n155));
Q_AD01HF U141 ( .A0(internal_state_value[34]), .B0(n155), .S(n156), .CO(n157));
Q_AD01HF U142 ( .A0(internal_state_value[35]), .B0(n157), .S(n158), .CO(n159));
Q_AD01HF U143 ( .A0(internal_state_value[36]), .B0(n159), .S(n160), .CO(n161));
Q_AD01HF U144 ( .A0(internal_state_value[37]), .B0(n161), .S(n162), .CO(n163));
Q_AD01HF U145 ( .A0(internal_state_value[38]), .B0(n163), .S(n164), .CO(n165));
Q_AD01HF U146 ( .A0(internal_state_value[39]), .B0(n165), .S(n166), .CO(n167));
Q_AD01HF U147 ( .A0(internal_state_value[40]), .B0(n167), .S(n168), .CO(n169));
Q_AD01HF U148 ( .A0(internal_state_value[41]), .B0(n169), .S(n170), .CO(n171));
Q_AD01HF U149 ( .A0(internal_state_value[42]), .B0(n171), .S(n172), .CO(n173));
Q_AD01HF U150 ( .A0(internal_state_value[43]), .B0(n173), .S(n174), .CO(n175));
Q_AD01HF U151 ( .A0(internal_state_value[44]), .B0(n175), .S(n176), .CO(n177));
Q_AD01HF U152 ( .A0(internal_state_value[45]), .B0(n177), .S(n178), .CO(n179));
Q_AD01HF U153 ( .A0(internal_state_value[46]), .B0(n179), .S(n180), .CO(n181));
Q_AD01HF U154 ( .A0(internal_state_value[47]), .B0(n181), .S(n182), .CO(n183));
Q_AD01HF U155 ( .A0(internal_state_value[48]), .B0(n183), .S(n184), .CO(n185));
Q_AD01HF U156 ( .A0(internal_state_value[49]), .B0(n185), .S(n186), .CO(n187));
Q_AD01HF U157 ( .A0(internal_state_value[50]), .B0(n187), .S(n188), .CO(n189));
Q_AD01HF U158 ( .A0(internal_state_value[51]), .B0(n189), .S(n190), .CO(n191));
Q_AD01HF U159 ( .A0(internal_state_value[52]), .B0(n191), .S(n192), .CO(n193));
Q_AD01HF U160 ( .A0(internal_state_value[53]), .B0(n193), .S(n194), .CO(n195));
Q_AD01HF U161 ( .A0(internal_state_value[54]), .B0(n195), .S(n196), .CO(n197));
Q_AD01HF U162 ( .A0(internal_state_value[55]), .B0(n197), .S(n198), .CO(n199));
Q_AD01HF U163 ( .A0(internal_state_value[56]), .B0(n199), .S(n200), .CO(n201));
Q_AD01HF U164 ( .A0(internal_state_value[57]), .B0(n201), .S(n202), .CO(n203));
Q_AD01HF U165 ( .A0(internal_state_value[58]), .B0(n203), .S(n204), .CO(n205));
Q_AD01HF U166 ( .A0(internal_state_value[59]), .B0(n205), .S(n206), .CO(n207));
Q_AD01HF U167 ( .A0(internal_state_value[60]), .B0(n207), .S(n208), .CO(n209));
Q_AD01HF U168 ( .A0(internal_state_value[61]), .B0(n209), .S(n210), .CO(n211));
Q_AD01HF U169 ( .A0(internal_state_value[62]), .B0(n211), .S(n212), .CO(n213));
Q_AD01HF U170 ( .A0(internal_state_value[63]), .B0(n213), .S(n214), .CO(n215));
Q_AD01HF U171 ( .A0(internal_state_value[64]), .B0(n215), .S(n216), .CO(n217));
Q_AD01HF U172 ( .A0(internal_state_value[65]), .B0(n217), .S(n218), .CO(n219));
Q_AD01HF U173 ( .A0(internal_state_value[66]), .B0(n219), .S(n220), .CO(n221));
Q_AD01HF U174 ( .A0(internal_state_value[67]), .B0(n221), .S(n222), .CO(n223));
Q_AD01HF U175 ( .A0(internal_state_value[68]), .B0(n223), .S(n224), .CO(n225));
Q_AD01HF U176 ( .A0(internal_state_value[69]), .B0(n225), .S(n226), .CO(n227));
Q_AD01HF U177 ( .A0(internal_state_value[70]), .B0(n227), .S(n228), .CO(n229));
Q_AD01HF U178 ( .A0(internal_state_value[71]), .B0(n229), .S(n230), .CO(n231));
Q_AD01HF U179 ( .A0(internal_state_value[72]), .B0(n231), .S(n232), .CO(n233));
Q_AD01HF U180 ( .A0(internal_state_value[73]), .B0(n233), .S(n234), .CO(n235));
Q_AD01HF U181 ( .A0(internal_state_value[74]), .B0(n235), .S(n236), .CO(n237));
Q_AD01HF U182 ( .A0(internal_state_value[75]), .B0(n237), .S(n238), .CO(n239));
Q_AD01HF U183 ( .A0(internal_state_value[76]), .B0(n239), .S(n240), .CO(n241));
Q_AD01HF U184 ( .A0(internal_state_value[77]), .B0(n241), .S(n242), .CO(n243));
Q_AD01HF U185 ( .A0(internal_state_value[78]), .B0(n243), .S(n244), .CO(n245));
Q_AD01HF U186 ( .A0(internal_state_value[79]), .B0(n245), .S(n246), .CO(n247));
Q_AD01HF U187 ( .A0(internal_state_value[80]), .B0(n247), .S(n248), .CO(n249));
Q_AD01HF U188 ( .A0(internal_state_value[81]), .B0(n249), .S(n250), .CO(n251));
Q_AD01HF U189 ( .A0(internal_state_value[82]), .B0(n251), .S(n252), .CO(n253));
Q_AD01HF U190 ( .A0(internal_state_value[83]), .B0(n253), .S(n254), .CO(n255));
Q_AD01HF U191 ( .A0(internal_state_value[84]), .B0(n255), .S(n256), .CO(n257));
Q_AD01HF U192 ( .A0(internal_state_value[85]), .B0(n257), .S(n258), .CO(n259));
Q_AD01HF U193 ( .A0(internal_state_value[86]), .B0(n259), .S(n260), .CO(n261));
Q_AD01HF U194 ( .A0(internal_state_value[87]), .B0(n261), .S(n262), .CO(n263));
Q_AD01HF U195 ( .A0(internal_state_value[88]), .B0(n263), .S(n264), .CO(n265));
Q_AD01HF U196 ( .A0(internal_state_value[89]), .B0(n265), .S(n266), .CO(n267));
Q_AD01HF U197 ( .A0(internal_state_value[90]), .B0(n267), .S(n268), .CO(n269));
Q_AD01HF U198 ( .A0(internal_state_value[91]), .B0(n269), .S(n270), .CO(n271));
Q_AD01HF U199 ( .A0(internal_state_value[92]), .B0(n271), .S(n272), .CO(n273));
Q_AD01HF U200 ( .A0(internal_state_value[93]), .B0(n273), .S(n274), .CO(n275));
Q_AD01HF U201 ( .A0(internal_state_value[94]), .B0(n275), .S(n276), .CO(n277));
Q_AD01HF U202 ( .A0(internal_state_value[95]), .B0(n277), .S(n278), .CO(n279));
Q_AD01HF U203 ( .A0(internal_state_value[96]), .B0(n279), .S(n280), .CO(n281));
Q_AD01HF U204 ( .A0(internal_state_value[97]), .B0(n281), .S(n282), .CO(n283));
Q_AD01HF U205 ( .A0(internal_state_value[98]), .B0(n283), .S(n284), .CO(n285));
Q_AD01HF U206 ( .A0(internal_state_value[99]), .B0(n285), .S(n286), .CO(n287));
Q_AD01HF U207 ( .A0(internal_state_value[100]), .B0(n287), .S(n288), .CO(n289));
Q_AD01HF U208 ( .A0(internal_state_value[101]), .B0(n289), .S(n290), .CO(n291));
Q_AD01HF U209 ( .A0(internal_state_value[102]), .B0(n291), .S(n292), .CO(n293));
Q_AD01HF U210 ( .A0(internal_state_value[103]), .B0(n293), .S(n294), .CO(n295));
Q_AD01HF U211 ( .A0(internal_state_value[104]), .B0(n295), .S(n296), .CO(n297));
Q_AD01HF U212 ( .A0(internal_state_value[105]), .B0(n297), .S(n298), .CO(n299));
Q_AD01HF U213 ( .A0(internal_state_value[106]), .B0(n299), .S(n300), .CO(n301));
Q_AD01HF U214 ( .A0(internal_state_value[107]), .B0(n301), .S(n302), .CO(n303));
Q_AD01HF U215 ( .A0(internal_state_value[108]), .B0(n303), .S(n304), .CO(n305));
Q_AD01HF U216 ( .A0(internal_state_value[109]), .B0(n305), .S(n306), .CO(n307));
Q_AD01HF U217 ( .A0(internal_state_value[110]), .B0(n307), .S(n308), .CO(n309));
Q_AD01HF U218 ( .A0(internal_state_value[111]), .B0(n309), .S(n310), .CO(n311));
Q_AD01HF U219 ( .A0(internal_state_value[112]), .B0(n311), .S(n312), .CO(n313));
Q_AD01HF U220 ( .A0(internal_state_value[113]), .B0(n313), .S(n314), .CO(n315));
Q_AD01HF U221 ( .A0(internal_state_value[114]), .B0(n315), .S(n316), .CO(n317));
Q_AD01HF U222 ( .A0(internal_state_value[115]), .B0(n317), .S(n318), .CO(n319));
Q_AD01HF U223 ( .A0(internal_state_value[116]), .B0(n319), .S(n320), .CO(n321));
Q_AD01HF U224 ( .A0(internal_state_value[117]), .B0(n321), .S(n322), .CO(n323));
Q_AD01HF U225 ( .A0(internal_state_value[118]), .B0(n323), .S(n324), .CO(n325));
Q_AD01HF U226 ( .A0(internal_state_value[119]), .B0(n325), .S(n326), .CO(n327));
Q_AD01HF U227 ( .A0(internal_state_value[120]), .B0(n327), .S(n328), .CO(n329));
Q_AD01HF U228 ( .A0(internal_state_value[121]), .B0(n329), .S(n330), .CO(n331));
Q_AD01HF U229 ( .A0(internal_state_value[122]), .B0(n331), .S(n332), .CO(n333));
Q_AD01HF U230 ( .A0(internal_state_value[123]), .B0(n333), .S(n334), .CO(n335));
Q_AD01HF U231 ( .A0(internal_state_value[124]), .B0(n335), .S(n336), .CO(n337));
Q_AD01HF U232 ( .A0(internal_state_value[125]), .B0(n337), .S(n338), .CO(n339));
Q_AD01HF U233 ( .A0(internal_state_value[126]), .B0(n339), .S(n340), .CO(n341));
Q_XOR2 U234 ( .A0(internal_state_value[127]), .A1(n341), .Z(n342));
Q_AN02 U235 ( .A0(fifo_in_valid), .A1(AesCiphOutR[0]), .Z(fifo_in[0]));
Q_AN02 U236 ( .A0(fifo_in_valid), .A1(AesCiphOutR[1]), .Z(fifo_in[1]));
Q_AN02 U237 ( .A0(fifo_in_valid), .A1(AesCiphOutR[2]), .Z(fifo_in[2]));
Q_AN02 U238 ( .A0(fifo_in_valid), .A1(AesCiphOutR[3]), .Z(fifo_in[3]));
Q_AN02 U239 ( .A0(fifo_in_valid), .A1(AesCiphOutR[4]), .Z(fifo_in[4]));
Q_AN02 U240 ( .A0(fifo_in_valid), .A1(AesCiphOutR[5]), .Z(fifo_in[5]));
Q_AN02 U241 ( .A0(fifo_in_valid), .A1(AesCiphOutR[6]), .Z(fifo_in[6]));
Q_AN02 U242 ( .A0(fifo_in_valid), .A1(AesCiphOutR[7]), .Z(fifo_in[7]));
Q_AN02 U243 ( .A0(fifo_in_valid), .A1(AesCiphOutR[8]), .Z(fifo_in[8]));
Q_AN02 U244 ( .A0(fifo_in_valid), .A1(AesCiphOutR[9]), .Z(fifo_in[9]));
Q_AN02 U245 ( .A0(fifo_in_valid), .A1(AesCiphOutR[10]), .Z(fifo_in[10]));
Q_AN02 U246 ( .A0(fifo_in_valid), .A1(AesCiphOutR[11]), .Z(fifo_in[11]));
Q_AN02 U247 ( .A0(fifo_in_valid), .A1(AesCiphOutR[12]), .Z(fifo_in[12]));
Q_AN02 U248 ( .A0(fifo_in_valid), .A1(AesCiphOutR[13]), .Z(fifo_in[13]));
Q_AN02 U249 ( .A0(fifo_in_valid), .A1(AesCiphOutR[14]), .Z(fifo_in[14]));
Q_AN02 U250 ( .A0(fifo_in_valid), .A1(AesCiphOutR[15]), .Z(fifo_in[15]));
Q_AN02 U251 ( .A0(fifo_in_valid), .A1(AesCiphOutR[16]), .Z(fifo_in[16]));
Q_AN02 U252 ( .A0(fifo_in_valid), .A1(AesCiphOutR[17]), .Z(fifo_in[17]));
Q_AN02 U253 ( .A0(fifo_in_valid), .A1(AesCiphOutR[18]), .Z(fifo_in[18]));
Q_AN02 U254 ( .A0(fifo_in_valid), .A1(AesCiphOutR[19]), .Z(fifo_in[19]));
Q_AN02 U255 ( .A0(fifo_in_valid), .A1(AesCiphOutR[20]), .Z(fifo_in[20]));
Q_AN02 U256 ( .A0(fifo_in_valid), .A1(AesCiphOutR[21]), .Z(fifo_in[21]));
Q_AN02 U257 ( .A0(fifo_in_valid), .A1(AesCiphOutR[22]), .Z(fifo_in[22]));
Q_AN02 U258 ( .A0(fifo_in_valid), .A1(AesCiphOutR[23]), .Z(fifo_in[23]));
Q_AN02 U259 ( .A0(fifo_in_valid), .A1(AesCiphOutR[24]), .Z(fifo_in[24]));
Q_AN02 U260 ( .A0(fifo_in_valid), .A1(AesCiphOutR[25]), .Z(fifo_in[25]));
Q_AN02 U261 ( .A0(fifo_in_valid), .A1(AesCiphOutR[26]), .Z(fifo_in[26]));
Q_AN02 U262 ( .A0(fifo_in_valid), .A1(AesCiphOutR[27]), .Z(fifo_in[27]));
Q_AN02 U263 ( .A0(fifo_in_valid), .A1(AesCiphOutR[28]), .Z(fifo_in[28]));
Q_AN02 U264 ( .A0(fifo_in_valid), .A1(AesCiphOutR[29]), .Z(fifo_in[29]));
Q_AN02 U265 ( .A0(fifo_in_valid), .A1(AesCiphOutR[30]), .Z(fifo_in[30]));
Q_AN02 U266 ( .A0(fifo_in_valid), .A1(AesCiphOutR[31]), .Z(fifo_in[31]));
Q_AN02 U267 ( .A0(fifo_in_valid), .A1(AesCiphOutR[32]), .Z(fifo_in[32]));
Q_AN02 U268 ( .A0(fifo_in_valid), .A1(AesCiphOutR[33]), .Z(fifo_in[33]));
Q_AN02 U269 ( .A0(fifo_in_valid), .A1(AesCiphOutR[34]), .Z(fifo_in[34]));
Q_AN02 U270 ( .A0(fifo_in_valid), .A1(AesCiphOutR[35]), .Z(fifo_in[35]));
Q_AN02 U271 ( .A0(fifo_in_valid), .A1(AesCiphOutR[36]), .Z(fifo_in[36]));
Q_AN02 U272 ( .A0(fifo_in_valid), .A1(AesCiphOutR[37]), .Z(fifo_in[37]));
Q_AN02 U273 ( .A0(fifo_in_valid), .A1(AesCiphOutR[38]), .Z(fifo_in[38]));
Q_AN02 U274 ( .A0(fifo_in_valid), .A1(AesCiphOutR[39]), .Z(fifo_in[39]));
Q_AN02 U275 ( .A0(fifo_in_valid), .A1(AesCiphOutR[40]), .Z(fifo_in[40]));
Q_AN02 U276 ( .A0(fifo_in_valid), .A1(AesCiphOutR[41]), .Z(fifo_in[41]));
Q_AN02 U277 ( .A0(fifo_in_valid), .A1(AesCiphOutR[42]), .Z(fifo_in[42]));
Q_AN02 U278 ( .A0(fifo_in_valid), .A1(AesCiphOutR[43]), .Z(fifo_in[43]));
Q_AN02 U279 ( .A0(fifo_in_valid), .A1(AesCiphOutR[44]), .Z(fifo_in[44]));
Q_AN02 U280 ( .A0(fifo_in_valid), .A1(AesCiphOutR[45]), .Z(fifo_in[45]));
Q_AN02 U281 ( .A0(fifo_in_valid), .A1(AesCiphOutR[46]), .Z(fifo_in[46]));
Q_AN02 U282 ( .A0(fifo_in_valid), .A1(AesCiphOutR[47]), .Z(fifo_in[47]));
Q_AN02 U283 ( .A0(fifo_in_valid), .A1(AesCiphOutR[48]), .Z(fifo_in[48]));
Q_AN02 U284 ( .A0(fifo_in_valid), .A1(AesCiphOutR[49]), .Z(fifo_in[49]));
Q_AN02 U285 ( .A0(fifo_in_valid), .A1(AesCiphOutR[50]), .Z(fifo_in[50]));
Q_AN02 U286 ( .A0(fifo_in_valid), .A1(AesCiphOutR[51]), .Z(fifo_in[51]));
Q_AN02 U287 ( .A0(fifo_in_valid), .A1(AesCiphOutR[52]), .Z(fifo_in[52]));
Q_AN02 U288 ( .A0(fifo_in_valid), .A1(AesCiphOutR[53]), .Z(fifo_in[53]));
Q_AN02 U289 ( .A0(fifo_in_valid), .A1(AesCiphOutR[54]), .Z(fifo_in[54]));
Q_AN02 U290 ( .A0(fifo_in_valid), .A1(AesCiphOutR[55]), .Z(fifo_in[55]));
Q_AN02 U291 ( .A0(fifo_in_valid), .A1(AesCiphOutR[56]), .Z(fifo_in[56]));
Q_AN02 U292 ( .A0(fifo_in_valid), .A1(AesCiphOutR[57]), .Z(fifo_in[57]));
Q_AN02 U293 ( .A0(fifo_in_valid), .A1(AesCiphOutR[58]), .Z(fifo_in[58]));
Q_AN02 U294 ( .A0(fifo_in_valid), .A1(AesCiphOutR[59]), .Z(fifo_in[59]));
Q_AN02 U295 ( .A0(fifo_in_valid), .A1(AesCiphOutR[60]), .Z(fifo_in[60]));
Q_AN02 U296 ( .A0(fifo_in_valid), .A1(AesCiphOutR[61]), .Z(fifo_in[61]));
Q_AN02 U297 ( .A0(fifo_in_valid), .A1(AesCiphOutR[62]), .Z(fifo_in[62]));
Q_AN02 U298 ( .A0(fifo_in_valid), .A1(AesCiphOutR[63]), .Z(fifo_in[63]));
Q_AN02 U299 ( .A0(fifo_in_valid), .A1(AesCiphOutR[64]), .Z(fifo_in[64]));
Q_AN02 U300 ( .A0(fifo_in_valid), .A1(AesCiphOutR[65]), .Z(fifo_in[65]));
Q_AN02 U301 ( .A0(fifo_in_valid), .A1(AesCiphOutR[66]), .Z(fifo_in[66]));
Q_AN02 U302 ( .A0(fifo_in_valid), .A1(AesCiphOutR[67]), .Z(fifo_in[67]));
Q_AN02 U303 ( .A0(fifo_in_valid), .A1(AesCiphOutR[68]), .Z(fifo_in[68]));
Q_AN02 U304 ( .A0(fifo_in_valid), .A1(AesCiphOutR[69]), .Z(fifo_in[69]));
Q_AN02 U305 ( .A0(fifo_in_valid), .A1(AesCiphOutR[70]), .Z(fifo_in[70]));
Q_AN02 U306 ( .A0(fifo_in_valid), .A1(AesCiphOutR[71]), .Z(fifo_in[71]));
Q_AN02 U307 ( .A0(fifo_in_valid), .A1(AesCiphOutR[72]), .Z(fifo_in[72]));
Q_AN02 U308 ( .A0(fifo_in_valid), .A1(AesCiphOutR[73]), .Z(fifo_in[73]));
Q_AN02 U309 ( .A0(fifo_in_valid), .A1(AesCiphOutR[74]), .Z(fifo_in[74]));
Q_AN02 U310 ( .A0(fifo_in_valid), .A1(AesCiphOutR[75]), .Z(fifo_in[75]));
Q_AN02 U311 ( .A0(fifo_in_valid), .A1(AesCiphOutR[76]), .Z(fifo_in[76]));
Q_AN02 U312 ( .A0(fifo_in_valid), .A1(AesCiphOutR[77]), .Z(fifo_in[77]));
Q_AN02 U313 ( .A0(fifo_in_valid), .A1(AesCiphOutR[78]), .Z(fifo_in[78]));
Q_AN02 U314 ( .A0(fifo_in_valid), .A1(AesCiphOutR[79]), .Z(fifo_in[79]));
Q_AN02 U315 ( .A0(fifo_in_valid), .A1(AesCiphOutR[80]), .Z(fifo_in[80]));
Q_AN02 U316 ( .A0(fifo_in_valid), .A1(AesCiphOutR[81]), .Z(fifo_in[81]));
Q_AN02 U317 ( .A0(fifo_in_valid), .A1(AesCiphOutR[82]), .Z(fifo_in[82]));
Q_AN02 U318 ( .A0(fifo_in_valid), .A1(AesCiphOutR[83]), .Z(fifo_in[83]));
Q_AN02 U319 ( .A0(fifo_in_valid), .A1(AesCiphOutR[84]), .Z(fifo_in[84]));
Q_AN02 U320 ( .A0(fifo_in_valid), .A1(AesCiphOutR[85]), .Z(fifo_in[85]));
Q_AN02 U321 ( .A0(fifo_in_valid), .A1(AesCiphOutR[86]), .Z(fifo_in[86]));
Q_AN02 U322 ( .A0(fifo_in_valid), .A1(AesCiphOutR[87]), .Z(fifo_in[87]));
Q_AN02 U323 ( .A0(fifo_in_valid), .A1(AesCiphOutR[88]), .Z(fifo_in[88]));
Q_AN02 U324 ( .A0(fifo_in_valid), .A1(AesCiphOutR[89]), .Z(fifo_in[89]));
Q_AN02 U325 ( .A0(fifo_in_valid), .A1(AesCiphOutR[90]), .Z(fifo_in[90]));
Q_AN02 U326 ( .A0(fifo_in_valid), .A1(AesCiphOutR[91]), .Z(fifo_in[91]));
Q_AN02 U327 ( .A0(fifo_in_valid), .A1(AesCiphOutR[92]), .Z(fifo_in[92]));
Q_AN02 U328 ( .A0(fifo_in_valid), .A1(AesCiphOutR[93]), .Z(fifo_in[93]));
Q_AN02 U329 ( .A0(fifo_in_valid), .A1(AesCiphOutR[94]), .Z(fifo_in[94]));
Q_AN02 U330 ( .A0(fifo_in_valid), .A1(AesCiphOutR[95]), .Z(fifo_in[95]));
Q_AN02 U331 ( .A0(fifo_in_valid), .A1(AesCiphOutR[96]), .Z(fifo_in[96]));
Q_AN02 U332 ( .A0(fifo_in_valid), .A1(AesCiphOutR[97]), .Z(fifo_in[97]));
Q_AN02 U333 ( .A0(fifo_in_valid), .A1(AesCiphOutR[98]), .Z(fifo_in[98]));
Q_AN02 U334 ( .A0(fifo_in_valid), .A1(AesCiphOutR[99]), .Z(fifo_in[99]));
Q_AN02 U335 ( .A0(fifo_in_valid), .A1(AesCiphOutR[100]), .Z(fifo_in[100]));
Q_AN02 U336 ( .A0(fifo_in_valid), .A1(AesCiphOutR[101]), .Z(fifo_in[101]));
Q_AN02 U337 ( .A0(fifo_in_valid), .A1(AesCiphOutR[102]), .Z(fifo_in[102]));
Q_AN02 U338 ( .A0(fifo_in_valid), .A1(AesCiphOutR[103]), .Z(fifo_in[103]));
Q_AN02 U339 ( .A0(fifo_in_valid), .A1(AesCiphOutR[104]), .Z(fifo_in[104]));
Q_AN02 U340 ( .A0(fifo_in_valid), .A1(AesCiphOutR[105]), .Z(fifo_in[105]));
Q_AN02 U341 ( .A0(fifo_in_valid), .A1(AesCiphOutR[106]), .Z(fifo_in[106]));
Q_AN02 U342 ( .A0(fifo_in_valid), .A1(AesCiphOutR[107]), .Z(fifo_in[107]));
Q_AN02 U343 ( .A0(fifo_in_valid), .A1(AesCiphOutR[108]), .Z(fifo_in[108]));
Q_AN02 U344 ( .A0(fifo_in_valid), .A1(AesCiphOutR[109]), .Z(fifo_in[109]));
Q_AN02 U345 ( .A0(fifo_in_valid), .A1(AesCiphOutR[110]), .Z(fifo_in[110]));
Q_AN02 U346 ( .A0(fifo_in_valid), .A1(AesCiphOutR[111]), .Z(fifo_in[111]));
Q_AN02 U347 ( .A0(fifo_in_valid), .A1(AesCiphOutR[112]), .Z(fifo_in[112]));
Q_AN02 U348 ( .A0(fifo_in_valid), .A1(AesCiphOutR[113]), .Z(fifo_in[113]));
Q_AN02 U349 ( .A0(fifo_in_valid), .A1(AesCiphOutR[114]), .Z(fifo_in[114]));
Q_AN02 U350 ( .A0(fifo_in_valid), .A1(AesCiphOutR[115]), .Z(fifo_in[115]));
Q_AN02 U351 ( .A0(fifo_in_valid), .A1(AesCiphOutR[116]), .Z(fifo_in[116]));
Q_AN02 U352 ( .A0(fifo_in_valid), .A1(AesCiphOutR[117]), .Z(fifo_in[117]));
Q_AN02 U353 ( .A0(fifo_in_valid), .A1(AesCiphOutR[118]), .Z(fifo_in[118]));
Q_AN02 U354 ( .A0(fifo_in_valid), .A1(AesCiphOutR[119]), .Z(fifo_in[119]));
Q_AN02 U355 ( .A0(fifo_in_valid), .A1(AesCiphOutR[120]), .Z(fifo_in[120]));
Q_AN02 U356 ( .A0(fifo_in_valid), .A1(AesCiphOutR[121]), .Z(fifo_in[121]));
Q_AN02 U357 ( .A0(fifo_in_valid), .A1(AesCiphOutR[122]), .Z(fifo_in[122]));
Q_AN02 U358 ( .A0(fifo_in_valid), .A1(AesCiphOutR[123]), .Z(fifo_in[123]));
Q_AN02 U359 ( .A0(fifo_in_valid), .A1(AesCiphOutR[124]), .Z(fifo_in[124]));
Q_AN02 U360 ( .A0(fifo_in_valid), .A1(AesCiphOutR[125]), .Z(fifo_in[125]));
Q_AN02 U361 ( .A0(fifo_in_valid), .A1(AesCiphOutR[126]), .Z(fifo_in[126]));
Q_AN02 U362 ( .A0(fifo_in_valid), .A1(AesCiphOutR[127]), .Z(fifo_in[127]));
Q_AN02 U363 ( .A0(KeyInVld), .A1(internal_state_key[0]), .Z(KeyIn[0]));
Q_AN02 U364 ( .A0(KeyInVld), .A1(internal_state_key[1]), .Z(KeyIn[1]));
Q_AN02 U365 ( .A0(KeyInVld), .A1(internal_state_key[2]), .Z(KeyIn[2]));
Q_AN02 U366 ( .A0(KeyInVld), .A1(internal_state_key[3]), .Z(KeyIn[3]));
Q_AN02 U367 ( .A0(KeyInVld), .A1(internal_state_key[4]), .Z(KeyIn[4]));
Q_AN02 U368 ( .A0(KeyInVld), .A1(internal_state_key[5]), .Z(KeyIn[5]));
Q_AN02 U369 ( .A0(KeyInVld), .A1(internal_state_key[6]), .Z(KeyIn[6]));
Q_AN02 U370 ( .A0(KeyInVld), .A1(internal_state_key[7]), .Z(KeyIn[7]));
Q_AN02 U371 ( .A0(KeyInVld), .A1(internal_state_key[8]), .Z(KeyIn[8]));
Q_AN02 U372 ( .A0(KeyInVld), .A1(internal_state_key[9]), .Z(KeyIn[9]));
Q_AN02 U373 ( .A0(KeyInVld), .A1(internal_state_key[10]), .Z(KeyIn[10]));
Q_AN02 U374 ( .A0(KeyInVld), .A1(internal_state_key[11]), .Z(KeyIn[11]));
Q_AN02 U375 ( .A0(KeyInVld), .A1(internal_state_key[12]), .Z(KeyIn[12]));
Q_AN02 U376 ( .A0(KeyInVld), .A1(internal_state_key[13]), .Z(KeyIn[13]));
Q_AN02 U377 ( .A0(KeyInVld), .A1(internal_state_key[14]), .Z(KeyIn[14]));
Q_AN02 U378 ( .A0(KeyInVld), .A1(internal_state_key[15]), .Z(KeyIn[15]));
Q_AN02 U379 ( .A0(KeyInVld), .A1(internal_state_key[16]), .Z(KeyIn[16]));
Q_AN02 U380 ( .A0(KeyInVld), .A1(internal_state_key[17]), .Z(KeyIn[17]));
Q_AN02 U381 ( .A0(KeyInVld), .A1(internal_state_key[18]), .Z(KeyIn[18]));
Q_AN02 U382 ( .A0(KeyInVld), .A1(internal_state_key[19]), .Z(KeyIn[19]));
Q_AN02 U383 ( .A0(KeyInVld), .A1(internal_state_key[20]), .Z(KeyIn[20]));
Q_AN02 U384 ( .A0(KeyInVld), .A1(internal_state_key[21]), .Z(KeyIn[21]));
Q_AN02 U385 ( .A0(KeyInVld), .A1(internal_state_key[22]), .Z(KeyIn[22]));
Q_AN02 U386 ( .A0(KeyInVld), .A1(internal_state_key[23]), .Z(KeyIn[23]));
Q_AN02 U387 ( .A0(KeyInVld), .A1(internal_state_key[24]), .Z(KeyIn[24]));
Q_AN02 U388 ( .A0(KeyInVld), .A1(internal_state_key[25]), .Z(KeyIn[25]));
Q_AN02 U389 ( .A0(KeyInVld), .A1(internal_state_key[26]), .Z(KeyIn[26]));
Q_AN02 U390 ( .A0(KeyInVld), .A1(internal_state_key[27]), .Z(KeyIn[27]));
Q_AN02 U391 ( .A0(KeyInVld), .A1(internal_state_key[28]), .Z(KeyIn[28]));
Q_AN02 U392 ( .A0(KeyInVld), .A1(internal_state_key[29]), .Z(KeyIn[29]));
Q_AN02 U393 ( .A0(KeyInVld), .A1(internal_state_key[30]), .Z(KeyIn[30]));
Q_AN02 U394 ( .A0(KeyInVld), .A1(internal_state_key[31]), .Z(KeyIn[31]));
Q_AN02 U395 ( .A0(KeyInVld), .A1(internal_state_key[32]), .Z(KeyIn[32]));
Q_AN02 U396 ( .A0(KeyInVld), .A1(internal_state_key[33]), .Z(KeyIn[33]));
Q_AN02 U397 ( .A0(KeyInVld), .A1(internal_state_key[34]), .Z(KeyIn[34]));
Q_AN02 U398 ( .A0(KeyInVld), .A1(internal_state_key[35]), .Z(KeyIn[35]));
Q_AN02 U399 ( .A0(KeyInVld), .A1(internal_state_key[36]), .Z(KeyIn[36]));
Q_AN02 U400 ( .A0(KeyInVld), .A1(internal_state_key[37]), .Z(KeyIn[37]));
Q_AN02 U401 ( .A0(KeyInVld), .A1(internal_state_key[38]), .Z(KeyIn[38]));
Q_AN02 U402 ( .A0(KeyInVld), .A1(internal_state_key[39]), .Z(KeyIn[39]));
Q_AN02 U403 ( .A0(KeyInVld), .A1(internal_state_key[40]), .Z(KeyIn[40]));
Q_AN02 U404 ( .A0(KeyInVld), .A1(internal_state_key[41]), .Z(KeyIn[41]));
Q_AN02 U405 ( .A0(KeyInVld), .A1(internal_state_key[42]), .Z(KeyIn[42]));
Q_AN02 U406 ( .A0(KeyInVld), .A1(internal_state_key[43]), .Z(KeyIn[43]));
Q_AN02 U407 ( .A0(KeyInVld), .A1(internal_state_key[44]), .Z(KeyIn[44]));
Q_AN02 U408 ( .A0(KeyInVld), .A1(internal_state_key[45]), .Z(KeyIn[45]));
Q_AN02 U409 ( .A0(KeyInVld), .A1(internal_state_key[46]), .Z(KeyIn[46]));
Q_AN02 U410 ( .A0(KeyInVld), .A1(internal_state_key[47]), .Z(KeyIn[47]));
Q_AN02 U411 ( .A0(KeyInVld), .A1(internal_state_key[48]), .Z(KeyIn[48]));
Q_AN02 U412 ( .A0(KeyInVld), .A1(internal_state_key[49]), .Z(KeyIn[49]));
Q_AN02 U413 ( .A0(KeyInVld), .A1(internal_state_key[50]), .Z(KeyIn[50]));
Q_AN02 U414 ( .A0(KeyInVld), .A1(internal_state_key[51]), .Z(KeyIn[51]));
Q_AN02 U415 ( .A0(KeyInVld), .A1(internal_state_key[52]), .Z(KeyIn[52]));
Q_AN02 U416 ( .A0(KeyInVld), .A1(internal_state_key[53]), .Z(KeyIn[53]));
Q_AN02 U417 ( .A0(KeyInVld), .A1(internal_state_key[54]), .Z(KeyIn[54]));
Q_AN02 U418 ( .A0(KeyInVld), .A1(internal_state_key[55]), .Z(KeyIn[55]));
Q_AN02 U419 ( .A0(KeyInVld), .A1(internal_state_key[56]), .Z(KeyIn[56]));
Q_AN02 U420 ( .A0(KeyInVld), .A1(internal_state_key[57]), .Z(KeyIn[57]));
Q_AN02 U421 ( .A0(KeyInVld), .A1(internal_state_key[58]), .Z(KeyIn[58]));
Q_AN02 U422 ( .A0(KeyInVld), .A1(internal_state_key[59]), .Z(KeyIn[59]));
Q_AN02 U423 ( .A0(KeyInVld), .A1(internal_state_key[60]), .Z(KeyIn[60]));
Q_AN02 U424 ( .A0(KeyInVld), .A1(internal_state_key[61]), .Z(KeyIn[61]));
Q_AN02 U425 ( .A0(KeyInVld), .A1(internal_state_key[62]), .Z(KeyIn[62]));
Q_AN02 U426 ( .A0(KeyInVld), .A1(internal_state_key[63]), .Z(KeyIn[63]));
Q_AN02 U427 ( .A0(KeyInVld), .A1(internal_state_key[64]), .Z(KeyIn[64]));
Q_AN02 U428 ( .A0(KeyInVld), .A1(internal_state_key[65]), .Z(KeyIn[65]));
Q_AN02 U429 ( .A0(KeyInVld), .A1(internal_state_key[66]), .Z(KeyIn[66]));
Q_AN02 U430 ( .A0(KeyInVld), .A1(internal_state_key[67]), .Z(KeyIn[67]));
Q_AN02 U431 ( .A0(KeyInVld), .A1(internal_state_key[68]), .Z(KeyIn[68]));
Q_AN02 U432 ( .A0(KeyInVld), .A1(internal_state_key[69]), .Z(KeyIn[69]));
Q_AN02 U433 ( .A0(KeyInVld), .A1(internal_state_key[70]), .Z(KeyIn[70]));
Q_AN02 U434 ( .A0(KeyInVld), .A1(internal_state_key[71]), .Z(KeyIn[71]));
Q_AN02 U435 ( .A0(KeyInVld), .A1(internal_state_key[72]), .Z(KeyIn[72]));
Q_AN02 U436 ( .A0(KeyInVld), .A1(internal_state_key[73]), .Z(KeyIn[73]));
Q_AN02 U437 ( .A0(KeyInVld), .A1(internal_state_key[74]), .Z(KeyIn[74]));
Q_AN02 U438 ( .A0(KeyInVld), .A1(internal_state_key[75]), .Z(KeyIn[75]));
Q_AN02 U439 ( .A0(KeyInVld), .A1(internal_state_key[76]), .Z(KeyIn[76]));
Q_AN02 U440 ( .A0(KeyInVld), .A1(internal_state_key[77]), .Z(KeyIn[77]));
Q_AN02 U441 ( .A0(KeyInVld), .A1(internal_state_key[78]), .Z(KeyIn[78]));
Q_AN02 U442 ( .A0(KeyInVld), .A1(internal_state_key[79]), .Z(KeyIn[79]));
Q_AN02 U443 ( .A0(KeyInVld), .A1(internal_state_key[80]), .Z(KeyIn[80]));
Q_AN02 U444 ( .A0(KeyInVld), .A1(internal_state_key[81]), .Z(KeyIn[81]));
Q_AN02 U445 ( .A0(KeyInVld), .A1(internal_state_key[82]), .Z(KeyIn[82]));
Q_AN02 U446 ( .A0(KeyInVld), .A1(internal_state_key[83]), .Z(KeyIn[83]));
Q_AN02 U447 ( .A0(KeyInVld), .A1(internal_state_key[84]), .Z(KeyIn[84]));
Q_AN02 U448 ( .A0(KeyInVld), .A1(internal_state_key[85]), .Z(KeyIn[85]));
Q_AN02 U449 ( .A0(KeyInVld), .A1(internal_state_key[86]), .Z(KeyIn[86]));
Q_AN02 U450 ( .A0(KeyInVld), .A1(internal_state_key[87]), .Z(KeyIn[87]));
Q_AN02 U451 ( .A0(KeyInVld), .A1(internal_state_key[88]), .Z(KeyIn[88]));
Q_AN02 U452 ( .A0(KeyInVld), .A1(internal_state_key[89]), .Z(KeyIn[89]));
Q_AN02 U453 ( .A0(KeyInVld), .A1(internal_state_key[90]), .Z(KeyIn[90]));
Q_AN02 U454 ( .A0(KeyInVld), .A1(internal_state_key[91]), .Z(KeyIn[91]));
Q_AN02 U455 ( .A0(KeyInVld), .A1(internal_state_key[92]), .Z(KeyIn[92]));
Q_AN02 U456 ( .A0(KeyInVld), .A1(internal_state_key[93]), .Z(KeyIn[93]));
Q_AN02 U457 ( .A0(KeyInVld), .A1(internal_state_key[94]), .Z(KeyIn[94]));
Q_AN02 U458 ( .A0(KeyInVld), .A1(internal_state_key[95]), .Z(KeyIn[95]));
Q_AN02 U459 ( .A0(KeyInVld), .A1(internal_state_key[96]), .Z(KeyIn[96]));
Q_AN02 U460 ( .A0(KeyInVld), .A1(internal_state_key[97]), .Z(KeyIn[97]));
Q_AN02 U461 ( .A0(KeyInVld), .A1(internal_state_key[98]), .Z(KeyIn[98]));
Q_AN02 U462 ( .A0(KeyInVld), .A1(internal_state_key[99]), .Z(KeyIn[99]));
Q_AN02 U463 ( .A0(KeyInVld), .A1(internal_state_key[100]), .Z(KeyIn[100]));
Q_AN02 U464 ( .A0(KeyInVld), .A1(internal_state_key[101]), .Z(KeyIn[101]));
Q_AN02 U465 ( .A0(KeyInVld), .A1(internal_state_key[102]), .Z(KeyIn[102]));
Q_AN02 U466 ( .A0(KeyInVld), .A1(internal_state_key[103]), .Z(KeyIn[103]));
Q_AN02 U467 ( .A0(KeyInVld), .A1(internal_state_key[104]), .Z(KeyIn[104]));
Q_AN02 U468 ( .A0(KeyInVld), .A1(internal_state_key[105]), .Z(KeyIn[105]));
Q_AN02 U469 ( .A0(KeyInVld), .A1(internal_state_key[106]), .Z(KeyIn[106]));
Q_AN02 U470 ( .A0(KeyInVld), .A1(internal_state_key[107]), .Z(KeyIn[107]));
Q_AN02 U471 ( .A0(KeyInVld), .A1(internal_state_key[108]), .Z(KeyIn[108]));
Q_AN02 U472 ( .A0(KeyInVld), .A1(internal_state_key[109]), .Z(KeyIn[109]));
Q_AN02 U473 ( .A0(KeyInVld), .A1(internal_state_key[110]), .Z(KeyIn[110]));
Q_AN02 U474 ( .A0(KeyInVld), .A1(internal_state_key[111]), .Z(KeyIn[111]));
Q_AN02 U475 ( .A0(KeyInVld), .A1(internal_state_key[112]), .Z(KeyIn[112]));
Q_AN02 U476 ( .A0(KeyInVld), .A1(internal_state_key[113]), .Z(KeyIn[113]));
Q_AN02 U477 ( .A0(KeyInVld), .A1(internal_state_key[114]), .Z(KeyIn[114]));
Q_AN02 U478 ( .A0(KeyInVld), .A1(internal_state_key[115]), .Z(KeyIn[115]));
Q_AN02 U479 ( .A0(KeyInVld), .A1(internal_state_key[116]), .Z(KeyIn[116]));
Q_AN02 U480 ( .A0(KeyInVld), .A1(internal_state_key[117]), .Z(KeyIn[117]));
Q_AN02 U481 ( .A0(KeyInVld), .A1(internal_state_key[118]), .Z(KeyIn[118]));
Q_AN02 U482 ( .A0(KeyInVld), .A1(internal_state_key[119]), .Z(KeyIn[119]));
Q_AN02 U483 ( .A0(KeyInVld), .A1(internal_state_key[120]), .Z(KeyIn[120]));
Q_AN02 U484 ( .A0(KeyInVld), .A1(internal_state_key[121]), .Z(KeyIn[121]));
Q_AN02 U485 ( .A0(KeyInVld), .A1(internal_state_key[122]), .Z(KeyIn[122]));
Q_AN02 U486 ( .A0(KeyInVld), .A1(internal_state_key[123]), .Z(KeyIn[123]));
Q_AN02 U487 ( .A0(KeyInVld), .A1(internal_state_key[124]), .Z(KeyIn[124]));
Q_AN02 U488 ( .A0(KeyInVld), .A1(internal_state_key[125]), .Z(KeyIn[125]));
Q_AN02 U489 ( .A0(KeyInVld), .A1(internal_state_key[126]), .Z(KeyIn[126]));
Q_AN02 U490 ( .A0(KeyInVld), .A1(internal_state_key[127]), .Z(KeyIn[127]));
Q_AN02 U491 ( .A0(KeyInVld), .A1(internal_state_key[128]), .Z(KeyIn[128]));
Q_AN02 U492 ( .A0(KeyInVld), .A1(internal_state_key[129]), .Z(KeyIn[129]));
Q_AN02 U493 ( .A0(KeyInVld), .A1(internal_state_key[130]), .Z(KeyIn[130]));
Q_AN02 U494 ( .A0(KeyInVld), .A1(internal_state_key[131]), .Z(KeyIn[131]));
Q_AN02 U495 ( .A0(KeyInVld), .A1(internal_state_key[132]), .Z(KeyIn[132]));
Q_AN02 U496 ( .A0(KeyInVld), .A1(internal_state_key[133]), .Z(KeyIn[133]));
Q_AN02 U497 ( .A0(KeyInVld), .A1(internal_state_key[134]), .Z(KeyIn[134]));
Q_AN02 U498 ( .A0(KeyInVld), .A1(internal_state_key[135]), .Z(KeyIn[135]));
Q_AN02 U499 ( .A0(KeyInVld), .A1(internal_state_key[136]), .Z(KeyIn[136]));
Q_AN02 U500 ( .A0(KeyInVld), .A1(internal_state_key[137]), .Z(KeyIn[137]));
Q_AN02 U501 ( .A0(KeyInVld), .A1(internal_state_key[138]), .Z(KeyIn[138]));
Q_AN02 U502 ( .A0(KeyInVld), .A1(internal_state_key[139]), .Z(KeyIn[139]));
Q_AN02 U503 ( .A0(KeyInVld), .A1(internal_state_key[140]), .Z(KeyIn[140]));
Q_AN02 U504 ( .A0(KeyInVld), .A1(internal_state_key[141]), .Z(KeyIn[141]));
Q_AN02 U505 ( .A0(KeyInVld), .A1(internal_state_key[142]), .Z(KeyIn[142]));
Q_AN02 U506 ( .A0(KeyInVld), .A1(internal_state_key[143]), .Z(KeyIn[143]));
Q_AN02 U507 ( .A0(KeyInVld), .A1(internal_state_key[144]), .Z(KeyIn[144]));
Q_AN02 U508 ( .A0(KeyInVld), .A1(internal_state_key[145]), .Z(KeyIn[145]));
Q_AN02 U509 ( .A0(KeyInVld), .A1(internal_state_key[146]), .Z(KeyIn[146]));
Q_AN02 U510 ( .A0(KeyInVld), .A1(internal_state_key[147]), .Z(KeyIn[147]));
Q_AN02 U511 ( .A0(KeyInVld), .A1(internal_state_key[148]), .Z(KeyIn[148]));
Q_AN02 U512 ( .A0(KeyInVld), .A1(internal_state_key[149]), .Z(KeyIn[149]));
Q_AN02 U513 ( .A0(KeyInVld), .A1(internal_state_key[150]), .Z(KeyIn[150]));
Q_AN02 U514 ( .A0(KeyInVld), .A1(internal_state_key[151]), .Z(KeyIn[151]));
Q_AN02 U515 ( .A0(KeyInVld), .A1(internal_state_key[152]), .Z(KeyIn[152]));
Q_AN02 U516 ( .A0(KeyInVld), .A1(internal_state_key[153]), .Z(KeyIn[153]));
Q_AN02 U517 ( .A0(KeyInVld), .A1(internal_state_key[154]), .Z(KeyIn[154]));
Q_AN02 U518 ( .A0(KeyInVld), .A1(internal_state_key[155]), .Z(KeyIn[155]));
Q_AN02 U519 ( .A0(KeyInVld), .A1(internal_state_key[156]), .Z(KeyIn[156]));
Q_AN02 U520 ( .A0(KeyInVld), .A1(internal_state_key[157]), .Z(KeyIn[157]));
Q_AN02 U521 ( .A0(KeyInVld), .A1(internal_state_key[158]), .Z(KeyIn[158]));
Q_AN02 U522 ( .A0(KeyInVld), .A1(internal_state_key[159]), .Z(KeyIn[159]));
Q_AN02 U523 ( .A0(KeyInVld), .A1(internal_state_key[160]), .Z(KeyIn[160]));
Q_AN02 U524 ( .A0(KeyInVld), .A1(internal_state_key[161]), .Z(KeyIn[161]));
Q_AN02 U525 ( .A0(KeyInVld), .A1(internal_state_key[162]), .Z(KeyIn[162]));
Q_AN02 U526 ( .A0(KeyInVld), .A1(internal_state_key[163]), .Z(KeyIn[163]));
Q_AN02 U527 ( .A0(KeyInVld), .A1(internal_state_key[164]), .Z(KeyIn[164]));
Q_AN02 U528 ( .A0(KeyInVld), .A1(internal_state_key[165]), .Z(KeyIn[165]));
Q_AN02 U529 ( .A0(KeyInVld), .A1(internal_state_key[166]), .Z(KeyIn[166]));
Q_AN02 U530 ( .A0(KeyInVld), .A1(internal_state_key[167]), .Z(KeyIn[167]));
Q_AN02 U531 ( .A0(KeyInVld), .A1(internal_state_key[168]), .Z(KeyIn[168]));
Q_AN02 U532 ( .A0(KeyInVld), .A1(internal_state_key[169]), .Z(KeyIn[169]));
Q_AN02 U533 ( .A0(KeyInVld), .A1(internal_state_key[170]), .Z(KeyIn[170]));
Q_AN02 U534 ( .A0(KeyInVld), .A1(internal_state_key[171]), .Z(KeyIn[171]));
Q_AN02 U535 ( .A0(KeyInVld), .A1(internal_state_key[172]), .Z(KeyIn[172]));
Q_AN02 U536 ( .A0(KeyInVld), .A1(internal_state_key[173]), .Z(KeyIn[173]));
Q_AN02 U537 ( .A0(KeyInVld), .A1(internal_state_key[174]), .Z(KeyIn[174]));
Q_AN02 U538 ( .A0(KeyInVld), .A1(internal_state_key[175]), .Z(KeyIn[175]));
Q_AN02 U539 ( .A0(KeyInVld), .A1(internal_state_key[176]), .Z(KeyIn[176]));
Q_AN02 U540 ( .A0(KeyInVld), .A1(internal_state_key[177]), .Z(KeyIn[177]));
Q_AN02 U541 ( .A0(KeyInVld), .A1(internal_state_key[178]), .Z(KeyIn[178]));
Q_AN02 U542 ( .A0(KeyInVld), .A1(internal_state_key[179]), .Z(KeyIn[179]));
Q_AN02 U543 ( .A0(KeyInVld), .A1(internal_state_key[180]), .Z(KeyIn[180]));
Q_AN02 U544 ( .A0(KeyInVld), .A1(internal_state_key[181]), .Z(KeyIn[181]));
Q_AN02 U545 ( .A0(KeyInVld), .A1(internal_state_key[182]), .Z(KeyIn[182]));
Q_AN02 U546 ( .A0(KeyInVld), .A1(internal_state_key[183]), .Z(KeyIn[183]));
Q_AN02 U547 ( .A0(KeyInVld), .A1(internal_state_key[184]), .Z(KeyIn[184]));
Q_AN02 U548 ( .A0(KeyInVld), .A1(internal_state_key[185]), .Z(KeyIn[185]));
Q_AN02 U549 ( .A0(KeyInVld), .A1(internal_state_key[186]), .Z(KeyIn[186]));
Q_AN02 U550 ( .A0(KeyInVld), .A1(internal_state_key[187]), .Z(KeyIn[187]));
Q_AN02 U551 ( .A0(KeyInVld), .A1(internal_state_key[188]), .Z(KeyIn[188]));
Q_AN02 U552 ( .A0(KeyInVld), .A1(internal_state_key[189]), .Z(KeyIn[189]));
Q_AN02 U553 ( .A0(KeyInVld), .A1(internal_state_key[190]), .Z(KeyIn[190]));
Q_AN02 U554 ( .A0(KeyInVld), .A1(internal_state_key[191]), .Z(KeyIn[191]));
Q_AN02 U555 ( .A0(KeyInVld), .A1(internal_state_key[192]), .Z(KeyIn[192]));
Q_AN02 U556 ( .A0(KeyInVld), .A1(internal_state_key[193]), .Z(KeyIn[193]));
Q_AN02 U557 ( .A0(KeyInVld), .A1(internal_state_key[194]), .Z(KeyIn[194]));
Q_AN02 U558 ( .A0(KeyInVld), .A1(internal_state_key[195]), .Z(KeyIn[195]));
Q_AN02 U559 ( .A0(KeyInVld), .A1(internal_state_key[196]), .Z(KeyIn[196]));
Q_AN02 U560 ( .A0(KeyInVld), .A1(internal_state_key[197]), .Z(KeyIn[197]));
Q_AN02 U561 ( .A0(KeyInVld), .A1(internal_state_key[198]), .Z(KeyIn[198]));
Q_AN02 U562 ( .A0(KeyInVld), .A1(internal_state_key[199]), .Z(KeyIn[199]));
Q_AN02 U563 ( .A0(KeyInVld), .A1(internal_state_key[200]), .Z(KeyIn[200]));
Q_AN02 U564 ( .A0(KeyInVld), .A1(internal_state_key[201]), .Z(KeyIn[201]));
Q_AN02 U565 ( .A0(KeyInVld), .A1(internal_state_key[202]), .Z(KeyIn[202]));
Q_AN02 U566 ( .A0(KeyInVld), .A1(internal_state_key[203]), .Z(KeyIn[203]));
Q_AN02 U567 ( .A0(KeyInVld), .A1(internal_state_key[204]), .Z(KeyIn[204]));
Q_AN02 U568 ( .A0(KeyInVld), .A1(internal_state_key[205]), .Z(KeyIn[205]));
Q_AN02 U569 ( .A0(KeyInVld), .A1(internal_state_key[206]), .Z(KeyIn[206]));
Q_AN02 U570 ( .A0(KeyInVld), .A1(internal_state_key[207]), .Z(KeyIn[207]));
Q_AN02 U571 ( .A0(KeyInVld), .A1(internal_state_key[208]), .Z(KeyIn[208]));
Q_AN02 U572 ( .A0(KeyInVld), .A1(internal_state_key[209]), .Z(KeyIn[209]));
Q_AN02 U573 ( .A0(KeyInVld), .A1(internal_state_key[210]), .Z(KeyIn[210]));
Q_AN02 U574 ( .A0(KeyInVld), .A1(internal_state_key[211]), .Z(KeyIn[211]));
Q_AN02 U575 ( .A0(KeyInVld), .A1(internal_state_key[212]), .Z(KeyIn[212]));
Q_AN02 U576 ( .A0(KeyInVld), .A1(internal_state_key[213]), .Z(KeyIn[213]));
Q_AN02 U577 ( .A0(KeyInVld), .A1(internal_state_key[214]), .Z(KeyIn[214]));
Q_AN02 U578 ( .A0(KeyInVld), .A1(internal_state_key[215]), .Z(KeyIn[215]));
Q_AN02 U579 ( .A0(KeyInVld), .A1(internal_state_key[216]), .Z(KeyIn[216]));
Q_AN02 U580 ( .A0(KeyInVld), .A1(internal_state_key[217]), .Z(KeyIn[217]));
Q_AN02 U581 ( .A0(KeyInVld), .A1(internal_state_key[218]), .Z(KeyIn[218]));
Q_AN02 U582 ( .A0(KeyInVld), .A1(internal_state_key[219]), .Z(KeyIn[219]));
Q_AN02 U583 ( .A0(KeyInVld), .A1(internal_state_key[220]), .Z(KeyIn[220]));
Q_AN02 U584 ( .A0(KeyInVld), .A1(internal_state_key[221]), .Z(KeyIn[221]));
Q_AN02 U585 ( .A0(KeyInVld), .A1(internal_state_key[222]), .Z(KeyIn[222]));
Q_AN02 U586 ( .A0(KeyInVld), .A1(internal_state_key[223]), .Z(KeyIn[223]));
Q_AN02 U587 ( .A0(KeyInVld), .A1(internal_state_key[224]), .Z(KeyIn[224]));
Q_AN02 U588 ( .A0(KeyInVld), .A1(internal_state_key[225]), .Z(KeyIn[225]));
Q_AN02 U589 ( .A0(KeyInVld), .A1(internal_state_key[226]), .Z(KeyIn[226]));
Q_AN02 U590 ( .A0(KeyInVld), .A1(internal_state_key[227]), .Z(KeyIn[227]));
Q_AN02 U591 ( .A0(KeyInVld), .A1(internal_state_key[228]), .Z(KeyIn[228]));
Q_AN02 U592 ( .A0(KeyInVld), .A1(internal_state_key[229]), .Z(KeyIn[229]));
Q_AN02 U593 ( .A0(KeyInVld), .A1(internal_state_key[230]), .Z(KeyIn[230]));
Q_AN02 U594 ( .A0(KeyInVld), .A1(internal_state_key[231]), .Z(KeyIn[231]));
Q_AN02 U595 ( .A0(KeyInVld), .A1(internal_state_key[232]), .Z(KeyIn[232]));
Q_AN02 U596 ( .A0(KeyInVld), .A1(internal_state_key[233]), .Z(KeyIn[233]));
Q_AN02 U597 ( .A0(KeyInVld), .A1(internal_state_key[234]), .Z(KeyIn[234]));
Q_AN02 U598 ( .A0(KeyInVld), .A1(internal_state_key[235]), .Z(KeyIn[235]));
Q_AN02 U599 ( .A0(KeyInVld), .A1(internal_state_key[236]), .Z(KeyIn[236]));
Q_AN02 U600 ( .A0(KeyInVld), .A1(internal_state_key[237]), .Z(KeyIn[237]));
Q_AN02 U601 ( .A0(KeyInVld), .A1(internal_state_key[238]), .Z(KeyIn[238]));
Q_AN02 U602 ( .A0(KeyInVld), .A1(internal_state_key[239]), .Z(KeyIn[239]));
Q_AN02 U603 ( .A0(KeyInVld), .A1(internal_state_key[240]), .Z(KeyIn[240]));
Q_AN02 U604 ( .A0(KeyInVld), .A1(internal_state_key[241]), .Z(KeyIn[241]));
Q_AN02 U605 ( .A0(KeyInVld), .A1(internal_state_key[242]), .Z(KeyIn[242]));
Q_AN02 U606 ( .A0(KeyInVld), .A1(internal_state_key[243]), .Z(KeyIn[243]));
Q_AN02 U607 ( .A0(KeyInVld), .A1(internal_state_key[244]), .Z(KeyIn[244]));
Q_AN02 U608 ( .A0(KeyInVld), .A1(internal_state_key[245]), .Z(KeyIn[245]));
Q_AN02 U609 ( .A0(KeyInVld), .A1(internal_state_key[246]), .Z(KeyIn[246]));
Q_AN02 U610 ( .A0(KeyInVld), .A1(internal_state_key[247]), .Z(KeyIn[247]));
Q_AN02 U611 ( .A0(KeyInVld), .A1(internal_state_key[248]), .Z(KeyIn[248]));
Q_AN02 U612 ( .A0(KeyInVld), .A1(internal_state_key[249]), .Z(KeyIn[249]));
Q_AN02 U613 ( .A0(KeyInVld), .A1(internal_state_key[250]), .Z(KeyIn[250]));
Q_AN02 U614 ( .A0(KeyInVld), .A1(internal_state_key[251]), .Z(KeyIn[251]));
Q_AN02 U615 ( .A0(KeyInVld), .A1(internal_state_key[252]), .Z(KeyIn[252]));
Q_AN02 U616 ( .A0(KeyInVld), .A1(internal_state_key[253]), .Z(KeyIn[253]));
Q_AN02 U617 ( .A0(KeyInVld), .A1(internal_state_key[254]), .Z(KeyIn[254]));
Q_AN02 U618 ( .A0(KeyInVld), .A1(internal_state_key[255]), .Z(KeyIn[255]));
Q_AN02 U619 ( .A0(CiphInVldR), .A1(n89), .Z(CiphIn[0]));
Q_AN02 U620 ( .A0(CiphInVldR), .A1(n91), .Z(CiphIn[1]));
Q_AN02 U621 ( .A0(CiphInVldR), .A1(n92), .Z(CiphIn[2]));
Q_AN02 U622 ( .A0(CiphInVldR), .A1(n94), .Z(CiphIn[3]));
Q_AN02 U623 ( .A0(CiphInVldR), .A1(n96), .Z(CiphIn[4]));
Q_AN02 U624 ( .A0(CiphInVldR), .A1(n98), .Z(CiphIn[5]));
Q_AN02 U625 ( .A0(CiphInVldR), .A1(n100), .Z(CiphIn[6]));
Q_AN02 U626 ( .A0(CiphInVldR), .A1(n102), .Z(CiphIn[7]));
Q_AN02 U627 ( .A0(CiphInVldR), .A1(n104), .Z(CiphIn[8]));
Q_AN02 U628 ( .A0(CiphInVldR), .A1(n106), .Z(CiphIn[9]));
Q_AN02 U629 ( .A0(CiphInVldR), .A1(n108), .Z(CiphIn[10]));
Q_AN02 U630 ( .A0(CiphInVldR), .A1(n110), .Z(CiphIn[11]));
Q_AN02 U631 ( .A0(CiphInVldR), .A1(n112), .Z(CiphIn[12]));
Q_AN02 U632 ( .A0(CiphInVldR), .A1(n114), .Z(CiphIn[13]));
Q_AN02 U633 ( .A0(CiphInVldR), .A1(n116), .Z(CiphIn[14]));
Q_AN02 U634 ( .A0(CiphInVldR), .A1(n118), .Z(CiphIn[15]));
Q_AN02 U635 ( .A0(CiphInVldR), .A1(n120), .Z(CiphIn[16]));
Q_AN02 U636 ( .A0(CiphInVldR), .A1(n122), .Z(CiphIn[17]));
Q_AN02 U637 ( .A0(CiphInVldR), .A1(n124), .Z(CiphIn[18]));
Q_AN02 U638 ( .A0(CiphInVldR), .A1(n126), .Z(CiphIn[19]));
Q_AN02 U639 ( .A0(CiphInVldR), .A1(n128), .Z(CiphIn[20]));
Q_AN02 U640 ( .A0(CiphInVldR), .A1(n130), .Z(CiphIn[21]));
Q_AN02 U641 ( .A0(CiphInVldR), .A1(n132), .Z(CiphIn[22]));
Q_AN02 U642 ( .A0(CiphInVldR), .A1(n134), .Z(CiphIn[23]));
Q_AN02 U643 ( .A0(CiphInVldR), .A1(n136), .Z(CiphIn[24]));
Q_AN02 U644 ( .A0(CiphInVldR), .A1(n138), .Z(CiphIn[25]));
Q_AN02 U645 ( .A0(CiphInVldR), .A1(n140), .Z(CiphIn[26]));
Q_AN02 U646 ( .A0(CiphInVldR), .A1(n142), .Z(CiphIn[27]));
Q_AN02 U647 ( .A0(CiphInVldR), .A1(n144), .Z(CiphIn[28]));
Q_AN02 U648 ( .A0(CiphInVldR), .A1(n146), .Z(CiphIn[29]));
Q_AN02 U649 ( .A0(CiphInVldR), .A1(n148), .Z(CiphIn[30]));
Q_AN02 U650 ( .A0(CiphInVldR), .A1(n150), .Z(CiphIn[31]));
Q_AN02 U651 ( .A0(CiphInVldR), .A1(n152), .Z(CiphIn[32]));
Q_AN02 U652 ( .A0(CiphInVldR), .A1(n154), .Z(CiphIn[33]));
Q_AN02 U653 ( .A0(CiphInVldR), .A1(n156), .Z(CiphIn[34]));
Q_AN02 U654 ( .A0(CiphInVldR), .A1(n158), .Z(CiphIn[35]));
Q_AN02 U655 ( .A0(CiphInVldR), .A1(n160), .Z(CiphIn[36]));
Q_AN02 U656 ( .A0(CiphInVldR), .A1(n162), .Z(CiphIn[37]));
Q_AN02 U657 ( .A0(CiphInVldR), .A1(n164), .Z(CiphIn[38]));
Q_AN02 U658 ( .A0(CiphInVldR), .A1(n166), .Z(CiphIn[39]));
Q_AN02 U659 ( .A0(CiphInVldR), .A1(n168), .Z(CiphIn[40]));
Q_AN02 U660 ( .A0(CiphInVldR), .A1(n170), .Z(CiphIn[41]));
Q_AN02 U661 ( .A0(CiphInVldR), .A1(n172), .Z(CiphIn[42]));
Q_AN02 U662 ( .A0(CiphInVldR), .A1(n174), .Z(CiphIn[43]));
Q_AN02 U663 ( .A0(CiphInVldR), .A1(n176), .Z(CiphIn[44]));
Q_AN02 U664 ( .A0(CiphInVldR), .A1(n178), .Z(CiphIn[45]));
Q_AN02 U665 ( .A0(CiphInVldR), .A1(n180), .Z(CiphIn[46]));
Q_AN02 U666 ( .A0(CiphInVldR), .A1(n182), .Z(CiphIn[47]));
Q_AN02 U667 ( .A0(CiphInVldR), .A1(n184), .Z(CiphIn[48]));
Q_AN02 U668 ( .A0(CiphInVldR), .A1(n186), .Z(CiphIn[49]));
Q_AN02 U669 ( .A0(CiphInVldR), .A1(n188), .Z(CiphIn[50]));
Q_AN02 U670 ( .A0(CiphInVldR), .A1(n190), .Z(CiphIn[51]));
Q_AN02 U671 ( .A0(CiphInVldR), .A1(n192), .Z(CiphIn[52]));
Q_AN02 U672 ( .A0(CiphInVldR), .A1(n194), .Z(CiphIn[53]));
Q_AN02 U673 ( .A0(CiphInVldR), .A1(n196), .Z(CiphIn[54]));
Q_AN02 U674 ( .A0(CiphInVldR), .A1(n198), .Z(CiphIn[55]));
Q_AN02 U675 ( .A0(CiphInVldR), .A1(n200), .Z(CiphIn[56]));
Q_AN02 U676 ( .A0(CiphInVldR), .A1(n202), .Z(CiphIn[57]));
Q_AN02 U677 ( .A0(CiphInVldR), .A1(n204), .Z(CiphIn[58]));
Q_AN02 U678 ( .A0(CiphInVldR), .A1(n206), .Z(CiphIn[59]));
Q_AN02 U679 ( .A0(CiphInVldR), .A1(n208), .Z(CiphIn[60]));
Q_AN02 U680 ( .A0(CiphInVldR), .A1(n210), .Z(CiphIn[61]));
Q_AN02 U681 ( .A0(CiphInVldR), .A1(n212), .Z(CiphIn[62]));
Q_AN02 U682 ( .A0(CiphInVldR), .A1(n214), .Z(CiphIn[63]));
Q_AN02 U683 ( .A0(CiphInVldR), .A1(n216), .Z(CiphIn[64]));
Q_AN02 U684 ( .A0(CiphInVldR), .A1(n218), .Z(CiphIn[65]));
Q_AN02 U685 ( .A0(CiphInVldR), .A1(n220), .Z(CiphIn[66]));
Q_AN02 U686 ( .A0(CiphInVldR), .A1(n222), .Z(CiphIn[67]));
Q_AN02 U687 ( .A0(CiphInVldR), .A1(n224), .Z(CiphIn[68]));
Q_AN02 U688 ( .A0(CiphInVldR), .A1(n226), .Z(CiphIn[69]));
Q_AN02 U689 ( .A0(CiphInVldR), .A1(n228), .Z(CiphIn[70]));
Q_AN02 U690 ( .A0(CiphInVldR), .A1(n230), .Z(CiphIn[71]));
Q_AN02 U691 ( .A0(CiphInVldR), .A1(n232), .Z(CiphIn[72]));
Q_AN02 U692 ( .A0(CiphInVldR), .A1(n234), .Z(CiphIn[73]));
Q_AN02 U693 ( .A0(CiphInVldR), .A1(n236), .Z(CiphIn[74]));
Q_AN02 U694 ( .A0(CiphInVldR), .A1(n238), .Z(CiphIn[75]));
Q_AN02 U695 ( .A0(CiphInVldR), .A1(n240), .Z(CiphIn[76]));
Q_AN02 U696 ( .A0(CiphInVldR), .A1(n242), .Z(CiphIn[77]));
Q_AN02 U697 ( .A0(CiphInVldR), .A1(n244), .Z(CiphIn[78]));
Q_AN02 U698 ( .A0(CiphInVldR), .A1(n246), .Z(CiphIn[79]));
Q_AN02 U699 ( .A0(CiphInVldR), .A1(n248), .Z(CiphIn[80]));
Q_AN02 U700 ( .A0(CiphInVldR), .A1(n250), .Z(CiphIn[81]));
Q_AN02 U701 ( .A0(CiphInVldR), .A1(n252), .Z(CiphIn[82]));
Q_AN02 U702 ( .A0(CiphInVldR), .A1(n254), .Z(CiphIn[83]));
Q_AN02 U703 ( .A0(CiphInVldR), .A1(n256), .Z(CiphIn[84]));
Q_AN02 U704 ( .A0(CiphInVldR), .A1(n258), .Z(CiphIn[85]));
Q_AN02 U705 ( .A0(CiphInVldR), .A1(n260), .Z(CiphIn[86]));
Q_AN02 U706 ( .A0(CiphInVldR), .A1(n262), .Z(CiphIn[87]));
Q_AN02 U707 ( .A0(CiphInVldR), .A1(n264), .Z(CiphIn[88]));
Q_AN02 U708 ( .A0(CiphInVldR), .A1(n266), .Z(CiphIn[89]));
Q_AN02 U709 ( .A0(CiphInVldR), .A1(n268), .Z(CiphIn[90]));
Q_AN02 U710 ( .A0(CiphInVldR), .A1(n270), .Z(CiphIn[91]));
Q_AN02 U711 ( .A0(CiphInVldR), .A1(n272), .Z(CiphIn[92]));
Q_AN02 U712 ( .A0(CiphInVldR), .A1(n274), .Z(CiphIn[93]));
Q_AN02 U713 ( .A0(CiphInVldR), .A1(n276), .Z(CiphIn[94]));
Q_AN02 U714 ( .A0(CiphInVldR), .A1(n278), .Z(CiphIn[95]));
Q_AN02 U715 ( .A0(CiphInVldR), .A1(n280), .Z(CiphIn[96]));
Q_AN02 U716 ( .A0(CiphInVldR), .A1(n282), .Z(CiphIn[97]));
Q_AN02 U717 ( .A0(CiphInVldR), .A1(n284), .Z(CiphIn[98]));
Q_AN02 U718 ( .A0(CiphInVldR), .A1(n286), .Z(CiphIn[99]));
Q_AN02 U719 ( .A0(CiphInVldR), .A1(n288), .Z(CiphIn[100]));
Q_AN02 U720 ( .A0(CiphInVldR), .A1(n290), .Z(CiphIn[101]));
Q_AN02 U721 ( .A0(CiphInVldR), .A1(n292), .Z(CiphIn[102]));
Q_AN02 U722 ( .A0(CiphInVldR), .A1(n294), .Z(CiphIn[103]));
Q_AN02 U723 ( .A0(CiphInVldR), .A1(n296), .Z(CiphIn[104]));
Q_AN02 U724 ( .A0(CiphInVldR), .A1(n298), .Z(CiphIn[105]));
Q_AN02 U725 ( .A0(CiphInVldR), .A1(n300), .Z(CiphIn[106]));
Q_AN02 U726 ( .A0(CiphInVldR), .A1(n302), .Z(CiphIn[107]));
Q_AN02 U727 ( .A0(CiphInVldR), .A1(n304), .Z(CiphIn[108]));
Q_AN02 U728 ( .A0(CiphInVldR), .A1(n306), .Z(CiphIn[109]));
Q_AN02 U729 ( .A0(CiphInVldR), .A1(n308), .Z(CiphIn[110]));
Q_AN02 U730 ( .A0(CiphInVldR), .A1(n310), .Z(CiphIn[111]));
Q_AN02 U731 ( .A0(CiphInVldR), .A1(n312), .Z(CiphIn[112]));
Q_AN02 U732 ( .A0(CiphInVldR), .A1(n314), .Z(CiphIn[113]));
Q_AN02 U733 ( .A0(CiphInVldR), .A1(n316), .Z(CiphIn[114]));
Q_AN02 U734 ( .A0(CiphInVldR), .A1(n318), .Z(CiphIn[115]));
Q_AN02 U735 ( .A0(CiphInVldR), .A1(n320), .Z(CiphIn[116]));
Q_AN02 U736 ( .A0(CiphInVldR), .A1(n322), .Z(CiphIn[117]));
Q_AN02 U737 ( .A0(CiphInVldR), .A1(n324), .Z(CiphIn[118]));
Q_AN02 U738 ( .A0(CiphInVldR), .A1(n326), .Z(CiphIn[119]));
Q_AN02 U739 ( .A0(CiphInVldR), .A1(n328), .Z(CiphIn[120]));
Q_AN02 U740 ( .A0(CiphInVldR), .A1(n330), .Z(CiphIn[121]));
Q_AN02 U741 ( .A0(CiphInVldR), .A1(n332), .Z(CiphIn[122]));
Q_AN02 U742 ( .A0(CiphInVldR), .A1(n334), .Z(CiphIn[123]));
Q_AN02 U743 ( .A0(CiphInVldR), .A1(n336), .Z(CiphIn[124]));
Q_AN02 U744 ( .A0(CiphInVldR), .A1(n338), .Z(CiphIn[125]));
Q_AN02 U745 ( .A0(CiphInVldR), .A1(n340), .Z(CiphIn[126]));
Q_AN02 U746 ( .A0(CiphInVldR), .A1(n342), .Z(CiphIn[127]));
Q_AN03 U747 ( .A0(n344), .A1(n345), .A2(n343), .Z(fifo_in_valid));
Q_AN02 U748 ( .A0(AesCiphOutVldR), .A1(n3), .Z(n343));
Q_AN02 U749 ( .A0(cur_state[1]), .A1(cur_state[0]), .Z(n344));
Q_AN02 U750 ( .A0(n346), .A1(n347), .Z(KeyInVld));
Q_INV U751 ( .A(KeyInStall), .Z(n347));
Q_AN02 U752 ( .A0(n79), .A1(cur_state[0]), .Z(n346));
Q_AN03 U753 ( .A0(n348), .A1(n349), .A2(n88), .Z(CiphInLastR));
Q_AN02 U754 ( .A0(n348), .A1(n350), .Z(CiphInVldR));
Q_ND02 U755 ( .A0(fifo_in_stall), .A1(n351), .Z(n350));
Q_INV U756 ( .A(n351), .Z(n349));
Q_AO21 U757 ( .A0(n348), .A1(n352), .B0(seed_expired), .Z(drng_idle));
Q_INV U758 ( .A(n350), .Z(n352));
Q_NR02 U759 ( .A0(in_count[2]), .A1(in_count[1]), .Z(n351));
Q_INV U760 ( .A(CiphInStall), .Z(n353));
Q_AN03 U761 ( .A0(cur_state[1]), .A1(n80), .A2(n353), .Z(n348));
Q_AD01HF U762 ( .A0(reseed_counter[1]), .B0(reseed_counter[0]), .S(n354), .CO(n355));
Q_AD01HF U763 ( .A0(reseed_counter[2]), .B0(n355), .S(n356), .CO(n357));
Q_AD01HF U764 ( .A0(reseed_counter[3]), .B0(n357), .S(n358), .CO(n359));
Q_AD01HF U765 ( .A0(reseed_counter[4]), .B0(n359), .S(n360), .CO(n361));
Q_AD01HF U766 ( .A0(reseed_counter[5]), .B0(n361), .S(n362), .CO(n363));
Q_AD01HF U767 ( .A0(reseed_counter[6]), .B0(n363), .S(n364), .CO(n365));
Q_AD01HF U768 ( .A0(reseed_counter[7]), .B0(n365), .S(n366), .CO(n367));
Q_AD01HF U769 ( .A0(reseed_counter[8]), .B0(n367), .S(n368), .CO(n369));
Q_AD01HF U770 ( .A0(reseed_counter[9]), .B0(n369), .S(n370), .CO(n371));
Q_AD01HF U771 ( .A0(reseed_counter[10]), .B0(n371), .S(n372), .CO(n373));
Q_AD01HF U772 ( .A0(reseed_counter[11]), .B0(n373), .S(n374), .CO(n375));
Q_AD01HF U773 ( .A0(reseed_counter[12]), .B0(n375), .S(n376), .CO(n377));
Q_AD01HF U774 ( .A0(reseed_counter[13]), .B0(n377), .S(n378), .CO(n379));
Q_AD01HF U775 ( .A0(reseed_counter[14]), .B0(n379), .S(n380), .CO(n381));
Q_AD01HF U776 ( .A0(reseed_counter[15]), .B0(n381), .S(n382), .CO(n383));
Q_AD01HF U777 ( .A0(reseed_counter[16]), .B0(n383), .S(n384), .CO(n385));
Q_AD01HF U778 ( .A0(reseed_counter[17]), .B0(n385), .S(n386), .CO(n387));
Q_AD01HF U779 ( .A0(reseed_counter[18]), .B0(n387), .S(n388), .CO(n389));
Q_AD01HF U780 ( .A0(reseed_counter[19]), .B0(n389), .S(n390), .CO(n391));
Q_AD01HF U781 ( .A0(reseed_counter[20]), .B0(n391), .S(n392), .CO(n393));
Q_AD01HF U782 ( .A0(reseed_counter[21]), .B0(n393), .S(n394), .CO(n395));
Q_AD01HF U783 ( .A0(reseed_counter[22]), .B0(n395), .S(n396), .CO(n397));
Q_AD01HF U784 ( .A0(reseed_counter[23]), .B0(n397), .S(n398), .CO(n399));
Q_AD01HF U785 ( .A0(reseed_counter[24]), .B0(n399), .S(n400), .CO(n401));
Q_AD01HF U786 ( .A0(reseed_counter[25]), .B0(n401), .S(n402), .CO(n403));
Q_AD01HF U787 ( .A0(reseed_counter[26]), .B0(n403), .S(n404), .CO(n405));
Q_AD01HF U788 ( .A0(reseed_counter[27]), .B0(n405), .S(n406), .CO(n407));
Q_AD01HF U789 ( .A0(reseed_counter[28]), .B0(n407), .S(n408), .CO(n409));
Q_AD01HF U790 ( .A0(reseed_counter[29]), .B0(n409), .S(n410), .CO(n411));
Q_AD01HF U791 ( .A0(reseed_counter[30]), .B0(n411), .S(n412), .CO(n413));
Q_AD01HF U792 ( .A0(reseed_counter[31]), .B0(n413), .S(n414), .CO(n415));
Q_AD01HF U793 ( .A0(reseed_counter[32]), .B0(n415), .S(n416), .CO(n417));
Q_AD01HF U794 ( .A0(reseed_counter[33]), .B0(n417), .S(n418), .CO(n419));
Q_AD01HF U795 ( .A0(reseed_counter[34]), .B0(n419), .S(n420), .CO(n421));
Q_AD01HF U796 ( .A0(reseed_counter[35]), .B0(n421), .S(n422), .CO(n423));
Q_AD01HF U797 ( .A0(reseed_counter[36]), .B0(n423), .S(n424), .CO(n425));
Q_AD01HF U798 ( .A0(reseed_counter[37]), .B0(n425), .S(n426), .CO(n427));
Q_AD01HF U799 ( .A0(reseed_counter[38]), .B0(n427), .S(n428), .CO(n429));
Q_AD01HF U800 ( .A0(reseed_counter[39]), .B0(n429), .S(n430), .CO(n431));
Q_AD01HF U801 ( .A0(reseed_counter[40]), .B0(n431), .S(n432), .CO(n433));
Q_AD01HF U802 ( .A0(reseed_counter[41]), .B0(n433), .S(n434), .CO(n435));
Q_AD01HF U803 ( .A0(reseed_counter[42]), .B0(n435), .S(n436), .CO(n437));
Q_AD01HF U804 ( .A0(reseed_counter[43]), .B0(n437), .S(n438), .CO(n439));
Q_AD01HF U805 ( .A0(reseed_counter[44]), .B0(n439), .S(n440), .CO(n441));
Q_AD01HF U806 ( .A0(reseed_counter[45]), .B0(n441), .S(n442), .CO(n443));
Q_AD01HF U807 ( .A0(reseed_counter[46]), .B0(n443), .S(n444), .CO(n445));
Q_XOR2 U808 ( .A0(reseed_counter[47]), .A1(n445), .Z(n446));
Q_NR02 U809 ( .A0(n497), .A1(reseed_counter[0]), .Z(n447));
Q_AN02 U810 ( .A0(n496), .A1(n354), .Z(n448));
Q_AN02 U811 ( .A0(n496), .A1(n356), .Z(n449));
Q_AN02 U812 ( .A0(n496), .A1(n358), .Z(n450));
Q_AN02 U813 ( .A0(n496), .A1(n360), .Z(n451));
Q_AN02 U814 ( .A0(n496), .A1(n362), .Z(n452));
Q_AN02 U815 ( .A0(n496), .A1(n364), .Z(n453));
Q_AN02 U816 ( .A0(n496), .A1(n366), .Z(n454));
Q_AN02 U817 ( .A0(n496), .A1(n368), .Z(n455));
Q_AN02 U818 ( .A0(n496), .A1(n370), .Z(n456));
Q_AN02 U819 ( .A0(n496), .A1(n372), .Z(n457));
Q_AN02 U820 ( .A0(n496), .A1(n374), .Z(n458));
Q_AN02 U821 ( .A0(n496), .A1(n376), .Z(n459));
Q_AN02 U822 ( .A0(n496), .A1(n378), .Z(n460));
Q_AN02 U823 ( .A0(n496), .A1(n380), .Z(n461));
Q_AN02 U824 ( .A0(n496), .A1(n382), .Z(n462));
Q_AN02 U825 ( .A0(n496), .A1(n384), .Z(n463));
Q_AN02 U826 ( .A0(n496), .A1(n386), .Z(n464));
Q_AN02 U827 ( .A0(n496), .A1(n388), .Z(n465));
Q_AN02 U828 ( .A0(n496), .A1(n390), .Z(n466));
Q_AN02 U829 ( .A0(n496), .A1(n392), .Z(n467));
Q_AN02 U830 ( .A0(n496), .A1(n394), .Z(n468));
Q_AN02 U831 ( .A0(n496), .A1(n396), .Z(n469));
Q_AN02 U832 ( .A0(n496), .A1(n398), .Z(n470));
Q_AN02 U833 ( .A0(n496), .A1(n400), .Z(n471));
Q_AN02 U834 ( .A0(n496), .A1(n402), .Z(n472));
Q_AN02 U835 ( .A0(n496), .A1(n404), .Z(n473));
Q_AN02 U836 ( .A0(n496), .A1(n406), .Z(n474));
Q_AN02 U837 ( .A0(n496), .A1(n408), .Z(n475));
Q_AN02 U838 ( .A0(n496), .A1(n410), .Z(n476));
Q_AN02 U839 ( .A0(n496), .A1(n412), .Z(n477));
Q_AN02 U840 ( .A0(n496), .A1(n414), .Z(n478));
Q_AN02 U841 ( .A0(n496), .A1(n416), .Z(n479));
Q_AN02 U842 ( .A0(n496), .A1(n418), .Z(n480));
Q_AN02 U843 ( .A0(n496), .A1(n420), .Z(n481));
Q_AN02 U844 ( .A0(n496), .A1(n422), .Z(n482));
Q_AN02 U845 ( .A0(n496), .A1(n424), .Z(n483));
Q_AN02 U846 ( .A0(n496), .A1(n426), .Z(n484));
Q_AN02 U847 ( .A0(n496), .A1(n428), .Z(n485));
Q_AN02 U848 ( .A0(n496), .A1(n430), .Z(n486));
Q_AN02 U849 ( .A0(n496), .A1(n432), .Z(n487));
Q_AN02 U850 ( .A0(n496), .A1(n434), .Z(n488));
Q_AN02 U851 ( .A0(n496), .A1(n436), .Z(n489));
Q_AN02 U852 ( .A0(n496), .A1(n438), .Z(n490));
Q_AN02 U853 ( .A0(n496), .A1(n440), .Z(n491));
Q_AN02 U854 ( .A0(n496), .A1(n442), .Z(n492));
Q_AN02 U855 ( .A0(n496), .A1(n444), .Z(n493));
Q_AN02 U856 ( .A0(n496), .A1(n446), .Z(n494));
Q_OR02 U857 ( .A0(CiphInLastR), .A1(n497), .Z(n495));
Q_INV U858 ( .A(n497), .Z(n496));
Q_NR02 U859 ( .A0(cur_state[1]), .A1(cur_state[0]), .Z(n497));
Q_MX02 U860 ( .S(n497), .A0(AesCiphOutR[0]), .A1(seed[128]), .Z(n498));
Q_MX02 U861 ( .S(n497), .A0(AesCiphOutR[1]), .A1(seed[129]), .Z(n499));
Q_MX02 U862 ( .S(n497), .A0(AesCiphOutR[2]), .A1(seed[130]), .Z(n500));
Q_MX02 U863 ( .S(n497), .A0(AesCiphOutR[3]), .A1(seed[131]), .Z(n501));
Q_MX02 U864 ( .S(n497), .A0(AesCiphOutR[4]), .A1(seed[132]), .Z(n502));
Q_MX02 U865 ( .S(n497), .A0(AesCiphOutR[5]), .A1(seed[133]), .Z(n503));
Q_MX02 U866 ( .S(n497), .A0(AesCiphOutR[6]), .A1(seed[134]), .Z(n504));
Q_MX02 U867 ( .S(n497), .A0(AesCiphOutR[7]), .A1(seed[135]), .Z(n505));
Q_MX02 U868 ( .S(n497), .A0(AesCiphOutR[8]), .A1(seed[136]), .Z(n506));
Q_MX02 U869 ( .S(n497), .A0(AesCiphOutR[9]), .A1(seed[137]), .Z(n507));
Q_MX02 U870 ( .S(n497), .A0(AesCiphOutR[10]), .A1(seed[138]), .Z(n508));
Q_MX02 U871 ( .S(n497), .A0(AesCiphOutR[11]), .A1(seed[139]), .Z(n509));
Q_MX02 U872 ( .S(n497), .A0(AesCiphOutR[12]), .A1(seed[140]), .Z(n510));
Q_MX02 U873 ( .S(n497), .A0(AesCiphOutR[13]), .A1(seed[141]), .Z(n511));
Q_MX02 U874 ( .S(n497), .A0(AesCiphOutR[14]), .A1(seed[142]), .Z(n512));
Q_MX02 U875 ( .S(n497), .A0(AesCiphOutR[15]), .A1(seed[143]), .Z(n513));
Q_MX02 U876 ( .S(n497), .A0(AesCiphOutR[16]), .A1(seed[144]), .Z(n514));
Q_MX02 U877 ( .S(n497), .A0(AesCiphOutR[17]), .A1(seed[145]), .Z(n515));
Q_MX02 U878 ( .S(n497), .A0(AesCiphOutR[18]), .A1(seed[146]), .Z(n516));
Q_MX02 U879 ( .S(n497), .A0(AesCiphOutR[19]), .A1(seed[147]), .Z(n517));
Q_MX02 U880 ( .S(n497), .A0(AesCiphOutR[20]), .A1(seed[148]), .Z(n518));
Q_MX02 U881 ( .S(n497), .A0(AesCiphOutR[21]), .A1(seed[149]), .Z(n519));
Q_MX02 U882 ( .S(n497), .A0(AesCiphOutR[22]), .A1(seed[150]), .Z(n520));
Q_MX02 U883 ( .S(n497), .A0(AesCiphOutR[23]), .A1(seed[151]), .Z(n521));
Q_MX02 U884 ( .S(n497), .A0(AesCiphOutR[24]), .A1(seed[152]), .Z(n522));
Q_MX02 U885 ( .S(n497), .A0(AesCiphOutR[25]), .A1(seed[153]), .Z(n523));
Q_MX02 U886 ( .S(n497), .A0(AesCiphOutR[26]), .A1(seed[154]), .Z(n524));
Q_MX02 U887 ( .S(n497), .A0(AesCiphOutR[27]), .A1(seed[155]), .Z(n525));
Q_MX02 U888 ( .S(n497), .A0(AesCiphOutR[28]), .A1(seed[156]), .Z(n526));
Q_MX02 U889 ( .S(n497), .A0(AesCiphOutR[29]), .A1(seed[157]), .Z(n527));
Q_MX02 U890 ( .S(n497), .A0(AesCiphOutR[30]), .A1(seed[158]), .Z(n528));
Q_MX02 U891 ( .S(n497), .A0(AesCiphOutR[31]), .A1(seed[159]), .Z(n529));
Q_MX02 U892 ( .S(n497), .A0(AesCiphOutR[32]), .A1(seed[160]), .Z(n530));
Q_MX02 U893 ( .S(n497), .A0(AesCiphOutR[33]), .A1(seed[161]), .Z(n531));
Q_MX02 U894 ( .S(n497), .A0(AesCiphOutR[34]), .A1(seed[162]), .Z(n532));
Q_MX02 U895 ( .S(n497), .A0(AesCiphOutR[35]), .A1(seed[163]), .Z(n533));
Q_MX02 U896 ( .S(n497), .A0(AesCiphOutR[36]), .A1(seed[164]), .Z(n534));
Q_MX02 U897 ( .S(n497), .A0(AesCiphOutR[37]), .A1(seed[165]), .Z(n535));
Q_MX02 U898 ( .S(n497), .A0(AesCiphOutR[38]), .A1(seed[166]), .Z(n536));
Q_MX02 U899 ( .S(n497), .A0(AesCiphOutR[39]), .A1(seed[167]), .Z(n537));
Q_MX02 U900 ( .S(n497), .A0(AesCiphOutR[40]), .A1(seed[168]), .Z(n538));
Q_MX02 U901 ( .S(n497), .A0(AesCiphOutR[41]), .A1(seed[169]), .Z(n539));
Q_MX02 U902 ( .S(n497), .A0(AesCiphOutR[42]), .A1(seed[170]), .Z(n540));
Q_MX02 U903 ( .S(n497), .A0(AesCiphOutR[43]), .A1(seed[171]), .Z(n541));
Q_MX02 U904 ( .S(n497), .A0(AesCiphOutR[44]), .A1(seed[172]), .Z(n542));
Q_MX02 U905 ( .S(n497), .A0(AesCiphOutR[45]), .A1(seed[173]), .Z(n543));
Q_MX02 U906 ( .S(n497), .A0(AesCiphOutR[46]), .A1(seed[174]), .Z(n544));
Q_MX02 U907 ( .S(n497), .A0(AesCiphOutR[47]), .A1(seed[175]), .Z(n545));
Q_MX02 U908 ( .S(n497), .A0(AesCiphOutR[48]), .A1(seed[176]), .Z(n546));
Q_MX02 U909 ( .S(n497), .A0(AesCiphOutR[49]), .A1(seed[177]), .Z(n547));
Q_MX02 U910 ( .S(n497), .A0(AesCiphOutR[50]), .A1(seed[178]), .Z(n548));
Q_MX02 U911 ( .S(n497), .A0(AesCiphOutR[51]), .A1(seed[179]), .Z(n549));
Q_MX02 U912 ( .S(n497), .A0(AesCiphOutR[52]), .A1(seed[180]), .Z(n550));
Q_MX02 U913 ( .S(n497), .A0(AesCiphOutR[53]), .A1(seed[181]), .Z(n551));
Q_MX02 U914 ( .S(n497), .A0(AesCiphOutR[54]), .A1(seed[182]), .Z(n552));
Q_MX02 U915 ( .S(n497), .A0(AesCiphOutR[55]), .A1(seed[183]), .Z(n553));
Q_MX02 U916 ( .S(n497), .A0(AesCiphOutR[56]), .A1(seed[184]), .Z(n554));
Q_MX02 U917 ( .S(n497), .A0(AesCiphOutR[57]), .A1(seed[185]), .Z(n555));
Q_MX02 U918 ( .S(n497), .A0(AesCiphOutR[58]), .A1(seed[186]), .Z(n556));
Q_MX02 U919 ( .S(n497), .A0(AesCiphOutR[59]), .A1(seed[187]), .Z(n557));
Q_MX02 U920 ( .S(n497), .A0(AesCiphOutR[60]), .A1(seed[188]), .Z(n558));
Q_MX02 U921 ( .S(n497), .A0(AesCiphOutR[61]), .A1(seed[189]), .Z(n559));
Q_MX02 U922 ( .S(n497), .A0(AesCiphOutR[62]), .A1(seed[190]), .Z(n560));
Q_MX02 U923 ( .S(n497), .A0(AesCiphOutR[63]), .A1(seed[191]), .Z(n561));
Q_MX02 U924 ( .S(n497), .A0(AesCiphOutR[64]), .A1(seed[192]), .Z(n562));
Q_MX02 U925 ( .S(n497), .A0(AesCiphOutR[65]), .A1(seed[193]), .Z(n563));
Q_MX02 U926 ( .S(n497), .A0(AesCiphOutR[66]), .A1(seed[194]), .Z(n564));
Q_MX02 U927 ( .S(n497), .A0(AesCiphOutR[67]), .A1(seed[195]), .Z(n565));
Q_MX02 U928 ( .S(n497), .A0(AesCiphOutR[68]), .A1(seed[196]), .Z(n566));
Q_MX02 U929 ( .S(n497), .A0(AesCiphOutR[69]), .A1(seed[197]), .Z(n567));
Q_MX02 U930 ( .S(n497), .A0(AesCiphOutR[70]), .A1(seed[198]), .Z(n568));
Q_MX02 U931 ( .S(n497), .A0(AesCiphOutR[71]), .A1(seed[199]), .Z(n569));
Q_MX02 U932 ( .S(n497), .A0(AesCiphOutR[72]), .A1(seed[200]), .Z(n570));
Q_MX02 U933 ( .S(n497), .A0(AesCiphOutR[73]), .A1(seed[201]), .Z(n571));
Q_MX02 U934 ( .S(n497), .A0(AesCiphOutR[74]), .A1(seed[202]), .Z(n572));
Q_MX02 U935 ( .S(n497), .A0(AesCiphOutR[75]), .A1(seed[203]), .Z(n573));
Q_MX02 U936 ( .S(n497), .A0(AesCiphOutR[76]), .A1(seed[204]), .Z(n574));
Q_MX02 U937 ( .S(n497), .A0(AesCiphOutR[77]), .A1(seed[205]), .Z(n575));
Q_MX02 U938 ( .S(n497), .A0(AesCiphOutR[78]), .A1(seed[206]), .Z(n576));
Q_MX02 U939 ( .S(n497), .A0(AesCiphOutR[79]), .A1(seed[207]), .Z(n577));
Q_MX02 U940 ( .S(n497), .A0(AesCiphOutR[80]), .A1(seed[208]), .Z(n578));
Q_MX02 U941 ( .S(n497), .A0(AesCiphOutR[81]), .A1(seed[209]), .Z(n579));
Q_MX02 U942 ( .S(n497), .A0(AesCiphOutR[82]), .A1(seed[210]), .Z(n580));
Q_MX02 U943 ( .S(n497), .A0(AesCiphOutR[83]), .A1(seed[211]), .Z(n581));
Q_MX02 U944 ( .S(n497), .A0(AesCiphOutR[84]), .A1(seed[212]), .Z(n582));
Q_MX02 U945 ( .S(n497), .A0(AesCiphOutR[85]), .A1(seed[213]), .Z(n583));
Q_MX02 U946 ( .S(n497), .A0(AesCiphOutR[86]), .A1(seed[214]), .Z(n584));
Q_MX02 U947 ( .S(n497), .A0(AesCiphOutR[87]), .A1(seed[215]), .Z(n585));
Q_MX02 U948 ( .S(n497), .A0(AesCiphOutR[88]), .A1(seed[216]), .Z(n586));
Q_MX02 U949 ( .S(n497), .A0(AesCiphOutR[89]), .A1(seed[217]), .Z(n587));
Q_MX02 U950 ( .S(n497), .A0(AesCiphOutR[90]), .A1(seed[218]), .Z(n588));
Q_MX02 U951 ( .S(n497), .A0(AesCiphOutR[91]), .A1(seed[219]), .Z(n589));
Q_MX02 U952 ( .S(n497), .A0(AesCiphOutR[92]), .A1(seed[220]), .Z(n590));
Q_MX02 U953 ( .S(n497), .A0(AesCiphOutR[93]), .A1(seed[221]), .Z(n591));
Q_MX02 U954 ( .S(n497), .A0(AesCiphOutR[94]), .A1(seed[222]), .Z(n592));
Q_MX02 U955 ( .S(n497), .A0(AesCiphOutR[95]), .A1(seed[223]), .Z(n593));
Q_MX02 U956 ( .S(n497), .A0(AesCiphOutR[96]), .A1(seed[224]), .Z(n594));
Q_MX02 U957 ( .S(n497), .A0(AesCiphOutR[97]), .A1(seed[225]), .Z(n595));
Q_MX02 U958 ( .S(n497), .A0(AesCiphOutR[98]), .A1(seed[226]), .Z(n596));
Q_MX02 U959 ( .S(n497), .A0(AesCiphOutR[99]), .A1(seed[227]), .Z(n597));
Q_MX02 U960 ( .S(n497), .A0(AesCiphOutR[100]), .A1(seed[228]), .Z(n598));
Q_MX02 U961 ( .S(n497), .A0(AesCiphOutR[101]), .A1(seed[229]), .Z(n599));
Q_MX02 U962 ( .S(n497), .A0(AesCiphOutR[102]), .A1(seed[230]), .Z(n600));
Q_MX02 U963 ( .S(n497), .A0(AesCiphOutR[103]), .A1(seed[231]), .Z(n601));
Q_MX02 U964 ( .S(n497), .A0(AesCiphOutR[104]), .A1(seed[232]), .Z(n602));
Q_MX02 U965 ( .S(n497), .A0(AesCiphOutR[105]), .A1(seed[233]), .Z(n603));
Q_MX02 U966 ( .S(n497), .A0(AesCiphOutR[106]), .A1(seed[234]), .Z(n604));
Q_MX02 U967 ( .S(n497), .A0(AesCiphOutR[107]), .A1(seed[235]), .Z(n605));
Q_MX02 U968 ( .S(n497), .A0(AesCiphOutR[108]), .A1(seed[236]), .Z(n606));
Q_MX02 U969 ( .S(n497), .A0(AesCiphOutR[109]), .A1(seed[237]), .Z(n607));
Q_MX02 U970 ( .S(n497), .A0(AesCiphOutR[110]), .A1(seed[238]), .Z(n608));
Q_MX02 U971 ( .S(n497), .A0(AesCiphOutR[111]), .A1(seed[239]), .Z(n609));
Q_MX02 U972 ( .S(n497), .A0(AesCiphOutR[112]), .A1(seed[240]), .Z(n610));
Q_MX02 U973 ( .S(n497), .A0(AesCiphOutR[113]), .A1(seed[241]), .Z(n611));
Q_MX02 U974 ( .S(n497), .A0(AesCiphOutR[114]), .A1(seed[242]), .Z(n612));
Q_MX02 U975 ( .S(n497), .A0(AesCiphOutR[115]), .A1(seed[243]), .Z(n613));
Q_MX02 U976 ( .S(n497), .A0(AesCiphOutR[116]), .A1(seed[244]), .Z(n614));
Q_MX02 U977 ( .S(n497), .A0(AesCiphOutR[117]), .A1(seed[245]), .Z(n615));
Q_MX02 U978 ( .S(n497), .A0(AesCiphOutR[118]), .A1(seed[246]), .Z(n616));
Q_MX02 U979 ( .S(n497), .A0(AesCiphOutR[119]), .A1(seed[247]), .Z(n617));
Q_MX02 U980 ( .S(n497), .A0(AesCiphOutR[120]), .A1(seed[248]), .Z(n618));
Q_MX02 U981 ( .S(n497), .A0(AesCiphOutR[121]), .A1(seed[249]), .Z(n619));
Q_MX02 U982 ( .S(n497), .A0(AesCiphOutR[122]), .A1(seed[250]), .Z(n620));
Q_MX02 U983 ( .S(n497), .A0(AesCiphOutR[123]), .A1(seed[251]), .Z(n621));
Q_MX02 U984 ( .S(n497), .A0(AesCiphOutR[124]), .A1(seed[252]), .Z(n622));
Q_MX02 U985 ( .S(n497), .A0(AesCiphOutR[125]), .A1(seed[253]), .Z(n623));
Q_MX02 U986 ( .S(n497), .A0(AesCiphOutR[126]), .A1(seed[254]), .Z(n624));
Q_MX02 U987 ( .S(n497), .A0(AesCiphOutR[127]), .A1(seed[255]), .Z(n625));
Q_MX02 U988 ( .S(n497), .A0(AesCiphOutR[0]), .A1(seed[256]), .Z(n626));
Q_MX02 U989 ( .S(n497), .A0(AesCiphOutR[1]), .A1(seed[257]), .Z(n627));
Q_MX02 U990 ( .S(n497), .A0(AesCiphOutR[2]), .A1(seed[258]), .Z(n628));
Q_MX02 U991 ( .S(n497), .A0(AesCiphOutR[3]), .A1(seed[259]), .Z(n629));
Q_MX02 U992 ( .S(n497), .A0(AesCiphOutR[4]), .A1(seed[260]), .Z(n630));
Q_MX02 U993 ( .S(n497), .A0(AesCiphOutR[5]), .A1(seed[261]), .Z(n631));
Q_MX02 U994 ( .S(n497), .A0(AesCiphOutR[6]), .A1(seed[262]), .Z(n632));
Q_MX02 U995 ( .S(n497), .A0(AesCiphOutR[7]), .A1(seed[263]), .Z(n633));
Q_MX02 U996 ( .S(n497), .A0(AesCiphOutR[8]), .A1(seed[264]), .Z(n634));
Q_MX02 U997 ( .S(n497), .A0(AesCiphOutR[9]), .A1(seed[265]), .Z(n635));
Q_MX02 U998 ( .S(n497), .A0(AesCiphOutR[10]), .A1(seed[266]), .Z(n636));
Q_MX02 U999 ( .S(n497), .A0(AesCiphOutR[11]), .A1(seed[267]), .Z(n637));
Q_MX02 U1000 ( .S(n497), .A0(AesCiphOutR[12]), .A1(seed[268]), .Z(n638));
Q_MX02 U1001 ( .S(n497), .A0(AesCiphOutR[13]), .A1(seed[269]), .Z(n639));
Q_MX02 U1002 ( .S(n497), .A0(AesCiphOutR[14]), .A1(seed[270]), .Z(n640));
Q_MX02 U1003 ( .S(n497), .A0(AesCiphOutR[15]), .A1(seed[271]), .Z(n641));
Q_MX02 U1004 ( .S(n497), .A0(AesCiphOutR[16]), .A1(seed[272]), .Z(n642));
Q_MX02 U1005 ( .S(n497), .A0(AesCiphOutR[17]), .A1(seed[273]), .Z(n643));
Q_MX02 U1006 ( .S(n497), .A0(AesCiphOutR[18]), .A1(seed[274]), .Z(n644));
Q_MX02 U1007 ( .S(n497), .A0(AesCiphOutR[19]), .A1(seed[275]), .Z(n645));
Q_MX02 U1008 ( .S(n497), .A0(AesCiphOutR[20]), .A1(seed[276]), .Z(n646));
Q_MX02 U1009 ( .S(n497), .A0(AesCiphOutR[21]), .A1(seed[277]), .Z(n647));
Q_MX02 U1010 ( .S(n497), .A0(AesCiphOutR[22]), .A1(seed[278]), .Z(n648));
Q_MX02 U1011 ( .S(n497), .A0(AesCiphOutR[23]), .A1(seed[279]), .Z(n649));
Q_MX02 U1012 ( .S(n497), .A0(AesCiphOutR[24]), .A1(seed[280]), .Z(n650));
Q_MX02 U1013 ( .S(n497), .A0(AesCiphOutR[25]), .A1(seed[281]), .Z(n651));
Q_MX02 U1014 ( .S(n497), .A0(AesCiphOutR[26]), .A1(seed[282]), .Z(n652));
Q_MX02 U1015 ( .S(n497), .A0(AesCiphOutR[27]), .A1(seed[283]), .Z(n653));
Q_MX02 U1016 ( .S(n497), .A0(AesCiphOutR[28]), .A1(seed[284]), .Z(n654));
Q_MX02 U1017 ( .S(n497), .A0(AesCiphOutR[29]), .A1(seed[285]), .Z(n655));
Q_MX02 U1018 ( .S(n497), .A0(AesCiphOutR[30]), .A1(seed[286]), .Z(n656));
Q_MX02 U1019 ( .S(n497), .A0(AesCiphOutR[31]), .A1(seed[287]), .Z(n657));
Q_MX02 U1020 ( .S(n497), .A0(AesCiphOutR[32]), .A1(seed[288]), .Z(n658));
Q_MX02 U1021 ( .S(n497), .A0(AesCiphOutR[33]), .A1(seed[289]), .Z(n659));
Q_MX02 U1022 ( .S(n497), .A0(AesCiphOutR[34]), .A1(seed[290]), .Z(n660));
Q_MX02 U1023 ( .S(n497), .A0(AesCiphOutR[35]), .A1(seed[291]), .Z(n661));
Q_MX02 U1024 ( .S(n497), .A0(AesCiphOutR[36]), .A1(seed[292]), .Z(n662));
Q_MX02 U1025 ( .S(n497), .A0(AesCiphOutR[37]), .A1(seed[293]), .Z(n663));
Q_MX02 U1026 ( .S(n497), .A0(AesCiphOutR[38]), .A1(seed[294]), .Z(n664));
Q_MX02 U1027 ( .S(n497), .A0(AesCiphOutR[39]), .A1(seed[295]), .Z(n665));
Q_MX02 U1028 ( .S(n497), .A0(AesCiphOutR[40]), .A1(seed[296]), .Z(n666));
Q_MX02 U1029 ( .S(n497), .A0(AesCiphOutR[41]), .A1(seed[297]), .Z(n667));
Q_MX02 U1030 ( .S(n497), .A0(AesCiphOutR[42]), .A1(seed[298]), .Z(n668));
Q_MX02 U1031 ( .S(n497), .A0(AesCiphOutR[43]), .A1(seed[299]), .Z(n669));
Q_MX02 U1032 ( .S(n497), .A0(AesCiphOutR[44]), .A1(seed[300]), .Z(n670));
Q_MX02 U1033 ( .S(n497), .A0(AesCiphOutR[45]), .A1(seed[301]), .Z(n671));
Q_MX02 U1034 ( .S(n497), .A0(AesCiphOutR[46]), .A1(seed[302]), .Z(n672));
Q_MX02 U1035 ( .S(n497), .A0(AesCiphOutR[47]), .A1(seed[303]), .Z(n673));
Q_MX02 U1036 ( .S(n497), .A0(AesCiphOutR[48]), .A1(seed[304]), .Z(n674));
Q_MX02 U1037 ( .S(n497), .A0(AesCiphOutR[49]), .A1(seed[305]), .Z(n675));
Q_MX02 U1038 ( .S(n497), .A0(AesCiphOutR[50]), .A1(seed[306]), .Z(n676));
Q_MX02 U1039 ( .S(n497), .A0(AesCiphOutR[51]), .A1(seed[307]), .Z(n677));
Q_MX02 U1040 ( .S(n497), .A0(AesCiphOutR[52]), .A1(seed[308]), .Z(n678));
Q_MX02 U1041 ( .S(n497), .A0(AesCiphOutR[53]), .A1(seed[309]), .Z(n679));
Q_MX02 U1042 ( .S(n497), .A0(AesCiphOutR[54]), .A1(seed[310]), .Z(n680));
Q_MX02 U1043 ( .S(n497), .A0(AesCiphOutR[55]), .A1(seed[311]), .Z(n681));
Q_MX02 U1044 ( .S(n497), .A0(AesCiphOutR[56]), .A1(seed[312]), .Z(n682));
Q_MX02 U1045 ( .S(n497), .A0(AesCiphOutR[57]), .A1(seed[313]), .Z(n683));
Q_MX02 U1046 ( .S(n497), .A0(AesCiphOutR[58]), .A1(seed[314]), .Z(n684));
Q_MX02 U1047 ( .S(n497), .A0(AesCiphOutR[59]), .A1(seed[315]), .Z(n685));
Q_MX02 U1048 ( .S(n497), .A0(AesCiphOutR[60]), .A1(seed[316]), .Z(n686));
Q_MX02 U1049 ( .S(n497), .A0(AesCiphOutR[61]), .A1(seed[317]), .Z(n687));
Q_MX02 U1050 ( .S(n497), .A0(AesCiphOutR[62]), .A1(seed[318]), .Z(n688));
Q_MX02 U1051 ( .S(n497), .A0(AesCiphOutR[63]), .A1(seed[319]), .Z(n689));
Q_MX02 U1052 ( .S(n497), .A0(AesCiphOutR[64]), .A1(seed[320]), .Z(n690));
Q_MX02 U1053 ( .S(n497), .A0(AesCiphOutR[65]), .A1(seed[321]), .Z(n691));
Q_MX02 U1054 ( .S(n497), .A0(AesCiphOutR[66]), .A1(seed[322]), .Z(n692));
Q_MX02 U1055 ( .S(n497), .A0(AesCiphOutR[67]), .A1(seed[323]), .Z(n693));
Q_MX02 U1056 ( .S(n497), .A0(AesCiphOutR[68]), .A1(seed[324]), .Z(n694));
Q_MX02 U1057 ( .S(n497), .A0(AesCiphOutR[69]), .A1(seed[325]), .Z(n695));
Q_MX02 U1058 ( .S(n497), .A0(AesCiphOutR[70]), .A1(seed[326]), .Z(n696));
Q_MX02 U1059 ( .S(n497), .A0(AesCiphOutR[71]), .A1(seed[327]), .Z(n697));
Q_MX02 U1060 ( .S(n497), .A0(AesCiphOutR[72]), .A1(seed[328]), .Z(n698));
Q_MX02 U1061 ( .S(n497), .A0(AesCiphOutR[73]), .A1(seed[329]), .Z(n699));
Q_MX02 U1062 ( .S(n497), .A0(AesCiphOutR[74]), .A1(seed[330]), .Z(n700));
Q_MX02 U1063 ( .S(n497), .A0(AesCiphOutR[75]), .A1(seed[331]), .Z(n701));
Q_MX02 U1064 ( .S(n497), .A0(AesCiphOutR[76]), .A1(seed[332]), .Z(n702));
Q_MX02 U1065 ( .S(n497), .A0(AesCiphOutR[77]), .A1(seed[333]), .Z(n703));
Q_MX02 U1066 ( .S(n497), .A0(AesCiphOutR[78]), .A1(seed[334]), .Z(n704));
Q_MX02 U1067 ( .S(n497), .A0(AesCiphOutR[79]), .A1(seed[335]), .Z(n705));
Q_MX02 U1068 ( .S(n497), .A0(AesCiphOutR[80]), .A1(seed[336]), .Z(n706));
Q_MX02 U1069 ( .S(n497), .A0(AesCiphOutR[81]), .A1(seed[337]), .Z(n707));
Q_MX02 U1070 ( .S(n497), .A0(AesCiphOutR[82]), .A1(seed[338]), .Z(n708));
Q_MX02 U1071 ( .S(n497), .A0(AesCiphOutR[83]), .A1(seed[339]), .Z(n709));
Q_MX02 U1072 ( .S(n497), .A0(AesCiphOutR[84]), .A1(seed[340]), .Z(n710));
Q_MX02 U1073 ( .S(n497), .A0(AesCiphOutR[85]), .A1(seed[341]), .Z(n711));
Q_MX02 U1074 ( .S(n497), .A0(AesCiphOutR[86]), .A1(seed[342]), .Z(n712));
Q_MX02 U1075 ( .S(n497), .A0(AesCiphOutR[87]), .A1(seed[343]), .Z(n713));
Q_MX02 U1076 ( .S(n497), .A0(AesCiphOutR[88]), .A1(seed[344]), .Z(n714));
Q_MX02 U1077 ( .S(n497), .A0(AesCiphOutR[89]), .A1(seed[345]), .Z(n715));
Q_MX02 U1078 ( .S(n497), .A0(AesCiphOutR[90]), .A1(seed[346]), .Z(n716));
Q_MX02 U1079 ( .S(n497), .A0(AesCiphOutR[91]), .A1(seed[347]), .Z(n717));
Q_MX02 U1080 ( .S(n497), .A0(AesCiphOutR[92]), .A1(seed[348]), .Z(n718));
Q_MX02 U1081 ( .S(n497), .A0(AesCiphOutR[93]), .A1(seed[349]), .Z(n719));
Q_MX02 U1082 ( .S(n497), .A0(AesCiphOutR[94]), .A1(seed[350]), .Z(n720));
Q_MX02 U1083 ( .S(n497), .A0(AesCiphOutR[95]), .A1(seed[351]), .Z(n721));
Q_MX02 U1084 ( .S(n497), .A0(AesCiphOutR[96]), .A1(seed[352]), .Z(n722));
Q_MX02 U1085 ( .S(n497), .A0(AesCiphOutR[97]), .A1(seed[353]), .Z(n723));
Q_MX02 U1086 ( .S(n497), .A0(AesCiphOutR[98]), .A1(seed[354]), .Z(n724));
Q_MX02 U1087 ( .S(n497), .A0(AesCiphOutR[99]), .A1(seed[355]), .Z(n725));
Q_MX02 U1088 ( .S(n497), .A0(AesCiphOutR[100]), .A1(seed[356]), .Z(n726));
Q_MX02 U1089 ( .S(n497), .A0(AesCiphOutR[101]), .A1(seed[357]), .Z(n727));
Q_MX02 U1090 ( .S(n497), .A0(AesCiphOutR[102]), .A1(seed[358]), .Z(n728));
Q_MX02 U1091 ( .S(n497), .A0(AesCiphOutR[103]), .A1(seed[359]), .Z(n729));
Q_MX02 U1092 ( .S(n497), .A0(AesCiphOutR[104]), .A1(seed[360]), .Z(n730));
Q_MX02 U1093 ( .S(n497), .A0(AesCiphOutR[105]), .A1(seed[361]), .Z(n731));
Q_MX02 U1094 ( .S(n497), .A0(AesCiphOutR[106]), .A1(seed[362]), .Z(n732));
Q_MX02 U1095 ( .S(n497), .A0(AesCiphOutR[107]), .A1(seed[363]), .Z(n733));
Q_MX02 U1096 ( .S(n497), .A0(AesCiphOutR[108]), .A1(seed[364]), .Z(n734));
Q_MX02 U1097 ( .S(n497), .A0(AesCiphOutR[109]), .A1(seed[365]), .Z(n735));
Q_MX02 U1098 ( .S(n497), .A0(AesCiphOutR[110]), .A1(seed[366]), .Z(n736));
Q_MX02 U1099 ( .S(n497), .A0(AesCiphOutR[111]), .A1(seed[367]), .Z(n737));
Q_MX02 U1100 ( .S(n497), .A0(AesCiphOutR[112]), .A1(seed[368]), .Z(n738));
Q_MX02 U1101 ( .S(n497), .A0(AesCiphOutR[113]), .A1(seed[369]), .Z(n739));
Q_MX02 U1102 ( .S(n497), .A0(AesCiphOutR[114]), .A1(seed[370]), .Z(n740));
Q_MX02 U1103 ( .S(n497), .A0(AesCiphOutR[115]), .A1(seed[371]), .Z(n741));
Q_MX02 U1104 ( .S(n497), .A0(AesCiphOutR[116]), .A1(seed[372]), .Z(n742));
Q_MX02 U1105 ( .S(n497), .A0(AesCiphOutR[117]), .A1(seed[373]), .Z(n743));
Q_MX02 U1106 ( .S(n497), .A0(AesCiphOutR[118]), .A1(seed[374]), .Z(n744));
Q_MX02 U1107 ( .S(n497), .A0(AesCiphOutR[119]), .A1(seed[375]), .Z(n745));
Q_MX02 U1108 ( .S(n497), .A0(AesCiphOutR[120]), .A1(seed[376]), .Z(n746));
Q_MX02 U1109 ( .S(n497), .A0(AesCiphOutR[121]), .A1(seed[377]), .Z(n747));
Q_MX02 U1110 ( .S(n497), .A0(AesCiphOutR[122]), .A1(seed[378]), .Z(n748));
Q_MX02 U1111 ( .S(n497), .A0(AesCiphOutR[123]), .A1(seed[379]), .Z(n749));
Q_MX02 U1112 ( .S(n497), .A0(AesCiphOutR[124]), .A1(seed[380]), .Z(n750));
Q_MX02 U1113 ( .S(n497), .A0(AesCiphOutR[125]), .A1(seed[381]), .Z(n751));
Q_MX02 U1114 ( .S(n497), .A0(AesCiphOutR[126]), .A1(seed[382]), .Z(n752));
Q_MX02 U1115 ( .S(n497), .A0(AesCiphOutR[127]), .A1(seed[383]), .Z(n753));
Q_AO21 U1116 ( .A0(n343), .A1(n754), .B0(n497), .Z(n757));
Q_AN02 U1117 ( .A0(out_count[1]), .A1(n755), .Z(n754));
Q_AO21 U1118 ( .A0(n343), .A1(n756), .B0(n497), .Z(n758));
Q_AN02 U1119 ( .A0(out_count[1]), .A1(out_count[0]), .Z(n756));
Q_AD01HF U1120 ( .A0(internal_state_value[1]), .B0(internal_state_value[0]), .S(n760), .CO(n761));
Q_AD01HF U1121 ( .A0(internal_state_value[2]), .B0(n761), .S(n762), .CO(n763));
Q_AD01HF U1122 ( .A0(internal_state_value[3]), .B0(n763), .S(n764), .CO(n765));
Q_AD01HF U1123 ( .A0(internal_state_value[4]), .B0(n765), .S(n766), .CO(n767));
Q_AD01HF U1124 ( .A0(internal_state_value[5]), .B0(n767), .S(n768), .CO(n769));
Q_AD01HF U1125 ( .A0(internal_state_value[6]), .B0(n769), .S(n770), .CO(n771));
Q_AD01HF U1126 ( .A0(internal_state_value[7]), .B0(n771), .S(n772), .CO(n773));
Q_AD01HF U1127 ( .A0(internal_state_value[8]), .B0(n773), .S(n774), .CO(n775));
Q_AD01HF U1128 ( .A0(internal_state_value[9]), .B0(n775), .S(n776), .CO(n777));
Q_AD01HF U1129 ( .A0(internal_state_value[10]), .B0(n777), .S(n778), .CO(n779));
Q_AD01HF U1130 ( .A0(internal_state_value[11]), .B0(n779), .S(n780), .CO(n781));
Q_AD01HF U1131 ( .A0(internal_state_value[12]), .B0(n781), .S(n782), .CO(n783));
Q_AD01HF U1132 ( .A0(internal_state_value[13]), .B0(n783), .S(n784), .CO(n785));
Q_AD01HF U1133 ( .A0(internal_state_value[14]), .B0(n785), .S(n786), .CO(n787));
Q_AD01HF U1134 ( .A0(internal_state_value[15]), .B0(n787), .S(n788), .CO(n789));
Q_AD01HF U1135 ( .A0(internal_state_value[16]), .B0(n789), .S(n790), .CO(n791));
Q_AD01HF U1136 ( .A0(internal_state_value[17]), .B0(n791), .S(n792), .CO(n793));
Q_AD01HF U1137 ( .A0(internal_state_value[18]), .B0(n793), .S(n794), .CO(n795));
Q_AD01HF U1138 ( .A0(internal_state_value[19]), .B0(n795), .S(n796), .CO(n797));
Q_AD01HF U1139 ( .A0(internal_state_value[20]), .B0(n797), .S(n798), .CO(n799));
Q_AD01HF U1140 ( .A0(internal_state_value[21]), .B0(n799), .S(n800), .CO(n801));
Q_AD01HF U1141 ( .A0(internal_state_value[22]), .B0(n801), .S(n802), .CO(n803));
Q_AD01HF U1142 ( .A0(internal_state_value[23]), .B0(n803), .S(n804), .CO(n805));
Q_AD01HF U1143 ( .A0(internal_state_value[24]), .B0(n805), .S(n806), .CO(n807));
Q_AD01HF U1144 ( .A0(internal_state_value[25]), .B0(n807), .S(n808), .CO(n809));
Q_AD01HF U1145 ( .A0(internal_state_value[26]), .B0(n809), .S(n810), .CO(n811));
Q_AD01HF U1146 ( .A0(internal_state_value[27]), .B0(n811), .S(n812), .CO(n813));
Q_AD01HF U1147 ( .A0(internal_state_value[28]), .B0(n813), .S(n814), .CO(n815));
Q_AD01HF U1148 ( .A0(internal_state_value[29]), .B0(n815), .S(n816), .CO(n817));
Q_AD01HF U1149 ( .A0(internal_state_value[30]), .B0(n817), .S(n818), .CO(n819));
Q_AD01HF U1150 ( .A0(internal_state_value[31]), .B0(n819), .S(n820), .CO(n821));
Q_AD01HF U1151 ( .A0(internal_state_value[32]), .B0(n821), .S(n822), .CO(n823));
Q_AD01HF U1152 ( .A0(internal_state_value[33]), .B0(n823), .S(n824), .CO(n825));
Q_AD01HF U1153 ( .A0(internal_state_value[34]), .B0(n825), .S(n826), .CO(n827));
Q_AD01HF U1154 ( .A0(internal_state_value[35]), .B0(n827), .S(n828), .CO(n829));
Q_AD01HF U1155 ( .A0(internal_state_value[36]), .B0(n829), .S(n830), .CO(n831));
Q_AD01HF U1156 ( .A0(internal_state_value[37]), .B0(n831), .S(n832), .CO(n833));
Q_AD01HF U1157 ( .A0(internal_state_value[38]), .B0(n833), .S(n834), .CO(n835));
Q_AD01HF U1158 ( .A0(internal_state_value[39]), .B0(n835), .S(n836), .CO(n837));
Q_AD01HF U1159 ( .A0(internal_state_value[40]), .B0(n837), .S(n838), .CO(n839));
Q_AD01HF U1160 ( .A0(internal_state_value[41]), .B0(n839), .S(n840), .CO(n841));
Q_AD01HF U1161 ( .A0(internal_state_value[42]), .B0(n841), .S(n842), .CO(n843));
Q_AD01HF U1162 ( .A0(internal_state_value[43]), .B0(n843), .S(n844), .CO(n845));
Q_AD01HF U1163 ( .A0(internal_state_value[44]), .B0(n845), .S(n846), .CO(n847));
Q_AD01HF U1164 ( .A0(internal_state_value[45]), .B0(n847), .S(n848), .CO(n849));
Q_AD01HF U1165 ( .A0(internal_state_value[46]), .B0(n849), .S(n850), .CO(n851));
Q_AD01HF U1166 ( .A0(internal_state_value[47]), .B0(n851), .S(n852), .CO(n853));
Q_AD01HF U1167 ( .A0(internal_state_value[48]), .B0(n853), .S(n854), .CO(n855));
Q_AD01HF U1168 ( .A0(internal_state_value[49]), .B0(n855), .S(n856), .CO(n857));
Q_AD01HF U1169 ( .A0(internal_state_value[50]), .B0(n857), .S(n858), .CO(n859));
Q_AD01HF U1170 ( .A0(internal_state_value[51]), .B0(n859), .S(n860), .CO(n861));
Q_AD01HF U1171 ( .A0(internal_state_value[52]), .B0(n861), .S(n862), .CO(n863));
Q_AD01HF U1172 ( .A0(internal_state_value[53]), .B0(n863), .S(n864), .CO(n865));
Q_AD01HF U1173 ( .A0(internal_state_value[54]), .B0(n865), .S(n866), .CO(n867));
Q_AD01HF U1174 ( .A0(internal_state_value[55]), .B0(n867), .S(n868), .CO(n869));
Q_AD01HF U1175 ( .A0(internal_state_value[56]), .B0(n869), .S(n870), .CO(n871));
Q_AD01HF U1176 ( .A0(internal_state_value[57]), .B0(n871), .S(n872), .CO(n873));
Q_AD01HF U1177 ( .A0(internal_state_value[58]), .B0(n873), .S(n874), .CO(n875));
Q_AD01HF U1178 ( .A0(internal_state_value[59]), .B0(n875), .S(n876), .CO(n877));
Q_AD01HF U1179 ( .A0(internal_state_value[60]), .B0(n877), .S(n878), .CO(n879));
Q_AD01HF U1180 ( .A0(internal_state_value[61]), .B0(n879), .S(n880), .CO(n881));
Q_AD01HF U1181 ( .A0(internal_state_value[62]), .B0(n881), .S(n882), .CO(n883));
Q_AD01HF U1182 ( .A0(internal_state_value[63]), .B0(n883), .S(n884), .CO(n885));
Q_AD01HF U1183 ( .A0(internal_state_value[64]), .B0(n885), .S(n886), .CO(n887));
Q_AD01HF U1184 ( .A0(internal_state_value[65]), .B0(n887), .S(n888), .CO(n889));
Q_AD01HF U1185 ( .A0(internal_state_value[66]), .B0(n889), .S(n890), .CO(n891));
Q_AD01HF U1186 ( .A0(internal_state_value[67]), .B0(n891), .S(n892), .CO(n893));
Q_AD01HF U1187 ( .A0(internal_state_value[68]), .B0(n893), .S(n894), .CO(n895));
Q_AD01HF U1188 ( .A0(internal_state_value[69]), .B0(n895), .S(n896), .CO(n897));
Q_AD01HF U1189 ( .A0(internal_state_value[70]), .B0(n897), .S(n898), .CO(n899));
Q_AD01HF U1190 ( .A0(internal_state_value[71]), .B0(n899), .S(n900), .CO(n901));
Q_AD01HF U1191 ( .A0(internal_state_value[72]), .B0(n901), .S(n902), .CO(n903));
Q_AD01HF U1192 ( .A0(internal_state_value[73]), .B0(n903), .S(n904), .CO(n905));
Q_AD01HF U1193 ( .A0(internal_state_value[74]), .B0(n905), .S(n906), .CO(n907));
Q_AD01HF U1194 ( .A0(internal_state_value[75]), .B0(n907), .S(n908), .CO(n909));
Q_AD01HF U1195 ( .A0(internal_state_value[76]), .B0(n909), .S(n910), .CO(n911));
Q_AD01HF U1196 ( .A0(internal_state_value[77]), .B0(n911), .S(n912), .CO(n913));
Q_AD01HF U1197 ( .A0(internal_state_value[78]), .B0(n913), .S(n914), .CO(n915));
Q_AD01HF U1198 ( .A0(internal_state_value[79]), .B0(n915), .S(n916), .CO(n917));
Q_AD01HF U1199 ( .A0(internal_state_value[80]), .B0(n917), .S(n918), .CO(n919));
Q_AD01HF U1200 ( .A0(internal_state_value[81]), .B0(n919), .S(n920), .CO(n921));
Q_AD01HF U1201 ( .A0(internal_state_value[82]), .B0(n921), .S(n922), .CO(n923));
Q_AD01HF U1202 ( .A0(internal_state_value[83]), .B0(n923), .S(n924), .CO(n925));
Q_AD01HF U1203 ( .A0(internal_state_value[84]), .B0(n925), .S(n926), .CO(n927));
Q_AD01HF U1204 ( .A0(internal_state_value[85]), .B0(n927), .S(n928), .CO(n929));
Q_AD01HF U1205 ( .A0(internal_state_value[86]), .B0(n929), .S(n930), .CO(n931));
Q_AD01HF U1206 ( .A0(internal_state_value[87]), .B0(n931), .S(n932), .CO(n933));
Q_AD01HF U1207 ( .A0(internal_state_value[88]), .B0(n933), .S(n934), .CO(n935));
Q_AD01HF U1208 ( .A0(internal_state_value[89]), .B0(n935), .S(n936), .CO(n937));
Q_AD01HF U1209 ( .A0(internal_state_value[90]), .B0(n937), .S(n938), .CO(n939));
Q_AD01HF U1210 ( .A0(internal_state_value[91]), .B0(n939), .S(n940), .CO(n941));
Q_AD01HF U1211 ( .A0(internal_state_value[92]), .B0(n941), .S(n942), .CO(n943));
Q_AD01HF U1212 ( .A0(internal_state_value[93]), .B0(n943), .S(n944), .CO(n945));
Q_AD01HF U1213 ( .A0(internal_state_value[94]), .B0(n945), .S(n946), .CO(n947));
Q_AD01HF U1214 ( .A0(internal_state_value[95]), .B0(n947), .S(n948), .CO(n949));
Q_AD01HF U1215 ( .A0(internal_state_value[96]), .B0(n949), .S(n950), .CO(n951));
Q_AD01HF U1216 ( .A0(internal_state_value[97]), .B0(n951), .S(n952), .CO(n953));
Q_AD01HF U1217 ( .A0(internal_state_value[98]), .B0(n953), .S(n954), .CO(n955));
Q_AD01HF U1218 ( .A0(internal_state_value[99]), .B0(n955), .S(n956), .CO(n957));
Q_AD01HF U1219 ( .A0(internal_state_value[100]), .B0(n957), .S(n958), .CO(n959));
Q_AD01HF U1220 ( .A0(internal_state_value[101]), .B0(n959), .S(n960), .CO(n961));
Q_AD01HF U1221 ( .A0(internal_state_value[102]), .B0(n961), .S(n962), .CO(n963));
Q_AD01HF U1222 ( .A0(internal_state_value[103]), .B0(n963), .S(n964), .CO(n965));
Q_AD01HF U1223 ( .A0(internal_state_value[104]), .B0(n965), .S(n966), .CO(n967));
Q_AD01HF U1224 ( .A0(internal_state_value[105]), .B0(n967), .S(n968), .CO(n969));
Q_AD01HF U1225 ( .A0(internal_state_value[106]), .B0(n969), .S(n970), .CO(n971));
Q_AD01HF U1226 ( .A0(internal_state_value[107]), .B0(n971), .S(n972), .CO(n973));
Q_AD01HF U1227 ( .A0(internal_state_value[108]), .B0(n973), .S(n974), .CO(n975));
Q_AD01HF U1228 ( .A0(internal_state_value[109]), .B0(n975), .S(n976), .CO(n977));
Q_AD01HF U1229 ( .A0(internal_state_value[110]), .B0(n977), .S(n978), .CO(n979));
Q_AD01HF U1230 ( .A0(internal_state_value[111]), .B0(n979), .S(n980), .CO(n981));
Q_AD01HF U1231 ( .A0(internal_state_value[112]), .B0(n981), .S(n982), .CO(n983));
Q_AD01HF U1232 ( .A0(internal_state_value[113]), .B0(n983), .S(n984), .CO(n985));
Q_AD01HF U1233 ( .A0(internal_state_value[114]), .B0(n985), .S(n986), .CO(n987));
Q_AD01HF U1234 ( .A0(internal_state_value[115]), .B0(n987), .S(n988), .CO(n989));
Q_AD01HF U1235 ( .A0(internal_state_value[116]), .B0(n989), .S(n990), .CO(n991));
Q_AD01HF U1236 ( .A0(internal_state_value[117]), .B0(n991), .S(n992), .CO(n993));
Q_AD01HF U1237 ( .A0(internal_state_value[118]), .B0(n993), .S(n994), .CO(n995));
Q_AD01HF U1238 ( .A0(internal_state_value[119]), .B0(n995), .S(n996), .CO(n997));
Q_AD01HF U1239 ( .A0(internal_state_value[120]), .B0(n997), .S(n998), .CO(n999));
Q_AD01HF U1240 ( .A0(internal_state_value[121]), .B0(n999), .S(n1000), .CO(n1001));
Q_AD01HF U1241 ( .A0(internal_state_value[122]), .B0(n1001), .S(n1002), .CO(n1003));
Q_AD01HF U1242 ( .A0(internal_state_value[123]), .B0(n1003), .S(n1004), .CO(n1005));
Q_AD01HF U1243 ( .A0(internal_state_value[124]), .B0(n1005), .S(n1006), .CO(n1007));
Q_AD01HF U1244 ( .A0(internal_state_value[125]), .B0(n1007), .S(n1008), .CO(n1009));
Q_AD01HF U1245 ( .A0(internal_state_value[126]), .B0(n1009), .S(n1010), .CO(n1011));
Q_XOR2 U1246 ( .A0(internal_state_value[127]), .A1(n1011), .Z(n1012));
Q_MX03 U1247 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[0]), .A1(seed[0]), .A2(n759), .Z(n1013));
Q_MX03 U1248 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[1]), .A1(seed[1]), .A2(n760), .Z(n1014));
Q_MX03 U1249 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[2]), .A1(seed[2]), .A2(n762), .Z(n1015));
Q_MX03 U1250 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[3]), .A1(seed[3]), .A2(n764), .Z(n1016));
Q_MX03 U1251 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[4]), .A1(seed[4]), .A2(n766), .Z(n1017));
Q_MX03 U1252 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[5]), .A1(seed[5]), .A2(n768), .Z(n1018));
Q_MX03 U1253 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[6]), .A1(seed[6]), .A2(n770), .Z(n1019));
Q_MX03 U1254 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[7]), .A1(seed[7]), .A2(n772), .Z(n1020));
Q_MX03 U1255 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[8]), .A1(seed[8]), .A2(n774), .Z(n1021));
Q_MX03 U1256 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[9]), .A1(seed[9]), .A2(n776), .Z(n1022));
Q_MX03 U1257 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[10]), .A1(seed[10]), .A2(n778), .Z(n1023));
Q_MX03 U1258 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[11]), .A1(seed[11]), .A2(n780), .Z(n1024));
Q_MX03 U1259 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[12]), .A1(seed[12]), .A2(n782), .Z(n1025));
Q_MX03 U1260 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[13]), .A1(seed[13]), .A2(n784), .Z(n1026));
Q_MX03 U1261 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[14]), .A1(seed[14]), .A2(n786), .Z(n1027));
Q_MX03 U1262 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[15]), .A1(seed[15]), .A2(n788), .Z(n1028));
Q_MX03 U1263 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[16]), .A1(seed[16]), .A2(n790), .Z(n1029));
Q_MX03 U1264 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[17]), .A1(seed[17]), .A2(n792), .Z(n1030));
Q_MX03 U1265 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[18]), .A1(seed[18]), .A2(n794), .Z(n1031));
Q_MX03 U1266 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[19]), .A1(seed[19]), .A2(n796), .Z(n1032));
Q_MX03 U1267 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[20]), .A1(seed[20]), .A2(n798), .Z(n1033));
Q_MX03 U1268 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[21]), .A1(seed[21]), .A2(n800), .Z(n1034));
Q_MX03 U1269 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[22]), .A1(seed[22]), .A2(n802), .Z(n1035));
Q_MX03 U1270 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[23]), .A1(seed[23]), .A2(n804), .Z(n1036));
Q_MX03 U1271 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[24]), .A1(seed[24]), .A2(n806), .Z(n1037));
Q_MX03 U1272 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[25]), .A1(seed[25]), .A2(n808), .Z(n1038));
Q_MX03 U1273 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[26]), .A1(seed[26]), .A2(n810), .Z(n1039));
Q_MX03 U1274 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[27]), .A1(seed[27]), .A2(n812), .Z(n1040));
Q_MX03 U1275 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[28]), .A1(seed[28]), .A2(n814), .Z(n1041));
Q_MX03 U1276 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[29]), .A1(seed[29]), .A2(n816), .Z(n1042));
Q_MX03 U1277 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[30]), .A1(seed[30]), .A2(n818), .Z(n1043));
Q_MX03 U1278 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[31]), .A1(seed[31]), .A2(n820), .Z(n1044));
Q_MX03 U1279 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[32]), .A1(seed[32]), .A2(n822), .Z(n1045));
Q_MX03 U1280 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[33]), .A1(seed[33]), .A2(n824), .Z(n1046));
Q_MX03 U1281 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[34]), .A1(seed[34]), .A2(n826), .Z(n1047));
Q_MX03 U1282 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[35]), .A1(seed[35]), .A2(n828), .Z(n1048));
Q_MX03 U1283 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[36]), .A1(seed[36]), .A2(n830), .Z(n1049));
Q_MX03 U1284 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[37]), .A1(seed[37]), .A2(n832), .Z(n1050));
Q_MX03 U1285 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[38]), .A1(seed[38]), .A2(n834), .Z(n1051));
Q_MX03 U1286 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[39]), .A1(seed[39]), .A2(n836), .Z(n1052));
Q_MX03 U1287 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[40]), .A1(seed[40]), .A2(n838), .Z(n1053));
Q_MX03 U1288 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[41]), .A1(seed[41]), .A2(n840), .Z(n1054));
Q_MX03 U1289 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[42]), .A1(seed[42]), .A2(n842), .Z(n1055));
Q_MX03 U1290 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[43]), .A1(seed[43]), .A2(n844), .Z(n1056));
Q_MX03 U1291 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[44]), .A1(seed[44]), .A2(n846), .Z(n1057));
Q_MX03 U1292 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[45]), .A1(seed[45]), .A2(n848), .Z(n1058));
Q_MX03 U1293 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[46]), .A1(seed[46]), .A2(n850), .Z(n1059));
Q_MX03 U1294 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[47]), .A1(seed[47]), .A2(n852), .Z(n1060));
Q_MX03 U1295 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[48]), .A1(seed[48]), .A2(n854), .Z(n1061));
Q_MX03 U1296 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[49]), .A1(seed[49]), .A2(n856), .Z(n1062));
Q_MX03 U1297 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[50]), .A1(seed[50]), .A2(n858), .Z(n1063));
Q_MX03 U1298 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[51]), .A1(seed[51]), .A2(n860), .Z(n1064));
Q_MX03 U1299 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[52]), .A1(seed[52]), .A2(n862), .Z(n1065));
Q_MX03 U1300 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[53]), .A1(seed[53]), .A2(n864), .Z(n1066));
Q_MX03 U1301 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[54]), .A1(seed[54]), .A2(n866), .Z(n1067));
Q_MX03 U1302 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[55]), .A1(seed[55]), .A2(n868), .Z(n1068));
Q_MX03 U1303 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[56]), .A1(seed[56]), .A2(n870), .Z(n1069));
Q_MX03 U1304 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[57]), .A1(seed[57]), .A2(n872), .Z(n1070));
Q_MX03 U1305 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[58]), .A1(seed[58]), .A2(n874), .Z(n1071));
Q_MX03 U1306 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[59]), .A1(seed[59]), .A2(n876), .Z(n1072));
Q_MX03 U1307 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[60]), .A1(seed[60]), .A2(n878), .Z(n1073));
Q_MX03 U1308 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[61]), .A1(seed[61]), .A2(n880), .Z(n1074));
Q_MX03 U1309 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[62]), .A1(seed[62]), .A2(n882), .Z(n1075));
Q_MX03 U1310 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[63]), .A1(seed[63]), .A2(n884), .Z(n1076));
Q_MX03 U1311 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[64]), .A1(seed[64]), .A2(n886), .Z(n1077));
Q_MX03 U1312 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[65]), .A1(seed[65]), .A2(n888), .Z(n1078));
Q_MX03 U1313 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[66]), .A1(seed[66]), .A2(n890), .Z(n1079));
Q_MX03 U1314 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[67]), .A1(seed[67]), .A2(n892), .Z(n1080));
Q_MX03 U1315 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[68]), .A1(seed[68]), .A2(n894), .Z(n1081));
Q_MX03 U1316 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[69]), .A1(seed[69]), .A2(n896), .Z(n1082));
Q_MX03 U1317 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[70]), .A1(seed[70]), .A2(n898), .Z(n1083));
Q_MX03 U1318 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[71]), .A1(seed[71]), .A2(n900), .Z(n1084));
Q_MX03 U1319 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[72]), .A1(seed[72]), .A2(n902), .Z(n1085));
Q_MX03 U1320 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[73]), .A1(seed[73]), .A2(n904), .Z(n1086));
Q_MX03 U1321 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[74]), .A1(seed[74]), .A2(n906), .Z(n1087));
Q_MX03 U1322 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[75]), .A1(seed[75]), .A2(n908), .Z(n1088));
Q_MX03 U1323 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[76]), .A1(seed[76]), .A2(n910), .Z(n1089));
Q_MX03 U1324 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[77]), .A1(seed[77]), .A2(n912), .Z(n1090));
Q_MX03 U1325 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[78]), .A1(seed[78]), .A2(n914), .Z(n1091));
Q_MX03 U1326 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[79]), .A1(seed[79]), .A2(n916), .Z(n1092));
Q_MX03 U1327 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[80]), .A1(seed[80]), .A2(n918), .Z(n1093));
Q_MX03 U1328 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[81]), .A1(seed[81]), .A2(n920), .Z(n1094));
Q_MX03 U1329 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[82]), .A1(seed[82]), .A2(n922), .Z(n1095));
Q_MX03 U1330 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[83]), .A1(seed[83]), .A2(n924), .Z(n1096));
Q_MX03 U1331 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[84]), .A1(seed[84]), .A2(n926), .Z(n1097));
Q_MX03 U1332 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[85]), .A1(seed[85]), .A2(n928), .Z(n1098));
Q_MX03 U1333 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[86]), .A1(seed[86]), .A2(n930), .Z(n1099));
Q_MX03 U1334 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[87]), .A1(seed[87]), .A2(n932), .Z(n1100));
Q_MX03 U1335 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[88]), .A1(seed[88]), .A2(n934), .Z(n1101));
Q_MX03 U1336 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[89]), .A1(seed[89]), .A2(n936), .Z(n1102));
Q_MX03 U1337 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[90]), .A1(seed[90]), .A2(n938), .Z(n1103));
Q_MX03 U1338 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[91]), .A1(seed[91]), .A2(n940), .Z(n1104));
Q_MX03 U1339 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[92]), .A1(seed[92]), .A2(n942), .Z(n1105));
Q_MX03 U1340 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[93]), .A1(seed[93]), .A2(n944), .Z(n1106));
Q_MX03 U1341 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[94]), .A1(seed[94]), .A2(n946), .Z(n1107));
Q_MX03 U1342 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[95]), .A1(seed[95]), .A2(n948), .Z(n1108));
Q_MX03 U1343 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[96]), .A1(seed[96]), .A2(n950), .Z(n1109));
Q_MX03 U1344 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[97]), .A1(seed[97]), .A2(n952), .Z(n1110));
Q_MX03 U1345 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[98]), .A1(seed[98]), .A2(n954), .Z(n1111));
Q_MX03 U1346 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[99]), .A1(seed[99]), .A2(n956), .Z(n1112));
Q_MX03 U1347 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[100]), .A1(seed[100]), .A2(n958), .Z(n1113));
Q_MX03 U1348 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[101]), .A1(seed[101]), .A2(n960), .Z(n1114));
Q_MX03 U1349 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[102]), .A1(seed[102]), .A2(n962), .Z(n1115));
Q_MX03 U1350 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[103]), .A1(seed[103]), .A2(n964), .Z(n1116));
Q_MX03 U1351 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[104]), .A1(seed[104]), .A2(n966), .Z(n1117));
Q_MX03 U1352 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[105]), .A1(seed[105]), .A2(n968), .Z(n1118));
Q_MX03 U1353 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[106]), .A1(seed[106]), .A2(n970), .Z(n1119));
Q_MX03 U1354 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[107]), .A1(seed[107]), .A2(n972), .Z(n1120));
Q_MX03 U1355 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[108]), .A1(seed[108]), .A2(n974), .Z(n1121));
Q_MX03 U1356 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[109]), .A1(seed[109]), .A2(n976), .Z(n1122));
Q_MX03 U1357 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[110]), .A1(seed[110]), .A2(n978), .Z(n1123));
Q_MX03 U1358 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[111]), .A1(seed[111]), .A2(n980), .Z(n1124));
Q_MX03 U1359 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[112]), .A1(seed[112]), .A2(n982), .Z(n1125));
Q_MX03 U1360 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[113]), .A1(seed[113]), .A2(n984), .Z(n1126));
Q_MX03 U1361 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[114]), .A1(seed[114]), .A2(n986), .Z(n1127));
Q_MX03 U1362 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[115]), .A1(seed[115]), .A2(n988), .Z(n1128));
Q_MX03 U1363 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[116]), .A1(seed[116]), .A2(n990), .Z(n1129));
Q_MX03 U1364 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[117]), .A1(seed[117]), .A2(n992), .Z(n1130));
Q_MX03 U1365 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[118]), .A1(seed[118]), .A2(n994), .Z(n1131));
Q_MX03 U1366 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[119]), .A1(seed[119]), .A2(n996), .Z(n1132));
Q_MX03 U1367 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[120]), .A1(seed[120]), .A2(n998), .Z(n1133));
Q_MX03 U1368 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[121]), .A1(seed[121]), .A2(n1000), .Z(n1134));
Q_MX03 U1369 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[122]), .A1(seed[122]), .A2(n1002), .Z(n1135));
Q_MX03 U1370 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[123]), .A1(seed[123]), .A2(n1004), .Z(n1136));
Q_MX03 U1371 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[124]), .A1(seed[124]), .A2(n1006), .Z(n1137));
Q_MX03 U1372 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[125]), .A1(seed[125]), .A2(n1008), .Z(n1138));
Q_MX03 U1373 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[126]), .A1(seed[126]), .A2(n1010), .Z(n1139));
Q_MX03 U1374 ( .S0(n497), .S1(n1144), .A0(AesCiphOutR[127]), .A1(seed[127]), .A2(n1012), .Z(n1140));
Q_AN02 U1375 ( .A0(KeyInVld), .A1(n496), .Z(n1144));
Q_OR02 U1376 ( .A0(n497), .A1(KeyInVld), .Z(n1141));
Q_AO21 U1377 ( .A0(n1142), .A1(n1143), .B0(n1141), .Z(n1145));
Q_AN02 U1378 ( .A0(AesCiphOutVldR), .A1(n755), .Z(n1143));
Q_AN02 U1379 ( .A0(out_count[2]), .A1(n345), .Z(n1142));
Q_AD01HF U1380 ( .A0(in_count[1]), .B0(in_count[0]), .S(n1147), .CO(n1148));
Q_XOR2 U1381 ( .A0(in_count[2]), .A1(n1148), .Z(n1149));
Q_AN03 U1382 ( .A0(n87), .A1(n1146), .A2(n1160), .Z(n1155));
Q_AN03 U1383 ( .A0(n87), .A1(n1147), .A2(n1160), .Z(n1156));
Q_AN03 U1384 ( .A0(n87), .A1(n1149), .A2(n1160), .Z(n1157));
Q_XOR2 U1385 ( .A0(out_count[2]), .A1(n756), .Z(n1151));
Q_AN03 U1386 ( .A0(n4), .A1(n755), .A2(n1160), .Z(n1152));
Q_AN03 U1387 ( .A0(n4), .A1(n1150), .A2(n1160), .Z(n1153));
Q_AN03 U1388 ( .A0(n4), .A1(n1151), .A2(n1160), .Z(n1154));
Q_OR02 U1389 ( .A0(CiphInVldR), .A1(n346), .Z(n1158));
Q_OR02 U1390 ( .A0(AesCiphOutVldR), .A1(n346), .Z(n1159));
Q_INV U1391 ( .A(n346), .Z(n1160));
Q_FDP4EP \out_count_REG[0] ( .CK(clk), .CE(n1159), .R(n1161), .D(n1152), .Q(out_count[0]));
Q_INV U1393 ( .A(rst_n), .Z(n1161));
Q_INV U1394 ( .A(out_count[0]), .Z(n755));
Q_FDP4EP \out_count_REG[1] ( .CK(clk), .CE(n1159), .R(n1161), .D(n1153), .Q(out_count[1]));
Q_INV U1396 ( .A(out_count[1]), .Z(n345));
Q_FDP4EP \out_count_REG[2] ( .CK(clk), .CE(n1159), .R(n1161), .D(n1154), .Q(out_count[2]));
Q_INV U1398 ( .A(out_count[2]), .Z(n3));
Q_FDP4EP \in_count_REG[0] ( .CK(clk), .CE(n1158), .R(n1161), .D(n1155), .Q(in_count[0]));
Q_INV U1400 ( .A(in_count[0]), .Z(n1146));
Q_FDP4EP \in_count_REG[1] ( .CK(clk), .CE(n1158), .R(n1161), .D(n1156), .Q(in_count[1]));
Q_FDP4EP \in_count_REG[2] ( .CK(clk), .CE(n1158), .R(n1161), .D(n1157), .Q(in_count[2]));
Q_INV U1403 ( .A(in_count[2]), .Z(n86));
Q_FDP4EP \internal_state_value_REG[0] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1013), .Q(internal_state_value[0]));
Q_INV U1405 ( .A(internal_state_value[0]), .Z(n759));
Q_FDP4EP \internal_state_value_REG[1] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1014), .Q(internal_state_value[1]));
Q_FDP4EP \internal_state_value_REG[2] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1015), .Q(internal_state_value[2]));
Q_FDP4EP \internal_state_value_REG[3] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1016), .Q(internal_state_value[3]));
Q_FDP4EP \internal_state_value_REG[4] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1017), .Q(internal_state_value[4]));
Q_FDP4EP \internal_state_value_REG[5] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1018), .Q(internal_state_value[5]));
Q_FDP4EP \internal_state_value_REG[6] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1019), .Q(internal_state_value[6]));
Q_FDP4EP \internal_state_value_REG[7] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1020), .Q(internal_state_value[7]));
Q_FDP4EP \internal_state_value_REG[8] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1021), .Q(internal_state_value[8]));
Q_FDP4EP \internal_state_value_REG[9] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1022), .Q(internal_state_value[9]));
Q_FDP4EP \internal_state_value_REG[10] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1023), .Q(internal_state_value[10]));
Q_FDP4EP \internal_state_value_REG[11] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1024), .Q(internal_state_value[11]));
Q_FDP4EP \internal_state_value_REG[12] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1025), .Q(internal_state_value[12]));
Q_FDP4EP \internal_state_value_REG[13] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1026), .Q(internal_state_value[13]));
Q_FDP4EP \internal_state_value_REG[14] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1027), .Q(internal_state_value[14]));
Q_FDP4EP \internal_state_value_REG[15] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1028), .Q(internal_state_value[15]));
Q_FDP4EP \internal_state_value_REG[16] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1029), .Q(internal_state_value[16]));
Q_FDP4EP \internal_state_value_REG[17] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1030), .Q(internal_state_value[17]));
Q_FDP4EP \internal_state_value_REG[18] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1031), .Q(internal_state_value[18]));
Q_FDP4EP \internal_state_value_REG[19] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1032), .Q(internal_state_value[19]));
Q_FDP4EP \internal_state_value_REG[20] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1033), .Q(internal_state_value[20]));
Q_FDP4EP \internal_state_value_REG[21] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1034), .Q(internal_state_value[21]));
Q_FDP4EP \internal_state_value_REG[22] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1035), .Q(internal_state_value[22]));
Q_FDP4EP \internal_state_value_REG[23] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1036), .Q(internal_state_value[23]));
Q_FDP4EP \internal_state_value_REG[24] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1037), .Q(internal_state_value[24]));
Q_FDP4EP \internal_state_value_REG[25] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1038), .Q(internal_state_value[25]));
Q_FDP4EP \internal_state_value_REG[26] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1039), .Q(internal_state_value[26]));
Q_FDP4EP \internal_state_value_REG[27] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1040), .Q(internal_state_value[27]));
Q_FDP4EP \internal_state_value_REG[28] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1041), .Q(internal_state_value[28]));
Q_FDP4EP \internal_state_value_REG[29] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1042), .Q(internal_state_value[29]));
Q_FDP4EP \internal_state_value_REG[30] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1043), .Q(internal_state_value[30]));
Q_FDP4EP \internal_state_value_REG[31] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1044), .Q(internal_state_value[31]));
Q_FDP4EP \internal_state_value_REG[32] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1045), .Q(internal_state_value[32]));
Q_FDP4EP \internal_state_value_REG[33] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1046), .Q(internal_state_value[33]));
Q_FDP4EP \internal_state_value_REG[34] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1047), .Q(internal_state_value[34]));
Q_FDP4EP \internal_state_value_REG[35] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1048), .Q(internal_state_value[35]));
Q_FDP4EP \internal_state_value_REG[36] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1049), .Q(internal_state_value[36]));
Q_FDP4EP \internal_state_value_REG[37] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1050), .Q(internal_state_value[37]));
Q_FDP4EP \internal_state_value_REG[38] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1051), .Q(internal_state_value[38]));
Q_FDP4EP \internal_state_value_REG[39] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1052), .Q(internal_state_value[39]));
Q_FDP4EP \internal_state_value_REG[40] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1053), .Q(internal_state_value[40]));
Q_FDP4EP \internal_state_value_REG[41] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1054), .Q(internal_state_value[41]));
Q_FDP4EP \internal_state_value_REG[42] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1055), .Q(internal_state_value[42]));
Q_FDP4EP \internal_state_value_REG[43] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1056), .Q(internal_state_value[43]));
Q_FDP4EP \internal_state_value_REG[44] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1057), .Q(internal_state_value[44]));
Q_FDP4EP \internal_state_value_REG[45] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1058), .Q(internal_state_value[45]));
Q_FDP4EP \internal_state_value_REG[46] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1059), .Q(internal_state_value[46]));
Q_FDP4EP \internal_state_value_REG[47] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1060), .Q(internal_state_value[47]));
Q_FDP4EP \internal_state_value_REG[48] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1061), .Q(internal_state_value[48]));
Q_FDP4EP \internal_state_value_REG[49] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1062), .Q(internal_state_value[49]));
Q_FDP4EP \internal_state_value_REG[50] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1063), .Q(internal_state_value[50]));
Q_FDP4EP \internal_state_value_REG[51] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1064), .Q(internal_state_value[51]));
Q_FDP4EP \internal_state_value_REG[52] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1065), .Q(internal_state_value[52]));
Q_FDP4EP \internal_state_value_REG[53] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1066), .Q(internal_state_value[53]));
Q_FDP4EP \internal_state_value_REG[54] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1067), .Q(internal_state_value[54]));
Q_FDP4EP \internal_state_value_REG[55] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1068), .Q(internal_state_value[55]));
Q_FDP4EP \internal_state_value_REG[56] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1069), .Q(internal_state_value[56]));
Q_FDP4EP \internal_state_value_REG[57] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1070), .Q(internal_state_value[57]));
Q_FDP4EP \internal_state_value_REG[58] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1071), .Q(internal_state_value[58]));
Q_FDP4EP \internal_state_value_REG[59] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1072), .Q(internal_state_value[59]));
Q_FDP4EP \internal_state_value_REG[60] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1073), .Q(internal_state_value[60]));
Q_FDP4EP \internal_state_value_REG[61] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1074), .Q(internal_state_value[61]));
Q_FDP4EP \internal_state_value_REG[62] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1075), .Q(internal_state_value[62]));
Q_FDP4EP \internal_state_value_REG[63] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1076), .Q(internal_state_value[63]));
Q_FDP4EP \internal_state_value_REG[64] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1077), .Q(internal_state_value[64]));
Q_FDP4EP \internal_state_value_REG[65] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1078), .Q(internal_state_value[65]));
Q_FDP4EP \internal_state_value_REG[66] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1079), .Q(internal_state_value[66]));
Q_FDP4EP \internal_state_value_REG[67] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1080), .Q(internal_state_value[67]));
Q_FDP4EP \internal_state_value_REG[68] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1081), .Q(internal_state_value[68]));
Q_FDP4EP \internal_state_value_REG[69] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1082), .Q(internal_state_value[69]));
Q_FDP4EP \internal_state_value_REG[70] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1083), .Q(internal_state_value[70]));
Q_FDP4EP \internal_state_value_REG[71] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1084), .Q(internal_state_value[71]));
Q_FDP4EP \internal_state_value_REG[72] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1085), .Q(internal_state_value[72]));
Q_FDP4EP \internal_state_value_REG[73] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1086), .Q(internal_state_value[73]));
Q_FDP4EP \internal_state_value_REG[74] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1087), .Q(internal_state_value[74]));
Q_FDP4EP \internal_state_value_REG[75] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1088), .Q(internal_state_value[75]));
Q_FDP4EP \internal_state_value_REG[76] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1089), .Q(internal_state_value[76]));
Q_FDP4EP \internal_state_value_REG[77] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1090), .Q(internal_state_value[77]));
Q_FDP4EP \internal_state_value_REG[78] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1091), .Q(internal_state_value[78]));
Q_FDP4EP \internal_state_value_REG[79] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1092), .Q(internal_state_value[79]));
Q_FDP4EP \internal_state_value_REG[80] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1093), .Q(internal_state_value[80]));
Q_FDP4EP \internal_state_value_REG[81] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1094), .Q(internal_state_value[81]));
Q_FDP4EP \internal_state_value_REG[82] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1095), .Q(internal_state_value[82]));
Q_FDP4EP \internal_state_value_REG[83] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1096), .Q(internal_state_value[83]));
Q_FDP4EP \internal_state_value_REG[84] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1097), .Q(internal_state_value[84]));
Q_FDP4EP \internal_state_value_REG[85] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1098), .Q(internal_state_value[85]));
Q_FDP4EP \internal_state_value_REG[86] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1099), .Q(internal_state_value[86]));
Q_FDP4EP \internal_state_value_REG[87] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1100), .Q(internal_state_value[87]));
Q_FDP4EP \internal_state_value_REG[88] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1101), .Q(internal_state_value[88]));
Q_FDP4EP \internal_state_value_REG[89] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1102), .Q(internal_state_value[89]));
Q_FDP4EP \internal_state_value_REG[90] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1103), .Q(internal_state_value[90]));
Q_FDP4EP \internal_state_value_REG[91] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1104), .Q(internal_state_value[91]));
Q_FDP4EP \internal_state_value_REG[92] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1105), .Q(internal_state_value[92]));
Q_FDP4EP \internal_state_value_REG[93] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1106), .Q(internal_state_value[93]));
Q_FDP4EP \internal_state_value_REG[94] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1107), .Q(internal_state_value[94]));
Q_FDP4EP \internal_state_value_REG[95] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1108), .Q(internal_state_value[95]));
Q_FDP4EP \internal_state_value_REG[96] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1109), .Q(internal_state_value[96]));
Q_FDP4EP \internal_state_value_REG[97] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1110), .Q(internal_state_value[97]));
Q_FDP4EP \internal_state_value_REG[98] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1111), .Q(internal_state_value[98]));
Q_FDP4EP \internal_state_value_REG[99] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1112), .Q(internal_state_value[99]));
Q_FDP4EP \internal_state_value_REG[100] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1113), .Q(internal_state_value[100]));
Q_FDP4EP \internal_state_value_REG[101] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1114), .Q(internal_state_value[101]));
Q_FDP4EP \internal_state_value_REG[102] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1115), .Q(internal_state_value[102]));
Q_FDP4EP \internal_state_value_REG[103] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1116), .Q(internal_state_value[103]));
Q_FDP4EP \internal_state_value_REG[104] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1117), .Q(internal_state_value[104]));
Q_FDP4EP \internal_state_value_REG[105] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1118), .Q(internal_state_value[105]));
Q_FDP4EP \internal_state_value_REG[106] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1119), .Q(internal_state_value[106]));
Q_FDP4EP \internal_state_value_REG[107] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1120), .Q(internal_state_value[107]));
Q_FDP4EP \internal_state_value_REG[108] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1121), .Q(internal_state_value[108]));
Q_FDP4EP \internal_state_value_REG[109] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1122), .Q(internal_state_value[109]));
Q_FDP4EP \internal_state_value_REG[110] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1123), .Q(internal_state_value[110]));
Q_FDP4EP \internal_state_value_REG[111] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1124), .Q(internal_state_value[111]));
Q_FDP4EP \internal_state_value_REG[112] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1125), .Q(internal_state_value[112]));
Q_FDP4EP \internal_state_value_REG[113] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1126), .Q(internal_state_value[113]));
Q_FDP4EP \internal_state_value_REG[114] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1127), .Q(internal_state_value[114]));
Q_FDP4EP \internal_state_value_REG[115] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1128), .Q(internal_state_value[115]));
Q_FDP4EP \internal_state_value_REG[116] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1129), .Q(internal_state_value[116]));
Q_FDP4EP \internal_state_value_REG[117] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1130), .Q(internal_state_value[117]));
Q_FDP4EP \internal_state_value_REG[118] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1131), .Q(internal_state_value[118]));
Q_FDP4EP \internal_state_value_REG[119] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1132), .Q(internal_state_value[119]));
Q_FDP4EP \internal_state_value_REG[120] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1133), .Q(internal_state_value[120]));
Q_FDP4EP \internal_state_value_REG[121] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1134), .Q(internal_state_value[121]));
Q_FDP4EP \internal_state_value_REG[122] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1135), .Q(internal_state_value[122]));
Q_FDP4EP \internal_state_value_REG[123] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1136), .Q(internal_state_value[123]));
Q_FDP4EP \internal_state_value_REG[124] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1137), .Q(internal_state_value[124]));
Q_FDP4EP \internal_state_value_REG[125] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1138), .Q(internal_state_value[125]));
Q_FDP4EP \internal_state_value_REG[126] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1139), .Q(internal_state_value[126]));
Q_FDP4EP \internal_state_value_REG[127] ( .CK(clk), .CE(n1145), .R(n1161), .D(n1140), .Q(internal_state_value[127]));
Q_FDP4EP \internal_state_key_REG[0] ( .CK(clk), .CE(n758), .R(n1161), .D(n498), .Q(internal_state_key[0]));
Q_FDP4EP \internal_state_key_REG[1] ( .CK(clk), .CE(n758), .R(n1161), .D(n499), .Q(internal_state_key[1]));
Q_FDP4EP \internal_state_key_REG[2] ( .CK(clk), .CE(n758), .R(n1161), .D(n500), .Q(internal_state_key[2]));
Q_FDP4EP \internal_state_key_REG[3] ( .CK(clk), .CE(n758), .R(n1161), .D(n501), .Q(internal_state_key[3]));
Q_FDP4EP \internal_state_key_REG[4] ( .CK(clk), .CE(n758), .R(n1161), .D(n502), .Q(internal_state_key[4]));
Q_FDP4EP \internal_state_key_REG[5] ( .CK(clk), .CE(n758), .R(n1161), .D(n503), .Q(internal_state_key[5]));
Q_FDP4EP \internal_state_key_REG[6] ( .CK(clk), .CE(n758), .R(n1161), .D(n504), .Q(internal_state_key[6]));
Q_FDP4EP \internal_state_key_REG[7] ( .CK(clk), .CE(n758), .R(n1161), .D(n505), .Q(internal_state_key[7]));
Q_FDP4EP \internal_state_key_REG[8] ( .CK(clk), .CE(n758), .R(n1161), .D(n506), .Q(internal_state_key[8]));
Q_FDP4EP \internal_state_key_REG[9] ( .CK(clk), .CE(n758), .R(n1161), .D(n507), .Q(internal_state_key[9]));
Q_FDP4EP \internal_state_key_REG[10] ( .CK(clk), .CE(n758), .R(n1161), .D(n508), .Q(internal_state_key[10]));
Q_FDP4EP \internal_state_key_REG[11] ( .CK(clk), .CE(n758), .R(n1161), .D(n509), .Q(internal_state_key[11]));
Q_FDP4EP \internal_state_key_REG[12] ( .CK(clk), .CE(n758), .R(n1161), .D(n510), .Q(internal_state_key[12]));
Q_FDP4EP \internal_state_key_REG[13] ( .CK(clk), .CE(n758), .R(n1161), .D(n511), .Q(internal_state_key[13]));
Q_FDP4EP \internal_state_key_REG[14] ( .CK(clk), .CE(n758), .R(n1161), .D(n512), .Q(internal_state_key[14]));
Q_FDP4EP \internal_state_key_REG[15] ( .CK(clk), .CE(n758), .R(n1161), .D(n513), .Q(internal_state_key[15]));
Q_FDP4EP \internal_state_key_REG[16] ( .CK(clk), .CE(n758), .R(n1161), .D(n514), .Q(internal_state_key[16]));
Q_FDP4EP \internal_state_key_REG[17] ( .CK(clk), .CE(n758), .R(n1161), .D(n515), .Q(internal_state_key[17]));
Q_FDP4EP \internal_state_key_REG[18] ( .CK(clk), .CE(n758), .R(n1161), .D(n516), .Q(internal_state_key[18]));
Q_FDP4EP \internal_state_key_REG[19] ( .CK(clk), .CE(n758), .R(n1161), .D(n517), .Q(internal_state_key[19]));
Q_FDP4EP \internal_state_key_REG[20] ( .CK(clk), .CE(n758), .R(n1161), .D(n518), .Q(internal_state_key[20]));
Q_FDP4EP \internal_state_key_REG[21] ( .CK(clk), .CE(n758), .R(n1161), .D(n519), .Q(internal_state_key[21]));
Q_FDP4EP \internal_state_key_REG[22] ( .CK(clk), .CE(n758), .R(n1161), .D(n520), .Q(internal_state_key[22]));
Q_FDP4EP \internal_state_key_REG[23] ( .CK(clk), .CE(n758), .R(n1161), .D(n521), .Q(internal_state_key[23]));
Q_FDP4EP \internal_state_key_REG[24] ( .CK(clk), .CE(n758), .R(n1161), .D(n522), .Q(internal_state_key[24]));
Q_FDP4EP \internal_state_key_REG[25] ( .CK(clk), .CE(n758), .R(n1161), .D(n523), .Q(internal_state_key[25]));
Q_FDP4EP \internal_state_key_REG[26] ( .CK(clk), .CE(n758), .R(n1161), .D(n524), .Q(internal_state_key[26]));
Q_FDP4EP \internal_state_key_REG[27] ( .CK(clk), .CE(n758), .R(n1161), .D(n525), .Q(internal_state_key[27]));
Q_FDP4EP \internal_state_key_REG[28] ( .CK(clk), .CE(n758), .R(n1161), .D(n526), .Q(internal_state_key[28]));
Q_FDP4EP \internal_state_key_REG[29] ( .CK(clk), .CE(n758), .R(n1161), .D(n527), .Q(internal_state_key[29]));
Q_FDP4EP \internal_state_key_REG[30] ( .CK(clk), .CE(n758), .R(n1161), .D(n528), .Q(internal_state_key[30]));
Q_FDP4EP \internal_state_key_REG[31] ( .CK(clk), .CE(n758), .R(n1161), .D(n529), .Q(internal_state_key[31]));
Q_FDP4EP \internal_state_key_REG[32] ( .CK(clk), .CE(n758), .R(n1161), .D(n530), .Q(internal_state_key[32]));
Q_FDP4EP \internal_state_key_REG[33] ( .CK(clk), .CE(n758), .R(n1161), .D(n531), .Q(internal_state_key[33]));
Q_FDP4EP \internal_state_key_REG[34] ( .CK(clk), .CE(n758), .R(n1161), .D(n532), .Q(internal_state_key[34]));
Q_FDP4EP \internal_state_key_REG[35] ( .CK(clk), .CE(n758), .R(n1161), .D(n533), .Q(internal_state_key[35]));
Q_FDP4EP \internal_state_key_REG[36] ( .CK(clk), .CE(n758), .R(n1161), .D(n534), .Q(internal_state_key[36]));
Q_FDP4EP \internal_state_key_REG[37] ( .CK(clk), .CE(n758), .R(n1161), .D(n535), .Q(internal_state_key[37]));
Q_FDP4EP \internal_state_key_REG[38] ( .CK(clk), .CE(n758), .R(n1161), .D(n536), .Q(internal_state_key[38]));
Q_FDP4EP \internal_state_key_REG[39] ( .CK(clk), .CE(n758), .R(n1161), .D(n537), .Q(internal_state_key[39]));
Q_FDP4EP \internal_state_key_REG[40] ( .CK(clk), .CE(n758), .R(n1161), .D(n538), .Q(internal_state_key[40]));
Q_FDP4EP \internal_state_key_REG[41] ( .CK(clk), .CE(n758), .R(n1161), .D(n539), .Q(internal_state_key[41]));
Q_FDP4EP \internal_state_key_REG[42] ( .CK(clk), .CE(n758), .R(n1161), .D(n540), .Q(internal_state_key[42]));
Q_FDP4EP \internal_state_key_REG[43] ( .CK(clk), .CE(n758), .R(n1161), .D(n541), .Q(internal_state_key[43]));
Q_FDP4EP \internal_state_key_REG[44] ( .CK(clk), .CE(n758), .R(n1161), .D(n542), .Q(internal_state_key[44]));
Q_FDP4EP \internal_state_key_REG[45] ( .CK(clk), .CE(n758), .R(n1161), .D(n543), .Q(internal_state_key[45]));
Q_FDP4EP \internal_state_key_REG[46] ( .CK(clk), .CE(n758), .R(n1161), .D(n544), .Q(internal_state_key[46]));
Q_FDP4EP \internal_state_key_REG[47] ( .CK(clk), .CE(n758), .R(n1161), .D(n545), .Q(internal_state_key[47]));
Q_FDP4EP \internal_state_key_REG[48] ( .CK(clk), .CE(n758), .R(n1161), .D(n546), .Q(internal_state_key[48]));
Q_FDP4EP \internal_state_key_REG[49] ( .CK(clk), .CE(n758), .R(n1161), .D(n547), .Q(internal_state_key[49]));
Q_FDP4EP \internal_state_key_REG[50] ( .CK(clk), .CE(n758), .R(n1161), .D(n548), .Q(internal_state_key[50]));
Q_FDP4EP \internal_state_key_REG[51] ( .CK(clk), .CE(n758), .R(n1161), .D(n549), .Q(internal_state_key[51]));
Q_FDP4EP \internal_state_key_REG[52] ( .CK(clk), .CE(n758), .R(n1161), .D(n550), .Q(internal_state_key[52]));
Q_FDP4EP \internal_state_key_REG[53] ( .CK(clk), .CE(n758), .R(n1161), .D(n551), .Q(internal_state_key[53]));
Q_FDP4EP \internal_state_key_REG[54] ( .CK(clk), .CE(n758), .R(n1161), .D(n552), .Q(internal_state_key[54]));
Q_FDP4EP \internal_state_key_REG[55] ( .CK(clk), .CE(n758), .R(n1161), .D(n553), .Q(internal_state_key[55]));
Q_FDP4EP \internal_state_key_REG[56] ( .CK(clk), .CE(n758), .R(n1161), .D(n554), .Q(internal_state_key[56]));
Q_FDP4EP \internal_state_key_REG[57] ( .CK(clk), .CE(n758), .R(n1161), .D(n555), .Q(internal_state_key[57]));
Q_FDP4EP \internal_state_key_REG[58] ( .CK(clk), .CE(n758), .R(n1161), .D(n556), .Q(internal_state_key[58]));
Q_FDP4EP \internal_state_key_REG[59] ( .CK(clk), .CE(n758), .R(n1161), .D(n557), .Q(internal_state_key[59]));
Q_FDP4EP \internal_state_key_REG[60] ( .CK(clk), .CE(n758), .R(n1161), .D(n558), .Q(internal_state_key[60]));
Q_FDP4EP \internal_state_key_REG[61] ( .CK(clk), .CE(n758), .R(n1161), .D(n559), .Q(internal_state_key[61]));
Q_FDP4EP \internal_state_key_REG[62] ( .CK(clk), .CE(n758), .R(n1161), .D(n560), .Q(internal_state_key[62]));
Q_FDP4EP \internal_state_key_REG[63] ( .CK(clk), .CE(n758), .R(n1161), .D(n561), .Q(internal_state_key[63]));
Q_FDP4EP \internal_state_key_REG[64] ( .CK(clk), .CE(n758), .R(n1161), .D(n562), .Q(internal_state_key[64]));
Q_FDP4EP \internal_state_key_REG[65] ( .CK(clk), .CE(n758), .R(n1161), .D(n563), .Q(internal_state_key[65]));
Q_FDP4EP \internal_state_key_REG[66] ( .CK(clk), .CE(n758), .R(n1161), .D(n564), .Q(internal_state_key[66]));
Q_FDP4EP \internal_state_key_REG[67] ( .CK(clk), .CE(n758), .R(n1161), .D(n565), .Q(internal_state_key[67]));
Q_FDP4EP \internal_state_key_REG[68] ( .CK(clk), .CE(n758), .R(n1161), .D(n566), .Q(internal_state_key[68]));
Q_FDP4EP \internal_state_key_REG[69] ( .CK(clk), .CE(n758), .R(n1161), .D(n567), .Q(internal_state_key[69]));
Q_FDP4EP \internal_state_key_REG[70] ( .CK(clk), .CE(n758), .R(n1161), .D(n568), .Q(internal_state_key[70]));
Q_FDP4EP \internal_state_key_REG[71] ( .CK(clk), .CE(n758), .R(n1161), .D(n569), .Q(internal_state_key[71]));
Q_FDP4EP \internal_state_key_REG[72] ( .CK(clk), .CE(n758), .R(n1161), .D(n570), .Q(internal_state_key[72]));
Q_FDP4EP \internal_state_key_REG[73] ( .CK(clk), .CE(n758), .R(n1161), .D(n571), .Q(internal_state_key[73]));
Q_FDP4EP \internal_state_key_REG[74] ( .CK(clk), .CE(n758), .R(n1161), .D(n572), .Q(internal_state_key[74]));
Q_FDP4EP \internal_state_key_REG[75] ( .CK(clk), .CE(n758), .R(n1161), .D(n573), .Q(internal_state_key[75]));
Q_FDP4EP \internal_state_key_REG[76] ( .CK(clk), .CE(n758), .R(n1161), .D(n574), .Q(internal_state_key[76]));
Q_FDP4EP \internal_state_key_REG[77] ( .CK(clk), .CE(n758), .R(n1161), .D(n575), .Q(internal_state_key[77]));
Q_FDP4EP \internal_state_key_REG[78] ( .CK(clk), .CE(n758), .R(n1161), .D(n576), .Q(internal_state_key[78]));
Q_FDP4EP \internal_state_key_REG[79] ( .CK(clk), .CE(n758), .R(n1161), .D(n577), .Q(internal_state_key[79]));
Q_FDP4EP \internal_state_key_REG[80] ( .CK(clk), .CE(n758), .R(n1161), .D(n578), .Q(internal_state_key[80]));
Q_FDP4EP \internal_state_key_REG[81] ( .CK(clk), .CE(n758), .R(n1161), .D(n579), .Q(internal_state_key[81]));
Q_FDP4EP \internal_state_key_REG[82] ( .CK(clk), .CE(n758), .R(n1161), .D(n580), .Q(internal_state_key[82]));
Q_FDP4EP \internal_state_key_REG[83] ( .CK(clk), .CE(n758), .R(n1161), .D(n581), .Q(internal_state_key[83]));
Q_FDP4EP \internal_state_key_REG[84] ( .CK(clk), .CE(n758), .R(n1161), .D(n582), .Q(internal_state_key[84]));
Q_FDP4EP \internal_state_key_REG[85] ( .CK(clk), .CE(n758), .R(n1161), .D(n583), .Q(internal_state_key[85]));
Q_FDP4EP \internal_state_key_REG[86] ( .CK(clk), .CE(n758), .R(n1161), .D(n584), .Q(internal_state_key[86]));
Q_FDP4EP \internal_state_key_REG[87] ( .CK(clk), .CE(n758), .R(n1161), .D(n585), .Q(internal_state_key[87]));
Q_FDP4EP \internal_state_key_REG[88] ( .CK(clk), .CE(n758), .R(n1161), .D(n586), .Q(internal_state_key[88]));
Q_FDP4EP \internal_state_key_REG[89] ( .CK(clk), .CE(n758), .R(n1161), .D(n587), .Q(internal_state_key[89]));
Q_FDP4EP \internal_state_key_REG[90] ( .CK(clk), .CE(n758), .R(n1161), .D(n588), .Q(internal_state_key[90]));
Q_FDP4EP \internal_state_key_REG[91] ( .CK(clk), .CE(n758), .R(n1161), .D(n589), .Q(internal_state_key[91]));
Q_FDP4EP \internal_state_key_REG[92] ( .CK(clk), .CE(n758), .R(n1161), .D(n590), .Q(internal_state_key[92]));
Q_FDP4EP \internal_state_key_REG[93] ( .CK(clk), .CE(n758), .R(n1161), .D(n591), .Q(internal_state_key[93]));
Q_FDP4EP \internal_state_key_REG[94] ( .CK(clk), .CE(n758), .R(n1161), .D(n592), .Q(internal_state_key[94]));
Q_FDP4EP \internal_state_key_REG[95] ( .CK(clk), .CE(n758), .R(n1161), .D(n593), .Q(internal_state_key[95]));
Q_FDP4EP \internal_state_key_REG[96] ( .CK(clk), .CE(n758), .R(n1161), .D(n594), .Q(internal_state_key[96]));
Q_FDP4EP \internal_state_key_REG[97] ( .CK(clk), .CE(n758), .R(n1161), .D(n595), .Q(internal_state_key[97]));
Q_FDP4EP \internal_state_key_REG[98] ( .CK(clk), .CE(n758), .R(n1161), .D(n596), .Q(internal_state_key[98]));
Q_FDP4EP \internal_state_key_REG[99] ( .CK(clk), .CE(n758), .R(n1161), .D(n597), .Q(internal_state_key[99]));
Q_FDP4EP \internal_state_key_REG[100] ( .CK(clk), .CE(n758), .R(n1161), .D(n598), .Q(internal_state_key[100]));
Q_FDP4EP \internal_state_key_REG[101] ( .CK(clk), .CE(n758), .R(n1161), .D(n599), .Q(internal_state_key[101]));
Q_FDP4EP \internal_state_key_REG[102] ( .CK(clk), .CE(n758), .R(n1161), .D(n600), .Q(internal_state_key[102]));
Q_FDP4EP \internal_state_key_REG[103] ( .CK(clk), .CE(n758), .R(n1161), .D(n601), .Q(internal_state_key[103]));
Q_FDP4EP \internal_state_key_REG[104] ( .CK(clk), .CE(n758), .R(n1161), .D(n602), .Q(internal_state_key[104]));
Q_FDP4EP \internal_state_key_REG[105] ( .CK(clk), .CE(n758), .R(n1161), .D(n603), .Q(internal_state_key[105]));
Q_FDP4EP \internal_state_key_REG[106] ( .CK(clk), .CE(n758), .R(n1161), .D(n604), .Q(internal_state_key[106]));
Q_FDP4EP \internal_state_key_REG[107] ( .CK(clk), .CE(n758), .R(n1161), .D(n605), .Q(internal_state_key[107]));
Q_FDP4EP \internal_state_key_REG[108] ( .CK(clk), .CE(n758), .R(n1161), .D(n606), .Q(internal_state_key[108]));
Q_FDP4EP \internal_state_key_REG[109] ( .CK(clk), .CE(n758), .R(n1161), .D(n607), .Q(internal_state_key[109]));
Q_FDP4EP \internal_state_key_REG[110] ( .CK(clk), .CE(n758), .R(n1161), .D(n608), .Q(internal_state_key[110]));
Q_FDP4EP \internal_state_key_REG[111] ( .CK(clk), .CE(n758), .R(n1161), .D(n609), .Q(internal_state_key[111]));
Q_FDP4EP \internal_state_key_REG[112] ( .CK(clk), .CE(n758), .R(n1161), .D(n610), .Q(internal_state_key[112]));
Q_FDP4EP \internal_state_key_REG[113] ( .CK(clk), .CE(n758), .R(n1161), .D(n611), .Q(internal_state_key[113]));
Q_FDP4EP \internal_state_key_REG[114] ( .CK(clk), .CE(n758), .R(n1161), .D(n612), .Q(internal_state_key[114]));
Q_FDP4EP \internal_state_key_REG[115] ( .CK(clk), .CE(n758), .R(n1161), .D(n613), .Q(internal_state_key[115]));
Q_FDP4EP \internal_state_key_REG[116] ( .CK(clk), .CE(n758), .R(n1161), .D(n614), .Q(internal_state_key[116]));
Q_FDP4EP \internal_state_key_REG[117] ( .CK(clk), .CE(n758), .R(n1161), .D(n615), .Q(internal_state_key[117]));
Q_FDP4EP \internal_state_key_REG[118] ( .CK(clk), .CE(n758), .R(n1161), .D(n616), .Q(internal_state_key[118]));
Q_FDP4EP \internal_state_key_REG[119] ( .CK(clk), .CE(n758), .R(n1161), .D(n617), .Q(internal_state_key[119]));
Q_FDP4EP \internal_state_key_REG[120] ( .CK(clk), .CE(n758), .R(n1161), .D(n618), .Q(internal_state_key[120]));
Q_FDP4EP \internal_state_key_REG[121] ( .CK(clk), .CE(n758), .R(n1161), .D(n619), .Q(internal_state_key[121]));
Q_FDP4EP \internal_state_key_REG[122] ( .CK(clk), .CE(n758), .R(n1161), .D(n620), .Q(internal_state_key[122]));
Q_FDP4EP \internal_state_key_REG[123] ( .CK(clk), .CE(n758), .R(n1161), .D(n621), .Q(internal_state_key[123]));
Q_FDP4EP \internal_state_key_REG[124] ( .CK(clk), .CE(n758), .R(n1161), .D(n622), .Q(internal_state_key[124]));
Q_FDP4EP \internal_state_key_REG[125] ( .CK(clk), .CE(n758), .R(n1161), .D(n623), .Q(internal_state_key[125]));
Q_FDP4EP \internal_state_key_REG[126] ( .CK(clk), .CE(n758), .R(n1161), .D(n624), .Q(internal_state_key[126]));
Q_FDP4EP \internal_state_key_REG[127] ( .CK(clk), .CE(n758), .R(n1161), .D(n625), .Q(internal_state_key[127]));
Q_FDP4EP \internal_state_key_REG[128] ( .CK(clk), .CE(n757), .R(n1161), .D(n626), .Q(internal_state_key[128]));
Q_FDP4EP \internal_state_key_REG[129] ( .CK(clk), .CE(n757), .R(n1161), .D(n627), .Q(internal_state_key[129]));
Q_FDP4EP \internal_state_key_REG[130] ( .CK(clk), .CE(n757), .R(n1161), .D(n628), .Q(internal_state_key[130]));
Q_FDP4EP \internal_state_key_REG[131] ( .CK(clk), .CE(n757), .R(n1161), .D(n629), .Q(internal_state_key[131]));
Q_FDP4EP \internal_state_key_REG[132] ( .CK(clk), .CE(n757), .R(n1161), .D(n630), .Q(internal_state_key[132]));
Q_FDP4EP \internal_state_key_REG[133] ( .CK(clk), .CE(n757), .R(n1161), .D(n631), .Q(internal_state_key[133]));
Q_FDP4EP \internal_state_key_REG[134] ( .CK(clk), .CE(n757), .R(n1161), .D(n632), .Q(internal_state_key[134]));
Q_FDP4EP \internal_state_key_REG[135] ( .CK(clk), .CE(n757), .R(n1161), .D(n633), .Q(internal_state_key[135]));
Q_FDP4EP \internal_state_key_REG[136] ( .CK(clk), .CE(n757), .R(n1161), .D(n634), .Q(internal_state_key[136]));
Q_FDP4EP \internal_state_key_REG[137] ( .CK(clk), .CE(n757), .R(n1161), .D(n635), .Q(internal_state_key[137]));
Q_FDP4EP \internal_state_key_REG[138] ( .CK(clk), .CE(n757), .R(n1161), .D(n636), .Q(internal_state_key[138]));
Q_FDP4EP \internal_state_key_REG[139] ( .CK(clk), .CE(n757), .R(n1161), .D(n637), .Q(internal_state_key[139]));
Q_FDP4EP \internal_state_key_REG[140] ( .CK(clk), .CE(n757), .R(n1161), .D(n638), .Q(internal_state_key[140]));
Q_FDP4EP \internal_state_key_REG[141] ( .CK(clk), .CE(n757), .R(n1161), .D(n639), .Q(internal_state_key[141]));
Q_FDP4EP \internal_state_key_REG[142] ( .CK(clk), .CE(n757), .R(n1161), .D(n640), .Q(internal_state_key[142]));
Q_FDP4EP \internal_state_key_REG[143] ( .CK(clk), .CE(n757), .R(n1161), .D(n641), .Q(internal_state_key[143]));
Q_FDP4EP \internal_state_key_REG[144] ( .CK(clk), .CE(n757), .R(n1161), .D(n642), .Q(internal_state_key[144]));
Q_FDP4EP \internal_state_key_REG[145] ( .CK(clk), .CE(n757), .R(n1161), .D(n643), .Q(internal_state_key[145]));
Q_FDP4EP \internal_state_key_REG[146] ( .CK(clk), .CE(n757), .R(n1161), .D(n644), .Q(internal_state_key[146]));
Q_FDP4EP \internal_state_key_REG[147] ( .CK(clk), .CE(n757), .R(n1161), .D(n645), .Q(internal_state_key[147]));
Q_FDP4EP \internal_state_key_REG[148] ( .CK(clk), .CE(n757), .R(n1161), .D(n646), .Q(internal_state_key[148]));
Q_FDP4EP \internal_state_key_REG[149] ( .CK(clk), .CE(n757), .R(n1161), .D(n647), .Q(internal_state_key[149]));
Q_FDP4EP \internal_state_key_REG[150] ( .CK(clk), .CE(n757), .R(n1161), .D(n648), .Q(internal_state_key[150]));
Q_FDP4EP \internal_state_key_REG[151] ( .CK(clk), .CE(n757), .R(n1161), .D(n649), .Q(internal_state_key[151]));
Q_FDP4EP \internal_state_key_REG[152] ( .CK(clk), .CE(n757), .R(n1161), .D(n650), .Q(internal_state_key[152]));
Q_FDP4EP \internal_state_key_REG[153] ( .CK(clk), .CE(n757), .R(n1161), .D(n651), .Q(internal_state_key[153]));
Q_FDP4EP \internal_state_key_REG[154] ( .CK(clk), .CE(n757), .R(n1161), .D(n652), .Q(internal_state_key[154]));
Q_FDP4EP \internal_state_key_REG[155] ( .CK(clk), .CE(n757), .R(n1161), .D(n653), .Q(internal_state_key[155]));
Q_FDP4EP \internal_state_key_REG[156] ( .CK(clk), .CE(n757), .R(n1161), .D(n654), .Q(internal_state_key[156]));
Q_FDP4EP \internal_state_key_REG[157] ( .CK(clk), .CE(n757), .R(n1161), .D(n655), .Q(internal_state_key[157]));
Q_FDP4EP \internal_state_key_REG[158] ( .CK(clk), .CE(n757), .R(n1161), .D(n656), .Q(internal_state_key[158]));
Q_FDP4EP \internal_state_key_REG[159] ( .CK(clk), .CE(n757), .R(n1161), .D(n657), .Q(internal_state_key[159]));
Q_FDP4EP \internal_state_key_REG[160] ( .CK(clk), .CE(n757), .R(n1161), .D(n658), .Q(internal_state_key[160]));
Q_FDP4EP \internal_state_key_REG[161] ( .CK(clk), .CE(n757), .R(n1161), .D(n659), .Q(internal_state_key[161]));
Q_FDP4EP \internal_state_key_REG[162] ( .CK(clk), .CE(n757), .R(n1161), .D(n660), .Q(internal_state_key[162]));
Q_FDP4EP \internal_state_key_REG[163] ( .CK(clk), .CE(n757), .R(n1161), .D(n661), .Q(internal_state_key[163]));
Q_FDP4EP \internal_state_key_REG[164] ( .CK(clk), .CE(n757), .R(n1161), .D(n662), .Q(internal_state_key[164]));
Q_FDP4EP \internal_state_key_REG[165] ( .CK(clk), .CE(n757), .R(n1161), .D(n663), .Q(internal_state_key[165]));
Q_FDP4EP \internal_state_key_REG[166] ( .CK(clk), .CE(n757), .R(n1161), .D(n664), .Q(internal_state_key[166]));
Q_FDP4EP \internal_state_key_REG[167] ( .CK(clk), .CE(n757), .R(n1161), .D(n665), .Q(internal_state_key[167]));
Q_FDP4EP \internal_state_key_REG[168] ( .CK(clk), .CE(n757), .R(n1161), .D(n666), .Q(internal_state_key[168]));
Q_FDP4EP \internal_state_key_REG[169] ( .CK(clk), .CE(n757), .R(n1161), .D(n667), .Q(internal_state_key[169]));
Q_FDP4EP \internal_state_key_REG[170] ( .CK(clk), .CE(n757), .R(n1161), .D(n668), .Q(internal_state_key[170]));
Q_FDP4EP \internal_state_key_REG[171] ( .CK(clk), .CE(n757), .R(n1161), .D(n669), .Q(internal_state_key[171]));
Q_FDP4EP \internal_state_key_REG[172] ( .CK(clk), .CE(n757), .R(n1161), .D(n670), .Q(internal_state_key[172]));
Q_FDP4EP \internal_state_key_REG[173] ( .CK(clk), .CE(n757), .R(n1161), .D(n671), .Q(internal_state_key[173]));
Q_FDP4EP \internal_state_key_REG[174] ( .CK(clk), .CE(n757), .R(n1161), .D(n672), .Q(internal_state_key[174]));
Q_FDP4EP \internal_state_key_REG[175] ( .CK(clk), .CE(n757), .R(n1161), .D(n673), .Q(internal_state_key[175]));
Q_FDP4EP \internal_state_key_REG[176] ( .CK(clk), .CE(n757), .R(n1161), .D(n674), .Q(internal_state_key[176]));
Q_FDP4EP \internal_state_key_REG[177] ( .CK(clk), .CE(n757), .R(n1161), .D(n675), .Q(internal_state_key[177]));
Q_FDP4EP \internal_state_key_REG[178] ( .CK(clk), .CE(n757), .R(n1161), .D(n676), .Q(internal_state_key[178]));
Q_FDP4EP \internal_state_key_REG[179] ( .CK(clk), .CE(n757), .R(n1161), .D(n677), .Q(internal_state_key[179]));
Q_FDP4EP \internal_state_key_REG[180] ( .CK(clk), .CE(n757), .R(n1161), .D(n678), .Q(internal_state_key[180]));
Q_FDP4EP \internal_state_key_REG[181] ( .CK(clk), .CE(n757), .R(n1161), .D(n679), .Q(internal_state_key[181]));
Q_FDP4EP \internal_state_key_REG[182] ( .CK(clk), .CE(n757), .R(n1161), .D(n680), .Q(internal_state_key[182]));
Q_FDP4EP \internal_state_key_REG[183] ( .CK(clk), .CE(n757), .R(n1161), .D(n681), .Q(internal_state_key[183]));
Q_FDP4EP \internal_state_key_REG[184] ( .CK(clk), .CE(n757), .R(n1161), .D(n682), .Q(internal_state_key[184]));
Q_FDP4EP \internal_state_key_REG[185] ( .CK(clk), .CE(n757), .R(n1161), .D(n683), .Q(internal_state_key[185]));
Q_FDP4EP \internal_state_key_REG[186] ( .CK(clk), .CE(n757), .R(n1161), .D(n684), .Q(internal_state_key[186]));
Q_FDP4EP \internal_state_key_REG[187] ( .CK(clk), .CE(n757), .R(n1161), .D(n685), .Q(internal_state_key[187]));
Q_FDP4EP \internal_state_key_REG[188] ( .CK(clk), .CE(n757), .R(n1161), .D(n686), .Q(internal_state_key[188]));
Q_FDP4EP \internal_state_key_REG[189] ( .CK(clk), .CE(n757), .R(n1161), .D(n687), .Q(internal_state_key[189]));
Q_FDP4EP \internal_state_key_REG[190] ( .CK(clk), .CE(n757), .R(n1161), .D(n688), .Q(internal_state_key[190]));
Q_FDP4EP \internal_state_key_REG[191] ( .CK(clk), .CE(n757), .R(n1161), .D(n689), .Q(internal_state_key[191]));
Q_FDP4EP \internal_state_key_REG[192] ( .CK(clk), .CE(n757), .R(n1161), .D(n690), .Q(internal_state_key[192]));
Q_FDP4EP \internal_state_key_REG[193] ( .CK(clk), .CE(n757), .R(n1161), .D(n691), .Q(internal_state_key[193]));
Q_FDP4EP \internal_state_key_REG[194] ( .CK(clk), .CE(n757), .R(n1161), .D(n692), .Q(internal_state_key[194]));
Q_FDP4EP \internal_state_key_REG[195] ( .CK(clk), .CE(n757), .R(n1161), .D(n693), .Q(internal_state_key[195]));
Q_FDP4EP \internal_state_key_REG[196] ( .CK(clk), .CE(n757), .R(n1161), .D(n694), .Q(internal_state_key[196]));
Q_FDP4EP \internal_state_key_REG[197] ( .CK(clk), .CE(n757), .R(n1161), .D(n695), .Q(internal_state_key[197]));
Q_FDP4EP \internal_state_key_REG[198] ( .CK(clk), .CE(n757), .R(n1161), .D(n696), .Q(internal_state_key[198]));
Q_FDP4EP \internal_state_key_REG[199] ( .CK(clk), .CE(n757), .R(n1161), .D(n697), .Q(internal_state_key[199]));
Q_FDP4EP \internal_state_key_REG[200] ( .CK(clk), .CE(n757), .R(n1161), .D(n698), .Q(internal_state_key[200]));
Q_FDP4EP \internal_state_key_REG[201] ( .CK(clk), .CE(n757), .R(n1161), .D(n699), .Q(internal_state_key[201]));
Q_FDP4EP \internal_state_key_REG[202] ( .CK(clk), .CE(n757), .R(n1161), .D(n700), .Q(internal_state_key[202]));
Q_FDP4EP \internal_state_key_REG[203] ( .CK(clk), .CE(n757), .R(n1161), .D(n701), .Q(internal_state_key[203]));
Q_FDP4EP \internal_state_key_REG[204] ( .CK(clk), .CE(n757), .R(n1161), .D(n702), .Q(internal_state_key[204]));
Q_FDP4EP \internal_state_key_REG[205] ( .CK(clk), .CE(n757), .R(n1161), .D(n703), .Q(internal_state_key[205]));
Q_FDP4EP \internal_state_key_REG[206] ( .CK(clk), .CE(n757), .R(n1161), .D(n704), .Q(internal_state_key[206]));
Q_FDP4EP \internal_state_key_REG[207] ( .CK(clk), .CE(n757), .R(n1161), .D(n705), .Q(internal_state_key[207]));
Q_FDP4EP \internal_state_key_REG[208] ( .CK(clk), .CE(n757), .R(n1161), .D(n706), .Q(internal_state_key[208]));
Q_FDP4EP \internal_state_key_REG[209] ( .CK(clk), .CE(n757), .R(n1161), .D(n707), .Q(internal_state_key[209]));
Q_FDP4EP \internal_state_key_REG[210] ( .CK(clk), .CE(n757), .R(n1161), .D(n708), .Q(internal_state_key[210]));
Q_FDP4EP \internal_state_key_REG[211] ( .CK(clk), .CE(n757), .R(n1161), .D(n709), .Q(internal_state_key[211]));
Q_FDP4EP \internal_state_key_REG[212] ( .CK(clk), .CE(n757), .R(n1161), .D(n710), .Q(internal_state_key[212]));
Q_FDP4EP \internal_state_key_REG[213] ( .CK(clk), .CE(n757), .R(n1161), .D(n711), .Q(internal_state_key[213]));
Q_FDP4EP \internal_state_key_REG[214] ( .CK(clk), .CE(n757), .R(n1161), .D(n712), .Q(internal_state_key[214]));
Q_FDP4EP \internal_state_key_REG[215] ( .CK(clk), .CE(n757), .R(n1161), .D(n713), .Q(internal_state_key[215]));
Q_FDP4EP \internal_state_key_REG[216] ( .CK(clk), .CE(n757), .R(n1161), .D(n714), .Q(internal_state_key[216]));
Q_FDP4EP \internal_state_key_REG[217] ( .CK(clk), .CE(n757), .R(n1161), .D(n715), .Q(internal_state_key[217]));
Q_FDP4EP \internal_state_key_REG[218] ( .CK(clk), .CE(n757), .R(n1161), .D(n716), .Q(internal_state_key[218]));
Q_FDP4EP \internal_state_key_REG[219] ( .CK(clk), .CE(n757), .R(n1161), .D(n717), .Q(internal_state_key[219]));
Q_FDP4EP \internal_state_key_REG[220] ( .CK(clk), .CE(n757), .R(n1161), .D(n718), .Q(internal_state_key[220]));
Q_FDP4EP \internal_state_key_REG[221] ( .CK(clk), .CE(n757), .R(n1161), .D(n719), .Q(internal_state_key[221]));
Q_FDP4EP \internal_state_key_REG[222] ( .CK(clk), .CE(n757), .R(n1161), .D(n720), .Q(internal_state_key[222]));
Q_FDP4EP \internal_state_key_REG[223] ( .CK(clk), .CE(n757), .R(n1161), .D(n721), .Q(internal_state_key[223]));
Q_FDP4EP \internal_state_key_REG[224] ( .CK(clk), .CE(n757), .R(n1161), .D(n722), .Q(internal_state_key[224]));
Q_FDP4EP \internal_state_key_REG[225] ( .CK(clk), .CE(n757), .R(n1161), .D(n723), .Q(internal_state_key[225]));
Q_FDP4EP \internal_state_key_REG[226] ( .CK(clk), .CE(n757), .R(n1161), .D(n724), .Q(internal_state_key[226]));
Q_FDP4EP \internal_state_key_REG[227] ( .CK(clk), .CE(n757), .R(n1161), .D(n725), .Q(internal_state_key[227]));
Q_FDP4EP \internal_state_key_REG[228] ( .CK(clk), .CE(n757), .R(n1161), .D(n726), .Q(internal_state_key[228]));
Q_FDP4EP \internal_state_key_REG[229] ( .CK(clk), .CE(n757), .R(n1161), .D(n727), .Q(internal_state_key[229]));
Q_FDP4EP \internal_state_key_REG[230] ( .CK(clk), .CE(n757), .R(n1161), .D(n728), .Q(internal_state_key[230]));
Q_FDP4EP \internal_state_key_REG[231] ( .CK(clk), .CE(n757), .R(n1161), .D(n729), .Q(internal_state_key[231]));
Q_FDP4EP \internal_state_key_REG[232] ( .CK(clk), .CE(n757), .R(n1161), .D(n730), .Q(internal_state_key[232]));
Q_FDP4EP \internal_state_key_REG[233] ( .CK(clk), .CE(n757), .R(n1161), .D(n731), .Q(internal_state_key[233]));
Q_FDP4EP \internal_state_key_REG[234] ( .CK(clk), .CE(n757), .R(n1161), .D(n732), .Q(internal_state_key[234]));
Q_FDP4EP \internal_state_key_REG[235] ( .CK(clk), .CE(n757), .R(n1161), .D(n733), .Q(internal_state_key[235]));
Q_FDP4EP \internal_state_key_REG[236] ( .CK(clk), .CE(n757), .R(n1161), .D(n734), .Q(internal_state_key[236]));
Q_FDP4EP \internal_state_key_REG[237] ( .CK(clk), .CE(n757), .R(n1161), .D(n735), .Q(internal_state_key[237]));
Q_FDP4EP \internal_state_key_REG[238] ( .CK(clk), .CE(n757), .R(n1161), .D(n736), .Q(internal_state_key[238]));
Q_FDP4EP \internal_state_key_REG[239] ( .CK(clk), .CE(n757), .R(n1161), .D(n737), .Q(internal_state_key[239]));
Q_FDP4EP \internal_state_key_REG[240] ( .CK(clk), .CE(n757), .R(n1161), .D(n738), .Q(internal_state_key[240]));
Q_FDP4EP \internal_state_key_REG[241] ( .CK(clk), .CE(n757), .R(n1161), .D(n739), .Q(internal_state_key[241]));
Q_FDP4EP \internal_state_key_REG[242] ( .CK(clk), .CE(n757), .R(n1161), .D(n740), .Q(internal_state_key[242]));
Q_FDP4EP \internal_state_key_REG[243] ( .CK(clk), .CE(n757), .R(n1161), .D(n741), .Q(internal_state_key[243]));
Q_FDP4EP \internal_state_key_REG[244] ( .CK(clk), .CE(n757), .R(n1161), .D(n742), .Q(internal_state_key[244]));
Q_FDP4EP \internal_state_key_REG[245] ( .CK(clk), .CE(n757), .R(n1161), .D(n743), .Q(internal_state_key[245]));
Q_FDP4EP \internal_state_key_REG[246] ( .CK(clk), .CE(n757), .R(n1161), .D(n744), .Q(internal_state_key[246]));
Q_FDP4EP \internal_state_key_REG[247] ( .CK(clk), .CE(n757), .R(n1161), .D(n745), .Q(internal_state_key[247]));
Q_FDP4EP \internal_state_key_REG[248] ( .CK(clk), .CE(n757), .R(n1161), .D(n746), .Q(internal_state_key[248]));
Q_FDP4EP \internal_state_key_REG[249] ( .CK(clk), .CE(n757), .R(n1161), .D(n747), .Q(internal_state_key[249]));
Q_FDP4EP \internal_state_key_REG[250] ( .CK(clk), .CE(n757), .R(n1161), .D(n748), .Q(internal_state_key[250]));
Q_FDP4EP \internal_state_key_REG[251] ( .CK(clk), .CE(n757), .R(n1161), .D(n749), .Q(internal_state_key[251]));
Q_FDP4EP \internal_state_key_REG[252] ( .CK(clk), .CE(n757), .R(n1161), .D(n750), .Q(internal_state_key[252]));
Q_FDP4EP \internal_state_key_REG[253] ( .CK(clk), .CE(n757), .R(n1161), .D(n751), .Q(internal_state_key[253]));
Q_FDP4EP \internal_state_key_REG[254] ( .CK(clk), .CE(n757), .R(n1161), .D(n752), .Q(internal_state_key[254]));
Q_FDP4EP \internal_state_key_REG[255] ( .CK(clk), .CE(n757), .R(n1161), .D(n753), .Q(internal_state_key[255]));
Q_FDP4EP \reseed_counter_REG[0] ( .CK(clk), .CE(n495), .R(n1161), .D(n447), .Q(reseed_counter[0]));
Q_FDP4EP \reseed_counter_REG[1] ( .CK(clk), .CE(n495), .R(n1161), .D(n448), .Q(reseed_counter[1]));
Q_FDP4EP \reseed_counter_REG[2] ( .CK(clk), .CE(n495), .R(n1161), .D(n449), .Q(reseed_counter[2]));
Q_FDP4EP \reseed_counter_REG[3] ( .CK(clk), .CE(n495), .R(n1161), .D(n450), .Q(reseed_counter[3]));
Q_FDP4EP \reseed_counter_REG[4] ( .CK(clk), .CE(n495), .R(n1161), .D(n451), .Q(reseed_counter[4]));
Q_FDP4EP \reseed_counter_REG[5] ( .CK(clk), .CE(n495), .R(n1161), .D(n452), .Q(reseed_counter[5]));
Q_FDP4EP \reseed_counter_REG[6] ( .CK(clk), .CE(n495), .R(n1161), .D(n453), .Q(reseed_counter[6]));
Q_FDP4EP \reseed_counter_REG[7] ( .CK(clk), .CE(n495), .R(n1161), .D(n454), .Q(reseed_counter[7]));
Q_FDP4EP \reseed_counter_REG[8] ( .CK(clk), .CE(n495), .R(n1161), .D(n455), .Q(reseed_counter[8]));
Q_FDP4EP \reseed_counter_REG[9] ( .CK(clk), .CE(n495), .R(n1161), .D(n456), .Q(reseed_counter[9]));
Q_FDP4EP \reseed_counter_REG[10] ( .CK(clk), .CE(n495), .R(n1161), .D(n457), .Q(reseed_counter[10]));
Q_FDP4EP \reseed_counter_REG[11] ( .CK(clk), .CE(n495), .R(n1161), .D(n458), .Q(reseed_counter[11]));
Q_FDP4EP \reseed_counter_REG[12] ( .CK(clk), .CE(n495), .R(n1161), .D(n459), .Q(reseed_counter[12]));
Q_FDP4EP \reseed_counter_REG[13] ( .CK(clk), .CE(n495), .R(n1161), .D(n460), .Q(reseed_counter[13]));
Q_FDP4EP \reseed_counter_REG[14] ( .CK(clk), .CE(n495), .R(n1161), .D(n461), .Q(reseed_counter[14]));
Q_FDP4EP \reseed_counter_REG[15] ( .CK(clk), .CE(n495), .R(n1161), .D(n462), .Q(reseed_counter[15]));
Q_FDP4EP \reseed_counter_REG[16] ( .CK(clk), .CE(n495), .R(n1161), .D(n463), .Q(reseed_counter[16]));
Q_FDP4EP \reseed_counter_REG[17] ( .CK(clk), .CE(n495), .R(n1161), .D(n464), .Q(reseed_counter[17]));
Q_FDP4EP \reseed_counter_REG[18] ( .CK(clk), .CE(n495), .R(n1161), .D(n465), .Q(reseed_counter[18]));
Q_FDP4EP \reseed_counter_REG[19] ( .CK(clk), .CE(n495), .R(n1161), .D(n466), .Q(reseed_counter[19]));
Q_FDP4EP \reseed_counter_REG[20] ( .CK(clk), .CE(n495), .R(n1161), .D(n467), .Q(reseed_counter[20]));
Q_FDP4EP \reseed_counter_REG[21] ( .CK(clk), .CE(n495), .R(n1161), .D(n468), .Q(reseed_counter[21]));
Q_FDP4EP \reseed_counter_REG[22] ( .CK(clk), .CE(n495), .R(n1161), .D(n469), .Q(reseed_counter[22]));
Q_FDP4EP \reseed_counter_REG[23] ( .CK(clk), .CE(n495), .R(n1161), .D(n470), .Q(reseed_counter[23]));
Q_FDP4EP \reseed_counter_REG[24] ( .CK(clk), .CE(n495), .R(n1161), .D(n471), .Q(reseed_counter[24]));
Q_FDP4EP \reseed_counter_REG[25] ( .CK(clk), .CE(n495), .R(n1161), .D(n472), .Q(reseed_counter[25]));
Q_FDP4EP \reseed_counter_REG[26] ( .CK(clk), .CE(n495), .R(n1161), .D(n473), .Q(reseed_counter[26]));
Q_FDP4EP \reseed_counter_REG[27] ( .CK(clk), .CE(n495), .R(n1161), .D(n474), .Q(reseed_counter[27]));
Q_FDP4EP \reseed_counter_REG[28] ( .CK(clk), .CE(n495), .R(n1161), .D(n475), .Q(reseed_counter[28]));
Q_FDP4EP \reseed_counter_REG[29] ( .CK(clk), .CE(n495), .R(n1161), .D(n476), .Q(reseed_counter[29]));
Q_FDP4EP \reseed_counter_REG[30] ( .CK(clk), .CE(n495), .R(n1161), .D(n477), .Q(reseed_counter[30]));
Q_FDP4EP \reseed_counter_REG[31] ( .CK(clk), .CE(n495), .R(n1161), .D(n478), .Q(reseed_counter[31]));
Q_FDP4EP \reseed_counter_REG[32] ( .CK(clk), .CE(n495), .R(n1161), .D(n479), .Q(reseed_counter[32]));
Q_FDP4EP \reseed_counter_REG[33] ( .CK(clk), .CE(n495), .R(n1161), .D(n480), .Q(reseed_counter[33]));
Q_FDP4EP \reseed_counter_REG[34] ( .CK(clk), .CE(n495), .R(n1161), .D(n481), .Q(reseed_counter[34]));
Q_FDP4EP \reseed_counter_REG[35] ( .CK(clk), .CE(n495), .R(n1161), .D(n482), .Q(reseed_counter[35]));
Q_FDP4EP \reseed_counter_REG[36] ( .CK(clk), .CE(n495), .R(n1161), .D(n483), .Q(reseed_counter[36]));
Q_FDP4EP \reseed_counter_REG[37] ( .CK(clk), .CE(n495), .R(n1161), .D(n484), .Q(reseed_counter[37]));
Q_FDP4EP \reseed_counter_REG[38] ( .CK(clk), .CE(n495), .R(n1161), .D(n485), .Q(reseed_counter[38]));
Q_FDP4EP \reseed_counter_REG[39] ( .CK(clk), .CE(n495), .R(n1161), .D(n486), .Q(reseed_counter[39]));
Q_FDP4EP \reseed_counter_REG[40] ( .CK(clk), .CE(n495), .R(n1161), .D(n487), .Q(reseed_counter[40]));
Q_FDP4EP \reseed_counter_REG[41] ( .CK(clk), .CE(n495), .R(n1161), .D(n488), .Q(reseed_counter[41]));
Q_FDP4EP \reseed_counter_REG[42] ( .CK(clk), .CE(n495), .R(n1161), .D(n489), .Q(reseed_counter[42]));
Q_FDP4EP \reseed_counter_REG[43] ( .CK(clk), .CE(n495), .R(n1161), .D(n490), .Q(reseed_counter[43]));
Q_FDP4EP \reseed_counter_REG[44] ( .CK(clk), .CE(n495), .R(n1161), .D(n491), .Q(reseed_counter[44]));
Q_FDP4EP \reseed_counter_REG[45] ( .CK(clk), .CE(n495), .R(n1161), .D(n492), .Q(reseed_counter[45]));
Q_FDP4EP \reseed_counter_REG[46] ( .CK(clk), .CE(n495), .R(n1161), .D(n493), .Q(reseed_counter[46]));
Q_FDP4EP \reseed_counter_REG[47] ( .CK(clk), .CE(n495), .R(n1161), .D(n494), .Q(reseed_counter[47]));
Q_FDP4EP \reseed_counter_limit_REG[0] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[0]), .Q(reseed_counter_limit[0]));
Q_FDP4EP \reseed_counter_limit_REG[1] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[1]), .Q(reseed_counter_limit[1]));
Q_FDP4EP \reseed_counter_limit_REG[2] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[2]), .Q(reseed_counter_limit[2]));
Q_FDP4EP \reseed_counter_limit_REG[3] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[3]), .Q(reseed_counter_limit[3]));
Q_FDP4EP \reseed_counter_limit_REG[4] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[4]), .Q(reseed_counter_limit[4]));
Q_FDP4EP \reseed_counter_limit_REG[5] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[5]), .Q(reseed_counter_limit[5]));
Q_FDP4EP \reseed_counter_limit_REG[6] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[6]), .Q(reseed_counter_limit[6]));
Q_FDP4EP \reseed_counter_limit_REG[7] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[7]), .Q(reseed_counter_limit[7]));
Q_FDP4EP \reseed_counter_limit_REG[8] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[8]), .Q(reseed_counter_limit[8]));
Q_FDP4EP \reseed_counter_limit_REG[9] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[9]), .Q(reseed_counter_limit[9]));
Q_FDP4EP \reseed_counter_limit_REG[10] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[10]), .Q(reseed_counter_limit[10]));
Q_FDP4EP \reseed_counter_limit_REG[11] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[11]), .Q(reseed_counter_limit[11]));
Q_FDP4EP \reseed_counter_limit_REG[12] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[12]), .Q(reseed_counter_limit[12]));
Q_FDP4EP \reseed_counter_limit_REG[13] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[13]), .Q(reseed_counter_limit[13]));
Q_FDP4EP \reseed_counter_limit_REG[14] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[14]), .Q(reseed_counter_limit[14]));
Q_FDP4EP \reseed_counter_limit_REG[15] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[15]), .Q(reseed_counter_limit[15]));
Q_FDP4EP \reseed_counter_limit_REG[16] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[16]), .Q(reseed_counter_limit[16]));
Q_FDP4EP \reseed_counter_limit_REG[17] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[17]), .Q(reseed_counter_limit[17]));
Q_FDP4EP \reseed_counter_limit_REG[18] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[18]), .Q(reseed_counter_limit[18]));
Q_FDP4EP \reseed_counter_limit_REG[19] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[19]), .Q(reseed_counter_limit[19]));
Q_FDP4EP \reseed_counter_limit_REG[20] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[20]), .Q(reseed_counter_limit[20]));
Q_FDP4EP \reseed_counter_limit_REG[21] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[21]), .Q(reseed_counter_limit[21]));
Q_FDP4EP \reseed_counter_limit_REG[22] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[22]), .Q(reseed_counter_limit[22]));
Q_FDP4EP \reseed_counter_limit_REG[23] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[23]), .Q(reseed_counter_limit[23]));
Q_FDP4EP \reseed_counter_limit_REG[24] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[24]), .Q(reseed_counter_limit[24]));
Q_FDP4EP \reseed_counter_limit_REG[25] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[25]), .Q(reseed_counter_limit[25]));
Q_FDP4EP \reseed_counter_limit_REG[26] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[26]), .Q(reseed_counter_limit[26]));
Q_FDP4EP \reseed_counter_limit_REG[27] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[27]), .Q(reseed_counter_limit[27]));
Q_FDP4EP \reseed_counter_limit_REG[28] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[28]), .Q(reseed_counter_limit[28]));
Q_FDP4EP \reseed_counter_limit_REG[29] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[29]), .Q(reseed_counter_limit[29]));
Q_FDP4EP \reseed_counter_limit_REG[30] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[30]), .Q(reseed_counter_limit[30]));
Q_FDP4EP \reseed_counter_limit_REG[31] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[31]), .Q(reseed_counter_limit[31]));
Q_FDP4EP \reseed_counter_limit_REG[32] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[32]), .Q(reseed_counter_limit[32]));
Q_FDP4EP \reseed_counter_limit_REG[33] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[33]), .Q(reseed_counter_limit[33]));
Q_FDP4EP \reseed_counter_limit_REG[34] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[34]), .Q(reseed_counter_limit[34]));
Q_FDP4EP \reseed_counter_limit_REG[35] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[35]), .Q(reseed_counter_limit[35]));
Q_FDP4EP \reseed_counter_limit_REG[36] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[36]), .Q(reseed_counter_limit[36]));
Q_FDP4EP \reseed_counter_limit_REG[37] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[37]), .Q(reseed_counter_limit[37]));
Q_FDP4EP \reseed_counter_limit_REG[38] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[38]), .Q(reseed_counter_limit[38]));
Q_FDP4EP \reseed_counter_limit_REG[39] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[39]), .Q(reseed_counter_limit[39]));
Q_FDP4EP \reseed_counter_limit_REG[40] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[40]), .Q(reseed_counter_limit[40]));
Q_FDP4EP \reseed_counter_limit_REG[41] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[41]), .Q(reseed_counter_limit[41]));
Q_FDP4EP \reseed_counter_limit_REG[42] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[42]), .Q(reseed_counter_limit[42]));
Q_FDP4EP \reseed_counter_limit_REG[43] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[43]), .Q(reseed_counter_limit[43]));
Q_FDP4EP \reseed_counter_limit_REG[44] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[44]), .Q(reseed_counter_limit[44]));
Q_FDP4EP \reseed_counter_limit_REG[45] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[45]), .Q(reseed_counter_limit[45]));
Q_FDP4EP \reseed_counter_limit_REG[46] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[46]), .Q(reseed_counter_limit[46]));
Q_FDP4EP \reseed_counter_limit_REG[47] ( .CK(clk), .CE(n497), .R(n1161), .D(seed_life[47]), .Q(reseed_counter_limit[47]));
endmodule
