
module ASSERTION ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire FAILURE;
Q_OR02 U0 ( .A0(xc_top.stop2), .A1(_ixc_isc.assertUCF), .Z(FAILURE));
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
endmodule
