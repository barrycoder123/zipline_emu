architecture module of axis_busreg is
  -- quickturn CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
  component Q_BRP
    port(Z : out std_logic) ;
  end component ;

begin
  _UnNamed_Inst_29 : Q_BRP port map (z) ;
end module;
