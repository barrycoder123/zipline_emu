
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
`_2_ (* upf_always_on = 1 *) 
module xc_top_1 ;
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
wire fclk;
wire uClk;
wire _ET3_COMPILER_RESERVED_NAME_DUTPI_APPLY_;
wire _ET3_COMPILER_RESERVED_NAME_LBRKER_ON_;
wire [63:0] _ET3_COMPILER_RESERVED_NAME_QT_CURR_EMUL_CYCLE_;
wire xc1xEcm;
wire callEmuPI;
wire [63:0] evalStepPI;
wire ckgHoldPI;
wire tbcHoldPI;
wire noOutputPI;
wire stopEmuPI;
wire oneStepPI;
wire stop1;
wire stop2;
wire stop4;
wire GFbusy;
wire svGFbusy;
wire otbGFbusy;
wire asyncCall;
wire svAsyncCall;
wire otbAsyncCall;
wire isfWait;
wire osfWait;
wire gfifoWait;
wire ecmHoldBusy;
wire sdlStop;
wire cpfStop;
wire eClk;
wire clockMCInit;
wire hasSFIFO;
wire hasGFIFO1;
wire hasGFIFO2;
wire hasPTX;
wire bpWait;
wire bWait;
wire xpHold;
wire mpEnable;
wire ixcHoldClk;
wire cakeCcEnable;
wire ptxBusy;
wire holdEcm;
wire bpHalt;
wire acHalt;
wire lockTrace;
wire [63:0] mioPOW_0;
wire [63:0] mioPOW_2;
wire mioPICnt;
wire [63:0] evalStepPIi;
wire callEmuPIi;
wire ckgHoldPIi;
wire stopEmuPIi;
wire oneStepPIi;
wire callEmuEv;
wire eventOn;
wire APPLY_PI;
wire APPLY_DUTPI;
wire lbrOnAll;
wire anyStop;
wire GFLBfull;
wire GFGBfull;
wire GFBw;
wire GFAck;
wire stopCond;
wire [12:0] GF2LevelMask;
wire bClk;
wire sampleXpChg;
wire bClkRH;
wire bClkHold;
wire it_endBuf;
wire it_newBuf;
wire _zz_xmr0;
wire dummyW;
wire syncEn;
wire ecmOn;
wire ecmSync;
wire ecmNotSync;
wire holdEcmTb;
wire ptxHoldEcm;
wire [31:0] mcDelta;
wire mcp;
`_2_ wire _ET3_COMPILER_RESERVED_NAME_ORION_INTERRUPT_;
`_2_ wire _ET3_COMPILER_RESERVED_NAME_DBI_APPLY_;
`_2_ wire _ET3_COMPILER_RESERVED_NAME_DBO_SAMPLE_;
`_2_ wire hotSwapOnPI;
`_2_ wire hssReset;
`_2_ wire sendPO;
`_2_ wire tbcPO;
`_2_ wire tbcPOd;
`_2_ wire stop1PO;
`_2_ wire stop1POd;
`_2_ wire stop2PO;
`_2_ wire stop2POd;
`_2_ wire stop4PO;
`_2_ wire stop4POd;
`_2_ wire stop3PO;
`_2_ wire stop3POd;
`_2_ wire it_newBufPO;
`_2_ wire stopSDLPO;
`_2_ wire stopEmuPO;
`_2_ wire stopCPFPO;
`_2_ wire [63:0] remStepPO;
`_2_ wire GFReset;
`_2_ wire stop3;
`_2_ wire stop1R;
`_2_ wire stop2R;
`_2_ wire stop4R;
`_2_ wire stopSDL;
`_2_ wire sdlStopRply;
`_2_ wire sdlStopRplyD;
`_2_ wire sdlEnable;
`_2_ wire sdlHaltHwClk;
`_2_ wire GFbusyW;
`_2_ wire FTcallW;
`_2_ wire FvSimple2;
`_2_ wire [7:0] DccFrameCycle;
`_2_ wire [7:0] DccFrameMark;
`_2_ wire [7:0] dccFrameFill;
`_2_ wire noHoldOn;
`_2_ wire tbcEnable;
`_2_ wire hwClkEnable;
`_2_ wire hwClkDbgEn;
`_2_ wire hwClkDbg;
`_2_ wire hwClkDbgOn;
`_2_ wire hwClkDbgTime;
`_2_ wire [63:0] hwSimTime;
`_2_ wire [63:0] ixcSimTime;
`_2_ wire [31:0] hwClkDelay;
`_2_ wire bpOn;
`_2_ wire bpOnD;
`_2_ wire mpOn;
`_2_ wire ecmOne;
`_2_ wire [7:0] fclkPerEval;
`_2_ wire tbcHold;
`_2_ wire stopT;
`_2_ wire stopTL;
`_2_ wire stopTLd;
`_2_ wire clockMC;
`_2_ wire eClkR;
`_2_ wire evalOn;
`_2_ wire evalOnOrig;
`_2_ wire sfifoSyncMode;
`_2_ wire syncOtbChannels;
`_2_ wire [7:0] gfPushDly;
`_2_ wire [3:0] gfPushFill;
`_2_ wire bWaitExtend;
`_2_ wire lastDelta;
`_2_ wire callEmu;
`_2_ wire callEmuPre;
`_2_ wire callEmuR;
`_2_ wire evalOnC;
`_2_ wire evalOnD;
`_2_ wire [2:0] fcnt;
`_2_ wire [7:0] evalOnDExt;
`_2_ wire [7:0] evalOnDCtl;
`_2_ wire simTimeOn;
`_2_ wire nextTime;
`_2_ wire [63:0] eCount;
`_2_ wire [63:0] evfCount;
`_2_ wire [63:0] bCount;
`_2_ wire [63:0] bpCount;
`_2_ wire [63:0] nbaCount;
`_2_ wire [31:0] aCount;
`_2_ wire [63:0] ixcHoldClkCnt;
`_2_ wire [63:0] ixcHoldSyncCnt;
`_2_ wire [63:0] ixcHoldEcmCnt;
`_2_ wire [63:0] fvSCount;
`_2_ wire [63:0] simTime;
`_2_ wire simTimeEnable;
`_2_ wire cakeUcEnable;
`_2_ wire initClock;
`_2_ wire holdEcmC;
`_2_ wire holdEcmD;
`_2_ wire xcReplayOn;
`_2_ wire xcRecordOn;
`_2_ wire evalOnSync;
`_2_ wire evalOnInt;
`_2_ wire [2:0] evalOnIntR;
`_2_ wire evalOnIntD;
`_2_ wire forceAbort;
`_2_ wire [15:0] bHaltCnt;
`_2_ wire [15:0] maxBpCycle;
`_2_ wire [15:0] aHaltCnt;
`_2_ wire [15:0] maxAcCycle;
`_2_ wire [3:0] lockTraceC;
`_2_ wire lockTraceOn;
`_2_ wire [63:0] lockTraceTime;
`_2_ wire xc_mioOn;
`_2_ wire xc_mioOnS;
`_2_ wire mioPOCnt;
`_2_ wire tbcPOmio;
`_2_ wire [63:0] mioPIW_0;
`_2_ wire [63:0] mioPIW_1;
`_2_ wire mioPICntd;
`_2_ wire [63:0] evalStepPImio;
`_2_ wire callEmuPImio;
`_2_ wire ckgHoldPImio;
`_2_ wire oneStepPImio;
`_2_ wire [63:0] nextDutTimeS;
`_2_ wire callEmuWaitC;
`_2_ wire callEmuWait;
`_2_ wire callEmuWaitN;
`_2_ wire callEmuPreD;
`_2_ wire applyPiR;
`_2_ wire dbiEvent;
`_2_ wire dbiEventD;
`_2_ wire FvUseOnly;
`_2_ wire FvUseOnlyR;
`_2_ wire eventOnR;
`_2_ wire eventOnRI;
`_2_ wire mpSampleOv;
`_2_ wire lbrOn;
`_2_ wire gfifoOff;
`_2_ wire gfifoAsyncOff;
`_2_ wire GFLock1;
`_2_ wire GFLock2;
`_2_ wire GFGBfullBw;
`_2_ wire GFGBfullBwD;
`_2_ wire GFLBfullD;
`_2_ wire tbcPOReg;
`_2_ wire xcReplayOnReg;
`_2_ wire GFLock2R;
`_2_ wire SFIFOLock;
`_2_ wire [7:0] gfifoAckWait;
`_2_ wire [2:0] mpSt;
`_2_ wire active;
`_2_ wire asyncBusy;
`_2_ wire GFbusyD;
`_2_ wire GFbusyD2;
`_2_ wire [12:0] tbcPODly;
`_2_ wire tbcPORdy;
`_2_ wire [1:0] tbcPOState;
`_2_ wire [1:0] tbcPOStateN;
`_2_ wire SFIFOLock2;
`_2_ wire bClkR;
`_2_ wire sampleXpV;
`_2_ wire [1:0] bpSt;
`_2_ wire bClkHoldD;
`_2_ wire ixcHoldClkR;
`_2_ wire intr;
`_2_ wire it_capture;
`_2_ wire it_replay;
`_2_ wire dummyR;
`_2_ wire hwClkHalt;
`_2_ wire sdlHaltHwClkR;
`_2_ wire [63:0] gfifoGBfullCnt;
`_2_ wire [63:0] gfifoLBfullCnt;
`_2_ wire [63:0] gfifoTBsyncCnt;
`_2_ wire [15:0] maxFck2Sync;
`_2_ wire [15:0] maxGfifo2Sync;
`_2_ wire [15:0] Fck2Sync;
`_2_ wire [15:0] Gfifo2Sync;
`_2_ wire ptxStop;
`_2_ wire ecmOnD;
`_2_ wire ecmNotSyncD;
`_2_ wire holdEcmPtxOn;
`_2_ wire holdEcmSync;
`_2_ wire dccState;
`_2_ wire [63:0] nextDutTimeP;
`_2_ wire [63:0] fclkCntr;
`_2_ wire [63:0] uClkCntr;
`_2_ wire [63:0] uClkErrTime;
supply1 n2504;
supply0 n3717;
supply1 n3718;
supply0 n3719;
supply1 n3720;
Q_BUF U0 ( .A(n2504), .Z(xc1xEcm));
Q_BUF U1 ( .A(n3717), .Z(mioPOW_2[63]));
Q_BUF U2 ( .A(n3717), .Z(mioPOW_2[62]));
Q_BUF U3 ( .A(n3717), .Z(mioPOW_2[61]));
Q_BUF U4 ( .A(n3717), .Z(mioPOW_2[60]));
Q_BUF U5 ( .A(n3717), .Z(mioPOW_2[59]));
Q_BUF U6 ( .A(n3717), .Z(mioPOW_2[58]));
Q_BUF U7 ( .A(n3717), .Z(mioPOW_2[57]));
Q_BUF U8 ( .A(n3717), .Z(mioPOW_2[56]));
Q_BUF U9 ( .A(n3717), .Z(mioPOW_2[55]));
Q_BUF U10 ( .A(n3717), .Z(mioPOW_2[54]));
Q_BUF U11 ( .A(n3717), .Z(mioPOW_2[53]));
Q_BUF U12 ( .A(n3717), .Z(mioPOW_2[52]));
Q_BUF U13 ( .A(n3717), .Z(mioPOW_2[51]));
Q_BUF U14 ( .A(n3717), .Z(mioPOW_2[50]));
Q_BUF U15 ( .A(n3717), .Z(mioPOW_2[49]));
Q_BUF U16 ( .A(n3717), .Z(mioPOW_2[48]));
Q_BUF U17 ( .A(n3717), .Z(mioPOW_2[47]));
Q_BUF U18 ( .A(n3717), .Z(mioPOW_2[46]));
Q_BUF U19 ( .A(n3717), .Z(mioPOW_2[45]));
Q_BUF U20 ( .A(n3717), .Z(mioPOW_2[44]));
Q_BUF U21 ( .A(n3717), .Z(mioPOW_2[43]));
Q_BUF U22 ( .A(n3717), .Z(mioPOW_2[42]));
Q_BUF U23 ( .A(n3717), .Z(mioPOW_2[41]));
Q_BUF U24 ( .A(n3717), .Z(mioPOW_2[40]));
Q_BUF U25 ( .A(n3717), .Z(mioPOW_2[39]));
Q_BUF U26 ( .A(n3717), .Z(mioPOW_2[38]));
Q_BUF U27 ( .A(n3717), .Z(mioPOW_2[37]));
Q_BUF U28 ( .A(n3717), .Z(mioPOW_2[36]));
Q_BUF U29 ( .A(n3717), .Z(mioPOW_2[35]));
Q_BUF U30 ( .A(n3717), .Z(mioPOW_2[34]));
Q_BUF U31 ( .A(n3717), .Z(mioPOW_2[33]));
Q_BUF U32 ( .A(n3717), .Z(mioPOW_2[32]));
Q_BUF U33 ( .A(n3717), .Z(mioPOW_2[31]));
Q_BUF U34 ( .A(n3717), .Z(mioPOW_2[30]));
Q_BUF U35 ( .A(n3717), .Z(mioPOW_2[29]));
Q_BUF U36 ( .A(n3717), .Z(mioPOW_2[28]));
Q_BUF U37 ( .A(n3717), .Z(mioPOW_2[27]));
Q_BUF U38 ( .A(n3717), .Z(mioPOW_2[26]));
Q_BUF U39 ( .A(n3717), .Z(mioPOW_2[25]));
Q_BUF U40 ( .A(n3717), .Z(mioPOW_2[24]));
Q_BUF U41 ( .A(n3717), .Z(mioPOW_2[23]));
Q_BUF U42 ( .A(n3717), .Z(mioPOW_2[22]));
Q_BUF U43 ( .A(n3717), .Z(mioPOW_2[21]));
Q_BUF U44 ( .A(n3717), .Z(mioPOW_2[20]));
Q_BUF U45 ( .A(n3717), .Z(mioPOW_2[19]));
Q_BUF U46 ( .A(n3717), .Z(mioPOW_2[18]));
Q_BUF U47 ( .A(n3717), .Z(mioPOW_2[17]));
Q_BUF U48 ( .A(n3717), .Z(mioPOW_2[16]));
Q_BUF U49 ( .A(n3717), .Z(mioPOW_2[15]));
Q_BUF U50 ( .A(n3717), .Z(mioPOW_2[14]));
Q_BUF U51 ( .A(n3717), .Z(mioPOW_2[13]));
Q_BUF U52 ( .A(n3717), .Z(mioPOW_2[12]));
Q_BUF U53 ( .A(n3717), .Z(mioPOW_2[11]));
Q_BUF U54 ( .A(n3717), .Z(mioPOW_2[10]));
Q_BUF U55 ( .A(n3717), .Z(mioPOW_2[9]));
Q_BUF U56 ( .A(lockTraceC[3]), .Z(lockTrace));
Q_BUF U57 ( .A(mioPOCnt), .Z(mioPOW_0[63]));
Q_BUF U58 ( .A(evalStepPIi[63]), .Z(ixc_time.nextTbTime[63]));
Q_BUF U59 ( .A(evalStepPIi[62]), .Z(ixc_time.nextTbTime[62]));
Q_BUF U60 ( .A(evalStepPIi[61]), .Z(ixc_time.nextTbTime[61]));
Q_BUF U61 ( .A(evalStepPIi[60]), .Z(ixc_time.nextTbTime[60]));
Q_BUF U62 ( .A(evalStepPIi[59]), .Z(ixc_time.nextTbTime[59]));
Q_BUF U63 ( .A(evalStepPIi[58]), .Z(ixc_time.nextTbTime[58]));
Q_BUF U64 ( .A(evalStepPIi[57]), .Z(ixc_time.nextTbTime[57]));
Q_BUF U65 ( .A(evalStepPIi[56]), .Z(ixc_time.nextTbTime[56]));
Q_BUF U66 ( .A(evalStepPIi[55]), .Z(ixc_time.nextTbTime[55]));
Q_BUF U67 ( .A(evalStepPIi[54]), .Z(ixc_time.nextTbTime[54]));
Q_BUF U68 ( .A(evalStepPIi[53]), .Z(ixc_time.nextTbTime[53]));
Q_BUF U69 ( .A(evalStepPIi[52]), .Z(ixc_time.nextTbTime[52]));
Q_BUF U70 ( .A(evalStepPIi[51]), .Z(ixc_time.nextTbTime[51]));
Q_BUF U71 ( .A(evalStepPIi[50]), .Z(ixc_time.nextTbTime[50]));
Q_BUF U72 ( .A(evalStepPIi[49]), .Z(ixc_time.nextTbTime[49]));
Q_BUF U73 ( .A(evalStepPIi[48]), .Z(ixc_time.nextTbTime[48]));
Q_BUF U74 ( .A(evalStepPIi[47]), .Z(ixc_time.nextTbTime[47]));
Q_BUF U75 ( .A(evalStepPIi[46]), .Z(ixc_time.nextTbTime[46]));
Q_BUF U76 ( .A(evalStepPIi[45]), .Z(ixc_time.nextTbTime[45]));
Q_BUF U77 ( .A(evalStepPIi[44]), .Z(ixc_time.nextTbTime[44]));
Q_BUF U78 ( .A(evalStepPIi[43]), .Z(ixc_time.nextTbTime[43]));
Q_BUF U79 ( .A(evalStepPIi[42]), .Z(ixc_time.nextTbTime[42]));
Q_BUF U80 ( .A(evalStepPIi[41]), .Z(ixc_time.nextTbTime[41]));
Q_BUF U81 ( .A(evalStepPIi[40]), .Z(ixc_time.nextTbTime[40]));
Q_BUF U82 ( .A(evalStepPIi[39]), .Z(ixc_time.nextTbTime[39]));
Q_BUF U83 ( .A(evalStepPIi[38]), .Z(ixc_time.nextTbTime[38]));
Q_BUF U84 ( .A(evalStepPIi[37]), .Z(ixc_time.nextTbTime[37]));
Q_BUF U85 ( .A(evalStepPIi[36]), .Z(ixc_time.nextTbTime[36]));
Q_BUF U86 ( .A(evalStepPIi[35]), .Z(ixc_time.nextTbTime[35]));
Q_BUF U87 ( .A(evalStepPIi[34]), .Z(ixc_time.nextTbTime[34]));
Q_BUF U88 ( .A(evalStepPIi[33]), .Z(ixc_time.nextTbTime[33]));
Q_BUF U89 ( .A(evalStepPIi[32]), .Z(ixc_time.nextTbTime[32]));
Q_BUF U90 ( .A(evalStepPIi[31]), .Z(ixc_time.nextTbTime[31]));
Q_BUF U91 ( .A(evalStepPIi[30]), .Z(ixc_time.nextTbTime[30]));
Q_BUF U92 ( .A(evalStepPIi[29]), .Z(ixc_time.nextTbTime[29]));
Q_BUF U93 ( .A(evalStepPIi[28]), .Z(ixc_time.nextTbTime[28]));
Q_BUF U94 ( .A(evalStepPIi[27]), .Z(ixc_time.nextTbTime[27]));
Q_BUF U95 ( .A(evalStepPIi[26]), .Z(ixc_time.nextTbTime[26]));
Q_BUF U96 ( .A(evalStepPIi[25]), .Z(ixc_time.nextTbTime[25]));
Q_BUF U97 ( .A(evalStepPIi[24]), .Z(ixc_time.nextTbTime[24]));
Q_BUF U98 ( .A(evalStepPIi[23]), .Z(ixc_time.nextTbTime[23]));
Q_BUF U99 ( .A(evalStepPIi[22]), .Z(ixc_time.nextTbTime[22]));
Q_BUF U100 ( .A(evalStepPIi[21]), .Z(ixc_time.nextTbTime[21]));
Q_BUF U101 ( .A(evalStepPIi[20]), .Z(ixc_time.nextTbTime[20]));
Q_BUF U102 ( .A(evalStepPIi[19]), .Z(ixc_time.nextTbTime[19]));
Q_BUF U103 ( .A(evalStepPIi[18]), .Z(ixc_time.nextTbTime[18]));
Q_BUF U104 ( .A(evalStepPIi[17]), .Z(ixc_time.nextTbTime[17]));
Q_BUF U105 ( .A(evalStepPIi[16]), .Z(ixc_time.nextTbTime[16]));
Q_BUF U106 ( .A(evalStepPIi[15]), .Z(ixc_time.nextTbTime[15]));
Q_BUF U107 ( .A(evalStepPIi[14]), .Z(ixc_time.nextTbTime[14]));
Q_BUF U108 ( .A(evalStepPIi[13]), .Z(ixc_time.nextTbTime[13]));
Q_BUF U109 ( .A(evalStepPIi[12]), .Z(ixc_time.nextTbTime[12]));
Q_BUF U110 ( .A(evalStepPIi[11]), .Z(ixc_time.nextTbTime[11]));
Q_BUF U111 ( .A(evalStepPIi[10]), .Z(ixc_time.nextTbTime[10]));
Q_BUF U112 ( .A(evalStepPIi[9]), .Z(ixc_time.nextTbTime[9]));
Q_BUF U113 ( .A(evalStepPIi[8]), .Z(ixc_time.nextTbTime[8]));
Q_BUF U114 ( .A(evalStepPIi[7]), .Z(ixc_time.nextTbTime[7]));
Q_BUF U115 ( .A(evalStepPIi[6]), .Z(ixc_time.nextTbTime[6]));
Q_BUF U116 ( .A(evalStepPIi[5]), .Z(ixc_time.nextTbTime[5]));
Q_BUF U117 ( .A(evalStepPIi[4]), .Z(ixc_time.nextTbTime[4]));
Q_BUF U118 ( .A(evalStepPIi[3]), .Z(ixc_time.nextTbTime[3]));
Q_BUF U119 ( .A(evalStepPIi[2]), .Z(ixc_time.nextTbTime[2]));
Q_BUF U120 ( .A(evalStepPIi[1]), .Z(ixc_time.nextTbTime[1]));
Q_BUF U121 ( .A(evalStepPIi[0]), .Z(ixc_time.nextTbTime[0]));
Q_BUF U122 ( .A(sendPO), .Z(mioPOW_2[0]));
Q_BUF U123 ( .A(eventOnRI), .Z(eventOn));
Q_BUF U124 ( .A(stopSDLPO), .Z(mioPOW_2[7]));
Q_BUF U125 ( .A(stopCPFPO), .Z(mioPOW_2[8]));
Q_BUF U126 ( .A(stop1PO), .Z(mioPOW_2[2]));
Q_BUF U127 ( .A(stop2PO), .Z(mioPOW_2[3]));
Q_BUF U128 ( .A(stop4PO), .Z(mioPOW_2[5]));
Q_BUF U129 ( .A(stop3PO), .Z(mioPOW_2[4]));
Q_BUF U130 ( .A(stopEmuPIi), .Z(stopEmuPO));
Q_BUF U131 ( .A(remStepPO[62]), .Z(mioPOW_0[62]));
Q_BUF U132 ( .A(remStepPO[61]), .Z(mioPOW_0[61]));
Q_BUF U133 ( .A(remStepPO[60]), .Z(mioPOW_0[60]));
Q_BUF U134 ( .A(remStepPO[59]), .Z(mioPOW_0[59]));
Q_BUF U135 ( .A(remStepPO[58]), .Z(mioPOW_0[58]));
Q_BUF U136 ( .A(remStepPO[57]), .Z(mioPOW_0[57]));
Q_BUF U137 ( .A(remStepPO[56]), .Z(mioPOW_0[56]));
Q_BUF U138 ( .A(remStepPO[55]), .Z(mioPOW_0[55]));
Q_BUF U139 ( .A(remStepPO[54]), .Z(mioPOW_0[54]));
Q_BUF U140 ( .A(remStepPO[53]), .Z(mioPOW_0[53]));
Q_BUF U141 ( .A(remStepPO[52]), .Z(mioPOW_0[52]));
Q_BUF U142 ( .A(remStepPO[51]), .Z(mioPOW_0[51]));
Q_BUF U143 ( .A(remStepPO[50]), .Z(mioPOW_0[50]));
Q_BUF U144 ( .A(remStepPO[49]), .Z(mioPOW_0[49]));
Q_BUF U145 ( .A(remStepPO[48]), .Z(mioPOW_0[48]));
Q_BUF U146 ( .A(remStepPO[47]), .Z(mioPOW_0[47]));
Q_BUF U147 ( .A(remStepPO[46]), .Z(mioPOW_0[46]));
Q_BUF U148 ( .A(remStepPO[45]), .Z(mioPOW_0[45]));
Q_BUF U149 ( .A(remStepPO[44]), .Z(mioPOW_0[44]));
Q_BUF U150 ( .A(remStepPO[43]), .Z(mioPOW_0[43]));
Q_BUF U151 ( .A(remStepPO[42]), .Z(mioPOW_0[42]));
Q_BUF U152 ( .A(remStepPO[41]), .Z(mioPOW_0[41]));
Q_BUF U153 ( .A(remStepPO[40]), .Z(mioPOW_0[40]));
Q_BUF U154 ( .A(remStepPO[39]), .Z(mioPOW_0[39]));
Q_BUF U155 ( .A(remStepPO[38]), .Z(mioPOW_0[38]));
Q_BUF U156 ( .A(remStepPO[37]), .Z(mioPOW_0[37]));
Q_BUF U157 ( .A(remStepPO[36]), .Z(mioPOW_0[36]));
Q_BUF U158 ( .A(remStepPO[35]), .Z(mioPOW_0[35]));
Q_BUF U159 ( .A(remStepPO[34]), .Z(mioPOW_0[34]));
Q_BUF U160 ( .A(remStepPO[33]), .Z(mioPOW_0[33]));
Q_BUF U161 ( .A(remStepPO[32]), .Z(mioPOW_0[32]));
Q_BUF U162 ( .A(remStepPO[31]), .Z(mioPOW_0[31]));
Q_BUF U163 ( .A(remStepPO[30]), .Z(mioPOW_0[30]));
Q_BUF U164 ( .A(remStepPO[29]), .Z(mioPOW_0[29]));
Q_BUF U165 ( .A(remStepPO[28]), .Z(mioPOW_0[28]));
Q_BUF U166 ( .A(remStepPO[27]), .Z(mioPOW_0[27]));
Q_BUF U167 ( .A(remStepPO[26]), .Z(mioPOW_0[26]));
Q_BUF U168 ( .A(remStepPO[25]), .Z(mioPOW_0[25]));
Q_BUF U169 ( .A(remStepPO[24]), .Z(mioPOW_0[24]));
Q_BUF U170 ( .A(remStepPO[23]), .Z(mioPOW_0[23]));
Q_BUF U171 ( .A(remStepPO[22]), .Z(mioPOW_0[22]));
Q_BUF U172 ( .A(remStepPO[21]), .Z(mioPOW_0[21]));
Q_BUF U173 ( .A(remStepPO[20]), .Z(mioPOW_0[20]));
Q_BUF U174 ( .A(remStepPO[19]), .Z(mioPOW_0[19]));
Q_BUF U175 ( .A(remStepPO[18]), .Z(mioPOW_0[18]));
Q_BUF U176 ( .A(remStepPO[17]), .Z(mioPOW_0[17]));
Q_BUF U177 ( .A(remStepPO[16]), .Z(mioPOW_0[16]));
Q_BUF U178 ( .A(remStepPO[15]), .Z(mioPOW_0[15]));
Q_BUF U179 ( .A(remStepPO[14]), .Z(mioPOW_0[14]));
Q_BUF U180 ( .A(remStepPO[13]), .Z(mioPOW_0[13]));
Q_BUF U181 ( .A(remStepPO[12]), .Z(mioPOW_0[12]));
Q_BUF U182 ( .A(remStepPO[11]), .Z(mioPOW_0[11]));
Q_BUF U183 ( .A(remStepPO[10]), .Z(mioPOW_0[10]));
Q_BUF U184 ( .A(remStepPO[9]), .Z(mioPOW_0[9]));
Q_BUF U185 ( .A(remStepPO[8]), .Z(mioPOW_0[8]));
Q_BUF U186 ( .A(remStepPO[7]), .Z(mioPOW_0[7]));
Q_BUF U187 ( .A(remStepPO[6]), .Z(mioPOW_0[6]));
Q_BUF U188 ( .A(remStepPO[5]), .Z(mioPOW_0[5]));
Q_BUF U189 ( .A(remStepPO[4]), .Z(mioPOW_0[4]));
Q_BUF U190 ( .A(remStepPO[3]), .Z(mioPOW_0[3]));
Q_BUF U191 ( .A(remStepPO[2]), .Z(mioPOW_0[2]));
Q_BUF U192 ( .A(remStepPO[1]), .Z(mioPOW_0[1]));
Q_BUF U193 ( .A(remStepPO[0]), .Z(mioPOW_0[0]));
Q_BUF U194 ( .A(tbcPO), .Z(mioPOW_2[1]));
Q_BUF U195 ( .A(it_newBufPO), .Z(mioPOW_2[6]));
Q_ASSIGN U196 ( .B(mioPIW_1[0]), .A(mioPICnt));
Q_BUF U197 ( .A(GFBw), .Z(bClkHold));
Q_BUF U198 ( .A(n3717), .Z(n1));
Q_AN02 U199 ( .A0(n2999), .A1(n2997), .Z(n2));
Q_AN02 U200 ( .A0(n2748), .A1(n2621), .Z(n3));
Q_AN02 U201 ( .A0(n2624), .A1(evalOn), .Z(n4));
Q_AN02 U202 ( .A0(n2414), .A1(initClock), .Z(n5));
Q_AN02 U203 ( .A0(n1972), .A1(n1524), .Z(n6));
Q_AN02 U204 ( .A0(n1848), .A1(n1523), .Z(n7));
Q_AN02 U205 ( .A0(n1724), .A1(n1522), .Z(n8));
Q_AN02 U206 ( .A0(n1462), .A1(n1427), .Z(n9));
Q_AN02 U207 ( .A0(n1264), .A1(hwClkDbgOn), .Z(n10));
Q_AN02 U208 ( .A0(n664), .A1(n401), .Z(n11));
Q_AN02 U209 ( .A0(n1036), .A1(n400), .Z(n12));
Q_AN02 U210 ( .A0(n912), .A1(n399), .Z(n13));
Q_AN02 U211 ( .A0(n788), .A1(n398), .Z(n14));
Q_AN02 U212 ( .A0(n81), .A1(initClock), .Z(n15));
Q_XNR3 U213 ( .A0(n3669), .A1(ixc_time.nextDutTime[31]), .A2(nextDutTimeP[31]), .Z(mcDelta[31]));
Q_XOR2 U214 ( .A0(initClock), .A1(fclkCntr[0]), .Z(n17));
Q_FDP0UA U215 ( .D(n17), .QTFCLK( ), .Q(fclkCntr[0]));
Q_MX02 U216 ( .S(initClock), .A0(fclkCntr[1]), .A1(n204), .Z(n18));
Q_FDP0UA U217 ( .D(n18), .QTFCLK( ), .Q(fclkCntr[1]));
Q_MX02 U218 ( .S(initClock), .A0(fclkCntr[2]), .A1(n202), .Z(n19));
Q_FDP0UA U219 ( .D(n19), .QTFCLK( ), .Q(fclkCntr[2]));
Q_MX02 U220 ( .S(initClock), .A0(fclkCntr[3]), .A1(n200), .Z(n20));
Q_FDP0UA U221 ( .D(n20), .QTFCLK( ), .Q(fclkCntr[3]));
Q_MX02 U222 ( .S(initClock), .A0(fclkCntr[4]), .A1(n198), .Z(n21));
Q_FDP0UA U223 ( .D(n21), .QTFCLK( ), .Q(fclkCntr[4]));
Q_MX02 U224 ( .S(initClock), .A0(fclkCntr[5]), .A1(n196), .Z(n22));
Q_FDP0UA U225 ( .D(n22), .QTFCLK( ), .Q(fclkCntr[5]));
Q_MX02 U226 ( .S(initClock), .A0(fclkCntr[6]), .A1(n194), .Z(n23));
Q_FDP0UA U227 ( .D(n23), .QTFCLK( ), .Q(fclkCntr[6]));
Q_MX02 U228 ( .S(initClock), .A0(fclkCntr[7]), .A1(n192), .Z(n24));
Q_FDP0UA U229 ( .D(n24), .QTFCLK( ), .Q(fclkCntr[7]));
Q_MX02 U230 ( .S(initClock), .A0(fclkCntr[8]), .A1(n190), .Z(n25));
Q_FDP0UA U231 ( .D(n25), .QTFCLK( ), .Q(fclkCntr[8]));
Q_MX02 U232 ( .S(initClock), .A0(fclkCntr[9]), .A1(n188), .Z(n26));
Q_FDP0UA U233 ( .D(n26), .QTFCLK( ), .Q(fclkCntr[9]));
Q_MX02 U234 ( .S(initClock), .A0(fclkCntr[10]), .A1(n186), .Z(n27));
Q_FDP0UA U235 ( .D(n27), .QTFCLK( ), .Q(fclkCntr[10]));
Q_MX02 U236 ( .S(initClock), .A0(fclkCntr[11]), .A1(n184), .Z(n28));
Q_FDP0UA U237 ( .D(n28), .QTFCLK( ), .Q(fclkCntr[11]));
Q_MX02 U238 ( .S(initClock), .A0(fclkCntr[12]), .A1(n182), .Z(n29));
Q_FDP0UA U239 ( .D(n29), .QTFCLK( ), .Q(fclkCntr[12]));
Q_MX02 U240 ( .S(initClock), .A0(fclkCntr[13]), .A1(n180), .Z(n30));
Q_FDP0UA U241 ( .D(n30), .QTFCLK( ), .Q(fclkCntr[13]));
Q_MX02 U242 ( .S(initClock), .A0(fclkCntr[14]), .A1(n178), .Z(n31));
Q_FDP0UA U243 ( .D(n31), .QTFCLK( ), .Q(fclkCntr[14]));
Q_MX02 U244 ( .S(initClock), .A0(fclkCntr[15]), .A1(n176), .Z(n32));
Q_FDP0UA U245 ( .D(n32), .QTFCLK( ), .Q(fclkCntr[15]));
Q_MX02 U246 ( .S(initClock), .A0(fclkCntr[16]), .A1(n174), .Z(n33));
Q_FDP0UA U247 ( .D(n33), .QTFCLK( ), .Q(fclkCntr[16]));
Q_MX02 U248 ( .S(initClock), .A0(fclkCntr[17]), .A1(n172), .Z(n34));
Q_FDP0UA U249 ( .D(n34), .QTFCLK( ), .Q(fclkCntr[17]));
Q_MX02 U250 ( .S(initClock), .A0(fclkCntr[18]), .A1(n170), .Z(n35));
Q_FDP0UA U251 ( .D(n35), .QTFCLK( ), .Q(fclkCntr[18]));
Q_MX02 U252 ( .S(initClock), .A0(fclkCntr[19]), .A1(n168), .Z(n36));
Q_FDP0UA U253 ( .D(n36), .QTFCLK( ), .Q(fclkCntr[19]));
Q_MX02 U254 ( .S(initClock), .A0(fclkCntr[20]), .A1(n166), .Z(n37));
Q_FDP0UA U255 ( .D(n37), .QTFCLK( ), .Q(fclkCntr[20]));
Q_MX02 U256 ( .S(initClock), .A0(fclkCntr[21]), .A1(n164), .Z(n38));
Q_FDP0UA U257 ( .D(n38), .QTFCLK( ), .Q(fclkCntr[21]));
Q_MX02 U258 ( .S(initClock), .A0(fclkCntr[22]), .A1(n162), .Z(n39));
Q_FDP0UA U259 ( .D(n39), .QTFCLK( ), .Q(fclkCntr[22]));
Q_MX02 U260 ( .S(initClock), .A0(fclkCntr[23]), .A1(n160), .Z(n40));
Q_FDP0UA U261 ( .D(n40), .QTFCLK( ), .Q(fclkCntr[23]));
Q_MX02 U262 ( .S(initClock), .A0(fclkCntr[24]), .A1(n158), .Z(n41));
Q_FDP0UA U263 ( .D(n41), .QTFCLK( ), .Q(fclkCntr[24]));
Q_MX02 U264 ( .S(initClock), .A0(fclkCntr[25]), .A1(n156), .Z(n42));
Q_FDP0UA U265 ( .D(n42), .QTFCLK( ), .Q(fclkCntr[25]));
Q_MX02 U266 ( .S(initClock), .A0(fclkCntr[26]), .A1(n154), .Z(n43));
Q_FDP0UA U267 ( .D(n43), .QTFCLK( ), .Q(fclkCntr[26]));
Q_MX02 U268 ( .S(initClock), .A0(fclkCntr[27]), .A1(n152), .Z(n44));
Q_FDP0UA U269 ( .D(n44), .QTFCLK( ), .Q(fclkCntr[27]));
Q_MX02 U270 ( .S(initClock), .A0(fclkCntr[28]), .A1(n150), .Z(n45));
Q_FDP0UA U271 ( .D(n45), .QTFCLK( ), .Q(fclkCntr[28]));
Q_MX02 U272 ( .S(initClock), .A0(fclkCntr[29]), .A1(n148), .Z(n46));
Q_FDP0UA U273 ( .D(n46), .QTFCLK( ), .Q(fclkCntr[29]));
Q_MX02 U274 ( .S(initClock), .A0(fclkCntr[30]), .A1(n146), .Z(n47));
Q_FDP0UA U275 ( .D(n47), .QTFCLK( ), .Q(fclkCntr[30]));
Q_MX02 U276 ( .S(initClock), .A0(fclkCntr[31]), .A1(n144), .Z(n48));
Q_FDP0UA U277 ( .D(n48), .QTFCLK( ), .Q(fclkCntr[31]));
Q_MX02 U278 ( .S(initClock), .A0(fclkCntr[32]), .A1(n142), .Z(n49));
Q_FDP0UA U279 ( .D(n49), .QTFCLK( ), .Q(fclkCntr[32]));
Q_MX02 U280 ( .S(initClock), .A0(fclkCntr[33]), .A1(n140), .Z(n50));
Q_FDP0UA U281 ( .D(n50), .QTFCLK( ), .Q(fclkCntr[33]));
Q_MX02 U282 ( .S(initClock), .A0(fclkCntr[34]), .A1(n138), .Z(n51));
Q_FDP0UA U283 ( .D(n51), .QTFCLK( ), .Q(fclkCntr[34]));
Q_MX02 U284 ( .S(initClock), .A0(fclkCntr[35]), .A1(n136), .Z(n52));
Q_FDP0UA U285 ( .D(n52), .QTFCLK( ), .Q(fclkCntr[35]));
Q_MX02 U286 ( .S(initClock), .A0(fclkCntr[36]), .A1(n134), .Z(n53));
Q_FDP0UA U287 ( .D(n53), .QTFCLK( ), .Q(fclkCntr[36]));
Q_MX02 U288 ( .S(initClock), .A0(fclkCntr[37]), .A1(n132), .Z(n54));
Q_FDP0UA U289 ( .D(n54), .QTFCLK( ), .Q(fclkCntr[37]));
Q_MX02 U290 ( .S(initClock), .A0(fclkCntr[38]), .A1(n130), .Z(n55));
Q_FDP0UA U291 ( .D(n55), .QTFCLK( ), .Q(fclkCntr[38]));
Q_MX02 U292 ( .S(initClock), .A0(fclkCntr[39]), .A1(n128), .Z(n56));
Q_FDP0UA U293 ( .D(n56), .QTFCLK( ), .Q(fclkCntr[39]));
Q_MX02 U294 ( .S(initClock), .A0(fclkCntr[40]), .A1(n126), .Z(n57));
Q_FDP0UA U295 ( .D(n57), .QTFCLK( ), .Q(fclkCntr[40]));
Q_MX02 U296 ( .S(initClock), .A0(fclkCntr[41]), .A1(n124), .Z(n58));
Q_FDP0UA U297 ( .D(n58), .QTFCLK( ), .Q(fclkCntr[41]));
Q_MX02 U298 ( .S(initClock), .A0(fclkCntr[42]), .A1(n122), .Z(n59));
Q_FDP0UA U299 ( .D(n59), .QTFCLK( ), .Q(fclkCntr[42]));
Q_MX02 U300 ( .S(initClock), .A0(fclkCntr[43]), .A1(n120), .Z(n60));
Q_FDP0UA U301 ( .D(n60), .QTFCLK( ), .Q(fclkCntr[43]));
Q_MX02 U302 ( .S(initClock), .A0(fclkCntr[44]), .A1(n118), .Z(n61));
Q_FDP0UA U303 ( .D(n61), .QTFCLK( ), .Q(fclkCntr[44]));
Q_MX02 U304 ( .S(initClock), .A0(fclkCntr[45]), .A1(n116), .Z(n62));
Q_FDP0UA U305 ( .D(n62), .QTFCLK( ), .Q(fclkCntr[45]));
Q_MX02 U306 ( .S(initClock), .A0(fclkCntr[46]), .A1(n114), .Z(n63));
Q_FDP0UA U307 ( .D(n63), .QTFCLK( ), .Q(fclkCntr[46]));
Q_MX02 U308 ( .S(initClock), .A0(fclkCntr[47]), .A1(n112), .Z(n64));
Q_FDP0UA U309 ( .D(n64), .QTFCLK( ), .Q(fclkCntr[47]));
Q_MX02 U310 ( .S(initClock), .A0(fclkCntr[48]), .A1(n110), .Z(n65));
Q_FDP0UA U311 ( .D(n65), .QTFCLK( ), .Q(fclkCntr[48]));
Q_MX02 U312 ( .S(initClock), .A0(fclkCntr[49]), .A1(n108), .Z(n66));
Q_FDP0UA U313 ( .D(n66), .QTFCLK( ), .Q(fclkCntr[49]));
Q_MX02 U314 ( .S(initClock), .A0(fclkCntr[50]), .A1(n106), .Z(n67));
Q_FDP0UA U315 ( .D(n67), .QTFCLK( ), .Q(fclkCntr[50]));
Q_MX02 U316 ( .S(initClock), .A0(fclkCntr[51]), .A1(n104), .Z(n68));
Q_FDP0UA U317 ( .D(n68), .QTFCLK( ), .Q(fclkCntr[51]));
Q_MX02 U318 ( .S(initClock), .A0(fclkCntr[52]), .A1(n102), .Z(n69));
Q_FDP0UA U319 ( .D(n69), .QTFCLK( ), .Q(fclkCntr[52]));
Q_MX02 U320 ( .S(initClock), .A0(fclkCntr[53]), .A1(n100), .Z(n70));
Q_FDP0UA U321 ( .D(n70), .QTFCLK( ), .Q(fclkCntr[53]));
Q_MX02 U322 ( .S(initClock), .A0(fclkCntr[54]), .A1(n98), .Z(n71));
Q_FDP0UA U323 ( .D(n71), .QTFCLK( ), .Q(fclkCntr[54]));
Q_MX02 U324 ( .S(initClock), .A0(fclkCntr[55]), .A1(n96), .Z(n72));
Q_FDP0UA U325 ( .D(n72), .QTFCLK( ), .Q(fclkCntr[55]));
Q_MX02 U326 ( .S(initClock), .A0(fclkCntr[56]), .A1(n94), .Z(n73));
Q_FDP0UA U327 ( .D(n73), .QTFCLK( ), .Q(fclkCntr[56]));
Q_MX02 U328 ( .S(initClock), .A0(fclkCntr[57]), .A1(n92), .Z(n74));
Q_FDP0UA U329 ( .D(n74), .QTFCLK( ), .Q(fclkCntr[57]));
Q_MX02 U330 ( .S(initClock), .A0(fclkCntr[58]), .A1(n90), .Z(n75));
Q_FDP0UA U331 ( .D(n75), .QTFCLK( ), .Q(fclkCntr[58]));
Q_MX02 U332 ( .S(initClock), .A0(fclkCntr[59]), .A1(n88), .Z(n76));
Q_FDP0UA U333 ( .D(n76), .QTFCLK( ), .Q(fclkCntr[59]));
Q_MX02 U334 ( .S(initClock), .A0(fclkCntr[60]), .A1(n86), .Z(n77));
Q_FDP0UA U335 ( .D(n77), .QTFCLK( ), .Q(fclkCntr[60]));
Q_MX02 U336 ( .S(initClock), .A0(fclkCntr[61]), .A1(n84), .Z(n78));
Q_FDP0UA U337 ( .D(n78), .QTFCLK( ), .Q(fclkCntr[61]));
Q_MX02 U338 ( .S(initClock), .A0(fclkCntr[62]), .A1(n82), .Z(n79));
Q_FDP0UA U339 ( .D(n79), .QTFCLK( ), .Q(fclkCntr[62]));
Q_FDP0UA U340 ( .D(n80), .QTFCLK( ), .Q(fclkCntr[63]));
Q_XOR2 U341 ( .A0(fclkCntr[63]), .A1(n15), .Z(n80));
Q_AD01HF U342 ( .A0(fclkCntr[62]), .B0(n83), .S(n82), .CO(n81));
Q_AD01HF U343 ( .A0(fclkCntr[61]), .B0(n85), .S(n84), .CO(n83));
Q_AD01HF U344 ( .A0(fclkCntr[60]), .B0(n87), .S(n86), .CO(n85));
Q_AD01HF U345 ( .A0(fclkCntr[59]), .B0(n89), .S(n88), .CO(n87));
Q_AD01HF U346 ( .A0(fclkCntr[58]), .B0(n91), .S(n90), .CO(n89));
Q_AD01HF U347 ( .A0(fclkCntr[57]), .B0(n93), .S(n92), .CO(n91));
Q_AD01HF U348 ( .A0(fclkCntr[56]), .B0(n95), .S(n94), .CO(n93));
Q_AD01HF U349 ( .A0(fclkCntr[55]), .B0(n97), .S(n96), .CO(n95));
Q_AD01HF U350 ( .A0(fclkCntr[54]), .B0(n99), .S(n98), .CO(n97));
Q_AD01HF U351 ( .A0(fclkCntr[53]), .B0(n101), .S(n100), .CO(n99));
Q_AD01HF U352 ( .A0(fclkCntr[52]), .B0(n103), .S(n102), .CO(n101));
Q_AD01HF U353 ( .A0(fclkCntr[51]), .B0(n105), .S(n104), .CO(n103));
Q_AD01HF U354 ( .A0(fclkCntr[50]), .B0(n107), .S(n106), .CO(n105));
Q_AD01HF U355 ( .A0(fclkCntr[49]), .B0(n109), .S(n108), .CO(n107));
Q_AD01HF U356 ( .A0(fclkCntr[48]), .B0(n111), .S(n110), .CO(n109));
Q_AD01HF U357 ( .A0(fclkCntr[47]), .B0(n113), .S(n112), .CO(n111));
Q_AD01HF U358 ( .A0(fclkCntr[46]), .B0(n115), .S(n114), .CO(n113));
Q_AD01HF U359 ( .A0(fclkCntr[45]), .B0(n117), .S(n116), .CO(n115));
Q_AD01HF U360 ( .A0(fclkCntr[44]), .B0(n119), .S(n118), .CO(n117));
Q_AD01HF U361 ( .A0(fclkCntr[43]), .B0(n121), .S(n120), .CO(n119));
Q_AD01HF U362 ( .A0(fclkCntr[42]), .B0(n123), .S(n122), .CO(n121));
Q_AD01HF U363 ( .A0(fclkCntr[41]), .B0(n125), .S(n124), .CO(n123));
Q_AD01HF U364 ( .A0(fclkCntr[40]), .B0(n127), .S(n126), .CO(n125));
Q_AD01HF U365 ( .A0(fclkCntr[39]), .B0(n129), .S(n128), .CO(n127));
Q_AD01HF U366 ( .A0(fclkCntr[38]), .B0(n131), .S(n130), .CO(n129));
Q_AD01HF U367 ( .A0(fclkCntr[37]), .B0(n133), .S(n132), .CO(n131));
Q_AD01HF U368 ( .A0(fclkCntr[36]), .B0(n135), .S(n134), .CO(n133));
Q_AD01HF U369 ( .A0(fclkCntr[35]), .B0(n137), .S(n136), .CO(n135));
Q_AD01HF U370 ( .A0(fclkCntr[34]), .B0(n139), .S(n138), .CO(n137));
Q_AD01HF U371 ( .A0(fclkCntr[33]), .B0(n141), .S(n140), .CO(n139));
Q_AD01HF U372 ( .A0(fclkCntr[32]), .B0(n143), .S(n142), .CO(n141));
Q_AD01HF U373 ( .A0(fclkCntr[31]), .B0(n145), .S(n144), .CO(n143));
Q_AD01HF U374 ( .A0(fclkCntr[30]), .B0(n147), .S(n146), .CO(n145));
Q_AD01HF U375 ( .A0(fclkCntr[29]), .B0(n149), .S(n148), .CO(n147));
Q_AD01HF U376 ( .A0(fclkCntr[28]), .B0(n151), .S(n150), .CO(n149));
Q_AD01HF U377 ( .A0(fclkCntr[27]), .B0(n153), .S(n152), .CO(n151));
Q_AD01HF U378 ( .A0(fclkCntr[26]), .B0(n155), .S(n154), .CO(n153));
Q_AD01HF U379 ( .A0(fclkCntr[25]), .B0(n157), .S(n156), .CO(n155));
Q_AD01HF U380 ( .A0(fclkCntr[24]), .B0(n159), .S(n158), .CO(n157));
Q_AD01HF U381 ( .A0(fclkCntr[23]), .B0(n161), .S(n160), .CO(n159));
Q_AD01HF U382 ( .A0(fclkCntr[22]), .B0(n163), .S(n162), .CO(n161));
Q_AD01HF U383 ( .A0(fclkCntr[21]), .B0(n165), .S(n164), .CO(n163));
Q_AD01HF U384 ( .A0(fclkCntr[20]), .B0(n167), .S(n166), .CO(n165));
Q_AD01HF U385 ( .A0(fclkCntr[19]), .B0(n169), .S(n168), .CO(n167));
Q_AD01HF U386 ( .A0(fclkCntr[18]), .B0(n171), .S(n170), .CO(n169));
Q_AD01HF U387 ( .A0(fclkCntr[17]), .B0(n173), .S(n172), .CO(n171));
Q_AD01HF U388 ( .A0(fclkCntr[16]), .B0(n175), .S(n174), .CO(n173));
Q_AD01HF U389 ( .A0(fclkCntr[15]), .B0(n177), .S(n176), .CO(n175));
Q_AD01HF U390 ( .A0(fclkCntr[14]), .B0(n179), .S(n178), .CO(n177));
Q_AD01HF U391 ( .A0(fclkCntr[13]), .B0(n181), .S(n180), .CO(n179));
Q_AD01HF U392 ( .A0(fclkCntr[12]), .B0(n183), .S(n182), .CO(n181));
Q_AD01HF U393 ( .A0(fclkCntr[11]), .B0(n185), .S(n184), .CO(n183));
Q_AD01HF U394 ( .A0(fclkCntr[10]), .B0(n187), .S(n186), .CO(n185));
Q_AD01HF U395 ( .A0(fclkCntr[9]), .B0(n189), .S(n188), .CO(n187));
Q_AD01HF U396 ( .A0(fclkCntr[8]), .B0(n191), .S(n190), .CO(n189));
Q_AD01HF U397 ( .A0(fclkCntr[7]), .B0(n193), .S(n192), .CO(n191));
Q_AD01HF U398 ( .A0(fclkCntr[6]), .B0(n195), .S(n194), .CO(n193));
Q_AD01HF U399 ( .A0(fclkCntr[5]), .B0(n197), .S(n196), .CO(n195));
Q_AD01HF U400 ( .A0(fclkCntr[4]), .B0(n199), .S(n198), .CO(n197));
Q_AD01HF U401 ( .A0(fclkCntr[3]), .B0(n201), .S(n200), .CO(n199));
Q_AD01HF U402 ( .A0(fclkCntr[2]), .B0(n203), .S(n202), .CO(n201));
Q_AD01HF U403 ( .A0(fclkCntr[1]), .B0(fclkCntr[0]), .S(n204), .CO(n203));
Q_OA21 U404 ( .A0(n206), .A1(n205), .B0(n299), .Z(n16));
Q_OR03 U405 ( .A0(n209), .A1(n208), .A2(n207), .Z(n205));
Q_OR03 U406 ( .A0(n212), .A1(n211), .A2(n210), .Z(n206));
Q_OR03 U407 ( .A0(n215), .A1(n214), .A2(n213), .Z(n207));
Q_OR03 U408 ( .A0(n218), .A1(n217), .A2(n216), .Z(n208));
Q_OR03 U409 ( .A0(n221), .A1(n220), .A2(n219), .Z(n209));
Q_OR03 U410 ( .A0(n224), .A1(n223), .A2(n222), .Z(n210));
Q_OR03 U411 ( .A0(n227), .A1(n226), .A2(n225), .Z(n211));
Q_OR03 U412 ( .A0(n230), .A1(n229), .A2(n228), .Z(n212));
Q_OR03 U413 ( .A0(n233), .A1(n232), .A2(n231), .Z(n213));
Q_OR03 U414 ( .A0(n298), .A1(n235), .A2(n234), .Z(n214));
Q_OR03 U415 ( .A0(n295), .A1(n296), .A2(n297), .Z(n215));
Q_OR03 U416 ( .A0(n292), .A1(n293), .A2(n294), .Z(n216));
Q_OR03 U417 ( .A0(n289), .A1(n290), .A2(n291), .Z(n217));
Q_OR03 U418 ( .A0(n286), .A1(n287), .A2(n288), .Z(n218));
Q_OR03 U419 ( .A0(n283), .A1(n284), .A2(n285), .Z(n219));
Q_OR03 U420 ( .A0(n280), .A1(n281), .A2(n282), .Z(n220));
Q_OR03 U421 ( .A0(n277), .A1(n278), .A2(n279), .Z(n221));
Q_OR03 U422 ( .A0(n274), .A1(n275), .A2(n276), .Z(n222));
Q_OR03 U423 ( .A0(n271), .A1(n272), .A2(n273), .Z(n223));
Q_OR03 U424 ( .A0(n268), .A1(n269), .A2(n270), .Z(n224));
Q_OR03 U425 ( .A0(n265), .A1(n266), .A2(n267), .Z(n225));
Q_OR03 U426 ( .A0(n262), .A1(n263), .A2(n264), .Z(n226));
Q_OR03 U427 ( .A0(n259), .A1(n260), .A2(n261), .Z(n227));
Q_OR03 U428 ( .A0(n256), .A1(n257), .A2(n258), .Z(n228));
Q_OR03 U429 ( .A0(n253), .A1(n254), .A2(n255), .Z(n229));
Q_OR03 U430 ( .A0(n250), .A1(n251), .A2(n252), .Z(n230));
Q_OR03 U431 ( .A0(n247), .A1(n248), .A2(n249), .Z(n231));
Q_OR03 U432 ( .A0(n244), .A1(n245), .A2(n246), .Z(n232));
Q_OR03 U433 ( .A0(n241), .A1(n242), .A2(n243), .Z(n233));
Q_OR03 U434 ( .A0(n238), .A1(n239), .A2(n240), .Z(n234));
Q_OR03 U435 ( .A0(uClkCntr[63]), .A1(n236), .A2(n237), .Z(n235));
Q_XOR2 U436 ( .A0(fclkCntr[63]), .A1(uClkCntr[62]), .Z(n236));
Q_XOR2 U437 ( .A0(fclkCntr[62]), .A1(uClkCntr[61]), .Z(n237));
Q_XOR2 U438 ( .A0(fclkCntr[61]), .A1(uClkCntr[60]), .Z(n238));
Q_XOR2 U439 ( .A0(fclkCntr[60]), .A1(uClkCntr[59]), .Z(n239));
Q_XOR2 U440 ( .A0(fclkCntr[59]), .A1(uClkCntr[58]), .Z(n240));
Q_XOR2 U441 ( .A0(fclkCntr[58]), .A1(uClkCntr[57]), .Z(n241));
Q_XOR2 U442 ( .A0(fclkCntr[57]), .A1(uClkCntr[56]), .Z(n242));
Q_XOR2 U443 ( .A0(fclkCntr[56]), .A1(uClkCntr[55]), .Z(n243));
Q_XOR2 U444 ( .A0(fclkCntr[55]), .A1(uClkCntr[54]), .Z(n244));
Q_XOR2 U445 ( .A0(fclkCntr[54]), .A1(uClkCntr[53]), .Z(n245));
Q_XOR2 U446 ( .A0(fclkCntr[53]), .A1(uClkCntr[52]), .Z(n246));
Q_XOR2 U447 ( .A0(fclkCntr[52]), .A1(uClkCntr[51]), .Z(n247));
Q_XOR2 U448 ( .A0(fclkCntr[51]), .A1(uClkCntr[50]), .Z(n248));
Q_XOR2 U449 ( .A0(fclkCntr[50]), .A1(uClkCntr[49]), .Z(n249));
Q_XOR2 U450 ( .A0(fclkCntr[49]), .A1(uClkCntr[48]), .Z(n250));
Q_XOR2 U451 ( .A0(fclkCntr[48]), .A1(uClkCntr[47]), .Z(n251));
Q_XOR2 U452 ( .A0(fclkCntr[47]), .A1(uClkCntr[46]), .Z(n252));
Q_XOR2 U453 ( .A0(fclkCntr[46]), .A1(uClkCntr[45]), .Z(n253));
Q_XOR2 U454 ( .A0(fclkCntr[45]), .A1(uClkCntr[44]), .Z(n254));
Q_XOR2 U455 ( .A0(fclkCntr[44]), .A1(uClkCntr[43]), .Z(n255));
Q_XOR2 U456 ( .A0(fclkCntr[43]), .A1(uClkCntr[42]), .Z(n256));
Q_XOR2 U457 ( .A0(fclkCntr[42]), .A1(uClkCntr[41]), .Z(n257));
Q_XOR2 U458 ( .A0(fclkCntr[41]), .A1(uClkCntr[40]), .Z(n258));
Q_XOR2 U459 ( .A0(fclkCntr[40]), .A1(uClkCntr[39]), .Z(n259));
Q_XOR2 U460 ( .A0(fclkCntr[39]), .A1(uClkCntr[38]), .Z(n260));
Q_XOR2 U461 ( .A0(fclkCntr[38]), .A1(uClkCntr[37]), .Z(n261));
Q_XOR2 U462 ( .A0(fclkCntr[37]), .A1(uClkCntr[36]), .Z(n262));
Q_XOR2 U463 ( .A0(fclkCntr[36]), .A1(uClkCntr[35]), .Z(n263));
Q_XOR2 U464 ( .A0(fclkCntr[35]), .A1(uClkCntr[34]), .Z(n264));
Q_XOR2 U465 ( .A0(fclkCntr[34]), .A1(uClkCntr[33]), .Z(n265));
Q_XOR2 U466 ( .A0(fclkCntr[33]), .A1(uClkCntr[32]), .Z(n266));
Q_XOR2 U467 ( .A0(fclkCntr[32]), .A1(uClkCntr[31]), .Z(n267));
Q_XOR2 U468 ( .A0(fclkCntr[31]), .A1(uClkCntr[30]), .Z(n268));
Q_XOR2 U469 ( .A0(fclkCntr[30]), .A1(uClkCntr[29]), .Z(n269));
Q_XOR2 U470 ( .A0(fclkCntr[29]), .A1(uClkCntr[28]), .Z(n270));
Q_XOR2 U471 ( .A0(fclkCntr[28]), .A1(uClkCntr[27]), .Z(n271));
Q_XOR2 U472 ( .A0(fclkCntr[27]), .A1(uClkCntr[26]), .Z(n272));
Q_XOR2 U473 ( .A0(fclkCntr[26]), .A1(uClkCntr[25]), .Z(n273));
Q_XOR2 U474 ( .A0(fclkCntr[25]), .A1(uClkCntr[24]), .Z(n274));
Q_XOR2 U475 ( .A0(fclkCntr[24]), .A1(uClkCntr[23]), .Z(n275));
Q_XOR2 U476 ( .A0(fclkCntr[23]), .A1(uClkCntr[22]), .Z(n276));
Q_XOR2 U477 ( .A0(fclkCntr[22]), .A1(uClkCntr[21]), .Z(n277));
Q_XOR2 U478 ( .A0(fclkCntr[21]), .A1(uClkCntr[20]), .Z(n278));
Q_XOR2 U479 ( .A0(fclkCntr[20]), .A1(uClkCntr[19]), .Z(n279));
Q_XOR2 U480 ( .A0(fclkCntr[19]), .A1(uClkCntr[18]), .Z(n280));
Q_XOR2 U481 ( .A0(fclkCntr[18]), .A1(uClkCntr[17]), .Z(n281));
Q_XOR2 U482 ( .A0(fclkCntr[17]), .A1(uClkCntr[16]), .Z(n282));
Q_XOR2 U483 ( .A0(fclkCntr[16]), .A1(uClkCntr[15]), .Z(n283));
Q_XOR2 U484 ( .A0(fclkCntr[15]), .A1(uClkCntr[14]), .Z(n284));
Q_XOR2 U485 ( .A0(fclkCntr[14]), .A1(uClkCntr[13]), .Z(n285));
Q_XOR2 U486 ( .A0(fclkCntr[13]), .A1(uClkCntr[12]), .Z(n286));
Q_XOR2 U487 ( .A0(fclkCntr[12]), .A1(uClkCntr[11]), .Z(n287));
Q_XOR2 U488 ( .A0(fclkCntr[11]), .A1(uClkCntr[10]), .Z(n288));
Q_XOR2 U489 ( .A0(fclkCntr[10]), .A1(uClkCntr[9]), .Z(n289));
Q_XOR2 U490 ( .A0(fclkCntr[9]), .A1(uClkCntr[8]), .Z(n290));
Q_XOR2 U491 ( .A0(fclkCntr[8]), .A1(uClkCntr[7]), .Z(n291));
Q_XOR2 U492 ( .A0(fclkCntr[7]), .A1(uClkCntr[6]), .Z(n292));
Q_XOR2 U493 ( .A0(fclkCntr[6]), .A1(uClkCntr[5]), .Z(n293));
Q_XOR2 U494 ( .A0(fclkCntr[5]), .A1(uClkCntr[4]), .Z(n294));
Q_XOR2 U495 ( .A0(fclkCntr[4]), .A1(uClkCntr[3]), .Z(n295));
Q_XOR2 U496 ( .A0(fclkCntr[3]), .A1(uClkCntr[2]), .Z(n296));
Q_XOR2 U497 ( .A0(fclkCntr[2]), .A1(uClkCntr[1]), .Z(n297));
Q_XOR2 U498 ( .A0(fclkCntr[1]), .A1(uClkCntr[0]), .Z(n298));
Q_NR02 U499 ( .A0(n301), .A1(n300), .Z(n299));
Q_OR03 U500 ( .A0(n304), .A1(n303), .A2(n302), .Z(n300));
Q_OR03 U501 ( .A0(n307), .A1(n306), .A2(n305), .Z(n301));
Q_OR03 U502 ( .A0(n310), .A1(n309), .A2(n308), .Z(n302));
Q_OR03 U503 ( .A0(n313), .A1(n312), .A2(n311), .Z(n303));
Q_OR03 U504 ( .A0(n316), .A1(n315), .A2(n314), .Z(n304));
Q_OR03 U505 ( .A0(n319), .A1(n318), .A2(n317), .Z(n305));
Q_OR03 U506 ( .A0(n322), .A1(n321), .A2(n320), .Z(n306));
Q_OR03 U507 ( .A0(n325), .A1(n324), .A2(n323), .Z(n307));
Q_OR03 U508 ( .A0(n328), .A1(n327), .A2(n326), .Z(n308));
Q_OR03 U509 ( .A0(uClkErrTime[0]), .A1(n330), .A2(n329), .Z(n309));
Q_OR03 U510 ( .A0(uClkErrTime[3]), .A1(uClkErrTime[2]), .A2(uClkErrTime[1]), .Z(n310));
Q_OR03 U511 ( .A0(uClkErrTime[6]), .A1(uClkErrTime[5]), .A2(uClkErrTime[4]), .Z(n311));
Q_OR03 U512 ( .A0(uClkErrTime[9]), .A1(uClkErrTime[8]), .A2(uClkErrTime[7]), .Z(n312));
Q_OR03 U513 ( .A0(uClkErrTime[12]), .A1(uClkErrTime[11]), .A2(uClkErrTime[10]), .Z(n313));
Q_OR03 U514 ( .A0(uClkErrTime[15]), .A1(uClkErrTime[14]), .A2(uClkErrTime[13]), .Z(n314));
Q_OR03 U515 ( .A0(uClkErrTime[18]), .A1(uClkErrTime[17]), .A2(uClkErrTime[16]), .Z(n315));
Q_OR03 U516 ( .A0(uClkErrTime[21]), .A1(uClkErrTime[20]), .A2(uClkErrTime[19]), .Z(n316));
Q_OR03 U517 ( .A0(uClkErrTime[24]), .A1(uClkErrTime[23]), .A2(uClkErrTime[22]), .Z(n317));
Q_OR03 U518 ( .A0(uClkErrTime[27]), .A1(uClkErrTime[26]), .A2(uClkErrTime[25]), .Z(n318));
Q_OR03 U519 ( .A0(uClkErrTime[30]), .A1(uClkErrTime[29]), .A2(uClkErrTime[28]), .Z(n319));
Q_OR03 U520 ( .A0(uClkErrTime[33]), .A1(uClkErrTime[32]), .A2(uClkErrTime[31]), .Z(n320));
Q_OR03 U521 ( .A0(uClkErrTime[36]), .A1(uClkErrTime[35]), .A2(uClkErrTime[34]), .Z(n321));
Q_OR03 U522 ( .A0(uClkErrTime[39]), .A1(uClkErrTime[38]), .A2(uClkErrTime[37]), .Z(n322));
Q_OR03 U523 ( .A0(uClkErrTime[42]), .A1(uClkErrTime[41]), .A2(uClkErrTime[40]), .Z(n323));
Q_OR03 U524 ( .A0(uClkErrTime[45]), .A1(uClkErrTime[44]), .A2(uClkErrTime[43]), .Z(n324));
Q_OR03 U525 ( .A0(uClkErrTime[48]), .A1(uClkErrTime[47]), .A2(uClkErrTime[46]), .Z(n325));
Q_OR03 U526 ( .A0(uClkErrTime[51]), .A1(uClkErrTime[50]), .A2(uClkErrTime[49]), .Z(n326));
Q_OR03 U527 ( .A0(uClkErrTime[54]), .A1(uClkErrTime[53]), .A2(uClkErrTime[52]), .Z(n327));
Q_OR03 U528 ( .A0(uClkErrTime[57]), .A1(uClkErrTime[56]), .A2(uClkErrTime[55]), .Z(n328));
Q_OR03 U529 ( .A0(uClkErrTime[60]), .A1(uClkErrTime[59]), .A2(uClkErrTime[58]), .Z(n329));
Q_OR03 U530 ( .A0(uClkErrTime[63]), .A1(uClkErrTime[62]), .A2(uClkErrTime[61]), .Z(n330));
Q_MX02 U531 ( .S(n16), .A0(uClkErrTime[0]), .A1(simTime[0]), .Z(n331));
Q_FDP0UA U532 ( .D(n331), .QTFCLK( ), .Q(uClkErrTime[0]));
Q_MX02 U533 ( .S(n16), .A0(uClkErrTime[1]), .A1(simTime[1]), .Z(n332));
Q_FDP0UA U534 ( .D(n332), .QTFCLK( ), .Q(uClkErrTime[1]));
Q_MX02 U535 ( .S(n16), .A0(uClkErrTime[2]), .A1(simTime[2]), .Z(n333));
Q_FDP0UA U536 ( .D(n333), .QTFCLK( ), .Q(uClkErrTime[2]));
Q_MX02 U537 ( .S(n16), .A0(uClkErrTime[3]), .A1(simTime[3]), .Z(n334));
Q_FDP0UA U538 ( .D(n334), .QTFCLK( ), .Q(uClkErrTime[3]));
Q_MX02 U539 ( .S(n16), .A0(uClkErrTime[4]), .A1(simTime[4]), .Z(n335));
Q_FDP0UA U540 ( .D(n335), .QTFCLK( ), .Q(uClkErrTime[4]));
Q_MX02 U541 ( .S(n16), .A0(uClkErrTime[5]), .A1(simTime[5]), .Z(n336));
Q_FDP0UA U542 ( .D(n336), .QTFCLK( ), .Q(uClkErrTime[5]));
Q_MX02 U543 ( .S(n16), .A0(uClkErrTime[6]), .A1(simTime[6]), .Z(n337));
Q_FDP0UA U544 ( .D(n337), .QTFCLK( ), .Q(uClkErrTime[6]));
Q_MX02 U545 ( .S(n16), .A0(uClkErrTime[7]), .A1(simTime[7]), .Z(n338));
Q_FDP0UA U546 ( .D(n338), .QTFCLK( ), .Q(uClkErrTime[7]));
Q_MX02 U547 ( .S(n16), .A0(uClkErrTime[8]), .A1(simTime[8]), .Z(n339));
Q_FDP0UA U548 ( .D(n339), .QTFCLK( ), .Q(uClkErrTime[8]));
Q_MX02 U549 ( .S(n16), .A0(uClkErrTime[9]), .A1(simTime[9]), .Z(n340));
Q_FDP0UA U550 ( .D(n340), .QTFCLK( ), .Q(uClkErrTime[9]));
Q_MX02 U551 ( .S(n16), .A0(uClkErrTime[10]), .A1(simTime[10]), .Z(n341));
Q_FDP0UA U552 ( .D(n341), .QTFCLK( ), .Q(uClkErrTime[10]));
Q_MX02 U553 ( .S(n16), .A0(uClkErrTime[11]), .A1(simTime[11]), .Z(n342));
Q_FDP0UA U554 ( .D(n342), .QTFCLK( ), .Q(uClkErrTime[11]));
Q_MX02 U555 ( .S(n16), .A0(uClkErrTime[12]), .A1(simTime[12]), .Z(n343));
Q_FDP0UA U556 ( .D(n343), .QTFCLK( ), .Q(uClkErrTime[12]));
Q_MX02 U557 ( .S(n16), .A0(uClkErrTime[13]), .A1(simTime[13]), .Z(n344));
Q_FDP0UA U558 ( .D(n344), .QTFCLK( ), .Q(uClkErrTime[13]));
Q_MX02 U559 ( .S(n16), .A0(uClkErrTime[14]), .A1(simTime[14]), .Z(n345));
Q_FDP0UA U560 ( .D(n345), .QTFCLK( ), .Q(uClkErrTime[14]));
Q_MX02 U561 ( .S(n16), .A0(uClkErrTime[15]), .A1(simTime[15]), .Z(n346));
Q_FDP0UA U562 ( .D(n346), .QTFCLK( ), .Q(uClkErrTime[15]));
Q_MX02 U563 ( .S(n16), .A0(uClkErrTime[16]), .A1(simTime[16]), .Z(n347));
Q_FDP0UA U564 ( .D(n347), .QTFCLK( ), .Q(uClkErrTime[16]));
Q_MX02 U565 ( .S(n16), .A0(uClkErrTime[17]), .A1(simTime[17]), .Z(n348));
Q_FDP0UA U566 ( .D(n348), .QTFCLK( ), .Q(uClkErrTime[17]));
Q_MX02 U567 ( .S(n16), .A0(uClkErrTime[18]), .A1(simTime[18]), .Z(n349));
Q_FDP0UA U568 ( .D(n349), .QTFCLK( ), .Q(uClkErrTime[18]));
Q_MX02 U569 ( .S(n16), .A0(uClkErrTime[19]), .A1(simTime[19]), .Z(n350));
Q_FDP0UA U570 ( .D(n350), .QTFCLK( ), .Q(uClkErrTime[19]));
Q_MX02 U571 ( .S(n16), .A0(uClkErrTime[20]), .A1(simTime[20]), .Z(n351));
Q_FDP0UA U572 ( .D(n351), .QTFCLK( ), .Q(uClkErrTime[20]));
Q_MX02 U573 ( .S(n16), .A0(uClkErrTime[21]), .A1(simTime[21]), .Z(n352));
Q_FDP0UA U574 ( .D(n352), .QTFCLK( ), .Q(uClkErrTime[21]));
Q_MX02 U575 ( .S(n16), .A0(uClkErrTime[22]), .A1(simTime[22]), .Z(n353));
Q_FDP0UA U576 ( .D(n353), .QTFCLK( ), .Q(uClkErrTime[22]));
Q_MX02 U577 ( .S(n16), .A0(uClkErrTime[23]), .A1(simTime[23]), .Z(n354));
Q_FDP0UA U578 ( .D(n354), .QTFCLK( ), .Q(uClkErrTime[23]));
Q_MX02 U579 ( .S(n16), .A0(uClkErrTime[24]), .A1(simTime[24]), .Z(n355));
Q_FDP0UA U580 ( .D(n355), .QTFCLK( ), .Q(uClkErrTime[24]));
Q_MX02 U581 ( .S(n16), .A0(uClkErrTime[25]), .A1(simTime[25]), .Z(n356));
Q_FDP0UA U582 ( .D(n356), .QTFCLK( ), .Q(uClkErrTime[25]));
Q_MX02 U583 ( .S(n16), .A0(uClkErrTime[26]), .A1(simTime[26]), .Z(n357));
Q_FDP0UA U584 ( .D(n357), .QTFCLK( ), .Q(uClkErrTime[26]));
Q_MX02 U585 ( .S(n16), .A0(uClkErrTime[27]), .A1(simTime[27]), .Z(n358));
Q_FDP0UA U586 ( .D(n358), .QTFCLK( ), .Q(uClkErrTime[27]));
Q_MX02 U587 ( .S(n16), .A0(uClkErrTime[28]), .A1(simTime[28]), .Z(n359));
Q_FDP0UA U588 ( .D(n359), .QTFCLK( ), .Q(uClkErrTime[28]));
Q_MX02 U589 ( .S(n16), .A0(uClkErrTime[29]), .A1(simTime[29]), .Z(n360));
Q_FDP0UA U590 ( .D(n360), .QTFCLK( ), .Q(uClkErrTime[29]));
Q_MX02 U591 ( .S(n16), .A0(uClkErrTime[30]), .A1(simTime[30]), .Z(n361));
Q_FDP0UA U592 ( .D(n361), .QTFCLK( ), .Q(uClkErrTime[30]));
Q_MX02 U593 ( .S(n16), .A0(uClkErrTime[31]), .A1(simTime[31]), .Z(n362));
Q_FDP0UA U594 ( .D(n362), .QTFCLK( ), .Q(uClkErrTime[31]));
Q_MX02 U595 ( .S(n16), .A0(uClkErrTime[32]), .A1(simTime[32]), .Z(n363));
Q_FDP0UA U596 ( .D(n363), .QTFCLK( ), .Q(uClkErrTime[32]));
Q_MX02 U597 ( .S(n16), .A0(uClkErrTime[33]), .A1(simTime[33]), .Z(n364));
Q_FDP0UA U598 ( .D(n364), .QTFCLK( ), .Q(uClkErrTime[33]));
Q_MX02 U599 ( .S(n16), .A0(uClkErrTime[34]), .A1(simTime[34]), .Z(n365));
Q_FDP0UA U600 ( .D(n365), .QTFCLK( ), .Q(uClkErrTime[34]));
Q_MX02 U601 ( .S(n16), .A0(uClkErrTime[35]), .A1(simTime[35]), .Z(n366));
Q_FDP0UA U602 ( .D(n366), .QTFCLK( ), .Q(uClkErrTime[35]));
Q_MX02 U603 ( .S(n16), .A0(uClkErrTime[36]), .A1(simTime[36]), .Z(n367));
Q_FDP0UA U604 ( .D(n367), .QTFCLK( ), .Q(uClkErrTime[36]));
Q_MX02 U605 ( .S(n16), .A0(uClkErrTime[37]), .A1(simTime[37]), .Z(n368));
Q_FDP0UA U606 ( .D(n368), .QTFCLK( ), .Q(uClkErrTime[37]));
Q_MX02 U607 ( .S(n16), .A0(uClkErrTime[38]), .A1(simTime[38]), .Z(n369));
Q_FDP0UA U608 ( .D(n369), .QTFCLK( ), .Q(uClkErrTime[38]));
Q_MX02 U609 ( .S(n16), .A0(uClkErrTime[39]), .A1(simTime[39]), .Z(n370));
Q_FDP0UA U610 ( .D(n370), .QTFCLK( ), .Q(uClkErrTime[39]));
Q_MX02 U611 ( .S(n16), .A0(uClkErrTime[40]), .A1(simTime[40]), .Z(n371));
Q_FDP0UA U612 ( .D(n371), .QTFCLK( ), .Q(uClkErrTime[40]));
Q_MX02 U613 ( .S(n16), .A0(uClkErrTime[41]), .A1(simTime[41]), .Z(n372));
Q_FDP0UA U614 ( .D(n372), .QTFCLK( ), .Q(uClkErrTime[41]));
Q_MX02 U615 ( .S(n16), .A0(uClkErrTime[42]), .A1(simTime[42]), .Z(n373));
Q_FDP0UA U616 ( .D(n373), .QTFCLK( ), .Q(uClkErrTime[42]));
Q_MX02 U617 ( .S(n16), .A0(uClkErrTime[43]), .A1(simTime[43]), .Z(n374));
Q_FDP0UA U618 ( .D(n374), .QTFCLK( ), .Q(uClkErrTime[43]));
Q_MX02 U619 ( .S(n16), .A0(uClkErrTime[44]), .A1(simTime[44]), .Z(n375));
Q_FDP0UA U620 ( .D(n375), .QTFCLK( ), .Q(uClkErrTime[44]));
Q_MX02 U621 ( .S(n16), .A0(uClkErrTime[45]), .A1(simTime[45]), .Z(n376));
Q_FDP0UA U622 ( .D(n376), .QTFCLK( ), .Q(uClkErrTime[45]));
Q_MX02 U623 ( .S(n16), .A0(uClkErrTime[46]), .A1(simTime[46]), .Z(n377));
Q_FDP0UA U624 ( .D(n377), .QTFCLK( ), .Q(uClkErrTime[46]));
Q_MX02 U625 ( .S(n16), .A0(uClkErrTime[47]), .A1(simTime[47]), .Z(n378));
Q_FDP0UA U626 ( .D(n378), .QTFCLK( ), .Q(uClkErrTime[47]));
Q_MX02 U627 ( .S(n16), .A0(uClkErrTime[48]), .A1(simTime[48]), .Z(n379));
Q_FDP0UA U628 ( .D(n379), .QTFCLK( ), .Q(uClkErrTime[48]));
Q_MX02 U629 ( .S(n16), .A0(uClkErrTime[49]), .A1(simTime[49]), .Z(n380));
Q_FDP0UA U630 ( .D(n380), .QTFCLK( ), .Q(uClkErrTime[49]));
Q_MX02 U631 ( .S(n16), .A0(uClkErrTime[50]), .A1(simTime[50]), .Z(n381));
Q_FDP0UA U632 ( .D(n381), .QTFCLK( ), .Q(uClkErrTime[50]));
Q_MX02 U633 ( .S(n16), .A0(uClkErrTime[51]), .A1(simTime[51]), .Z(n382));
Q_FDP0UA U634 ( .D(n382), .QTFCLK( ), .Q(uClkErrTime[51]));
Q_MX02 U635 ( .S(n16), .A0(uClkErrTime[52]), .A1(simTime[52]), .Z(n383));
Q_FDP0UA U636 ( .D(n383), .QTFCLK( ), .Q(uClkErrTime[52]));
Q_MX02 U637 ( .S(n16), .A0(uClkErrTime[53]), .A1(simTime[53]), .Z(n384));
Q_FDP0UA U638 ( .D(n384), .QTFCLK( ), .Q(uClkErrTime[53]));
Q_MX02 U639 ( .S(n16), .A0(uClkErrTime[54]), .A1(simTime[54]), .Z(n385));
Q_FDP0UA U640 ( .D(n385), .QTFCLK( ), .Q(uClkErrTime[54]));
Q_MX02 U641 ( .S(n16), .A0(uClkErrTime[55]), .A1(simTime[55]), .Z(n386));
Q_FDP0UA U642 ( .D(n386), .QTFCLK( ), .Q(uClkErrTime[55]));
Q_MX02 U643 ( .S(n16), .A0(uClkErrTime[56]), .A1(simTime[56]), .Z(n387));
Q_FDP0UA U644 ( .D(n387), .QTFCLK( ), .Q(uClkErrTime[56]));
Q_MX02 U645 ( .S(n16), .A0(uClkErrTime[57]), .A1(simTime[57]), .Z(n388));
Q_FDP0UA U646 ( .D(n388), .QTFCLK( ), .Q(uClkErrTime[57]));
Q_MX02 U647 ( .S(n16), .A0(uClkErrTime[58]), .A1(simTime[58]), .Z(n389));
Q_FDP0UA U648 ( .D(n389), .QTFCLK( ), .Q(uClkErrTime[58]));
Q_MX02 U649 ( .S(n16), .A0(uClkErrTime[59]), .A1(simTime[59]), .Z(n390));
Q_FDP0UA U650 ( .D(n390), .QTFCLK( ), .Q(uClkErrTime[59]));
Q_MX02 U651 ( .S(n16), .A0(uClkErrTime[60]), .A1(simTime[60]), .Z(n391));
Q_FDP0UA U652 ( .D(n391), .QTFCLK( ), .Q(uClkErrTime[60]));
Q_MX02 U653 ( .S(n16), .A0(uClkErrTime[61]), .A1(simTime[61]), .Z(n392));
Q_FDP0UA U654 ( .D(n392), .QTFCLK( ), .Q(uClkErrTime[61]));
Q_MX02 U655 ( .S(n16), .A0(uClkErrTime[62]), .A1(simTime[62]), .Z(n393));
Q_FDP0UA U656 ( .D(n393), .QTFCLK( ), .Q(uClkErrTime[62]));
Q_MX02 U657 ( .S(n16), .A0(uClkErrTime[63]), .A1(simTime[63]), .Z(n394));
Q_FDP0UA U658 ( .D(n394), .QTFCLK( ), .Q(uClkErrTime[63]));
Q_INV U659 ( .A(holdEcmTb), .Z(n395));
Q_AN02 U660 ( .A0(n395), .A1(n3667), .Z(n396));
Q_MX02 U661 ( .S(n396), .A0(holdEcmTb), .A1(holdEcmSync), .Z(n397));
Q_FDP0UA U662 ( .D(n397), .QTFCLK( ), .Q(holdEcmSync));
Q_FDP0UA U663 ( .D(ecmNotSync), .QTFCLK( ), .Q(ecmNotSyncD));
Q_FDP0UA U664 ( .D(ecmOn), .QTFCLK( ), .Q(ecmOnD));
Q_FDP0UA U665 ( .D(anyStop), .QTFCLK( ), .Q(ptxStop));
Q_FDP0UA U666 ( .D(maxFck2Sync[15]), .QTFCLK( ), .Q(maxFck2Sync[15]));
Q_FDP0UA U667 ( .D(maxFck2Sync[14]), .QTFCLK( ), .Q(maxFck2Sync[14]));
Q_FDP0UA U668 ( .D(maxFck2Sync[13]), .QTFCLK( ), .Q(maxFck2Sync[13]));
Q_FDP0UA U669 ( .D(maxFck2Sync[12]), .QTFCLK( ), .Q(maxFck2Sync[12]));
Q_FDP0UA U670 ( .D(maxFck2Sync[11]), .QTFCLK( ), .Q(maxFck2Sync[11]));
Q_FDP0UA U671 ( .D(maxFck2Sync[10]), .QTFCLK( ), .Q(maxFck2Sync[10]));
Q_FDP0UA U672 ( .D(maxFck2Sync[9]), .QTFCLK( ), .Q(maxFck2Sync[9]));
Q_FDP0UA U673 ( .D(maxFck2Sync[8]), .QTFCLK( ), .Q(maxFck2Sync[8]));
Q_FDP0UA U674 ( .D(maxFck2Sync[7]), .QTFCLK( ), .Q(maxFck2Sync[7]));
Q_FDP0UA U675 ( .D(maxFck2Sync[6]), .QTFCLK( ), .Q(maxFck2Sync[6]));
Q_FDP0UA U676 ( .D(maxFck2Sync[5]), .QTFCLK( ), .Q(maxFck2Sync[5]));
Q_FDP0UA U677 ( .D(maxFck2Sync[4]), .QTFCLK( ), .Q(maxFck2Sync[4]));
Q_FDP0UA U678 ( .D(maxFck2Sync[3]), .QTFCLK( ), .Q(maxFck2Sync[3]));
Q_FDP0UA U679 ( .D(maxFck2Sync[2]), .QTFCLK( ), .Q(maxFck2Sync[2]));
Q_FDP0UA U680 ( .D(maxFck2Sync[1]), .QTFCLK( ), .Q(maxFck2Sync[1]));
Q_FDP0UA U681 ( .D(maxFck2Sync[0]), .QTFCLK( ), .Q(maxFck2Sync[0]));
Q_FDP0UA U682 ( .D(maxGfifo2Sync[15]), .QTFCLK( ), .Q(maxGfifo2Sync[15]));
Q_FDP0UA U683 ( .D(maxGfifo2Sync[14]), .QTFCLK( ), .Q(maxGfifo2Sync[14]));
Q_FDP0UA U684 ( .D(maxGfifo2Sync[13]), .QTFCLK( ), .Q(maxGfifo2Sync[13]));
Q_FDP0UA U685 ( .D(maxGfifo2Sync[12]), .QTFCLK( ), .Q(maxGfifo2Sync[12]));
Q_FDP0UA U686 ( .D(maxGfifo2Sync[11]), .QTFCLK( ), .Q(maxGfifo2Sync[11]));
Q_FDP0UA U687 ( .D(maxGfifo2Sync[10]), .QTFCLK( ), .Q(maxGfifo2Sync[10]));
Q_FDP0UA U688 ( .D(maxGfifo2Sync[9]), .QTFCLK( ), .Q(maxGfifo2Sync[9]));
Q_FDP0UA U689 ( .D(maxGfifo2Sync[8]), .QTFCLK( ), .Q(maxGfifo2Sync[8]));
Q_FDP0UA U690 ( .D(maxGfifo2Sync[7]), .QTFCLK( ), .Q(maxGfifo2Sync[7]));
Q_FDP0UA U691 ( .D(maxGfifo2Sync[6]), .QTFCLK( ), .Q(maxGfifo2Sync[6]));
Q_FDP0UA U692 ( .D(maxGfifo2Sync[5]), .QTFCLK( ), .Q(maxGfifo2Sync[5]));
Q_FDP0UA U693 ( .D(maxGfifo2Sync[4]), .QTFCLK( ), .Q(maxGfifo2Sync[4]));
Q_FDP0UA U694 ( .D(maxGfifo2Sync[3]), .QTFCLK( ), .Q(maxGfifo2Sync[3]));
Q_FDP0UA U695 ( .D(maxGfifo2Sync[2]), .QTFCLK( ), .Q(maxGfifo2Sync[2]));
Q_FDP0UA U696 ( .D(maxGfifo2Sync[1]), .QTFCLK( ), .Q(maxGfifo2Sync[1]));
Q_FDP0UA U697 ( .D(maxGfifo2Sync[0]), .QTFCLK( ), .Q(maxGfifo2Sync[0]));
Q_NR02 U698 ( .A0(GFGBfullBw), .A1(GFGBfullBwD), .Z(n406));
Q_NR02 U699 ( .A0(GFLBfull), .A1(GFLBfullD), .Z(n404));
Q_AN02 U700 ( .A0(n406), .A1(n404), .Z(n403));
Q_INV U701 ( .A(evalOnC), .Z(n402));
Q_AN03 U702 ( .A0(GFbusy), .A1(n402), .A2(n403), .Z(n398));
Q_INV U703 ( .A(n404), .Z(n405));
Q_AN02 U704 ( .A0(n406), .A1(n405), .Z(n399));
Q_INV U705 ( .A(n406), .Z(n400));
Q_NR02 U706 ( .A0(holdEcm), .A1(holdEcmD), .Z(n407));
Q_INV U707 ( .A(n407), .Z(n401));
Q_XOR2 U708 ( .A0(n398), .A1(gfifoTBsyncCnt[0]), .Z(n408));
Q_FDP0UA U709 ( .D(n408), .QTFCLK( ), .Q(gfifoTBsyncCnt[0]));
Q_MX02 U710 ( .S(n398), .A0(gfifoTBsyncCnt[1]), .A1(n911), .Z(n409));
Q_FDP0UA U711 ( .D(n409), .QTFCLK( ), .Q(gfifoTBsyncCnt[1]));
Q_MX02 U712 ( .S(n398), .A0(gfifoTBsyncCnt[2]), .A1(n909), .Z(n410));
Q_FDP0UA U713 ( .D(n410), .QTFCLK( ), .Q(gfifoTBsyncCnt[2]));
Q_MX02 U714 ( .S(n398), .A0(gfifoTBsyncCnt[3]), .A1(n907), .Z(n411));
Q_FDP0UA U715 ( .D(n411), .QTFCLK( ), .Q(gfifoTBsyncCnt[3]));
Q_MX02 U716 ( .S(n398), .A0(gfifoTBsyncCnt[4]), .A1(n905), .Z(n412));
Q_FDP0UA U717 ( .D(n412), .QTFCLK( ), .Q(gfifoTBsyncCnt[4]));
Q_MX02 U718 ( .S(n398), .A0(gfifoTBsyncCnt[5]), .A1(n903), .Z(n413));
Q_FDP0UA U719 ( .D(n413), .QTFCLK( ), .Q(gfifoTBsyncCnt[5]));
Q_MX02 U720 ( .S(n398), .A0(gfifoTBsyncCnt[6]), .A1(n901), .Z(n414));
Q_FDP0UA U721 ( .D(n414), .QTFCLK( ), .Q(gfifoTBsyncCnt[6]));
Q_MX02 U722 ( .S(n398), .A0(gfifoTBsyncCnt[7]), .A1(n899), .Z(n415));
Q_FDP0UA U723 ( .D(n415), .QTFCLK( ), .Q(gfifoTBsyncCnt[7]));
Q_MX02 U724 ( .S(n398), .A0(gfifoTBsyncCnt[8]), .A1(n897), .Z(n416));
Q_FDP0UA U725 ( .D(n416), .QTFCLK( ), .Q(gfifoTBsyncCnt[8]));
Q_MX02 U726 ( .S(n398), .A0(gfifoTBsyncCnt[9]), .A1(n895), .Z(n417));
Q_FDP0UA U727 ( .D(n417), .QTFCLK( ), .Q(gfifoTBsyncCnt[9]));
Q_MX02 U728 ( .S(n398), .A0(gfifoTBsyncCnt[10]), .A1(n893), .Z(n418));
Q_FDP0UA U729 ( .D(n418), .QTFCLK( ), .Q(gfifoTBsyncCnt[10]));
Q_MX02 U730 ( .S(n398), .A0(gfifoTBsyncCnt[11]), .A1(n891), .Z(n419));
Q_FDP0UA U731 ( .D(n419), .QTFCLK( ), .Q(gfifoTBsyncCnt[11]));
Q_MX02 U732 ( .S(n398), .A0(gfifoTBsyncCnt[12]), .A1(n889), .Z(n420));
Q_FDP0UA U733 ( .D(n420), .QTFCLK( ), .Q(gfifoTBsyncCnt[12]));
Q_MX02 U734 ( .S(n398), .A0(gfifoTBsyncCnt[13]), .A1(n887), .Z(n421));
Q_FDP0UA U735 ( .D(n421), .QTFCLK( ), .Q(gfifoTBsyncCnt[13]));
Q_MX02 U736 ( .S(n398), .A0(gfifoTBsyncCnt[14]), .A1(n885), .Z(n422));
Q_FDP0UA U737 ( .D(n422), .QTFCLK( ), .Q(gfifoTBsyncCnt[14]));
Q_MX02 U738 ( .S(n398), .A0(gfifoTBsyncCnt[15]), .A1(n883), .Z(n423));
Q_FDP0UA U739 ( .D(n423), .QTFCLK( ), .Q(gfifoTBsyncCnt[15]));
Q_MX02 U740 ( .S(n398), .A0(gfifoTBsyncCnt[16]), .A1(n881), .Z(n424));
Q_FDP0UA U741 ( .D(n424), .QTFCLK( ), .Q(gfifoTBsyncCnt[16]));
Q_MX02 U742 ( .S(n398), .A0(gfifoTBsyncCnt[17]), .A1(n879), .Z(n425));
Q_FDP0UA U743 ( .D(n425), .QTFCLK( ), .Q(gfifoTBsyncCnt[17]));
Q_MX02 U744 ( .S(n398), .A0(gfifoTBsyncCnt[18]), .A1(n877), .Z(n426));
Q_FDP0UA U745 ( .D(n426), .QTFCLK( ), .Q(gfifoTBsyncCnt[18]));
Q_MX02 U746 ( .S(n398), .A0(gfifoTBsyncCnt[19]), .A1(n875), .Z(n427));
Q_FDP0UA U747 ( .D(n427), .QTFCLK( ), .Q(gfifoTBsyncCnt[19]));
Q_MX02 U748 ( .S(n398), .A0(gfifoTBsyncCnt[20]), .A1(n873), .Z(n428));
Q_FDP0UA U749 ( .D(n428), .QTFCLK( ), .Q(gfifoTBsyncCnt[20]));
Q_MX02 U750 ( .S(n398), .A0(gfifoTBsyncCnt[21]), .A1(n871), .Z(n429));
Q_FDP0UA U751 ( .D(n429), .QTFCLK( ), .Q(gfifoTBsyncCnt[21]));
Q_MX02 U752 ( .S(n398), .A0(gfifoTBsyncCnt[22]), .A1(n869), .Z(n430));
Q_FDP0UA U753 ( .D(n430), .QTFCLK( ), .Q(gfifoTBsyncCnt[22]));
Q_MX02 U754 ( .S(n398), .A0(gfifoTBsyncCnt[23]), .A1(n867), .Z(n431));
Q_FDP0UA U755 ( .D(n431), .QTFCLK( ), .Q(gfifoTBsyncCnt[23]));
Q_MX02 U756 ( .S(n398), .A0(gfifoTBsyncCnt[24]), .A1(n865), .Z(n432));
Q_FDP0UA U757 ( .D(n432), .QTFCLK( ), .Q(gfifoTBsyncCnt[24]));
Q_MX02 U758 ( .S(n398), .A0(gfifoTBsyncCnt[25]), .A1(n863), .Z(n433));
Q_FDP0UA U759 ( .D(n433), .QTFCLK( ), .Q(gfifoTBsyncCnt[25]));
Q_MX02 U760 ( .S(n398), .A0(gfifoTBsyncCnt[26]), .A1(n861), .Z(n434));
Q_FDP0UA U761 ( .D(n434), .QTFCLK( ), .Q(gfifoTBsyncCnt[26]));
Q_MX02 U762 ( .S(n398), .A0(gfifoTBsyncCnt[27]), .A1(n859), .Z(n435));
Q_FDP0UA U763 ( .D(n435), .QTFCLK( ), .Q(gfifoTBsyncCnt[27]));
Q_MX02 U764 ( .S(n398), .A0(gfifoTBsyncCnt[28]), .A1(n857), .Z(n436));
Q_FDP0UA U765 ( .D(n436), .QTFCLK( ), .Q(gfifoTBsyncCnt[28]));
Q_MX02 U766 ( .S(n398), .A0(gfifoTBsyncCnt[29]), .A1(n855), .Z(n437));
Q_FDP0UA U767 ( .D(n437), .QTFCLK( ), .Q(gfifoTBsyncCnt[29]));
Q_MX02 U768 ( .S(n398), .A0(gfifoTBsyncCnt[30]), .A1(n853), .Z(n438));
Q_FDP0UA U769 ( .D(n438), .QTFCLK( ), .Q(gfifoTBsyncCnt[30]));
Q_MX02 U770 ( .S(n398), .A0(gfifoTBsyncCnt[31]), .A1(n851), .Z(n439));
Q_FDP0UA U771 ( .D(n439), .QTFCLK( ), .Q(gfifoTBsyncCnt[31]));
Q_MX02 U772 ( .S(n398), .A0(gfifoTBsyncCnt[32]), .A1(n849), .Z(n440));
Q_FDP0UA U773 ( .D(n440), .QTFCLK( ), .Q(gfifoTBsyncCnt[32]));
Q_MX02 U774 ( .S(n398), .A0(gfifoTBsyncCnt[33]), .A1(n847), .Z(n441));
Q_FDP0UA U775 ( .D(n441), .QTFCLK( ), .Q(gfifoTBsyncCnt[33]));
Q_MX02 U776 ( .S(n398), .A0(gfifoTBsyncCnt[34]), .A1(n845), .Z(n442));
Q_FDP0UA U777 ( .D(n442), .QTFCLK( ), .Q(gfifoTBsyncCnt[34]));
Q_MX02 U778 ( .S(n398), .A0(gfifoTBsyncCnt[35]), .A1(n843), .Z(n443));
Q_FDP0UA U779 ( .D(n443), .QTFCLK( ), .Q(gfifoTBsyncCnt[35]));
Q_MX02 U780 ( .S(n398), .A0(gfifoTBsyncCnt[36]), .A1(n841), .Z(n444));
Q_FDP0UA U781 ( .D(n444), .QTFCLK( ), .Q(gfifoTBsyncCnt[36]));
Q_MX02 U782 ( .S(n398), .A0(gfifoTBsyncCnt[37]), .A1(n839), .Z(n445));
Q_FDP0UA U783 ( .D(n445), .QTFCLK( ), .Q(gfifoTBsyncCnt[37]));
Q_MX02 U784 ( .S(n398), .A0(gfifoTBsyncCnt[38]), .A1(n837), .Z(n446));
Q_FDP0UA U785 ( .D(n446), .QTFCLK( ), .Q(gfifoTBsyncCnt[38]));
Q_MX02 U786 ( .S(n398), .A0(gfifoTBsyncCnt[39]), .A1(n835), .Z(n447));
Q_FDP0UA U787 ( .D(n447), .QTFCLK( ), .Q(gfifoTBsyncCnt[39]));
Q_MX02 U788 ( .S(n398), .A0(gfifoTBsyncCnt[40]), .A1(n833), .Z(n448));
Q_FDP0UA U789 ( .D(n448), .QTFCLK( ), .Q(gfifoTBsyncCnt[40]));
Q_MX02 U790 ( .S(n398), .A0(gfifoTBsyncCnt[41]), .A1(n831), .Z(n449));
Q_FDP0UA U791 ( .D(n449), .QTFCLK( ), .Q(gfifoTBsyncCnt[41]));
Q_MX02 U792 ( .S(n398), .A0(gfifoTBsyncCnt[42]), .A1(n829), .Z(n450));
Q_FDP0UA U793 ( .D(n450), .QTFCLK( ), .Q(gfifoTBsyncCnt[42]));
Q_MX02 U794 ( .S(n398), .A0(gfifoTBsyncCnt[43]), .A1(n827), .Z(n451));
Q_FDP0UA U795 ( .D(n451), .QTFCLK( ), .Q(gfifoTBsyncCnt[43]));
Q_MX02 U796 ( .S(n398), .A0(gfifoTBsyncCnt[44]), .A1(n825), .Z(n452));
Q_FDP0UA U797 ( .D(n452), .QTFCLK( ), .Q(gfifoTBsyncCnt[44]));
Q_MX02 U798 ( .S(n398), .A0(gfifoTBsyncCnt[45]), .A1(n823), .Z(n453));
Q_FDP0UA U799 ( .D(n453), .QTFCLK( ), .Q(gfifoTBsyncCnt[45]));
Q_MX02 U800 ( .S(n398), .A0(gfifoTBsyncCnt[46]), .A1(n821), .Z(n454));
Q_FDP0UA U801 ( .D(n454), .QTFCLK( ), .Q(gfifoTBsyncCnt[46]));
Q_MX02 U802 ( .S(n398), .A0(gfifoTBsyncCnt[47]), .A1(n819), .Z(n455));
Q_FDP0UA U803 ( .D(n455), .QTFCLK( ), .Q(gfifoTBsyncCnt[47]));
Q_MX02 U804 ( .S(n398), .A0(gfifoTBsyncCnt[48]), .A1(n817), .Z(n456));
Q_FDP0UA U805 ( .D(n456), .QTFCLK( ), .Q(gfifoTBsyncCnt[48]));
Q_MX02 U806 ( .S(n398), .A0(gfifoTBsyncCnt[49]), .A1(n815), .Z(n457));
Q_FDP0UA U807 ( .D(n457), .QTFCLK( ), .Q(gfifoTBsyncCnt[49]));
Q_MX02 U808 ( .S(n398), .A0(gfifoTBsyncCnt[50]), .A1(n813), .Z(n458));
Q_FDP0UA U809 ( .D(n458), .QTFCLK( ), .Q(gfifoTBsyncCnt[50]));
Q_MX02 U810 ( .S(n398), .A0(gfifoTBsyncCnt[51]), .A1(n811), .Z(n459));
Q_FDP0UA U811 ( .D(n459), .QTFCLK( ), .Q(gfifoTBsyncCnt[51]));
Q_MX02 U812 ( .S(n398), .A0(gfifoTBsyncCnt[52]), .A1(n809), .Z(n460));
Q_FDP0UA U813 ( .D(n460), .QTFCLK( ), .Q(gfifoTBsyncCnt[52]));
Q_MX02 U814 ( .S(n398), .A0(gfifoTBsyncCnt[53]), .A1(n807), .Z(n461));
Q_FDP0UA U815 ( .D(n461), .QTFCLK( ), .Q(gfifoTBsyncCnt[53]));
Q_MX02 U816 ( .S(n398), .A0(gfifoTBsyncCnt[54]), .A1(n805), .Z(n462));
Q_FDP0UA U817 ( .D(n462), .QTFCLK( ), .Q(gfifoTBsyncCnt[54]));
Q_MX02 U818 ( .S(n398), .A0(gfifoTBsyncCnt[55]), .A1(n803), .Z(n463));
Q_FDP0UA U819 ( .D(n463), .QTFCLK( ), .Q(gfifoTBsyncCnt[55]));
Q_MX02 U820 ( .S(n398), .A0(gfifoTBsyncCnt[56]), .A1(n801), .Z(n464));
Q_FDP0UA U821 ( .D(n464), .QTFCLK( ), .Q(gfifoTBsyncCnt[56]));
Q_MX02 U822 ( .S(n398), .A0(gfifoTBsyncCnt[57]), .A1(n799), .Z(n465));
Q_FDP0UA U823 ( .D(n465), .QTFCLK( ), .Q(gfifoTBsyncCnt[57]));
Q_MX02 U824 ( .S(n398), .A0(gfifoTBsyncCnt[58]), .A1(n797), .Z(n466));
Q_FDP0UA U825 ( .D(n466), .QTFCLK( ), .Q(gfifoTBsyncCnt[58]));
Q_MX02 U826 ( .S(n398), .A0(gfifoTBsyncCnt[59]), .A1(n795), .Z(n467));
Q_FDP0UA U827 ( .D(n467), .QTFCLK( ), .Q(gfifoTBsyncCnt[59]));
Q_MX02 U828 ( .S(n398), .A0(gfifoTBsyncCnt[60]), .A1(n793), .Z(n468));
Q_FDP0UA U829 ( .D(n468), .QTFCLK( ), .Q(gfifoTBsyncCnt[60]));
Q_MX02 U830 ( .S(n398), .A0(gfifoTBsyncCnt[61]), .A1(n791), .Z(n469));
Q_FDP0UA U831 ( .D(n469), .QTFCLK( ), .Q(gfifoTBsyncCnt[61]));
Q_MX02 U832 ( .S(n398), .A0(gfifoTBsyncCnt[62]), .A1(n789), .Z(n470));
Q_FDP0UA U833 ( .D(n470), .QTFCLK( ), .Q(gfifoTBsyncCnt[62]));
Q_FDP0UA U834 ( .D(n471), .QTFCLK( ), .Q(gfifoTBsyncCnt[63]));
Q_XOR2 U835 ( .A0(n399), .A1(gfifoLBfullCnt[0]), .Z(n472));
Q_FDP0UA U836 ( .D(n472), .QTFCLK( ), .Q(gfifoLBfullCnt[0]));
Q_MX02 U837 ( .S(n399), .A0(gfifoLBfullCnt[1]), .A1(n1035), .Z(n473));
Q_FDP0UA U838 ( .D(n473), .QTFCLK( ), .Q(gfifoLBfullCnt[1]));
Q_MX02 U839 ( .S(n399), .A0(gfifoLBfullCnt[2]), .A1(n1033), .Z(n474));
Q_FDP0UA U840 ( .D(n474), .QTFCLK( ), .Q(gfifoLBfullCnt[2]));
Q_MX02 U841 ( .S(n399), .A0(gfifoLBfullCnt[3]), .A1(n1031), .Z(n475));
Q_FDP0UA U842 ( .D(n475), .QTFCLK( ), .Q(gfifoLBfullCnt[3]));
Q_MX02 U843 ( .S(n399), .A0(gfifoLBfullCnt[4]), .A1(n1029), .Z(n476));
Q_FDP0UA U844 ( .D(n476), .QTFCLK( ), .Q(gfifoLBfullCnt[4]));
Q_MX02 U845 ( .S(n399), .A0(gfifoLBfullCnt[5]), .A1(n1027), .Z(n477));
Q_FDP0UA U846 ( .D(n477), .QTFCLK( ), .Q(gfifoLBfullCnt[5]));
Q_MX02 U847 ( .S(n399), .A0(gfifoLBfullCnt[6]), .A1(n1025), .Z(n478));
Q_FDP0UA U848 ( .D(n478), .QTFCLK( ), .Q(gfifoLBfullCnt[6]));
Q_MX02 U849 ( .S(n399), .A0(gfifoLBfullCnt[7]), .A1(n1023), .Z(n479));
Q_FDP0UA U850 ( .D(n479), .QTFCLK( ), .Q(gfifoLBfullCnt[7]));
Q_MX02 U851 ( .S(n399), .A0(gfifoLBfullCnt[8]), .A1(n1021), .Z(n480));
Q_FDP0UA U852 ( .D(n480), .QTFCLK( ), .Q(gfifoLBfullCnt[8]));
Q_MX02 U853 ( .S(n399), .A0(gfifoLBfullCnt[9]), .A1(n1019), .Z(n481));
Q_FDP0UA U854 ( .D(n481), .QTFCLK( ), .Q(gfifoLBfullCnt[9]));
Q_MX02 U855 ( .S(n399), .A0(gfifoLBfullCnt[10]), .A1(n1017), .Z(n482));
Q_FDP0UA U856 ( .D(n482), .QTFCLK( ), .Q(gfifoLBfullCnt[10]));
Q_MX02 U857 ( .S(n399), .A0(gfifoLBfullCnt[11]), .A1(n1015), .Z(n483));
Q_FDP0UA U858 ( .D(n483), .QTFCLK( ), .Q(gfifoLBfullCnt[11]));
Q_MX02 U859 ( .S(n399), .A0(gfifoLBfullCnt[12]), .A1(n1013), .Z(n484));
Q_FDP0UA U860 ( .D(n484), .QTFCLK( ), .Q(gfifoLBfullCnt[12]));
Q_MX02 U861 ( .S(n399), .A0(gfifoLBfullCnt[13]), .A1(n1011), .Z(n485));
Q_FDP0UA U862 ( .D(n485), .QTFCLK( ), .Q(gfifoLBfullCnt[13]));
Q_MX02 U863 ( .S(n399), .A0(gfifoLBfullCnt[14]), .A1(n1009), .Z(n486));
Q_FDP0UA U864 ( .D(n486), .QTFCLK( ), .Q(gfifoLBfullCnt[14]));
Q_MX02 U865 ( .S(n399), .A0(gfifoLBfullCnt[15]), .A1(n1007), .Z(n487));
Q_FDP0UA U866 ( .D(n487), .QTFCLK( ), .Q(gfifoLBfullCnt[15]));
Q_MX02 U867 ( .S(n399), .A0(gfifoLBfullCnt[16]), .A1(n1005), .Z(n488));
Q_FDP0UA U868 ( .D(n488), .QTFCLK( ), .Q(gfifoLBfullCnt[16]));
Q_MX02 U869 ( .S(n399), .A0(gfifoLBfullCnt[17]), .A1(n1003), .Z(n489));
Q_FDP0UA U870 ( .D(n489), .QTFCLK( ), .Q(gfifoLBfullCnt[17]));
Q_MX02 U871 ( .S(n399), .A0(gfifoLBfullCnt[18]), .A1(n1001), .Z(n490));
Q_FDP0UA U872 ( .D(n490), .QTFCLK( ), .Q(gfifoLBfullCnt[18]));
Q_MX02 U873 ( .S(n399), .A0(gfifoLBfullCnt[19]), .A1(n999), .Z(n491));
Q_FDP0UA U874 ( .D(n491), .QTFCLK( ), .Q(gfifoLBfullCnt[19]));
Q_MX02 U875 ( .S(n399), .A0(gfifoLBfullCnt[20]), .A1(n997), .Z(n492));
Q_FDP0UA U876 ( .D(n492), .QTFCLK( ), .Q(gfifoLBfullCnt[20]));
Q_MX02 U877 ( .S(n399), .A0(gfifoLBfullCnt[21]), .A1(n995), .Z(n493));
Q_FDP0UA U878 ( .D(n493), .QTFCLK( ), .Q(gfifoLBfullCnt[21]));
Q_MX02 U879 ( .S(n399), .A0(gfifoLBfullCnt[22]), .A1(n993), .Z(n494));
Q_FDP0UA U880 ( .D(n494), .QTFCLK( ), .Q(gfifoLBfullCnt[22]));
Q_MX02 U881 ( .S(n399), .A0(gfifoLBfullCnt[23]), .A1(n991), .Z(n495));
Q_FDP0UA U882 ( .D(n495), .QTFCLK( ), .Q(gfifoLBfullCnt[23]));
Q_MX02 U883 ( .S(n399), .A0(gfifoLBfullCnt[24]), .A1(n989), .Z(n496));
Q_FDP0UA U884 ( .D(n496), .QTFCLK( ), .Q(gfifoLBfullCnt[24]));
Q_MX02 U885 ( .S(n399), .A0(gfifoLBfullCnt[25]), .A1(n987), .Z(n497));
Q_FDP0UA U886 ( .D(n497), .QTFCLK( ), .Q(gfifoLBfullCnt[25]));
Q_MX02 U887 ( .S(n399), .A0(gfifoLBfullCnt[26]), .A1(n985), .Z(n498));
Q_FDP0UA U888 ( .D(n498), .QTFCLK( ), .Q(gfifoLBfullCnt[26]));
Q_MX02 U889 ( .S(n399), .A0(gfifoLBfullCnt[27]), .A1(n983), .Z(n499));
Q_FDP0UA U890 ( .D(n499), .QTFCLK( ), .Q(gfifoLBfullCnt[27]));
Q_MX02 U891 ( .S(n399), .A0(gfifoLBfullCnt[28]), .A1(n981), .Z(n500));
Q_FDP0UA U892 ( .D(n500), .QTFCLK( ), .Q(gfifoLBfullCnt[28]));
Q_MX02 U893 ( .S(n399), .A0(gfifoLBfullCnt[29]), .A1(n979), .Z(n501));
Q_FDP0UA U894 ( .D(n501), .QTFCLK( ), .Q(gfifoLBfullCnt[29]));
Q_MX02 U895 ( .S(n399), .A0(gfifoLBfullCnt[30]), .A1(n977), .Z(n502));
Q_FDP0UA U896 ( .D(n502), .QTFCLK( ), .Q(gfifoLBfullCnt[30]));
Q_MX02 U897 ( .S(n399), .A0(gfifoLBfullCnt[31]), .A1(n975), .Z(n503));
Q_FDP0UA U898 ( .D(n503), .QTFCLK( ), .Q(gfifoLBfullCnt[31]));
Q_MX02 U899 ( .S(n399), .A0(gfifoLBfullCnt[32]), .A1(n973), .Z(n504));
Q_FDP0UA U900 ( .D(n504), .QTFCLK( ), .Q(gfifoLBfullCnt[32]));
Q_MX02 U901 ( .S(n399), .A0(gfifoLBfullCnt[33]), .A1(n971), .Z(n505));
Q_FDP0UA U902 ( .D(n505), .QTFCLK( ), .Q(gfifoLBfullCnt[33]));
Q_MX02 U903 ( .S(n399), .A0(gfifoLBfullCnt[34]), .A1(n969), .Z(n506));
Q_FDP0UA U904 ( .D(n506), .QTFCLK( ), .Q(gfifoLBfullCnt[34]));
Q_MX02 U905 ( .S(n399), .A0(gfifoLBfullCnt[35]), .A1(n967), .Z(n507));
Q_FDP0UA U906 ( .D(n507), .QTFCLK( ), .Q(gfifoLBfullCnt[35]));
Q_MX02 U907 ( .S(n399), .A0(gfifoLBfullCnt[36]), .A1(n965), .Z(n508));
Q_FDP0UA U908 ( .D(n508), .QTFCLK( ), .Q(gfifoLBfullCnt[36]));
Q_MX02 U909 ( .S(n399), .A0(gfifoLBfullCnt[37]), .A1(n963), .Z(n509));
Q_FDP0UA U910 ( .D(n509), .QTFCLK( ), .Q(gfifoLBfullCnt[37]));
Q_MX02 U911 ( .S(n399), .A0(gfifoLBfullCnt[38]), .A1(n961), .Z(n510));
Q_FDP0UA U912 ( .D(n510), .QTFCLK( ), .Q(gfifoLBfullCnt[38]));
Q_MX02 U913 ( .S(n399), .A0(gfifoLBfullCnt[39]), .A1(n959), .Z(n511));
Q_FDP0UA U914 ( .D(n511), .QTFCLK( ), .Q(gfifoLBfullCnt[39]));
Q_MX02 U915 ( .S(n399), .A0(gfifoLBfullCnt[40]), .A1(n957), .Z(n512));
Q_FDP0UA U916 ( .D(n512), .QTFCLK( ), .Q(gfifoLBfullCnt[40]));
Q_MX02 U917 ( .S(n399), .A0(gfifoLBfullCnt[41]), .A1(n955), .Z(n513));
Q_FDP0UA U918 ( .D(n513), .QTFCLK( ), .Q(gfifoLBfullCnt[41]));
Q_MX02 U919 ( .S(n399), .A0(gfifoLBfullCnt[42]), .A1(n953), .Z(n514));
Q_FDP0UA U920 ( .D(n514), .QTFCLK( ), .Q(gfifoLBfullCnt[42]));
Q_MX02 U921 ( .S(n399), .A0(gfifoLBfullCnt[43]), .A1(n951), .Z(n515));
Q_FDP0UA U922 ( .D(n515), .QTFCLK( ), .Q(gfifoLBfullCnt[43]));
Q_MX02 U923 ( .S(n399), .A0(gfifoLBfullCnt[44]), .A1(n949), .Z(n516));
Q_FDP0UA U924 ( .D(n516), .QTFCLK( ), .Q(gfifoLBfullCnt[44]));
Q_MX02 U925 ( .S(n399), .A0(gfifoLBfullCnt[45]), .A1(n947), .Z(n517));
Q_FDP0UA U926 ( .D(n517), .QTFCLK( ), .Q(gfifoLBfullCnt[45]));
Q_MX02 U927 ( .S(n399), .A0(gfifoLBfullCnt[46]), .A1(n945), .Z(n518));
Q_FDP0UA U928 ( .D(n518), .QTFCLK( ), .Q(gfifoLBfullCnt[46]));
Q_MX02 U929 ( .S(n399), .A0(gfifoLBfullCnt[47]), .A1(n943), .Z(n519));
Q_FDP0UA U930 ( .D(n519), .QTFCLK( ), .Q(gfifoLBfullCnt[47]));
Q_MX02 U931 ( .S(n399), .A0(gfifoLBfullCnt[48]), .A1(n941), .Z(n520));
Q_FDP0UA U932 ( .D(n520), .QTFCLK( ), .Q(gfifoLBfullCnt[48]));
Q_MX02 U933 ( .S(n399), .A0(gfifoLBfullCnt[49]), .A1(n939), .Z(n521));
Q_FDP0UA U934 ( .D(n521), .QTFCLK( ), .Q(gfifoLBfullCnt[49]));
Q_MX02 U935 ( .S(n399), .A0(gfifoLBfullCnt[50]), .A1(n937), .Z(n522));
Q_FDP0UA U936 ( .D(n522), .QTFCLK( ), .Q(gfifoLBfullCnt[50]));
Q_MX02 U937 ( .S(n399), .A0(gfifoLBfullCnt[51]), .A1(n935), .Z(n523));
Q_FDP0UA U938 ( .D(n523), .QTFCLK( ), .Q(gfifoLBfullCnt[51]));
Q_MX02 U939 ( .S(n399), .A0(gfifoLBfullCnt[52]), .A1(n933), .Z(n524));
Q_FDP0UA U940 ( .D(n524), .QTFCLK( ), .Q(gfifoLBfullCnt[52]));
Q_MX02 U941 ( .S(n399), .A0(gfifoLBfullCnt[53]), .A1(n931), .Z(n525));
Q_FDP0UA U942 ( .D(n525), .QTFCLK( ), .Q(gfifoLBfullCnt[53]));
Q_MX02 U943 ( .S(n399), .A0(gfifoLBfullCnt[54]), .A1(n929), .Z(n526));
Q_FDP0UA U944 ( .D(n526), .QTFCLK( ), .Q(gfifoLBfullCnt[54]));
Q_MX02 U945 ( .S(n399), .A0(gfifoLBfullCnt[55]), .A1(n927), .Z(n527));
Q_FDP0UA U946 ( .D(n527), .QTFCLK( ), .Q(gfifoLBfullCnt[55]));
Q_MX02 U947 ( .S(n399), .A0(gfifoLBfullCnt[56]), .A1(n925), .Z(n528));
Q_FDP0UA U948 ( .D(n528), .QTFCLK( ), .Q(gfifoLBfullCnt[56]));
Q_MX02 U949 ( .S(n399), .A0(gfifoLBfullCnt[57]), .A1(n923), .Z(n529));
Q_FDP0UA U950 ( .D(n529), .QTFCLK( ), .Q(gfifoLBfullCnt[57]));
Q_MX02 U951 ( .S(n399), .A0(gfifoLBfullCnt[58]), .A1(n921), .Z(n530));
Q_FDP0UA U952 ( .D(n530), .QTFCLK( ), .Q(gfifoLBfullCnt[58]));
Q_MX02 U953 ( .S(n399), .A0(gfifoLBfullCnt[59]), .A1(n919), .Z(n531));
Q_FDP0UA U954 ( .D(n531), .QTFCLK( ), .Q(gfifoLBfullCnt[59]));
Q_MX02 U955 ( .S(n399), .A0(gfifoLBfullCnt[60]), .A1(n917), .Z(n532));
Q_FDP0UA U956 ( .D(n532), .QTFCLK( ), .Q(gfifoLBfullCnt[60]));
Q_MX02 U957 ( .S(n399), .A0(gfifoLBfullCnt[61]), .A1(n915), .Z(n533));
Q_FDP0UA U958 ( .D(n533), .QTFCLK( ), .Q(gfifoLBfullCnt[61]));
Q_MX02 U959 ( .S(n399), .A0(gfifoLBfullCnt[62]), .A1(n913), .Z(n534));
Q_FDP0UA U960 ( .D(n534), .QTFCLK( ), .Q(gfifoLBfullCnt[62]));
Q_FDP0UA U961 ( .D(n535), .QTFCLK( ), .Q(gfifoLBfullCnt[63]));
Q_XOR2 U962 ( .A0(n400), .A1(gfifoGBfullCnt[0]), .Z(n536));
Q_FDP0UA U963 ( .D(n536), .QTFCLK( ), .Q(gfifoGBfullCnt[0]));
Q_MX02 U964 ( .S(n406), .A0(n1159), .A1(gfifoGBfullCnt[1]), .Z(n537));
Q_FDP0UA U965 ( .D(n537), .QTFCLK( ), .Q(gfifoGBfullCnt[1]));
Q_MX02 U966 ( .S(n406), .A0(n1157), .A1(gfifoGBfullCnt[2]), .Z(n538));
Q_FDP0UA U967 ( .D(n538), .QTFCLK( ), .Q(gfifoGBfullCnt[2]));
Q_MX02 U968 ( .S(n406), .A0(n1155), .A1(gfifoGBfullCnt[3]), .Z(n539));
Q_FDP0UA U969 ( .D(n539), .QTFCLK( ), .Q(gfifoGBfullCnt[3]));
Q_MX02 U970 ( .S(n406), .A0(n1153), .A1(gfifoGBfullCnt[4]), .Z(n540));
Q_FDP0UA U971 ( .D(n540), .QTFCLK( ), .Q(gfifoGBfullCnt[4]));
Q_MX02 U972 ( .S(n406), .A0(n1151), .A1(gfifoGBfullCnt[5]), .Z(n541));
Q_FDP0UA U973 ( .D(n541), .QTFCLK( ), .Q(gfifoGBfullCnt[5]));
Q_MX02 U974 ( .S(n406), .A0(n1149), .A1(gfifoGBfullCnt[6]), .Z(n542));
Q_FDP0UA U975 ( .D(n542), .QTFCLK( ), .Q(gfifoGBfullCnt[6]));
Q_MX02 U976 ( .S(n406), .A0(n1147), .A1(gfifoGBfullCnt[7]), .Z(n543));
Q_FDP0UA U977 ( .D(n543), .QTFCLK( ), .Q(gfifoGBfullCnt[7]));
Q_MX02 U978 ( .S(n406), .A0(n1145), .A1(gfifoGBfullCnt[8]), .Z(n544));
Q_FDP0UA U979 ( .D(n544), .QTFCLK( ), .Q(gfifoGBfullCnt[8]));
Q_MX02 U980 ( .S(n406), .A0(n1143), .A1(gfifoGBfullCnt[9]), .Z(n545));
Q_FDP0UA U981 ( .D(n545), .QTFCLK( ), .Q(gfifoGBfullCnt[9]));
Q_MX02 U982 ( .S(n406), .A0(n1141), .A1(gfifoGBfullCnt[10]), .Z(n546));
Q_FDP0UA U983 ( .D(n546), .QTFCLK( ), .Q(gfifoGBfullCnt[10]));
Q_MX02 U984 ( .S(n406), .A0(n1139), .A1(gfifoGBfullCnt[11]), .Z(n547));
Q_FDP0UA U985 ( .D(n547), .QTFCLK( ), .Q(gfifoGBfullCnt[11]));
Q_MX02 U986 ( .S(n406), .A0(n1137), .A1(gfifoGBfullCnt[12]), .Z(n548));
Q_FDP0UA U987 ( .D(n548), .QTFCLK( ), .Q(gfifoGBfullCnt[12]));
Q_MX02 U988 ( .S(n406), .A0(n1135), .A1(gfifoGBfullCnt[13]), .Z(n549));
Q_FDP0UA U989 ( .D(n549), .QTFCLK( ), .Q(gfifoGBfullCnt[13]));
Q_MX02 U990 ( .S(n406), .A0(n1133), .A1(gfifoGBfullCnt[14]), .Z(n550));
Q_FDP0UA U991 ( .D(n550), .QTFCLK( ), .Q(gfifoGBfullCnt[14]));
Q_MX02 U992 ( .S(n406), .A0(n1131), .A1(gfifoGBfullCnt[15]), .Z(n551));
Q_FDP0UA U993 ( .D(n551), .QTFCLK( ), .Q(gfifoGBfullCnt[15]));
Q_MX02 U994 ( .S(n406), .A0(n1129), .A1(gfifoGBfullCnt[16]), .Z(n552));
Q_FDP0UA U995 ( .D(n552), .QTFCLK( ), .Q(gfifoGBfullCnt[16]));
Q_MX02 U996 ( .S(n406), .A0(n1127), .A1(gfifoGBfullCnt[17]), .Z(n553));
Q_FDP0UA U997 ( .D(n553), .QTFCLK( ), .Q(gfifoGBfullCnt[17]));
Q_MX02 U998 ( .S(n406), .A0(n1125), .A1(gfifoGBfullCnt[18]), .Z(n554));
Q_FDP0UA U999 ( .D(n554), .QTFCLK( ), .Q(gfifoGBfullCnt[18]));
Q_MX02 U1000 ( .S(n406), .A0(n1123), .A1(gfifoGBfullCnt[19]), .Z(n555));
Q_FDP0UA U1001 ( .D(n555), .QTFCLK( ), .Q(gfifoGBfullCnt[19]));
Q_MX02 U1002 ( .S(n406), .A0(n1121), .A1(gfifoGBfullCnt[20]), .Z(n556));
Q_FDP0UA U1003 ( .D(n556), .QTFCLK( ), .Q(gfifoGBfullCnt[20]));
Q_MX02 U1004 ( .S(n406), .A0(n1119), .A1(gfifoGBfullCnt[21]), .Z(n557));
Q_FDP0UA U1005 ( .D(n557), .QTFCLK( ), .Q(gfifoGBfullCnt[21]));
Q_MX02 U1006 ( .S(n406), .A0(n1117), .A1(gfifoGBfullCnt[22]), .Z(n558));
Q_FDP0UA U1007 ( .D(n558), .QTFCLK( ), .Q(gfifoGBfullCnt[22]));
Q_MX02 U1008 ( .S(n406), .A0(n1115), .A1(gfifoGBfullCnt[23]), .Z(n559));
Q_FDP0UA U1009 ( .D(n559), .QTFCLK( ), .Q(gfifoGBfullCnt[23]));
Q_MX02 U1010 ( .S(n406), .A0(n1113), .A1(gfifoGBfullCnt[24]), .Z(n560));
Q_FDP0UA U1011 ( .D(n560), .QTFCLK( ), .Q(gfifoGBfullCnt[24]));
Q_MX02 U1012 ( .S(n406), .A0(n1111), .A1(gfifoGBfullCnt[25]), .Z(n561));
Q_FDP0UA U1013 ( .D(n561), .QTFCLK( ), .Q(gfifoGBfullCnt[25]));
Q_MX02 U1014 ( .S(n406), .A0(n1109), .A1(gfifoGBfullCnt[26]), .Z(n562));
Q_FDP0UA U1015 ( .D(n562), .QTFCLK( ), .Q(gfifoGBfullCnt[26]));
Q_MX02 U1016 ( .S(n406), .A0(n1107), .A1(gfifoGBfullCnt[27]), .Z(n563));
Q_FDP0UA U1017 ( .D(n563), .QTFCLK( ), .Q(gfifoGBfullCnt[27]));
Q_MX02 U1018 ( .S(n406), .A0(n1105), .A1(gfifoGBfullCnt[28]), .Z(n564));
Q_FDP0UA U1019 ( .D(n564), .QTFCLK( ), .Q(gfifoGBfullCnt[28]));
Q_MX02 U1020 ( .S(n406), .A0(n1103), .A1(gfifoGBfullCnt[29]), .Z(n565));
Q_FDP0UA U1021 ( .D(n565), .QTFCLK( ), .Q(gfifoGBfullCnt[29]));
Q_MX02 U1022 ( .S(n406), .A0(n1101), .A1(gfifoGBfullCnt[30]), .Z(n566));
Q_FDP0UA U1023 ( .D(n566), .QTFCLK( ), .Q(gfifoGBfullCnt[30]));
Q_MX02 U1024 ( .S(n406), .A0(n1099), .A1(gfifoGBfullCnt[31]), .Z(n567));
Q_FDP0UA U1025 ( .D(n567), .QTFCLK( ), .Q(gfifoGBfullCnt[31]));
Q_MX02 U1026 ( .S(n406), .A0(n1097), .A1(gfifoGBfullCnt[32]), .Z(n568));
Q_FDP0UA U1027 ( .D(n568), .QTFCLK( ), .Q(gfifoGBfullCnt[32]));
Q_MX02 U1028 ( .S(n406), .A0(n1095), .A1(gfifoGBfullCnt[33]), .Z(n569));
Q_FDP0UA U1029 ( .D(n569), .QTFCLK( ), .Q(gfifoGBfullCnt[33]));
Q_MX02 U1030 ( .S(n406), .A0(n1093), .A1(gfifoGBfullCnt[34]), .Z(n570));
Q_FDP0UA U1031 ( .D(n570), .QTFCLK( ), .Q(gfifoGBfullCnt[34]));
Q_MX02 U1032 ( .S(n406), .A0(n1091), .A1(gfifoGBfullCnt[35]), .Z(n571));
Q_FDP0UA U1033 ( .D(n571), .QTFCLK( ), .Q(gfifoGBfullCnt[35]));
Q_MX02 U1034 ( .S(n406), .A0(n1089), .A1(gfifoGBfullCnt[36]), .Z(n572));
Q_FDP0UA U1035 ( .D(n572), .QTFCLK( ), .Q(gfifoGBfullCnt[36]));
Q_MX02 U1036 ( .S(n406), .A0(n1087), .A1(gfifoGBfullCnt[37]), .Z(n573));
Q_FDP0UA U1037 ( .D(n573), .QTFCLK( ), .Q(gfifoGBfullCnt[37]));
Q_MX02 U1038 ( .S(n406), .A0(n1085), .A1(gfifoGBfullCnt[38]), .Z(n574));
Q_FDP0UA U1039 ( .D(n574), .QTFCLK( ), .Q(gfifoGBfullCnt[38]));
Q_MX02 U1040 ( .S(n406), .A0(n1083), .A1(gfifoGBfullCnt[39]), .Z(n575));
Q_FDP0UA U1041 ( .D(n575), .QTFCLK( ), .Q(gfifoGBfullCnt[39]));
Q_MX02 U1042 ( .S(n406), .A0(n1081), .A1(gfifoGBfullCnt[40]), .Z(n576));
Q_FDP0UA U1043 ( .D(n576), .QTFCLK( ), .Q(gfifoGBfullCnt[40]));
Q_MX02 U1044 ( .S(n406), .A0(n1079), .A1(gfifoGBfullCnt[41]), .Z(n577));
Q_FDP0UA U1045 ( .D(n577), .QTFCLK( ), .Q(gfifoGBfullCnt[41]));
Q_MX02 U1046 ( .S(n406), .A0(n1077), .A1(gfifoGBfullCnt[42]), .Z(n578));
Q_FDP0UA U1047 ( .D(n578), .QTFCLK( ), .Q(gfifoGBfullCnt[42]));
Q_MX02 U1048 ( .S(n406), .A0(n1075), .A1(gfifoGBfullCnt[43]), .Z(n579));
Q_FDP0UA U1049 ( .D(n579), .QTFCLK( ), .Q(gfifoGBfullCnt[43]));
Q_MX02 U1050 ( .S(n406), .A0(n1073), .A1(gfifoGBfullCnt[44]), .Z(n580));
Q_FDP0UA U1051 ( .D(n580), .QTFCLK( ), .Q(gfifoGBfullCnt[44]));
Q_MX02 U1052 ( .S(n406), .A0(n1071), .A1(gfifoGBfullCnt[45]), .Z(n581));
Q_FDP0UA U1053 ( .D(n581), .QTFCLK( ), .Q(gfifoGBfullCnt[45]));
Q_MX02 U1054 ( .S(n406), .A0(n1069), .A1(gfifoGBfullCnt[46]), .Z(n582));
Q_FDP0UA U1055 ( .D(n582), .QTFCLK( ), .Q(gfifoGBfullCnt[46]));
Q_MX02 U1056 ( .S(n406), .A0(n1067), .A1(gfifoGBfullCnt[47]), .Z(n583));
Q_FDP0UA U1057 ( .D(n583), .QTFCLK( ), .Q(gfifoGBfullCnt[47]));
Q_MX02 U1058 ( .S(n406), .A0(n1065), .A1(gfifoGBfullCnt[48]), .Z(n584));
Q_FDP0UA U1059 ( .D(n584), .QTFCLK( ), .Q(gfifoGBfullCnt[48]));
Q_MX02 U1060 ( .S(n406), .A0(n1063), .A1(gfifoGBfullCnt[49]), .Z(n585));
Q_FDP0UA U1061 ( .D(n585), .QTFCLK( ), .Q(gfifoGBfullCnt[49]));
Q_MX02 U1062 ( .S(n406), .A0(n1061), .A1(gfifoGBfullCnt[50]), .Z(n586));
Q_FDP0UA U1063 ( .D(n586), .QTFCLK( ), .Q(gfifoGBfullCnt[50]));
Q_MX02 U1064 ( .S(n406), .A0(n1059), .A1(gfifoGBfullCnt[51]), .Z(n587));
Q_FDP0UA U1065 ( .D(n587), .QTFCLK( ), .Q(gfifoGBfullCnt[51]));
Q_MX02 U1066 ( .S(n406), .A0(n1057), .A1(gfifoGBfullCnt[52]), .Z(n588));
Q_FDP0UA U1067 ( .D(n588), .QTFCLK( ), .Q(gfifoGBfullCnt[52]));
Q_MX02 U1068 ( .S(n406), .A0(n1055), .A1(gfifoGBfullCnt[53]), .Z(n589));
Q_FDP0UA U1069 ( .D(n589), .QTFCLK( ), .Q(gfifoGBfullCnt[53]));
Q_MX02 U1070 ( .S(n406), .A0(n1053), .A1(gfifoGBfullCnt[54]), .Z(n590));
Q_FDP0UA U1071 ( .D(n590), .QTFCLK( ), .Q(gfifoGBfullCnt[54]));
Q_MX02 U1072 ( .S(n406), .A0(n1051), .A1(gfifoGBfullCnt[55]), .Z(n591));
Q_FDP0UA U1073 ( .D(n591), .QTFCLK( ), .Q(gfifoGBfullCnt[55]));
Q_MX02 U1074 ( .S(n406), .A0(n1049), .A1(gfifoGBfullCnt[56]), .Z(n592));
Q_FDP0UA U1075 ( .D(n592), .QTFCLK( ), .Q(gfifoGBfullCnt[56]));
Q_MX02 U1076 ( .S(n406), .A0(n1047), .A1(gfifoGBfullCnt[57]), .Z(n593));
Q_FDP0UA U1077 ( .D(n593), .QTFCLK( ), .Q(gfifoGBfullCnt[57]));
Q_MX02 U1078 ( .S(n406), .A0(n1045), .A1(gfifoGBfullCnt[58]), .Z(n594));
Q_FDP0UA U1079 ( .D(n594), .QTFCLK( ), .Q(gfifoGBfullCnt[58]));
Q_MX02 U1080 ( .S(n406), .A0(n1043), .A1(gfifoGBfullCnt[59]), .Z(n595));
Q_FDP0UA U1081 ( .D(n595), .QTFCLK( ), .Q(gfifoGBfullCnt[59]));
Q_MX02 U1082 ( .S(n406), .A0(n1041), .A1(gfifoGBfullCnt[60]), .Z(n596));
Q_FDP0UA U1083 ( .D(n596), .QTFCLK( ), .Q(gfifoGBfullCnt[60]));
Q_MX02 U1084 ( .S(n406), .A0(n1039), .A1(gfifoGBfullCnt[61]), .Z(n597));
Q_FDP0UA U1085 ( .D(n597), .QTFCLK( ), .Q(gfifoGBfullCnt[61]));
Q_MX02 U1086 ( .S(n406), .A0(n1037), .A1(gfifoGBfullCnt[62]), .Z(n598));
Q_FDP0UA U1087 ( .D(n598), .QTFCLK( ), .Q(gfifoGBfullCnt[62]));
Q_FDP0UA U1088 ( .D(n599), .QTFCLK( ), .Q(gfifoGBfullCnt[63]));
Q_XOR2 U1089 ( .A0(n401), .A1(ixcHoldEcmCnt[0]), .Z(n600));
Q_FDP0UA U1090 ( .D(n600), .QTFCLK( ), .Q(ixcHoldEcmCnt[0]));
Q_MX02 U1091 ( .S(n407), .A0(n787), .A1(ixcHoldEcmCnt[1]), .Z(n601));
Q_FDP0UA U1092 ( .D(n601), .QTFCLK( ), .Q(ixcHoldEcmCnt[1]));
Q_MX02 U1093 ( .S(n407), .A0(n785), .A1(ixcHoldEcmCnt[2]), .Z(n602));
Q_FDP0UA U1094 ( .D(n602), .QTFCLK( ), .Q(ixcHoldEcmCnt[2]));
Q_MX02 U1095 ( .S(n407), .A0(n783), .A1(ixcHoldEcmCnt[3]), .Z(n603));
Q_FDP0UA U1096 ( .D(n603), .QTFCLK( ), .Q(ixcHoldEcmCnt[3]));
Q_MX02 U1097 ( .S(n407), .A0(n781), .A1(ixcHoldEcmCnt[4]), .Z(n604));
Q_FDP0UA U1098 ( .D(n604), .QTFCLK( ), .Q(ixcHoldEcmCnt[4]));
Q_MX02 U1099 ( .S(n407), .A0(n779), .A1(ixcHoldEcmCnt[5]), .Z(n605));
Q_FDP0UA U1100 ( .D(n605), .QTFCLK( ), .Q(ixcHoldEcmCnt[5]));
Q_MX02 U1101 ( .S(n407), .A0(n777), .A1(ixcHoldEcmCnt[6]), .Z(n606));
Q_FDP0UA U1102 ( .D(n606), .QTFCLK( ), .Q(ixcHoldEcmCnt[6]));
Q_MX02 U1103 ( .S(n407), .A0(n775), .A1(ixcHoldEcmCnt[7]), .Z(n607));
Q_FDP0UA U1104 ( .D(n607), .QTFCLK( ), .Q(ixcHoldEcmCnt[7]));
Q_MX02 U1105 ( .S(n407), .A0(n773), .A1(ixcHoldEcmCnt[8]), .Z(n608));
Q_FDP0UA U1106 ( .D(n608), .QTFCLK( ), .Q(ixcHoldEcmCnt[8]));
Q_MX02 U1107 ( .S(n407), .A0(n771), .A1(ixcHoldEcmCnt[9]), .Z(n609));
Q_FDP0UA U1108 ( .D(n609), .QTFCLK( ), .Q(ixcHoldEcmCnt[9]));
Q_MX02 U1109 ( .S(n407), .A0(n769), .A1(ixcHoldEcmCnt[10]), .Z(n610));
Q_FDP0UA U1110 ( .D(n610), .QTFCLK( ), .Q(ixcHoldEcmCnt[10]));
Q_MX02 U1111 ( .S(n407), .A0(n767), .A1(ixcHoldEcmCnt[11]), .Z(n611));
Q_FDP0UA U1112 ( .D(n611), .QTFCLK( ), .Q(ixcHoldEcmCnt[11]));
Q_MX02 U1113 ( .S(n407), .A0(n765), .A1(ixcHoldEcmCnt[12]), .Z(n612));
Q_FDP0UA U1114 ( .D(n612), .QTFCLK( ), .Q(ixcHoldEcmCnt[12]));
Q_MX02 U1115 ( .S(n407), .A0(n763), .A1(ixcHoldEcmCnt[13]), .Z(n613));
Q_FDP0UA U1116 ( .D(n613), .QTFCLK( ), .Q(ixcHoldEcmCnt[13]));
Q_MX02 U1117 ( .S(n407), .A0(n761), .A1(ixcHoldEcmCnt[14]), .Z(n614));
Q_FDP0UA U1118 ( .D(n614), .QTFCLK( ), .Q(ixcHoldEcmCnt[14]));
Q_MX02 U1119 ( .S(n407), .A0(n759), .A1(ixcHoldEcmCnt[15]), .Z(n615));
Q_FDP0UA U1120 ( .D(n615), .QTFCLK( ), .Q(ixcHoldEcmCnt[15]));
Q_MX02 U1121 ( .S(n407), .A0(n757), .A1(ixcHoldEcmCnt[16]), .Z(n616));
Q_FDP0UA U1122 ( .D(n616), .QTFCLK( ), .Q(ixcHoldEcmCnt[16]));
Q_MX02 U1123 ( .S(n407), .A0(n755), .A1(ixcHoldEcmCnt[17]), .Z(n617));
Q_FDP0UA U1124 ( .D(n617), .QTFCLK( ), .Q(ixcHoldEcmCnt[17]));
Q_MX02 U1125 ( .S(n407), .A0(n753), .A1(ixcHoldEcmCnt[18]), .Z(n618));
Q_FDP0UA U1126 ( .D(n618), .QTFCLK( ), .Q(ixcHoldEcmCnt[18]));
Q_MX02 U1127 ( .S(n407), .A0(n751), .A1(ixcHoldEcmCnt[19]), .Z(n619));
Q_FDP0UA U1128 ( .D(n619), .QTFCLK( ), .Q(ixcHoldEcmCnt[19]));
Q_MX02 U1129 ( .S(n407), .A0(n749), .A1(ixcHoldEcmCnt[20]), .Z(n620));
Q_FDP0UA U1130 ( .D(n620), .QTFCLK( ), .Q(ixcHoldEcmCnt[20]));
Q_MX02 U1131 ( .S(n407), .A0(n747), .A1(ixcHoldEcmCnt[21]), .Z(n621));
Q_FDP0UA U1132 ( .D(n621), .QTFCLK( ), .Q(ixcHoldEcmCnt[21]));
Q_MX02 U1133 ( .S(n407), .A0(n745), .A1(ixcHoldEcmCnt[22]), .Z(n622));
Q_FDP0UA U1134 ( .D(n622), .QTFCLK( ), .Q(ixcHoldEcmCnt[22]));
Q_MX02 U1135 ( .S(n407), .A0(n743), .A1(ixcHoldEcmCnt[23]), .Z(n623));
Q_FDP0UA U1136 ( .D(n623), .QTFCLK( ), .Q(ixcHoldEcmCnt[23]));
Q_MX02 U1137 ( .S(n407), .A0(n741), .A1(ixcHoldEcmCnt[24]), .Z(n624));
Q_FDP0UA U1138 ( .D(n624), .QTFCLK( ), .Q(ixcHoldEcmCnt[24]));
Q_MX02 U1139 ( .S(n407), .A0(n739), .A1(ixcHoldEcmCnt[25]), .Z(n625));
Q_FDP0UA U1140 ( .D(n625), .QTFCLK( ), .Q(ixcHoldEcmCnt[25]));
Q_MX02 U1141 ( .S(n407), .A0(n737), .A1(ixcHoldEcmCnt[26]), .Z(n626));
Q_FDP0UA U1142 ( .D(n626), .QTFCLK( ), .Q(ixcHoldEcmCnt[26]));
Q_MX02 U1143 ( .S(n407), .A0(n735), .A1(ixcHoldEcmCnt[27]), .Z(n627));
Q_FDP0UA U1144 ( .D(n627), .QTFCLK( ), .Q(ixcHoldEcmCnt[27]));
Q_MX02 U1145 ( .S(n407), .A0(n733), .A1(ixcHoldEcmCnt[28]), .Z(n628));
Q_FDP0UA U1146 ( .D(n628), .QTFCLK( ), .Q(ixcHoldEcmCnt[28]));
Q_MX02 U1147 ( .S(n407), .A0(n731), .A1(ixcHoldEcmCnt[29]), .Z(n629));
Q_FDP0UA U1148 ( .D(n629), .QTFCLK( ), .Q(ixcHoldEcmCnt[29]));
Q_MX02 U1149 ( .S(n407), .A0(n729), .A1(ixcHoldEcmCnt[30]), .Z(n630));
Q_FDP0UA U1150 ( .D(n630), .QTFCLK( ), .Q(ixcHoldEcmCnt[30]));
Q_MX02 U1151 ( .S(n407), .A0(n727), .A1(ixcHoldEcmCnt[31]), .Z(n631));
Q_FDP0UA U1152 ( .D(n631), .QTFCLK( ), .Q(ixcHoldEcmCnt[31]));
Q_MX02 U1153 ( .S(n407), .A0(n725), .A1(ixcHoldEcmCnt[32]), .Z(n632));
Q_FDP0UA U1154 ( .D(n632), .QTFCLK( ), .Q(ixcHoldEcmCnt[32]));
Q_MX02 U1155 ( .S(n407), .A0(n723), .A1(ixcHoldEcmCnt[33]), .Z(n633));
Q_FDP0UA U1156 ( .D(n633), .QTFCLK( ), .Q(ixcHoldEcmCnt[33]));
Q_MX02 U1157 ( .S(n407), .A0(n721), .A1(ixcHoldEcmCnt[34]), .Z(n634));
Q_FDP0UA U1158 ( .D(n634), .QTFCLK( ), .Q(ixcHoldEcmCnt[34]));
Q_MX02 U1159 ( .S(n407), .A0(n719), .A1(ixcHoldEcmCnt[35]), .Z(n635));
Q_FDP0UA U1160 ( .D(n635), .QTFCLK( ), .Q(ixcHoldEcmCnt[35]));
Q_MX02 U1161 ( .S(n407), .A0(n717), .A1(ixcHoldEcmCnt[36]), .Z(n636));
Q_FDP0UA U1162 ( .D(n636), .QTFCLK( ), .Q(ixcHoldEcmCnt[36]));
Q_MX02 U1163 ( .S(n407), .A0(n715), .A1(ixcHoldEcmCnt[37]), .Z(n637));
Q_FDP0UA U1164 ( .D(n637), .QTFCLK( ), .Q(ixcHoldEcmCnt[37]));
Q_MX02 U1165 ( .S(n407), .A0(n713), .A1(ixcHoldEcmCnt[38]), .Z(n638));
Q_FDP0UA U1166 ( .D(n638), .QTFCLK( ), .Q(ixcHoldEcmCnt[38]));
Q_MX02 U1167 ( .S(n407), .A0(n711), .A1(ixcHoldEcmCnt[39]), .Z(n639));
Q_FDP0UA U1168 ( .D(n639), .QTFCLK( ), .Q(ixcHoldEcmCnt[39]));
Q_MX02 U1169 ( .S(n407), .A0(n709), .A1(ixcHoldEcmCnt[40]), .Z(n640));
Q_FDP0UA U1170 ( .D(n640), .QTFCLK( ), .Q(ixcHoldEcmCnt[40]));
Q_MX02 U1171 ( .S(n407), .A0(n707), .A1(ixcHoldEcmCnt[41]), .Z(n641));
Q_FDP0UA U1172 ( .D(n641), .QTFCLK( ), .Q(ixcHoldEcmCnt[41]));
Q_MX02 U1173 ( .S(n407), .A0(n705), .A1(ixcHoldEcmCnt[42]), .Z(n642));
Q_FDP0UA U1174 ( .D(n642), .QTFCLK( ), .Q(ixcHoldEcmCnt[42]));
Q_MX02 U1175 ( .S(n407), .A0(n703), .A1(ixcHoldEcmCnt[43]), .Z(n643));
Q_FDP0UA U1176 ( .D(n643), .QTFCLK( ), .Q(ixcHoldEcmCnt[43]));
Q_MX02 U1177 ( .S(n407), .A0(n701), .A1(ixcHoldEcmCnt[44]), .Z(n644));
Q_FDP0UA U1178 ( .D(n644), .QTFCLK( ), .Q(ixcHoldEcmCnt[44]));
Q_MX02 U1179 ( .S(n407), .A0(n699), .A1(ixcHoldEcmCnt[45]), .Z(n645));
Q_FDP0UA U1180 ( .D(n645), .QTFCLK( ), .Q(ixcHoldEcmCnt[45]));
Q_MX02 U1181 ( .S(n407), .A0(n697), .A1(ixcHoldEcmCnt[46]), .Z(n646));
Q_FDP0UA U1182 ( .D(n646), .QTFCLK( ), .Q(ixcHoldEcmCnt[46]));
Q_MX02 U1183 ( .S(n407), .A0(n695), .A1(ixcHoldEcmCnt[47]), .Z(n647));
Q_FDP0UA U1184 ( .D(n647), .QTFCLK( ), .Q(ixcHoldEcmCnt[47]));
Q_MX02 U1185 ( .S(n407), .A0(n693), .A1(ixcHoldEcmCnt[48]), .Z(n648));
Q_FDP0UA U1186 ( .D(n648), .QTFCLK( ), .Q(ixcHoldEcmCnt[48]));
Q_MX02 U1187 ( .S(n407), .A0(n691), .A1(ixcHoldEcmCnt[49]), .Z(n649));
Q_FDP0UA U1188 ( .D(n649), .QTFCLK( ), .Q(ixcHoldEcmCnt[49]));
Q_MX02 U1189 ( .S(n407), .A0(n689), .A1(ixcHoldEcmCnt[50]), .Z(n650));
Q_FDP0UA U1190 ( .D(n650), .QTFCLK( ), .Q(ixcHoldEcmCnt[50]));
Q_MX02 U1191 ( .S(n407), .A0(n687), .A1(ixcHoldEcmCnt[51]), .Z(n651));
Q_FDP0UA U1192 ( .D(n651), .QTFCLK( ), .Q(ixcHoldEcmCnt[51]));
Q_MX02 U1193 ( .S(n407), .A0(n685), .A1(ixcHoldEcmCnt[52]), .Z(n652));
Q_FDP0UA U1194 ( .D(n652), .QTFCLK( ), .Q(ixcHoldEcmCnt[52]));
Q_MX02 U1195 ( .S(n407), .A0(n683), .A1(ixcHoldEcmCnt[53]), .Z(n653));
Q_FDP0UA U1196 ( .D(n653), .QTFCLK( ), .Q(ixcHoldEcmCnt[53]));
Q_MX02 U1197 ( .S(n407), .A0(n681), .A1(ixcHoldEcmCnt[54]), .Z(n654));
Q_FDP0UA U1198 ( .D(n654), .QTFCLK( ), .Q(ixcHoldEcmCnt[54]));
Q_MX02 U1199 ( .S(n407), .A0(n679), .A1(ixcHoldEcmCnt[55]), .Z(n655));
Q_FDP0UA U1200 ( .D(n655), .QTFCLK( ), .Q(ixcHoldEcmCnt[55]));
Q_MX02 U1201 ( .S(n407), .A0(n677), .A1(ixcHoldEcmCnt[56]), .Z(n656));
Q_FDP0UA U1202 ( .D(n656), .QTFCLK( ), .Q(ixcHoldEcmCnt[56]));
Q_MX02 U1203 ( .S(n407), .A0(n675), .A1(ixcHoldEcmCnt[57]), .Z(n657));
Q_FDP0UA U1204 ( .D(n657), .QTFCLK( ), .Q(ixcHoldEcmCnt[57]));
Q_MX02 U1205 ( .S(n407), .A0(n673), .A1(ixcHoldEcmCnt[58]), .Z(n658));
Q_FDP0UA U1206 ( .D(n658), .QTFCLK( ), .Q(ixcHoldEcmCnt[58]));
Q_MX02 U1207 ( .S(n407), .A0(n671), .A1(ixcHoldEcmCnt[59]), .Z(n659));
Q_FDP0UA U1208 ( .D(n659), .QTFCLK( ), .Q(ixcHoldEcmCnt[59]));
Q_MX02 U1209 ( .S(n407), .A0(n669), .A1(ixcHoldEcmCnt[60]), .Z(n660));
Q_FDP0UA U1210 ( .D(n660), .QTFCLK( ), .Q(ixcHoldEcmCnt[60]));
Q_MX02 U1211 ( .S(n407), .A0(n667), .A1(ixcHoldEcmCnt[61]), .Z(n661));
Q_FDP0UA U1212 ( .D(n661), .QTFCLK( ), .Q(ixcHoldEcmCnt[61]));
Q_MX02 U1213 ( .S(n407), .A0(n665), .A1(ixcHoldEcmCnt[62]), .Z(n662));
Q_FDP0UA U1214 ( .D(n662), .QTFCLK( ), .Q(ixcHoldEcmCnt[62]));
Q_FDP0UA U1215 ( .D(n663), .QTFCLK( ), .Q(ixcHoldEcmCnt[63]));
Q_XOR2 U1216 ( .A0(ixcHoldEcmCnt[63]), .A1(n11), .Z(n663));
Q_AD01HF U1217 ( .A0(ixcHoldEcmCnt[62]), .B0(n666), .S(n665), .CO(n664));
Q_AD01HF U1218 ( .A0(ixcHoldEcmCnt[61]), .B0(n668), .S(n667), .CO(n666));
Q_AD01HF U1219 ( .A0(ixcHoldEcmCnt[60]), .B0(n670), .S(n669), .CO(n668));
Q_AD01HF U1220 ( .A0(ixcHoldEcmCnt[59]), .B0(n672), .S(n671), .CO(n670));
Q_AD01HF U1221 ( .A0(ixcHoldEcmCnt[58]), .B0(n674), .S(n673), .CO(n672));
Q_AD01HF U1222 ( .A0(ixcHoldEcmCnt[57]), .B0(n676), .S(n675), .CO(n674));
Q_AD01HF U1223 ( .A0(ixcHoldEcmCnt[56]), .B0(n678), .S(n677), .CO(n676));
Q_AD01HF U1224 ( .A0(ixcHoldEcmCnt[55]), .B0(n680), .S(n679), .CO(n678));
Q_AD01HF U1225 ( .A0(ixcHoldEcmCnt[54]), .B0(n682), .S(n681), .CO(n680));
Q_AD01HF U1226 ( .A0(ixcHoldEcmCnt[53]), .B0(n684), .S(n683), .CO(n682));
Q_AD01HF U1227 ( .A0(ixcHoldEcmCnt[52]), .B0(n686), .S(n685), .CO(n684));
Q_AD01HF U1228 ( .A0(ixcHoldEcmCnt[51]), .B0(n688), .S(n687), .CO(n686));
Q_AD01HF U1229 ( .A0(ixcHoldEcmCnt[50]), .B0(n690), .S(n689), .CO(n688));
Q_AD01HF U1230 ( .A0(ixcHoldEcmCnt[49]), .B0(n692), .S(n691), .CO(n690));
Q_AD01HF U1231 ( .A0(ixcHoldEcmCnt[48]), .B0(n694), .S(n693), .CO(n692));
Q_AD01HF U1232 ( .A0(ixcHoldEcmCnt[47]), .B0(n696), .S(n695), .CO(n694));
Q_AD01HF U1233 ( .A0(ixcHoldEcmCnt[46]), .B0(n698), .S(n697), .CO(n696));
Q_AD01HF U1234 ( .A0(ixcHoldEcmCnt[45]), .B0(n700), .S(n699), .CO(n698));
Q_AD01HF U1235 ( .A0(ixcHoldEcmCnt[44]), .B0(n702), .S(n701), .CO(n700));
Q_AD01HF U1236 ( .A0(ixcHoldEcmCnt[43]), .B0(n704), .S(n703), .CO(n702));
Q_AD01HF U1237 ( .A0(ixcHoldEcmCnt[42]), .B0(n706), .S(n705), .CO(n704));
Q_AD01HF U1238 ( .A0(ixcHoldEcmCnt[41]), .B0(n708), .S(n707), .CO(n706));
Q_AD01HF U1239 ( .A0(ixcHoldEcmCnt[40]), .B0(n710), .S(n709), .CO(n708));
Q_AD01HF U1240 ( .A0(ixcHoldEcmCnt[39]), .B0(n712), .S(n711), .CO(n710));
Q_AD01HF U1241 ( .A0(ixcHoldEcmCnt[38]), .B0(n714), .S(n713), .CO(n712));
Q_AD01HF U1242 ( .A0(ixcHoldEcmCnt[37]), .B0(n716), .S(n715), .CO(n714));
Q_AD01HF U1243 ( .A0(ixcHoldEcmCnt[36]), .B0(n718), .S(n717), .CO(n716));
Q_AD01HF U1244 ( .A0(ixcHoldEcmCnt[35]), .B0(n720), .S(n719), .CO(n718));
Q_AD01HF U1245 ( .A0(ixcHoldEcmCnt[34]), .B0(n722), .S(n721), .CO(n720));
Q_AD01HF U1246 ( .A0(ixcHoldEcmCnt[33]), .B0(n724), .S(n723), .CO(n722));
Q_AD01HF U1247 ( .A0(ixcHoldEcmCnt[32]), .B0(n726), .S(n725), .CO(n724));
Q_AD01HF U1248 ( .A0(ixcHoldEcmCnt[31]), .B0(n728), .S(n727), .CO(n726));
Q_AD01HF U1249 ( .A0(ixcHoldEcmCnt[30]), .B0(n730), .S(n729), .CO(n728));
Q_AD01HF U1250 ( .A0(ixcHoldEcmCnt[29]), .B0(n732), .S(n731), .CO(n730));
Q_AD01HF U1251 ( .A0(ixcHoldEcmCnt[28]), .B0(n734), .S(n733), .CO(n732));
Q_AD01HF U1252 ( .A0(ixcHoldEcmCnt[27]), .B0(n736), .S(n735), .CO(n734));
Q_AD01HF U1253 ( .A0(ixcHoldEcmCnt[26]), .B0(n738), .S(n737), .CO(n736));
Q_AD01HF U1254 ( .A0(ixcHoldEcmCnt[25]), .B0(n740), .S(n739), .CO(n738));
Q_AD01HF U1255 ( .A0(ixcHoldEcmCnt[24]), .B0(n742), .S(n741), .CO(n740));
Q_AD01HF U1256 ( .A0(ixcHoldEcmCnt[23]), .B0(n744), .S(n743), .CO(n742));
Q_AD01HF U1257 ( .A0(ixcHoldEcmCnt[22]), .B0(n746), .S(n745), .CO(n744));
Q_AD01HF U1258 ( .A0(ixcHoldEcmCnt[21]), .B0(n748), .S(n747), .CO(n746));
Q_AD01HF U1259 ( .A0(ixcHoldEcmCnt[20]), .B0(n750), .S(n749), .CO(n748));
Q_AD01HF U1260 ( .A0(ixcHoldEcmCnt[19]), .B0(n752), .S(n751), .CO(n750));
Q_AD01HF U1261 ( .A0(ixcHoldEcmCnt[18]), .B0(n754), .S(n753), .CO(n752));
Q_AD01HF U1262 ( .A0(ixcHoldEcmCnt[17]), .B0(n756), .S(n755), .CO(n754));
Q_AD01HF U1263 ( .A0(ixcHoldEcmCnt[16]), .B0(n758), .S(n757), .CO(n756));
Q_AD01HF U1264 ( .A0(ixcHoldEcmCnt[15]), .B0(n760), .S(n759), .CO(n758));
Q_AD01HF U1265 ( .A0(ixcHoldEcmCnt[14]), .B0(n762), .S(n761), .CO(n760));
Q_AD01HF U1266 ( .A0(ixcHoldEcmCnt[13]), .B0(n764), .S(n763), .CO(n762));
Q_AD01HF U1267 ( .A0(ixcHoldEcmCnt[12]), .B0(n766), .S(n765), .CO(n764));
Q_AD01HF U1268 ( .A0(ixcHoldEcmCnt[11]), .B0(n768), .S(n767), .CO(n766));
Q_AD01HF U1269 ( .A0(ixcHoldEcmCnt[10]), .B0(n770), .S(n769), .CO(n768));
Q_AD01HF U1270 ( .A0(ixcHoldEcmCnt[9]), .B0(n772), .S(n771), .CO(n770));
Q_AD01HF U1271 ( .A0(ixcHoldEcmCnt[8]), .B0(n774), .S(n773), .CO(n772));
Q_AD01HF U1272 ( .A0(ixcHoldEcmCnt[7]), .B0(n776), .S(n775), .CO(n774));
Q_AD01HF U1273 ( .A0(ixcHoldEcmCnt[6]), .B0(n778), .S(n777), .CO(n776));
Q_AD01HF U1274 ( .A0(ixcHoldEcmCnt[5]), .B0(n780), .S(n779), .CO(n778));
Q_AD01HF U1275 ( .A0(ixcHoldEcmCnt[4]), .B0(n782), .S(n781), .CO(n780));
Q_AD01HF U1276 ( .A0(ixcHoldEcmCnt[3]), .B0(n784), .S(n783), .CO(n782));
Q_AD01HF U1277 ( .A0(ixcHoldEcmCnt[2]), .B0(n786), .S(n785), .CO(n784));
Q_AD01HF U1278 ( .A0(ixcHoldEcmCnt[1]), .B0(ixcHoldEcmCnt[0]), .S(n787), .CO(n786));
Q_XOR2 U1279 ( .A0(gfifoTBsyncCnt[63]), .A1(n14), .Z(n471));
Q_AD01HF U1280 ( .A0(gfifoTBsyncCnt[62]), .B0(n790), .S(n789), .CO(n788));
Q_AD01HF U1281 ( .A0(gfifoTBsyncCnt[61]), .B0(n792), .S(n791), .CO(n790));
Q_AD01HF U1282 ( .A0(gfifoTBsyncCnt[60]), .B0(n794), .S(n793), .CO(n792));
Q_AD01HF U1283 ( .A0(gfifoTBsyncCnt[59]), .B0(n796), .S(n795), .CO(n794));
Q_AD01HF U1284 ( .A0(gfifoTBsyncCnt[58]), .B0(n798), .S(n797), .CO(n796));
Q_AD01HF U1285 ( .A0(gfifoTBsyncCnt[57]), .B0(n800), .S(n799), .CO(n798));
Q_AD01HF U1286 ( .A0(gfifoTBsyncCnt[56]), .B0(n802), .S(n801), .CO(n800));
Q_AD01HF U1287 ( .A0(gfifoTBsyncCnt[55]), .B0(n804), .S(n803), .CO(n802));
Q_AD01HF U1288 ( .A0(gfifoTBsyncCnt[54]), .B0(n806), .S(n805), .CO(n804));
Q_AD01HF U1289 ( .A0(gfifoTBsyncCnt[53]), .B0(n808), .S(n807), .CO(n806));
Q_AD01HF U1290 ( .A0(gfifoTBsyncCnt[52]), .B0(n810), .S(n809), .CO(n808));
Q_AD01HF U1291 ( .A0(gfifoTBsyncCnt[51]), .B0(n812), .S(n811), .CO(n810));
Q_AD01HF U1292 ( .A0(gfifoTBsyncCnt[50]), .B0(n814), .S(n813), .CO(n812));
Q_AD01HF U1293 ( .A0(gfifoTBsyncCnt[49]), .B0(n816), .S(n815), .CO(n814));
Q_AD01HF U1294 ( .A0(gfifoTBsyncCnt[48]), .B0(n818), .S(n817), .CO(n816));
Q_AD01HF U1295 ( .A0(gfifoTBsyncCnt[47]), .B0(n820), .S(n819), .CO(n818));
Q_AD01HF U1296 ( .A0(gfifoTBsyncCnt[46]), .B0(n822), .S(n821), .CO(n820));
Q_AD01HF U1297 ( .A0(gfifoTBsyncCnt[45]), .B0(n824), .S(n823), .CO(n822));
Q_AD01HF U1298 ( .A0(gfifoTBsyncCnt[44]), .B0(n826), .S(n825), .CO(n824));
Q_AD01HF U1299 ( .A0(gfifoTBsyncCnt[43]), .B0(n828), .S(n827), .CO(n826));
Q_AD01HF U1300 ( .A0(gfifoTBsyncCnt[42]), .B0(n830), .S(n829), .CO(n828));
Q_AD01HF U1301 ( .A0(gfifoTBsyncCnt[41]), .B0(n832), .S(n831), .CO(n830));
Q_AD01HF U1302 ( .A0(gfifoTBsyncCnt[40]), .B0(n834), .S(n833), .CO(n832));
Q_AD01HF U1303 ( .A0(gfifoTBsyncCnt[39]), .B0(n836), .S(n835), .CO(n834));
Q_AD01HF U1304 ( .A0(gfifoTBsyncCnt[38]), .B0(n838), .S(n837), .CO(n836));
Q_AD01HF U1305 ( .A0(gfifoTBsyncCnt[37]), .B0(n840), .S(n839), .CO(n838));
Q_AD01HF U1306 ( .A0(gfifoTBsyncCnt[36]), .B0(n842), .S(n841), .CO(n840));
Q_AD01HF U1307 ( .A0(gfifoTBsyncCnt[35]), .B0(n844), .S(n843), .CO(n842));
Q_AD01HF U1308 ( .A0(gfifoTBsyncCnt[34]), .B0(n846), .S(n845), .CO(n844));
Q_AD01HF U1309 ( .A0(gfifoTBsyncCnt[33]), .B0(n848), .S(n847), .CO(n846));
Q_AD01HF U1310 ( .A0(gfifoTBsyncCnt[32]), .B0(n850), .S(n849), .CO(n848));
Q_AD01HF U1311 ( .A0(gfifoTBsyncCnt[31]), .B0(n852), .S(n851), .CO(n850));
Q_AD01HF U1312 ( .A0(gfifoTBsyncCnt[30]), .B0(n854), .S(n853), .CO(n852));
Q_AD01HF U1313 ( .A0(gfifoTBsyncCnt[29]), .B0(n856), .S(n855), .CO(n854));
Q_AD01HF U1314 ( .A0(gfifoTBsyncCnt[28]), .B0(n858), .S(n857), .CO(n856));
Q_AD01HF U1315 ( .A0(gfifoTBsyncCnt[27]), .B0(n860), .S(n859), .CO(n858));
Q_AD01HF U1316 ( .A0(gfifoTBsyncCnt[26]), .B0(n862), .S(n861), .CO(n860));
Q_AD01HF U1317 ( .A0(gfifoTBsyncCnt[25]), .B0(n864), .S(n863), .CO(n862));
Q_AD01HF U1318 ( .A0(gfifoTBsyncCnt[24]), .B0(n866), .S(n865), .CO(n864));
Q_AD01HF U1319 ( .A0(gfifoTBsyncCnt[23]), .B0(n868), .S(n867), .CO(n866));
Q_AD01HF U1320 ( .A0(gfifoTBsyncCnt[22]), .B0(n870), .S(n869), .CO(n868));
Q_AD01HF U1321 ( .A0(gfifoTBsyncCnt[21]), .B0(n872), .S(n871), .CO(n870));
Q_AD01HF U1322 ( .A0(gfifoTBsyncCnt[20]), .B0(n874), .S(n873), .CO(n872));
Q_AD01HF U1323 ( .A0(gfifoTBsyncCnt[19]), .B0(n876), .S(n875), .CO(n874));
Q_AD01HF U1324 ( .A0(gfifoTBsyncCnt[18]), .B0(n878), .S(n877), .CO(n876));
Q_AD01HF U1325 ( .A0(gfifoTBsyncCnt[17]), .B0(n880), .S(n879), .CO(n878));
Q_AD01HF U1326 ( .A0(gfifoTBsyncCnt[16]), .B0(n882), .S(n881), .CO(n880));
Q_AD01HF U1327 ( .A0(gfifoTBsyncCnt[15]), .B0(n884), .S(n883), .CO(n882));
Q_AD01HF U1328 ( .A0(gfifoTBsyncCnt[14]), .B0(n886), .S(n885), .CO(n884));
Q_AD01HF U1329 ( .A0(gfifoTBsyncCnt[13]), .B0(n888), .S(n887), .CO(n886));
Q_AD01HF U1330 ( .A0(gfifoTBsyncCnt[12]), .B0(n890), .S(n889), .CO(n888));
Q_AD01HF U1331 ( .A0(gfifoTBsyncCnt[11]), .B0(n892), .S(n891), .CO(n890));
Q_AD01HF U1332 ( .A0(gfifoTBsyncCnt[10]), .B0(n894), .S(n893), .CO(n892));
Q_AD01HF U1333 ( .A0(gfifoTBsyncCnt[9]), .B0(n896), .S(n895), .CO(n894));
Q_AD01HF U1334 ( .A0(gfifoTBsyncCnt[8]), .B0(n898), .S(n897), .CO(n896));
Q_AD01HF U1335 ( .A0(gfifoTBsyncCnt[7]), .B0(n900), .S(n899), .CO(n898));
Q_AD01HF U1336 ( .A0(gfifoTBsyncCnt[6]), .B0(n902), .S(n901), .CO(n900));
Q_AD01HF U1337 ( .A0(gfifoTBsyncCnt[5]), .B0(n904), .S(n903), .CO(n902));
Q_AD01HF U1338 ( .A0(gfifoTBsyncCnt[4]), .B0(n906), .S(n905), .CO(n904));
Q_AD01HF U1339 ( .A0(gfifoTBsyncCnt[3]), .B0(n908), .S(n907), .CO(n906));
Q_AD01HF U1340 ( .A0(gfifoTBsyncCnt[2]), .B0(n910), .S(n909), .CO(n908));
Q_AD01HF U1341 ( .A0(gfifoTBsyncCnt[1]), .B0(gfifoTBsyncCnt[0]), .S(n911), .CO(n910));
Q_XOR2 U1342 ( .A0(gfifoLBfullCnt[63]), .A1(n13), .Z(n535));
Q_AD01HF U1343 ( .A0(gfifoLBfullCnt[62]), .B0(n914), .S(n913), .CO(n912));
Q_AD01HF U1344 ( .A0(gfifoLBfullCnt[61]), .B0(n916), .S(n915), .CO(n914));
Q_AD01HF U1345 ( .A0(gfifoLBfullCnt[60]), .B0(n918), .S(n917), .CO(n916));
Q_AD01HF U1346 ( .A0(gfifoLBfullCnt[59]), .B0(n920), .S(n919), .CO(n918));
Q_AD01HF U1347 ( .A0(gfifoLBfullCnt[58]), .B0(n922), .S(n921), .CO(n920));
Q_AD01HF U1348 ( .A0(gfifoLBfullCnt[57]), .B0(n924), .S(n923), .CO(n922));
Q_AD01HF U1349 ( .A0(gfifoLBfullCnt[56]), .B0(n926), .S(n925), .CO(n924));
Q_AD01HF U1350 ( .A0(gfifoLBfullCnt[55]), .B0(n928), .S(n927), .CO(n926));
Q_AD01HF U1351 ( .A0(gfifoLBfullCnt[54]), .B0(n930), .S(n929), .CO(n928));
Q_AD01HF U1352 ( .A0(gfifoLBfullCnt[53]), .B0(n932), .S(n931), .CO(n930));
Q_AD01HF U1353 ( .A0(gfifoLBfullCnt[52]), .B0(n934), .S(n933), .CO(n932));
Q_AD01HF U1354 ( .A0(gfifoLBfullCnt[51]), .B0(n936), .S(n935), .CO(n934));
Q_AD01HF U1355 ( .A0(gfifoLBfullCnt[50]), .B0(n938), .S(n937), .CO(n936));
Q_AD01HF U1356 ( .A0(gfifoLBfullCnt[49]), .B0(n940), .S(n939), .CO(n938));
Q_AD01HF U1357 ( .A0(gfifoLBfullCnt[48]), .B0(n942), .S(n941), .CO(n940));
Q_AD01HF U1358 ( .A0(gfifoLBfullCnt[47]), .B0(n944), .S(n943), .CO(n942));
Q_AD01HF U1359 ( .A0(gfifoLBfullCnt[46]), .B0(n946), .S(n945), .CO(n944));
Q_AD01HF U1360 ( .A0(gfifoLBfullCnt[45]), .B0(n948), .S(n947), .CO(n946));
Q_AD01HF U1361 ( .A0(gfifoLBfullCnt[44]), .B0(n950), .S(n949), .CO(n948));
Q_AD01HF U1362 ( .A0(gfifoLBfullCnt[43]), .B0(n952), .S(n951), .CO(n950));
Q_AD01HF U1363 ( .A0(gfifoLBfullCnt[42]), .B0(n954), .S(n953), .CO(n952));
Q_AD01HF U1364 ( .A0(gfifoLBfullCnt[41]), .B0(n956), .S(n955), .CO(n954));
Q_AD01HF U1365 ( .A0(gfifoLBfullCnt[40]), .B0(n958), .S(n957), .CO(n956));
Q_AD01HF U1366 ( .A0(gfifoLBfullCnt[39]), .B0(n960), .S(n959), .CO(n958));
Q_AD01HF U1367 ( .A0(gfifoLBfullCnt[38]), .B0(n962), .S(n961), .CO(n960));
Q_AD01HF U1368 ( .A0(gfifoLBfullCnt[37]), .B0(n964), .S(n963), .CO(n962));
Q_AD01HF U1369 ( .A0(gfifoLBfullCnt[36]), .B0(n966), .S(n965), .CO(n964));
Q_AD01HF U1370 ( .A0(gfifoLBfullCnt[35]), .B0(n968), .S(n967), .CO(n966));
Q_AD01HF U1371 ( .A0(gfifoLBfullCnt[34]), .B0(n970), .S(n969), .CO(n968));
Q_AD01HF U1372 ( .A0(gfifoLBfullCnt[33]), .B0(n972), .S(n971), .CO(n970));
Q_AD01HF U1373 ( .A0(gfifoLBfullCnt[32]), .B0(n974), .S(n973), .CO(n972));
Q_AD01HF U1374 ( .A0(gfifoLBfullCnt[31]), .B0(n976), .S(n975), .CO(n974));
Q_AD01HF U1375 ( .A0(gfifoLBfullCnt[30]), .B0(n978), .S(n977), .CO(n976));
Q_AD01HF U1376 ( .A0(gfifoLBfullCnt[29]), .B0(n980), .S(n979), .CO(n978));
Q_AD01HF U1377 ( .A0(gfifoLBfullCnt[28]), .B0(n982), .S(n981), .CO(n980));
Q_AD01HF U1378 ( .A0(gfifoLBfullCnt[27]), .B0(n984), .S(n983), .CO(n982));
Q_AD01HF U1379 ( .A0(gfifoLBfullCnt[26]), .B0(n986), .S(n985), .CO(n984));
Q_AD01HF U1380 ( .A0(gfifoLBfullCnt[25]), .B0(n988), .S(n987), .CO(n986));
Q_AD01HF U1381 ( .A0(gfifoLBfullCnt[24]), .B0(n990), .S(n989), .CO(n988));
Q_AD01HF U1382 ( .A0(gfifoLBfullCnt[23]), .B0(n992), .S(n991), .CO(n990));
Q_AD01HF U1383 ( .A0(gfifoLBfullCnt[22]), .B0(n994), .S(n993), .CO(n992));
Q_AD01HF U1384 ( .A0(gfifoLBfullCnt[21]), .B0(n996), .S(n995), .CO(n994));
Q_AD01HF U1385 ( .A0(gfifoLBfullCnt[20]), .B0(n998), .S(n997), .CO(n996));
Q_AD01HF U1386 ( .A0(gfifoLBfullCnt[19]), .B0(n1000), .S(n999), .CO(n998));
Q_AD01HF U1387 ( .A0(gfifoLBfullCnt[18]), .B0(n1002), .S(n1001), .CO(n1000));
Q_AD01HF U1388 ( .A0(gfifoLBfullCnt[17]), .B0(n1004), .S(n1003), .CO(n1002));
Q_AD01HF U1389 ( .A0(gfifoLBfullCnt[16]), .B0(n1006), .S(n1005), .CO(n1004));
Q_AD01HF U1390 ( .A0(gfifoLBfullCnt[15]), .B0(n1008), .S(n1007), .CO(n1006));
Q_AD01HF U1391 ( .A0(gfifoLBfullCnt[14]), .B0(n1010), .S(n1009), .CO(n1008));
Q_AD01HF U1392 ( .A0(gfifoLBfullCnt[13]), .B0(n1012), .S(n1011), .CO(n1010));
Q_AD01HF U1393 ( .A0(gfifoLBfullCnt[12]), .B0(n1014), .S(n1013), .CO(n1012));
Q_AD01HF U1394 ( .A0(gfifoLBfullCnt[11]), .B0(n1016), .S(n1015), .CO(n1014));
Q_AD01HF U1395 ( .A0(gfifoLBfullCnt[10]), .B0(n1018), .S(n1017), .CO(n1016));
Q_AD01HF U1396 ( .A0(gfifoLBfullCnt[9]), .B0(n1020), .S(n1019), .CO(n1018));
Q_AD01HF U1397 ( .A0(gfifoLBfullCnt[8]), .B0(n1022), .S(n1021), .CO(n1020));
Q_AD01HF U1398 ( .A0(gfifoLBfullCnt[7]), .B0(n1024), .S(n1023), .CO(n1022));
Q_AD01HF U1399 ( .A0(gfifoLBfullCnt[6]), .B0(n1026), .S(n1025), .CO(n1024));
Q_AD01HF U1400 ( .A0(gfifoLBfullCnt[5]), .B0(n1028), .S(n1027), .CO(n1026));
Q_AD01HF U1401 ( .A0(gfifoLBfullCnt[4]), .B0(n1030), .S(n1029), .CO(n1028));
Q_AD01HF U1402 ( .A0(gfifoLBfullCnt[3]), .B0(n1032), .S(n1031), .CO(n1030));
Q_AD01HF U1403 ( .A0(gfifoLBfullCnt[2]), .B0(n1034), .S(n1033), .CO(n1032));
Q_AD01HF U1404 ( .A0(gfifoLBfullCnt[1]), .B0(gfifoLBfullCnt[0]), .S(n1035), .CO(n1034));
Q_XOR2 U1405 ( .A0(gfifoGBfullCnt[63]), .A1(n12), .Z(n599));
Q_AD01HF U1406 ( .A0(gfifoGBfullCnt[62]), .B0(n1038), .S(n1037), .CO(n1036));
Q_AD01HF U1407 ( .A0(gfifoGBfullCnt[61]), .B0(n1040), .S(n1039), .CO(n1038));
Q_AD01HF U1408 ( .A0(gfifoGBfullCnt[60]), .B0(n1042), .S(n1041), .CO(n1040));
Q_AD01HF U1409 ( .A0(gfifoGBfullCnt[59]), .B0(n1044), .S(n1043), .CO(n1042));
Q_AD01HF U1410 ( .A0(gfifoGBfullCnt[58]), .B0(n1046), .S(n1045), .CO(n1044));
Q_AD01HF U1411 ( .A0(gfifoGBfullCnt[57]), .B0(n1048), .S(n1047), .CO(n1046));
Q_AD01HF U1412 ( .A0(gfifoGBfullCnt[56]), .B0(n1050), .S(n1049), .CO(n1048));
Q_AD01HF U1413 ( .A0(gfifoGBfullCnt[55]), .B0(n1052), .S(n1051), .CO(n1050));
Q_AD01HF U1414 ( .A0(gfifoGBfullCnt[54]), .B0(n1054), .S(n1053), .CO(n1052));
Q_AD01HF U1415 ( .A0(gfifoGBfullCnt[53]), .B0(n1056), .S(n1055), .CO(n1054));
Q_AD01HF U1416 ( .A0(gfifoGBfullCnt[52]), .B0(n1058), .S(n1057), .CO(n1056));
Q_AD01HF U1417 ( .A0(gfifoGBfullCnt[51]), .B0(n1060), .S(n1059), .CO(n1058));
Q_AD01HF U1418 ( .A0(gfifoGBfullCnt[50]), .B0(n1062), .S(n1061), .CO(n1060));
Q_AD01HF U1419 ( .A0(gfifoGBfullCnt[49]), .B0(n1064), .S(n1063), .CO(n1062));
Q_AD01HF U1420 ( .A0(gfifoGBfullCnt[48]), .B0(n1066), .S(n1065), .CO(n1064));
Q_AD01HF U1421 ( .A0(gfifoGBfullCnt[47]), .B0(n1068), .S(n1067), .CO(n1066));
Q_AD01HF U1422 ( .A0(gfifoGBfullCnt[46]), .B0(n1070), .S(n1069), .CO(n1068));
Q_AD01HF U1423 ( .A0(gfifoGBfullCnt[45]), .B0(n1072), .S(n1071), .CO(n1070));
Q_AD01HF U1424 ( .A0(gfifoGBfullCnt[44]), .B0(n1074), .S(n1073), .CO(n1072));
Q_AD01HF U1425 ( .A0(gfifoGBfullCnt[43]), .B0(n1076), .S(n1075), .CO(n1074));
Q_AD01HF U1426 ( .A0(gfifoGBfullCnt[42]), .B0(n1078), .S(n1077), .CO(n1076));
Q_AD01HF U1427 ( .A0(gfifoGBfullCnt[41]), .B0(n1080), .S(n1079), .CO(n1078));
Q_AD01HF U1428 ( .A0(gfifoGBfullCnt[40]), .B0(n1082), .S(n1081), .CO(n1080));
Q_AD01HF U1429 ( .A0(gfifoGBfullCnt[39]), .B0(n1084), .S(n1083), .CO(n1082));
Q_AD01HF U1430 ( .A0(gfifoGBfullCnt[38]), .B0(n1086), .S(n1085), .CO(n1084));
Q_AD01HF U1431 ( .A0(gfifoGBfullCnt[37]), .B0(n1088), .S(n1087), .CO(n1086));
Q_AD01HF U1432 ( .A0(gfifoGBfullCnt[36]), .B0(n1090), .S(n1089), .CO(n1088));
Q_AD01HF U1433 ( .A0(gfifoGBfullCnt[35]), .B0(n1092), .S(n1091), .CO(n1090));
Q_AD01HF U1434 ( .A0(gfifoGBfullCnt[34]), .B0(n1094), .S(n1093), .CO(n1092));
Q_AD01HF U1435 ( .A0(gfifoGBfullCnt[33]), .B0(n1096), .S(n1095), .CO(n1094));
Q_AD01HF U1436 ( .A0(gfifoGBfullCnt[32]), .B0(n1098), .S(n1097), .CO(n1096));
Q_AD01HF U1437 ( .A0(gfifoGBfullCnt[31]), .B0(n1100), .S(n1099), .CO(n1098));
Q_AD01HF U1438 ( .A0(gfifoGBfullCnt[30]), .B0(n1102), .S(n1101), .CO(n1100));
Q_AD01HF U1439 ( .A0(gfifoGBfullCnt[29]), .B0(n1104), .S(n1103), .CO(n1102));
Q_AD01HF U1440 ( .A0(gfifoGBfullCnt[28]), .B0(n1106), .S(n1105), .CO(n1104));
Q_AD01HF U1441 ( .A0(gfifoGBfullCnt[27]), .B0(n1108), .S(n1107), .CO(n1106));
Q_AD01HF U1442 ( .A0(gfifoGBfullCnt[26]), .B0(n1110), .S(n1109), .CO(n1108));
Q_AD01HF U1443 ( .A0(gfifoGBfullCnt[25]), .B0(n1112), .S(n1111), .CO(n1110));
Q_AD01HF U1444 ( .A0(gfifoGBfullCnt[24]), .B0(n1114), .S(n1113), .CO(n1112));
Q_AD01HF U1445 ( .A0(gfifoGBfullCnt[23]), .B0(n1116), .S(n1115), .CO(n1114));
Q_AD01HF U1446 ( .A0(gfifoGBfullCnt[22]), .B0(n1118), .S(n1117), .CO(n1116));
Q_AD01HF U1447 ( .A0(gfifoGBfullCnt[21]), .B0(n1120), .S(n1119), .CO(n1118));
Q_AD01HF U1448 ( .A0(gfifoGBfullCnt[20]), .B0(n1122), .S(n1121), .CO(n1120));
Q_AD01HF U1449 ( .A0(gfifoGBfullCnt[19]), .B0(n1124), .S(n1123), .CO(n1122));
Q_AD01HF U1450 ( .A0(gfifoGBfullCnt[18]), .B0(n1126), .S(n1125), .CO(n1124));
Q_AD01HF U1451 ( .A0(gfifoGBfullCnt[17]), .B0(n1128), .S(n1127), .CO(n1126));
Q_AD01HF U1452 ( .A0(gfifoGBfullCnt[16]), .B0(n1130), .S(n1129), .CO(n1128));
Q_AD01HF U1453 ( .A0(gfifoGBfullCnt[15]), .B0(n1132), .S(n1131), .CO(n1130));
Q_AD01HF U1454 ( .A0(gfifoGBfullCnt[14]), .B0(n1134), .S(n1133), .CO(n1132));
Q_AD01HF U1455 ( .A0(gfifoGBfullCnt[13]), .B0(n1136), .S(n1135), .CO(n1134));
Q_AD01HF U1456 ( .A0(gfifoGBfullCnt[12]), .B0(n1138), .S(n1137), .CO(n1136));
Q_AD01HF U1457 ( .A0(gfifoGBfullCnt[11]), .B0(n1140), .S(n1139), .CO(n1138));
Q_AD01HF U1458 ( .A0(gfifoGBfullCnt[10]), .B0(n1142), .S(n1141), .CO(n1140));
Q_AD01HF U1459 ( .A0(gfifoGBfullCnt[9]), .B0(n1144), .S(n1143), .CO(n1142));
Q_AD01HF U1460 ( .A0(gfifoGBfullCnt[8]), .B0(n1146), .S(n1145), .CO(n1144));
Q_AD01HF U1461 ( .A0(gfifoGBfullCnt[7]), .B0(n1148), .S(n1147), .CO(n1146));
Q_AD01HF U1462 ( .A0(gfifoGBfullCnt[6]), .B0(n1150), .S(n1149), .CO(n1148));
Q_AD01HF U1463 ( .A0(gfifoGBfullCnt[5]), .B0(n1152), .S(n1151), .CO(n1150));
Q_AD01HF U1464 ( .A0(gfifoGBfullCnt[4]), .B0(n1154), .S(n1153), .CO(n1152));
Q_AD01HF U1465 ( .A0(gfifoGBfullCnt[3]), .B0(n1156), .S(n1155), .CO(n1154));
Q_AD01HF U1466 ( .A0(gfifoGBfullCnt[2]), .B0(n1158), .S(n1157), .CO(n1156));
Q_AD01HF U1467 ( .A0(gfifoGBfullCnt[1]), .B0(gfifoGBfullCnt[0]), .S(n1159), .CO(n1158));
Q_INV U1468 ( .A(sdlHaltHwClk), .Z(n1161));
Q_INV U1469 ( .A(sdlStop), .Z(n1160));
Q_AO21 U1470 ( .A0(sdlHaltHwClkR), .A1(n1160), .B0(n1161), .Z(n1163));
Q_INV U1471 ( .A(callEmu), .Z(n1162));
Q_NR02 U1472 ( .A0(callEmu), .A1(evalOnC), .Z(n1165));
Q_AN02 U1473 ( .A0(n1165), .A1(n1163), .Z(n1164));
Q_MX02 U1474 ( .S(n1164), .A0(n1167), .A1(hwClkHalt), .Z(n1166));
Q_FDP0UA U1475 ( .D(n1166), .QTFCLK( ), .Q(hwClkHalt));
Q_AO21 U1476 ( .A0(sdlStop), .A1(sdlHaltHwClk), .B0(n1165), .Z(n1167));
Q_FDP0UA U1477 ( .D(sdlHaltHwClk), .QTFCLK( ), .Q(sdlHaltHwClkR));
Q_MX02 U1478 ( .S(hwClkDbgOn), .A0(hwClkDelay[0]), .A1(n1406), .Z(n1168));
Q_FDP0UA U1479 ( .D(n1168), .QTFCLK( ), .Q(hwClkDelay[0]));
Q_MX02 U1480 ( .S(hwClkDbgOn), .A0(hwClkDelay[1]), .A1(n1405), .Z(n1169));
Q_FDP0UA U1481 ( .D(n1169), .QTFCLK( ), .Q(hwClkDelay[1]));
Q_MX02 U1482 ( .S(hwClkDbgOn), .A0(hwClkDelay[2]), .A1(n1404), .Z(n1170));
Q_FDP0UA U1483 ( .D(n1170), .QTFCLK( ), .Q(hwClkDelay[2]));
Q_MX02 U1484 ( .S(hwClkDbgOn), .A0(hwClkDelay[3]), .A1(n1403), .Z(n1171));
Q_FDP0UA U1485 ( .D(n1171), .QTFCLK( ), .Q(hwClkDelay[3]));
Q_MX02 U1486 ( .S(hwClkDbgOn), .A0(hwClkDelay[4]), .A1(n1402), .Z(n1172));
Q_FDP0UA U1487 ( .D(n1172), .QTFCLK( ), .Q(hwClkDelay[4]));
Q_MX02 U1488 ( .S(hwClkDbgOn), .A0(hwClkDelay[5]), .A1(n1401), .Z(n1173));
Q_FDP0UA U1489 ( .D(n1173), .QTFCLK( ), .Q(hwClkDelay[5]));
Q_MX02 U1490 ( .S(hwClkDbgOn), .A0(hwClkDelay[6]), .A1(n1400), .Z(n1174));
Q_FDP0UA U1491 ( .D(n1174), .QTFCLK( ), .Q(hwClkDelay[6]));
Q_MX02 U1492 ( .S(hwClkDbgOn), .A0(hwClkDelay[7]), .A1(n1399), .Z(n1175));
Q_FDP0UA U1493 ( .D(n1175), .QTFCLK( ), .Q(hwClkDelay[7]));
Q_MX02 U1494 ( .S(hwClkDbgOn), .A0(hwClkDelay[8]), .A1(n1398), .Z(n1176));
Q_FDP0UA U1495 ( .D(n1176), .QTFCLK( ), .Q(hwClkDelay[8]));
Q_MX02 U1496 ( .S(hwClkDbgOn), .A0(hwClkDelay[9]), .A1(n1397), .Z(n1177));
Q_FDP0UA U1497 ( .D(n1177), .QTFCLK( ), .Q(hwClkDelay[9]));
Q_MX02 U1498 ( .S(hwClkDbgOn), .A0(hwClkDelay[10]), .A1(n1396), .Z(n1178));
Q_FDP0UA U1499 ( .D(n1178), .QTFCLK( ), .Q(hwClkDelay[10]));
Q_MX02 U1500 ( .S(hwClkDbgOn), .A0(hwClkDelay[11]), .A1(n1395), .Z(n1179));
Q_FDP0UA U1501 ( .D(n1179), .QTFCLK( ), .Q(hwClkDelay[11]));
Q_MX02 U1502 ( .S(hwClkDbgOn), .A0(hwClkDelay[12]), .A1(n1394), .Z(n1180));
Q_FDP0UA U1503 ( .D(n1180), .QTFCLK( ), .Q(hwClkDelay[12]));
Q_MX02 U1504 ( .S(hwClkDbgOn), .A0(hwClkDelay[13]), .A1(n1393), .Z(n1181));
Q_FDP0UA U1505 ( .D(n1181), .QTFCLK( ), .Q(hwClkDelay[13]));
Q_MX02 U1506 ( .S(hwClkDbgOn), .A0(hwClkDelay[14]), .A1(n1392), .Z(n1182));
Q_FDP0UA U1507 ( .D(n1182), .QTFCLK( ), .Q(hwClkDelay[14]));
Q_MX02 U1508 ( .S(hwClkDbgOn), .A0(hwClkDelay[15]), .A1(n1391), .Z(n1183));
Q_FDP0UA U1509 ( .D(n1183), .QTFCLK( ), .Q(hwClkDelay[15]));
Q_MX02 U1510 ( .S(hwClkDbgOn), .A0(hwClkDelay[16]), .A1(n1390), .Z(n1184));
Q_FDP0UA U1511 ( .D(n1184), .QTFCLK( ), .Q(hwClkDelay[16]));
Q_MX02 U1512 ( .S(hwClkDbgOn), .A0(hwClkDelay[17]), .A1(n1389), .Z(n1185));
Q_FDP0UA U1513 ( .D(n1185), .QTFCLK( ), .Q(hwClkDelay[17]));
Q_MX02 U1514 ( .S(hwClkDbgOn), .A0(hwClkDelay[18]), .A1(n1388), .Z(n1186));
Q_FDP0UA U1515 ( .D(n1186), .QTFCLK( ), .Q(hwClkDelay[18]));
Q_MX02 U1516 ( .S(hwClkDbgOn), .A0(hwClkDelay[19]), .A1(n1387), .Z(n1187));
Q_FDP0UA U1517 ( .D(n1187), .QTFCLK( ), .Q(hwClkDelay[19]));
Q_MX02 U1518 ( .S(hwClkDbgOn), .A0(hwClkDelay[20]), .A1(n1386), .Z(n1188));
Q_FDP0UA U1519 ( .D(n1188), .QTFCLK( ), .Q(hwClkDelay[20]));
Q_MX02 U1520 ( .S(hwClkDbgOn), .A0(hwClkDelay[21]), .A1(n1385), .Z(n1189));
Q_FDP0UA U1521 ( .D(n1189), .QTFCLK( ), .Q(hwClkDelay[21]));
Q_MX02 U1522 ( .S(hwClkDbgOn), .A0(hwClkDelay[22]), .A1(n1384), .Z(n1190));
Q_FDP0UA U1523 ( .D(n1190), .QTFCLK( ), .Q(hwClkDelay[22]));
Q_MX02 U1524 ( .S(hwClkDbgOn), .A0(hwClkDelay[23]), .A1(n1383), .Z(n1191));
Q_FDP0UA U1525 ( .D(n1191), .QTFCLK( ), .Q(hwClkDelay[23]));
Q_MX02 U1526 ( .S(hwClkDbgOn), .A0(hwClkDelay[24]), .A1(n1382), .Z(n1192));
Q_FDP0UA U1527 ( .D(n1192), .QTFCLK( ), .Q(hwClkDelay[24]));
Q_MX02 U1528 ( .S(hwClkDbgOn), .A0(hwClkDelay[25]), .A1(n1381), .Z(n1193));
Q_FDP0UA U1529 ( .D(n1193), .QTFCLK( ), .Q(hwClkDelay[25]));
Q_MX02 U1530 ( .S(hwClkDbgOn), .A0(hwClkDelay[26]), .A1(n1380), .Z(n1194));
Q_FDP0UA U1531 ( .D(n1194), .QTFCLK( ), .Q(hwClkDelay[26]));
Q_MX02 U1532 ( .S(hwClkDbgOn), .A0(hwClkDelay[27]), .A1(n1379), .Z(n1195));
Q_FDP0UA U1533 ( .D(n1195), .QTFCLK( ), .Q(hwClkDelay[27]));
Q_MX02 U1534 ( .S(hwClkDbgOn), .A0(hwClkDelay[28]), .A1(n1378), .Z(n1196));
Q_FDP0UA U1535 ( .D(n1196), .QTFCLK( ), .Q(hwClkDelay[28]));
Q_MX02 U1536 ( .S(hwClkDbgOn), .A0(hwClkDelay[29]), .A1(n1377), .Z(n1197));
Q_FDP0UA U1537 ( .D(n1197), .QTFCLK( ), .Q(hwClkDelay[29]));
Q_MX02 U1538 ( .S(hwClkDbgOn), .A0(hwClkDelay[30]), .A1(n1376), .Z(n1198));
Q_FDP0UA U1539 ( .D(n1198), .QTFCLK( ), .Q(hwClkDelay[30]));
Q_MX02 U1540 ( .S(hwClkDbgOn), .A0(hwClkDelay[31]), .A1(n1375), .Z(n1199));
Q_FDP0UA U1541 ( .D(n1199), .QTFCLK( ), .Q(hwClkDelay[31]));
Q_MX02 U1542 ( .S(hwClkDbgOn), .A0(hwSimTime[0]), .A1(n1374), .Z(n1200));
Q_FDP0UA U1543 ( .D(n1200), .QTFCLK( ), .Q(hwSimTime[0]));
Q_MX02 U1544 ( .S(hwClkDbgOn), .A0(hwSimTime[1]), .A1(n1372), .Z(n1201));
Q_FDP0UA U1545 ( .D(n1201), .QTFCLK( ), .Q(hwSimTime[1]));
Q_MX02 U1546 ( .S(hwClkDbgOn), .A0(hwSimTime[2]), .A1(n1370), .Z(n1202));
Q_FDP0UA U1547 ( .D(n1202), .QTFCLK( ), .Q(hwSimTime[2]));
Q_MX02 U1548 ( .S(hwClkDbgOn), .A0(hwSimTime[3]), .A1(n1369), .Z(n1203));
Q_FDP0UA U1549 ( .D(n1203), .QTFCLK( ), .Q(hwSimTime[3]));
Q_MX02 U1550 ( .S(hwClkDbgOn), .A0(hwSimTime[4]), .A1(n1367), .Z(n1204));
Q_FDP0UA U1551 ( .D(n1204), .QTFCLK( ), .Q(hwSimTime[4]));
Q_MX02 U1552 ( .S(hwClkDbgOn), .A0(hwSimTime[5]), .A1(n1366), .Z(n1205));
Q_FDP0UA U1553 ( .D(n1205), .QTFCLK( ), .Q(hwSimTime[5]));
Q_MX02 U1554 ( .S(hwClkDbgOn), .A0(hwSimTime[6]), .A1(n1364), .Z(n1206));
Q_FDP0UA U1555 ( .D(n1206), .QTFCLK( ), .Q(hwSimTime[6]));
Q_MX02 U1556 ( .S(hwClkDbgOn), .A0(hwSimTime[7]), .A1(n1363), .Z(n1207));
Q_FDP0UA U1557 ( .D(n1207), .QTFCLK( ), .Q(hwSimTime[7]));
Q_MX02 U1558 ( .S(hwClkDbgOn), .A0(hwSimTime[8]), .A1(n1361), .Z(n1208));
Q_FDP0UA U1559 ( .D(n1208), .QTFCLK( ), .Q(hwSimTime[8]));
Q_MX02 U1560 ( .S(hwClkDbgOn), .A0(hwSimTime[9]), .A1(n1360), .Z(n1209));
Q_FDP0UA U1561 ( .D(n1209), .QTFCLK( ), .Q(hwSimTime[9]));
Q_MX02 U1562 ( .S(hwClkDbgOn), .A0(hwSimTime[10]), .A1(n1358), .Z(n1210));
Q_FDP0UA U1563 ( .D(n1210), .QTFCLK( ), .Q(hwSimTime[10]));
Q_MX02 U1564 ( .S(hwClkDbgOn), .A0(hwSimTime[11]), .A1(n1357), .Z(n1211));
Q_FDP0UA U1565 ( .D(n1211), .QTFCLK( ), .Q(hwSimTime[11]));
Q_MX02 U1566 ( .S(hwClkDbgOn), .A0(hwSimTime[12]), .A1(n1355), .Z(n1212));
Q_FDP0UA U1567 ( .D(n1212), .QTFCLK( ), .Q(hwSimTime[12]));
Q_MX02 U1568 ( .S(hwClkDbgOn), .A0(hwSimTime[13]), .A1(n1354), .Z(n1213));
Q_FDP0UA U1569 ( .D(n1213), .QTFCLK( ), .Q(hwSimTime[13]));
Q_MX02 U1570 ( .S(hwClkDbgOn), .A0(hwSimTime[14]), .A1(n1352), .Z(n1214));
Q_FDP0UA U1571 ( .D(n1214), .QTFCLK( ), .Q(hwSimTime[14]));
Q_MX02 U1572 ( .S(hwClkDbgOn), .A0(hwSimTime[15]), .A1(n1351), .Z(n1215));
Q_FDP0UA U1573 ( .D(n1215), .QTFCLK( ), .Q(hwSimTime[15]));
Q_MX02 U1574 ( .S(hwClkDbgOn), .A0(hwSimTime[16]), .A1(n1349), .Z(n1216));
Q_FDP0UA U1575 ( .D(n1216), .QTFCLK( ), .Q(hwSimTime[16]));
Q_MX02 U1576 ( .S(hwClkDbgOn), .A0(hwSimTime[17]), .A1(n1348), .Z(n1217));
Q_FDP0UA U1577 ( .D(n1217), .QTFCLK( ), .Q(hwSimTime[17]));
Q_MX02 U1578 ( .S(hwClkDbgOn), .A0(hwSimTime[18]), .A1(n1346), .Z(n1218));
Q_FDP0UA U1579 ( .D(n1218), .QTFCLK( ), .Q(hwSimTime[18]));
Q_MX02 U1580 ( .S(hwClkDbgOn), .A0(hwSimTime[19]), .A1(n1345), .Z(n1219));
Q_FDP0UA U1581 ( .D(n1219), .QTFCLK( ), .Q(hwSimTime[19]));
Q_MX02 U1582 ( .S(hwClkDbgOn), .A0(hwSimTime[20]), .A1(n1343), .Z(n1220));
Q_FDP0UA U1583 ( .D(n1220), .QTFCLK( ), .Q(hwSimTime[20]));
Q_MX02 U1584 ( .S(hwClkDbgOn), .A0(hwSimTime[21]), .A1(n1342), .Z(n1221));
Q_FDP0UA U1585 ( .D(n1221), .QTFCLK( ), .Q(hwSimTime[21]));
Q_MX02 U1586 ( .S(hwClkDbgOn), .A0(hwSimTime[22]), .A1(n1340), .Z(n1222));
Q_FDP0UA U1587 ( .D(n1222), .QTFCLK( ), .Q(hwSimTime[22]));
Q_MX02 U1588 ( .S(hwClkDbgOn), .A0(hwSimTime[23]), .A1(n1339), .Z(n1223));
Q_FDP0UA U1589 ( .D(n1223), .QTFCLK( ), .Q(hwSimTime[23]));
Q_MX02 U1590 ( .S(hwClkDbgOn), .A0(hwSimTime[24]), .A1(n1337), .Z(n1224));
Q_FDP0UA U1591 ( .D(n1224), .QTFCLK( ), .Q(hwSimTime[24]));
Q_MX02 U1592 ( .S(hwClkDbgOn), .A0(hwSimTime[25]), .A1(n1336), .Z(n1225));
Q_FDP0UA U1593 ( .D(n1225), .QTFCLK( ), .Q(hwSimTime[25]));
Q_MX02 U1594 ( .S(hwClkDbgOn), .A0(hwSimTime[26]), .A1(n1334), .Z(n1226));
Q_FDP0UA U1595 ( .D(n1226), .QTFCLK( ), .Q(hwSimTime[26]));
Q_MX02 U1596 ( .S(hwClkDbgOn), .A0(hwSimTime[27]), .A1(n1333), .Z(n1227));
Q_FDP0UA U1597 ( .D(n1227), .QTFCLK( ), .Q(hwSimTime[27]));
Q_MX02 U1598 ( .S(hwClkDbgOn), .A0(hwSimTime[28]), .A1(n1331), .Z(n1228));
Q_FDP0UA U1599 ( .D(n1228), .QTFCLK( ), .Q(hwSimTime[28]));
Q_MX02 U1600 ( .S(hwClkDbgOn), .A0(hwSimTime[29]), .A1(n1330), .Z(n1229));
Q_FDP0UA U1601 ( .D(n1229), .QTFCLK( ), .Q(hwSimTime[29]));
Q_MX02 U1602 ( .S(hwClkDbgOn), .A0(hwSimTime[30]), .A1(n1328), .Z(n1230));
Q_FDP0UA U1603 ( .D(n1230), .QTFCLK( ), .Q(hwSimTime[30]));
Q_MX02 U1604 ( .S(hwClkDbgOn), .A0(hwSimTime[31]), .A1(n1327), .Z(n1231));
Q_FDP0UA U1605 ( .D(n1231), .QTFCLK( ), .Q(hwSimTime[31]));
Q_MX02 U1606 ( .S(hwClkDbgOn), .A0(hwSimTime[32]), .A1(n1325), .Z(n1232));
Q_FDP0UA U1607 ( .D(n1232), .QTFCLK( ), .Q(hwSimTime[32]));
Q_MX02 U1608 ( .S(hwClkDbgOn), .A0(hwSimTime[33]), .A1(n1323), .Z(n1233));
Q_FDP0UA U1609 ( .D(n1233), .QTFCLK( ), .Q(hwSimTime[33]));
Q_MX02 U1610 ( .S(hwClkDbgOn), .A0(hwSimTime[34]), .A1(n1321), .Z(n1234));
Q_FDP0UA U1611 ( .D(n1234), .QTFCLK( ), .Q(hwSimTime[34]));
Q_MX02 U1612 ( .S(hwClkDbgOn), .A0(hwSimTime[35]), .A1(n1319), .Z(n1235));
Q_FDP0UA U1613 ( .D(n1235), .QTFCLK( ), .Q(hwSimTime[35]));
Q_MX02 U1614 ( .S(hwClkDbgOn), .A0(hwSimTime[36]), .A1(n1317), .Z(n1236));
Q_FDP0UA U1615 ( .D(n1236), .QTFCLK( ), .Q(hwSimTime[36]));
Q_MX02 U1616 ( .S(hwClkDbgOn), .A0(hwSimTime[37]), .A1(n1315), .Z(n1237));
Q_FDP0UA U1617 ( .D(n1237), .QTFCLK( ), .Q(hwSimTime[37]));
Q_MX02 U1618 ( .S(hwClkDbgOn), .A0(hwSimTime[38]), .A1(n1313), .Z(n1238));
Q_FDP0UA U1619 ( .D(n1238), .QTFCLK( ), .Q(hwSimTime[38]));
Q_MX02 U1620 ( .S(hwClkDbgOn), .A0(hwSimTime[39]), .A1(n1311), .Z(n1239));
Q_FDP0UA U1621 ( .D(n1239), .QTFCLK( ), .Q(hwSimTime[39]));
Q_MX02 U1622 ( .S(hwClkDbgOn), .A0(hwSimTime[40]), .A1(n1309), .Z(n1240));
Q_FDP0UA U1623 ( .D(n1240), .QTFCLK( ), .Q(hwSimTime[40]));
Q_MX02 U1624 ( .S(hwClkDbgOn), .A0(hwSimTime[41]), .A1(n1307), .Z(n1241));
Q_FDP0UA U1625 ( .D(n1241), .QTFCLK( ), .Q(hwSimTime[41]));
Q_MX02 U1626 ( .S(hwClkDbgOn), .A0(hwSimTime[42]), .A1(n1305), .Z(n1242));
Q_FDP0UA U1627 ( .D(n1242), .QTFCLK( ), .Q(hwSimTime[42]));
Q_MX02 U1628 ( .S(hwClkDbgOn), .A0(hwSimTime[43]), .A1(n1303), .Z(n1243));
Q_FDP0UA U1629 ( .D(n1243), .QTFCLK( ), .Q(hwSimTime[43]));
Q_MX02 U1630 ( .S(hwClkDbgOn), .A0(hwSimTime[44]), .A1(n1301), .Z(n1244));
Q_FDP0UA U1631 ( .D(n1244), .QTFCLK( ), .Q(hwSimTime[44]));
Q_MX02 U1632 ( .S(hwClkDbgOn), .A0(hwSimTime[45]), .A1(n1299), .Z(n1245));
Q_FDP0UA U1633 ( .D(n1245), .QTFCLK( ), .Q(hwSimTime[45]));
Q_MX02 U1634 ( .S(hwClkDbgOn), .A0(hwSimTime[46]), .A1(n1297), .Z(n1246));
Q_FDP0UA U1635 ( .D(n1246), .QTFCLK( ), .Q(hwSimTime[46]));
Q_MX02 U1636 ( .S(hwClkDbgOn), .A0(hwSimTime[47]), .A1(n1295), .Z(n1247));
Q_FDP0UA U1637 ( .D(n1247), .QTFCLK( ), .Q(hwSimTime[47]));
Q_MX02 U1638 ( .S(hwClkDbgOn), .A0(hwSimTime[48]), .A1(n1293), .Z(n1248));
Q_FDP0UA U1639 ( .D(n1248), .QTFCLK( ), .Q(hwSimTime[48]));
Q_MX02 U1640 ( .S(hwClkDbgOn), .A0(hwSimTime[49]), .A1(n1291), .Z(n1249));
Q_FDP0UA U1641 ( .D(n1249), .QTFCLK( ), .Q(hwSimTime[49]));
Q_MX02 U1642 ( .S(hwClkDbgOn), .A0(hwSimTime[50]), .A1(n1289), .Z(n1250));
Q_FDP0UA U1643 ( .D(n1250), .QTFCLK( ), .Q(hwSimTime[50]));
Q_MX02 U1644 ( .S(hwClkDbgOn), .A0(hwSimTime[51]), .A1(n1287), .Z(n1251));
Q_FDP0UA U1645 ( .D(n1251), .QTFCLK( ), .Q(hwSimTime[51]));
Q_MX02 U1646 ( .S(hwClkDbgOn), .A0(hwSimTime[52]), .A1(n1285), .Z(n1252));
Q_FDP0UA U1647 ( .D(n1252), .QTFCLK( ), .Q(hwSimTime[52]));
Q_MX02 U1648 ( .S(hwClkDbgOn), .A0(hwSimTime[53]), .A1(n1283), .Z(n1253));
Q_FDP0UA U1649 ( .D(n1253), .QTFCLK( ), .Q(hwSimTime[53]));
Q_MX02 U1650 ( .S(hwClkDbgOn), .A0(hwSimTime[54]), .A1(n1281), .Z(n1254));
Q_FDP0UA U1651 ( .D(n1254), .QTFCLK( ), .Q(hwSimTime[54]));
Q_MX02 U1652 ( .S(hwClkDbgOn), .A0(hwSimTime[55]), .A1(n1279), .Z(n1255));
Q_FDP0UA U1653 ( .D(n1255), .QTFCLK( ), .Q(hwSimTime[55]));
Q_MX02 U1654 ( .S(hwClkDbgOn), .A0(hwSimTime[56]), .A1(n1277), .Z(n1256));
Q_FDP0UA U1655 ( .D(n1256), .QTFCLK( ), .Q(hwSimTime[56]));
Q_MX02 U1656 ( .S(hwClkDbgOn), .A0(hwSimTime[57]), .A1(n1275), .Z(n1257));
Q_FDP0UA U1657 ( .D(n1257), .QTFCLK( ), .Q(hwSimTime[57]));
Q_MX02 U1658 ( .S(hwClkDbgOn), .A0(hwSimTime[58]), .A1(n1273), .Z(n1258));
Q_FDP0UA U1659 ( .D(n1258), .QTFCLK( ), .Q(hwSimTime[58]));
Q_MX02 U1660 ( .S(hwClkDbgOn), .A0(hwSimTime[59]), .A1(n1271), .Z(n1259));
Q_FDP0UA U1661 ( .D(n1259), .QTFCLK( ), .Q(hwSimTime[59]));
Q_MX02 U1662 ( .S(hwClkDbgOn), .A0(hwSimTime[60]), .A1(n1269), .Z(n1260));
Q_FDP0UA U1663 ( .D(n1260), .QTFCLK( ), .Q(hwSimTime[60]));
Q_MX02 U1664 ( .S(hwClkDbgOn), .A0(hwSimTime[61]), .A1(n1267), .Z(n1261));
Q_FDP0UA U1665 ( .D(n1261), .QTFCLK( ), .Q(hwSimTime[61]));
Q_MX02 U1666 ( .S(hwClkDbgOn), .A0(hwSimTime[62]), .A1(n1265), .Z(n1262));
Q_FDP0UA U1667 ( .D(n1262), .QTFCLK( ), .Q(hwSimTime[62]));
Q_FDP0UA U1668 ( .D(n1263), .QTFCLK( ), .Q(hwSimTime[63]));
Q_XOR2 U1669 ( .A0(hwSimTime[63]), .A1(n10), .Z(n1263));
Q_AD01HF U1670 ( .A0(hwSimTime[62]), .B0(n1266), .S(n1265), .CO(n1264));
Q_AD01HF U1671 ( .A0(hwSimTime[61]), .B0(n1268), .S(n1267), .CO(n1266));
Q_AD01HF U1672 ( .A0(hwSimTime[60]), .B0(n1270), .S(n1269), .CO(n1268));
Q_AD01HF U1673 ( .A0(hwSimTime[59]), .B0(n1272), .S(n1271), .CO(n1270));
Q_AD01HF U1674 ( .A0(hwSimTime[58]), .B0(n1274), .S(n1273), .CO(n1272));
Q_AD01HF U1675 ( .A0(hwSimTime[57]), .B0(n1276), .S(n1275), .CO(n1274));
Q_AD01HF U1676 ( .A0(hwSimTime[56]), .B0(n1278), .S(n1277), .CO(n1276));
Q_AD01HF U1677 ( .A0(hwSimTime[55]), .B0(n1280), .S(n1279), .CO(n1278));
Q_AD01HF U1678 ( .A0(hwSimTime[54]), .B0(n1282), .S(n1281), .CO(n1280));
Q_AD01HF U1679 ( .A0(hwSimTime[53]), .B0(n1284), .S(n1283), .CO(n1282));
Q_AD01HF U1680 ( .A0(hwSimTime[52]), .B0(n1286), .S(n1285), .CO(n1284));
Q_AD01HF U1681 ( .A0(hwSimTime[51]), .B0(n1288), .S(n1287), .CO(n1286));
Q_AD01HF U1682 ( .A0(hwSimTime[50]), .B0(n1290), .S(n1289), .CO(n1288));
Q_AD01HF U1683 ( .A0(hwSimTime[49]), .B0(n1292), .S(n1291), .CO(n1290));
Q_AD01HF U1684 ( .A0(hwSimTime[48]), .B0(n1294), .S(n1293), .CO(n1292));
Q_AD01HF U1685 ( .A0(hwSimTime[47]), .B0(n1296), .S(n1295), .CO(n1294));
Q_AD01HF U1686 ( .A0(hwSimTime[46]), .B0(n1298), .S(n1297), .CO(n1296));
Q_AD01HF U1687 ( .A0(hwSimTime[45]), .B0(n1300), .S(n1299), .CO(n1298));
Q_AD01HF U1688 ( .A0(hwSimTime[44]), .B0(n1302), .S(n1301), .CO(n1300));
Q_AD01HF U1689 ( .A0(hwSimTime[43]), .B0(n1304), .S(n1303), .CO(n1302));
Q_AD01HF U1690 ( .A0(hwSimTime[42]), .B0(n1306), .S(n1305), .CO(n1304));
Q_AD01HF U1691 ( .A0(hwSimTime[41]), .B0(n1308), .S(n1307), .CO(n1306));
Q_AD01HF U1692 ( .A0(hwSimTime[40]), .B0(n1310), .S(n1309), .CO(n1308));
Q_AD01HF U1693 ( .A0(hwSimTime[39]), .B0(n1312), .S(n1311), .CO(n1310));
Q_AD01HF U1694 ( .A0(hwSimTime[38]), .B0(n1314), .S(n1313), .CO(n1312));
Q_AD01HF U1695 ( .A0(hwSimTime[37]), .B0(n1316), .S(n1315), .CO(n1314));
Q_AD01HF U1696 ( .A0(hwSimTime[36]), .B0(n1318), .S(n1317), .CO(n1316));
Q_AD01HF U1697 ( .A0(hwSimTime[35]), .B0(n1320), .S(n1319), .CO(n1318));
Q_AD01HF U1698 ( .A0(hwSimTime[34]), .B0(n1322), .S(n1321), .CO(n1320));
Q_AD01HF U1699 ( .A0(hwSimTime[33]), .B0(n1324), .S(n1323), .CO(n1322));
Q_AD01HF U1700 ( .A0(hwSimTime[32]), .B0(n1326), .S(n1325), .CO(n1324));
Q_AD02 U1701 ( .CI(n1329), .A0(hwSimTime[30]), .A1(hwSimTime[31]), .B0(n1376), .B1(n1375), .S0(n1328), .S1(n1327), .CO(n1326));
Q_AD02 U1702 ( .CI(n1332), .A0(hwSimTime[28]), .A1(hwSimTime[29]), .B0(n1378), .B1(n1377), .S0(n1331), .S1(n1330), .CO(n1329));
Q_AD02 U1703 ( .CI(n1335), .A0(hwSimTime[26]), .A1(hwSimTime[27]), .B0(n1380), .B1(n1379), .S0(n1334), .S1(n1333), .CO(n1332));
Q_AD02 U1704 ( .CI(n1338), .A0(hwSimTime[24]), .A1(hwSimTime[25]), .B0(n1382), .B1(n1381), .S0(n1337), .S1(n1336), .CO(n1335));
Q_AD02 U1705 ( .CI(n1341), .A0(hwSimTime[22]), .A1(hwSimTime[23]), .B0(n1384), .B1(n1383), .S0(n1340), .S1(n1339), .CO(n1338));
Q_AD02 U1706 ( .CI(n1344), .A0(hwSimTime[20]), .A1(hwSimTime[21]), .B0(n1386), .B1(n1385), .S0(n1343), .S1(n1342), .CO(n1341));
Q_AD02 U1707 ( .CI(n1347), .A0(hwSimTime[18]), .A1(hwSimTime[19]), .B0(n1388), .B1(n1387), .S0(n1346), .S1(n1345), .CO(n1344));
Q_AD02 U1708 ( .CI(n1350), .A0(hwSimTime[16]), .A1(hwSimTime[17]), .B0(n1390), .B1(n1389), .S0(n1349), .S1(n1348), .CO(n1347));
Q_AD02 U1709 ( .CI(n1353), .A0(hwSimTime[14]), .A1(hwSimTime[15]), .B0(n1392), .B1(n1391), .S0(n1352), .S1(n1351), .CO(n1350));
Q_AD02 U1710 ( .CI(n1356), .A0(hwSimTime[12]), .A1(hwSimTime[13]), .B0(n1394), .B1(n1393), .S0(n1355), .S1(n1354), .CO(n1353));
Q_AD02 U1711 ( .CI(n1359), .A0(hwSimTime[10]), .A1(hwSimTime[11]), .B0(n1396), .B1(n1395), .S0(n1358), .S1(n1357), .CO(n1356));
Q_AD02 U1712 ( .CI(n1362), .A0(hwSimTime[8]), .A1(hwSimTime[9]), .B0(n1398), .B1(n1397), .S0(n1361), .S1(n1360), .CO(n1359));
Q_AD02 U1713 ( .CI(n1365), .A0(hwSimTime[6]), .A1(hwSimTime[7]), .B0(n1400), .B1(n1399), .S0(n1364), .S1(n1363), .CO(n1362));
Q_AD02 U1714 ( .CI(n1368), .A0(hwSimTime[4]), .A1(hwSimTime[5]), .B0(n1402), .B1(n1401), .S0(n1367), .S1(n1366), .CO(n1365));
Q_AD02 U1715 ( .CI(n1371), .A0(hwSimTime[2]), .A1(hwSimTime[3]), .B0(n1404), .B1(n1403), .S0(n1370), .S1(n1369), .CO(n1368));
Q_AD01 U1716 ( .CI(n1405), .A0(hwSimTime[1]), .B0(n1373), .S(n1372), .CO(n1371));
Q_AD01HF U1717 ( .A0(hwSimTime[0]), .B0(n1406), .S(n1374), .CO(n1373));
Q_AN02 U1718 ( .A0(n1408), .A1(hwClkDelay[31]), .Z(n1375));
Q_AN02 U1719 ( .A0(n1408), .A1(hwClkDelay[30]), .Z(n1376));
Q_AN02 U1720 ( .A0(n1408), .A1(hwClkDelay[29]), .Z(n1377));
Q_AN02 U1721 ( .A0(n1408), .A1(hwClkDelay[28]), .Z(n1378));
Q_AN02 U1722 ( .A0(n1408), .A1(hwClkDelay[27]), .Z(n1379));
Q_AN02 U1723 ( .A0(n1408), .A1(hwClkDelay[26]), .Z(n1380));
Q_AN02 U1724 ( .A0(n1408), .A1(hwClkDelay[25]), .Z(n1381));
Q_AN02 U1725 ( .A0(n1408), .A1(hwClkDelay[24]), .Z(n1382));
Q_AN02 U1726 ( .A0(n1408), .A1(hwClkDelay[23]), .Z(n1383));
Q_AN02 U1727 ( .A0(n1408), .A1(hwClkDelay[22]), .Z(n1384));
Q_AN02 U1728 ( .A0(n1408), .A1(hwClkDelay[21]), .Z(n1385));
Q_AN02 U1729 ( .A0(n1408), .A1(hwClkDelay[20]), .Z(n1386));
Q_AN02 U1730 ( .A0(n1408), .A1(hwClkDelay[19]), .Z(n1387));
Q_AN02 U1731 ( .A0(n1408), .A1(hwClkDelay[18]), .Z(n1388));
Q_AN02 U1732 ( .A0(n1408), .A1(hwClkDelay[17]), .Z(n1389));
Q_AN02 U1733 ( .A0(n1408), .A1(hwClkDelay[16]), .Z(n1390));
Q_AN02 U1734 ( .A0(n1408), .A1(hwClkDelay[15]), .Z(n1391));
Q_AN02 U1735 ( .A0(n1408), .A1(hwClkDelay[14]), .Z(n1392));
Q_AN02 U1736 ( .A0(n1408), .A1(hwClkDelay[13]), .Z(n1393));
Q_AN02 U1737 ( .A0(n1408), .A1(hwClkDelay[12]), .Z(n1394));
Q_AN02 U1738 ( .A0(n1408), .A1(hwClkDelay[11]), .Z(n1395));
Q_AN02 U1739 ( .A0(n1408), .A1(hwClkDelay[10]), .Z(n1396));
Q_AN02 U1740 ( .A0(n1408), .A1(hwClkDelay[9]), .Z(n1397));
Q_AN02 U1741 ( .A0(n1408), .A1(hwClkDelay[8]), .Z(n1398));
Q_AN02 U1742 ( .A0(n1408), .A1(hwClkDelay[7]), .Z(n1399));
Q_AN02 U1743 ( .A0(n1408), .A1(hwClkDelay[6]), .Z(n1400));
Q_AN02 U1744 ( .A0(n1408), .A1(hwClkDelay[5]), .Z(n1401));
Q_AN02 U1745 ( .A0(n1408), .A1(hwClkDelay[4]), .Z(n1402));
Q_AN02 U1746 ( .A0(n1408), .A1(hwClkDelay[3]), .Z(n1403));
Q_AN02 U1747 ( .A0(n1408), .A1(hwClkDelay[2]), .Z(n1404));
Q_AN02 U1748 ( .A0(n1408), .A1(hwClkDelay[1]), .Z(n1405));
Q_OR02 U1749 ( .A0(n1407), .A1(hwClkDelay[0]), .Z(n1406));
Q_INV U1750 ( .A(n1408), .Z(n1407));
Q_OR02 U1751 ( .A0(n1410), .A1(n1409), .Z(n1408));
Q_OR03 U1752 ( .A0(n1413), .A1(n1412), .A2(n1411), .Z(n1409));
Q_OR03 U1753 ( .A0(n1416), .A1(n1415), .A2(n1414), .Z(n1410));
Q_OR03 U1754 ( .A0(n1419), .A1(n1418), .A2(n1417), .Z(n1411));
Q_OR03 U1755 ( .A0(n1422), .A1(n1421), .A2(n1420), .Z(n1412));
Q_OR03 U1756 ( .A0(hwClkDelay[1]), .A1(hwClkDelay[0]), .A2(n1423), .Z(n1413));
Q_OR03 U1757 ( .A0(hwClkDelay[4]), .A1(hwClkDelay[3]), .A2(hwClkDelay[2]), .Z(n1414));
Q_OR03 U1758 ( .A0(hwClkDelay[7]), .A1(hwClkDelay[6]), .A2(hwClkDelay[5]), .Z(n1415));
Q_OR03 U1759 ( .A0(hwClkDelay[10]), .A1(hwClkDelay[9]), .A2(hwClkDelay[8]), .Z(n1416));
Q_OR03 U1760 ( .A0(hwClkDelay[13]), .A1(hwClkDelay[12]), .A2(hwClkDelay[11]), .Z(n1417));
Q_OR03 U1761 ( .A0(hwClkDelay[16]), .A1(hwClkDelay[15]), .A2(hwClkDelay[14]), .Z(n1418));
Q_OR03 U1762 ( .A0(hwClkDelay[19]), .A1(hwClkDelay[18]), .A2(hwClkDelay[17]), .Z(n1419));
Q_OR03 U1763 ( .A0(hwClkDelay[22]), .A1(hwClkDelay[21]), .A2(hwClkDelay[20]), .Z(n1420));
Q_OR03 U1764 ( .A0(hwClkDelay[25]), .A1(hwClkDelay[24]), .A2(hwClkDelay[23]), .Z(n1421));
Q_OR03 U1765 ( .A0(hwClkDelay[28]), .A1(hwClkDelay[27]), .A2(hwClkDelay[26]), .Z(n1422));
Q_OR03 U1766 ( .A0(hwClkDelay[31]), .A1(hwClkDelay[30]), .A2(hwClkDelay[29]), .Z(n1423));
Q_AO21 U1767 ( .A0(ckgHoldPIi), .A1(oneStepPIi), .B0(n1162), .Z(n1425));
Q_INV U1768 ( .A(n1425), .Z(n1424));
Q_OR02 U1769 ( .A0(n1424), .A1(hwClkEnable), .Z(n1426));
Q_FDP0UA U1770 ( .D(n1426), .QTFCLK( ), .Q(hwClkEnable));
Q_FDP0UA U1771 ( .D(dummyW), .QTFCLK( ), .Q(dummyR));
Q_FDP0UA U1772 ( .D(it_capture), .QTFCLK( ), .Q(it_capture));
Q_FDP0UA U1773 ( .D(it_replay), .QTFCLK( ), .Q(it_replay));
Q_INV U1774 ( .A(acHalt), .Z(n1428));
Q_AN02 U1775 ( .A0(asyncCall), .A1(n1428), .Z(n1429));
Q_AN02 U1776 ( .A0(n1429), .A1(n402), .Z(n1427));
Q_XOR2 U1777 ( .A0(n1427), .A1(aCount[0]), .Z(n1430));
Q_FDP0UA U1778 ( .D(n1430), .QTFCLK( ), .Q(aCount[0]));
Q_MX02 U1779 ( .S(n1427), .A0(aCount[1]), .A1(n1521), .Z(n1431));
Q_FDP0UA U1780 ( .D(n1431), .QTFCLK( ), .Q(aCount[1]));
Q_MX02 U1781 ( .S(n1427), .A0(aCount[2]), .A1(n1519), .Z(n1432));
Q_FDP0UA U1782 ( .D(n1432), .QTFCLK( ), .Q(aCount[2]));
Q_MX02 U1783 ( .S(n1427), .A0(aCount[3]), .A1(n1517), .Z(n1433));
Q_FDP0UA U1784 ( .D(n1433), .QTFCLK( ), .Q(aCount[3]));
Q_MX02 U1785 ( .S(n1427), .A0(aCount[4]), .A1(n1515), .Z(n1434));
Q_FDP0UA U1786 ( .D(n1434), .QTFCLK( ), .Q(aCount[4]));
Q_MX02 U1787 ( .S(n1427), .A0(aCount[5]), .A1(n1513), .Z(n1435));
Q_FDP0UA U1788 ( .D(n1435), .QTFCLK( ), .Q(aCount[5]));
Q_MX02 U1789 ( .S(n1427), .A0(aCount[6]), .A1(n1511), .Z(n1436));
Q_FDP0UA U1790 ( .D(n1436), .QTFCLK( ), .Q(aCount[6]));
Q_MX02 U1791 ( .S(n1427), .A0(aCount[7]), .A1(n1509), .Z(n1437));
Q_FDP0UA U1792 ( .D(n1437), .QTFCLK( ), .Q(aCount[7]));
Q_MX02 U1793 ( .S(n1427), .A0(aCount[8]), .A1(n1507), .Z(n1438));
Q_FDP0UA U1794 ( .D(n1438), .QTFCLK( ), .Q(aCount[8]));
Q_MX02 U1795 ( .S(n1427), .A0(aCount[9]), .A1(n1505), .Z(n1439));
Q_FDP0UA U1796 ( .D(n1439), .QTFCLK( ), .Q(aCount[9]));
Q_MX02 U1797 ( .S(n1427), .A0(aCount[10]), .A1(n1503), .Z(n1440));
Q_FDP0UA U1798 ( .D(n1440), .QTFCLK( ), .Q(aCount[10]));
Q_MX02 U1799 ( .S(n1427), .A0(aCount[11]), .A1(n1501), .Z(n1441));
Q_FDP0UA U1800 ( .D(n1441), .QTFCLK( ), .Q(aCount[11]));
Q_MX02 U1801 ( .S(n1427), .A0(aCount[12]), .A1(n1499), .Z(n1442));
Q_FDP0UA U1802 ( .D(n1442), .QTFCLK( ), .Q(aCount[12]));
Q_MX02 U1803 ( .S(n1427), .A0(aCount[13]), .A1(n1497), .Z(n1443));
Q_FDP0UA U1804 ( .D(n1443), .QTFCLK( ), .Q(aCount[13]));
Q_MX02 U1805 ( .S(n1427), .A0(aCount[14]), .A1(n1495), .Z(n1444));
Q_FDP0UA U1806 ( .D(n1444), .QTFCLK( ), .Q(aCount[14]));
Q_MX02 U1807 ( .S(n1427), .A0(aCount[15]), .A1(n1493), .Z(n1445));
Q_FDP0UA U1808 ( .D(n1445), .QTFCLK( ), .Q(aCount[15]));
Q_MX02 U1809 ( .S(n1427), .A0(aCount[16]), .A1(n1491), .Z(n1446));
Q_FDP0UA U1810 ( .D(n1446), .QTFCLK( ), .Q(aCount[16]));
Q_MX02 U1811 ( .S(n1427), .A0(aCount[17]), .A1(n1489), .Z(n1447));
Q_FDP0UA U1812 ( .D(n1447), .QTFCLK( ), .Q(aCount[17]));
Q_MX02 U1813 ( .S(n1427), .A0(aCount[18]), .A1(n1487), .Z(n1448));
Q_FDP0UA U1814 ( .D(n1448), .QTFCLK( ), .Q(aCount[18]));
Q_MX02 U1815 ( .S(n1427), .A0(aCount[19]), .A1(n1485), .Z(n1449));
Q_FDP0UA U1816 ( .D(n1449), .QTFCLK( ), .Q(aCount[19]));
Q_MX02 U1817 ( .S(n1427), .A0(aCount[20]), .A1(n1483), .Z(n1450));
Q_FDP0UA U1818 ( .D(n1450), .QTFCLK( ), .Q(aCount[20]));
Q_MX02 U1819 ( .S(n1427), .A0(aCount[21]), .A1(n1481), .Z(n1451));
Q_FDP0UA U1820 ( .D(n1451), .QTFCLK( ), .Q(aCount[21]));
Q_MX02 U1821 ( .S(n1427), .A0(aCount[22]), .A1(n1479), .Z(n1452));
Q_FDP0UA U1822 ( .D(n1452), .QTFCLK( ), .Q(aCount[22]));
Q_MX02 U1823 ( .S(n1427), .A0(aCount[23]), .A1(n1477), .Z(n1453));
Q_FDP0UA U1824 ( .D(n1453), .QTFCLK( ), .Q(aCount[23]));
Q_MX02 U1825 ( .S(n1427), .A0(aCount[24]), .A1(n1475), .Z(n1454));
Q_FDP0UA U1826 ( .D(n1454), .QTFCLK( ), .Q(aCount[24]));
Q_MX02 U1827 ( .S(n1427), .A0(aCount[25]), .A1(n1473), .Z(n1455));
Q_FDP0UA U1828 ( .D(n1455), .QTFCLK( ), .Q(aCount[25]));
Q_MX02 U1829 ( .S(n1427), .A0(aCount[26]), .A1(n1471), .Z(n1456));
Q_FDP0UA U1830 ( .D(n1456), .QTFCLK( ), .Q(aCount[26]));
Q_MX02 U1831 ( .S(n1427), .A0(aCount[27]), .A1(n1469), .Z(n1457));
Q_FDP0UA U1832 ( .D(n1457), .QTFCLK( ), .Q(aCount[27]));
Q_MX02 U1833 ( .S(n1427), .A0(aCount[28]), .A1(n1467), .Z(n1458));
Q_FDP0UA U1834 ( .D(n1458), .QTFCLK( ), .Q(aCount[28]));
Q_MX02 U1835 ( .S(n1427), .A0(aCount[29]), .A1(n1465), .Z(n1459));
Q_FDP0UA U1836 ( .D(n1459), .QTFCLK( ), .Q(aCount[29]));
Q_MX02 U1837 ( .S(n1427), .A0(aCount[30]), .A1(n1463), .Z(n1460));
Q_FDP0UA U1838 ( .D(n1460), .QTFCLK( ), .Q(aCount[30]));
Q_FDP0UA U1839 ( .D(n1461), .QTFCLK( ), .Q(aCount[31]));
Q_XOR2 U1840 ( .A0(aCount[31]), .A1(n9), .Z(n1461));
Q_AD01HF U1841 ( .A0(aCount[30]), .B0(n1464), .S(n1463), .CO(n1462));
Q_AD01HF U1842 ( .A0(aCount[29]), .B0(n1466), .S(n1465), .CO(n1464));
Q_AD01HF U1843 ( .A0(aCount[28]), .B0(n1468), .S(n1467), .CO(n1466));
Q_AD01HF U1844 ( .A0(aCount[27]), .B0(n1470), .S(n1469), .CO(n1468));
Q_AD01HF U1845 ( .A0(aCount[26]), .B0(n1472), .S(n1471), .CO(n1470));
Q_AD01HF U1846 ( .A0(aCount[25]), .B0(n1474), .S(n1473), .CO(n1472));
Q_AD01HF U1847 ( .A0(aCount[24]), .B0(n1476), .S(n1475), .CO(n1474));
Q_AD01HF U1848 ( .A0(aCount[23]), .B0(n1478), .S(n1477), .CO(n1476));
Q_AD01HF U1849 ( .A0(aCount[22]), .B0(n1480), .S(n1479), .CO(n1478));
Q_AD01HF U1850 ( .A0(aCount[21]), .B0(n1482), .S(n1481), .CO(n1480));
Q_AD01HF U1851 ( .A0(aCount[20]), .B0(n1484), .S(n1483), .CO(n1482));
Q_AD01HF U1852 ( .A0(aCount[19]), .B0(n1486), .S(n1485), .CO(n1484));
Q_AD01HF U1853 ( .A0(aCount[18]), .B0(n1488), .S(n1487), .CO(n1486));
Q_AD01HF U1854 ( .A0(aCount[17]), .B0(n1490), .S(n1489), .CO(n1488));
Q_AD01HF U1855 ( .A0(aCount[16]), .B0(n1492), .S(n1491), .CO(n1490));
Q_AD01HF U1856 ( .A0(aCount[15]), .B0(n1494), .S(n1493), .CO(n1492));
Q_AD01HF U1857 ( .A0(aCount[14]), .B0(n1496), .S(n1495), .CO(n1494));
Q_AD01HF U1858 ( .A0(aCount[13]), .B0(n1498), .S(n1497), .CO(n1496));
Q_AD01HF U1859 ( .A0(aCount[12]), .B0(n1500), .S(n1499), .CO(n1498));
Q_AD01HF U1860 ( .A0(aCount[11]), .B0(n1502), .S(n1501), .CO(n1500));
Q_AD01HF U1861 ( .A0(aCount[10]), .B0(n1504), .S(n1503), .CO(n1502));
Q_AD01HF U1862 ( .A0(aCount[9]), .B0(n1506), .S(n1505), .CO(n1504));
Q_AD01HF U1863 ( .A0(aCount[8]), .B0(n1508), .S(n1507), .CO(n1506));
Q_AD01HF U1864 ( .A0(aCount[7]), .B0(n1510), .S(n1509), .CO(n1508));
Q_AD01HF U1865 ( .A0(aCount[6]), .B0(n1512), .S(n1511), .CO(n1510));
Q_AD01HF U1866 ( .A0(aCount[5]), .B0(n1514), .S(n1513), .CO(n1512));
Q_AD01HF U1867 ( .A0(aCount[4]), .B0(n1516), .S(n1515), .CO(n1514));
Q_AD01HF U1868 ( .A0(aCount[3]), .B0(n1518), .S(n1517), .CO(n1516));
Q_AD01HF U1869 ( .A0(aCount[2]), .B0(n1520), .S(n1519), .CO(n1518));
Q_AD01HF U1870 ( .A0(aCount[1]), .B0(aCount[0]), .S(n1521), .CO(n1520));
Q_OR02 U1871 ( .A0(xpHold), .A1(bpWait), .Z(n1525));
Q_NR02 U1872 ( .A0(sampleXpChg), .A1(n1525), .Z(n1526));
Q_OR02 U1873 ( .A0(bClkHold), .A1(n1526), .Z(n1531));
Q_INV U1874 ( .A(ixcHoldClk), .Z(n1527));
Q_OR02 U1875 ( .A0(n1527), .A1(n1531), .Z(n1528));
Q_INV U1876 ( .A(n1528), .Z(n1522));
Q_INV U1877 ( .A(sampleXpChg), .Z(n1529));
Q_OR03 U1878 ( .A0(n1529), .A1(bpWait), .A2(bClkHold), .Z(n1530));
Q_INV U1879 ( .A(n1530), .Z(n1523));
Q_INV U1880 ( .A(n1531), .Z(n1524));
Q_XOR2 U1881 ( .A0(n1522), .A1(ixcHoldClkCnt[0]), .Z(n1532));
Q_FDP0UA U1882 ( .D(n1532), .QTFCLK( ), .Q(ixcHoldClkCnt[0]));
Q_MX02 U1883 ( .S(n1528), .A0(n1847), .A1(ixcHoldClkCnt[1]), .Z(n1533));
Q_FDP0UA U1884 ( .D(n1533), .QTFCLK( ), .Q(ixcHoldClkCnt[1]));
Q_MX02 U1885 ( .S(n1528), .A0(n1845), .A1(ixcHoldClkCnt[2]), .Z(n1534));
Q_FDP0UA U1886 ( .D(n1534), .QTFCLK( ), .Q(ixcHoldClkCnt[2]));
Q_MX02 U1887 ( .S(n1528), .A0(n1843), .A1(ixcHoldClkCnt[3]), .Z(n1535));
Q_FDP0UA U1888 ( .D(n1535), .QTFCLK( ), .Q(ixcHoldClkCnt[3]));
Q_MX02 U1889 ( .S(n1528), .A0(n1841), .A1(ixcHoldClkCnt[4]), .Z(n1536));
Q_FDP0UA U1890 ( .D(n1536), .QTFCLK( ), .Q(ixcHoldClkCnt[4]));
Q_MX02 U1891 ( .S(n1528), .A0(n1839), .A1(ixcHoldClkCnt[5]), .Z(n1537));
Q_FDP0UA U1892 ( .D(n1537), .QTFCLK( ), .Q(ixcHoldClkCnt[5]));
Q_MX02 U1893 ( .S(n1528), .A0(n1837), .A1(ixcHoldClkCnt[6]), .Z(n1538));
Q_FDP0UA U1894 ( .D(n1538), .QTFCLK( ), .Q(ixcHoldClkCnt[6]));
Q_MX02 U1895 ( .S(n1528), .A0(n1835), .A1(ixcHoldClkCnt[7]), .Z(n1539));
Q_FDP0UA U1896 ( .D(n1539), .QTFCLK( ), .Q(ixcHoldClkCnt[7]));
Q_MX02 U1897 ( .S(n1528), .A0(n1833), .A1(ixcHoldClkCnt[8]), .Z(n1540));
Q_FDP0UA U1898 ( .D(n1540), .QTFCLK( ), .Q(ixcHoldClkCnt[8]));
Q_MX02 U1899 ( .S(n1528), .A0(n1831), .A1(ixcHoldClkCnt[9]), .Z(n1541));
Q_FDP0UA U1900 ( .D(n1541), .QTFCLK( ), .Q(ixcHoldClkCnt[9]));
Q_MX02 U1901 ( .S(n1528), .A0(n1829), .A1(ixcHoldClkCnt[10]), .Z(n1542));
Q_FDP0UA U1902 ( .D(n1542), .QTFCLK( ), .Q(ixcHoldClkCnt[10]));
Q_MX02 U1903 ( .S(n1528), .A0(n1827), .A1(ixcHoldClkCnt[11]), .Z(n1543));
Q_FDP0UA U1904 ( .D(n1543), .QTFCLK( ), .Q(ixcHoldClkCnt[11]));
Q_MX02 U1905 ( .S(n1528), .A0(n1825), .A1(ixcHoldClkCnt[12]), .Z(n1544));
Q_FDP0UA U1906 ( .D(n1544), .QTFCLK( ), .Q(ixcHoldClkCnt[12]));
Q_MX02 U1907 ( .S(n1528), .A0(n1823), .A1(ixcHoldClkCnt[13]), .Z(n1545));
Q_FDP0UA U1908 ( .D(n1545), .QTFCLK( ), .Q(ixcHoldClkCnt[13]));
Q_MX02 U1909 ( .S(n1528), .A0(n1821), .A1(ixcHoldClkCnt[14]), .Z(n1546));
Q_FDP0UA U1910 ( .D(n1546), .QTFCLK( ), .Q(ixcHoldClkCnt[14]));
Q_MX02 U1911 ( .S(n1528), .A0(n1819), .A1(ixcHoldClkCnt[15]), .Z(n1547));
Q_FDP0UA U1912 ( .D(n1547), .QTFCLK( ), .Q(ixcHoldClkCnt[15]));
Q_MX02 U1913 ( .S(n1528), .A0(n1817), .A1(ixcHoldClkCnt[16]), .Z(n1548));
Q_FDP0UA U1914 ( .D(n1548), .QTFCLK( ), .Q(ixcHoldClkCnt[16]));
Q_MX02 U1915 ( .S(n1528), .A0(n1815), .A1(ixcHoldClkCnt[17]), .Z(n1549));
Q_FDP0UA U1916 ( .D(n1549), .QTFCLK( ), .Q(ixcHoldClkCnt[17]));
Q_MX02 U1917 ( .S(n1528), .A0(n1813), .A1(ixcHoldClkCnt[18]), .Z(n1550));
Q_FDP0UA U1918 ( .D(n1550), .QTFCLK( ), .Q(ixcHoldClkCnt[18]));
Q_MX02 U1919 ( .S(n1528), .A0(n1811), .A1(ixcHoldClkCnt[19]), .Z(n1551));
Q_FDP0UA U1920 ( .D(n1551), .QTFCLK( ), .Q(ixcHoldClkCnt[19]));
Q_MX02 U1921 ( .S(n1528), .A0(n1809), .A1(ixcHoldClkCnt[20]), .Z(n1552));
Q_FDP0UA U1922 ( .D(n1552), .QTFCLK( ), .Q(ixcHoldClkCnt[20]));
Q_MX02 U1923 ( .S(n1528), .A0(n1807), .A1(ixcHoldClkCnt[21]), .Z(n1553));
Q_FDP0UA U1924 ( .D(n1553), .QTFCLK( ), .Q(ixcHoldClkCnt[21]));
Q_MX02 U1925 ( .S(n1528), .A0(n1805), .A1(ixcHoldClkCnt[22]), .Z(n1554));
Q_FDP0UA U1926 ( .D(n1554), .QTFCLK( ), .Q(ixcHoldClkCnt[22]));
Q_MX02 U1927 ( .S(n1528), .A0(n1803), .A1(ixcHoldClkCnt[23]), .Z(n1555));
Q_FDP0UA U1928 ( .D(n1555), .QTFCLK( ), .Q(ixcHoldClkCnt[23]));
Q_MX02 U1929 ( .S(n1528), .A0(n1801), .A1(ixcHoldClkCnt[24]), .Z(n1556));
Q_FDP0UA U1930 ( .D(n1556), .QTFCLK( ), .Q(ixcHoldClkCnt[24]));
Q_MX02 U1931 ( .S(n1528), .A0(n1799), .A1(ixcHoldClkCnt[25]), .Z(n1557));
Q_FDP0UA U1932 ( .D(n1557), .QTFCLK( ), .Q(ixcHoldClkCnt[25]));
Q_MX02 U1933 ( .S(n1528), .A0(n1797), .A1(ixcHoldClkCnt[26]), .Z(n1558));
Q_FDP0UA U1934 ( .D(n1558), .QTFCLK( ), .Q(ixcHoldClkCnt[26]));
Q_MX02 U1935 ( .S(n1528), .A0(n1795), .A1(ixcHoldClkCnt[27]), .Z(n1559));
Q_FDP0UA U1936 ( .D(n1559), .QTFCLK( ), .Q(ixcHoldClkCnt[27]));
Q_MX02 U1937 ( .S(n1528), .A0(n1793), .A1(ixcHoldClkCnt[28]), .Z(n1560));
Q_FDP0UA U1938 ( .D(n1560), .QTFCLK( ), .Q(ixcHoldClkCnt[28]));
Q_MX02 U1939 ( .S(n1528), .A0(n1791), .A1(ixcHoldClkCnt[29]), .Z(n1561));
Q_FDP0UA U1940 ( .D(n1561), .QTFCLK( ), .Q(ixcHoldClkCnt[29]));
Q_MX02 U1941 ( .S(n1528), .A0(n1789), .A1(ixcHoldClkCnt[30]), .Z(n1562));
Q_FDP0UA U1942 ( .D(n1562), .QTFCLK( ), .Q(ixcHoldClkCnt[30]));
Q_MX02 U1943 ( .S(n1528), .A0(n1787), .A1(ixcHoldClkCnt[31]), .Z(n1563));
Q_FDP0UA U1944 ( .D(n1563), .QTFCLK( ), .Q(ixcHoldClkCnt[31]));
Q_MX02 U1945 ( .S(n1528), .A0(n1785), .A1(ixcHoldClkCnt[32]), .Z(n1564));
Q_FDP0UA U1946 ( .D(n1564), .QTFCLK( ), .Q(ixcHoldClkCnt[32]));
Q_MX02 U1947 ( .S(n1528), .A0(n1783), .A1(ixcHoldClkCnt[33]), .Z(n1565));
Q_FDP0UA U1948 ( .D(n1565), .QTFCLK( ), .Q(ixcHoldClkCnt[33]));
Q_MX02 U1949 ( .S(n1528), .A0(n1781), .A1(ixcHoldClkCnt[34]), .Z(n1566));
Q_FDP0UA U1950 ( .D(n1566), .QTFCLK( ), .Q(ixcHoldClkCnt[34]));
Q_MX02 U1951 ( .S(n1528), .A0(n1779), .A1(ixcHoldClkCnt[35]), .Z(n1567));
Q_FDP0UA U1952 ( .D(n1567), .QTFCLK( ), .Q(ixcHoldClkCnt[35]));
Q_MX02 U1953 ( .S(n1528), .A0(n1777), .A1(ixcHoldClkCnt[36]), .Z(n1568));
Q_FDP0UA U1954 ( .D(n1568), .QTFCLK( ), .Q(ixcHoldClkCnt[36]));
Q_MX02 U1955 ( .S(n1528), .A0(n1775), .A1(ixcHoldClkCnt[37]), .Z(n1569));
Q_FDP0UA U1956 ( .D(n1569), .QTFCLK( ), .Q(ixcHoldClkCnt[37]));
Q_MX02 U1957 ( .S(n1528), .A0(n1773), .A1(ixcHoldClkCnt[38]), .Z(n1570));
Q_FDP0UA U1958 ( .D(n1570), .QTFCLK( ), .Q(ixcHoldClkCnt[38]));
Q_MX02 U1959 ( .S(n1528), .A0(n1771), .A1(ixcHoldClkCnt[39]), .Z(n1571));
Q_FDP0UA U1960 ( .D(n1571), .QTFCLK( ), .Q(ixcHoldClkCnt[39]));
Q_MX02 U1961 ( .S(n1528), .A0(n1769), .A1(ixcHoldClkCnt[40]), .Z(n1572));
Q_FDP0UA U1962 ( .D(n1572), .QTFCLK( ), .Q(ixcHoldClkCnt[40]));
Q_MX02 U1963 ( .S(n1528), .A0(n1767), .A1(ixcHoldClkCnt[41]), .Z(n1573));
Q_FDP0UA U1964 ( .D(n1573), .QTFCLK( ), .Q(ixcHoldClkCnt[41]));
Q_MX02 U1965 ( .S(n1528), .A0(n1765), .A1(ixcHoldClkCnt[42]), .Z(n1574));
Q_FDP0UA U1966 ( .D(n1574), .QTFCLK( ), .Q(ixcHoldClkCnt[42]));
Q_MX02 U1967 ( .S(n1528), .A0(n1763), .A1(ixcHoldClkCnt[43]), .Z(n1575));
Q_FDP0UA U1968 ( .D(n1575), .QTFCLK( ), .Q(ixcHoldClkCnt[43]));
Q_MX02 U1969 ( .S(n1528), .A0(n1761), .A1(ixcHoldClkCnt[44]), .Z(n1576));
Q_FDP0UA U1970 ( .D(n1576), .QTFCLK( ), .Q(ixcHoldClkCnt[44]));
Q_MX02 U1971 ( .S(n1528), .A0(n1759), .A1(ixcHoldClkCnt[45]), .Z(n1577));
Q_FDP0UA U1972 ( .D(n1577), .QTFCLK( ), .Q(ixcHoldClkCnt[45]));
Q_MX02 U1973 ( .S(n1528), .A0(n1757), .A1(ixcHoldClkCnt[46]), .Z(n1578));
Q_FDP0UA U1974 ( .D(n1578), .QTFCLK( ), .Q(ixcHoldClkCnt[46]));
Q_MX02 U1975 ( .S(n1528), .A0(n1755), .A1(ixcHoldClkCnt[47]), .Z(n1579));
Q_FDP0UA U1976 ( .D(n1579), .QTFCLK( ), .Q(ixcHoldClkCnt[47]));
Q_MX02 U1977 ( .S(n1528), .A0(n1753), .A1(ixcHoldClkCnt[48]), .Z(n1580));
Q_FDP0UA U1978 ( .D(n1580), .QTFCLK( ), .Q(ixcHoldClkCnt[48]));
Q_MX02 U1979 ( .S(n1528), .A0(n1751), .A1(ixcHoldClkCnt[49]), .Z(n1581));
Q_FDP0UA U1980 ( .D(n1581), .QTFCLK( ), .Q(ixcHoldClkCnt[49]));
Q_MX02 U1981 ( .S(n1528), .A0(n1749), .A1(ixcHoldClkCnt[50]), .Z(n1582));
Q_FDP0UA U1982 ( .D(n1582), .QTFCLK( ), .Q(ixcHoldClkCnt[50]));
Q_MX02 U1983 ( .S(n1528), .A0(n1747), .A1(ixcHoldClkCnt[51]), .Z(n1583));
Q_FDP0UA U1984 ( .D(n1583), .QTFCLK( ), .Q(ixcHoldClkCnt[51]));
Q_MX02 U1985 ( .S(n1528), .A0(n1745), .A1(ixcHoldClkCnt[52]), .Z(n1584));
Q_FDP0UA U1986 ( .D(n1584), .QTFCLK( ), .Q(ixcHoldClkCnt[52]));
Q_MX02 U1987 ( .S(n1528), .A0(n1743), .A1(ixcHoldClkCnt[53]), .Z(n1585));
Q_FDP0UA U1988 ( .D(n1585), .QTFCLK( ), .Q(ixcHoldClkCnt[53]));
Q_MX02 U1989 ( .S(n1528), .A0(n1741), .A1(ixcHoldClkCnt[54]), .Z(n1586));
Q_FDP0UA U1990 ( .D(n1586), .QTFCLK( ), .Q(ixcHoldClkCnt[54]));
Q_MX02 U1991 ( .S(n1528), .A0(n1739), .A1(ixcHoldClkCnt[55]), .Z(n1587));
Q_FDP0UA U1992 ( .D(n1587), .QTFCLK( ), .Q(ixcHoldClkCnt[55]));
Q_MX02 U1993 ( .S(n1528), .A0(n1737), .A1(ixcHoldClkCnt[56]), .Z(n1588));
Q_FDP0UA U1994 ( .D(n1588), .QTFCLK( ), .Q(ixcHoldClkCnt[56]));
Q_MX02 U1995 ( .S(n1528), .A0(n1735), .A1(ixcHoldClkCnt[57]), .Z(n1589));
Q_FDP0UA U1996 ( .D(n1589), .QTFCLK( ), .Q(ixcHoldClkCnt[57]));
Q_MX02 U1997 ( .S(n1528), .A0(n1733), .A1(ixcHoldClkCnt[58]), .Z(n1590));
Q_FDP0UA U1998 ( .D(n1590), .QTFCLK( ), .Q(ixcHoldClkCnt[58]));
Q_MX02 U1999 ( .S(n1528), .A0(n1731), .A1(ixcHoldClkCnt[59]), .Z(n1591));
Q_FDP0UA U2000 ( .D(n1591), .QTFCLK( ), .Q(ixcHoldClkCnt[59]));
Q_MX02 U2001 ( .S(n1528), .A0(n1729), .A1(ixcHoldClkCnt[60]), .Z(n1592));
Q_FDP0UA U2002 ( .D(n1592), .QTFCLK( ), .Q(ixcHoldClkCnt[60]));
Q_MX02 U2003 ( .S(n1528), .A0(n1727), .A1(ixcHoldClkCnt[61]), .Z(n1593));
Q_FDP0UA U2004 ( .D(n1593), .QTFCLK( ), .Q(ixcHoldClkCnt[61]));
Q_MX02 U2005 ( .S(n1528), .A0(n1725), .A1(ixcHoldClkCnt[62]), .Z(n1594));
Q_FDP0UA U2006 ( .D(n1594), .QTFCLK( ), .Q(ixcHoldClkCnt[62]));
Q_FDP0UA U2007 ( .D(n1595), .QTFCLK( ), .Q(ixcHoldClkCnt[63]));
Q_XOR2 U2008 ( .A0(n1523), .A1(nbaCount[0]), .Z(n1596));
Q_FDP0UA U2009 ( .D(n1596), .QTFCLK( ), .Q(nbaCount[0]));
Q_MX02 U2010 ( .S(n1530), .A0(n1971), .A1(nbaCount[1]), .Z(n1597));
Q_FDP0UA U2011 ( .D(n1597), .QTFCLK( ), .Q(nbaCount[1]));
Q_MX02 U2012 ( .S(n1530), .A0(n1969), .A1(nbaCount[2]), .Z(n1598));
Q_FDP0UA U2013 ( .D(n1598), .QTFCLK( ), .Q(nbaCount[2]));
Q_MX02 U2014 ( .S(n1530), .A0(n1967), .A1(nbaCount[3]), .Z(n1599));
Q_FDP0UA U2015 ( .D(n1599), .QTFCLK( ), .Q(nbaCount[3]));
Q_MX02 U2016 ( .S(n1530), .A0(n1965), .A1(nbaCount[4]), .Z(n1600));
Q_FDP0UA U2017 ( .D(n1600), .QTFCLK( ), .Q(nbaCount[4]));
Q_MX02 U2018 ( .S(n1530), .A0(n1963), .A1(nbaCount[5]), .Z(n1601));
Q_FDP0UA U2019 ( .D(n1601), .QTFCLK( ), .Q(nbaCount[5]));
Q_MX02 U2020 ( .S(n1530), .A0(n1961), .A1(nbaCount[6]), .Z(n1602));
Q_FDP0UA U2021 ( .D(n1602), .QTFCLK( ), .Q(nbaCount[6]));
Q_MX02 U2022 ( .S(n1530), .A0(n1959), .A1(nbaCount[7]), .Z(n1603));
Q_FDP0UA U2023 ( .D(n1603), .QTFCLK( ), .Q(nbaCount[7]));
Q_MX02 U2024 ( .S(n1530), .A0(n1957), .A1(nbaCount[8]), .Z(n1604));
Q_FDP0UA U2025 ( .D(n1604), .QTFCLK( ), .Q(nbaCount[8]));
Q_MX02 U2026 ( .S(n1530), .A0(n1955), .A1(nbaCount[9]), .Z(n1605));
Q_FDP0UA U2027 ( .D(n1605), .QTFCLK( ), .Q(nbaCount[9]));
Q_MX02 U2028 ( .S(n1530), .A0(n1953), .A1(nbaCount[10]), .Z(n1606));
Q_FDP0UA U2029 ( .D(n1606), .QTFCLK( ), .Q(nbaCount[10]));
Q_MX02 U2030 ( .S(n1530), .A0(n1951), .A1(nbaCount[11]), .Z(n1607));
Q_FDP0UA U2031 ( .D(n1607), .QTFCLK( ), .Q(nbaCount[11]));
Q_MX02 U2032 ( .S(n1530), .A0(n1949), .A1(nbaCount[12]), .Z(n1608));
Q_FDP0UA U2033 ( .D(n1608), .QTFCLK( ), .Q(nbaCount[12]));
Q_MX02 U2034 ( .S(n1530), .A0(n1947), .A1(nbaCount[13]), .Z(n1609));
Q_FDP0UA U2035 ( .D(n1609), .QTFCLK( ), .Q(nbaCount[13]));
Q_MX02 U2036 ( .S(n1530), .A0(n1945), .A1(nbaCount[14]), .Z(n1610));
Q_FDP0UA U2037 ( .D(n1610), .QTFCLK( ), .Q(nbaCount[14]));
Q_MX02 U2038 ( .S(n1530), .A0(n1943), .A1(nbaCount[15]), .Z(n1611));
Q_FDP0UA U2039 ( .D(n1611), .QTFCLK( ), .Q(nbaCount[15]));
Q_MX02 U2040 ( .S(n1530), .A0(n1941), .A1(nbaCount[16]), .Z(n1612));
Q_FDP0UA U2041 ( .D(n1612), .QTFCLK( ), .Q(nbaCount[16]));
Q_MX02 U2042 ( .S(n1530), .A0(n1939), .A1(nbaCount[17]), .Z(n1613));
Q_FDP0UA U2043 ( .D(n1613), .QTFCLK( ), .Q(nbaCount[17]));
Q_MX02 U2044 ( .S(n1530), .A0(n1937), .A1(nbaCount[18]), .Z(n1614));
Q_FDP0UA U2045 ( .D(n1614), .QTFCLK( ), .Q(nbaCount[18]));
Q_MX02 U2046 ( .S(n1530), .A0(n1935), .A1(nbaCount[19]), .Z(n1615));
Q_FDP0UA U2047 ( .D(n1615), .QTFCLK( ), .Q(nbaCount[19]));
Q_MX02 U2048 ( .S(n1530), .A0(n1933), .A1(nbaCount[20]), .Z(n1616));
Q_FDP0UA U2049 ( .D(n1616), .QTFCLK( ), .Q(nbaCount[20]));
Q_MX02 U2050 ( .S(n1530), .A0(n1931), .A1(nbaCount[21]), .Z(n1617));
Q_FDP0UA U2051 ( .D(n1617), .QTFCLK( ), .Q(nbaCount[21]));
Q_MX02 U2052 ( .S(n1530), .A0(n1929), .A1(nbaCount[22]), .Z(n1618));
Q_FDP0UA U2053 ( .D(n1618), .QTFCLK( ), .Q(nbaCount[22]));
Q_MX02 U2054 ( .S(n1530), .A0(n1927), .A1(nbaCount[23]), .Z(n1619));
Q_FDP0UA U2055 ( .D(n1619), .QTFCLK( ), .Q(nbaCount[23]));
Q_MX02 U2056 ( .S(n1530), .A0(n1925), .A1(nbaCount[24]), .Z(n1620));
Q_FDP0UA U2057 ( .D(n1620), .QTFCLK( ), .Q(nbaCount[24]));
Q_MX02 U2058 ( .S(n1530), .A0(n1923), .A1(nbaCount[25]), .Z(n1621));
Q_FDP0UA U2059 ( .D(n1621), .QTFCLK( ), .Q(nbaCount[25]));
Q_MX02 U2060 ( .S(n1530), .A0(n1921), .A1(nbaCount[26]), .Z(n1622));
Q_FDP0UA U2061 ( .D(n1622), .QTFCLK( ), .Q(nbaCount[26]));
Q_MX02 U2062 ( .S(n1530), .A0(n1919), .A1(nbaCount[27]), .Z(n1623));
Q_FDP0UA U2063 ( .D(n1623), .QTFCLK( ), .Q(nbaCount[27]));
Q_MX02 U2064 ( .S(n1530), .A0(n1917), .A1(nbaCount[28]), .Z(n1624));
Q_FDP0UA U2065 ( .D(n1624), .QTFCLK( ), .Q(nbaCount[28]));
Q_MX02 U2066 ( .S(n1530), .A0(n1915), .A1(nbaCount[29]), .Z(n1625));
Q_FDP0UA U2067 ( .D(n1625), .QTFCLK( ), .Q(nbaCount[29]));
Q_MX02 U2068 ( .S(n1530), .A0(n1913), .A1(nbaCount[30]), .Z(n1626));
Q_FDP0UA U2069 ( .D(n1626), .QTFCLK( ), .Q(nbaCount[30]));
Q_MX02 U2070 ( .S(n1530), .A0(n1911), .A1(nbaCount[31]), .Z(n1627));
Q_FDP0UA U2071 ( .D(n1627), .QTFCLK( ), .Q(nbaCount[31]));
Q_MX02 U2072 ( .S(n1530), .A0(n1909), .A1(nbaCount[32]), .Z(n1628));
Q_FDP0UA U2073 ( .D(n1628), .QTFCLK( ), .Q(nbaCount[32]));
Q_MX02 U2074 ( .S(n1530), .A0(n1907), .A1(nbaCount[33]), .Z(n1629));
Q_FDP0UA U2075 ( .D(n1629), .QTFCLK( ), .Q(nbaCount[33]));
Q_MX02 U2076 ( .S(n1530), .A0(n1905), .A1(nbaCount[34]), .Z(n1630));
Q_FDP0UA U2077 ( .D(n1630), .QTFCLK( ), .Q(nbaCount[34]));
Q_MX02 U2078 ( .S(n1530), .A0(n1903), .A1(nbaCount[35]), .Z(n1631));
Q_FDP0UA U2079 ( .D(n1631), .QTFCLK( ), .Q(nbaCount[35]));
Q_MX02 U2080 ( .S(n1530), .A0(n1901), .A1(nbaCount[36]), .Z(n1632));
Q_FDP0UA U2081 ( .D(n1632), .QTFCLK( ), .Q(nbaCount[36]));
Q_MX02 U2082 ( .S(n1530), .A0(n1899), .A1(nbaCount[37]), .Z(n1633));
Q_FDP0UA U2083 ( .D(n1633), .QTFCLK( ), .Q(nbaCount[37]));
Q_MX02 U2084 ( .S(n1530), .A0(n1897), .A1(nbaCount[38]), .Z(n1634));
Q_FDP0UA U2085 ( .D(n1634), .QTFCLK( ), .Q(nbaCount[38]));
Q_MX02 U2086 ( .S(n1530), .A0(n1895), .A1(nbaCount[39]), .Z(n1635));
Q_FDP0UA U2087 ( .D(n1635), .QTFCLK( ), .Q(nbaCount[39]));
Q_MX02 U2088 ( .S(n1530), .A0(n1893), .A1(nbaCount[40]), .Z(n1636));
Q_FDP0UA U2089 ( .D(n1636), .QTFCLK( ), .Q(nbaCount[40]));
Q_MX02 U2090 ( .S(n1530), .A0(n1891), .A1(nbaCount[41]), .Z(n1637));
Q_FDP0UA U2091 ( .D(n1637), .QTFCLK( ), .Q(nbaCount[41]));
Q_MX02 U2092 ( .S(n1530), .A0(n1889), .A1(nbaCount[42]), .Z(n1638));
Q_FDP0UA U2093 ( .D(n1638), .QTFCLK( ), .Q(nbaCount[42]));
Q_MX02 U2094 ( .S(n1530), .A0(n1887), .A1(nbaCount[43]), .Z(n1639));
Q_FDP0UA U2095 ( .D(n1639), .QTFCLK( ), .Q(nbaCount[43]));
Q_MX02 U2096 ( .S(n1530), .A0(n1885), .A1(nbaCount[44]), .Z(n1640));
Q_FDP0UA U2097 ( .D(n1640), .QTFCLK( ), .Q(nbaCount[44]));
Q_MX02 U2098 ( .S(n1530), .A0(n1883), .A1(nbaCount[45]), .Z(n1641));
Q_FDP0UA U2099 ( .D(n1641), .QTFCLK( ), .Q(nbaCount[45]));
Q_MX02 U2100 ( .S(n1530), .A0(n1881), .A1(nbaCount[46]), .Z(n1642));
Q_FDP0UA U2101 ( .D(n1642), .QTFCLK( ), .Q(nbaCount[46]));
Q_MX02 U2102 ( .S(n1530), .A0(n1879), .A1(nbaCount[47]), .Z(n1643));
Q_FDP0UA U2103 ( .D(n1643), .QTFCLK( ), .Q(nbaCount[47]));
Q_MX02 U2104 ( .S(n1530), .A0(n1877), .A1(nbaCount[48]), .Z(n1644));
Q_FDP0UA U2105 ( .D(n1644), .QTFCLK( ), .Q(nbaCount[48]));
Q_MX02 U2106 ( .S(n1530), .A0(n1875), .A1(nbaCount[49]), .Z(n1645));
Q_FDP0UA U2107 ( .D(n1645), .QTFCLK( ), .Q(nbaCount[49]));
Q_MX02 U2108 ( .S(n1530), .A0(n1873), .A1(nbaCount[50]), .Z(n1646));
Q_FDP0UA U2109 ( .D(n1646), .QTFCLK( ), .Q(nbaCount[50]));
Q_MX02 U2110 ( .S(n1530), .A0(n1871), .A1(nbaCount[51]), .Z(n1647));
Q_FDP0UA U2111 ( .D(n1647), .QTFCLK( ), .Q(nbaCount[51]));
Q_MX02 U2112 ( .S(n1530), .A0(n1869), .A1(nbaCount[52]), .Z(n1648));
Q_FDP0UA U2113 ( .D(n1648), .QTFCLK( ), .Q(nbaCount[52]));
Q_MX02 U2114 ( .S(n1530), .A0(n1867), .A1(nbaCount[53]), .Z(n1649));
Q_FDP0UA U2115 ( .D(n1649), .QTFCLK( ), .Q(nbaCount[53]));
Q_MX02 U2116 ( .S(n1530), .A0(n1865), .A1(nbaCount[54]), .Z(n1650));
Q_FDP0UA U2117 ( .D(n1650), .QTFCLK( ), .Q(nbaCount[54]));
Q_MX02 U2118 ( .S(n1530), .A0(n1863), .A1(nbaCount[55]), .Z(n1651));
Q_FDP0UA U2119 ( .D(n1651), .QTFCLK( ), .Q(nbaCount[55]));
Q_MX02 U2120 ( .S(n1530), .A0(n1861), .A1(nbaCount[56]), .Z(n1652));
Q_FDP0UA U2121 ( .D(n1652), .QTFCLK( ), .Q(nbaCount[56]));
Q_MX02 U2122 ( .S(n1530), .A0(n1859), .A1(nbaCount[57]), .Z(n1653));
Q_FDP0UA U2123 ( .D(n1653), .QTFCLK( ), .Q(nbaCount[57]));
Q_MX02 U2124 ( .S(n1530), .A0(n1857), .A1(nbaCount[58]), .Z(n1654));
Q_FDP0UA U2125 ( .D(n1654), .QTFCLK( ), .Q(nbaCount[58]));
Q_MX02 U2126 ( .S(n1530), .A0(n1855), .A1(nbaCount[59]), .Z(n1655));
Q_FDP0UA U2127 ( .D(n1655), .QTFCLK( ), .Q(nbaCount[59]));
Q_MX02 U2128 ( .S(n1530), .A0(n1853), .A1(nbaCount[60]), .Z(n1656));
Q_FDP0UA U2129 ( .D(n1656), .QTFCLK( ), .Q(nbaCount[60]));
Q_MX02 U2130 ( .S(n1530), .A0(n1851), .A1(nbaCount[61]), .Z(n1657));
Q_FDP0UA U2131 ( .D(n1657), .QTFCLK( ), .Q(nbaCount[61]));
Q_MX02 U2132 ( .S(n1530), .A0(n1849), .A1(nbaCount[62]), .Z(n1658));
Q_FDP0UA U2133 ( .D(n1658), .QTFCLK( ), .Q(nbaCount[62]));
Q_FDP0UA U2134 ( .D(n1659), .QTFCLK( ), .Q(nbaCount[63]));
Q_XOR2 U2135 ( .A0(n1524), .A1(bCount[0]), .Z(n1660));
Q_FDP0UA U2136 ( .D(n1660), .QTFCLK( ), .Q(bCount[0]));
Q_MX02 U2137 ( .S(n1531), .A0(n2095), .A1(bCount[1]), .Z(n1661));
Q_FDP0UA U2138 ( .D(n1661), .QTFCLK( ), .Q(bCount[1]));
Q_MX02 U2139 ( .S(n1531), .A0(n2093), .A1(bCount[2]), .Z(n1662));
Q_FDP0UA U2140 ( .D(n1662), .QTFCLK( ), .Q(bCount[2]));
Q_MX02 U2141 ( .S(n1531), .A0(n2091), .A1(bCount[3]), .Z(n1663));
Q_FDP0UA U2142 ( .D(n1663), .QTFCLK( ), .Q(bCount[3]));
Q_MX02 U2143 ( .S(n1531), .A0(n2089), .A1(bCount[4]), .Z(n1664));
Q_FDP0UA U2144 ( .D(n1664), .QTFCLK( ), .Q(bCount[4]));
Q_MX02 U2145 ( .S(n1531), .A0(n2087), .A1(bCount[5]), .Z(n1665));
Q_FDP0UA U2146 ( .D(n1665), .QTFCLK( ), .Q(bCount[5]));
Q_MX02 U2147 ( .S(n1531), .A0(n2085), .A1(bCount[6]), .Z(n1666));
Q_FDP0UA U2148 ( .D(n1666), .QTFCLK( ), .Q(bCount[6]));
Q_MX02 U2149 ( .S(n1531), .A0(n2083), .A1(bCount[7]), .Z(n1667));
Q_FDP0UA U2150 ( .D(n1667), .QTFCLK( ), .Q(bCount[7]));
Q_MX02 U2151 ( .S(n1531), .A0(n2081), .A1(bCount[8]), .Z(n1668));
Q_FDP0UA U2152 ( .D(n1668), .QTFCLK( ), .Q(bCount[8]));
Q_MX02 U2153 ( .S(n1531), .A0(n2079), .A1(bCount[9]), .Z(n1669));
Q_FDP0UA U2154 ( .D(n1669), .QTFCLK( ), .Q(bCount[9]));
Q_MX02 U2155 ( .S(n1531), .A0(n2077), .A1(bCount[10]), .Z(n1670));
Q_FDP0UA U2156 ( .D(n1670), .QTFCLK( ), .Q(bCount[10]));
Q_MX02 U2157 ( .S(n1531), .A0(n2075), .A1(bCount[11]), .Z(n1671));
Q_FDP0UA U2158 ( .D(n1671), .QTFCLK( ), .Q(bCount[11]));
Q_MX02 U2159 ( .S(n1531), .A0(n2073), .A1(bCount[12]), .Z(n1672));
Q_FDP0UA U2160 ( .D(n1672), .QTFCLK( ), .Q(bCount[12]));
Q_MX02 U2161 ( .S(n1531), .A0(n2071), .A1(bCount[13]), .Z(n1673));
Q_FDP0UA U2162 ( .D(n1673), .QTFCLK( ), .Q(bCount[13]));
Q_MX02 U2163 ( .S(n1531), .A0(n2069), .A1(bCount[14]), .Z(n1674));
Q_FDP0UA U2164 ( .D(n1674), .QTFCLK( ), .Q(bCount[14]));
Q_MX02 U2165 ( .S(n1531), .A0(n2067), .A1(bCount[15]), .Z(n1675));
Q_FDP0UA U2166 ( .D(n1675), .QTFCLK( ), .Q(bCount[15]));
Q_MX02 U2167 ( .S(n1531), .A0(n2065), .A1(bCount[16]), .Z(n1676));
Q_FDP0UA U2168 ( .D(n1676), .QTFCLK( ), .Q(bCount[16]));
Q_MX02 U2169 ( .S(n1531), .A0(n2063), .A1(bCount[17]), .Z(n1677));
Q_FDP0UA U2170 ( .D(n1677), .QTFCLK( ), .Q(bCount[17]));
Q_MX02 U2171 ( .S(n1531), .A0(n2061), .A1(bCount[18]), .Z(n1678));
Q_FDP0UA U2172 ( .D(n1678), .QTFCLK( ), .Q(bCount[18]));
Q_MX02 U2173 ( .S(n1531), .A0(n2059), .A1(bCount[19]), .Z(n1679));
Q_FDP0UA U2174 ( .D(n1679), .QTFCLK( ), .Q(bCount[19]));
Q_MX02 U2175 ( .S(n1531), .A0(n2057), .A1(bCount[20]), .Z(n1680));
Q_FDP0UA U2176 ( .D(n1680), .QTFCLK( ), .Q(bCount[20]));
Q_MX02 U2177 ( .S(n1531), .A0(n2055), .A1(bCount[21]), .Z(n1681));
Q_FDP0UA U2178 ( .D(n1681), .QTFCLK( ), .Q(bCount[21]));
Q_MX02 U2179 ( .S(n1531), .A0(n2053), .A1(bCount[22]), .Z(n1682));
Q_FDP0UA U2180 ( .D(n1682), .QTFCLK( ), .Q(bCount[22]));
Q_MX02 U2181 ( .S(n1531), .A0(n2051), .A1(bCount[23]), .Z(n1683));
Q_FDP0UA U2182 ( .D(n1683), .QTFCLK( ), .Q(bCount[23]));
Q_MX02 U2183 ( .S(n1531), .A0(n2049), .A1(bCount[24]), .Z(n1684));
Q_FDP0UA U2184 ( .D(n1684), .QTFCLK( ), .Q(bCount[24]));
Q_MX02 U2185 ( .S(n1531), .A0(n2047), .A1(bCount[25]), .Z(n1685));
Q_FDP0UA U2186 ( .D(n1685), .QTFCLK( ), .Q(bCount[25]));
Q_MX02 U2187 ( .S(n1531), .A0(n2045), .A1(bCount[26]), .Z(n1686));
Q_FDP0UA U2188 ( .D(n1686), .QTFCLK( ), .Q(bCount[26]));
Q_MX02 U2189 ( .S(n1531), .A0(n2043), .A1(bCount[27]), .Z(n1687));
Q_FDP0UA U2190 ( .D(n1687), .QTFCLK( ), .Q(bCount[27]));
Q_MX02 U2191 ( .S(n1531), .A0(n2041), .A1(bCount[28]), .Z(n1688));
Q_FDP0UA U2192 ( .D(n1688), .QTFCLK( ), .Q(bCount[28]));
Q_MX02 U2193 ( .S(n1531), .A0(n2039), .A1(bCount[29]), .Z(n1689));
Q_FDP0UA U2194 ( .D(n1689), .QTFCLK( ), .Q(bCount[29]));
Q_MX02 U2195 ( .S(n1531), .A0(n2037), .A1(bCount[30]), .Z(n1690));
Q_FDP0UA U2196 ( .D(n1690), .QTFCLK( ), .Q(bCount[30]));
Q_MX02 U2197 ( .S(n1531), .A0(n2035), .A1(bCount[31]), .Z(n1691));
Q_FDP0UA U2198 ( .D(n1691), .QTFCLK( ), .Q(bCount[31]));
Q_MX02 U2199 ( .S(n1531), .A0(n2033), .A1(bCount[32]), .Z(n1692));
Q_FDP0UA U2200 ( .D(n1692), .QTFCLK( ), .Q(bCount[32]));
Q_MX02 U2201 ( .S(n1531), .A0(n2031), .A1(bCount[33]), .Z(n1693));
Q_FDP0UA U2202 ( .D(n1693), .QTFCLK( ), .Q(bCount[33]));
Q_MX02 U2203 ( .S(n1531), .A0(n2029), .A1(bCount[34]), .Z(n1694));
Q_FDP0UA U2204 ( .D(n1694), .QTFCLK( ), .Q(bCount[34]));
Q_MX02 U2205 ( .S(n1531), .A0(n2027), .A1(bCount[35]), .Z(n1695));
Q_FDP0UA U2206 ( .D(n1695), .QTFCLK( ), .Q(bCount[35]));
Q_MX02 U2207 ( .S(n1531), .A0(n2025), .A1(bCount[36]), .Z(n1696));
Q_FDP0UA U2208 ( .D(n1696), .QTFCLK( ), .Q(bCount[36]));
Q_MX02 U2209 ( .S(n1531), .A0(n2023), .A1(bCount[37]), .Z(n1697));
Q_FDP0UA U2210 ( .D(n1697), .QTFCLK( ), .Q(bCount[37]));
Q_MX02 U2211 ( .S(n1531), .A0(n2021), .A1(bCount[38]), .Z(n1698));
Q_FDP0UA U2212 ( .D(n1698), .QTFCLK( ), .Q(bCount[38]));
Q_MX02 U2213 ( .S(n1531), .A0(n2019), .A1(bCount[39]), .Z(n1699));
Q_FDP0UA U2214 ( .D(n1699), .QTFCLK( ), .Q(bCount[39]));
Q_MX02 U2215 ( .S(n1531), .A0(n2017), .A1(bCount[40]), .Z(n1700));
Q_FDP0UA U2216 ( .D(n1700), .QTFCLK( ), .Q(bCount[40]));
Q_MX02 U2217 ( .S(n1531), .A0(n2015), .A1(bCount[41]), .Z(n1701));
Q_FDP0UA U2218 ( .D(n1701), .QTFCLK( ), .Q(bCount[41]));
Q_MX02 U2219 ( .S(n1531), .A0(n2013), .A1(bCount[42]), .Z(n1702));
Q_FDP0UA U2220 ( .D(n1702), .QTFCLK( ), .Q(bCount[42]));
Q_MX02 U2221 ( .S(n1531), .A0(n2011), .A1(bCount[43]), .Z(n1703));
Q_FDP0UA U2222 ( .D(n1703), .QTFCLK( ), .Q(bCount[43]));
Q_MX02 U2223 ( .S(n1531), .A0(n2009), .A1(bCount[44]), .Z(n1704));
Q_FDP0UA U2224 ( .D(n1704), .QTFCLK( ), .Q(bCount[44]));
Q_MX02 U2225 ( .S(n1531), .A0(n2007), .A1(bCount[45]), .Z(n1705));
Q_FDP0UA U2226 ( .D(n1705), .QTFCLK( ), .Q(bCount[45]));
Q_MX02 U2227 ( .S(n1531), .A0(n2005), .A1(bCount[46]), .Z(n1706));
Q_FDP0UA U2228 ( .D(n1706), .QTFCLK( ), .Q(bCount[46]));
Q_MX02 U2229 ( .S(n1531), .A0(n2003), .A1(bCount[47]), .Z(n1707));
Q_FDP0UA U2230 ( .D(n1707), .QTFCLK( ), .Q(bCount[47]));
Q_MX02 U2231 ( .S(n1531), .A0(n2001), .A1(bCount[48]), .Z(n1708));
Q_FDP0UA U2232 ( .D(n1708), .QTFCLK( ), .Q(bCount[48]));
Q_MX02 U2233 ( .S(n1531), .A0(n1999), .A1(bCount[49]), .Z(n1709));
Q_FDP0UA U2234 ( .D(n1709), .QTFCLK( ), .Q(bCount[49]));
Q_MX02 U2235 ( .S(n1531), .A0(n1997), .A1(bCount[50]), .Z(n1710));
Q_FDP0UA U2236 ( .D(n1710), .QTFCLK( ), .Q(bCount[50]));
Q_MX02 U2237 ( .S(n1531), .A0(n1995), .A1(bCount[51]), .Z(n1711));
Q_FDP0UA U2238 ( .D(n1711), .QTFCLK( ), .Q(bCount[51]));
Q_MX02 U2239 ( .S(n1531), .A0(n1993), .A1(bCount[52]), .Z(n1712));
Q_FDP0UA U2240 ( .D(n1712), .QTFCLK( ), .Q(bCount[52]));
Q_MX02 U2241 ( .S(n1531), .A0(n1991), .A1(bCount[53]), .Z(n1713));
Q_FDP0UA U2242 ( .D(n1713), .QTFCLK( ), .Q(bCount[53]));
Q_MX02 U2243 ( .S(n1531), .A0(n1989), .A1(bCount[54]), .Z(n1714));
Q_FDP0UA U2244 ( .D(n1714), .QTFCLK( ), .Q(bCount[54]));
Q_MX02 U2245 ( .S(n1531), .A0(n1987), .A1(bCount[55]), .Z(n1715));
Q_FDP0UA U2246 ( .D(n1715), .QTFCLK( ), .Q(bCount[55]));
Q_MX02 U2247 ( .S(n1531), .A0(n1985), .A1(bCount[56]), .Z(n1716));
Q_FDP0UA U2248 ( .D(n1716), .QTFCLK( ), .Q(bCount[56]));
Q_MX02 U2249 ( .S(n1531), .A0(n1983), .A1(bCount[57]), .Z(n1717));
Q_FDP0UA U2250 ( .D(n1717), .QTFCLK( ), .Q(bCount[57]));
Q_MX02 U2251 ( .S(n1531), .A0(n1981), .A1(bCount[58]), .Z(n1718));
Q_FDP0UA U2252 ( .D(n1718), .QTFCLK( ), .Q(bCount[58]));
Q_MX02 U2253 ( .S(n1531), .A0(n1979), .A1(bCount[59]), .Z(n1719));
Q_FDP0UA U2254 ( .D(n1719), .QTFCLK( ), .Q(bCount[59]));
Q_MX02 U2255 ( .S(n1531), .A0(n1977), .A1(bCount[60]), .Z(n1720));
Q_FDP0UA U2256 ( .D(n1720), .QTFCLK( ), .Q(bCount[60]));
Q_MX02 U2257 ( .S(n1531), .A0(n1975), .A1(bCount[61]), .Z(n1721));
Q_FDP0UA U2258 ( .D(n1721), .QTFCLK( ), .Q(bCount[61]));
Q_MX02 U2259 ( .S(n1531), .A0(n1973), .A1(bCount[62]), .Z(n1722));
Q_FDP0UA U2260 ( .D(n1722), .QTFCLK( ), .Q(bCount[62]));
Q_FDP0UA U2261 ( .D(n1723), .QTFCLK( ), .Q(bCount[63]));
Q_XOR2 U2262 ( .A0(ixcHoldClkCnt[63]), .A1(n8), .Z(n1595));
Q_AD01HF U2263 ( .A0(ixcHoldClkCnt[62]), .B0(n1726), .S(n1725), .CO(n1724));
Q_AD01HF U2264 ( .A0(ixcHoldClkCnt[61]), .B0(n1728), .S(n1727), .CO(n1726));
Q_AD01HF U2265 ( .A0(ixcHoldClkCnt[60]), .B0(n1730), .S(n1729), .CO(n1728));
Q_AD01HF U2266 ( .A0(ixcHoldClkCnt[59]), .B0(n1732), .S(n1731), .CO(n1730));
Q_AD01HF U2267 ( .A0(ixcHoldClkCnt[58]), .B0(n1734), .S(n1733), .CO(n1732));
Q_AD01HF U2268 ( .A0(ixcHoldClkCnt[57]), .B0(n1736), .S(n1735), .CO(n1734));
Q_AD01HF U2269 ( .A0(ixcHoldClkCnt[56]), .B0(n1738), .S(n1737), .CO(n1736));
Q_AD01HF U2270 ( .A0(ixcHoldClkCnt[55]), .B0(n1740), .S(n1739), .CO(n1738));
Q_AD01HF U2271 ( .A0(ixcHoldClkCnt[54]), .B0(n1742), .S(n1741), .CO(n1740));
Q_AD01HF U2272 ( .A0(ixcHoldClkCnt[53]), .B0(n1744), .S(n1743), .CO(n1742));
Q_AD01HF U2273 ( .A0(ixcHoldClkCnt[52]), .B0(n1746), .S(n1745), .CO(n1744));
Q_AD01HF U2274 ( .A0(ixcHoldClkCnt[51]), .B0(n1748), .S(n1747), .CO(n1746));
Q_AD01HF U2275 ( .A0(ixcHoldClkCnt[50]), .B0(n1750), .S(n1749), .CO(n1748));
Q_AD01HF U2276 ( .A0(ixcHoldClkCnt[49]), .B0(n1752), .S(n1751), .CO(n1750));
Q_AD01HF U2277 ( .A0(ixcHoldClkCnt[48]), .B0(n1754), .S(n1753), .CO(n1752));
Q_AD01HF U2278 ( .A0(ixcHoldClkCnt[47]), .B0(n1756), .S(n1755), .CO(n1754));
Q_AD01HF U2279 ( .A0(ixcHoldClkCnt[46]), .B0(n1758), .S(n1757), .CO(n1756));
Q_AD01HF U2280 ( .A0(ixcHoldClkCnt[45]), .B0(n1760), .S(n1759), .CO(n1758));
Q_AD01HF U2281 ( .A0(ixcHoldClkCnt[44]), .B0(n1762), .S(n1761), .CO(n1760));
Q_AD01HF U2282 ( .A0(ixcHoldClkCnt[43]), .B0(n1764), .S(n1763), .CO(n1762));
Q_AD01HF U2283 ( .A0(ixcHoldClkCnt[42]), .B0(n1766), .S(n1765), .CO(n1764));
Q_AD01HF U2284 ( .A0(ixcHoldClkCnt[41]), .B0(n1768), .S(n1767), .CO(n1766));
Q_AD01HF U2285 ( .A0(ixcHoldClkCnt[40]), .B0(n1770), .S(n1769), .CO(n1768));
Q_AD01HF U2286 ( .A0(ixcHoldClkCnt[39]), .B0(n1772), .S(n1771), .CO(n1770));
Q_AD01HF U2287 ( .A0(ixcHoldClkCnt[38]), .B0(n1774), .S(n1773), .CO(n1772));
Q_AD01HF U2288 ( .A0(ixcHoldClkCnt[37]), .B0(n1776), .S(n1775), .CO(n1774));
Q_AD01HF U2289 ( .A0(ixcHoldClkCnt[36]), .B0(n1778), .S(n1777), .CO(n1776));
Q_AD01HF U2290 ( .A0(ixcHoldClkCnt[35]), .B0(n1780), .S(n1779), .CO(n1778));
Q_AD01HF U2291 ( .A0(ixcHoldClkCnt[34]), .B0(n1782), .S(n1781), .CO(n1780));
Q_AD01HF U2292 ( .A0(ixcHoldClkCnt[33]), .B0(n1784), .S(n1783), .CO(n1782));
Q_AD01HF U2293 ( .A0(ixcHoldClkCnt[32]), .B0(n1786), .S(n1785), .CO(n1784));
Q_AD01HF U2294 ( .A0(ixcHoldClkCnt[31]), .B0(n1788), .S(n1787), .CO(n1786));
Q_AD01HF U2295 ( .A0(ixcHoldClkCnt[30]), .B0(n1790), .S(n1789), .CO(n1788));
Q_AD01HF U2296 ( .A0(ixcHoldClkCnt[29]), .B0(n1792), .S(n1791), .CO(n1790));
Q_AD01HF U2297 ( .A0(ixcHoldClkCnt[28]), .B0(n1794), .S(n1793), .CO(n1792));
Q_AD01HF U2298 ( .A0(ixcHoldClkCnt[27]), .B0(n1796), .S(n1795), .CO(n1794));
Q_AD01HF U2299 ( .A0(ixcHoldClkCnt[26]), .B0(n1798), .S(n1797), .CO(n1796));
Q_AD01HF U2300 ( .A0(ixcHoldClkCnt[25]), .B0(n1800), .S(n1799), .CO(n1798));
Q_AD01HF U2301 ( .A0(ixcHoldClkCnt[24]), .B0(n1802), .S(n1801), .CO(n1800));
Q_AD01HF U2302 ( .A0(ixcHoldClkCnt[23]), .B0(n1804), .S(n1803), .CO(n1802));
Q_AD01HF U2303 ( .A0(ixcHoldClkCnt[22]), .B0(n1806), .S(n1805), .CO(n1804));
Q_AD01HF U2304 ( .A0(ixcHoldClkCnt[21]), .B0(n1808), .S(n1807), .CO(n1806));
Q_AD01HF U2305 ( .A0(ixcHoldClkCnt[20]), .B0(n1810), .S(n1809), .CO(n1808));
Q_AD01HF U2306 ( .A0(ixcHoldClkCnt[19]), .B0(n1812), .S(n1811), .CO(n1810));
Q_AD01HF U2307 ( .A0(ixcHoldClkCnt[18]), .B0(n1814), .S(n1813), .CO(n1812));
Q_AD01HF U2308 ( .A0(ixcHoldClkCnt[17]), .B0(n1816), .S(n1815), .CO(n1814));
Q_AD01HF U2309 ( .A0(ixcHoldClkCnt[16]), .B0(n1818), .S(n1817), .CO(n1816));
Q_AD01HF U2310 ( .A0(ixcHoldClkCnt[15]), .B0(n1820), .S(n1819), .CO(n1818));
Q_AD01HF U2311 ( .A0(ixcHoldClkCnt[14]), .B0(n1822), .S(n1821), .CO(n1820));
Q_AD01HF U2312 ( .A0(ixcHoldClkCnt[13]), .B0(n1824), .S(n1823), .CO(n1822));
Q_AD01HF U2313 ( .A0(ixcHoldClkCnt[12]), .B0(n1826), .S(n1825), .CO(n1824));
Q_AD01HF U2314 ( .A0(ixcHoldClkCnt[11]), .B0(n1828), .S(n1827), .CO(n1826));
Q_AD01HF U2315 ( .A0(ixcHoldClkCnt[10]), .B0(n1830), .S(n1829), .CO(n1828));
Q_AD01HF U2316 ( .A0(ixcHoldClkCnt[9]), .B0(n1832), .S(n1831), .CO(n1830));
Q_AD01HF U2317 ( .A0(ixcHoldClkCnt[8]), .B0(n1834), .S(n1833), .CO(n1832));
Q_AD01HF U2318 ( .A0(ixcHoldClkCnt[7]), .B0(n1836), .S(n1835), .CO(n1834));
Q_AD01HF U2319 ( .A0(ixcHoldClkCnt[6]), .B0(n1838), .S(n1837), .CO(n1836));
Q_AD01HF U2320 ( .A0(ixcHoldClkCnt[5]), .B0(n1840), .S(n1839), .CO(n1838));
Q_AD01HF U2321 ( .A0(ixcHoldClkCnt[4]), .B0(n1842), .S(n1841), .CO(n1840));
Q_AD01HF U2322 ( .A0(ixcHoldClkCnt[3]), .B0(n1844), .S(n1843), .CO(n1842));
Q_AD01HF U2323 ( .A0(ixcHoldClkCnt[2]), .B0(n1846), .S(n1845), .CO(n1844));
Q_AD01HF U2324 ( .A0(ixcHoldClkCnt[1]), .B0(ixcHoldClkCnt[0]), .S(n1847), .CO(n1846));
Q_XOR2 U2325 ( .A0(nbaCount[63]), .A1(n7), .Z(n1659));
Q_AD01HF U2326 ( .A0(nbaCount[62]), .B0(n1850), .S(n1849), .CO(n1848));
Q_AD01HF U2327 ( .A0(nbaCount[61]), .B0(n1852), .S(n1851), .CO(n1850));
Q_AD01HF U2328 ( .A0(nbaCount[60]), .B0(n1854), .S(n1853), .CO(n1852));
Q_AD01HF U2329 ( .A0(nbaCount[59]), .B0(n1856), .S(n1855), .CO(n1854));
Q_AD01HF U2330 ( .A0(nbaCount[58]), .B0(n1858), .S(n1857), .CO(n1856));
Q_AD01HF U2331 ( .A0(nbaCount[57]), .B0(n1860), .S(n1859), .CO(n1858));
Q_AD01HF U2332 ( .A0(nbaCount[56]), .B0(n1862), .S(n1861), .CO(n1860));
Q_AD01HF U2333 ( .A0(nbaCount[55]), .B0(n1864), .S(n1863), .CO(n1862));
Q_AD01HF U2334 ( .A0(nbaCount[54]), .B0(n1866), .S(n1865), .CO(n1864));
Q_AD01HF U2335 ( .A0(nbaCount[53]), .B0(n1868), .S(n1867), .CO(n1866));
Q_AD01HF U2336 ( .A0(nbaCount[52]), .B0(n1870), .S(n1869), .CO(n1868));
Q_AD01HF U2337 ( .A0(nbaCount[51]), .B0(n1872), .S(n1871), .CO(n1870));
Q_AD01HF U2338 ( .A0(nbaCount[50]), .B0(n1874), .S(n1873), .CO(n1872));
Q_AD01HF U2339 ( .A0(nbaCount[49]), .B0(n1876), .S(n1875), .CO(n1874));
Q_AD01HF U2340 ( .A0(nbaCount[48]), .B0(n1878), .S(n1877), .CO(n1876));
Q_AD01HF U2341 ( .A0(nbaCount[47]), .B0(n1880), .S(n1879), .CO(n1878));
Q_AD01HF U2342 ( .A0(nbaCount[46]), .B0(n1882), .S(n1881), .CO(n1880));
Q_AD01HF U2343 ( .A0(nbaCount[45]), .B0(n1884), .S(n1883), .CO(n1882));
Q_AD01HF U2344 ( .A0(nbaCount[44]), .B0(n1886), .S(n1885), .CO(n1884));
Q_AD01HF U2345 ( .A0(nbaCount[43]), .B0(n1888), .S(n1887), .CO(n1886));
Q_AD01HF U2346 ( .A0(nbaCount[42]), .B0(n1890), .S(n1889), .CO(n1888));
Q_AD01HF U2347 ( .A0(nbaCount[41]), .B0(n1892), .S(n1891), .CO(n1890));
Q_AD01HF U2348 ( .A0(nbaCount[40]), .B0(n1894), .S(n1893), .CO(n1892));
Q_AD01HF U2349 ( .A0(nbaCount[39]), .B0(n1896), .S(n1895), .CO(n1894));
Q_AD01HF U2350 ( .A0(nbaCount[38]), .B0(n1898), .S(n1897), .CO(n1896));
Q_AD01HF U2351 ( .A0(nbaCount[37]), .B0(n1900), .S(n1899), .CO(n1898));
Q_AD01HF U2352 ( .A0(nbaCount[36]), .B0(n1902), .S(n1901), .CO(n1900));
Q_AD01HF U2353 ( .A0(nbaCount[35]), .B0(n1904), .S(n1903), .CO(n1902));
Q_AD01HF U2354 ( .A0(nbaCount[34]), .B0(n1906), .S(n1905), .CO(n1904));
Q_AD01HF U2355 ( .A0(nbaCount[33]), .B0(n1908), .S(n1907), .CO(n1906));
Q_AD01HF U2356 ( .A0(nbaCount[32]), .B0(n1910), .S(n1909), .CO(n1908));
Q_AD01HF U2357 ( .A0(nbaCount[31]), .B0(n1912), .S(n1911), .CO(n1910));
Q_AD01HF U2358 ( .A0(nbaCount[30]), .B0(n1914), .S(n1913), .CO(n1912));
Q_AD01HF U2359 ( .A0(nbaCount[29]), .B0(n1916), .S(n1915), .CO(n1914));
Q_AD01HF U2360 ( .A0(nbaCount[28]), .B0(n1918), .S(n1917), .CO(n1916));
Q_AD01HF U2361 ( .A0(nbaCount[27]), .B0(n1920), .S(n1919), .CO(n1918));
Q_AD01HF U2362 ( .A0(nbaCount[26]), .B0(n1922), .S(n1921), .CO(n1920));
Q_AD01HF U2363 ( .A0(nbaCount[25]), .B0(n1924), .S(n1923), .CO(n1922));
Q_AD01HF U2364 ( .A0(nbaCount[24]), .B0(n1926), .S(n1925), .CO(n1924));
Q_AD01HF U2365 ( .A0(nbaCount[23]), .B0(n1928), .S(n1927), .CO(n1926));
Q_AD01HF U2366 ( .A0(nbaCount[22]), .B0(n1930), .S(n1929), .CO(n1928));
Q_AD01HF U2367 ( .A0(nbaCount[21]), .B0(n1932), .S(n1931), .CO(n1930));
Q_AD01HF U2368 ( .A0(nbaCount[20]), .B0(n1934), .S(n1933), .CO(n1932));
Q_AD01HF U2369 ( .A0(nbaCount[19]), .B0(n1936), .S(n1935), .CO(n1934));
Q_AD01HF U2370 ( .A0(nbaCount[18]), .B0(n1938), .S(n1937), .CO(n1936));
Q_AD01HF U2371 ( .A0(nbaCount[17]), .B0(n1940), .S(n1939), .CO(n1938));
Q_AD01HF U2372 ( .A0(nbaCount[16]), .B0(n1942), .S(n1941), .CO(n1940));
Q_AD01HF U2373 ( .A0(nbaCount[15]), .B0(n1944), .S(n1943), .CO(n1942));
Q_AD01HF U2374 ( .A0(nbaCount[14]), .B0(n1946), .S(n1945), .CO(n1944));
Q_AD01HF U2375 ( .A0(nbaCount[13]), .B0(n1948), .S(n1947), .CO(n1946));
Q_AD01HF U2376 ( .A0(nbaCount[12]), .B0(n1950), .S(n1949), .CO(n1948));
Q_AD01HF U2377 ( .A0(nbaCount[11]), .B0(n1952), .S(n1951), .CO(n1950));
Q_AD01HF U2378 ( .A0(nbaCount[10]), .B0(n1954), .S(n1953), .CO(n1952));
Q_AD01HF U2379 ( .A0(nbaCount[9]), .B0(n1956), .S(n1955), .CO(n1954));
Q_AD01HF U2380 ( .A0(nbaCount[8]), .B0(n1958), .S(n1957), .CO(n1956));
Q_AD01HF U2381 ( .A0(nbaCount[7]), .B0(n1960), .S(n1959), .CO(n1958));
Q_AD01HF U2382 ( .A0(nbaCount[6]), .B0(n1962), .S(n1961), .CO(n1960));
Q_AD01HF U2383 ( .A0(nbaCount[5]), .B0(n1964), .S(n1963), .CO(n1962));
Q_AD01HF U2384 ( .A0(nbaCount[4]), .B0(n1966), .S(n1965), .CO(n1964));
Q_AD01HF U2385 ( .A0(nbaCount[3]), .B0(n1968), .S(n1967), .CO(n1966));
Q_AD01HF U2386 ( .A0(nbaCount[2]), .B0(n1970), .S(n1969), .CO(n1968));
Q_AD01HF U2387 ( .A0(nbaCount[1]), .B0(nbaCount[0]), .S(n1971), .CO(n1970));
Q_XOR2 U2388 ( .A0(bCount[63]), .A1(n6), .Z(n1723));
Q_AD01HF U2389 ( .A0(bCount[62]), .B0(n1974), .S(n1973), .CO(n1972));
Q_AD01HF U2390 ( .A0(bCount[61]), .B0(n1976), .S(n1975), .CO(n1974));
Q_AD01HF U2391 ( .A0(bCount[60]), .B0(n1978), .S(n1977), .CO(n1976));
Q_AD01HF U2392 ( .A0(bCount[59]), .B0(n1980), .S(n1979), .CO(n1978));
Q_AD01HF U2393 ( .A0(bCount[58]), .B0(n1982), .S(n1981), .CO(n1980));
Q_AD01HF U2394 ( .A0(bCount[57]), .B0(n1984), .S(n1983), .CO(n1982));
Q_AD01HF U2395 ( .A0(bCount[56]), .B0(n1986), .S(n1985), .CO(n1984));
Q_AD01HF U2396 ( .A0(bCount[55]), .B0(n1988), .S(n1987), .CO(n1986));
Q_AD01HF U2397 ( .A0(bCount[54]), .B0(n1990), .S(n1989), .CO(n1988));
Q_AD01HF U2398 ( .A0(bCount[53]), .B0(n1992), .S(n1991), .CO(n1990));
Q_AD01HF U2399 ( .A0(bCount[52]), .B0(n1994), .S(n1993), .CO(n1992));
Q_AD01HF U2400 ( .A0(bCount[51]), .B0(n1996), .S(n1995), .CO(n1994));
Q_AD01HF U2401 ( .A0(bCount[50]), .B0(n1998), .S(n1997), .CO(n1996));
Q_AD01HF U2402 ( .A0(bCount[49]), .B0(n2000), .S(n1999), .CO(n1998));
Q_AD01HF U2403 ( .A0(bCount[48]), .B0(n2002), .S(n2001), .CO(n2000));
Q_AD01HF U2404 ( .A0(bCount[47]), .B0(n2004), .S(n2003), .CO(n2002));
Q_AD01HF U2405 ( .A0(bCount[46]), .B0(n2006), .S(n2005), .CO(n2004));
Q_AD01HF U2406 ( .A0(bCount[45]), .B0(n2008), .S(n2007), .CO(n2006));
Q_AD01HF U2407 ( .A0(bCount[44]), .B0(n2010), .S(n2009), .CO(n2008));
Q_AD01HF U2408 ( .A0(bCount[43]), .B0(n2012), .S(n2011), .CO(n2010));
Q_AD01HF U2409 ( .A0(bCount[42]), .B0(n2014), .S(n2013), .CO(n2012));
Q_AD01HF U2410 ( .A0(bCount[41]), .B0(n2016), .S(n2015), .CO(n2014));
Q_AD01HF U2411 ( .A0(bCount[40]), .B0(n2018), .S(n2017), .CO(n2016));
Q_AD01HF U2412 ( .A0(bCount[39]), .B0(n2020), .S(n2019), .CO(n2018));
Q_AD01HF U2413 ( .A0(bCount[38]), .B0(n2022), .S(n2021), .CO(n2020));
Q_AD01HF U2414 ( .A0(bCount[37]), .B0(n2024), .S(n2023), .CO(n2022));
Q_AD01HF U2415 ( .A0(bCount[36]), .B0(n2026), .S(n2025), .CO(n2024));
Q_AD01HF U2416 ( .A0(bCount[35]), .B0(n2028), .S(n2027), .CO(n2026));
Q_AD01HF U2417 ( .A0(bCount[34]), .B0(n2030), .S(n2029), .CO(n2028));
Q_AD01HF U2418 ( .A0(bCount[33]), .B0(n2032), .S(n2031), .CO(n2030));
Q_AD01HF U2419 ( .A0(bCount[32]), .B0(n2034), .S(n2033), .CO(n2032));
Q_AD01HF U2420 ( .A0(bCount[31]), .B0(n2036), .S(n2035), .CO(n2034));
Q_AD01HF U2421 ( .A0(bCount[30]), .B0(n2038), .S(n2037), .CO(n2036));
Q_AD01HF U2422 ( .A0(bCount[29]), .B0(n2040), .S(n2039), .CO(n2038));
Q_AD01HF U2423 ( .A0(bCount[28]), .B0(n2042), .S(n2041), .CO(n2040));
Q_AD01HF U2424 ( .A0(bCount[27]), .B0(n2044), .S(n2043), .CO(n2042));
Q_AD01HF U2425 ( .A0(bCount[26]), .B0(n2046), .S(n2045), .CO(n2044));
Q_AD01HF U2426 ( .A0(bCount[25]), .B0(n2048), .S(n2047), .CO(n2046));
Q_AD01HF U2427 ( .A0(bCount[24]), .B0(n2050), .S(n2049), .CO(n2048));
Q_AD01HF U2428 ( .A0(bCount[23]), .B0(n2052), .S(n2051), .CO(n2050));
Q_AD01HF U2429 ( .A0(bCount[22]), .B0(n2054), .S(n2053), .CO(n2052));
Q_AD01HF U2430 ( .A0(bCount[21]), .B0(n2056), .S(n2055), .CO(n2054));
Q_AD01HF U2431 ( .A0(bCount[20]), .B0(n2058), .S(n2057), .CO(n2056));
Q_AD01HF U2432 ( .A0(bCount[19]), .B0(n2060), .S(n2059), .CO(n2058));
Q_AD01HF U2433 ( .A0(bCount[18]), .B0(n2062), .S(n2061), .CO(n2060));
Q_AD01HF U2434 ( .A0(bCount[17]), .B0(n2064), .S(n2063), .CO(n2062));
Q_AD01HF U2435 ( .A0(bCount[16]), .B0(n2066), .S(n2065), .CO(n2064));
Q_AD01HF U2436 ( .A0(bCount[15]), .B0(n2068), .S(n2067), .CO(n2066));
Q_AD01HF U2437 ( .A0(bCount[14]), .B0(n2070), .S(n2069), .CO(n2068));
Q_AD01HF U2438 ( .A0(bCount[13]), .B0(n2072), .S(n2071), .CO(n2070));
Q_AD01HF U2439 ( .A0(bCount[12]), .B0(n2074), .S(n2073), .CO(n2072));
Q_AD01HF U2440 ( .A0(bCount[11]), .B0(n2076), .S(n2075), .CO(n2074));
Q_AD01HF U2441 ( .A0(bCount[10]), .B0(n2078), .S(n2077), .CO(n2076));
Q_AD01HF U2442 ( .A0(bCount[9]), .B0(n2080), .S(n2079), .CO(n2078));
Q_AD01HF U2443 ( .A0(bCount[8]), .B0(n2082), .S(n2081), .CO(n2080));
Q_AD01HF U2444 ( .A0(bCount[7]), .B0(n2084), .S(n2083), .CO(n2082));
Q_AD01HF U2445 ( .A0(bCount[6]), .B0(n2086), .S(n2085), .CO(n2084));
Q_AD01HF U2446 ( .A0(bCount[5]), .B0(n2088), .S(n2087), .CO(n2086));
Q_AD01HF U2447 ( .A0(bCount[4]), .B0(n2090), .S(n2089), .CO(n2088));
Q_AD01HF U2448 ( .A0(bCount[3]), .B0(n2092), .S(n2091), .CO(n2090));
Q_AD01HF U2449 ( .A0(bCount[2]), .B0(n2094), .S(n2093), .CO(n2092));
Q_AD01HF U2450 ( .A0(bCount[1]), .B0(bCount[0]), .S(n2095), .CO(n2094));
Q_OR02 U2451 ( .A0(bpWait), .A1(bpSt[1]), .Z(n2097));
Q_OR02 U2452 ( .A0(bpSt[1]), .A1(mpOn), .Z(n2106));
Q_INV U2453 ( .A(bpSt[1]), .Z(n2107));
Q_OR02 U2454 ( .A0(sampleXpChg), .A1(n2096), .Z(n2108));
Q_AN02 U2455 ( .A0(mpOn), .A1(sampleXpChg), .Z(n2109));
Q_INV U2456 ( .A(n2109), .Z(n2098));
Q_OA21 U2457 ( .A0(n2098), .A1(bpSt[1]), .B0(n2110), .Z(n2099));
Q_INV U2458 ( .A(n2099), .Z(n2100));
Q_MX02 U2459 ( .S(bpWait), .A0(n2100), .A1(n2106), .Z(n2101));
Q_INV U2460 ( .A(n2101), .Z(n2102));
Q_MX02 U2461 ( .S(bpSt[0]), .A0(n2102), .A1(n2097), .Z(n2103));
Q_INV U2462 ( .A(n2108), .Z(n2116));
Q_OR02 U2463 ( .A0(bpSt[1]), .A1(n2116), .Z(n2104));
Q_MX02 U2464 ( .S(bpWait), .A0(n2104), .A1(bpSt[1]), .Z(n2105));
Q_OR02 U2465 ( .A0(n2108), .A1(n2107), .Z(n2110));
Q_OA21 U2466 ( .A0(n2109), .A1(bpSt[1]), .B0(n2110), .Z(n2111));
Q_MX02 U2467 ( .S(bpWait), .A0(n2111), .A1(n2106), .Z(n2112));
Q_INV U2468 ( .A(n2112), .Z(n2113));
Q_MX02 U2469 ( .S(bpSt[0]), .A0(n2113), .A1(n2105), .Z(n2114));
Q_OR02 U2470 ( .A0(bClkHold), .A1(n2114), .Z(n2115));
Q_NR02 U2471 ( .A0(bpWait), .A1(n2116), .Z(n2117));
Q_MX02 U2472 ( .S(n2103), .A0(bpWait), .A1(bpSt[0]), .Z(n2118));
Q_FDP0UA U2473 ( .D(n2118), .QTFCLK( ), .Q(bpSt[0]));
Q_MX02 U2474 ( .S(n2103), .A0(n2117), .A1(bpSt[1]), .Z(n2119));
Q_FDP0UA U2475 ( .D(n2119), .QTFCLK( ), .Q(bpSt[1]));
Q_XNR2 U2476 ( .A0(n2115), .A1(bClkR), .Z(n2120));
Q_FDP0UA U2477 ( .D(n2120), .QTFCLK( ), .Q(bClkR));
Q_INV U2478 ( .A(n2121), .Z(n2096));
Q_XNR2 U2479 ( .A0(uClk), .A1(clockMC), .Z(n2121));
Q_FDP0UA U2480 ( .D(bClkHold), .QTFCLK( ), .Q(bClkHoldD));
Q_FDP0UA U2481 ( .D(holdEcm), .QTFCLK( ), .Q(holdEcmD));
Q_FDP0UA U2482 ( .D(tbcPOStateN[1]), .QTFCLK( ), .Q(tbcPOState[1]));
Q_FDP0UA U2483 ( .D(tbcPOStateN[0]), .QTFCLK( ), .Q(tbcPOState[0]));
Q_INV U2484 ( .A(GF2LevelMask[0]), .Z(n2122));
Q_INV U2485 ( .A(GF2LevelMask[1]), .Z(n2123));
Q_INV U2486 ( .A(GF2LevelMask[2]), .Z(n2124));
Q_INV U2487 ( .A(GF2LevelMask[3]), .Z(n2125));
Q_INV U2488 ( .A(GF2LevelMask[4]), .Z(n2126));
Q_INV U2489 ( .A(GF2LevelMask[5]), .Z(n2127));
Q_INV U2490 ( .A(GF2LevelMask[6]), .Z(n2128));
Q_INV U2491 ( .A(GF2LevelMask[7]), .Z(n2129));
Q_INV U2492 ( .A(GF2LevelMask[8]), .Z(n2130));
Q_INV U2493 ( .A(GF2LevelMask[9]), .Z(n2131));
Q_INV U2494 ( .A(GF2LevelMask[10]), .Z(n2132));
Q_INV U2495 ( .A(GF2LevelMask[11]), .Z(n2133));
Q_INV U2496 ( .A(GF2LevelMask[12]), .Z(n2134));
Q_OR02 U2497 ( .A0(tbcPOd), .A1(n2122), .Z(n2135));
Q_OR02 U2498 ( .A0(tbcPODly[0]), .A1(n2123), .Z(n2136));
Q_OR02 U2499 ( .A0(tbcPODly[1]), .A1(n2124), .Z(n2137));
Q_OR02 U2500 ( .A0(tbcPODly[2]), .A1(n2125), .Z(n2138));
Q_OR02 U2501 ( .A0(tbcPODly[3]), .A1(n2126), .Z(n2139));
Q_OR02 U2502 ( .A0(tbcPODly[4]), .A1(n2127), .Z(n2140));
Q_OR02 U2503 ( .A0(tbcPODly[5]), .A1(n2128), .Z(n2141));
Q_OR02 U2504 ( .A0(tbcPODly[6]), .A1(n2129), .Z(n2142));
Q_OR02 U2505 ( .A0(tbcPODly[7]), .A1(n2130), .Z(n2143));
Q_OR02 U2506 ( .A0(tbcPODly[8]), .A1(n2131), .Z(n2144));
Q_OR02 U2507 ( .A0(tbcPODly[9]), .A1(n2132), .Z(n2145));
Q_OR02 U2508 ( .A0(tbcPODly[10]), .A1(n2133), .Z(n2146));
Q_OR02 U2509 ( .A0(tbcPODly[11]), .A1(n2134), .Z(n2147));
Q_FDP0UA U2510 ( .D(n2147), .QTFCLK( ), .Q(tbcPODly[12]));
Q_FDP0UA U2511 ( .D(n2146), .QTFCLK( ), .Q(tbcPODly[11]));
Q_FDP0UA U2512 ( .D(n2145), .QTFCLK( ), .Q(tbcPODly[10]));
Q_FDP0UA U2513 ( .D(n2144), .QTFCLK( ), .Q(tbcPODly[9]));
Q_FDP0UA U2514 ( .D(n2143), .QTFCLK( ), .Q(tbcPODly[8]));
Q_FDP0UA U2515 ( .D(n2142), .QTFCLK( ), .Q(tbcPODly[7]));
Q_FDP0UA U2516 ( .D(n2141), .QTFCLK( ), .Q(tbcPODly[6]));
Q_FDP0UA U2517 ( .D(n2140), .QTFCLK( ), .Q(tbcPODly[5]));
Q_FDP0UA U2518 ( .D(n2139), .QTFCLK( ), .Q(tbcPODly[4]));
Q_FDP0UA U2519 ( .D(n2138), .QTFCLK( ), .Q(tbcPODly[3]));
Q_FDP0UA U2520 ( .D(n2137), .QTFCLK( ), .Q(tbcPODly[2]));
Q_FDP0UA U2521 ( .D(n2136), .QTFCLK( ), .Q(tbcPODly[1]));
Q_FDP0UA U2522 ( .D(n2135), .QTFCLK( ), .Q(tbcPODly[0]));
Q_FDP0UA U2523 ( .D(GFbusyD), .QTFCLK( ), .Q(GFbusyD2));
Q_FDP0UA U2524 ( .D(GFbusy), .QTFCLK( ), .Q(GFbusyD));
Q_INV U2525 ( .A(mpSt[2]), .Z(n2149));
Q_AN03 U2526 ( .A0(n2149), .A1(mpSt[1]), .A2(mpSt[0]), .Z(n2150));
Q_OR02 U2527 ( .A0(n2150), .A1(asyncBusy), .Z(n2148));
Q_MX02 U2528 ( .S(n2148), .A0(asyncBusy), .A1(n1429), .Z(n2151));
Q_FDP0UA U2529 ( .D(n2151), .QTFCLK( ), .Q(asyncBusy));
Q_INV U2530 ( .A(mpSt[1]), .Z(n2161));
Q_NR02 U2531 ( .A0(mpSt[1]), .A1(callEmu), .Z(n2164));
Q_INV U2532 ( .A(stopCond), .Z(n2197));
Q_AN02 U2533 ( .A0(mpSt[1]), .A1(n2197), .Z(n2179));
Q_OA21 U2534 ( .A0(n2164), .A1(n2179), .B0(n2191), .Z(n2167));
Q_INV U2535 ( .A(mpEnable), .Z(n2186));
Q_OA21 U2536 ( .A0(n2186), .A1(bpHalt), .B0(n2165), .Z(n2166));
Q_NR02 U2537 ( .A0(mpEnable), .A1(bpHalt), .Z(n2176));
Q_INV U2538 ( .A(stopEmuPO), .Z(n2165));
Q_OR02 U2539 ( .A0(n2176), .A1(n2166), .Z(n2182));
Q_INV U2540 ( .A(mpSt[0]), .Z(n2191));
Q_AN02 U2541 ( .A0(mpSt[1]), .A1(mpSt[0]), .Z(n2188));
Q_AO21 U2542 ( .A0(n2182), .A1(n2188), .B0(n2168), .Z(n2169));
Q_OR02 U2543 ( .A0(n2167), .A1(mpSt[2]), .Z(n2168));
Q_AN02 U2544 ( .A0(callEmu), .A1(n2121), .Z(n2170));
Q_OR02 U2545 ( .A0(mpSt[0]), .A1(n2170), .Z(n2196));
Q_NR02 U2546 ( .A0(mpSt[2]), .A1(mpSt[1]), .Z(n2172));
Q_INV U2547 ( .A(gfifoOff), .Z(n2171));
Q_AN02 U2548 ( .A0(n2172), .A1(n2171), .Z(n2173));
Q_AO21 U2549 ( .A0(n2173), .A1(n2196), .B0(initClock), .Z(n2209));
Q_AN02 U2550 ( .A0(n2197), .A1(mpEnable), .Z(n2192));
Q_OA21 U2551 ( .A0(n2192), .A1(mpSt[0]), .B0(mpSt[1]), .Z(n2175));
Q_AN03 U2552 ( .A0(n2161), .A1(callEmu), .A2(n2121), .Z(n2180));
Q_OA21 U2553 ( .A0(mpSt[0]), .A1(n2180), .B0(n2189), .Z(n2174));
Q_INV U2554 ( .A(ckgHoldPIi), .Z(n2189));
Q_OA21 U2555 ( .A0(n2175), .A1(n2174), .B0(n2149), .Z(n2152));
Q_INV U2556 ( .A(n2176), .Z(n2177));
Q_AN03 U2557 ( .A0(n2191), .A1(callEmu), .A2(n2161), .Z(n2184));
Q_AO21 U2558 ( .A0(n2177), .A1(n2188), .B0(n2184), .Z(n2178));
Q_AN02 U2559 ( .A0(n2149), .A1(n2178), .Z(n2153));
Q_OR03 U2560 ( .A0(n2179), .A1(mpSt[0]), .A2(n2180), .Z(n2181));
Q_AN02 U2561 ( .A0(n2149), .A1(n2181), .Z(n2154));
Q_INV U2562 ( .A(n2182), .Z(n2183));
Q_AO21 U2563 ( .A0(n2183), .A1(n2188), .B0(n2184), .Z(n2185));
Q_AN02 U2564 ( .A0(n2149), .A1(n2185), .Z(n2155));
Q_NR02 U2565 ( .A0(mpSt[1]), .A1(mpSt[0]), .Z(n2158));
Q_INV U2566 ( .A(n2158), .Z(n2156));
Q_OA21 U2567 ( .A0(n2186), .A1(mpSt[0]), .B0(mpSt[1]), .Z(n2187));
Q_INV U2568 ( .A(n2187), .Z(n2157));
Q_INV U2569 ( .A(n2188), .Z(n2159));
Q_NR02 U2570 ( .A0(mpSt[1]), .A1(ckgHoldPIi), .Z(n2190));
Q_AN02 U2571 ( .A0(n2196), .A1(n2190), .Z(n2193));
Q_AN02 U2572 ( .A0(mpSt[1]), .A1(n2191), .Z(n2198));
Q_AO21 U2573 ( .A0(n2198), .A1(n2192), .B0(n2193), .Z(n2194));
Q_AN02 U2574 ( .A0(n2149), .A1(n2194), .Z(n2160));
Q_OA21 U2575 ( .A0(n2121), .A1(mpSt[0]), .B0(n2161), .Z(n2195));
Q_OR02 U2576 ( .A0(n2198), .A1(n2195), .Z(n2162));
Q_AN02 U2577 ( .A0(n2196), .A1(n2161), .Z(n2199));
Q_AO21 U2578 ( .A0(n2198), .A1(n2197), .B0(n2199), .Z(n2200));
Q_AN02 U2579 ( .A0(n2149), .A1(n2200), .Z(n2163));
Q_FDP0UA U2580 ( .D(n2163), .QTFCLK( ), .Q(active));
Q_MX02 U2581 ( .S(n2169), .A0(n2208), .A1(mpSt[0]), .Z(n2201));
Q_FDP0UA U2582 ( .D(n2201), .QTFCLK( ), .Q(mpSt[0]));
Q_MX02 U2583 ( .S(n2169), .A0(n2162), .A1(mpSt[1]), .Z(n2202));
Q_FDP0UA U2584 ( .D(n2202), .QTFCLK( ), .Q(mpSt[1]));
Q_AN02 U2585 ( .A0(n2169), .A1(mpSt[2]), .Z(n2203));
Q_FDP0UA U2586 ( .D(n2203), .QTFCLK( ), .Q(mpSt[2]));
Q_FDP0UA U2587 ( .D(n2160), .QTFCLK( ), .Q(lbrOn));
Q_MX02 U2588 ( .S(n2152), .A0(simTimeOn), .A1(n2159), .Z(n2204));
Q_FDP0UA U2589 ( .D(n2204), .QTFCLK( ), .Q(simTimeOn));
Q_MX02 U2590 ( .S(n2153), .A0(evalOnC), .A1(n2158), .Z(n2205));
Q_FDP0UA U2591 ( .D(n2205), .QTFCLK( ), .Q(evalOnC));
Q_MX02 U2592 ( .S(n2154), .A0(mpOn), .A1(n2157), .Z(n2206));
Q_FDP0UA U2593 ( .D(n2206), .QTFCLK( ), .Q(mpOn));
Q_MX02 U2594 ( .S(n2155), .A0(tbcPOd), .A1(n2156), .Z(n2207));
Q_FDP0UA U2595 ( .D(n2207), .QTFCLK( ), .Q(tbcPOd));
Q_XNR2 U2596 ( .A0(n2162), .A1(mpSt[1]), .Z(n2208));
Q_FDP0UA U2597 ( .D(n2209), .QTFCLK( ), .Q(initClock));
Q_FDP0UA U2598 ( .D(n2210), .QTFCLK( ), .Q(eClkR));
Q_XOR2 U2599 ( .A0(simTimeEnable), .A1(eClkR), .Z(n2210));
Q_INV U2600 ( .A(hotSwapOnPI), .Z(n2211));
Q_NR02 U2601 ( .A0(hotSwapOnPI), .A1(cakeCcEnable), .Z(n2212));
Q_MX02 U2602 ( .S(n2212), .A0(n2214), .A1(clockMC), .Z(n2213));
Q_FDP0UA U2603 ( .D(n2213), .QTFCLK( ), .Q(clockMC));
Q_MX02 U2604 ( .S(hotSwapOnPI), .A0(n2215), .A1(clockMCInit), .Z(n2214));
Q_INV U2605 ( .A(clockMC), .Z(n2215));
Q_NR02 U2606 ( .A0(n2217), .A1(n2216), .Z(n2218));
Q_FDP0UA U2607 ( .D(evalOnInt), .QTFCLK( ), .Q(evalOnIntR[0]));
Q_FDP0UA U2608 ( .D(evalOnIntR[0]), .QTFCLK( ), .Q(evalOnIntR[1]));
Q_FDP0UA U2609 ( .D(evalOnIntR[1]), .QTFCLK( ), .Q(evalOnIntR[2]));
Q_FDP0UA U2610 ( .D(n2217), .QTFCLK( ), .Q(evalOnIntD));
Q_MX02 U2611 ( .S(n2218), .A0(n2234), .A1(evalOnDExt[0]), .Z(n2219));
Q_FDP0UA U2612 ( .D(n2219), .QTFCLK( ), .Q(evalOnDExt[0]));
Q_MX02 U2613 ( .S(n2218), .A0(n2233), .A1(evalOnDExt[1]), .Z(n2220));
Q_FDP0UA U2614 ( .D(n2220), .QTFCLK( ), .Q(evalOnDExt[1]));
Q_MX02 U2615 ( .S(n2218), .A0(n2232), .A1(evalOnDExt[2]), .Z(n2221));
Q_FDP0UA U2616 ( .D(n2221), .QTFCLK( ), .Q(evalOnDExt[2]));
Q_MX02 U2617 ( .S(n2218), .A0(n2231), .A1(evalOnDExt[3]), .Z(n2222));
Q_FDP0UA U2618 ( .D(n2222), .QTFCLK( ), .Q(evalOnDExt[3]));
Q_MX02 U2619 ( .S(n2218), .A0(n2230), .A1(evalOnDExt[4]), .Z(n2223));
Q_FDP0UA U2620 ( .D(n2223), .QTFCLK( ), .Q(evalOnDExt[4]));
Q_MX02 U2621 ( .S(n2218), .A0(n2229), .A1(evalOnDExt[5]), .Z(n2224));
Q_FDP0UA U2622 ( .D(n2224), .QTFCLK( ), .Q(evalOnDExt[5]));
Q_MX02 U2623 ( .S(n2218), .A0(n2228), .A1(evalOnDExt[6]), .Z(n2225));
Q_FDP0UA U2624 ( .D(n2225), .QTFCLK( ), .Q(evalOnDExt[6]));
Q_MX02 U2625 ( .S(n2218), .A0(n2227), .A1(evalOnDExt[7]), .Z(n2226));
Q_FDP0UA U2626 ( .D(n2226), .QTFCLK( ), .Q(evalOnDExt[7]));
Q_MX02 U2627 ( .S(n2217), .A0(n2235), .A1(evalOnDCtl[7]), .Z(n2227));
Q_MX02 U2628 ( .S(n2217), .A0(n2237), .A1(evalOnDCtl[6]), .Z(n2228));
Q_MX02 U2629 ( .S(n2217), .A0(n2239), .A1(evalOnDCtl[5]), .Z(n2229));
Q_MX02 U2630 ( .S(n2217), .A0(n2241), .A1(evalOnDCtl[4]), .Z(n2230));
Q_MX02 U2631 ( .S(n2217), .A0(n2243), .A1(evalOnDCtl[3]), .Z(n2231));
Q_MX02 U2632 ( .S(n2217), .A0(n2245), .A1(evalOnDCtl[2]), .Z(n2232));
Q_MX02 U2633 ( .S(n2217), .A0(n2247), .A1(evalOnDCtl[1]), .Z(n2233));
Q_MX02 U2634 ( .S(n2217), .A0(n2248), .A1(evalOnDCtl[0]), .Z(n2234));
Q_XNR2 U2635 ( .A0(evalOnDExt[7]), .A1(n2236), .Z(n2235));
Q_OR02 U2636 ( .A0(evalOnDExt[6]), .A1(n2238), .Z(n2236));
Q_XNR2 U2637 ( .A0(evalOnDExt[6]), .A1(n2238), .Z(n2237));
Q_OR02 U2638 ( .A0(evalOnDExt[5]), .A1(n2240), .Z(n2238));
Q_XNR2 U2639 ( .A0(evalOnDExt[5]), .A1(n2240), .Z(n2239));
Q_OR02 U2640 ( .A0(evalOnDExt[4]), .A1(n2242), .Z(n2240));
Q_XNR2 U2641 ( .A0(evalOnDExt[4]), .A1(n2242), .Z(n2241));
Q_OR02 U2642 ( .A0(evalOnDExt[3]), .A1(n2244), .Z(n2242));
Q_XNR2 U2643 ( .A0(evalOnDExt[3]), .A1(n2244), .Z(n2243));
Q_OR02 U2644 ( .A0(evalOnDExt[2]), .A1(n2246), .Z(n2244));
Q_XNR2 U2645 ( .A0(evalOnDExt[2]), .A1(n2246), .Z(n2245));
Q_OR02 U2646 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .Z(n2246));
Q_XNR2 U2647 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .Z(n2247));
Q_INV U2648 ( .A(evalOnDExt[0]), .Z(n2248));
Q_OR03 U2649 ( .A0(evalOnInt), .A1(evalOnIntR[0]), .A2(evalOnIntR[1]), .Z(n2217));
Q_OR02 U2650 ( .A0(n2250), .A1(n2249), .Z(n2216));
Q_OR03 U2651 ( .A0(evalOnDExt[1]), .A1(evalOnDExt[0]), .A2(n2251), .Z(n2249));
Q_OR03 U2652 ( .A0(evalOnDExt[4]), .A1(evalOnDExt[3]), .A2(evalOnDExt[2]), .Z(n2250));
Q_OR03 U2653 ( .A0(evalOnDExt[7]), .A1(evalOnDExt[6]), .A2(evalOnDExt[5]), .Z(n2251));
Q_FDP0UA U2654 ( .D(evalOnC), .QTFCLK( ), .Q(evalOnD));
Q_FDP0UA U2655 ( .D(stopTL), .QTFCLK( ), .Q(stopTLd));
Q_FDP0UA U2656 ( .D(mioPOW_2[4]), .QTFCLK( ), .Q(stop3POd));
Q_FDP0UA U2657 ( .D(mioPOW_2[5]), .QTFCLK( ), .Q(stop4POd));
Q_FDP0UA U2658 ( .D(mioPOW_2[3]), .QTFCLK( ), .Q(stop2POd));
Q_FDP0UA U2659 ( .D(mioPOW_2[2]), .QTFCLK( ), .Q(stop1POd));
Q_FDP0UA U2660 ( .D(sdlStopRply), .QTFCLK( ), .Q(sdlStopRplyD));
Q_INV U2661 ( .A(hasGFIFO2), .Z(n2253));
Q_NR02 U2662 ( .A0(hasGFIFO1), .A1(hasGFIFO2), .Z(n2254));
Q_INV U2663 ( .A(n2254), .Z(n2252));
Q_MX02 U2664 ( .S(n2254), .A0(GFAck), .A1(gfifoAckWait[0]), .Z(n2255));
Q_FDP0UA U2665 ( .D(n2255), .QTFCLK( ), .Q(gfifoAckWait[0]));
Q_MX02 U2666 ( .S(n2254), .A0(gfifoAckWait[0]), .A1(gfifoAckWait[1]), .Z(n2256));
Q_FDP0UA U2667 ( .D(n2256), .QTFCLK( ), .Q(gfifoAckWait[1]));
Q_MX02 U2668 ( .S(n2254), .A0(gfifoAckWait[1]), .A1(gfifoAckWait[2]), .Z(n2257));
Q_FDP0UA U2669 ( .D(n2257), .QTFCLK( ), .Q(gfifoAckWait[2]));
Q_MX02 U2670 ( .S(n2254), .A0(gfifoAckWait[2]), .A1(gfifoAckWait[3]), .Z(n2258));
Q_FDP0UA U2671 ( .D(n2258), .QTFCLK( ), .Q(gfifoAckWait[3]));
Q_MX02 U2672 ( .S(n2254), .A0(gfifoAckWait[3]), .A1(gfifoAckWait[4]), .Z(n2259));
Q_FDP0UA U2673 ( .D(n2259), .QTFCLK( ), .Q(gfifoAckWait[4]));
Q_MX02 U2674 ( .S(n2254), .A0(gfifoAckWait[4]), .A1(gfifoAckWait[5]), .Z(n2260));
Q_FDP0UA U2675 ( .D(n2260), .QTFCLK( ), .Q(gfifoAckWait[5]));
Q_MX02 U2676 ( .S(n2254), .A0(gfifoAckWait[5]), .A1(gfifoAckWait[6]), .Z(n2261));
Q_FDP0UA U2677 ( .D(n2261), .QTFCLK( ), .Q(gfifoAckWait[6]));
Q_MX02 U2678 ( .S(n2254), .A0(gfifoAckWait[6]), .A1(gfifoAckWait[7]), .Z(n2262));
Q_FDP0UA U2679 ( .D(n2262), .QTFCLK( ), .Q(gfifoAckWait[7]));
Q_FDP0UA U2680 ( .D(SFIFOLock), .QTFCLK( ), .Q(SFIFOLock));
Q_FDP0UA U2681 ( .D(GFLBfull), .QTFCLK( ), .Q(GFLBfullD));
Q_FDP0UA U2682 ( .D(GFGBfullBw), .QTFCLK( ), .Q(GFGBfullBwD));
Q_FDP0UA U2683 ( .D(gfifoOff), .QTFCLK( ), .Q(gfifoOff));
Q_FDP0UA U2684 ( .D(gfifoAsyncOff), .QTFCLK( ), .Q(gfifoAsyncOff));
Q_FDP0UA U2685 ( .D(dbiEvent), .QTFCLK( ), .Q(dbiEventD));
Q_FDP0UA U2686 ( .D(APPLY_PI), .QTFCLK( ), .Q(applyPiR));
Q_FDP0UA U2687 ( .D(FvUseOnly), .QTFCLK( ), .Q(FvUseOnlyR));
Q_FDP0UA U2688 ( .D(callEmuPIi), .QTFCLK( ), .Q(sendPO));
Q_FDP0UA U2689 ( .D(callEmuPre), .QTFCLK( ), .Q(callEmuPreD));
Q_FDP0UA U2690 ( .D(sfifoSyncMode), .QTFCLK( ), .Q(sfifoSyncMode));
Q_FDP0UA U2691 ( .D(syncOtbChannels), .QTFCLK( ), .Q(syncOtbChannels));
Q_FDP0UA U2692 ( .D(fclkPerEval[7]), .QTFCLK( ), .Q(fclkPerEval[7]));
Q_FDP0UA U2693 ( .D(fclkPerEval[6]), .QTFCLK( ), .Q(fclkPerEval[6]));
Q_FDP0UA U2694 ( .D(fclkPerEval[5]), .QTFCLK( ), .Q(fclkPerEval[5]));
Q_FDP0UA U2695 ( .D(fclkPerEval[4]), .QTFCLK( ), .Q(fclkPerEval[4]));
Q_FDP0UA U2696 ( .D(fclkPerEval[3]), .QTFCLK( ), .Q(fclkPerEval[3]));
Q_FDP0UA U2697 ( .D(fclkPerEval[2]), .QTFCLK( ), .Q(fclkPerEval[2]));
Q_FDP0UA U2698 ( .D(fclkPerEval[1]), .QTFCLK( ), .Q(fclkPerEval[1]));
Q_FDP0UA U2699 ( .D(fclkPerEval[0]), .QTFCLK( ), .Q(fclkPerEval[0]));
Q_FDP0UA U2700 ( .D(sdlEnable), .QTFCLK( ), .Q(sdlEnable));
Q_FDP0UA U2701 ( .D(tbcEnable), .QTFCLK( ), .Q(tbcEnable));
Q_FDP0UA U2702 ( .D(evalOnDCtl[7]), .QTFCLK( ), .Q(evalOnDCtl[7]));
Q_FDP0UA U2703 ( .D(evalOnDCtl[6]), .QTFCLK( ), .Q(evalOnDCtl[6]));
Q_FDP0UA U2704 ( .D(evalOnDCtl[5]), .QTFCLK( ), .Q(evalOnDCtl[5]));
Q_FDP0UA U2705 ( .D(evalOnDCtl[4]), .QTFCLK( ), .Q(evalOnDCtl[4]));
Q_FDP0UA U2706 ( .D(evalOnDCtl[3]), .QTFCLK( ), .Q(evalOnDCtl[3]));
Q_FDP0UA U2707 ( .D(evalOnDCtl[2]), .QTFCLK( ), .Q(evalOnDCtl[2]));
Q_FDP0UA U2708 ( .D(evalOnDCtl[1]), .QTFCLK( ), .Q(evalOnDCtl[1]));
Q_FDP0UA U2709 ( .D(evalOnDCtl[0]), .QTFCLK( ), .Q(evalOnDCtl[0]));
Q_FDP0UA U2710 ( .D(hwClkDbg), .QTFCLK( ), .Q(hwClkDbg));
Q_FDP0UA U2711 ( .D(hwClkDbgTime), .QTFCLK( ), .Q(hwClkDbgTime));
Q_FDP0UA U2712 ( .D(sdlHaltHwClk), .QTFCLK( ), .Q(sdlHaltHwClk));
Q_FDP0UA U2713 ( .D(forceAbort), .QTFCLK( ), .Q(forceAbort));
Q_FDP0UA U2714 ( .D(maxBpCycle[15]), .QTFCLK( ), .Q(maxBpCycle[15]));
Q_FDP0UA U2715 ( .D(maxBpCycle[14]), .QTFCLK( ), .Q(maxBpCycle[14]));
Q_FDP0UA U2716 ( .D(maxBpCycle[13]), .QTFCLK( ), .Q(maxBpCycle[13]));
Q_FDP0UA U2717 ( .D(maxBpCycle[12]), .QTFCLK( ), .Q(maxBpCycle[12]));
Q_FDP0UA U2718 ( .D(maxBpCycle[11]), .QTFCLK( ), .Q(maxBpCycle[11]));
Q_FDP0UA U2719 ( .D(maxBpCycle[10]), .QTFCLK( ), .Q(maxBpCycle[10]));
Q_FDP0UA U2720 ( .D(maxBpCycle[9]), .QTFCLK( ), .Q(maxBpCycle[9]));
Q_FDP0UA U2721 ( .D(maxBpCycle[8]), .QTFCLK( ), .Q(maxBpCycle[8]));
Q_FDP0UA U2722 ( .D(maxBpCycle[7]), .QTFCLK( ), .Q(maxBpCycle[7]));
Q_FDP0UA U2723 ( .D(maxBpCycle[6]), .QTFCLK( ), .Q(maxBpCycle[6]));
Q_FDP0UA U2724 ( .D(maxBpCycle[5]), .QTFCLK( ), .Q(maxBpCycle[5]));
Q_FDP0UA U2725 ( .D(maxBpCycle[4]), .QTFCLK( ), .Q(maxBpCycle[4]));
Q_FDP0UA U2726 ( .D(maxBpCycle[3]), .QTFCLK( ), .Q(maxBpCycle[3]));
Q_FDP0UA U2727 ( .D(maxBpCycle[2]), .QTFCLK( ), .Q(maxBpCycle[2]));
Q_FDP0UA U2728 ( .D(maxBpCycle[1]), .QTFCLK( ), .Q(maxBpCycle[1]));
Q_FDP0UA U2729 ( .D(maxBpCycle[0]), .QTFCLK( ), .Q(maxBpCycle[0]));
Q_FDP0UA U2730 ( .D(maxAcCycle[15]), .QTFCLK( ), .Q(maxAcCycle[15]));
Q_FDP0UA U2731 ( .D(maxAcCycle[14]), .QTFCLK( ), .Q(maxAcCycle[14]));
Q_FDP0UA U2732 ( .D(maxAcCycle[13]), .QTFCLK( ), .Q(maxAcCycle[13]));
Q_FDP0UA U2733 ( .D(maxAcCycle[12]), .QTFCLK( ), .Q(maxAcCycle[12]));
Q_FDP0UA U2734 ( .D(maxAcCycle[11]), .QTFCLK( ), .Q(maxAcCycle[11]));
Q_FDP0UA U2735 ( .D(maxAcCycle[10]), .QTFCLK( ), .Q(maxAcCycle[10]));
Q_FDP0UA U2736 ( .D(maxAcCycle[9]), .QTFCLK( ), .Q(maxAcCycle[9]));
Q_FDP0UA U2737 ( .D(maxAcCycle[8]), .QTFCLK( ), .Q(maxAcCycle[8]));
Q_FDP0UA U2738 ( .D(maxAcCycle[7]), .QTFCLK( ), .Q(maxAcCycle[7]));
Q_FDP0UA U2739 ( .D(maxAcCycle[6]), .QTFCLK( ), .Q(maxAcCycle[6]));
Q_FDP0UA U2740 ( .D(maxAcCycle[5]), .QTFCLK( ), .Q(maxAcCycle[5]));
Q_FDP0UA U2741 ( .D(maxAcCycle[4]), .QTFCLK( ), .Q(maxAcCycle[4]));
Q_FDP0UA U2742 ( .D(maxAcCycle[3]), .QTFCLK( ), .Q(maxAcCycle[3]));
Q_FDP0UA U2743 ( .D(maxAcCycle[2]), .QTFCLK( ), .Q(maxAcCycle[2]));
Q_FDP0UA U2744 ( .D(maxAcCycle[1]), .QTFCLK( ), .Q(maxAcCycle[1]));
Q_FDP0UA U2745 ( .D(maxAcCycle[0]), .QTFCLK( ), .Q(maxAcCycle[0]));
Q_FDP0UA U2746 ( .D(hssReset), .QTFCLK( ), .Q(hssReset));
Q_FDP0UA U2747 ( .D(FvSimple2), .QTFCLK( ), .Q(FvSimple2));
Q_FDP0UA U2748 ( .D(DccFrameCycle[7]), .QTFCLK( ), .Q(DccFrameCycle[7]));
Q_FDP0UA U2749 ( .D(DccFrameCycle[6]), .QTFCLK( ), .Q(DccFrameCycle[6]));
Q_FDP0UA U2750 ( .D(DccFrameCycle[5]), .QTFCLK( ), .Q(DccFrameCycle[5]));
Q_FDP0UA U2751 ( .D(DccFrameCycle[4]), .QTFCLK( ), .Q(DccFrameCycle[4]));
Q_FDP0UA U2752 ( .D(DccFrameCycle[3]), .QTFCLK( ), .Q(DccFrameCycle[3]));
Q_FDP0UA U2753 ( .D(DccFrameCycle[2]), .QTFCLK( ), .Q(DccFrameCycle[2]));
Q_FDP0UA U2754 ( .D(DccFrameCycle[1]), .QTFCLK( ), .Q(DccFrameCycle[1]));
Q_FDP0UA U2755 ( .D(DccFrameCycle[0]), .QTFCLK( ), .Q(DccFrameCycle[0]));
Q_FDP0UA U2756 ( .D(DccFrameMark[7]), .QTFCLK( ), .Q(DccFrameMark[7]));
Q_FDP0UA U2757 ( .D(DccFrameMark[6]), .QTFCLK( ), .Q(DccFrameMark[6]));
Q_FDP0UA U2758 ( .D(DccFrameMark[5]), .QTFCLK( ), .Q(DccFrameMark[5]));
Q_FDP0UA U2759 ( .D(DccFrameMark[4]), .QTFCLK( ), .Q(DccFrameMark[4]));
Q_FDP0UA U2760 ( .D(DccFrameMark[3]), .QTFCLK( ), .Q(DccFrameMark[3]));
Q_FDP0UA U2761 ( .D(DccFrameMark[2]), .QTFCLK( ), .Q(DccFrameMark[2]));
Q_FDP0UA U2762 ( .D(DccFrameMark[1]), .QTFCLK( ), .Q(DccFrameMark[1]));
Q_FDP0UA U2763 ( .D(DccFrameMark[0]), .QTFCLK( ), .Q(DccFrameMark[0]));
Q_FDP0UA U2764 ( .D(xcReplayOn), .QTFCLK( ), .Q(xcReplayOn));
Q_FDP0UA U2765 ( .D(xcRecordOn), .QTFCLK( ), .Q(xcRecordOn));
Q_FDP0UA U2766 ( .D(xc_mioOn), .QTFCLK( ), .Q(xc_mioOn));
Q_FDP0UA U2767 ( .D(gfPushDly[7]), .QTFCLK( ), .Q(gfPushDly[7]));
Q_FDP0UA U2768 ( .D(gfPushDly[6]), .QTFCLK( ), .Q(gfPushDly[6]));
Q_FDP0UA U2769 ( .D(gfPushDly[5]), .QTFCLK( ), .Q(gfPushDly[5]));
Q_FDP0UA U2770 ( .D(gfPushDly[4]), .QTFCLK( ), .Q(gfPushDly[4]));
Q_FDP0UA U2771 ( .D(gfPushDly[3]), .QTFCLK( ), .Q(gfPushDly[3]));
Q_FDP0UA U2772 ( .D(gfPushDly[2]), .QTFCLK( ), .Q(gfPushDly[2]));
Q_FDP0UA U2773 ( .D(gfPushDly[1]), .QTFCLK( ), .Q(gfPushDly[1]));
Q_FDP0UA U2774 ( .D(gfPushDly[0]), .QTFCLK( ), .Q(gfPushDly[0]));
Q_FDP0UA U2775 ( .D(gfPushFill[3]), .QTFCLK( ), .Q(gfPushFill[3]));
Q_FDP0UA U2776 ( .D(gfPushFill[2]), .QTFCLK( ), .Q(gfPushFill[2]));
Q_FDP0UA U2777 ( .D(gfPushFill[1]), .QTFCLK( ), .Q(gfPushFill[1]));
Q_FDP0UA U2778 ( .D(gfPushFill[0]), .QTFCLK( ), .Q(gfPushFill[0]));
Q_AN02 U2779 ( .A0(holdEcm), .A1(active), .Z(holdEcmC));
Q_NR02 U2780 ( .A0(mpSt[2]), .A1(mpSt[0]), .Z(n2264));
Q_MX02 U2781 ( .S(n2172), .A0(n2265), .A1(n2266), .Z(simTimeEnable));
Q_AN02 U2782 ( .A0(n2264), .A1(n2192), .Z(n2265));
Q_MX02 U2783 ( .S(n2264), .A0(n2189), .A1(n2267), .Z(n2266));
Q_AN03 U2784 ( .A0(callEmu), .A1(n2121), .A2(n2189), .Z(n2267));
Q_INV U2785 ( .A(stopSDL), .Z(n2268));
Q_ND02 U2786 ( .A0(n3285), .A1(n2268), .Z(n2269));
Q_INV U2787 ( .A(cpfStop), .Z(n2270));
Q_LSN01 U2788 ( .S(n2270), .R(n3285), .Q(stopCPFPO), .QN( ));
Q_OR03 U2789 ( .A0(mioPOW_2[7]), .A1(stopEmuPO), .A2(n2271), .Z(stop3));
Q_OR03 U2790 ( .A0(bpHalt), .A1(mioPOW_2[6]), .A2(mioPOW_2[8]), .Z(n2271));
Q_LDP0 stopSDLPO_REG  ( .G(n2269), .D(stopSDL), .Q(stopSDLPO), .QN( ));
Q_MX02 U2792 ( .S(oneStepPIi), .A0(ixc_time.stopEcm), .A1(mpOn), .Z(stopT));
Q_AO21 U2793 ( .A0(lastDelta), .A1(evalOnC), .B0(hotSwapOnPI), .Z(mpSampleOv));
Q_AN02 U2794 ( .A0(dbiEvent), .A1(n2616), .Z(FvUseOnly));
Q_OR03 U2795 ( .A0(evalOnInt), .A1(n2272), .A2(n2216), .Z(evalOn));
Q_AN02 U2796 ( .A0(evalOnIntD), .A1(n2288), .Z(n2272));
Q_AN03 U2797 ( .A0(sdlEnable), .A1(sdlStop), .A2(xcReplayOn), .Z(sdlStopRply));
Q_AN03 U2798 ( .A0(sdlEnable), .A1(sdlStop), .A2(n2273), .Z(stopSDL));
Q_INV U2799 ( .A(xcReplayOn), .Z(n2273));
Q_AN02 U2800 ( .A0(stop4), .A1(tbcEnable), .Z(stop4R));
Q_AN02 U2801 ( .A0(stop2), .A1(tbcEnable), .Z(stop2R));
Q_AN02 U2802 ( .A0(stop1), .A1(tbcEnable), .Z(stop1R));
Q_AN02 U2803 ( .A0(n2275), .A1(n2274), .Z(evalOnInt));
Q_OR03 U2804 ( .A0(FTcallW), .A1(evalOnSync), .A2(lockTraceOn), .Z(n2274));
Q_INV U2805 ( .A(sdlStopRplyD), .Z(n2276));
Q_OA21 U2806 ( .A0(evalOnOrig), .A1(GFbusyW), .B0(n2276), .Z(evalOnSync));
Q_OR03 U2807 ( .A0(hwClkDbgOn), .A1(eventOnR), .A2(callEmuPre), .Z(n2277));
Q_AO21 U2808 ( .A0(tbcPOd), .A1(n2278), .B0(n2277), .Z(evalOnOrig));
Q_INV U2809 ( .A(mioPOW_2[1]), .Z(n2278));
Q_AN02 U2810 ( .A0(n2279), .A1(n2288), .Z(GFbusyW));
Q_OR03 U2811 ( .A0(dbiEvent), .A1(n2281), .A2(n2280), .Z(n2279));
Q_OR03 U2812 ( .A0(isfWait), .A1(gfifoWait), .A2(ptxBusy), .Z(n2280));
Q_OR03 U2813 ( .A0(callEmuWait), .A1(callEmuEv), .A2(osfWait), .Z(n2281));
Q_AN03 U2814 ( .A0(n2282), .A1(APPLY_PI), .A2(n2211), .Z(dbiEvent));
Q_INV U2815 ( .A(applyPiR), .Z(n2282));
Q_OR03 U2816 ( .A0(svAsyncCall), .A1(n2283), .A2(n2284), .Z(FTcallW));
Q_OR03 U2817 ( .A0(ecmHoldBusy), .A1(GFAck), .A2(otbAsyncCall), .Z(n2283));
Q_OR02 U2818 ( .A0(n2286), .A1(n2285), .Z(n2284));
Q_OR03 U2819 ( .A0(gfifoAckWait[1]), .A1(gfifoAckWait[0]), .A2(n2287), .Z(n2285));
Q_OR03 U2820 ( .A0(gfifoAckWait[4]), .A1(gfifoAckWait[3]), .A2(gfifoAckWait[2]), .Z(n2286));
Q_OR03 U2821 ( .A0(gfifoAckWait[7]), .A1(gfifoAckWait[6]), .A2(gfifoAckWait[5]), .Z(n2287));
Q_INV U2822 ( .A(FvSimple2), .Z(n2288));
Q_FDP0 callEmuWait_REG  ( .CK(uClk), .D(callEmuWaitN), .Q(callEmuWait), .QN( ));
Q_AO21 U2824 ( .A0(asyncCall), .A1(sfifoSyncMode), .B0(n2289), .Z(n2290));
Q_OR03 U2825 ( .A0(holdEcm), .A1(ptxBusy), .A2(isfWait), .Z(n2289));
Q_FDP0 callEmuWaitC_REG  ( .CK(uClk), .D(n2290), .Q(callEmuWaitC), .QN( ));
Q_AD01HF U2827 ( .A0(uClkCntr[1]), .B0(uClkCntr[0]), .S(n2291), .CO(n2292));
Q_AD01HF U2828 ( .A0(uClkCntr[2]), .B0(n2292), .S(n2293), .CO(n2294));
Q_AD01HF U2829 ( .A0(uClkCntr[3]), .B0(n2294), .S(n2295), .CO(n2296));
Q_AD01HF U2830 ( .A0(uClkCntr[4]), .B0(n2296), .S(n2297), .CO(n2298));
Q_AD01HF U2831 ( .A0(uClkCntr[5]), .B0(n2298), .S(n2299), .CO(n2300));
Q_AD01HF U2832 ( .A0(uClkCntr[6]), .B0(n2300), .S(n2301), .CO(n2302));
Q_AD01HF U2833 ( .A0(uClkCntr[7]), .B0(n2302), .S(n2303), .CO(n2304));
Q_AD01HF U2834 ( .A0(uClkCntr[8]), .B0(n2304), .S(n2305), .CO(n2306));
Q_AD01HF U2835 ( .A0(uClkCntr[9]), .B0(n2306), .S(n2307), .CO(n2308));
Q_AD01HF U2836 ( .A0(uClkCntr[10]), .B0(n2308), .S(n2309), .CO(n2310));
Q_AD01HF U2837 ( .A0(uClkCntr[11]), .B0(n2310), .S(n2311), .CO(n2312));
Q_AD01HF U2838 ( .A0(uClkCntr[12]), .B0(n2312), .S(n2313), .CO(n2314));
Q_AD01HF U2839 ( .A0(uClkCntr[13]), .B0(n2314), .S(n2315), .CO(n2316));
Q_AD01HF U2840 ( .A0(uClkCntr[14]), .B0(n2316), .S(n2317), .CO(n2318));
Q_AD01HF U2841 ( .A0(uClkCntr[15]), .B0(n2318), .S(n2319), .CO(n2320));
Q_AD01HF U2842 ( .A0(uClkCntr[16]), .B0(n2320), .S(n2321), .CO(n2322));
Q_AD01HF U2843 ( .A0(uClkCntr[17]), .B0(n2322), .S(n2323), .CO(n2324));
Q_AD01HF U2844 ( .A0(uClkCntr[18]), .B0(n2324), .S(n2325), .CO(n2326));
Q_AD01HF U2845 ( .A0(uClkCntr[19]), .B0(n2326), .S(n2327), .CO(n2328));
Q_AD01HF U2846 ( .A0(uClkCntr[20]), .B0(n2328), .S(n2329), .CO(n2330));
Q_AD01HF U2847 ( .A0(uClkCntr[21]), .B0(n2330), .S(n2331), .CO(n2332));
Q_AD01HF U2848 ( .A0(uClkCntr[22]), .B0(n2332), .S(n2333), .CO(n2334));
Q_AD01HF U2849 ( .A0(uClkCntr[23]), .B0(n2334), .S(n2335), .CO(n2336));
Q_AD01HF U2850 ( .A0(uClkCntr[24]), .B0(n2336), .S(n2337), .CO(n2338));
Q_AD01HF U2851 ( .A0(uClkCntr[25]), .B0(n2338), .S(n2339), .CO(n2340));
Q_AD01HF U2852 ( .A0(uClkCntr[26]), .B0(n2340), .S(n2341), .CO(n2342));
Q_AD01HF U2853 ( .A0(uClkCntr[27]), .B0(n2342), .S(n2343), .CO(n2344));
Q_AD01HF U2854 ( .A0(uClkCntr[28]), .B0(n2344), .S(n2345), .CO(n2346));
Q_AD01HF U2855 ( .A0(uClkCntr[29]), .B0(n2346), .S(n2347), .CO(n2348));
Q_AD01HF U2856 ( .A0(uClkCntr[30]), .B0(n2348), .S(n2349), .CO(n2350));
Q_AD01HF U2857 ( .A0(uClkCntr[31]), .B0(n2350), .S(n2351), .CO(n2352));
Q_AD01HF U2858 ( .A0(uClkCntr[32]), .B0(n2352), .S(n2353), .CO(n2354));
Q_AD01HF U2859 ( .A0(uClkCntr[33]), .B0(n2354), .S(n2355), .CO(n2356));
Q_AD01HF U2860 ( .A0(uClkCntr[34]), .B0(n2356), .S(n2357), .CO(n2358));
Q_AD01HF U2861 ( .A0(uClkCntr[35]), .B0(n2358), .S(n2359), .CO(n2360));
Q_AD01HF U2862 ( .A0(uClkCntr[36]), .B0(n2360), .S(n2361), .CO(n2362));
Q_AD01HF U2863 ( .A0(uClkCntr[37]), .B0(n2362), .S(n2363), .CO(n2364));
Q_AD01HF U2864 ( .A0(uClkCntr[38]), .B0(n2364), .S(n2365), .CO(n2366));
Q_AD01HF U2865 ( .A0(uClkCntr[39]), .B0(n2366), .S(n2367), .CO(n2368));
Q_AD01HF U2866 ( .A0(uClkCntr[40]), .B0(n2368), .S(n2369), .CO(n2370));
Q_AD01HF U2867 ( .A0(uClkCntr[41]), .B0(n2370), .S(n2371), .CO(n2372));
Q_AD01HF U2868 ( .A0(uClkCntr[42]), .B0(n2372), .S(n2373), .CO(n2374));
Q_AD01HF U2869 ( .A0(uClkCntr[43]), .B0(n2374), .S(n2375), .CO(n2376));
Q_AD01HF U2870 ( .A0(uClkCntr[44]), .B0(n2376), .S(n2377), .CO(n2378));
Q_AD01HF U2871 ( .A0(uClkCntr[45]), .B0(n2378), .S(n2379), .CO(n2380));
Q_AD01HF U2872 ( .A0(uClkCntr[46]), .B0(n2380), .S(n2381), .CO(n2382));
Q_AD01HF U2873 ( .A0(uClkCntr[47]), .B0(n2382), .S(n2383), .CO(n2384));
Q_AD01HF U2874 ( .A0(uClkCntr[48]), .B0(n2384), .S(n2385), .CO(n2386));
Q_AD01HF U2875 ( .A0(uClkCntr[49]), .B0(n2386), .S(n2387), .CO(n2388));
Q_AD01HF U2876 ( .A0(uClkCntr[50]), .B0(n2388), .S(n2389), .CO(n2390));
Q_AD01HF U2877 ( .A0(uClkCntr[51]), .B0(n2390), .S(n2391), .CO(n2392));
Q_AD01HF U2878 ( .A0(uClkCntr[52]), .B0(n2392), .S(n2393), .CO(n2394));
Q_AD01HF U2879 ( .A0(uClkCntr[53]), .B0(n2394), .S(n2395), .CO(n2396));
Q_AD01HF U2880 ( .A0(uClkCntr[54]), .B0(n2396), .S(n2397), .CO(n2398));
Q_AD01HF U2881 ( .A0(uClkCntr[55]), .B0(n2398), .S(n2399), .CO(n2400));
Q_AD01HF U2882 ( .A0(uClkCntr[56]), .B0(n2400), .S(n2401), .CO(n2402));
Q_AD01HF U2883 ( .A0(uClkCntr[57]), .B0(n2402), .S(n2403), .CO(n2404));
Q_AD01HF U2884 ( .A0(uClkCntr[58]), .B0(n2404), .S(n2405), .CO(n2406));
Q_AD01HF U2885 ( .A0(uClkCntr[59]), .B0(n2406), .S(n2407), .CO(n2408));
Q_AD01HF U2886 ( .A0(uClkCntr[60]), .B0(n2408), .S(n2409), .CO(n2410));
Q_AD01HF U2887 ( .A0(uClkCntr[61]), .B0(n2410), .S(n2411), .CO(n2412));
Q_AD01HF U2888 ( .A0(uClkCntr[62]), .B0(n2412), .S(n2413), .CO(n2414));
Q_FDP0 \nextDutTimeP_REG[63] ( .CK(mcp), .D(ixc_time.nextDutTime[63]), .Q(nextDutTimeP[63]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[62] ( .CK(mcp), .D(ixc_time.nextDutTime[62]), .Q(nextDutTimeP[62]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[61] ( .CK(mcp), .D(ixc_time.nextDutTime[61]), .Q(nextDutTimeP[61]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[60] ( .CK(mcp), .D(ixc_time.nextDutTime[60]), .Q(nextDutTimeP[60]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[59] ( .CK(mcp), .D(ixc_time.nextDutTime[59]), .Q(nextDutTimeP[59]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[58] ( .CK(mcp), .D(ixc_time.nextDutTime[58]), .Q(nextDutTimeP[58]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[57] ( .CK(mcp), .D(ixc_time.nextDutTime[57]), .Q(nextDutTimeP[57]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[56] ( .CK(mcp), .D(ixc_time.nextDutTime[56]), .Q(nextDutTimeP[56]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[55] ( .CK(mcp), .D(ixc_time.nextDutTime[55]), .Q(nextDutTimeP[55]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[54] ( .CK(mcp), .D(ixc_time.nextDutTime[54]), .Q(nextDutTimeP[54]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[53] ( .CK(mcp), .D(ixc_time.nextDutTime[53]), .Q(nextDutTimeP[53]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[52] ( .CK(mcp), .D(ixc_time.nextDutTime[52]), .Q(nextDutTimeP[52]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[51] ( .CK(mcp), .D(ixc_time.nextDutTime[51]), .Q(nextDutTimeP[51]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[50] ( .CK(mcp), .D(ixc_time.nextDutTime[50]), .Q(nextDutTimeP[50]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[49] ( .CK(mcp), .D(ixc_time.nextDutTime[49]), .Q(nextDutTimeP[49]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[48] ( .CK(mcp), .D(ixc_time.nextDutTime[48]), .Q(nextDutTimeP[48]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[47] ( .CK(mcp), .D(ixc_time.nextDutTime[47]), .Q(nextDutTimeP[47]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[46] ( .CK(mcp), .D(ixc_time.nextDutTime[46]), .Q(nextDutTimeP[46]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[45] ( .CK(mcp), .D(ixc_time.nextDutTime[45]), .Q(nextDutTimeP[45]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[44] ( .CK(mcp), .D(ixc_time.nextDutTime[44]), .Q(nextDutTimeP[44]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[43] ( .CK(mcp), .D(ixc_time.nextDutTime[43]), .Q(nextDutTimeP[43]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[42] ( .CK(mcp), .D(ixc_time.nextDutTime[42]), .Q(nextDutTimeP[42]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[41] ( .CK(mcp), .D(ixc_time.nextDutTime[41]), .Q(nextDutTimeP[41]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[40] ( .CK(mcp), .D(ixc_time.nextDutTime[40]), .Q(nextDutTimeP[40]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[39] ( .CK(mcp), .D(ixc_time.nextDutTime[39]), .Q(nextDutTimeP[39]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[38] ( .CK(mcp), .D(ixc_time.nextDutTime[38]), .Q(nextDutTimeP[38]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[37] ( .CK(mcp), .D(ixc_time.nextDutTime[37]), .Q(nextDutTimeP[37]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[36] ( .CK(mcp), .D(ixc_time.nextDutTime[36]), .Q(nextDutTimeP[36]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[35] ( .CK(mcp), .D(ixc_time.nextDutTime[35]), .Q(nextDutTimeP[35]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[34] ( .CK(mcp), .D(ixc_time.nextDutTime[34]), .Q(nextDutTimeP[34]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[33] ( .CK(mcp), .D(ixc_time.nextDutTime[33]), .Q(nextDutTimeP[33]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[32] ( .CK(mcp), .D(ixc_time.nextDutTime[32]), .Q(nextDutTimeP[32]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[31] ( .CK(mcp), .D(ixc_time.nextDutTime[31]), .Q(nextDutTimeP[31]), .QN( ));
Q_FDP0 \nextDutTimeP_REG[30] ( .CK(mcp), .D(ixc_time.nextDutTime[30]), .Q(nextDutTimeP[30]), .QN(n3685));
Q_FDP0 \nextDutTimeP_REG[29] ( .CK(mcp), .D(ixc_time.nextDutTime[29]), .Q(nextDutTimeP[29]), .QN(n3686));
Q_FDP0 \nextDutTimeP_REG[28] ( .CK(mcp), .D(ixc_time.nextDutTime[28]), .Q(nextDutTimeP[28]), .QN(n3687));
Q_FDP0 \nextDutTimeP_REG[27] ( .CK(mcp), .D(ixc_time.nextDutTime[27]), .Q(nextDutTimeP[27]), .QN(n3688));
Q_FDP0 \nextDutTimeP_REG[26] ( .CK(mcp), .D(ixc_time.nextDutTime[26]), .Q(nextDutTimeP[26]), .QN(n3689));
Q_FDP0 \nextDutTimeP_REG[25] ( .CK(mcp), .D(ixc_time.nextDutTime[25]), .Q(nextDutTimeP[25]), .QN(n3690));
Q_FDP0 \nextDutTimeP_REG[24] ( .CK(mcp), .D(ixc_time.nextDutTime[24]), .Q(nextDutTimeP[24]), .QN(n3691));
Q_FDP0 \nextDutTimeP_REG[23] ( .CK(mcp), .D(ixc_time.nextDutTime[23]), .Q(nextDutTimeP[23]), .QN(n3692));
Q_FDP0 \nextDutTimeP_REG[22] ( .CK(mcp), .D(ixc_time.nextDutTime[22]), .Q(nextDutTimeP[22]), .QN(n3693));
Q_FDP0 \nextDutTimeP_REG[21] ( .CK(mcp), .D(ixc_time.nextDutTime[21]), .Q(nextDutTimeP[21]), .QN(n3694));
Q_FDP0 \nextDutTimeP_REG[20] ( .CK(mcp), .D(ixc_time.nextDutTime[20]), .Q(nextDutTimeP[20]), .QN(n3695));
Q_FDP0 \nextDutTimeP_REG[19] ( .CK(mcp), .D(ixc_time.nextDutTime[19]), .Q(nextDutTimeP[19]), .QN(n3696));
Q_FDP0 \nextDutTimeP_REG[18] ( .CK(mcp), .D(ixc_time.nextDutTime[18]), .Q(nextDutTimeP[18]), .QN(n3697));
Q_FDP0 \nextDutTimeP_REG[17] ( .CK(mcp), .D(ixc_time.nextDutTime[17]), .Q(nextDutTimeP[17]), .QN(n3698));
Q_FDP0 \nextDutTimeP_REG[16] ( .CK(mcp), .D(ixc_time.nextDutTime[16]), .Q(nextDutTimeP[16]), .QN(n3699));
Q_FDP0 \nextDutTimeP_REG[15] ( .CK(mcp), .D(ixc_time.nextDutTime[15]), .Q(nextDutTimeP[15]), .QN(n3700));
Q_FDP0 \nextDutTimeP_REG[14] ( .CK(mcp), .D(ixc_time.nextDutTime[14]), .Q(nextDutTimeP[14]), .QN(n3701));
Q_FDP0 \nextDutTimeP_REG[13] ( .CK(mcp), .D(ixc_time.nextDutTime[13]), .Q(nextDutTimeP[13]), .QN(n3702));
Q_FDP0 \nextDutTimeP_REG[12] ( .CK(mcp), .D(ixc_time.nextDutTime[12]), .Q(nextDutTimeP[12]), .QN(n3703));
Q_FDP0 \nextDutTimeP_REG[11] ( .CK(mcp), .D(ixc_time.nextDutTime[11]), .Q(nextDutTimeP[11]), .QN(n3704));
Q_FDP0 \nextDutTimeP_REG[10] ( .CK(mcp), .D(ixc_time.nextDutTime[10]), .Q(nextDutTimeP[10]), .QN(n3705));
Q_FDP0 \nextDutTimeP_REG[9] ( .CK(mcp), .D(ixc_time.nextDutTime[9]), .Q(nextDutTimeP[9]), .QN(n3706));
Q_FDP0 \nextDutTimeP_REG[8] ( .CK(mcp), .D(ixc_time.nextDutTime[8]), .Q(nextDutTimeP[8]), .QN(n3707));
Q_FDP0 \nextDutTimeP_REG[7] ( .CK(mcp), .D(ixc_time.nextDutTime[7]), .Q(nextDutTimeP[7]), .QN(n3708));
Q_FDP0 \nextDutTimeP_REG[6] ( .CK(mcp), .D(ixc_time.nextDutTime[6]), .Q(nextDutTimeP[6]), .QN(n3709));
Q_FDP0 \nextDutTimeP_REG[5] ( .CK(mcp), .D(ixc_time.nextDutTime[5]), .Q(nextDutTimeP[5]), .QN(n3710));
Q_FDP0 \nextDutTimeP_REG[4] ( .CK(mcp), .D(ixc_time.nextDutTime[4]), .Q(nextDutTimeP[4]), .QN(n3711));
Q_FDP0 \nextDutTimeP_REG[3] ( .CK(mcp), .D(ixc_time.nextDutTime[3]), .Q(nextDutTimeP[3]), .QN(n3712));
Q_FDP0 \nextDutTimeP_REG[2] ( .CK(mcp), .D(ixc_time.nextDutTime[2]), .Q(nextDutTimeP[2]), .QN(n3713));
Q_FDP0 \nextDutTimeP_REG[1] ( .CK(mcp), .D(ixc_time.nextDutTime[1]), .Q(nextDutTimeP[1]), .QN(n3714));
Q_FDP0 \nextDutTimeP_REG[0] ( .CK(mcp), .D(ixc_time.nextDutTime[0]), .Q(nextDutTimeP[0]), .QN(n3715));
Q_AO21 U2953 ( .A0(n2464), .A1(n1525), .B0(lbrOn), .Z(n2419));
Q_AO21 U2954 ( .A0(n2419), .A1(dccState), .B0(n2420), .Z(n2421));
Q_INV U2955 ( .A(n2424), .Z(n2420));
Q_INV U2956 ( .A(n2416), .Z(n2422));
Q_OR02 U2957 ( .A0(n2422), .A1(n2421), .Z(n2423));
Q_OR02 U2958 ( .A0(dccState), .A1(lbrOn), .Z(n2424));
Q_AN02 U2959 ( .A0(n2416), .A1(n2424), .Z(n2417));
Q_INV U2960 ( .A(n2415), .Z(n2418));
Q_AN02 U2961 ( .A0(dccState), .A1(n2468), .Z(n2425));
Q_AN02 U2962 ( .A0(dccState), .A1(n2469), .Z(n2426));
Q_AN02 U2963 ( .A0(dccState), .A1(n2470), .Z(n2427));
Q_AN02 U2964 ( .A0(dccState), .A1(n2471), .Z(n2428));
Q_AN02 U2965 ( .A0(dccState), .A1(n2472), .Z(n2429));
Q_AN02 U2966 ( .A0(dccState), .A1(n2473), .Z(n2430));
Q_AN02 U2967 ( .A0(dccState), .A1(n2474), .Z(n2431));
Q_OR02 U2968 ( .A0(n2433), .A1(n2475), .Z(n2432));
Q_AN03 U2969 ( .A0(n1525), .A1(n2435), .A2(dccState), .Z(n2434));
Q_AO21 U2970 ( .A0(n2450), .A1(n2436), .B0(n2451), .Z(n2435));
Q_OR03 U2971 ( .A0(n2448), .A1(n2437), .A2(n2438), .Z(n2436));
Q_AO21 U2972 ( .A0(n2440), .A1(n2444), .B0(n2439), .Z(n2438));
Q_AN03 U2973 ( .A0(n2440), .A1(n2443), .A2(n2441), .Z(n2439));
Q_AN02 U2974 ( .A0(n2475), .A1(n2442), .Z(n2441));
Q_INV U2975 ( .A(DccFrameMark[0]), .Z(n2442));
Q_OR02 U2976 ( .A0(n2474), .A1(n2445), .Z(n2443));
Q_AN02 U2977 ( .A0(n2474), .A1(n2445), .Z(n2444));
Q_INV U2978 ( .A(DccFrameMark[1]), .Z(n2445));
Q_OA21 U2979 ( .A0(n2473), .A1(n2446), .B0(n2447), .Z(n2440));
Q_AN03 U2980 ( .A0(n2473), .A1(n2446), .A2(n2447), .Z(n2437));
Q_INV U2981 ( .A(DccFrameMark[2]), .Z(n2446));
Q_OR02 U2982 ( .A0(n2472), .A1(n2449), .Z(n2447));
Q_AN02 U2983 ( .A0(n2472), .A1(n2449), .Z(n2448));
Q_INV U2984 ( .A(DccFrameMark[3]), .Z(n2449));
Q_OR03 U2985 ( .A0(n2462), .A1(n2452), .A2(n2453), .Z(n2451));
Q_AO21 U2986 ( .A0(n2456), .A1(n2458), .B0(n2454), .Z(n2453));
Q_OA21 U2987 ( .A0(n2471), .A1(n2457), .B0(n2455), .Z(n2450));
Q_AN03 U2988 ( .A0(n2471), .A1(n2457), .A2(n2455), .Z(n2454));
Q_INV U2989 ( .A(DccFrameMark[4]), .Z(n2457));
Q_OA21 U2990 ( .A0(n2470), .A1(n2459), .B0(n2456), .Z(n2455));
Q_AN02 U2991 ( .A0(n2470), .A1(n2459), .Z(n2458));
Q_INV U2992 ( .A(DccFrameMark[5]), .Z(n2459));
Q_OA21 U2993 ( .A0(n2469), .A1(n2460), .B0(n2461), .Z(n2456));
Q_AN03 U2994 ( .A0(n2469), .A1(n2460), .A2(n2461), .Z(n2452));
Q_INV U2995 ( .A(DccFrameMark[6]), .Z(n2460));
Q_OR02 U2996 ( .A0(n2468), .A1(n2463), .Z(n2461));
Q_AN02 U2997 ( .A0(n2468), .A1(n2463), .Z(n2462));
Q_INV U2998 ( .A(DccFrameMark[7]), .Z(n2463));
Q_OR02 U2999 ( .A0(n2466), .A1(n2465), .Z(n2464));
Q_OR03 U3000 ( .A0(n2469), .A1(n2468), .A2(n2467), .Z(n2465));
Q_OR03 U3001 ( .A0(n2472), .A1(n2471), .A2(n2470), .Z(n2466));
Q_OR03 U3002 ( .A0(n2475), .A1(n2474), .A2(n2473), .Z(n2467));
Q_AN02 U3003 ( .A0(n2418), .A1(n2487), .Z(n2468));
Q_AN02 U3004 ( .A0(n2418), .A1(n2489), .Z(n2469));
Q_AN02 U3005 ( .A0(n2418), .A1(n2491), .Z(n2470));
Q_AN02 U3006 ( .A0(n2418), .A1(n2493), .Z(n2471));
Q_AN02 U3007 ( .A0(n2418), .A1(n2495), .Z(n2472));
Q_AN02 U3008 ( .A0(n2418), .A1(n2497), .Z(n2473));
Q_AN02 U3009 ( .A0(n2418), .A1(n2499), .Z(n2474));
Q_NR02 U3010 ( .A0(n2415), .A1(dccFrameFill[0]), .Z(n2475));
Q_AN02 U3011 ( .A0(n2477), .A1(n2476), .Z(n2415));
Q_AN03 U3012 ( .A0(n2480), .A1(n2479), .A2(n2478), .Z(n2476));
Q_AN03 U3013 ( .A0(n2483), .A1(n2482), .A2(n2481), .Z(n2477));
Q_AN03 U3014 ( .A0(n2486), .A1(n2485), .A2(n2484), .Z(n2478));
Q_XNR2 U3015 ( .A0(n2487), .A1(DccFrameCycle[7]), .Z(n2479));
Q_XNR2 U3016 ( .A0(n2489), .A1(DccFrameCycle[6]), .Z(n2480));
Q_XNR2 U3017 ( .A0(n2491), .A1(DccFrameCycle[5]), .Z(n2481));
Q_XNR2 U3018 ( .A0(n2493), .A1(DccFrameCycle[4]), .Z(n2482));
Q_XNR2 U3019 ( .A0(n2495), .A1(DccFrameCycle[3]), .Z(n2483));
Q_XNR2 U3020 ( .A0(n2497), .A1(DccFrameCycle[2]), .Z(n2484));
Q_XNR2 U3021 ( .A0(n2499), .A1(DccFrameCycle[1]), .Z(n2485));
Q_XOR2 U3022 ( .A0(dccFrameFill[0]), .A1(DccFrameCycle[0]), .Z(n2486));
Q_XOR2 U3023 ( .A0(dccFrameFill[7]), .A1(n2488), .Z(n2487));
Q_AD01HF U3024 ( .A0(dccFrameFill[6]), .B0(n2490), .S(n2489), .CO(n2488));
Q_AD01HF U3025 ( .A0(dccFrameFill[5]), .B0(n2492), .S(n2491), .CO(n2490));
Q_AD01HF U3026 ( .A0(dccFrameFill[4]), .B0(n2494), .S(n2493), .CO(n2492));
Q_AD01HF U3027 ( .A0(dccFrameFill[3]), .B0(n2496), .S(n2495), .CO(n2494));
Q_AD01HF U3028 ( .A0(dccFrameFill[2]), .B0(n2498), .S(n2497), .CO(n2496));
Q_AD01HF U3029 ( .A0(dccFrameFill[1]), .B0(dccFrameFill[0]), .S(n2499), .CO(n2498));
Q_OR02 U3030 ( .A0(n2501), .A1(n2500), .Z(n2416));
Q_OR03 U3031 ( .A0(DccFrameCycle[1]), .A1(DccFrameCycle[0]), .A2(n2502), .Z(n2500));
Q_OR03 U3032 ( .A0(DccFrameCycle[4]), .A1(DccFrameCycle[3]), .A2(DccFrameCycle[2]), .Z(n2501));
Q_OR03 U3033 ( .A0(DccFrameCycle[7]), .A1(DccFrameCycle[6]), .A2(DccFrameCycle[5]), .Z(n2502));
Q_AN02 U3034 ( .A0(ptxHoldEcm), .A1(xcRecordOn), .Z(n2503));
Q_FDP0 holdEcmPtxOn_REG  ( .CK(uClk), .D(n2503), .Q(holdEcmPtxOn), .QN( ));
Q_BUFZP U3036 ( .OE(syncEn), .A(n2504), .Z(stop1));
Q_OR02 U3037 ( .A0(GFbusy), .A1(n402), .Z(n2507));
Q_MX02 U3038 ( .S(evalOnC), .A0(maxFck2Sync[15]), .A1(n2570), .Z(n2508));
Q_MX02 U3039 ( .S(evalOnC), .A0(maxFck2Sync[14]), .A1(n2572), .Z(n2509));
Q_MX02 U3040 ( .S(evalOnC), .A0(maxFck2Sync[13]), .A1(n2574), .Z(n2510));
Q_MX02 U3041 ( .S(evalOnC), .A0(maxFck2Sync[12]), .A1(n2576), .Z(n2511));
Q_MX02 U3042 ( .S(evalOnC), .A0(maxFck2Sync[11]), .A1(n2578), .Z(n2512));
Q_MX02 U3043 ( .S(evalOnC), .A0(maxFck2Sync[10]), .A1(n2580), .Z(n2513));
Q_MX02 U3044 ( .S(evalOnC), .A0(maxFck2Sync[9]), .A1(n2582), .Z(n2514));
Q_MX02 U3045 ( .S(evalOnC), .A0(maxFck2Sync[8]), .A1(n2584), .Z(n2515));
Q_MX02 U3046 ( .S(evalOnC), .A0(maxFck2Sync[7]), .A1(n2586), .Z(n2516));
Q_MX02 U3047 ( .S(evalOnC), .A0(maxFck2Sync[6]), .A1(n2588), .Z(n2517));
Q_MX02 U3048 ( .S(evalOnC), .A0(maxFck2Sync[5]), .A1(n2590), .Z(n2518));
Q_MX02 U3049 ( .S(evalOnC), .A0(maxFck2Sync[4]), .A1(n2592), .Z(n2519));
Q_MX02 U3050 ( .S(evalOnC), .A0(maxFck2Sync[3]), .A1(n2594), .Z(n2520));
Q_MX02 U3051 ( .S(evalOnC), .A0(maxFck2Sync[2]), .A1(n2596), .Z(n2521));
Q_MX02 U3052 ( .S(evalOnC), .A0(maxFck2Sync[1]), .A1(n2598), .Z(n2522));
Q_MX02 U3053 ( .S(evalOnC), .A0(maxFck2Sync[0]), .A1(n2599), .Z(n2523));
Q_MX02 U3054 ( .S(n2507), .A0(n2540), .A1(maxGfifo2Sync[15]), .Z(n2524));
Q_MX02 U3055 ( .S(n2507), .A0(n2542), .A1(maxGfifo2Sync[14]), .Z(n2525));
Q_MX02 U3056 ( .S(n2507), .A0(n2544), .A1(maxGfifo2Sync[13]), .Z(n2526));
Q_MX02 U3057 ( .S(n2507), .A0(n2546), .A1(maxGfifo2Sync[12]), .Z(n2527));
Q_MX02 U3058 ( .S(n2507), .A0(n2548), .A1(maxGfifo2Sync[11]), .Z(n2528));
Q_MX02 U3059 ( .S(n2507), .A0(n2550), .A1(maxGfifo2Sync[10]), .Z(n2529));
Q_MX02 U3060 ( .S(n2507), .A0(n2552), .A1(maxGfifo2Sync[9]), .Z(n2530));
Q_MX02 U3061 ( .S(n2507), .A0(n2554), .A1(maxGfifo2Sync[8]), .Z(n2531));
Q_MX02 U3062 ( .S(n2507), .A0(n2556), .A1(maxGfifo2Sync[7]), .Z(n2532));
Q_MX02 U3063 ( .S(n2507), .A0(n2558), .A1(maxGfifo2Sync[6]), .Z(n2533));
Q_MX02 U3064 ( .S(n2507), .A0(n2560), .A1(maxGfifo2Sync[5]), .Z(n2534));
Q_MX02 U3065 ( .S(n2507), .A0(n2562), .A1(maxGfifo2Sync[4]), .Z(n2535));
Q_MX02 U3066 ( .S(n2507), .A0(n2564), .A1(maxGfifo2Sync[3]), .Z(n2536));
Q_MX02 U3067 ( .S(n2507), .A0(n2566), .A1(maxGfifo2Sync[2]), .Z(n2537));
Q_MX02 U3068 ( .S(n2507), .A0(n2568), .A1(maxGfifo2Sync[1]), .Z(n2538));
Q_MX02 U3069 ( .S(n2507), .A0(n2569), .A1(maxGfifo2Sync[0]), .Z(n2539));
Q_XNR2 U3070 ( .A0(Gfifo2Sync[15]), .A1(n2541), .Z(n2540));
Q_OR02 U3071 ( .A0(Gfifo2Sync[14]), .A1(n2543), .Z(n2541));
Q_XNR2 U3072 ( .A0(Gfifo2Sync[14]), .A1(n2543), .Z(n2542));
Q_OR02 U3073 ( .A0(Gfifo2Sync[13]), .A1(n2545), .Z(n2543));
Q_XNR2 U3074 ( .A0(Gfifo2Sync[13]), .A1(n2545), .Z(n2544));
Q_OR02 U3075 ( .A0(Gfifo2Sync[12]), .A1(n2547), .Z(n2545));
Q_XNR2 U3076 ( .A0(Gfifo2Sync[12]), .A1(n2547), .Z(n2546));
Q_OR02 U3077 ( .A0(Gfifo2Sync[11]), .A1(n2549), .Z(n2547));
Q_XNR2 U3078 ( .A0(Gfifo2Sync[11]), .A1(n2549), .Z(n2548));
Q_OR02 U3079 ( .A0(Gfifo2Sync[10]), .A1(n2551), .Z(n2549));
Q_XNR2 U3080 ( .A0(Gfifo2Sync[10]), .A1(n2551), .Z(n2550));
Q_OR02 U3081 ( .A0(Gfifo2Sync[9]), .A1(n2553), .Z(n2551));
Q_XNR2 U3082 ( .A0(Gfifo2Sync[9]), .A1(n2553), .Z(n2552));
Q_OR02 U3083 ( .A0(Gfifo2Sync[8]), .A1(n2555), .Z(n2553));
Q_XNR2 U3084 ( .A0(Gfifo2Sync[8]), .A1(n2555), .Z(n2554));
Q_OR02 U3085 ( .A0(Gfifo2Sync[7]), .A1(n2557), .Z(n2555));
Q_XNR2 U3086 ( .A0(Gfifo2Sync[7]), .A1(n2557), .Z(n2556));
Q_OR02 U3087 ( .A0(Gfifo2Sync[6]), .A1(n2559), .Z(n2557));
Q_XNR2 U3088 ( .A0(Gfifo2Sync[6]), .A1(n2559), .Z(n2558));
Q_OR02 U3089 ( .A0(Gfifo2Sync[5]), .A1(n2561), .Z(n2559));
Q_XNR2 U3090 ( .A0(Gfifo2Sync[5]), .A1(n2561), .Z(n2560));
Q_OR02 U3091 ( .A0(Gfifo2Sync[4]), .A1(n2563), .Z(n2561));
Q_XNR2 U3092 ( .A0(Gfifo2Sync[4]), .A1(n2563), .Z(n2562));
Q_OR02 U3093 ( .A0(Gfifo2Sync[3]), .A1(n2565), .Z(n2563));
Q_XNR2 U3094 ( .A0(Gfifo2Sync[3]), .A1(n2565), .Z(n2564));
Q_OR02 U3095 ( .A0(Gfifo2Sync[2]), .A1(n2567), .Z(n2565));
Q_XNR2 U3096 ( .A0(Gfifo2Sync[2]), .A1(n2567), .Z(n2566));
Q_OR02 U3097 ( .A0(Gfifo2Sync[1]), .A1(Gfifo2Sync[0]), .Z(n2567));
Q_XNR2 U3098 ( .A0(Gfifo2Sync[1]), .A1(Gfifo2Sync[0]), .Z(n2568));
Q_XNR2 U3099 ( .A0(Fck2Sync[15]), .A1(n2571), .Z(n2570));
Q_OR02 U3100 ( .A0(Fck2Sync[14]), .A1(n2573), .Z(n2571));
Q_XNR2 U3101 ( .A0(Fck2Sync[14]), .A1(n2573), .Z(n2572));
Q_OR02 U3102 ( .A0(Fck2Sync[13]), .A1(n2575), .Z(n2573));
Q_XNR2 U3103 ( .A0(Fck2Sync[13]), .A1(n2575), .Z(n2574));
Q_OR02 U3104 ( .A0(Fck2Sync[12]), .A1(n2577), .Z(n2575));
Q_XNR2 U3105 ( .A0(Fck2Sync[12]), .A1(n2577), .Z(n2576));
Q_OR02 U3106 ( .A0(Fck2Sync[11]), .A1(n2579), .Z(n2577));
Q_XNR2 U3107 ( .A0(Fck2Sync[11]), .A1(n2579), .Z(n2578));
Q_OR02 U3108 ( .A0(Fck2Sync[10]), .A1(n2581), .Z(n2579));
Q_XNR2 U3109 ( .A0(Fck2Sync[10]), .A1(n2581), .Z(n2580));
Q_OR02 U3110 ( .A0(Fck2Sync[9]), .A1(n2583), .Z(n2581));
Q_XNR2 U3111 ( .A0(Fck2Sync[9]), .A1(n2583), .Z(n2582));
Q_OR02 U3112 ( .A0(Fck2Sync[8]), .A1(n2585), .Z(n2583));
Q_XNR2 U3113 ( .A0(Fck2Sync[8]), .A1(n2585), .Z(n2584));
Q_OR02 U3114 ( .A0(Fck2Sync[7]), .A1(n2587), .Z(n2585));
Q_XNR2 U3115 ( .A0(Fck2Sync[7]), .A1(n2587), .Z(n2586));
Q_OR02 U3116 ( .A0(Fck2Sync[6]), .A1(n2589), .Z(n2587));
Q_XNR2 U3117 ( .A0(Fck2Sync[6]), .A1(n2589), .Z(n2588));
Q_OR02 U3118 ( .A0(Fck2Sync[5]), .A1(n2591), .Z(n2589));
Q_XNR2 U3119 ( .A0(Fck2Sync[5]), .A1(n2591), .Z(n2590));
Q_OR02 U3120 ( .A0(Fck2Sync[4]), .A1(n2593), .Z(n2591));
Q_XNR2 U3121 ( .A0(Fck2Sync[4]), .A1(n2593), .Z(n2592));
Q_OR02 U3122 ( .A0(Fck2Sync[3]), .A1(n2595), .Z(n2593));
Q_XNR2 U3123 ( .A0(Fck2Sync[3]), .A1(n2595), .Z(n2594));
Q_OR02 U3124 ( .A0(Fck2Sync[2]), .A1(n2597), .Z(n2595));
Q_XNR2 U3125 ( .A0(Fck2Sync[2]), .A1(n2597), .Z(n2596));
Q_OR02 U3126 ( .A0(Fck2Sync[1]), .A1(Fck2Sync[0]), .Z(n2597));
Q_XNR2 U3127 ( .A0(Fck2Sync[1]), .A1(Fck2Sync[0]), .Z(n2598));
Q_OR03 U3128 ( .A0(n2601), .A1(n2600), .A2(n2507), .Z(n2505));
Q_OR03 U3129 ( .A0(n2604), .A1(n2603), .A2(n2602), .Z(n2600));
Q_OR03 U3130 ( .A0(Gfifo2Sync[0]), .A1(n2606), .A2(n2605), .Z(n2601));
Q_OR03 U3131 ( .A0(Gfifo2Sync[3]), .A1(Gfifo2Sync[2]), .A2(Gfifo2Sync[1]), .Z(n2602));
Q_OR03 U3132 ( .A0(Gfifo2Sync[6]), .A1(Gfifo2Sync[5]), .A2(Gfifo2Sync[4]), .Z(n2603));
Q_OR03 U3133 ( .A0(Gfifo2Sync[9]), .A1(Gfifo2Sync[8]), .A2(Gfifo2Sync[7]), .Z(n2604));
Q_OR03 U3134 ( .A0(Gfifo2Sync[12]), .A1(Gfifo2Sync[11]), .A2(Gfifo2Sync[10]), .Z(n2605));
Q_OR03 U3135 ( .A0(Gfifo2Sync[15]), .A1(Gfifo2Sync[14]), .A2(Gfifo2Sync[13]), .Z(n2606));
Q_OR03 U3136 ( .A0(n2608), .A1(n2607), .A2(n402), .Z(n2506));
Q_OR03 U3137 ( .A0(n2611), .A1(n2610), .A2(n2609), .Z(n2607));
Q_OR03 U3138 ( .A0(Fck2Sync[0]), .A1(n2613), .A2(n2612), .Z(n2608));
Q_OR03 U3139 ( .A0(Fck2Sync[3]), .A1(Fck2Sync[2]), .A2(Fck2Sync[1]), .Z(n2609));
Q_OR03 U3140 ( .A0(Fck2Sync[6]), .A1(Fck2Sync[5]), .A2(Fck2Sync[4]), .Z(n2610));
Q_OR03 U3141 ( .A0(Fck2Sync[9]), .A1(Fck2Sync[8]), .A2(Fck2Sync[7]), .Z(n2611));
Q_OR03 U3142 ( .A0(Fck2Sync[12]), .A1(Fck2Sync[11]), .A2(Fck2Sync[10]), .Z(n2612));
Q_OR03 U3143 ( .A0(Fck2Sync[15]), .A1(Fck2Sync[14]), .A2(Fck2Sync[13]), .Z(n2613));
Q_OA21 U3144 ( .A0(hwClkDbgEn), .A1(cakeUcEnable), .B0(hwClkDbg), .Z(hwClkDbgOn));
Q_INV U3145 ( .A(it_newBuf), .Z(n2614));
Q_LSN01 U3146 ( .S(n2614), .R(n1162), .Q(it_newBufPO), .QN( ));
Q_INV U3147 ( .A(callEmuEv), .Z(n2616));
Q_NR02 U3148 ( .A0(callEmuEv), .A1(hasGFIFO1), .Z(n2618));
Q_NR02 U3149 ( .A0(hasGFIFO2), .A1(hasSFIFO), .Z(n2619));
Q_INV U3150 ( .A(hasPTX), .Z(n2617));
Q_AN03 U3151 ( .A0(n2618), .A1(n2617), .A2(n2619), .Z(n2615));
Q_NR02 U3152 ( .A0(n2615), .A1(callEmuEv), .Z(n2620));
Q_MX02 U3153 ( .S(n2615), .A0(n2620), .A1(mioPOW_2[1]), .Z(intr));
Q_INV U3154 ( .A(evalOnD), .Z(n2622));
Q_AN02 U3155 ( .A0(n1165), .A1(n2622), .Z(n2623));
Q_INV U3156 ( .A(n2623), .Z(n2621));
Q_AD01HF U3157 ( .A0(fvSCount[62]), .B0(n2626), .S(n2625), .CO(n2624));
Q_AD01HF U3158 ( .A0(fvSCount[61]), .B0(n2628), .S(n2627), .CO(n2626));
Q_AD01HF U3159 ( .A0(fvSCount[60]), .B0(n2630), .S(n2629), .CO(n2628));
Q_AD01HF U3160 ( .A0(fvSCount[59]), .B0(n2632), .S(n2631), .CO(n2630));
Q_AD01HF U3161 ( .A0(fvSCount[58]), .B0(n2634), .S(n2633), .CO(n2632));
Q_AD01HF U3162 ( .A0(fvSCount[57]), .B0(n2636), .S(n2635), .CO(n2634));
Q_AD01HF U3163 ( .A0(fvSCount[56]), .B0(n2638), .S(n2637), .CO(n2636));
Q_AD01HF U3164 ( .A0(fvSCount[55]), .B0(n2640), .S(n2639), .CO(n2638));
Q_AD01HF U3165 ( .A0(fvSCount[54]), .B0(n2642), .S(n2641), .CO(n2640));
Q_AD01HF U3166 ( .A0(fvSCount[53]), .B0(n2644), .S(n2643), .CO(n2642));
Q_AD01HF U3167 ( .A0(fvSCount[52]), .B0(n2646), .S(n2645), .CO(n2644));
Q_AD01HF U3168 ( .A0(fvSCount[51]), .B0(n2648), .S(n2647), .CO(n2646));
Q_AD01HF U3169 ( .A0(fvSCount[50]), .B0(n2650), .S(n2649), .CO(n2648));
Q_AD01HF U3170 ( .A0(fvSCount[49]), .B0(n2652), .S(n2651), .CO(n2650));
Q_AD01HF U3171 ( .A0(fvSCount[48]), .B0(n2654), .S(n2653), .CO(n2652));
Q_AD01HF U3172 ( .A0(fvSCount[47]), .B0(n2656), .S(n2655), .CO(n2654));
Q_AD01HF U3173 ( .A0(fvSCount[46]), .B0(n2658), .S(n2657), .CO(n2656));
Q_AD01HF U3174 ( .A0(fvSCount[45]), .B0(n2660), .S(n2659), .CO(n2658));
Q_AD01HF U3175 ( .A0(fvSCount[44]), .B0(n2662), .S(n2661), .CO(n2660));
Q_AD01HF U3176 ( .A0(fvSCount[43]), .B0(n2664), .S(n2663), .CO(n2662));
Q_AD01HF U3177 ( .A0(fvSCount[42]), .B0(n2666), .S(n2665), .CO(n2664));
Q_AD01HF U3178 ( .A0(fvSCount[41]), .B0(n2668), .S(n2667), .CO(n2666));
Q_AD01HF U3179 ( .A0(fvSCount[40]), .B0(n2670), .S(n2669), .CO(n2668));
Q_AD01HF U3180 ( .A0(fvSCount[39]), .B0(n2672), .S(n2671), .CO(n2670));
Q_AD01HF U3181 ( .A0(fvSCount[38]), .B0(n2674), .S(n2673), .CO(n2672));
Q_AD01HF U3182 ( .A0(fvSCount[37]), .B0(n2676), .S(n2675), .CO(n2674));
Q_AD01HF U3183 ( .A0(fvSCount[36]), .B0(n2678), .S(n2677), .CO(n2676));
Q_AD01HF U3184 ( .A0(fvSCount[35]), .B0(n2680), .S(n2679), .CO(n2678));
Q_AD01HF U3185 ( .A0(fvSCount[34]), .B0(n2682), .S(n2681), .CO(n2680));
Q_AD01HF U3186 ( .A0(fvSCount[33]), .B0(n2684), .S(n2683), .CO(n2682));
Q_AD01HF U3187 ( .A0(fvSCount[32]), .B0(n2686), .S(n2685), .CO(n2684));
Q_AD01HF U3188 ( .A0(fvSCount[31]), .B0(n2688), .S(n2687), .CO(n2686));
Q_AD01HF U3189 ( .A0(fvSCount[30]), .B0(n2690), .S(n2689), .CO(n2688));
Q_AD01HF U3190 ( .A0(fvSCount[29]), .B0(n2692), .S(n2691), .CO(n2690));
Q_AD01HF U3191 ( .A0(fvSCount[28]), .B0(n2694), .S(n2693), .CO(n2692));
Q_AD01HF U3192 ( .A0(fvSCount[27]), .B0(n2696), .S(n2695), .CO(n2694));
Q_AD01HF U3193 ( .A0(fvSCount[26]), .B0(n2698), .S(n2697), .CO(n2696));
Q_AD01HF U3194 ( .A0(fvSCount[25]), .B0(n2700), .S(n2699), .CO(n2698));
Q_AD01HF U3195 ( .A0(fvSCount[24]), .B0(n2702), .S(n2701), .CO(n2700));
Q_AD01HF U3196 ( .A0(fvSCount[23]), .B0(n2704), .S(n2703), .CO(n2702));
Q_AD01HF U3197 ( .A0(fvSCount[22]), .B0(n2706), .S(n2705), .CO(n2704));
Q_AD01HF U3198 ( .A0(fvSCount[21]), .B0(n2708), .S(n2707), .CO(n2706));
Q_AD01HF U3199 ( .A0(fvSCount[20]), .B0(n2710), .S(n2709), .CO(n2708));
Q_AD01HF U3200 ( .A0(fvSCount[19]), .B0(n2712), .S(n2711), .CO(n2710));
Q_AD01HF U3201 ( .A0(fvSCount[18]), .B0(n2714), .S(n2713), .CO(n2712));
Q_AD01HF U3202 ( .A0(fvSCount[17]), .B0(n2716), .S(n2715), .CO(n2714));
Q_AD01HF U3203 ( .A0(fvSCount[16]), .B0(n2718), .S(n2717), .CO(n2716));
Q_AD01HF U3204 ( .A0(fvSCount[15]), .B0(n2720), .S(n2719), .CO(n2718));
Q_AD01HF U3205 ( .A0(fvSCount[14]), .B0(n2722), .S(n2721), .CO(n2720));
Q_AD01HF U3206 ( .A0(fvSCount[13]), .B0(n2724), .S(n2723), .CO(n2722));
Q_AD01HF U3207 ( .A0(fvSCount[12]), .B0(n2726), .S(n2725), .CO(n2724));
Q_AD01HF U3208 ( .A0(fvSCount[11]), .B0(n2728), .S(n2727), .CO(n2726));
Q_AD01HF U3209 ( .A0(fvSCount[10]), .B0(n2730), .S(n2729), .CO(n2728));
Q_AD01HF U3210 ( .A0(fvSCount[9]), .B0(n2732), .S(n2731), .CO(n2730));
Q_AD01HF U3211 ( .A0(fvSCount[8]), .B0(n2734), .S(n2733), .CO(n2732));
Q_AD01HF U3212 ( .A0(fvSCount[7]), .B0(n2736), .S(n2735), .CO(n2734));
Q_AD01HF U3213 ( .A0(fvSCount[6]), .B0(n2738), .S(n2737), .CO(n2736));
Q_AD01HF U3214 ( .A0(fvSCount[5]), .B0(n2740), .S(n2739), .CO(n2738));
Q_AD01HF U3215 ( .A0(fvSCount[4]), .B0(n2742), .S(n2741), .CO(n2740));
Q_AD01HF U3216 ( .A0(fvSCount[3]), .B0(n2744), .S(n2743), .CO(n2742));
Q_AD01HF U3217 ( .A0(fvSCount[2]), .B0(n2746), .S(n2745), .CO(n2744));
Q_AD01HF U3218 ( .A0(fvSCount[1]), .B0(fvSCount[0]), .S(n2747), .CO(n2746));
Q_AD01HF U3219 ( .A0(evfCount[62]), .B0(n2750), .S(n2749), .CO(n2748));
Q_AD01HF U3220 ( .A0(evfCount[61]), .B0(n2752), .S(n2751), .CO(n2750));
Q_AD01HF U3221 ( .A0(evfCount[60]), .B0(n2754), .S(n2753), .CO(n2752));
Q_AD01HF U3222 ( .A0(evfCount[59]), .B0(n2756), .S(n2755), .CO(n2754));
Q_AD01HF U3223 ( .A0(evfCount[58]), .B0(n2758), .S(n2757), .CO(n2756));
Q_AD01HF U3224 ( .A0(evfCount[57]), .B0(n2760), .S(n2759), .CO(n2758));
Q_AD01HF U3225 ( .A0(evfCount[56]), .B0(n2762), .S(n2761), .CO(n2760));
Q_AD01HF U3226 ( .A0(evfCount[55]), .B0(n2764), .S(n2763), .CO(n2762));
Q_AD01HF U3227 ( .A0(evfCount[54]), .B0(n2766), .S(n2765), .CO(n2764));
Q_AD01HF U3228 ( .A0(evfCount[53]), .B0(n2768), .S(n2767), .CO(n2766));
Q_AD01HF U3229 ( .A0(evfCount[52]), .B0(n2770), .S(n2769), .CO(n2768));
Q_AD01HF U3230 ( .A0(evfCount[51]), .B0(n2772), .S(n2771), .CO(n2770));
Q_AD01HF U3231 ( .A0(evfCount[50]), .B0(n2774), .S(n2773), .CO(n2772));
Q_AD01HF U3232 ( .A0(evfCount[49]), .B0(n2776), .S(n2775), .CO(n2774));
Q_AD01HF U3233 ( .A0(evfCount[48]), .B0(n2778), .S(n2777), .CO(n2776));
Q_AD01HF U3234 ( .A0(evfCount[47]), .B0(n2780), .S(n2779), .CO(n2778));
Q_AD01HF U3235 ( .A0(evfCount[46]), .B0(n2782), .S(n2781), .CO(n2780));
Q_AD01HF U3236 ( .A0(evfCount[45]), .B0(n2784), .S(n2783), .CO(n2782));
Q_AD01HF U3237 ( .A0(evfCount[44]), .B0(n2786), .S(n2785), .CO(n2784));
Q_AD01HF U3238 ( .A0(evfCount[43]), .B0(n2788), .S(n2787), .CO(n2786));
Q_AD01HF U3239 ( .A0(evfCount[42]), .B0(n2790), .S(n2789), .CO(n2788));
Q_AD01HF U3240 ( .A0(evfCount[41]), .B0(n2792), .S(n2791), .CO(n2790));
Q_AD01HF U3241 ( .A0(evfCount[40]), .B0(n2794), .S(n2793), .CO(n2792));
Q_AD01HF U3242 ( .A0(evfCount[39]), .B0(n2796), .S(n2795), .CO(n2794));
Q_AD01HF U3243 ( .A0(evfCount[38]), .B0(n2798), .S(n2797), .CO(n2796));
Q_AD01HF U3244 ( .A0(evfCount[37]), .B0(n2800), .S(n2799), .CO(n2798));
Q_AD01HF U3245 ( .A0(evfCount[36]), .B0(n2802), .S(n2801), .CO(n2800));
Q_AD01HF U3246 ( .A0(evfCount[35]), .B0(n2804), .S(n2803), .CO(n2802));
Q_AD01HF U3247 ( .A0(evfCount[34]), .B0(n2806), .S(n2805), .CO(n2804));
Q_AD01HF U3248 ( .A0(evfCount[33]), .B0(n2808), .S(n2807), .CO(n2806));
Q_AD01HF U3249 ( .A0(evfCount[32]), .B0(n2810), .S(n2809), .CO(n2808));
Q_AD01HF U3250 ( .A0(evfCount[31]), .B0(n2812), .S(n2811), .CO(n2810));
Q_AD01HF U3251 ( .A0(evfCount[30]), .B0(n2814), .S(n2813), .CO(n2812));
Q_AD01HF U3252 ( .A0(evfCount[29]), .B0(n2816), .S(n2815), .CO(n2814));
Q_AD01HF U3253 ( .A0(evfCount[28]), .B0(n2818), .S(n2817), .CO(n2816));
Q_AD01HF U3254 ( .A0(evfCount[27]), .B0(n2820), .S(n2819), .CO(n2818));
Q_AD01HF U3255 ( .A0(evfCount[26]), .B0(n2822), .S(n2821), .CO(n2820));
Q_AD01HF U3256 ( .A0(evfCount[25]), .B0(n2824), .S(n2823), .CO(n2822));
Q_AD01HF U3257 ( .A0(evfCount[24]), .B0(n2826), .S(n2825), .CO(n2824));
Q_AD01HF U3258 ( .A0(evfCount[23]), .B0(n2828), .S(n2827), .CO(n2826));
Q_AD01HF U3259 ( .A0(evfCount[22]), .B0(n2830), .S(n2829), .CO(n2828));
Q_AD01HF U3260 ( .A0(evfCount[21]), .B0(n2832), .S(n2831), .CO(n2830));
Q_AD01HF U3261 ( .A0(evfCount[20]), .B0(n2834), .S(n2833), .CO(n2832));
Q_AD01HF U3262 ( .A0(evfCount[19]), .B0(n2836), .S(n2835), .CO(n2834));
Q_AD01HF U3263 ( .A0(evfCount[18]), .B0(n2838), .S(n2837), .CO(n2836));
Q_AD01HF U3264 ( .A0(evfCount[17]), .B0(n2840), .S(n2839), .CO(n2838));
Q_AD01HF U3265 ( .A0(evfCount[16]), .B0(n2842), .S(n2841), .CO(n2840));
Q_AD01HF U3266 ( .A0(evfCount[15]), .B0(n2844), .S(n2843), .CO(n2842));
Q_AD01HF U3267 ( .A0(evfCount[14]), .B0(n2846), .S(n2845), .CO(n2844));
Q_AD01HF U3268 ( .A0(evfCount[13]), .B0(n2848), .S(n2847), .CO(n2846));
Q_AD01HF U3269 ( .A0(evfCount[12]), .B0(n2850), .S(n2849), .CO(n2848));
Q_AD01HF U3270 ( .A0(evfCount[11]), .B0(n2852), .S(n2851), .CO(n2850));
Q_AD01HF U3271 ( .A0(evfCount[10]), .B0(n2854), .S(n2853), .CO(n2852));
Q_AD01HF U3272 ( .A0(evfCount[9]), .B0(n2856), .S(n2855), .CO(n2854));
Q_AD01HF U3273 ( .A0(evfCount[8]), .B0(n2858), .S(n2857), .CO(n2856));
Q_AD01HF U3274 ( .A0(evfCount[7]), .B0(n2860), .S(n2859), .CO(n2858));
Q_AD01HF U3275 ( .A0(evfCount[6]), .B0(n2862), .S(n2861), .CO(n2860));
Q_AD01HF U3276 ( .A0(evfCount[5]), .B0(n2864), .S(n2863), .CO(n2862));
Q_AD01HF U3277 ( .A0(evfCount[4]), .B0(n2866), .S(n2865), .CO(n2864));
Q_AD01HF U3278 ( .A0(evfCount[3]), .B0(n2868), .S(n2867), .CO(n2866));
Q_AD01HF U3279 ( .A0(evfCount[2]), .B0(n2870), .S(n2869), .CO(n2868));
Q_AD01HF U3280 ( .A0(evfCount[1]), .B0(evfCount[0]), .S(n2871), .CO(n2870));
Q_AD01HF U3281 ( .A0(eCount[1]), .B0(eCount[0]), .S(n2873), .CO(n2874));
Q_AD01HF U3282 ( .A0(eCount[2]), .B0(n2874), .S(n2875), .CO(n2876));
Q_AD01HF U3283 ( .A0(eCount[3]), .B0(n2876), .S(n2877), .CO(n2878));
Q_AD01HF U3284 ( .A0(eCount[4]), .B0(n2878), .S(n2879), .CO(n2880));
Q_AD01HF U3285 ( .A0(eCount[5]), .B0(n2880), .S(n2881), .CO(n2882));
Q_AD01HF U3286 ( .A0(eCount[6]), .B0(n2882), .S(n2883), .CO(n2884));
Q_AD01HF U3287 ( .A0(eCount[7]), .B0(n2884), .S(n2885), .CO(n2886));
Q_AD01HF U3288 ( .A0(eCount[8]), .B0(n2886), .S(n2887), .CO(n2888));
Q_AD01HF U3289 ( .A0(eCount[9]), .B0(n2888), .S(n2889), .CO(n2890));
Q_AD01HF U3290 ( .A0(eCount[10]), .B0(n2890), .S(n2891), .CO(n2892));
Q_AD01HF U3291 ( .A0(eCount[11]), .B0(n2892), .S(n2893), .CO(n2894));
Q_AD01HF U3292 ( .A0(eCount[12]), .B0(n2894), .S(n2895), .CO(n2896));
Q_AD01HF U3293 ( .A0(eCount[13]), .B0(n2896), .S(n2897), .CO(n2898));
Q_AD01HF U3294 ( .A0(eCount[14]), .B0(n2898), .S(n2899), .CO(n2900));
Q_AD01HF U3295 ( .A0(eCount[15]), .B0(n2900), .S(n2901), .CO(n2902));
Q_AD01HF U3296 ( .A0(eCount[16]), .B0(n2902), .S(n2903), .CO(n2904));
Q_AD01HF U3297 ( .A0(eCount[17]), .B0(n2904), .S(n2905), .CO(n2906));
Q_AD01HF U3298 ( .A0(eCount[18]), .B0(n2906), .S(n2907), .CO(n2908));
Q_AD01HF U3299 ( .A0(eCount[19]), .B0(n2908), .S(n2909), .CO(n2910));
Q_AD01HF U3300 ( .A0(eCount[20]), .B0(n2910), .S(n2911), .CO(n2912));
Q_AD01HF U3301 ( .A0(eCount[21]), .B0(n2912), .S(n2913), .CO(n2914));
Q_AD01HF U3302 ( .A0(eCount[22]), .B0(n2914), .S(n2915), .CO(n2916));
Q_AD01HF U3303 ( .A0(eCount[23]), .B0(n2916), .S(n2917), .CO(n2918));
Q_AD01HF U3304 ( .A0(eCount[24]), .B0(n2918), .S(n2919), .CO(n2920));
Q_AD01HF U3305 ( .A0(eCount[25]), .B0(n2920), .S(n2921), .CO(n2922));
Q_AD01HF U3306 ( .A0(eCount[26]), .B0(n2922), .S(n2923), .CO(n2924));
Q_AD01HF U3307 ( .A0(eCount[27]), .B0(n2924), .S(n2925), .CO(n2926));
Q_AD01HF U3308 ( .A0(eCount[28]), .B0(n2926), .S(n2927), .CO(n2928));
Q_AD01HF U3309 ( .A0(eCount[29]), .B0(n2928), .S(n2929), .CO(n2930));
Q_AD01HF U3310 ( .A0(eCount[30]), .B0(n2930), .S(n2931), .CO(n2932));
Q_AD01HF U3311 ( .A0(eCount[31]), .B0(n2932), .S(n2933), .CO(n2934));
Q_AD01HF U3312 ( .A0(eCount[32]), .B0(n2934), .S(n2935), .CO(n2936));
Q_AD01HF U3313 ( .A0(eCount[33]), .B0(n2936), .S(n2937), .CO(n2938));
Q_AD01HF U3314 ( .A0(eCount[34]), .B0(n2938), .S(n2939), .CO(n2940));
Q_AD01HF U3315 ( .A0(eCount[35]), .B0(n2940), .S(n2941), .CO(n2942));
Q_AD01HF U3316 ( .A0(eCount[36]), .B0(n2942), .S(n2943), .CO(n2944));
Q_AD01HF U3317 ( .A0(eCount[37]), .B0(n2944), .S(n2945), .CO(n2946));
Q_AD01HF U3318 ( .A0(eCount[38]), .B0(n2946), .S(n2947), .CO(n2948));
Q_AD01HF U3319 ( .A0(eCount[39]), .B0(n2948), .S(n2949), .CO(n2950));
Q_AD01HF U3320 ( .A0(eCount[40]), .B0(n2950), .S(n2951), .CO(n2952));
Q_AD01HF U3321 ( .A0(eCount[41]), .B0(n2952), .S(n2953), .CO(n2954));
Q_AD01HF U3322 ( .A0(eCount[42]), .B0(n2954), .S(n2955), .CO(n2956));
Q_AD01HF U3323 ( .A0(eCount[43]), .B0(n2956), .S(n2957), .CO(n2958));
Q_AD01HF U3324 ( .A0(eCount[44]), .B0(n2958), .S(n2959), .CO(n2960));
Q_AD01HF U3325 ( .A0(eCount[45]), .B0(n2960), .S(n2961), .CO(n2962));
Q_AD01HF U3326 ( .A0(eCount[46]), .B0(n2962), .S(n2963), .CO(n2964));
Q_AD01HF U3327 ( .A0(eCount[47]), .B0(n2964), .S(n2965), .CO(n2966));
Q_AD01HF U3328 ( .A0(eCount[48]), .B0(n2966), .S(n2967), .CO(n2968));
Q_AD01HF U3329 ( .A0(eCount[49]), .B0(n2968), .S(n2969), .CO(n2970));
Q_AD01HF U3330 ( .A0(eCount[50]), .B0(n2970), .S(n2971), .CO(n2972));
Q_AD01HF U3331 ( .A0(eCount[51]), .B0(n2972), .S(n2973), .CO(n2974));
Q_AD01HF U3332 ( .A0(eCount[52]), .B0(n2974), .S(n2975), .CO(n2976));
Q_AD01HF U3333 ( .A0(eCount[53]), .B0(n2976), .S(n2977), .CO(n2978));
Q_AD01HF U3334 ( .A0(eCount[54]), .B0(n2978), .S(n2979), .CO(n2980));
Q_AD01HF U3335 ( .A0(eCount[55]), .B0(n2980), .S(n2981), .CO(n2982));
Q_AD01HF U3336 ( .A0(eCount[56]), .B0(n2982), .S(n2983), .CO(n2984));
Q_AD01HF U3337 ( .A0(eCount[57]), .B0(n2984), .S(n2985), .CO(n2986));
Q_AD01HF U3338 ( .A0(eCount[58]), .B0(n2986), .S(n2987), .CO(n2988));
Q_AD01HF U3339 ( .A0(eCount[59]), .B0(n2988), .S(n2989), .CO(n2990));
Q_AD01HF U3340 ( .A0(eCount[60]), .B0(n2990), .S(n2991), .CO(n2992));
Q_AD01HF U3341 ( .A0(eCount[61]), .B0(n2992), .S(n2993), .CO(n2994));
Q_AD01HF U3342 ( .A0(eCount[62]), .B0(n2994), .S(n2995), .CO(n2996));
Q_FDP0 \eCount_REG[62] ( .CK(eClk), .D(n2995), .Q(eCount[62]), .QN( ));
Q_FDP0 \eCount_REG[61] ( .CK(eClk), .D(n2993), .Q(eCount[61]), .QN( ));
Q_FDP0 \eCount_REG[60] ( .CK(eClk), .D(n2991), .Q(eCount[60]), .QN( ));
Q_FDP0 \eCount_REG[59] ( .CK(eClk), .D(n2989), .Q(eCount[59]), .QN( ));
Q_FDP0 \eCount_REG[58] ( .CK(eClk), .D(n2987), .Q(eCount[58]), .QN( ));
Q_FDP0 \eCount_REG[57] ( .CK(eClk), .D(n2985), .Q(eCount[57]), .QN( ));
Q_FDP0 \eCount_REG[56] ( .CK(eClk), .D(n2983), .Q(eCount[56]), .QN( ));
Q_FDP0 \eCount_REG[55] ( .CK(eClk), .D(n2981), .Q(eCount[55]), .QN( ));
Q_FDP0 \eCount_REG[54] ( .CK(eClk), .D(n2979), .Q(eCount[54]), .QN( ));
Q_FDP0 \eCount_REG[53] ( .CK(eClk), .D(n2977), .Q(eCount[53]), .QN( ));
Q_FDP0 \eCount_REG[52] ( .CK(eClk), .D(n2975), .Q(eCount[52]), .QN( ));
Q_FDP0 \eCount_REG[51] ( .CK(eClk), .D(n2973), .Q(eCount[51]), .QN( ));
Q_FDP0 \eCount_REG[50] ( .CK(eClk), .D(n2971), .Q(eCount[50]), .QN( ));
Q_FDP0 \eCount_REG[49] ( .CK(eClk), .D(n2969), .Q(eCount[49]), .QN( ));
Q_FDP0 \eCount_REG[48] ( .CK(eClk), .D(n2967), .Q(eCount[48]), .QN( ));
Q_FDP0 \eCount_REG[47] ( .CK(eClk), .D(n2965), .Q(eCount[47]), .QN( ));
Q_FDP0 \eCount_REG[46] ( .CK(eClk), .D(n2963), .Q(eCount[46]), .QN( ));
Q_FDP0 \eCount_REG[45] ( .CK(eClk), .D(n2961), .Q(eCount[45]), .QN( ));
Q_FDP0 \eCount_REG[44] ( .CK(eClk), .D(n2959), .Q(eCount[44]), .QN( ));
Q_FDP0 \eCount_REG[43] ( .CK(eClk), .D(n2957), .Q(eCount[43]), .QN( ));
Q_FDP0 \eCount_REG[42] ( .CK(eClk), .D(n2955), .Q(eCount[42]), .QN( ));
Q_FDP0 \eCount_REG[41] ( .CK(eClk), .D(n2953), .Q(eCount[41]), .QN( ));
Q_FDP0 \eCount_REG[40] ( .CK(eClk), .D(n2951), .Q(eCount[40]), .QN( ));
Q_FDP0 \eCount_REG[39] ( .CK(eClk), .D(n2949), .Q(eCount[39]), .QN( ));
Q_FDP0 \eCount_REG[38] ( .CK(eClk), .D(n2947), .Q(eCount[38]), .QN( ));
Q_FDP0 \eCount_REG[37] ( .CK(eClk), .D(n2945), .Q(eCount[37]), .QN( ));
Q_FDP0 \eCount_REG[36] ( .CK(eClk), .D(n2943), .Q(eCount[36]), .QN( ));
Q_FDP0 \eCount_REG[35] ( .CK(eClk), .D(n2941), .Q(eCount[35]), .QN( ));
Q_FDP0 \eCount_REG[34] ( .CK(eClk), .D(n2939), .Q(eCount[34]), .QN( ));
Q_FDP0 \eCount_REG[33] ( .CK(eClk), .D(n2937), .Q(eCount[33]), .QN( ));
Q_FDP0 \eCount_REG[32] ( .CK(eClk), .D(n2935), .Q(eCount[32]), .QN( ));
Q_FDP0 \eCount_REG[31] ( .CK(eClk), .D(n2933), .Q(eCount[31]), .QN( ));
Q_FDP0 \eCount_REG[30] ( .CK(eClk), .D(n2931), .Q(eCount[30]), .QN( ));
Q_FDP0 \eCount_REG[29] ( .CK(eClk), .D(n2929), .Q(eCount[29]), .QN( ));
Q_FDP0 \eCount_REG[28] ( .CK(eClk), .D(n2927), .Q(eCount[28]), .QN( ));
Q_FDP0 \eCount_REG[27] ( .CK(eClk), .D(n2925), .Q(eCount[27]), .QN( ));
Q_FDP0 \eCount_REG[26] ( .CK(eClk), .D(n2923), .Q(eCount[26]), .QN( ));
Q_FDP0 \eCount_REG[25] ( .CK(eClk), .D(n2921), .Q(eCount[25]), .QN( ));
Q_FDP0 \eCount_REG[24] ( .CK(eClk), .D(n2919), .Q(eCount[24]), .QN( ));
Q_FDP0 \eCount_REG[23] ( .CK(eClk), .D(n2917), .Q(eCount[23]), .QN( ));
Q_FDP0 \eCount_REG[22] ( .CK(eClk), .D(n2915), .Q(eCount[22]), .QN( ));
Q_FDP0 \eCount_REG[21] ( .CK(eClk), .D(n2913), .Q(eCount[21]), .QN( ));
Q_FDP0 \eCount_REG[20] ( .CK(eClk), .D(n2911), .Q(eCount[20]), .QN( ));
Q_FDP0 \eCount_REG[19] ( .CK(eClk), .D(n2909), .Q(eCount[19]), .QN( ));
Q_FDP0 \eCount_REG[18] ( .CK(eClk), .D(n2907), .Q(eCount[18]), .QN( ));
Q_FDP0 \eCount_REG[17] ( .CK(eClk), .D(n2905), .Q(eCount[17]), .QN( ));
Q_FDP0 \eCount_REG[16] ( .CK(eClk), .D(n2903), .Q(eCount[16]), .QN( ));
Q_FDP0 \eCount_REG[15] ( .CK(eClk), .D(n2901), .Q(eCount[15]), .QN( ));
Q_FDP0 \eCount_REG[14] ( .CK(eClk), .D(n2899), .Q(eCount[14]), .QN( ));
Q_FDP0 \eCount_REG[13] ( .CK(eClk), .D(n2897), .Q(eCount[13]), .QN( ));
Q_FDP0 \eCount_REG[12] ( .CK(eClk), .D(n2895), .Q(eCount[12]), .QN( ));
Q_FDP0 \eCount_REG[11] ( .CK(eClk), .D(n2893), .Q(eCount[11]), .QN( ));
Q_FDP0 \eCount_REG[10] ( .CK(eClk), .D(n2891), .Q(eCount[10]), .QN( ));
Q_FDP0 \eCount_REG[9] ( .CK(eClk), .D(n2889), .Q(eCount[9]), .QN( ));
Q_FDP0 \eCount_REG[8] ( .CK(eClk), .D(n2887), .Q(eCount[8]), .QN( ));
Q_FDP0 \eCount_REG[7] ( .CK(eClk), .D(n2885), .Q(eCount[7]), .QN( ));
Q_FDP0 \eCount_REG[6] ( .CK(eClk), .D(n2883), .Q(eCount[6]), .QN( ));
Q_FDP0 \eCount_REG[5] ( .CK(eClk), .D(n2881), .Q(eCount[5]), .QN( ));
Q_FDP0 \eCount_REG[4] ( .CK(eClk), .D(n2879), .Q(eCount[4]), .QN( ));
Q_FDP0 \eCount_REG[3] ( .CK(eClk), .D(n2877), .Q(eCount[3]), .QN( ));
Q_FDP0 \eCount_REG[2] ( .CK(eClk), .D(n2875), .Q(eCount[2]), .QN( ));
Q_FDP0 \eCount_REG[1] ( .CK(eClk), .D(n2873), .Q(eCount[1]), .QN( ));
Q_FDP0 \eCount_REG[0] ( .CK(eClk), .D(n2872), .Q(eCount[0]), .QN(n2872));
Q_AN02 U3406 ( .A0(ixcHoldClk), .A1(n2998), .Z(n2997));
Q_AD01HF U3407 ( .A0(ixcHoldSyncCnt[62]), .B0(n3001), .S(n3000), .CO(n2999));
Q_AD01HF U3408 ( .A0(ixcHoldSyncCnt[61]), .B0(n3003), .S(n3002), .CO(n3001));
Q_AD01HF U3409 ( .A0(ixcHoldSyncCnt[60]), .B0(n3005), .S(n3004), .CO(n3003));
Q_AD01HF U3410 ( .A0(ixcHoldSyncCnt[59]), .B0(n3007), .S(n3006), .CO(n3005));
Q_AD01HF U3411 ( .A0(ixcHoldSyncCnt[58]), .B0(n3009), .S(n3008), .CO(n3007));
Q_AD01HF U3412 ( .A0(ixcHoldSyncCnt[57]), .B0(n3011), .S(n3010), .CO(n3009));
Q_AD01HF U3413 ( .A0(ixcHoldSyncCnt[56]), .B0(n3013), .S(n3012), .CO(n3011));
Q_AD01HF U3414 ( .A0(ixcHoldSyncCnt[55]), .B0(n3015), .S(n3014), .CO(n3013));
Q_AD01HF U3415 ( .A0(ixcHoldSyncCnt[54]), .B0(n3017), .S(n3016), .CO(n3015));
Q_AD01HF U3416 ( .A0(ixcHoldSyncCnt[53]), .B0(n3019), .S(n3018), .CO(n3017));
Q_AD01HF U3417 ( .A0(ixcHoldSyncCnt[52]), .B0(n3021), .S(n3020), .CO(n3019));
Q_AD01HF U3418 ( .A0(ixcHoldSyncCnt[51]), .B0(n3023), .S(n3022), .CO(n3021));
Q_AD01HF U3419 ( .A0(ixcHoldSyncCnt[50]), .B0(n3025), .S(n3024), .CO(n3023));
Q_AD01HF U3420 ( .A0(ixcHoldSyncCnt[49]), .B0(n3027), .S(n3026), .CO(n3025));
Q_AD01HF U3421 ( .A0(ixcHoldSyncCnt[48]), .B0(n3029), .S(n3028), .CO(n3027));
Q_AD01HF U3422 ( .A0(ixcHoldSyncCnt[47]), .B0(n3031), .S(n3030), .CO(n3029));
Q_AD01HF U3423 ( .A0(ixcHoldSyncCnt[46]), .B0(n3033), .S(n3032), .CO(n3031));
Q_AD01HF U3424 ( .A0(ixcHoldSyncCnt[45]), .B0(n3035), .S(n3034), .CO(n3033));
Q_AD01HF U3425 ( .A0(ixcHoldSyncCnt[44]), .B0(n3037), .S(n3036), .CO(n3035));
Q_AD01HF U3426 ( .A0(ixcHoldSyncCnt[43]), .B0(n3039), .S(n3038), .CO(n3037));
Q_AD01HF U3427 ( .A0(ixcHoldSyncCnt[42]), .B0(n3041), .S(n3040), .CO(n3039));
Q_AD01HF U3428 ( .A0(ixcHoldSyncCnt[41]), .B0(n3043), .S(n3042), .CO(n3041));
Q_AD01HF U3429 ( .A0(ixcHoldSyncCnt[40]), .B0(n3045), .S(n3044), .CO(n3043));
Q_AD01HF U3430 ( .A0(ixcHoldSyncCnt[39]), .B0(n3047), .S(n3046), .CO(n3045));
Q_AD01HF U3431 ( .A0(ixcHoldSyncCnt[38]), .B0(n3049), .S(n3048), .CO(n3047));
Q_AD01HF U3432 ( .A0(ixcHoldSyncCnt[37]), .B0(n3051), .S(n3050), .CO(n3049));
Q_AD01HF U3433 ( .A0(ixcHoldSyncCnt[36]), .B0(n3053), .S(n3052), .CO(n3051));
Q_AD01HF U3434 ( .A0(ixcHoldSyncCnt[35]), .B0(n3055), .S(n3054), .CO(n3053));
Q_AD01HF U3435 ( .A0(ixcHoldSyncCnt[34]), .B0(n3057), .S(n3056), .CO(n3055));
Q_AD01HF U3436 ( .A0(ixcHoldSyncCnt[33]), .B0(n3059), .S(n3058), .CO(n3057));
Q_AD01HF U3437 ( .A0(ixcHoldSyncCnt[32]), .B0(n3061), .S(n3060), .CO(n3059));
Q_AD01HF U3438 ( .A0(ixcHoldSyncCnt[31]), .B0(n3063), .S(n3062), .CO(n3061));
Q_AD01HF U3439 ( .A0(ixcHoldSyncCnt[30]), .B0(n3065), .S(n3064), .CO(n3063));
Q_AD01HF U3440 ( .A0(ixcHoldSyncCnt[29]), .B0(n3067), .S(n3066), .CO(n3065));
Q_AD01HF U3441 ( .A0(ixcHoldSyncCnt[28]), .B0(n3069), .S(n3068), .CO(n3067));
Q_AD01HF U3442 ( .A0(ixcHoldSyncCnt[27]), .B0(n3071), .S(n3070), .CO(n3069));
Q_AD01HF U3443 ( .A0(ixcHoldSyncCnt[26]), .B0(n3073), .S(n3072), .CO(n3071));
Q_AD01HF U3444 ( .A0(ixcHoldSyncCnt[25]), .B0(n3075), .S(n3074), .CO(n3073));
Q_AD01HF U3445 ( .A0(ixcHoldSyncCnt[24]), .B0(n3077), .S(n3076), .CO(n3075));
Q_AD01HF U3446 ( .A0(ixcHoldSyncCnt[23]), .B0(n3079), .S(n3078), .CO(n3077));
Q_AD01HF U3447 ( .A0(ixcHoldSyncCnt[22]), .B0(n3081), .S(n3080), .CO(n3079));
Q_AD01HF U3448 ( .A0(ixcHoldSyncCnt[21]), .B0(n3083), .S(n3082), .CO(n3081));
Q_AD01HF U3449 ( .A0(ixcHoldSyncCnt[20]), .B0(n3085), .S(n3084), .CO(n3083));
Q_AD01HF U3450 ( .A0(ixcHoldSyncCnt[19]), .B0(n3087), .S(n3086), .CO(n3085));
Q_AD01HF U3451 ( .A0(ixcHoldSyncCnt[18]), .B0(n3089), .S(n3088), .CO(n3087));
Q_AD01HF U3452 ( .A0(ixcHoldSyncCnt[17]), .B0(n3091), .S(n3090), .CO(n3089));
Q_AD01HF U3453 ( .A0(ixcHoldSyncCnt[16]), .B0(n3093), .S(n3092), .CO(n3091));
Q_AD01HF U3454 ( .A0(ixcHoldSyncCnt[15]), .B0(n3095), .S(n3094), .CO(n3093));
Q_AD01HF U3455 ( .A0(ixcHoldSyncCnt[14]), .B0(n3097), .S(n3096), .CO(n3095));
Q_AD01HF U3456 ( .A0(ixcHoldSyncCnt[13]), .B0(n3099), .S(n3098), .CO(n3097));
Q_AD01HF U3457 ( .A0(ixcHoldSyncCnt[12]), .B0(n3101), .S(n3100), .CO(n3099));
Q_AD01HF U3458 ( .A0(ixcHoldSyncCnt[11]), .B0(n3103), .S(n3102), .CO(n3101));
Q_AD01HF U3459 ( .A0(ixcHoldSyncCnt[10]), .B0(n3105), .S(n3104), .CO(n3103));
Q_AD01HF U3460 ( .A0(ixcHoldSyncCnt[9]), .B0(n3107), .S(n3106), .CO(n3105));
Q_AD01HF U3461 ( .A0(ixcHoldSyncCnt[8]), .B0(n3109), .S(n3108), .CO(n3107));
Q_AD01HF U3462 ( .A0(ixcHoldSyncCnt[7]), .B0(n3111), .S(n3110), .CO(n3109));
Q_AD01HF U3463 ( .A0(ixcHoldSyncCnt[6]), .B0(n3113), .S(n3112), .CO(n3111));
Q_AD01HF U3464 ( .A0(ixcHoldSyncCnt[5]), .B0(n3115), .S(n3114), .CO(n3113));
Q_AD01HF U3465 ( .A0(ixcHoldSyncCnt[4]), .B0(n3117), .S(n3116), .CO(n3115));
Q_AD01HF U3466 ( .A0(ixcHoldSyncCnt[3]), .B0(n3119), .S(n3118), .CO(n3117));
Q_AD01HF U3467 ( .A0(ixcHoldSyncCnt[2]), .B0(n3121), .S(n3120), .CO(n3119));
Q_AD01HF U3468 ( .A0(ixcHoldSyncCnt[1]), .B0(ixcHoldSyncCnt[0]), .S(n3122), .CO(n3121));
Q_FDP0 ixcHoldClkR_REG  ( .CK(uClk), .D(ixcHoldClk), .Q(ixcHoldClkR), .QN(n2998));
Q_AD01HF U3470 ( .A0(bpCount[1]), .B0(bpCount[0]), .S(n3124), .CO(n3125));
Q_AD01HF U3471 ( .A0(bpCount[2]), .B0(n3125), .S(n3126), .CO(n3127));
Q_AD01HF U3472 ( .A0(bpCount[3]), .B0(n3127), .S(n3128), .CO(n3129));
Q_AD01HF U3473 ( .A0(bpCount[4]), .B0(n3129), .S(n3130), .CO(n3131));
Q_AD01HF U3474 ( .A0(bpCount[5]), .B0(n3131), .S(n3132), .CO(n3133));
Q_AD01HF U3475 ( .A0(bpCount[6]), .B0(n3133), .S(n3134), .CO(n3135));
Q_AD01HF U3476 ( .A0(bpCount[7]), .B0(n3135), .S(n3136), .CO(n3137));
Q_AD01HF U3477 ( .A0(bpCount[8]), .B0(n3137), .S(n3138), .CO(n3139));
Q_AD01HF U3478 ( .A0(bpCount[9]), .B0(n3139), .S(n3140), .CO(n3141));
Q_AD01HF U3479 ( .A0(bpCount[10]), .B0(n3141), .S(n3142), .CO(n3143));
Q_AD01HF U3480 ( .A0(bpCount[11]), .B0(n3143), .S(n3144), .CO(n3145));
Q_AD01HF U3481 ( .A0(bpCount[12]), .B0(n3145), .S(n3146), .CO(n3147));
Q_AD01HF U3482 ( .A0(bpCount[13]), .B0(n3147), .S(n3148), .CO(n3149));
Q_AD01HF U3483 ( .A0(bpCount[14]), .B0(n3149), .S(n3150), .CO(n3151));
Q_AD01HF U3484 ( .A0(bpCount[15]), .B0(n3151), .S(n3152), .CO(n3153));
Q_AD01HF U3485 ( .A0(bpCount[16]), .B0(n3153), .S(n3154), .CO(n3155));
Q_AD01HF U3486 ( .A0(bpCount[17]), .B0(n3155), .S(n3156), .CO(n3157));
Q_AD01HF U3487 ( .A0(bpCount[18]), .B0(n3157), .S(n3158), .CO(n3159));
Q_AD01HF U3488 ( .A0(bpCount[19]), .B0(n3159), .S(n3160), .CO(n3161));
Q_AD01HF U3489 ( .A0(bpCount[20]), .B0(n3161), .S(n3162), .CO(n3163));
Q_AD01HF U3490 ( .A0(bpCount[21]), .B0(n3163), .S(n3164), .CO(n3165));
Q_AD01HF U3491 ( .A0(bpCount[22]), .B0(n3165), .S(n3166), .CO(n3167));
Q_AD01HF U3492 ( .A0(bpCount[23]), .B0(n3167), .S(n3168), .CO(n3169));
Q_AD01HF U3493 ( .A0(bpCount[24]), .B0(n3169), .S(n3170), .CO(n3171));
Q_AD01HF U3494 ( .A0(bpCount[25]), .B0(n3171), .S(n3172), .CO(n3173));
Q_AD01HF U3495 ( .A0(bpCount[26]), .B0(n3173), .S(n3174), .CO(n3175));
Q_AD01HF U3496 ( .A0(bpCount[27]), .B0(n3175), .S(n3176), .CO(n3177));
Q_AD01HF U3497 ( .A0(bpCount[28]), .B0(n3177), .S(n3178), .CO(n3179));
Q_AD01HF U3498 ( .A0(bpCount[29]), .B0(n3179), .S(n3180), .CO(n3181));
Q_AD01HF U3499 ( .A0(bpCount[30]), .B0(n3181), .S(n3182), .CO(n3183));
Q_AD01HF U3500 ( .A0(bpCount[31]), .B0(n3183), .S(n3184), .CO(n3185));
Q_AD01HF U3501 ( .A0(bpCount[32]), .B0(n3185), .S(n3186), .CO(n3187));
Q_AD01HF U3502 ( .A0(bpCount[33]), .B0(n3187), .S(n3188), .CO(n3189));
Q_AD01HF U3503 ( .A0(bpCount[34]), .B0(n3189), .S(n3190), .CO(n3191));
Q_AD01HF U3504 ( .A0(bpCount[35]), .B0(n3191), .S(n3192), .CO(n3193));
Q_AD01HF U3505 ( .A0(bpCount[36]), .B0(n3193), .S(n3194), .CO(n3195));
Q_AD01HF U3506 ( .A0(bpCount[37]), .B0(n3195), .S(n3196), .CO(n3197));
Q_AD01HF U3507 ( .A0(bpCount[38]), .B0(n3197), .S(n3198), .CO(n3199));
Q_AD01HF U3508 ( .A0(bpCount[39]), .B0(n3199), .S(n3200), .CO(n3201));
Q_AD01HF U3509 ( .A0(bpCount[40]), .B0(n3201), .S(n3202), .CO(n3203));
Q_AD01HF U3510 ( .A0(bpCount[41]), .B0(n3203), .S(n3204), .CO(n3205));
Q_AD01HF U3511 ( .A0(bpCount[42]), .B0(n3205), .S(n3206), .CO(n3207));
Q_AD01HF U3512 ( .A0(bpCount[43]), .B0(n3207), .S(n3208), .CO(n3209));
Q_AD01HF U3513 ( .A0(bpCount[44]), .B0(n3209), .S(n3210), .CO(n3211));
Q_AD01HF U3514 ( .A0(bpCount[45]), .B0(n3211), .S(n3212), .CO(n3213));
Q_AD01HF U3515 ( .A0(bpCount[46]), .B0(n3213), .S(n3214), .CO(n3215));
Q_AD01HF U3516 ( .A0(bpCount[47]), .B0(n3215), .S(n3216), .CO(n3217));
Q_AD01HF U3517 ( .A0(bpCount[48]), .B0(n3217), .S(n3218), .CO(n3219));
Q_AD01HF U3518 ( .A0(bpCount[49]), .B0(n3219), .S(n3220), .CO(n3221));
Q_AD01HF U3519 ( .A0(bpCount[50]), .B0(n3221), .S(n3222), .CO(n3223));
Q_AD01HF U3520 ( .A0(bpCount[51]), .B0(n3223), .S(n3224), .CO(n3225));
Q_AD01HF U3521 ( .A0(bpCount[52]), .B0(n3225), .S(n3226), .CO(n3227));
Q_AD01HF U3522 ( .A0(bpCount[53]), .B0(n3227), .S(n3228), .CO(n3229));
Q_AD01HF U3523 ( .A0(bpCount[54]), .B0(n3229), .S(n3230), .CO(n3231));
Q_AD01HF U3524 ( .A0(bpCount[55]), .B0(n3231), .S(n3232), .CO(n3233));
Q_AD01HF U3525 ( .A0(bpCount[56]), .B0(n3233), .S(n3234), .CO(n3235));
Q_AD01HF U3526 ( .A0(bpCount[57]), .B0(n3235), .S(n3236), .CO(n3237));
Q_AD01HF U3527 ( .A0(bpCount[58]), .B0(n3237), .S(n3238), .CO(n3239));
Q_AD01HF U3528 ( .A0(bpCount[59]), .B0(n3239), .S(n3240), .CO(n3241));
Q_AD01HF U3529 ( .A0(bpCount[60]), .B0(n3241), .S(n3242), .CO(n3243));
Q_AD01HF U3530 ( .A0(bpCount[61]), .B0(n3243), .S(n3244), .CO(n3245));
Q_AD01HF U3531 ( .A0(bpCount[62]), .B0(n3245), .S(n3246), .CO(n3247));
Q_FDP0 \bpCount_REG[62] ( .CK(bClk), .D(n3246), .Q(bpCount[62]), .QN( ));
Q_FDP0 \bpCount_REG[61] ( .CK(bClk), .D(n3244), .Q(bpCount[61]), .QN( ));
Q_FDP0 \bpCount_REG[60] ( .CK(bClk), .D(n3242), .Q(bpCount[60]), .QN( ));
Q_FDP0 \bpCount_REG[59] ( .CK(bClk), .D(n3240), .Q(bpCount[59]), .QN( ));
Q_FDP0 \bpCount_REG[58] ( .CK(bClk), .D(n3238), .Q(bpCount[58]), .QN( ));
Q_FDP0 \bpCount_REG[57] ( .CK(bClk), .D(n3236), .Q(bpCount[57]), .QN( ));
Q_FDP0 \bpCount_REG[56] ( .CK(bClk), .D(n3234), .Q(bpCount[56]), .QN( ));
Q_FDP0 \bpCount_REG[55] ( .CK(bClk), .D(n3232), .Q(bpCount[55]), .QN( ));
Q_FDP0 \bpCount_REG[54] ( .CK(bClk), .D(n3230), .Q(bpCount[54]), .QN( ));
Q_FDP0 \bpCount_REG[53] ( .CK(bClk), .D(n3228), .Q(bpCount[53]), .QN( ));
Q_FDP0 \bpCount_REG[52] ( .CK(bClk), .D(n3226), .Q(bpCount[52]), .QN( ));
Q_FDP0 \bpCount_REG[51] ( .CK(bClk), .D(n3224), .Q(bpCount[51]), .QN( ));
Q_FDP0 \bpCount_REG[50] ( .CK(bClk), .D(n3222), .Q(bpCount[50]), .QN( ));
Q_FDP0 \bpCount_REG[49] ( .CK(bClk), .D(n3220), .Q(bpCount[49]), .QN( ));
Q_FDP0 \bpCount_REG[48] ( .CK(bClk), .D(n3218), .Q(bpCount[48]), .QN( ));
Q_FDP0 \bpCount_REG[47] ( .CK(bClk), .D(n3216), .Q(bpCount[47]), .QN( ));
Q_FDP0 \bpCount_REG[46] ( .CK(bClk), .D(n3214), .Q(bpCount[46]), .QN( ));
Q_FDP0 \bpCount_REG[45] ( .CK(bClk), .D(n3212), .Q(bpCount[45]), .QN( ));
Q_FDP0 \bpCount_REG[44] ( .CK(bClk), .D(n3210), .Q(bpCount[44]), .QN( ));
Q_FDP0 \bpCount_REG[43] ( .CK(bClk), .D(n3208), .Q(bpCount[43]), .QN( ));
Q_FDP0 \bpCount_REG[42] ( .CK(bClk), .D(n3206), .Q(bpCount[42]), .QN( ));
Q_FDP0 \bpCount_REG[41] ( .CK(bClk), .D(n3204), .Q(bpCount[41]), .QN( ));
Q_FDP0 \bpCount_REG[40] ( .CK(bClk), .D(n3202), .Q(bpCount[40]), .QN( ));
Q_FDP0 \bpCount_REG[39] ( .CK(bClk), .D(n3200), .Q(bpCount[39]), .QN( ));
Q_FDP0 \bpCount_REG[38] ( .CK(bClk), .D(n3198), .Q(bpCount[38]), .QN( ));
Q_FDP0 \bpCount_REG[37] ( .CK(bClk), .D(n3196), .Q(bpCount[37]), .QN( ));
Q_FDP0 \bpCount_REG[36] ( .CK(bClk), .D(n3194), .Q(bpCount[36]), .QN( ));
Q_FDP0 \bpCount_REG[35] ( .CK(bClk), .D(n3192), .Q(bpCount[35]), .QN( ));
Q_FDP0 \bpCount_REG[34] ( .CK(bClk), .D(n3190), .Q(bpCount[34]), .QN( ));
Q_FDP0 \bpCount_REG[33] ( .CK(bClk), .D(n3188), .Q(bpCount[33]), .QN( ));
Q_FDP0 \bpCount_REG[32] ( .CK(bClk), .D(n3186), .Q(bpCount[32]), .QN( ));
Q_FDP0 \bpCount_REG[31] ( .CK(bClk), .D(n3184), .Q(bpCount[31]), .QN( ));
Q_FDP0 \bpCount_REG[30] ( .CK(bClk), .D(n3182), .Q(bpCount[30]), .QN( ));
Q_FDP0 \bpCount_REG[29] ( .CK(bClk), .D(n3180), .Q(bpCount[29]), .QN( ));
Q_FDP0 \bpCount_REG[28] ( .CK(bClk), .D(n3178), .Q(bpCount[28]), .QN( ));
Q_FDP0 \bpCount_REG[27] ( .CK(bClk), .D(n3176), .Q(bpCount[27]), .QN( ));
Q_FDP0 \bpCount_REG[26] ( .CK(bClk), .D(n3174), .Q(bpCount[26]), .QN( ));
Q_FDP0 \bpCount_REG[25] ( .CK(bClk), .D(n3172), .Q(bpCount[25]), .QN( ));
Q_FDP0 \bpCount_REG[24] ( .CK(bClk), .D(n3170), .Q(bpCount[24]), .QN( ));
Q_FDP0 \bpCount_REG[23] ( .CK(bClk), .D(n3168), .Q(bpCount[23]), .QN( ));
Q_FDP0 \bpCount_REG[22] ( .CK(bClk), .D(n3166), .Q(bpCount[22]), .QN( ));
Q_FDP0 \bpCount_REG[21] ( .CK(bClk), .D(n3164), .Q(bpCount[21]), .QN( ));
Q_FDP0 \bpCount_REG[20] ( .CK(bClk), .D(n3162), .Q(bpCount[20]), .QN( ));
Q_FDP0 \bpCount_REG[19] ( .CK(bClk), .D(n3160), .Q(bpCount[19]), .QN( ));
Q_FDP0 \bpCount_REG[18] ( .CK(bClk), .D(n3158), .Q(bpCount[18]), .QN( ));
Q_FDP0 \bpCount_REG[17] ( .CK(bClk), .D(n3156), .Q(bpCount[17]), .QN( ));
Q_FDP0 \bpCount_REG[16] ( .CK(bClk), .D(n3154), .Q(bpCount[16]), .QN( ));
Q_FDP0 \bpCount_REG[15] ( .CK(bClk), .D(n3152), .Q(bpCount[15]), .QN( ));
Q_FDP0 \bpCount_REG[14] ( .CK(bClk), .D(n3150), .Q(bpCount[14]), .QN( ));
Q_FDP0 \bpCount_REG[13] ( .CK(bClk), .D(n3148), .Q(bpCount[13]), .QN( ));
Q_FDP0 \bpCount_REG[12] ( .CK(bClk), .D(n3146), .Q(bpCount[12]), .QN( ));
Q_FDP0 \bpCount_REG[11] ( .CK(bClk), .D(n3144), .Q(bpCount[11]), .QN( ));
Q_FDP0 \bpCount_REG[10] ( .CK(bClk), .D(n3142), .Q(bpCount[10]), .QN( ));
Q_FDP0 \bpCount_REG[9] ( .CK(bClk), .D(n3140), .Q(bpCount[9]), .QN( ));
Q_FDP0 \bpCount_REG[8] ( .CK(bClk), .D(n3138), .Q(bpCount[8]), .QN( ));
Q_FDP0 \bpCount_REG[7] ( .CK(bClk), .D(n3136), .Q(bpCount[7]), .QN( ));
Q_FDP0 \bpCount_REG[6] ( .CK(bClk), .D(n3134), .Q(bpCount[6]), .QN( ));
Q_FDP0 \bpCount_REG[5] ( .CK(bClk), .D(n3132), .Q(bpCount[5]), .QN( ));
Q_FDP0 \bpCount_REG[4] ( .CK(bClk), .D(n3130), .Q(bpCount[4]), .QN( ));
Q_FDP0 \bpCount_REG[3] ( .CK(bClk), .D(n3128), .Q(bpCount[3]), .QN( ));
Q_FDP0 \bpCount_REG[2] ( .CK(bClk), .D(n3126), .Q(bpCount[2]), .QN( ));
Q_FDP0 \bpCount_REG[1] ( .CK(bClk), .D(n3124), .Q(bpCount[1]), .QN( ));
Q_FDP0 \bpCount_REG[0] ( .CK(bClk), .D(n3123), .Q(bpCount[0]), .QN(n3123));
Q_NR02 U3595 ( .A0(bpSt[1]), .A1(bpSt[0]), .Z(n3248));
Q_MX02 U3596 ( .S(n3248), .A0(n3249), .A1(n3251), .Z(lastDelta));
Q_NR03 U3597 ( .A0(n3248), .A1(bpHalt), .A2(bClkHoldD), .Z(bpOn));
Q_AN02 U3598 ( .A0(n3250), .A1(n2121), .Z(n3249));
Q_INV U3599 ( .A(sampleXpV), .Z(n3250));
Q_ND02 U3600 ( .A0(sampleXpV), .A1(mpOn), .Z(n3251));
Q_OR02 U3601 ( .A0(bpWait), .A1(sampleXpChg), .Z(sampleXpV));
Q_FDP0 SFIFOLock2_REG  ( .CK(uClk), .D(SFIFOLock), .Q(SFIFOLock2), .QN( ));
Q_AO21 U3603 ( .A0(callEmuEv), .A1(tbcPOState[0]), .B0(n3258), .Z(n3253));
Q_AO21 U3604 ( .A0(tbcPOd), .A1(tbcPORdy), .B0(tbcPOState[0]), .Z(n3257));
Q_OR02 U3605 ( .A0(tbcPOState[1]), .A1(n3253), .Z(n3260));
Q_INV U3606 ( .A(n3260), .Z(n3254));
Q_OR02 U3607 ( .A0(forceAbort), .A1(n3254), .Z(tbcPO));
Q_INV U3608 ( .A(tbcPOd), .Z(n3255));
Q_OR02 U3609 ( .A0(tbcPOState[0]), .A1(n3255), .Z(n3256));
Q_INV U3610 ( .A(n3257), .Z(n3258));
Q_MX02 U3611 ( .S(tbcPOState[1]), .A0(n3258), .A1(n3256), .Z(n3259));
Q_OR02 U3612 ( .A0(forceAbort), .A1(n3259), .Z(n3252));
Q_OR02 U3613 ( .A0(forceAbort), .A1(n3260), .Z(n3261));
Q_INV U3614 ( .A(n3261), .Z(tbcPOStateN[0]));
Q_XOR2 U3615 ( .A0(n3261), .A1(n3252), .Z(tbcPOStateN[1]));
Q_AN03 U3616 ( .A0(tbcPODly[12]), .A1(tbcPODly[11]), .A2(tbcPODly[10]), .Z(n3262));
Q_AN03 U3617 ( .A0(tbcPODly[9]), .A1(tbcPODly[8]), .A2(tbcPODly[7]), .Z(n3263));
Q_AN03 U3618 ( .A0(tbcPODly[6]), .A1(tbcPODly[5]), .A2(tbcPODly[4]), .Z(n3264));
Q_AN03 U3619 ( .A0(tbcPODly[3]), .A1(tbcPODly[2]), .A2(tbcPODly[1]), .Z(n3265));
Q_AN03 U3620 ( .A0(tbcPODly[0]), .A1(n3262), .A2(n3263), .Z(n3266));
Q_AN03 U3621 ( .A0(n3264), .A1(n3265), .A2(n3266), .Z(n3267));
Q_OR02 U3622 ( .A0(n3267), .A1(n2253), .Z(n3268));
Q_INV U3623 ( .A(gfifoWait), .Z(n3269));
Q_NR03 U3624 ( .A0(osfWait), .A1(asyncBusy), .A2(ptxBusy), .Z(n3270));
Q_AN03 U3625 ( .A0(n3269), .A1(n3270), .A2(n3268), .Z(tbcPORdy));
Q_INV U3626 ( .A(stop3), .Z(n3278));
Q_AN02 U3627 ( .A0(n3285), .A1(n3278), .Z(n3271));
Q_AN02 U3628 ( .A0(n3285), .A1(stop3), .Z(n3272));
Q_INV U3629 ( .A(stopT), .Z(n3279));
Q_AN02 U3630 ( .A0(n3285), .A1(n3279), .Z(n3273));
Q_AN02 U3631 ( .A0(n3285), .A1(stopT), .Z(n3274));
Q_MX02 U3632 ( .S(n3271), .A0(n3272), .A1(stop3POd), .Z(stop3PO));
Q_MX02 U3633 ( .S(oneStepPIi), .A0(ixcSimTime[63]), .A1(evfCount[63]), .Z(remStepPO[63]));
Q_MX02 U3634 ( .S(oneStepPIi), .A0(ixcSimTime[62]), .A1(evfCount[62]), .Z(remStepPO[62]));
Q_MX02 U3635 ( .S(oneStepPIi), .A0(ixcSimTime[61]), .A1(evfCount[61]), .Z(remStepPO[61]));
Q_MX02 U3636 ( .S(oneStepPIi), .A0(ixcSimTime[60]), .A1(evfCount[60]), .Z(remStepPO[60]));
Q_MX02 U3637 ( .S(oneStepPIi), .A0(ixcSimTime[59]), .A1(evfCount[59]), .Z(remStepPO[59]));
Q_MX02 U3638 ( .S(oneStepPIi), .A0(ixcSimTime[58]), .A1(evfCount[58]), .Z(remStepPO[58]));
Q_MX02 U3639 ( .S(oneStepPIi), .A0(ixcSimTime[57]), .A1(evfCount[57]), .Z(remStepPO[57]));
Q_MX02 U3640 ( .S(oneStepPIi), .A0(ixcSimTime[56]), .A1(evfCount[56]), .Z(remStepPO[56]));
Q_MX02 U3641 ( .S(oneStepPIi), .A0(ixcSimTime[55]), .A1(evfCount[55]), .Z(remStepPO[55]));
Q_MX02 U3642 ( .S(oneStepPIi), .A0(ixcSimTime[54]), .A1(evfCount[54]), .Z(remStepPO[54]));
Q_MX02 U3643 ( .S(oneStepPIi), .A0(ixcSimTime[53]), .A1(evfCount[53]), .Z(remStepPO[53]));
Q_MX02 U3644 ( .S(oneStepPIi), .A0(ixcSimTime[52]), .A1(evfCount[52]), .Z(remStepPO[52]));
Q_MX02 U3645 ( .S(oneStepPIi), .A0(ixcSimTime[51]), .A1(evfCount[51]), .Z(remStepPO[51]));
Q_MX02 U3646 ( .S(oneStepPIi), .A0(ixcSimTime[50]), .A1(evfCount[50]), .Z(remStepPO[50]));
Q_MX02 U3647 ( .S(oneStepPIi), .A0(ixcSimTime[49]), .A1(evfCount[49]), .Z(remStepPO[49]));
Q_MX02 U3648 ( .S(oneStepPIi), .A0(ixcSimTime[48]), .A1(evfCount[48]), .Z(remStepPO[48]));
Q_MX02 U3649 ( .S(oneStepPIi), .A0(ixcSimTime[47]), .A1(evfCount[47]), .Z(remStepPO[47]));
Q_MX02 U3650 ( .S(oneStepPIi), .A0(ixcSimTime[46]), .A1(evfCount[46]), .Z(remStepPO[46]));
Q_MX02 U3651 ( .S(oneStepPIi), .A0(ixcSimTime[45]), .A1(evfCount[45]), .Z(remStepPO[45]));
Q_MX02 U3652 ( .S(oneStepPIi), .A0(ixcSimTime[44]), .A1(evfCount[44]), .Z(remStepPO[44]));
Q_MX02 U3653 ( .S(oneStepPIi), .A0(ixcSimTime[43]), .A1(evfCount[43]), .Z(remStepPO[43]));
Q_MX02 U3654 ( .S(oneStepPIi), .A0(ixcSimTime[42]), .A1(evfCount[42]), .Z(remStepPO[42]));
Q_MX02 U3655 ( .S(oneStepPIi), .A0(ixcSimTime[41]), .A1(evfCount[41]), .Z(remStepPO[41]));
Q_MX02 U3656 ( .S(oneStepPIi), .A0(ixcSimTime[40]), .A1(evfCount[40]), .Z(remStepPO[40]));
Q_MX02 U3657 ( .S(oneStepPIi), .A0(ixcSimTime[39]), .A1(evfCount[39]), .Z(remStepPO[39]));
Q_MX02 U3658 ( .S(oneStepPIi), .A0(ixcSimTime[38]), .A1(evfCount[38]), .Z(remStepPO[38]));
Q_MX02 U3659 ( .S(oneStepPIi), .A0(ixcSimTime[37]), .A1(evfCount[37]), .Z(remStepPO[37]));
Q_MX02 U3660 ( .S(oneStepPIi), .A0(ixcSimTime[36]), .A1(evfCount[36]), .Z(remStepPO[36]));
Q_MX02 U3661 ( .S(oneStepPIi), .A0(ixcSimTime[35]), .A1(evfCount[35]), .Z(remStepPO[35]));
Q_MX02 U3662 ( .S(oneStepPIi), .A0(ixcSimTime[34]), .A1(evfCount[34]), .Z(remStepPO[34]));
Q_MX02 U3663 ( .S(oneStepPIi), .A0(ixcSimTime[33]), .A1(evfCount[33]), .Z(remStepPO[33]));
Q_MX02 U3664 ( .S(oneStepPIi), .A0(ixcSimTime[32]), .A1(evfCount[32]), .Z(remStepPO[32]));
Q_MX02 U3665 ( .S(oneStepPIi), .A0(ixcSimTime[31]), .A1(evfCount[31]), .Z(remStepPO[31]));
Q_MX02 U3666 ( .S(oneStepPIi), .A0(ixcSimTime[30]), .A1(evfCount[30]), .Z(remStepPO[30]));
Q_MX02 U3667 ( .S(oneStepPIi), .A0(ixcSimTime[29]), .A1(evfCount[29]), .Z(remStepPO[29]));
Q_MX02 U3668 ( .S(oneStepPIi), .A0(ixcSimTime[28]), .A1(evfCount[28]), .Z(remStepPO[28]));
Q_MX02 U3669 ( .S(oneStepPIi), .A0(ixcSimTime[27]), .A1(evfCount[27]), .Z(remStepPO[27]));
Q_MX02 U3670 ( .S(oneStepPIi), .A0(ixcSimTime[26]), .A1(evfCount[26]), .Z(remStepPO[26]));
Q_MX02 U3671 ( .S(oneStepPIi), .A0(ixcSimTime[25]), .A1(evfCount[25]), .Z(remStepPO[25]));
Q_MX02 U3672 ( .S(oneStepPIi), .A0(ixcSimTime[24]), .A1(evfCount[24]), .Z(remStepPO[24]));
Q_MX02 U3673 ( .S(oneStepPIi), .A0(ixcSimTime[23]), .A1(evfCount[23]), .Z(remStepPO[23]));
Q_MX02 U3674 ( .S(oneStepPIi), .A0(ixcSimTime[22]), .A1(evfCount[22]), .Z(remStepPO[22]));
Q_MX02 U3675 ( .S(oneStepPIi), .A0(ixcSimTime[21]), .A1(evfCount[21]), .Z(remStepPO[21]));
Q_MX02 U3676 ( .S(oneStepPIi), .A0(ixcSimTime[20]), .A1(evfCount[20]), .Z(remStepPO[20]));
Q_MX02 U3677 ( .S(oneStepPIi), .A0(ixcSimTime[19]), .A1(evfCount[19]), .Z(remStepPO[19]));
Q_MX02 U3678 ( .S(oneStepPIi), .A0(ixcSimTime[18]), .A1(evfCount[18]), .Z(remStepPO[18]));
Q_MX02 U3679 ( .S(oneStepPIi), .A0(ixcSimTime[17]), .A1(evfCount[17]), .Z(remStepPO[17]));
Q_MX02 U3680 ( .S(oneStepPIi), .A0(ixcSimTime[16]), .A1(evfCount[16]), .Z(remStepPO[16]));
Q_MX02 U3681 ( .S(oneStepPIi), .A0(ixcSimTime[15]), .A1(evfCount[15]), .Z(remStepPO[15]));
Q_MX02 U3682 ( .S(oneStepPIi), .A0(ixcSimTime[14]), .A1(evfCount[14]), .Z(remStepPO[14]));
Q_MX02 U3683 ( .S(oneStepPIi), .A0(ixcSimTime[13]), .A1(evfCount[13]), .Z(remStepPO[13]));
Q_MX02 U3684 ( .S(oneStepPIi), .A0(ixcSimTime[12]), .A1(evfCount[12]), .Z(remStepPO[12]));
Q_MX02 U3685 ( .S(oneStepPIi), .A0(ixcSimTime[11]), .A1(evfCount[11]), .Z(remStepPO[11]));
Q_MX02 U3686 ( .S(oneStepPIi), .A0(ixcSimTime[10]), .A1(evfCount[10]), .Z(remStepPO[10]));
Q_MX02 U3687 ( .S(oneStepPIi), .A0(ixcSimTime[9]), .A1(evfCount[9]), .Z(remStepPO[9]));
Q_MX02 U3688 ( .S(oneStepPIi), .A0(ixcSimTime[8]), .A1(evfCount[8]), .Z(remStepPO[8]));
Q_MX02 U3689 ( .S(oneStepPIi), .A0(ixcSimTime[7]), .A1(evfCount[7]), .Z(remStepPO[7]));
Q_MX02 U3690 ( .S(oneStepPIi), .A0(ixcSimTime[6]), .A1(evfCount[6]), .Z(remStepPO[6]));
Q_MX02 U3691 ( .S(oneStepPIi), .A0(ixcSimTime[5]), .A1(evfCount[5]), .Z(remStepPO[5]));
Q_MX02 U3692 ( .S(oneStepPIi), .A0(ixcSimTime[4]), .A1(evfCount[4]), .Z(remStepPO[4]));
Q_MX02 U3693 ( .S(oneStepPIi), .A0(ixcSimTime[3]), .A1(evfCount[3]), .Z(remStepPO[3]));
Q_MX02 U3694 ( .S(oneStepPIi), .A0(ixcSimTime[2]), .A1(evfCount[2]), .Z(remStepPO[2]));
Q_MX02 U3695 ( .S(oneStepPIi), .A0(ixcSimTime[1]), .A1(evfCount[1]), .Z(remStepPO[1]));
Q_MX02 U3696 ( .S(oneStepPIi), .A0(ixcSimTime[0]), .A1(evfCount[0]), .Z(remStepPO[0]));
Q_MX02 U3697 ( .S(n3273), .A0(n3274), .A1(stopTLd), .Z(stopTL));
Q_MX02 U3698 ( .S(n3275), .A0(stop4POd), .A1(stop4R), .Z(stop4PO));
Q_MX02 U3699 ( .S(n3276), .A0(stop2POd), .A1(stop2R), .Z(stop2PO));
Q_MX02 U3700 ( .S(n3277), .A0(stop1POd), .A1(stop1R), .Z(stop1PO));
Q_OR02 U3701 ( .A0(callEmuPre), .A1(stop4R), .Z(n3275));
Q_OR02 U3702 ( .A0(callEmuPre), .A1(stop2R), .Z(n3276));
Q_OR02 U3703 ( .A0(callEmuPre), .A1(stop1R), .Z(n3277));
Q_OR02 U3704 ( .A0(callEmuPre), .A1(evalOnC), .Z(n3280));
Q_FDP0 eventOnR_REG  ( .CK(uClk), .D(n3280), .Q(eventOnR), .QN( ));
Q_OR03 U3706 ( .A0(callEmuPre), .A1(evalOnC), .A2(hotSwapOnPI), .Z(n3281));
Q_FDP0 eventOnRI_REG  ( .CK(uClk), .D(n3281), .Q(eventOnRI), .QN( ));
Q_AO21 U3708 ( .A0(n2616), .A1(tbcPOReg), .B0(GFLock1), .Z(GFLock2R));
Q_OA21 U3709 ( .A0(GFLock2R), .A1(xcReplayOnReg), .B0(n2252), .Z(GFLock2));
Q_FDP0 tbcPOReg_REG  ( .CK(uClk), .D(mioPOW_2[1]), .Q(tbcPOReg), .QN( ));
Q_FDP0 xcReplayOnReg_REG  ( .CK(uClk), .D(xcReplayOn), .Q(xcReplayOnReg), .QN( ));
Q_OA21 U3712 ( .A0(gfifoOff), .A1(hotSwapOnPI), .B0(n2252), .Z(n3282));
Q_FDP0 GFLock1_REG  ( .CK(uClk), .D(n3282), .Q(GFLock1), .QN( ));
Q_INV U3714 ( .A(gfifoAsyncOff), .Z(n3283));
Q_AN02 U3715 ( .A0(GFGBfull), .A1(n3283), .Z(n3284));
Q_FDP0 GFGBfullBw_REG  ( .CK(uClk), .D(n3284), .Q(GFGBfullBw), .QN( ));
Q_AN02 U3717 ( .A0(callEmuPreD), .A1(callEmuPre), .Z(callEmu));
Q_NR02 U3718 ( .A0(callEmuEv), .A1(callEmuWait), .Z(n3286));
Q_OR02 U3719 ( .A0(n3286), .A1(callEmuWaitC), .Z(n3285));
Q_INV U3720 ( .A(n3285), .Z(callEmuPre));
Q_INV U3721 ( .A(n3286), .Z(n3287));
Q_AN02 U3722 ( .A0(callEmuWaitC), .A1(n3287), .Z(callEmuWaitN));
Q_OR02 U3723 ( .A0(hotSwapOnPI), .A1(callEmu), .Z(n3288));
Q_FDP0 callEmuR_REG  ( .CK(uClk), .D(callEmuPIi), .Q(callEmuR), .QN( ));
Q_OR02 U3725 ( .A0(oneStepPIi), .A1(n2189), .Z(n3292));
Q_MX02 U3726 ( .S(callEmuEv), .A0(simTimeOn), .A1(n3292), .Z(n3293));
Q_OR03 U3727 ( .A0(hwClkDbgTime), .A1(lockTraceOn), .A2(n3293), .Z(n3289));
Q_OR03 U3728 ( .A0(lockTraceOn), .A1(callEmuEv), .A2(hwClkDbgTime), .Z(n3294));
Q_OR02 U3729 ( .A0(n2616), .A1(oneStepPIi), .Z(n3297));
Q_AO21 U3730 ( .A0(n3295), .A1(n3297), .B0(hwClkDbgTime), .Z(n3296));
Q_INV U3731 ( .A(n3296), .Z(n3290));
Q_NR02 U3732 ( .A0(lockTraceOn), .A1(n3297), .Z(n3298));
Q_OR02 U3733 ( .A0(hwClkDbgTime), .A1(n3298), .Z(n3291));
Q_LDP0 \simTime_REG[0] ( .G(n3289), .D(n3425), .Q(simTime[0]), .QN( ));
Q_LDP0 \simTime_REG[1] ( .G(n3289), .D(n3423), .Q(simTime[1]), .QN( ));
Q_LDP0 \simTime_REG[2] ( .G(n3289), .D(n3421), .Q(simTime[2]), .QN(n3569));
Q_LDP0 \simTime_REG[3] ( .G(n3289), .D(n3419), .Q(simTime[3]), .QN( ));
Q_LDP0 \simTime_REG[4] ( .G(n3289), .D(n3417), .Q(simTime[4]), .QN( ));
Q_LDP0 \simTime_REG[5] ( .G(n3289), .D(n3415), .Q(simTime[5]), .QN( ));
Q_LDP0 \simTime_REG[6] ( .G(n3289), .D(n3413), .Q(simTime[6]), .QN( ));
Q_LDP0 \simTime_REG[7] ( .G(n3289), .D(n3411), .Q(simTime[7]), .QN( ));
Q_LDP0 \simTime_REG[8] ( .G(n3289), .D(n3409), .Q(simTime[8]), .QN( ));
Q_LDP0 \simTime_REG[9] ( .G(n3289), .D(n3407), .Q(simTime[9]), .QN( ));
Q_LDP0 \simTime_REG[10] ( .G(n3289), .D(n3405), .Q(simTime[10]), .QN( ));
Q_LDP0 \simTime_REG[11] ( .G(n3289), .D(n3403), .Q(simTime[11]), .QN( ));
Q_LDP0 \simTime_REG[12] ( .G(n3289), .D(n3401), .Q(simTime[12]), .QN( ));
Q_LDP0 \simTime_REG[13] ( .G(n3289), .D(n3399), .Q(simTime[13]), .QN( ));
Q_LDP0 \simTime_REG[14] ( .G(n3289), .D(n3397), .Q(simTime[14]), .QN( ));
Q_LDP0 \simTime_REG[15] ( .G(n3289), .D(n3395), .Q(simTime[15]), .QN( ));
Q_LDP0 \simTime_REG[16] ( .G(n3289), .D(n3393), .Q(simTime[16]), .QN( ));
Q_LDP0 \simTime_REG[17] ( .G(n3289), .D(n3391), .Q(simTime[17]), .QN( ));
Q_LDP0 \simTime_REG[18] ( .G(n3289), .D(n3389), .Q(simTime[18]), .QN( ));
Q_LDP0 \simTime_REG[19] ( .G(n3289), .D(n3387), .Q(simTime[19]), .QN( ));
Q_LDP0 \simTime_REG[20] ( .G(n3289), .D(n3385), .Q(simTime[20]), .QN( ));
Q_LDP0 \simTime_REG[21] ( .G(n3289), .D(n3383), .Q(simTime[21]), .QN( ));
Q_LDP0 \simTime_REG[22] ( .G(n3289), .D(n3381), .Q(simTime[22]), .QN( ));
Q_LDP0 \simTime_REG[23] ( .G(n3289), .D(n3379), .Q(simTime[23]), .QN( ));
Q_LDP0 \simTime_REG[24] ( .G(n3289), .D(n3377), .Q(simTime[24]), .QN( ));
Q_LDP0 \simTime_REG[25] ( .G(n3289), .D(n3375), .Q(simTime[25]), .QN( ));
Q_LDP0 \simTime_REG[26] ( .G(n3289), .D(n3373), .Q(simTime[26]), .QN( ));
Q_LDP0 \simTime_REG[27] ( .G(n3289), .D(n3371), .Q(simTime[27]), .QN( ));
Q_LDP0 \simTime_REG[28] ( .G(n3289), .D(n3369), .Q(simTime[28]), .QN( ));
Q_LDP0 \simTime_REG[29] ( .G(n3289), .D(n3367), .Q(simTime[29]), .QN( ));
Q_LDP0 \simTime_REG[30] ( .G(n3289), .D(n3365), .Q(simTime[30]), .QN( ));
Q_LDP0 \simTime_REG[31] ( .G(n3289), .D(n3363), .Q(simTime[31]), .QN( ));
Q_LDP0 \simTime_REG[32] ( .G(n3289), .D(n3361), .Q(simTime[32]), .QN( ));
Q_LDP0 \simTime_REG[33] ( .G(n3289), .D(n3359), .Q(simTime[33]), .QN( ));
Q_LDP0 \simTime_REG[34] ( .G(n3289), .D(n3357), .Q(simTime[34]), .QN( ));
Q_LDP0 \simTime_REG[35] ( .G(n3289), .D(n3355), .Q(simTime[35]), .QN( ));
Q_LDP0 \simTime_REG[36] ( .G(n3289), .D(n3353), .Q(simTime[36]), .QN( ));
Q_LDP0 \simTime_REG[37] ( .G(n3289), .D(n3351), .Q(simTime[37]), .QN( ));
Q_LDP0 \simTime_REG[38] ( .G(n3289), .D(n3349), .Q(simTime[38]), .QN( ));
Q_LDP0 \simTime_REG[39] ( .G(n3289), .D(n3347), .Q(simTime[39]), .QN( ));
Q_LDP0 \simTime_REG[40] ( .G(n3289), .D(n3345), .Q(simTime[40]), .QN( ));
Q_LDP0 \simTime_REG[41] ( .G(n3289), .D(n3343), .Q(simTime[41]), .QN( ));
Q_LDP0 \simTime_REG[42] ( .G(n3289), .D(n3341), .Q(simTime[42]), .QN( ));
Q_LDP0 \simTime_REG[43] ( .G(n3289), .D(n3339), .Q(simTime[43]), .QN( ));
Q_LDP0 \simTime_REG[44] ( .G(n3289), .D(n3337), .Q(simTime[44]), .QN( ));
Q_LDP0 \simTime_REG[45] ( .G(n3289), .D(n3335), .Q(simTime[45]), .QN( ));
Q_LDP0 \simTime_REG[46] ( .G(n3289), .D(n3333), .Q(simTime[46]), .QN( ));
Q_LDP0 \simTime_REG[47] ( .G(n3289), .D(n3331), .Q(simTime[47]), .QN( ));
Q_LDP0 \simTime_REG[48] ( .G(n3289), .D(n3329), .Q(simTime[48]), .QN( ));
Q_LDP0 \simTime_REG[49] ( .G(n3289), .D(n3327), .Q(simTime[49]), .QN( ));
Q_LDP0 \simTime_REG[50] ( .G(n3289), .D(n3325), .Q(simTime[50]), .QN( ));
Q_LDP0 \simTime_REG[51] ( .G(n3289), .D(n3323), .Q(simTime[51]), .QN( ));
Q_LDP0 \simTime_REG[52] ( .G(n3289), .D(n3321), .Q(simTime[52]), .QN( ));
Q_LDP0 \simTime_REG[53] ( .G(n3289), .D(n3319), .Q(simTime[53]), .QN( ));
Q_LDP0 \simTime_REG[54] ( .G(n3289), .D(n3317), .Q(simTime[54]), .QN( ));
Q_LDP0 \simTime_REG[55] ( .G(n3289), .D(n3315), .Q(simTime[55]), .QN( ));
Q_LDP0 \simTime_REG[56] ( .G(n3289), .D(n3313), .Q(simTime[56]), .QN( ));
Q_LDP0 \simTime_REG[57] ( .G(n3289), .D(n3311), .Q(simTime[57]), .QN( ));
Q_LDP0 \simTime_REG[58] ( .G(n3289), .D(n3309), .Q(simTime[58]), .QN( ));
Q_LDP0 \simTime_REG[59] ( .G(n3289), .D(n3307), .Q(simTime[59]), .QN( ));
Q_LDP0 \simTime_REG[60] ( .G(n3289), .D(n3305), .Q(simTime[60]), .QN( ));
Q_LDP0 \simTime_REG[61] ( .G(n3289), .D(n3303), .Q(simTime[61]), .QN( ));
Q_LDP0 \simTime_REG[62] ( .G(n3289), .D(n3301), .Q(simTime[62]), .QN( ));
Q_LDP0 \simTime_REG[63] ( .G(n3289), .D(n3299), .Q(simTime[63]), .QN( ));
Q_MX02 U3798 ( .S(n3294), .A0(ixcSimTime[63]), .A1(n3300), .Z(n3299));
Q_MX04 U3799 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[63]), .A1(hwSimTime[63]), .A2(lockTraceTime[63]), .A3(nextDutTimeS[63]), .Z(n3300));
Q_MX02 U3800 ( .S(n3294), .A0(ixcSimTime[62]), .A1(n3302), .Z(n3301));
Q_MX04 U3801 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[62]), .A1(hwSimTime[62]), .A2(lockTraceTime[62]), .A3(nextDutTimeS[62]), .Z(n3302));
Q_MX02 U3802 ( .S(n3294), .A0(ixcSimTime[61]), .A1(n3304), .Z(n3303));
Q_MX04 U3803 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[61]), .A1(hwSimTime[61]), .A2(lockTraceTime[61]), .A3(nextDutTimeS[61]), .Z(n3304));
Q_MX02 U3804 ( .S(n3294), .A0(ixcSimTime[60]), .A1(n3306), .Z(n3305));
Q_MX04 U3805 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[60]), .A1(hwSimTime[60]), .A2(lockTraceTime[60]), .A3(nextDutTimeS[60]), .Z(n3306));
Q_MX02 U3806 ( .S(n3294), .A0(ixcSimTime[59]), .A1(n3308), .Z(n3307));
Q_MX04 U3807 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[59]), .A1(hwSimTime[59]), .A2(lockTraceTime[59]), .A3(nextDutTimeS[59]), .Z(n3308));
Q_MX02 U3808 ( .S(n3294), .A0(ixcSimTime[58]), .A1(n3310), .Z(n3309));
Q_MX04 U3809 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[58]), .A1(hwSimTime[58]), .A2(lockTraceTime[58]), .A3(nextDutTimeS[58]), .Z(n3310));
Q_MX02 U3810 ( .S(n3294), .A0(ixcSimTime[57]), .A1(n3312), .Z(n3311));
Q_MX04 U3811 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[57]), .A1(hwSimTime[57]), .A2(lockTraceTime[57]), .A3(nextDutTimeS[57]), .Z(n3312));
Q_MX02 U3812 ( .S(n3294), .A0(ixcSimTime[56]), .A1(n3314), .Z(n3313));
Q_MX04 U3813 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[56]), .A1(hwSimTime[56]), .A2(lockTraceTime[56]), .A3(nextDutTimeS[56]), .Z(n3314));
Q_MX02 U3814 ( .S(n3294), .A0(ixcSimTime[55]), .A1(n3316), .Z(n3315));
Q_MX04 U3815 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[55]), .A1(hwSimTime[55]), .A2(lockTraceTime[55]), .A3(nextDutTimeS[55]), .Z(n3316));
Q_MX02 U3816 ( .S(n3294), .A0(ixcSimTime[54]), .A1(n3318), .Z(n3317));
Q_MX04 U3817 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[54]), .A1(hwSimTime[54]), .A2(lockTraceTime[54]), .A3(nextDutTimeS[54]), .Z(n3318));
Q_MX02 U3818 ( .S(n3294), .A0(ixcSimTime[53]), .A1(n3320), .Z(n3319));
Q_MX04 U3819 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[53]), .A1(hwSimTime[53]), .A2(lockTraceTime[53]), .A3(nextDutTimeS[53]), .Z(n3320));
Q_MX02 U3820 ( .S(n3294), .A0(ixcSimTime[52]), .A1(n3322), .Z(n3321));
Q_MX04 U3821 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[52]), .A1(hwSimTime[52]), .A2(lockTraceTime[52]), .A3(nextDutTimeS[52]), .Z(n3322));
Q_MX02 U3822 ( .S(n3294), .A0(ixcSimTime[51]), .A1(n3324), .Z(n3323));
Q_MX04 U3823 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[51]), .A1(hwSimTime[51]), .A2(lockTraceTime[51]), .A3(nextDutTimeS[51]), .Z(n3324));
Q_MX02 U3824 ( .S(n3294), .A0(ixcSimTime[50]), .A1(n3326), .Z(n3325));
Q_MX04 U3825 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[50]), .A1(hwSimTime[50]), .A2(lockTraceTime[50]), .A3(nextDutTimeS[50]), .Z(n3326));
Q_MX02 U3826 ( .S(n3294), .A0(ixcSimTime[49]), .A1(n3328), .Z(n3327));
Q_MX04 U3827 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[49]), .A1(hwSimTime[49]), .A2(lockTraceTime[49]), .A3(nextDutTimeS[49]), .Z(n3328));
Q_MX02 U3828 ( .S(n3294), .A0(ixcSimTime[48]), .A1(n3330), .Z(n3329));
Q_MX04 U3829 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[48]), .A1(hwSimTime[48]), .A2(lockTraceTime[48]), .A3(nextDutTimeS[48]), .Z(n3330));
Q_MX02 U3830 ( .S(n3294), .A0(ixcSimTime[47]), .A1(n3332), .Z(n3331));
Q_MX04 U3831 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[47]), .A1(hwSimTime[47]), .A2(lockTraceTime[47]), .A3(nextDutTimeS[47]), .Z(n3332));
Q_MX02 U3832 ( .S(n3294), .A0(ixcSimTime[46]), .A1(n3334), .Z(n3333));
Q_MX04 U3833 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[46]), .A1(hwSimTime[46]), .A2(lockTraceTime[46]), .A3(nextDutTimeS[46]), .Z(n3334));
Q_MX02 U3834 ( .S(n3294), .A0(ixcSimTime[45]), .A1(n3336), .Z(n3335));
Q_MX04 U3835 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[45]), .A1(hwSimTime[45]), .A2(lockTraceTime[45]), .A3(nextDutTimeS[45]), .Z(n3336));
Q_MX02 U3836 ( .S(n3294), .A0(ixcSimTime[44]), .A1(n3338), .Z(n3337));
Q_MX04 U3837 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[44]), .A1(hwSimTime[44]), .A2(lockTraceTime[44]), .A3(nextDutTimeS[44]), .Z(n3338));
Q_MX02 U3838 ( .S(n3294), .A0(ixcSimTime[43]), .A1(n3340), .Z(n3339));
Q_MX04 U3839 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[43]), .A1(hwSimTime[43]), .A2(lockTraceTime[43]), .A3(nextDutTimeS[43]), .Z(n3340));
Q_MX02 U3840 ( .S(n3294), .A0(ixcSimTime[42]), .A1(n3342), .Z(n3341));
Q_MX04 U3841 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[42]), .A1(hwSimTime[42]), .A2(lockTraceTime[42]), .A3(nextDutTimeS[42]), .Z(n3342));
Q_MX02 U3842 ( .S(n3294), .A0(ixcSimTime[41]), .A1(n3344), .Z(n3343));
Q_MX04 U3843 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[41]), .A1(hwSimTime[41]), .A2(lockTraceTime[41]), .A3(nextDutTimeS[41]), .Z(n3344));
Q_MX02 U3844 ( .S(n3294), .A0(ixcSimTime[40]), .A1(n3346), .Z(n3345));
Q_MX04 U3845 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[40]), .A1(hwSimTime[40]), .A2(lockTraceTime[40]), .A3(nextDutTimeS[40]), .Z(n3346));
Q_MX02 U3846 ( .S(n3294), .A0(ixcSimTime[39]), .A1(n3348), .Z(n3347));
Q_MX04 U3847 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[39]), .A1(hwSimTime[39]), .A2(lockTraceTime[39]), .A3(nextDutTimeS[39]), .Z(n3348));
Q_MX02 U3848 ( .S(n3294), .A0(ixcSimTime[38]), .A1(n3350), .Z(n3349));
Q_MX04 U3849 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[38]), .A1(hwSimTime[38]), .A2(lockTraceTime[38]), .A3(nextDutTimeS[38]), .Z(n3350));
Q_MX02 U3850 ( .S(n3294), .A0(ixcSimTime[37]), .A1(n3352), .Z(n3351));
Q_MX04 U3851 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[37]), .A1(hwSimTime[37]), .A2(lockTraceTime[37]), .A3(nextDutTimeS[37]), .Z(n3352));
Q_MX02 U3852 ( .S(n3294), .A0(ixcSimTime[36]), .A1(n3354), .Z(n3353));
Q_MX04 U3853 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[36]), .A1(hwSimTime[36]), .A2(lockTraceTime[36]), .A3(nextDutTimeS[36]), .Z(n3354));
Q_MX02 U3854 ( .S(n3294), .A0(ixcSimTime[35]), .A1(n3356), .Z(n3355));
Q_MX04 U3855 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[35]), .A1(hwSimTime[35]), .A2(lockTraceTime[35]), .A3(nextDutTimeS[35]), .Z(n3356));
Q_MX02 U3856 ( .S(n3294), .A0(ixcSimTime[34]), .A1(n3358), .Z(n3357));
Q_MX04 U3857 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[34]), .A1(hwSimTime[34]), .A2(lockTraceTime[34]), .A3(nextDutTimeS[34]), .Z(n3358));
Q_MX02 U3858 ( .S(n3294), .A0(ixcSimTime[33]), .A1(n3360), .Z(n3359));
Q_MX04 U3859 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[33]), .A1(hwSimTime[33]), .A2(lockTraceTime[33]), .A3(nextDutTimeS[33]), .Z(n3360));
Q_MX02 U3860 ( .S(n3294), .A0(ixcSimTime[32]), .A1(n3362), .Z(n3361));
Q_MX04 U3861 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[32]), .A1(hwSimTime[32]), .A2(lockTraceTime[32]), .A3(nextDutTimeS[32]), .Z(n3362));
Q_MX02 U3862 ( .S(n3294), .A0(ixcSimTime[31]), .A1(n3364), .Z(n3363));
Q_MX04 U3863 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[31]), .A1(hwSimTime[31]), .A2(lockTraceTime[31]), .A3(nextDutTimeS[31]), .Z(n3364));
Q_MX02 U3864 ( .S(n3294), .A0(ixcSimTime[30]), .A1(n3366), .Z(n3365));
Q_MX04 U3865 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[30]), .A1(hwSimTime[30]), .A2(lockTraceTime[30]), .A3(nextDutTimeS[30]), .Z(n3366));
Q_MX02 U3866 ( .S(n3294), .A0(ixcSimTime[29]), .A1(n3368), .Z(n3367));
Q_MX04 U3867 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[29]), .A1(hwSimTime[29]), .A2(lockTraceTime[29]), .A3(nextDutTimeS[29]), .Z(n3368));
Q_MX02 U3868 ( .S(n3294), .A0(ixcSimTime[28]), .A1(n3370), .Z(n3369));
Q_MX04 U3869 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[28]), .A1(hwSimTime[28]), .A2(lockTraceTime[28]), .A3(nextDutTimeS[28]), .Z(n3370));
Q_MX02 U3870 ( .S(n3294), .A0(ixcSimTime[27]), .A1(n3372), .Z(n3371));
Q_MX04 U3871 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[27]), .A1(hwSimTime[27]), .A2(lockTraceTime[27]), .A3(nextDutTimeS[27]), .Z(n3372));
Q_MX02 U3872 ( .S(n3294), .A0(ixcSimTime[26]), .A1(n3374), .Z(n3373));
Q_MX04 U3873 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[26]), .A1(hwSimTime[26]), .A2(lockTraceTime[26]), .A3(nextDutTimeS[26]), .Z(n3374));
Q_MX02 U3874 ( .S(n3294), .A0(ixcSimTime[25]), .A1(n3376), .Z(n3375));
Q_MX04 U3875 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[25]), .A1(hwSimTime[25]), .A2(lockTraceTime[25]), .A3(nextDutTimeS[25]), .Z(n3376));
Q_MX02 U3876 ( .S(n3294), .A0(ixcSimTime[24]), .A1(n3378), .Z(n3377));
Q_MX04 U3877 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[24]), .A1(hwSimTime[24]), .A2(lockTraceTime[24]), .A3(nextDutTimeS[24]), .Z(n3378));
Q_MX02 U3878 ( .S(n3294), .A0(ixcSimTime[23]), .A1(n3380), .Z(n3379));
Q_MX04 U3879 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[23]), .A1(hwSimTime[23]), .A2(lockTraceTime[23]), .A3(nextDutTimeS[23]), .Z(n3380));
Q_MX02 U3880 ( .S(n3294), .A0(ixcSimTime[22]), .A1(n3382), .Z(n3381));
Q_MX04 U3881 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[22]), .A1(hwSimTime[22]), .A2(lockTraceTime[22]), .A3(nextDutTimeS[22]), .Z(n3382));
Q_MX02 U3882 ( .S(n3294), .A0(ixcSimTime[21]), .A1(n3384), .Z(n3383));
Q_MX04 U3883 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[21]), .A1(hwSimTime[21]), .A2(lockTraceTime[21]), .A3(nextDutTimeS[21]), .Z(n3384));
Q_MX02 U3884 ( .S(n3294), .A0(ixcSimTime[20]), .A1(n3386), .Z(n3385));
Q_MX04 U3885 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[20]), .A1(hwSimTime[20]), .A2(lockTraceTime[20]), .A3(nextDutTimeS[20]), .Z(n3386));
Q_MX02 U3886 ( .S(n3294), .A0(ixcSimTime[19]), .A1(n3388), .Z(n3387));
Q_MX04 U3887 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[19]), .A1(hwSimTime[19]), .A2(lockTraceTime[19]), .A3(nextDutTimeS[19]), .Z(n3388));
Q_MX02 U3888 ( .S(n3294), .A0(ixcSimTime[18]), .A1(n3390), .Z(n3389));
Q_MX04 U3889 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[18]), .A1(hwSimTime[18]), .A2(lockTraceTime[18]), .A3(nextDutTimeS[18]), .Z(n3390));
Q_MX02 U3890 ( .S(n3294), .A0(ixcSimTime[17]), .A1(n3392), .Z(n3391));
Q_MX04 U3891 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[17]), .A1(hwSimTime[17]), .A2(lockTraceTime[17]), .A3(nextDutTimeS[17]), .Z(n3392));
Q_MX02 U3892 ( .S(n3294), .A0(ixcSimTime[16]), .A1(n3394), .Z(n3393));
Q_MX04 U3893 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[16]), .A1(hwSimTime[16]), .A2(lockTraceTime[16]), .A3(nextDutTimeS[16]), .Z(n3394));
Q_MX02 U3894 ( .S(n3294), .A0(ixcSimTime[15]), .A1(n3396), .Z(n3395));
Q_MX04 U3895 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[15]), .A1(hwSimTime[15]), .A2(lockTraceTime[15]), .A3(nextDutTimeS[15]), .Z(n3396));
Q_MX02 U3896 ( .S(n3294), .A0(ixcSimTime[14]), .A1(n3398), .Z(n3397));
Q_MX04 U3897 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[14]), .A1(hwSimTime[14]), .A2(lockTraceTime[14]), .A3(nextDutTimeS[14]), .Z(n3398));
Q_MX02 U3898 ( .S(n3294), .A0(ixcSimTime[13]), .A1(n3400), .Z(n3399));
Q_MX04 U3899 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[13]), .A1(hwSimTime[13]), .A2(lockTraceTime[13]), .A3(nextDutTimeS[13]), .Z(n3400));
Q_MX02 U3900 ( .S(n3294), .A0(ixcSimTime[12]), .A1(n3402), .Z(n3401));
Q_MX04 U3901 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[12]), .A1(hwSimTime[12]), .A2(lockTraceTime[12]), .A3(nextDutTimeS[12]), .Z(n3402));
Q_MX02 U3902 ( .S(n3294), .A0(ixcSimTime[11]), .A1(n3404), .Z(n3403));
Q_MX04 U3903 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[11]), .A1(hwSimTime[11]), .A2(lockTraceTime[11]), .A3(nextDutTimeS[11]), .Z(n3404));
Q_MX02 U3904 ( .S(n3294), .A0(ixcSimTime[10]), .A1(n3406), .Z(n3405));
Q_MX04 U3905 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[10]), .A1(hwSimTime[10]), .A2(lockTraceTime[10]), .A3(nextDutTimeS[10]), .Z(n3406));
Q_MX02 U3906 ( .S(n3294), .A0(ixcSimTime[9]), .A1(n3408), .Z(n3407));
Q_MX04 U3907 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[9]), .A1(hwSimTime[9]), .A2(lockTraceTime[9]), .A3(nextDutTimeS[9]), .Z(n3408));
Q_MX02 U3908 ( .S(n3294), .A0(ixcSimTime[8]), .A1(n3410), .Z(n3409));
Q_MX04 U3909 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[8]), .A1(hwSimTime[8]), .A2(lockTraceTime[8]), .A3(nextDutTimeS[8]), .Z(n3410));
Q_MX02 U3910 ( .S(n3294), .A0(ixcSimTime[7]), .A1(n3412), .Z(n3411));
Q_MX04 U3911 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[7]), .A1(hwSimTime[7]), .A2(lockTraceTime[7]), .A3(nextDutTimeS[7]), .Z(n3412));
Q_MX02 U3912 ( .S(n3294), .A0(ixcSimTime[6]), .A1(n3414), .Z(n3413));
Q_MX04 U3913 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[6]), .A1(hwSimTime[6]), .A2(lockTraceTime[6]), .A3(nextDutTimeS[6]), .Z(n3414));
Q_MX02 U3914 ( .S(n3294), .A0(ixcSimTime[5]), .A1(n3416), .Z(n3415));
Q_MX04 U3915 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[5]), .A1(hwSimTime[5]), .A2(lockTraceTime[5]), .A3(nextDutTimeS[5]), .Z(n3416));
Q_MX02 U3916 ( .S(n3294), .A0(ixcSimTime[4]), .A1(n3418), .Z(n3417));
Q_MX04 U3917 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[4]), .A1(hwSimTime[4]), .A2(lockTraceTime[4]), .A3(nextDutTimeS[4]), .Z(n3418));
Q_MX02 U3918 ( .S(n3294), .A0(ixcSimTime[3]), .A1(n3420), .Z(n3419));
Q_MX04 U3919 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[3]), .A1(hwSimTime[3]), .A2(lockTraceTime[3]), .A3(nextDutTimeS[3]), .Z(n3420));
Q_MX02 U3920 ( .S(n3294), .A0(ixcSimTime[2]), .A1(n3422), .Z(n3421));
Q_MX04 U3921 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[2]), .A1(hwSimTime[2]), .A2(lockTraceTime[2]), .A3(nextDutTimeS[2]), .Z(n3422));
Q_MX02 U3922 ( .S(n3294), .A0(ixcSimTime[1]), .A1(n3424), .Z(n3423));
Q_MX04 U3923 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[1]), .A1(hwSimTime[1]), .A2(lockTraceTime[1]), .A3(nextDutTimeS[1]), .Z(n3424));
Q_MX02 U3924 ( .S(n3294), .A0(ixcSimTime[0]), .A1(n3426), .Z(n3425));
Q_MX04 U3925 ( .S0(n3291), .S1(n3290), .A0(ixc_time.nextTbTime[0]), .A1(hwSimTime[0]), .A2(lockTraceTime[0]), .A3(nextDutTimeS[0]), .Z(n3426));
Q_MX02 U3926 ( .S(oneStepPIi), .A0(ixc_time.simTime[63]), .A1(ixc_time.nextTbTime[63]), .Z(ixcSimTime[63]));
Q_MX02 U3927 ( .S(oneStepPIi), .A0(ixc_time.simTime[62]), .A1(ixc_time.nextTbTime[62]), .Z(ixcSimTime[62]));
Q_MX02 U3928 ( .S(oneStepPIi), .A0(ixc_time.simTime[61]), .A1(ixc_time.nextTbTime[61]), .Z(ixcSimTime[61]));
Q_MX02 U3929 ( .S(oneStepPIi), .A0(ixc_time.simTime[60]), .A1(ixc_time.nextTbTime[60]), .Z(ixcSimTime[60]));
Q_MX02 U3930 ( .S(oneStepPIi), .A0(ixc_time.simTime[59]), .A1(ixc_time.nextTbTime[59]), .Z(ixcSimTime[59]));
Q_MX02 U3931 ( .S(oneStepPIi), .A0(ixc_time.simTime[58]), .A1(ixc_time.nextTbTime[58]), .Z(ixcSimTime[58]));
Q_MX02 U3932 ( .S(oneStepPIi), .A0(ixc_time.simTime[57]), .A1(ixc_time.nextTbTime[57]), .Z(ixcSimTime[57]));
Q_MX02 U3933 ( .S(oneStepPIi), .A0(ixc_time.simTime[56]), .A1(ixc_time.nextTbTime[56]), .Z(ixcSimTime[56]));
Q_MX02 U3934 ( .S(oneStepPIi), .A0(ixc_time.simTime[55]), .A1(ixc_time.nextTbTime[55]), .Z(ixcSimTime[55]));
Q_MX02 U3935 ( .S(oneStepPIi), .A0(ixc_time.simTime[54]), .A1(ixc_time.nextTbTime[54]), .Z(ixcSimTime[54]));
Q_MX02 U3936 ( .S(oneStepPIi), .A0(ixc_time.simTime[53]), .A1(ixc_time.nextTbTime[53]), .Z(ixcSimTime[53]));
Q_MX02 U3937 ( .S(oneStepPIi), .A0(ixc_time.simTime[52]), .A1(ixc_time.nextTbTime[52]), .Z(ixcSimTime[52]));
Q_MX02 U3938 ( .S(oneStepPIi), .A0(ixc_time.simTime[51]), .A1(ixc_time.nextTbTime[51]), .Z(ixcSimTime[51]));
Q_MX02 U3939 ( .S(oneStepPIi), .A0(ixc_time.simTime[50]), .A1(ixc_time.nextTbTime[50]), .Z(ixcSimTime[50]));
Q_MX02 U3940 ( .S(oneStepPIi), .A0(ixc_time.simTime[49]), .A1(ixc_time.nextTbTime[49]), .Z(ixcSimTime[49]));
Q_MX02 U3941 ( .S(oneStepPIi), .A0(ixc_time.simTime[48]), .A1(ixc_time.nextTbTime[48]), .Z(ixcSimTime[48]));
Q_MX02 U3942 ( .S(oneStepPIi), .A0(ixc_time.simTime[47]), .A1(ixc_time.nextTbTime[47]), .Z(ixcSimTime[47]));
Q_MX02 U3943 ( .S(oneStepPIi), .A0(ixc_time.simTime[46]), .A1(ixc_time.nextTbTime[46]), .Z(ixcSimTime[46]));
Q_MX02 U3944 ( .S(oneStepPIi), .A0(ixc_time.simTime[45]), .A1(ixc_time.nextTbTime[45]), .Z(ixcSimTime[45]));
Q_MX02 U3945 ( .S(oneStepPIi), .A0(ixc_time.simTime[44]), .A1(ixc_time.nextTbTime[44]), .Z(ixcSimTime[44]));
Q_MX02 U3946 ( .S(oneStepPIi), .A0(ixc_time.simTime[43]), .A1(ixc_time.nextTbTime[43]), .Z(ixcSimTime[43]));
Q_MX02 U3947 ( .S(oneStepPIi), .A0(ixc_time.simTime[42]), .A1(ixc_time.nextTbTime[42]), .Z(ixcSimTime[42]));
Q_MX02 U3948 ( .S(oneStepPIi), .A0(ixc_time.simTime[41]), .A1(ixc_time.nextTbTime[41]), .Z(ixcSimTime[41]));
Q_MX02 U3949 ( .S(oneStepPIi), .A0(ixc_time.simTime[40]), .A1(ixc_time.nextTbTime[40]), .Z(ixcSimTime[40]));
Q_MX02 U3950 ( .S(oneStepPIi), .A0(ixc_time.simTime[39]), .A1(ixc_time.nextTbTime[39]), .Z(ixcSimTime[39]));
Q_MX02 U3951 ( .S(oneStepPIi), .A0(ixc_time.simTime[38]), .A1(ixc_time.nextTbTime[38]), .Z(ixcSimTime[38]));
Q_MX02 U3952 ( .S(oneStepPIi), .A0(ixc_time.simTime[37]), .A1(ixc_time.nextTbTime[37]), .Z(ixcSimTime[37]));
Q_MX02 U3953 ( .S(oneStepPIi), .A0(ixc_time.simTime[36]), .A1(ixc_time.nextTbTime[36]), .Z(ixcSimTime[36]));
Q_MX02 U3954 ( .S(oneStepPIi), .A0(ixc_time.simTime[35]), .A1(ixc_time.nextTbTime[35]), .Z(ixcSimTime[35]));
Q_MX02 U3955 ( .S(oneStepPIi), .A0(ixc_time.simTime[34]), .A1(ixc_time.nextTbTime[34]), .Z(ixcSimTime[34]));
Q_MX02 U3956 ( .S(oneStepPIi), .A0(ixc_time.simTime[33]), .A1(ixc_time.nextTbTime[33]), .Z(ixcSimTime[33]));
Q_MX02 U3957 ( .S(oneStepPIi), .A0(ixc_time.simTime[32]), .A1(ixc_time.nextTbTime[32]), .Z(ixcSimTime[32]));
Q_MX02 U3958 ( .S(oneStepPIi), .A0(ixc_time.simTime[31]), .A1(ixc_time.nextTbTime[31]), .Z(ixcSimTime[31]));
Q_MX02 U3959 ( .S(oneStepPIi), .A0(ixc_time.simTime[30]), .A1(ixc_time.nextTbTime[30]), .Z(ixcSimTime[30]));
Q_MX02 U3960 ( .S(oneStepPIi), .A0(ixc_time.simTime[29]), .A1(ixc_time.nextTbTime[29]), .Z(ixcSimTime[29]));
Q_MX02 U3961 ( .S(oneStepPIi), .A0(ixc_time.simTime[28]), .A1(ixc_time.nextTbTime[28]), .Z(ixcSimTime[28]));
Q_MX02 U3962 ( .S(oneStepPIi), .A0(ixc_time.simTime[27]), .A1(ixc_time.nextTbTime[27]), .Z(ixcSimTime[27]));
Q_MX02 U3963 ( .S(oneStepPIi), .A0(ixc_time.simTime[26]), .A1(ixc_time.nextTbTime[26]), .Z(ixcSimTime[26]));
Q_MX02 U3964 ( .S(oneStepPIi), .A0(ixc_time.simTime[25]), .A1(ixc_time.nextTbTime[25]), .Z(ixcSimTime[25]));
Q_MX02 U3965 ( .S(oneStepPIi), .A0(ixc_time.simTime[24]), .A1(ixc_time.nextTbTime[24]), .Z(ixcSimTime[24]));
Q_MX02 U3966 ( .S(oneStepPIi), .A0(ixc_time.simTime[23]), .A1(ixc_time.nextTbTime[23]), .Z(ixcSimTime[23]));
Q_MX02 U3967 ( .S(oneStepPIi), .A0(ixc_time.simTime[22]), .A1(ixc_time.nextTbTime[22]), .Z(ixcSimTime[22]));
Q_MX02 U3968 ( .S(oneStepPIi), .A0(ixc_time.simTime[21]), .A1(ixc_time.nextTbTime[21]), .Z(ixcSimTime[21]));
Q_MX02 U3969 ( .S(oneStepPIi), .A0(ixc_time.simTime[20]), .A1(ixc_time.nextTbTime[20]), .Z(ixcSimTime[20]));
Q_MX02 U3970 ( .S(oneStepPIi), .A0(ixc_time.simTime[19]), .A1(ixc_time.nextTbTime[19]), .Z(ixcSimTime[19]));
Q_MX02 U3971 ( .S(oneStepPIi), .A0(ixc_time.simTime[18]), .A1(ixc_time.nextTbTime[18]), .Z(ixcSimTime[18]));
Q_MX02 U3972 ( .S(oneStepPIi), .A0(ixc_time.simTime[17]), .A1(ixc_time.nextTbTime[17]), .Z(ixcSimTime[17]));
Q_MX02 U3973 ( .S(oneStepPIi), .A0(ixc_time.simTime[16]), .A1(ixc_time.nextTbTime[16]), .Z(ixcSimTime[16]));
Q_MX02 U3974 ( .S(oneStepPIi), .A0(ixc_time.simTime[15]), .A1(ixc_time.nextTbTime[15]), .Z(ixcSimTime[15]));
Q_MX02 U3975 ( .S(oneStepPIi), .A0(ixc_time.simTime[14]), .A1(ixc_time.nextTbTime[14]), .Z(ixcSimTime[14]));
Q_MX02 U3976 ( .S(oneStepPIi), .A0(ixc_time.simTime[13]), .A1(ixc_time.nextTbTime[13]), .Z(ixcSimTime[13]));
Q_MX02 U3977 ( .S(oneStepPIi), .A0(ixc_time.simTime[12]), .A1(ixc_time.nextTbTime[12]), .Z(ixcSimTime[12]));
Q_MX02 U3978 ( .S(oneStepPIi), .A0(ixc_time.simTime[11]), .A1(ixc_time.nextTbTime[11]), .Z(ixcSimTime[11]));
Q_MX02 U3979 ( .S(oneStepPIi), .A0(ixc_time.simTime[10]), .A1(ixc_time.nextTbTime[10]), .Z(ixcSimTime[10]));
Q_MX02 U3980 ( .S(oneStepPIi), .A0(ixc_time.simTime[9]), .A1(ixc_time.nextTbTime[9]), .Z(ixcSimTime[9]));
Q_MX02 U3981 ( .S(oneStepPIi), .A0(ixc_time.simTime[8]), .A1(ixc_time.nextTbTime[8]), .Z(ixcSimTime[8]));
Q_MX02 U3982 ( .S(oneStepPIi), .A0(ixc_time.simTime[7]), .A1(ixc_time.nextTbTime[7]), .Z(ixcSimTime[7]));
Q_MX02 U3983 ( .S(oneStepPIi), .A0(ixc_time.simTime[6]), .A1(ixc_time.nextTbTime[6]), .Z(ixcSimTime[6]));
Q_MX02 U3984 ( .S(oneStepPIi), .A0(ixc_time.simTime[5]), .A1(ixc_time.nextTbTime[5]), .Z(ixcSimTime[5]));
Q_MX02 U3985 ( .S(oneStepPIi), .A0(ixc_time.simTime[4]), .A1(ixc_time.nextTbTime[4]), .Z(ixcSimTime[4]));
Q_MX02 U3986 ( .S(oneStepPIi), .A0(ixc_time.simTime[3]), .A1(ixc_time.nextTbTime[3]), .Z(ixcSimTime[3]));
Q_MX02 U3987 ( .S(oneStepPIi), .A0(ixc_time.simTime[2]), .A1(ixc_time.nextTbTime[2]), .Z(ixcSimTime[2]));
Q_MX02 U3988 ( .S(oneStepPIi), .A0(ixc_time.simTime[1]), .A1(ixc_time.nextTbTime[1]), .Z(ixcSimTime[1]));
Q_MX02 U3989 ( .S(oneStepPIi), .A0(ixc_time.simTime[0]), .A1(ixc_time.nextTbTime[0]), .Z(ixcSimTime[0]));
Q_FDP0 \nextDutTimeS_REG[63] ( .CK(uClk), .D(ixc_time.nextDutTime[63]), .Q(nextDutTimeS[63]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[62] ( .CK(uClk), .D(ixc_time.nextDutTime[62]), .Q(nextDutTimeS[62]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[61] ( .CK(uClk), .D(ixc_time.nextDutTime[61]), .Q(nextDutTimeS[61]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[60] ( .CK(uClk), .D(ixc_time.nextDutTime[60]), .Q(nextDutTimeS[60]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[59] ( .CK(uClk), .D(ixc_time.nextDutTime[59]), .Q(nextDutTimeS[59]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[58] ( .CK(uClk), .D(ixc_time.nextDutTime[58]), .Q(nextDutTimeS[58]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[57] ( .CK(uClk), .D(ixc_time.nextDutTime[57]), .Q(nextDutTimeS[57]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[56] ( .CK(uClk), .D(ixc_time.nextDutTime[56]), .Q(nextDutTimeS[56]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[55] ( .CK(uClk), .D(ixc_time.nextDutTime[55]), .Q(nextDutTimeS[55]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[54] ( .CK(uClk), .D(ixc_time.nextDutTime[54]), .Q(nextDutTimeS[54]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[53] ( .CK(uClk), .D(ixc_time.nextDutTime[53]), .Q(nextDutTimeS[53]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[52] ( .CK(uClk), .D(ixc_time.nextDutTime[52]), .Q(nextDutTimeS[52]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[51] ( .CK(uClk), .D(ixc_time.nextDutTime[51]), .Q(nextDutTimeS[51]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[50] ( .CK(uClk), .D(ixc_time.nextDutTime[50]), .Q(nextDutTimeS[50]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[49] ( .CK(uClk), .D(ixc_time.nextDutTime[49]), .Q(nextDutTimeS[49]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[48] ( .CK(uClk), .D(ixc_time.nextDutTime[48]), .Q(nextDutTimeS[48]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[47] ( .CK(uClk), .D(ixc_time.nextDutTime[47]), .Q(nextDutTimeS[47]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[46] ( .CK(uClk), .D(ixc_time.nextDutTime[46]), .Q(nextDutTimeS[46]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[45] ( .CK(uClk), .D(ixc_time.nextDutTime[45]), .Q(nextDutTimeS[45]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[44] ( .CK(uClk), .D(ixc_time.nextDutTime[44]), .Q(nextDutTimeS[44]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[43] ( .CK(uClk), .D(ixc_time.nextDutTime[43]), .Q(nextDutTimeS[43]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[42] ( .CK(uClk), .D(ixc_time.nextDutTime[42]), .Q(nextDutTimeS[42]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[41] ( .CK(uClk), .D(ixc_time.nextDutTime[41]), .Q(nextDutTimeS[41]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[40] ( .CK(uClk), .D(ixc_time.nextDutTime[40]), .Q(nextDutTimeS[40]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[39] ( .CK(uClk), .D(ixc_time.nextDutTime[39]), .Q(nextDutTimeS[39]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[38] ( .CK(uClk), .D(ixc_time.nextDutTime[38]), .Q(nextDutTimeS[38]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[37] ( .CK(uClk), .D(ixc_time.nextDutTime[37]), .Q(nextDutTimeS[37]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[36] ( .CK(uClk), .D(ixc_time.nextDutTime[36]), .Q(nextDutTimeS[36]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[35] ( .CK(uClk), .D(ixc_time.nextDutTime[35]), .Q(nextDutTimeS[35]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[34] ( .CK(uClk), .D(ixc_time.nextDutTime[34]), .Q(nextDutTimeS[34]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[33] ( .CK(uClk), .D(ixc_time.nextDutTime[33]), .Q(nextDutTimeS[33]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[32] ( .CK(uClk), .D(ixc_time.nextDutTime[32]), .Q(nextDutTimeS[32]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[31] ( .CK(uClk), .D(ixc_time.nextDutTime[31]), .Q(nextDutTimeS[31]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[30] ( .CK(uClk), .D(ixc_time.nextDutTime[30]), .Q(nextDutTimeS[30]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[29] ( .CK(uClk), .D(ixc_time.nextDutTime[29]), .Q(nextDutTimeS[29]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[28] ( .CK(uClk), .D(ixc_time.nextDutTime[28]), .Q(nextDutTimeS[28]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[27] ( .CK(uClk), .D(ixc_time.nextDutTime[27]), .Q(nextDutTimeS[27]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[26] ( .CK(uClk), .D(ixc_time.nextDutTime[26]), .Q(nextDutTimeS[26]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[25] ( .CK(uClk), .D(ixc_time.nextDutTime[25]), .Q(nextDutTimeS[25]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[24] ( .CK(uClk), .D(ixc_time.nextDutTime[24]), .Q(nextDutTimeS[24]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[23] ( .CK(uClk), .D(ixc_time.nextDutTime[23]), .Q(nextDutTimeS[23]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[22] ( .CK(uClk), .D(ixc_time.nextDutTime[22]), .Q(nextDutTimeS[22]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[21] ( .CK(uClk), .D(ixc_time.nextDutTime[21]), .Q(nextDutTimeS[21]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[20] ( .CK(uClk), .D(ixc_time.nextDutTime[20]), .Q(nextDutTimeS[20]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[19] ( .CK(uClk), .D(ixc_time.nextDutTime[19]), .Q(nextDutTimeS[19]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[18] ( .CK(uClk), .D(ixc_time.nextDutTime[18]), .Q(nextDutTimeS[18]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[17] ( .CK(uClk), .D(ixc_time.nextDutTime[17]), .Q(nextDutTimeS[17]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[16] ( .CK(uClk), .D(ixc_time.nextDutTime[16]), .Q(nextDutTimeS[16]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[15] ( .CK(uClk), .D(ixc_time.nextDutTime[15]), .Q(nextDutTimeS[15]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[14] ( .CK(uClk), .D(ixc_time.nextDutTime[14]), .Q(nextDutTimeS[14]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[13] ( .CK(uClk), .D(ixc_time.nextDutTime[13]), .Q(nextDutTimeS[13]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[12] ( .CK(uClk), .D(ixc_time.nextDutTime[12]), .Q(nextDutTimeS[12]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[11] ( .CK(uClk), .D(ixc_time.nextDutTime[11]), .Q(nextDutTimeS[11]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[10] ( .CK(uClk), .D(ixc_time.nextDutTime[10]), .Q(nextDutTimeS[10]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[9] ( .CK(uClk), .D(ixc_time.nextDutTime[9]), .Q(nextDutTimeS[9]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[8] ( .CK(uClk), .D(ixc_time.nextDutTime[8]), .Q(nextDutTimeS[8]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[7] ( .CK(uClk), .D(ixc_time.nextDutTime[7]), .Q(nextDutTimeS[7]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[6] ( .CK(uClk), .D(ixc_time.nextDutTime[6]), .Q(nextDutTimeS[6]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[5] ( .CK(uClk), .D(ixc_time.nextDutTime[5]), .Q(nextDutTimeS[5]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[4] ( .CK(uClk), .D(ixc_time.nextDutTime[4]), .Q(nextDutTimeS[4]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[3] ( .CK(uClk), .D(ixc_time.nextDutTime[3]), .Q(nextDutTimeS[3]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[2] ( .CK(uClk), .D(ixc_time.nextDutTime[2]), .Q(nextDutTimeS[2]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[1] ( .CK(uClk), .D(ixc_time.nextDutTime[1]), .Q(nextDutTimeS[1]), .QN( ));
Q_FDP0 \nextDutTimeS_REG[0] ( .CK(uClk), .D(ixc_time.nextDutTime[0]), .Q(nextDutTimeS[0]), .QN( ));
Q_LDP0 oneStepPImio_REG  ( .G(n3427), .D(mioPIW_1[4]), .Q(oneStepPImio), .QN( ));
Q_LDP0 ckgHoldPImio_REG  ( .G(n3427), .D(mioPIW_1[2]), .Q(ckgHoldPImio), .QN( ));
Q_LDP0 callEmuPImio_REG  ( .G(n3427), .D(mioPIW_1[1]), .Q(callEmuPImio), .QN( ));
Q_LDP0 \evalStepPImio_REG[0] ( .G(n3427), .D(mioPIW_0[0]), .Q(evalStepPImio[0]), .QN( ));
Q_LDP0 \evalStepPImio_REG[1] ( .G(n3427), .D(mioPIW_0[1]), .Q(evalStepPImio[1]), .QN( ));
Q_LDP0 \evalStepPImio_REG[2] ( .G(n3427), .D(mioPIW_0[2]), .Q(evalStepPImio[2]), .QN( ));
Q_LDP0 \evalStepPImio_REG[3] ( .G(n3427), .D(mioPIW_0[3]), .Q(evalStepPImio[3]), .QN( ));
Q_LDP0 \evalStepPImio_REG[4] ( .G(n3427), .D(mioPIW_0[4]), .Q(evalStepPImio[4]), .QN( ));
Q_LDP0 \evalStepPImio_REG[5] ( .G(n3427), .D(mioPIW_0[5]), .Q(evalStepPImio[5]), .QN( ));
Q_LDP0 \evalStepPImio_REG[6] ( .G(n3427), .D(mioPIW_0[6]), .Q(evalStepPImio[6]), .QN( ));
Q_LDP0 \evalStepPImio_REG[7] ( .G(n3427), .D(mioPIW_0[7]), .Q(evalStepPImio[7]), .QN( ));
Q_LDP0 \evalStepPImio_REG[8] ( .G(n3427), .D(mioPIW_0[8]), .Q(evalStepPImio[8]), .QN( ));
Q_LDP0 \evalStepPImio_REG[9] ( .G(n3427), .D(mioPIW_0[9]), .Q(evalStepPImio[9]), .QN( ));
Q_LDP0 \evalStepPImio_REG[10] ( .G(n3427), .D(mioPIW_0[10]), .Q(evalStepPImio[10]), .QN( ));
Q_LDP0 \evalStepPImio_REG[11] ( .G(n3427), .D(mioPIW_0[11]), .Q(evalStepPImio[11]), .QN( ));
Q_LDP0 \evalStepPImio_REG[12] ( .G(n3427), .D(mioPIW_0[12]), .Q(evalStepPImio[12]), .QN( ));
Q_LDP0 \evalStepPImio_REG[13] ( .G(n3427), .D(mioPIW_0[13]), .Q(evalStepPImio[13]), .QN( ));
Q_LDP0 \evalStepPImio_REG[14] ( .G(n3427), .D(mioPIW_0[14]), .Q(evalStepPImio[14]), .QN( ));
Q_LDP0 \evalStepPImio_REG[15] ( .G(n3427), .D(mioPIW_0[15]), .Q(evalStepPImio[15]), .QN( ));
Q_LDP0 \evalStepPImio_REG[16] ( .G(n3427), .D(mioPIW_0[16]), .Q(evalStepPImio[16]), .QN( ));
Q_LDP0 \evalStepPImio_REG[17] ( .G(n3427), .D(mioPIW_0[17]), .Q(evalStepPImio[17]), .QN( ));
Q_LDP0 \evalStepPImio_REG[18] ( .G(n3427), .D(mioPIW_0[18]), .Q(evalStepPImio[18]), .QN( ));
Q_LDP0 \evalStepPImio_REG[19] ( .G(n3427), .D(mioPIW_0[19]), .Q(evalStepPImio[19]), .QN( ));
Q_LDP0 \evalStepPImio_REG[20] ( .G(n3427), .D(mioPIW_0[20]), .Q(evalStepPImio[20]), .QN( ));
Q_LDP0 \evalStepPImio_REG[21] ( .G(n3427), .D(mioPIW_0[21]), .Q(evalStepPImio[21]), .QN( ));
Q_LDP0 \evalStepPImio_REG[22] ( .G(n3427), .D(mioPIW_0[22]), .Q(evalStepPImio[22]), .QN( ));
Q_LDP0 \evalStepPImio_REG[23] ( .G(n3427), .D(mioPIW_0[23]), .Q(evalStepPImio[23]), .QN( ));
Q_LDP0 \evalStepPImio_REG[24] ( .G(n3427), .D(mioPIW_0[24]), .Q(evalStepPImio[24]), .QN( ));
Q_LDP0 \evalStepPImio_REG[25] ( .G(n3427), .D(mioPIW_0[25]), .Q(evalStepPImio[25]), .QN( ));
Q_LDP0 \evalStepPImio_REG[26] ( .G(n3427), .D(mioPIW_0[26]), .Q(evalStepPImio[26]), .QN( ));
Q_LDP0 \evalStepPImio_REG[27] ( .G(n3427), .D(mioPIW_0[27]), .Q(evalStepPImio[27]), .QN( ));
Q_LDP0 \evalStepPImio_REG[28] ( .G(n3427), .D(mioPIW_0[28]), .Q(evalStepPImio[28]), .QN( ));
Q_LDP0 \evalStepPImio_REG[29] ( .G(n3427), .D(mioPIW_0[29]), .Q(evalStepPImio[29]), .QN( ));
Q_LDP0 \evalStepPImio_REG[30] ( .G(n3427), .D(mioPIW_0[30]), .Q(evalStepPImio[30]), .QN( ));
Q_LDP0 \evalStepPImio_REG[31] ( .G(n3427), .D(mioPIW_0[31]), .Q(evalStepPImio[31]), .QN( ));
Q_LDP0 \evalStepPImio_REG[32] ( .G(n3427), .D(mioPIW_0[32]), .Q(evalStepPImio[32]), .QN( ));
Q_LDP0 \evalStepPImio_REG[33] ( .G(n3427), .D(mioPIW_0[33]), .Q(evalStepPImio[33]), .QN( ));
Q_LDP0 \evalStepPImio_REG[34] ( .G(n3427), .D(mioPIW_0[34]), .Q(evalStepPImio[34]), .QN( ));
Q_LDP0 \evalStepPImio_REG[35] ( .G(n3427), .D(mioPIW_0[35]), .Q(evalStepPImio[35]), .QN( ));
Q_LDP0 \evalStepPImio_REG[36] ( .G(n3427), .D(mioPIW_0[36]), .Q(evalStepPImio[36]), .QN( ));
Q_LDP0 \evalStepPImio_REG[37] ( .G(n3427), .D(mioPIW_0[37]), .Q(evalStepPImio[37]), .QN( ));
Q_LDP0 \evalStepPImio_REG[38] ( .G(n3427), .D(mioPIW_0[38]), .Q(evalStepPImio[38]), .QN( ));
Q_LDP0 \evalStepPImio_REG[39] ( .G(n3427), .D(mioPIW_0[39]), .Q(evalStepPImio[39]), .QN( ));
Q_LDP0 \evalStepPImio_REG[40] ( .G(n3427), .D(mioPIW_0[40]), .Q(evalStepPImio[40]), .QN( ));
Q_LDP0 \evalStepPImio_REG[41] ( .G(n3427), .D(mioPIW_0[41]), .Q(evalStepPImio[41]), .QN( ));
Q_LDP0 \evalStepPImio_REG[42] ( .G(n3427), .D(mioPIW_0[42]), .Q(evalStepPImio[42]), .QN( ));
Q_LDP0 \evalStepPImio_REG[43] ( .G(n3427), .D(mioPIW_0[43]), .Q(evalStepPImio[43]), .QN( ));
Q_LDP0 \evalStepPImio_REG[44] ( .G(n3427), .D(mioPIW_0[44]), .Q(evalStepPImio[44]), .QN( ));
Q_LDP0 \evalStepPImio_REG[45] ( .G(n3427), .D(mioPIW_0[45]), .Q(evalStepPImio[45]), .QN( ));
Q_LDP0 \evalStepPImio_REG[46] ( .G(n3427), .D(mioPIW_0[46]), .Q(evalStepPImio[46]), .QN( ));
Q_LDP0 \evalStepPImio_REG[47] ( .G(n3427), .D(mioPIW_0[47]), .Q(evalStepPImio[47]), .QN( ));
Q_LDP0 \evalStepPImio_REG[48] ( .G(n3427), .D(mioPIW_0[48]), .Q(evalStepPImio[48]), .QN( ));
Q_LDP0 \evalStepPImio_REG[49] ( .G(n3427), .D(mioPIW_0[49]), .Q(evalStepPImio[49]), .QN( ));
Q_LDP0 \evalStepPImio_REG[50] ( .G(n3427), .D(mioPIW_0[50]), .Q(evalStepPImio[50]), .QN( ));
Q_LDP0 \evalStepPImio_REG[51] ( .G(n3427), .D(mioPIW_0[51]), .Q(evalStepPImio[51]), .QN( ));
Q_LDP0 \evalStepPImio_REG[52] ( .G(n3427), .D(mioPIW_0[52]), .Q(evalStepPImio[52]), .QN( ));
Q_LDP0 \evalStepPImio_REG[53] ( .G(n3427), .D(mioPIW_0[53]), .Q(evalStepPImio[53]), .QN( ));
Q_LDP0 \evalStepPImio_REG[54] ( .G(n3427), .D(mioPIW_0[54]), .Q(evalStepPImio[54]), .QN( ));
Q_LDP0 \evalStepPImio_REG[55] ( .G(n3427), .D(mioPIW_0[55]), .Q(evalStepPImio[55]), .QN( ));
Q_LDP0 \evalStepPImio_REG[56] ( .G(n3427), .D(mioPIW_0[56]), .Q(evalStepPImio[56]), .QN( ));
Q_LDP0 \evalStepPImio_REG[57] ( .G(n3427), .D(mioPIW_0[57]), .Q(evalStepPImio[57]), .QN( ));
Q_LDP0 \evalStepPImio_REG[58] ( .G(n3427), .D(mioPIW_0[58]), .Q(evalStepPImio[58]), .QN( ));
Q_LDP0 \evalStepPImio_REG[59] ( .G(n3427), .D(mioPIW_0[59]), .Q(evalStepPImio[59]), .QN( ));
Q_LDP0 \evalStepPImio_REG[60] ( .G(n3427), .D(mioPIW_0[60]), .Q(evalStepPImio[60]), .QN( ));
Q_LDP0 \evalStepPImio_REG[61] ( .G(n3427), .D(mioPIW_0[61]), .Q(evalStepPImio[61]), .QN( ));
Q_LDP0 \evalStepPImio_REG[62] ( .G(n3427), .D(mioPIW_0[62]), .Q(evalStepPImio[62]), .QN( ));
Q_LDP0 \evalStepPImio_REG[63] ( .G(n3427), .D(mioPIW_0[63]), .Q(evalStepPImio[63]), .QN( ));
Q_XOR2 U4121 ( .A0(mioPICnt), .A1(mioPICntd), .Z(n3427));
Q_AN03 U4122 ( .A0(xc_mioOnS), .A1(n3429), .A2(mioPOW_2[1]), .Z(n3428));
Q_FDP0 tbcPOmio_REG  ( .CK(uClk), .D(mioPOW_2[1]), .Q(tbcPOmio), .QN(n3429));
Q_FDP0 xc_mioOnS_REG  ( .CK(uClk), .D(xc_mioOn), .Q(xc_mioOnS), .QN( ));
Q_OR03 U4125 ( .A0(bpHalt), .A1(acHalt), .A2(forceAbort), .Z(n3435));
Q_NR02 U4126 ( .A0(lockTrace), .A1(lockTraceC[2]), .Z(n3434));
Q_NR02 U4127 ( .A0(lockTraceC[1]), .A1(lockTraceC[0]), .Z(n3433));
Q_AN02 U4128 ( .A0(n3434), .A1(n3433), .Z(n3437));
Q_AN02 U4129 ( .A0(n3437), .A1(n3435), .Z(n3430));
Q_INV U4130 ( .A(n3437), .Z(n3431));
Q_INV U4131 ( .A(n3435), .Z(n3436));
Q_MX02 U4132 ( .S(n3437), .A0(lockTrace), .A1(n3436), .Z(n3438));
Q_AN02 U4133 ( .A0(n3431), .A1(n3443), .Z(n3439));
Q_AN02 U4134 ( .A0(n3431), .A1(n3445), .Z(n3440));
Q_AN02 U4135 ( .A0(n3431), .A1(n3447), .Z(n3441));
Q_OR02 U4136 ( .A0(n3437), .A1(n3432), .Z(n3442));
Q_XOR2 U4137 ( .A0(lockTrace), .A1(n3444), .Z(n3443));
Q_AD01HF U4138 ( .A0(lockTraceC[2]), .B0(n3446), .S(n3445), .CO(n3444));
Q_AD01HF U4139 ( .A0(lockTraceC[1]), .B0(lockTraceC[0]), .S(n3447), .CO(n3446));
Q_XOR2 U4140 ( .A0(simTime[63]), .A1(n3449), .Z(n3448));
Q_AD01HF U4141 ( .A0(simTime[62]), .B0(n3451), .S(n3450), .CO(n3449));
Q_AD01HF U4142 ( .A0(simTime[61]), .B0(n3453), .S(n3452), .CO(n3451));
Q_AD01HF U4143 ( .A0(simTime[60]), .B0(n3455), .S(n3454), .CO(n3453));
Q_AD01HF U4144 ( .A0(simTime[59]), .B0(n3457), .S(n3456), .CO(n3455));
Q_AD01HF U4145 ( .A0(simTime[58]), .B0(n3459), .S(n3458), .CO(n3457));
Q_AD01HF U4146 ( .A0(simTime[57]), .B0(n3461), .S(n3460), .CO(n3459));
Q_AD01HF U4147 ( .A0(simTime[56]), .B0(n3463), .S(n3462), .CO(n3461));
Q_AD01HF U4148 ( .A0(simTime[55]), .B0(n3465), .S(n3464), .CO(n3463));
Q_AD01HF U4149 ( .A0(simTime[54]), .B0(n3467), .S(n3466), .CO(n3465));
Q_AD01HF U4150 ( .A0(simTime[53]), .B0(n3469), .S(n3468), .CO(n3467));
Q_AD01HF U4151 ( .A0(simTime[52]), .B0(n3471), .S(n3470), .CO(n3469));
Q_AD01HF U4152 ( .A0(simTime[51]), .B0(n3473), .S(n3472), .CO(n3471));
Q_AD01HF U4153 ( .A0(simTime[50]), .B0(n3475), .S(n3474), .CO(n3473));
Q_AD01HF U4154 ( .A0(simTime[49]), .B0(n3477), .S(n3476), .CO(n3475));
Q_AD01HF U4155 ( .A0(simTime[48]), .B0(n3479), .S(n3478), .CO(n3477));
Q_AD01HF U4156 ( .A0(simTime[47]), .B0(n3481), .S(n3480), .CO(n3479));
Q_AD01HF U4157 ( .A0(simTime[46]), .B0(n3483), .S(n3482), .CO(n3481));
Q_AD01HF U4158 ( .A0(simTime[45]), .B0(n3485), .S(n3484), .CO(n3483));
Q_AD01HF U4159 ( .A0(simTime[44]), .B0(n3487), .S(n3486), .CO(n3485));
Q_AD01HF U4160 ( .A0(simTime[43]), .B0(n3489), .S(n3488), .CO(n3487));
Q_AD01HF U4161 ( .A0(simTime[42]), .B0(n3491), .S(n3490), .CO(n3489));
Q_AD01HF U4162 ( .A0(simTime[41]), .B0(n3493), .S(n3492), .CO(n3491));
Q_AD01HF U4163 ( .A0(simTime[40]), .B0(n3495), .S(n3494), .CO(n3493));
Q_AD01HF U4164 ( .A0(simTime[39]), .B0(n3497), .S(n3496), .CO(n3495));
Q_AD01HF U4165 ( .A0(simTime[38]), .B0(n3499), .S(n3498), .CO(n3497));
Q_AD01HF U4166 ( .A0(simTime[37]), .B0(n3501), .S(n3500), .CO(n3499));
Q_AD01HF U4167 ( .A0(simTime[36]), .B0(n3503), .S(n3502), .CO(n3501));
Q_AD01HF U4168 ( .A0(simTime[35]), .B0(n3505), .S(n3504), .CO(n3503));
Q_AD01HF U4169 ( .A0(simTime[34]), .B0(n3507), .S(n3506), .CO(n3505));
Q_AD01HF U4170 ( .A0(simTime[33]), .B0(n3509), .S(n3508), .CO(n3507));
Q_AD01HF U4171 ( .A0(simTime[32]), .B0(n3511), .S(n3510), .CO(n3509));
Q_AD01HF U4172 ( .A0(simTime[31]), .B0(n3513), .S(n3512), .CO(n3511));
Q_AD01HF U4173 ( .A0(simTime[30]), .B0(n3515), .S(n3514), .CO(n3513));
Q_AD01HF U4174 ( .A0(simTime[29]), .B0(n3517), .S(n3516), .CO(n3515));
Q_AD01HF U4175 ( .A0(simTime[28]), .B0(n3519), .S(n3518), .CO(n3517));
Q_AD01HF U4176 ( .A0(simTime[27]), .B0(n3521), .S(n3520), .CO(n3519));
Q_AD01HF U4177 ( .A0(simTime[26]), .B0(n3523), .S(n3522), .CO(n3521));
Q_AD01HF U4178 ( .A0(simTime[25]), .B0(n3525), .S(n3524), .CO(n3523));
Q_AD01HF U4179 ( .A0(simTime[24]), .B0(n3527), .S(n3526), .CO(n3525));
Q_AD01HF U4180 ( .A0(simTime[23]), .B0(n3529), .S(n3528), .CO(n3527));
Q_AD01HF U4181 ( .A0(simTime[22]), .B0(n3531), .S(n3530), .CO(n3529));
Q_AD01HF U4182 ( .A0(simTime[21]), .B0(n3533), .S(n3532), .CO(n3531));
Q_AD01HF U4183 ( .A0(simTime[20]), .B0(n3535), .S(n3534), .CO(n3533));
Q_AD01HF U4184 ( .A0(simTime[19]), .B0(n3537), .S(n3536), .CO(n3535));
Q_AD01HF U4185 ( .A0(simTime[18]), .B0(n3539), .S(n3538), .CO(n3537));
Q_AD01HF U4186 ( .A0(simTime[17]), .B0(n3541), .S(n3540), .CO(n3539));
Q_AD01HF U4187 ( .A0(simTime[16]), .B0(n3543), .S(n3542), .CO(n3541));
Q_AD01HF U4188 ( .A0(simTime[15]), .B0(n3545), .S(n3544), .CO(n3543));
Q_AD01HF U4189 ( .A0(simTime[14]), .B0(n3547), .S(n3546), .CO(n3545));
Q_AD01HF U4190 ( .A0(simTime[13]), .B0(n3549), .S(n3548), .CO(n3547));
Q_AD01HF U4191 ( .A0(simTime[12]), .B0(n3551), .S(n3550), .CO(n3549));
Q_AD01HF U4192 ( .A0(simTime[11]), .B0(n3553), .S(n3552), .CO(n3551));
Q_AD01HF U4193 ( .A0(simTime[10]), .B0(n3555), .S(n3554), .CO(n3553));
Q_AD01HF U4194 ( .A0(simTime[9]), .B0(n3557), .S(n3556), .CO(n3555));
Q_AD01HF U4195 ( .A0(simTime[8]), .B0(n3559), .S(n3558), .CO(n3557));
Q_AD01HF U4196 ( .A0(simTime[7]), .B0(n3561), .S(n3560), .CO(n3559));
Q_AD01HF U4197 ( .A0(simTime[6]), .B0(n3563), .S(n3562), .CO(n3561));
Q_AD01HF U4198 ( .A0(simTime[5]), .B0(n3565), .S(n3564), .CO(n3563));
Q_AD01HF U4199 ( .A0(simTime[4]), .B0(n3567), .S(n3566), .CO(n3565));
Q_AD01HF U4200 ( .A0(simTime[3]), .B0(simTime[2]), .S(n3568), .CO(n3567));
Q_AN02 U4201 ( .A0(asyncCall), .A1(acHalt), .Z(n3570));
Q_AN02 U4202 ( .A0(asyncCall), .A1(n3587), .Z(n3571));
Q_AN02 U4203 ( .A0(asyncCall), .A1(n3589), .Z(n3572));
Q_AN02 U4204 ( .A0(asyncCall), .A1(n3591), .Z(n3573));
Q_AN02 U4205 ( .A0(asyncCall), .A1(n3593), .Z(n3574));
Q_AN02 U4206 ( .A0(asyncCall), .A1(n3595), .Z(n3575));
Q_AN02 U4207 ( .A0(asyncCall), .A1(n3597), .Z(n3576));
Q_AN02 U4208 ( .A0(asyncCall), .A1(n3599), .Z(n3577));
Q_AN02 U4209 ( .A0(asyncCall), .A1(n3601), .Z(n3578));
Q_AN02 U4210 ( .A0(asyncCall), .A1(n3603), .Z(n3579));
Q_AN02 U4211 ( .A0(asyncCall), .A1(n3605), .Z(n3580));
Q_AN02 U4212 ( .A0(asyncCall), .A1(n3607), .Z(n3581));
Q_AN02 U4213 ( .A0(asyncCall), .A1(n3609), .Z(n3582));
Q_AN02 U4214 ( .A0(asyncCall), .A1(n3611), .Z(n3583));
Q_AN02 U4215 ( .A0(asyncCall), .A1(n3613), .Z(n3584));
Q_AN02 U4216 ( .A0(asyncCall), .A1(n3615), .Z(n3585));
Q_AN02 U4217 ( .A0(asyncCall), .A1(n3616), .Z(n3586));
Q_XOR2 U4218 ( .A0(aHaltCnt[15]), .A1(n3588), .Z(n3587));
Q_AD01HF U4219 ( .A0(aHaltCnt[14]), .B0(n3590), .S(n3589), .CO(n3588));
Q_AD01HF U4220 ( .A0(aHaltCnt[13]), .B0(n3592), .S(n3591), .CO(n3590));
Q_AD01HF U4221 ( .A0(aHaltCnt[12]), .B0(n3594), .S(n3593), .CO(n3592));
Q_AD01HF U4222 ( .A0(aHaltCnt[11]), .B0(n3596), .S(n3595), .CO(n3594));
Q_AD01HF U4223 ( .A0(aHaltCnt[10]), .B0(n3598), .S(n3597), .CO(n3596));
Q_AD01HF U4224 ( .A0(aHaltCnt[9]), .B0(n3600), .S(n3599), .CO(n3598));
Q_AD01HF U4225 ( .A0(aHaltCnt[8]), .B0(n3602), .S(n3601), .CO(n3600));
Q_AD01HF U4226 ( .A0(aHaltCnt[7]), .B0(n3604), .S(n3603), .CO(n3602));
Q_AD01HF U4227 ( .A0(aHaltCnt[6]), .B0(n3606), .S(n3605), .CO(n3604));
Q_AD01HF U4228 ( .A0(aHaltCnt[5]), .B0(n3608), .S(n3607), .CO(n3606));
Q_AD01HF U4229 ( .A0(aHaltCnt[4]), .B0(n3610), .S(n3609), .CO(n3608));
Q_AD01HF U4230 ( .A0(aHaltCnt[3]), .B0(n3612), .S(n3611), .CO(n3610));
Q_AD01HF U4231 ( .A0(aHaltCnt[2]), .B0(n3614), .S(n3613), .CO(n3612));
Q_AD01HF U4232 ( .A0(aHaltCnt[1]), .B0(aHaltCnt[0]), .S(n3615), .CO(n3614));
Q_INV U4233 ( .A(evalOnInt), .Z(n3618));
Q_OA21 U4234 ( .A0(n3618), .A1(bpHalt), .B0(n3617), .Z(n3619));
Q_INV U4235 ( .A(mpOn), .Z(n3617));
Q_AN02 U4236 ( .A0(n3617), .A1(n3636), .Z(n3620));
Q_AN02 U4237 ( .A0(n3617), .A1(n3638), .Z(n3621));
Q_AN02 U4238 ( .A0(n3617), .A1(n3640), .Z(n3622));
Q_AN02 U4239 ( .A0(n3617), .A1(n3642), .Z(n3623));
Q_AN02 U4240 ( .A0(n3617), .A1(n3644), .Z(n3624));
Q_AN02 U4241 ( .A0(n3617), .A1(n3646), .Z(n3625));
Q_AN02 U4242 ( .A0(n3617), .A1(n3648), .Z(n3626));
Q_AN02 U4243 ( .A0(n3617), .A1(n3650), .Z(n3627));
Q_AN02 U4244 ( .A0(n3617), .A1(n3652), .Z(n3628));
Q_AN02 U4245 ( .A0(n3617), .A1(n3654), .Z(n3629));
Q_AN02 U4246 ( .A0(n3617), .A1(n3656), .Z(n3630));
Q_AN02 U4247 ( .A0(n3617), .A1(n3658), .Z(n3631));
Q_AN02 U4248 ( .A0(n3617), .A1(n3660), .Z(n3632));
Q_AN02 U4249 ( .A0(n3617), .A1(n3662), .Z(n3633));
Q_AN02 U4250 ( .A0(n3617), .A1(n3664), .Z(n3634));
Q_NR02 U4251 ( .A0(mpOn), .A1(bHaltCnt[0]), .Z(n3635));
Q_XOR2 U4252 ( .A0(bHaltCnt[15]), .A1(n3637), .Z(n3636));
Q_AD01HF U4253 ( .A0(bHaltCnt[14]), .B0(n3639), .S(n3638), .CO(n3637));
Q_AD01HF U4254 ( .A0(bHaltCnt[13]), .B0(n3641), .S(n3640), .CO(n3639));
Q_AD01HF U4255 ( .A0(bHaltCnt[12]), .B0(n3643), .S(n3642), .CO(n3641));
Q_AD01HF U4256 ( .A0(bHaltCnt[11]), .B0(n3645), .S(n3644), .CO(n3643));
Q_AD01HF U4257 ( .A0(bHaltCnt[10]), .B0(n3647), .S(n3646), .CO(n3645));
Q_AD01HF U4258 ( .A0(bHaltCnt[9]), .B0(n3649), .S(n3648), .CO(n3647));
Q_AD01HF U4259 ( .A0(bHaltCnt[8]), .B0(n3651), .S(n3650), .CO(n3649));
Q_AD01HF U4260 ( .A0(bHaltCnt[7]), .B0(n3653), .S(n3652), .CO(n3651));
Q_AD01HF U4261 ( .A0(bHaltCnt[6]), .B0(n3655), .S(n3654), .CO(n3653));
Q_AD01HF U4262 ( .A0(bHaltCnt[5]), .B0(n3657), .S(n3656), .CO(n3655));
Q_AD01HF U4263 ( .A0(bHaltCnt[4]), .B0(n3659), .S(n3658), .CO(n3657));
Q_AD01HF U4264 ( .A0(bHaltCnt[3]), .B0(n3661), .S(n3660), .CO(n3659));
Q_AD01HF U4265 ( .A0(bHaltCnt[2]), .B0(n3663), .S(n3662), .CO(n3661));
Q_AD01HF U4266 ( .A0(bHaltCnt[1]), .B0(bHaltCnt[0]), .S(n3664), .CO(n3663));
Q_INV U4267 ( .A(uClk), .Z(n3665));
Q_OR02 U4268 ( .A0(hssReset), .A1(hotSwapOnPI), .Z(n3666));
Q_FDP0 GFReset_REG  ( .CK(uClk), .D(n3666), .Q(GFReset), .QN( ));
Q_MX02 U4270 ( .S(xc_mioOnS), .A0(oneStepPI), .A1(oneStepPImio), .Z(oneStepPIi));
Q_MX02 U4271 ( .S(xc_mioOnS), .A0(stopEmuPI), .A1(mioPIW_1[3]), .Z(stopEmuPIi));
Q_MX02 U4272 ( .S(xc_mioOnS), .A0(ckgHoldPI), .A1(ckgHoldPImio), .Z(ckgHoldPIi));
Q_MX02 U4273 ( .S(xc_mioOnS), .A0(callEmuPI), .A1(callEmuPImio), .Z(callEmuPIi));
Q_MX02 U4274 ( .S(xc_mioOnS), .A0(evalStepPI[63]), .A1(evalStepPImio[63]), .Z(evalStepPIi[63]));
Q_MX02 U4275 ( .S(xc_mioOnS), .A0(evalStepPI[62]), .A1(evalStepPImio[62]), .Z(evalStepPIi[62]));
Q_MX02 U4276 ( .S(xc_mioOnS), .A0(evalStepPI[61]), .A1(evalStepPImio[61]), .Z(evalStepPIi[61]));
Q_MX02 U4277 ( .S(xc_mioOnS), .A0(evalStepPI[60]), .A1(evalStepPImio[60]), .Z(evalStepPIi[60]));
Q_MX02 U4278 ( .S(xc_mioOnS), .A0(evalStepPI[59]), .A1(evalStepPImio[59]), .Z(evalStepPIi[59]));
Q_MX02 U4279 ( .S(xc_mioOnS), .A0(evalStepPI[58]), .A1(evalStepPImio[58]), .Z(evalStepPIi[58]));
Q_MX02 U4280 ( .S(xc_mioOnS), .A0(evalStepPI[57]), .A1(evalStepPImio[57]), .Z(evalStepPIi[57]));
Q_MX02 U4281 ( .S(xc_mioOnS), .A0(evalStepPI[56]), .A1(evalStepPImio[56]), .Z(evalStepPIi[56]));
Q_MX02 U4282 ( .S(xc_mioOnS), .A0(evalStepPI[55]), .A1(evalStepPImio[55]), .Z(evalStepPIi[55]));
Q_MX02 U4283 ( .S(xc_mioOnS), .A0(evalStepPI[54]), .A1(evalStepPImio[54]), .Z(evalStepPIi[54]));
Q_MX02 U4284 ( .S(xc_mioOnS), .A0(evalStepPI[53]), .A1(evalStepPImio[53]), .Z(evalStepPIi[53]));
Q_MX02 U4285 ( .S(xc_mioOnS), .A0(evalStepPI[52]), .A1(evalStepPImio[52]), .Z(evalStepPIi[52]));
Q_MX02 U4286 ( .S(xc_mioOnS), .A0(evalStepPI[51]), .A1(evalStepPImio[51]), .Z(evalStepPIi[51]));
Q_MX02 U4287 ( .S(xc_mioOnS), .A0(evalStepPI[50]), .A1(evalStepPImio[50]), .Z(evalStepPIi[50]));
Q_MX02 U4288 ( .S(xc_mioOnS), .A0(evalStepPI[49]), .A1(evalStepPImio[49]), .Z(evalStepPIi[49]));
Q_MX02 U4289 ( .S(xc_mioOnS), .A0(evalStepPI[48]), .A1(evalStepPImio[48]), .Z(evalStepPIi[48]));
Q_MX02 U4290 ( .S(xc_mioOnS), .A0(evalStepPI[47]), .A1(evalStepPImio[47]), .Z(evalStepPIi[47]));
Q_MX02 U4291 ( .S(xc_mioOnS), .A0(evalStepPI[46]), .A1(evalStepPImio[46]), .Z(evalStepPIi[46]));
Q_MX02 U4292 ( .S(xc_mioOnS), .A0(evalStepPI[45]), .A1(evalStepPImio[45]), .Z(evalStepPIi[45]));
Q_MX02 U4293 ( .S(xc_mioOnS), .A0(evalStepPI[44]), .A1(evalStepPImio[44]), .Z(evalStepPIi[44]));
Q_MX02 U4294 ( .S(xc_mioOnS), .A0(evalStepPI[43]), .A1(evalStepPImio[43]), .Z(evalStepPIi[43]));
Q_MX02 U4295 ( .S(xc_mioOnS), .A0(evalStepPI[42]), .A1(evalStepPImio[42]), .Z(evalStepPIi[42]));
Q_MX02 U4296 ( .S(xc_mioOnS), .A0(evalStepPI[41]), .A1(evalStepPImio[41]), .Z(evalStepPIi[41]));
Q_MX02 U4297 ( .S(xc_mioOnS), .A0(evalStepPI[40]), .A1(evalStepPImio[40]), .Z(evalStepPIi[40]));
Q_MX02 U4298 ( .S(xc_mioOnS), .A0(evalStepPI[39]), .A1(evalStepPImio[39]), .Z(evalStepPIi[39]));
Q_MX02 U4299 ( .S(xc_mioOnS), .A0(evalStepPI[38]), .A1(evalStepPImio[38]), .Z(evalStepPIi[38]));
Q_MX02 U4300 ( .S(xc_mioOnS), .A0(evalStepPI[37]), .A1(evalStepPImio[37]), .Z(evalStepPIi[37]));
Q_MX02 U4301 ( .S(xc_mioOnS), .A0(evalStepPI[36]), .A1(evalStepPImio[36]), .Z(evalStepPIi[36]));
Q_MX02 U4302 ( .S(xc_mioOnS), .A0(evalStepPI[35]), .A1(evalStepPImio[35]), .Z(evalStepPIi[35]));
Q_MX02 U4303 ( .S(xc_mioOnS), .A0(evalStepPI[34]), .A1(evalStepPImio[34]), .Z(evalStepPIi[34]));
Q_MX02 U4304 ( .S(xc_mioOnS), .A0(evalStepPI[33]), .A1(evalStepPImio[33]), .Z(evalStepPIi[33]));
Q_MX02 U4305 ( .S(xc_mioOnS), .A0(evalStepPI[32]), .A1(evalStepPImio[32]), .Z(evalStepPIi[32]));
Q_MX02 U4306 ( .S(xc_mioOnS), .A0(evalStepPI[31]), .A1(evalStepPImio[31]), .Z(evalStepPIi[31]));
Q_MX02 U4307 ( .S(xc_mioOnS), .A0(evalStepPI[30]), .A1(evalStepPImio[30]), .Z(evalStepPIi[30]));
Q_MX02 U4308 ( .S(xc_mioOnS), .A0(evalStepPI[29]), .A1(evalStepPImio[29]), .Z(evalStepPIi[29]));
Q_MX02 U4309 ( .S(xc_mioOnS), .A0(evalStepPI[28]), .A1(evalStepPImio[28]), .Z(evalStepPIi[28]));
Q_MX02 U4310 ( .S(xc_mioOnS), .A0(evalStepPI[27]), .A1(evalStepPImio[27]), .Z(evalStepPIi[27]));
Q_MX02 U4311 ( .S(xc_mioOnS), .A0(evalStepPI[26]), .A1(evalStepPImio[26]), .Z(evalStepPIi[26]));
Q_MX02 U4312 ( .S(xc_mioOnS), .A0(evalStepPI[25]), .A1(evalStepPImio[25]), .Z(evalStepPIi[25]));
Q_MX02 U4313 ( .S(xc_mioOnS), .A0(evalStepPI[24]), .A1(evalStepPImio[24]), .Z(evalStepPIi[24]));
Q_MX02 U4314 ( .S(xc_mioOnS), .A0(evalStepPI[23]), .A1(evalStepPImio[23]), .Z(evalStepPIi[23]));
Q_MX02 U4315 ( .S(xc_mioOnS), .A0(evalStepPI[22]), .A1(evalStepPImio[22]), .Z(evalStepPIi[22]));
Q_MX02 U4316 ( .S(xc_mioOnS), .A0(evalStepPI[21]), .A1(evalStepPImio[21]), .Z(evalStepPIi[21]));
Q_MX02 U4317 ( .S(xc_mioOnS), .A0(evalStepPI[20]), .A1(evalStepPImio[20]), .Z(evalStepPIi[20]));
Q_MX02 U4318 ( .S(xc_mioOnS), .A0(evalStepPI[19]), .A1(evalStepPImio[19]), .Z(evalStepPIi[19]));
Q_MX02 U4319 ( .S(xc_mioOnS), .A0(evalStepPI[18]), .A1(evalStepPImio[18]), .Z(evalStepPIi[18]));
Q_MX02 U4320 ( .S(xc_mioOnS), .A0(evalStepPI[17]), .A1(evalStepPImio[17]), .Z(evalStepPIi[17]));
Q_MX02 U4321 ( .S(xc_mioOnS), .A0(evalStepPI[16]), .A1(evalStepPImio[16]), .Z(evalStepPIi[16]));
Q_MX02 U4322 ( .S(xc_mioOnS), .A0(evalStepPI[15]), .A1(evalStepPImio[15]), .Z(evalStepPIi[15]));
Q_MX02 U4323 ( .S(xc_mioOnS), .A0(evalStepPI[14]), .A1(evalStepPImio[14]), .Z(evalStepPIi[14]));
Q_MX02 U4324 ( .S(xc_mioOnS), .A0(evalStepPI[13]), .A1(evalStepPImio[13]), .Z(evalStepPIi[13]));
Q_MX02 U4325 ( .S(xc_mioOnS), .A0(evalStepPI[12]), .A1(evalStepPImio[12]), .Z(evalStepPIi[12]));
Q_MX02 U4326 ( .S(xc_mioOnS), .A0(evalStepPI[11]), .A1(evalStepPImio[11]), .Z(evalStepPIi[11]));
Q_MX02 U4327 ( .S(xc_mioOnS), .A0(evalStepPI[10]), .A1(evalStepPImio[10]), .Z(evalStepPIi[10]));
Q_MX02 U4328 ( .S(xc_mioOnS), .A0(evalStepPI[9]), .A1(evalStepPImio[9]), .Z(evalStepPIi[9]));
Q_MX02 U4329 ( .S(xc_mioOnS), .A0(evalStepPI[8]), .A1(evalStepPImio[8]), .Z(evalStepPIi[8]));
Q_MX02 U4330 ( .S(xc_mioOnS), .A0(evalStepPI[7]), .A1(evalStepPImio[7]), .Z(evalStepPIi[7]));
Q_MX02 U4331 ( .S(xc_mioOnS), .A0(evalStepPI[6]), .A1(evalStepPImio[6]), .Z(evalStepPIi[6]));
Q_MX02 U4332 ( .S(xc_mioOnS), .A0(evalStepPI[5]), .A1(evalStepPImio[5]), .Z(evalStepPIi[5]));
Q_MX02 U4333 ( .S(xc_mioOnS), .A0(evalStepPI[4]), .A1(evalStepPImio[4]), .Z(evalStepPIi[4]));
Q_MX02 U4334 ( .S(xc_mioOnS), .A0(evalStepPI[3]), .A1(evalStepPImio[3]), .Z(evalStepPIi[3]));
Q_MX02 U4335 ( .S(xc_mioOnS), .A0(evalStepPI[2]), .A1(evalStepPImio[2]), .Z(evalStepPIi[2]));
Q_MX02 U4336 ( .S(xc_mioOnS), .A0(evalStepPI[1]), .A1(evalStepPImio[1]), .Z(evalStepPIi[1]));
Q_MX02 U4337 ( .S(xc_mioOnS), .A0(evalStepPI[0]), .A1(evalStepPImio[0]), .Z(evalStepPIi[0]));
Q_RDN U4338 ( .Z(ixcHoldClk));
Q_RDN U4339 ( .Z(ptxBusy));
Q_INV U4340 ( .A(maxBpCycle[15]), .Z(n3864));
Q_AN02 U4341 ( .A0(bHaltCnt[15]), .A1(n3864), .Z(n3863));
Q_OR02 U4342 ( .A0(bHaltCnt[15]), .A1(n3864), .Z(n3862));
Q_INV U4343 ( .A(maxBpCycle[14]), .Z(n3861));
Q_AN03 U4344 ( .A0(bHaltCnt[14]), .A1(n3861), .A2(n3862), .Z(n3853));
Q_OA21 U4345 ( .A0(bHaltCnt[14]), .A1(n3861), .B0(n3862), .Z(n3857));
Q_INV U4346 ( .A(maxBpCycle[13]), .Z(n3860));
Q_AN02 U4347 ( .A0(bHaltCnt[13]), .A1(n3860), .Z(n3859));
Q_OA21 U4348 ( .A0(bHaltCnt[13]), .A1(n3860), .B0(n3857), .Z(n3856));
Q_INV U4349 ( .A(maxBpCycle[12]), .Z(n3858));
Q_AN03 U4350 ( .A0(bHaltCnt[12]), .A1(n3858), .A2(n3856), .Z(n3855));
Q_OA21 U4351 ( .A0(bHaltCnt[12]), .A1(n3858), .B0(n3856), .Z(n3851));
Q_AO21 U4352 ( .A0(n3857), .A1(n3859), .B0(n3855), .Z(n3854));
Q_OR03 U4353 ( .A0(n3863), .A1(n3853), .A2(n3854), .Z(n3852));
Q_INV U4354 ( .A(maxBpCycle[11]), .Z(n3850));
Q_AN02 U4355 ( .A0(bHaltCnt[11]), .A1(n3850), .Z(n3849));
Q_OR02 U4356 ( .A0(bHaltCnt[11]), .A1(n3850), .Z(n3848));
Q_INV U4357 ( .A(maxBpCycle[10]), .Z(n3847));
Q_AN02 U4358 ( .A0(bHaltCnt[10]), .A1(n3847), .Z(n3846));
Q_OA21 U4359 ( .A0(bHaltCnt[10]), .A1(n3847), .B0(n3848), .Z(n3841));
Q_INV U4360 ( .A(maxBpCycle[9]), .Z(n3845));
Q_AN02 U4361 ( .A0(bHaltCnt[9]), .A1(n3845), .Z(n3844));
Q_OA21 U4362 ( .A0(bHaltCnt[9]), .A1(n3845), .B0(n3841), .Z(n3840));
Q_INV U4363 ( .A(maxBpCycle[8]), .Z(n3843));
Q_AN03 U4364 ( .A0(bHaltCnt[8]), .A1(n3843), .A2(n3840), .Z(n3839));
Q_OR02 U4365 ( .A0(bHaltCnt[8]), .A1(n3843), .Z(n3842));
Q_AO21 U4366 ( .A0(n3841), .A1(n3844), .B0(n3839), .Z(n3838));
Q_AO21 U4367 ( .A0(n3848), .A1(n3846), .B0(n3849), .Z(n3837));
Q_OA21 U4368 ( .A0(n3837), .A1(n3838), .B0(n3851), .Z(n3805));
Q_AN03 U4369 ( .A0(n3840), .A1(n3842), .A2(n3851), .Z(n3808));
Q_INV U4370 ( .A(maxBpCycle[7]), .Z(n3836));
Q_AN02 U4371 ( .A0(bHaltCnt[7]), .A1(n3836), .Z(n3835));
Q_OR02 U4372 ( .A0(bHaltCnt[7]), .A1(n3836), .Z(n3834));
Q_INV U4373 ( .A(maxBpCycle[6]), .Z(n3833));
Q_AN03 U4374 ( .A0(bHaltCnt[6]), .A1(n3833), .A2(n3834), .Z(n3825));
Q_OA21 U4375 ( .A0(bHaltCnt[6]), .A1(n3833), .B0(n3834), .Z(n3829));
Q_INV U4376 ( .A(maxBpCycle[5]), .Z(n3832));
Q_AN02 U4377 ( .A0(bHaltCnt[5]), .A1(n3832), .Z(n3831));
Q_OA21 U4378 ( .A0(bHaltCnt[5]), .A1(n3832), .B0(n3829), .Z(n3828));
Q_INV U4379 ( .A(maxBpCycle[4]), .Z(n3830));
Q_AN03 U4380 ( .A0(bHaltCnt[4]), .A1(n3830), .A2(n3828), .Z(n3827));
Q_OA21 U4381 ( .A0(bHaltCnt[4]), .A1(n3830), .B0(n3828), .Z(n3823));
Q_AO21 U4382 ( .A0(n3829), .A1(n3831), .B0(n3827), .Z(n3826));
Q_OR03 U4383 ( .A0(n3835), .A1(n3825), .A2(n3826), .Z(n3824));
Q_INV U4384 ( .A(maxBpCycle[3]), .Z(n3822));
Q_AN02 U4385 ( .A0(bHaltCnt[3]), .A1(n3822), .Z(n3821));
Q_OR02 U4386 ( .A0(bHaltCnt[3]), .A1(n3822), .Z(n3820));
Q_INV U4387 ( .A(maxBpCycle[2]), .Z(n3819));
Q_AN03 U4388 ( .A0(bHaltCnt[2]), .A1(n3819), .A2(n3820), .Z(n3810));
Q_OA21 U4389 ( .A0(bHaltCnt[2]), .A1(n3819), .B0(n3820), .Z(n3813));
Q_INV U4390 ( .A(maxBpCycle[1]), .Z(n3818));
Q_AN02 U4391 ( .A0(bHaltCnt[1]), .A1(n3818), .Z(n3817));
Q_OR02 U4392 ( .A0(bHaltCnt[1]), .A1(n3818), .Z(n3816));
Q_INV U4393 ( .A(maxBpCycle[0]), .Z(n3815));
Q_AN02 U4394 ( .A0(bHaltCnt[0]), .A1(n3815), .Z(n3814));
Q_AN03 U4395 ( .A0(n3813), .A1(n3816), .A2(n3814), .Z(n3812));
Q_AO21 U4396 ( .A0(n3813), .A1(n3817), .B0(n3812), .Z(n3811));
Q_OR03 U4397 ( .A0(n3821), .A1(n3810), .A2(n3811), .Z(n3809));
Q_AN03 U4398 ( .A0(n3808), .A1(n3823), .A2(n3809), .Z(n3807));
Q_AO21 U4399 ( .A0(n3808), .A1(n3824), .B0(n3807), .Z(n3806));
Q_OR03 U4400 ( .A0(n3852), .A1(n3805), .A2(n3806), .Z(n3804));
Q_OR03 U4401 ( .A0(maxBpCycle[15]), .A1(maxBpCycle[14]), .A2(maxBpCycle[13]), .Z(n3803));
Q_OR03 U4402 ( .A0(maxBpCycle[12]), .A1(maxBpCycle[11]), .A2(maxBpCycle[10]), .Z(n3802));
Q_OR03 U4403 ( .A0(maxBpCycle[9]), .A1(maxBpCycle[8]), .A2(maxBpCycle[7]), .Z(n3801));
Q_OR03 U4404 ( .A0(maxBpCycle[6]), .A1(maxBpCycle[5]), .A2(maxBpCycle[4]), .Z(n3800));
Q_OR03 U4405 ( .A0(maxBpCycle[3]), .A1(maxBpCycle[2]), .A2(maxBpCycle[1]), .Z(n3799));
Q_OR03 U4406 ( .A0(maxBpCycle[0]), .A1(n3803), .A2(n3802), .Z(n3798));
Q_OR03 U4407 ( .A0(n3801), .A1(n3800), .A2(n3799), .Z(n3797));
Q_OA21 U4408 ( .A0(n3798), .A1(n3797), .B0(n3804), .Z(bpHalt));
Q_INV U4409 ( .A(maxAcCycle[15]), .Z(n3796));
Q_AN02 U4410 ( .A0(aHaltCnt[15]), .A1(n3796), .Z(n3795));
Q_OR02 U4411 ( .A0(aHaltCnt[15]), .A1(n3796), .Z(n3794));
Q_INV U4412 ( .A(maxAcCycle[14]), .Z(n3793));
Q_AN03 U4413 ( .A0(aHaltCnt[14]), .A1(n3793), .A2(n3794), .Z(n3785));
Q_OA21 U4414 ( .A0(aHaltCnt[14]), .A1(n3793), .B0(n3794), .Z(n3789));
Q_INV U4415 ( .A(maxAcCycle[13]), .Z(n3792));
Q_AN02 U4416 ( .A0(aHaltCnt[13]), .A1(n3792), .Z(n3791));
Q_OA21 U4417 ( .A0(aHaltCnt[13]), .A1(n3792), .B0(n3789), .Z(n3788));
Q_INV U4418 ( .A(maxAcCycle[12]), .Z(n3790));
Q_AN03 U4419 ( .A0(aHaltCnt[12]), .A1(n3790), .A2(n3788), .Z(n3787));
Q_OA21 U4420 ( .A0(aHaltCnt[12]), .A1(n3790), .B0(n3788), .Z(n3783));
Q_AO21 U4421 ( .A0(n3789), .A1(n3791), .B0(n3787), .Z(n3786));
Q_OR03 U4422 ( .A0(n3795), .A1(n3785), .A2(n3786), .Z(n3784));
Q_INV U4423 ( .A(maxAcCycle[11]), .Z(n3782));
Q_AN02 U4424 ( .A0(aHaltCnt[11]), .A1(n3782), .Z(n3781));
Q_OR02 U4425 ( .A0(aHaltCnt[11]), .A1(n3782), .Z(n3780));
Q_INV U4426 ( .A(maxAcCycle[10]), .Z(n3779));
Q_AN02 U4427 ( .A0(aHaltCnt[10]), .A1(n3779), .Z(n3778));
Q_OA21 U4428 ( .A0(aHaltCnt[10]), .A1(n3779), .B0(n3780), .Z(n3773));
Q_INV U4429 ( .A(maxAcCycle[9]), .Z(n3777));
Q_AN02 U4430 ( .A0(aHaltCnt[9]), .A1(n3777), .Z(n3776));
Q_OA21 U4431 ( .A0(aHaltCnt[9]), .A1(n3777), .B0(n3773), .Z(n3772));
Q_INV U4432 ( .A(maxAcCycle[8]), .Z(n3775));
Q_AN03 U4433 ( .A0(aHaltCnt[8]), .A1(n3775), .A2(n3772), .Z(n3771));
Q_OR02 U4434 ( .A0(aHaltCnt[8]), .A1(n3775), .Z(n3774));
Q_AO21 U4435 ( .A0(n3773), .A1(n3776), .B0(n3771), .Z(n3770));
Q_AO21 U4436 ( .A0(n3780), .A1(n3778), .B0(n3781), .Z(n3769));
Q_OA21 U4437 ( .A0(n3769), .A1(n3770), .B0(n3783), .Z(n3737));
Q_AN03 U4438 ( .A0(n3772), .A1(n3774), .A2(n3783), .Z(n3740));
Q_INV U4439 ( .A(maxAcCycle[7]), .Z(n3768));
Q_AN02 U4440 ( .A0(aHaltCnt[7]), .A1(n3768), .Z(n3767));
Q_OR02 U4441 ( .A0(aHaltCnt[7]), .A1(n3768), .Z(n3766));
Q_INV U4442 ( .A(maxAcCycle[6]), .Z(n3765));
Q_AN03 U4443 ( .A0(aHaltCnt[6]), .A1(n3765), .A2(n3766), .Z(n3757));
Q_OA21 U4444 ( .A0(aHaltCnt[6]), .A1(n3765), .B0(n3766), .Z(n3761));
Q_INV U4445 ( .A(maxAcCycle[5]), .Z(n3764));
Q_AN02 U4446 ( .A0(aHaltCnt[5]), .A1(n3764), .Z(n3763));
Q_OA21 U4447 ( .A0(aHaltCnt[5]), .A1(n3764), .B0(n3761), .Z(n3760));
Q_INV U4448 ( .A(maxAcCycle[4]), .Z(n3762));
Q_AN03 U4449 ( .A0(aHaltCnt[4]), .A1(n3762), .A2(n3760), .Z(n3759));
Q_OA21 U4450 ( .A0(aHaltCnt[4]), .A1(n3762), .B0(n3760), .Z(n3755));
Q_AO21 U4451 ( .A0(n3761), .A1(n3763), .B0(n3759), .Z(n3758));
Q_OR03 U4452 ( .A0(n3767), .A1(n3757), .A2(n3758), .Z(n3756));
Q_INV U4453 ( .A(maxAcCycle[3]), .Z(n3754));
Q_AN02 U4454 ( .A0(aHaltCnt[3]), .A1(n3754), .Z(n3753));
Q_OR02 U4455 ( .A0(aHaltCnt[3]), .A1(n3754), .Z(n3752));
Q_INV U4456 ( .A(maxAcCycle[2]), .Z(n3751));
Q_AN03 U4457 ( .A0(aHaltCnt[2]), .A1(n3751), .A2(n3752), .Z(n3742));
Q_OA21 U4458 ( .A0(aHaltCnt[2]), .A1(n3751), .B0(n3752), .Z(n3745));
Q_INV U4459 ( .A(maxAcCycle[1]), .Z(n3750));
Q_AN02 U4460 ( .A0(aHaltCnt[1]), .A1(n3750), .Z(n3749));
Q_OR02 U4461 ( .A0(aHaltCnt[1]), .A1(n3750), .Z(n3748));
Q_INV U4462 ( .A(maxAcCycle[0]), .Z(n3747));
Q_AN02 U4463 ( .A0(aHaltCnt[0]), .A1(n3747), .Z(n3746));
Q_AN03 U4464 ( .A0(n3745), .A1(n3748), .A2(n3746), .Z(n3744));
Q_AO21 U4465 ( .A0(n3745), .A1(n3749), .B0(n3744), .Z(n3743));
Q_OR03 U4466 ( .A0(n3753), .A1(n3742), .A2(n3743), .Z(n3741));
Q_AN03 U4467 ( .A0(n3740), .A1(n3755), .A2(n3741), .Z(n3739));
Q_AO21 U4468 ( .A0(n3740), .A1(n3756), .B0(n3739), .Z(n3738));
Q_OR03 U4469 ( .A0(n3784), .A1(n3737), .A2(n3738), .Z(n3736));
Q_OR03 U4470 ( .A0(maxAcCycle[15]), .A1(maxAcCycle[14]), .A2(maxAcCycle[13]), .Z(n3735));
Q_OR03 U4471 ( .A0(maxAcCycle[12]), .A1(maxAcCycle[11]), .A2(maxAcCycle[10]), .Z(n3734));
Q_OR03 U4472 ( .A0(maxAcCycle[9]), .A1(maxAcCycle[8]), .A2(maxAcCycle[7]), .Z(n3733));
Q_OR03 U4473 ( .A0(maxAcCycle[6]), .A1(maxAcCycle[5]), .A2(maxAcCycle[4]), .Z(n3732));
Q_OR03 U4474 ( .A0(maxAcCycle[3]), .A1(maxAcCycle[2]), .A2(maxAcCycle[1]), .Z(n3731));
Q_OR03 U4475 ( .A0(maxAcCycle[0]), .A1(n3735), .A2(n3734), .Z(n3730));
Q_OR03 U4476 ( .A0(n3733), .A1(n3732), .A2(n3731), .Z(n3729));
Q_OA21 U4477 ( .A0(n3730), .A1(n3729), .B0(n3736), .Z(acHalt));
Q_XOR2 U4478 ( .A0(callEmuPIi), .A1(callEmuR), .Z(callEmuEv));
Q_OR02 U4479 ( .A0(lbrOn), .A1(hotSwapOnPI), .Z(lbrOnAll));
Q_OR02 U4480 ( .A0(GFLBfull), .A1(GFGBfullBw), .Z(GFBw));
Q_RDN U4481 ( .Z(GFAck));
Q_OR03 U4482 ( .A0(stop3), .A1(stopT), .A2(mioPOW_2[5]), .Z(n3728));
Q_OR03 U4483 ( .A0(mioPOW_2[3]), .A1(mioPOW_2[2]), .A2(n3728), .Z(stopCond));
Q_OR02 U4484 ( .A0(bClkR), .A1(bpHalt), .Z(bClkRH));
Q_OR03 U4485 ( .A0(n2599), .A1(n2613), .A2(n2612), .Z(n3727));
Q_OR02 U4486 ( .A0(n3727), .A1(n2607), .Z(n3726));
Q_OR03 U4487 ( .A0(n2569), .A1(n2606), .A2(n2605), .Z(n3725));
Q_OR02 U4488 ( .A0(n3725), .A1(n2600), .Z(n3724));
Q_ND02 U4489 ( .A0(n3726), .A1(n3724), .Z(syncEn));
Q_RDN U4490 ( .Z(svGFbusy));
Q_RDN U4491 ( .Z(otbGFbusy));
Q_RDN U4492 ( .Z(svAsyncCall));
Q_RDN U4493 ( .Z(otbAsyncCall));
Q_RDN U4494 ( .Z(ecmHoldBusy));
Q_EV_WOR qstp1 ( .A(stop1));
Q_EV_WOR qstp2 ( .A(stop2));
Q_EV_WOR qstp4 ( .A(stop4));
Q_RDN U4498 ( .Z(stop1));
Q_RDN U4499 ( .Z(stop2));
Q_RDN U4500 ( .Z(stop4));
Q_AO21 U4501 ( .A0(otbGFbusy), .A1(hasGFIFO1), .B0(svGFbusy), .Z(GFbusy));
Q_AO21 U4502 ( .A0(otbAsyncCall), .A1(syncOtbChannels), .B0(svAsyncCall), .Z(asyncCall));
Q_RDN U4503 ( .Z(isfWait));
Q_RDN U4504 ( .Z(osfWait));
Q_MPCLK uc ( .uClk(uClk));
Q_AN02 U4506 ( .A0(ixc_time.runClk), .A1(simTimeEnable), .Z(cakeCcEnable));
Q_PULSE U4507 ( .A(eClkR), .Z(eClk));
Q_BUF U4508 ( .A(_ET3_COMPILER_RESERVED_NAME_DBI_APPLY_), .Z(APPLY_PI));
Q_BUF U4509 ( .A(lbrOnAll), .Z(_ET3_COMPILER_RESERVED_NAME_LBRKER_ON_));
Q_RDN U4510 ( .Z(GFLBfull));
Q_RDN U4511 ( .Z(GFGBfull));
Q_EV_WOR_START gbf ( .A(GFGBfullBw));
Q_NR03 U4513 ( .A0(n2191), .A1(mpSt[1]), .A2(mpSt[2]), .Z(n3723));
Q_OR03 U4514 ( .A0(n2170), .A1(n3723), .A2(hotSwapOnPI), .Z(APPLY_DUTPI));
Q_MPCLK1P mc1pi ( .clk(clockMC));
Q_CLKSRC mcsi ( .clk(clockMC));
Q_OR03 U4517 ( .A0(GFbusy), .A1(GFbusyD), .A2(GFbusyD2), .Z(gfifoWait));
Q_RDN U4518 ( .Z(bpWait));
Q_RDN U4519 ( .Z(bWait));
Q_RDN U4520 ( .Z(sampleXpChg));
Q_EV_WOR qbwi ( .A(bpWait));
Q_EV_WOR qxci ( .A(sampleXpChg));
Q_PULSE U4523 ( .A(bClkRH), .Z(bClk));
Q_OR03 U4524 ( .A0(bWait), .A1(bWaitExtend), .A2(holdEcmC), .Z(n3722));
Q_OR03 U4525 ( .A0(bClkHoldD), .A1(ixcHoldClk), .A2(bClkHold), .Z(n3721));
Q_OR02 U4526 ( .A0(n3722), .A1(n3721), .Z(xpHold));
Q_EV_WOR_START bkh ( .A(bClkHoldD));
Q_EV_WOR_START hec ( .A(holdEcmC));
Q_BUF intrBuf ( .A(intr), .Z(_ET3_COMPILER_RESERVED_NAME_ORION_INTERRUPT_));
Q_RDN U4530 ( .Z(it_endBuf));
Q_OA21 U4531 ( .A0(it_capture), .A1(it_replay), .B0(it_endBuf), .Z(it_newBuf));
Q_RBUFZN  dum1 ( dummyW, n3720, n3719);
Q_RBUFZP  dum2 ( dummyW, n3718, n1);
Q_OR03 U4534 ( .A0(mioPOW_2[4]), .A1(stopTL), .A2(mioPOW_2[5]), .Z(n3716));
Q_OR03 U4535 ( .A0(mioPOW_2[3]), .A1(mioPOW_2[2]), .A2(n3716), .Z(anyStop));
Q_EV_WOR_START qsynci ( .A(syncEn));
Q_OR02 U4537 ( .A0(callEmu), .A1(simTimeEnable), .Z(ecmOn));
Q_OR03 U4538 ( .A0(svAsyncCall), .A1(otbAsyncCall), .A2(ptxBusy), .Z(ecmNotSync));
Q_RDN U4539 ( .Z(holdEcmTb));
Q_RDN U4540 ( .Z(ptxHoldEcm));
Q_OR03 U4541 ( .A0(holdEcmTb), .A1(holdEcmPtxOn), .A2(holdEcmSync), .Z(holdEcm));
Q_PULSE U4542 ( .A(clockMC), .Z(mcp));
Q_XNR2 U4543 ( .A0(ixc_time.nextDutTime[0]), .A1(n3715), .Z(mcDelta[0]));
Q_OR02 U4544 ( .A0(ixc_time.nextDutTime[0]), .A1(n3715), .Z(n3684));
Q_AD02 U4545 ( .CI(n3684), .A0(ixc_time.nextDutTime[1]), .A1(ixc_time.nextDutTime[2]), .B0(n3714), .B1(n3713), .S0(mcDelta[1]), .S1(mcDelta[2]), .CO(n3683));
Q_AD02 U4546 ( .CI(n3683), .A0(ixc_time.nextDutTime[3]), .A1(ixc_time.nextDutTime[4]), .B0(n3712), .B1(n3711), .S0(mcDelta[3]), .S1(mcDelta[4]), .CO(n3682));
Q_AD02 U4547 ( .CI(n3682), .A0(ixc_time.nextDutTime[5]), .A1(ixc_time.nextDutTime[6]), .B0(n3710), .B1(n3709), .S0(mcDelta[5]), .S1(mcDelta[6]), .CO(n3681));
Q_AD02 U4548 ( .CI(n3681), .A0(ixc_time.nextDutTime[7]), .A1(ixc_time.nextDutTime[8]), .B0(n3708), .B1(n3707), .S0(mcDelta[7]), .S1(mcDelta[8]), .CO(n3680));
Q_AD02 U4549 ( .CI(n3680), .A0(ixc_time.nextDutTime[9]), .A1(ixc_time.nextDutTime[10]), .B0(n3706), .B1(n3705), .S0(mcDelta[9]), .S1(mcDelta[10]), .CO(n3679));
Q_AD02 U4550 ( .CI(n3679), .A0(ixc_time.nextDutTime[11]), .A1(ixc_time.nextDutTime[12]), .B0(n3704), .B1(n3703), .S0(mcDelta[11]), .S1(mcDelta[12]), .CO(n3678));
Q_AD02 U4551 ( .CI(n3678), .A0(ixc_time.nextDutTime[13]), .A1(ixc_time.nextDutTime[14]), .B0(n3702), .B1(n3701), .S0(mcDelta[13]), .S1(mcDelta[14]), .CO(n3677));
Q_AD02 U4552 ( .CI(n3677), .A0(ixc_time.nextDutTime[15]), .A1(ixc_time.nextDutTime[16]), .B0(n3700), .B1(n3699), .S0(mcDelta[15]), .S1(mcDelta[16]), .CO(n3676));
Q_AD02 U4553 ( .CI(n3676), .A0(ixc_time.nextDutTime[17]), .A1(ixc_time.nextDutTime[18]), .B0(n3698), .B1(n3697), .S0(mcDelta[17]), .S1(mcDelta[18]), .CO(n3675));
Q_AD02 U4554 ( .CI(n3675), .A0(ixc_time.nextDutTime[19]), .A1(ixc_time.nextDutTime[20]), .B0(n3696), .B1(n3695), .S0(mcDelta[19]), .S1(mcDelta[20]), .CO(n3674));
Q_AD02 U4555 ( .CI(n3674), .A0(ixc_time.nextDutTime[21]), .A1(ixc_time.nextDutTime[22]), .B0(n3694), .B1(n3693), .S0(mcDelta[21]), .S1(mcDelta[22]), .CO(n3673));
Q_AD02 U4556 ( .CI(n3673), .A0(ixc_time.nextDutTime[23]), .A1(ixc_time.nextDutTime[24]), .B0(n3692), .B1(n3691), .S0(mcDelta[23]), .S1(mcDelta[24]), .CO(n3672));
Q_AD02 U4557 ( .CI(n3672), .A0(ixc_time.nextDutTime[25]), .A1(ixc_time.nextDutTime[26]), .B0(n3690), .B1(n3689), .S0(mcDelta[25]), .S1(mcDelta[26]), .CO(n3671));
Q_AD02 U4558 ( .CI(n3671), .A0(ixc_time.nextDutTime[27]), .A1(ixc_time.nextDutTime[28]), .B0(n3688), .B1(n3687), .S0(mcDelta[27]), .S1(mcDelta[28]), .CO(n3670));
Q_AD02 U4559 ( .CI(n3670), .A0(ixc_time.nextDutTime[29]), .A1(ixc_time.nextDutTime[30]), .B0(n3686), .B1(n3685), .S0(mcDelta[29]), .S1(mcDelta[30]), .CO(n3669));
Q_NOT_TOUCH _zzqnthw ( .sig());
Q_INV U4561 ( .A(xpHold), .Z(n3668));
Q_AN03 U4562 ( .A0(lastDelta), .A1(n3668), .A2(n2121), .Z(mpEnable));
Q_BUF U4563 ( .A(APPLY_DUTPI), .Z(_ET3_COMPILER_RESERVED_NAME_DUTPI_APPLY_));
Q_EV_WOR qxhi ( .A(xpHold));
Q_OR02 U4565 ( .A0(ecmNotSync), .A1(ecmNotSyncD), .Z(n3667));
Q_INV U4566 ( .A(n3667), .Z(ecmSync));
Q_FDP4EP cakeUcEnable_REG  ( .CK(n3665), .CE(simTimeEnable), .R(n3717), .D(n2504), .Q(cakeUcEnable));
Q_INV U4568 ( .A(n3619), .Z(n4773));
Q_FDP4EP \bHaltCnt_REG[15] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3620), .Q(bHaltCnt[15]));
Q_FDP4EP \bHaltCnt_REG[14] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3621), .Q(bHaltCnt[14]));
Q_FDP4EP \bHaltCnt_REG[13] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3622), .Q(bHaltCnt[13]));
Q_FDP4EP \bHaltCnt_REG[12] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3623), .Q(bHaltCnt[12]));
Q_FDP4EP \bHaltCnt_REG[11] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3624), .Q(bHaltCnt[11]));
Q_FDP4EP \bHaltCnt_REG[10] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3625), .Q(bHaltCnt[10]));
Q_FDP4EP \bHaltCnt_REG[9] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3626), .Q(bHaltCnt[9]));
Q_FDP4EP \bHaltCnt_REG[8] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3627), .Q(bHaltCnt[8]));
Q_FDP4EP \bHaltCnt_REG[7] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3628), .Q(bHaltCnt[7]));
Q_FDP4EP \bHaltCnt_REG[6] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3629), .Q(bHaltCnt[6]));
Q_FDP4EP \bHaltCnt_REG[5] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3630), .Q(bHaltCnt[5]));
Q_FDP4EP \bHaltCnt_REG[4] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3631), .Q(bHaltCnt[4]));
Q_FDP4EP \bHaltCnt_REG[3] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3632), .Q(bHaltCnt[3]));
Q_FDP4EP \bHaltCnt_REG[2] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3633), .Q(bHaltCnt[2]));
Q_FDP4EP \bHaltCnt_REG[1] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3634), .Q(bHaltCnt[1]));
Q_FDP4EP \bHaltCnt_REG[0] ( .CK(uClk), .CE(n4773), .R(n3717), .D(n3635), .Q(bHaltCnt[0]));
Q_INV U4585 ( .A(n3570), .Z(n4774));
Q_FDP4EP \aHaltCnt_REG[15] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3571), .Q(aHaltCnt[15]));
Q_FDP4EP \aHaltCnt_REG[14] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3572), .Q(aHaltCnt[14]));
Q_FDP4EP \aHaltCnt_REG[13] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3573), .Q(aHaltCnt[13]));
Q_FDP4EP \aHaltCnt_REG[12] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3574), .Q(aHaltCnt[12]));
Q_FDP4EP \aHaltCnt_REG[11] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3575), .Q(aHaltCnt[11]));
Q_FDP4EP \aHaltCnt_REG[10] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3576), .Q(aHaltCnt[10]));
Q_FDP4EP \aHaltCnt_REG[9] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3577), .Q(aHaltCnt[9]));
Q_FDP4EP \aHaltCnt_REG[8] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3578), .Q(aHaltCnt[8]));
Q_FDP4EP \aHaltCnt_REG[7] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3579), .Q(aHaltCnt[7]));
Q_FDP4EP \aHaltCnt_REG[6] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3580), .Q(aHaltCnt[6]));
Q_FDP4EP \aHaltCnt_REG[5] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3581), .Q(aHaltCnt[5]));
Q_FDP4EP \aHaltCnt_REG[4] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3582), .Q(aHaltCnt[4]));
Q_FDP4EP \aHaltCnt_REG[3] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3583), .Q(aHaltCnt[3]));
Q_FDP4EP \aHaltCnt_REG[2] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3584), .Q(aHaltCnt[2]));
Q_FDP4EP \aHaltCnt_REG[1] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3585), .Q(aHaltCnt[1]));
Q_FDP4EP \aHaltCnt_REG[0] ( .CK(uClk), .CE(n4774), .R(n3717), .D(n3586), .Q(aHaltCnt[0]));
Q_INV U4602 ( .A(aHaltCnt[0]), .Z(n3616));
Q_FDP4EP lockTraceOn_REG  ( .CK(uClk), .CE(n3430), .R(n3717), .D(n2504), .Q(lockTraceOn));
Q_INV U4604 ( .A(lockTraceOn), .Z(n3295));
Q_INV U4605 ( .A(n3438), .Z(n4775));
Q_FDP4EP \lockTraceC_REG[3] ( .CK(uClk), .CE(n4775), .R(n3717), .D(n3439), .Q(lockTraceC[3]));
Q_INV U4607 ( .A(lockTrace), .Z(n2275));
Q_FDP4EP \lockTraceC_REG[2] ( .CK(uClk), .CE(n4775), .R(n3717), .D(n3440), .Q(lockTraceC[2]));
Q_FDP4EP \lockTraceC_REG[1] ( .CK(uClk), .CE(n4775), .R(n3717), .D(n3441), .Q(lockTraceC[1]));
Q_FDP4EP \lockTraceC_REG[0] ( .CK(uClk), .CE(n4775), .R(n3717), .D(n3442), .Q(lockTraceC[0]));
Q_INV U4611 ( .A(lockTraceC[0]), .Z(n3432));
Q_FDP4EP \lockTraceTime_REG[63] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3448), .Q(lockTraceTime[63]));
Q_FDP4EP \lockTraceTime_REG[62] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3450), .Q(lockTraceTime[62]));
Q_FDP4EP \lockTraceTime_REG[61] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3452), .Q(lockTraceTime[61]));
Q_FDP4EP \lockTraceTime_REG[60] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3454), .Q(lockTraceTime[60]));
Q_FDP4EP \lockTraceTime_REG[59] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3456), .Q(lockTraceTime[59]));
Q_FDP4EP \lockTraceTime_REG[58] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3458), .Q(lockTraceTime[58]));
Q_FDP4EP \lockTraceTime_REG[57] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3460), .Q(lockTraceTime[57]));
Q_FDP4EP \lockTraceTime_REG[56] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3462), .Q(lockTraceTime[56]));
Q_FDP4EP \lockTraceTime_REG[55] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3464), .Q(lockTraceTime[55]));
Q_FDP4EP \lockTraceTime_REG[54] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3466), .Q(lockTraceTime[54]));
Q_FDP4EP \lockTraceTime_REG[53] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3468), .Q(lockTraceTime[53]));
Q_FDP4EP \lockTraceTime_REG[52] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3470), .Q(lockTraceTime[52]));
Q_FDP4EP \lockTraceTime_REG[51] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3472), .Q(lockTraceTime[51]));
Q_FDP4EP \lockTraceTime_REG[50] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3474), .Q(lockTraceTime[50]));
Q_FDP4EP \lockTraceTime_REG[49] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3476), .Q(lockTraceTime[49]));
Q_FDP4EP \lockTraceTime_REG[48] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3478), .Q(lockTraceTime[48]));
Q_FDP4EP \lockTraceTime_REG[47] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3480), .Q(lockTraceTime[47]));
Q_FDP4EP \lockTraceTime_REG[46] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3482), .Q(lockTraceTime[46]));
Q_FDP4EP \lockTraceTime_REG[45] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3484), .Q(lockTraceTime[45]));
Q_FDP4EP \lockTraceTime_REG[44] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3486), .Q(lockTraceTime[44]));
Q_FDP4EP \lockTraceTime_REG[43] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3488), .Q(lockTraceTime[43]));
Q_FDP4EP \lockTraceTime_REG[42] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3490), .Q(lockTraceTime[42]));
Q_FDP4EP \lockTraceTime_REG[41] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3492), .Q(lockTraceTime[41]));
Q_FDP4EP \lockTraceTime_REG[40] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3494), .Q(lockTraceTime[40]));
Q_FDP4EP \lockTraceTime_REG[39] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3496), .Q(lockTraceTime[39]));
Q_FDP4EP \lockTraceTime_REG[38] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3498), .Q(lockTraceTime[38]));
Q_FDP4EP \lockTraceTime_REG[37] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3500), .Q(lockTraceTime[37]));
Q_FDP4EP \lockTraceTime_REG[36] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3502), .Q(lockTraceTime[36]));
Q_FDP4EP \lockTraceTime_REG[35] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3504), .Q(lockTraceTime[35]));
Q_FDP4EP \lockTraceTime_REG[34] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3506), .Q(lockTraceTime[34]));
Q_FDP4EP \lockTraceTime_REG[33] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3508), .Q(lockTraceTime[33]));
Q_FDP4EP \lockTraceTime_REG[32] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3510), .Q(lockTraceTime[32]));
Q_FDP4EP \lockTraceTime_REG[31] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3512), .Q(lockTraceTime[31]));
Q_FDP4EP \lockTraceTime_REG[30] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3514), .Q(lockTraceTime[30]));
Q_FDP4EP \lockTraceTime_REG[29] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3516), .Q(lockTraceTime[29]));
Q_FDP4EP \lockTraceTime_REG[28] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3518), .Q(lockTraceTime[28]));
Q_FDP4EP \lockTraceTime_REG[27] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3520), .Q(lockTraceTime[27]));
Q_FDP4EP \lockTraceTime_REG[26] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3522), .Q(lockTraceTime[26]));
Q_FDP4EP \lockTraceTime_REG[25] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3524), .Q(lockTraceTime[25]));
Q_FDP4EP \lockTraceTime_REG[24] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3526), .Q(lockTraceTime[24]));
Q_FDP4EP \lockTraceTime_REG[23] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3528), .Q(lockTraceTime[23]));
Q_FDP4EP \lockTraceTime_REG[22] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3530), .Q(lockTraceTime[22]));
Q_FDP4EP \lockTraceTime_REG[21] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3532), .Q(lockTraceTime[21]));
Q_FDP4EP \lockTraceTime_REG[20] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3534), .Q(lockTraceTime[20]));
Q_FDP4EP \lockTraceTime_REG[19] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3536), .Q(lockTraceTime[19]));
Q_FDP4EP \lockTraceTime_REG[18] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3538), .Q(lockTraceTime[18]));
Q_FDP4EP \lockTraceTime_REG[17] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3540), .Q(lockTraceTime[17]));
Q_FDP4EP \lockTraceTime_REG[16] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3542), .Q(lockTraceTime[16]));
Q_FDP4EP \lockTraceTime_REG[15] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3544), .Q(lockTraceTime[15]));
Q_FDP4EP \lockTraceTime_REG[14] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3546), .Q(lockTraceTime[14]));
Q_FDP4EP \lockTraceTime_REG[13] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3548), .Q(lockTraceTime[13]));
Q_FDP4EP \lockTraceTime_REG[12] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3550), .Q(lockTraceTime[12]));
Q_FDP4EP \lockTraceTime_REG[11] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3552), .Q(lockTraceTime[11]));
Q_FDP4EP \lockTraceTime_REG[10] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3554), .Q(lockTraceTime[10]));
Q_FDP4EP \lockTraceTime_REG[9] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3556), .Q(lockTraceTime[9]));
Q_FDP4EP \lockTraceTime_REG[8] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3558), .Q(lockTraceTime[8]));
Q_FDP4EP \lockTraceTime_REG[7] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3560), .Q(lockTraceTime[7]));
Q_FDP4EP \lockTraceTime_REG[6] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3562), .Q(lockTraceTime[6]));
Q_FDP4EP \lockTraceTime_REG[5] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3564), .Q(lockTraceTime[5]));
Q_FDP4EP \lockTraceTime_REG[4] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3566), .Q(lockTraceTime[4]));
Q_FDP4EP \lockTraceTime_REG[3] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3568), .Q(lockTraceTime[3]));
Q_FDP4EP \lockTraceTime_REG[2] ( .CK(uClk), .CE(n3430), .R(n3717), .D(n3569), .Q(lockTraceTime[2]));
Q_FDP4EP \lockTraceTime_REG[1] ( .CK(uClk), .CE(n3430), .R(n3717), .D(simTime[1]), .Q(lockTraceTime[1]));
Q_FDP4EP \lockTraceTime_REG[0] ( .CK(uClk), .CE(n3430), .R(n3717), .D(simTime[0]), .Q(lockTraceTime[0]));
Q_INV U4676 ( .A(mioPOW_0[63]), .Z(n4776));
Q_FDP4EP mioPOCnt_REG  ( .CK(uClk), .CE(n3428), .R(n3717), .D(n4776), .Q(mioPOCnt));
Q_FDP4EP mioPICntd_REG  ( .CK(uClk), .CE(xc_mioOnS), .R(n3717), .D(mioPICnt), .Q(mioPICntd));
Q_FDP4EP ecmOne_REG  ( .CK(uClk), .CE(n3288), .R(n3717), .D(n2504), .Q(ecmOne));
Q_INV U4680 ( .A(bpCount[63]), .Z(n4777));
Q_FDP4EP \bpCount_REG[63] ( .CK(bClk), .CE(n3247), .R(n3717), .D(n4777), .Q(bpCount[63]));
Q_INV U4682 ( .A(ixcHoldSyncCnt[63]), .Z(n4778));
Q_FDP4EP \ixcHoldSyncCnt_REG[63] ( .CK(uClk), .CE(n2), .R(n3717), .D(n4778), .Q(ixcHoldSyncCnt[63]));
Q_FDP4EP \ixcHoldSyncCnt_REG[62] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3000), .Q(ixcHoldSyncCnt[62]));
Q_FDP4EP \ixcHoldSyncCnt_REG[61] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3002), .Q(ixcHoldSyncCnt[61]));
Q_FDP4EP \ixcHoldSyncCnt_REG[60] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3004), .Q(ixcHoldSyncCnt[60]));
Q_FDP4EP \ixcHoldSyncCnt_REG[59] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3006), .Q(ixcHoldSyncCnt[59]));
Q_FDP4EP \ixcHoldSyncCnt_REG[58] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3008), .Q(ixcHoldSyncCnt[58]));
Q_FDP4EP \ixcHoldSyncCnt_REG[57] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3010), .Q(ixcHoldSyncCnt[57]));
Q_FDP4EP \ixcHoldSyncCnt_REG[56] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3012), .Q(ixcHoldSyncCnt[56]));
Q_FDP4EP \ixcHoldSyncCnt_REG[55] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3014), .Q(ixcHoldSyncCnt[55]));
Q_FDP4EP \ixcHoldSyncCnt_REG[54] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3016), .Q(ixcHoldSyncCnt[54]));
Q_FDP4EP \ixcHoldSyncCnt_REG[53] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3018), .Q(ixcHoldSyncCnt[53]));
Q_FDP4EP \ixcHoldSyncCnt_REG[52] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3020), .Q(ixcHoldSyncCnt[52]));
Q_FDP4EP \ixcHoldSyncCnt_REG[51] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3022), .Q(ixcHoldSyncCnt[51]));
Q_FDP4EP \ixcHoldSyncCnt_REG[50] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3024), .Q(ixcHoldSyncCnt[50]));
Q_FDP4EP \ixcHoldSyncCnt_REG[49] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3026), .Q(ixcHoldSyncCnt[49]));
Q_FDP4EP \ixcHoldSyncCnt_REG[48] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3028), .Q(ixcHoldSyncCnt[48]));
Q_FDP4EP \ixcHoldSyncCnt_REG[47] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3030), .Q(ixcHoldSyncCnt[47]));
Q_FDP4EP \ixcHoldSyncCnt_REG[46] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3032), .Q(ixcHoldSyncCnt[46]));
Q_FDP4EP \ixcHoldSyncCnt_REG[45] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3034), .Q(ixcHoldSyncCnt[45]));
Q_FDP4EP \ixcHoldSyncCnt_REG[44] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3036), .Q(ixcHoldSyncCnt[44]));
Q_FDP4EP \ixcHoldSyncCnt_REG[43] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3038), .Q(ixcHoldSyncCnt[43]));
Q_FDP4EP \ixcHoldSyncCnt_REG[42] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3040), .Q(ixcHoldSyncCnt[42]));
Q_FDP4EP \ixcHoldSyncCnt_REG[41] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3042), .Q(ixcHoldSyncCnt[41]));
Q_FDP4EP \ixcHoldSyncCnt_REG[40] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3044), .Q(ixcHoldSyncCnt[40]));
Q_FDP4EP \ixcHoldSyncCnt_REG[39] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3046), .Q(ixcHoldSyncCnt[39]));
Q_FDP4EP \ixcHoldSyncCnt_REG[38] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3048), .Q(ixcHoldSyncCnt[38]));
Q_FDP4EP \ixcHoldSyncCnt_REG[37] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3050), .Q(ixcHoldSyncCnt[37]));
Q_FDP4EP \ixcHoldSyncCnt_REG[36] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3052), .Q(ixcHoldSyncCnt[36]));
Q_FDP4EP \ixcHoldSyncCnt_REG[35] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3054), .Q(ixcHoldSyncCnt[35]));
Q_FDP4EP \ixcHoldSyncCnt_REG[34] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3056), .Q(ixcHoldSyncCnt[34]));
Q_FDP4EP \ixcHoldSyncCnt_REG[33] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3058), .Q(ixcHoldSyncCnt[33]));
Q_FDP4EP \ixcHoldSyncCnt_REG[32] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3060), .Q(ixcHoldSyncCnt[32]));
Q_FDP4EP \ixcHoldSyncCnt_REG[31] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3062), .Q(ixcHoldSyncCnt[31]));
Q_FDP4EP \ixcHoldSyncCnt_REG[30] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3064), .Q(ixcHoldSyncCnt[30]));
Q_FDP4EP \ixcHoldSyncCnt_REG[29] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3066), .Q(ixcHoldSyncCnt[29]));
Q_FDP4EP \ixcHoldSyncCnt_REG[28] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3068), .Q(ixcHoldSyncCnt[28]));
Q_FDP4EP \ixcHoldSyncCnt_REG[27] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3070), .Q(ixcHoldSyncCnt[27]));
Q_FDP4EP \ixcHoldSyncCnt_REG[26] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3072), .Q(ixcHoldSyncCnt[26]));
Q_FDP4EP \ixcHoldSyncCnt_REG[25] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3074), .Q(ixcHoldSyncCnt[25]));
Q_FDP4EP \ixcHoldSyncCnt_REG[24] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3076), .Q(ixcHoldSyncCnt[24]));
Q_FDP4EP \ixcHoldSyncCnt_REG[23] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3078), .Q(ixcHoldSyncCnt[23]));
Q_FDP4EP \ixcHoldSyncCnt_REG[22] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3080), .Q(ixcHoldSyncCnt[22]));
Q_FDP4EP \ixcHoldSyncCnt_REG[21] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3082), .Q(ixcHoldSyncCnt[21]));
Q_FDP4EP \ixcHoldSyncCnt_REG[20] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3084), .Q(ixcHoldSyncCnt[20]));
Q_FDP4EP \ixcHoldSyncCnt_REG[19] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3086), .Q(ixcHoldSyncCnt[19]));
Q_FDP4EP \ixcHoldSyncCnt_REG[18] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3088), .Q(ixcHoldSyncCnt[18]));
Q_FDP4EP \ixcHoldSyncCnt_REG[17] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3090), .Q(ixcHoldSyncCnt[17]));
Q_FDP4EP \ixcHoldSyncCnt_REG[16] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3092), .Q(ixcHoldSyncCnt[16]));
Q_FDP4EP \ixcHoldSyncCnt_REG[15] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3094), .Q(ixcHoldSyncCnt[15]));
Q_FDP4EP \ixcHoldSyncCnt_REG[14] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3096), .Q(ixcHoldSyncCnt[14]));
Q_FDP4EP \ixcHoldSyncCnt_REG[13] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3098), .Q(ixcHoldSyncCnt[13]));
Q_FDP4EP \ixcHoldSyncCnt_REG[12] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3100), .Q(ixcHoldSyncCnt[12]));
Q_FDP4EP \ixcHoldSyncCnt_REG[11] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3102), .Q(ixcHoldSyncCnt[11]));
Q_FDP4EP \ixcHoldSyncCnt_REG[10] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3104), .Q(ixcHoldSyncCnt[10]));
Q_FDP4EP \ixcHoldSyncCnt_REG[9] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3106), .Q(ixcHoldSyncCnt[9]));
Q_FDP4EP \ixcHoldSyncCnt_REG[8] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3108), .Q(ixcHoldSyncCnt[8]));
Q_FDP4EP \ixcHoldSyncCnt_REG[7] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3110), .Q(ixcHoldSyncCnt[7]));
Q_FDP4EP \ixcHoldSyncCnt_REG[6] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3112), .Q(ixcHoldSyncCnt[6]));
Q_FDP4EP \ixcHoldSyncCnt_REG[5] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3114), .Q(ixcHoldSyncCnt[5]));
Q_FDP4EP \ixcHoldSyncCnt_REG[4] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3116), .Q(ixcHoldSyncCnt[4]));
Q_FDP4EP \ixcHoldSyncCnt_REG[3] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3118), .Q(ixcHoldSyncCnt[3]));
Q_FDP4EP \ixcHoldSyncCnt_REG[2] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3120), .Q(ixcHoldSyncCnt[2]));
Q_FDP4EP \ixcHoldSyncCnt_REG[1] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n3122), .Q(ixcHoldSyncCnt[1]));
Q_INV U4746 ( .A(ixcHoldSyncCnt[0]), .Z(n4779));
Q_FDP4EP \ixcHoldSyncCnt_REG[0] ( .CK(uClk), .CE(n2997), .R(n3717), .D(n4779), .Q(ixcHoldSyncCnt[0]));
Q_INV U4748 ( .A(eCount[63]), .Z(n4780));
Q_FDP4EP \eCount_REG[63] ( .CK(eClk), .CE(n2996), .R(n3717), .D(n4780), .Q(eCount[63]));
Q_INV U4750 ( .A(evfCount[63]), .Z(n4781));
Q_FDP4EP \evfCount_REG[63] ( .CK(uClk), .CE(n3), .R(n3717), .D(n4781), .Q(evfCount[63]));
Q_FDP4EP \evfCount_REG[62] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2749), .Q(evfCount[62]));
Q_FDP4EP \evfCount_REG[61] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2751), .Q(evfCount[61]));
Q_FDP4EP \evfCount_REG[60] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2753), .Q(evfCount[60]));
Q_FDP4EP \evfCount_REG[59] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2755), .Q(evfCount[59]));
Q_FDP4EP \evfCount_REG[58] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2757), .Q(evfCount[58]));
Q_FDP4EP \evfCount_REG[57] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2759), .Q(evfCount[57]));
Q_FDP4EP \evfCount_REG[56] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2761), .Q(evfCount[56]));
Q_FDP4EP \evfCount_REG[55] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2763), .Q(evfCount[55]));
Q_FDP4EP \evfCount_REG[54] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2765), .Q(evfCount[54]));
Q_FDP4EP \evfCount_REG[53] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2767), .Q(evfCount[53]));
Q_FDP4EP \evfCount_REG[52] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2769), .Q(evfCount[52]));
Q_FDP4EP \evfCount_REG[51] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2771), .Q(evfCount[51]));
Q_FDP4EP \evfCount_REG[50] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2773), .Q(evfCount[50]));
Q_FDP4EP \evfCount_REG[49] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2775), .Q(evfCount[49]));
Q_FDP4EP \evfCount_REG[48] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2777), .Q(evfCount[48]));
Q_FDP4EP \evfCount_REG[47] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2779), .Q(evfCount[47]));
Q_FDP4EP \evfCount_REG[46] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2781), .Q(evfCount[46]));
Q_FDP4EP \evfCount_REG[45] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2783), .Q(evfCount[45]));
Q_FDP4EP \evfCount_REG[44] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2785), .Q(evfCount[44]));
Q_FDP4EP \evfCount_REG[43] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2787), .Q(evfCount[43]));
Q_FDP4EP \evfCount_REG[42] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2789), .Q(evfCount[42]));
Q_FDP4EP \evfCount_REG[41] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2791), .Q(evfCount[41]));
Q_FDP4EP \evfCount_REG[40] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2793), .Q(evfCount[40]));
Q_FDP4EP \evfCount_REG[39] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2795), .Q(evfCount[39]));
Q_FDP4EP \evfCount_REG[38] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2797), .Q(evfCount[38]));
Q_FDP4EP \evfCount_REG[37] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2799), .Q(evfCount[37]));
Q_FDP4EP \evfCount_REG[36] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2801), .Q(evfCount[36]));
Q_FDP4EP \evfCount_REG[35] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2803), .Q(evfCount[35]));
Q_FDP4EP \evfCount_REG[34] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2805), .Q(evfCount[34]));
Q_FDP4EP \evfCount_REG[33] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2807), .Q(evfCount[33]));
Q_FDP4EP \evfCount_REG[32] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2809), .Q(evfCount[32]));
Q_FDP4EP \evfCount_REG[31] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2811), .Q(evfCount[31]));
Q_FDP4EP \evfCount_REG[30] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2813), .Q(evfCount[30]));
Q_FDP4EP \evfCount_REG[29] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2815), .Q(evfCount[29]));
Q_FDP4EP \evfCount_REG[28] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2817), .Q(evfCount[28]));
Q_FDP4EP \evfCount_REG[27] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2819), .Q(evfCount[27]));
Q_FDP4EP \evfCount_REG[26] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2821), .Q(evfCount[26]));
Q_FDP4EP \evfCount_REG[25] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2823), .Q(evfCount[25]));
Q_FDP4EP \evfCount_REG[24] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2825), .Q(evfCount[24]));
Q_FDP4EP \evfCount_REG[23] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2827), .Q(evfCount[23]));
Q_FDP4EP \evfCount_REG[22] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2829), .Q(evfCount[22]));
Q_FDP4EP \evfCount_REG[21] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2831), .Q(evfCount[21]));
Q_FDP4EP \evfCount_REG[20] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2833), .Q(evfCount[20]));
Q_FDP4EP \evfCount_REG[19] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2835), .Q(evfCount[19]));
Q_FDP4EP \evfCount_REG[18] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2837), .Q(evfCount[18]));
Q_FDP4EP \evfCount_REG[17] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2839), .Q(evfCount[17]));
Q_FDP4EP \evfCount_REG[16] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2841), .Q(evfCount[16]));
Q_FDP4EP \evfCount_REG[15] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2843), .Q(evfCount[15]));
Q_FDP4EP \evfCount_REG[14] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2845), .Q(evfCount[14]));
Q_FDP4EP \evfCount_REG[13] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2847), .Q(evfCount[13]));
Q_FDP4EP \evfCount_REG[12] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2849), .Q(evfCount[12]));
Q_FDP4EP \evfCount_REG[11] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2851), .Q(evfCount[11]));
Q_FDP4EP \evfCount_REG[10] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2853), .Q(evfCount[10]));
Q_FDP4EP \evfCount_REG[9] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2855), .Q(evfCount[9]));
Q_FDP4EP \evfCount_REG[8] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2857), .Q(evfCount[8]));
Q_FDP4EP \evfCount_REG[7] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2859), .Q(evfCount[7]));
Q_FDP4EP \evfCount_REG[6] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2861), .Q(evfCount[6]));
Q_FDP4EP \evfCount_REG[5] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2863), .Q(evfCount[5]));
Q_FDP4EP \evfCount_REG[4] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2865), .Q(evfCount[4]));
Q_FDP4EP \evfCount_REG[3] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2867), .Q(evfCount[3]));
Q_FDP4EP \evfCount_REG[2] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2869), .Q(evfCount[2]));
Q_FDP4EP \evfCount_REG[1] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n2871), .Q(evfCount[1]));
Q_INV U4814 ( .A(evfCount[0]), .Z(n4782));
Q_FDP4EP \evfCount_REG[0] ( .CK(uClk), .CE(n2621), .R(n3717), .D(n4782), .Q(evfCount[0]));
Q_INV U4816 ( .A(fvSCount[63]), .Z(n4783));
Q_FDP4EP \fvSCount_REG[63] ( .CK(uClk), .CE(n4), .R(n3717), .D(n4783), .Q(fvSCount[63]));
Q_FDP4EP \fvSCount_REG[62] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2625), .Q(fvSCount[62]));
Q_FDP4EP \fvSCount_REG[61] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2627), .Q(fvSCount[61]));
Q_FDP4EP \fvSCount_REG[60] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2629), .Q(fvSCount[60]));
Q_FDP4EP \fvSCount_REG[59] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2631), .Q(fvSCount[59]));
Q_FDP4EP \fvSCount_REG[58] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2633), .Q(fvSCount[58]));
Q_FDP4EP \fvSCount_REG[57] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2635), .Q(fvSCount[57]));
Q_FDP4EP \fvSCount_REG[56] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2637), .Q(fvSCount[56]));
Q_FDP4EP \fvSCount_REG[55] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2639), .Q(fvSCount[55]));
Q_FDP4EP \fvSCount_REG[54] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2641), .Q(fvSCount[54]));
Q_FDP4EP \fvSCount_REG[53] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2643), .Q(fvSCount[53]));
Q_FDP4EP \fvSCount_REG[52] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2645), .Q(fvSCount[52]));
Q_FDP4EP \fvSCount_REG[51] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2647), .Q(fvSCount[51]));
Q_FDP4EP \fvSCount_REG[50] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2649), .Q(fvSCount[50]));
Q_FDP4EP \fvSCount_REG[49] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2651), .Q(fvSCount[49]));
Q_FDP4EP \fvSCount_REG[48] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2653), .Q(fvSCount[48]));
Q_FDP4EP \fvSCount_REG[47] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2655), .Q(fvSCount[47]));
Q_FDP4EP \fvSCount_REG[46] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2657), .Q(fvSCount[46]));
Q_FDP4EP \fvSCount_REG[45] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2659), .Q(fvSCount[45]));
Q_FDP4EP \fvSCount_REG[44] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2661), .Q(fvSCount[44]));
Q_FDP4EP \fvSCount_REG[43] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2663), .Q(fvSCount[43]));
Q_FDP4EP \fvSCount_REG[42] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2665), .Q(fvSCount[42]));
Q_FDP4EP \fvSCount_REG[41] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2667), .Q(fvSCount[41]));
Q_FDP4EP \fvSCount_REG[40] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2669), .Q(fvSCount[40]));
Q_FDP4EP \fvSCount_REG[39] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2671), .Q(fvSCount[39]));
Q_FDP4EP \fvSCount_REG[38] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2673), .Q(fvSCount[38]));
Q_FDP4EP \fvSCount_REG[37] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2675), .Q(fvSCount[37]));
Q_FDP4EP \fvSCount_REG[36] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2677), .Q(fvSCount[36]));
Q_FDP4EP \fvSCount_REG[35] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2679), .Q(fvSCount[35]));
Q_FDP4EP \fvSCount_REG[34] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2681), .Q(fvSCount[34]));
Q_FDP4EP \fvSCount_REG[33] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2683), .Q(fvSCount[33]));
Q_FDP4EP \fvSCount_REG[32] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2685), .Q(fvSCount[32]));
Q_FDP4EP \fvSCount_REG[31] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2687), .Q(fvSCount[31]));
Q_FDP4EP \fvSCount_REG[30] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2689), .Q(fvSCount[30]));
Q_FDP4EP \fvSCount_REG[29] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2691), .Q(fvSCount[29]));
Q_FDP4EP \fvSCount_REG[28] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2693), .Q(fvSCount[28]));
Q_FDP4EP \fvSCount_REG[27] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2695), .Q(fvSCount[27]));
Q_FDP4EP \fvSCount_REG[26] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2697), .Q(fvSCount[26]));
Q_FDP4EP \fvSCount_REG[25] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2699), .Q(fvSCount[25]));
Q_FDP4EP \fvSCount_REG[24] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2701), .Q(fvSCount[24]));
Q_FDP4EP \fvSCount_REG[23] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2703), .Q(fvSCount[23]));
Q_FDP4EP \fvSCount_REG[22] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2705), .Q(fvSCount[22]));
Q_FDP4EP \fvSCount_REG[21] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2707), .Q(fvSCount[21]));
Q_FDP4EP \fvSCount_REG[20] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2709), .Q(fvSCount[20]));
Q_FDP4EP \fvSCount_REG[19] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2711), .Q(fvSCount[19]));
Q_FDP4EP \fvSCount_REG[18] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2713), .Q(fvSCount[18]));
Q_FDP4EP \fvSCount_REG[17] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2715), .Q(fvSCount[17]));
Q_FDP4EP \fvSCount_REG[16] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2717), .Q(fvSCount[16]));
Q_FDP4EP \fvSCount_REG[15] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2719), .Q(fvSCount[15]));
Q_FDP4EP \fvSCount_REG[14] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2721), .Q(fvSCount[14]));
Q_FDP4EP \fvSCount_REG[13] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2723), .Q(fvSCount[13]));
Q_FDP4EP \fvSCount_REG[12] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2725), .Q(fvSCount[12]));
Q_FDP4EP \fvSCount_REG[11] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2727), .Q(fvSCount[11]));
Q_FDP4EP \fvSCount_REG[10] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2729), .Q(fvSCount[10]));
Q_FDP4EP \fvSCount_REG[9] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2731), .Q(fvSCount[9]));
Q_FDP4EP \fvSCount_REG[8] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2733), .Q(fvSCount[8]));
Q_FDP4EP \fvSCount_REG[7] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2735), .Q(fvSCount[7]));
Q_FDP4EP \fvSCount_REG[6] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2737), .Q(fvSCount[6]));
Q_FDP4EP \fvSCount_REG[5] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2739), .Q(fvSCount[5]));
Q_FDP4EP \fvSCount_REG[4] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2741), .Q(fvSCount[4]));
Q_FDP4EP \fvSCount_REG[3] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2743), .Q(fvSCount[3]));
Q_FDP4EP \fvSCount_REG[2] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2745), .Q(fvSCount[2]));
Q_FDP4EP \fvSCount_REG[1] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n2747), .Q(fvSCount[1]));
Q_INV U4880 ( .A(fvSCount[0]), .Z(n4784));
Q_FDP4EP \fvSCount_REG[0] ( .CK(uClk), .CE(evalOn), .R(n3717), .D(n4784), .Q(fvSCount[0]));
Q_FDP4EP \Fck2Sync_REG[15] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2508), .Q(Fck2Sync[15]));
Q_FDP4EP \Fck2Sync_REG[14] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2509), .Q(Fck2Sync[14]));
Q_FDP4EP \Fck2Sync_REG[13] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2510), .Q(Fck2Sync[13]));
Q_FDP4EP \Fck2Sync_REG[12] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2511), .Q(Fck2Sync[12]));
Q_FDP4EP \Fck2Sync_REG[11] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2512), .Q(Fck2Sync[11]));
Q_FDP4EP \Fck2Sync_REG[10] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2513), .Q(Fck2Sync[10]));
Q_FDP4EP \Fck2Sync_REG[9] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2514), .Q(Fck2Sync[9]));
Q_FDP4EP \Fck2Sync_REG[8] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2515), .Q(Fck2Sync[8]));
Q_FDP4EP \Fck2Sync_REG[7] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2516), .Q(Fck2Sync[7]));
Q_FDP4EP \Fck2Sync_REG[6] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2517), .Q(Fck2Sync[6]));
Q_FDP4EP \Fck2Sync_REG[5] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2518), .Q(Fck2Sync[5]));
Q_FDP4EP \Fck2Sync_REG[4] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2519), .Q(Fck2Sync[4]));
Q_FDP4EP \Fck2Sync_REG[3] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2520), .Q(Fck2Sync[3]));
Q_FDP4EP \Fck2Sync_REG[2] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2521), .Q(Fck2Sync[2]));
Q_FDP4EP \Fck2Sync_REG[1] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2522), .Q(Fck2Sync[1]));
Q_FDP4EP \Fck2Sync_REG[0] ( .CK(uClk), .CE(n2506), .R(n3717), .D(n2523), .Q(Fck2Sync[0]));
Q_INV U4898 ( .A(Fck2Sync[0]), .Z(n2599));
Q_FDP4EP \Gfifo2Sync_REG[15] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2524), .Q(Gfifo2Sync[15]));
Q_FDP4EP \Gfifo2Sync_REG[14] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2525), .Q(Gfifo2Sync[14]));
Q_FDP4EP \Gfifo2Sync_REG[13] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2526), .Q(Gfifo2Sync[13]));
Q_FDP4EP \Gfifo2Sync_REG[12] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2527), .Q(Gfifo2Sync[12]));
Q_FDP4EP \Gfifo2Sync_REG[11] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2528), .Q(Gfifo2Sync[11]));
Q_FDP4EP \Gfifo2Sync_REG[10] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2529), .Q(Gfifo2Sync[10]));
Q_FDP4EP \Gfifo2Sync_REG[9] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2530), .Q(Gfifo2Sync[9]));
Q_FDP4EP \Gfifo2Sync_REG[8] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2531), .Q(Gfifo2Sync[8]));
Q_FDP4EP \Gfifo2Sync_REG[7] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2532), .Q(Gfifo2Sync[7]));
Q_FDP4EP \Gfifo2Sync_REG[6] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2533), .Q(Gfifo2Sync[6]));
Q_FDP4EP \Gfifo2Sync_REG[5] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2534), .Q(Gfifo2Sync[5]));
Q_FDP4EP \Gfifo2Sync_REG[4] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2535), .Q(Gfifo2Sync[4]));
Q_FDP4EP \Gfifo2Sync_REG[3] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2536), .Q(Gfifo2Sync[3]));
Q_FDP4EP \Gfifo2Sync_REG[2] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2537), .Q(Gfifo2Sync[2]));
Q_FDP4EP \Gfifo2Sync_REG[1] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2538), .Q(Gfifo2Sync[1]));
Q_FDP4EP \Gfifo2Sync_REG[0] ( .CK(uClk), .CE(n2505), .R(n3717), .D(n2539), .Q(Gfifo2Sync[0]));
Q_INV U4915 ( .A(Gfifo2Sync[0]), .Z(n2569));
Q_FDP4EP bWaitExtend_REG  ( .CK(uClk), .CE(n2416), .R(n3717), .D(n2434), .Q(bWaitExtend));
Q_FDP4EP \dccFrameFill_REG[7] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2425), .Q(dccFrameFill[7]));
Q_FDP4EP \dccFrameFill_REG[6] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2426), .Q(dccFrameFill[6]));
Q_FDP4EP \dccFrameFill_REG[5] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2427), .Q(dccFrameFill[5]));
Q_FDP4EP \dccFrameFill_REG[4] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2428), .Q(dccFrameFill[4]));
Q_FDP4EP \dccFrameFill_REG[3] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2429), .Q(dccFrameFill[3]));
Q_FDP4EP \dccFrameFill_REG[2] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2430), .Q(dccFrameFill[2]));
Q_FDP4EP \dccFrameFill_REG[1] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2431), .Q(dccFrameFill[1]));
Q_FDP4EP \dccFrameFill_REG[0] ( .CK(uClk), .CE(n2417), .R(n3717), .D(n2432), .Q(dccFrameFill[0]));
Q_INV U4925 ( .A(n2423), .Z(n4785));
Q_FDP4EP dccState_REG  ( .CK(uClk), .CE(n4785), .R(n3717), .D(lbrOn), .Q(dccState));
Q_INV U4927 ( .A(dccState), .Z(n2433));
Q_INV U4928 ( .A(uClkCntr[0]), .Z(n4786));
Q_FDP4EP \uClkCntr_REG[0] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n4786), .Q(uClkCntr[0]));
Q_FDP4EP \uClkCntr_REG[1] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2291), .Q(uClkCntr[1]));
Q_FDP4EP \uClkCntr_REG[2] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2293), .Q(uClkCntr[2]));
Q_FDP4EP \uClkCntr_REG[3] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2295), .Q(uClkCntr[3]));
Q_FDP4EP \uClkCntr_REG[4] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2297), .Q(uClkCntr[4]));
Q_FDP4EP \uClkCntr_REG[5] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2299), .Q(uClkCntr[5]));
Q_FDP4EP \uClkCntr_REG[6] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2301), .Q(uClkCntr[6]));
Q_FDP4EP \uClkCntr_REG[7] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2303), .Q(uClkCntr[7]));
Q_FDP4EP \uClkCntr_REG[8] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2305), .Q(uClkCntr[8]));
Q_FDP4EP \uClkCntr_REG[9] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2307), .Q(uClkCntr[9]));
Q_FDP4EP \uClkCntr_REG[10] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2309), .Q(uClkCntr[10]));
Q_FDP4EP \uClkCntr_REG[11] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2311), .Q(uClkCntr[11]));
Q_FDP4EP \uClkCntr_REG[12] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2313), .Q(uClkCntr[12]));
Q_FDP4EP \uClkCntr_REG[13] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2315), .Q(uClkCntr[13]));
Q_FDP4EP \uClkCntr_REG[14] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2317), .Q(uClkCntr[14]));
Q_FDP4EP \uClkCntr_REG[15] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2319), .Q(uClkCntr[15]));
Q_FDP4EP \uClkCntr_REG[16] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2321), .Q(uClkCntr[16]));
Q_FDP4EP \uClkCntr_REG[17] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2323), .Q(uClkCntr[17]));
Q_FDP4EP \uClkCntr_REG[18] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2325), .Q(uClkCntr[18]));
Q_FDP4EP \uClkCntr_REG[19] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2327), .Q(uClkCntr[19]));
Q_FDP4EP \uClkCntr_REG[20] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2329), .Q(uClkCntr[20]));
Q_FDP4EP \uClkCntr_REG[21] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2331), .Q(uClkCntr[21]));
Q_FDP4EP \uClkCntr_REG[22] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2333), .Q(uClkCntr[22]));
Q_FDP4EP \uClkCntr_REG[23] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2335), .Q(uClkCntr[23]));
Q_FDP4EP \uClkCntr_REG[24] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2337), .Q(uClkCntr[24]));
Q_FDP4EP \uClkCntr_REG[25] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2339), .Q(uClkCntr[25]));
Q_FDP4EP \uClkCntr_REG[26] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2341), .Q(uClkCntr[26]));
Q_FDP4EP \uClkCntr_REG[27] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2343), .Q(uClkCntr[27]));
Q_FDP4EP \uClkCntr_REG[28] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2345), .Q(uClkCntr[28]));
Q_FDP4EP \uClkCntr_REG[29] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2347), .Q(uClkCntr[29]));
Q_FDP4EP \uClkCntr_REG[30] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2349), .Q(uClkCntr[30]));
Q_FDP4EP \uClkCntr_REG[31] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2351), .Q(uClkCntr[31]));
Q_FDP4EP \uClkCntr_REG[32] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2353), .Q(uClkCntr[32]));
Q_FDP4EP \uClkCntr_REG[33] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2355), .Q(uClkCntr[33]));
Q_FDP4EP \uClkCntr_REG[34] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2357), .Q(uClkCntr[34]));
Q_FDP4EP \uClkCntr_REG[35] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2359), .Q(uClkCntr[35]));
Q_FDP4EP \uClkCntr_REG[36] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2361), .Q(uClkCntr[36]));
Q_FDP4EP \uClkCntr_REG[37] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2363), .Q(uClkCntr[37]));
Q_FDP4EP \uClkCntr_REG[38] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2365), .Q(uClkCntr[38]));
Q_FDP4EP \uClkCntr_REG[39] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2367), .Q(uClkCntr[39]));
Q_FDP4EP \uClkCntr_REG[40] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2369), .Q(uClkCntr[40]));
Q_FDP4EP \uClkCntr_REG[41] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2371), .Q(uClkCntr[41]));
Q_FDP4EP \uClkCntr_REG[42] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2373), .Q(uClkCntr[42]));
Q_FDP4EP \uClkCntr_REG[43] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2375), .Q(uClkCntr[43]));
Q_FDP4EP \uClkCntr_REG[44] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2377), .Q(uClkCntr[44]));
Q_FDP4EP \uClkCntr_REG[45] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2379), .Q(uClkCntr[45]));
Q_FDP4EP \uClkCntr_REG[46] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2381), .Q(uClkCntr[46]));
Q_FDP4EP \uClkCntr_REG[47] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2383), .Q(uClkCntr[47]));
Q_FDP4EP \uClkCntr_REG[48] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2385), .Q(uClkCntr[48]));
Q_FDP4EP \uClkCntr_REG[49] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2387), .Q(uClkCntr[49]));
Q_FDP4EP \uClkCntr_REG[50] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2389), .Q(uClkCntr[50]));
Q_FDP4EP \uClkCntr_REG[51] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2391), .Q(uClkCntr[51]));
Q_FDP4EP \uClkCntr_REG[52] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2393), .Q(uClkCntr[52]));
Q_FDP4EP \uClkCntr_REG[53] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2395), .Q(uClkCntr[53]));
Q_FDP4EP \uClkCntr_REG[54] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2397), .Q(uClkCntr[54]));
Q_FDP4EP \uClkCntr_REG[55] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2399), .Q(uClkCntr[55]));
Q_FDP4EP \uClkCntr_REG[56] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2401), .Q(uClkCntr[56]));
Q_FDP4EP \uClkCntr_REG[57] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2403), .Q(uClkCntr[57]));
Q_FDP4EP \uClkCntr_REG[58] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2405), .Q(uClkCntr[58]));
Q_FDP4EP \uClkCntr_REG[59] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2407), .Q(uClkCntr[59]));
Q_FDP4EP \uClkCntr_REG[60] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2409), .Q(uClkCntr[60]));
Q_FDP4EP \uClkCntr_REG[61] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2411), .Q(uClkCntr[61]));
Q_FDP4EP \uClkCntr_REG[62] ( .CK(uClk), .CE(initClock), .R(n3717), .D(n2413), .Q(uClkCntr[62]));
Q_INV U4992 ( .A(uClkCntr[63]), .Z(n4787));
Q_FDP4EP \uClkCntr_REG[63] ( .CK(uClk), .CE(n5), .R(n3717), .D(n4787), .Q(uClkCntr[63]));
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE "xc_top"
// pragma CVASTRPROP MODULE HDLICE HDL_TEMPLATE_LIB "IXCOM_TEMP_LIBRARY"
// pragma CVASTRPROP MODULE HDLICE PROP_IXCOM_MOD TRUE
// pragma CVASTRPROP MODULE HDLICE PROP_RANOFF TRUE
// pragma CVASTRPROP MODULE HDLICE ALWAYS_ON TRUE
endmodule
