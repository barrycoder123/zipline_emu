
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_xcm118 ( clk, rst_n, wr_stb, reg_addr, cmnd_op, 
	cmnd_addr, cmnd_table_id, stat_code, stat_datawords, stat_addr, 
	stat_table_id, capability_lst, capability_type, enable, .addr_limit( {
	\addr_limit[0][8] , \addr_limit[0][7] , \addr_limit[0][6] , 
	\addr_limit[0][5] , \addr_limit[0][4] , \addr_limit[0][3] , 
	\addr_limit[0][2] , \addr_limit[0][1] , \addr_limit[0][0] } ), 
	wr_dat, rd_dat, sw_cs, sw_ce, sw_we, sw_add, sw_wdat, sw_rdat, 
	sw_match, sw_aindex, grant, yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [8:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [8:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][8] ;
input \addr_limit[0][7] ;
input \addr_limit[0][6] ;
input \addr_limit[0][5] ;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [95:0] wr_dat;
output [95:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [8:0] sw_add;
output [95:0] sw_wdat;
input [95:0] sw_rdat;
input sw_match;
input [7:0] sw_aindex;
input grant;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:8] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:95] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:8] _zy_simnet_sw_add_11_w$;
wire [0:95] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [8:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [5:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [8:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(n1), .Z(stat_datawords[0]));
Q_BUF U1 ( .A(n2), .Z(stat_datawords[1]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U5 ( .A(n1), .Z(capability_type[0]));
Q_BUF U6 ( .A(n1), .Z(capability_type[1]));
Q_BUF U7 ( .A(n1), .Z(capability_type[2]));
Q_BUF U8 ( .A(n1), .Z(capability_type[3]));
Q_BUF U9 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[2]));
Q_BUF U12 ( .A(n2), .Z(capability_lst[3]));
Q_BUF U13 ( .A(n2), .Z(capability_lst[4]));
Q_BUF U14 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[6]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U17 ( .A(n2), .Z(capability_lst[8]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U23 ( .A(n2), .Z(capability_lst[14]));
Q_BUF U24 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U25 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_or_ini_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_96 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:95], sw_wdat[95:0]);
ixc_assign_9 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:8], sw_add[8:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_96 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:95], rd_dat[95:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n1, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n2, 
	n1, n1, n1, n1, n1, n2, n1, n2, n2, n2, n2, n2, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_9 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:8], stat_addr[8:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n2, n1});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_9 _zz_strnp_6 ( stat_addr[8:0], maxaddr[8:0]);
Q_AN02 U46 ( .A0(n36), .A1(grant), .Z(igrant));
Q_AN02 U47 ( .A0(cmnd_issued), .A1(n35), .Z(badaddr));
Q_OR03 U48 ( .A0(n16), .A1(n34), .A2(n33), .Z(n35));
Q_AN02 U49 ( .A0(n17), .A1(n29), .Z(n34));
Q_AN02 U50 ( .A0(n17), .A1(n30), .Z(n32));
Q_AN03 U51 ( .A0(cmnd_addr[0]), .A1(n31), .A2(n32), .Z(n33));
Q_INV U52 ( .A(maxaddr[0]), .Z(n31));
Q_OR03 U53 ( .A0(n26), .A1(n25), .A2(n28), .Z(n29));
Q_OA21 U54 ( .A0(cmnd_addr[1]), .A1(n22), .B0(n24), .Z(n30));
Q_AN03 U55 ( .A0(cmnd_addr[1]), .A1(n22), .A2(n24), .Z(n25));
Q_INV U56 ( .A(maxaddr[1]), .Z(n22));
Q_OA21 U57 ( .A0(cmnd_addr[2]), .A1(n21), .B0(n23), .Z(n24));
Q_AN03 U58 ( .A0(cmnd_addr[2]), .A1(n21), .A2(n23), .Z(n26));
Q_INV U59 ( .A(maxaddr[2]), .Z(n21));
Q_OA21 U60 ( .A0(cmnd_addr[3]), .A1(n20), .B0(n19), .Z(n23));
Q_AN03 U61 ( .A0(cmnd_addr[3]), .A1(n20), .A2(n19), .Z(n27));
Q_INV U62 ( .A(maxaddr[3]), .Z(n20));
Q_OR02 U63 ( .A0(cmnd_addr[4]), .A1(n18), .Z(n19));
Q_AO21 U64 ( .A0(cmnd_addr[4]), .A1(n18), .B0(n27), .Z(n28));
Q_INV U65 ( .A(maxaddr[4]), .Z(n18));
Q_OR03 U66 ( .A0(n13), .A1(n12), .A2(n15), .Z(n16));
Q_OA21 U67 ( .A0(cmnd_addr[5]), .A1(n9), .B0(n11), .Z(n17));
Q_AN03 U68 ( .A0(cmnd_addr[5]), .A1(n9), .A2(n11), .Z(n12));
Q_INV U69 ( .A(maxaddr[5]), .Z(n9));
Q_OA21 U70 ( .A0(cmnd_addr[6]), .A1(n8), .B0(n10), .Z(n11));
Q_AN03 U71 ( .A0(cmnd_addr[6]), .A1(n8), .A2(n10), .Z(n13));
Q_INV U72 ( .A(maxaddr[6]), .Z(n8));
Q_OA21 U73 ( .A0(cmnd_addr[7]), .A1(n7), .B0(n6), .Z(n10));
Q_AN03 U74 ( .A0(cmnd_addr[7]), .A1(n7), .A2(n6), .Z(n14));
Q_INV U75 ( .A(maxaddr[7]), .Z(n7));
Q_OR02 U76 ( .A0(cmnd_addr[8]), .A1(n5), .Z(n6));
Q_AO21 U77 ( .A0(cmnd_addr[8]), .A1(n5), .B0(n14), .Z(n15));
Q_INV U78 ( .A(maxaddr[8]), .Z(n5));
Q_AN02 U79 ( .A0(n3), .A1(n4), .Z(timeout));
Q_AN03 U80 ( .A0(timer_r[2]), .A1(timer_r[1]), .A2(timer_r[0]), .Z(n4));
Q_AN03 U81 ( .A0(timer_r[5]), .A1(timer_r[4]), .A2(timer_r[3]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timer_r[5]);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U86 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U87 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U88 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U89 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U90 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_MX02 U91 ( .S(rst_or_ini_r), .A0(cmnd_addr[5]), .A1(rst_addr_r[5]), .Z(sw_add[5]));
Q_MX02 U92 ( .S(rst_or_ini_r), .A0(cmnd_addr[6]), .A1(rst_addr_r[6]), .Z(sw_add[6]));
Q_MX02 U93 ( .S(rst_or_ini_r), .A0(cmnd_addr[7]), .A1(rst_addr_r[7]), .Z(sw_add[7]));
Q_MX02 U94 ( .S(rst_or_ini_r), .A0(cmnd_addr[8]), .A1(rst_addr_r[8]), .Z(sw_add[8]));
Q_AN02 U95 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U96 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U97 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U98 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U99 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_AN02 U100 ( .A0(enable), .A1(\addr_limit[0][5] ), .Z(maxaddr[5]));
Q_AN02 U101 ( .A0(enable), .A1(\addr_limit[0][6] ), .Z(maxaddr[6]));
Q_AN02 U102 ( .A0(enable), .A1(\addr_limit[0][7] ), .Z(maxaddr[7]));
Q_AN02 U103 ( .A0(enable), .A1(\addr_limit[0][8] ), .Z(maxaddr[8]));
Q_INV U104 ( .A(reg_addr[4]), .Z(n37));
Q_INV U105 ( .A(reg_addr[5]), .Z(n38));
Q_INV U106 ( .A(reg_addr[7]), .Z(n39));
Q_OR03 U107 ( .A0(reg_addr[10]), .A1(reg_addr[9]), .A2(reg_addr[8]), .Z(n40));
Q_OR03 U108 ( .A0(n39), .A1(reg_addr[6]), .A2(n38), .Z(n41));
Q_OR03 U109 ( .A0(n37), .A1(reg_addr[3]), .A2(reg_addr[2]), .Z(n42));
Q_OR03 U110 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n40), .Z(n43));
Q_NR03 U111 ( .A0(n41), .A1(n42), .A2(n43), .Z(n44));
Q_AN02 U112 ( .A0(wr_stb), .A1(n44), .Z(n68));
Q_INV U113 ( .A(n63), .Z(cmnd_issued));
Q_INV U114 ( .A(unsupported_op), .Z(n62));
Q_OA21 U115 ( .A0(n46), .A1(n47), .B0(n45), .Z(unsupported_op));
Q_AN02 U116 ( .A0(n45), .A1(n48), .Z(ack_error));
Q_AO21 U117 ( .A0(n50), .A1(n51), .B0(n49), .Z(n63));
Q_INV U118 ( .A(n68), .Z(n49));
Q_MX02 U119 ( .S(cmnd[3]), .A0(n54), .A1(n52), .Z(n50));
Q_INV U120 ( .A(cmnd_cmp_stb), .Z(n64));
Q_AN02 U121 ( .A0(n45), .A1(n55), .Z(cmnd_cmp_stb));
Q_AN02 U122 ( .A0(n45), .A1(n56), .Z(cmnd_tmo_stb));
Q_AN03 U123 ( .A0(n45), .A1(n51), .A2(n54), .Z(cmnd_sis_stb));
Q_AN02 U124 ( .A0(n68), .A1(cmnd[3]), .Z(n45));
Q_AN02 U125 ( .A0(n57), .A1(n48), .Z(cmnd_inc_stb));
Q_AN02 U126 ( .A0(n52), .A1(cmnd[0]), .Z(n48));
Q_AN02 U127 ( .A0(n57), .A1(n56), .Z(cmnd_ini_stb));
Q_AN02 U128 ( .A0(n52), .A1(n51), .Z(n56));
Q_AN02 U129 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n52));
Q_INV U130 ( .A(cmnd_rst_stb), .Z(n65));
Q_AN02 U131 ( .A0(n47), .A1(n58), .Z(cmnd_rst_stb));
Q_AN02 U132 ( .A0(n57), .A1(cmnd[0]), .Z(n58));
Q_AN02 U133 ( .A0(n47), .A1(n59), .Z(cmnd_dis_stb));
Q_AN02 U134 ( .A0(n57), .A1(n51), .Z(n59));
Q_AN02 U135 ( .A0(cmnd[2]), .A1(n60), .Z(n47));
Q_AN02 U136 ( .A0(n46), .A1(n58), .Z(cmnd_ena_stb));
Q_INV U137 ( .A(cmnd_wr_stb), .Z(n66));
Q_AN02 U138 ( .A0(n46), .A1(n59), .Z(cmnd_wr_stb));
Q_INV U139 ( .A(cmnd[0]), .Z(n51));
Q_AN02 U140 ( .A0(n61), .A1(cmnd[1]), .Z(n46));
Q_INV U141 ( .A(cmnd_rd_stb), .Z(n67));
Q_AN02 U142 ( .A0(n57), .A1(n55), .Z(cmnd_rd_stb));
Q_AN02 U143 ( .A0(n54), .A1(cmnd[0]), .Z(n55));
Q_NR02 U144 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n54));
Q_INV U145 ( .A(cmnd[1]), .Z(n60));
Q_INV U146 ( .A(cmnd[2]), .Z(n61));
Q_AN02 U147 ( .A0(n68), .A1(n53), .Z(n57));
Q_INV U148 ( .A(cmnd[3]), .Z(n53));
Q_OR02 U149 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n516));
Q_XNR2 U150 ( .A0(rst_addr_r[0]), .A1(maxaddr[0]), .Z(n69));
Q_XNR2 U151 ( .A0(rst_addr_r[1]), .A1(maxaddr[1]), .Z(n70));
Q_XNR2 U152 ( .A0(rst_addr_r[2]), .A1(maxaddr[2]), .Z(n71));
Q_XNR2 U153 ( .A0(rst_addr_r[3]), .A1(maxaddr[3]), .Z(n72));
Q_XNR2 U154 ( .A0(rst_addr_r[4]), .A1(maxaddr[4]), .Z(n73));
Q_XNR2 U155 ( .A0(rst_addr_r[5]), .A1(maxaddr[5]), .Z(n74));
Q_XNR2 U156 ( .A0(rst_addr_r[6]), .A1(maxaddr[6]), .Z(n75));
Q_XNR2 U157 ( .A0(rst_addr_r[7]), .A1(maxaddr[7]), .Z(n76));
Q_XNR2 U158 ( .A0(rst_addr_r[8]), .A1(maxaddr[8]), .Z(n77));
Q_AN03 U159 ( .A0(n77), .A1(n76), .A2(n75), .Z(n78));
Q_AN03 U160 ( .A0(n74), .A1(n73), .A2(n72), .Z(n79));
Q_AN03 U161 ( .A0(n71), .A1(n70), .A2(n69), .Z(n80));
Q_AN03 U162 ( .A0(n78), .A1(n79), .A2(n80), .Z(n517));
Q_XNR2 U163 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n81));
Q_XNR2 U164 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n82));
Q_XNR2 U165 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n83));
Q_XNR2 U166 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n84));
Q_XNR2 U167 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n85));
Q_XNR2 U168 ( .A0(rst_addr_r[5]), .A1(cmnd_addr[5]), .Z(n86));
Q_XNR2 U169 ( .A0(rst_addr_r[6]), .A1(cmnd_addr[6]), .Z(n87));
Q_XNR2 U170 ( .A0(rst_addr_r[7]), .A1(cmnd_addr[7]), .Z(n88));
Q_XNR2 U171 ( .A0(rst_addr_r[8]), .A1(cmnd_addr[8]), .Z(n89));
Q_AN03 U172 ( .A0(n89), .A1(n88), .A2(n87), .Z(n90));
Q_AN03 U173 ( .A0(n86), .A1(n85), .A2(n84), .Z(n91));
Q_AN03 U174 ( .A0(n83), .A1(n82), .A2(n81), .Z(n92));
Q_AN03 U175 ( .A0(n90), .A1(n91), .A2(n92), .Z(n518));
Q_AN02 U176 ( .A0(init_inc_r), .A1(igrant), .Z(n93));
Q_XOR2 U177 ( .A0(inc_r[0]), .A1(n93), .Z(n94));
Q_AD01HF U178 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n95), .CO(n96));
Q_AD01HF U179 ( .A0(rst_addr_r[1]), .B0(n96), .S(n97), .CO(n98));
Q_AD01HF U180 ( .A0(rst_addr_r[2]), .B0(n98), .S(n99), .CO(n100));
Q_AD01HF U181 ( .A0(rst_addr_r[3]), .B0(n100), .S(n101), .CO(n102));
Q_AD01HF U182 ( .A0(rst_addr_r[4]), .B0(n102), .S(n103), .CO(n104));
Q_AD01HF U183 ( .A0(rst_addr_r[5]), .B0(n104), .S(n105), .CO(n106));
Q_AD01HF U184 ( .A0(rst_addr_r[6]), .B0(n106), .S(n107), .CO(n108));
Q_AD01HF U185 ( .A0(rst_addr_r[7]), .B0(n108), .S(n109), .CO(n110));
Q_XOR2 U186 ( .A0(rst_addr_r[8]), .A1(n110), .Z(n111));
Q_AD01HF U187 ( .A0(timer_r[1]), .B0(timer_r[0]), .S(n113), .CO(n114));
Q_AD01HF U188 ( .A0(timer_r[2]), .B0(n114), .S(n115), .CO(n116));
Q_AD01HF U189 ( .A0(timer_r[3]), .B0(n116), .S(n117), .CO(n118));
Q_AD01HF U190 ( .A0(timer_r[4]), .B0(n118), .S(n119), .CO(n120));
Q_XOR2 U191 ( .A0(timer_r[5]), .A1(n120), .Z(n121));
Q_MX02 U192 ( .S(n435), .A0(n127), .A1(n123), .Z(n122));
Q_ND02 U193 ( .A0(n124), .A1(n125), .Z(n123));
Q_ND02 U194 ( .A0(n493), .A1(n399), .Z(n125));
Q_OR02 U195 ( .A0(n126), .A1(n399), .Z(n124));
Q_OR02 U196 ( .A0(n399), .A1(n495), .Z(n127));
Q_INV U197 ( .A(n128), .Z(n129));
Q_MX02 U198 ( .S(n435), .A0(n124), .A1(n130), .Z(n128));
Q_INV U199 ( .A(n131), .Z(n130));
Q_INV U200 ( .A(n132), .Z(n133));
Q_MX02 U201 ( .S(n435), .A0(n139), .A1(n134), .Z(n132));
Q_INV U202 ( .A(n135), .Z(n134));
Q_MX02 U203 ( .S(n399), .A0(n131), .A1(n136), .Z(n135));
Q_INV U204 ( .A(n137), .Z(n136));
Q_XOR2 U205 ( .A0(n493), .A1(n138), .Z(n131));
Q_OR02 U206 ( .A0(n494), .A1(n126), .Z(n139));
Q_OR02 U207 ( .A0(n493), .A1(n495), .Z(n126));
Q_NR02 U208 ( .A0(n496), .A1(n141), .Z(n140));
Q_MX02 U209 ( .S(n399), .A0(n137), .A1(n495), .Z(n141));
Q_OR02 U210 ( .A0(n493), .A1(n138), .Z(n137));
Q_INV U211 ( .A(n495), .Z(n138));
Q_AN03 U212 ( .A0(n494), .A1(n493), .A2(n496), .Z(n142));
Q_AO21 U213 ( .A0(n142), .A1(state_r[3]), .B0(n140), .Z(n522));
Q_AO21 U214 ( .A0(n142), .A1(state_r[2]), .B0(n133), .Z(n521));
Q_AO21 U215 ( .A0(n142), .A1(state_r[1]), .B0(n129), .Z(n520));
Q_AO21 U216 ( .A0(n142), .A1(state_r[0]), .B0(n122), .Z(n519));
Q_AN02 U217 ( .A0(n497), .A1(n112), .Z(n143));
Q_AN02 U218 ( .A0(n497), .A1(n113), .Z(n144));
Q_AN02 U219 ( .A0(n497), .A1(n115), .Z(n145));
Q_AN02 U220 ( .A0(n497), .A1(n117), .Z(n146));
Q_AN02 U221 ( .A0(n497), .A1(n119), .Z(n147));
Q_AN02 U222 ( .A0(n497), .A1(n121), .Z(n148));
Q_AN02 U223 ( .A0(n499), .A1(cmnd_addr[0]), .Z(n149));
Q_MX02 U224 ( .S(n500), .A0(n149), .A1(n95), .Z(n150));
Q_AN02 U225 ( .A0(n499), .A1(cmnd_addr[1]), .Z(n151));
Q_MX02 U226 ( .S(n500), .A0(n151), .A1(n97), .Z(n152));
Q_AN02 U227 ( .A0(n499), .A1(cmnd_addr[2]), .Z(n153));
Q_MX02 U228 ( .S(n500), .A0(n153), .A1(n99), .Z(n154));
Q_AN02 U229 ( .A0(n499), .A1(cmnd_addr[3]), .Z(n155));
Q_MX02 U230 ( .S(n500), .A0(n155), .A1(n101), .Z(n156));
Q_AN02 U231 ( .A0(n499), .A1(cmnd_addr[4]), .Z(n157));
Q_MX02 U232 ( .S(n500), .A0(n157), .A1(n103), .Z(n158));
Q_AN02 U233 ( .A0(n499), .A1(cmnd_addr[5]), .Z(n159));
Q_MX02 U234 ( .S(n500), .A0(n159), .A1(n105), .Z(n160));
Q_AN02 U235 ( .A0(n499), .A1(cmnd_addr[6]), .Z(n161));
Q_MX02 U236 ( .S(n500), .A0(n161), .A1(n107), .Z(n162));
Q_AN02 U237 ( .A0(n499), .A1(cmnd_addr[7]), .Z(n163));
Q_MX02 U238 ( .S(n500), .A0(n163), .A1(n109), .Z(n164));
Q_AN02 U239 ( .A0(n499), .A1(cmnd_addr[8]), .Z(n165));
Q_MX02 U240 ( .S(n500), .A0(n165), .A1(n111), .Z(n166));
Q_AN02 U241 ( .A0(n505), .A1(n94), .Z(n167));
Q_MX03 U242 ( .S0(n507), .S1(n508), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n168));
Q_MX03 U243 ( .S0(n507), .S1(n508), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n169));
Q_MX03 U244 ( .S0(n507), .S1(n508), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n170));
Q_MX03 U245 ( .S0(n507), .S1(n508), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n171));
Q_MX03 U246 ( .S0(n507), .S1(n508), .A0(sw_aindex[4]), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n172));
Q_MX03 U247 ( .S0(n507), .S1(n508), .A0(sw_aindex[5]), .A1(wr_dat[5]), .A2(sw_rdat[5]), .Z(n173));
Q_MX03 U248 ( .S0(n507), .S1(n508), .A0(sw_aindex[6]), .A1(wr_dat[6]), .A2(sw_rdat[6]), .Z(n174));
Q_MX03 U249 ( .S0(n507), .S1(n508), .A0(sw_aindex[7]), .A1(wr_dat[7]), .A2(sw_rdat[7]), .Z(n175));
Q_MX03 U250 ( .S0(n507), .S1(n508), .A0(sw_match), .A1(wr_dat[8]), .A2(sw_rdat[8]), .Z(n176));
Q_AN02 U251 ( .A0(n507), .A1(wr_dat[9]), .Z(n177));
Q_MX02 U252 ( .S(n508), .A0(n177), .A1(sw_rdat[9]), .Z(n178));
Q_AN02 U253 ( .A0(n507), .A1(wr_dat[10]), .Z(n179));
Q_MX02 U254 ( .S(n508), .A0(n179), .A1(sw_rdat[10]), .Z(n180));
Q_AN02 U255 ( .A0(n507), .A1(wr_dat[11]), .Z(n181));
Q_MX02 U256 ( .S(n508), .A0(n181), .A1(sw_rdat[11]), .Z(n182));
Q_AN02 U257 ( .A0(n507), .A1(wr_dat[12]), .Z(n183));
Q_MX02 U258 ( .S(n508), .A0(n183), .A1(sw_rdat[12]), .Z(n184));
Q_AN02 U259 ( .A0(n507), .A1(wr_dat[13]), .Z(n185));
Q_MX02 U260 ( .S(n508), .A0(n185), .A1(sw_rdat[13]), .Z(n186));
Q_AN02 U261 ( .A0(n507), .A1(wr_dat[14]), .Z(n187));
Q_MX02 U262 ( .S(n508), .A0(n187), .A1(sw_rdat[14]), .Z(n188));
Q_AN02 U263 ( .A0(n507), .A1(wr_dat[15]), .Z(n189));
Q_MX02 U264 ( .S(n508), .A0(n189), .A1(sw_rdat[15]), .Z(n190));
Q_AN02 U265 ( .A0(n507), .A1(wr_dat[16]), .Z(n191));
Q_MX02 U266 ( .S(n508), .A0(n191), .A1(sw_rdat[16]), .Z(n192));
Q_AN02 U267 ( .A0(n507), .A1(wr_dat[17]), .Z(n193));
Q_MX02 U268 ( .S(n508), .A0(n193), .A1(sw_rdat[17]), .Z(n194));
Q_AN02 U269 ( .A0(n507), .A1(wr_dat[18]), .Z(n195));
Q_MX02 U270 ( .S(n508), .A0(n195), .A1(sw_rdat[18]), .Z(n196));
Q_AN02 U271 ( .A0(n507), .A1(wr_dat[19]), .Z(n197));
Q_MX02 U272 ( .S(n508), .A0(n197), .A1(sw_rdat[19]), .Z(n198));
Q_AN02 U273 ( .A0(n507), .A1(wr_dat[20]), .Z(n199));
Q_MX02 U274 ( .S(n508), .A0(n199), .A1(sw_rdat[20]), .Z(n200));
Q_AN02 U275 ( .A0(n507), .A1(wr_dat[21]), .Z(n201));
Q_MX02 U276 ( .S(n508), .A0(n201), .A1(sw_rdat[21]), .Z(n202));
Q_AN02 U277 ( .A0(n507), .A1(wr_dat[22]), .Z(n203));
Q_MX02 U278 ( .S(n508), .A0(n203), .A1(sw_rdat[22]), .Z(n204));
Q_AN02 U279 ( .A0(n507), .A1(wr_dat[23]), .Z(n205));
Q_MX02 U280 ( .S(n508), .A0(n205), .A1(sw_rdat[23]), .Z(n206));
Q_AN02 U281 ( .A0(n507), .A1(wr_dat[24]), .Z(n207));
Q_MX02 U282 ( .S(n508), .A0(n207), .A1(sw_rdat[24]), .Z(n208));
Q_AN02 U283 ( .A0(n507), .A1(wr_dat[25]), .Z(n209));
Q_MX02 U284 ( .S(n508), .A0(n209), .A1(sw_rdat[25]), .Z(n210));
Q_AN02 U285 ( .A0(n507), .A1(wr_dat[26]), .Z(n211));
Q_MX02 U286 ( .S(n508), .A0(n211), .A1(sw_rdat[26]), .Z(n212));
Q_AN02 U287 ( .A0(n507), .A1(wr_dat[27]), .Z(n213));
Q_MX02 U288 ( .S(n508), .A0(n213), .A1(sw_rdat[27]), .Z(n214));
Q_AN02 U289 ( .A0(n507), .A1(wr_dat[28]), .Z(n215));
Q_MX02 U290 ( .S(n508), .A0(n215), .A1(sw_rdat[28]), .Z(n216));
Q_AN02 U291 ( .A0(n507), .A1(wr_dat[29]), .Z(n217));
Q_MX02 U292 ( .S(n508), .A0(n217), .A1(sw_rdat[29]), .Z(n218));
Q_AN02 U293 ( .A0(n507), .A1(wr_dat[30]), .Z(n219));
Q_MX02 U294 ( .S(n508), .A0(n219), .A1(sw_rdat[30]), .Z(n220));
Q_AN02 U295 ( .A0(n507), .A1(wr_dat[31]), .Z(n221));
Q_MX02 U296 ( .S(n508), .A0(n221), .A1(sw_rdat[31]), .Z(n222));
Q_AN02 U297 ( .A0(n507), .A1(wr_dat[32]), .Z(n223));
Q_MX02 U298 ( .S(n508), .A0(n223), .A1(sw_rdat[32]), .Z(n224));
Q_AN02 U299 ( .A0(n507), .A1(wr_dat[33]), .Z(n225));
Q_MX02 U300 ( .S(n508), .A0(n225), .A1(sw_rdat[33]), .Z(n226));
Q_AN02 U301 ( .A0(n507), .A1(wr_dat[34]), .Z(n227));
Q_MX02 U302 ( .S(n508), .A0(n227), .A1(sw_rdat[34]), .Z(n228));
Q_AN02 U303 ( .A0(n507), .A1(wr_dat[35]), .Z(n229));
Q_MX02 U304 ( .S(n508), .A0(n229), .A1(sw_rdat[35]), .Z(n230));
Q_AN02 U305 ( .A0(n507), .A1(wr_dat[36]), .Z(n231));
Q_MX02 U306 ( .S(n508), .A0(n231), .A1(sw_rdat[36]), .Z(n232));
Q_AN02 U307 ( .A0(n507), .A1(wr_dat[37]), .Z(n233));
Q_MX02 U308 ( .S(n508), .A0(n233), .A1(sw_rdat[37]), .Z(n234));
Q_AN02 U309 ( .A0(n507), .A1(wr_dat[38]), .Z(n235));
Q_MX02 U310 ( .S(n508), .A0(n235), .A1(sw_rdat[38]), .Z(n236));
Q_AN02 U311 ( .A0(n507), .A1(wr_dat[39]), .Z(n237));
Q_MX02 U312 ( .S(n508), .A0(n237), .A1(sw_rdat[39]), .Z(n238));
Q_AN02 U313 ( .A0(n507), .A1(wr_dat[40]), .Z(n239));
Q_MX02 U314 ( .S(n508), .A0(n239), .A1(sw_rdat[40]), .Z(n240));
Q_AN02 U315 ( .A0(n507), .A1(wr_dat[41]), .Z(n241));
Q_MX02 U316 ( .S(n508), .A0(n241), .A1(sw_rdat[41]), .Z(n242));
Q_AN02 U317 ( .A0(n507), .A1(wr_dat[42]), .Z(n243));
Q_MX02 U318 ( .S(n508), .A0(n243), .A1(sw_rdat[42]), .Z(n244));
Q_AN02 U319 ( .A0(n507), .A1(wr_dat[43]), .Z(n245));
Q_MX02 U320 ( .S(n508), .A0(n245), .A1(sw_rdat[43]), .Z(n246));
Q_AN02 U321 ( .A0(n507), .A1(wr_dat[44]), .Z(n247));
Q_MX02 U322 ( .S(n508), .A0(n247), .A1(sw_rdat[44]), .Z(n248));
Q_AN02 U323 ( .A0(n507), .A1(wr_dat[45]), .Z(n249));
Q_MX02 U324 ( .S(n508), .A0(n249), .A1(sw_rdat[45]), .Z(n250));
Q_AN02 U325 ( .A0(n507), .A1(wr_dat[46]), .Z(n251));
Q_MX02 U326 ( .S(n508), .A0(n251), .A1(sw_rdat[46]), .Z(n252));
Q_AN02 U327 ( .A0(n507), .A1(wr_dat[47]), .Z(n253));
Q_MX02 U328 ( .S(n508), .A0(n253), .A1(sw_rdat[47]), .Z(n254));
Q_AN02 U329 ( .A0(n507), .A1(wr_dat[48]), .Z(n255));
Q_MX02 U330 ( .S(n508), .A0(n255), .A1(sw_rdat[48]), .Z(n256));
Q_AN02 U331 ( .A0(n507), .A1(wr_dat[49]), .Z(n257));
Q_MX02 U332 ( .S(n508), .A0(n257), .A1(sw_rdat[49]), .Z(n258));
Q_AN02 U333 ( .A0(n507), .A1(wr_dat[50]), .Z(n259));
Q_MX02 U334 ( .S(n508), .A0(n259), .A1(sw_rdat[50]), .Z(n260));
Q_AN02 U335 ( .A0(n507), .A1(wr_dat[51]), .Z(n261));
Q_MX02 U336 ( .S(n508), .A0(n261), .A1(sw_rdat[51]), .Z(n262));
Q_AN02 U337 ( .A0(n507), .A1(wr_dat[52]), .Z(n263));
Q_MX02 U338 ( .S(n508), .A0(n263), .A1(sw_rdat[52]), .Z(n264));
Q_AN02 U339 ( .A0(n507), .A1(wr_dat[53]), .Z(n265));
Q_MX02 U340 ( .S(n508), .A0(n265), .A1(sw_rdat[53]), .Z(n266));
Q_AN02 U341 ( .A0(n507), .A1(wr_dat[54]), .Z(n267));
Q_MX02 U342 ( .S(n508), .A0(n267), .A1(sw_rdat[54]), .Z(n268));
Q_AN02 U343 ( .A0(n507), .A1(wr_dat[55]), .Z(n269));
Q_MX02 U344 ( .S(n508), .A0(n269), .A1(sw_rdat[55]), .Z(n270));
Q_AN02 U345 ( .A0(n507), .A1(wr_dat[56]), .Z(n271));
Q_MX02 U346 ( .S(n508), .A0(n271), .A1(sw_rdat[56]), .Z(n272));
Q_AN02 U347 ( .A0(n507), .A1(wr_dat[57]), .Z(n273));
Q_MX02 U348 ( .S(n508), .A0(n273), .A1(sw_rdat[57]), .Z(n274));
Q_AN02 U349 ( .A0(n507), .A1(wr_dat[58]), .Z(n275));
Q_MX02 U350 ( .S(n508), .A0(n275), .A1(sw_rdat[58]), .Z(n276));
Q_AN02 U351 ( .A0(n507), .A1(wr_dat[59]), .Z(n277));
Q_MX02 U352 ( .S(n508), .A0(n277), .A1(sw_rdat[59]), .Z(n278));
Q_AN02 U353 ( .A0(n507), .A1(wr_dat[60]), .Z(n279));
Q_MX02 U354 ( .S(n508), .A0(n279), .A1(sw_rdat[60]), .Z(n280));
Q_AN02 U355 ( .A0(n507), .A1(wr_dat[61]), .Z(n281));
Q_MX02 U356 ( .S(n508), .A0(n281), .A1(sw_rdat[61]), .Z(n282));
Q_AN02 U357 ( .A0(n507), .A1(wr_dat[62]), .Z(n283));
Q_MX02 U358 ( .S(n508), .A0(n283), .A1(sw_rdat[62]), .Z(n284));
Q_AN02 U359 ( .A0(n507), .A1(wr_dat[63]), .Z(n285));
Q_MX02 U360 ( .S(n508), .A0(n285), .A1(sw_rdat[63]), .Z(n286));
Q_AN02 U361 ( .A0(n507), .A1(wr_dat[64]), .Z(n287));
Q_MX02 U362 ( .S(n508), .A0(n287), .A1(sw_rdat[64]), .Z(n288));
Q_AN02 U363 ( .A0(n507), .A1(wr_dat[65]), .Z(n289));
Q_MX02 U364 ( .S(n508), .A0(n289), .A1(sw_rdat[65]), .Z(n290));
Q_AN02 U365 ( .A0(n507), .A1(wr_dat[66]), .Z(n291));
Q_MX02 U366 ( .S(n508), .A0(n291), .A1(sw_rdat[66]), .Z(n292));
Q_AN02 U367 ( .A0(n507), .A1(wr_dat[67]), .Z(n293));
Q_MX02 U368 ( .S(n508), .A0(n293), .A1(sw_rdat[67]), .Z(n294));
Q_AN02 U369 ( .A0(n507), .A1(wr_dat[68]), .Z(n295));
Q_MX02 U370 ( .S(n508), .A0(n295), .A1(sw_rdat[68]), .Z(n296));
Q_AN02 U371 ( .A0(n507), .A1(wr_dat[69]), .Z(n297));
Q_MX02 U372 ( .S(n508), .A0(n297), .A1(sw_rdat[69]), .Z(n298));
Q_AN02 U373 ( .A0(n507), .A1(wr_dat[70]), .Z(n299));
Q_MX02 U374 ( .S(n508), .A0(n299), .A1(sw_rdat[70]), .Z(n300));
Q_AN02 U375 ( .A0(n507), .A1(wr_dat[71]), .Z(n301));
Q_MX02 U376 ( .S(n508), .A0(n301), .A1(sw_rdat[71]), .Z(n302));
Q_AN02 U377 ( .A0(n507), .A1(wr_dat[72]), .Z(n303));
Q_MX02 U378 ( .S(n508), .A0(n303), .A1(sw_rdat[72]), .Z(n304));
Q_AN02 U379 ( .A0(n507), .A1(wr_dat[73]), .Z(n305));
Q_MX02 U380 ( .S(n508), .A0(n305), .A1(sw_rdat[73]), .Z(n306));
Q_AN02 U381 ( .A0(n507), .A1(wr_dat[74]), .Z(n307));
Q_MX02 U382 ( .S(n508), .A0(n307), .A1(sw_rdat[74]), .Z(n308));
Q_AN02 U383 ( .A0(n507), .A1(wr_dat[75]), .Z(n309));
Q_MX02 U384 ( .S(n508), .A0(n309), .A1(sw_rdat[75]), .Z(n310));
Q_AN02 U385 ( .A0(n507), .A1(wr_dat[76]), .Z(n311));
Q_MX02 U386 ( .S(n508), .A0(n311), .A1(sw_rdat[76]), .Z(n312));
Q_AN02 U387 ( .A0(n507), .A1(wr_dat[77]), .Z(n313));
Q_MX02 U388 ( .S(n508), .A0(n313), .A1(sw_rdat[77]), .Z(n314));
Q_AN02 U389 ( .A0(n507), .A1(wr_dat[78]), .Z(n315));
Q_MX02 U390 ( .S(n508), .A0(n315), .A1(sw_rdat[78]), .Z(n316));
Q_AN02 U391 ( .A0(n507), .A1(wr_dat[79]), .Z(n317));
Q_MX02 U392 ( .S(n508), .A0(n317), .A1(sw_rdat[79]), .Z(n318));
Q_AN02 U393 ( .A0(n507), .A1(wr_dat[80]), .Z(n319));
Q_MX02 U394 ( .S(n508), .A0(n319), .A1(sw_rdat[80]), .Z(n320));
Q_AN02 U395 ( .A0(n507), .A1(wr_dat[81]), .Z(n321));
Q_MX02 U396 ( .S(n508), .A0(n321), .A1(sw_rdat[81]), .Z(n322));
Q_AN02 U397 ( .A0(n507), .A1(wr_dat[82]), .Z(n323));
Q_MX02 U398 ( .S(n508), .A0(n323), .A1(sw_rdat[82]), .Z(n324));
Q_AN02 U399 ( .A0(n507), .A1(wr_dat[83]), .Z(n325));
Q_MX02 U400 ( .S(n508), .A0(n325), .A1(sw_rdat[83]), .Z(n326));
Q_AN02 U401 ( .A0(n507), .A1(wr_dat[84]), .Z(n327));
Q_MX02 U402 ( .S(n508), .A0(n327), .A1(sw_rdat[84]), .Z(n328));
Q_AN02 U403 ( .A0(n507), .A1(wr_dat[85]), .Z(n329));
Q_MX02 U404 ( .S(n508), .A0(n329), .A1(sw_rdat[85]), .Z(n330));
Q_AN02 U405 ( .A0(n507), .A1(wr_dat[86]), .Z(n331));
Q_MX02 U406 ( .S(n508), .A0(n331), .A1(sw_rdat[86]), .Z(n332));
Q_AN02 U407 ( .A0(n507), .A1(wr_dat[87]), .Z(n333));
Q_MX02 U408 ( .S(n508), .A0(n333), .A1(sw_rdat[87]), .Z(n334));
Q_AN02 U409 ( .A0(n507), .A1(wr_dat[88]), .Z(n335));
Q_MX02 U410 ( .S(n508), .A0(n335), .A1(sw_rdat[88]), .Z(n336));
Q_AN02 U411 ( .A0(n507), .A1(wr_dat[89]), .Z(n337));
Q_MX02 U412 ( .S(n508), .A0(n337), .A1(sw_rdat[89]), .Z(n338));
Q_AN02 U413 ( .A0(n507), .A1(wr_dat[90]), .Z(n339));
Q_MX02 U414 ( .S(n508), .A0(n339), .A1(sw_rdat[90]), .Z(n340));
Q_AN02 U415 ( .A0(n507), .A1(wr_dat[91]), .Z(n341));
Q_MX02 U416 ( .S(n508), .A0(n341), .A1(sw_rdat[91]), .Z(n342));
Q_AN02 U417 ( .A0(n507), .A1(wr_dat[92]), .Z(n343));
Q_MX02 U418 ( .S(n508), .A0(n343), .A1(sw_rdat[92]), .Z(n344));
Q_AN02 U419 ( .A0(n507), .A1(wr_dat[93]), .Z(n345));
Q_MX02 U420 ( .S(n508), .A0(n345), .A1(sw_rdat[93]), .Z(n346));
Q_AN02 U421 ( .A0(n507), .A1(wr_dat[94]), .Z(n347));
Q_MX02 U422 ( .S(n508), .A0(n347), .A1(sw_rdat[94]), .Z(n348));
Q_AN02 U423 ( .A0(n507), .A1(wr_dat[95]), .Z(n349));
Q_MX02 U424 ( .S(n508), .A0(n349), .A1(sw_rdat[95]), .Z(n350));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n522), .Q(state_r[3]), .QN(n408));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n521), .Q(state_r[2]), .QN(n409));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n520), .Q(state_r[1]), .QN(n411));
Q_FDP1 \state_r_REG[0] ( .CK(clk), .R(rst_n), .D(n519), .Q(state_r[0]), .QN(n380));
Q_FDP1 \timer_r_REG[5] ( .CK(clk), .R(rst_n), .D(n148), .Q(timer_r[5]), .QN( ));
Q_FDP1 \timer_r_REG[4] ( .CK(clk), .R(rst_n), .D(n147), .Q(timer_r[4]), .QN( ));
Q_FDP1 \timer_r_REG[3] ( .CK(clk), .R(rst_n), .D(n146), .Q(timer_r[3]), .QN( ));
Q_FDP1 \timer_r_REG[2] ( .CK(clk), .R(rst_n), .D(n145), .Q(timer_r[2]), .QN( ));
Q_FDP1 \timer_r_REG[1] ( .CK(clk), .R(rst_n), .D(n144), .Q(timer_r[1]), .QN( ));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n143), .Q(timer_r[0]), .QN(n112));
Q_ND02 U435 ( .A0(n352), .A1(n353), .Z(n351));
Q_ND02 U436 ( .A0(n354), .A1(n466), .Z(n353));
Q_OR02 U437 ( .A0(n355), .A1(n510), .Z(n354));
Q_INV U438 ( .A(n509), .Z(n355));
Q_ND02 U439 ( .A0(n352), .A1(n357), .Z(n356));
Q_ND02 U440 ( .A0(n509), .A1(n466), .Z(n357));
Q_OR03 U441 ( .A0(n509), .A1(n510), .A2(n466), .Z(n352));
Q_MX02 U442 ( .S(n466), .A0(n509), .A1(n510), .Z(n358));
Q_FDP2 \stat_code_REG[2] ( .CK(clk), .S(rst_n), .D(n359), .Q(stat_code[2]), .QN( ));
Q_MX02 U444 ( .S(n481), .A0(stat_code[2]), .A1(n358), .Z(n359));
Q_FDP2 \stat_code_REG[1] ( .CK(clk), .S(rst_n), .D(n360), .Q(stat_code[1]), .QN( ));
Q_MX02 U446 ( .S(n481), .A0(stat_code[1]), .A1(n356), .Z(n360));
Q_FDP2 \stat_code_REG[0] ( .CK(clk), .S(rst_n), .D(n361), .Q(stat_code[0]), .QN( ));
Q_MX02 U448 ( .S(n481), .A0(stat_code[0]), .A1(n351), .Z(n361));
Q_FDP2 init_r_REG  ( .CK(clk), .S(rst_n), .D(n362), .Q(init_r), .QN(enable));
Q_MX02 U450 ( .S(n512), .A0(init_r), .A1(n506), .Z(n362));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n504), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n503), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n502), .Q(rst_r), .QN(n523));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n501), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n498), .Q(sw_we_r), .QN( ));
Q_OA21 U456 ( .A0(n364), .A1(n365), .B0(n363), .Z(n493));
Q_OR03 U457 ( .A0(n367), .A1(n368), .A2(n366), .Z(n365));
Q_AN03 U458 ( .A0(state_r[0]), .A1(n371), .A2(n369), .Z(n370));
Q_AN02 U459 ( .A0(n66), .A1(cmnd_rd_stb), .Z(n371));
Q_AN02 U460 ( .A0(n374), .A1(n63), .Z(n375));
Q_AN03 U461 ( .A0(n376), .A1(n375), .A2(n372), .Z(n373));
Q_AN02 U462 ( .A0(n377), .A1(state_r[0]), .Z(n376));
Q_OR03 U463 ( .A0(n373), .A1(n378), .A2(n370), .Z(n368));
Q_AN02 U464 ( .A0(n369), .A1(n379), .Z(n378));
Q_NR02 U465 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n379));
Q_OA21 U466 ( .A0(n382), .A1(n383), .B0(n381), .Z(n367));
Q_AN02 U467 ( .A0(n384), .A1(n385), .Z(n383));
Q_NR02 U468 ( .A0(state_r[0]), .A1(igrant), .Z(n385));
Q_OA21 U469 ( .A0(n388), .A1(n389), .B0(n387), .Z(n382));
Q_AN02 U470 ( .A0(n390), .A1(n386), .Z(n389));
Q_NR02 U471 ( .A0(n391), .A1(n518), .Z(n388));
Q_INV U472 ( .A(n392), .Z(n374));
Q_AN03 U473 ( .A0(cmnd_rst_stb), .A1(n369), .A2(n394), .Z(n395));
Q_OR03 U474 ( .A0(n396), .A1(n395), .A2(n393), .Z(n364));
Q_AN03 U475 ( .A0(n380), .A1(n398), .A2(n397), .Z(n396));
Q_INV U476 ( .A(n399), .Z(n494));
Q_OA21 U477 ( .A0(n400), .A1(n366), .B0(n363), .Z(n399));
Q_AO21 U478 ( .A0(n369), .A1(n403), .B0(n402), .Z(n400));
Q_AN02 U479 ( .A0(state_r[0]), .A1(cmnd_wr_stb), .Z(n403));
Q_AN03 U480 ( .A0(n407), .A1(n380), .A2(n405), .Z(n406));
Q_NR02 U481 ( .A0(state_r[3]), .A1(state_r[2]), .Z(n407));
Q_MX02 U482 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n410), .Z(n405));
Q_OR03 U483 ( .A0(n412), .A1(n406), .A2(n404), .Z(n366));
Q_AN02 U484 ( .A0(n413), .A1(n381), .Z(n404));
Q_AN02 U485 ( .A0(n377), .A1(n63), .Z(n381));
Q_AN02 U486 ( .A0(n414), .A1(n415), .Z(n412));
Q_NR02 U487 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n415));
Q_MX02 U488 ( .S(state_r[3]), .A0(n417), .A1(n416), .Z(n413));
Q_AN02 U489 ( .A0(n452), .A1(n410), .Z(n418));
Q_AN02 U490 ( .A0(ack_error), .A1(enable), .Z(n410));
Q_AO21 U491 ( .A0(n419), .A1(n380), .B0(n418), .Z(n416));
Q_AN02 U492 ( .A0(state_r[2]), .A1(igrant), .Z(n421));
Q_AO21 U493 ( .A0(n422), .A1(n423), .B0(n420), .Z(n417));
Q_OA21 U494 ( .A0(state_r[0]), .A1(n424), .B0(n421), .Z(n420));
Q_AN02 U495 ( .A0(n411), .A1(n518), .Z(n424));
Q_OR02 U496 ( .A0(state_r[2]), .A1(n392), .Z(n422));
Q_AN02 U497 ( .A0(igrant), .A1(n517), .Z(n392));
Q_OA21 U498 ( .A0(n425), .A1(n426), .B0(n401), .Z(n402));
Q_AN03 U499 ( .A0(n427), .A1(n408), .A2(n394), .Z(n426));
Q_AN02 U500 ( .A0(n428), .A1(n429), .Z(n425));
Q_AN03 U501 ( .A0(n431), .A1(n432), .A2(n430), .Z(n495));
Q_AO21 U502 ( .A0(n427), .A1(n434), .B0(n433), .Z(n430));
Q_INV U503 ( .A(n433), .Z(n434));
Q_INV U504 ( .A(n435), .Z(n496));
Q_OA21 U505 ( .A0(n436), .A1(n393), .B0(n363), .Z(n435));
Q_AN03 U506 ( .A0(n433), .A1(n432), .A2(n369), .Z(n437));
Q_AN02 U507 ( .A0(state_r[0]), .A1(n66), .Z(n432));
Q_AO21 U508 ( .A0(n67), .A1(cmnd_cmp_stb), .B0(cmnd_rd_stb), .Z(n433));
Q_AN03 U509 ( .A0(n427), .A1(n369), .A2(n394), .Z(n438));
Q_AN02 U510 ( .A0(n439), .A1(n64), .Z(n394));
Q_AO21 U511 ( .A0(n65), .A1(n516), .B0(cmnd_rst_stb), .Z(n427));
Q_AN03 U512 ( .A0(n428), .A1(n63), .A2(n397), .Z(n441));
Q_AN02 U513 ( .A0(n377), .A1(n384), .Z(n397));
Q_AN02 U514 ( .A0(state_r[3]), .A1(n401), .Z(n384));
Q_OR03 U515 ( .A0(n441), .A1(n440), .A2(n437), .Z(n436));
Q_AO21 U516 ( .A0(n442), .A1(n443), .B0(n438), .Z(n440));
Q_AN02 U517 ( .A0(igrant), .A1(n63), .Z(n398));
Q_AN02 U518 ( .A0(n444), .A1(n398), .Z(n442));
Q_NR02 U519 ( .A0(timeout), .A1(state_r[0]), .Z(n444));
Q_AN02 U520 ( .A0(ack_error), .A1(init_r), .Z(n446));
Q_AO21 U521 ( .A0(n414), .A1(cmnd_dis_stb), .B0(n445), .Z(n393));
Q_AN02 U522 ( .A0(n439), .A1(n448), .Z(n447));
Q_NR02 U523 ( .A0(cmnd_cmp_stb), .A1(n516), .Z(n448));
Q_AN02 U524 ( .A0(state_r[0]), .A1(n449), .Z(n439));
Q_NR02 U525 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n449));
Q_AN03 U526 ( .A0(n65), .A1(n369), .A2(n447), .Z(n414));
Q_OA21 U527 ( .A0(n450), .A1(n451), .B0(n446), .Z(n445));
Q_AN02 U528 ( .A0(n452), .A1(n429), .Z(n450));
Q_AN03 U529 ( .A0(n377), .A1(state_r[3]), .A2(n63), .Z(n429));
Q_INV U530 ( .A(n390), .Z(n423));
Q_AO21 U531 ( .A0(n380), .A1(igrant), .B0(state_r[0]), .Z(n428));
Q_AN02 U532 ( .A0(n386), .A1(n504), .Z(n497));
Q_INV U533 ( .A(igrant), .Z(n386));
Q_OA21 U534 ( .A0(n454), .A1(n455), .B0(n453), .Z(n498));
Q_AN02 U535 ( .A0(n521), .A1(n456), .Z(n455));
Q_AN02 U536 ( .A0(cmnd_sis_stb), .A1(n457), .Z(n499));
Q_INV U537 ( .A(n500), .Z(n457));
Q_ND02 U538 ( .A0(n390), .A1(n409), .Z(n452));
Q_OR02 U539 ( .A0(state_r[0]), .A1(state_r[1]), .Z(n391));
Q_ND02 U540 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n390));
Q_OA21 U541 ( .A0(n454), .A1(n458), .B0(n453), .Z(n501));
Q_AN02 U542 ( .A0(n521), .A1(n459), .Z(n458));
Q_AN02 U543 ( .A0(n460), .A1(n461), .Z(n454));
Q_AN02 U544 ( .A0(n462), .A1(n461), .Z(n502));
Q_OR03 U545 ( .A0(n463), .A1(n503), .A2(n502), .Z(n504));
Q_AN03 U546 ( .A0(n522), .A1(n460), .A2(n459), .Z(n503));
Q_AN03 U547 ( .A0(n453), .A1(n521), .A2(n464), .Z(n463));
Q_INV U548 ( .A(n461), .Z(n464));
Q_INV U549 ( .A(n465), .Z(n505));
Q_AN02 U550 ( .A0(n443), .A1(state_r[0]), .Z(n508));
Q_AN03 U551 ( .A0(state_r[2]), .A1(state_r[1]), .A2(n408), .Z(n443));
Q_AN02 U552 ( .A0(n468), .A1(n469), .Z(n470));
Q_INV U553 ( .A(n471), .Z(n468));
Q_OR03 U554 ( .A0(n472), .A1(n470), .A2(n467), .Z(n466));
Q_AN03 U555 ( .A0(n474), .A1(n62), .A2(n473), .Z(n467));
Q_OR02 U556 ( .A0(n461), .A1(n475), .Z(n472));
Q_AN02 U557 ( .A0(n520), .A1(n519), .Z(n461));
Q_INV U558 ( .A(n462), .Z(n475));
Q_AN02 U559 ( .A0(n462), .A1(n476), .Z(n469));
Q_OA21 U560 ( .A0(n477), .A1(n456), .B0(n469), .Z(n509));
Q_AN02 U561 ( .A0(n62), .A1(n520), .Z(n471));
Q_OA21 U562 ( .A0(n474), .A1(badaddr), .B0(n471), .Z(n477));
Q_AN02 U563 ( .A0(timeout), .A1(n363), .Z(n474));
Q_OA21 U564 ( .A0(n478), .A1(n479), .B0(n462), .Z(n510));
Q_AO21 U565 ( .A0(n456), .A1(n519), .B0(n459), .Z(n479));
Q_AN02 U566 ( .A0(unsupported_op), .A1(n480), .Z(n478));
Q_ND02 U567 ( .A0(n451), .A1(n473), .Z(n481));
Q_AN02 U568 ( .A0(n462), .A1(n480), .Z(n473));
Q_AN02 U569 ( .A0(n520), .A1(n476), .Z(n480));
Q_AN02 U570 ( .A0(n372), .A1(n380), .Z(n451));
Q_AN02 U571 ( .A0(n408), .A1(n419), .Z(n372));
Q_OA21 U572 ( .A0(n507), .A1(n482), .B0(n363), .Z(n511));
Q_AN02 U573 ( .A0(n483), .A1(state_r[1]), .Z(n482));
Q_INV U574 ( .A(n506), .Z(n507));
Q_AN02 U575 ( .A0(n408), .A1(n401), .Z(n369));
Q_MX02 U576 ( .S(state_r[0]), .A0(n484), .A1(n387), .Z(n483));
Q_AN02 U577 ( .A0(state_r[3]), .A1(n409), .Z(n484));
Q_AN02 U578 ( .A0(n408), .A1(state_r[2]), .Z(n387));
Q_AN03 U579 ( .A0(n462), .A1(n459), .A2(n506), .Z(n485));
Q_NR02 U580 ( .A0(n520), .A1(n519), .Z(n459));
Q_INV U581 ( .A(n519), .Z(n476));
Q_INV U582 ( .A(n520), .Z(n456));
Q_NR02 U583 ( .A0(n522), .A1(n521), .Z(n462));
Q_INV U584 ( .A(n521), .Z(n460));
Q_INV U585 ( .A(n522), .Z(n453));
Q_AO21 U586 ( .A0(n431), .A1(n486), .B0(n485), .Z(n512));
Q_AN02 U587 ( .A0(n380), .A1(cmnd_ena_stb), .Z(n486));
Q_OR02 U588 ( .A0(state_r[3]), .A1(state_r[1]), .Z(n487));
Q_OR03 U589 ( .A0(state_r[2]), .A1(state_r[0]), .A2(n487), .Z(n506));
Q_AN03 U590 ( .A0(n489), .A1(n411), .A2(n488), .Z(n513));
Q_AO21 U591 ( .A0(state_r[2]), .A1(n380), .B0(n465), .Z(n488));
Q_AN02 U592 ( .A0(n409), .A1(state_r[0]), .Z(n465));
Q_ND02 U593 ( .A0(n431), .A1(state_r[0]), .Z(n514));
Q_AN02 U594 ( .A0(n489), .A1(n401), .Z(n431));
Q_NR02 U595 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n401));
Q_AN02 U596 ( .A0(n490), .A1(n489), .Z(n500));
Q_NR02 U597 ( .A0(badaddr), .A1(state_r[3]), .Z(n489));
Q_INV U598 ( .A(badaddr), .Z(n363));
Q_OR03 U599 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n500), .Z(n515));
Q_MX02 U600 ( .S(state_r[0]), .A0(n491), .A1(n419), .Z(n490));
Q_AN02 U601 ( .A0(state_r[2]), .A1(n411), .Z(n491));
Q_AN02 U602 ( .A0(n409), .A1(state_r[1]), .Z(n419));
Q_OR02 U603 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n492));
Q_INV U604 ( .A(timeout), .Z(n377));
Q_AN02 U605 ( .A0(n523), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U606 ( .A0(n523), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U607 ( .A0(n523), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U608 ( .A0(n523), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U609 ( .A0(n523), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U610 ( .A0(n523), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U611 ( .A0(n523), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U612 ( .A0(n523), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U613 ( .A0(n523), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U614 ( .A0(n523), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U615 ( .A0(n523), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U616 ( .A0(n523), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U617 ( .A0(n523), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U618 ( .A0(n523), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U619 ( .A0(n523), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U620 ( .A0(n523), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U621 ( .A0(n523), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U622 ( .A0(n523), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U623 ( .A0(n523), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U624 ( .A0(n523), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U625 ( .A0(n523), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U626 ( .A0(n523), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U627 ( .A0(n523), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U628 ( .A0(n523), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U629 ( .A0(n523), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U630 ( .A0(n523), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U631 ( .A0(n523), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U632 ( .A0(n523), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U633 ( .A0(n523), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U634 ( .A0(n523), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U635 ( .A0(n523), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U636 ( .A0(n523), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_AN02 U637 ( .A0(n523), .A1(wr_dat[32]), .Z(sw_wdat[32]));
Q_AN02 U638 ( .A0(n523), .A1(wr_dat[33]), .Z(sw_wdat[33]));
Q_AN02 U639 ( .A0(n523), .A1(wr_dat[34]), .Z(sw_wdat[34]));
Q_AN02 U640 ( .A0(n523), .A1(wr_dat[35]), .Z(sw_wdat[35]));
Q_AN02 U641 ( .A0(n523), .A1(wr_dat[36]), .Z(sw_wdat[36]));
Q_AN02 U642 ( .A0(n523), .A1(wr_dat[37]), .Z(sw_wdat[37]));
Q_AN02 U643 ( .A0(n523), .A1(wr_dat[38]), .Z(sw_wdat[38]));
Q_AN02 U644 ( .A0(n523), .A1(wr_dat[39]), .Z(sw_wdat[39]));
Q_AN02 U645 ( .A0(n523), .A1(wr_dat[40]), .Z(sw_wdat[40]));
Q_AN02 U646 ( .A0(n523), .A1(wr_dat[41]), .Z(sw_wdat[41]));
Q_AN02 U647 ( .A0(n523), .A1(wr_dat[42]), .Z(sw_wdat[42]));
Q_AN02 U648 ( .A0(n523), .A1(wr_dat[43]), .Z(sw_wdat[43]));
Q_AN02 U649 ( .A0(n523), .A1(wr_dat[44]), .Z(sw_wdat[44]));
Q_AN02 U650 ( .A0(n523), .A1(wr_dat[45]), .Z(sw_wdat[45]));
Q_AN02 U651 ( .A0(n523), .A1(wr_dat[46]), .Z(sw_wdat[46]));
Q_AN02 U652 ( .A0(n523), .A1(wr_dat[47]), .Z(sw_wdat[47]));
Q_AN02 U653 ( .A0(n523), .A1(wr_dat[48]), .Z(sw_wdat[48]));
Q_AN02 U654 ( .A0(n523), .A1(wr_dat[49]), .Z(sw_wdat[49]));
Q_AN02 U655 ( .A0(n523), .A1(wr_dat[50]), .Z(sw_wdat[50]));
Q_AN02 U656 ( .A0(n523), .A1(wr_dat[51]), .Z(sw_wdat[51]));
Q_AN02 U657 ( .A0(n523), .A1(wr_dat[52]), .Z(sw_wdat[52]));
Q_AN02 U658 ( .A0(n523), .A1(wr_dat[53]), .Z(sw_wdat[53]));
Q_AN02 U659 ( .A0(n523), .A1(wr_dat[54]), .Z(sw_wdat[54]));
Q_AN02 U660 ( .A0(n523), .A1(wr_dat[55]), .Z(sw_wdat[55]));
Q_AN02 U661 ( .A0(n523), .A1(wr_dat[56]), .Z(sw_wdat[56]));
Q_AN02 U662 ( .A0(n523), .A1(wr_dat[57]), .Z(sw_wdat[57]));
Q_AN02 U663 ( .A0(n523), .A1(wr_dat[58]), .Z(sw_wdat[58]));
Q_AN02 U664 ( .A0(n523), .A1(wr_dat[59]), .Z(sw_wdat[59]));
Q_AN02 U665 ( .A0(n523), .A1(wr_dat[60]), .Z(sw_wdat[60]));
Q_AN02 U666 ( .A0(n523), .A1(wr_dat[61]), .Z(sw_wdat[61]));
Q_AN02 U667 ( .A0(n523), .A1(wr_dat[62]), .Z(sw_wdat[62]));
Q_AN02 U668 ( .A0(n523), .A1(wr_dat[63]), .Z(sw_wdat[63]));
Q_AN02 U669 ( .A0(n523), .A1(wr_dat[64]), .Z(sw_wdat[64]));
Q_AN02 U670 ( .A0(n523), .A1(wr_dat[65]), .Z(sw_wdat[65]));
Q_AN02 U671 ( .A0(n523), .A1(wr_dat[66]), .Z(sw_wdat[66]));
Q_AN02 U672 ( .A0(n523), .A1(wr_dat[67]), .Z(sw_wdat[67]));
Q_AN02 U673 ( .A0(n523), .A1(wr_dat[68]), .Z(sw_wdat[68]));
Q_AN02 U674 ( .A0(n523), .A1(wr_dat[69]), .Z(sw_wdat[69]));
Q_AN02 U675 ( .A0(n523), .A1(wr_dat[70]), .Z(sw_wdat[70]));
Q_AN02 U676 ( .A0(n523), .A1(wr_dat[71]), .Z(sw_wdat[71]));
Q_AN02 U677 ( .A0(n523), .A1(wr_dat[72]), .Z(sw_wdat[72]));
Q_AN02 U678 ( .A0(n523), .A1(wr_dat[73]), .Z(sw_wdat[73]));
Q_AN02 U679 ( .A0(n523), .A1(wr_dat[74]), .Z(sw_wdat[74]));
Q_AN02 U680 ( .A0(n523), .A1(wr_dat[75]), .Z(sw_wdat[75]));
Q_AN02 U681 ( .A0(n523), .A1(wr_dat[76]), .Z(sw_wdat[76]));
Q_AN02 U682 ( .A0(n523), .A1(wr_dat[77]), .Z(sw_wdat[77]));
Q_AN02 U683 ( .A0(n523), .A1(wr_dat[78]), .Z(sw_wdat[78]));
Q_AN02 U684 ( .A0(n523), .A1(wr_dat[79]), .Z(sw_wdat[79]));
Q_AN02 U685 ( .A0(n523), .A1(wr_dat[80]), .Z(sw_wdat[80]));
Q_AN02 U686 ( .A0(n523), .A1(wr_dat[81]), .Z(sw_wdat[81]));
Q_AN02 U687 ( .A0(n523), .A1(wr_dat[82]), .Z(sw_wdat[82]));
Q_AN02 U688 ( .A0(n523), .A1(wr_dat[83]), .Z(sw_wdat[83]));
Q_AN02 U689 ( .A0(n523), .A1(wr_dat[84]), .Z(sw_wdat[84]));
Q_AN02 U690 ( .A0(n523), .A1(wr_dat[85]), .Z(sw_wdat[85]));
Q_AN02 U691 ( .A0(n523), .A1(wr_dat[86]), .Z(sw_wdat[86]));
Q_AN02 U692 ( .A0(n523), .A1(wr_dat[87]), .Z(sw_wdat[87]));
Q_AN02 U693 ( .A0(n523), .A1(wr_dat[88]), .Z(sw_wdat[88]));
Q_AN02 U694 ( .A0(n523), .A1(wr_dat[89]), .Z(sw_wdat[89]));
Q_AN02 U695 ( .A0(n523), .A1(wr_dat[90]), .Z(sw_wdat[90]));
Q_AN02 U696 ( .A0(n523), .A1(wr_dat[91]), .Z(sw_wdat[91]));
Q_AN02 U697 ( .A0(n523), .A1(wr_dat[92]), .Z(sw_wdat[92]));
Q_AN02 U698 ( .A0(n523), .A1(wr_dat[93]), .Z(sw_wdat[93]));
Q_AN02 U699 ( .A0(n523), .A1(wr_dat[94]), .Z(sw_wdat[94]));
Q_AN02 U700 ( .A0(n523), .A1(wr_dat[95]), .Z(sw_wdat[95]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n492), .R(n524), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U702 ( .A(rst_n), .Z(n524));
Q_INV U703 ( .A(sim_tmo_r), .Z(n36));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n515), .R(n524), .D(n150), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n515), .R(n524), .D(n152), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n515), .R(n524), .D(n154), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n515), .R(n524), .D(n156), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n515), .R(n524), .D(n158), .Q(rst_addr_r[4]));
Q_FDP4EP \rst_addr_r_REG[5] ( .CK(clk), .CE(n515), .R(n524), .D(n160), .Q(rst_addr_r[5]));
Q_FDP4EP \rst_addr_r_REG[6] ( .CK(clk), .CE(n515), .R(n524), .D(n162), .Q(rst_addr_r[6]));
Q_FDP4EP \rst_addr_r_REG[7] ( .CK(clk), .CE(n515), .R(n524), .D(n164), .Q(rst_addr_r[7]));
Q_FDP4EP \rst_addr_r_REG[8] ( .CK(clk), .CE(n515), .R(n524), .D(n166), .Q(rst_addr_r[8]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n513), .R(n524), .D(n167), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n511), .R(n524), .D(n168), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n511), .R(n524), .D(n169), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n511), .R(n524), .D(n170), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n511), .R(n524), .D(n171), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n511), .R(n524), .D(n172), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n511), .R(n524), .D(n173), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n511), .R(n524), .D(n174), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n511), .R(n524), .D(n175), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n511), .R(n524), .D(n176), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n511), .R(n524), .D(n178), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n511), .R(n524), .D(n180), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n511), .R(n524), .D(n182), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n511), .R(n524), .D(n184), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n511), .R(n524), .D(n186), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n511), .R(n524), .D(n188), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n511), .R(n524), .D(n190), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n511), .R(n524), .D(n192), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n511), .R(n524), .D(n194), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n511), .R(n524), .D(n196), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n511), .R(n524), .D(n198), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n511), .R(n524), .D(n200), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n511), .R(n524), .D(n202), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n511), .R(n524), .D(n204), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n511), .R(n524), .D(n206), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n511), .R(n524), .D(n208), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n511), .R(n524), .D(n210), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n511), .R(n524), .D(n212), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n511), .R(n524), .D(n214), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n511), .R(n524), .D(n216), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n511), .R(n524), .D(n218), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n511), .R(n524), .D(n220), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n511), .R(n524), .D(n222), .Q(rd_dat[31]));
Q_FDP4EP \rd_dat_REG[32] ( .CK(clk), .CE(n511), .R(n524), .D(n224), .Q(rd_dat[32]));
Q_FDP4EP \rd_dat_REG[33] ( .CK(clk), .CE(n511), .R(n524), .D(n226), .Q(rd_dat[33]));
Q_FDP4EP \rd_dat_REG[34] ( .CK(clk), .CE(n511), .R(n524), .D(n228), .Q(rd_dat[34]));
Q_FDP4EP \rd_dat_REG[35] ( .CK(clk), .CE(n511), .R(n524), .D(n230), .Q(rd_dat[35]));
Q_FDP4EP \rd_dat_REG[36] ( .CK(clk), .CE(n511), .R(n524), .D(n232), .Q(rd_dat[36]));
Q_FDP4EP \rd_dat_REG[37] ( .CK(clk), .CE(n511), .R(n524), .D(n234), .Q(rd_dat[37]));
Q_FDP4EP \rd_dat_REG[38] ( .CK(clk), .CE(n511), .R(n524), .D(n236), .Q(rd_dat[38]));
Q_FDP4EP \rd_dat_REG[39] ( .CK(clk), .CE(n511), .R(n524), .D(n238), .Q(rd_dat[39]));
Q_FDP4EP \rd_dat_REG[40] ( .CK(clk), .CE(n511), .R(n524), .D(n240), .Q(rd_dat[40]));
Q_FDP4EP \rd_dat_REG[41] ( .CK(clk), .CE(n511), .R(n524), .D(n242), .Q(rd_dat[41]));
Q_FDP4EP \rd_dat_REG[42] ( .CK(clk), .CE(n511), .R(n524), .D(n244), .Q(rd_dat[42]));
Q_FDP4EP \rd_dat_REG[43] ( .CK(clk), .CE(n511), .R(n524), .D(n246), .Q(rd_dat[43]));
Q_FDP4EP \rd_dat_REG[44] ( .CK(clk), .CE(n511), .R(n524), .D(n248), .Q(rd_dat[44]));
Q_FDP4EP \rd_dat_REG[45] ( .CK(clk), .CE(n511), .R(n524), .D(n250), .Q(rd_dat[45]));
Q_FDP4EP \rd_dat_REG[46] ( .CK(clk), .CE(n511), .R(n524), .D(n252), .Q(rd_dat[46]));
Q_FDP4EP \rd_dat_REG[47] ( .CK(clk), .CE(n511), .R(n524), .D(n254), .Q(rd_dat[47]));
Q_FDP4EP \rd_dat_REG[48] ( .CK(clk), .CE(n511), .R(n524), .D(n256), .Q(rd_dat[48]));
Q_FDP4EP \rd_dat_REG[49] ( .CK(clk), .CE(n511), .R(n524), .D(n258), .Q(rd_dat[49]));
Q_FDP4EP \rd_dat_REG[50] ( .CK(clk), .CE(n511), .R(n524), .D(n260), .Q(rd_dat[50]));
Q_FDP4EP \rd_dat_REG[51] ( .CK(clk), .CE(n511), .R(n524), .D(n262), .Q(rd_dat[51]));
Q_FDP4EP \rd_dat_REG[52] ( .CK(clk), .CE(n511), .R(n524), .D(n264), .Q(rd_dat[52]));
Q_FDP4EP \rd_dat_REG[53] ( .CK(clk), .CE(n511), .R(n524), .D(n266), .Q(rd_dat[53]));
Q_FDP4EP \rd_dat_REG[54] ( .CK(clk), .CE(n511), .R(n524), .D(n268), .Q(rd_dat[54]));
Q_FDP4EP \rd_dat_REG[55] ( .CK(clk), .CE(n511), .R(n524), .D(n270), .Q(rd_dat[55]));
Q_FDP4EP \rd_dat_REG[56] ( .CK(clk), .CE(n511), .R(n524), .D(n272), .Q(rd_dat[56]));
Q_FDP4EP \rd_dat_REG[57] ( .CK(clk), .CE(n511), .R(n524), .D(n274), .Q(rd_dat[57]));
Q_FDP4EP \rd_dat_REG[58] ( .CK(clk), .CE(n511), .R(n524), .D(n276), .Q(rd_dat[58]));
Q_FDP4EP \rd_dat_REG[59] ( .CK(clk), .CE(n511), .R(n524), .D(n278), .Q(rd_dat[59]));
Q_FDP4EP \rd_dat_REG[60] ( .CK(clk), .CE(n511), .R(n524), .D(n280), .Q(rd_dat[60]));
Q_FDP4EP \rd_dat_REG[61] ( .CK(clk), .CE(n511), .R(n524), .D(n282), .Q(rd_dat[61]));
Q_FDP4EP \rd_dat_REG[62] ( .CK(clk), .CE(n511), .R(n524), .D(n284), .Q(rd_dat[62]));
Q_FDP4EP \rd_dat_REG[63] ( .CK(clk), .CE(n511), .R(n524), .D(n286), .Q(rd_dat[63]));
Q_FDP4EP \rd_dat_REG[64] ( .CK(clk), .CE(n511), .R(n524), .D(n288), .Q(rd_dat[64]));
Q_FDP4EP \rd_dat_REG[65] ( .CK(clk), .CE(n511), .R(n524), .D(n290), .Q(rd_dat[65]));
Q_FDP4EP \rd_dat_REG[66] ( .CK(clk), .CE(n511), .R(n524), .D(n292), .Q(rd_dat[66]));
Q_FDP4EP \rd_dat_REG[67] ( .CK(clk), .CE(n511), .R(n524), .D(n294), .Q(rd_dat[67]));
Q_FDP4EP \rd_dat_REG[68] ( .CK(clk), .CE(n511), .R(n524), .D(n296), .Q(rd_dat[68]));
Q_FDP4EP \rd_dat_REG[69] ( .CK(clk), .CE(n511), .R(n524), .D(n298), .Q(rd_dat[69]));
Q_FDP4EP \rd_dat_REG[70] ( .CK(clk), .CE(n511), .R(n524), .D(n300), .Q(rd_dat[70]));
Q_FDP4EP \rd_dat_REG[71] ( .CK(clk), .CE(n511), .R(n524), .D(n302), .Q(rd_dat[71]));
Q_FDP4EP \rd_dat_REG[72] ( .CK(clk), .CE(n511), .R(n524), .D(n304), .Q(rd_dat[72]));
Q_FDP4EP \rd_dat_REG[73] ( .CK(clk), .CE(n511), .R(n524), .D(n306), .Q(rd_dat[73]));
Q_FDP4EP \rd_dat_REG[74] ( .CK(clk), .CE(n511), .R(n524), .D(n308), .Q(rd_dat[74]));
Q_FDP4EP \rd_dat_REG[75] ( .CK(clk), .CE(n511), .R(n524), .D(n310), .Q(rd_dat[75]));
Q_FDP4EP \rd_dat_REG[76] ( .CK(clk), .CE(n511), .R(n524), .D(n312), .Q(rd_dat[76]));
Q_FDP4EP \rd_dat_REG[77] ( .CK(clk), .CE(n511), .R(n524), .D(n314), .Q(rd_dat[77]));
Q_FDP4EP \rd_dat_REG[78] ( .CK(clk), .CE(n511), .R(n524), .D(n316), .Q(rd_dat[78]));
Q_FDP4EP \rd_dat_REG[79] ( .CK(clk), .CE(n511), .R(n524), .D(n318), .Q(rd_dat[79]));
Q_FDP4EP \rd_dat_REG[80] ( .CK(clk), .CE(n511), .R(n524), .D(n320), .Q(rd_dat[80]));
Q_FDP4EP \rd_dat_REG[81] ( .CK(clk), .CE(n511), .R(n524), .D(n322), .Q(rd_dat[81]));
Q_FDP4EP \rd_dat_REG[82] ( .CK(clk), .CE(n511), .R(n524), .D(n324), .Q(rd_dat[82]));
Q_FDP4EP \rd_dat_REG[83] ( .CK(clk), .CE(n511), .R(n524), .D(n326), .Q(rd_dat[83]));
Q_FDP4EP \rd_dat_REG[84] ( .CK(clk), .CE(n511), .R(n524), .D(n328), .Q(rd_dat[84]));
Q_FDP4EP \rd_dat_REG[85] ( .CK(clk), .CE(n511), .R(n524), .D(n330), .Q(rd_dat[85]));
Q_FDP4EP \rd_dat_REG[86] ( .CK(clk), .CE(n511), .R(n524), .D(n332), .Q(rd_dat[86]));
Q_FDP4EP \rd_dat_REG[87] ( .CK(clk), .CE(n511), .R(n524), .D(n334), .Q(rd_dat[87]));
Q_FDP4EP \rd_dat_REG[88] ( .CK(clk), .CE(n511), .R(n524), .D(n336), .Q(rd_dat[88]));
Q_FDP4EP \rd_dat_REG[89] ( .CK(clk), .CE(n511), .R(n524), .D(n338), .Q(rd_dat[89]));
Q_FDP4EP \rd_dat_REG[90] ( .CK(clk), .CE(n511), .R(n524), .D(n340), .Q(rd_dat[90]));
Q_FDP4EP \rd_dat_REG[91] ( .CK(clk), .CE(n511), .R(n524), .D(n342), .Q(rd_dat[91]));
Q_FDP4EP \rd_dat_REG[92] ( .CK(clk), .CE(n511), .R(n524), .D(n344), .Q(rd_dat[92]));
Q_FDP4EP \rd_dat_REG[93] ( .CK(clk), .CE(n511), .R(n524), .D(n346), .Q(rd_dat[93]));
Q_FDP4EP \rd_dat_REG[94] ( .CK(clk), .CE(n511), .R(n524), .D(n348), .Q(rd_dat[94]));
Q_FDP4EP \rd_dat_REG[95] ( .CK(clk), .CE(n511), .R(n524), .D(n350), .Q(rd_dat[95]));
Q_INV U810 ( .A(n514), .Z(n525));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n525), .R(n524), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 8 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
