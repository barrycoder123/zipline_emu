
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif

module cr_crc ( crc, clk, rst_n, data_in, data_valid, data_vbytes, enable, 
	init_value, init);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
output [31:0] crc;
input clk;
input rst_n;
input [63:0] data_in;
input data_valid;
input [7:0] data_vbytes;
input enable;
input [31:0] init_value;
input init;
wire [0:31] _zy_simnet_crc_0_w$;
wire [31:0] crc_r;
wire [7:0] data_vbits;
supply0 n1;
Q_BUF U0 ( .A(n1), .Z(data_vbits[0]));
Q_BUF U1 ( .A(n1), .Z(data_vbits[1]));
Q_BUF U2 ( .A(n1), .Z(data_vbits[2]));
Q_BUF U3 ( .A(n1), .Z(data_vbits[7]));
ixc_assign_32 _zz_strnp_0 ( _zy_simnet_crc_0_w$[0:31], crc[31:0]);
Q_AN02 U5 ( .A0(enable), .A1(n2), .Z(crc[31]));
Q_AN02 U6 ( .A0(enable), .A1(n3), .Z(crc[30]));
Q_AN02 U7 ( .A0(enable), .A1(n4), .Z(crc[29]));
Q_AN02 U8 ( .A0(enable), .A1(n5), .Z(crc[28]));
Q_AN02 U9 ( .A0(enable), .A1(n6), .Z(crc[27]));
Q_AN02 U10 ( .A0(enable), .A1(n7), .Z(crc[26]));
Q_AN02 U11 ( .A0(enable), .A1(n8), .Z(crc[25]));
Q_AN02 U12 ( .A0(enable), .A1(n9), .Z(crc[24]));
Q_AN02 U13 ( .A0(enable), .A1(n10), .Z(crc[23]));
Q_AN02 U14 ( .A0(enable), .A1(n11), .Z(crc[22]));
Q_AN02 U15 ( .A0(enable), .A1(n12), .Z(crc[21]));
Q_AN02 U16 ( .A0(enable), .A1(n13), .Z(crc[20]));
Q_AN02 U17 ( .A0(enable), .A1(n14), .Z(crc[19]));
Q_AN02 U18 ( .A0(enable), .A1(n15), .Z(crc[18]));
Q_AN02 U19 ( .A0(enable), .A1(n16), .Z(crc[17]));
Q_AN02 U20 ( .A0(enable), .A1(n17), .Z(crc[16]));
Q_AN02 U21 ( .A0(enable), .A1(n18), .Z(crc[15]));
Q_AN02 U22 ( .A0(enable), .A1(n19), .Z(crc[14]));
Q_AN02 U23 ( .A0(enable), .A1(n20), .Z(crc[13]));
Q_AN02 U24 ( .A0(enable), .A1(n21), .Z(crc[12]));
Q_AN02 U25 ( .A0(enable), .A1(n22), .Z(crc[11]));
Q_AN02 U26 ( .A0(enable), .A1(n23), .Z(crc[10]));
Q_AN02 U27 ( .A0(enable), .A1(n24), .Z(crc[9]));
Q_AN02 U28 ( .A0(enable), .A1(n25), .Z(crc[8]));
Q_AN02 U29 ( .A0(enable), .A1(n26), .Z(crc[7]));
Q_AN02 U30 ( .A0(enable), .A1(n27), .Z(crc[6]));
Q_AN02 U31 ( .A0(enable), .A1(n28), .Z(crc[5]));
Q_AN02 U32 ( .A0(enable), .A1(n29), .Z(crc[4]));
Q_AN02 U33 ( .A0(enable), .A1(n30), .Z(crc[3]));
Q_AN02 U34 ( .A0(enable), .A1(n31), .Z(crc[2]));
Q_AN02 U35 ( .A0(enable), .A1(n32), .Z(crc[1]));
Q_AN02 U36 ( .A0(enable), .A1(n33), .Z(crc[0]));
Q_AN02 U37 ( .A0(data_vbytes[7]), .A1(data_vbytes[6]), .Z(n34));
Q_AN02 U38 ( .A0(data_vbytes[5]), .A1(data_vbytes[4]), .Z(n41));
Q_AN03 U39 ( .A0(n34), .A1(n41), .A2(n37), .Z(data_vbits[6]));
Q_AN02 U40 ( .A0(data_vbytes[3]), .A1(data_vbytes[2]), .Z(n49));
Q_AN02 U41 ( .A0(data_vbytes[1]), .A1(data_vbytes[0]), .Z(n42));
Q_AN02 U42 ( .A0(n49), .A1(n42), .Z(n37));
Q_INV U43 ( .A(data_vbytes[6]), .Z(n44));
Q_AN02 U44 ( .A0(data_vbytes[6]), .A1(data_vbytes[5]), .Z(n45));
Q_OR02 U45 ( .A0(n44), .A1(n45), .Z(n36));
Q_NR02 U46 ( .A0(data_vbytes[5]), .A1(data_vbytes[4]), .Z(n35));
Q_AN02 U47 ( .A0(n44), .A1(n35), .Z(n40));
Q_AO21 U48 ( .A0(n36), .A1(data_vbytes[4]), .B0(n40), .Z(n38));
Q_INV U49 ( .A(data_vbytes[7]), .Z(n52));
Q_AN03 U50 ( .A0(n52), .A1(n37), .A2(n38), .Z(data_vbits[5]));
Q_INV U51 ( .A(data_vbytes[3]), .Z(n39));
Q_AN02 U52 ( .A0(n40), .A1(n39), .Z(n47));
Q_AO21 U53 ( .A0(n41), .A1(n49), .B0(n47), .Z(n43));
Q_AN03 U54 ( .A0(n52), .A1(n42), .A2(n43), .Z(data_vbits[4]));
Q_NR02 U55 ( .A0(data_vbytes[6]), .A1(data_vbytes[5]), .Z(n46));
Q_OA21 U56 ( .A0(n46), .A1(n45), .B0(n50), .Z(n51));
Q_AO21 U57 ( .A0(n48), .A1(n47), .B0(n51), .Z(n53));
Q_AN03 U58 ( .A0(data_vbytes[4]), .A1(data_vbytes[1]), .A2(n49), .Z(n50));
Q_AN03 U59 ( .A0(n52), .A1(data_vbytes[0]), .A2(n53), .Z(data_vbits[3]));
Q_XOR2 U60 ( .A0(data_in[0]), .A1(crc_r[0]), .Z(n54));
Q_XOR2 U61 ( .A0(data_in[1]), .A1(crc_r[1]), .Z(n55));
Q_XOR2 U62 ( .A0(data_in[2]), .A1(crc_r[2]), .Z(n56));
Q_XOR2 U63 ( .A0(data_in[3]), .A1(crc_r[3]), .Z(n57));
Q_XOR2 U64 ( .A0(data_in[4]), .A1(crc_r[4]), .Z(n58));
Q_XOR2 U65 ( .A0(data_in[5]), .A1(crc_r[5]), .Z(n59));
Q_XOR2 U66 ( .A0(data_in[6]), .A1(crc_r[6]), .Z(n60));
Q_XOR2 U67 ( .A0(data_in[7]), .A1(crc_r[7]), .Z(n61));
Q_XOR2 U68 ( .A0(data_in[8]), .A1(crc_r[8]), .Z(n62));
Q_XOR2 U69 ( .A0(data_in[9]), .A1(crc_r[9]), .Z(n63));
Q_XOR2 U70 ( .A0(data_in[10]), .A1(crc_r[10]), .Z(n64));
Q_XOR2 U71 ( .A0(data_in[11]), .A1(crc_r[11]), .Z(n65));
Q_XOR2 U72 ( .A0(data_in[12]), .A1(crc_r[12]), .Z(n66));
Q_XOR2 U73 ( .A0(data_in[13]), .A1(crc_r[13]), .Z(n67));
Q_XOR2 U74 ( .A0(data_in[14]), .A1(crc_r[14]), .Z(n68));
Q_XOR2 U75 ( .A0(data_in[15]), .A1(crc_r[15]), .Z(n69));
Q_XOR2 U76 ( .A0(data_in[16]), .A1(crc_r[16]), .Z(n70));
Q_XOR2 U77 ( .A0(data_in[17]), .A1(crc_r[17]), .Z(n71));
Q_XOR2 U78 ( .A0(data_in[18]), .A1(crc_r[18]), .Z(n72));
Q_XOR2 U79 ( .A0(data_in[19]), .A1(crc_r[19]), .Z(n73));
Q_XOR2 U80 ( .A0(data_in[20]), .A1(crc_r[20]), .Z(n74));
Q_XOR2 U81 ( .A0(data_in[21]), .A1(crc_r[21]), .Z(n75));
Q_XOR2 U82 ( .A0(data_in[22]), .A1(crc_r[22]), .Z(n76));
Q_XOR2 U83 ( .A0(data_in[23]), .A1(crc_r[23]), .Z(n77));
Q_XOR2 U84 ( .A0(data_in[24]), .A1(crc_r[24]), .Z(n78));
Q_XOR2 U85 ( .A0(data_in[25]), .A1(crc_r[25]), .Z(n79));
Q_XOR2 U86 ( .A0(data_in[26]), .A1(crc_r[26]), .Z(n80));
Q_XOR2 U87 ( .A0(data_in[27]), .A1(crc_r[27]), .Z(n81));
Q_XOR2 U88 ( .A0(data_in[28]), .A1(crc_r[28]), .Z(n82));
Q_XOR2 U89 ( .A0(data_in[29]), .A1(crc_r[29]), .Z(n83));
Q_XOR2 U90 ( .A0(data_in[30]), .A1(crc_r[30]), .Z(n84));
Q_XOR2 U91 ( .A0(data_in[31]), .A1(crc_r[31]), .Z(n85));
Q_MX02 U92 ( .S(data_vbits[3]), .A0(data_in[56]), .A1(n54), .Z(n86));
Q_MX02 U93 ( .S(data_vbits[3]), .A0(data_in[57]), .A1(n55), .Z(n87));
Q_MX02 U94 ( .S(data_vbits[3]), .A0(data_in[58]), .A1(n56), .Z(n88));
Q_MX02 U95 ( .S(data_vbits[3]), .A0(data_in[59]), .A1(n57), .Z(n89));
Q_MX02 U96 ( .S(data_vbits[3]), .A0(data_in[60]), .A1(n58), .Z(n90));
Q_MX02 U97 ( .S(data_vbits[3]), .A0(data_in[61]), .A1(n59), .Z(n91));
Q_MX02 U98 ( .S(data_vbits[3]), .A0(data_in[62]), .A1(n60), .Z(n92));
Q_MX02 U99 ( .S(data_vbits[3]), .A0(data_in[63]), .A1(n61), .Z(n93));
Q_MX02 U100 ( .S(data_vbits[3]), .A0(n54), .A1(n62), .Z(n94));
Q_MX02 U101 ( .S(data_vbits[3]), .A0(n55), .A1(n63), .Z(n95));
Q_MX02 U102 ( .S(data_vbits[3]), .A0(n56), .A1(n64), .Z(n96));
Q_MX02 U103 ( .S(data_vbits[3]), .A0(n57), .A1(n65), .Z(n97));
Q_MX02 U104 ( .S(data_vbits[3]), .A0(n58), .A1(n66), .Z(n98));
Q_MX02 U105 ( .S(data_vbits[3]), .A0(n59), .A1(n67), .Z(n99));
Q_MX02 U106 ( .S(data_vbits[3]), .A0(n60), .A1(n68), .Z(n100));
Q_MX02 U107 ( .S(data_vbits[3]), .A0(n61), .A1(n69), .Z(n101));
Q_MX02 U108 ( .S(data_vbits[3]), .A0(n62), .A1(n70), .Z(n102));
Q_MX02 U109 ( .S(data_vbits[3]), .A0(n63), .A1(n71), .Z(n103));
Q_MX02 U110 ( .S(data_vbits[3]), .A0(n64), .A1(n72), .Z(n104));
Q_MX02 U111 ( .S(data_vbits[3]), .A0(n65), .A1(n73), .Z(n105));
Q_MX02 U112 ( .S(data_vbits[3]), .A0(n66), .A1(n74), .Z(n106));
Q_MX02 U113 ( .S(data_vbits[3]), .A0(n67), .A1(n75), .Z(n107));
Q_MX02 U114 ( .S(data_vbits[3]), .A0(n68), .A1(n76), .Z(n108));
Q_MX02 U115 ( .S(data_vbits[3]), .A0(n69), .A1(n77), .Z(n109));
Q_MX02 U116 ( .S(data_vbits[3]), .A0(n70), .A1(n78), .Z(n110));
Q_MX02 U117 ( .S(data_vbits[3]), .A0(n71), .A1(n79), .Z(n111));
Q_MX02 U118 ( .S(data_vbits[3]), .A0(n72), .A1(n80), .Z(n112));
Q_MX02 U119 ( .S(data_vbits[3]), .A0(n73), .A1(n81), .Z(n113));
Q_MX02 U120 ( .S(data_vbits[3]), .A0(n74), .A1(n82), .Z(n114));
Q_MX02 U121 ( .S(data_vbits[3]), .A0(n75), .A1(n83), .Z(n115));
Q_MX02 U122 ( .S(data_vbits[3]), .A0(n76), .A1(n84), .Z(n116));
Q_MX02 U123 ( .S(data_vbits[3]), .A0(n77), .A1(n85), .Z(n117));
Q_MX02 U124 ( .S(data_vbits[3]), .A0(n78), .A1(data_in[32]), .Z(n118));
Q_MX02 U125 ( .S(data_vbits[3]), .A0(n79), .A1(data_in[33]), .Z(n119));
Q_MX02 U126 ( .S(data_vbits[3]), .A0(n80), .A1(data_in[34]), .Z(n120));
Q_MX02 U127 ( .S(data_vbits[3]), .A0(n81), .A1(data_in[35]), .Z(n121));
Q_MX02 U128 ( .S(data_vbits[3]), .A0(n82), .A1(data_in[36]), .Z(n122));
Q_MX02 U129 ( .S(data_vbits[3]), .A0(n83), .A1(data_in[37]), .Z(n123));
Q_MX02 U130 ( .S(data_vbits[3]), .A0(n84), .A1(data_in[38]), .Z(n124));
Q_MX02 U131 ( .S(data_vbits[3]), .A0(n85), .A1(data_in[39]), .Z(n125));
Q_MX02 U132 ( .S(data_vbits[3]), .A0(data_in[32]), .A1(data_in[40]), .Z(n126));
Q_MX02 U133 ( .S(data_vbits[3]), .A0(data_in[33]), .A1(data_in[41]), .Z(n127));
Q_MX02 U134 ( .S(data_vbits[3]), .A0(data_in[34]), .A1(data_in[42]), .Z(n128));
Q_MX02 U135 ( .S(data_vbits[3]), .A0(data_in[35]), .A1(data_in[43]), .Z(n129));
Q_MX02 U136 ( .S(data_vbits[3]), .A0(data_in[36]), .A1(data_in[44]), .Z(n130));
Q_MX02 U137 ( .S(data_vbits[3]), .A0(data_in[37]), .A1(data_in[45]), .Z(n131));
Q_MX02 U138 ( .S(data_vbits[3]), .A0(data_in[38]), .A1(data_in[46]), .Z(n132));
Q_MX02 U139 ( .S(data_vbits[3]), .A0(data_in[39]), .A1(data_in[47]), .Z(n133));
Q_MX02 U140 ( .S(data_vbits[3]), .A0(data_in[40]), .A1(data_in[48]), .Z(n134));
Q_MX02 U141 ( .S(data_vbits[3]), .A0(data_in[41]), .A1(data_in[49]), .Z(n135));
Q_MX02 U142 ( .S(data_vbits[3]), .A0(data_in[42]), .A1(data_in[50]), .Z(n136));
Q_MX02 U143 ( .S(data_vbits[3]), .A0(data_in[43]), .A1(data_in[51]), .Z(n137));
Q_MX02 U144 ( .S(data_vbits[3]), .A0(data_in[44]), .A1(data_in[52]), .Z(n138));
Q_MX02 U145 ( .S(data_vbits[3]), .A0(data_in[45]), .A1(data_in[53]), .Z(n139));
Q_MX02 U146 ( .S(data_vbits[3]), .A0(data_in[46]), .A1(data_in[54]), .Z(n140));
Q_MX02 U147 ( .S(data_vbits[3]), .A0(data_in[47]), .A1(data_in[55]), .Z(n141));
Q_MX02 U148 ( .S(data_vbits[3]), .A0(data_in[48]), .A1(data_in[56]), .Z(n142));
Q_MX02 U149 ( .S(data_vbits[3]), .A0(data_in[49]), .A1(data_in[57]), .Z(n143));
Q_MX02 U150 ( .S(data_vbits[3]), .A0(data_in[50]), .A1(data_in[58]), .Z(n144));
Q_MX02 U151 ( .S(data_vbits[3]), .A0(data_in[51]), .A1(data_in[59]), .Z(n145));
Q_MX02 U152 ( .S(data_vbits[3]), .A0(data_in[52]), .A1(data_in[60]), .Z(n146));
Q_MX02 U153 ( .S(data_vbits[3]), .A0(data_in[53]), .A1(data_in[61]), .Z(n147));
Q_MX02 U154 ( .S(data_vbits[3]), .A0(data_in[54]), .A1(data_in[62]), .Z(n148));
Q_MX02 U155 ( .S(data_vbits[3]), .A0(data_in[55]), .A1(data_in[63]), .Z(n149));
Q_INV U156 ( .A(data_vbits[3]), .Z(n342));
Q_AN02 U157 ( .A0(n342), .A1(data_in[56]), .Z(n150));
Q_AN02 U158 ( .A0(n342), .A1(data_in[57]), .Z(n151));
Q_AN02 U159 ( .A0(n342), .A1(data_in[58]), .Z(n152));
Q_AN02 U160 ( .A0(n342), .A1(data_in[59]), .Z(n153));
Q_AN02 U161 ( .A0(n342), .A1(data_in[60]), .Z(n154));
Q_AN02 U162 ( .A0(n342), .A1(data_in[61]), .Z(n155));
Q_AN02 U163 ( .A0(n342), .A1(data_in[62]), .Z(n156));
Q_AN02 U164 ( .A0(n342), .A1(data_in[63]), .Z(n157));
Q_MX02 U165 ( .S(data_vbits[4]), .A0(n134), .A1(n86), .Z(n158));
Q_MX02 U166 ( .S(data_vbits[4]), .A0(n135), .A1(n87), .Z(n159));
Q_MX02 U167 ( .S(data_vbits[4]), .A0(n136), .A1(n88), .Z(n160));
Q_MX02 U168 ( .S(data_vbits[4]), .A0(n137), .A1(n89), .Z(n161));
Q_MX02 U169 ( .S(data_vbits[4]), .A0(n138), .A1(n90), .Z(n162));
Q_MX02 U170 ( .S(data_vbits[4]), .A0(n139), .A1(n91), .Z(n163));
Q_MX02 U171 ( .S(data_vbits[4]), .A0(n140), .A1(n92), .Z(n164));
Q_MX02 U172 ( .S(data_vbits[4]), .A0(n141), .A1(n93), .Z(n165));
Q_MX02 U173 ( .S(data_vbits[4]), .A0(n142), .A1(n94), .Z(n166));
Q_MX02 U174 ( .S(data_vbits[4]), .A0(n143), .A1(n95), .Z(n167));
Q_MX02 U175 ( .S(data_vbits[4]), .A0(n144), .A1(n96), .Z(n168));
Q_MX02 U176 ( .S(data_vbits[4]), .A0(n145), .A1(n97), .Z(n169));
Q_MX02 U177 ( .S(data_vbits[4]), .A0(n146), .A1(n98), .Z(n170));
Q_MX02 U178 ( .S(data_vbits[4]), .A0(n147), .A1(n99), .Z(n171));
Q_MX02 U179 ( .S(data_vbits[4]), .A0(n148), .A1(n100), .Z(n172));
Q_MX02 U180 ( .S(data_vbits[4]), .A0(n149), .A1(n101), .Z(n173));
Q_MX02 U181 ( .S(data_vbits[4]), .A0(n86), .A1(n102), .Z(n174));
Q_MX02 U182 ( .S(data_vbits[4]), .A0(n87), .A1(n103), .Z(n175));
Q_MX02 U183 ( .S(data_vbits[4]), .A0(n88), .A1(n104), .Z(n176));
Q_MX02 U184 ( .S(data_vbits[4]), .A0(n89), .A1(n105), .Z(n177));
Q_MX02 U185 ( .S(data_vbits[4]), .A0(n90), .A1(n106), .Z(n178));
Q_MX02 U186 ( .S(data_vbits[4]), .A0(n91), .A1(n107), .Z(n179));
Q_MX02 U187 ( .S(data_vbits[4]), .A0(n92), .A1(n108), .Z(n180));
Q_MX02 U188 ( .S(data_vbits[4]), .A0(n93), .A1(n109), .Z(n181));
Q_MX02 U189 ( .S(data_vbits[4]), .A0(n94), .A1(n110), .Z(n182));
Q_MX02 U190 ( .S(data_vbits[4]), .A0(n95), .A1(n111), .Z(n183));
Q_MX02 U191 ( .S(data_vbits[4]), .A0(n96), .A1(n112), .Z(n184));
Q_MX02 U192 ( .S(data_vbits[4]), .A0(n97), .A1(n113), .Z(n185));
Q_MX02 U193 ( .S(data_vbits[4]), .A0(n98), .A1(n114), .Z(n186));
Q_MX02 U194 ( .S(data_vbits[4]), .A0(n99), .A1(n115), .Z(n187));
Q_MX02 U195 ( .S(data_vbits[4]), .A0(n100), .A1(n116), .Z(n188));
Q_MX02 U196 ( .S(data_vbits[4]), .A0(n101), .A1(n117), .Z(n189));
Q_MX02 U197 ( .S(data_vbits[4]), .A0(n102), .A1(n118), .Z(n190));
Q_MX02 U198 ( .S(data_vbits[4]), .A0(n103), .A1(n119), .Z(n191));
Q_MX02 U199 ( .S(data_vbits[4]), .A0(n104), .A1(n120), .Z(n192));
Q_MX02 U200 ( .S(data_vbits[4]), .A0(n105), .A1(n121), .Z(n193));
Q_MX02 U201 ( .S(data_vbits[4]), .A0(n106), .A1(n122), .Z(n194));
Q_MX02 U202 ( .S(data_vbits[4]), .A0(n107), .A1(n123), .Z(n195));
Q_MX02 U203 ( .S(data_vbits[4]), .A0(n108), .A1(n124), .Z(n196));
Q_MX02 U204 ( .S(data_vbits[4]), .A0(n109), .A1(n125), .Z(n197));
Q_MX02 U205 ( .S(data_vbits[4]), .A0(n110), .A1(n126), .Z(n198));
Q_MX02 U206 ( .S(data_vbits[4]), .A0(n111), .A1(n127), .Z(n199));
Q_MX02 U207 ( .S(data_vbits[4]), .A0(n112), .A1(n128), .Z(n200));
Q_MX02 U208 ( .S(data_vbits[4]), .A0(n113), .A1(n129), .Z(n201));
Q_MX02 U209 ( .S(data_vbits[4]), .A0(n114), .A1(n130), .Z(n202));
Q_MX02 U210 ( .S(data_vbits[4]), .A0(n115), .A1(n131), .Z(n203));
Q_MX02 U211 ( .S(data_vbits[4]), .A0(n116), .A1(n132), .Z(n204));
Q_MX02 U212 ( .S(data_vbits[4]), .A0(n117), .A1(n133), .Z(n205));
Q_MX02 U213 ( .S(data_vbits[4]), .A0(n118), .A1(n134), .Z(n206));
Q_MX02 U214 ( .S(data_vbits[4]), .A0(n119), .A1(n135), .Z(n207));
Q_MX02 U215 ( .S(data_vbits[4]), .A0(n120), .A1(n136), .Z(n208));
Q_MX02 U216 ( .S(data_vbits[4]), .A0(n121), .A1(n137), .Z(n209));
Q_MX02 U217 ( .S(data_vbits[4]), .A0(n122), .A1(n138), .Z(n210));
Q_MX02 U218 ( .S(data_vbits[4]), .A0(n123), .A1(n139), .Z(n211));
Q_MX02 U219 ( .S(data_vbits[4]), .A0(n124), .A1(n140), .Z(n212));
Q_MX02 U220 ( .S(data_vbits[4]), .A0(n125), .A1(n141), .Z(n213));
Q_MX02 U221 ( .S(data_vbits[4]), .A0(n126), .A1(n142), .Z(n214));
Q_MX02 U222 ( .S(data_vbits[4]), .A0(n127), .A1(n143), .Z(n215));
Q_MX02 U223 ( .S(data_vbits[4]), .A0(n128), .A1(n144), .Z(n216));
Q_MX02 U224 ( .S(data_vbits[4]), .A0(n129), .A1(n145), .Z(n217));
Q_MX02 U225 ( .S(data_vbits[4]), .A0(n130), .A1(n146), .Z(n218));
Q_MX02 U226 ( .S(data_vbits[4]), .A0(n131), .A1(n147), .Z(n219));
Q_MX02 U227 ( .S(data_vbits[4]), .A0(n132), .A1(n148), .Z(n220));
Q_MX02 U228 ( .S(data_vbits[4]), .A0(n133), .A1(n149), .Z(n221));
Q_MX02 U229 ( .S(data_vbits[4]), .A0(n134), .A1(n150), .Z(n222));
Q_MX02 U230 ( .S(data_vbits[4]), .A0(n135), .A1(n151), .Z(n223));
Q_MX02 U231 ( .S(data_vbits[4]), .A0(n136), .A1(n152), .Z(n224));
Q_MX02 U232 ( .S(data_vbits[4]), .A0(n137), .A1(n153), .Z(n225));
Q_MX02 U233 ( .S(data_vbits[4]), .A0(n138), .A1(n154), .Z(n226));
Q_MX02 U234 ( .S(data_vbits[4]), .A0(n139), .A1(n155), .Z(n227));
Q_MX02 U235 ( .S(data_vbits[4]), .A0(n140), .A1(n156), .Z(n228));
Q_MX02 U236 ( .S(data_vbits[4]), .A0(n141), .A1(n157), .Z(n229));
Q_INV U237 ( .A(data_vbits[4]), .Z(n343));
Q_AN02 U238 ( .A0(n343), .A1(n142), .Z(n230));
Q_AN02 U239 ( .A0(n343), .A1(n143), .Z(n231));
Q_AN02 U240 ( .A0(n343), .A1(n144), .Z(n232));
Q_AN02 U241 ( .A0(n343), .A1(n145), .Z(n233));
Q_AN02 U242 ( .A0(n343), .A1(n146), .Z(n234));
Q_AN02 U243 ( .A0(n343), .A1(n147), .Z(n235));
Q_AN02 U244 ( .A0(n343), .A1(n148), .Z(n236));
Q_AN02 U245 ( .A0(n343), .A1(n149), .Z(n237));
Q_AN02 U246 ( .A0(n343), .A1(n150), .Z(n238));
Q_AN02 U247 ( .A0(n343), .A1(n151), .Z(n239));
Q_AN02 U248 ( .A0(n343), .A1(n152), .Z(n240));
Q_AN02 U249 ( .A0(n343), .A1(n153), .Z(n241));
Q_AN02 U250 ( .A0(n343), .A1(n154), .Z(n242));
Q_AN02 U251 ( .A0(n343), .A1(n155), .Z(n243));
Q_AN02 U252 ( .A0(n343), .A1(n156), .Z(n244));
Q_AN02 U253 ( .A0(n343), .A1(n157), .Z(n245));
Q_MX02 U254 ( .S(data_vbits[5]), .A0(n182), .A1(n214), .Z(n246));
Q_MX02 U255 ( .S(data_vbits[5]), .A0(n183), .A1(n215), .Z(n247));
Q_MX02 U256 ( .S(data_vbits[5]), .A0(n184), .A1(n216), .Z(n248));
Q_MX02 U257 ( .S(data_vbits[5]), .A0(n185), .A1(n217), .Z(n249));
Q_MX02 U258 ( .S(data_vbits[5]), .A0(n186), .A1(n218), .Z(n250));
Q_MX02 U259 ( .S(data_vbits[5]), .A0(n187), .A1(n219), .Z(n251));
Q_MX02 U260 ( .S(data_vbits[5]), .A0(n188), .A1(n220), .Z(n252));
Q_MX02 U261 ( .S(data_vbits[5]), .A0(n189), .A1(n221), .Z(n253));
Q_INV U262 ( .A(data_vbits[5]), .Z(n347));
Q_AN02 U263 ( .A0(n347), .A1(n214), .Z(n254));
Q_AN02 U264 ( .A0(n347), .A1(n215), .Z(n255));
Q_AN02 U265 ( .A0(n347), .A1(n216), .Z(n256));
Q_AN02 U266 ( .A0(n347), .A1(n217), .Z(n257));
Q_AN02 U267 ( .A0(n347), .A1(n218), .Z(n258));
Q_AN02 U268 ( .A0(n347), .A1(n219), .Z(n259));
Q_AN02 U269 ( .A0(n347), .A1(n220), .Z(n260));
Q_AN02 U270 ( .A0(n347), .A1(n221), .Z(n261));
Q_AN02 U271 ( .A0(n347), .A1(n222), .Z(n262));
Q_AN02 U272 ( .A0(n347), .A1(n223), .Z(n263));
Q_AN02 U273 ( .A0(n347), .A1(n224), .Z(n264));
Q_AN02 U274 ( .A0(n347), .A1(n225), .Z(n265));
Q_AN02 U275 ( .A0(n347), .A1(n226), .Z(n266));
Q_AN02 U276 ( .A0(n347), .A1(n227), .Z(n267));
Q_AN02 U277 ( .A0(n347), .A1(n228), .Z(n268));
Q_AN02 U278 ( .A0(n347), .A1(n229), .Z(n269));
Q_AN02 U279 ( .A0(n347), .A1(n230), .Z(n270));
Q_AN02 U280 ( .A0(n347), .A1(n231), .Z(n271));
Q_AN02 U281 ( .A0(n347), .A1(n232), .Z(n272));
Q_AN02 U282 ( .A0(n347), .A1(n233), .Z(n273));
Q_AN02 U283 ( .A0(n347), .A1(n234), .Z(n274));
Q_AN02 U284 ( .A0(n347), .A1(n235), .Z(n275));
Q_AN02 U285 ( .A0(n347), .A1(n236), .Z(n276));
Q_AN02 U286 ( .A0(n347), .A1(n237), .Z(n277));
Q_AN02 U287 ( .A0(n347), .A1(n238), .Z(n278));
Q_AN02 U288 ( .A0(n347), .A1(n239), .Z(n279));
Q_AN02 U289 ( .A0(n347), .A1(n240), .Z(n280));
Q_AN02 U290 ( .A0(n347), .A1(n241), .Z(n281));
Q_AN02 U291 ( .A0(n347), .A1(n242), .Z(n282));
Q_AN02 U292 ( .A0(n347), .A1(n243), .Z(n283));
Q_AN02 U293 ( .A0(n347), .A1(n244), .Z(n284));
Q_AN02 U294 ( .A0(n347), .A1(n245), .Z(n285));
Q_MX03 U295 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n214), .A1(n182), .A2(n254), .Z(n310));
Q_MX03 U296 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n215), .A1(n183), .A2(n255), .Z(n311));
Q_MX03 U297 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n216), .A1(n184), .A2(n256), .Z(n312));
Q_MX03 U298 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n217), .A1(n185), .A2(n257), .Z(n313));
Q_MX03 U299 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n218), .A1(n186), .A2(n258), .Z(n314));
Q_MX03 U300 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n219), .A1(n187), .A2(n259), .Z(n315));
Q_MX03 U301 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n220), .A1(n188), .A2(n260), .Z(n316));
Q_MX03 U302 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n221), .A1(n189), .A2(n261), .Z(n317));
Q_MX03 U303 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n158), .A1(n190), .A2(n262), .Z(n318));
Q_MX03 U304 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n159), .A1(n191), .A2(n263), .Z(n319));
Q_MX03 U305 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n160), .A1(n192), .A2(n264), .Z(n320));
Q_MX03 U306 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n161), .A1(n193), .A2(n265), .Z(n321));
Q_MX03 U307 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n162), .A1(n194), .A2(n266), .Z(n322));
Q_MX03 U308 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n163), .A1(n195), .A2(n267), .Z(n323));
Q_MX03 U309 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n164), .A1(n196), .A2(n268), .Z(n324));
Q_MX03 U310 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n165), .A1(n197), .A2(n269), .Z(n325));
Q_MX03 U311 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n166), .A1(n198), .A2(n270), .Z(n326));
Q_MX03 U312 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n167), .A1(n199), .A2(n271), .Z(n327));
Q_MX03 U313 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n168), .A1(n200), .A2(n272), .Z(n328));
Q_MX03 U314 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n169), .A1(n201), .A2(n273), .Z(n329));
Q_MX03 U315 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n170), .A1(n202), .A2(n274), .Z(n330));
Q_MX03 U316 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n171), .A1(n203), .A2(n275), .Z(n331));
Q_MX03 U317 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n172), .A1(n204), .A2(n276), .Z(n332));
Q_MX03 U318 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n173), .A1(n205), .A2(n277), .Z(n333));
Q_MX03 U319 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n174), .A1(n206), .A2(n278), .Z(n334));
Q_MX03 U320 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n175), .A1(n207), .A2(n279), .Z(n335));
Q_MX03 U321 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n176), .A1(n208), .A2(n280), .Z(n336));
Q_MX03 U322 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n177), .A1(n209), .A2(n281), .Z(n337));
Q_MX03 U323 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n178), .A1(n210), .A2(n282), .Z(n338));
Q_MX03 U324 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n179), .A1(n211), .A2(n283), .Z(n339));
Q_MX03 U325 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n180), .A1(n212), .A2(n284), .Z(n340));
Q_MX03 U326 ( .S0(data_vbits[5]), .S1(data_vbits[6]), .A0(n181), .A1(n213), .A2(n285), .Z(n341));
Q_INV U327 ( .A(data_vbits[6]), .Z(n349));
Q_OR02 U328 ( .A0(n347), .A1(n508), .Z(n344));
Q_ND02 U329 ( .A0(data_vbits[5]), .A1(data_vbits[4]), .Z(n345));
Q_OR02 U330 ( .A0(n347), .A1(n509), .Z(n346));
Q_ND03 U331 ( .A0(n347), .A1(n508), .A2(n349), .Z(n353));
Q_NR02 U332 ( .A0(data_vbits[5]), .A1(data_vbits[4]), .Z(n348));
Q_ND03 U333 ( .A0(n347), .A1(n509), .A2(n349), .Z(n355));
Q_ND02 U334 ( .A0(n349), .A1(n344), .Z(n350));
Q_ND02 U335 ( .A0(n349), .A1(n345), .Z(n351));
Q_ND02 U336 ( .A0(n349), .A1(n346), .Z(n352));
Q_ND02 U337 ( .A0(n349), .A1(n348), .Z(n354));
Q_AN02 U338 ( .A0(n246), .A1(data_vbits[6]), .Z(n356));
Q_AN02 U339 ( .A0(n247), .A1(data_vbits[6]), .Z(n357));
Q_AN02 U340 ( .A0(n248), .A1(data_vbits[6]), .Z(n358));
Q_AN02 U341 ( .A0(n249), .A1(data_vbits[6]), .Z(n359));
Q_AN02 U342 ( .A0(n250), .A1(data_vbits[6]), .Z(n360));
Q_AN02 U343 ( .A0(n251), .A1(data_vbits[6]), .Z(n361));
Q_AN02 U344 ( .A0(n252), .A1(data_vbits[6]), .Z(n362));
Q_AN02 U345 ( .A0(n253), .A1(data_vbits[6]), .Z(n363));
Q_AN02 U346 ( .A0(n286), .A1(n350), .Z(n364));
Q_AN02 U347 ( .A0(n287), .A1(n350), .Z(n365));
Q_AN02 U348 ( .A0(n288), .A1(n350), .Z(n366));
Q_AN02 U349 ( .A0(n289), .A1(n350), .Z(n367));
Q_AN02 U350 ( .A0(n290), .A1(n350), .Z(n368));
Q_AN02 U351 ( .A0(n291), .A1(n350), .Z(n369));
Q_AN02 U352 ( .A0(n292), .A1(n350), .Z(n370));
Q_AN02 U353 ( .A0(n293), .A1(n350), .Z(n371));
Q_AN02 U354 ( .A0(n294), .A1(n351), .Z(n372));
Q_AN02 U355 ( .A0(n295), .A1(n351), .Z(n373));
Q_AN02 U356 ( .A0(n296), .A1(n351), .Z(n374));
Q_AN02 U357 ( .A0(n297), .A1(n351), .Z(n375));
Q_AN02 U358 ( .A0(n298), .A1(n351), .Z(n376));
Q_AN02 U359 ( .A0(n299), .A1(n351), .Z(n377));
Q_AN02 U360 ( .A0(n300), .A1(n351), .Z(n378));
Q_AN02 U361 ( .A0(n301), .A1(n351), .Z(n379));
Q_AN02 U362 ( .A0(n302), .A1(n352), .Z(n380));
Q_AN02 U363 ( .A0(n303), .A1(n352), .Z(n381));
Q_AN02 U364 ( .A0(n304), .A1(n352), .Z(n382));
Q_AN02 U365 ( .A0(n305), .A1(n352), .Z(n383));
Q_AN02 U366 ( .A0(n306), .A1(n352), .Z(n384));
Q_AN02 U367 ( .A0(n307), .A1(n352), .Z(n385));
Q_AN02 U368 ( .A0(n308), .A1(n352), .Z(n386));
Q_AN02 U369 ( .A0(n309), .A1(n352), .Z(n387));
Q_AN02 U370 ( .A0(n310), .A1(n510), .Z(n388));
Q_AN02 U371 ( .A0(n311), .A1(n510), .Z(n389));
Q_AN02 U372 ( .A0(n312), .A1(n510), .Z(n390));
Q_AN02 U373 ( .A0(n313), .A1(n510), .Z(n391));
Q_AN02 U374 ( .A0(n314), .A1(n510), .Z(n392));
Q_AN02 U375 ( .A0(n315), .A1(n510), .Z(n393));
Q_AN02 U376 ( .A0(n316), .A1(n510), .Z(n394));
Q_AN02 U377 ( .A0(n317), .A1(n510), .Z(n395));
Q_AN02 U378 ( .A0(n318), .A1(n353), .Z(n396));
Q_AN02 U379 ( .A0(n319), .A1(n353), .Z(n397));
Q_AN02 U380 ( .A0(n320), .A1(n353), .Z(n398));
Q_AN02 U381 ( .A0(n321), .A1(n353), .Z(n399));
Q_AN02 U382 ( .A0(n322), .A1(n353), .Z(n400));
Q_AN02 U383 ( .A0(n323), .A1(n353), .Z(n401));
Q_AN02 U384 ( .A0(n324), .A1(n353), .Z(n402));
Q_AN02 U385 ( .A0(n325), .A1(n353), .Z(n403));
Q_AN02 U386 ( .A0(n326), .A1(n354), .Z(n404));
Q_AN02 U387 ( .A0(n327), .A1(n354), .Z(n405));
Q_AN02 U388 ( .A0(n328), .A1(n354), .Z(n406));
Q_AN02 U389 ( .A0(n329), .A1(n354), .Z(n407));
Q_AN02 U390 ( .A0(n330), .A1(n354), .Z(n408));
Q_AN02 U391 ( .A0(n331), .A1(n354), .Z(n409));
Q_AN02 U392 ( .A0(n332), .A1(n354), .Z(n410));
Q_AN02 U393 ( .A0(n333), .A1(n354), .Z(n411));
Q_AN02 U394 ( .A0(n334), .A1(n355), .Z(n412));
Q_AN02 U395 ( .A0(n335), .A1(n355), .Z(n413));
Q_AN02 U396 ( .A0(n336), .A1(n355), .Z(n414));
Q_AN02 U397 ( .A0(n337), .A1(n355), .Z(n415));
Q_AN02 U398 ( .A0(n338), .A1(n355), .Z(n416));
Q_AN02 U399 ( .A0(n339), .A1(n355), .Z(n417));
Q_AN02 U400 ( .A0(n340), .A1(n355), .Z(n418));
Q_AN02 U401 ( .A0(n341), .A1(n355), .Z(n419));
Q_MX02 U402 ( .S(data_vbits[3]), .A0(crc_r[24]), .A1(crc_r[0]), .Z(n420));
Q_MX02 U403 ( .S(data_vbits[3]), .A0(crc_r[25]), .A1(crc_r[1]), .Z(n421));
Q_MX02 U404 ( .S(data_vbits[3]), .A0(crc_r[26]), .A1(crc_r[2]), .Z(n422));
Q_MX02 U405 ( .S(data_vbits[3]), .A0(crc_r[27]), .A1(crc_r[3]), .Z(n423));
Q_MX02 U406 ( .S(data_vbits[3]), .A0(crc_r[28]), .A1(crc_r[4]), .Z(n424));
Q_MX02 U407 ( .S(data_vbits[3]), .A0(crc_r[29]), .A1(crc_r[5]), .Z(n425));
Q_MX02 U408 ( .S(data_vbits[3]), .A0(crc_r[30]), .A1(crc_r[6]), .Z(n426));
Q_MX02 U409 ( .S(data_vbits[3]), .A0(crc_r[31]), .A1(crc_r[7]), .Z(n427));
Q_MX02 U410 ( .S(data_vbits[3]), .A0(crc_r[0]), .A1(crc_r[8]), .Z(n428));
Q_MX02 U411 ( .S(data_vbits[3]), .A0(crc_r[1]), .A1(crc_r[9]), .Z(n429));
Q_MX02 U412 ( .S(data_vbits[3]), .A0(crc_r[2]), .A1(crc_r[10]), .Z(n430));
Q_MX02 U413 ( .S(data_vbits[3]), .A0(crc_r[3]), .A1(crc_r[11]), .Z(n431));
Q_MX02 U414 ( .S(data_vbits[3]), .A0(crc_r[4]), .A1(crc_r[12]), .Z(n432));
Q_MX02 U415 ( .S(data_vbits[3]), .A0(crc_r[5]), .A1(crc_r[13]), .Z(n433));
Q_MX02 U416 ( .S(data_vbits[3]), .A0(crc_r[6]), .A1(crc_r[14]), .Z(n434));
Q_MX02 U417 ( .S(data_vbits[3]), .A0(crc_r[7]), .A1(crc_r[15]), .Z(n435));
Q_MX02 U418 ( .S(data_vbits[3]), .A0(crc_r[8]), .A1(crc_r[16]), .Z(n436));
Q_MX02 U419 ( .S(data_vbits[3]), .A0(crc_r[9]), .A1(crc_r[17]), .Z(n437));
Q_MX02 U420 ( .S(data_vbits[3]), .A0(crc_r[10]), .A1(crc_r[18]), .Z(n438));
Q_MX02 U421 ( .S(data_vbits[3]), .A0(crc_r[11]), .A1(crc_r[19]), .Z(n439));
Q_MX02 U422 ( .S(data_vbits[3]), .A0(crc_r[12]), .A1(crc_r[20]), .Z(n440));
Q_MX02 U423 ( .S(data_vbits[3]), .A0(crc_r[13]), .A1(crc_r[21]), .Z(n441));
Q_MX02 U424 ( .S(data_vbits[3]), .A0(crc_r[14]), .A1(crc_r[22]), .Z(n442));
Q_MX02 U425 ( .S(data_vbits[3]), .A0(crc_r[15]), .A1(crc_r[23]), .Z(n443));
Q_MX02 U426 ( .S(data_vbits[3]), .A0(crc_r[16]), .A1(crc_r[24]), .Z(n444));
Q_MX02 U427 ( .S(data_vbits[3]), .A0(crc_r[17]), .A1(crc_r[25]), .Z(n445));
Q_MX02 U428 ( .S(data_vbits[3]), .A0(crc_r[18]), .A1(crc_r[26]), .Z(n446));
Q_MX02 U429 ( .S(data_vbits[3]), .A0(crc_r[19]), .A1(crc_r[27]), .Z(n447));
Q_MX02 U430 ( .S(data_vbits[3]), .A0(crc_r[20]), .A1(crc_r[28]), .Z(n448));
Q_MX02 U431 ( .S(data_vbits[3]), .A0(crc_r[21]), .A1(crc_r[29]), .Z(n449));
Q_MX02 U432 ( .S(data_vbits[3]), .A0(crc_r[22]), .A1(crc_r[30]), .Z(n450));
Q_MX02 U433 ( .S(data_vbits[3]), .A0(crc_r[23]), .A1(crc_r[31]), .Z(n451));
Q_AN02 U434 ( .A0(n342), .A1(crc_r[24]), .Z(n452));
Q_AN02 U435 ( .A0(n342), .A1(crc_r[25]), .Z(n453));
Q_AN02 U436 ( .A0(n342), .A1(crc_r[26]), .Z(n454));
Q_AN02 U437 ( .A0(n342), .A1(crc_r[27]), .Z(n455));
Q_AN02 U438 ( .A0(n342), .A1(crc_r[28]), .Z(n456));
Q_AN02 U439 ( .A0(n342), .A1(crc_r[29]), .Z(n457));
Q_AN02 U440 ( .A0(n342), .A1(crc_r[30]), .Z(n458));
Q_AN02 U441 ( .A0(n342), .A1(crc_r[31]), .Z(n459));
Q_MX02 U442 ( .S(data_vbits[4]), .A0(n428), .A1(n444), .Z(n460));
Q_MX02 U443 ( .S(data_vbits[4]), .A0(n429), .A1(n445), .Z(n461));
Q_MX02 U444 ( .S(data_vbits[4]), .A0(n430), .A1(n446), .Z(n462));
Q_MX02 U445 ( .S(data_vbits[4]), .A0(n431), .A1(n447), .Z(n463));
Q_MX02 U446 ( .S(data_vbits[4]), .A0(n432), .A1(n448), .Z(n464));
Q_MX02 U447 ( .S(data_vbits[4]), .A0(n433), .A1(n449), .Z(n465));
Q_MX02 U448 ( .S(data_vbits[4]), .A0(n434), .A1(n450), .Z(n466));
Q_MX02 U449 ( .S(data_vbits[4]), .A0(n435), .A1(n451), .Z(n467));
Q_AN02 U450 ( .A0(n343), .A1(n444), .Z(n468));
Q_AN02 U451 ( .A0(n343), .A1(n445), .Z(n469));
Q_AN02 U452 ( .A0(n343), .A1(n446), .Z(n470));
Q_AN02 U453 ( .A0(n343), .A1(n447), .Z(n471));
Q_AN02 U454 ( .A0(n343), .A1(n448), .Z(n472));
Q_AN02 U455 ( .A0(n343), .A1(n449), .Z(n473));
Q_AN02 U456 ( .A0(n343), .A1(n450), .Z(n474));
Q_AN02 U457 ( .A0(n343), .A1(n451), .Z(n475));
Q_AN02 U458 ( .A0(n343), .A1(n452), .Z(n476));
Q_AN02 U459 ( .A0(n343), .A1(n453), .Z(n477));
Q_AN02 U460 ( .A0(n343), .A1(n454), .Z(n478));
Q_AN02 U461 ( .A0(n343), .A1(n455), .Z(n479));
Q_AN02 U462 ( .A0(n343), .A1(n456), .Z(n480));
Q_AN02 U463 ( .A0(n343), .A1(n457), .Z(n481));
Q_AN02 U464 ( .A0(n343), .A1(n458), .Z(n482));
Q_AN02 U465 ( .A0(n343), .A1(n459), .Z(n483));
Q_MX03 U466 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n444), .A1(n428), .A2(n468), .Z(n492));
Q_MX03 U467 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n445), .A1(n429), .A2(n469), .Z(n493));
Q_MX03 U468 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n446), .A1(n430), .A2(n470), .Z(n494));
Q_MX03 U469 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n447), .A1(n431), .A2(n471), .Z(n495));
Q_MX03 U470 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n448), .A1(n432), .A2(n472), .Z(n496));
Q_MX03 U471 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n449), .A1(n433), .A2(n473), .Z(n497));
Q_MX03 U472 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n450), .A1(n434), .A2(n474), .Z(n498));
Q_MX03 U473 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n451), .A1(n435), .A2(n475), .Z(n499));
Q_MX03 U474 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n420), .A1(n436), .A2(n476), .Z(n500));
Q_MX03 U475 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n421), .A1(n437), .A2(n477), .Z(n501));
Q_MX03 U476 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n422), .A1(n438), .A2(n478), .Z(n502));
Q_MX03 U477 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n423), .A1(n439), .A2(n479), .Z(n503));
Q_MX03 U478 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n424), .A1(n440), .A2(n480), .Z(n504));
Q_MX03 U479 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n425), .A1(n441), .A2(n481), .Z(n505));
Q_MX03 U480 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n426), .A1(n442), .A2(n482), .Z(n506));
Q_MX03 U481 ( .S0(data_vbits[4]), .S1(data_vbits[5]), .A0(n427), .A1(n443), .A2(n483), .Z(n507));
Q_AN03 U482 ( .A0(n349), .A1(n460), .A2(n511), .Z(n515));
Q_AN03 U483 ( .A0(n349), .A1(n461), .A2(n511), .Z(n516));
Q_AN03 U484 ( .A0(n349), .A1(n462), .A2(n511), .Z(n517));
Q_AN03 U485 ( .A0(n349), .A1(n463), .A2(n511), .Z(n518));
Q_AN03 U486 ( .A0(n349), .A1(n464), .A2(n511), .Z(n519));
Q_AN03 U487 ( .A0(n349), .A1(n465), .A2(n511), .Z(n520));
Q_AN03 U488 ( .A0(n349), .A1(n466), .A2(n511), .Z(n521));
Q_AN03 U489 ( .A0(n349), .A1(n467), .A2(n511), .Z(n522));
Q_AN03 U490 ( .A0(n349), .A1(n484), .A2(n512), .Z(n523));
Q_AN03 U491 ( .A0(n349), .A1(n485), .A2(n512), .Z(n524));
Q_AN03 U492 ( .A0(n349), .A1(n486), .A2(n512), .Z(n525));
Q_AN03 U493 ( .A0(n349), .A1(n487), .A2(n512), .Z(n526));
Q_AN03 U494 ( .A0(n349), .A1(n488), .A2(n512), .Z(n527));
Q_AN03 U495 ( .A0(n349), .A1(n489), .A2(n512), .Z(n528));
Q_AN03 U496 ( .A0(n349), .A1(n490), .A2(n512), .Z(n529));
Q_AN03 U497 ( .A0(n349), .A1(n491), .A2(n512), .Z(n530));
Q_AN03 U498 ( .A0(n349), .A1(n492), .A2(n513), .Z(n531));
Q_AN03 U499 ( .A0(n349), .A1(n493), .A2(n513), .Z(n532));
Q_AN03 U500 ( .A0(n349), .A1(n494), .A2(n513), .Z(n533));
Q_AN03 U501 ( .A0(n349), .A1(n495), .A2(n513), .Z(n534));
Q_AN03 U502 ( .A0(n349), .A1(n496), .A2(n513), .Z(n535));
Q_AN03 U503 ( .A0(n349), .A1(n497), .A2(n513), .Z(n536));
Q_AN03 U504 ( .A0(n349), .A1(n498), .A2(n513), .Z(n537));
Q_AN03 U505 ( .A0(n349), .A1(n499), .A2(n513), .Z(n538));
Q_AN03 U506 ( .A0(n349), .A1(n500), .A2(n514), .Z(n539));
Q_AN03 U507 ( .A0(n349), .A1(n501), .A2(n514), .Z(n540));
Q_AN03 U508 ( .A0(n349), .A1(n502), .A2(n514), .Z(n541));
Q_AN03 U509 ( .A0(n349), .A1(n503), .A2(n514), .Z(n542));
Q_AN03 U510 ( .A0(n349), .A1(n504), .A2(n514), .Z(n543));
Q_AN03 U511 ( .A0(n349), .A1(n505), .A2(n514), .Z(n544));
Q_AN03 U512 ( .A0(n349), .A1(n506), .A2(n514), .Z(n545));
Q_AN03 U513 ( .A0(n349), .A1(n507), .A2(n514), .Z(n546));
Q_ND02 U514 ( .A0(data_vbits[4]), .A1(data_vbits[3]), .Z(n508));
Q_NR02 U515 ( .A0(data_vbits[4]), .A1(data_vbits[3]), .Z(n509));
Q_OR02 U516 ( .A0(data_vbits[5]), .A1(data_vbits[6]), .Z(n510));
Q_INV U517 ( .A(n510), .Z(n511));
Q_AN02 U518 ( .A0(n511), .A1(n508), .Z(n512));
Q_NR02 U519 ( .A0(n510), .A1(data_vbits[4]), .Z(n513));
Q_AN02 U520 ( .A0(n511), .A1(n509), .Z(n514));
Q_XOR3 U521 ( .A0(n515), .A1(n416), .A2(n415), .Z(n547));
Q_XOR3 U522 ( .A0(n411), .A1(n408), .A2(n404), .Z(n548));
Q_XOR3 U523 ( .A0(n403), .A1(n402), .A2(n399), .Z(n549));
Q_XOR3 U524 ( .A0(n393), .A1(n392), .A2(n390), .Z(n550));
Q_XOR3 U525 ( .A0(n389), .A1(n385), .A2(n384), .Z(n551));
Q_XOR3 U526 ( .A0(n383), .A1(n378), .A2(n377), .Z(n552));
Q_XOR3 U527 ( .A0(n372), .A1(n369), .A2(n367), .Z(n553));
Q_XOR3 U528 ( .A0(n366), .A1(n361), .A2(n358), .Z(n554));
Q_XOR3 U529 ( .A0(n356), .A1(n547), .A2(n996), .Z(n555));
Q_XOR3 U530 ( .A0(n548), .A1(n549), .A2(n902), .Z(n556));
Q_XOR3 U531 ( .A0(n550), .A1(n551), .A2(n552), .Z(n557));
Q_XOR3 U532 ( .A0(n811), .A1(n553), .A2(n554), .Z(n558));
Q_XOR3 U533 ( .A0(n555), .A1(n556), .A2(n557), .Z(n559));
Q_XOR2 U534 ( .A0(n558), .A1(n559), .Z(n560));
Q_XOR3 U535 ( .A0(n516), .A1(n417), .A2(n416), .Z(n561));
Q_XOR3 U536 ( .A0(n412), .A1(n409), .A2(n405), .Z(n562));
Q_XOR3 U537 ( .A0(n404), .A1(n403), .A2(n400), .Z(n563));
Q_XOR3 U538 ( .A0(n394), .A1(n393), .A2(n391), .Z(n564));
Q_XOR3 U539 ( .A0(n390), .A1(n386), .A2(n385), .Z(n565));
Q_XOR3 U540 ( .A0(n384), .A1(n379), .A2(n378), .Z(n566));
Q_XOR3 U541 ( .A0(n373), .A1(n370), .A2(n368), .Z(n567));
Q_XOR3 U542 ( .A0(n367), .A1(n362), .A2(n359), .Z(n568));
Q_XOR3 U543 ( .A0(n357), .A1(n356), .A2(n561), .Z(n569));
Q_XOR3 U544 ( .A0(n719), .A1(n562), .A2(n563), .Z(n570));
Q_XOR3 U545 ( .A0(n608), .A1(n564), .A2(n565), .Z(n571));
Q_XOR3 U546 ( .A0(n566), .A1(n725), .A2(n567), .Z(n572));
Q_XOR3 U547 ( .A0(n568), .A1(n569), .A2(n570), .Z(n573));
Q_XOR3 U548 ( .A0(n571), .A1(n572), .A2(n573), .Z(n574));
Q_XOR3 U549 ( .A0(n517), .A1(n418), .A2(n417), .Z(n575));
Q_XOR3 U550 ( .A0(n413), .A1(n410), .A2(n406), .Z(n576));
Q_XOR3 U551 ( .A0(n405), .A1(n404), .A2(n401), .Z(n577));
Q_XOR3 U552 ( .A0(n395), .A1(n394), .A2(n392), .Z(n578));
Q_XOR3 U553 ( .A0(n391), .A1(n387), .A2(n386), .Z(n579));
Q_XOR3 U554 ( .A0(n385), .A1(n380), .A2(n379), .Z(n580));
Q_XOR3 U555 ( .A0(n377), .A1(n376), .A2(n375), .Z(n581));
Q_XOR3 U556 ( .A0(n374), .A1(n371), .A2(n369), .Z(n582));
Q_XOR3 U557 ( .A0(n368), .A1(n363), .A2(n360), .Z(n583));
Q_XOR3 U558 ( .A0(n575), .A1(n820), .A2(n576), .Z(n584));
Q_XOR3 U559 ( .A0(n577), .A1(n682), .A2(n578), .Z(n585));
Q_XOR3 U560 ( .A0(n579), .A1(n580), .A2(n581), .Z(n586));
Q_XOR3 U561 ( .A0(n582), .A1(n583), .A2(n826), .Z(n587));
Q_XOR3 U562 ( .A0(n584), .A1(n585), .A2(n586), .Z(n588));
Q_XOR2 U563 ( .A0(n587), .A1(n588), .Z(n589));
Q_XOR3 U564 ( .A0(n518), .A1(n419), .A2(n418), .Z(n590));
Q_XOR3 U565 ( .A0(n414), .A1(n411), .A2(n407), .Z(n591));
Q_XOR3 U566 ( .A0(n400), .A1(n398), .A2(n397), .Z(n592));
Q_XOR3 U567 ( .A0(n396), .A1(n395), .A2(n393), .Z(n593));
Q_XOR3 U568 ( .A0(n392), .A1(n388), .A2(n387), .Z(n594));
Q_XOR3 U569 ( .A0(n386), .A1(n381), .A2(n380), .Z(n595));
Q_XOR3 U570 ( .A0(n375), .A1(n372), .A2(n370), .Z(n596));
Q_XOR3 U571 ( .A0(n369), .A1(n364), .A2(n361), .Z(n597));
Q_XOR3 U572 ( .A0(n590), .A1(n832), .A2(n591), .Z(n598));
Q_XOR3 U573 ( .A0(n916), .A1(n592), .A2(n593), .Z(n599));
Q_XOR3 U574 ( .A0(n594), .A1(n595), .A2(n810), .Z(n600));
Q_XOR3 U575 ( .A0(n596), .A1(n597), .A2(n838), .Z(n601));
Q_XOR3 U576 ( .A0(n598), .A1(n599), .A2(n600), .Z(n602));
Q_XOR2 U577 ( .A0(n601), .A1(n602), .Z(n603));
Q_XOR3 U578 ( .A0(n519), .A1(n419), .A2(n418), .Z(n604));
Q_XOR3 U579 ( .A0(n417), .A1(n414), .A2(n413), .Z(n605));
Q_XOR3 U580 ( .A0(n411), .A1(n407), .A2(n406), .Z(n606));
Q_XOR3 U581 ( .A0(n404), .A1(n402), .A2(n401), .Z(n607));
Q_XOR3 U582 ( .A0(n398), .A1(n396), .A2(n395), .Z(n608));
Q_XOR3 U583 ( .A0(n392), .A1(n390), .A2(n388), .Z(n609));
Q_XOR3 U584 ( .A0(n387), .A1(n385), .A2(n384), .Z(n610));
Q_XOR3 U585 ( .A0(n383), .A1(n382), .A2(n381), .Z(n611));
Q_XOR3 U586 ( .A0(n379), .A1(n376), .A2(n375), .Z(n612));
Q_XOR3 U587 ( .A0(n370), .A1(n369), .A2(n367), .Z(n613));
Q_XOR3 U588 ( .A0(n366), .A1(n365), .A2(n362), .Z(n614));
Q_XOR3 U589 ( .A0(n361), .A1(n360), .A2(n359), .Z(n615));
Q_XOR3 U590 ( .A0(n604), .A1(n605), .A2(n606), .Z(n616));
Q_XOR3 U591 ( .A0(n607), .A1(n608), .A2(n609), .Z(n617));
Q_XOR3 U592 ( .A0(n610), .A1(n611), .A2(n612), .Z(n618));
Q_XOR3 U593 ( .A0(n970), .A1(n613), .A2(n614), .Z(n619));
Q_XOR3 U594 ( .A0(n615), .A1(n616), .A2(n617), .Z(n620));
Q_XOR3 U595 ( .A0(n618), .A1(n619), .A2(n620), .Z(n621));
Q_XOR3 U596 ( .A0(n520), .A1(n419), .A2(n418), .Z(n622));
Q_XOR3 U597 ( .A0(n416), .A1(n413), .A2(n411), .Z(n623));
Q_XOR3 U598 ( .A0(n407), .A1(n405), .A2(n404), .Z(n624));
Q_XOR3 U599 ( .A0(n396), .A1(n395), .A2(n394), .Z(n625));
Q_XOR3 U600 ( .A0(n388), .A1(n386), .A2(n382), .Z(n626));
Q_XOR3 U601 ( .A0(n380), .A1(n378), .A2(n376), .Z(n627));
Q_XOR3 U602 ( .A0(n374), .A1(n371), .A2(n370), .Z(n628));
Q_XOR3 U603 ( .A0(n369), .A1(n368), .A2(n363), .Z(n629));
Q_XOR3 U604 ( .A0(n362), .A1(n360), .A2(n358), .Z(n630));
Q_XOR3 U605 ( .A0(n356), .A1(n622), .A2(n623), .Z(n631));
Q_XOR3 U606 ( .A0(n624), .A1(n625), .A2(n983), .Z(n632));
Q_XOR3 U607 ( .A0(n626), .A1(n627), .A2(n628), .Z(n633));
Q_XOR3 U608 ( .A0(n629), .A1(n630), .A2(n631), .Z(n634));
Q_XOR3 U609 ( .A0(n632), .A1(n633), .A2(n634), .Z(n635));
Q_XOR3 U610 ( .A0(n521), .A1(n419), .A2(n417), .Z(n636));
Q_XOR3 U611 ( .A0(n416), .A1(n415), .A2(n413), .Z(n637));
Q_XOR3 U612 ( .A0(n411), .A1(n406), .A2(n405), .Z(n638));
Q_XOR3 U613 ( .A0(n399), .A1(n396), .A2(n394), .Z(n639));
Q_XOR3 U614 ( .A0(n391), .A1(n390), .A2(n387), .Z(n640));
Q_XOR3 U615 ( .A0(n385), .A1(n384), .A2(n381), .Z(n641));
Q_XOR3 U616 ( .A0(n379), .A1(n378), .A2(n374), .Z(n642));
Q_XOR3 U617 ( .A0(n367), .A1(n366), .A2(n364), .Z(n643));
Q_XOR3 U618 ( .A0(n363), .A1(n359), .A2(n358), .Z(n644));
Q_XOR3 U619 ( .A0(n357), .A1(n636), .A2(n637), .Z(n645));
Q_XOR3 U620 ( .A0(n638), .A1(n845), .A2(n639), .Z(n646));
Q_XOR3 U621 ( .A0(n640), .A1(n641), .A2(n642), .Z(n647));
Q_XOR3 U622 ( .A0(n954), .A1(n643), .A2(n644), .Z(n648));
Q_XOR3 U623 ( .A0(n645), .A1(n646), .A2(n647), .Z(n649));
Q_XOR2 U624 ( .A0(n648), .A1(n649), .Z(n650));
Q_XOR3 U625 ( .A0(n522), .A1(n418), .A2(n417), .Z(n651));
Q_XOR3 U626 ( .A0(n415), .A1(n413), .A2(n411), .Z(n652));
Q_XOR3 U627 ( .A0(n408), .A1(n407), .A2(n406), .Z(n653));
Q_XOR3 U628 ( .A0(n405), .A1(n402), .A2(n400), .Z(n654));
Q_XOR3 U629 ( .A0(n399), .A1(n394), .A2(n393), .Z(n655));
Q_XOR3 U630 ( .A0(n388), .A1(n386), .A2(n384), .Z(n656));
Q_XOR3 U631 ( .A0(n383), .A1(n382), .A2(n380), .Z(n657));
Q_XOR3 U632 ( .A0(n368), .A1(n366), .A2(n365), .Z(n658));
Q_XOR3 U633 ( .A0(n364), .A1(n361), .A2(n360), .Z(n659));
Q_XOR3 U634 ( .A0(n359), .A1(n651), .A2(n652), .Z(n660));
Q_XOR3 U635 ( .A0(n653), .A1(n654), .A2(n655), .Z(n661));
Q_XOR3 U636 ( .A0(n967), .A1(n656), .A2(n657), .Z(n662));
Q_XOR3 U637 ( .A0(n724), .A1(n824), .A2(n658), .Z(n663));
Q_XOR3 U638 ( .A0(n659), .A1(n660), .A2(n661), .Z(n664));
Q_XOR3 U639 ( .A0(n662), .A1(n663), .A2(n664), .Z(n665));
Q_XOR3 U640 ( .A0(n523), .A1(n419), .A2(n418), .Z(n666));
Q_XOR3 U641 ( .A0(n400), .A1(n395), .A2(n394), .Z(n667));
Q_XOR3 U642 ( .A0(n389), .A1(n387), .A2(n385), .Z(n668));
Q_XOR3 U643 ( .A0(n384), .A1(n383), .A2(n381), .Z(n669));
Q_XOR3 U644 ( .A0(n380), .A1(n379), .A2(n378), .Z(n670));
Q_XOR3 U645 ( .A0(n369), .A1(n367), .A2(n366), .Z(n671));
Q_XOR3 U646 ( .A0(n360), .A1(n356), .A2(n666), .Z(n672));
Q_XOR3 U647 ( .A0(n680), .A1(n915), .A2(n749), .Z(n673));
Q_XOR3 U648 ( .A0(n667), .A1(n983), .A2(n668), .Z(n674));
Q_XOR3 U649 ( .A0(n669), .A1(n670), .A2(n836), .Z(n675));
Q_XOR3 U650 ( .A0(n671), .A1(n754), .A2(n672), .Z(n676));
Q_XOR3 U651 ( .A0(n673), .A1(n674), .A2(n675), .Z(n677));
Q_XOR2 U652 ( .A0(n676), .A1(n677), .Z(n678));
Q_XOR3 U653 ( .A0(n524), .A1(n419), .A2(n417), .Z(n679));
Q_XOR3 U654 ( .A0(n416), .A1(n414), .A2(n412), .Z(n680));
Q_XOR3 U655 ( .A0(n407), .A1(n403), .A2(n401), .Z(n681));
Q_XOR3 U656 ( .A0(n399), .A1(n397), .A2(n396), .Z(n682));
Q_XOR3 U657 ( .A0(n394), .A1(n391), .A2(n389), .Z(n683));
Q_XOR3 U658 ( .A0(n363), .A1(n362), .A2(n358), .Z(n684));
Q_XOR3 U659 ( .A0(n357), .A1(n679), .A2(n680), .Z(n685));
Q_XOR3 U660 ( .A0(n947), .A1(n681), .A2(n682), .Z(n686));
Q_XOR3 U661 ( .A0(n683), .A1(n864), .A2(n708), .Z(n687));
Q_XOR3 U662 ( .A0(n724), .A1(n970), .A2(n781), .Z(n688));
Q_XOR3 U663 ( .A0(n684), .A1(n685), .A2(n686), .Z(n689));
Q_XOR3 U664 ( .A0(n687), .A1(n688), .A2(n689), .Z(n690));
Q_XOR3 U665 ( .A0(n525), .A1(n418), .A2(n417), .Z(n691));
Q_XOR3 U666 ( .A0(n416), .A1(n414), .A2(n410), .Z(n692));
Q_XOR3 U667 ( .A0(n403), .A1(n400), .A2(n399), .Z(n693));
Q_XOR3 U668 ( .A0(n398), .A1(n394), .A2(n393), .Z(n694));
Q_XOR3 U669 ( .A0(n381), .A1(n380), .A2(n379), .Z(n695));
Q_XOR3 U670 ( .A0(n377), .A1(n374), .A2(n371), .Z(n696));
Q_XOR3 U671 ( .A0(n370), .A1(n367), .A2(n366), .Z(n697));
Q_XOR3 U672 ( .A0(n364), .A1(n363), .A2(n361), .Z(n698));
Q_XOR3 U673 ( .A0(n359), .A1(n356), .A2(n691), .Z(n699));
Q_XOR3 U674 ( .A0(n692), .A1(n693), .A2(n694), .Z(n700));
Q_XOR3 U675 ( .A0(n765), .A1(n695), .A2(n696), .Z(n701));
Q_XOR3 U676 ( .A0(n697), .A1(n698), .A2(n699), .Z(n702));
Q_XOR3 U677 ( .A0(n700), .A1(n701), .A2(n702), .Z(n703));
Q_XOR3 U678 ( .A0(n526), .A1(n419), .A2(n418), .Z(n704));
Q_XOR3 U679 ( .A0(n417), .A1(n415), .A2(n411), .Z(n705));
Q_XOR3 U680 ( .A0(n404), .A1(n401), .A2(n400), .Z(n706));
Q_XOR3 U681 ( .A0(n399), .A1(n395), .A2(n394), .Z(n707));
Q_XOR3 U682 ( .A0(n382), .A1(n381), .A2(n380), .Z(n708));
Q_XOR3 U683 ( .A0(n378), .A1(n375), .A2(n372), .Z(n709));
Q_XOR3 U684 ( .A0(n371), .A1(n368), .A2(n367), .Z(n710));
Q_XOR3 U685 ( .A0(n365), .A1(n364), .A2(n362), .Z(n711));
Q_XOR3 U686 ( .A0(n360), .A1(n357), .A2(n356), .Z(n712));
Q_XOR3 U687 ( .A0(n704), .A1(n705), .A2(n706), .Z(n713));
Q_XOR3 U688 ( .A0(n707), .A1(n864), .A2(n708), .Z(n714));
Q_XOR3 U689 ( .A0(n709), .A1(n710), .A2(n711), .Z(n715));
Q_XOR3 U690 ( .A0(n712), .A1(n713), .A2(n714), .Z(n716));
Q_XOR2 U691 ( .A0(n715), .A1(n716), .Z(n717));
Q_XOR3 U692 ( .A0(n527), .A1(n419), .A2(n418), .Z(n718));
Q_XOR3 U693 ( .A0(n415), .A1(n414), .A2(n413), .Z(n719));
Q_XOR3 U694 ( .A0(n404), .A1(n403), .A2(n401), .Z(n720));
Q_XOR3 U695 ( .A0(n400), .A1(n399), .A2(n397), .Z(n721));
Q_XOR3 U696 ( .A0(n392), .A1(n390), .A2(n387), .Z(n722));
Q_XOR3 U697 ( .A0(n385), .A1(n382), .A2(n381), .Z(n723));
Q_XOR3 U698 ( .A0(n379), .A1(n378), .A2(n377), .Z(n724));
Q_XOR3 U699 ( .A0(n376), .A1(n375), .A2(n374), .Z(n725));
Q_XOR3 U700 ( .A0(n368), .A1(n367), .A2(n365), .Z(n726));
Q_XOR3 U701 ( .A0(n363), .A1(n357), .A2(n356), .Z(n727));
Q_XOR3 U702 ( .A0(n718), .A1(n719), .A2(n861), .Z(n728));
Q_XOR3 U703 ( .A0(n720), .A1(n721), .A2(n886), .Z(n729));
Q_XOR3 U704 ( .A0(n722), .A1(n723), .A2(n724), .Z(n730));
Q_XOR3 U705 ( .A0(n725), .A1(n726), .A2(n727), .Z(n731));
Q_XOR3 U706 ( .A0(n728), .A1(n729), .A2(n730), .Z(n732));
Q_XOR2 U707 ( .A0(n731), .A1(n732), .Z(n733));
Q_XOR3 U708 ( .A0(n528), .A1(n419), .A2(n413), .Z(n734));
Q_XOR3 U709 ( .A0(n411), .A1(n409), .A2(n408), .Z(n735));
Q_XOR3 U710 ( .A0(n406), .A1(n405), .A2(n403), .Z(n736));
Q_XOR3 U711 ( .A0(n398), .A1(n392), .A2(n391), .Z(n737));
Q_XOR3 U712 ( .A0(n386), .A1(n385), .A2(n384), .Z(n738));
Q_XOR3 U713 ( .A0(n382), .A1(n380), .A2(n379), .Z(n739));
Q_XOR3 U714 ( .A0(n372), .A1(n368), .A2(n367), .Z(n740));
Q_XOR3 U715 ( .A0(n364), .A1(n361), .A2(n357), .Z(n741));
Q_XOR3 U716 ( .A0(n356), .A1(n734), .A2(n735), .Z(n742));
Q_XOR3 U717 ( .A0(n736), .A1(n965), .A2(n737), .Z(n743));
Q_XOR3 U718 ( .A0(n951), .A1(n738), .A2(n739), .Z(n744));
Q_XOR3 U719 ( .A0(n1003), .A1(n740), .A2(n741), .Z(n745));
Q_XOR3 U720 ( .A0(n742), .A1(n743), .A2(n744), .Z(n746));
Q_XOR2 U721 ( .A0(n745), .A1(n746), .Z(n747));
Q_XOR3 U722 ( .A0(n529), .A1(n416), .A2(n415), .Z(n748));
Q_XOR3 U723 ( .A0(n406), .A1(n403), .A2(n401), .Z(n749));
Q_XOR3 U724 ( .A0(n394), .A1(n391), .A2(n387), .Z(n750));
Q_XOR3 U725 ( .A0(n386), .A1(n384), .A2(n381), .Z(n751));
Q_XOR3 U726 ( .A0(n380), .A1(n378), .A2(n372), .Z(n752));
Q_XOR3 U727 ( .A0(n368), .A1(n367), .A2(n366), .Z(n753));
Q_XOR3 U728 ( .A0(n365), .A1(n362), .A2(n361), .Z(n754));
Q_XOR3 U729 ( .A0(n357), .A1(n356), .A2(n748), .Z(n755));
Q_XOR3 U730 ( .A0(n883), .A1(n915), .A2(n749), .Z(n756));
Q_XOR3 U731 ( .A0(n846), .A1(n750), .A2(n751), .Z(n757));
Q_XOR3 U732 ( .A0(n752), .A1(n753), .A2(n754), .Z(n758));
Q_XOR3 U733 ( .A0(n755), .A1(n756), .A2(n757), .Z(n759));
Q_XOR2 U734 ( .A0(n758), .A1(n759), .Z(n760));
Q_XOR3 U735 ( .A0(n530), .A1(n417), .A2(n416), .Z(n761));
Q_XOR3 U736 ( .A0(n407), .A1(n404), .A2(n402), .Z(n762));
Q_XOR3 U737 ( .A0(n401), .A1(n398), .A2(n396), .Z(n763));
Q_XOR3 U738 ( .A0(n395), .A1(n392), .A2(n388), .Z(n764));
Q_XOR3 U739 ( .A0(n387), .A1(n385), .A2(n382), .Z(n765));
Q_XOR3 U740 ( .A0(n381), .A1(n379), .A2(n373), .Z(n766));
Q_XOR3 U741 ( .A0(n369), .A1(n368), .A2(n367), .Z(n767));
Q_XOR3 U742 ( .A0(n366), .A1(n363), .A2(n362), .Z(n768));
Q_XOR3 U743 ( .A0(n358), .A1(n357), .A2(n761), .Z(n769));
Q_XOR3 U744 ( .A0(n899), .A1(n931), .A2(n762), .Z(n770));
Q_XOR3 U745 ( .A0(n763), .A1(n764), .A2(n765), .Z(n771));
Q_XOR3 U746 ( .A0(n766), .A1(n767), .A2(n768), .Z(n772));
Q_XOR3 U747 ( .A0(n769), .A1(n770), .A2(n771), .Z(n773));
Q_XOR2 U748 ( .A0(n772), .A1(n773), .Z(n774));
Q_XOR3 U749 ( .A0(n531), .A1(n418), .A2(n417), .Z(n775));
Q_XOR3 U750 ( .A0(n415), .A1(n413), .A2(n412), .Z(n776));
Q_XOR3 U751 ( .A0(n408), .A1(n405), .A2(n403), .Z(n777));
Q_XOR3 U752 ( .A0(n402), .A1(n399), .A2(n397), .Z(n778));
Q_XOR3 U753 ( .A0(n396), .A1(n393), .A2(n389), .Z(n779));
Q_XOR3 U754 ( .A0(n382), .A1(n380), .A2(n374), .Z(n780));
Q_XOR3 U755 ( .A0(n370), .A1(n369), .A2(n368), .Z(n781));
Q_XOR3 U756 ( .A0(n367), .A1(n364), .A2(n363), .Z(n782));
Q_XOR3 U757 ( .A0(n359), .A1(n358), .A2(n775), .Z(n783));
Q_XOR3 U758 ( .A0(n776), .A1(n947), .A2(n777), .Z(n784));
Q_XOR3 U759 ( .A0(n778), .A1(n779), .A2(n864), .Z(n785));
Q_XOR3 U760 ( .A0(n780), .A1(n781), .A2(n782), .Z(n786));
Q_XOR3 U761 ( .A0(n783), .A1(n784), .A2(n785), .Z(n787));
Q_XOR2 U762 ( .A0(n786), .A1(n787), .Z(n788));
Q_XOR3 U763 ( .A0(n532), .A1(n419), .A2(n418), .Z(n789));
Q_XOR3 U764 ( .A0(n416), .A1(n414), .A2(n413), .Z(n790));
Q_XOR3 U765 ( .A0(n409), .A1(n406), .A2(n404), .Z(n791));
Q_XOR3 U766 ( .A0(n403), .A1(n400), .A2(n398), .Z(n792));
Q_XOR3 U767 ( .A0(n397), .A1(n394), .A2(n390), .Z(n793));
Q_XOR3 U768 ( .A0(n389), .A1(n387), .A2(n384), .Z(n794));
Q_XOR3 U769 ( .A0(n383), .A1(n381), .A2(n375), .Z(n795));
Q_XOR3 U770 ( .A0(n371), .A1(n370), .A2(n369), .Z(n796));
Q_XOR3 U771 ( .A0(n368), .A1(n365), .A2(n364), .Z(n797));
Q_XOR3 U772 ( .A0(n360), .A1(n359), .A2(n789), .Z(n798));
Q_XOR3 U773 ( .A0(n790), .A1(n963), .A2(n791), .Z(n799));
Q_XOR3 U774 ( .A0(n792), .A1(n793), .A2(n794), .Z(n800));
Q_XOR3 U775 ( .A0(n795), .A1(n796), .A2(n797), .Z(n801));
Q_XOR3 U776 ( .A0(n798), .A1(n799), .A2(n800), .Z(n802));
Q_XOR2 U777 ( .A0(n801), .A1(n802), .Z(n803));
Q_XOR3 U778 ( .A0(n533), .A1(n419), .A2(n417), .Z(n804));
Q_XOR3 U779 ( .A0(n416), .A1(n410), .A2(n408), .Z(n805));
Q_XOR3 U780 ( .A0(n407), .A1(n405), .A2(n403), .Z(n806));
Q_XOR3 U781 ( .A0(n402), .A1(n401), .A2(n398), .Z(n807));
Q_XOR3 U782 ( .A0(n397), .A1(n394), .A2(n393), .Z(n808));
Q_XOR3 U783 ( .A0(n388), .A1(n383), .A2(n382), .Z(n809));
Q_XOR3 U784 ( .A0(n378), .A1(n377), .A2(n376), .Z(n810));
Q_XOR3 U785 ( .A0(n375), .A1(n374), .A2(n373), .Z(n811));
Q_XOR3 U786 ( .A0(n365), .A1(n360), .A2(n358), .Z(n812));
Q_XOR3 U787 ( .A0(n356), .A1(n804), .A2(n805), .Z(n813));
Q_XOR3 U788 ( .A0(n806), .A1(n807), .A2(n808), .Z(n814));
Q_XOR3 U789 ( .A0(n863), .A1(n809), .A2(n810), .Z(n815));
Q_XOR3 U790 ( .A0(n811), .A1(n987), .A2(n812), .Z(n816));
Q_XOR3 U791 ( .A0(n813), .A1(n814), .A2(n815), .Z(n817));
Q_XOR2 U792 ( .A0(n816), .A1(n817), .Z(n818));
Q_XOR3 U793 ( .A0(n534), .A1(n418), .A2(n417), .Z(n819));
Q_XOR3 U794 ( .A0(n416), .A1(n415), .A2(n414), .Z(n820));
Q_XOR3 U795 ( .A0(n413), .A1(n412), .A2(n409), .Z(n821));
Q_XOR3 U796 ( .A0(n406), .A1(n398), .A2(n397), .Z(n822));
Q_XOR3 U797 ( .A0(n385), .A1(n379), .A2(n376), .Z(n823));
Q_XOR3 U798 ( .A0(n373), .A1(n371), .A2(n369), .Z(n824));
Q_XOR3 U799 ( .A0(n368), .A1(n367), .A2(n359), .Z(n825));
Q_XOR3 U800 ( .A0(n358), .A1(n357), .A2(n356), .Z(n826));
Q_XOR3 U801 ( .A0(n819), .A1(n820), .A2(n821), .Z(n827));
Q_XOR3 U802 ( .A0(n822), .A1(n823), .A2(n824), .Z(n828));
Q_XOR3 U803 ( .A0(n825), .A1(n826), .A2(n827), .Z(n829));
Q_XOR2 U804 ( .A0(n828), .A1(n829), .Z(n830));
Q_XOR3 U805 ( .A0(n535), .A1(n419), .A2(n418), .Z(n831));
Q_XOR3 U806 ( .A0(n417), .A1(n416), .A2(n415), .Z(n832));
Q_XOR3 U807 ( .A0(n414), .A1(n413), .A2(n410), .Z(n833));
Q_XOR3 U808 ( .A0(n407), .A1(n399), .A2(n398), .Z(n834));
Q_XOR3 U809 ( .A0(n386), .A1(n380), .A2(n377), .Z(n835));
Q_XOR3 U810 ( .A0(n374), .A1(n372), .A2(n370), .Z(n836));
Q_XOR3 U811 ( .A0(n369), .A1(n368), .A2(n360), .Z(n837));
Q_XOR3 U812 ( .A0(n359), .A1(n358), .A2(n357), .Z(n838));
Q_XOR3 U813 ( .A0(n356), .A1(n831), .A2(n832), .Z(n839));
Q_XOR3 U814 ( .A0(n833), .A1(n834), .A2(n835), .Z(n840));
Q_XOR3 U815 ( .A0(n836), .A1(n837), .A2(n838), .Z(n841));
Q_XOR3 U816 ( .A0(n839), .A1(n840), .A2(n841), .Z(n842));
Q_XOR3 U817 ( .A0(n536), .A1(n419), .A2(n418), .Z(n843));
Q_XOR3 U818 ( .A0(n417), .A1(n413), .A2(n412), .Z(n844));
Q_XOR3 U819 ( .A0(n404), .A1(n403), .A2(n402), .Z(n845));
Q_XOR3 U820 ( .A0(n400), .A1(n397), .A2(n395), .Z(n846));
Q_XOR3 U821 ( .A0(n394), .A1(n393), .A2(n392), .Z(n847));
Q_XOR3 U822 ( .A0(n390), .A1(n389), .A2(n387), .Z(n848));
Q_XOR3 U823 ( .A0(n385), .A1(n384), .A2(n383), .Z(n849));
Q_XOR3 U824 ( .A0(n381), .A1(n377), .A2(n374), .Z(n850));
Q_XOR3 U825 ( .A0(n372), .A1(n371), .A2(n370), .Z(n851));
Q_XOR3 U826 ( .A0(n367), .A1(n366), .A2(n360), .Z(n852));
Q_XOR3 U827 ( .A0(n359), .A1(n357), .A2(n356), .Z(n853));
Q_XOR3 U828 ( .A0(n843), .A1(n844), .A2(n845), .Z(n854));
Q_XOR3 U829 ( .A0(n846), .A1(n847), .A2(n848), .Z(n855));
Q_XOR3 U830 ( .A0(n849), .A1(n850), .A2(n851), .Z(n856));
Q_XOR3 U831 ( .A0(n852), .A1(n853), .A2(n854), .Z(n857));
Q_XOR3 U832 ( .A0(n855), .A1(n856), .A2(n857), .Z(n858));
Q_XOR3 U833 ( .A0(n537), .A1(n419), .A2(n418), .Z(n859));
Q_XOR3 U834 ( .A0(n416), .A1(n415), .A2(n412), .Z(n860));
Q_XOR3 U835 ( .A0(n411), .A1(n408), .A2(n405), .Z(n861));
Q_XOR3 U836 ( .A0(n402), .A1(n401), .A2(n399), .Z(n862));
Q_XOR3 U837 ( .A0(n392), .A1(n391), .A2(n389), .Z(n863));
Q_XOR3 U838 ( .A0(n388), .A1(n386), .A2(n383), .Z(n864));
Q_XOR3 U839 ( .A0(n382), .A1(n377), .A2(n374), .Z(n865));
Q_XOR3 U840 ( .A0(n366), .A1(n360), .A2(n357), .Z(n866));
Q_XOR3 U841 ( .A0(n859), .A1(n860), .A2(n861), .Z(n867));
Q_XOR3 U842 ( .A0(n862), .A1(n917), .A2(n863), .Z(n868));
Q_XOR3 U843 ( .A0(n864), .A1(n865), .A2(n922), .Z(n869));
Q_XOR3 U844 ( .A0(n866), .A1(n867), .A2(n868), .Z(n870));
Q_XOR2 U845 ( .A0(n869), .A1(n870), .Z(n871));
Q_XOR3 U846 ( .A0(n538), .A1(n419), .A2(n417), .Z(n872));
Q_XOR3 U847 ( .A0(n415), .A1(n414), .A2(n411), .Z(n873));
Q_XOR3 U848 ( .A0(n409), .A1(n408), .A2(n406), .Z(n874));
Q_XOR3 U849 ( .A0(n404), .A1(n400), .A2(n398), .Z(n875));
Q_XOR3 U850 ( .A0(n395), .A1(n394), .A2(n387), .Z(n876));
Q_XOR3 U851 ( .A0(n385), .A1(n377), .A2(n374), .Z(n877));
Q_XOR3 U852 ( .A0(n373), .A1(n370), .A2(n366), .Z(n878));
Q_XOR3 U853 ( .A0(n872), .A1(n873), .A2(n874), .Z(n879));
Q_XOR3 U854 ( .A0(n875), .A1(n876), .A2(n877), .Z(n880));
Q_XOR3 U855 ( .A0(n878), .A1(n879), .A2(n880), .Z(n881));
Q_XOR3 U856 ( .A0(n539), .A1(n418), .A2(n414), .Z(n882));
Q_XOR3 U857 ( .A0(n413), .A1(n411), .A2(n410), .Z(n883));
Q_XOR3 U858 ( .A0(n405), .A1(n404), .A2(n403), .Z(n884));
Q_XOR3 U859 ( .A0(n402), .A1(n401), .A2(n397), .Z(n885));
Q_XOR3 U860 ( .A0(n396), .A1(n394), .A2(n393), .Z(n886));
Q_XOR3 U861 ( .A0(n392), .A1(n390), .A2(n389), .Z(n887));
Q_XOR3 U862 ( .A0(n388), .A1(n386), .A2(n385), .Z(n888));
Q_XOR3 U863 ( .A0(n384), .A1(n383), .A2(n377), .Z(n889));
Q_XOR3 U864 ( .A0(n373), .A1(n372), .A2(n371), .Z(n890));
Q_XOR3 U865 ( .A0(n369), .A1(n366), .A2(n361), .Z(n891));
Q_XOR3 U866 ( .A0(n358), .A1(n356), .A2(n882), .Z(n892));
Q_XOR3 U867 ( .A0(n883), .A1(n915), .A2(n884), .Z(n893));
Q_XOR3 U868 ( .A0(n885), .A1(n886), .A2(n887), .Z(n894));
Q_XOR3 U869 ( .A0(n888), .A1(n889), .A2(n890), .Z(n895));
Q_XOR3 U870 ( .A0(n891), .A1(n892), .A2(n893), .Z(n896));
Q_XOR3 U871 ( .A0(n894), .A1(n895), .A2(n896), .Z(n897));
Q_XOR3 U872 ( .A0(n540), .A1(n419), .A2(n415), .Z(n898));
Q_XOR3 U873 ( .A0(n414), .A1(n412), .A2(n411), .Z(n899));
Q_XOR3 U874 ( .A0(n406), .A1(n405), .A2(n404), .Z(n900));
Q_XOR3 U875 ( .A0(n403), .A1(n402), .A2(n398), .Z(n901));
Q_XOR3 U876 ( .A0(n397), .A1(n395), .A2(n394), .Z(n902));
Q_XOR3 U877 ( .A0(n393), .A1(n391), .A2(n390), .Z(n903));
Q_XOR3 U878 ( .A0(n389), .A1(n387), .A2(n386), .Z(n904));
Q_XOR3 U879 ( .A0(n385), .A1(n384), .A2(n378), .Z(n905));
Q_XOR3 U880 ( .A0(n374), .A1(n373), .A2(n372), .Z(n906));
Q_XOR3 U881 ( .A0(n370), .A1(n367), .A2(n362), .Z(n907));
Q_XOR3 U882 ( .A0(n359), .A1(n357), .A2(n898), .Z(n908));
Q_XOR3 U883 ( .A0(n899), .A1(n931), .A2(n900), .Z(n909));
Q_XOR3 U884 ( .A0(n901), .A1(n902), .A2(n903), .Z(n910));
Q_XOR3 U885 ( .A0(n904), .A1(n905), .A2(n906), .Z(n911));
Q_XOR3 U886 ( .A0(n907), .A1(n908), .A2(n909), .Z(n912));
Q_XOR3 U887 ( .A0(n910), .A1(n911), .A2(n912), .Z(n913));
Q_XOR3 U888 ( .A0(n541), .A1(n414), .A2(n410), .Z(n914));
Q_XOR3 U889 ( .A0(n409), .A1(n408), .A2(n407), .Z(n915));
Q_XOR3 U890 ( .A0(n406), .A1(n405), .A2(n402), .Z(n916));
Q_XOR3 U891 ( .A0(n398), .A1(n397), .A2(n396), .Z(n917));
Q_XOR3 U892 ( .A0(n393), .A1(n391), .A2(n389), .Z(n918));
Q_XOR3 U893 ( .A0(n388), .A1(n387), .A2(n386), .Z(n919));
Q_XOR3 U894 ( .A0(n384), .A1(n383), .A2(n379), .Z(n920));
Q_XOR3 U895 ( .A0(n378), .A1(n377), .A2(n372), .Z(n921));
Q_XOR3 U896 ( .A0(n371), .A1(n369), .A2(n368), .Z(n922));
Q_XOR3 U897 ( .A0(n367), .A1(n366), .A2(n363), .Z(n923));
Q_XOR3 U898 ( .A0(n361), .A1(n360), .A2(n914), .Z(n924));
Q_XOR3 U899 ( .A0(n915), .A1(n916), .A2(n917), .Z(n925));
Q_XOR3 U900 ( .A0(n918), .A1(n919), .A2(n920), .Z(n926));
Q_XOR3 U901 ( .A0(n921), .A1(n922), .A2(n923), .Z(n927));
Q_XOR3 U902 ( .A0(n924), .A1(n925), .A2(n926), .Z(n928));
Q_XOR2 U903 ( .A0(n927), .A1(n928), .Z(n929));
Q_XOR3 U904 ( .A0(n542), .A1(n415), .A2(n411), .Z(n930));
Q_XOR3 U905 ( .A0(n410), .A1(n409), .A2(n408), .Z(n931));
Q_XOR3 U906 ( .A0(n407), .A1(n406), .A2(n403), .Z(n932));
Q_XOR3 U907 ( .A0(n399), .A1(n398), .A2(n397), .Z(n933));
Q_XOR3 U908 ( .A0(n394), .A1(n392), .A2(n390), .Z(n934));
Q_XOR3 U909 ( .A0(n389), .A1(n388), .A2(n387), .Z(n935));
Q_XOR3 U910 ( .A0(n385), .A1(n384), .A2(n380), .Z(n936));
Q_XOR3 U911 ( .A0(n379), .A1(n378), .A2(n373), .Z(n937));
Q_XOR3 U912 ( .A0(n372), .A1(n370), .A2(n369), .Z(n938));
Q_XOR3 U913 ( .A0(n368), .A1(n367), .A2(n364), .Z(n939));
Q_XOR3 U914 ( .A0(n362), .A1(n361), .A2(n356), .Z(n940));
Q_XOR3 U915 ( .A0(n930), .A1(n931), .A2(n932), .Z(n941));
Q_XOR3 U916 ( .A0(n933), .A1(n934), .A2(n935), .Z(n942));
Q_XOR3 U917 ( .A0(n936), .A1(n937), .A2(n938), .Z(n943));
Q_XOR3 U918 ( .A0(n939), .A1(n940), .A2(n941), .Z(n944));
Q_XOR3 U919 ( .A0(n942), .A1(n943), .A2(n944), .Z(n945));
Q_XOR3 U920 ( .A0(n543), .A1(n416), .A2(n412), .Z(n946));
Q_XOR3 U921 ( .A0(n411), .A1(n410), .A2(n409), .Z(n947));
Q_XOR3 U922 ( .A0(n408), .A1(n407), .A2(n404), .Z(n948));
Q_XOR3 U923 ( .A0(n400), .A1(n399), .A2(n398), .Z(n949));
Q_XOR3 U924 ( .A0(n395), .A1(n393), .A2(n391), .Z(n950));
Q_XOR3 U925 ( .A0(n390), .A1(n389), .A2(n388), .Z(n951));
Q_XOR3 U926 ( .A0(n386), .A1(n385), .A2(n381), .Z(n952));
Q_XOR3 U927 ( .A0(n380), .A1(n379), .A2(n374), .Z(n953));
Q_XOR3 U928 ( .A0(n373), .A1(n371), .A2(n370), .Z(n954));
Q_XOR3 U929 ( .A0(n369), .A1(n368), .A2(n365), .Z(n955));
Q_XOR3 U930 ( .A0(n363), .A1(n362), .A2(n357), .Z(n956));
Q_XOR3 U931 ( .A0(n946), .A1(n947), .A2(n948), .Z(n957));
Q_XOR3 U932 ( .A0(n949), .A1(n950), .A2(n951), .Z(n958));
Q_XOR3 U933 ( .A0(n952), .A1(n953), .A2(n954), .Z(n959));
Q_XOR3 U934 ( .A0(n955), .A1(n956), .A2(n957), .Z(n960));
Q_XOR3 U935 ( .A0(n958), .A1(n959), .A2(n960), .Z(n961));
Q_XOR3 U936 ( .A0(n544), .A1(n417), .A2(n413), .Z(n962));
Q_XOR3 U937 ( .A0(n412), .A1(n411), .A2(n410), .Z(n963));
Q_XOR3 U938 ( .A0(n409), .A1(n408), .A2(n405), .Z(n964));
Q_XOR3 U939 ( .A0(n401), .A1(n400), .A2(n399), .Z(n965));
Q_XOR3 U940 ( .A0(n396), .A1(n394), .A2(n392), .Z(n966));
Q_XOR3 U941 ( .A0(n391), .A1(n390), .A2(n389), .Z(n967));
Q_XOR3 U942 ( .A0(n387), .A1(n386), .A2(n382), .Z(n968));
Q_XOR3 U943 ( .A0(n381), .A1(n380), .A2(n375), .Z(n969));
Q_XOR3 U944 ( .A0(n374), .A1(n372), .A2(n371), .Z(n970));
Q_XOR3 U945 ( .A0(n370), .A1(n369), .A2(n366), .Z(n971));
Q_XOR3 U946 ( .A0(n364), .A1(n363), .A2(n358), .Z(n972));
Q_XOR3 U947 ( .A0(n962), .A1(n963), .A2(n964), .Z(n973));
Q_XOR3 U948 ( .A0(n965), .A1(n966), .A2(n967), .Z(n974));
Q_XOR3 U949 ( .A0(n968), .A1(n969), .A2(n970), .Z(n975));
Q_XOR3 U950 ( .A0(n971), .A1(n972), .A2(n973), .Z(n976));
Q_XOR3 U951 ( .A0(n974), .A1(n975), .A2(n976), .Z(n977));
Q_XOR3 U952 ( .A0(n545), .A1(n418), .A2(n414), .Z(n978));
Q_XOR3 U953 ( .A0(n413), .A1(n412), .A2(n411), .Z(n979));
Q_XOR3 U954 ( .A0(n410), .A1(n409), .A2(n406), .Z(n980));
Q_XOR3 U955 ( .A0(n402), .A1(n401), .A2(n400), .Z(n981));
Q_XOR3 U956 ( .A0(n397), .A1(n395), .A2(n393), .Z(n982));
Q_XOR3 U957 ( .A0(n392), .A1(n391), .A2(n390), .Z(n983));
Q_XOR3 U958 ( .A0(n388), .A1(n387), .A2(n383), .Z(n984));
Q_XOR3 U959 ( .A0(n382), .A1(n381), .A2(n376), .Z(n985));
Q_XOR3 U960 ( .A0(n375), .A1(n373), .A2(n372), .Z(n986));
Q_XOR3 U961 ( .A0(n371), .A1(n370), .A2(n367), .Z(n987));
Q_XOR3 U962 ( .A0(n365), .A1(n364), .A2(n359), .Z(n988));
Q_XOR3 U963 ( .A0(n356), .A1(n978), .A2(n979), .Z(n989));
Q_XOR3 U964 ( .A0(n980), .A1(n981), .A2(n982), .Z(n990));
Q_XOR3 U965 ( .A0(n983), .A1(n984), .A2(n985), .Z(n991));
Q_XOR3 U966 ( .A0(n986), .A1(n987), .A2(n988), .Z(n992));
Q_XOR3 U967 ( .A0(n989), .A1(n990), .A2(n991), .Z(n993));
Q_XOR2 U968 ( .A0(n992), .A1(n993), .Z(n994));
Q_XOR3 U969 ( .A0(n546), .A1(n419), .A2(n415), .Z(n995));
Q_XOR3 U970 ( .A0(n414), .A1(n413), .A2(n412), .Z(n996));
Q_XOR3 U971 ( .A0(n411), .A1(n410), .A2(n407), .Z(n997));
Q_XOR3 U972 ( .A0(n403), .A1(n402), .A2(n401), .Z(n998));
Q_XOR3 U973 ( .A0(n398), .A1(n396), .A2(n394), .Z(n999));
Q_XOR3 U974 ( .A0(n393), .A1(n392), .A2(n391), .Z(n1000));
Q_XOR3 U975 ( .A0(n389), .A1(n388), .A2(n384), .Z(n1001));
Q_XOR3 U976 ( .A0(n383), .A1(n382), .A2(n377), .Z(n1002));
Q_XOR3 U977 ( .A0(n376), .A1(n374), .A2(n373), .Z(n1003));
Q_XOR3 U978 ( .A0(n372), .A1(n371), .A2(n368), .Z(n1004));
Q_XOR3 U979 ( .A0(n366), .A1(n365), .A2(n360), .Z(n1005));
Q_XOR3 U980 ( .A0(n357), .A1(n995), .A2(n996), .Z(n1006));
Q_XOR3 U981 ( .A0(n997), .A1(n998), .A2(n999), .Z(n1007));
Q_XOR3 U982 ( .A0(n1000), .A1(n1001), .A2(n1002), .Z(n1008));
Q_XOR3 U983 ( .A0(n1003), .A1(n1004), .A2(n1005), .Z(n1009));
Q_XOR3 U984 ( .A0(n1006), .A1(n1007), .A2(n1008), .Z(n1010));
Q_XOR2 U985 ( .A0(n1009), .A1(n1010), .Z(n1011));
Q_FDP1 \crc_r_REG[31] ( .CK(clk), .R(rst_n), .D(n1012), .Q(crc_r[31]), .QN(n2));
Q_MX03 U987 ( .S0(init), .S1(n1044), .A0(n1011), .A1(init_value[31]), .A2(crc_r[31]), .Z(n1012));
Q_FDP1 \crc_r_REG[30] ( .CK(clk), .R(rst_n), .D(n1013), .Q(crc_r[30]), .QN(n3));
Q_MX03 U989 ( .S0(init), .S1(n1044), .A0(n994), .A1(init_value[30]), .A2(crc_r[30]), .Z(n1013));
Q_FDP1 \crc_r_REG[29] ( .CK(clk), .R(rst_n), .D(n1014), .Q(crc_r[29]), .QN(n4));
Q_MX03 U991 ( .S0(init), .S1(n1044), .A0(n977), .A1(init_value[29]), .A2(crc_r[29]), .Z(n1014));
Q_FDP1 \crc_r_REG[28] ( .CK(clk), .R(rst_n), .D(n1015), .Q(crc_r[28]), .QN(n5));
Q_MX03 U993 ( .S0(init), .S1(n1044), .A0(n961), .A1(init_value[28]), .A2(crc_r[28]), .Z(n1015));
Q_FDP1 \crc_r_REG[27] ( .CK(clk), .R(rst_n), .D(n1016), .Q(crc_r[27]), .QN(n6));
Q_MX03 U995 ( .S0(init), .S1(n1044), .A0(n945), .A1(init_value[27]), .A2(crc_r[27]), .Z(n1016));
Q_FDP1 \crc_r_REG[26] ( .CK(clk), .R(rst_n), .D(n1017), .Q(crc_r[26]), .QN(n7));
Q_MX03 U997 ( .S0(init), .S1(n1044), .A0(n929), .A1(init_value[26]), .A2(crc_r[26]), .Z(n1017));
Q_FDP1 \crc_r_REG[25] ( .CK(clk), .R(rst_n), .D(n1018), .Q(crc_r[25]), .QN(n8));
Q_MX03 U999 ( .S0(init), .S1(n1044), .A0(n913), .A1(init_value[25]), .A2(crc_r[25]), .Z(n1018));
Q_FDP1 \crc_r_REG[24] ( .CK(clk), .R(rst_n), .D(n1019), .Q(crc_r[24]), .QN(n9));
Q_MX03 U1001 ( .S0(init), .S1(n1044), .A0(n897), .A1(init_value[24]), .A2(crc_r[24]), .Z(n1019));
Q_FDP1 \crc_r_REG[23] ( .CK(clk), .R(rst_n), .D(n1020), .Q(crc_r[23]), .QN(n10));
Q_MX03 U1003 ( .S0(init), .S1(n1044), .A0(n881), .A1(init_value[23]), .A2(crc_r[23]), .Z(n1020));
Q_FDP1 \crc_r_REG[22] ( .CK(clk), .R(rst_n), .D(n1021), .Q(crc_r[22]), .QN(n11));
Q_MX03 U1005 ( .S0(init), .S1(n1044), .A0(n871), .A1(init_value[22]), .A2(crc_r[22]), .Z(n1021));
Q_FDP1 \crc_r_REG[21] ( .CK(clk), .R(rst_n), .D(n1022), .Q(crc_r[21]), .QN(n12));
Q_MX03 U1007 ( .S0(init), .S1(n1044), .A0(n858), .A1(init_value[21]), .A2(crc_r[21]), .Z(n1022));
Q_FDP1 \crc_r_REG[20] ( .CK(clk), .R(rst_n), .D(n1023), .Q(crc_r[20]), .QN(n13));
Q_MX03 U1009 ( .S0(init), .S1(n1044), .A0(n842), .A1(init_value[20]), .A2(crc_r[20]), .Z(n1023));
Q_FDP1 \crc_r_REG[19] ( .CK(clk), .R(rst_n), .D(n1024), .Q(crc_r[19]), .QN(n14));
Q_MX03 U1011 ( .S0(init), .S1(n1044), .A0(n830), .A1(init_value[19]), .A2(crc_r[19]), .Z(n1024));
Q_FDP1 \crc_r_REG[18] ( .CK(clk), .R(rst_n), .D(n1025), .Q(crc_r[18]), .QN(n15));
Q_MX03 U1013 ( .S0(init), .S1(n1044), .A0(n818), .A1(init_value[18]), .A2(crc_r[18]), .Z(n1025));
Q_FDP1 \crc_r_REG[17] ( .CK(clk), .R(rst_n), .D(n1026), .Q(crc_r[17]), .QN(n16));
Q_MX03 U1015 ( .S0(init), .S1(n1044), .A0(n803), .A1(init_value[17]), .A2(crc_r[17]), .Z(n1026));
Q_FDP1 \crc_r_REG[16] ( .CK(clk), .R(rst_n), .D(n1027), .Q(crc_r[16]), .QN(n17));
Q_MX03 U1017 ( .S0(init), .S1(n1044), .A0(n788), .A1(init_value[16]), .A2(crc_r[16]), .Z(n1027));
Q_FDP1 \crc_r_REG[15] ( .CK(clk), .R(rst_n), .D(n1028), .Q(crc_r[15]), .QN(n18));
Q_MX03 U1019 ( .S0(init), .S1(n1044), .A0(n774), .A1(init_value[15]), .A2(crc_r[15]), .Z(n1028));
Q_FDP1 \crc_r_REG[14] ( .CK(clk), .R(rst_n), .D(n1029), .Q(crc_r[14]), .QN(n19));
Q_MX03 U1021 ( .S0(init), .S1(n1044), .A0(n760), .A1(init_value[14]), .A2(crc_r[14]), .Z(n1029));
Q_FDP1 \crc_r_REG[13] ( .CK(clk), .R(rst_n), .D(n1030), .Q(crc_r[13]), .QN(n20));
Q_MX03 U1023 ( .S0(init), .S1(n1044), .A0(n747), .A1(init_value[13]), .A2(crc_r[13]), .Z(n1030));
Q_FDP1 \crc_r_REG[12] ( .CK(clk), .R(rst_n), .D(n1031), .Q(crc_r[12]), .QN(n21));
Q_MX03 U1025 ( .S0(init), .S1(n1044), .A0(n733), .A1(init_value[12]), .A2(crc_r[12]), .Z(n1031));
Q_FDP1 \crc_r_REG[11] ( .CK(clk), .R(rst_n), .D(n1032), .Q(crc_r[11]), .QN(n22));
Q_MX03 U1027 ( .S0(init), .S1(n1044), .A0(n717), .A1(init_value[11]), .A2(crc_r[11]), .Z(n1032));
Q_FDP1 \crc_r_REG[10] ( .CK(clk), .R(rst_n), .D(n1033), .Q(crc_r[10]), .QN(n23));
Q_MX03 U1029 ( .S0(init), .S1(n1044), .A0(n703), .A1(init_value[10]), .A2(crc_r[10]), .Z(n1033));
Q_FDP1 \crc_r_REG[9] ( .CK(clk), .R(rst_n), .D(n1034), .Q(crc_r[9]), .QN(n24));
Q_MX03 U1031 ( .S0(init), .S1(n1044), .A0(n690), .A1(init_value[9]), .A2(crc_r[9]), .Z(n1034));
Q_FDP1 \crc_r_REG[8] ( .CK(clk), .R(rst_n), .D(n1035), .Q(crc_r[8]), .QN(n25));
Q_MX03 U1033 ( .S0(init), .S1(n1044), .A0(n678), .A1(init_value[8]), .A2(crc_r[8]), .Z(n1035));
Q_FDP1 \crc_r_REG[7] ( .CK(clk), .R(rst_n), .D(n1036), .Q(crc_r[7]), .QN(n26));
Q_MX03 U1035 ( .S0(init), .S1(n1044), .A0(n665), .A1(init_value[7]), .A2(crc_r[7]), .Z(n1036));
Q_FDP1 \crc_r_REG[6] ( .CK(clk), .R(rst_n), .D(n1037), .Q(crc_r[6]), .QN(n27));
Q_MX03 U1037 ( .S0(init), .S1(n1044), .A0(n650), .A1(init_value[6]), .A2(crc_r[6]), .Z(n1037));
Q_FDP1 \crc_r_REG[5] ( .CK(clk), .R(rst_n), .D(n1038), .Q(crc_r[5]), .QN(n28));
Q_MX03 U1039 ( .S0(init), .S1(n1044), .A0(n635), .A1(init_value[5]), .A2(crc_r[5]), .Z(n1038));
Q_FDP1 \crc_r_REG[4] ( .CK(clk), .R(rst_n), .D(n1039), .Q(crc_r[4]), .QN(n29));
Q_MX03 U1041 ( .S0(init), .S1(n1044), .A0(n621), .A1(init_value[4]), .A2(crc_r[4]), .Z(n1039));
Q_FDP1 \crc_r_REG[3] ( .CK(clk), .R(rst_n), .D(n1040), .Q(crc_r[3]), .QN(n30));
Q_MX03 U1043 ( .S0(init), .S1(n1044), .A0(n603), .A1(init_value[3]), .A2(crc_r[3]), .Z(n1040));
Q_FDP1 \crc_r_REG[2] ( .CK(clk), .R(rst_n), .D(n1041), .Q(crc_r[2]), .QN(n31));
Q_MX03 U1045 ( .S0(init), .S1(n1044), .A0(n589), .A1(init_value[2]), .A2(crc_r[2]), .Z(n1041));
Q_FDP1 \crc_r_REG[1] ( .CK(clk), .R(rst_n), .D(n1042), .Q(crc_r[1]), .QN(n32));
Q_MX03 U1047 ( .S0(init), .S1(n1044), .A0(n574), .A1(init_value[1]), .A2(crc_r[1]), .Z(n1042));
Q_FDP1 \crc_r_REG[0] ( .CK(clk), .R(rst_n), .D(n1043), .Q(crc_r[0]), .QN(n33));
Q_MX03 U1049 ( .S0(init), .S1(n1044), .A0(n560), .A1(init_value[0]), .A2(crc_r[0]), .Z(n1043));
Q_NR02 U1050 ( .A0(init), .A1(data_valid), .Z(n1044));
Q_MX02 U1051 ( .S(data_vbits[5]), .A0(n427), .A1(n459), .Z(n1045));
Q_MX02 U1052 ( .S(data_vbits[4]), .A0(n443), .A1(n1045), .Z(n491));
Q_MX02 U1053 ( .S(data_vbits[5]), .A0(n426), .A1(n458), .Z(n1046));
Q_MX02 U1054 ( .S(data_vbits[4]), .A0(n442), .A1(n1046), .Z(n490));
Q_MX02 U1055 ( .S(data_vbits[5]), .A0(n425), .A1(n457), .Z(n1047));
Q_MX02 U1056 ( .S(data_vbits[4]), .A0(n441), .A1(n1047), .Z(n489));
Q_MX02 U1057 ( .S(data_vbits[5]), .A0(n424), .A1(n456), .Z(n1048));
Q_MX02 U1058 ( .S(data_vbits[4]), .A0(n440), .A1(n1048), .Z(n488));
Q_MX02 U1059 ( .S(data_vbits[5]), .A0(n423), .A1(n455), .Z(n1049));
Q_MX02 U1060 ( .S(data_vbits[4]), .A0(n439), .A1(n1049), .Z(n487));
Q_MX02 U1061 ( .S(data_vbits[5]), .A0(n422), .A1(n454), .Z(n1050));
Q_MX02 U1062 ( .S(data_vbits[4]), .A0(n438), .A1(n1050), .Z(n486));
Q_MX02 U1063 ( .S(data_vbits[5]), .A0(n421), .A1(n453), .Z(n1051));
Q_MX02 U1064 ( .S(data_vbits[4]), .A0(n437), .A1(n1051), .Z(n485));
Q_MX02 U1065 ( .S(data_vbits[5]), .A0(n420), .A1(n452), .Z(n1052));
Q_MX02 U1066 ( .S(data_vbits[4]), .A0(n436), .A1(n1052), .Z(n484));
Q_MX02 U1067 ( .S(data_vbits[6]), .A0(n181), .A1(n245), .Z(n1053));
Q_MX02 U1068 ( .S(data_vbits[5]), .A0(n213), .A1(n1053), .Z(n309));
Q_MX02 U1069 ( .S(data_vbits[6]), .A0(n180), .A1(n244), .Z(n1054));
Q_MX02 U1070 ( .S(data_vbits[5]), .A0(n212), .A1(n1054), .Z(n308));
Q_MX02 U1071 ( .S(data_vbits[6]), .A0(n179), .A1(n243), .Z(n1055));
Q_MX02 U1072 ( .S(data_vbits[5]), .A0(n211), .A1(n1055), .Z(n307));
Q_MX02 U1073 ( .S(data_vbits[6]), .A0(n178), .A1(n242), .Z(n1056));
Q_MX02 U1074 ( .S(data_vbits[5]), .A0(n210), .A1(n1056), .Z(n306));
Q_MX02 U1075 ( .S(data_vbits[6]), .A0(n177), .A1(n241), .Z(n1057));
Q_MX02 U1076 ( .S(data_vbits[5]), .A0(n209), .A1(n1057), .Z(n305));
Q_MX02 U1077 ( .S(data_vbits[6]), .A0(n176), .A1(n240), .Z(n1058));
Q_MX02 U1078 ( .S(data_vbits[5]), .A0(n208), .A1(n1058), .Z(n304));
Q_MX02 U1079 ( .S(data_vbits[6]), .A0(n175), .A1(n239), .Z(n1059));
Q_MX02 U1080 ( .S(data_vbits[5]), .A0(n207), .A1(n1059), .Z(n303));
Q_MX02 U1081 ( .S(data_vbits[6]), .A0(n174), .A1(n238), .Z(n1060));
Q_MX02 U1082 ( .S(data_vbits[5]), .A0(n206), .A1(n1060), .Z(n302));
Q_MX02 U1083 ( .S(data_vbits[6]), .A0(n173), .A1(n237), .Z(n1061));
Q_MX02 U1084 ( .S(data_vbits[5]), .A0(n205), .A1(n1061), .Z(n301));
Q_MX02 U1085 ( .S(data_vbits[6]), .A0(n172), .A1(n236), .Z(n1062));
Q_MX02 U1086 ( .S(data_vbits[5]), .A0(n204), .A1(n1062), .Z(n300));
Q_MX02 U1087 ( .S(data_vbits[6]), .A0(n171), .A1(n235), .Z(n1063));
Q_MX02 U1088 ( .S(data_vbits[5]), .A0(n203), .A1(n1063), .Z(n299));
Q_MX02 U1089 ( .S(data_vbits[6]), .A0(n170), .A1(n234), .Z(n1064));
Q_MX02 U1090 ( .S(data_vbits[5]), .A0(n202), .A1(n1064), .Z(n298));
Q_MX02 U1091 ( .S(data_vbits[6]), .A0(n169), .A1(n233), .Z(n1065));
Q_MX02 U1092 ( .S(data_vbits[5]), .A0(n201), .A1(n1065), .Z(n297));
Q_MX02 U1093 ( .S(data_vbits[6]), .A0(n168), .A1(n232), .Z(n1066));
Q_MX02 U1094 ( .S(data_vbits[5]), .A0(n200), .A1(n1066), .Z(n296));
Q_MX02 U1095 ( .S(data_vbits[6]), .A0(n167), .A1(n231), .Z(n1067));
Q_MX02 U1096 ( .S(data_vbits[5]), .A0(n199), .A1(n1067), .Z(n295));
Q_MX02 U1097 ( .S(data_vbits[6]), .A0(n166), .A1(n230), .Z(n1068));
Q_MX02 U1098 ( .S(data_vbits[5]), .A0(n198), .A1(n1068), .Z(n294));
Q_MX02 U1099 ( .S(data_vbits[6]), .A0(n165), .A1(n229), .Z(n1069));
Q_MX02 U1100 ( .S(data_vbits[5]), .A0(n197), .A1(n1069), .Z(n293));
Q_MX02 U1101 ( .S(data_vbits[6]), .A0(n164), .A1(n228), .Z(n1070));
Q_MX02 U1102 ( .S(data_vbits[5]), .A0(n196), .A1(n1070), .Z(n292));
Q_MX02 U1103 ( .S(data_vbits[6]), .A0(n163), .A1(n227), .Z(n1071));
Q_MX02 U1104 ( .S(data_vbits[5]), .A0(n195), .A1(n1071), .Z(n291));
Q_MX02 U1105 ( .S(data_vbits[6]), .A0(n162), .A1(n226), .Z(n1072));
Q_MX02 U1106 ( .S(data_vbits[5]), .A0(n194), .A1(n1072), .Z(n290));
Q_MX02 U1107 ( .S(data_vbits[6]), .A0(n161), .A1(n225), .Z(n1073));
Q_MX02 U1108 ( .S(data_vbits[5]), .A0(n193), .A1(n1073), .Z(n289));
Q_MX02 U1109 ( .S(data_vbits[6]), .A0(n160), .A1(n224), .Z(n1074));
Q_MX02 U1110 ( .S(data_vbits[5]), .A0(n192), .A1(n1074), .Z(n288));
Q_MX02 U1111 ( .S(data_vbits[6]), .A0(n159), .A1(n223), .Z(n1075));
Q_MX02 U1112 ( .S(data_vbits[5]), .A0(n191), .A1(n1075), .Z(n287));
Q_MX02 U1113 ( .S(data_vbits[6]), .A0(n158), .A1(n222), .Z(n1076));
Q_MX02 U1114 ( .S(data_vbits[5]), .A0(n190), .A1(n1076), .Z(n286));
Q_XNR2 U1115 ( .A0(data_vbytes[2]), .A1(data_vbytes[1]), .Z(n48));
endmodule
