architecture module of ixc_sfifo_bind_512_2 is

begin
end module;
