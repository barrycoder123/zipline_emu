
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_indirect_access_cntrl_v2_xcm126 ( clk, rst_n, wr_stb, reg_addr, 
	cmnd_op, cmnd_addr, cmnd_table_id, stat_code, stat_datawords, 
	stat_addr, stat_table_id, capability_lst, capability_type, enable, 
	.addr_limit( {\addr_limit[0][14] , \addr_limit[0][13] , 
	\addr_limit[0][12] , \addr_limit[0][11] , \addr_limit[0][10] , 
	\addr_limit[0][9] , \addr_limit[0][8] , \addr_limit[0][7] , 
	\addr_limit[0][6] , \addr_limit[0][5] , \addr_limit[0][4] , 
	\addr_limit[0][3] , \addr_limit[0][2] , \addr_limit[0][1] , 
	\addr_limit[0][0] } ), wr_dat, rd_dat, sw_cs, sw_ce, sw_we, sw_add, 
	sw_wdat, sw_rdat, sw_match, sw_aindex, grant, rsp, yield, reset);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input wr_stb;
input [10:0] reg_addr;
input [3:0] cmnd_op;
input [14:0] cmnd_addr;
input [0:0] cmnd_table_id;
output [2:0] stat_code;
output [4:0] stat_datawords;
output [14:0] stat_addr;
output [0:0] stat_table_id;
output [15:0] capability_lst;
output [3:0] capability_type;
output enable;
input \addr_limit[0][14] ;
input \addr_limit[0][13] ;
input \addr_limit[0][12] ;
input \addr_limit[0][11] ;
input \addr_limit[0][10] ;
input \addr_limit[0][9] ;
input \addr_limit[0][8] ;
input \addr_limit[0][7] ;
input \addr_limit[0][6] ;
input \addr_limit[0][5] ;
input \addr_limit[0][4] ;
input \addr_limit[0][3] ;
input \addr_limit[0][2] ;
input \addr_limit[0][1] ;
input \addr_limit[0][0] ;
input [63:0] wr_dat;
output [63:0] rd_dat;
output sw_cs;
output sw_ce;
output sw_we;
output [14:0] sw_add;
output [63:0] sw_wdat;
input [63:0] sw_rdat;
input sw_match;
input [13:0] sw_aindex;
input grant;
input rsp;
output yield;
output reset;
wire [0:2] _zy_simnet_stat_code_0_w$;
wire [0:4] _zy_simnet_stat_datawords_1_w$;
wire [0:14] _zy_simnet_stat_addr_2_w$;
wire _zy_simnet_stat_table_id_3_w$;
wire [0:15] _zy_simnet_capability_lst_4_w$;
wire [0:3] _zy_simnet_capability_type_5_w$;
wire _zy_simnet_enable_6_w$;
wire [0:63] _zy_simnet_rd_dat_7_w$;
wire _zy_simnet_sw_cs_8_w$;
wire _zy_simnet_sw_ce_9_w$;
wire _zy_simnet_sw_we_10_w$;
wire [0:14] _zy_simnet_sw_add_11_w$;
wire [0:63] _zy_simnet_sw_wdat_12_w$;
wire _zy_simnet_yield_13_w$;
wire _zy_simnet_reset_14_w$;
wire [3:0] cmnd;
wire init_r;
wire [0:0] inc_r;
wire init_inc_r;
wire sw_cs_r;
wire sw_ce_r;
wire rst_r;
wire rst_or_ini_r;
wire [14:0] rst_addr_r;
wire sw_we_r;
wire cmnd_rd_stb;
wire cmnd_wr_stb;
wire cmnd_ena_stb;
wire cmnd_dis_stb;
wire cmnd_rst_stb;
wire cmnd_ini_stb;
wire cmnd_inc_stb;
wire cmnd_sis_stb;
wire cmnd_tmo_stb;
wire cmnd_cmp_stb;
wire cmnd_issued;
wire ack_error;
wire unsupported_op;
wire [3:0] state_r;
wire [5:0] timer_r;
wire timeout;
wire sim_tmo_r;
wire [14:0] maxaddr;
wire badaddr;
wire igrant;
wire [2:0] stat;
supply0 n1;
supply1 n2;
Q_BUF U0 ( .A(n2), .Z(stat_datawords[0]));
Q_BUF U1 ( .A(n1), .Z(stat_datawords[1]));
Q_BUF U2 ( .A(n1), .Z(stat_datawords[2]));
Q_BUF U3 ( .A(n1), .Z(stat_datawords[3]));
Q_BUF U4 ( .A(n1), .Z(stat_datawords[4]));
Q_BUF U5 ( .A(n1), .Z(capability_type[0]));
Q_BUF U6 ( .A(n1), .Z(capability_type[1]));
Q_BUF U7 ( .A(n1), .Z(capability_type[2]));
Q_BUF U8 ( .A(n1), .Z(capability_type[3]));
Q_BUF U9 ( .A(n2), .Z(capability_lst[0]));
Q_BUF U10 ( .A(n2), .Z(capability_lst[1]));
Q_BUF U11 ( .A(n2), .Z(capability_lst[2]));
Q_BUF U12 ( .A(n2), .Z(capability_lst[3]));
Q_BUF U13 ( .A(n2), .Z(capability_lst[4]));
Q_BUF U14 ( .A(n2), .Z(capability_lst[5]));
Q_BUF U15 ( .A(n2), .Z(capability_lst[6]));
Q_BUF U16 ( .A(n1), .Z(capability_lst[7]));
Q_BUF U17 ( .A(n2), .Z(capability_lst[8]));
Q_BUF U18 ( .A(n1), .Z(capability_lst[9]));
Q_BUF U19 ( .A(n1), .Z(capability_lst[10]));
Q_BUF U20 ( .A(n1), .Z(capability_lst[11]));
Q_BUF U21 ( .A(n1), .Z(capability_lst[12]));
Q_BUF U22 ( .A(n1), .Z(capability_lst[13]));
Q_BUF U23 ( .A(n2), .Z(capability_lst[14]));
Q_BUF U24 ( .A(n2), .Z(capability_lst[15]));
Q_BUF U25 ( .A(n1), .Z(stat_table_id[0]));
ixc_assign_3 _zz_strnp_7 ( stat[2:0], stat_code[2:0]);
ixc_assign_4 _zz_strnp_1 ( cmnd[3:0], cmnd_op[3:0]);
ixc_assign \genblk1._zz_strnp_0 ( reset, rst_or_ini_r);
ixc_context_read_6 _zzixc_ctxrd_0 ( { stat_code[2], stat_code[1], 
	stat_code[0], stat[2], stat[1], stat[0]});
ixc_assign _zz_strnp_22 ( _zy_simnet_reset_14_w$, reset);
ixc_assign _zz_strnp_21 ( _zy_simnet_yield_13_w$, yield);
ixc_assign_64 _zz_strnp_20 ( _zy_simnet_sw_wdat_12_w$[0:63], sw_wdat[63:0]);
ixc_assign_15 _zz_strnp_19 ( _zy_simnet_sw_add_11_w$[0:14], sw_add[14:0]);
ixc_assign _zz_strnp_18 ( _zy_simnet_sw_we_10_w$, sw_we);
ixc_assign _zz_strnp_17 ( _zy_simnet_sw_ce_9_w$, sw_ce);
ixc_assign _zz_strnp_16 ( _zy_simnet_sw_cs_8_w$, sw_cs);
ixc_assign_64 _zz_strnp_15 ( _zy_simnet_rd_dat_7_w$[0:63], rd_dat[63:0]);
ixc_assign _zz_strnp_14 ( _zy_simnet_enable_6_w$, enable);
ixc_assign_4 _zz_strnp_13 ( _zy_simnet_capability_type_5_w$[0:3], { n1, n1, 
	n1, n1});
ixc_assign_16 _zz_strnp_12 ( _zy_simnet_capability_lst_4_w$[0:15], { n2, n2, 
	n1, n1, n1, n1, n1, n2, n1, n2, n2, n2, n2, n2, n2, n2});
ixc_assign _zz_strnp_11 ( _zy_simnet_stat_table_id_3_w$, n1);
ixc_assign_15 _zz_strnp_10 ( _zy_simnet_stat_addr_2_w$[0:14], stat_addr[14:0]);
ixc_assign_5 _zz_strnp_9 ( _zy_simnet_stat_datawords_1_w$[0:4], { n1, n1, n1, 
	n1, n2});
ixc_assign_3 _zz_strnp_8 ( _zy_simnet_stat_code_0_w$[0:2], stat_code[2:0]);
ixc_assign_15 _zz_strnp_6 ( stat_addr[14:0], maxaddr[14:0]);
Q_AN02 U46 ( .A0(n57), .A1(grant), .Z(igrant));
Q_OA21 U47 ( .A0(n56), .A1(n55), .B0(cmnd_issued), .Z(badaddr));
Q_AO21 U48 ( .A0(n17), .A1(n29), .B0(n16), .Z(n56));
Q_AO21 U49 ( .A0(n53), .A1(n42), .B0(n54), .Z(n55));
Q_AN03 U50 ( .A0(n53), .A1(n43), .A2(n52), .Z(n54));
Q_AN02 U51 ( .A0(n17), .A1(n30), .Z(n53));
Q_OR03 U52 ( .A0(n45), .A1(n51), .A2(n50), .Z(n52));
Q_AN03 U53 ( .A0(cmnd_addr[0]), .A1(n48), .A2(n49), .Z(n50));
Q_INV U54 ( .A(maxaddr[0]), .Z(n48));
Q_OA21 U55 ( .A0(cmnd_addr[1]), .A1(n47), .B0(n46), .Z(n49));
Q_AN03 U56 ( .A0(cmnd_addr[1]), .A1(n47), .A2(n46), .Z(n51));
Q_INV U57 ( .A(maxaddr[1]), .Z(n47));
Q_OR02 U58 ( .A0(cmnd_addr[2]), .A1(n44), .Z(n46));
Q_AN02 U59 ( .A0(cmnd_addr[2]), .A1(n44), .Z(n45));
Q_INV U60 ( .A(maxaddr[2]), .Z(n44));
Q_OR03 U61 ( .A0(n39), .A1(n38), .A2(n41), .Z(n42));
Q_OA21 U62 ( .A0(cmnd_addr[3]), .A1(n35), .B0(n37), .Z(n43));
Q_AN03 U63 ( .A0(cmnd_addr[3]), .A1(n35), .A2(n37), .Z(n38));
Q_INV U64 ( .A(maxaddr[3]), .Z(n35));
Q_OA21 U65 ( .A0(cmnd_addr[4]), .A1(n34), .B0(n36), .Z(n37));
Q_AN03 U66 ( .A0(cmnd_addr[4]), .A1(n34), .A2(n36), .Z(n39));
Q_INV U67 ( .A(maxaddr[4]), .Z(n34));
Q_OA21 U68 ( .A0(cmnd_addr[5]), .A1(n33), .B0(n32), .Z(n36));
Q_AN03 U69 ( .A0(cmnd_addr[5]), .A1(n33), .A2(n32), .Z(n40));
Q_INV U70 ( .A(maxaddr[5]), .Z(n33));
Q_OR02 U71 ( .A0(cmnd_addr[6]), .A1(n31), .Z(n32));
Q_AO21 U72 ( .A0(cmnd_addr[6]), .A1(n31), .B0(n40), .Z(n41));
Q_INV U73 ( .A(maxaddr[6]), .Z(n31));
Q_OR03 U74 ( .A0(n26), .A1(n25), .A2(n28), .Z(n29));
Q_OA21 U75 ( .A0(cmnd_addr[7]), .A1(n22), .B0(n24), .Z(n30));
Q_AN03 U76 ( .A0(cmnd_addr[7]), .A1(n22), .A2(n24), .Z(n25));
Q_INV U77 ( .A(maxaddr[7]), .Z(n22));
Q_OA21 U78 ( .A0(cmnd_addr[8]), .A1(n21), .B0(n23), .Z(n24));
Q_AN03 U79 ( .A0(cmnd_addr[8]), .A1(n21), .A2(n23), .Z(n26));
Q_INV U80 ( .A(maxaddr[8]), .Z(n21));
Q_OA21 U81 ( .A0(cmnd_addr[9]), .A1(n20), .B0(n19), .Z(n23));
Q_AN03 U82 ( .A0(cmnd_addr[9]), .A1(n20), .A2(n19), .Z(n27));
Q_INV U83 ( .A(maxaddr[9]), .Z(n20));
Q_OR02 U84 ( .A0(cmnd_addr[10]), .A1(n18), .Z(n19));
Q_AO21 U85 ( .A0(cmnd_addr[10]), .A1(n18), .B0(n27), .Z(n28));
Q_INV U86 ( .A(maxaddr[10]), .Z(n18));
Q_OR03 U87 ( .A0(n13), .A1(n12), .A2(n15), .Z(n16));
Q_OA21 U88 ( .A0(cmnd_addr[11]), .A1(n9), .B0(n11), .Z(n17));
Q_AN03 U89 ( .A0(cmnd_addr[11]), .A1(n9), .A2(n11), .Z(n12));
Q_INV U90 ( .A(maxaddr[11]), .Z(n9));
Q_OA21 U91 ( .A0(cmnd_addr[12]), .A1(n8), .B0(n10), .Z(n11));
Q_AN03 U92 ( .A0(cmnd_addr[12]), .A1(n8), .A2(n10), .Z(n13));
Q_INV U93 ( .A(maxaddr[12]), .Z(n8));
Q_OA21 U94 ( .A0(cmnd_addr[13]), .A1(n7), .B0(n6), .Z(n10));
Q_AN03 U95 ( .A0(cmnd_addr[13]), .A1(n7), .A2(n6), .Z(n14));
Q_INV U96 ( .A(maxaddr[13]), .Z(n7));
Q_OR02 U97 ( .A0(cmnd_addr[14]), .A1(n5), .Z(n6));
Q_AO21 U98 ( .A0(cmnd_addr[14]), .A1(n5), .B0(n14), .Z(n15));
Q_INV U99 ( .A(maxaddr[14]), .Z(n5));
Q_AN02 U100 ( .A0(n3), .A1(n4), .Z(timeout));
Q_AN03 U101 ( .A0(timer_r[2]), .A1(timer_r[1]), .A2(timer_r[0]), .Z(n4));
Q_AN03 U102 ( .A0(timer_r[5]), .A1(timer_r[4]), .A2(timer_r[3]), .Z(n3));
ixc_assign _zz_strnp_5 ( yield, timer_r[5]);
ixc_assign _zz_strnp_4 ( sw_we, sw_we_r);
ixc_assign _zz_strnp_3 ( sw_ce, sw_ce_r);
ixc_assign _zz_strnp_2 ( sw_cs, sw_cs_r);
Q_MX02 U107 ( .S(rst_or_ini_r), .A0(cmnd_addr[0]), .A1(rst_addr_r[0]), .Z(sw_add[0]));
Q_MX02 U108 ( .S(rst_or_ini_r), .A0(cmnd_addr[1]), .A1(rst_addr_r[1]), .Z(sw_add[1]));
Q_MX02 U109 ( .S(rst_or_ini_r), .A0(cmnd_addr[2]), .A1(rst_addr_r[2]), .Z(sw_add[2]));
Q_MX02 U110 ( .S(rst_or_ini_r), .A0(cmnd_addr[3]), .A1(rst_addr_r[3]), .Z(sw_add[3]));
Q_MX02 U111 ( .S(rst_or_ini_r), .A0(cmnd_addr[4]), .A1(rst_addr_r[4]), .Z(sw_add[4]));
Q_MX02 U112 ( .S(rst_or_ini_r), .A0(cmnd_addr[5]), .A1(rst_addr_r[5]), .Z(sw_add[5]));
Q_MX02 U113 ( .S(rst_or_ini_r), .A0(cmnd_addr[6]), .A1(rst_addr_r[6]), .Z(sw_add[6]));
Q_MX02 U114 ( .S(rst_or_ini_r), .A0(cmnd_addr[7]), .A1(rst_addr_r[7]), .Z(sw_add[7]));
Q_MX02 U115 ( .S(rst_or_ini_r), .A0(cmnd_addr[8]), .A1(rst_addr_r[8]), .Z(sw_add[8]));
Q_MX02 U116 ( .S(rst_or_ini_r), .A0(cmnd_addr[9]), .A1(rst_addr_r[9]), .Z(sw_add[9]));
Q_MX02 U117 ( .S(rst_or_ini_r), .A0(cmnd_addr[10]), .A1(rst_addr_r[10]), .Z(sw_add[10]));
Q_MX02 U118 ( .S(rst_or_ini_r), .A0(cmnd_addr[11]), .A1(rst_addr_r[11]), .Z(sw_add[11]));
Q_MX02 U119 ( .S(rst_or_ini_r), .A0(cmnd_addr[12]), .A1(rst_addr_r[12]), .Z(sw_add[12]));
Q_MX02 U120 ( .S(rst_or_ini_r), .A0(cmnd_addr[13]), .A1(rst_addr_r[13]), .Z(sw_add[13]));
Q_MX02 U121 ( .S(rst_or_ini_r), .A0(cmnd_addr[14]), .A1(rst_addr_r[14]), .Z(sw_add[14]));
Q_AN02 U122 ( .A0(enable), .A1(\addr_limit[0][0] ), .Z(maxaddr[0]));
Q_AN02 U123 ( .A0(enable), .A1(\addr_limit[0][1] ), .Z(maxaddr[1]));
Q_AN02 U124 ( .A0(enable), .A1(\addr_limit[0][2] ), .Z(maxaddr[2]));
Q_AN02 U125 ( .A0(enable), .A1(\addr_limit[0][3] ), .Z(maxaddr[3]));
Q_AN02 U126 ( .A0(enable), .A1(\addr_limit[0][4] ), .Z(maxaddr[4]));
Q_AN02 U127 ( .A0(enable), .A1(\addr_limit[0][5] ), .Z(maxaddr[5]));
Q_AN02 U128 ( .A0(enable), .A1(\addr_limit[0][6] ), .Z(maxaddr[6]));
Q_AN02 U129 ( .A0(enable), .A1(\addr_limit[0][7] ), .Z(maxaddr[7]));
Q_AN02 U130 ( .A0(enable), .A1(\addr_limit[0][8] ), .Z(maxaddr[8]));
Q_AN02 U131 ( .A0(enable), .A1(\addr_limit[0][9] ), .Z(maxaddr[9]));
Q_AN02 U132 ( .A0(enable), .A1(\addr_limit[0][10] ), .Z(maxaddr[10]));
Q_AN02 U133 ( .A0(enable), .A1(\addr_limit[0][11] ), .Z(maxaddr[11]));
Q_AN02 U134 ( .A0(enable), .A1(\addr_limit[0][12] ), .Z(maxaddr[12]));
Q_AN02 U135 ( .A0(enable), .A1(\addr_limit[0][13] ), .Z(maxaddr[13]));
Q_AN02 U136 ( .A0(enable), .A1(\addr_limit[0][14] ), .Z(maxaddr[14]));
Q_INV U137 ( .A(reg_addr[7]), .Z(n58));
Q_INV U138 ( .A(reg_addr[8]), .Z(n59));
Q_OR03 U139 ( .A0(reg_addr[10]), .A1(reg_addr[9]), .A2(n59), .Z(n60));
Q_OR03 U140 ( .A0(n58), .A1(reg_addr[6]), .A2(reg_addr[5]), .Z(n61));
Q_ND03 U141 ( .A0(reg_addr[4]), .A1(reg_addr[3]), .A2(reg_addr[2]), .Z(n62));
Q_OR03 U142 ( .A0(reg_addr[1]), .A1(reg_addr[0]), .A2(n60), .Z(n63));
Q_NR03 U143 ( .A0(n61), .A1(n62), .A2(n63), .Z(n64));
Q_AN02 U144 ( .A0(wr_stb), .A1(n64), .Z(n87));
Q_INV U145 ( .A(n83), .Z(cmnd_issued));
Q_INV U146 ( .A(unsupported_op), .Z(n82));
Q_OA21 U147 ( .A0(n66), .A1(n67), .B0(n65), .Z(unsupported_op));
Q_AN02 U148 ( .A0(n65), .A1(n68), .Z(ack_error));
Q_AO21 U149 ( .A0(n70), .A1(n71), .B0(n69), .Z(n83));
Q_INV U150 ( .A(n87), .Z(n69));
Q_MX02 U151 ( .S(cmnd[3]), .A0(n74), .A1(n72), .Z(n70));
Q_INV U152 ( .A(cmnd_cmp_stb), .Z(n84));
Q_AN02 U153 ( .A0(n65), .A1(n75), .Z(cmnd_cmp_stb));
Q_AN02 U154 ( .A0(n65), .A1(n76), .Z(cmnd_tmo_stb));
Q_AN03 U155 ( .A0(n65), .A1(n71), .A2(n74), .Z(cmnd_sis_stb));
Q_AN02 U156 ( .A0(n87), .A1(cmnd[3]), .Z(n65));
Q_AN02 U157 ( .A0(n77), .A1(n68), .Z(cmnd_inc_stb));
Q_AN02 U158 ( .A0(n72), .A1(cmnd[0]), .Z(n68));
Q_AN02 U159 ( .A0(n77), .A1(n76), .Z(cmnd_ini_stb));
Q_AN02 U160 ( .A0(n72), .A1(n71), .Z(n76));
Q_AN02 U161 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n72));
Q_INV U162 ( .A(cmnd_rst_stb), .Z(n85));
Q_AN02 U163 ( .A0(n67), .A1(n78), .Z(cmnd_rst_stb));
Q_AN02 U164 ( .A0(n77), .A1(cmnd[0]), .Z(n78));
Q_AN02 U165 ( .A0(n67), .A1(n79), .Z(cmnd_dis_stb));
Q_AN02 U166 ( .A0(n77), .A1(n71), .Z(n79));
Q_AN02 U167 ( .A0(cmnd[2]), .A1(n80), .Z(n67));
Q_AN02 U168 ( .A0(n66), .A1(n78), .Z(cmnd_ena_stb));
Q_INV U169 ( .A(cmnd_wr_stb), .Z(n86));
Q_AN02 U170 ( .A0(n66), .A1(n79), .Z(cmnd_wr_stb));
Q_INV U171 ( .A(cmnd[0]), .Z(n71));
Q_AN02 U172 ( .A0(n81), .A1(cmnd[1]), .Z(n66));
Q_AN02 U173 ( .A0(n77), .A1(n75), .Z(cmnd_rd_stb));
Q_AN02 U174 ( .A0(n74), .A1(cmnd[0]), .Z(n75));
Q_NR02 U175 ( .A0(cmnd[2]), .A1(cmnd[1]), .Z(n74));
Q_INV U176 ( .A(cmnd[1]), .Z(n80));
Q_INV U177 ( .A(cmnd[2]), .Z(n81));
Q_AN02 U178 ( .A0(n87), .A1(n73), .Z(n77));
Q_INV U179 ( .A(cmnd[3]), .Z(n73));
Q_OR02 U180 ( .A0(cmnd_ini_stb), .A1(cmnd_inc_stb), .Z(n493));
Q_XNR2 U181 ( .A0(rst_addr_r[0]), .A1(maxaddr[0]), .Z(n88));
Q_XNR2 U182 ( .A0(rst_addr_r[1]), .A1(maxaddr[1]), .Z(n89));
Q_XNR2 U183 ( .A0(rst_addr_r[2]), .A1(maxaddr[2]), .Z(n90));
Q_XNR2 U184 ( .A0(rst_addr_r[3]), .A1(maxaddr[3]), .Z(n91));
Q_XNR2 U185 ( .A0(rst_addr_r[4]), .A1(maxaddr[4]), .Z(n92));
Q_XNR2 U186 ( .A0(rst_addr_r[5]), .A1(maxaddr[5]), .Z(n93));
Q_XNR2 U187 ( .A0(rst_addr_r[6]), .A1(maxaddr[6]), .Z(n94));
Q_XNR2 U188 ( .A0(rst_addr_r[7]), .A1(maxaddr[7]), .Z(n95));
Q_XNR2 U189 ( .A0(rst_addr_r[8]), .A1(maxaddr[8]), .Z(n96));
Q_XNR2 U190 ( .A0(rst_addr_r[9]), .A1(maxaddr[9]), .Z(n97));
Q_XNR2 U191 ( .A0(rst_addr_r[10]), .A1(maxaddr[10]), .Z(n98));
Q_XNR2 U192 ( .A0(rst_addr_r[11]), .A1(maxaddr[11]), .Z(n99));
Q_XNR2 U193 ( .A0(rst_addr_r[12]), .A1(maxaddr[12]), .Z(n100));
Q_XNR2 U194 ( .A0(rst_addr_r[13]), .A1(maxaddr[13]), .Z(n101));
Q_XNR2 U195 ( .A0(rst_addr_r[14]), .A1(maxaddr[14]), .Z(n102));
Q_AN03 U196 ( .A0(n102), .A1(n101), .A2(n100), .Z(n103));
Q_AN03 U197 ( .A0(n99), .A1(n98), .A2(n97), .Z(n104));
Q_AN03 U198 ( .A0(n96), .A1(n95), .A2(n94), .Z(n105));
Q_AN03 U199 ( .A0(n93), .A1(n92), .A2(n91), .Z(n106));
Q_AN03 U200 ( .A0(n90), .A1(n89), .A2(n88), .Z(n107));
Q_AN03 U201 ( .A0(n103), .A1(n104), .A2(n105), .Z(n108));
Q_AN03 U202 ( .A0(n106), .A1(n107), .A2(n108), .Z(n494));
Q_XNR2 U203 ( .A0(rst_addr_r[0]), .A1(cmnd_addr[0]), .Z(n109));
Q_XNR2 U204 ( .A0(rst_addr_r[1]), .A1(cmnd_addr[1]), .Z(n110));
Q_XNR2 U205 ( .A0(rst_addr_r[2]), .A1(cmnd_addr[2]), .Z(n111));
Q_XNR2 U206 ( .A0(rst_addr_r[3]), .A1(cmnd_addr[3]), .Z(n112));
Q_XNR2 U207 ( .A0(rst_addr_r[4]), .A1(cmnd_addr[4]), .Z(n113));
Q_XNR2 U208 ( .A0(rst_addr_r[5]), .A1(cmnd_addr[5]), .Z(n114));
Q_XNR2 U209 ( .A0(rst_addr_r[6]), .A1(cmnd_addr[6]), .Z(n115));
Q_XNR2 U210 ( .A0(rst_addr_r[7]), .A1(cmnd_addr[7]), .Z(n116));
Q_XNR2 U211 ( .A0(rst_addr_r[8]), .A1(cmnd_addr[8]), .Z(n117));
Q_XNR2 U212 ( .A0(rst_addr_r[9]), .A1(cmnd_addr[9]), .Z(n118));
Q_XNR2 U213 ( .A0(rst_addr_r[10]), .A1(cmnd_addr[10]), .Z(n119));
Q_XNR2 U214 ( .A0(rst_addr_r[11]), .A1(cmnd_addr[11]), .Z(n120));
Q_XNR2 U215 ( .A0(rst_addr_r[12]), .A1(cmnd_addr[12]), .Z(n121));
Q_XNR2 U216 ( .A0(rst_addr_r[13]), .A1(cmnd_addr[13]), .Z(n122));
Q_XNR2 U217 ( .A0(rst_addr_r[14]), .A1(cmnd_addr[14]), .Z(n123));
Q_AN03 U218 ( .A0(n123), .A1(n122), .A2(n121), .Z(n124));
Q_AN03 U219 ( .A0(n120), .A1(n119), .A2(n118), .Z(n125));
Q_AN03 U220 ( .A0(n117), .A1(n116), .A2(n115), .Z(n126));
Q_AN03 U221 ( .A0(n114), .A1(n113), .A2(n112), .Z(n127));
Q_AN03 U222 ( .A0(n111), .A1(n110), .A2(n109), .Z(n128));
Q_AN03 U223 ( .A0(n124), .A1(n125), .A2(n126), .Z(n129));
Q_AN03 U224 ( .A0(n127), .A1(n128), .A2(n129), .Z(n495));
Q_AN02 U225 ( .A0(init_inc_r), .A1(igrant), .Z(n130));
Q_XOR2 U226 ( .A0(inc_r[0]), .A1(n130), .Z(n131));
Q_AD01HF U227 ( .A0(rst_addr_r[0]), .B0(igrant), .S(n132), .CO(n133));
Q_AD01HF U228 ( .A0(rst_addr_r[1]), .B0(n133), .S(n134), .CO(n135));
Q_AD01HF U229 ( .A0(rst_addr_r[2]), .B0(n135), .S(n136), .CO(n137));
Q_AD01HF U230 ( .A0(rst_addr_r[3]), .B0(n137), .S(n138), .CO(n139));
Q_AD01HF U231 ( .A0(rst_addr_r[4]), .B0(n139), .S(n140), .CO(n141));
Q_AD01HF U232 ( .A0(rst_addr_r[5]), .B0(n141), .S(n142), .CO(n143));
Q_AD01HF U233 ( .A0(rst_addr_r[6]), .B0(n143), .S(n144), .CO(n145));
Q_AD01HF U234 ( .A0(rst_addr_r[7]), .B0(n145), .S(n146), .CO(n147));
Q_AD01HF U235 ( .A0(rst_addr_r[8]), .B0(n147), .S(n148), .CO(n149));
Q_AD01HF U236 ( .A0(rst_addr_r[9]), .B0(n149), .S(n150), .CO(n151));
Q_AD01HF U237 ( .A0(rst_addr_r[10]), .B0(n151), .S(n152), .CO(n153));
Q_AD01HF U238 ( .A0(rst_addr_r[11]), .B0(n153), .S(n154), .CO(n155));
Q_AD01HF U239 ( .A0(rst_addr_r[12]), .B0(n155), .S(n156), .CO(n157));
Q_AD01HF U240 ( .A0(rst_addr_r[13]), .B0(n157), .S(n158), .CO(n159));
Q_XOR2 U241 ( .A0(rst_addr_r[14]), .A1(n159), .Z(n160));
Q_AD01HF U242 ( .A0(timer_r[1]), .B0(timer_r[0]), .S(n162), .CO(n163));
Q_AD01HF U243 ( .A0(timer_r[2]), .B0(n163), .S(n164), .CO(n165));
Q_AD01HF U244 ( .A0(timer_r[3]), .B0(n165), .S(n166), .CO(n167));
Q_AD01HF U245 ( .A0(timer_r[4]), .B0(n167), .S(n168), .CO(n169));
Q_XOR2 U246 ( .A0(timer_r[5]), .A1(n169), .Z(n170));
Q_INV U247 ( .A(n171), .Z(n172));
Q_MX02 U248 ( .S(n416), .A0(n175), .A1(n173), .Z(n171));
Q_XOR2 U249 ( .A0(n471), .A1(n174), .Z(n173));
Q_AN02 U250 ( .A0(n470), .A1(n472), .Z(n174));
Q_OR02 U251 ( .A0(n471), .A1(n176), .Z(n175));
Q_INV U252 ( .A(n177), .Z(n178));
Q_MX02 U253 ( .S(n471), .A0(n179), .A1(n180), .Z(n177));
Q_ND02 U254 ( .A0(n349), .A1(n472), .Z(n180));
Q_AN02 U255 ( .A0(n416), .A1(n182), .Z(n181));
Q_MX02 U256 ( .S(n471), .A0(n183), .A1(n176), .Z(n182));
Q_NR02 U257 ( .A0(n349), .A1(n472), .Z(n183));
Q_OR02 U258 ( .A0(n470), .A1(n472), .Z(n176));
Q_NR03 U259 ( .A0(n473), .A1(n471), .A2(n185), .Z(n184));
Q_INV U260 ( .A(n179), .Z(n185));
Q_XOR2 U261 ( .A0(n349), .A1(n472), .Z(n179));
Q_AN02 U262 ( .A0(n473), .A1(n471), .Z(n186));
Q_AO21 U263 ( .A0(n186), .A1(state_r[3]), .B0(n184), .Z(n499));
Q_AO21 U264 ( .A0(n186), .A1(state_r[2]), .B0(n181), .Z(n498));
Q_AO21 U265 ( .A0(n186), .A1(state_r[1]), .B0(n178), .Z(n497));
Q_AO21 U266 ( .A0(n186), .A1(state_r[0]), .B0(n172), .Z(n496));
Q_AN02 U267 ( .A0(n474), .A1(n161), .Z(n187));
Q_AN02 U268 ( .A0(n474), .A1(n162), .Z(n188));
Q_AN02 U269 ( .A0(n474), .A1(n164), .Z(n189));
Q_AN02 U270 ( .A0(n474), .A1(n166), .Z(n190));
Q_AN02 U271 ( .A0(n474), .A1(n168), .Z(n191));
Q_AN02 U272 ( .A0(n474), .A1(n170), .Z(n192));
Q_AN02 U273 ( .A0(n476), .A1(cmnd_addr[0]), .Z(n193));
Q_MX02 U274 ( .S(n477), .A0(n193), .A1(n132), .Z(n194));
Q_AN02 U275 ( .A0(n476), .A1(cmnd_addr[1]), .Z(n195));
Q_MX02 U276 ( .S(n477), .A0(n195), .A1(n134), .Z(n196));
Q_AN02 U277 ( .A0(n476), .A1(cmnd_addr[2]), .Z(n197));
Q_MX02 U278 ( .S(n477), .A0(n197), .A1(n136), .Z(n198));
Q_AN02 U279 ( .A0(n476), .A1(cmnd_addr[3]), .Z(n199));
Q_MX02 U280 ( .S(n477), .A0(n199), .A1(n138), .Z(n200));
Q_AN02 U281 ( .A0(n476), .A1(cmnd_addr[4]), .Z(n201));
Q_MX02 U282 ( .S(n477), .A0(n201), .A1(n140), .Z(n202));
Q_AN02 U283 ( .A0(n476), .A1(cmnd_addr[5]), .Z(n203));
Q_MX02 U284 ( .S(n477), .A0(n203), .A1(n142), .Z(n204));
Q_AN02 U285 ( .A0(n476), .A1(cmnd_addr[6]), .Z(n205));
Q_MX02 U286 ( .S(n477), .A0(n205), .A1(n144), .Z(n206));
Q_AN02 U287 ( .A0(n476), .A1(cmnd_addr[7]), .Z(n207));
Q_MX02 U288 ( .S(n477), .A0(n207), .A1(n146), .Z(n208));
Q_AN02 U289 ( .A0(n476), .A1(cmnd_addr[8]), .Z(n209));
Q_MX02 U290 ( .S(n477), .A0(n209), .A1(n148), .Z(n210));
Q_AN02 U291 ( .A0(n476), .A1(cmnd_addr[9]), .Z(n211));
Q_MX02 U292 ( .S(n477), .A0(n211), .A1(n150), .Z(n212));
Q_AN02 U293 ( .A0(n476), .A1(cmnd_addr[10]), .Z(n213));
Q_MX02 U294 ( .S(n477), .A0(n213), .A1(n152), .Z(n214));
Q_AN02 U295 ( .A0(n476), .A1(cmnd_addr[11]), .Z(n215));
Q_MX02 U296 ( .S(n477), .A0(n215), .A1(n154), .Z(n216));
Q_AN02 U297 ( .A0(n476), .A1(cmnd_addr[12]), .Z(n217));
Q_MX02 U298 ( .S(n477), .A0(n217), .A1(n156), .Z(n218));
Q_AN02 U299 ( .A0(n476), .A1(cmnd_addr[13]), .Z(n219));
Q_MX02 U300 ( .S(n477), .A0(n219), .A1(n158), .Z(n220));
Q_AN02 U301 ( .A0(n476), .A1(cmnd_addr[14]), .Z(n221));
Q_MX02 U302 ( .S(n477), .A0(n221), .A1(n160), .Z(n222));
Q_AN02 U303 ( .A0(n482), .A1(n131), .Z(n223));
Q_MX03 U304 ( .S0(n484), .S1(n485), .A0(sw_aindex[0]), .A1(wr_dat[0]), .A2(sw_rdat[0]), .Z(n224));
Q_MX03 U305 ( .S0(n484), .S1(n485), .A0(sw_aindex[1]), .A1(wr_dat[1]), .A2(sw_rdat[1]), .Z(n225));
Q_MX03 U306 ( .S0(n484), .S1(n485), .A0(sw_aindex[2]), .A1(wr_dat[2]), .A2(sw_rdat[2]), .Z(n226));
Q_MX03 U307 ( .S0(n484), .S1(n485), .A0(sw_aindex[3]), .A1(wr_dat[3]), .A2(sw_rdat[3]), .Z(n227));
Q_MX03 U308 ( .S0(n484), .S1(n485), .A0(sw_aindex[4]), .A1(wr_dat[4]), .A2(sw_rdat[4]), .Z(n228));
Q_MX03 U309 ( .S0(n484), .S1(n485), .A0(sw_aindex[5]), .A1(wr_dat[5]), .A2(sw_rdat[5]), .Z(n229));
Q_MX03 U310 ( .S0(n484), .S1(n485), .A0(sw_aindex[6]), .A1(wr_dat[6]), .A2(sw_rdat[6]), .Z(n230));
Q_MX03 U311 ( .S0(n484), .S1(n485), .A0(sw_aindex[7]), .A1(wr_dat[7]), .A2(sw_rdat[7]), .Z(n231));
Q_MX03 U312 ( .S0(n484), .S1(n485), .A0(sw_aindex[8]), .A1(wr_dat[8]), .A2(sw_rdat[8]), .Z(n232));
Q_MX03 U313 ( .S0(n484), .S1(n485), .A0(sw_aindex[9]), .A1(wr_dat[9]), .A2(sw_rdat[9]), .Z(n233));
Q_MX03 U314 ( .S0(n484), .S1(n485), .A0(sw_aindex[10]), .A1(wr_dat[10]), .A2(sw_rdat[10]), .Z(n234));
Q_MX03 U315 ( .S0(n484), .S1(n485), .A0(sw_aindex[11]), .A1(wr_dat[11]), .A2(sw_rdat[11]), .Z(n235));
Q_MX03 U316 ( .S0(n484), .S1(n485), .A0(sw_aindex[12]), .A1(wr_dat[12]), .A2(sw_rdat[12]), .Z(n236));
Q_MX03 U317 ( .S0(n484), .S1(n485), .A0(sw_aindex[13]), .A1(wr_dat[13]), .A2(sw_rdat[13]), .Z(n237));
Q_MX03 U318 ( .S0(n484), .S1(n485), .A0(sw_match), .A1(wr_dat[14]), .A2(sw_rdat[14]), .Z(n238));
Q_AN02 U319 ( .A0(n484), .A1(wr_dat[15]), .Z(n239));
Q_MX02 U320 ( .S(n485), .A0(n239), .A1(sw_rdat[15]), .Z(n240));
Q_AN02 U321 ( .A0(n484), .A1(wr_dat[16]), .Z(n241));
Q_MX02 U322 ( .S(n485), .A0(n241), .A1(sw_rdat[16]), .Z(n242));
Q_AN02 U323 ( .A0(n484), .A1(wr_dat[17]), .Z(n243));
Q_MX02 U324 ( .S(n485), .A0(n243), .A1(sw_rdat[17]), .Z(n244));
Q_AN02 U325 ( .A0(n484), .A1(wr_dat[18]), .Z(n245));
Q_MX02 U326 ( .S(n485), .A0(n245), .A1(sw_rdat[18]), .Z(n246));
Q_AN02 U327 ( .A0(n484), .A1(wr_dat[19]), .Z(n247));
Q_MX02 U328 ( .S(n485), .A0(n247), .A1(sw_rdat[19]), .Z(n248));
Q_AN02 U329 ( .A0(n484), .A1(wr_dat[20]), .Z(n249));
Q_MX02 U330 ( .S(n485), .A0(n249), .A1(sw_rdat[20]), .Z(n250));
Q_AN02 U331 ( .A0(n484), .A1(wr_dat[21]), .Z(n251));
Q_MX02 U332 ( .S(n485), .A0(n251), .A1(sw_rdat[21]), .Z(n252));
Q_AN02 U333 ( .A0(n484), .A1(wr_dat[22]), .Z(n253));
Q_MX02 U334 ( .S(n485), .A0(n253), .A1(sw_rdat[22]), .Z(n254));
Q_AN02 U335 ( .A0(n484), .A1(wr_dat[23]), .Z(n255));
Q_MX02 U336 ( .S(n485), .A0(n255), .A1(sw_rdat[23]), .Z(n256));
Q_AN02 U337 ( .A0(n484), .A1(wr_dat[24]), .Z(n257));
Q_MX02 U338 ( .S(n485), .A0(n257), .A1(sw_rdat[24]), .Z(n258));
Q_AN02 U339 ( .A0(n484), .A1(wr_dat[25]), .Z(n259));
Q_MX02 U340 ( .S(n485), .A0(n259), .A1(sw_rdat[25]), .Z(n260));
Q_AN02 U341 ( .A0(n484), .A1(wr_dat[26]), .Z(n261));
Q_MX02 U342 ( .S(n485), .A0(n261), .A1(sw_rdat[26]), .Z(n262));
Q_AN02 U343 ( .A0(n484), .A1(wr_dat[27]), .Z(n263));
Q_MX02 U344 ( .S(n485), .A0(n263), .A1(sw_rdat[27]), .Z(n264));
Q_AN02 U345 ( .A0(n484), .A1(wr_dat[28]), .Z(n265));
Q_MX02 U346 ( .S(n485), .A0(n265), .A1(sw_rdat[28]), .Z(n266));
Q_AN02 U347 ( .A0(n484), .A1(wr_dat[29]), .Z(n267));
Q_MX02 U348 ( .S(n485), .A0(n267), .A1(sw_rdat[29]), .Z(n268));
Q_AN02 U349 ( .A0(n484), .A1(wr_dat[30]), .Z(n269));
Q_MX02 U350 ( .S(n485), .A0(n269), .A1(sw_rdat[30]), .Z(n270));
Q_AN02 U351 ( .A0(n484), .A1(wr_dat[31]), .Z(n271));
Q_MX02 U352 ( .S(n485), .A0(n271), .A1(sw_rdat[31]), .Z(n272));
Q_AN02 U353 ( .A0(n484), .A1(wr_dat[32]), .Z(n273));
Q_MX02 U354 ( .S(n485), .A0(n273), .A1(sw_rdat[32]), .Z(n274));
Q_AN02 U355 ( .A0(n484), .A1(wr_dat[33]), .Z(n275));
Q_MX02 U356 ( .S(n485), .A0(n275), .A1(sw_rdat[33]), .Z(n276));
Q_AN02 U357 ( .A0(n484), .A1(wr_dat[34]), .Z(n277));
Q_MX02 U358 ( .S(n485), .A0(n277), .A1(sw_rdat[34]), .Z(n278));
Q_AN02 U359 ( .A0(n484), .A1(wr_dat[35]), .Z(n279));
Q_MX02 U360 ( .S(n485), .A0(n279), .A1(sw_rdat[35]), .Z(n280));
Q_AN02 U361 ( .A0(n484), .A1(wr_dat[36]), .Z(n281));
Q_MX02 U362 ( .S(n485), .A0(n281), .A1(sw_rdat[36]), .Z(n282));
Q_AN02 U363 ( .A0(n484), .A1(wr_dat[37]), .Z(n283));
Q_MX02 U364 ( .S(n485), .A0(n283), .A1(sw_rdat[37]), .Z(n284));
Q_AN02 U365 ( .A0(n484), .A1(wr_dat[38]), .Z(n285));
Q_MX02 U366 ( .S(n485), .A0(n285), .A1(sw_rdat[38]), .Z(n286));
Q_AN02 U367 ( .A0(n484), .A1(wr_dat[39]), .Z(n287));
Q_MX02 U368 ( .S(n485), .A0(n287), .A1(sw_rdat[39]), .Z(n288));
Q_AN02 U369 ( .A0(n484), .A1(wr_dat[40]), .Z(n289));
Q_MX02 U370 ( .S(n485), .A0(n289), .A1(sw_rdat[40]), .Z(n290));
Q_AN02 U371 ( .A0(n484), .A1(wr_dat[41]), .Z(n291));
Q_MX02 U372 ( .S(n485), .A0(n291), .A1(sw_rdat[41]), .Z(n292));
Q_AN02 U373 ( .A0(n484), .A1(wr_dat[42]), .Z(n293));
Q_MX02 U374 ( .S(n485), .A0(n293), .A1(sw_rdat[42]), .Z(n294));
Q_AN02 U375 ( .A0(n484), .A1(wr_dat[43]), .Z(n295));
Q_MX02 U376 ( .S(n485), .A0(n295), .A1(sw_rdat[43]), .Z(n296));
Q_AN02 U377 ( .A0(n484), .A1(wr_dat[44]), .Z(n297));
Q_MX02 U378 ( .S(n485), .A0(n297), .A1(sw_rdat[44]), .Z(n298));
Q_AN02 U379 ( .A0(n484), .A1(wr_dat[45]), .Z(n299));
Q_MX02 U380 ( .S(n485), .A0(n299), .A1(sw_rdat[45]), .Z(n300));
Q_AN02 U381 ( .A0(n484), .A1(wr_dat[46]), .Z(n301));
Q_MX02 U382 ( .S(n485), .A0(n301), .A1(sw_rdat[46]), .Z(n302));
Q_AN02 U383 ( .A0(n484), .A1(wr_dat[47]), .Z(n303));
Q_MX02 U384 ( .S(n485), .A0(n303), .A1(sw_rdat[47]), .Z(n304));
Q_AN02 U385 ( .A0(n484), .A1(wr_dat[48]), .Z(n305));
Q_MX02 U386 ( .S(n485), .A0(n305), .A1(sw_rdat[48]), .Z(n306));
Q_AN02 U387 ( .A0(n484), .A1(wr_dat[49]), .Z(n307));
Q_MX02 U388 ( .S(n485), .A0(n307), .A1(sw_rdat[49]), .Z(n308));
Q_AN02 U389 ( .A0(n484), .A1(wr_dat[50]), .Z(n309));
Q_MX02 U390 ( .S(n485), .A0(n309), .A1(sw_rdat[50]), .Z(n310));
Q_AN02 U391 ( .A0(n484), .A1(wr_dat[51]), .Z(n311));
Q_MX02 U392 ( .S(n485), .A0(n311), .A1(sw_rdat[51]), .Z(n312));
Q_AN02 U393 ( .A0(n484), .A1(wr_dat[52]), .Z(n313));
Q_MX02 U394 ( .S(n485), .A0(n313), .A1(sw_rdat[52]), .Z(n314));
Q_AN02 U395 ( .A0(n484), .A1(wr_dat[53]), .Z(n315));
Q_MX02 U396 ( .S(n485), .A0(n315), .A1(sw_rdat[53]), .Z(n316));
Q_AN02 U397 ( .A0(n484), .A1(wr_dat[54]), .Z(n317));
Q_MX02 U398 ( .S(n485), .A0(n317), .A1(sw_rdat[54]), .Z(n318));
Q_AN02 U399 ( .A0(n484), .A1(wr_dat[55]), .Z(n319));
Q_MX02 U400 ( .S(n485), .A0(n319), .A1(sw_rdat[55]), .Z(n320));
Q_AN02 U401 ( .A0(n484), .A1(wr_dat[56]), .Z(n321));
Q_MX02 U402 ( .S(n485), .A0(n321), .A1(sw_rdat[56]), .Z(n322));
Q_AN02 U403 ( .A0(n484), .A1(wr_dat[57]), .Z(n323));
Q_MX02 U404 ( .S(n485), .A0(n323), .A1(sw_rdat[57]), .Z(n324));
Q_AN02 U405 ( .A0(n484), .A1(wr_dat[58]), .Z(n325));
Q_MX02 U406 ( .S(n485), .A0(n325), .A1(sw_rdat[58]), .Z(n326));
Q_AN02 U407 ( .A0(n484), .A1(wr_dat[59]), .Z(n327));
Q_MX02 U408 ( .S(n485), .A0(n327), .A1(sw_rdat[59]), .Z(n328));
Q_AN02 U409 ( .A0(n484), .A1(wr_dat[60]), .Z(n329));
Q_MX02 U410 ( .S(n485), .A0(n329), .A1(sw_rdat[60]), .Z(n330));
Q_AN02 U411 ( .A0(n484), .A1(wr_dat[61]), .Z(n331));
Q_MX02 U412 ( .S(n485), .A0(n331), .A1(sw_rdat[61]), .Z(n332));
Q_AN02 U413 ( .A0(n484), .A1(wr_dat[62]), .Z(n333));
Q_MX02 U414 ( .S(n485), .A0(n333), .A1(sw_rdat[62]), .Z(n334));
Q_AN02 U415 ( .A0(n484), .A1(wr_dat[63]), .Z(n335));
Q_MX02 U416 ( .S(n485), .A0(n335), .A1(sw_rdat[63]), .Z(n336));
Q_FDP1 \state_r_REG[3] ( .CK(clk), .R(rst_n), .D(n499), .Q(state_r[3]), .QN(n364));
Q_FDP1 \state_r_REG[2] ( .CK(clk), .R(rst_n), .D(n498), .Q(state_r[2]), .QN(n365));
Q_FDP1 \state_r_REG[1] ( .CK(clk), .R(rst_n), .D(n497), .Q(state_r[1]), .QN(n367));
Q_FDP1 \state_r_REG[0] ( .CK(clk), .R(rst_n), .D(n496), .Q(state_r[0]), .QN(n363));
Q_FDP1 \timer_r_REG[5] ( .CK(clk), .R(rst_n), .D(n192), .Q(timer_r[5]), .QN( ));
Q_FDP1 \timer_r_REG[4] ( .CK(clk), .R(rst_n), .D(n191), .Q(timer_r[4]), .QN( ));
Q_FDP1 \timer_r_REG[3] ( .CK(clk), .R(rst_n), .D(n190), .Q(timer_r[3]), .QN( ));
Q_FDP1 \timer_r_REG[2] ( .CK(clk), .R(rst_n), .D(n189), .Q(timer_r[2]), .QN( ));
Q_FDP1 \timer_r_REG[1] ( .CK(clk), .R(rst_n), .D(n188), .Q(timer_r[1]), .QN( ));
Q_FDP1 \timer_r_REG[0] ( .CK(clk), .R(rst_n), .D(n187), .Q(timer_r[0]), .QN(n161));
Q_ND02 U427 ( .A0(n338), .A1(n339), .Z(n337));
Q_ND02 U428 ( .A0(n340), .A1(n442), .Z(n339));
Q_OR02 U429 ( .A0(n341), .A1(n487), .Z(n340));
Q_INV U430 ( .A(n486), .Z(n341));
Q_ND02 U431 ( .A0(n338), .A1(n343), .Z(n342));
Q_ND02 U432 ( .A0(n486), .A1(n442), .Z(n343));
Q_OR03 U433 ( .A0(n486), .A1(n487), .A2(n442), .Z(n338));
Q_MX02 U434 ( .S(n442), .A0(n486), .A1(n487), .Z(n344));
Q_FDP2 \stat_code_REG[2] ( .CK(clk), .S(rst_n), .D(n345), .Q(stat_code[2]), .QN( ));
Q_MX02 U436 ( .S(n457), .A0(stat_code[2]), .A1(n344), .Z(n345));
Q_FDP2 \stat_code_REG[1] ( .CK(clk), .S(rst_n), .D(n346), .Q(stat_code[1]), .QN( ));
Q_MX02 U438 ( .S(n457), .A0(stat_code[1]), .A1(n342), .Z(n346));
Q_FDP2 \stat_code_REG[0] ( .CK(clk), .S(rst_n), .D(n347), .Q(stat_code[0]), .QN( ));
Q_MX02 U440 ( .S(n457), .A0(stat_code[0]), .A1(n337), .Z(n347));
Q_FDP2 init_r_REG  ( .CK(clk), .S(rst_n), .D(n348), .Q(init_r), .QN(enable));
Q_MX02 U442 ( .S(n489), .A0(init_r), .A1(n483), .Z(n348));
Q_FDP1 sw_cs_r_REG  ( .CK(clk), .R(rst_n), .D(n481), .Q(sw_cs_r), .QN( ));
Q_FDP1 sw_ce_r_REG  ( .CK(clk), .R(rst_n), .D(n480), .Q(sw_ce_r), .QN( ));
Q_FDP1 rst_r_REG  ( .CK(clk), .R(rst_n), .D(n479), .Q(rst_r), .QN(n500));
Q_FDP1 rst_or_ini_r_REG  ( .CK(clk), .R(rst_n), .D(n478), .Q(rst_or_ini_r), .QN( ));
Q_FDP1 sw_we_r_REG  ( .CK(clk), .R(rst_n), .D(n475), .Q(sw_we_r), .QN( ));
Q_INV U448 ( .A(n349), .Z(n470));
Q_OA21 U449 ( .A0(n351), .A1(n352), .B0(n350), .Z(n349));
Q_AN03 U450 ( .A0(state_r[0]), .A1(n356), .A2(n354), .Z(n355));
Q_OR03 U451 ( .A0(n358), .A1(n359), .A2(n353), .Z(n352));
Q_AO21 U452 ( .A0(n360), .A1(n361), .B0(n355), .Z(n357));
Q_AN02 U453 ( .A0(n362), .A1(n363), .Z(n361));
Q_NR02 U454 ( .A0(state_r[3]), .A1(state_r[2]), .Z(n362));
Q_MX02 U455 ( .S(state_r[1]), .A0(cmnd_ena_stb), .A1(n366), .Z(n360));
Q_AN02 U456 ( .A0(n369), .A1(n83), .Z(n368));
Q_AO21 U457 ( .A0(n370), .A1(n371), .B0(n357), .Z(n358));
Q_NR02 U458 ( .A0(cmnd_dis_stb), .A1(unsupported_op), .Z(n371));
Q_OA21 U459 ( .A0(n372), .A1(n373), .B0(n368), .Z(n359));
Q_AN03 U460 ( .A0(n375), .A1(state_r[3]), .A2(n366), .Z(n374));
Q_AN02 U461 ( .A0(ack_error), .A1(enable), .Z(n366));
Q_OR02 U462 ( .A0(n376), .A1(n374), .Z(n373));
Q_AN02 U463 ( .A0(n364), .A1(igrant), .Z(n377));
Q_OA21 U464 ( .A0(n378), .A1(n379), .B0(n377), .Z(n372));
Q_AN02 U465 ( .A0(n381), .A1(n494), .Z(n378));
Q_OA21 U466 ( .A0(state_r[0]), .A1(n495), .B0(n380), .Z(n379));
Q_AN02 U467 ( .A0(n385), .A1(n84), .Z(n383));
Q_AN03 U468 ( .A0(cmnd_rst_stb), .A1(n354), .A2(n383), .Z(n384));
Q_OR03 U469 ( .A0(n386), .A1(n384), .A2(n382), .Z(n351));
Q_AN02 U470 ( .A0(n387), .A1(n388), .Z(n386));
Q_NR02 U471 ( .A0(timeout), .A1(state_r[0]), .Z(n389));
Q_OA21 U472 ( .A0(n390), .A1(n353), .B0(n350), .Z(n471));
Q_OR02 U473 ( .A0(n391), .A1(n392), .Z(n390));
Q_AO21 U474 ( .A0(n395), .A1(n396), .B0(n393), .Z(n353));
Q_AN02 U475 ( .A0(n397), .A1(n83), .Z(n396));
Q_NR02 U476 ( .A0(timeout), .A1(state_r[3]), .Z(n397));
Q_OA21 U477 ( .A0(n398), .A1(n399), .B0(n394), .Z(n393));
Q_AN02 U478 ( .A0(n364), .A1(n400), .Z(n399));
Q_NR02 U479 ( .A0(state_r[0]), .A1(cmnd_ena_stb), .Z(n400));
Q_AN02 U480 ( .A0(n401), .A1(n402), .Z(n398));
Q_MX02 U481 ( .S(state_r[0]), .A0(n404), .A1(n403), .Z(n401));
Q_AO21 U482 ( .A0(n406), .A1(n381), .B0(n405), .Z(n395));
Q_OA21 U483 ( .A0(n407), .A1(n408), .B0(state_r[2]), .Z(n405));
Q_NR02 U484 ( .A0(n409), .A1(rsp), .Z(n408));
Q_INV U485 ( .A(rsp), .Z(n403));
Q_AO21 U486 ( .A0(n409), .A1(n404), .B0(n410), .Z(n407));
Q_NR02 U487 ( .A0(n411), .A1(n495), .Z(n410));
Q_ND02 U488 ( .A0(igrant), .A1(n494), .Z(n406));
Q_OA21 U489 ( .A0(n412), .A1(n413), .B0(n491), .Z(n472));
Q_AN02 U490 ( .A0(n414), .A1(n415), .Z(n412));
Q_INV U491 ( .A(n416), .Z(n473));
Q_OA21 U492 ( .A0(n417), .A1(n391), .B0(n350), .Z(n416));
Q_AN03 U493 ( .A0(n413), .A1(state_r[0]), .A2(n354), .Z(n392));
Q_INV U494 ( .A(n415), .Z(n413));
Q_AN02 U495 ( .A0(n86), .A1(cmnd_rd_stb), .Z(n356));
Q_AN03 U496 ( .A0(n354), .A1(n385), .A2(n414), .Z(n418));
Q_AO21 U497 ( .A0(cmnd_rst_stb), .A1(n84), .B0(cmnd_cmp_stb), .Z(n414));
Q_OR03 U498 ( .A0(n419), .A1(n418), .A2(n392), .Z(n417));
Q_AN02 U499 ( .A0(n420), .A1(n387), .Z(n419));
Q_AN03 U500 ( .A0(igrant), .A1(n83), .A2(n389), .Z(n387));
Q_AO21 U501 ( .A0(n421), .A1(n422), .B0(n382), .Z(n391));
Q_AN03 U502 ( .A0(n84), .A1(n493), .A2(n385), .Z(n422));
Q_AN02 U503 ( .A0(ack_error), .A1(init_r), .Z(n424));
Q_AO21 U504 ( .A0(n370), .A1(cmnd_dis_stb), .B0(n423), .Z(n382));
Q_AN03 U505 ( .A0(n385), .A1(n425), .A2(n421), .Z(n370));
Q_NR02 U506 ( .A0(cmnd_cmp_stb), .A1(n493), .Z(n425));
Q_AN02 U507 ( .A0(state_r[0]), .A1(n415), .Z(n385));
Q_NR02 U508 ( .A0(cmnd_wr_stb), .A1(cmnd_rd_stb), .Z(n415));
Q_AN02 U509 ( .A0(n85), .A1(n354), .Z(n421));
Q_OA21 U510 ( .A0(n426), .A1(n427), .B0(n424), .Z(n423));
Q_AN02 U511 ( .A0(n375), .A1(n402), .Z(n426));
Q_AN03 U512 ( .A0(n369), .A1(state_r[3]), .A2(n83), .Z(n402));
Q_INV U513 ( .A(n394), .Z(n375));
Q_AN02 U514 ( .A0(n404), .A1(n481), .Z(n474));
Q_INV U515 ( .A(igrant), .Z(n404));
Q_OA21 U516 ( .A0(n429), .A1(n430), .B0(n428), .Z(n475));
Q_AN02 U517 ( .A0(cmnd_sis_stb), .A1(n431), .Z(n476));
Q_INV U518 ( .A(n477), .Z(n431));
Q_OR02 U519 ( .A0(state_r[0]), .A1(state_r[1]), .Z(n411));
Q_ND02 U520 ( .A0(state_r[1]), .A1(state_r[0]), .Z(n409));
Q_OA21 U521 ( .A0(n429), .A1(n432), .B0(n428), .Z(n478));
Q_AN02 U522 ( .A0(n430), .A1(n433), .Z(n432));
Q_AN02 U523 ( .A0(n498), .A1(n434), .Z(n430));
Q_AN02 U524 ( .A0(n428), .A1(n429), .Z(n479));
Q_AN02 U525 ( .A0(n435), .A1(n496), .Z(n429));
Q_OR03 U526 ( .A0(n479), .A1(n436), .A2(n480), .Z(n481));
Q_AN02 U527 ( .A0(n499), .A1(n437), .Z(n480));
Q_AN03 U528 ( .A0(n428), .A1(n498), .A2(n438), .Z(n436));
Q_INV U529 ( .A(n439), .Z(n438));
Q_INV U530 ( .A(n440), .Z(n482));
Q_AN02 U531 ( .A0(n441), .A1(state_r[0]), .Z(n485));
Q_AN02 U532 ( .A0(n444), .A1(n445), .Z(n446));
Q_INV U533 ( .A(n447), .Z(n444));
Q_OR03 U534 ( .A0(n448), .A1(n446), .A2(n443), .Z(n442));
Q_AN03 U535 ( .A0(n450), .A1(n82), .A2(n449), .Z(n443));
Q_OR02 U536 ( .A0(n439), .A1(n451), .Z(n448));
Q_AN02 U537 ( .A0(n497), .A1(n496), .Z(n439));
Q_INV U538 ( .A(n452), .Z(n451));
Q_AN02 U539 ( .A0(n428), .A1(n453), .Z(n445));
Q_NR02 U540 ( .A0(n498), .A1(n496), .Z(n453));
Q_OA21 U541 ( .A0(n455), .A1(n434), .B0(n445), .Z(n486));
Q_AN02 U542 ( .A0(n82), .A1(n497), .Z(n447));
Q_OA21 U543 ( .A0(n450), .A1(badaddr), .B0(n447), .Z(n455));
Q_AN02 U544 ( .A0(timeout), .A1(n350), .Z(n450));
Q_NR02 U545 ( .A0(n499), .A1(n498), .Z(n452));
Q_OA21 U546 ( .A0(n456), .A1(n434), .B0(n452), .Z(n487));
Q_AN03 U547 ( .A0(n497), .A1(n433), .A2(unsupported_op), .Z(n456));
Q_ND02 U548 ( .A0(n427), .A1(n449), .Z(n457));
Q_AN02 U549 ( .A0(n435), .A1(n458), .Z(n449));
Q_NR02 U550 ( .A0(n499), .A1(n496), .Z(n458));
Q_AN02 U551 ( .A0(n454), .A1(n497), .Z(n435));
Q_AN02 U552 ( .A0(n459), .A1(n460), .Z(n427));
Q_NR02 U553 ( .A0(state_r[3]), .A1(state_r[0]), .Z(n459));
Q_OA21 U554 ( .A0(n484), .A1(n376), .B0(n350), .Z(n488));
Q_AN03 U555 ( .A0(state_r[0]), .A1(rsp), .A2(n420), .Z(n376));
Q_INV U556 ( .A(n483), .Z(n484));
Q_AN02 U557 ( .A0(n364), .A1(n394), .Z(n354));
Q_OR02 U558 ( .A0(n441), .A1(n388), .Z(n420));
Q_AN02 U559 ( .A0(state_r[3]), .A1(n394), .Z(n388));
Q_AN03 U560 ( .A0(state_r[2]), .A1(state_r[1]), .A2(n364), .Z(n441));
Q_AN03 U561 ( .A0(n483), .A1(n428), .A2(n437), .Z(n461));
Q_AN02 U562 ( .A0(n462), .A1(n433), .Z(n437));
Q_INV U563 ( .A(n496), .Z(n433));
Q_NR02 U564 ( .A0(n498), .A1(n497), .Z(n462));
Q_INV U565 ( .A(n497), .Z(n434));
Q_INV U566 ( .A(n498), .Z(n454));
Q_INV U567 ( .A(n499), .Z(n428));
Q_AO21 U568 ( .A0(n463), .A1(n464), .B0(n461), .Z(n489));
Q_AN02 U569 ( .A0(n363), .A1(cmnd_ena_stb), .Z(n464));
Q_OR02 U570 ( .A0(state_r[3]), .A1(state_r[1]), .Z(n465));
Q_OR03 U571 ( .A0(state_r[2]), .A1(state_r[0]), .A2(n465), .Z(n483));
Q_AN03 U572 ( .A0(n467), .A1(n367), .A2(n466), .Z(n490));
Q_AO21 U573 ( .A0(state_r[2]), .A1(n363), .B0(n440), .Z(n466));
Q_AN02 U574 ( .A0(n365), .A1(state_r[0]), .Z(n440));
Q_AN02 U575 ( .A0(n463), .A1(state_r[0]), .Z(n491));
Q_AN02 U576 ( .A0(n467), .A1(n394), .Z(n463));
Q_NR02 U577 ( .A0(state_r[2]), .A1(state_r[1]), .Z(n394));
Q_NR02 U578 ( .A0(badaddr), .A1(state_r[3]), .Z(n467));
Q_INV U579 ( .A(badaddr), .Z(n350));
Q_OR03 U580 ( .A0(cmnd_rst_stb), .A1(cmnd_sis_stb), .A2(n477), .Z(n492));
Q_OA21 U581 ( .A0(n381), .A1(n468), .B0(n467), .Z(n477));
Q_AN02 U582 ( .A0(n380), .A1(n363), .Z(n468));
Q_AN02 U583 ( .A0(state_r[2]), .A1(n367), .Z(n380));
Q_AN02 U584 ( .A0(n460), .A1(state_r[0]), .Z(n381));
Q_AN02 U585 ( .A0(n365), .A1(state_r[1]), .Z(n460));
Q_OR02 U586 ( .A0(cmnd_tmo_stb), .A1(timeout), .Z(n469));
Q_INV U587 ( .A(timeout), .Z(n369));
Q_AN02 U588 ( .A0(n500), .A1(wr_dat[0]), .Z(sw_wdat[0]));
Q_AN02 U589 ( .A0(n500), .A1(wr_dat[1]), .Z(sw_wdat[1]));
Q_AN02 U590 ( .A0(n500), .A1(wr_dat[2]), .Z(sw_wdat[2]));
Q_AN02 U591 ( .A0(n500), .A1(wr_dat[3]), .Z(sw_wdat[3]));
Q_AN02 U592 ( .A0(n500), .A1(wr_dat[4]), .Z(sw_wdat[4]));
Q_AN02 U593 ( .A0(n500), .A1(wr_dat[5]), .Z(sw_wdat[5]));
Q_AN02 U594 ( .A0(n500), .A1(wr_dat[6]), .Z(sw_wdat[6]));
Q_AN02 U595 ( .A0(n500), .A1(wr_dat[7]), .Z(sw_wdat[7]));
Q_AN02 U596 ( .A0(n500), .A1(wr_dat[8]), .Z(sw_wdat[8]));
Q_AN02 U597 ( .A0(n500), .A1(wr_dat[9]), .Z(sw_wdat[9]));
Q_AN02 U598 ( .A0(n500), .A1(wr_dat[10]), .Z(sw_wdat[10]));
Q_AN02 U599 ( .A0(n500), .A1(wr_dat[11]), .Z(sw_wdat[11]));
Q_AN02 U600 ( .A0(n500), .A1(wr_dat[12]), .Z(sw_wdat[12]));
Q_AN02 U601 ( .A0(n500), .A1(wr_dat[13]), .Z(sw_wdat[13]));
Q_AN02 U602 ( .A0(n500), .A1(wr_dat[14]), .Z(sw_wdat[14]));
Q_AN02 U603 ( .A0(n500), .A1(wr_dat[15]), .Z(sw_wdat[15]));
Q_AN02 U604 ( .A0(n500), .A1(wr_dat[16]), .Z(sw_wdat[16]));
Q_AN02 U605 ( .A0(n500), .A1(wr_dat[17]), .Z(sw_wdat[17]));
Q_AN02 U606 ( .A0(n500), .A1(wr_dat[18]), .Z(sw_wdat[18]));
Q_AN02 U607 ( .A0(n500), .A1(wr_dat[19]), .Z(sw_wdat[19]));
Q_AN02 U608 ( .A0(n500), .A1(wr_dat[20]), .Z(sw_wdat[20]));
Q_AN02 U609 ( .A0(n500), .A1(wr_dat[21]), .Z(sw_wdat[21]));
Q_AN02 U610 ( .A0(n500), .A1(wr_dat[22]), .Z(sw_wdat[22]));
Q_AN02 U611 ( .A0(n500), .A1(wr_dat[23]), .Z(sw_wdat[23]));
Q_AN02 U612 ( .A0(n500), .A1(wr_dat[24]), .Z(sw_wdat[24]));
Q_AN02 U613 ( .A0(n500), .A1(wr_dat[25]), .Z(sw_wdat[25]));
Q_AN02 U614 ( .A0(n500), .A1(wr_dat[26]), .Z(sw_wdat[26]));
Q_AN02 U615 ( .A0(n500), .A1(wr_dat[27]), .Z(sw_wdat[27]));
Q_AN02 U616 ( .A0(n500), .A1(wr_dat[28]), .Z(sw_wdat[28]));
Q_AN02 U617 ( .A0(n500), .A1(wr_dat[29]), .Z(sw_wdat[29]));
Q_AN02 U618 ( .A0(n500), .A1(wr_dat[30]), .Z(sw_wdat[30]));
Q_AN02 U619 ( .A0(n500), .A1(wr_dat[31]), .Z(sw_wdat[31]));
Q_AN02 U620 ( .A0(n500), .A1(wr_dat[32]), .Z(sw_wdat[32]));
Q_AN02 U621 ( .A0(n500), .A1(wr_dat[33]), .Z(sw_wdat[33]));
Q_AN02 U622 ( .A0(n500), .A1(wr_dat[34]), .Z(sw_wdat[34]));
Q_AN02 U623 ( .A0(n500), .A1(wr_dat[35]), .Z(sw_wdat[35]));
Q_AN02 U624 ( .A0(n500), .A1(wr_dat[36]), .Z(sw_wdat[36]));
Q_AN02 U625 ( .A0(n500), .A1(wr_dat[37]), .Z(sw_wdat[37]));
Q_AN02 U626 ( .A0(n500), .A1(wr_dat[38]), .Z(sw_wdat[38]));
Q_AN02 U627 ( .A0(n500), .A1(wr_dat[39]), .Z(sw_wdat[39]));
Q_AN02 U628 ( .A0(n500), .A1(wr_dat[40]), .Z(sw_wdat[40]));
Q_AN02 U629 ( .A0(n500), .A1(wr_dat[41]), .Z(sw_wdat[41]));
Q_AN02 U630 ( .A0(n500), .A1(wr_dat[42]), .Z(sw_wdat[42]));
Q_AN02 U631 ( .A0(n500), .A1(wr_dat[43]), .Z(sw_wdat[43]));
Q_AN02 U632 ( .A0(n500), .A1(wr_dat[44]), .Z(sw_wdat[44]));
Q_AN02 U633 ( .A0(n500), .A1(wr_dat[45]), .Z(sw_wdat[45]));
Q_AN02 U634 ( .A0(n500), .A1(wr_dat[46]), .Z(sw_wdat[46]));
Q_AN02 U635 ( .A0(n500), .A1(wr_dat[47]), .Z(sw_wdat[47]));
Q_AN02 U636 ( .A0(n500), .A1(wr_dat[48]), .Z(sw_wdat[48]));
Q_AN02 U637 ( .A0(n500), .A1(wr_dat[49]), .Z(sw_wdat[49]));
Q_AN02 U638 ( .A0(n500), .A1(wr_dat[50]), .Z(sw_wdat[50]));
Q_AN02 U639 ( .A0(n500), .A1(wr_dat[51]), .Z(sw_wdat[51]));
Q_AN02 U640 ( .A0(n500), .A1(wr_dat[52]), .Z(sw_wdat[52]));
Q_AN02 U641 ( .A0(n500), .A1(wr_dat[53]), .Z(sw_wdat[53]));
Q_AN02 U642 ( .A0(n500), .A1(wr_dat[54]), .Z(sw_wdat[54]));
Q_AN02 U643 ( .A0(n500), .A1(wr_dat[55]), .Z(sw_wdat[55]));
Q_AN02 U644 ( .A0(n500), .A1(wr_dat[56]), .Z(sw_wdat[56]));
Q_AN02 U645 ( .A0(n500), .A1(wr_dat[57]), .Z(sw_wdat[57]));
Q_AN02 U646 ( .A0(n500), .A1(wr_dat[58]), .Z(sw_wdat[58]));
Q_AN02 U647 ( .A0(n500), .A1(wr_dat[59]), .Z(sw_wdat[59]));
Q_AN02 U648 ( .A0(n500), .A1(wr_dat[60]), .Z(sw_wdat[60]));
Q_AN02 U649 ( .A0(n500), .A1(wr_dat[61]), .Z(sw_wdat[61]));
Q_AN02 U650 ( .A0(n500), .A1(wr_dat[62]), .Z(sw_wdat[62]));
Q_AN02 U651 ( .A0(n500), .A1(wr_dat[63]), .Z(sw_wdat[63]));
Q_FDP4EP sim_tmo_r_REG  ( .CK(clk), .CE(n469), .R(n501), .D(cmnd_tmo_stb), .Q(sim_tmo_r));
Q_INV U653 ( .A(rst_n), .Z(n501));
Q_INV U654 ( .A(sim_tmo_r), .Z(n57));
Q_FDP4EP \rst_addr_r_REG[0] ( .CK(clk), .CE(n492), .R(n501), .D(n194), .Q(rst_addr_r[0]));
Q_FDP4EP \rst_addr_r_REG[1] ( .CK(clk), .CE(n492), .R(n501), .D(n196), .Q(rst_addr_r[1]));
Q_FDP4EP \rst_addr_r_REG[2] ( .CK(clk), .CE(n492), .R(n501), .D(n198), .Q(rst_addr_r[2]));
Q_FDP4EP \rst_addr_r_REG[3] ( .CK(clk), .CE(n492), .R(n501), .D(n200), .Q(rst_addr_r[3]));
Q_FDP4EP \rst_addr_r_REG[4] ( .CK(clk), .CE(n492), .R(n501), .D(n202), .Q(rst_addr_r[4]));
Q_FDP4EP \rst_addr_r_REG[5] ( .CK(clk), .CE(n492), .R(n501), .D(n204), .Q(rst_addr_r[5]));
Q_FDP4EP \rst_addr_r_REG[6] ( .CK(clk), .CE(n492), .R(n501), .D(n206), .Q(rst_addr_r[6]));
Q_FDP4EP \rst_addr_r_REG[7] ( .CK(clk), .CE(n492), .R(n501), .D(n208), .Q(rst_addr_r[7]));
Q_FDP4EP \rst_addr_r_REG[8] ( .CK(clk), .CE(n492), .R(n501), .D(n210), .Q(rst_addr_r[8]));
Q_FDP4EP \rst_addr_r_REG[9] ( .CK(clk), .CE(n492), .R(n501), .D(n212), .Q(rst_addr_r[9]));
Q_FDP4EP \rst_addr_r_REG[10] ( .CK(clk), .CE(n492), .R(n501), .D(n214), .Q(rst_addr_r[10]));
Q_FDP4EP \rst_addr_r_REG[11] ( .CK(clk), .CE(n492), .R(n501), .D(n216), .Q(rst_addr_r[11]));
Q_FDP4EP \rst_addr_r_REG[12] ( .CK(clk), .CE(n492), .R(n501), .D(n218), .Q(rst_addr_r[12]));
Q_FDP4EP \rst_addr_r_REG[13] ( .CK(clk), .CE(n492), .R(n501), .D(n220), .Q(rst_addr_r[13]));
Q_FDP4EP \rst_addr_r_REG[14] ( .CK(clk), .CE(n492), .R(n501), .D(n222), .Q(rst_addr_r[14]));
Q_FDP4EP \inc_r_REG[0] ( .CK(clk), .CE(n490), .R(n501), .D(n223), .Q(inc_r[0]));
Q_FDP4EP \rd_dat_REG[0] ( .CK(clk), .CE(n488), .R(n501), .D(n224), .Q(rd_dat[0]));
Q_FDP4EP \rd_dat_REG[1] ( .CK(clk), .CE(n488), .R(n501), .D(n225), .Q(rd_dat[1]));
Q_FDP4EP \rd_dat_REG[2] ( .CK(clk), .CE(n488), .R(n501), .D(n226), .Q(rd_dat[2]));
Q_FDP4EP \rd_dat_REG[3] ( .CK(clk), .CE(n488), .R(n501), .D(n227), .Q(rd_dat[3]));
Q_FDP4EP \rd_dat_REG[4] ( .CK(clk), .CE(n488), .R(n501), .D(n228), .Q(rd_dat[4]));
Q_FDP4EP \rd_dat_REG[5] ( .CK(clk), .CE(n488), .R(n501), .D(n229), .Q(rd_dat[5]));
Q_FDP4EP \rd_dat_REG[6] ( .CK(clk), .CE(n488), .R(n501), .D(n230), .Q(rd_dat[6]));
Q_FDP4EP \rd_dat_REG[7] ( .CK(clk), .CE(n488), .R(n501), .D(n231), .Q(rd_dat[7]));
Q_FDP4EP \rd_dat_REG[8] ( .CK(clk), .CE(n488), .R(n501), .D(n232), .Q(rd_dat[8]));
Q_FDP4EP \rd_dat_REG[9] ( .CK(clk), .CE(n488), .R(n501), .D(n233), .Q(rd_dat[9]));
Q_FDP4EP \rd_dat_REG[10] ( .CK(clk), .CE(n488), .R(n501), .D(n234), .Q(rd_dat[10]));
Q_FDP4EP \rd_dat_REG[11] ( .CK(clk), .CE(n488), .R(n501), .D(n235), .Q(rd_dat[11]));
Q_FDP4EP \rd_dat_REG[12] ( .CK(clk), .CE(n488), .R(n501), .D(n236), .Q(rd_dat[12]));
Q_FDP4EP \rd_dat_REG[13] ( .CK(clk), .CE(n488), .R(n501), .D(n237), .Q(rd_dat[13]));
Q_FDP4EP \rd_dat_REG[14] ( .CK(clk), .CE(n488), .R(n501), .D(n238), .Q(rd_dat[14]));
Q_FDP4EP \rd_dat_REG[15] ( .CK(clk), .CE(n488), .R(n501), .D(n240), .Q(rd_dat[15]));
Q_FDP4EP \rd_dat_REG[16] ( .CK(clk), .CE(n488), .R(n501), .D(n242), .Q(rd_dat[16]));
Q_FDP4EP \rd_dat_REG[17] ( .CK(clk), .CE(n488), .R(n501), .D(n244), .Q(rd_dat[17]));
Q_FDP4EP \rd_dat_REG[18] ( .CK(clk), .CE(n488), .R(n501), .D(n246), .Q(rd_dat[18]));
Q_FDP4EP \rd_dat_REG[19] ( .CK(clk), .CE(n488), .R(n501), .D(n248), .Q(rd_dat[19]));
Q_FDP4EP \rd_dat_REG[20] ( .CK(clk), .CE(n488), .R(n501), .D(n250), .Q(rd_dat[20]));
Q_FDP4EP \rd_dat_REG[21] ( .CK(clk), .CE(n488), .R(n501), .D(n252), .Q(rd_dat[21]));
Q_FDP4EP \rd_dat_REG[22] ( .CK(clk), .CE(n488), .R(n501), .D(n254), .Q(rd_dat[22]));
Q_FDP4EP \rd_dat_REG[23] ( .CK(clk), .CE(n488), .R(n501), .D(n256), .Q(rd_dat[23]));
Q_FDP4EP \rd_dat_REG[24] ( .CK(clk), .CE(n488), .R(n501), .D(n258), .Q(rd_dat[24]));
Q_FDP4EP \rd_dat_REG[25] ( .CK(clk), .CE(n488), .R(n501), .D(n260), .Q(rd_dat[25]));
Q_FDP4EP \rd_dat_REG[26] ( .CK(clk), .CE(n488), .R(n501), .D(n262), .Q(rd_dat[26]));
Q_FDP4EP \rd_dat_REG[27] ( .CK(clk), .CE(n488), .R(n501), .D(n264), .Q(rd_dat[27]));
Q_FDP4EP \rd_dat_REG[28] ( .CK(clk), .CE(n488), .R(n501), .D(n266), .Q(rd_dat[28]));
Q_FDP4EP \rd_dat_REG[29] ( .CK(clk), .CE(n488), .R(n501), .D(n268), .Q(rd_dat[29]));
Q_FDP4EP \rd_dat_REG[30] ( .CK(clk), .CE(n488), .R(n501), .D(n270), .Q(rd_dat[30]));
Q_FDP4EP \rd_dat_REG[31] ( .CK(clk), .CE(n488), .R(n501), .D(n272), .Q(rd_dat[31]));
Q_FDP4EP \rd_dat_REG[32] ( .CK(clk), .CE(n488), .R(n501), .D(n274), .Q(rd_dat[32]));
Q_FDP4EP \rd_dat_REG[33] ( .CK(clk), .CE(n488), .R(n501), .D(n276), .Q(rd_dat[33]));
Q_FDP4EP \rd_dat_REG[34] ( .CK(clk), .CE(n488), .R(n501), .D(n278), .Q(rd_dat[34]));
Q_FDP4EP \rd_dat_REG[35] ( .CK(clk), .CE(n488), .R(n501), .D(n280), .Q(rd_dat[35]));
Q_FDP4EP \rd_dat_REG[36] ( .CK(clk), .CE(n488), .R(n501), .D(n282), .Q(rd_dat[36]));
Q_FDP4EP \rd_dat_REG[37] ( .CK(clk), .CE(n488), .R(n501), .D(n284), .Q(rd_dat[37]));
Q_FDP4EP \rd_dat_REG[38] ( .CK(clk), .CE(n488), .R(n501), .D(n286), .Q(rd_dat[38]));
Q_FDP4EP \rd_dat_REG[39] ( .CK(clk), .CE(n488), .R(n501), .D(n288), .Q(rd_dat[39]));
Q_FDP4EP \rd_dat_REG[40] ( .CK(clk), .CE(n488), .R(n501), .D(n290), .Q(rd_dat[40]));
Q_FDP4EP \rd_dat_REG[41] ( .CK(clk), .CE(n488), .R(n501), .D(n292), .Q(rd_dat[41]));
Q_FDP4EP \rd_dat_REG[42] ( .CK(clk), .CE(n488), .R(n501), .D(n294), .Q(rd_dat[42]));
Q_FDP4EP \rd_dat_REG[43] ( .CK(clk), .CE(n488), .R(n501), .D(n296), .Q(rd_dat[43]));
Q_FDP4EP \rd_dat_REG[44] ( .CK(clk), .CE(n488), .R(n501), .D(n298), .Q(rd_dat[44]));
Q_FDP4EP \rd_dat_REG[45] ( .CK(clk), .CE(n488), .R(n501), .D(n300), .Q(rd_dat[45]));
Q_FDP4EP \rd_dat_REG[46] ( .CK(clk), .CE(n488), .R(n501), .D(n302), .Q(rd_dat[46]));
Q_FDP4EP \rd_dat_REG[47] ( .CK(clk), .CE(n488), .R(n501), .D(n304), .Q(rd_dat[47]));
Q_FDP4EP \rd_dat_REG[48] ( .CK(clk), .CE(n488), .R(n501), .D(n306), .Q(rd_dat[48]));
Q_FDP4EP \rd_dat_REG[49] ( .CK(clk), .CE(n488), .R(n501), .D(n308), .Q(rd_dat[49]));
Q_FDP4EP \rd_dat_REG[50] ( .CK(clk), .CE(n488), .R(n501), .D(n310), .Q(rd_dat[50]));
Q_FDP4EP \rd_dat_REG[51] ( .CK(clk), .CE(n488), .R(n501), .D(n312), .Q(rd_dat[51]));
Q_FDP4EP \rd_dat_REG[52] ( .CK(clk), .CE(n488), .R(n501), .D(n314), .Q(rd_dat[52]));
Q_FDP4EP \rd_dat_REG[53] ( .CK(clk), .CE(n488), .R(n501), .D(n316), .Q(rd_dat[53]));
Q_FDP4EP \rd_dat_REG[54] ( .CK(clk), .CE(n488), .R(n501), .D(n318), .Q(rd_dat[54]));
Q_FDP4EP \rd_dat_REG[55] ( .CK(clk), .CE(n488), .R(n501), .D(n320), .Q(rd_dat[55]));
Q_FDP4EP \rd_dat_REG[56] ( .CK(clk), .CE(n488), .R(n501), .D(n322), .Q(rd_dat[56]));
Q_FDP4EP \rd_dat_REG[57] ( .CK(clk), .CE(n488), .R(n501), .D(n324), .Q(rd_dat[57]));
Q_FDP4EP \rd_dat_REG[58] ( .CK(clk), .CE(n488), .R(n501), .D(n326), .Q(rd_dat[58]));
Q_FDP4EP \rd_dat_REG[59] ( .CK(clk), .CE(n488), .R(n501), .D(n328), .Q(rd_dat[59]));
Q_FDP4EP \rd_dat_REG[60] ( .CK(clk), .CE(n488), .R(n501), .D(n330), .Q(rd_dat[60]));
Q_FDP4EP \rd_dat_REG[61] ( .CK(clk), .CE(n488), .R(n501), .D(n332), .Q(rd_dat[61]));
Q_FDP4EP \rd_dat_REG[62] ( .CK(clk), .CE(n488), .R(n501), .D(n334), .Q(rd_dat[62]));
Q_FDP4EP \rd_dat_REG[63] ( .CK(clk), .CE(n488), .R(n501), .D(n336), .Q(rd_dat[63]));
Q_FDP4EP init_inc_r_REG  ( .CK(clk), .CE(n491), .R(n501), .D(n1), .Q(init_inc_r));
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_m1 "addr_limit (2,0) 1 14 0 0 0"
// pragma CVASTRPROP MODULE HDLICE HDL_UCDB_MDARRAY_DECL_NUM "1"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "-1 genblk2  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 genblk1  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk2"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "genblk1"
endmodule
