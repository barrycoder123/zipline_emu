
`ifndef _2_                      
`ifdef CBV                      
`define _2_                      
`else                      
`define _2_ (* _2_state_ *)                      
`endif                      
`endif
(* celldefine = 1 *) 
module nx_ram_1rw_xcm108 ( clk, rst_n, ovstb, lvm, mlvm, mrdten, bimc_rst_n, 
	bimc_isync, bimc_idat, bimc_odat, bimc_osync, 
	ro_uncorrectable_ecc_error, bwe, din, add, cs, we, dout);
// pragma CVASTRPROP MODULE HDLICE HDL_MODULE_ATTRIBUTE "0 vlog"
input clk;
input rst_n;
input ovstb;
input lvm;
input mlvm;
input mrdten;
input bimc_rst_n;
input bimc_isync;
input bimc_idat;
output bimc_odat;
output bimc_osync;
output ro_uncorrectable_ecc_error;
input [37:0] bwe;
input [37:0] din;
input [13:0] add;
input cs;
input we;
output [37:0] dout;
wire _zy_simnet_bimc_odat_0_w$;
wire _zy_simnet_bimc_osync_1_w$;
wire _zy_simnet_ro_uncorrectable_ecc_error_2_w$;
wire bimc_iclk;
wire bimc_irstn;
wire rst_clk_n;
wire p_mode_disable_ecc_mem;
wire byp;
wire se;
wire rds;
wire [1:0] ecc_corrupt;
wire rst_rclk_n;
wire sew;
wire web;
wire ro_mem_ecc_error_ev;
wire ro_mem_ecc_corrected;
wire [13:0] ro_mem_ecc_error_addr;
wire [37:0] \g.dout_i ;
wire [37:0] \g.dat_r ;
wire [37:0] \g.din_i ;
wire [16383:0] \g.we_clk ;
wire [31:0] \g.u_ram._zyictd_sysfunc_11_L263_10 ;
wire [16383:0] \g.we_gate ;
wire [13:0] \g.add_r ;
supply0 n138;
Q_BUF U0 ( .A(n138), .Z(p_mode_disable_ecc_mem));
Q_BUF U1 ( .A(n138), .Z(byp));
Q_BUF U2 ( .A(n138), .Z(se));
Q_BUF U3 ( .A(n138), .Z(rds));
Q_BUF U4 ( .A(n138), .Z(ecc_corrupt[1]));
Q_BUF U5 ( .A(n138), .Z(ecc_corrupt[0]));
Q_BUF U6 ( .A(n138), .Z(sew));
Q_ASSIGN U7 ( .B(clk), .A(\g.we_clk [16383]));
Q_ASSIGN U8 ( .B(clk), .A(\g.we_clk [16382]));
Q_ASSIGN U9 ( .B(clk), .A(\g.we_clk [16381]));
Q_ASSIGN U10 ( .B(clk), .A(\g.we_clk [16380]));
Q_ASSIGN U11 ( .B(clk), .A(\g.we_clk [16379]));
Q_ASSIGN U12 ( .B(clk), .A(\g.we_clk [16378]));
Q_ASSIGN U13 ( .B(clk), .A(\g.we_clk [16377]));
Q_ASSIGN U14 ( .B(clk), .A(\g.we_clk [16376]));
Q_ASSIGN U15 ( .B(clk), .A(\g.we_clk [16375]));
Q_ASSIGN U16 ( .B(clk), .A(\g.we_clk [16374]));
Q_ASSIGN U17 ( .B(clk), .A(\g.we_clk [16373]));
Q_ASSIGN U18 ( .B(clk), .A(\g.we_clk [16372]));
Q_ASSIGN U19 ( .B(clk), .A(\g.we_clk [16371]));
Q_ASSIGN U20 ( .B(clk), .A(\g.we_clk [16370]));
Q_ASSIGN U21 ( .B(clk), .A(\g.we_clk [16369]));
Q_ASSIGN U22 ( .B(clk), .A(\g.we_clk [16368]));
Q_ASSIGN U23 ( .B(clk), .A(\g.we_clk [16367]));
Q_ASSIGN U24 ( .B(clk), .A(\g.we_clk [16366]));
Q_ASSIGN U25 ( .B(clk), .A(\g.we_clk [16365]));
Q_ASSIGN U26 ( .B(clk), .A(\g.we_clk [16364]));
Q_ASSIGN U27 ( .B(clk), .A(\g.we_clk [16363]));
Q_ASSIGN U28 ( .B(clk), .A(\g.we_clk [16362]));
Q_ASSIGN U29 ( .B(clk), .A(\g.we_clk [16361]));
Q_ASSIGN U30 ( .B(clk), .A(\g.we_clk [16360]));
Q_ASSIGN U31 ( .B(clk), .A(\g.we_clk [16359]));
Q_ASSIGN U32 ( .B(clk), .A(\g.we_clk [16358]));
Q_ASSIGN U33 ( .B(clk), .A(\g.we_clk [16357]));
Q_ASSIGN U34 ( .B(clk), .A(\g.we_clk [16356]));
Q_ASSIGN U35 ( .B(clk), .A(\g.we_clk [16355]));
Q_ASSIGN U36 ( .B(clk), .A(\g.we_clk [16354]));
Q_ASSIGN U37 ( .B(clk), .A(\g.we_clk [16353]));
Q_ASSIGN U38 ( .B(clk), .A(\g.we_clk [16352]));
Q_ASSIGN U39 ( .B(clk), .A(\g.we_clk [16351]));
Q_ASSIGN U40 ( .B(clk), .A(\g.we_clk [16350]));
Q_ASSIGN U41 ( .B(clk), .A(\g.we_clk [16349]));
Q_ASSIGN U42 ( .B(clk), .A(\g.we_clk [16348]));
Q_ASSIGN U43 ( .B(clk), .A(\g.we_clk [16347]));
Q_ASSIGN U44 ( .B(clk), .A(\g.we_clk [16346]));
Q_ASSIGN U45 ( .B(clk), .A(\g.we_clk [16345]));
Q_ASSIGN U46 ( .B(clk), .A(\g.we_clk [16344]));
Q_ASSIGN U47 ( .B(clk), .A(\g.we_clk [16343]));
Q_ASSIGN U48 ( .B(clk), .A(\g.we_clk [16342]));
Q_ASSIGN U49 ( .B(clk), .A(\g.we_clk [16341]));
Q_ASSIGN U50 ( .B(clk), .A(\g.we_clk [16340]));
Q_ASSIGN U51 ( .B(clk), .A(\g.we_clk [16339]));
Q_ASSIGN U52 ( .B(clk), .A(\g.we_clk [16338]));
Q_ASSIGN U53 ( .B(clk), .A(\g.we_clk [16337]));
Q_ASSIGN U54 ( .B(clk), .A(\g.we_clk [16336]));
Q_ASSIGN U55 ( .B(clk), .A(\g.we_clk [16335]));
Q_ASSIGN U56 ( .B(clk), .A(\g.we_clk [16334]));
Q_ASSIGN U57 ( .B(clk), .A(\g.we_clk [16333]));
Q_ASSIGN U58 ( .B(clk), .A(\g.we_clk [16332]));
Q_ASSIGN U59 ( .B(clk), .A(\g.we_clk [16331]));
Q_ASSIGN U60 ( .B(clk), .A(\g.we_clk [16330]));
Q_ASSIGN U61 ( .B(clk), .A(\g.we_clk [16329]));
Q_ASSIGN U62 ( .B(clk), .A(\g.we_clk [16328]));
Q_ASSIGN U63 ( .B(clk), .A(\g.we_clk [16327]));
Q_ASSIGN U64 ( .B(clk), .A(\g.we_clk [16326]));
Q_ASSIGN U65 ( .B(clk), .A(\g.we_clk [16325]));
Q_ASSIGN U66 ( .B(clk), .A(\g.we_clk [16324]));
Q_ASSIGN U67 ( .B(clk), .A(\g.we_clk [16323]));
Q_ASSIGN U68 ( .B(clk), .A(\g.we_clk [16322]));
Q_ASSIGN U69 ( .B(clk), .A(\g.we_clk [16321]));
Q_ASSIGN U70 ( .B(clk), .A(\g.we_clk [16320]));
Q_ASSIGN U71 ( .B(clk), .A(\g.we_clk [16319]));
Q_ASSIGN U72 ( .B(clk), .A(\g.we_clk [16318]));
Q_ASSIGN U73 ( .B(clk), .A(\g.we_clk [16317]));
Q_ASSIGN U74 ( .B(clk), .A(\g.we_clk [16316]));
Q_ASSIGN U75 ( .B(clk), .A(\g.we_clk [16315]));
Q_ASSIGN U76 ( .B(clk), .A(\g.we_clk [16314]));
Q_ASSIGN U77 ( .B(clk), .A(\g.we_clk [16313]));
Q_ASSIGN U78 ( .B(clk), .A(\g.we_clk [16312]));
Q_ASSIGN U79 ( .B(clk), .A(\g.we_clk [16311]));
Q_ASSIGN U80 ( .B(clk), .A(\g.we_clk [16310]));
Q_ASSIGN U81 ( .B(clk), .A(\g.we_clk [16309]));
Q_ASSIGN U82 ( .B(clk), .A(\g.we_clk [16308]));
Q_ASSIGN U83 ( .B(clk), .A(\g.we_clk [16307]));
Q_ASSIGN U84 ( .B(clk), .A(\g.we_clk [16306]));
Q_ASSIGN U85 ( .B(clk), .A(\g.we_clk [16305]));
Q_ASSIGN U86 ( .B(clk), .A(\g.we_clk [16304]));
Q_ASSIGN U87 ( .B(clk), .A(\g.we_clk [16303]));
Q_ASSIGN U88 ( .B(clk), .A(\g.we_clk [16302]));
Q_ASSIGN U89 ( .B(clk), .A(\g.we_clk [16301]));
Q_ASSIGN U90 ( .B(clk), .A(\g.we_clk [16300]));
Q_ASSIGN U91 ( .B(clk), .A(\g.we_clk [16299]));
Q_ASSIGN U92 ( .B(clk), .A(\g.we_clk [16298]));
Q_ASSIGN U93 ( .B(clk), .A(\g.we_clk [16297]));
Q_ASSIGN U94 ( .B(clk), .A(\g.we_clk [16296]));
Q_ASSIGN U95 ( .B(clk), .A(\g.we_clk [16295]));
Q_ASSIGN U96 ( .B(clk), .A(\g.we_clk [16294]));
Q_ASSIGN U97 ( .B(clk), .A(\g.we_clk [16293]));
Q_ASSIGN U98 ( .B(clk), .A(\g.we_clk [16292]));
Q_ASSIGN U99 ( .B(clk), .A(\g.we_clk [16291]));
Q_ASSIGN U100 ( .B(clk), .A(\g.we_clk [16290]));
Q_ASSIGN U101 ( .B(clk), .A(\g.we_clk [16289]));
Q_ASSIGN U102 ( .B(clk), .A(\g.we_clk [16288]));
Q_ASSIGN U103 ( .B(clk), .A(\g.we_clk [16287]));
Q_ASSIGN U104 ( .B(clk), .A(\g.we_clk [16286]));
Q_ASSIGN U105 ( .B(clk), .A(\g.we_clk [16285]));
Q_ASSIGN U106 ( .B(clk), .A(\g.we_clk [16284]));
Q_ASSIGN U107 ( .B(clk), .A(\g.we_clk [16283]));
Q_ASSIGN U108 ( .B(clk), .A(\g.we_clk [16282]));
Q_ASSIGN U109 ( .B(clk), .A(\g.we_clk [16281]));
Q_ASSIGN U110 ( .B(clk), .A(\g.we_clk [16280]));
Q_ASSIGN U111 ( .B(clk), .A(\g.we_clk [16279]));
Q_ASSIGN U112 ( .B(clk), .A(\g.we_clk [16278]));
Q_ASSIGN U113 ( .B(clk), .A(\g.we_clk [16277]));
Q_ASSIGN U114 ( .B(clk), .A(\g.we_clk [16276]));
Q_ASSIGN U115 ( .B(clk), .A(\g.we_clk [16275]));
Q_ASSIGN U116 ( .B(clk), .A(\g.we_clk [16274]));
Q_ASSIGN U117 ( .B(clk), .A(\g.we_clk [16273]));
Q_ASSIGN U118 ( .B(clk), .A(\g.we_clk [16272]));
Q_ASSIGN U119 ( .B(clk), .A(\g.we_clk [16271]));
Q_ASSIGN U120 ( .B(clk), .A(\g.we_clk [16270]));
Q_ASSIGN U121 ( .B(clk), .A(\g.we_clk [16269]));
Q_ASSIGN U122 ( .B(clk), .A(\g.we_clk [16268]));
Q_ASSIGN U123 ( .B(clk), .A(\g.we_clk [16267]));
Q_ASSIGN U124 ( .B(clk), .A(\g.we_clk [16266]));
Q_ASSIGN U125 ( .B(clk), .A(\g.we_clk [16265]));
Q_ASSIGN U126 ( .B(clk), .A(\g.we_clk [16264]));
Q_ASSIGN U127 ( .B(clk), .A(\g.we_clk [16263]));
Q_ASSIGN U128 ( .B(clk), .A(\g.we_clk [16262]));
Q_ASSIGN U129 ( .B(clk), .A(\g.we_clk [16261]));
Q_ASSIGN U130 ( .B(clk), .A(\g.we_clk [16260]));
Q_ASSIGN U131 ( .B(clk), .A(\g.we_clk [16259]));
Q_ASSIGN U132 ( .B(clk), .A(\g.we_clk [16258]));
Q_ASSIGN U133 ( .B(clk), .A(\g.we_clk [16257]));
Q_ASSIGN U134 ( .B(clk), .A(\g.we_clk [16256]));
Q_ASSIGN U135 ( .B(clk), .A(\g.we_clk [16255]));
Q_ASSIGN U136 ( .B(clk), .A(\g.we_clk [16254]));
Q_ASSIGN U137 ( .B(clk), .A(\g.we_clk [16253]));
Q_ASSIGN U138 ( .B(clk), .A(\g.we_clk [16252]));
Q_ASSIGN U139 ( .B(clk), .A(\g.we_clk [16251]));
Q_ASSIGN U140 ( .B(clk), .A(\g.we_clk [16250]));
Q_ASSIGN U141 ( .B(clk), .A(\g.we_clk [16249]));
Q_ASSIGN U142 ( .B(clk), .A(\g.we_clk [16248]));
Q_ASSIGN U143 ( .B(clk), .A(\g.we_clk [16247]));
Q_ASSIGN U144 ( .B(clk), .A(\g.we_clk [16246]));
Q_ASSIGN U145 ( .B(clk), .A(\g.we_clk [16245]));
Q_ASSIGN U146 ( .B(clk), .A(\g.we_clk [16244]));
Q_ASSIGN U147 ( .B(clk), .A(\g.we_clk [16243]));
Q_ASSIGN U148 ( .B(clk), .A(\g.we_clk [16242]));
Q_ASSIGN U149 ( .B(clk), .A(\g.we_clk [16241]));
Q_ASSIGN U150 ( .B(clk), .A(\g.we_clk [16240]));
Q_ASSIGN U151 ( .B(clk), .A(\g.we_clk [16239]));
Q_ASSIGN U152 ( .B(clk), .A(\g.we_clk [16238]));
Q_ASSIGN U153 ( .B(clk), .A(\g.we_clk [16237]));
Q_ASSIGN U154 ( .B(clk), .A(\g.we_clk [16236]));
Q_ASSIGN U155 ( .B(clk), .A(\g.we_clk [16235]));
Q_ASSIGN U156 ( .B(clk), .A(\g.we_clk [16234]));
Q_ASSIGN U157 ( .B(clk), .A(\g.we_clk [16233]));
Q_ASSIGN U158 ( .B(clk), .A(\g.we_clk [16232]));
Q_ASSIGN U159 ( .B(clk), .A(\g.we_clk [16231]));
Q_ASSIGN U160 ( .B(clk), .A(\g.we_clk [16230]));
Q_ASSIGN U161 ( .B(clk), .A(\g.we_clk [16229]));
Q_ASSIGN U162 ( .B(clk), .A(\g.we_clk [16228]));
Q_ASSIGN U163 ( .B(clk), .A(\g.we_clk [16227]));
Q_ASSIGN U164 ( .B(clk), .A(\g.we_clk [16226]));
Q_ASSIGN U165 ( .B(clk), .A(\g.we_clk [16225]));
Q_ASSIGN U166 ( .B(clk), .A(\g.we_clk [16224]));
Q_ASSIGN U167 ( .B(clk), .A(\g.we_clk [16223]));
Q_ASSIGN U168 ( .B(clk), .A(\g.we_clk [16222]));
Q_ASSIGN U169 ( .B(clk), .A(\g.we_clk [16221]));
Q_ASSIGN U170 ( .B(clk), .A(\g.we_clk [16220]));
Q_ASSIGN U171 ( .B(clk), .A(\g.we_clk [16219]));
Q_ASSIGN U172 ( .B(clk), .A(\g.we_clk [16218]));
Q_ASSIGN U173 ( .B(clk), .A(\g.we_clk [16217]));
Q_ASSIGN U174 ( .B(clk), .A(\g.we_clk [16216]));
Q_ASSIGN U175 ( .B(clk), .A(\g.we_clk [16215]));
Q_ASSIGN U176 ( .B(clk), .A(\g.we_clk [16214]));
Q_ASSIGN U177 ( .B(clk), .A(\g.we_clk [16213]));
Q_ASSIGN U178 ( .B(clk), .A(\g.we_clk [16212]));
Q_ASSIGN U179 ( .B(clk), .A(\g.we_clk [16211]));
Q_ASSIGN U180 ( .B(clk), .A(\g.we_clk [16210]));
Q_ASSIGN U181 ( .B(clk), .A(\g.we_clk [16209]));
Q_ASSIGN U182 ( .B(clk), .A(\g.we_clk [16208]));
Q_ASSIGN U183 ( .B(clk), .A(\g.we_clk [16207]));
Q_ASSIGN U184 ( .B(clk), .A(\g.we_clk [16206]));
Q_ASSIGN U185 ( .B(clk), .A(\g.we_clk [16205]));
Q_ASSIGN U186 ( .B(clk), .A(\g.we_clk [16204]));
Q_ASSIGN U187 ( .B(clk), .A(\g.we_clk [16203]));
Q_ASSIGN U188 ( .B(clk), .A(\g.we_clk [16202]));
Q_ASSIGN U189 ( .B(clk), .A(\g.we_clk [16201]));
Q_ASSIGN U190 ( .B(clk), .A(\g.we_clk [16200]));
Q_ASSIGN U191 ( .B(clk), .A(\g.we_clk [16199]));
Q_ASSIGN U192 ( .B(clk), .A(\g.we_clk [16198]));
Q_ASSIGN U193 ( .B(clk), .A(\g.we_clk [16197]));
Q_ASSIGN U194 ( .B(clk), .A(\g.we_clk [16196]));
Q_ASSIGN U195 ( .B(clk), .A(\g.we_clk [16195]));
Q_ASSIGN U196 ( .B(clk), .A(\g.we_clk [16194]));
Q_ASSIGN U197 ( .B(clk), .A(\g.we_clk [16193]));
Q_ASSIGN U198 ( .B(clk), .A(\g.we_clk [16192]));
Q_ASSIGN U199 ( .B(clk), .A(\g.we_clk [16191]));
Q_ASSIGN U200 ( .B(clk), .A(\g.we_clk [16190]));
Q_ASSIGN U201 ( .B(clk), .A(\g.we_clk [16189]));
Q_ASSIGN U202 ( .B(clk), .A(\g.we_clk [16188]));
Q_ASSIGN U203 ( .B(clk), .A(\g.we_clk [16187]));
Q_ASSIGN U204 ( .B(clk), .A(\g.we_clk [16186]));
Q_ASSIGN U205 ( .B(clk), .A(\g.we_clk [16185]));
Q_ASSIGN U206 ( .B(clk), .A(\g.we_clk [16184]));
Q_ASSIGN U207 ( .B(clk), .A(\g.we_clk [16183]));
Q_ASSIGN U208 ( .B(clk), .A(\g.we_clk [16182]));
Q_ASSIGN U209 ( .B(clk), .A(\g.we_clk [16181]));
Q_ASSIGN U210 ( .B(clk), .A(\g.we_clk [16180]));
Q_ASSIGN U211 ( .B(clk), .A(\g.we_clk [16179]));
Q_ASSIGN U212 ( .B(clk), .A(\g.we_clk [16178]));
Q_ASSIGN U213 ( .B(clk), .A(\g.we_clk [16177]));
Q_ASSIGN U214 ( .B(clk), .A(\g.we_clk [16176]));
Q_ASSIGN U215 ( .B(clk), .A(\g.we_clk [16175]));
Q_ASSIGN U216 ( .B(clk), .A(\g.we_clk [16174]));
Q_ASSIGN U217 ( .B(clk), .A(\g.we_clk [16173]));
Q_ASSIGN U218 ( .B(clk), .A(\g.we_clk [16172]));
Q_ASSIGN U219 ( .B(clk), .A(\g.we_clk [16171]));
Q_ASSIGN U220 ( .B(clk), .A(\g.we_clk [16170]));
Q_ASSIGN U221 ( .B(clk), .A(\g.we_clk [16169]));
Q_ASSIGN U222 ( .B(clk), .A(\g.we_clk [16168]));
Q_ASSIGN U223 ( .B(clk), .A(\g.we_clk [16167]));
Q_ASSIGN U224 ( .B(clk), .A(\g.we_clk [16166]));
Q_ASSIGN U225 ( .B(clk), .A(\g.we_clk [16165]));
Q_ASSIGN U226 ( .B(clk), .A(\g.we_clk [16164]));
Q_ASSIGN U227 ( .B(clk), .A(\g.we_clk [16163]));
Q_ASSIGN U228 ( .B(clk), .A(\g.we_clk [16162]));
Q_ASSIGN U229 ( .B(clk), .A(\g.we_clk [16161]));
Q_ASSIGN U230 ( .B(clk), .A(\g.we_clk [16160]));
Q_ASSIGN U231 ( .B(clk), .A(\g.we_clk [16159]));
Q_ASSIGN U232 ( .B(clk), .A(\g.we_clk [16158]));
Q_ASSIGN U233 ( .B(clk), .A(\g.we_clk [16157]));
Q_ASSIGN U234 ( .B(clk), .A(\g.we_clk [16156]));
Q_ASSIGN U235 ( .B(clk), .A(\g.we_clk [16155]));
Q_ASSIGN U236 ( .B(clk), .A(\g.we_clk [16154]));
Q_ASSIGN U237 ( .B(clk), .A(\g.we_clk [16153]));
Q_ASSIGN U238 ( .B(clk), .A(\g.we_clk [16152]));
Q_ASSIGN U239 ( .B(clk), .A(\g.we_clk [16151]));
Q_ASSIGN U240 ( .B(clk), .A(\g.we_clk [16150]));
Q_ASSIGN U241 ( .B(clk), .A(\g.we_clk [16149]));
Q_ASSIGN U242 ( .B(clk), .A(\g.we_clk [16148]));
Q_ASSIGN U243 ( .B(clk), .A(\g.we_clk [16147]));
Q_ASSIGN U244 ( .B(clk), .A(\g.we_clk [16146]));
Q_ASSIGN U245 ( .B(clk), .A(\g.we_clk [16145]));
Q_ASSIGN U246 ( .B(clk), .A(\g.we_clk [16144]));
Q_ASSIGN U247 ( .B(clk), .A(\g.we_clk [16143]));
Q_ASSIGN U248 ( .B(clk), .A(\g.we_clk [16142]));
Q_ASSIGN U249 ( .B(clk), .A(\g.we_clk [16141]));
Q_ASSIGN U250 ( .B(clk), .A(\g.we_clk [16140]));
Q_ASSIGN U251 ( .B(clk), .A(\g.we_clk [16139]));
Q_ASSIGN U252 ( .B(clk), .A(\g.we_clk [16138]));
Q_ASSIGN U253 ( .B(clk), .A(\g.we_clk [16137]));
Q_ASSIGN U254 ( .B(clk), .A(\g.we_clk [16136]));
Q_ASSIGN U255 ( .B(clk), .A(\g.we_clk [16135]));
Q_ASSIGN U256 ( .B(clk), .A(\g.we_clk [16134]));
Q_ASSIGN U257 ( .B(clk), .A(\g.we_clk [16133]));
Q_ASSIGN U258 ( .B(clk), .A(\g.we_clk [16132]));
Q_ASSIGN U259 ( .B(clk), .A(\g.we_clk [16131]));
Q_ASSIGN U260 ( .B(clk), .A(\g.we_clk [16130]));
Q_ASSIGN U261 ( .B(clk), .A(\g.we_clk [16129]));
Q_ASSIGN U262 ( .B(clk), .A(\g.we_clk [16128]));
Q_ASSIGN U263 ( .B(clk), .A(\g.we_clk [16127]));
Q_ASSIGN U264 ( .B(clk), .A(\g.we_clk [16126]));
Q_ASSIGN U265 ( .B(clk), .A(\g.we_clk [16125]));
Q_ASSIGN U266 ( .B(clk), .A(\g.we_clk [16124]));
Q_ASSIGN U267 ( .B(clk), .A(\g.we_clk [16123]));
Q_ASSIGN U268 ( .B(clk), .A(\g.we_clk [16122]));
Q_ASSIGN U269 ( .B(clk), .A(\g.we_clk [16121]));
Q_ASSIGN U270 ( .B(clk), .A(\g.we_clk [16120]));
Q_ASSIGN U271 ( .B(clk), .A(\g.we_clk [16119]));
Q_ASSIGN U272 ( .B(clk), .A(\g.we_clk [16118]));
Q_ASSIGN U273 ( .B(clk), .A(\g.we_clk [16117]));
Q_ASSIGN U274 ( .B(clk), .A(\g.we_clk [16116]));
Q_ASSIGN U275 ( .B(clk), .A(\g.we_clk [16115]));
Q_ASSIGN U276 ( .B(clk), .A(\g.we_clk [16114]));
Q_ASSIGN U277 ( .B(clk), .A(\g.we_clk [16113]));
Q_ASSIGN U278 ( .B(clk), .A(\g.we_clk [16112]));
Q_ASSIGN U279 ( .B(clk), .A(\g.we_clk [16111]));
Q_ASSIGN U280 ( .B(clk), .A(\g.we_clk [16110]));
Q_ASSIGN U281 ( .B(clk), .A(\g.we_clk [16109]));
Q_ASSIGN U282 ( .B(clk), .A(\g.we_clk [16108]));
Q_ASSIGN U283 ( .B(clk), .A(\g.we_clk [16107]));
Q_ASSIGN U284 ( .B(clk), .A(\g.we_clk [16106]));
Q_ASSIGN U285 ( .B(clk), .A(\g.we_clk [16105]));
Q_ASSIGN U286 ( .B(clk), .A(\g.we_clk [16104]));
Q_ASSIGN U287 ( .B(clk), .A(\g.we_clk [16103]));
Q_ASSIGN U288 ( .B(clk), .A(\g.we_clk [16102]));
Q_ASSIGN U289 ( .B(clk), .A(\g.we_clk [16101]));
Q_ASSIGN U290 ( .B(clk), .A(\g.we_clk [16100]));
Q_ASSIGN U291 ( .B(clk), .A(\g.we_clk [16099]));
Q_ASSIGN U292 ( .B(clk), .A(\g.we_clk [16098]));
Q_ASSIGN U293 ( .B(clk), .A(\g.we_clk [16097]));
Q_ASSIGN U294 ( .B(clk), .A(\g.we_clk [16096]));
Q_ASSIGN U295 ( .B(clk), .A(\g.we_clk [16095]));
Q_ASSIGN U296 ( .B(clk), .A(\g.we_clk [16094]));
Q_ASSIGN U297 ( .B(clk), .A(\g.we_clk [16093]));
Q_ASSIGN U298 ( .B(clk), .A(\g.we_clk [16092]));
Q_ASSIGN U299 ( .B(clk), .A(\g.we_clk [16091]));
Q_ASSIGN U300 ( .B(clk), .A(\g.we_clk [16090]));
Q_ASSIGN U301 ( .B(clk), .A(\g.we_clk [16089]));
Q_ASSIGN U302 ( .B(clk), .A(\g.we_clk [16088]));
Q_ASSIGN U303 ( .B(clk), .A(\g.we_clk [16087]));
Q_ASSIGN U304 ( .B(clk), .A(\g.we_clk [16086]));
Q_ASSIGN U305 ( .B(clk), .A(\g.we_clk [16085]));
Q_ASSIGN U306 ( .B(clk), .A(\g.we_clk [16084]));
Q_ASSIGN U307 ( .B(clk), .A(\g.we_clk [16083]));
Q_ASSIGN U308 ( .B(clk), .A(\g.we_clk [16082]));
Q_ASSIGN U309 ( .B(clk), .A(\g.we_clk [16081]));
Q_ASSIGN U310 ( .B(clk), .A(\g.we_clk [16080]));
Q_ASSIGN U311 ( .B(clk), .A(\g.we_clk [16079]));
Q_ASSIGN U312 ( .B(clk), .A(\g.we_clk [16078]));
Q_ASSIGN U313 ( .B(clk), .A(\g.we_clk [16077]));
Q_ASSIGN U314 ( .B(clk), .A(\g.we_clk [16076]));
Q_ASSIGN U315 ( .B(clk), .A(\g.we_clk [16075]));
Q_ASSIGN U316 ( .B(clk), .A(\g.we_clk [16074]));
Q_ASSIGN U317 ( .B(clk), .A(\g.we_clk [16073]));
Q_ASSIGN U318 ( .B(clk), .A(\g.we_clk [16072]));
Q_ASSIGN U319 ( .B(clk), .A(\g.we_clk [16071]));
Q_ASSIGN U320 ( .B(clk), .A(\g.we_clk [16070]));
Q_ASSIGN U321 ( .B(clk), .A(\g.we_clk [16069]));
Q_ASSIGN U322 ( .B(clk), .A(\g.we_clk [16068]));
Q_ASSIGN U323 ( .B(clk), .A(\g.we_clk [16067]));
Q_ASSIGN U324 ( .B(clk), .A(\g.we_clk [16066]));
Q_ASSIGN U325 ( .B(clk), .A(\g.we_clk [16065]));
Q_ASSIGN U326 ( .B(clk), .A(\g.we_clk [16064]));
Q_ASSIGN U327 ( .B(clk), .A(\g.we_clk [16063]));
Q_ASSIGN U328 ( .B(clk), .A(\g.we_clk [16062]));
Q_ASSIGN U329 ( .B(clk), .A(\g.we_clk [16061]));
Q_ASSIGN U330 ( .B(clk), .A(\g.we_clk [16060]));
Q_ASSIGN U331 ( .B(clk), .A(\g.we_clk [16059]));
Q_ASSIGN U332 ( .B(clk), .A(\g.we_clk [16058]));
Q_ASSIGN U333 ( .B(clk), .A(\g.we_clk [16057]));
Q_ASSIGN U334 ( .B(clk), .A(\g.we_clk [16056]));
Q_ASSIGN U335 ( .B(clk), .A(\g.we_clk [16055]));
Q_ASSIGN U336 ( .B(clk), .A(\g.we_clk [16054]));
Q_ASSIGN U337 ( .B(clk), .A(\g.we_clk [16053]));
Q_ASSIGN U338 ( .B(clk), .A(\g.we_clk [16052]));
Q_ASSIGN U339 ( .B(clk), .A(\g.we_clk [16051]));
Q_ASSIGN U340 ( .B(clk), .A(\g.we_clk [16050]));
Q_ASSIGN U341 ( .B(clk), .A(\g.we_clk [16049]));
Q_ASSIGN U342 ( .B(clk), .A(\g.we_clk [16048]));
Q_ASSIGN U343 ( .B(clk), .A(\g.we_clk [16047]));
Q_ASSIGN U344 ( .B(clk), .A(\g.we_clk [16046]));
Q_ASSIGN U345 ( .B(clk), .A(\g.we_clk [16045]));
Q_ASSIGN U346 ( .B(clk), .A(\g.we_clk [16044]));
Q_ASSIGN U347 ( .B(clk), .A(\g.we_clk [16043]));
Q_ASSIGN U348 ( .B(clk), .A(\g.we_clk [16042]));
Q_ASSIGN U349 ( .B(clk), .A(\g.we_clk [16041]));
Q_ASSIGN U350 ( .B(clk), .A(\g.we_clk [16040]));
Q_ASSIGN U351 ( .B(clk), .A(\g.we_clk [16039]));
Q_ASSIGN U352 ( .B(clk), .A(\g.we_clk [16038]));
Q_ASSIGN U353 ( .B(clk), .A(\g.we_clk [16037]));
Q_ASSIGN U354 ( .B(clk), .A(\g.we_clk [16036]));
Q_ASSIGN U355 ( .B(clk), .A(\g.we_clk [16035]));
Q_ASSIGN U356 ( .B(clk), .A(\g.we_clk [16034]));
Q_ASSIGN U357 ( .B(clk), .A(\g.we_clk [16033]));
Q_ASSIGN U358 ( .B(clk), .A(\g.we_clk [16032]));
Q_ASSIGN U359 ( .B(clk), .A(\g.we_clk [16031]));
Q_ASSIGN U360 ( .B(clk), .A(\g.we_clk [16030]));
Q_ASSIGN U361 ( .B(clk), .A(\g.we_clk [16029]));
Q_ASSIGN U362 ( .B(clk), .A(\g.we_clk [16028]));
Q_ASSIGN U363 ( .B(clk), .A(\g.we_clk [16027]));
Q_ASSIGN U364 ( .B(clk), .A(\g.we_clk [16026]));
Q_ASSIGN U365 ( .B(clk), .A(\g.we_clk [16025]));
Q_ASSIGN U366 ( .B(clk), .A(\g.we_clk [16024]));
Q_ASSIGN U367 ( .B(clk), .A(\g.we_clk [16023]));
Q_ASSIGN U368 ( .B(clk), .A(\g.we_clk [16022]));
Q_ASSIGN U369 ( .B(clk), .A(\g.we_clk [16021]));
Q_ASSIGN U370 ( .B(clk), .A(\g.we_clk [16020]));
Q_ASSIGN U371 ( .B(clk), .A(\g.we_clk [16019]));
Q_ASSIGN U372 ( .B(clk), .A(\g.we_clk [16018]));
Q_ASSIGN U373 ( .B(clk), .A(\g.we_clk [16017]));
Q_ASSIGN U374 ( .B(clk), .A(\g.we_clk [16016]));
Q_ASSIGN U375 ( .B(clk), .A(\g.we_clk [16015]));
Q_ASSIGN U376 ( .B(clk), .A(\g.we_clk [16014]));
Q_ASSIGN U377 ( .B(clk), .A(\g.we_clk [16013]));
Q_ASSIGN U378 ( .B(clk), .A(\g.we_clk [16012]));
Q_ASSIGN U379 ( .B(clk), .A(\g.we_clk [16011]));
Q_ASSIGN U380 ( .B(clk), .A(\g.we_clk [16010]));
Q_ASSIGN U381 ( .B(clk), .A(\g.we_clk [16009]));
Q_ASSIGN U382 ( .B(clk), .A(\g.we_clk [16008]));
Q_ASSIGN U383 ( .B(clk), .A(\g.we_clk [16007]));
Q_ASSIGN U384 ( .B(clk), .A(\g.we_clk [16006]));
Q_ASSIGN U385 ( .B(clk), .A(\g.we_clk [16005]));
Q_ASSIGN U386 ( .B(clk), .A(\g.we_clk [16004]));
Q_ASSIGN U387 ( .B(clk), .A(\g.we_clk [16003]));
Q_ASSIGN U388 ( .B(clk), .A(\g.we_clk [16002]));
Q_ASSIGN U389 ( .B(clk), .A(\g.we_clk [16001]));
Q_ASSIGN U390 ( .B(clk), .A(\g.we_clk [16000]));
Q_ASSIGN U391 ( .B(clk), .A(\g.we_clk [15999]));
Q_ASSIGN U392 ( .B(clk), .A(\g.we_clk [15998]));
Q_ASSIGN U393 ( .B(clk), .A(\g.we_clk [15997]));
Q_ASSIGN U394 ( .B(clk), .A(\g.we_clk [15996]));
Q_ASSIGN U395 ( .B(clk), .A(\g.we_clk [15995]));
Q_ASSIGN U396 ( .B(clk), .A(\g.we_clk [15994]));
Q_ASSIGN U397 ( .B(clk), .A(\g.we_clk [15993]));
Q_ASSIGN U398 ( .B(clk), .A(\g.we_clk [15992]));
Q_ASSIGN U399 ( .B(clk), .A(\g.we_clk [15991]));
Q_ASSIGN U400 ( .B(clk), .A(\g.we_clk [15990]));
Q_ASSIGN U401 ( .B(clk), .A(\g.we_clk [15989]));
Q_ASSIGN U402 ( .B(clk), .A(\g.we_clk [15988]));
Q_ASSIGN U403 ( .B(clk), .A(\g.we_clk [15987]));
Q_ASSIGN U404 ( .B(clk), .A(\g.we_clk [15986]));
Q_ASSIGN U405 ( .B(clk), .A(\g.we_clk [15985]));
Q_ASSIGN U406 ( .B(clk), .A(\g.we_clk [15984]));
Q_ASSIGN U407 ( .B(clk), .A(\g.we_clk [15983]));
Q_ASSIGN U408 ( .B(clk), .A(\g.we_clk [15982]));
Q_ASSIGN U409 ( .B(clk), .A(\g.we_clk [15981]));
Q_ASSIGN U410 ( .B(clk), .A(\g.we_clk [15980]));
Q_ASSIGN U411 ( .B(clk), .A(\g.we_clk [15979]));
Q_ASSIGN U412 ( .B(clk), .A(\g.we_clk [15978]));
Q_ASSIGN U413 ( .B(clk), .A(\g.we_clk [15977]));
Q_ASSIGN U414 ( .B(clk), .A(\g.we_clk [15976]));
Q_ASSIGN U415 ( .B(clk), .A(\g.we_clk [15975]));
Q_ASSIGN U416 ( .B(clk), .A(\g.we_clk [15974]));
Q_ASSIGN U417 ( .B(clk), .A(\g.we_clk [15973]));
Q_ASSIGN U418 ( .B(clk), .A(\g.we_clk [15972]));
Q_ASSIGN U419 ( .B(clk), .A(\g.we_clk [15971]));
Q_ASSIGN U420 ( .B(clk), .A(\g.we_clk [15970]));
Q_ASSIGN U421 ( .B(clk), .A(\g.we_clk [15969]));
Q_ASSIGN U422 ( .B(clk), .A(\g.we_clk [15968]));
Q_ASSIGN U423 ( .B(clk), .A(\g.we_clk [15967]));
Q_ASSIGN U424 ( .B(clk), .A(\g.we_clk [15966]));
Q_ASSIGN U425 ( .B(clk), .A(\g.we_clk [15965]));
Q_ASSIGN U426 ( .B(clk), .A(\g.we_clk [15964]));
Q_ASSIGN U427 ( .B(clk), .A(\g.we_clk [15963]));
Q_ASSIGN U428 ( .B(clk), .A(\g.we_clk [15962]));
Q_ASSIGN U429 ( .B(clk), .A(\g.we_clk [15961]));
Q_ASSIGN U430 ( .B(clk), .A(\g.we_clk [15960]));
Q_ASSIGN U431 ( .B(clk), .A(\g.we_clk [15959]));
Q_ASSIGN U432 ( .B(clk), .A(\g.we_clk [15958]));
Q_ASSIGN U433 ( .B(clk), .A(\g.we_clk [15957]));
Q_ASSIGN U434 ( .B(clk), .A(\g.we_clk [15956]));
Q_ASSIGN U435 ( .B(clk), .A(\g.we_clk [15955]));
Q_ASSIGN U436 ( .B(clk), .A(\g.we_clk [15954]));
Q_ASSIGN U437 ( .B(clk), .A(\g.we_clk [15953]));
Q_ASSIGN U438 ( .B(clk), .A(\g.we_clk [15952]));
Q_ASSIGN U439 ( .B(clk), .A(\g.we_clk [15951]));
Q_ASSIGN U440 ( .B(clk), .A(\g.we_clk [15950]));
Q_ASSIGN U441 ( .B(clk), .A(\g.we_clk [15949]));
Q_ASSIGN U442 ( .B(clk), .A(\g.we_clk [15948]));
Q_ASSIGN U443 ( .B(clk), .A(\g.we_clk [15947]));
Q_ASSIGN U444 ( .B(clk), .A(\g.we_clk [15946]));
Q_ASSIGN U445 ( .B(clk), .A(\g.we_clk [15945]));
Q_ASSIGN U446 ( .B(clk), .A(\g.we_clk [15944]));
Q_ASSIGN U447 ( .B(clk), .A(\g.we_clk [15943]));
Q_ASSIGN U448 ( .B(clk), .A(\g.we_clk [15942]));
Q_ASSIGN U449 ( .B(clk), .A(\g.we_clk [15941]));
Q_ASSIGN U450 ( .B(clk), .A(\g.we_clk [15940]));
Q_ASSIGN U451 ( .B(clk), .A(\g.we_clk [15939]));
Q_ASSIGN U452 ( .B(clk), .A(\g.we_clk [15938]));
Q_ASSIGN U453 ( .B(clk), .A(\g.we_clk [15937]));
Q_ASSIGN U454 ( .B(clk), .A(\g.we_clk [15936]));
Q_ASSIGN U455 ( .B(clk), .A(\g.we_clk [15935]));
Q_ASSIGN U456 ( .B(clk), .A(\g.we_clk [15934]));
Q_ASSIGN U457 ( .B(clk), .A(\g.we_clk [15933]));
Q_ASSIGN U458 ( .B(clk), .A(\g.we_clk [15932]));
Q_ASSIGN U459 ( .B(clk), .A(\g.we_clk [15931]));
Q_ASSIGN U460 ( .B(clk), .A(\g.we_clk [15930]));
Q_ASSIGN U461 ( .B(clk), .A(\g.we_clk [15929]));
Q_ASSIGN U462 ( .B(clk), .A(\g.we_clk [15928]));
Q_ASSIGN U463 ( .B(clk), .A(\g.we_clk [15927]));
Q_ASSIGN U464 ( .B(clk), .A(\g.we_clk [15926]));
Q_ASSIGN U465 ( .B(clk), .A(\g.we_clk [15925]));
Q_ASSIGN U466 ( .B(clk), .A(\g.we_clk [15924]));
Q_ASSIGN U467 ( .B(clk), .A(\g.we_clk [15923]));
Q_ASSIGN U468 ( .B(clk), .A(\g.we_clk [15922]));
Q_ASSIGN U469 ( .B(clk), .A(\g.we_clk [15921]));
Q_ASSIGN U470 ( .B(clk), .A(\g.we_clk [15920]));
Q_ASSIGN U471 ( .B(clk), .A(\g.we_clk [15919]));
Q_ASSIGN U472 ( .B(clk), .A(\g.we_clk [15918]));
Q_ASSIGN U473 ( .B(clk), .A(\g.we_clk [15917]));
Q_ASSIGN U474 ( .B(clk), .A(\g.we_clk [15916]));
Q_ASSIGN U475 ( .B(clk), .A(\g.we_clk [15915]));
Q_ASSIGN U476 ( .B(clk), .A(\g.we_clk [15914]));
Q_ASSIGN U477 ( .B(clk), .A(\g.we_clk [15913]));
Q_ASSIGN U478 ( .B(clk), .A(\g.we_clk [15912]));
Q_ASSIGN U479 ( .B(clk), .A(\g.we_clk [15911]));
Q_ASSIGN U480 ( .B(clk), .A(\g.we_clk [15910]));
Q_ASSIGN U481 ( .B(clk), .A(\g.we_clk [15909]));
Q_ASSIGN U482 ( .B(clk), .A(\g.we_clk [15908]));
Q_ASSIGN U483 ( .B(clk), .A(\g.we_clk [15907]));
Q_ASSIGN U484 ( .B(clk), .A(\g.we_clk [15906]));
Q_ASSIGN U485 ( .B(clk), .A(\g.we_clk [15905]));
Q_ASSIGN U486 ( .B(clk), .A(\g.we_clk [15904]));
Q_ASSIGN U487 ( .B(clk), .A(\g.we_clk [15903]));
Q_ASSIGN U488 ( .B(clk), .A(\g.we_clk [15902]));
Q_ASSIGN U489 ( .B(clk), .A(\g.we_clk [15901]));
Q_ASSIGN U490 ( .B(clk), .A(\g.we_clk [15900]));
Q_ASSIGN U491 ( .B(clk), .A(\g.we_clk [15899]));
Q_ASSIGN U492 ( .B(clk), .A(\g.we_clk [15898]));
Q_ASSIGN U493 ( .B(clk), .A(\g.we_clk [15897]));
Q_ASSIGN U494 ( .B(clk), .A(\g.we_clk [15896]));
Q_ASSIGN U495 ( .B(clk), .A(\g.we_clk [15895]));
Q_ASSIGN U496 ( .B(clk), .A(\g.we_clk [15894]));
Q_ASSIGN U497 ( .B(clk), .A(\g.we_clk [15893]));
Q_ASSIGN U498 ( .B(clk), .A(\g.we_clk [15892]));
Q_ASSIGN U499 ( .B(clk), .A(\g.we_clk [15891]));
Q_ASSIGN U500 ( .B(clk), .A(\g.we_clk [15890]));
Q_ASSIGN U501 ( .B(clk), .A(\g.we_clk [15889]));
Q_ASSIGN U502 ( .B(clk), .A(\g.we_clk [15888]));
Q_ASSIGN U503 ( .B(clk), .A(\g.we_clk [15887]));
Q_ASSIGN U504 ( .B(clk), .A(\g.we_clk [15886]));
Q_ASSIGN U505 ( .B(clk), .A(\g.we_clk [15885]));
Q_ASSIGN U506 ( .B(clk), .A(\g.we_clk [15884]));
Q_ASSIGN U507 ( .B(clk), .A(\g.we_clk [15883]));
Q_ASSIGN U508 ( .B(clk), .A(\g.we_clk [15882]));
Q_ASSIGN U509 ( .B(clk), .A(\g.we_clk [15881]));
Q_ASSIGN U510 ( .B(clk), .A(\g.we_clk [15880]));
Q_ASSIGN U511 ( .B(clk), .A(\g.we_clk [15879]));
Q_ASSIGN U512 ( .B(clk), .A(\g.we_clk [15878]));
Q_ASSIGN U513 ( .B(clk), .A(\g.we_clk [15877]));
Q_ASSIGN U514 ( .B(clk), .A(\g.we_clk [15876]));
Q_ASSIGN U515 ( .B(clk), .A(\g.we_clk [15875]));
Q_ASSIGN U516 ( .B(clk), .A(\g.we_clk [15874]));
Q_ASSIGN U517 ( .B(clk), .A(\g.we_clk [15873]));
Q_ASSIGN U518 ( .B(clk), .A(\g.we_clk [15872]));
Q_ASSIGN U519 ( .B(clk), .A(\g.we_clk [15871]));
Q_ASSIGN U520 ( .B(clk), .A(\g.we_clk [15870]));
Q_ASSIGN U521 ( .B(clk), .A(\g.we_clk [15869]));
Q_ASSIGN U522 ( .B(clk), .A(\g.we_clk [15868]));
Q_ASSIGN U523 ( .B(clk), .A(\g.we_clk [15867]));
Q_ASSIGN U524 ( .B(clk), .A(\g.we_clk [15866]));
Q_ASSIGN U525 ( .B(clk), .A(\g.we_clk [15865]));
Q_ASSIGN U526 ( .B(clk), .A(\g.we_clk [15864]));
Q_ASSIGN U527 ( .B(clk), .A(\g.we_clk [15863]));
Q_ASSIGN U528 ( .B(clk), .A(\g.we_clk [15862]));
Q_ASSIGN U529 ( .B(clk), .A(\g.we_clk [15861]));
Q_ASSIGN U530 ( .B(clk), .A(\g.we_clk [15860]));
Q_ASSIGN U531 ( .B(clk), .A(\g.we_clk [15859]));
Q_ASSIGN U532 ( .B(clk), .A(\g.we_clk [15858]));
Q_ASSIGN U533 ( .B(clk), .A(\g.we_clk [15857]));
Q_ASSIGN U534 ( .B(clk), .A(\g.we_clk [15856]));
Q_ASSIGN U535 ( .B(clk), .A(\g.we_clk [15855]));
Q_ASSIGN U536 ( .B(clk), .A(\g.we_clk [15854]));
Q_ASSIGN U537 ( .B(clk), .A(\g.we_clk [15853]));
Q_ASSIGN U538 ( .B(clk), .A(\g.we_clk [15852]));
Q_ASSIGN U539 ( .B(clk), .A(\g.we_clk [15851]));
Q_ASSIGN U540 ( .B(clk), .A(\g.we_clk [15850]));
Q_ASSIGN U541 ( .B(clk), .A(\g.we_clk [15849]));
Q_ASSIGN U542 ( .B(clk), .A(\g.we_clk [15848]));
Q_ASSIGN U543 ( .B(clk), .A(\g.we_clk [15847]));
Q_ASSIGN U544 ( .B(clk), .A(\g.we_clk [15846]));
Q_ASSIGN U545 ( .B(clk), .A(\g.we_clk [15845]));
Q_ASSIGN U546 ( .B(clk), .A(\g.we_clk [15844]));
Q_ASSIGN U547 ( .B(clk), .A(\g.we_clk [15843]));
Q_ASSIGN U548 ( .B(clk), .A(\g.we_clk [15842]));
Q_ASSIGN U549 ( .B(clk), .A(\g.we_clk [15841]));
Q_ASSIGN U550 ( .B(clk), .A(\g.we_clk [15840]));
Q_ASSIGN U551 ( .B(clk), .A(\g.we_clk [15839]));
Q_ASSIGN U552 ( .B(clk), .A(\g.we_clk [15838]));
Q_ASSIGN U553 ( .B(clk), .A(\g.we_clk [15837]));
Q_ASSIGN U554 ( .B(clk), .A(\g.we_clk [15836]));
Q_ASSIGN U555 ( .B(clk), .A(\g.we_clk [15835]));
Q_ASSIGN U556 ( .B(clk), .A(\g.we_clk [15834]));
Q_ASSIGN U557 ( .B(clk), .A(\g.we_clk [15833]));
Q_ASSIGN U558 ( .B(clk), .A(\g.we_clk [15832]));
Q_ASSIGN U559 ( .B(clk), .A(\g.we_clk [15831]));
Q_ASSIGN U560 ( .B(clk), .A(\g.we_clk [15830]));
Q_ASSIGN U561 ( .B(clk), .A(\g.we_clk [15829]));
Q_ASSIGN U562 ( .B(clk), .A(\g.we_clk [15828]));
Q_ASSIGN U563 ( .B(clk), .A(\g.we_clk [15827]));
Q_ASSIGN U564 ( .B(clk), .A(\g.we_clk [15826]));
Q_ASSIGN U565 ( .B(clk), .A(\g.we_clk [15825]));
Q_ASSIGN U566 ( .B(clk), .A(\g.we_clk [15824]));
Q_ASSIGN U567 ( .B(clk), .A(\g.we_clk [15823]));
Q_ASSIGN U568 ( .B(clk), .A(\g.we_clk [15822]));
Q_ASSIGN U569 ( .B(clk), .A(\g.we_clk [15821]));
Q_ASSIGN U570 ( .B(clk), .A(\g.we_clk [15820]));
Q_ASSIGN U571 ( .B(clk), .A(\g.we_clk [15819]));
Q_ASSIGN U572 ( .B(clk), .A(\g.we_clk [15818]));
Q_ASSIGN U573 ( .B(clk), .A(\g.we_clk [15817]));
Q_ASSIGN U574 ( .B(clk), .A(\g.we_clk [15816]));
Q_ASSIGN U575 ( .B(clk), .A(\g.we_clk [15815]));
Q_ASSIGN U576 ( .B(clk), .A(\g.we_clk [15814]));
Q_ASSIGN U577 ( .B(clk), .A(\g.we_clk [15813]));
Q_ASSIGN U578 ( .B(clk), .A(\g.we_clk [15812]));
Q_ASSIGN U579 ( .B(clk), .A(\g.we_clk [15811]));
Q_ASSIGN U580 ( .B(clk), .A(\g.we_clk [15810]));
Q_ASSIGN U581 ( .B(clk), .A(\g.we_clk [15809]));
Q_ASSIGN U582 ( .B(clk), .A(\g.we_clk [15808]));
Q_ASSIGN U583 ( .B(clk), .A(\g.we_clk [15807]));
Q_ASSIGN U584 ( .B(clk), .A(\g.we_clk [15806]));
Q_ASSIGN U585 ( .B(clk), .A(\g.we_clk [15805]));
Q_ASSIGN U586 ( .B(clk), .A(\g.we_clk [15804]));
Q_ASSIGN U587 ( .B(clk), .A(\g.we_clk [15803]));
Q_ASSIGN U588 ( .B(clk), .A(\g.we_clk [15802]));
Q_ASSIGN U589 ( .B(clk), .A(\g.we_clk [15801]));
Q_ASSIGN U590 ( .B(clk), .A(\g.we_clk [15800]));
Q_ASSIGN U591 ( .B(clk), .A(\g.we_clk [15799]));
Q_ASSIGN U592 ( .B(clk), .A(\g.we_clk [15798]));
Q_ASSIGN U593 ( .B(clk), .A(\g.we_clk [15797]));
Q_ASSIGN U594 ( .B(clk), .A(\g.we_clk [15796]));
Q_ASSIGN U595 ( .B(clk), .A(\g.we_clk [15795]));
Q_ASSIGN U596 ( .B(clk), .A(\g.we_clk [15794]));
Q_ASSIGN U597 ( .B(clk), .A(\g.we_clk [15793]));
Q_ASSIGN U598 ( .B(clk), .A(\g.we_clk [15792]));
Q_ASSIGN U599 ( .B(clk), .A(\g.we_clk [15791]));
Q_ASSIGN U600 ( .B(clk), .A(\g.we_clk [15790]));
Q_ASSIGN U601 ( .B(clk), .A(\g.we_clk [15789]));
Q_ASSIGN U602 ( .B(clk), .A(\g.we_clk [15788]));
Q_ASSIGN U603 ( .B(clk), .A(\g.we_clk [15787]));
Q_ASSIGN U604 ( .B(clk), .A(\g.we_clk [15786]));
Q_ASSIGN U605 ( .B(clk), .A(\g.we_clk [15785]));
Q_ASSIGN U606 ( .B(clk), .A(\g.we_clk [15784]));
Q_ASSIGN U607 ( .B(clk), .A(\g.we_clk [15783]));
Q_ASSIGN U608 ( .B(clk), .A(\g.we_clk [15782]));
Q_ASSIGN U609 ( .B(clk), .A(\g.we_clk [15781]));
Q_ASSIGN U610 ( .B(clk), .A(\g.we_clk [15780]));
Q_ASSIGN U611 ( .B(clk), .A(\g.we_clk [15779]));
Q_ASSIGN U612 ( .B(clk), .A(\g.we_clk [15778]));
Q_ASSIGN U613 ( .B(clk), .A(\g.we_clk [15777]));
Q_ASSIGN U614 ( .B(clk), .A(\g.we_clk [15776]));
Q_ASSIGN U615 ( .B(clk), .A(\g.we_clk [15775]));
Q_ASSIGN U616 ( .B(clk), .A(\g.we_clk [15774]));
Q_ASSIGN U617 ( .B(clk), .A(\g.we_clk [15773]));
Q_ASSIGN U618 ( .B(clk), .A(\g.we_clk [15772]));
Q_ASSIGN U619 ( .B(clk), .A(\g.we_clk [15771]));
Q_ASSIGN U620 ( .B(clk), .A(\g.we_clk [15770]));
Q_ASSIGN U621 ( .B(clk), .A(\g.we_clk [15769]));
Q_ASSIGN U622 ( .B(clk), .A(\g.we_clk [15768]));
Q_ASSIGN U623 ( .B(clk), .A(\g.we_clk [15767]));
Q_ASSIGN U624 ( .B(clk), .A(\g.we_clk [15766]));
Q_ASSIGN U625 ( .B(clk), .A(\g.we_clk [15765]));
Q_ASSIGN U626 ( .B(clk), .A(\g.we_clk [15764]));
Q_ASSIGN U627 ( .B(clk), .A(\g.we_clk [15763]));
Q_ASSIGN U628 ( .B(clk), .A(\g.we_clk [15762]));
Q_ASSIGN U629 ( .B(clk), .A(\g.we_clk [15761]));
Q_ASSIGN U630 ( .B(clk), .A(\g.we_clk [15760]));
Q_ASSIGN U631 ( .B(clk), .A(\g.we_clk [15759]));
Q_ASSIGN U632 ( .B(clk), .A(\g.we_clk [15758]));
Q_ASSIGN U633 ( .B(clk), .A(\g.we_clk [15757]));
Q_ASSIGN U634 ( .B(clk), .A(\g.we_clk [15756]));
Q_ASSIGN U635 ( .B(clk), .A(\g.we_clk [15755]));
Q_ASSIGN U636 ( .B(clk), .A(\g.we_clk [15754]));
Q_ASSIGN U637 ( .B(clk), .A(\g.we_clk [15753]));
Q_ASSIGN U638 ( .B(clk), .A(\g.we_clk [15752]));
Q_ASSIGN U639 ( .B(clk), .A(\g.we_clk [15751]));
Q_ASSIGN U640 ( .B(clk), .A(\g.we_clk [15750]));
Q_ASSIGN U641 ( .B(clk), .A(\g.we_clk [15749]));
Q_ASSIGN U642 ( .B(clk), .A(\g.we_clk [15748]));
Q_ASSIGN U643 ( .B(clk), .A(\g.we_clk [15747]));
Q_ASSIGN U644 ( .B(clk), .A(\g.we_clk [15746]));
Q_ASSIGN U645 ( .B(clk), .A(\g.we_clk [15745]));
Q_ASSIGN U646 ( .B(clk), .A(\g.we_clk [15744]));
Q_ASSIGN U647 ( .B(clk), .A(\g.we_clk [15743]));
Q_ASSIGN U648 ( .B(clk), .A(\g.we_clk [15742]));
Q_ASSIGN U649 ( .B(clk), .A(\g.we_clk [15741]));
Q_ASSIGN U650 ( .B(clk), .A(\g.we_clk [15740]));
Q_ASSIGN U651 ( .B(clk), .A(\g.we_clk [15739]));
Q_ASSIGN U652 ( .B(clk), .A(\g.we_clk [15738]));
Q_ASSIGN U653 ( .B(clk), .A(\g.we_clk [15737]));
Q_ASSIGN U654 ( .B(clk), .A(\g.we_clk [15736]));
Q_ASSIGN U655 ( .B(clk), .A(\g.we_clk [15735]));
Q_ASSIGN U656 ( .B(clk), .A(\g.we_clk [15734]));
Q_ASSIGN U657 ( .B(clk), .A(\g.we_clk [15733]));
Q_ASSIGN U658 ( .B(clk), .A(\g.we_clk [15732]));
Q_ASSIGN U659 ( .B(clk), .A(\g.we_clk [15731]));
Q_ASSIGN U660 ( .B(clk), .A(\g.we_clk [15730]));
Q_ASSIGN U661 ( .B(clk), .A(\g.we_clk [15729]));
Q_ASSIGN U662 ( .B(clk), .A(\g.we_clk [15728]));
Q_ASSIGN U663 ( .B(clk), .A(\g.we_clk [15727]));
Q_ASSIGN U664 ( .B(clk), .A(\g.we_clk [15726]));
Q_ASSIGN U665 ( .B(clk), .A(\g.we_clk [15725]));
Q_ASSIGN U666 ( .B(clk), .A(\g.we_clk [15724]));
Q_ASSIGN U667 ( .B(clk), .A(\g.we_clk [15723]));
Q_ASSIGN U668 ( .B(clk), .A(\g.we_clk [15722]));
Q_ASSIGN U669 ( .B(clk), .A(\g.we_clk [15721]));
Q_ASSIGN U670 ( .B(clk), .A(\g.we_clk [15720]));
Q_ASSIGN U671 ( .B(clk), .A(\g.we_clk [15719]));
Q_ASSIGN U672 ( .B(clk), .A(\g.we_clk [15718]));
Q_ASSIGN U673 ( .B(clk), .A(\g.we_clk [15717]));
Q_ASSIGN U674 ( .B(clk), .A(\g.we_clk [15716]));
Q_ASSIGN U675 ( .B(clk), .A(\g.we_clk [15715]));
Q_ASSIGN U676 ( .B(clk), .A(\g.we_clk [15714]));
Q_ASSIGN U677 ( .B(clk), .A(\g.we_clk [15713]));
Q_ASSIGN U678 ( .B(clk), .A(\g.we_clk [15712]));
Q_ASSIGN U679 ( .B(clk), .A(\g.we_clk [15711]));
Q_ASSIGN U680 ( .B(clk), .A(\g.we_clk [15710]));
Q_ASSIGN U681 ( .B(clk), .A(\g.we_clk [15709]));
Q_ASSIGN U682 ( .B(clk), .A(\g.we_clk [15708]));
Q_ASSIGN U683 ( .B(clk), .A(\g.we_clk [15707]));
Q_ASSIGN U684 ( .B(clk), .A(\g.we_clk [15706]));
Q_ASSIGN U685 ( .B(clk), .A(\g.we_clk [15705]));
Q_ASSIGN U686 ( .B(clk), .A(\g.we_clk [15704]));
Q_ASSIGN U687 ( .B(clk), .A(\g.we_clk [15703]));
Q_ASSIGN U688 ( .B(clk), .A(\g.we_clk [15702]));
Q_ASSIGN U689 ( .B(clk), .A(\g.we_clk [15701]));
Q_ASSIGN U690 ( .B(clk), .A(\g.we_clk [15700]));
Q_ASSIGN U691 ( .B(clk), .A(\g.we_clk [15699]));
Q_ASSIGN U692 ( .B(clk), .A(\g.we_clk [15698]));
Q_ASSIGN U693 ( .B(clk), .A(\g.we_clk [15697]));
Q_ASSIGN U694 ( .B(clk), .A(\g.we_clk [15696]));
Q_ASSIGN U695 ( .B(clk), .A(\g.we_clk [15695]));
Q_ASSIGN U696 ( .B(clk), .A(\g.we_clk [15694]));
Q_ASSIGN U697 ( .B(clk), .A(\g.we_clk [15693]));
Q_ASSIGN U698 ( .B(clk), .A(\g.we_clk [15692]));
Q_ASSIGN U699 ( .B(clk), .A(\g.we_clk [15691]));
Q_ASSIGN U700 ( .B(clk), .A(\g.we_clk [15690]));
Q_ASSIGN U701 ( .B(clk), .A(\g.we_clk [15689]));
Q_ASSIGN U702 ( .B(clk), .A(\g.we_clk [15688]));
Q_ASSIGN U703 ( .B(clk), .A(\g.we_clk [15687]));
Q_ASSIGN U704 ( .B(clk), .A(\g.we_clk [15686]));
Q_ASSIGN U705 ( .B(clk), .A(\g.we_clk [15685]));
Q_ASSIGN U706 ( .B(clk), .A(\g.we_clk [15684]));
Q_ASSIGN U707 ( .B(clk), .A(\g.we_clk [15683]));
Q_ASSIGN U708 ( .B(clk), .A(\g.we_clk [15682]));
Q_ASSIGN U709 ( .B(clk), .A(\g.we_clk [15681]));
Q_ASSIGN U710 ( .B(clk), .A(\g.we_clk [15680]));
Q_ASSIGN U711 ( .B(clk), .A(\g.we_clk [15679]));
Q_ASSIGN U712 ( .B(clk), .A(\g.we_clk [15678]));
Q_ASSIGN U713 ( .B(clk), .A(\g.we_clk [15677]));
Q_ASSIGN U714 ( .B(clk), .A(\g.we_clk [15676]));
Q_ASSIGN U715 ( .B(clk), .A(\g.we_clk [15675]));
Q_ASSIGN U716 ( .B(clk), .A(\g.we_clk [15674]));
Q_ASSIGN U717 ( .B(clk), .A(\g.we_clk [15673]));
Q_ASSIGN U718 ( .B(clk), .A(\g.we_clk [15672]));
Q_ASSIGN U719 ( .B(clk), .A(\g.we_clk [15671]));
Q_ASSIGN U720 ( .B(clk), .A(\g.we_clk [15670]));
Q_ASSIGN U721 ( .B(clk), .A(\g.we_clk [15669]));
Q_ASSIGN U722 ( .B(clk), .A(\g.we_clk [15668]));
Q_ASSIGN U723 ( .B(clk), .A(\g.we_clk [15667]));
Q_ASSIGN U724 ( .B(clk), .A(\g.we_clk [15666]));
Q_ASSIGN U725 ( .B(clk), .A(\g.we_clk [15665]));
Q_ASSIGN U726 ( .B(clk), .A(\g.we_clk [15664]));
Q_ASSIGN U727 ( .B(clk), .A(\g.we_clk [15663]));
Q_ASSIGN U728 ( .B(clk), .A(\g.we_clk [15662]));
Q_ASSIGN U729 ( .B(clk), .A(\g.we_clk [15661]));
Q_ASSIGN U730 ( .B(clk), .A(\g.we_clk [15660]));
Q_ASSIGN U731 ( .B(clk), .A(\g.we_clk [15659]));
Q_ASSIGN U732 ( .B(clk), .A(\g.we_clk [15658]));
Q_ASSIGN U733 ( .B(clk), .A(\g.we_clk [15657]));
Q_ASSIGN U734 ( .B(clk), .A(\g.we_clk [15656]));
Q_ASSIGN U735 ( .B(clk), .A(\g.we_clk [15655]));
Q_ASSIGN U736 ( .B(clk), .A(\g.we_clk [15654]));
Q_ASSIGN U737 ( .B(clk), .A(\g.we_clk [15653]));
Q_ASSIGN U738 ( .B(clk), .A(\g.we_clk [15652]));
Q_ASSIGN U739 ( .B(clk), .A(\g.we_clk [15651]));
Q_ASSIGN U740 ( .B(clk), .A(\g.we_clk [15650]));
Q_ASSIGN U741 ( .B(clk), .A(\g.we_clk [15649]));
Q_ASSIGN U742 ( .B(clk), .A(\g.we_clk [15648]));
Q_ASSIGN U743 ( .B(clk), .A(\g.we_clk [15647]));
Q_ASSIGN U744 ( .B(clk), .A(\g.we_clk [15646]));
Q_ASSIGN U745 ( .B(clk), .A(\g.we_clk [15645]));
Q_ASSIGN U746 ( .B(clk), .A(\g.we_clk [15644]));
Q_ASSIGN U747 ( .B(clk), .A(\g.we_clk [15643]));
Q_ASSIGN U748 ( .B(clk), .A(\g.we_clk [15642]));
Q_ASSIGN U749 ( .B(clk), .A(\g.we_clk [15641]));
Q_ASSIGN U750 ( .B(clk), .A(\g.we_clk [15640]));
Q_ASSIGN U751 ( .B(clk), .A(\g.we_clk [15639]));
Q_ASSIGN U752 ( .B(clk), .A(\g.we_clk [15638]));
Q_ASSIGN U753 ( .B(clk), .A(\g.we_clk [15637]));
Q_ASSIGN U754 ( .B(clk), .A(\g.we_clk [15636]));
Q_ASSIGN U755 ( .B(clk), .A(\g.we_clk [15635]));
Q_ASSIGN U756 ( .B(clk), .A(\g.we_clk [15634]));
Q_ASSIGN U757 ( .B(clk), .A(\g.we_clk [15633]));
Q_ASSIGN U758 ( .B(clk), .A(\g.we_clk [15632]));
Q_ASSIGN U759 ( .B(clk), .A(\g.we_clk [15631]));
Q_ASSIGN U760 ( .B(clk), .A(\g.we_clk [15630]));
Q_ASSIGN U761 ( .B(clk), .A(\g.we_clk [15629]));
Q_ASSIGN U762 ( .B(clk), .A(\g.we_clk [15628]));
Q_ASSIGN U763 ( .B(clk), .A(\g.we_clk [15627]));
Q_ASSIGN U764 ( .B(clk), .A(\g.we_clk [15626]));
Q_ASSIGN U765 ( .B(clk), .A(\g.we_clk [15625]));
Q_ASSIGN U766 ( .B(clk), .A(\g.we_clk [15624]));
Q_ASSIGN U767 ( .B(clk), .A(\g.we_clk [15623]));
Q_ASSIGN U768 ( .B(clk), .A(\g.we_clk [15622]));
Q_ASSIGN U769 ( .B(clk), .A(\g.we_clk [15621]));
Q_ASSIGN U770 ( .B(clk), .A(\g.we_clk [15620]));
Q_ASSIGN U771 ( .B(clk), .A(\g.we_clk [15619]));
Q_ASSIGN U772 ( .B(clk), .A(\g.we_clk [15618]));
Q_ASSIGN U773 ( .B(clk), .A(\g.we_clk [15617]));
Q_ASSIGN U774 ( .B(clk), .A(\g.we_clk [15616]));
Q_ASSIGN U775 ( .B(clk), .A(\g.we_clk [15615]));
Q_ASSIGN U776 ( .B(clk), .A(\g.we_clk [15614]));
Q_ASSIGN U777 ( .B(clk), .A(\g.we_clk [15613]));
Q_ASSIGN U778 ( .B(clk), .A(\g.we_clk [15612]));
Q_ASSIGN U779 ( .B(clk), .A(\g.we_clk [15611]));
Q_ASSIGN U780 ( .B(clk), .A(\g.we_clk [15610]));
Q_ASSIGN U781 ( .B(clk), .A(\g.we_clk [15609]));
Q_ASSIGN U782 ( .B(clk), .A(\g.we_clk [15608]));
Q_ASSIGN U783 ( .B(clk), .A(\g.we_clk [15607]));
Q_ASSIGN U784 ( .B(clk), .A(\g.we_clk [15606]));
Q_ASSIGN U785 ( .B(clk), .A(\g.we_clk [15605]));
Q_ASSIGN U786 ( .B(clk), .A(\g.we_clk [15604]));
Q_ASSIGN U787 ( .B(clk), .A(\g.we_clk [15603]));
Q_ASSIGN U788 ( .B(clk), .A(\g.we_clk [15602]));
Q_ASSIGN U789 ( .B(clk), .A(\g.we_clk [15601]));
Q_ASSIGN U790 ( .B(clk), .A(\g.we_clk [15600]));
Q_ASSIGN U791 ( .B(clk), .A(\g.we_clk [15599]));
Q_ASSIGN U792 ( .B(clk), .A(\g.we_clk [15598]));
Q_ASSIGN U793 ( .B(clk), .A(\g.we_clk [15597]));
Q_ASSIGN U794 ( .B(clk), .A(\g.we_clk [15596]));
Q_ASSIGN U795 ( .B(clk), .A(\g.we_clk [15595]));
Q_ASSIGN U796 ( .B(clk), .A(\g.we_clk [15594]));
Q_ASSIGN U797 ( .B(clk), .A(\g.we_clk [15593]));
Q_ASSIGN U798 ( .B(clk), .A(\g.we_clk [15592]));
Q_ASSIGN U799 ( .B(clk), .A(\g.we_clk [15591]));
Q_ASSIGN U800 ( .B(clk), .A(\g.we_clk [15590]));
Q_ASSIGN U801 ( .B(clk), .A(\g.we_clk [15589]));
Q_ASSIGN U802 ( .B(clk), .A(\g.we_clk [15588]));
Q_ASSIGN U803 ( .B(clk), .A(\g.we_clk [15587]));
Q_ASSIGN U804 ( .B(clk), .A(\g.we_clk [15586]));
Q_ASSIGN U805 ( .B(clk), .A(\g.we_clk [15585]));
Q_ASSIGN U806 ( .B(clk), .A(\g.we_clk [15584]));
Q_ASSIGN U807 ( .B(clk), .A(\g.we_clk [15583]));
Q_ASSIGN U808 ( .B(clk), .A(\g.we_clk [15582]));
Q_ASSIGN U809 ( .B(clk), .A(\g.we_clk [15581]));
Q_ASSIGN U810 ( .B(clk), .A(\g.we_clk [15580]));
Q_ASSIGN U811 ( .B(clk), .A(\g.we_clk [15579]));
Q_ASSIGN U812 ( .B(clk), .A(\g.we_clk [15578]));
Q_ASSIGN U813 ( .B(clk), .A(\g.we_clk [15577]));
Q_ASSIGN U814 ( .B(clk), .A(\g.we_clk [15576]));
Q_ASSIGN U815 ( .B(clk), .A(\g.we_clk [15575]));
Q_ASSIGN U816 ( .B(clk), .A(\g.we_clk [15574]));
Q_ASSIGN U817 ( .B(clk), .A(\g.we_clk [15573]));
Q_ASSIGN U818 ( .B(clk), .A(\g.we_clk [15572]));
Q_ASSIGN U819 ( .B(clk), .A(\g.we_clk [15571]));
Q_ASSIGN U820 ( .B(clk), .A(\g.we_clk [15570]));
Q_ASSIGN U821 ( .B(clk), .A(\g.we_clk [15569]));
Q_ASSIGN U822 ( .B(clk), .A(\g.we_clk [15568]));
Q_ASSIGN U823 ( .B(clk), .A(\g.we_clk [15567]));
Q_ASSIGN U824 ( .B(clk), .A(\g.we_clk [15566]));
Q_ASSIGN U825 ( .B(clk), .A(\g.we_clk [15565]));
Q_ASSIGN U826 ( .B(clk), .A(\g.we_clk [15564]));
Q_ASSIGN U827 ( .B(clk), .A(\g.we_clk [15563]));
Q_ASSIGN U828 ( .B(clk), .A(\g.we_clk [15562]));
Q_ASSIGN U829 ( .B(clk), .A(\g.we_clk [15561]));
Q_ASSIGN U830 ( .B(clk), .A(\g.we_clk [15560]));
Q_ASSIGN U831 ( .B(clk), .A(\g.we_clk [15559]));
Q_ASSIGN U832 ( .B(clk), .A(\g.we_clk [15558]));
Q_ASSIGN U833 ( .B(clk), .A(\g.we_clk [15557]));
Q_ASSIGN U834 ( .B(clk), .A(\g.we_clk [15556]));
Q_ASSIGN U835 ( .B(clk), .A(\g.we_clk [15555]));
Q_ASSIGN U836 ( .B(clk), .A(\g.we_clk [15554]));
Q_ASSIGN U837 ( .B(clk), .A(\g.we_clk [15553]));
Q_ASSIGN U838 ( .B(clk), .A(\g.we_clk [15552]));
Q_ASSIGN U839 ( .B(clk), .A(\g.we_clk [15551]));
Q_ASSIGN U840 ( .B(clk), .A(\g.we_clk [15550]));
Q_ASSIGN U841 ( .B(clk), .A(\g.we_clk [15549]));
Q_ASSIGN U842 ( .B(clk), .A(\g.we_clk [15548]));
Q_ASSIGN U843 ( .B(clk), .A(\g.we_clk [15547]));
Q_ASSIGN U844 ( .B(clk), .A(\g.we_clk [15546]));
Q_ASSIGN U845 ( .B(clk), .A(\g.we_clk [15545]));
Q_ASSIGN U846 ( .B(clk), .A(\g.we_clk [15544]));
Q_ASSIGN U847 ( .B(clk), .A(\g.we_clk [15543]));
Q_ASSIGN U848 ( .B(clk), .A(\g.we_clk [15542]));
Q_ASSIGN U849 ( .B(clk), .A(\g.we_clk [15541]));
Q_ASSIGN U850 ( .B(clk), .A(\g.we_clk [15540]));
Q_ASSIGN U851 ( .B(clk), .A(\g.we_clk [15539]));
Q_ASSIGN U852 ( .B(clk), .A(\g.we_clk [15538]));
Q_ASSIGN U853 ( .B(clk), .A(\g.we_clk [15537]));
Q_ASSIGN U854 ( .B(clk), .A(\g.we_clk [15536]));
Q_ASSIGN U855 ( .B(clk), .A(\g.we_clk [15535]));
Q_ASSIGN U856 ( .B(clk), .A(\g.we_clk [15534]));
Q_ASSIGN U857 ( .B(clk), .A(\g.we_clk [15533]));
Q_ASSIGN U858 ( .B(clk), .A(\g.we_clk [15532]));
Q_ASSIGN U859 ( .B(clk), .A(\g.we_clk [15531]));
Q_ASSIGN U860 ( .B(clk), .A(\g.we_clk [15530]));
Q_ASSIGN U861 ( .B(clk), .A(\g.we_clk [15529]));
Q_ASSIGN U862 ( .B(clk), .A(\g.we_clk [15528]));
Q_ASSIGN U863 ( .B(clk), .A(\g.we_clk [15527]));
Q_ASSIGN U864 ( .B(clk), .A(\g.we_clk [15526]));
Q_ASSIGN U865 ( .B(clk), .A(\g.we_clk [15525]));
Q_ASSIGN U866 ( .B(clk), .A(\g.we_clk [15524]));
Q_ASSIGN U867 ( .B(clk), .A(\g.we_clk [15523]));
Q_ASSIGN U868 ( .B(clk), .A(\g.we_clk [15522]));
Q_ASSIGN U869 ( .B(clk), .A(\g.we_clk [15521]));
Q_ASSIGN U870 ( .B(clk), .A(\g.we_clk [15520]));
Q_ASSIGN U871 ( .B(clk), .A(\g.we_clk [15519]));
Q_ASSIGN U872 ( .B(clk), .A(\g.we_clk [15518]));
Q_ASSIGN U873 ( .B(clk), .A(\g.we_clk [15517]));
Q_ASSIGN U874 ( .B(clk), .A(\g.we_clk [15516]));
Q_ASSIGN U875 ( .B(clk), .A(\g.we_clk [15515]));
Q_ASSIGN U876 ( .B(clk), .A(\g.we_clk [15514]));
Q_ASSIGN U877 ( .B(clk), .A(\g.we_clk [15513]));
Q_ASSIGN U878 ( .B(clk), .A(\g.we_clk [15512]));
Q_ASSIGN U879 ( .B(clk), .A(\g.we_clk [15511]));
Q_ASSIGN U880 ( .B(clk), .A(\g.we_clk [15510]));
Q_ASSIGN U881 ( .B(clk), .A(\g.we_clk [15509]));
Q_ASSIGN U882 ( .B(clk), .A(\g.we_clk [15508]));
Q_ASSIGN U883 ( .B(clk), .A(\g.we_clk [15507]));
Q_ASSIGN U884 ( .B(clk), .A(\g.we_clk [15506]));
Q_ASSIGN U885 ( .B(clk), .A(\g.we_clk [15505]));
Q_ASSIGN U886 ( .B(clk), .A(\g.we_clk [15504]));
Q_ASSIGN U887 ( .B(clk), .A(\g.we_clk [15503]));
Q_ASSIGN U888 ( .B(clk), .A(\g.we_clk [15502]));
Q_ASSIGN U889 ( .B(clk), .A(\g.we_clk [15501]));
Q_ASSIGN U890 ( .B(clk), .A(\g.we_clk [15500]));
Q_ASSIGN U891 ( .B(clk), .A(\g.we_clk [15499]));
Q_ASSIGN U892 ( .B(clk), .A(\g.we_clk [15498]));
Q_ASSIGN U893 ( .B(clk), .A(\g.we_clk [15497]));
Q_ASSIGN U894 ( .B(clk), .A(\g.we_clk [15496]));
Q_ASSIGN U895 ( .B(clk), .A(\g.we_clk [15495]));
Q_ASSIGN U896 ( .B(clk), .A(\g.we_clk [15494]));
Q_ASSIGN U897 ( .B(clk), .A(\g.we_clk [15493]));
Q_ASSIGN U898 ( .B(clk), .A(\g.we_clk [15492]));
Q_ASSIGN U899 ( .B(clk), .A(\g.we_clk [15491]));
Q_ASSIGN U900 ( .B(clk), .A(\g.we_clk [15490]));
Q_ASSIGN U901 ( .B(clk), .A(\g.we_clk [15489]));
Q_ASSIGN U902 ( .B(clk), .A(\g.we_clk [15488]));
Q_ASSIGN U903 ( .B(clk), .A(\g.we_clk [15487]));
Q_ASSIGN U904 ( .B(clk), .A(\g.we_clk [15486]));
Q_ASSIGN U905 ( .B(clk), .A(\g.we_clk [15485]));
Q_ASSIGN U906 ( .B(clk), .A(\g.we_clk [15484]));
Q_ASSIGN U907 ( .B(clk), .A(\g.we_clk [15483]));
Q_ASSIGN U908 ( .B(clk), .A(\g.we_clk [15482]));
Q_ASSIGN U909 ( .B(clk), .A(\g.we_clk [15481]));
Q_ASSIGN U910 ( .B(clk), .A(\g.we_clk [15480]));
Q_ASSIGN U911 ( .B(clk), .A(\g.we_clk [15479]));
Q_ASSIGN U912 ( .B(clk), .A(\g.we_clk [15478]));
Q_ASSIGN U913 ( .B(clk), .A(\g.we_clk [15477]));
Q_ASSIGN U914 ( .B(clk), .A(\g.we_clk [15476]));
Q_ASSIGN U915 ( .B(clk), .A(\g.we_clk [15475]));
Q_ASSIGN U916 ( .B(clk), .A(\g.we_clk [15474]));
Q_ASSIGN U917 ( .B(clk), .A(\g.we_clk [15473]));
Q_ASSIGN U918 ( .B(clk), .A(\g.we_clk [15472]));
Q_ASSIGN U919 ( .B(clk), .A(\g.we_clk [15471]));
Q_ASSIGN U920 ( .B(clk), .A(\g.we_clk [15470]));
Q_ASSIGN U921 ( .B(clk), .A(\g.we_clk [15469]));
Q_ASSIGN U922 ( .B(clk), .A(\g.we_clk [15468]));
Q_ASSIGN U923 ( .B(clk), .A(\g.we_clk [15467]));
Q_ASSIGN U924 ( .B(clk), .A(\g.we_clk [15466]));
Q_ASSIGN U925 ( .B(clk), .A(\g.we_clk [15465]));
Q_ASSIGN U926 ( .B(clk), .A(\g.we_clk [15464]));
Q_ASSIGN U927 ( .B(clk), .A(\g.we_clk [15463]));
Q_ASSIGN U928 ( .B(clk), .A(\g.we_clk [15462]));
Q_ASSIGN U929 ( .B(clk), .A(\g.we_clk [15461]));
Q_ASSIGN U930 ( .B(clk), .A(\g.we_clk [15460]));
Q_ASSIGN U931 ( .B(clk), .A(\g.we_clk [15459]));
Q_ASSIGN U932 ( .B(clk), .A(\g.we_clk [15458]));
Q_ASSIGN U933 ( .B(clk), .A(\g.we_clk [15457]));
Q_ASSIGN U934 ( .B(clk), .A(\g.we_clk [15456]));
Q_ASSIGN U935 ( .B(clk), .A(\g.we_clk [15455]));
Q_ASSIGN U936 ( .B(clk), .A(\g.we_clk [15454]));
Q_ASSIGN U937 ( .B(clk), .A(\g.we_clk [15453]));
Q_ASSIGN U938 ( .B(clk), .A(\g.we_clk [15452]));
Q_ASSIGN U939 ( .B(clk), .A(\g.we_clk [15451]));
Q_ASSIGN U940 ( .B(clk), .A(\g.we_clk [15450]));
Q_ASSIGN U941 ( .B(clk), .A(\g.we_clk [15449]));
Q_ASSIGN U942 ( .B(clk), .A(\g.we_clk [15448]));
Q_ASSIGN U943 ( .B(clk), .A(\g.we_clk [15447]));
Q_ASSIGN U944 ( .B(clk), .A(\g.we_clk [15446]));
Q_ASSIGN U945 ( .B(clk), .A(\g.we_clk [15445]));
Q_ASSIGN U946 ( .B(clk), .A(\g.we_clk [15444]));
Q_ASSIGN U947 ( .B(clk), .A(\g.we_clk [15443]));
Q_ASSIGN U948 ( .B(clk), .A(\g.we_clk [15442]));
Q_ASSIGN U949 ( .B(clk), .A(\g.we_clk [15441]));
Q_ASSIGN U950 ( .B(clk), .A(\g.we_clk [15440]));
Q_ASSIGN U951 ( .B(clk), .A(\g.we_clk [15439]));
Q_ASSIGN U952 ( .B(clk), .A(\g.we_clk [15438]));
Q_ASSIGN U953 ( .B(clk), .A(\g.we_clk [15437]));
Q_ASSIGN U954 ( .B(clk), .A(\g.we_clk [15436]));
Q_ASSIGN U955 ( .B(clk), .A(\g.we_clk [15435]));
Q_ASSIGN U956 ( .B(clk), .A(\g.we_clk [15434]));
Q_ASSIGN U957 ( .B(clk), .A(\g.we_clk [15433]));
Q_ASSIGN U958 ( .B(clk), .A(\g.we_clk [15432]));
Q_ASSIGN U959 ( .B(clk), .A(\g.we_clk [15431]));
Q_ASSIGN U960 ( .B(clk), .A(\g.we_clk [15430]));
Q_ASSIGN U961 ( .B(clk), .A(\g.we_clk [15429]));
Q_ASSIGN U962 ( .B(clk), .A(\g.we_clk [15428]));
Q_ASSIGN U963 ( .B(clk), .A(\g.we_clk [15427]));
Q_ASSIGN U964 ( .B(clk), .A(\g.we_clk [15426]));
Q_ASSIGN U965 ( .B(clk), .A(\g.we_clk [15425]));
Q_ASSIGN U966 ( .B(clk), .A(\g.we_clk [15424]));
Q_ASSIGN U967 ( .B(clk), .A(\g.we_clk [15423]));
Q_ASSIGN U968 ( .B(clk), .A(\g.we_clk [15422]));
Q_ASSIGN U969 ( .B(clk), .A(\g.we_clk [15421]));
Q_ASSIGN U970 ( .B(clk), .A(\g.we_clk [15420]));
Q_ASSIGN U971 ( .B(clk), .A(\g.we_clk [15419]));
Q_ASSIGN U972 ( .B(clk), .A(\g.we_clk [15418]));
Q_ASSIGN U973 ( .B(clk), .A(\g.we_clk [15417]));
Q_ASSIGN U974 ( .B(clk), .A(\g.we_clk [15416]));
Q_ASSIGN U975 ( .B(clk), .A(\g.we_clk [15415]));
Q_ASSIGN U976 ( .B(clk), .A(\g.we_clk [15414]));
Q_ASSIGN U977 ( .B(clk), .A(\g.we_clk [15413]));
Q_ASSIGN U978 ( .B(clk), .A(\g.we_clk [15412]));
Q_ASSIGN U979 ( .B(clk), .A(\g.we_clk [15411]));
Q_ASSIGN U980 ( .B(clk), .A(\g.we_clk [15410]));
Q_ASSIGN U981 ( .B(clk), .A(\g.we_clk [15409]));
Q_ASSIGN U982 ( .B(clk), .A(\g.we_clk [15408]));
Q_ASSIGN U983 ( .B(clk), .A(\g.we_clk [15407]));
Q_ASSIGN U984 ( .B(clk), .A(\g.we_clk [15406]));
Q_ASSIGN U985 ( .B(clk), .A(\g.we_clk [15405]));
Q_ASSIGN U986 ( .B(clk), .A(\g.we_clk [15404]));
Q_ASSIGN U987 ( .B(clk), .A(\g.we_clk [15403]));
Q_ASSIGN U988 ( .B(clk), .A(\g.we_clk [15402]));
Q_ASSIGN U989 ( .B(clk), .A(\g.we_clk [15401]));
Q_ASSIGN U990 ( .B(clk), .A(\g.we_clk [15400]));
Q_ASSIGN U991 ( .B(clk), .A(\g.we_clk [15399]));
Q_ASSIGN U992 ( .B(clk), .A(\g.we_clk [15398]));
Q_ASSIGN U993 ( .B(clk), .A(\g.we_clk [15397]));
Q_ASSIGN U994 ( .B(clk), .A(\g.we_clk [15396]));
Q_ASSIGN U995 ( .B(clk), .A(\g.we_clk [15395]));
Q_ASSIGN U996 ( .B(clk), .A(\g.we_clk [15394]));
Q_ASSIGN U997 ( .B(clk), .A(\g.we_clk [15393]));
Q_ASSIGN U998 ( .B(clk), .A(\g.we_clk [15392]));
Q_ASSIGN U999 ( .B(clk), .A(\g.we_clk [15391]));
Q_ASSIGN U1000 ( .B(clk), .A(\g.we_clk [15390]));
Q_ASSIGN U1001 ( .B(clk), .A(\g.we_clk [15389]));
Q_ASSIGN U1002 ( .B(clk), .A(\g.we_clk [15388]));
Q_ASSIGN U1003 ( .B(clk), .A(\g.we_clk [15387]));
Q_ASSIGN U1004 ( .B(clk), .A(\g.we_clk [15386]));
Q_ASSIGN U1005 ( .B(clk), .A(\g.we_clk [15385]));
Q_ASSIGN U1006 ( .B(clk), .A(\g.we_clk [15384]));
Q_ASSIGN U1007 ( .B(clk), .A(\g.we_clk [15383]));
Q_ASSIGN U1008 ( .B(clk), .A(\g.we_clk [15382]));
Q_ASSIGN U1009 ( .B(clk), .A(\g.we_clk [15381]));
Q_ASSIGN U1010 ( .B(clk), .A(\g.we_clk [15380]));
Q_ASSIGN U1011 ( .B(clk), .A(\g.we_clk [15379]));
Q_ASSIGN U1012 ( .B(clk), .A(\g.we_clk [15378]));
Q_ASSIGN U1013 ( .B(clk), .A(\g.we_clk [15377]));
Q_ASSIGN U1014 ( .B(clk), .A(\g.we_clk [15376]));
Q_ASSIGN U1015 ( .B(clk), .A(\g.we_clk [15375]));
Q_ASSIGN U1016 ( .B(clk), .A(\g.we_clk [15374]));
Q_ASSIGN U1017 ( .B(clk), .A(\g.we_clk [15373]));
Q_ASSIGN U1018 ( .B(clk), .A(\g.we_clk [15372]));
Q_ASSIGN U1019 ( .B(clk), .A(\g.we_clk [15371]));
Q_ASSIGN U1020 ( .B(clk), .A(\g.we_clk [15370]));
Q_ASSIGN U1021 ( .B(clk), .A(\g.we_clk [15369]));
Q_ASSIGN U1022 ( .B(clk), .A(\g.we_clk [15368]));
Q_ASSIGN U1023 ( .B(clk), .A(\g.we_clk [15367]));
Q_ASSIGN U1024 ( .B(clk), .A(\g.we_clk [15366]));
Q_ASSIGN U1025 ( .B(clk), .A(\g.we_clk [15365]));
Q_ASSIGN U1026 ( .B(clk), .A(\g.we_clk [15364]));
Q_ASSIGN U1027 ( .B(clk), .A(\g.we_clk [15363]));
Q_ASSIGN U1028 ( .B(clk), .A(\g.we_clk [15362]));
Q_ASSIGN U1029 ( .B(clk), .A(\g.we_clk [15361]));
Q_ASSIGN U1030 ( .B(clk), .A(\g.we_clk [15360]));
Q_ASSIGN U1031 ( .B(clk), .A(\g.we_clk [15359]));
Q_ASSIGN U1032 ( .B(clk), .A(\g.we_clk [15358]));
Q_ASSIGN U1033 ( .B(clk), .A(\g.we_clk [15357]));
Q_ASSIGN U1034 ( .B(clk), .A(\g.we_clk [15356]));
Q_ASSIGN U1035 ( .B(clk), .A(\g.we_clk [15355]));
Q_ASSIGN U1036 ( .B(clk), .A(\g.we_clk [15354]));
Q_ASSIGN U1037 ( .B(clk), .A(\g.we_clk [15353]));
Q_ASSIGN U1038 ( .B(clk), .A(\g.we_clk [15352]));
Q_ASSIGN U1039 ( .B(clk), .A(\g.we_clk [15351]));
Q_ASSIGN U1040 ( .B(clk), .A(\g.we_clk [15350]));
Q_ASSIGN U1041 ( .B(clk), .A(\g.we_clk [15349]));
Q_ASSIGN U1042 ( .B(clk), .A(\g.we_clk [15348]));
Q_ASSIGN U1043 ( .B(clk), .A(\g.we_clk [15347]));
Q_ASSIGN U1044 ( .B(clk), .A(\g.we_clk [15346]));
Q_ASSIGN U1045 ( .B(clk), .A(\g.we_clk [15345]));
Q_ASSIGN U1046 ( .B(clk), .A(\g.we_clk [15344]));
Q_ASSIGN U1047 ( .B(clk), .A(\g.we_clk [15343]));
Q_ASSIGN U1048 ( .B(clk), .A(\g.we_clk [15342]));
Q_ASSIGN U1049 ( .B(clk), .A(\g.we_clk [15341]));
Q_ASSIGN U1050 ( .B(clk), .A(\g.we_clk [15340]));
Q_ASSIGN U1051 ( .B(clk), .A(\g.we_clk [15339]));
Q_ASSIGN U1052 ( .B(clk), .A(\g.we_clk [15338]));
Q_ASSIGN U1053 ( .B(clk), .A(\g.we_clk [15337]));
Q_ASSIGN U1054 ( .B(clk), .A(\g.we_clk [15336]));
Q_ASSIGN U1055 ( .B(clk), .A(\g.we_clk [15335]));
Q_ASSIGN U1056 ( .B(clk), .A(\g.we_clk [15334]));
Q_ASSIGN U1057 ( .B(clk), .A(\g.we_clk [15333]));
Q_ASSIGN U1058 ( .B(clk), .A(\g.we_clk [15332]));
Q_ASSIGN U1059 ( .B(clk), .A(\g.we_clk [15331]));
Q_ASSIGN U1060 ( .B(clk), .A(\g.we_clk [15330]));
Q_ASSIGN U1061 ( .B(clk), .A(\g.we_clk [15329]));
Q_ASSIGN U1062 ( .B(clk), .A(\g.we_clk [15328]));
Q_ASSIGN U1063 ( .B(clk), .A(\g.we_clk [15327]));
Q_ASSIGN U1064 ( .B(clk), .A(\g.we_clk [15326]));
Q_ASSIGN U1065 ( .B(clk), .A(\g.we_clk [15325]));
Q_ASSIGN U1066 ( .B(clk), .A(\g.we_clk [15324]));
Q_ASSIGN U1067 ( .B(clk), .A(\g.we_clk [15323]));
Q_ASSIGN U1068 ( .B(clk), .A(\g.we_clk [15322]));
Q_ASSIGN U1069 ( .B(clk), .A(\g.we_clk [15321]));
Q_ASSIGN U1070 ( .B(clk), .A(\g.we_clk [15320]));
Q_ASSIGN U1071 ( .B(clk), .A(\g.we_clk [15319]));
Q_ASSIGN U1072 ( .B(clk), .A(\g.we_clk [15318]));
Q_ASSIGN U1073 ( .B(clk), .A(\g.we_clk [15317]));
Q_ASSIGN U1074 ( .B(clk), .A(\g.we_clk [15316]));
Q_ASSIGN U1075 ( .B(clk), .A(\g.we_clk [15315]));
Q_ASSIGN U1076 ( .B(clk), .A(\g.we_clk [15314]));
Q_ASSIGN U1077 ( .B(clk), .A(\g.we_clk [15313]));
Q_ASSIGN U1078 ( .B(clk), .A(\g.we_clk [15312]));
Q_ASSIGN U1079 ( .B(clk), .A(\g.we_clk [15311]));
Q_ASSIGN U1080 ( .B(clk), .A(\g.we_clk [15310]));
Q_ASSIGN U1081 ( .B(clk), .A(\g.we_clk [15309]));
Q_ASSIGN U1082 ( .B(clk), .A(\g.we_clk [15308]));
Q_ASSIGN U1083 ( .B(clk), .A(\g.we_clk [15307]));
Q_ASSIGN U1084 ( .B(clk), .A(\g.we_clk [15306]));
Q_ASSIGN U1085 ( .B(clk), .A(\g.we_clk [15305]));
Q_ASSIGN U1086 ( .B(clk), .A(\g.we_clk [15304]));
Q_ASSIGN U1087 ( .B(clk), .A(\g.we_clk [15303]));
Q_ASSIGN U1088 ( .B(clk), .A(\g.we_clk [15302]));
Q_ASSIGN U1089 ( .B(clk), .A(\g.we_clk [15301]));
Q_ASSIGN U1090 ( .B(clk), .A(\g.we_clk [15300]));
Q_ASSIGN U1091 ( .B(clk), .A(\g.we_clk [15299]));
Q_ASSIGN U1092 ( .B(clk), .A(\g.we_clk [15298]));
Q_ASSIGN U1093 ( .B(clk), .A(\g.we_clk [15297]));
Q_ASSIGN U1094 ( .B(clk), .A(\g.we_clk [15296]));
Q_ASSIGN U1095 ( .B(clk), .A(\g.we_clk [15295]));
Q_ASSIGN U1096 ( .B(clk), .A(\g.we_clk [15294]));
Q_ASSIGN U1097 ( .B(clk), .A(\g.we_clk [15293]));
Q_ASSIGN U1098 ( .B(clk), .A(\g.we_clk [15292]));
Q_ASSIGN U1099 ( .B(clk), .A(\g.we_clk [15291]));
Q_ASSIGN U1100 ( .B(clk), .A(\g.we_clk [15290]));
Q_ASSIGN U1101 ( .B(clk), .A(\g.we_clk [15289]));
Q_ASSIGN U1102 ( .B(clk), .A(\g.we_clk [15288]));
Q_ASSIGN U1103 ( .B(clk), .A(\g.we_clk [15287]));
Q_ASSIGN U1104 ( .B(clk), .A(\g.we_clk [15286]));
Q_ASSIGN U1105 ( .B(clk), .A(\g.we_clk [15285]));
Q_ASSIGN U1106 ( .B(clk), .A(\g.we_clk [15284]));
Q_ASSIGN U1107 ( .B(clk), .A(\g.we_clk [15283]));
Q_ASSIGN U1108 ( .B(clk), .A(\g.we_clk [15282]));
Q_ASSIGN U1109 ( .B(clk), .A(\g.we_clk [15281]));
Q_ASSIGN U1110 ( .B(clk), .A(\g.we_clk [15280]));
Q_ASSIGN U1111 ( .B(clk), .A(\g.we_clk [15279]));
Q_ASSIGN U1112 ( .B(clk), .A(\g.we_clk [15278]));
Q_ASSIGN U1113 ( .B(clk), .A(\g.we_clk [15277]));
Q_ASSIGN U1114 ( .B(clk), .A(\g.we_clk [15276]));
Q_ASSIGN U1115 ( .B(clk), .A(\g.we_clk [15275]));
Q_ASSIGN U1116 ( .B(clk), .A(\g.we_clk [15274]));
Q_ASSIGN U1117 ( .B(clk), .A(\g.we_clk [15273]));
Q_ASSIGN U1118 ( .B(clk), .A(\g.we_clk [15272]));
Q_ASSIGN U1119 ( .B(clk), .A(\g.we_clk [15271]));
Q_ASSIGN U1120 ( .B(clk), .A(\g.we_clk [15270]));
Q_ASSIGN U1121 ( .B(clk), .A(\g.we_clk [15269]));
Q_ASSIGN U1122 ( .B(clk), .A(\g.we_clk [15268]));
Q_ASSIGN U1123 ( .B(clk), .A(\g.we_clk [15267]));
Q_ASSIGN U1124 ( .B(clk), .A(\g.we_clk [15266]));
Q_ASSIGN U1125 ( .B(clk), .A(\g.we_clk [15265]));
Q_ASSIGN U1126 ( .B(clk), .A(\g.we_clk [15264]));
Q_ASSIGN U1127 ( .B(clk), .A(\g.we_clk [15263]));
Q_ASSIGN U1128 ( .B(clk), .A(\g.we_clk [15262]));
Q_ASSIGN U1129 ( .B(clk), .A(\g.we_clk [15261]));
Q_ASSIGN U1130 ( .B(clk), .A(\g.we_clk [15260]));
Q_ASSIGN U1131 ( .B(clk), .A(\g.we_clk [15259]));
Q_ASSIGN U1132 ( .B(clk), .A(\g.we_clk [15258]));
Q_ASSIGN U1133 ( .B(clk), .A(\g.we_clk [15257]));
Q_ASSIGN U1134 ( .B(clk), .A(\g.we_clk [15256]));
Q_ASSIGN U1135 ( .B(clk), .A(\g.we_clk [15255]));
Q_ASSIGN U1136 ( .B(clk), .A(\g.we_clk [15254]));
Q_ASSIGN U1137 ( .B(clk), .A(\g.we_clk [15253]));
Q_ASSIGN U1138 ( .B(clk), .A(\g.we_clk [15252]));
Q_ASSIGN U1139 ( .B(clk), .A(\g.we_clk [15251]));
Q_ASSIGN U1140 ( .B(clk), .A(\g.we_clk [15250]));
Q_ASSIGN U1141 ( .B(clk), .A(\g.we_clk [15249]));
Q_ASSIGN U1142 ( .B(clk), .A(\g.we_clk [15248]));
Q_ASSIGN U1143 ( .B(clk), .A(\g.we_clk [15247]));
Q_ASSIGN U1144 ( .B(clk), .A(\g.we_clk [15246]));
Q_ASSIGN U1145 ( .B(clk), .A(\g.we_clk [15245]));
Q_ASSIGN U1146 ( .B(clk), .A(\g.we_clk [15244]));
Q_ASSIGN U1147 ( .B(clk), .A(\g.we_clk [15243]));
Q_ASSIGN U1148 ( .B(clk), .A(\g.we_clk [15242]));
Q_ASSIGN U1149 ( .B(clk), .A(\g.we_clk [15241]));
Q_ASSIGN U1150 ( .B(clk), .A(\g.we_clk [15240]));
Q_ASSIGN U1151 ( .B(clk), .A(\g.we_clk [15239]));
Q_ASSIGN U1152 ( .B(clk), .A(\g.we_clk [15238]));
Q_ASSIGN U1153 ( .B(clk), .A(\g.we_clk [15237]));
Q_ASSIGN U1154 ( .B(clk), .A(\g.we_clk [15236]));
Q_ASSIGN U1155 ( .B(clk), .A(\g.we_clk [15235]));
Q_ASSIGN U1156 ( .B(clk), .A(\g.we_clk [15234]));
Q_ASSIGN U1157 ( .B(clk), .A(\g.we_clk [15233]));
Q_ASSIGN U1158 ( .B(clk), .A(\g.we_clk [15232]));
Q_ASSIGN U1159 ( .B(clk), .A(\g.we_clk [15231]));
Q_ASSIGN U1160 ( .B(clk), .A(\g.we_clk [15230]));
Q_ASSIGN U1161 ( .B(clk), .A(\g.we_clk [15229]));
Q_ASSIGN U1162 ( .B(clk), .A(\g.we_clk [15228]));
Q_ASSIGN U1163 ( .B(clk), .A(\g.we_clk [15227]));
Q_ASSIGN U1164 ( .B(clk), .A(\g.we_clk [15226]));
Q_ASSIGN U1165 ( .B(clk), .A(\g.we_clk [15225]));
Q_ASSIGN U1166 ( .B(clk), .A(\g.we_clk [15224]));
Q_ASSIGN U1167 ( .B(clk), .A(\g.we_clk [15223]));
Q_ASSIGN U1168 ( .B(clk), .A(\g.we_clk [15222]));
Q_ASSIGN U1169 ( .B(clk), .A(\g.we_clk [15221]));
Q_ASSIGN U1170 ( .B(clk), .A(\g.we_clk [15220]));
Q_ASSIGN U1171 ( .B(clk), .A(\g.we_clk [15219]));
Q_ASSIGN U1172 ( .B(clk), .A(\g.we_clk [15218]));
Q_ASSIGN U1173 ( .B(clk), .A(\g.we_clk [15217]));
Q_ASSIGN U1174 ( .B(clk), .A(\g.we_clk [15216]));
Q_ASSIGN U1175 ( .B(clk), .A(\g.we_clk [15215]));
Q_ASSIGN U1176 ( .B(clk), .A(\g.we_clk [15214]));
Q_ASSIGN U1177 ( .B(clk), .A(\g.we_clk [15213]));
Q_ASSIGN U1178 ( .B(clk), .A(\g.we_clk [15212]));
Q_ASSIGN U1179 ( .B(clk), .A(\g.we_clk [15211]));
Q_ASSIGN U1180 ( .B(clk), .A(\g.we_clk [15210]));
Q_ASSIGN U1181 ( .B(clk), .A(\g.we_clk [15209]));
Q_ASSIGN U1182 ( .B(clk), .A(\g.we_clk [15208]));
Q_ASSIGN U1183 ( .B(clk), .A(\g.we_clk [15207]));
Q_ASSIGN U1184 ( .B(clk), .A(\g.we_clk [15206]));
Q_ASSIGN U1185 ( .B(clk), .A(\g.we_clk [15205]));
Q_ASSIGN U1186 ( .B(clk), .A(\g.we_clk [15204]));
Q_ASSIGN U1187 ( .B(clk), .A(\g.we_clk [15203]));
Q_ASSIGN U1188 ( .B(clk), .A(\g.we_clk [15202]));
Q_ASSIGN U1189 ( .B(clk), .A(\g.we_clk [15201]));
Q_ASSIGN U1190 ( .B(clk), .A(\g.we_clk [15200]));
Q_ASSIGN U1191 ( .B(clk), .A(\g.we_clk [15199]));
Q_ASSIGN U1192 ( .B(clk), .A(\g.we_clk [15198]));
Q_ASSIGN U1193 ( .B(clk), .A(\g.we_clk [15197]));
Q_ASSIGN U1194 ( .B(clk), .A(\g.we_clk [15196]));
Q_ASSIGN U1195 ( .B(clk), .A(\g.we_clk [15195]));
Q_ASSIGN U1196 ( .B(clk), .A(\g.we_clk [15194]));
Q_ASSIGN U1197 ( .B(clk), .A(\g.we_clk [15193]));
Q_ASSIGN U1198 ( .B(clk), .A(\g.we_clk [15192]));
Q_ASSIGN U1199 ( .B(clk), .A(\g.we_clk [15191]));
Q_ASSIGN U1200 ( .B(clk), .A(\g.we_clk [15190]));
Q_ASSIGN U1201 ( .B(clk), .A(\g.we_clk [15189]));
Q_ASSIGN U1202 ( .B(clk), .A(\g.we_clk [15188]));
Q_ASSIGN U1203 ( .B(clk), .A(\g.we_clk [15187]));
Q_ASSIGN U1204 ( .B(clk), .A(\g.we_clk [15186]));
Q_ASSIGN U1205 ( .B(clk), .A(\g.we_clk [15185]));
Q_ASSIGN U1206 ( .B(clk), .A(\g.we_clk [15184]));
Q_ASSIGN U1207 ( .B(clk), .A(\g.we_clk [15183]));
Q_ASSIGN U1208 ( .B(clk), .A(\g.we_clk [15182]));
Q_ASSIGN U1209 ( .B(clk), .A(\g.we_clk [15181]));
Q_ASSIGN U1210 ( .B(clk), .A(\g.we_clk [15180]));
Q_ASSIGN U1211 ( .B(clk), .A(\g.we_clk [15179]));
Q_ASSIGN U1212 ( .B(clk), .A(\g.we_clk [15178]));
Q_ASSIGN U1213 ( .B(clk), .A(\g.we_clk [15177]));
Q_ASSIGN U1214 ( .B(clk), .A(\g.we_clk [15176]));
Q_ASSIGN U1215 ( .B(clk), .A(\g.we_clk [15175]));
Q_ASSIGN U1216 ( .B(clk), .A(\g.we_clk [15174]));
Q_ASSIGN U1217 ( .B(clk), .A(\g.we_clk [15173]));
Q_ASSIGN U1218 ( .B(clk), .A(\g.we_clk [15172]));
Q_ASSIGN U1219 ( .B(clk), .A(\g.we_clk [15171]));
Q_ASSIGN U1220 ( .B(clk), .A(\g.we_clk [15170]));
Q_ASSIGN U1221 ( .B(clk), .A(\g.we_clk [15169]));
Q_ASSIGN U1222 ( .B(clk), .A(\g.we_clk [15168]));
Q_ASSIGN U1223 ( .B(clk), .A(\g.we_clk [15167]));
Q_ASSIGN U1224 ( .B(clk), .A(\g.we_clk [15166]));
Q_ASSIGN U1225 ( .B(clk), .A(\g.we_clk [15165]));
Q_ASSIGN U1226 ( .B(clk), .A(\g.we_clk [15164]));
Q_ASSIGN U1227 ( .B(clk), .A(\g.we_clk [15163]));
Q_ASSIGN U1228 ( .B(clk), .A(\g.we_clk [15162]));
Q_ASSIGN U1229 ( .B(clk), .A(\g.we_clk [15161]));
Q_ASSIGN U1230 ( .B(clk), .A(\g.we_clk [15160]));
Q_ASSIGN U1231 ( .B(clk), .A(\g.we_clk [15159]));
Q_ASSIGN U1232 ( .B(clk), .A(\g.we_clk [15158]));
Q_ASSIGN U1233 ( .B(clk), .A(\g.we_clk [15157]));
Q_ASSIGN U1234 ( .B(clk), .A(\g.we_clk [15156]));
Q_ASSIGN U1235 ( .B(clk), .A(\g.we_clk [15155]));
Q_ASSIGN U1236 ( .B(clk), .A(\g.we_clk [15154]));
Q_ASSIGN U1237 ( .B(clk), .A(\g.we_clk [15153]));
Q_ASSIGN U1238 ( .B(clk), .A(\g.we_clk [15152]));
Q_ASSIGN U1239 ( .B(clk), .A(\g.we_clk [15151]));
Q_ASSIGN U1240 ( .B(clk), .A(\g.we_clk [15150]));
Q_ASSIGN U1241 ( .B(clk), .A(\g.we_clk [15149]));
Q_ASSIGN U1242 ( .B(clk), .A(\g.we_clk [15148]));
Q_ASSIGN U1243 ( .B(clk), .A(\g.we_clk [15147]));
Q_ASSIGN U1244 ( .B(clk), .A(\g.we_clk [15146]));
Q_ASSIGN U1245 ( .B(clk), .A(\g.we_clk [15145]));
Q_ASSIGN U1246 ( .B(clk), .A(\g.we_clk [15144]));
Q_ASSIGN U1247 ( .B(clk), .A(\g.we_clk [15143]));
Q_ASSIGN U1248 ( .B(clk), .A(\g.we_clk [15142]));
Q_ASSIGN U1249 ( .B(clk), .A(\g.we_clk [15141]));
Q_ASSIGN U1250 ( .B(clk), .A(\g.we_clk [15140]));
Q_ASSIGN U1251 ( .B(clk), .A(\g.we_clk [15139]));
Q_ASSIGN U1252 ( .B(clk), .A(\g.we_clk [15138]));
Q_ASSIGN U1253 ( .B(clk), .A(\g.we_clk [15137]));
Q_ASSIGN U1254 ( .B(clk), .A(\g.we_clk [15136]));
Q_ASSIGN U1255 ( .B(clk), .A(\g.we_clk [15135]));
Q_ASSIGN U1256 ( .B(clk), .A(\g.we_clk [15134]));
Q_ASSIGN U1257 ( .B(clk), .A(\g.we_clk [15133]));
Q_ASSIGN U1258 ( .B(clk), .A(\g.we_clk [15132]));
Q_ASSIGN U1259 ( .B(clk), .A(\g.we_clk [15131]));
Q_ASSIGN U1260 ( .B(clk), .A(\g.we_clk [15130]));
Q_ASSIGN U1261 ( .B(clk), .A(\g.we_clk [15129]));
Q_ASSIGN U1262 ( .B(clk), .A(\g.we_clk [15128]));
Q_ASSIGN U1263 ( .B(clk), .A(\g.we_clk [15127]));
Q_ASSIGN U1264 ( .B(clk), .A(\g.we_clk [15126]));
Q_ASSIGN U1265 ( .B(clk), .A(\g.we_clk [15125]));
Q_ASSIGN U1266 ( .B(clk), .A(\g.we_clk [15124]));
Q_ASSIGN U1267 ( .B(clk), .A(\g.we_clk [15123]));
Q_ASSIGN U1268 ( .B(clk), .A(\g.we_clk [15122]));
Q_ASSIGN U1269 ( .B(clk), .A(\g.we_clk [15121]));
Q_ASSIGN U1270 ( .B(clk), .A(\g.we_clk [15120]));
Q_ASSIGN U1271 ( .B(clk), .A(\g.we_clk [15119]));
Q_ASSIGN U1272 ( .B(clk), .A(\g.we_clk [15118]));
Q_ASSIGN U1273 ( .B(clk), .A(\g.we_clk [15117]));
Q_ASSIGN U1274 ( .B(clk), .A(\g.we_clk [15116]));
Q_ASSIGN U1275 ( .B(clk), .A(\g.we_clk [15115]));
Q_ASSIGN U1276 ( .B(clk), .A(\g.we_clk [15114]));
Q_ASSIGN U1277 ( .B(clk), .A(\g.we_clk [15113]));
Q_ASSIGN U1278 ( .B(clk), .A(\g.we_clk [15112]));
Q_ASSIGN U1279 ( .B(clk), .A(\g.we_clk [15111]));
Q_ASSIGN U1280 ( .B(clk), .A(\g.we_clk [15110]));
Q_ASSIGN U1281 ( .B(clk), .A(\g.we_clk [15109]));
Q_ASSIGN U1282 ( .B(clk), .A(\g.we_clk [15108]));
Q_ASSIGN U1283 ( .B(clk), .A(\g.we_clk [15107]));
Q_ASSIGN U1284 ( .B(clk), .A(\g.we_clk [15106]));
Q_ASSIGN U1285 ( .B(clk), .A(\g.we_clk [15105]));
Q_ASSIGN U1286 ( .B(clk), .A(\g.we_clk [15104]));
Q_ASSIGN U1287 ( .B(clk), .A(\g.we_clk [15103]));
Q_ASSIGN U1288 ( .B(clk), .A(\g.we_clk [15102]));
Q_ASSIGN U1289 ( .B(clk), .A(\g.we_clk [15101]));
Q_ASSIGN U1290 ( .B(clk), .A(\g.we_clk [15100]));
Q_ASSIGN U1291 ( .B(clk), .A(\g.we_clk [15099]));
Q_ASSIGN U1292 ( .B(clk), .A(\g.we_clk [15098]));
Q_ASSIGN U1293 ( .B(clk), .A(\g.we_clk [15097]));
Q_ASSIGN U1294 ( .B(clk), .A(\g.we_clk [15096]));
Q_ASSIGN U1295 ( .B(clk), .A(\g.we_clk [15095]));
Q_ASSIGN U1296 ( .B(clk), .A(\g.we_clk [15094]));
Q_ASSIGN U1297 ( .B(clk), .A(\g.we_clk [15093]));
Q_ASSIGN U1298 ( .B(clk), .A(\g.we_clk [15092]));
Q_ASSIGN U1299 ( .B(clk), .A(\g.we_clk [15091]));
Q_ASSIGN U1300 ( .B(clk), .A(\g.we_clk [15090]));
Q_ASSIGN U1301 ( .B(clk), .A(\g.we_clk [15089]));
Q_ASSIGN U1302 ( .B(clk), .A(\g.we_clk [15088]));
Q_ASSIGN U1303 ( .B(clk), .A(\g.we_clk [15087]));
Q_ASSIGN U1304 ( .B(clk), .A(\g.we_clk [15086]));
Q_ASSIGN U1305 ( .B(clk), .A(\g.we_clk [15085]));
Q_ASSIGN U1306 ( .B(clk), .A(\g.we_clk [15084]));
Q_ASSIGN U1307 ( .B(clk), .A(\g.we_clk [15083]));
Q_ASSIGN U1308 ( .B(clk), .A(\g.we_clk [15082]));
Q_ASSIGN U1309 ( .B(clk), .A(\g.we_clk [15081]));
Q_ASSIGN U1310 ( .B(clk), .A(\g.we_clk [15080]));
Q_ASSIGN U1311 ( .B(clk), .A(\g.we_clk [15079]));
Q_ASSIGN U1312 ( .B(clk), .A(\g.we_clk [15078]));
Q_ASSIGN U1313 ( .B(clk), .A(\g.we_clk [15077]));
Q_ASSIGN U1314 ( .B(clk), .A(\g.we_clk [15076]));
Q_ASSIGN U1315 ( .B(clk), .A(\g.we_clk [15075]));
Q_ASSIGN U1316 ( .B(clk), .A(\g.we_clk [15074]));
Q_ASSIGN U1317 ( .B(clk), .A(\g.we_clk [15073]));
Q_ASSIGN U1318 ( .B(clk), .A(\g.we_clk [15072]));
Q_ASSIGN U1319 ( .B(clk), .A(\g.we_clk [15071]));
Q_ASSIGN U1320 ( .B(clk), .A(\g.we_clk [15070]));
Q_ASSIGN U1321 ( .B(clk), .A(\g.we_clk [15069]));
Q_ASSIGN U1322 ( .B(clk), .A(\g.we_clk [15068]));
Q_ASSIGN U1323 ( .B(clk), .A(\g.we_clk [15067]));
Q_ASSIGN U1324 ( .B(clk), .A(\g.we_clk [15066]));
Q_ASSIGN U1325 ( .B(clk), .A(\g.we_clk [15065]));
Q_ASSIGN U1326 ( .B(clk), .A(\g.we_clk [15064]));
Q_ASSIGN U1327 ( .B(clk), .A(\g.we_clk [15063]));
Q_ASSIGN U1328 ( .B(clk), .A(\g.we_clk [15062]));
Q_ASSIGN U1329 ( .B(clk), .A(\g.we_clk [15061]));
Q_ASSIGN U1330 ( .B(clk), .A(\g.we_clk [15060]));
Q_ASSIGN U1331 ( .B(clk), .A(\g.we_clk [15059]));
Q_ASSIGN U1332 ( .B(clk), .A(\g.we_clk [15058]));
Q_ASSIGN U1333 ( .B(clk), .A(\g.we_clk [15057]));
Q_ASSIGN U1334 ( .B(clk), .A(\g.we_clk [15056]));
Q_ASSIGN U1335 ( .B(clk), .A(\g.we_clk [15055]));
Q_ASSIGN U1336 ( .B(clk), .A(\g.we_clk [15054]));
Q_ASSIGN U1337 ( .B(clk), .A(\g.we_clk [15053]));
Q_ASSIGN U1338 ( .B(clk), .A(\g.we_clk [15052]));
Q_ASSIGN U1339 ( .B(clk), .A(\g.we_clk [15051]));
Q_ASSIGN U1340 ( .B(clk), .A(\g.we_clk [15050]));
Q_ASSIGN U1341 ( .B(clk), .A(\g.we_clk [15049]));
Q_ASSIGN U1342 ( .B(clk), .A(\g.we_clk [15048]));
Q_ASSIGN U1343 ( .B(clk), .A(\g.we_clk [15047]));
Q_ASSIGN U1344 ( .B(clk), .A(\g.we_clk [15046]));
Q_ASSIGN U1345 ( .B(clk), .A(\g.we_clk [15045]));
Q_ASSIGN U1346 ( .B(clk), .A(\g.we_clk [15044]));
Q_ASSIGN U1347 ( .B(clk), .A(\g.we_clk [15043]));
Q_ASSIGN U1348 ( .B(clk), .A(\g.we_clk [15042]));
Q_ASSIGN U1349 ( .B(clk), .A(\g.we_clk [15041]));
Q_ASSIGN U1350 ( .B(clk), .A(\g.we_clk [15040]));
Q_ASSIGN U1351 ( .B(clk), .A(\g.we_clk [15039]));
Q_ASSIGN U1352 ( .B(clk), .A(\g.we_clk [15038]));
Q_ASSIGN U1353 ( .B(clk), .A(\g.we_clk [15037]));
Q_ASSIGN U1354 ( .B(clk), .A(\g.we_clk [15036]));
Q_ASSIGN U1355 ( .B(clk), .A(\g.we_clk [15035]));
Q_ASSIGN U1356 ( .B(clk), .A(\g.we_clk [15034]));
Q_ASSIGN U1357 ( .B(clk), .A(\g.we_clk [15033]));
Q_ASSIGN U1358 ( .B(clk), .A(\g.we_clk [15032]));
Q_ASSIGN U1359 ( .B(clk), .A(\g.we_clk [15031]));
Q_ASSIGN U1360 ( .B(clk), .A(\g.we_clk [15030]));
Q_ASSIGN U1361 ( .B(clk), .A(\g.we_clk [15029]));
Q_ASSIGN U1362 ( .B(clk), .A(\g.we_clk [15028]));
Q_ASSIGN U1363 ( .B(clk), .A(\g.we_clk [15027]));
Q_ASSIGN U1364 ( .B(clk), .A(\g.we_clk [15026]));
Q_ASSIGN U1365 ( .B(clk), .A(\g.we_clk [15025]));
Q_ASSIGN U1366 ( .B(clk), .A(\g.we_clk [15024]));
Q_ASSIGN U1367 ( .B(clk), .A(\g.we_clk [15023]));
Q_ASSIGN U1368 ( .B(clk), .A(\g.we_clk [15022]));
Q_ASSIGN U1369 ( .B(clk), .A(\g.we_clk [15021]));
Q_ASSIGN U1370 ( .B(clk), .A(\g.we_clk [15020]));
Q_ASSIGN U1371 ( .B(clk), .A(\g.we_clk [15019]));
Q_ASSIGN U1372 ( .B(clk), .A(\g.we_clk [15018]));
Q_ASSIGN U1373 ( .B(clk), .A(\g.we_clk [15017]));
Q_ASSIGN U1374 ( .B(clk), .A(\g.we_clk [15016]));
Q_ASSIGN U1375 ( .B(clk), .A(\g.we_clk [15015]));
Q_ASSIGN U1376 ( .B(clk), .A(\g.we_clk [15014]));
Q_ASSIGN U1377 ( .B(clk), .A(\g.we_clk [15013]));
Q_ASSIGN U1378 ( .B(clk), .A(\g.we_clk [15012]));
Q_ASSIGN U1379 ( .B(clk), .A(\g.we_clk [15011]));
Q_ASSIGN U1380 ( .B(clk), .A(\g.we_clk [15010]));
Q_ASSIGN U1381 ( .B(clk), .A(\g.we_clk [15009]));
Q_ASSIGN U1382 ( .B(clk), .A(\g.we_clk [15008]));
Q_ASSIGN U1383 ( .B(clk), .A(\g.we_clk [15007]));
Q_ASSIGN U1384 ( .B(clk), .A(\g.we_clk [15006]));
Q_ASSIGN U1385 ( .B(clk), .A(\g.we_clk [15005]));
Q_ASSIGN U1386 ( .B(clk), .A(\g.we_clk [15004]));
Q_ASSIGN U1387 ( .B(clk), .A(\g.we_clk [15003]));
Q_ASSIGN U1388 ( .B(clk), .A(\g.we_clk [15002]));
Q_ASSIGN U1389 ( .B(clk), .A(\g.we_clk [15001]));
Q_ASSIGN U1390 ( .B(clk), .A(\g.we_clk [15000]));
Q_ASSIGN U1391 ( .B(clk), .A(\g.we_clk [14999]));
Q_ASSIGN U1392 ( .B(clk), .A(\g.we_clk [14998]));
Q_ASSIGN U1393 ( .B(clk), .A(\g.we_clk [14997]));
Q_ASSIGN U1394 ( .B(clk), .A(\g.we_clk [14996]));
Q_ASSIGN U1395 ( .B(clk), .A(\g.we_clk [14995]));
Q_ASSIGN U1396 ( .B(clk), .A(\g.we_clk [14994]));
Q_ASSIGN U1397 ( .B(clk), .A(\g.we_clk [14993]));
Q_ASSIGN U1398 ( .B(clk), .A(\g.we_clk [14992]));
Q_ASSIGN U1399 ( .B(clk), .A(\g.we_clk [14991]));
Q_ASSIGN U1400 ( .B(clk), .A(\g.we_clk [14990]));
Q_ASSIGN U1401 ( .B(clk), .A(\g.we_clk [14989]));
Q_ASSIGN U1402 ( .B(clk), .A(\g.we_clk [14988]));
Q_ASSIGN U1403 ( .B(clk), .A(\g.we_clk [14987]));
Q_ASSIGN U1404 ( .B(clk), .A(\g.we_clk [14986]));
Q_ASSIGN U1405 ( .B(clk), .A(\g.we_clk [14985]));
Q_ASSIGN U1406 ( .B(clk), .A(\g.we_clk [14984]));
Q_ASSIGN U1407 ( .B(clk), .A(\g.we_clk [14983]));
Q_ASSIGN U1408 ( .B(clk), .A(\g.we_clk [14982]));
Q_ASSIGN U1409 ( .B(clk), .A(\g.we_clk [14981]));
Q_ASSIGN U1410 ( .B(clk), .A(\g.we_clk [14980]));
Q_ASSIGN U1411 ( .B(clk), .A(\g.we_clk [14979]));
Q_ASSIGN U1412 ( .B(clk), .A(\g.we_clk [14978]));
Q_ASSIGN U1413 ( .B(clk), .A(\g.we_clk [14977]));
Q_ASSIGN U1414 ( .B(clk), .A(\g.we_clk [14976]));
Q_ASSIGN U1415 ( .B(clk), .A(\g.we_clk [14975]));
Q_ASSIGN U1416 ( .B(clk), .A(\g.we_clk [14974]));
Q_ASSIGN U1417 ( .B(clk), .A(\g.we_clk [14973]));
Q_ASSIGN U1418 ( .B(clk), .A(\g.we_clk [14972]));
Q_ASSIGN U1419 ( .B(clk), .A(\g.we_clk [14971]));
Q_ASSIGN U1420 ( .B(clk), .A(\g.we_clk [14970]));
Q_ASSIGN U1421 ( .B(clk), .A(\g.we_clk [14969]));
Q_ASSIGN U1422 ( .B(clk), .A(\g.we_clk [14968]));
Q_ASSIGN U1423 ( .B(clk), .A(\g.we_clk [14967]));
Q_ASSIGN U1424 ( .B(clk), .A(\g.we_clk [14966]));
Q_ASSIGN U1425 ( .B(clk), .A(\g.we_clk [14965]));
Q_ASSIGN U1426 ( .B(clk), .A(\g.we_clk [14964]));
Q_ASSIGN U1427 ( .B(clk), .A(\g.we_clk [14963]));
Q_ASSIGN U1428 ( .B(clk), .A(\g.we_clk [14962]));
Q_ASSIGN U1429 ( .B(clk), .A(\g.we_clk [14961]));
Q_ASSIGN U1430 ( .B(clk), .A(\g.we_clk [14960]));
Q_ASSIGN U1431 ( .B(clk), .A(\g.we_clk [14959]));
Q_ASSIGN U1432 ( .B(clk), .A(\g.we_clk [14958]));
Q_ASSIGN U1433 ( .B(clk), .A(\g.we_clk [14957]));
Q_ASSIGN U1434 ( .B(clk), .A(\g.we_clk [14956]));
Q_ASSIGN U1435 ( .B(clk), .A(\g.we_clk [14955]));
Q_ASSIGN U1436 ( .B(clk), .A(\g.we_clk [14954]));
Q_ASSIGN U1437 ( .B(clk), .A(\g.we_clk [14953]));
Q_ASSIGN U1438 ( .B(clk), .A(\g.we_clk [14952]));
Q_ASSIGN U1439 ( .B(clk), .A(\g.we_clk [14951]));
Q_ASSIGN U1440 ( .B(clk), .A(\g.we_clk [14950]));
Q_ASSIGN U1441 ( .B(clk), .A(\g.we_clk [14949]));
Q_ASSIGN U1442 ( .B(clk), .A(\g.we_clk [14948]));
Q_ASSIGN U1443 ( .B(clk), .A(\g.we_clk [14947]));
Q_ASSIGN U1444 ( .B(clk), .A(\g.we_clk [14946]));
Q_ASSIGN U1445 ( .B(clk), .A(\g.we_clk [14945]));
Q_ASSIGN U1446 ( .B(clk), .A(\g.we_clk [14944]));
Q_ASSIGN U1447 ( .B(clk), .A(\g.we_clk [14943]));
Q_ASSIGN U1448 ( .B(clk), .A(\g.we_clk [14942]));
Q_ASSIGN U1449 ( .B(clk), .A(\g.we_clk [14941]));
Q_ASSIGN U1450 ( .B(clk), .A(\g.we_clk [14940]));
Q_ASSIGN U1451 ( .B(clk), .A(\g.we_clk [14939]));
Q_ASSIGN U1452 ( .B(clk), .A(\g.we_clk [14938]));
Q_ASSIGN U1453 ( .B(clk), .A(\g.we_clk [14937]));
Q_ASSIGN U1454 ( .B(clk), .A(\g.we_clk [14936]));
Q_ASSIGN U1455 ( .B(clk), .A(\g.we_clk [14935]));
Q_ASSIGN U1456 ( .B(clk), .A(\g.we_clk [14934]));
Q_ASSIGN U1457 ( .B(clk), .A(\g.we_clk [14933]));
Q_ASSIGN U1458 ( .B(clk), .A(\g.we_clk [14932]));
Q_ASSIGN U1459 ( .B(clk), .A(\g.we_clk [14931]));
Q_ASSIGN U1460 ( .B(clk), .A(\g.we_clk [14930]));
Q_ASSIGN U1461 ( .B(clk), .A(\g.we_clk [14929]));
Q_ASSIGN U1462 ( .B(clk), .A(\g.we_clk [14928]));
Q_ASSIGN U1463 ( .B(clk), .A(\g.we_clk [14927]));
Q_ASSIGN U1464 ( .B(clk), .A(\g.we_clk [14926]));
Q_ASSIGN U1465 ( .B(clk), .A(\g.we_clk [14925]));
Q_ASSIGN U1466 ( .B(clk), .A(\g.we_clk [14924]));
Q_ASSIGN U1467 ( .B(clk), .A(\g.we_clk [14923]));
Q_ASSIGN U1468 ( .B(clk), .A(\g.we_clk [14922]));
Q_ASSIGN U1469 ( .B(clk), .A(\g.we_clk [14921]));
Q_ASSIGN U1470 ( .B(clk), .A(\g.we_clk [14920]));
Q_ASSIGN U1471 ( .B(clk), .A(\g.we_clk [14919]));
Q_ASSIGN U1472 ( .B(clk), .A(\g.we_clk [14918]));
Q_ASSIGN U1473 ( .B(clk), .A(\g.we_clk [14917]));
Q_ASSIGN U1474 ( .B(clk), .A(\g.we_clk [14916]));
Q_ASSIGN U1475 ( .B(clk), .A(\g.we_clk [14915]));
Q_ASSIGN U1476 ( .B(clk), .A(\g.we_clk [14914]));
Q_ASSIGN U1477 ( .B(clk), .A(\g.we_clk [14913]));
Q_ASSIGN U1478 ( .B(clk), .A(\g.we_clk [14912]));
Q_ASSIGN U1479 ( .B(clk), .A(\g.we_clk [14911]));
Q_ASSIGN U1480 ( .B(clk), .A(\g.we_clk [14910]));
Q_ASSIGN U1481 ( .B(clk), .A(\g.we_clk [14909]));
Q_ASSIGN U1482 ( .B(clk), .A(\g.we_clk [14908]));
Q_ASSIGN U1483 ( .B(clk), .A(\g.we_clk [14907]));
Q_ASSIGN U1484 ( .B(clk), .A(\g.we_clk [14906]));
Q_ASSIGN U1485 ( .B(clk), .A(\g.we_clk [14905]));
Q_ASSIGN U1486 ( .B(clk), .A(\g.we_clk [14904]));
Q_ASSIGN U1487 ( .B(clk), .A(\g.we_clk [14903]));
Q_ASSIGN U1488 ( .B(clk), .A(\g.we_clk [14902]));
Q_ASSIGN U1489 ( .B(clk), .A(\g.we_clk [14901]));
Q_ASSIGN U1490 ( .B(clk), .A(\g.we_clk [14900]));
Q_ASSIGN U1491 ( .B(clk), .A(\g.we_clk [14899]));
Q_ASSIGN U1492 ( .B(clk), .A(\g.we_clk [14898]));
Q_ASSIGN U1493 ( .B(clk), .A(\g.we_clk [14897]));
Q_ASSIGN U1494 ( .B(clk), .A(\g.we_clk [14896]));
Q_ASSIGN U1495 ( .B(clk), .A(\g.we_clk [14895]));
Q_ASSIGN U1496 ( .B(clk), .A(\g.we_clk [14894]));
Q_ASSIGN U1497 ( .B(clk), .A(\g.we_clk [14893]));
Q_ASSIGN U1498 ( .B(clk), .A(\g.we_clk [14892]));
Q_ASSIGN U1499 ( .B(clk), .A(\g.we_clk [14891]));
Q_ASSIGN U1500 ( .B(clk), .A(\g.we_clk [14890]));
Q_ASSIGN U1501 ( .B(clk), .A(\g.we_clk [14889]));
Q_ASSIGN U1502 ( .B(clk), .A(\g.we_clk [14888]));
Q_ASSIGN U1503 ( .B(clk), .A(\g.we_clk [14887]));
Q_ASSIGN U1504 ( .B(clk), .A(\g.we_clk [14886]));
Q_ASSIGN U1505 ( .B(clk), .A(\g.we_clk [14885]));
Q_ASSIGN U1506 ( .B(clk), .A(\g.we_clk [14884]));
Q_ASSIGN U1507 ( .B(clk), .A(\g.we_clk [14883]));
Q_ASSIGN U1508 ( .B(clk), .A(\g.we_clk [14882]));
Q_ASSIGN U1509 ( .B(clk), .A(\g.we_clk [14881]));
Q_ASSIGN U1510 ( .B(clk), .A(\g.we_clk [14880]));
Q_ASSIGN U1511 ( .B(clk), .A(\g.we_clk [14879]));
Q_ASSIGN U1512 ( .B(clk), .A(\g.we_clk [14878]));
Q_ASSIGN U1513 ( .B(clk), .A(\g.we_clk [14877]));
Q_ASSIGN U1514 ( .B(clk), .A(\g.we_clk [14876]));
Q_ASSIGN U1515 ( .B(clk), .A(\g.we_clk [14875]));
Q_ASSIGN U1516 ( .B(clk), .A(\g.we_clk [14874]));
Q_ASSIGN U1517 ( .B(clk), .A(\g.we_clk [14873]));
Q_ASSIGN U1518 ( .B(clk), .A(\g.we_clk [14872]));
Q_ASSIGN U1519 ( .B(clk), .A(\g.we_clk [14871]));
Q_ASSIGN U1520 ( .B(clk), .A(\g.we_clk [14870]));
Q_ASSIGN U1521 ( .B(clk), .A(\g.we_clk [14869]));
Q_ASSIGN U1522 ( .B(clk), .A(\g.we_clk [14868]));
Q_ASSIGN U1523 ( .B(clk), .A(\g.we_clk [14867]));
Q_ASSIGN U1524 ( .B(clk), .A(\g.we_clk [14866]));
Q_ASSIGN U1525 ( .B(clk), .A(\g.we_clk [14865]));
Q_ASSIGN U1526 ( .B(clk), .A(\g.we_clk [14864]));
Q_ASSIGN U1527 ( .B(clk), .A(\g.we_clk [14863]));
Q_ASSIGN U1528 ( .B(clk), .A(\g.we_clk [14862]));
Q_ASSIGN U1529 ( .B(clk), .A(\g.we_clk [14861]));
Q_ASSIGN U1530 ( .B(clk), .A(\g.we_clk [14860]));
Q_ASSIGN U1531 ( .B(clk), .A(\g.we_clk [14859]));
Q_ASSIGN U1532 ( .B(clk), .A(\g.we_clk [14858]));
Q_ASSIGN U1533 ( .B(clk), .A(\g.we_clk [14857]));
Q_ASSIGN U1534 ( .B(clk), .A(\g.we_clk [14856]));
Q_ASSIGN U1535 ( .B(clk), .A(\g.we_clk [14855]));
Q_ASSIGN U1536 ( .B(clk), .A(\g.we_clk [14854]));
Q_ASSIGN U1537 ( .B(clk), .A(\g.we_clk [14853]));
Q_ASSIGN U1538 ( .B(clk), .A(\g.we_clk [14852]));
Q_ASSIGN U1539 ( .B(clk), .A(\g.we_clk [14851]));
Q_ASSIGN U1540 ( .B(clk), .A(\g.we_clk [14850]));
Q_ASSIGN U1541 ( .B(clk), .A(\g.we_clk [14849]));
Q_ASSIGN U1542 ( .B(clk), .A(\g.we_clk [14848]));
Q_ASSIGN U1543 ( .B(clk), .A(\g.we_clk [14847]));
Q_ASSIGN U1544 ( .B(clk), .A(\g.we_clk [14846]));
Q_ASSIGN U1545 ( .B(clk), .A(\g.we_clk [14845]));
Q_ASSIGN U1546 ( .B(clk), .A(\g.we_clk [14844]));
Q_ASSIGN U1547 ( .B(clk), .A(\g.we_clk [14843]));
Q_ASSIGN U1548 ( .B(clk), .A(\g.we_clk [14842]));
Q_ASSIGN U1549 ( .B(clk), .A(\g.we_clk [14841]));
Q_ASSIGN U1550 ( .B(clk), .A(\g.we_clk [14840]));
Q_ASSIGN U1551 ( .B(clk), .A(\g.we_clk [14839]));
Q_ASSIGN U1552 ( .B(clk), .A(\g.we_clk [14838]));
Q_ASSIGN U1553 ( .B(clk), .A(\g.we_clk [14837]));
Q_ASSIGN U1554 ( .B(clk), .A(\g.we_clk [14836]));
Q_ASSIGN U1555 ( .B(clk), .A(\g.we_clk [14835]));
Q_ASSIGN U1556 ( .B(clk), .A(\g.we_clk [14834]));
Q_ASSIGN U1557 ( .B(clk), .A(\g.we_clk [14833]));
Q_ASSIGN U1558 ( .B(clk), .A(\g.we_clk [14832]));
Q_ASSIGN U1559 ( .B(clk), .A(\g.we_clk [14831]));
Q_ASSIGN U1560 ( .B(clk), .A(\g.we_clk [14830]));
Q_ASSIGN U1561 ( .B(clk), .A(\g.we_clk [14829]));
Q_ASSIGN U1562 ( .B(clk), .A(\g.we_clk [14828]));
Q_ASSIGN U1563 ( .B(clk), .A(\g.we_clk [14827]));
Q_ASSIGN U1564 ( .B(clk), .A(\g.we_clk [14826]));
Q_ASSIGN U1565 ( .B(clk), .A(\g.we_clk [14825]));
Q_ASSIGN U1566 ( .B(clk), .A(\g.we_clk [14824]));
Q_ASSIGN U1567 ( .B(clk), .A(\g.we_clk [14823]));
Q_ASSIGN U1568 ( .B(clk), .A(\g.we_clk [14822]));
Q_ASSIGN U1569 ( .B(clk), .A(\g.we_clk [14821]));
Q_ASSIGN U1570 ( .B(clk), .A(\g.we_clk [14820]));
Q_ASSIGN U1571 ( .B(clk), .A(\g.we_clk [14819]));
Q_ASSIGN U1572 ( .B(clk), .A(\g.we_clk [14818]));
Q_ASSIGN U1573 ( .B(clk), .A(\g.we_clk [14817]));
Q_ASSIGN U1574 ( .B(clk), .A(\g.we_clk [14816]));
Q_ASSIGN U1575 ( .B(clk), .A(\g.we_clk [14815]));
Q_ASSIGN U1576 ( .B(clk), .A(\g.we_clk [14814]));
Q_ASSIGN U1577 ( .B(clk), .A(\g.we_clk [14813]));
Q_ASSIGN U1578 ( .B(clk), .A(\g.we_clk [14812]));
Q_ASSIGN U1579 ( .B(clk), .A(\g.we_clk [14811]));
Q_ASSIGN U1580 ( .B(clk), .A(\g.we_clk [14810]));
Q_ASSIGN U1581 ( .B(clk), .A(\g.we_clk [14809]));
Q_ASSIGN U1582 ( .B(clk), .A(\g.we_clk [14808]));
Q_ASSIGN U1583 ( .B(clk), .A(\g.we_clk [14807]));
Q_ASSIGN U1584 ( .B(clk), .A(\g.we_clk [14806]));
Q_ASSIGN U1585 ( .B(clk), .A(\g.we_clk [14805]));
Q_ASSIGN U1586 ( .B(clk), .A(\g.we_clk [14804]));
Q_ASSIGN U1587 ( .B(clk), .A(\g.we_clk [14803]));
Q_ASSIGN U1588 ( .B(clk), .A(\g.we_clk [14802]));
Q_ASSIGN U1589 ( .B(clk), .A(\g.we_clk [14801]));
Q_ASSIGN U1590 ( .B(clk), .A(\g.we_clk [14800]));
Q_ASSIGN U1591 ( .B(clk), .A(\g.we_clk [14799]));
Q_ASSIGN U1592 ( .B(clk), .A(\g.we_clk [14798]));
Q_ASSIGN U1593 ( .B(clk), .A(\g.we_clk [14797]));
Q_ASSIGN U1594 ( .B(clk), .A(\g.we_clk [14796]));
Q_ASSIGN U1595 ( .B(clk), .A(\g.we_clk [14795]));
Q_ASSIGN U1596 ( .B(clk), .A(\g.we_clk [14794]));
Q_ASSIGN U1597 ( .B(clk), .A(\g.we_clk [14793]));
Q_ASSIGN U1598 ( .B(clk), .A(\g.we_clk [14792]));
Q_ASSIGN U1599 ( .B(clk), .A(\g.we_clk [14791]));
Q_ASSIGN U1600 ( .B(clk), .A(\g.we_clk [14790]));
Q_ASSIGN U1601 ( .B(clk), .A(\g.we_clk [14789]));
Q_ASSIGN U1602 ( .B(clk), .A(\g.we_clk [14788]));
Q_ASSIGN U1603 ( .B(clk), .A(\g.we_clk [14787]));
Q_ASSIGN U1604 ( .B(clk), .A(\g.we_clk [14786]));
Q_ASSIGN U1605 ( .B(clk), .A(\g.we_clk [14785]));
Q_ASSIGN U1606 ( .B(clk), .A(\g.we_clk [14784]));
Q_ASSIGN U1607 ( .B(clk), .A(\g.we_clk [14783]));
Q_ASSIGN U1608 ( .B(clk), .A(\g.we_clk [14782]));
Q_ASSIGN U1609 ( .B(clk), .A(\g.we_clk [14781]));
Q_ASSIGN U1610 ( .B(clk), .A(\g.we_clk [14780]));
Q_ASSIGN U1611 ( .B(clk), .A(\g.we_clk [14779]));
Q_ASSIGN U1612 ( .B(clk), .A(\g.we_clk [14778]));
Q_ASSIGN U1613 ( .B(clk), .A(\g.we_clk [14777]));
Q_ASSIGN U1614 ( .B(clk), .A(\g.we_clk [14776]));
Q_ASSIGN U1615 ( .B(clk), .A(\g.we_clk [14775]));
Q_ASSIGN U1616 ( .B(clk), .A(\g.we_clk [14774]));
Q_ASSIGN U1617 ( .B(clk), .A(\g.we_clk [14773]));
Q_ASSIGN U1618 ( .B(clk), .A(\g.we_clk [14772]));
Q_ASSIGN U1619 ( .B(clk), .A(\g.we_clk [14771]));
Q_ASSIGN U1620 ( .B(clk), .A(\g.we_clk [14770]));
Q_ASSIGN U1621 ( .B(clk), .A(\g.we_clk [14769]));
Q_ASSIGN U1622 ( .B(clk), .A(\g.we_clk [14768]));
Q_ASSIGN U1623 ( .B(clk), .A(\g.we_clk [14767]));
Q_ASSIGN U1624 ( .B(clk), .A(\g.we_clk [14766]));
Q_ASSIGN U1625 ( .B(clk), .A(\g.we_clk [14765]));
Q_ASSIGN U1626 ( .B(clk), .A(\g.we_clk [14764]));
Q_ASSIGN U1627 ( .B(clk), .A(\g.we_clk [14763]));
Q_ASSIGN U1628 ( .B(clk), .A(\g.we_clk [14762]));
Q_ASSIGN U1629 ( .B(clk), .A(\g.we_clk [14761]));
Q_ASSIGN U1630 ( .B(clk), .A(\g.we_clk [14760]));
Q_ASSIGN U1631 ( .B(clk), .A(\g.we_clk [14759]));
Q_ASSIGN U1632 ( .B(clk), .A(\g.we_clk [14758]));
Q_ASSIGN U1633 ( .B(clk), .A(\g.we_clk [14757]));
Q_ASSIGN U1634 ( .B(clk), .A(\g.we_clk [14756]));
Q_ASSIGN U1635 ( .B(clk), .A(\g.we_clk [14755]));
Q_ASSIGN U1636 ( .B(clk), .A(\g.we_clk [14754]));
Q_ASSIGN U1637 ( .B(clk), .A(\g.we_clk [14753]));
Q_ASSIGN U1638 ( .B(clk), .A(\g.we_clk [14752]));
Q_ASSIGN U1639 ( .B(clk), .A(\g.we_clk [14751]));
Q_ASSIGN U1640 ( .B(clk), .A(\g.we_clk [14750]));
Q_ASSIGN U1641 ( .B(clk), .A(\g.we_clk [14749]));
Q_ASSIGN U1642 ( .B(clk), .A(\g.we_clk [14748]));
Q_ASSIGN U1643 ( .B(clk), .A(\g.we_clk [14747]));
Q_ASSIGN U1644 ( .B(clk), .A(\g.we_clk [14746]));
Q_ASSIGN U1645 ( .B(clk), .A(\g.we_clk [14745]));
Q_ASSIGN U1646 ( .B(clk), .A(\g.we_clk [14744]));
Q_ASSIGN U1647 ( .B(clk), .A(\g.we_clk [14743]));
Q_ASSIGN U1648 ( .B(clk), .A(\g.we_clk [14742]));
Q_ASSIGN U1649 ( .B(clk), .A(\g.we_clk [14741]));
Q_ASSIGN U1650 ( .B(clk), .A(\g.we_clk [14740]));
Q_ASSIGN U1651 ( .B(clk), .A(\g.we_clk [14739]));
Q_ASSIGN U1652 ( .B(clk), .A(\g.we_clk [14738]));
Q_ASSIGN U1653 ( .B(clk), .A(\g.we_clk [14737]));
Q_ASSIGN U1654 ( .B(clk), .A(\g.we_clk [14736]));
Q_ASSIGN U1655 ( .B(clk), .A(\g.we_clk [14735]));
Q_ASSIGN U1656 ( .B(clk), .A(\g.we_clk [14734]));
Q_ASSIGN U1657 ( .B(clk), .A(\g.we_clk [14733]));
Q_ASSIGN U1658 ( .B(clk), .A(\g.we_clk [14732]));
Q_ASSIGN U1659 ( .B(clk), .A(\g.we_clk [14731]));
Q_ASSIGN U1660 ( .B(clk), .A(\g.we_clk [14730]));
Q_ASSIGN U1661 ( .B(clk), .A(\g.we_clk [14729]));
Q_ASSIGN U1662 ( .B(clk), .A(\g.we_clk [14728]));
Q_ASSIGN U1663 ( .B(clk), .A(\g.we_clk [14727]));
Q_ASSIGN U1664 ( .B(clk), .A(\g.we_clk [14726]));
Q_ASSIGN U1665 ( .B(clk), .A(\g.we_clk [14725]));
Q_ASSIGN U1666 ( .B(clk), .A(\g.we_clk [14724]));
Q_ASSIGN U1667 ( .B(clk), .A(\g.we_clk [14723]));
Q_ASSIGN U1668 ( .B(clk), .A(\g.we_clk [14722]));
Q_ASSIGN U1669 ( .B(clk), .A(\g.we_clk [14721]));
Q_ASSIGN U1670 ( .B(clk), .A(\g.we_clk [14720]));
Q_ASSIGN U1671 ( .B(clk), .A(\g.we_clk [14719]));
Q_ASSIGN U1672 ( .B(clk), .A(\g.we_clk [14718]));
Q_ASSIGN U1673 ( .B(clk), .A(\g.we_clk [14717]));
Q_ASSIGN U1674 ( .B(clk), .A(\g.we_clk [14716]));
Q_ASSIGN U1675 ( .B(clk), .A(\g.we_clk [14715]));
Q_ASSIGN U1676 ( .B(clk), .A(\g.we_clk [14714]));
Q_ASSIGN U1677 ( .B(clk), .A(\g.we_clk [14713]));
Q_ASSIGN U1678 ( .B(clk), .A(\g.we_clk [14712]));
Q_ASSIGN U1679 ( .B(clk), .A(\g.we_clk [14711]));
Q_ASSIGN U1680 ( .B(clk), .A(\g.we_clk [14710]));
Q_ASSIGN U1681 ( .B(clk), .A(\g.we_clk [14709]));
Q_ASSIGN U1682 ( .B(clk), .A(\g.we_clk [14708]));
Q_ASSIGN U1683 ( .B(clk), .A(\g.we_clk [14707]));
Q_ASSIGN U1684 ( .B(clk), .A(\g.we_clk [14706]));
Q_ASSIGN U1685 ( .B(clk), .A(\g.we_clk [14705]));
Q_ASSIGN U1686 ( .B(clk), .A(\g.we_clk [14704]));
Q_ASSIGN U1687 ( .B(clk), .A(\g.we_clk [14703]));
Q_ASSIGN U1688 ( .B(clk), .A(\g.we_clk [14702]));
Q_ASSIGN U1689 ( .B(clk), .A(\g.we_clk [14701]));
Q_ASSIGN U1690 ( .B(clk), .A(\g.we_clk [14700]));
Q_ASSIGN U1691 ( .B(clk), .A(\g.we_clk [14699]));
Q_ASSIGN U1692 ( .B(clk), .A(\g.we_clk [14698]));
Q_ASSIGN U1693 ( .B(clk), .A(\g.we_clk [14697]));
Q_ASSIGN U1694 ( .B(clk), .A(\g.we_clk [14696]));
Q_ASSIGN U1695 ( .B(clk), .A(\g.we_clk [14695]));
Q_ASSIGN U1696 ( .B(clk), .A(\g.we_clk [14694]));
Q_ASSIGN U1697 ( .B(clk), .A(\g.we_clk [14693]));
Q_ASSIGN U1698 ( .B(clk), .A(\g.we_clk [14692]));
Q_ASSIGN U1699 ( .B(clk), .A(\g.we_clk [14691]));
Q_ASSIGN U1700 ( .B(clk), .A(\g.we_clk [14690]));
Q_ASSIGN U1701 ( .B(clk), .A(\g.we_clk [14689]));
Q_ASSIGN U1702 ( .B(clk), .A(\g.we_clk [14688]));
Q_ASSIGN U1703 ( .B(clk), .A(\g.we_clk [14687]));
Q_ASSIGN U1704 ( .B(clk), .A(\g.we_clk [14686]));
Q_ASSIGN U1705 ( .B(clk), .A(\g.we_clk [14685]));
Q_ASSIGN U1706 ( .B(clk), .A(\g.we_clk [14684]));
Q_ASSIGN U1707 ( .B(clk), .A(\g.we_clk [14683]));
Q_ASSIGN U1708 ( .B(clk), .A(\g.we_clk [14682]));
Q_ASSIGN U1709 ( .B(clk), .A(\g.we_clk [14681]));
Q_ASSIGN U1710 ( .B(clk), .A(\g.we_clk [14680]));
Q_ASSIGN U1711 ( .B(clk), .A(\g.we_clk [14679]));
Q_ASSIGN U1712 ( .B(clk), .A(\g.we_clk [14678]));
Q_ASSIGN U1713 ( .B(clk), .A(\g.we_clk [14677]));
Q_ASSIGN U1714 ( .B(clk), .A(\g.we_clk [14676]));
Q_ASSIGN U1715 ( .B(clk), .A(\g.we_clk [14675]));
Q_ASSIGN U1716 ( .B(clk), .A(\g.we_clk [14674]));
Q_ASSIGN U1717 ( .B(clk), .A(\g.we_clk [14673]));
Q_ASSIGN U1718 ( .B(clk), .A(\g.we_clk [14672]));
Q_ASSIGN U1719 ( .B(clk), .A(\g.we_clk [14671]));
Q_ASSIGN U1720 ( .B(clk), .A(\g.we_clk [14670]));
Q_ASSIGN U1721 ( .B(clk), .A(\g.we_clk [14669]));
Q_ASSIGN U1722 ( .B(clk), .A(\g.we_clk [14668]));
Q_ASSIGN U1723 ( .B(clk), .A(\g.we_clk [14667]));
Q_ASSIGN U1724 ( .B(clk), .A(\g.we_clk [14666]));
Q_ASSIGN U1725 ( .B(clk), .A(\g.we_clk [14665]));
Q_ASSIGN U1726 ( .B(clk), .A(\g.we_clk [14664]));
Q_ASSIGN U1727 ( .B(clk), .A(\g.we_clk [14663]));
Q_ASSIGN U1728 ( .B(clk), .A(\g.we_clk [14662]));
Q_ASSIGN U1729 ( .B(clk), .A(\g.we_clk [14661]));
Q_ASSIGN U1730 ( .B(clk), .A(\g.we_clk [14660]));
Q_ASSIGN U1731 ( .B(clk), .A(\g.we_clk [14659]));
Q_ASSIGN U1732 ( .B(clk), .A(\g.we_clk [14658]));
Q_ASSIGN U1733 ( .B(clk), .A(\g.we_clk [14657]));
Q_ASSIGN U1734 ( .B(clk), .A(\g.we_clk [14656]));
Q_ASSIGN U1735 ( .B(clk), .A(\g.we_clk [14655]));
Q_ASSIGN U1736 ( .B(clk), .A(\g.we_clk [14654]));
Q_ASSIGN U1737 ( .B(clk), .A(\g.we_clk [14653]));
Q_ASSIGN U1738 ( .B(clk), .A(\g.we_clk [14652]));
Q_ASSIGN U1739 ( .B(clk), .A(\g.we_clk [14651]));
Q_ASSIGN U1740 ( .B(clk), .A(\g.we_clk [14650]));
Q_ASSIGN U1741 ( .B(clk), .A(\g.we_clk [14649]));
Q_ASSIGN U1742 ( .B(clk), .A(\g.we_clk [14648]));
Q_ASSIGN U1743 ( .B(clk), .A(\g.we_clk [14647]));
Q_ASSIGN U1744 ( .B(clk), .A(\g.we_clk [14646]));
Q_ASSIGN U1745 ( .B(clk), .A(\g.we_clk [14645]));
Q_ASSIGN U1746 ( .B(clk), .A(\g.we_clk [14644]));
Q_ASSIGN U1747 ( .B(clk), .A(\g.we_clk [14643]));
Q_ASSIGN U1748 ( .B(clk), .A(\g.we_clk [14642]));
Q_ASSIGN U1749 ( .B(clk), .A(\g.we_clk [14641]));
Q_ASSIGN U1750 ( .B(clk), .A(\g.we_clk [14640]));
Q_ASSIGN U1751 ( .B(clk), .A(\g.we_clk [14639]));
Q_ASSIGN U1752 ( .B(clk), .A(\g.we_clk [14638]));
Q_ASSIGN U1753 ( .B(clk), .A(\g.we_clk [14637]));
Q_ASSIGN U1754 ( .B(clk), .A(\g.we_clk [14636]));
Q_ASSIGN U1755 ( .B(clk), .A(\g.we_clk [14635]));
Q_ASSIGN U1756 ( .B(clk), .A(\g.we_clk [14634]));
Q_ASSIGN U1757 ( .B(clk), .A(\g.we_clk [14633]));
Q_ASSIGN U1758 ( .B(clk), .A(\g.we_clk [14632]));
Q_ASSIGN U1759 ( .B(clk), .A(\g.we_clk [14631]));
Q_ASSIGN U1760 ( .B(clk), .A(\g.we_clk [14630]));
Q_ASSIGN U1761 ( .B(clk), .A(\g.we_clk [14629]));
Q_ASSIGN U1762 ( .B(clk), .A(\g.we_clk [14628]));
Q_ASSIGN U1763 ( .B(clk), .A(\g.we_clk [14627]));
Q_ASSIGN U1764 ( .B(clk), .A(\g.we_clk [14626]));
Q_ASSIGN U1765 ( .B(clk), .A(\g.we_clk [14625]));
Q_ASSIGN U1766 ( .B(clk), .A(\g.we_clk [14624]));
Q_ASSIGN U1767 ( .B(clk), .A(\g.we_clk [14623]));
Q_ASSIGN U1768 ( .B(clk), .A(\g.we_clk [14622]));
Q_ASSIGN U1769 ( .B(clk), .A(\g.we_clk [14621]));
Q_ASSIGN U1770 ( .B(clk), .A(\g.we_clk [14620]));
Q_ASSIGN U1771 ( .B(clk), .A(\g.we_clk [14619]));
Q_ASSIGN U1772 ( .B(clk), .A(\g.we_clk [14618]));
Q_ASSIGN U1773 ( .B(clk), .A(\g.we_clk [14617]));
Q_ASSIGN U1774 ( .B(clk), .A(\g.we_clk [14616]));
Q_ASSIGN U1775 ( .B(clk), .A(\g.we_clk [14615]));
Q_ASSIGN U1776 ( .B(clk), .A(\g.we_clk [14614]));
Q_ASSIGN U1777 ( .B(clk), .A(\g.we_clk [14613]));
Q_ASSIGN U1778 ( .B(clk), .A(\g.we_clk [14612]));
Q_ASSIGN U1779 ( .B(clk), .A(\g.we_clk [14611]));
Q_ASSIGN U1780 ( .B(clk), .A(\g.we_clk [14610]));
Q_ASSIGN U1781 ( .B(clk), .A(\g.we_clk [14609]));
Q_ASSIGN U1782 ( .B(clk), .A(\g.we_clk [14608]));
Q_ASSIGN U1783 ( .B(clk), .A(\g.we_clk [14607]));
Q_ASSIGN U1784 ( .B(clk), .A(\g.we_clk [14606]));
Q_ASSIGN U1785 ( .B(clk), .A(\g.we_clk [14605]));
Q_ASSIGN U1786 ( .B(clk), .A(\g.we_clk [14604]));
Q_ASSIGN U1787 ( .B(clk), .A(\g.we_clk [14603]));
Q_ASSIGN U1788 ( .B(clk), .A(\g.we_clk [14602]));
Q_ASSIGN U1789 ( .B(clk), .A(\g.we_clk [14601]));
Q_ASSIGN U1790 ( .B(clk), .A(\g.we_clk [14600]));
Q_ASSIGN U1791 ( .B(clk), .A(\g.we_clk [14599]));
Q_ASSIGN U1792 ( .B(clk), .A(\g.we_clk [14598]));
Q_ASSIGN U1793 ( .B(clk), .A(\g.we_clk [14597]));
Q_ASSIGN U1794 ( .B(clk), .A(\g.we_clk [14596]));
Q_ASSIGN U1795 ( .B(clk), .A(\g.we_clk [14595]));
Q_ASSIGN U1796 ( .B(clk), .A(\g.we_clk [14594]));
Q_ASSIGN U1797 ( .B(clk), .A(\g.we_clk [14593]));
Q_ASSIGN U1798 ( .B(clk), .A(\g.we_clk [14592]));
Q_ASSIGN U1799 ( .B(clk), .A(\g.we_clk [14591]));
Q_ASSIGN U1800 ( .B(clk), .A(\g.we_clk [14590]));
Q_ASSIGN U1801 ( .B(clk), .A(\g.we_clk [14589]));
Q_ASSIGN U1802 ( .B(clk), .A(\g.we_clk [14588]));
Q_ASSIGN U1803 ( .B(clk), .A(\g.we_clk [14587]));
Q_ASSIGN U1804 ( .B(clk), .A(\g.we_clk [14586]));
Q_ASSIGN U1805 ( .B(clk), .A(\g.we_clk [14585]));
Q_ASSIGN U1806 ( .B(clk), .A(\g.we_clk [14584]));
Q_ASSIGN U1807 ( .B(clk), .A(\g.we_clk [14583]));
Q_ASSIGN U1808 ( .B(clk), .A(\g.we_clk [14582]));
Q_ASSIGN U1809 ( .B(clk), .A(\g.we_clk [14581]));
Q_ASSIGN U1810 ( .B(clk), .A(\g.we_clk [14580]));
Q_ASSIGN U1811 ( .B(clk), .A(\g.we_clk [14579]));
Q_ASSIGN U1812 ( .B(clk), .A(\g.we_clk [14578]));
Q_ASSIGN U1813 ( .B(clk), .A(\g.we_clk [14577]));
Q_ASSIGN U1814 ( .B(clk), .A(\g.we_clk [14576]));
Q_ASSIGN U1815 ( .B(clk), .A(\g.we_clk [14575]));
Q_ASSIGN U1816 ( .B(clk), .A(\g.we_clk [14574]));
Q_ASSIGN U1817 ( .B(clk), .A(\g.we_clk [14573]));
Q_ASSIGN U1818 ( .B(clk), .A(\g.we_clk [14572]));
Q_ASSIGN U1819 ( .B(clk), .A(\g.we_clk [14571]));
Q_ASSIGN U1820 ( .B(clk), .A(\g.we_clk [14570]));
Q_ASSIGN U1821 ( .B(clk), .A(\g.we_clk [14569]));
Q_ASSIGN U1822 ( .B(clk), .A(\g.we_clk [14568]));
Q_ASSIGN U1823 ( .B(clk), .A(\g.we_clk [14567]));
Q_ASSIGN U1824 ( .B(clk), .A(\g.we_clk [14566]));
Q_ASSIGN U1825 ( .B(clk), .A(\g.we_clk [14565]));
Q_ASSIGN U1826 ( .B(clk), .A(\g.we_clk [14564]));
Q_ASSIGN U1827 ( .B(clk), .A(\g.we_clk [14563]));
Q_ASSIGN U1828 ( .B(clk), .A(\g.we_clk [14562]));
Q_ASSIGN U1829 ( .B(clk), .A(\g.we_clk [14561]));
Q_ASSIGN U1830 ( .B(clk), .A(\g.we_clk [14560]));
Q_ASSIGN U1831 ( .B(clk), .A(\g.we_clk [14559]));
Q_ASSIGN U1832 ( .B(clk), .A(\g.we_clk [14558]));
Q_ASSIGN U1833 ( .B(clk), .A(\g.we_clk [14557]));
Q_ASSIGN U1834 ( .B(clk), .A(\g.we_clk [14556]));
Q_ASSIGN U1835 ( .B(clk), .A(\g.we_clk [14555]));
Q_ASSIGN U1836 ( .B(clk), .A(\g.we_clk [14554]));
Q_ASSIGN U1837 ( .B(clk), .A(\g.we_clk [14553]));
Q_ASSIGN U1838 ( .B(clk), .A(\g.we_clk [14552]));
Q_ASSIGN U1839 ( .B(clk), .A(\g.we_clk [14551]));
Q_ASSIGN U1840 ( .B(clk), .A(\g.we_clk [14550]));
Q_ASSIGN U1841 ( .B(clk), .A(\g.we_clk [14549]));
Q_ASSIGN U1842 ( .B(clk), .A(\g.we_clk [14548]));
Q_ASSIGN U1843 ( .B(clk), .A(\g.we_clk [14547]));
Q_ASSIGN U1844 ( .B(clk), .A(\g.we_clk [14546]));
Q_ASSIGN U1845 ( .B(clk), .A(\g.we_clk [14545]));
Q_ASSIGN U1846 ( .B(clk), .A(\g.we_clk [14544]));
Q_ASSIGN U1847 ( .B(clk), .A(\g.we_clk [14543]));
Q_ASSIGN U1848 ( .B(clk), .A(\g.we_clk [14542]));
Q_ASSIGN U1849 ( .B(clk), .A(\g.we_clk [14541]));
Q_ASSIGN U1850 ( .B(clk), .A(\g.we_clk [14540]));
Q_ASSIGN U1851 ( .B(clk), .A(\g.we_clk [14539]));
Q_ASSIGN U1852 ( .B(clk), .A(\g.we_clk [14538]));
Q_ASSIGN U1853 ( .B(clk), .A(\g.we_clk [14537]));
Q_ASSIGN U1854 ( .B(clk), .A(\g.we_clk [14536]));
Q_ASSIGN U1855 ( .B(clk), .A(\g.we_clk [14535]));
Q_ASSIGN U1856 ( .B(clk), .A(\g.we_clk [14534]));
Q_ASSIGN U1857 ( .B(clk), .A(\g.we_clk [14533]));
Q_ASSIGN U1858 ( .B(clk), .A(\g.we_clk [14532]));
Q_ASSIGN U1859 ( .B(clk), .A(\g.we_clk [14531]));
Q_ASSIGN U1860 ( .B(clk), .A(\g.we_clk [14530]));
Q_ASSIGN U1861 ( .B(clk), .A(\g.we_clk [14529]));
Q_ASSIGN U1862 ( .B(clk), .A(\g.we_clk [14528]));
Q_ASSIGN U1863 ( .B(clk), .A(\g.we_clk [14527]));
Q_ASSIGN U1864 ( .B(clk), .A(\g.we_clk [14526]));
Q_ASSIGN U1865 ( .B(clk), .A(\g.we_clk [14525]));
Q_ASSIGN U1866 ( .B(clk), .A(\g.we_clk [14524]));
Q_ASSIGN U1867 ( .B(clk), .A(\g.we_clk [14523]));
Q_ASSIGN U1868 ( .B(clk), .A(\g.we_clk [14522]));
Q_ASSIGN U1869 ( .B(clk), .A(\g.we_clk [14521]));
Q_ASSIGN U1870 ( .B(clk), .A(\g.we_clk [14520]));
Q_ASSIGN U1871 ( .B(clk), .A(\g.we_clk [14519]));
Q_ASSIGN U1872 ( .B(clk), .A(\g.we_clk [14518]));
Q_ASSIGN U1873 ( .B(clk), .A(\g.we_clk [14517]));
Q_ASSIGN U1874 ( .B(clk), .A(\g.we_clk [14516]));
Q_ASSIGN U1875 ( .B(clk), .A(\g.we_clk [14515]));
Q_ASSIGN U1876 ( .B(clk), .A(\g.we_clk [14514]));
Q_ASSIGN U1877 ( .B(clk), .A(\g.we_clk [14513]));
Q_ASSIGN U1878 ( .B(clk), .A(\g.we_clk [14512]));
Q_ASSIGN U1879 ( .B(clk), .A(\g.we_clk [14511]));
Q_ASSIGN U1880 ( .B(clk), .A(\g.we_clk [14510]));
Q_ASSIGN U1881 ( .B(clk), .A(\g.we_clk [14509]));
Q_ASSIGN U1882 ( .B(clk), .A(\g.we_clk [14508]));
Q_ASSIGN U1883 ( .B(clk), .A(\g.we_clk [14507]));
Q_ASSIGN U1884 ( .B(clk), .A(\g.we_clk [14506]));
Q_ASSIGN U1885 ( .B(clk), .A(\g.we_clk [14505]));
Q_ASSIGN U1886 ( .B(clk), .A(\g.we_clk [14504]));
Q_ASSIGN U1887 ( .B(clk), .A(\g.we_clk [14503]));
Q_ASSIGN U1888 ( .B(clk), .A(\g.we_clk [14502]));
Q_ASSIGN U1889 ( .B(clk), .A(\g.we_clk [14501]));
Q_ASSIGN U1890 ( .B(clk), .A(\g.we_clk [14500]));
Q_ASSIGN U1891 ( .B(clk), .A(\g.we_clk [14499]));
Q_ASSIGN U1892 ( .B(clk), .A(\g.we_clk [14498]));
Q_ASSIGN U1893 ( .B(clk), .A(\g.we_clk [14497]));
Q_ASSIGN U1894 ( .B(clk), .A(\g.we_clk [14496]));
Q_ASSIGN U1895 ( .B(clk), .A(\g.we_clk [14495]));
Q_ASSIGN U1896 ( .B(clk), .A(\g.we_clk [14494]));
Q_ASSIGN U1897 ( .B(clk), .A(\g.we_clk [14493]));
Q_ASSIGN U1898 ( .B(clk), .A(\g.we_clk [14492]));
Q_ASSIGN U1899 ( .B(clk), .A(\g.we_clk [14491]));
Q_ASSIGN U1900 ( .B(clk), .A(\g.we_clk [14490]));
Q_ASSIGN U1901 ( .B(clk), .A(\g.we_clk [14489]));
Q_ASSIGN U1902 ( .B(clk), .A(\g.we_clk [14488]));
Q_ASSIGN U1903 ( .B(clk), .A(\g.we_clk [14487]));
Q_ASSIGN U1904 ( .B(clk), .A(\g.we_clk [14486]));
Q_ASSIGN U1905 ( .B(clk), .A(\g.we_clk [14485]));
Q_ASSIGN U1906 ( .B(clk), .A(\g.we_clk [14484]));
Q_ASSIGN U1907 ( .B(clk), .A(\g.we_clk [14483]));
Q_ASSIGN U1908 ( .B(clk), .A(\g.we_clk [14482]));
Q_ASSIGN U1909 ( .B(clk), .A(\g.we_clk [14481]));
Q_ASSIGN U1910 ( .B(clk), .A(\g.we_clk [14480]));
Q_ASSIGN U1911 ( .B(clk), .A(\g.we_clk [14479]));
Q_ASSIGN U1912 ( .B(clk), .A(\g.we_clk [14478]));
Q_ASSIGN U1913 ( .B(clk), .A(\g.we_clk [14477]));
Q_ASSIGN U1914 ( .B(clk), .A(\g.we_clk [14476]));
Q_ASSIGN U1915 ( .B(clk), .A(\g.we_clk [14475]));
Q_ASSIGN U1916 ( .B(clk), .A(\g.we_clk [14474]));
Q_ASSIGN U1917 ( .B(clk), .A(\g.we_clk [14473]));
Q_ASSIGN U1918 ( .B(clk), .A(\g.we_clk [14472]));
Q_ASSIGN U1919 ( .B(clk), .A(\g.we_clk [14471]));
Q_ASSIGN U1920 ( .B(clk), .A(\g.we_clk [14470]));
Q_ASSIGN U1921 ( .B(clk), .A(\g.we_clk [14469]));
Q_ASSIGN U1922 ( .B(clk), .A(\g.we_clk [14468]));
Q_ASSIGN U1923 ( .B(clk), .A(\g.we_clk [14467]));
Q_ASSIGN U1924 ( .B(clk), .A(\g.we_clk [14466]));
Q_ASSIGN U1925 ( .B(clk), .A(\g.we_clk [14465]));
Q_ASSIGN U1926 ( .B(clk), .A(\g.we_clk [14464]));
Q_ASSIGN U1927 ( .B(clk), .A(\g.we_clk [14463]));
Q_ASSIGN U1928 ( .B(clk), .A(\g.we_clk [14462]));
Q_ASSIGN U1929 ( .B(clk), .A(\g.we_clk [14461]));
Q_ASSIGN U1930 ( .B(clk), .A(\g.we_clk [14460]));
Q_ASSIGN U1931 ( .B(clk), .A(\g.we_clk [14459]));
Q_ASSIGN U1932 ( .B(clk), .A(\g.we_clk [14458]));
Q_ASSIGN U1933 ( .B(clk), .A(\g.we_clk [14457]));
Q_ASSIGN U1934 ( .B(clk), .A(\g.we_clk [14456]));
Q_ASSIGN U1935 ( .B(clk), .A(\g.we_clk [14455]));
Q_ASSIGN U1936 ( .B(clk), .A(\g.we_clk [14454]));
Q_ASSIGN U1937 ( .B(clk), .A(\g.we_clk [14453]));
Q_ASSIGN U1938 ( .B(clk), .A(\g.we_clk [14452]));
Q_ASSIGN U1939 ( .B(clk), .A(\g.we_clk [14451]));
Q_ASSIGN U1940 ( .B(clk), .A(\g.we_clk [14450]));
Q_ASSIGN U1941 ( .B(clk), .A(\g.we_clk [14449]));
Q_ASSIGN U1942 ( .B(clk), .A(\g.we_clk [14448]));
Q_ASSIGN U1943 ( .B(clk), .A(\g.we_clk [14447]));
Q_ASSIGN U1944 ( .B(clk), .A(\g.we_clk [14446]));
Q_ASSIGN U1945 ( .B(clk), .A(\g.we_clk [14445]));
Q_ASSIGN U1946 ( .B(clk), .A(\g.we_clk [14444]));
Q_ASSIGN U1947 ( .B(clk), .A(\g.we_clk [14443]));
Q_ASSIGN U1948 ( .B(clk), .A(\g.we_clk [14442]));
Q_ASSIGN U1949 ( .B(clk), .A(\g.we_clk [14441]));
Q_ASSIGN U1950 ( .B(clk), .A(\g.we_clk [14440]));
Q_ASSIGN U1951 ( .B(clk), .A(\g.we_clk [14439]));
Q_ASSIGN U1952 ( .B(clk), .A(\g.we_clk [14438]));
Q_ASSIGN U1953 ( .B(clk), .A(\g.we_clk [14437]));
Q_ASSIGN U1954 ( .B(clk), .A(\g.we_clk [14436]));
Q_ASSIGN U1955 ( .B(clk), .A(\g.we_clk [14435]));
Q_ASSIGN U1956 ( .B(clk), .A(\g.we_clk [14434]));
Q_ASSIGN U1957 ( .B(clk), .A(\g.we_clk [14433]));
Q_ASSIGN U1958 ( .B(clk), .A(\g.we_clk [14432]));
Q_ASSIGN U1959 ( .B(clk), .A(\g.we_clk [14431]));
Q_ASSIGN U1960 ( .B(clk), .A(\g.we_clk [14430]));
Q_ASSIGN U1961 ( .B(clk), .A(\g.we_clk [14429]));
Q_ASSIGN U1962 ( .B(clk), .A(\g.we_clk [14428]));
Q_ASSIGN U1963 ( .B(clk), .A(\g.we_clk [14427]));
Q_ASSIGN U1964 ( .B(clk), .A(\g.we_clk [14426]));
Q_ASSIGN U1965 ( .B(clk), .A(\g.we_clk [14425]));
Q_ASSIGN U1966 ( .B(clk), .A(\g.we_clk [14424]));
Q_ASSIGN U1967 ( .B(clk), .A(\g.we_clk [14423]));
Q_ASSIGN U1968 ( .B(clk), .A(\g.we_clk [14422]));
Q_ASSIGN U1969 ( .B(clk), .A(\g.we_clk [14421]));
Q_ASSIGN U1970 ( .B(clk), .A(\g.we_clk [14420]));
Q_ASSIGN U1971 ( .B(clk), .A(\g.we_clk [14419]));
Q_ASSIGN U1972 ( .B(clk), .A(\g.we_clk [14418]));
Q_ASSIGN U1973 ( .B(clk), .A(\g.we_clk [14417]));
Q_ASSIGN U1974 ( .B(clk), .A(\g.we_clk [14416]));
Q_ASSIGN U1975 ( .B(clk), .A(\g.we_clk [14415]));
Q_ASSIGN U1976 ( .B(clk), .A(\g.we_clk [14414]));
Q_ASSIGN U1977 ( .B(clk), .A(\g.we_clk [14413]));
Q_ASSIGN U1978 ( .B(clk), .A(\g.we_clk [14412]));
Q_ASSIGN U1979 ( .B(clk), .A(\g.we_clk [14411]));
Q_ASSIGN U1980 ( .B(clk), .A(\g.we_clk [14410]));
Q_ASSIGN U1981 ( .B(clk), .A(\g.we_clk [14409]));
Q_ASSIGN U1982 ( .B(clk), .A(\g.we_clk [14408]));
Q_ASSIGN U1983 ( .B(clk), .A(\g.we_clk [14407]));
Q_ASSIGN U1984 ( .B(clk), .A(\g.we_clk [14406]));
Q_ASSIGN U1985 ( .B(clk), .A(\g.we_clk [14405]));
Q_ASSIGN U1986 ( .B(clk), .A(\g.we_clk [14404]));
Q_ASSIGN U1987 ( .B(clk), .A(\g.we_clk [14403]));
Q_ASSIGN U1988 ( .B(clk), .A(\g.we_clk [14402]));
Q_ASSIGN U1989 ( .B(clk), .A(\g.we_clk [14401]));
Q_ASSIGN U1990 ( .B(clk), .A(\g.we_clk [14400]));
Q_ASSIGN U1991 ( .B(clk), .A(\g.we_clk [14399]));
Q_ASSIGN U1992 ( .B(clk), .A(\g.we_clk [14398]));
Q_ASSIGN U1993 ( .B(clk), .A(\g.we_clk [14397]));
Q_ASSIGN U1994 ( .B(clk), .A(\g.we_clk [14396]));
Q_ASSIGN U1995 ( .B(clk), .A(\g.we_clk [14395]));
Q_ASSIGN U1996 ( .B(clk), .A(\g.we_clk [14394]));
Q_ASSIGN U1997 ( .B(clk), .A(\g.we_clk [14393]));
Q_ASSIGN U1998 ( .B(clk), .A(\g.we_clk [14392]));
Q_ASSIGN U1999 ( .B(clk), .A(\g.we_clk [14391]));
Q_ASSIGN U2000 ( .B(clk), .A(\g.we_clk [14390]));
Q_ASSIGN U2001 ( .B(clk), .A(\g.we_clk [14389]));
Q_ASSIGN U2002 ( .B(clk), .A(\g.we_clk [14388]));
Q_ASSIGN U2003 ( .B(clk), .A(\g.we_clk [14387]));
Q_ASSIGN U2004 ( .B(clk), .A(\g.we_clk [14386]));
Q_ASSIGN U2005 ( .B(clk), .A(\g.we_clk [14385]));
Q_ASSIGN U2006 ( .B(clk), .A(\g.we_clk [14384]));
Q_ASSIGN U2007 ( .B(clk), .A(\g.we_clk [14383]));
Q_ASSIGN U2008 ( .B(clk), .A(\g.we_clk [14382]));
Q_ASSIGN U2009 ( .B(clk), .A(\g.we_clk [14381]));
Q_ASSIGN U2010 ( .B(clk), .A(\g.we_clk [14380]));
Q_ASSIGN U2011 ( .B(clk), .A(\g.we_clk [14379]));
Q_ASSIGN U2012 ( .B(clk), .A(\g.we_clk [14378]));
Q_ASSIGN U2013 ( .B(clk), .A(\g.we_clk [14377]));
Q_ASSIGN U2014 ( .B(clk), .A(\g.we_clk [14376]));
Q_ASSIGN U2015 ( .B(clk), .A(\g.we_clk [14375]));
Q_ASSIGN U2016 ( .B(clk), .A(\g.we_clk [14374]));
Q_ASSIGN U2017 ( .B(clk), .A(\g.we_clk [14373]));
Q_ASSIGN U2018 ( .B(clk), .A(\g.we_clk [14372]));
Q_ASSIGN U2019 ( .B(clk), .A(\g.we_clk [14371]));
Q_ASSIGN U2020 ( .B(clk), .A(\g.we_clk [14370]));
Q_ASSIGN U2021 ( .B(clk), .A(\g.we_clk [14369]));
Q_ASSIGN U2022 ( .B(clk), .A(\g.we_clk [14368]));
Q_ASSIGN U2023 ( .B(clk), .A(\g.we_clk [14367]));
Q_ASSIGN U2024 ( .B(clk), .A(\g.we_clk [14366]));
Q_ASSIGN U2025 ( .B(clk), .A(\g.we_clk [14365]));
Q_ASSIGN U2026 ( .B(clk), .A(\g.we_clk [14364]));
Q_ASSIGN U2027 ( .B(clk), .A(\g.we_clk [14363]));
Q_ASSIGN U2028 ( .B(clk), .A(\g.we_clk [14362]));
Q_ASSIGN U2029 ( .B(clk), .A(\g.we_clk [14361]));
Q_ASSIGN U2030 ( .B(clk), .A(\g.we_clk [14360]));
Q_ASSIGN U2031 ( .B(clk), .A(\g.we_clk [14359]));
Q_ASSIGN U2032 ( .B(clk), .A(\g.we_clk [14358]));
Q_ASSIGN U2033 ( .B(clk), .A(\g.we_clk [14357]));
Q_ASSIGN U2034 ( .B(clk), .A(\g.we_clk [14356]));
Q_ASSIGN U2035 ( .B(clk), .A(\g.we_clk [14355]));
Q_ASSIGN U2036 ( .B(clk), .A(\g.we_clk [14354]));
Q_ASSIGN U2037 ( .B(clk), .A(\g.we_clk [14353]));
Q_ASSIGN U2038 ( .B(clk), .A(\g.we_clk [14352]));
Q_ASSIGN U2039 ( .B(clk), .A(\g.we_clk [14351]));
Q_ASSIGN U2040 ( .B(clk), .A(\g.we_clk [14350]));
Q_ASSIGN U2041 ( .B(clk), .A(\g.we_clk [14349]));
Q_ASSIGN U2042 ( .B(clk), .A(\g.we_clk [14348]));
Q_ASSIGN U2043 ( .B(clk), .A(\g.we_clk [14347]));
Q_ASSIGN U2044 ( .B(clk), .A(\g.we_clk [14346]));
Q_ASSIGN U2045 ( .B(clk), .A(\g.we_clk [14345]));
Q_ASSIGN U2046 ( .B(clk), .A(\g.we_clk [14344]));
Q_ASSIGN U2047 ( .B(clk), .A(\g.we_clk [14343]));
Q_ASSIGN U2048 ( .B(clk), .A(\g.we_clk [14342]));
Q_ASSIGN U2049 ( .B(clk), .A(\g.we_clk [14341]));
Q_ASSIGN U2050 ( .B(clk), .A(\g.we_clk [14340]));
Q_ASSIGN U2051 ( .B(clk), .A(\g.we_clk [14339]));
Q_ASSIGN U2052 ( .B(clk), .A(\g.we_clk [14338]));
Q_ASSIGN U2053 ( .B(clk), .A(\g.we_clk [14337]));
Q_ASSIGN U2054 ( .B(clk), .A(\g.we_clk [14336]));
Q_ASSIGN U2055 ( .B(clk), .A(\g.we_clk [14335]));
Q_ASSIGN U2056 ( .B(clk), .A(\g.we_clk [14334]));
Q_ASSIGN U2057 ( .B(clk), .A(\g.we_clk [14333]));
Q_ASSIGN U2058 ( .B(clk), .A(\g.we_clk [14332]));
Q_ASSIGN U2059 ( .B(clk), .A(\g.we_clk [14331]));
Q_ASSIGN U2060 ( .B(clk), .A(\g.we_clk [14330]));
Q_ASSIGN U2061 ( .B(clk), .A(\g.we_clk [14329]));
Q_ASSIGN U2062 ( .B(clk), .A(\g.we_clk [14328]));
Q_ASSIGN U2063 ( .B(clk), .A(\g.we_clk [14327]));
Q_ASSIGN U2064 ( .B(clk), .A(\g.we_clk [14326]));
Q_ASSIGN U2065 ( .B(clk), .A(\g.we_clk [14325]));
Q_ASSIGN U2066 ( .B(clk), .A(\g.we_clk [14324]));
Q_ASSIGN U2067 ( .B(clk), .A(\g.we_clk [14323]));
Q_ASSIGN U2068 ( .B(clk), .A(\g.we_clk [14322]));
Q_ASSIGN U2069 ( .B(clk), .A(\g.we_clk [14321]));
Q_ASSIGN U2070 ( .B(clk), .A(\g.we_clk [14320]));
Q_ASSIGN U2071 ( .B(clk), .A(\g.we_clk [14319]));
Q_ASSIGN U2072 ( .B(clk), .A(\g.we_clk [14318]));
Q_ASSIGN U2073 ( .B(clk), .A(\g.we_clk [14317]));
Q_ASSIGN U2074 ( .B(clk), .A(\g.we_clk [14316]));
Q_ASSIGN U2075 ( .B(clk), .A(\g.we_clk [14315]));
Q_ASSIGN U2076 ( .B(clk), .A(\g.we_clk [14314]));
Q_ASSIGN U2077 ( .B(clk), .A(\g.we_clk [14313]));
Q_ASSIGN U2078 ( .B(clk), .A(\g.we_clk [14312]));
Q_ASSIGN U2079 ( .B(clk), .A(\g.we_clk [14311]));
Q_ASSIGN U2080 ( .B(clk), .A(\g.we_clk [14310]));
Q_ASSIGN U2081 ( .B(clk), .A(\g.we_clk [14309]));
Q_ASSIGN U2082 ( .B(clk), .A(\g.we_clk [14308]));
Q_ASSIGN U2083 ( .B(clk), .A(\g.we_clk [14307]));
Q_ASSIGN U2084 ( .B(clk), .A(\g.we_clk [14306]));
Q_ASSIGN U2085 ( .B(clk), .A(\g.we_clk [14305]));
Q_ASSIGN U2086 ( .B(clk), .A(\g.we_clk [14304]));
Q_ASSIGN U2087 ( .B(clk), .A(\g.we_clk [14303]));
Q_ASSIGN U2088 ( .B(clk), .A(\g.we_clk [14302]));
Q_ASSIGN U2089 ( .B(clk), .A(\g.we_clk [14301]));
Q_ASSIGN U2090 ( .B(clk), .A(\g.we_clk [14300]));
Q_ASSIGN U2091 ( .B(clk), .A(\g.we_clk [14299]));
Q_ASSIGN U2092 ( .B(clk), .A(\g.we_clk [14298]));
Q_ASSIGN U2093 ( .B(clk), .A(\g.we_clk [14297]));
Q_ASSIGN U2094 ( .B(clk), .A(\g.we_clk [14296]));
Q_ASSIGN U2095 ( .B(clk), .A(\g.we_clk [14295]));
Q_ASSIGN U2096 ( .B(clk), .A(\g.we_clk [14294]));
Q_ASSIGN U2097 ( .B(clk), .A(\g.we_clk [14293]));
Q_ASSIGN U2098 ( .B(clk), .A(\g.we_clk [14292]));
Q_ASSIGN U2099 ( .B(clk), .A(\g.we_clk [14291]));
Q_ASSIGN U2100 ( .B(clk), .A(\g.we_clk [14290]));
Q_ASSIGN U2101 ( .B(clk), .A(\g.we_clk [14289]));
Q_ASSIGN U2102 ( .B(clk), .A(\g.we_clk [14288]));
Q_ASSIGN U2103 ( .B(clk), .A(\g.we_clk [14287]));
Q_ASSIGN U2104 ( .B(clk), .A(\g.we_clk [14286]));
Q_ASSIGN U2105 ( .B(clk), .A(\g.we_clk [14285]));
Q_ASSIGN U2106 ( .B(clk), .A(\g.we_clk [14284]));
Q_ASSIGN U2107 ( .B(clk), .A(\g.we_clk [14283]));
Q_ASSIGN U2108 ( .B(clk), .A(\g.we_clk [14282]));
Q_ASSIGN U2109 ( .B(clk), .A(\g.we_clk [14281]));
Q_ASSIGN U2110 ( .B(clk), .A(\g.we_clk [14280]));
Q_ASSIGN U2111 ( .B(clk), .A(\g.we_clk [14279]));
Q_ASSIGN U2112 ( .B(clk), .A(\g.we_clk [14278]));
Q_ASSIGN U2113 ( .B(clk), .A(\g.we_clk [14277]));
Q_ASSIGN U2114 ( .B(clk), .A(\g.we_clk [14276]));
Q_ASSIGN U2115 ( .B(clk), .A(\g.we_clk [14275]));
Q_ASSIGN U2116 ( .B(clk), .A(\g.we_clk [14274]));
Q_ASSIGN U2117 ( .B(clk), .A(\g.we_clk [14273]));
Q_ASSIGN U2118 ( .B(clk), .A(\g.we_clk [14272]));
Q_ASSIGN U2119 ( .B(clk), .A(\g.we_clk [14271]));
Q_ASSIGN U2120 ( .B(clk), .A(\g.we_clk [14270]));
Q_ASSIGN U2121 ( .B(clk), .A(\g.we_clk [14269]));
Q_ASSIGN U2122 ( .B(clk), .A(\g.we_clk [14268]));
Q_ASSIGN U2123 ( .B(clk), .A(\g.we_clk [14267]));
Q_ASSIGN U2124 ( .B(clk), .A(\g.we_clk [14266]));
Q_ASSIGN U2125 ( .B(clk), .A(\g.we_clk [14265]));
Q_ASSIGN U2126 ( .B(clk), .A(\g.we_clk [14264]));
Q_ASSIGN U2127 ( .B(clk), .A(\g.we_clk [14263]));
Q_ASSIGN U2128 ( .B(clk), .A(\g.we_clk [14262]));
Q_ASSIGN U2129 ( .B(clk), .A(\g.we_clk [14261]));
Q_ASSIGN U2130 ( .B(clk), .A(\g.we_clk [14260]));
Q_ASSIGN U2131 ( .B(clk), .A(\g.we_clk [14259]));
Q_ASSIGN U2132 ( .B(clk), .A(\g.we_clk [14258]));
Q_ASSIGN U2133 ( .B(clk), .A(\g.we_clk [14257]));
Q_ASSIGN U2134 ( .B(clk), .A(\g.we_clk [14256]));
Q_ASSIGN U2135 ( .B(clk), .A(\g.we_clk [14255]));
Q_ASSIGN U2136 ( .B(clk), .A(\g.we_clk [14254]));
Q_ASSIGN U2137 ( .B(clk), .A(\g.we_clk [14253]));
Q_ASSIGN U2138 ( .B(clk), .A(\g.we_clk [14252]));
Q_ASSIGN U2139 ( .B(clk), .A(\g.we_clk [14251]));
Q_ASSIGN U2140 ( .B(clk), .A(\g.we_clk [14250]));
Q_ASSIGN U2141 ( .B(clk), .A(\g.we_clk [14249]));
Q_ASSIGN U2142 ( .B(clk), .A(\g.we_clk [14248]));
Q_ASSIGN U2143 ( .B(clk), .A(\g.we_clk [14247]));
Q_ASSIGN U2144 ( .B(clk), .A(\g.we_clk [14246]));
Q_ASSIGN U2145 ( .B(clk), .A(\g.we_clk [14245]));
Q_ASSIGN U2146 ( .B(clk), .A(\g.we_clk [14244]));
Q_ASSIGN U2147 ( .B(clk), .A(\g.we_clk [14243]));
Q_ASSIGN U2148 ( .B(clk), .A(\g.we_clk [14242]));
Q_ASSIGN U2149 ( .B(clk), .A(\g.we_clk [14241]));
Q_ASSIGN U2150 ( .B(clk), .A(\g.we_clk [14240]));
Q_ASSIGN U2151 ( .B(clk), .A(\g.we_clk [14239]));
Q_ASSIGN U2152 ( .B(clk), .A(\g.we_clk [14238]));
Q_ASSIGN U2153 ( .B(clk), .A(\g.we_clk [14237]));
Q_ASSIGN U2154 ( .B(clk), .A(\g.we_clk [14236]));
Q_ASSIGN U2155 ( .B(clk), .A(\g.we_clk [14235]));
Q_ASSIGN U2156 ( .B(clk), .A(\g.we_clk [14234]));
Q_ASSIGN U2157 ( .B(clk), .A(\g.we_clk [14233]));
Q_ASSIGN U2158 ( .B(clk), .A(\g.we_clk [14232]));
Q_ASSIGN U2159 ( .B(clk), .A(\g.we_clk [14231]));
Q_ASSIGN U2160 ( .B(clk), .A(\g.we_clk [14230]));
Q_ASSIGN U2161 ( .B(clk), .A(\g.we_clk [14229]));
Q_ASSIGN U2162 ( .B(clk), .A(\g.we_clk [14228]));
Q_ASSIGN U2163 ( .B(clk), .A(\g.we_clk [14227]));
Q_ASSIGN U2164 ( .B(clk), .A(\g.we_clk [14226]));
Q_ASSIGN U2165 ( .B(clk), .A(\g.we_clk [14225]));
Q_ASSIGN U2166 ( .B(clk), .A(\g.we_clk [14224]));
Q_ASSIGN U2167 ( .B(clk), .A(\g.we_clk [14223]));
Q_ASSIGN U2168 ( .B(clk), .A(\g.we_clk [14222]));
Q_ASSIGN U2169 ( .B(clk), .A(\g.we_clk [14221]));
Q_ASSIGN U2170 ( .B(clk), .A(\g.we_clk [14220]));
Q_ASSIGN U2171 ( .B(clk), .A(\g.we_clk [14219]));
Q_ASSIGN U2172 ( .B(clk), .A(\g.we_clk [14218]));
Q_ASSIGN U2173 ( .B(clk), .A(\g.we_clk [14217]));
Q_ASSIGN U2174 ( .B(clk), .A(\g.we_clk [14216]));
Q_ASSIGN U2175 ( .B(clk), .A(\g.we_clk [14215]));
Q_ASSIGN U2176 ( .B(clk), .A(\g.we_clk [14214]));
Q_ASSIGN U2177 ( .B(clk), .A(\g.we_clk [14213]));
Q_ASSIGN U2178 ( .B(clk), .A(\g.we_clk [14212]));
Q_ASSIGN U2179 ( .B(clk), .A(\g.we_clk [14211]));
Q_ASSIGN U2180 ( .B(clk), .A(\g.we_clk [14210]));
Q_ASSIGN U2181 ( .B(clk), .A(\g.we_clk [14209]));
Q_ASSIGN U2182 ( .B(clk), .A(\g.we_clk [14208]));
Q_ASSIGN U2183 ( .B(clk), .A(\g.we_clk [14207]));
Q_ASSIGN U2184 ( .B(clk), .A(\g.we_clk [14206]));
Q_ASSIGN U2185 ( .B(clk), .A(\g.we_clk [14205]));
Q_ASSIGN U2186 ( .B(clk), .A(\g.we_clk [14204]));
Q_ASSIGN U2187 ( .B(clk), .A(\g.we_clk [14203]));
Q_ASSIGN U2188 ( .B(clk), .A(\g.we_clk [14202]));
Q_ASSIGN U2189 ( .B(clk), .A(\g.we_clk [14201]));
Q_ASSIGN U2190 ( .B(clk), .A(\g.we_clk [14200]));
Q_ASSIGN U2191 ( .B(clk), .A(\g.we_clk [14199]));
Q_ASSIGN U2192 ( .B(clk), .A(\g.we_clk [14198]));
Q_ASSIGN U2193 ( .B(clk), .A(\g.we_clk [14197]));
Q_ASSIGN U2194 ( .B(clk), .A(\g.we_clk [14196]));
Q_ASSIGN U2195 ( .B(clk), .A(\g.we_clk [14195]));
Q_ASSIGN U2196 ( .B(clk), .A(\g.we_clk [14194]));
Q_ASSIGN U2197 ( .B(clk), .A(\g.we_clk [14193]));
Q_ASSIGN U2198 ( .B(clk), .A(\g.we_clk [14192]));
Q_ASSIGN U2199 ( .B(clk), .A(\g.we_clk [14191]));
Q_ASSIGN U2200 ( .B(clk), .A(\g.we_clk [14190]));
Q_ASSIGN U2201 ( .B(clk), .A(\g.we_clk [14189]));
Q_ASSIGN U2202 ( .B(clk), .A(\g.we_clk [14188]));
Q_ASSIGN U2203 ( .B(clk), .A(\g.we_clk [14187]));
Q_ASSIGN U2204 ( .B(clk), .A(\g.we_clk [14186]));
Q_ASSIGN U2205 ( .B(clk), .A(\g.we_clk [14185]));
Q_ASSIGN U2206 ( .B(clk), .A(\g.we_clk [14184]));
Q_ASSIGN U2207 ( .B(clk), .A(\g.we_clk [14183]));
Q_ASSIGN U2208 ( .B(clk), .A(\g.we_clk [14182]));
Q_ASSIGN U2209 ( .B(clk), .A(\g.we_clk [14181]));
Q_ASSIGN U2210 ( .B(clk), .A(\g.we_clk [14180]));
Q_ASSIGN U2211 ( .B(clk), .A(\g.we_clk [14179]));
Q_ASSIGN U2212 ( .B(clk), .A(\g.we_clk [14178]));
Q_ASSIGN U2213 ( .B(clk), .A(\g.we_clk [14177]));
Q_ASSIGN U2214 ( .B(clk), .A(\g.we_clk [14176]));
Q_ASSIGN U2215 ( .B(clk), .A(\g.we_clk [14175]));
Q_ASSIGN U2216 ( .B(clk), .A(\g.we_clk [14174]));
Q_ASSIGN U2217 ( .B(clk), .A(\g.we_clk [14173]));
Q_ASSIGN U2218 ( .B(clk), .A(\g.we_clk [14172]));
Q_ASSIGN U2219 ( .B(clk), .A(\g.we_clk [14171]));
Q_ASSIGN U2220 ( .B(clk), .A(\g.we_clk [14170]));
Q_ASSIGN U2221 ( .B(clk), .A(\g.we_clk [14169]));
Q_ASSIGN U2222 ( .B(clk), .A(\g.we_clk [14168]));
Q_ASSIGN U2223 ( .B(clk), .A(\g.we_clk [14167]));
Q_ASSIGN U2224 ( .B(clk), .A(\g.we_clk [14166]));
Q_ASSIGN U2225 ( .B(clk), .A(\g.we_clk [14165]));
Q_ASSIGN U2226 ( .B(clk), .A(\g.we_clk [14164]));
Q_ASSIGN U2227 ( .B(clk), .A(\g.we_clk [14163]));
Q_ASSIGN U2228 ( .B(clk), .A(\g.we_clk [14162]));
Q_ASSIGN U2229 ( .B(clk), .A(\g.we_clk [14161]));
Q_ASSIGN U2230 ( .B(clk), .A(\g.we_clk [14160]));
Q_ASSIGN U2231 ( .B(clk), .A(\g.we_clk [14159]));
Q_ASSIGN U2232 ( .B(clk), .A(\g.we_clk [14158]));
Q_ASSIGN U2233 ( .B(clk), .A(\g.we_clk [14157]));
Q_ASSIGN U2234 ( .B(clk), .A(\g.we_clk [14156]));
Q_ASSIGN U2235 ( .B(clk), .A(\g.we_clk [14155]));
Q_ASSIGN U2236 ( .B(clk), .A(\g.we_clk [14154]));
Q_ASSIGN U2237 ( .B(clk), .A(\g.we_clk [14153]));
Q_ASSIGN U2238 ( .B(clk), .A(\g.we_clk [14152]));
Q_ASSIGN U2239 ( .B(clk), .A(\g.we_clk [14151]));
Q_ASSIGN U2240 ( .B(clk), .A(\g.we_clk [14150]));
Q_ASSIGN U2241 ( .B(clk), .A(\g.we_clk [14149]));
Q_ASSIGN U2242 ( .B(clk), .A(\g.we_clk [14148]));
Q_ASSIGN U2243 ( .B(clk), .A(\g.we_clk [14147]));
Q_ASSIGN U2244 ( .B(clk), .A(\g.we_clk [14146]));
Q_ASSIGN U2245 ( .B(clk), .A(\g.we_clk [14145]));
Q_ASSIGN U2246 ( .B(clk), .A(\g.we_clk [14144]));
Q_ASSIGN U2247 ( .B(clk), .A(\g.we_clk [14143]));
Q_ASSIGN U2248 ( .B(clk), .A(\g.we_clk [14142]));
Q_ASSIGN U2249 ( .B(clk), .A(\g.we_clk [14141]));
Q_ASSIGN U2250 ( .B(clk), .A(\g.we_clk [14140]));
Q_ASSIGN U2251 ( .B(clk), .A(\g.we_clk [14139]));
Q_ASSIGN U2252 ( .B(clk), .A(\g.we_clk [14138]));
Q_ASSIGN U2253 ( .B(clk), .A(\g.we_clk [14137]));
Q_ASSIGN U2254 ( .B(clk), .A(\g.we_clk [14136]));
Q_ASSIGN U2255 ( .B(clk), .A(\g.we_clk [14135]));
Q_ASSIGN U2256 ( .B(clk), .A(\g.we_clk [14134]));
Q_ASSIGN U2257 ( .B(clk), .A(\g.we_clk [14133]));
Q_ASSIGN U2258 ( .B(clk), .A(\g.we_clk [14132]));
Q_ASSIGN U2259 ( .B(clk), .A(\g.we_clk [14131]));
Q_ASSIGN U2260 ( .B(clk), .A(\g.we_clk [14130]));
Q_ASSIGN U2261 ( .B(clk), .A(\g.we_clk [14129]));
Q_ASSIGN U2262 ( .B(clk), .A(\g.we_clk [14128]));
Q_ASSIGN U2263 ( .B(clk), .A(\g.we_clk [14127]));
Q_ASSIGN U2264 ( .B(clk), .A(\g.we_clk [14126]));
Q_ASSIGN U2265 ( .B(clk), .A(\g.we_clk [14125]));
Q_ASSIGN U2266 ( .B(clk), .A(\g.we_clk [14124]));
Q_ASSIGN U2267 ( .B(clk), .A(\g.we_clk [14123]));
Q_ASSIGN U2268 ( .B(clk), .A(\g.we_clk [14122]));
Q_ASSIGN U2269 ( .B(clk), .A(\g.we_clk [14121]));
Q_ASSIGN U2270 ( .B(clk), .A(\g.we_clk [14120]));
Q_ASSIGN U2271 ( .B(clk), .A(\g.we_clk [14119]));
Q_ASSIGN U2272 ( .B(clk), .A(\g.we_clk [14118]));
Q_ASSIGN U2273 ( .B(clk), .A(\g.we_clk [14117]));
Q_ASSIGN U2274 ( .B(clk), .A(\g.we_clk [14116]));
Q_ASSIGN U2275 ( .B(clk), .A(\g.we_clk [14115]));
Q_ASSIGN U2276 ( .B(clk), .A(\g.we_clk [14114]));
Q_ASSIGN U2277 ( .B(clk), .A(\g.we_clk [14113]));
Q_ASSIGN U2278 ( .B(clk), .A(\g.we_clk [14112]));
Q_ASSIGN U2279 ( .B(clk), .A(\g.we_clk [14111]));
Q_ASSIGN U2280 ( .B(clk), .A(\g.we_clk [14110]));
Q_ASSIGN U2281 ( .B(clk), .A(\g.we_clk [14109]));
Q_ASSIGN U2282 ( .B(clk), .A(\g.we_clk [14108]));
Q_ASSIGN U2283 ( .B(clk), .A(\g.we_clk [14107]));
Q_ASSIGN U2284 ( .B(clk), .A(\g.we_clk [14106]));
Q_ASSIGN U2285 ( .B(clk), .A(\g.we_clk [14105]));
Q_ASSIGN U2286 ( .B(clk), .A(\g.we_clk [14104]));
Q_ASSIGN U2287 ( .B(clk), .A(\g.we_clk [14103]));
Q_ASSIGN U2288 ( .B(clk), .A(\g.we_clk [14102]));
Q_ASSIGN U2289 ( .B(clk), .A(\g.we_clk [14101]));
Q_ASSIGN U2290 ( .B(clk), .A(\g.we_clk [14100]));
Q_ASSIGN U2291 ( .B(clk), .A(\g.we_clk [14099]));
Q_ASSIGN U2292 ( .B(clk), .A(\g.we_clk [14098]));
Q_ASSIGN U2293 ( .B(clk), .A(\g.we_clk [14097]));
Q_ASSIGN U2294 ( .B(clk), .A(\g.we_clk [14096]));
Q_ASSIGN U2295 ( .B(clk), .A(\g.we_clk [14095]));
Q_ASSIGN U2296 ( .B(clk), .A(\g.we_clk [14094]));
Q_ASSIGN U2297 ( .B(clk), .A(\g.we_clk [14093]));
Q_ASSIGN U2298 ( .B(clk), .A(\g.we_clk [14092]));
Q_ASSIGN U2299 ( .B(clk), .A(\g.we_clk [14091]));
Q_ASSIGN U2300 ( .B(clk), .A(\g.we_clk [14090]));
Q_ASSIGN U2301 ( .B(clk), .A(\g.we_clk [14089]));
Q_ASSIGN U2302 ( .B(clk), .A(\g.we_clk [14088]));
Q_ASSIGN U2303 ( .B(clk), .A(\g.we_clk [14087]));
Q_ASSIGN U2304 ( .B(clk), .A(\g.we_clk [14086]));
Q_ASSIGN U2305 ( .B(clk), .A(\g.we_clk [14085]));
Q_ASSIGN U2306 ( .B(clk), .A(\g.we_clk [14084]));
Q_ASSIGN U2307 ( .B(clk), .A(\g.we_clk [14083]));
Q_ASSIGN U2308 ( .B(clk), .A(\g.we_clk [14082]));
Q_ASSIGN U2309 ( .B(clk), .A(\g.we_clk [14081]));
Q_ASSIGN U2310 ( .B(clk), .A(\g.we_clk [14080]));
Q_ASSIGN U2311 ( .B(clk), .A(\g.we_clk [14079]));
Q_ASSIGN U2312 ( .B(clk), .A(\g.we_clk [14078]));
Q_ASSIGN U2313 ( .B(clk), .A(\g.we_clk [14077]));
Q_ASSIGN U2314 ( .B(clk), .A(\g.we_clk [14076]));
Q_ASSIGN U2315 ( .B(clk), .A(\g.we_clk [14075]));
Q_ASSIGN U2316 ( .B(clk), .A(\g.we_clk [14074]));
Q_ASSIGN U2317 ( .B(clk), .A(\g.we_clk [14073]));
Q_ASSIGN U2318 ( .B(clk), .A(\g.we_clk [14072]));
Q_ASSIGN U2319 ( .B(clk), .A(\g.we_clk [14071]));
Q_ASSIGN U2320 ( .B(clk), .A(\g.we_clk [14070]));
Q_ASSIGN U2321 ( .B(clk), .A(\g.we_clk [14069]));
Q_ASSIGN U2322 ( .B(clk), .A(\g.we_clk [14068]));
Q_ASSIGN U2323 ( .B(clk), .A(\g.we_clk [14067]));
Q_ASSIGN U2324 ( .B(clk), .A(\g.we_clk [14066]));
Q_ASSIGN U2325 ( .B(clk), .A(\g.we_clk [14065]));
Q_ASSIGN U2326 ( .B(clk), .A(\g.we_clk [14064]));
Q_ASSIGN U2327 ( .B(clk), .A(\g.we_clk [14063]));
Q_ASSIGN U2328 ( .B(clk), .A(\g.we_clk [14062]));
Q_ASSIGN U2329 ( .B(clk), .A(\g.we_clk [14061]));
Q_ASSIGN U2330 ( .B(clk), .A(\g.we_clk [14060]));
Q_ASSIGN U2331 ( .B(clk), .A(\g.we_clk [14059]));
Q_ASSIGN U2332 ( .B(clk), .A(\g.we_clk [14058]));
Q_ASSIGN U2333 ( .B(clk), .A(\g.we_clk [14057]));
Q_ASSIGN U2334 ( .B(clk), .A(\g.we_clk [14056]));
Q_ASSIGN U2335 ( .B(clk), .A(\g.we_clk [14055]));
Q_ASSIGN U2336 ( .B(clk), .A(\g.we_clk [14054]));
Q_ASSIGN U2337 ( .B(clk), .A(\g.we_clk [14053]));
Q_ASSIGN U2338 ( .B(clk), .A(\g.we_clk [14052]));
Q_ASSIGN U2339 ( .B(clk), .A(\g.we_clk [14051]));
Q_ASSIGN U2340 ( .B(clk), .A(\g.we_clk [14050]));
Q_ASSIGN U2341 ( .B(clk), .A(\g.we_clk [14049]));
Q_ASSIGN U2342 ( .B(clk), .A(\g.we_clk [14048]));
Q_ASSIGN U2343 ( .B(clk), .A(\g.we_clk [14047]));
Q_ASSIGN U2344 ( .B(clk), .A(\g.we_clk [14046]));
Q_ASSIGN U2345 ( .B(clk), .A(\g.we_clk [14045]));
Q_ASSIGN U2346 ( .B(clk), .A(\g.we_clk [14044]));
Q_ASSIGN U2347 ( .B(clk), .A(\g.we_clk [14043]));
Q_ASSIGN U2348 ( .B(clk), .A(\g.we_clk [14042]));
Q_ASSIGN U2349 ( .B(clk), .A(\g.we_clk [14041]));
Q_ASSIGN U2350 ( .B(clk), .A(\g.we_clk [14040]));
Q_ASSIGN U2351 ( .B(clk), .A(\g.we_clk [14039]));
Q_ASSIGN U2352 ( .B(clk), .A(\g.we_clk [14038]));
Q_ASSIGN U2353 ( .B(clk), .A(\g.we_clk [14037]));
Q_ASSIGN U2354 ( .B(clk), .A(\g.we_clk [14036]));
Q_ASSIGN U2355 ( .B(clk), .A(\g.we_clk [14035]));
Q_ASSIGN U2356 ( .B(clk), .A(\g.we_clk [14034]));
Q_ASSIGN U2357 ( .B(clk), .A(\g.we_clk [14033]));
Q_ASSIGN U2358 ( .B(clk), .A(\g.we_clk [14032]));
Q_ASSIGN U2359 ( .B(clk), .A(\g.we_clk [14031]));
Q_ASSIGN U2360 ( .B(clk), .A(\g.we_clk [14030]));
Q_ASSIGN U2361 ( .B(clk), .A(\g.we_clk [14029]));
Q_ASSIGN U2362 ( .B(clk), .A(\g.we_clk [14028]));
Q_ASSIGN U2363 ( .B(clk), .A(\g.we_clk [14027]));
Q_ASSIGN U2364 ( .B(clk), .A(\g.we_clk [14026]));
Q_ASSIGN U2365 ( .B(clk), .A(\g.we_clk [14025]));
Q_ASSIGN U2366 ( .B(clk), .A(\g.we_clk [14024]));
Q_ASSIGN U2367 ( .B(clk), .A(\g.we_clk [14023]));
Q_ASSIGN U2368 ( .B(clk), .A(\g.we_clk [14022]));
Q_ASSIGN U2369 ( .B(clk), .A(\g.we_clk [14021]));
Q_ASSIGN U2370 ( .B(clk), .A(\g.we_clk [14020]));
Q_ASSIGN U2371 ( .B(clk), .A(\g.we_clk [14019]));
Q_ASSIGN U2372 ( .B(clk), .A(\g.we_clk [14018]));
Q_ASSIGN U2373 ( .B(clk), .A(\g.we_clk [14017]));
Q_ASSIGN U2374 ( .B(clk), .A(\g.we_clk [14016]));
Q_ASSIGN U2375 ( .B(clk), .A(\g.we_clk [14015]));
Q_ASSIGN U2376 ( .B(clk), .A(\g.we_clk [14014]));
Q_ASSIGN U2377 ( .B(clk), .A(\g.we_clk [14013]));
Q_ASSIGN U2378 ( .B(clk), .A(\g.we_clk [14012]));
Q_ASSIGN U2379 ( .B(clk), .A(\g.we_clk [14011]));
Q_ASSIGN U2380 ( .B(clk), .A(\g.we_clk [14010]));
Q_ASSIGN U2381 ( .B(clk), .A(\g.we_clk [14009]));
Q_ASSIGN U2382 ( .B(clk), .A(\g.we_clk [14008]));
Q_ASSIGN U2383 ( .B(clk), .A(\g.we_clk [14007]));
Q_ASSIGN U2384 ( .B(clk), .A(\g.we_clk [14006]));
Q_ASSIGN U2385 ( .B(clk), .A(\g.we_clk [14005]));
Q_ASSIGN U2386 ( .B(clk), .A(\g.we_clk [14004]));
Q_ASSIGN U2387 ( .B(clk), .A(\g.we_clk [14003]));
Q_ASSIGN U2388 ( .B(clk), .A(\g.we_clk [14002]));
Q_ASSIGN U2389 ( .B(clk), .A(\g.we_clk [14001]));
Q_ASSIGN U2390 ( .B(clk), .A(\g.we_clk [14000]));
Q_ASSIGN U2391 ( .B(clk), .A(\g.we_clk [13999]));
Q_ASSIGN U2392 ( .B(clk), .A(\g.we_clk [13998]));
Q_ASSIGN U2393 ( .B(clk), .A(\g.we_clk [13997]));
Q_ASSIGN U2394 ( .B(clk), .A(\g.we_clk [13996]));
Q_ASSIGN U2395 ( .B(clk), .A(\g.we_clk [13995]));
Q_ASSIGN U2396 ( .B(clk), .A(\g.we_clk [13994]));
Q_ASSIGN U2397 ( .B(clk), .A(\g.we_clk [13993]));
Q_ASSIGN U2398 ( .B(clk), .A(\g.we_clk [13992]));
Q_ASSIGN U2399 ( .B(clk), .A(\g.we_clk [13991]));
Q_ASSIGN U2400 ( .B(clk), .A(\g.we_clk [13990]));
Q_ASSIGN U2401 ( .B(clk), .A(\g.we_clk [13989]));
Q_ASSIGN U2402 ( .B(clk), .A(\g.we_clk [13988]));
Q_ASSIGN U2403 ( .B(clk), .A(\g.we_clk [13987]));
Q_ASSIGN U2404 ( .B(clk), .A(\g.we_clk [13986]));
Q_ASSIGN U2405 ( .B(clk), .A(\g.we_clk [13985]));
Q_ASSIGN U2406 ( .B(clk), .A(\g.we_clk [13984]));
Q_ASSIGN U2407 ( .B(clk), .A(\g.we_clk [13983]));
Q_ASSIGN U2408 ( .B(clk), .A(\g.we_clk [13982]));
Q_ASSIGN U2409 ( .B(clk), .A(\g.we_clk [13981]));
Q_ASSIGN U2410 ( .B(clk), .A(\g.we_clk [13980]));
Q_ASSIGN U2411 ( .B(clk), .A(\g.we_clk [13979]));
Q_ASSIGN U2412 ( .B(clk), .A(\g.we_clk [13978]));
Q_ASSIGN U2413 ( .B(clk), .A(\g.we_clk [13977]));
Q_ASSIGN U2414 ( .B(clk), .A(\g.we_clk [13976]));
Q_ASSIGN U2415 ( .B(clk), .A(\g.we_clk [13975]));
Q_ASSIGN U2416 ( .B(clk), .A(\g.we_clk [13974]));
Q_ASSIGN U2417 ( .B(clk), .A(\g.we_clk [13973]));
Q_ASSIGN U2418 ( .B(clk), .A(\g.we_clk [13972]));
Q_ASSIGN U2419 ( .B(clk), .A(\g.we_clk [13971]));
Q_ASSIGN U2420 ( .B(clk), .A(\g.we_clk [13970]));
Q_ASSIGN U2421 ( .B(clk), .A(\g.we_clk [13969]));
Q_ASSIGN U2422 ( .B(clk), .A(\g.we_clk [13968]));
Q_ASSIGN U2423 ( .B(clk), .A(\g.we_clk [13967]));
Q_ASSIGN U2424 ( .B(clk), .A(\g.we_clk [13966]));
Q_ASSIGN U2425 ( .B(clk), .A(\g.we_clk [13965]));
Q_ASSIGN U2426 ( .B(clk), .A(\g.we_clk [13964]));
Q_ASSIGN U2427 ( .B(clk), .A(\g.we_clk [13963]));
Q_ASSIGN U2428 ( .B(clk), .A(\g.we_clk [13962]));
Q_ASSIGN U2429 ( .B(clk), .A(\g.we_clk [13961]));
Q_ASSIGN U2430 ( .B(clk), .A(\g.we_clk [13960]));
Q_ASSIGN U2431 ( .B(clk), .A(\g.we_clk [13959]));
Q_ASSIGN U2432 ( .B(clk), .A(\g.we_clk [13958]));
Q_ASSIGN U2433 ( .B(clk), .A(\g.we_clk [13957]));
Q_ASSIGN U2434 ( .B(clk), .A(\g.we_clk [13956]));
Q_ASSIGN U2435 ( .B(clk), .A(\g.we_clk [13955]));
Q_ASSIGN U2436 ( .B(clk), .A(\g.we_clk [13954]));
Q_ASSIGN U2437 ( .B(clk), .A(\g.we_clk [13953]));
Q_ASSIGN U2438 ( .B(clk), .A(\g.we_clk [13952]));
Q_ASSIGN U2439 ( .B(clk), .A(\g.we_clk [13951]));
Q_ASSIGN U2440 ( .B(clk), .A(\g.we_clk [13950]));
Q_ASSIGN U2441 ( .B(clk), .A(\g.we_clk [13949]));
Q_ASSIGN U2442 ( .B(clk), .A(\g.we_clk [13948]));
Q_ASSIGN U2443 ( .B(clk), .A(\g.we_clk [13947]));
Q_ASSIGN U2444 ( .B(clk), .A(\g.we_clk [13946]));
Q_ASSIGN U2445 ( .B(clk), .A(\g.we_clk [13945]));
Q_ASSIGN U2446 ( .B(clk), .A(\g.we_clk [13944]));
Q_ASSIGN U2447 ( .B(clk), .A(\g.we_clk [13943]));
Q_ASSIGN U2448 ( .B(clk), .A(\g.we_clk [13942]));
Q_ASSIGN U2449 ( .B(clk), .A(\g.we_clk [13941]));
Q_ASSIGN U2450 ( .B(clk), .A(\g.we_clk [13940]));
Q_ASSIGN U2451 ( .B(clk), .A(\g.we_clk [13939]));
Q_ASSIGN U2452 ( .B(clk), .A(\g.we_clk [13938]));
Q_ASSIGN U2453 ( .B(clk), .A(\g.we_clk [13937]));
Q_ASSIGN U2454 ( .B(clk), .A(\g.we_clk [13936]));
Q_ASSIGN U2455 ( .B(clk), .A(\g.we_clk [13935]));
Q_ASSIGN U2456 ( .B(clk), .A(\g.we_clk [13934]));
Q_ASSIGN U2457 ( .B(clk), .A(\g.we_clk [13933]));
Q_ASSIGN U2458 ( .B(clk), .A(\g.we_clk [13932]));
Q_ASSIGN U2459 ( .B(clk), .A(\g.we_clk [13931]));
Q_ASSIGN U2460 ( .B(clk), .A(\g.we_clk [13930]));
Q_ASSIGN U2461 ( .B(clk), .A(\g.we_clk [13929]));
Q_ASSIGN U2462 ( .B(clk), .A(\g.we_clk [13928]));
Q_ASSIGN U2463 ( .B(clk), .A(\g.we_clk [13927]));
Q_ASSIGN U2464 ( .B(clk), .A(\g.we_clk [13926]));
Q_ASSIGN U2465 ( .B(clk), .A(\g.we_clk [13925]));
Q_ASSIGN U2466 ( .B(clk), .A(\g.we_clk [13924]));
Q_ASSIGN U2467 ( .B(clk), .A(\g.we_clk [13923]));
Q_ASSIGN U2468 ( .B(clk), .A(\g.we_clk [13922]));
Q_ASSIGN U2469 ( .B(clk), .A(\g.we_clk [13921]));
Q_ASSIGN U2470 ( .B(clk), .A(\g.we_clk [13920]));
Q_ASSIGN U2471 ( .B(clk), .A(\g.we_clk [13919]));
Q_ASSIGN U2472 ( .B(clk), .A(\g.we_clk [13918]));
Q_ASSIGN U2473 ( .B(clk), .A(\g.we_clk [13917]));
Q_ASSIGN U2474 ( .B(clk), .A(\g.we_clk [13916]));
Q_ASSIGN U2475 ( .B(clk), .A(\g.we_clk [13915]));
Q_ASSIGN U2476 ( .B(clk), .A(\g.we_clk [13914]));
Q_ASSIGN U2477 ( .B(clk), .A(\g.we_clk [13913]));
Q_ASSIGN U2478 ( .B(clk), .A(\g.we_clk [13912]));
Q_ASSIGN U2479 ( .B(clk), .A(\g.we_clk [13911]));
Q_ASSIGN U2480 ( .B(clk), .A(\g.we_clk [13910]));
Q_ASSIGN U2481 ( .B(clk), .A(\g.we_clk [13909]));
Q_ASSIGN U2482 ( .B(clk), .A(\g.we_clk [13908]));
Q_ASSIGN U2483 ( .B(clk), .A(\g.we_clk [13907]));
Q_ASSIGN U2484 ( .B(clk), .A(\g.we_clk [13906]));
Q_ASSIGN U2485 ( .B(clk), .A(\g.we_clk [13905]));
Q_ASSIGN U2486 ( .B(clk), .A(\g.we_clk [13904]));
Q_ASSIGN U2487 ( .B(clk), .A(\g.we_clk [13903]));
Q_ASSIGN U2488 ( .B(clk), .A(\g.we_clk [13902]));
Q_ASSIGN U2489 ( .B(clk), .A(\g.we_clk [13901]));
Q_ASSIGN U2490 ( .B(clk), .A(\g.we_clk [13900]));
Q_ASSIGN U2491 ( .B(clk), .A(\g.we_clk [13899]));
Q_ASSIGN U2492 ( .B(clk), .A(\g.we_clk [13898]));
Q_ASSIGN U2493 ( .B(clk), .A(\g.we_clk [13897]));
Q_ASSIGN U2494 ( .B(clk), .A(\g.we_clk [13896]));
Q_ASSIGN U2495 ( .B(clk), .A(\g.we_clk [13895]));
Q_ASSIGN U2496 ( .B(clk), .A(\g.we_clk [13894]));
Q_ASSIGN U2497 ( .B(clk), .A(\g.we_clk [13893]));
Q_ASSIGN U2498 ( .B(clk), .A(\g.we_clk [13892]));
Q_ASSIGN U2499 ( .B(clk), .A(\g.we_clk [13891]));
Q_ASSIGN U2500 ( .B(clk), .A(\g.we_clk [13890]));
Q_ASSIGN U2501 ( .B(clk), .A(\g.we_clk [13889]));
Q_ASSIGN U2502 ( .B(clk), .A(\g.we_clk [13888]));
Q_ASSIGN U2503 ( .B(clk), .A(\g.we_clk [13887]));
Q_ASSIGN U2504 ( .B(clk), .A(\g.we_clk [13886]));
Q_ASSIGN U2505 ( .B(clk), .A(\g.we_clk [13885]));
Q_ASSIGN U2506 ( .B(clk), .A(\g.we_clk [13884]));
Q_ASSIGN U2507 ( .B(clk), .A(\g.we_clk [13883]));
Q_ASSIGN U2508 ( .B(clk), .A(\g.we_clk [13882]));
Q_ASSIGN U2509 ( .B(clk), .A(\g.we_clk [13881]));
Q_ASSIGN U2510 ( .B(clk), .A(\g.we_clk [13880]));
Q_ASSIGN U2511 ( .B(clk), .A(\g.we_clk [13879]));
Q_ASSIGN U2512 ( .B(clk), .A(\g.we_clk [13878]));
Q_ASSIGN U2513 ( .B(clk), .A(\g.we_clk [13877]));
Q_ASSIGN U2514 ( .B(clk), .A(\g.we_clk [13876]));
Q_ASSIGN U2515 ( .B(clk), .A(\g.we_clk [13875]));
Q_ASSIGN U2516 ( .B(clk), .A(\g.we_clk [13874]));
Q_ASSIGN U2517 ( .B(clk), .A(\g.we_clk [13873]));
Q_ASSIGN U2518 ( .B(clk), .A(\g.we_clk [13872]));
Q_ASSIGN U2519 ( .B(clk), .A(\g.we_clk [13871]));
Q_ASSIGN U2520 ( .B(clk), .A(\g.we_clk [13870]));
Q_ASSIGN U2521 ( .B(clk), .A(\g.we_clk [13869]));
Q_ASSIGN U2522 ( .B(clk), .A(\g.we_clk [13868]));
Q_ASSIGN U2523 ( .B(clk), .A(\g.we_clk [13867]));
Q_ASSIGN U2524 ( .B(clk), .A(\g.we_clk [13866]));
Q_ASSIGN U2525 ( .B(clk), .A(\g.we_clk [13865]));
Q_ASSIGN U2526 ( .B(clk), .A(\g.we_clk [13864]));
Q_ASSIGN U2527 ( .B(clk), .A(\g.we_clk [13863]));
Q_ASSIGN U2528 ( .B(clk), .A(\g.we_clk [13862]));
Q_ASSIGN U2529 ( .B(clk), .A(\g.we_clk [13861]));
Q_ASSIGN U2530 ( .B(clk), .A(\g.we_clk [13860]));
Q_ASSIGN U2531 ( .B(clk), .A(\g.we_clk [13859]));
Q_ASSIGN U2532 ( .B(clk), .A(\g.we_clk [13858]));
Q_ASSIGN U2533 ( .B(clk), .A(\g.we_clk [13857]));
Q_ASSIGN U2534 ( .B(clk), .A(\g.we_clk [13856]));
Q_ASSIGN U2535 ( .B(clk), .A(\g.we_clk [13855]));
Q_ASSIGN U2536 ( .B(clk), .A(\g.we_clk [13854]));
Q_ASSIGN U2537 ( .B(clk), .A(\g.we_clk [13853]));
Q_ASSIGN U2538 ( .B(clk), .A(\g.we_clk [13852]));
Q_ASSIGN U2539 ( .B(clk), .A(\g.we_clk [13851]));
Q_ASSIGN U2540 ( .B(clk), .A(\g.we_clk [13850]));
Q_ASSIGN U2541 ( .B(clk), .A(\g.we_clk [13849]));
Q_ASSIGN U2542 ( .B(clk), .A(\g.we_clk [13848]));
Q_ASSIGN U2543 ( .B(clk), .A(\g.we_clk [13847]));
Q_ASSIGN U2544 ( .B(clk), .A(\g.we_clk [13846]));
Q_ASSIGN U2545 ( .B(clk), .A(\g.we_clk [13845]));
Q_ASSIGN U2546 ( .B(clk), .A(\g.we_clk [13844]));
Q_ASSIGN U2547 ( .B(clk), .A(\g.we_clk [13843]));
Q_ASSIGN U2548 ( .B(clk), .A(\g.we_clk [13842]));
Q_ASSIGN U2549 ( .B(clk), .A(\g.we_clk [13841]));
Q_ASSIGN U2550 ( .B(clk), .A(\g.we_clk [13840]));
Q_ASSIGN U2551 ( .B(clk), .A(\g.we_clk [13839]));
Q_ASSIGN U2552 ( .B(clk), .A(\g.we_clk [13838]));
Q_ASSIGN U2553 ( .B(clk), .A(\g.we_clk [13837]));
Q_ASSIGN U2554 ( .B(clk), .A(\g.we_clk [13836]));
Q_ASSIGN U2555 ( .B(clk), .A(\g.we_clk [13835]));
Q_ASSIGN U2556 ( .B(clk), .A(\g.we_clk [13834]));
Q_ASSIGN U2557 ( .B(clk), .A(\g.we_clk [13833]));
Q_ASSIGN U2558 ( .B(clk), .A(\g.we_clk [13832]));
Q_ASSIGN U2559 ( .B(clk), .A(\g.we_clk [13831]));
Q_ASSIGN U2560 ( .B(clk), .A(\g.we_clk [13830]));
Q_ASSIGN U2561 ( .B(clk), .A(\g.we_clk [13829]));
Q_ASSIGN U2562 ( .B(clk), .A(\g.we_clk [13828]));
Q_ASSIGN U2563 ( .B(clk), .A(\g.we_clk [13827]));
Q_ASSIGN U2564 ( .B(clk), .A(\g.we_clk [13826]));
Q_ASSIGN U2565 ( .B(clk), .A(\g.we_clk [13825]));
Q_ASSIGN U2566 ( .B(clk), .A(\g.we_clk [13824]));
Q_ASSIGN U2567 ( .B(clk), .A(\g.we_clk [13823]));
Q_ASSIGN U2568 ( .B(clk), .A(\g.we_clk [13822]));
Q_ASSIGN U2569 ( .B(clk), .A(\g.we_clk [13821]));
Q_ASSIGN U2570 ( .B(clk), .A(\g.we_clk [13820]));
Q_ASSIGN U2571 ( .B(clk), .A(\g.we_clk [13819]));
Q_ASSIGN U2572 ( .B(clk), .A(\g.we_clk [13818]));
Q_ASSIGN U2573 ( .B(clk), .A(\g.we_clk [13817]));
Q_ASSIGN U2574 ( .B(clk), .A(\g.we_clk [13816]));
Q_ASSIGN U2575 ( .B(clk), .A(\g.we_clk [13815]));
Q_ASSIGN U2576 ( .B(clk), .A(\g.we_clk [13814]));
Q_ASSIGN U2577 ( .B(clk), .A(\g.we_clk [13813]));
Q_ASSIGN U2578 ( .B(clk), .A(\g.we_clk [13812]));
Q_ASSIGN U2579 ( .B(clk), .A(\g.we_clk [13811]));
Q_ASSIGN U2580 ( .B(clk), .A(\g.we_clk [13810]));
Q_ASSIGN U2581 ( .B(clk), .A(\g.we_clk [13809]));
Q_ASSIGN U2582 ( .B(clk), .A(\g.we_clk [13808]));
Q_ASSIGN U2583 ( .B(clk), .A(\g.we_clk [13807]));
Q_ASSIGN U2584 ( .B(clk), .A(\g.we_clk [13806]));
Q_ASSIGN U2585 ( .B(clk), .A(\g.we_clk [13805]));
Q_ASSIGN U2586 ( .B(clk), .A(\g.we_clk [13804]));
Q_ASSIGN U2587 ( .B(clk), .A(\g.we_clk [13803]));
Q_ASSIGN U2588 ( .B(clk), .A(\g.we_clk [13802]));
Q_ASSIGN U2589 ( .B(clk), .A(\g.we_clk [13801]));
Q_ASSIGN U2590 ( .B(clk), .A(\g.we_clk [13800]));
Q_ASSIGN U2591 ( .B(clk), .A(\g.we_clk [13799]));
Q_ASSIGN U2592 ( .B(clk), .A(\g.we_clk [13798]));
Q_ASSIGN U2593 ( .B(clk), .A(\g.we_clk [13797]));
Q_ASSIGN U2594 ( .B(clk), .A(\g.we_clk [13796]));
Q_ASSIGN U2595 ( .B(clk), .A(\g.we_clk [13795]));
Q_ASSIGN U2596 ( .B(clk), .A(\g.we_clk [13794]));
Q_ASSIGN U2597 ( .B(clk), .A(\g.we_clk [13793]));
Q_ASSIGN U2598 ( .B(clk), .A(\g.we_clk [13792]));
Q_ASSIGN U2599 ( .B(clk), .A(\g.we_clk [13791]));
Q_ASSIGN U2600 ( .B(clk), .A(\g.we_clk [13790]));
Q_ASSIGN U2601 ( .B(clk), .A(\g.we_clk [13789]));
Q_ASSIGN U2602 ( .B(clk), .A(\g.we_clk [13788]));
Q_ASSIGN U2603 ( .B(clk), .A(\g.we_clk [13787]));
Q_ASSIGN U2604 ( .B(clk), .A(\g.we_clk [13786]));
Q_ASSIGN U2605 ( .B(clk), .A(\g.we_clk [13785]));
Q_ASSIGN U2606 ( .B(clk), .A(\g.we_clk [13784]));
Q_ASSIGN U2607 ( .B(clk), .A(\g.we_clk [13783]));
Q_ASSIGN U2608 ( .B(clk), .A(\g.we_clk [13782]));
Q_ASSIGN U2609 ( .B(clk), .A(\g.we_clk [13781]));
Q_ASSIGN U2610 ( .B(clk), .A(\g.we_clk [13780]));
Q_ASSIGN U2611 ( .B(clk), .A(\g.we_clk [13779]));
Q_ASSIGN U2612 ( .B(clk), .A(\g.we_clk [13778]));
Q_ASSIGN U2613 ( .B(clk), .A(\g.we_clk [13777]));
Q_ASSIGN U2614 ( .B(clk), .A(\g.we_clk [13776]));
Q_ASSIGN U2615 ( .B(clk), .A(\g.we_clk [13775]));
Q_ASSIGN U2616 ( .B(clk), .A(\g.we_clk [13774]));
Q_ASSIGN U2617 ( .B(clk), .A(\g.we_clk [13773]));
Q_ASSIGN U2618 ( .B(clk), .A(\g.we_clk [13772]));
Q_ASSIGN U2619 ( .B(clk), .A(\g.we_clk [13771]));
Q_ASSIGN U2620 ( .B(clk), .A(\g.we_clk [13770]));
Q_ASSIGN U2621 ( .B(clk), .A(\g.we_clk [13769]));
Q_ASSIGN U2622 ( .B(clk), .A(\g.we_clk [13768]));
Q_ASSIGN U2623 ( .B(clk), .A(\g.we_clk [13767]));
Q_ASSIGN U2624 ( .B(clk), .A(\g.we_clk [13766]));
Q_ASSIGN U2625 ( .B(clk), .A(\g.we_clk [13765]));
Q_ASSIGN U2626 ( .B(clk), .A(\g.we_clk [13764]));
Q_ASSIGN U2627 ( .B(clk), .A(\g.we_clk [13763]));
Q_ASSIGN U2628 ( .B(clk), .A(\g.we_clk [13762]));
Q_ASSIGN U2629 ( .B(clk), .A(\g.we_clk [13761]));
Q_ASSIGN U2630 ( .B(clk), .A(\g.we_clk [13760]));
Q_ASSIGN U2631 ( .B(clk), .A(\g.we_clk [13759]));
Q_ASSIGN U2632 ( .B(clk), .A(\g.we_clk [13758]));
Q_ASSIGN U2633 ( .B(clk), .A(\g.we_clk [13757]));
Q_ASSIGN U2634 ( .B(clk), .A(\g.we_clk [13756]));
Q_ASSIGN U2635 ( .B(clk), .A(\g.we_clk [13755]));
Q_ASSIGN U2636 ( .B(clk), .A(\g.we_clk [13754]));
Q_ASSIGN U2637 ( .B(clk), .A(\g.we_clk [13753]));
Q_ASSIGN U2638 ( .B(clk), .A(\g.we_clk [13752]));
Q_ASSIGN U2639 ( .B(clk), .A(\g.we_clk [13751]));
Q_ASSIGN U2640 ( .B(clk), .A(\g.we_clk [13750]));
Q_ASSIGN U2641 ( .B(clk), .A(\g.we_clk [13749]));
Q_ASSIGN U2642 ( .B(clk), .A(\g.we_clk [13748]));
Q_ASSIGN U2643 ( .B(clk), .A(\g.we_clk [13747]));
Q_ASSIGN U2644 ( .B(clk), .A(\g.we_clk [13746]));
Q_ASSIGN U2645 ( .B(clk), .A(\g.we_clk [13745]));
Q_ASSIGN U2646 ( .B(clk), .A(\g.we_clk [13744]));
Q_ASSIGN U2647 ( .B(clk), .A(\g.we_clk [13743]));
Q_ASSIGN U2648 ( .B(clk), .A(\g.we_clk [13742]));
Q_ASSIGN U2649 ( .B(clk), .A(\g.we_clk [13741]));
Q_ASSIGN U2650 ( .B(clk), .A(\g.we_clk [13740]));
Q_ASSIGN U2651 ( .B(clk), .A(\g.we_clk [13739]));
Q_ASSIGN U2652 ( .B(clk), .A(\g.we_clk [13738]));
Q_ASSIGN U2653 ( .B(clk), .A(\g.we_clk [13737]));
Q_ASSIGN U2654 ( .B(clk), .A(\g.we_clk [13736]));
Q_ASSIGN U2655 ( .B(clk), .A(\g.we_clk [13735]));
Q_ASSIGN U2656 ( .B(clk), .A(\g.we_clk [13734]));
Q_ASSIGN U2657 ( .B(clk), .A(\g.we_clk [13733]));
Q_ASSIGN U2658 ( .B(clk), .A(\g.we_clk [13732]));
Q_ASSIGN U2659 ( .B(clk), .A(\g.we_clk [13731]));
Q_ASSIGN U2660 ( .B(clk), .A(\g.we_clk [13730]));
Q_ASSIGN U2661 ( .B(clk), .A(\g.we_clk [13729]));
Q_ASSIGN U2662 ( .B(clk), .A(\g.we_clk [13728]));
Q_ASSIGN U2663 ( .B(clk), .A(\g.we_clk [13727]));
Q_ASSIGN U2664 ( .B(clk), .A(\g.we_clk [13726]));
Q_ASSIGN U2665 ( .B(clk), .A(\g.we_clk [13725]));
Q_ASSIGN U2666 ( .B(clk), .A(\g.we_clk [13724]));
Q_ASSIGN U2667 ( .B(clk), .A(\g.we_clk [13723]));
Q_ASSIGN U2668 ( .B(clk), .A(\g.we_clk [13722]));
Q_ASSIGN U2669 ( .B(clk), .A(\g.we_clk [13721]));
Q_ASSIGN U2670 ( .B(clk), .A(\g.we_clk [13720]));
Q_ASSIGN U2671 ( .B(clk), .A(\g.we_clk [13719]));
Q_ASSIGN U2672 ( .B(clk), .A(\g.we_clk [13718]));
Q_ASSIGN U2673 ( .B(clk), .A(\g.we_clk [13717]));
Q_ASSIGN U2674 ( .B(clk), .A(\g.we_clk [13716]));
Q_ASSIGN U2675 ( .B(clk), .A(\g.we_clk [13715]));
Q_ASSIGN U2676 ( .B(clk), .A(\g.we_clk [13714]));
Q_ASSIGN U2677 ( .B(clk), .A(\g.we_clk [13713]));
Q_ASSIGN U2678 ( .B(clk), .A(\g.we_clk [13712]));
Q_ASSIGN U2679 ( .B(clk), .A(\g.we_clk [13711]));
Q_ASSIGN U2680 ( .B(clk), .A(\g.we_clk [13710]));
Q_ASSIGN U2681 ( .B(clk), .A(\g.we_clk [13709]));
Q_ASSIGN U2682 ( .B(clk), .A(\g.we_clk [13708]));
Q_ASSIGN U2683 ( .B(clk), .A(\g.we_clk [13707]));
Q_ASSIGN U2684 ( .B(clk), .A(\g.we_clk [13706]));
Q_ASSIGN U2685 ( .B(clk), .A(\g.we_clk [13705]));
Q_ASSIGN U2686 ( .B(clk), .A(\g.we_clk [13704]));
Q_ASSIGN U2687 ( .B(clk), .A(\g.we_clk [13703]));
Q_ASSIGN U2688 ( .B(clk), .A(\g.we_clk [13702]));
Q_ASSIGN U2689 ( .B(clk), .A(\g.we_clk [13701]));
Q_ASSIGN U2690 ( .B(clk), .A(\g.we_clk [13700]));
Q_ASSIGN U2691 ( .B(clk), .A(\g.we_clk [13699]));
Q_ASSIGN U2692 ( .B(clk), .A(\g.we_clk [13698]));
Q_ASSIGN U2693 ( .B(clk), .A(\g.we_clk [13697]));
Q_ASSIGN U2694 ( .B(clk), .A(\g.we_clk [13696]));
Q_ASSIGN U2695 ( .B(clk), .A(\g.we_clk [13695]));
Q_ASSIGN U2696 ( .B(clk), .A(\g.we_clk [13694]));
Q_ASSIGN U2697 ( .B(clk), .A(\g.we_clk [13693]));
Q_ASSIGN U2698 ( .B(clk), .A(\g.we_clk [13692]));
Q_ASSIGN U2699 ( .B(clk), .A(\g.we_clk [13691]));
Q_ASSIGN U2700 ( .B(clk), .A(\g.we_clk [13690]));
Q_ASSIGN U2701 ( .B(clk), .A(\g.we_clk [13689]));
Q_ASSIGN U2702 ( .B(clk), .A(\g.we_clk [13688]));
Q_ASSIGN U2703 ( .B(clk), .A(\g.we_clk [13687]));
Q_ASSIGN U2704 ( .B(clk), .A(\g.we_clk [13686]));
Q_ASSIGN U2705 ( .B(clk), .A(\g.we_clk [13685]));
Q_ASSIGN U2706 ( .B(clk), .A(\g.we_clk [13684]));
Q_ASSIGN U2707 ( .B(clk), .A(\g.we_clk [13683]));
Q_ASSIGN U2708 ( .B(clk), .A(\g.we_clk [13682]));
Q_ASSIGN U2709 ( .B(clk), .A(\g.we_clk [13681]));
Q_ASSIGN U2710 ( .B(clk), .A(\g.we_clk [13680]));
Q_ASSIGN U2711 ( .B(clk), .A(\g.we_clk [13679]));
Q_ASSIGN U2712 ( .B(clk), .A(\g.we_clk [13678]));
Q_ASSIGN U2713 ( .B(clk), .A(\g.we_clk [13677]));
Q_ASSIGN U2714 ( .B(clk), .A(\g.we_clk [13676]));
Q_ASSIGN U2715 ( .B(clk), .A(\g.we_clk [13675]));
Q_ASSIGN U2716 ( .B(clk), .A(\g.we_clk [13674]));
Q_ASSIGN U2717 ( .B(clk), .A(\g.we_clk [13673]));
Q_ASSIGN U2718 ( .B(clk), .A(\g.we_clk [13672]));
Q_ASSIGN U2719 ( .B(clk), .A(\g.we_clk [13671]));
Q_ASSIGN U2720 ( .B(clk), .A(\g.we_clk [13670]));
Q_ASSIGN U2721 ( .B(clk), .A(\g.we_clk [13669]));
Q_ASSIGN U2722 ( .B(clk), .A(\g.we_clk [13668]));
Q_ASSIGN U2723 ( .B(clk), .A(\g.we_clk [13667]));
Q_ASSIGN U2724 ( .B(clk), .A(\g.we_clk [13666]));
Q_ASSIGN U2725 ( .B(clk), .A(\g.we_clk [13665]));
Q_ASSIGN U2726 ( .B(clk), .A(\g.we_clk [13664]));
Q_ASSIGN U2727 ( .B(clk), .A(\g.we_clk [13663]));
Q_ASSIGN U2728 ( .B(clk), .A(\g.we_clk [13662]));
Q_ASSIGN U2729 ( .B(clk), .A(\g.we_clk [13661]));
Q_ASSIGN U2730 ( .B(clk), .A(\g.we_clk [13660]));
Q_ASSIGN U2731 ( .B(clk), .A(\g.we_clk [13659]));
Q_ASSIGN U2732 ( .B(clk), .A(\g.we_clk [13658]));
Q_ASSIGN U2733 ( .B(clk), .A(\g.we_clk [13657]));
Q_ASSIGN U2734 ( .B(clk), .A(\g.we_clk [13656]));
Q_ASSIGN U2735 ( .B(clk), .A(\g.we_clk [13655]));
Q_ASSIGN U2736 ( .B(clk), .A(\g.we_clk [13654]));
Q_ASSIGN U2737 ( .B(clk), .A(\g.we_clk [13653]));
Q_ASSIGN U2738 ( .B(clk), .A(\g.we_clk [13652]));
Q_ASSIGN U2739 ( .B(clk), .A(\g.we_clk [13651]));
Q_ASSIGN U2740 ( .B(clk), .A(\g.we_clk [13650]));
Q_ASSIGN U2741 ( .B(clk), .A(\g.we_clk [13649]));
Q_ASSIGN U2742 ( .B(clk), .A(\g.we_clk [13648]));
Q_ASSIGN U2743 ( .B(clk), .A(\g.we_clk [13647]));
Q_ASSIGN U2744 ( .B(clk), .A(\g.we_clk [13646]));
Q_ASSIGN U2745 ( .B(clk), .A(\g.we_clk [13645]));
Q_ASSIGN U2746 ( .B(clk), .A(\g.we_clk [13644]));
Q_ASSIGN U2747 ( .B(clk), .A(\g.we_clk [13643]));
Q_ASSIGN U2748 ( .B(clk), .A(\g.we_clk [13642]));
Q_ASSIGN U2749 ( .B(clk), .A(\g.we_clk [13641]));
Q_ASSIGN U2750 ( .B(clk), .A(\g.we_clk [13640]));
Q_ASSIGN U2751 ( .B(clk), .A(\g.we_clk [13639]));
Q_ASSIGN U2752 ( .B(clk), .A(\g.we_clk [13638]));
Q_ASSIGN U2753 ( .B(clk), .A(\g.we_clk [13637]));
Q_ASSIGN U2754 ( .B(clk), .A(\g.we_clk [13636]));
Q_ASSIGN U2755 ( .B(clk), .A(\g.we_clk [13635]));
Q_ASSIGN U2756 ( .B(clk), .A(\g.we_clk [13634]));
Q_ASSIGN U2757 ( .B(clk), .A(\g.we_clk [13633]));
Q_ASSIGN U2758 ( .B(clk), .A(\g.we_clk [13632]));
Q_ASSIGN U2759 ( .B(clk), .A(\g.we_clk [13631]));
Q_ASSIGN U2760 ( .B(clk), .A(\g.we_clk [13630]));
Q_ASSIGN U2761 ( .B(clk), .A(\g.we_clk [13629]));
Q_ASSIGN U2762 ( .B(clk), .A(\g.we_clk [13628]));
Q_ASSIGN U2763 ( .B(clk), .A(\g.we_clk [13627]));
Q_ASSIGN U2764 ( .B(clk), .A(\g.we_clk [13626]));
Q_ASSIGN U2765 ( .B(clk), .A(\g.we_clk [13625]));
Q_ASSIGN U2766 ( .B(clk), .A(\g.we_clk [13624]));
Q_ASSIGN U2767 ( .B(clk), .A(\g.we_clk [13623]));
Q_ASSIGN U2768 ( .B(clk), .A(\g.we_clk [13622]));
Q_ASSIGN U2769 ( .B(clk), .A(\g.we_clk [13621]));
Q_ASSIGN U2770 ( .B(clk), .A(\g.we_clk [13620]));
Q_ASSIGN U2771 ( .B(clk), .A(\g.we_clk [13619]));
Q_ASSIGN U2772 ( .B(clk), .A(\g.we_clk [13618]));
Q_ASSIGN U2773 ( .B(clk), .A(\g.we_clk [13617]));
Q_ASSIGN U2774 ( .B(clk), .A(\g.we_clk [13616]));
Q_ASSIGN U2775 ( .B(clk), .A(\g.we_clk [13615]));
Q_ASSIGN U2776 ( .B(clk), .A(\g.we_clk [13614]));
Q_ASSIGN U2777 ( .B(clk), .A(\g.we_clk [13613]));
Q_ASSIGN U2778 ( .B(clk), .A(\g.we_clk [13612]));
Q_ASSIGN U2779 ( .B(clk), .A(\g.we_clk [13611]));
Q_ASSIGN U2780 ( .B(clk), .A(\g.we_clk [13610]));
Q_ASSIGN U2781 ( .B(clk), .A(\g.we_clk [13609]));
Q_ASSIGN U2782 ( .B(clk), .A(\g.we_clk [13608]));
Q_ASSIGN U2783 ( .B(clk), .A(\g.we_clk [13607]));
Q_ASSIGN U2784 ( .B(clk), .A(\g.we_clk [13606]));
Q_ASSIGN U2785 ( .B(clk), .A(\g.we_clk [13605]));
Q_ASSIGN U2786 ( .B(clk), .A(\g.we_clk [13604]));
Q_ASSIGN U2787 ( .B(clk), .A(\g.we_clk [13603]));
Q_ASSIGN U2788 ( .B(clk), .A(\g.we_clk [13602]));
Q_ASSIGN U2789 ( .B(clk), .A(\g.we_clk [13601]));
Q_ASSIGN U2790 ( .B(clk), .A(\g.we_clk [13600]));
Q_ASSIGN U2791 ( .B(clk), .A(\g.we_clk [13599]));
Q_ASSIGN U2792 ( .B(clk), .A(\g.we_clk [13598]));
Q_ASSIGN U2793 ( .B(clk), .A(\g.we_clk [13597]));
Q_ASSIGN U2794 ( .B(clk), .A(\g.we_clk [13596]));
Q_ASSIGN U2795 ( .B(clk), .A(\g.we_clk [13595]));
Q_ASSIGN U2796 ( .B(clk), .A(\g.we_clk [13594]));
Q_ASSIGN U2797 ( .B(clk), .A(\g.we_clk [13593]));
Q_ASSIGN U2798 ( .B(clk), .A(\g.we_clk [13592]));
Q_ASSIGN U2799 ( .B(clk), .A(\g.we_clk [13591]));
Q_ASSIGN U2800 ( .B(clk), .A(\g.we_clk [13590]));
Q_ASSIGN U2801 ( .B(clk), .A(\g.we_clk [13589]));
Q_ASSIGN U2802 ( .B(clk), .A(\g.we_clk [13588]));
Q_ASSIGN U2803 ( .B(clk), .A(\g.we_clk [13587]));
Q_ASSIGN U2804 ( .B(clk), .A(\g.we_clk [13586]));
Q_ASSIGN U2805 ( .B(clk), .A(\g.we_clk [13585]));
Q_ASSIGN U2806 ( .B(clk), .A(\g.we_clk [13584]));
Q_ASSIGN U2807 ( .B(clk), .A(\g.we_clk [13583]));
Q_ASSIGN U2808 ( .B(clk), .A(\g.we_clk [13582]));
Q_ASSIGN U2809 ( .B(clk), .A(\g.we_clk [13581]));
Q_ASSIGN U2810 ( .B(clk), .A(\g.we_clk [13580]));
Q_ASSIGN U2811 ( .B(clk), .A(\g.we_clk [13579]));
Q_ASSIGN U2812 ( .B(clk), .A(\g.we_clk [13578]));
Q_ASSIGN U2813 ( .B(clk), .A(\g.we_clk [13577]));
Q_ASSIGN U2814 ( .B(clk), .A(\g.we_clk [13576]));
Q_ASSIGN U2815 ( .B(clk), .A(\g.we_clk [13575]));
Q_ASSIGN U2816 ( .B(clk), .A(\g.we_clk [13574]));
Q_ASSIGN U2817 ( .B(clk), .A(\g.we_clk [13573]));
Q_ASSIGN U2818 ( .B(clk), .A(\g.we_clk [13572]));
Q_ASSIGN U2819 ( .B(clk), .A(\g.we_clk [13571]));
Q_ASSIGN U2820 ( .B(clk), .A(\g.we_clk [13570]));
Q_ASSIGN U2821 ( .B(clk), .A(\g.we_clk [13569]));
Q_ASSIGN U2822 ( .B(clk), .A(\g.we_clk [13568]));
Q_ASSIGN U2823 ( .B(clk), .A(\g.we_clk [13567]));
Q_ASSIGN U2824 ( .B(clk), .A(\g.we_clk [13566]));
Q_ASSIGN U2825 ( .B(clk), .A(\g.we_clk [13565]));
Q_ASSIGN U2826 ( .B(clk), .A(\g.we_clk [13564]));
Q_ASSIGN U2827 ( .B(clk), .A(\g.we_clk [13563]));
Q_ASSIGN U2828 ( .B(clk), .A(\g.we_clk [13562]));
Q_ASSIGN U2829 ( .B(clk), .A(\g.we_clk [13561]));
Q_ASSIGN U2830 ( .B(clk), .A(\g.we_clk [13560]));
Q_ASSIGN U2831 ( .B(clk), .A(\g.we_clk [13559]));
Q_ASSIGN U2832 ( .B(clk), .A(\g.we_clk [13558]));
Q_ASSIGN U2833 ( .B(clk), .A(\g.we_clk [13557]));
Q_ASSIGN U2834 ( .B(clk), .A(\g.we_clk [13556]));
Q_ASSIGN U2835 ( .B(clk), .A(\g.we_clk [13555]));
Q_ASSIGN U2836 ( .B(clk), .A(\g.we_clk [13554]));
Q_ASSIGN U2837 ( .B(clk), .A(\g.we_clk [13553]));
Q_ASSIGN U2838 ( .B(clk), .A(\g.we_clk [13552]));
Q_ASSIGN U2839 ( .B(clk), .A(\g.we_clk [13551]));
Q_ASSIGN U2840 ( .B(clk), .A(\g.we_clk [13550]));
Q_ASSIGN U2841 ( .B(clk), .A(\g.we_clk [13549]));
Q_ASSIGN U2842 ( .B(clk), .A(\g.we_clk [13548]));
Q_ASSIGN U2843 ( .B(clk), .A(\g.we_clk [13547]));
Q_ASSIGN U2844 ( .B(clk), .A(\g.we_clk [13546]));
Q_ASSIGN U2845 ( .B(clk), .A(\g.we_clk [13545]));
Q_ASSIGN U2846 ( .B(clk), .A(\g.we_clk [13544]));
Q_ASSIGN U2847 ( .B(clk), .A(\g.we_clk [13543]));
Q_ASSIGN U2848 ( .B(clk), .A(\g.we_clk [13542]));
Q_ASSIGN U2849 ( .B(clk), .A(\g.we_clk [13541]));
Q_ASSIGN U2850 ( .B(clk), .A(\g.we_clk [13540]));
Q_ASSIGN U2851 ( .B(clk), .A(\g.we_clk [13539]));
Q_ASSIGN U2852 ( .B(clk), .A(\g.we_clk [13538]));
Q_ASSIGN U2853 ( .B(clk), .A(\g.we_clk [13537]));
Q_ASSIGN U2854 ( .B(clk), .A(\g.we_clk [13536]));
Q_ASSIGN U2855 ( .B(clk), .A(\g.we_clk [13535]));
Q_ASSIGN U2856 ( .B(clk), .A(\g.we_clk [13534]));
Q_ASSIGN U2857 ( .B(clk), .A(\g.we_clk [13533]));
Q_ASSIGN U2858 ( .B(clk), .A(\g.we_clk [13532]));
Q_ASSIGN U2859 ( .B(clk), .A(\g.we_clk [13531]));
Q_ASSIGN U2860 ( .B(clk), .A(\g.we_clk [13530]));
Q_ASSIGN U2861 ( .B(clk), .A(\g.we_clk [13529]));
Q_ASSIGN U2862 ( .B(clk), .A(\g.we_clk [13528]));
Q_ASSIGN U2863 ( .B(clk), .A(\g.we_clk [13527]));
Q_ASSIGN U2864 ( .B(clk), .A(\g.we_clk [13526]));
Q_ASSIGN U2865 ( .B(clk), .A(\g.we_clk [13525]));
Q_ASSIGN U2866 ( .B(clk), .A(\g.we_clk [13524]));
Q_ASSIGN U2867 ( .B(clk), .A(\g.we_clk [13523]));
Q_ASSIGN U2868 ( .B(clk), .A(\g.we_clk [13522]));
Q_ASSIGN U2869 ( .B(clk), .A(\g.we_clk [13521]));
Q_ASSIGN U2870 ( .B(clk), .A(\g.we_clk [13520]));
Q_ASSIGN U2871 ( .B(clk), .A(\g.we_clk [13519]));
Q_ASSIGN U2872 ( .B(clk), .A(\g.we_clk [13518]));
Q_ASSIGN U2873 ( .B(clk), .A(\g.we_clk [13517]));
Q_ASSIGN U2874 ( .B(clk), .A(\g.we_clk [13516]));
Q_ASSIGN U2875 ( .B(clk), .A(\g.we_clk [13515]));
Q_ASSIGN U2876 ( .B(clk), .A(\g.we_clk [13514]));
Q_ASSIGN U2877 ( .B(clk), .A(\g.we_clk [13513]));
Q_ASSIGN U2878 ( .B(clk), .A(\g.we_clk [13512]));
Q_ASSIGN U2879 ( .B(clk), .A(\g.we_clk [13511]));
Q_ASSIGN U2880 ( .B(clk), .A(\g.we_clk [13510]));
Q_ASSIGN U2881 ( .B(clk), .A(\g.we_clk [13509]));
Q_ASSIGN U2882 ( .B(clk), .A(\g.we_clk [13508]));
Q_ASSIGN U2883 ( .B(clk), .A(\g.we_clk [13507]));
Q_ASSIGN U2884 ( .B(clk), .A(\g.we_clk [13506]));
Q_ASSIGN U2885 ( .B(clk), .A(\g.we_clk [13505]));
Q_ASSIGN U2886 ( .B(clk), .A(\g.we_clk [13504]));
Q_ASSIGN U2887 ( .B(clk), .A(\g.we_clk [13503]));
Q_ASSIGN U2888 ( .B(clk), .A(\g.we_clk [13502]));
Q_ASSIGN U2889 ( .B(clk), .A(\g.we_clk [13501]));
Q_ASSIGN U2890 ( .B(clk), .A(\g.we_clk [13500]));
Q_ASSIGN U2891 ( .B(clk), .A(\g.we_clk [13499]));
Q_ASSIGN U2892 ( .B(clk), .A(\g.we_clk [13498]));
Q_ASSIGN U2893 ( .B(clk), .A(\g.we_clk [13497]));
Q_ASSIGN U2894 ( .B(clk), .A(\g.we_clk [13496]));
Q_ASSIGN U2895 ( .B(clk), .A(\g.we_clk [13495]));
Q_ASSIGN U2896 ( .B(clk), .A(\g.we_clk [13494]));
Q_ASSIGN U2897 ( .B(clk), .A(\g.we_clk [13493]));
Q_ASSIGN U2898 ( .B(clk), .A(\g.we_clk [13492]));
Q_ASSIGN U2899 ( .B(clk), .A(\g.we_clk [13491]));
Q_ASSIGN U2900 ( .B(clk), .A(\g.we_clk [13490]));
Q_ASSIGN U2901 ( .B(clk), .A(\g.we_clk [13489]));
Q_ASSIGN U2902 ( .B(clk), .A(\g.we_clk [13488]));
Q_ASSIGN U2903 ( .B(clk), .A(\g.we_clk [13487]));
Q_ASSIGN U2904 ( .B(clk), .A(\g.we_clk [13486]));
Q_ASSIGN U2905 ( .B(clk), .A(\g.we_clk [13485]));
Q_ASSIGN U2906 ( .B(clk), .A(\g.we_clk [13484]));
Q_ASSIGN U2907 ( .B(clk), .A(\g.we_clk [13483]));
Q_ASSIGN U2908 ( .B(clk), .A(\g.we_clk [13482]));
Q_ASSIGN U2909 ( .B(clk), .A(\g.we_clk [13481]));
Q_ASSIGN U2910 ( .B(clk), .A(\g.we_clk [13480]));
Q_ASSIGN U2911 ( .B(clk), .A(\g.we_clk [13479]));
Q_ASSIGN U2912 ( .B(clk), .A(\g.we_clk [13478]));
Q_ASSIGN U2913 ( .B(clk), .A(\g.we_clk [13477]));
Q_ASSIGN U2914 ( .B(clk), .A(\g.we_clk [13476]));
Q_ASSIGN U2915 ( .B(clk), .A(\g.we_clk [13475]));
Q_ASSIGN U2916 ( .B(clk), .A(\g.we_clk [13474]));
Q_ASSIGN U2917 ( .B(clk), .A(\g.we_clk [13473]));
Q_ASSIGN U2918 ( .B(clk), .A(\g.we_clk [13472]));
Q_ASSIGN U2919 ( .B(clk), .A(\g.we_clk [13471]));
Q_ASSIGN U2920 ( .B(clk), .A(\g.we_clk [13470]));
Q_ASSIGN U2921 ( .B(clk), .A(\g.we_clk [13469]));
Q_ASSIGN U2922 ( .B(clk), .A(\g.we_clk [13468]));
Q_ASSIGN U2923 ( .B(clk), .A(\g.we_clk [13467]));
Q_ASSIGN U2924 ( .B(clk), .A(\g.we_clk [13466]));
Q_ASSIGN U2925 ( .B(clk), .A(\g.we_clk [13465]));
Q_ASSIGN U2926 ( .B(clk), .A(\g.we_clk [13464]));
Q_ASSIGN U2927 ( .B(clk), .A(\g.we_clk [13463]));
Q_ASSIGN U2928 ( .B(clk), .A(\g.we_clk [13462]));
Q_ASSIGN U2929 ( .B(clk), .A(\g.we_clk [13461]));
Q_ASSIGN U2930 ( .B(clk), .A(\g.we_clk [13460]));
Q_ASSIGN U2931 ( .B(clk), .A(\g.we_clk [13459]));
Q_ASSIGN U2932 ( .B(clk), .A(\g.we_clk [13458]));
Q_ASSIGN U2933 ( .B(clk), .A(\g.we_clk [13457]));
Q_ASSIGN U2934 ( .B(clk), .A(\g.we_clk [13456]));
Q_ASSIGN U2935 ( .B(clk), .A(\g.we_clk [13455]));
Q_ASSIGN U2936 ( .B(clk), .A(\g.we_clk [13454]));
Q_ASSIGN U2937 ( .B(clk), .A(\g.we_clk [13453]));
Q_ASSIGN U2938 ( .B(clk), .A(\g.we_clk [13452]));
Q_ASSIGN U2939 ( .B(clk), .A(\g.we_clk [13451]));
Q_ASSIGN U2940 ( .B(clk), .A(\g.we_clk [13450]));
Q_ASSIGN U2941 ( .B(clk), .A(\g.we_clk [13449]));
Q_ASSIGN U2942 ( .B(clk), .A(\g.we_clk [13448]));
Q_ASSIGN U2943 ( .B(clk), .A(\g.we_clk [13447]));
Q_ASSIGN U2944 ( .B(clk), .A(\g.we_clk [13446]));
Q_ASSIGN U2945 ( .B(clk), .A(\g.we_clk [13445]));
Q_ASSIGN U2946 ( .B(clk), .A(\g.we_clk [13444]));
Q_ASSIGN U2947 ( .B(clk), .A(\g.we_clk [13443]));
Q_ASSIGN U2948 ( .B(clk), .A(\g.we_clk [13442]));
Q_ASSIGN U2949 ( .B(clk), .A(\g.we_clk [13441]));
Q_ASSIGN U2950 ( .B(clk), .A(\g.we_clk [13440]));
Q_ASSIGN U2951 ( .B(clk), .A(\g.we_clk [13439]));
Q_ASSIGN U2952 ( .B(clk), .A(\g.we_clk [13438]));
Q_ASSIGN U2953 ( .B(clk), .A(\g.we_clk [13437]));
Q_ASSIGN U2954 ( .B(clk), .A(\g.we_clk [13436]));
Q_ASSIGN U2955 ( .B(clk), .A(\g.we_clk [13435]));
Q_ASSIGN U2956 ( .B(clk), .A(\g.we_clk [13434]));
Q_ASSIGN U2957 ( .B(clk), .A(\g.we_clk [13433]));
Q_ASSIGN U2958 ( .B(clk), .A(\g.we_clk [13432]));
Q_ASSIGN U2959 ( .B(clk), .A(\g.we_clk [13431]));
Q_ASSIGN U2960 ( .B(clk), .A(\g.we_clk [13430]));
Q_ASSIGN U2961 ( .B(clk), .A(\g.we_clk [13429]));
Q_ASSIGN U2962 ( .B(clk), .A(\g.we_clk [13428]));
Q_ASSIGN U2963 ( .B(clk), .A(\g.we_clk [13427]));
Q_ASSIGN U2964 ( .B(clk), .A(\g.we_clk [13426]));
Q_ASSIGN U2965 ( .B(clk), .A(\g.we_clk [13425]));
Q_ASSIGN U2966 ( .B(clk), .A(\g.we_clk [13424]));
Q_ASSIGN U2967 ( .B(clk), .A(\g.we_clk [13423]));
Q_ASSIGN U2968 ( .B(clk), .A(\g.we_clk [13422]));
Q_ASSIGN U2969 ( .B(clk), .A(\g.we_clk [13421]));
Q_ASSIGN U2970 ( .B(clk), .A(\g.we_clk [13420]));
Q_ASSIGN U2971 ( .B(clk), .A(\g.we_clk [13419]));
Q_ASSIGN U2972 ( .B(clk), .A(\g.we_clk [13418]));
Q_ASSIGN U2973 ( .B(clk), .A(\g.we_clk [13417]));
Q_ASSIGN U2974 ( .B(clk), .A(\g.we_clk [13416]));
Q_ASSIGN U2975 ( .B(clk), .A(\g.we_clk [13415]));
Q_ASSIGN U2976 ( .B(clk), .A(\g.we_clk [13414]));
Q_ASSIGN U2977 ( .B(clk), .A(\g.we_clk [13413]));
Q_ASSIGN U2978 ( .B(clk), .A(\g.we_clk [13412]));
Q_ASSIGN U2979 ( .B(clk), .A(\g.we_clk [13411]));
Q_ASSIGN U2980 ( .B(clk), .A(\g.we_clk [13410]));
Q_ASSIGN U2981 ( .B(clk), .A(\g.we_clk [13409]));
Q_ASSIGN U2982 ( .B(clk), .A(\g.we_clk [13408]));
Q_ASSIGN U2983 ( .B(clk), .A(\g.we_clk [13407]));
Q_ASSIGN U2984 ( .B(clk), .A(\g.we_clk [13406]));
Q_ASSIGN U2985 ( .B(clk), .A(\g.we_clk [13405]));
Q_ASSIGN U2986 ( .B(clk), .A(\g.we_clk [13404]));
Q_ASSIGN U2987 ( .B(clk), .A(\g.we_clk [13403]));
Q_ASSIGN U2988 ( .B(clk), .A(\g.we_clk [13402]));
Q_ASSIGN U2989 ( .B(clk), .A(\g.we_clk [13401]));
Q_ASSIGN U2990 ( .B(clk), .A(\g.we_clk [13400]));
Q_ASSIGN U2991 ( .B(clk), .A(\g.we_clk [13399]));
Q_ASSIGN U2992 ( .B(clk), .A(\g.we_clk [13398]));
Q_ASSIGN U2993 ( .B(clk), .A(\g.we_clk [13397]));
Q_ASSIGN U2994 ( .B(clk), .A(\g.we_clk [13396]));
Q_ASSIGN U2995 ( .B(clk), .A(\g.we_clk [13395]));
Q_ASSIGN U2996 ( .B(clk), .A(\g.we_clk [13394]));
Q_ASSIGN U2997 ( .B(clk), .A(\g.we_clk [13393]));
Q_ASSIGN U2998 ( .B(clk), .A(\g.we_clk [13392]));
Q_ASSIGN U2999 ( .B(clk), .A(\g.we_clk [13391]));
Q_ASSIGN U3000 ( .B(clk), .A(\g.we_clk [13390]));
Q_ASSIGN U3001 ( .B(clk), .A(\g.we_clk [13389]));
Q_ASSIGN U3002 ( .B(clk), .A(\g.we_clk [13388]));
Q_ASSIGN U3003 ( .B(clk), .A(\g.we_clk [13387]));
Q_ASSIGN U3004 ( .B(clk), .A(\g.we_clk [13386]));
Q_ASSIGN U3005 ( .B(clk), .A(\g.we_clk [13385]));
Q_ASSIGN U3006 ( .B(clk), .A(\g.we_clk [13384]));
Q_ASSIGN U3007 ( .B(clk), .A(\g.we_clk [13383]));
Q_ASSIGN U3008 ( .B(clk), .A(\g.we_clk [13382]));
Q_ASSIGN U3009 ( .B(clk), .A(\g.we_clk [13381]));
Q_ASSIGN U3010 ( .B(clk), .A(\g.we_clk [13380]));
Q_ASSIGN U3011 ( .B(clk), .A(\g.we_clk [13379]));
Q_ASSIGN U3012 ( .B(clk), .A(\g.we_clk [13378]));
Q_ASSIGN U3013 ( .B(clk), .A(\g.we_clk [13377]));
Q_ASSIGN U3014 ( .B(clk), .A(\g.we_clk [13376]));
Q_ASSIGN U3015 ( .B(clk), .A(\g.we_clk [13375]));
Q_ASSIGN U3016 ( .B(clk), .A(\g.we_clk [13374]));
Q_ASSIGN U3017 ( .B(clk), .A(\g.we_clk [13373]));
Q_ASSIGN U3018 ( .B(clk), .A(\g.we_clk [13372]));
Q_ASSIGN U3019 ( .B(clk), .A(\g.we_clk [13371]));
Q_ASSIGN U3020 ( .B(clk), .A(\g.we_clk [13370]));
Q_ASSIGN U3021 ( .B(clk), .A(\g.we_clk [13369]));
Q_ASSIGN U3022 ( .B(clk), .A(\g.we_clk [13368]));
Q_ASSIGN U3023 ( .B(clk), .A(\g.we_clk [13367]));
Q_ASSIGN U3024 ( .B(clk), .A(\g.we_clk [13366]));
Q_ASSIGN U3025 ( .B(clk), .A(\g.we_clk [13365]));
Q_ASSIGN U3026 ( .B(clk), .A(\g.we_clk [13364]));
Q_ASSIGN U3027 ( .B(clk), .A(\g.we_clk [13363]));
Q_ASSIGN U3028 ( .B(clk), .A(\g.we_clk [13362]));
Q_ASSIGN U3029 ( .B(clk), .A(\g.we_clk [13361]));
Q_ASSIGN U3030 ( .B(clk), .A(\g.we_clk [13360]));
Q_ASSIGN U3031 ( .B(clk), .A(\g.we_clk [13359]));
Q_ASSIGN U3032 ( .B(clk), .A(\g.we_clk [13358]));
Q_ASSIGN U3033 ( .B(clk), .A(\g.we_clk [13357]));
Q_ASSIGN U3034 ( .B(clk), .A(\g.we_clk [13356]));
Q_ASSIGN U3035 ( .B(clk), .A(\g.we_clk [13355]));
Q_ASSIGN U3036 ( .B(clk), .A(\g.we_clk [13354]));
Q_ASSIGN U3037 ( .B(clk), .A(\g.we_clk [13353]));
Q_ASSIGN U3038 ( .B(clk), .A(\g.we_clk [13352]));
Q_ASSIGN U3039 ( .B(clk), .A(\g.we_clk [13351]));
Q_ASSIGN U3040 ( .B(clk), .A(\g.we_clk [13350]));
Q_ASSIGN U3041 ( .B(clk), .A(\g.we_clk [13349]));
Q_ASSIGN U3042 ( .B(clk), .A(\g.we_clk [13348]));
Q_ASSIGN U3043 ( .B(clk), .A(\g.we_clk [13347]));
Q_ASSIGN U3044 ( .B(clk), .A(\g.we_clk [13346]));
Q_ASSIGN U3045 ( .B(clk), .A(\g.we_clk [13345]));
Q_ASSIGN U3046 ( .B(clk), .A(\g.we_clk [13344]));
Q_ASSIGN U3047 ( .B(clk), .A(\g.we_clk [13343]));
Q_ASSIGN U3048 ( .B(clk), .A(\g.we_clk [13342]));
Q_ASSIGN U3049 ( .B(clk), .A(\g.we_clk [13341]));
Q_ASSIGN U3050 ( .B(clk), .A(\g.we_clk [13340]));
Q_ASSIGN U3051 ( .B(clk), .A(\g.we_clk [13339]));
Q_ASSIGN U3052 ( .B(clk), .A(\g.we_clk [13338]));
Q_ASSIGN U3053 ( .B(clk), .A(\g.we_clk [13337]));
Q_ASSIGN U3054 ( .B(clk), .A(\g.we_clk [13336]));
Q_ASSIGN U3055 ( .B(clk), .A(\g.we_clk [13335]));
Q_ASSIGN U3056 ( .B(clk), .A(\g.we_clk [13334]));
Q_ASSIGN U3057 ( .B(clk), .A(\g.we_clk [13333]));
Q_ASSIGN U3058 ( .B(clk), .A(\g.we_clk [13332]));
Q_ASSIGN U3059 ( .B(clk), .A(\g.we_clk [13331]));
Q_ASSIGN U3060 ( .B(clk), .A(\g.we_clk [13330]));
Q_ASSIGN U3061 ( .B(clk), .A(\g.we_clk [13329]));
Q_ASSIGN U3062 ( .B(clk), .A(\g.we_clk [13328]));
Q_ASSIGN U3063 ( .B(clk), .A(\g.we_clk [13327]));
Q_ASSIGN U3064 ( .B(clk), .A(\g.we_clk [13326]));
Q_ASSIGN U3065 ( .B(clk), .A(\g.we_clk [13325]));
Q_ASSIGN U3066 ( .B(clk), .A(\g.we_clk [13324]));
Q_ASSIGN U3067 ( .B(clk), .A(\g.we_clk [13323]));
Q_ASSIGN U3068 ( .B(clk), .A(\g.we_clk [13322]));
Q_ASSIGN U3069 ( .B(clk), .A(\g.we_clk [13321]));
Q_ASSIGN U3070 ( .B(clk), .A(\g.we_clk [13320]));
Q_ASSIGN U3071 ( .B(clk), .A(\g.we_clk [13319]));
Q_ASSIGN U3072 ( .B(clk), .A(\g.we_clk [13318]));
Q_ASSIGN U3073 ( .B(clk), .A(\g.we_clk [13317]));
Q_ASSIGN U3074 ( .B(clk), .A(\g.we_clk [13316]));
Q_ASSIGN U3075 ( .B(clk), .A(\g.we_clk [13315]));
Q_ASSIGN U3076 ( .B(clk), .A(\g.we_clk [13314]));
Q_ASSIGN U3077 ( .B(clk), .A(\g.we_clk [13313]));
Q_ASSIGN U3078 ( .B(clk), .A(\g.we_clk [13312]));
Q_ASSIGN U3079 ( .B(clk), .A(\g.we_clk [13311]));
Q_ASSIGN U3080 ( .B(clk), .A(\g.we_clk [13310]));
Q_ASSIGN U3081 ( .B(clk), .A(\g.we_clk [13309]));
Q_ASSIGN U3082 ( .B(clk), .A(\g.we_clk [13308]));
Q_ASSIGN U3083 ( .B(clk), .A(\g.we_clk [13307]));
Q_ASSIGN U3084 ( .B(clk), .A(\g.we_clk [13306]));
Q_ASSIGN U3085 ( .B(clk), .A(\g.we_clk [13305]));
Q_ASSIGN U3086 ( .B(clk), .A(\g.we_clk [13304]));
Q_ASSIGN U3087 ( .B(clk), .A(\g.we_clk [13303]));
Q_ASSIGN U3088 ( .B(clk), .A(\g.we_clk [13302]));
Q_ASSIGN U3089 ( .B(clk), .A(\g.we_clk [13301]));
Q_ASSIGN U3090 ( .B(clk), .A(\g.we_clk [13300]));
Q_ASSIGN U3091 ( .B(clk), .A(\g.we_clk [13299]));
Q_ASSIGN U3092 ( .B(clk), .A(\g.we_clk [13298]));
Q_ASSIGN U3093 ( .B(clk), .A(\g.we_clk [13297]));
Q_ASSIGN U3094 ( .B(clk), .A(\g.we_clk [13296]));
Q_ASSIGN U3095 ( .B(clk), .A(\g.we_clk [13295]));
Q_ASSIGN U3096 ( .B(clk), .A(\g.we_clk [13294]));
Q_ASSIGN U3097 ( .B(clk), .A(\g.we_clk [13293]));
Q_ASSIGN U3098 ( .B(clk), .A(\g.we_clk [13292]));
Q_ASSIGN U3099 ( .B(clk), .A(\g.we_clk [13291]));
Q_ASSIGN U3100 ( .B(clk), .A(\g.we_clk [13290]));
Q_ASSIGN U3101 ( .B(clk), .A(\g.we_clk [13289]));
Q_ASSIGN U3102 ( .B(clk), .A(\g.we_clk [13288]));
Q_ASSIGN U3103 ( .B(clk), .A(\g.we_clk [13287]));
Q_ASSIGN U3104 ( .B(clk), .A(\g.we_clk [13286]));
Q_ASSIGN U3105 ( .B(clk), .A(\g.we_clk [13285]));
Q_ASSIGN U3106 ( .B(clk), .A(\g.we_clk [13284]));
Q_ASSIGN U3107 ( .B(clk), .A(\g.we_clk [13283]));
Q_ASSIGN U3108 ( .B(clk), .A(\g.we_clk [13282]));
Q_ASSIGN U3109 ( .B(clk), .A(\g.we_clk [13281]));
Q_ASSIGN U3110 ( .B(clk), .A(\g.we_clk [13280]));
Q_ASSIGN U3111 ( .B(clk), .A(\g.we_clk [13279]));
Q_ASSIGN U3112 ( .B(clk), .A(\g.we_clk [13278]));
Q_ASSIGN U3113 ( .B(clk), .A(\g.we_clk [13277]));
Q_ASSIGN U3114 ( .B(clk), .A(\g.we_clk [13276]));
Q_ASSIGN U3115 ( .B(clk), .A(\g.we_clk [13275]));
Q_ASSIGN U3116 ( .B(clk), .A(\g.we_clk [13274]));
Q_ASSIGN U3117 ( .B(clk), .A(\g.we_clk [13273]));
Q_ASSIGN U3118 ( .B(clk), .A(\g.we_clk [13272]));
Q_ASSIGN U3119 ( .B(clk), .A(\g.we_clk [13271]));
Q_ASSIGN U3120 ( .B(clk), .A(\g.we_clk [13270]));
Q_ASSIGN U3121 ( .B(clk), .A(\g.we_clk [13269]));
Q_ASSIGN U3122 ( .B(clk), .A(\g.we_clk [13268]));
Q_ASSIGN U3123 ( .B(clk), .A(\g.we_clk [13267]));
Q_ASSIGN U3124 ( .B(clk), .A(\g.we_clk [13266]));
Q_ASSIGN U3125 ( .B(clk), .A(\g.we_clk [13265]));
Q_ASSIGN U3126 ( .B(clk), .A(\g.we_clk [13264]));
Q_ASSIGN U3127 ( .B(clk), .A(\g.we_clk [13263]));
Q_ASSIGN U3128 ( .B(clk), .A(\g.we_clk [13262]));
Q_ASSIGN U3129 ( .B(clk), .A(\g.we_clk [13261]));
Q_ASSIGN U3130 ( .B(clk), .A(\g.we_clk [13260]));
Q_ASSIGN U3131 ( .B(clk), .A(\g.we_clk [13259]));
Q_ASSIGN U3132 ( .B(clk), .A(\g.we_clk [13258]));
Q_ASSIGN U3133 ( .B(clk), .A(\g.we_clk [13257]));
Q_ASSIGN U3134 ( .B(clk), .A(\g.we_clk [13256]));
Q_ASSIGN U3135 ( .B(clk), .A(\g.we_clk [13255]));
Q_ASSIGN U3136 ( .B(clk), .A(\g.we_clk [13254]));
Q_ASSIGN U3137 ( .B(clk), .A(\g.we_clk [13253]));
Q_ASSIGN U3138 ( .B(clk), .A(\g.we_clk [13252]));
Q_ASSIGN U3139 ( .B(clk), .A(\g.we_clk [13251]));
Q_ASSIGN U3140 ( .B(clk), .A(\g.we_clk [13250]));
Q_ASSIGN U3141 ( .B(clk), .A(\g.we_clk [13249]));
Q_ASSIGN U3142 ( .B(clk), .A(\g.we_clk [13248]));
Q_ASSIGN U3143 ( .B(clk), .A(\g.we_clk [13247]));
Q_ASSIGN U3144 ( .B(clk), .A(\g.we_clk [13246]));
Q_ASSIGN U3145 ( .B(clk), .A(\g.we_clk [13245]));
Q_ASSIGN U3146 ( .B(clk), .A(\g.we_clk [13244]));
Q_ASSIGN U3147 ( .B(clk), .A(\g.we_clk [13243]));
Q_ASSIGN U3148 ( .B(clk), .A(\g.we_clk [13242]));
Q_ASSIGN U3149 ( .B(clk), .A(\g.we_clk [13241]));
Q_ASSIGN U3150 ( .B(clk), .A(\g.we_clk [13240]));
Q_ASSIGN U3151 ( .B(clk), .A(\g.we_clk [13239]));
Q_ASSIGN U3152 ( .B(clk), .A(\g.we_clk [13238]));
Q_ASSIGN U3153 ( .B(clk), .A(\g.we_clk [13237]));
Q_ASSIGN U3154 ( .B(clk), .A(\g.we_clk [13236]));
Q_ASSIGN U3155 ( .B(clk), .A(\g.we_clk [13235]));
Q_ASSIGN U3156 ( .B(clk), .A(\g.we_clk [13234]));
Q_ASSIGN U3157 ( .B(clk), .A(\g.we_clk [13233]));
Q_ASSIGN U3158 ( .B(clk), .A(\g.we_clk [13232]));
Q_ASSIGN U3159 ( .B(clk), .A(\g.we_clk [13231]));
Q_ASSIGN U3160 ( .B(clk), .A(\g.we_clk [13230]));
Q_ASSIGN U3161 ( .B(clk), .A(\g.we_clk [13229]));
Q_ASSIGN U3162 ( .B(clk), .A(\g.we_clk [13228]));
Q_ASSIGN U3163 ( .B(clk), .A(\g.we_clk [13227]));
Q_ASSIGN U3164 ( .B(clk), .A(\g.we_clk [13226]));
Q_ASSIGN U3165 ( .B(clk), .A(\g.we_clk [13225]));
Q_ASSIGN U3166 ( .B(clk), .A(\g.we_clk [13224]));
Q_ASSIGN U3167 ( .B(clk), .A(\g.we_clk [13223]));
Q_ASSIGN U3168 ( .B(clk), .A(\g.we_clk [13222]));
Q_ASSIGN U3169 ( .B(clk), .A(\g.we_clk [13221]));
Q_ASSIGN U3170 ( .B(clk), .A(\g.we_clk [13220]));
Q_ASSIGN U3171 ( .B(clk), .A(\g.we_clk [13219]));
Q_ASSIGN U3172 ( .B(clk), .A(\g.we_clk [13218]));
Q_ASSIGN U3173 ( .B(clk), .A(\g.we_clk [13217]));
Q_ASSIGN U3174 ( .B(clk), .A(\g.we_clk [13216]));
Q_ASSIGN U3175 ( .B(clk), .A(\g.we_clk [13215]));
Q_ASSIGN U3176 ( .B(clk), .A(\g.we_clk [13214]));
Q_ASSIGN U3177 ( .B(clk), .A(\g.we_clk [13213]));
Q_ASSIGN U3178 ( .B(clk), .A(\g.we_clk [13212]));
Q_ASSIGN U3179 ( .B(clk), .A(\g.we_clk [13211]));
Q_ASSIGN U3180 ( .B(clk), .A(\g.we_clk [13210]));
Q_ASSIGN U3181 ( .B(clk), .A(\g.we_clk [13209]));
Q_ASSIGN U3182 ( .B(clk), .A(\g.we_clk [13208]));
Q_ASSIGN U3183 ( .B(clk), .A(\g.we_clk [13207]));
Q_ASSIGN U3184 ( .B(clk), .A(\g.we_clk [13206]));
Q_ASSIGN U3185 ( .B(clk), .A(\g.we_clk [13205]));
Q_ASSIGN U3186 ( .B(clk), .A(\g.we_clk [13204]));
Q_ASSIGN U3187 ( .B(clk), .A(\g.we_clk [13203]));
Q_ASSIGN U3188 ( .B(clk), .A(\g.we_clk [13202]));
Q_ASSIGN U3189 ( .B(clk), .A(\g.we_clk [13201]));
Q_ASSIGN U3190 ( .B(clk), .A(\g.we_clk [13200]));
Q_ASSIGN U3191 ( .B(clk), .A(\g.we_clk [13199]));
Q_ASSIGN U3192 ( .B(clk), .A(\g.we_clk [13198]));
Q_ASSIGN U3193 ( .B(clk), .A(\g.we_clk [13197]));
Q_ASSIGN U3194 ( .B(clk), .A(\g.we_clk [13196]));
Q_ASSIGN U3195 ( .B(clk), .A(\g.we_clk [13195]));
Q_ASSIGN U3196 ( .B(clk), .A(\g.we_clk [13194]));
Q_ASSIGN U3197 ( .B(clk), .A(\g.we_clk [13193]));
Q_ASSIGN U3198 ( .B(clk), .A(\g.we_clk [13192]));
Q_ASSIGN U3199 ( .B(clk), .A(\g.we_clk [13191]));
Q_ASSIGN U3200 ( .B(clk), .A(\g.we_clk [13190]));
Q_ASSIGN U3201 ( .B(clk), .A(\g.we_clk [13189]));
Q_ASSIGN U3202 ( .B(clk), .A(\g.we_clk [13188]));
Q_ASSIGN U3203 ( .B(clk), .A(\g.we_clk [13187]));
Q_ASSIGN U3204 ( .B(clk), .A(\g.we_clk [13186]));
Q_ASSIGN U3205 ( .B(clk), .A(\g.we_clk [13185]));
Q_ASSIGN U3206 ( .B(clk), .A(\g.we_clk [13184]));
Q_ASSIGN U3207 ( .B(clk), .A(\g.we_clk [13183]));
Q_ASSIGN U3208 ( .B(clk), .A(\g.we_clk [13182]));
Q_ASSIGN U3209 ( .B(clk), .A(\g.we_clk [13181]));
Q_ASSIGN U3210 ( .B(clk), .A(\g.we_clk [13180]));
Q_ASSIGN U3211 ( .B(clk), .A(\g.we_clk [13179]));
Q_ASSIGN U3212 ( .B(clk), .A(\g.we_clk [13178]));
Q_ASSIGN U3213 ( .B(clk), .A(\g.we_clk [13177]));
Q_ASSIGN U3214 ( .B(clk), .A(\g.we_clk [13176]));
Q_ASSIGN U3215 ( .B(clk), .A(\g.we_clk [13175]));
Q_ASSIGN U3216 ( .B(clk), .A(\g.we_clk [13174]));
Q_ASSIGN U3217 ( .B(clk), .A(\g.we_clk [13173]));
Q_ASSIGN U3218 ( .B(clk), .A(\g.we_clk [13172]));
Q_ASSIGN U3219 ( .B(clk), .A(\g.we_clk [13171]));
Q_ASSIGN U3220 ( .B(clk), .A(\g.we_clk [13170]));
Q_ASSIGN U3221 ( .B(clk), .A(\g.we_clk [13169]));
Q_ASSIGN U3222 ( .B(clk), .A(\g.we_clk [13168]));
Q_ASSIGN U3223 ( .B(clk), .A(\g.we_clk [13167]));
Q_ASSIGN U3224 ( .B(clk), .A(\g.we_clk [13166]));
Q_ASSIGN U3225 ( .B(clk), .A(\g.we_clk [13165]));
Q_ASSIGN U3226 ( .B(clk), .A(\g.we_clk [13164]));
Q_ASSIGN U3227 ( .B(clk), .A(\g.we_clk [13163]));
Q_ASSIGN U3228 ( .B(clk), .A(\g.we_clk [13162]));
Q_ASSIGN U3229 ( .B(clk), .A(\g.we_clk [13161]));
Q_ASSIGN U3230 ( .B(clk), .A(\g.we_clk [13160]));
Q_ASSIGN U3231 ( .B(clk), .A(\g.we_clk [13159]));
Q_ASSIGN U3232 ( .B(clk), .A(\g.we_clk [13158]));
Q_ASSIGN U3233 ( .B(clk), .A(\g.we_clk [13157]));
Q_ASSIGN U3234 ( .B(clk), .A(\g.we_clk [13156]));
Q_ASSIGN U3235 ( .B(clk), .A(\g.we_clk [13155]));
Q_ASSIGN U3236 ( .B(clk), .A(\g.we_clk [13154]));
Q_ASSIGN U3237 ( .B(clk), .A(\g.we_clk [13153]));
Q_ASSIGN U3238 ( .B(clk), .A(\g.we_clk [13152]));
Q_ASSIGN U3239 ( .B(clk), .A(\g.we_clk [13151]));
Q_ASSIGN U3240 ( .B(clk), .A(\g.we_clk [13150]));
Q_ASSIGN U3241 ( .B(clk), .A(\g.we_clk [13149]));
Q_ASSIGN U3242 ( .B(clk), .A(\g.we_clk [13148]));
Q_ASSIGN U3243 ( .B(clk), .A(\g.we_clk [13147]));
Q_ASSIGN U3244 ( .B(clk), .A(\g.we_clk [13146]));
Q_ASSIGN U3245 ( .B(clk), .A(\g.we_clk [13145]));
Q_ASSIGN U3246 ( .B(clk), .A(\g.we_clk [13144]));
Q_ASSIGN U3247 ( .B(clk), .A(\g.we_clk [13143]));
Q_ASSIGN U3248 ( .B(clk), .A(\g.we_clk [13142]));
Q_ASSIGN U3249 ( .B(clk), .A(\g.we_clk [13141]));
Q_ASSIGN U3250 ( .B(clk), .A(\g.we_clk [13140]));
Q_ASSIGN U3251 ( .B(clk), .A(\g.we_clk [13139]));
Q_ASSIGN U3252 ( .B(clk), .A(\g.we_clk [13138]));
Q_ASSIGN U3253 ( .B(clk), .A(\g.we_clk [13137]));
Q_ASSIGN U3254 ( .B(clk), .A(\g.we_clk [13136]));
Q_ASSIGN U3255 ( .B(clk), .A(\g.we_clk [13135]));
Q_ASSIGN U3256 ( .B(clk), .A(\g.we_clk [13134]));
Q_ASSIGN U3257 ( .B(clk), .A(\g.we_clk [13133]));
Q_ASSIGN U3258 ( .B(clk), .A(\g.we_clk [13132]));
Q_ASSIGN U3259 ( .B(clk), .A(\g.we_clk [13131]));
Q_ASSIGN U3260 ( .B(clk), .A(\g.we_clk [13130]));
Q_ASSIGN U3261 ( .B(clk), .A(\g.we_clk [13129]));
Q_ASSIGN U3262 ( .B(clk), .A(\g.we_clk [13128]));
Q_ASSIGN U3263 ( .B(clk), .A(\g.we_clk [13127]));
Q_ASSIGN U3264 ( .B(clk), .A(\g.we_clk [13126]));
Q_ASSIGN U3265 ( .B(clk), .A(\g.we_clk [13125]));
Q_ASSIGN U3266 ( .B(clk), .A(\g.we_clk [13124]));
Q_ASSIGN U3267 ( .B(clk), .A(\g.we_clk [13123]));
Q_ASSIGN U3268 ( .B(clk), .A(\g.we_clk [13122]));
Q_ASSIGN U3269 ( .B(clk), .A(\g.we_clk [13121]));
Q_ASSIGN U3270 ( .B(clk), .A(\g.we_clk [13120]));
Q_ASSIGN U3271 ( .B(clk), .A(\g.we_clk [13119]));
Q_ASSIGN U3272 ( .B(clk), .A(\g.we_clk [13118]));
Q_ASSIGN U3273 ( .B(clk), .A(\g.we_clk [13117]));
Q_ASSIGN U3274 ( .B(clk), .A(\g.we_clk [13116]));
Q_ASSIGN U3275 ( .B(clk), .A(\g.we_clk [13115]));
Q_ASSIGN U3276 ( .B(clk), .A(\g.we_clk [13114]));
Q_ASSIGN U3277 ( .B(clk), .A(\g.we_clk [13113]));
Q_ASSIGN U3278 ( .B(clk), .A(\g.we_clk [13112]));
Q_ASSIGN U3279 ( .B(clk), .A(\g.we_clk [13111]));
Q_ASSIGN U3280 ( .B(clk), .A(\g.we_clk [13110]));
Q_ASSIGN U3281 ( .B(clk), .A(\g.we_clk [13109]));
Q_ASSIGN U3282 ( .B(clk), .A(\g.we_clk [13108]));
Q_ASSIGN U3283 ( .B(clk), .A(\g.we_clk [13107]));
Q_ASSIGN U3284 ( .B(clk), .A(\g.we_clk [13106]));
Q_ASSIGN U3285 ( .B(clk), .A(\g.we_clk [13105]));
Q_ASSIGN U3286 ( .B(clk), .A(\g.we_clk [13104]));
Q_ASSIGN U3287 ( .B(clk), .A(\g.we_clk [13103]));
Q_ASSIGN U3288 ( .B(clk), .A(\g.we_clk [13102]));
Q_ASSIGN U3289 ( .B(clk), .A(\g.we_clk [13101]));
Q_ASSIGN U3290 ( .B(clk), .A(\g.we_clk [13100]));
Q_ASSIGN U3291 ( .B(clk), .A(\g.we_clk [13099]));
Q_ASSIGN U3292 ( .B(clk), .A(\g.we_clk [13098]));
Q_ASSIGN U3293 ( .B(clk), .A(\g.we_clk [13097]));
Q_ASSIGN U3294 ( .B(clk), .A(\g.we_clk [13096]));
Q_ASSIGN U3295 ( .B(clk), .A(\g.we_clk [13095]));
Q_ASSIGN U3296 ( .B(clk), .A(\g.we_clk [13094]));
Q_ASSIGN U3297 ( .B(clk), .A(\g.we_clk [13093]));
Q_ASSIGN U3298 ( .B(clk), .A(\g.we_clk [13092]));
Q_ASSIGN U3299 ( .B(clk), .A(\g.we_clk [13091]));
Q_ASSIGN U3300 ( .B(clk), .A(\g.we_clk [13090]));
Q_ASSIGN U3301 ( .B(clk), .A(\g.we_clk [13089]));
Q_ASSIGN U3302 ( .B(clk), .A(\g.we_clk [13088]));
Q_ASSIGN U3303 ( .B(clk), .A(\g.we_clk [13087]));
Q_ASSIGN U3304 ( .B(clk), .A(\g.we_clk [13086]));
Q_ASSIGN U3305 ( .B(clk), .A(\g.we_clk [13085]));
Q_ASSIGN U3306 ( .B(clk), .A(\g.we_clk [13084]));
Q_ASSIGN U3307 ( .B(clk), .A(\g.we_clk [13083]));
Q_ASSIGN U3308 ( .B(clk), .A(\g.we_clk [13082]));
Q_ASSIGN U3309 ( .B(clk), .A(\g.we_clk [13081]));
Q_ASSIGN U3310 ( .B(clk), .A(\g.we_clk [13080]));
Q_ASSIGN U3311 ( .B(clk), .A(\g.we_clk [13079]));
Q_ASSIGN U3312 ( .B(clk), .A(\g.we_clk [13078]));
Q_ASSIGN U3313 ( .B(clk), .A(\g.we_clk [13077]));
Q_ASSIGN U3314 ( .B(clk), .A(\g.we_clk [13076]));
Q_ASSIGN U3315 ( .B(clk), .A(\g.we_clk [13075]));
Q_ASSIGN U3316 ( .B(clk), .A(\g.we_clk [13074]));
Q_ASSIGN U3317 ( .B(clk), .A(\g.we_clk [13073]));
Q_ASSIGN U3318 ( .B(clk), .A(\g.we_clk [13072]));
Q_ASSIGN U3319 ( .B(clk), .A(\g.we_clk [13071]));
Q_ASSIGN U3320 ( .B(clk), .A(\g.we_clk [13070]));
Q_ASSIGN U3321 ( .B(clk), .A(\g.we_clk [13069]));
Q_ASSIGN U3322 ( .B(clk), .A(\g.we_clk [13068]));
Q_ASSIGN U3323 ( .B(clk), .A(\g.we_clk [13067]));
Q_ASSIGN U3324 ( .B(clk), .A(\g.we_clk [13066]));
Q_ASSIGN U3325 ( .B(clk), .A(\g.we_clk [13065]));
Q_ASSIGN U3326 ( .B(clk), .A(\g.we_clk [13064]));
Q_ASSIGN U3327 ( .B(clk), .A(\g.we_clk [13063]));
Q_ASSIGN U3328 ( .B(clk), .A(\g.we_clk [13062]));
Q_ASSIGN U3329 ( .B(clk), .A(\g.we_clk [13061]));
Q_ASSIGN U3330 ( .B(clk), .A(\g.we_clk [13060]));
Q_ASSIGN U3331 ( .B(clk), .A(\g.we_clk [13059]));
Q_ASSIGN U3332 ( .B(clk), .A(\g.we_clk [13058]));
Q_ASSIGN U3333 ( .B(clk), .A(\g.we_clk [13057]));
Q_ASSIGN U3334 ( .B(clk), .A(\g.we_clk [13056]));
Q_ASSIGN U3335 ( .B(clk), .A(\g.we_clk [13055]));
Q_ASSIGN U3336 ( .B(clk), .A(\g.we_clk [13054]));
Q_ASSIGN U3337 ( .B(clk), .A(\g.we_clk [13053]));
Q_ASSIGN U3338 ( .B(clk), .A(\g.we_clk [13052]));
Q_ASSIGN U3339 ( .B(clk), .A(\g.we_clk [13051]));
Q_ASSIGN U3340 ( .B(clk), .A(\g.we_clk [13050]));
Q_ASSIGN U3341 ( .B(clk), .A(\g.we_clk [13049]));
Q_ASSIGN U3342 ( .B(clk), .A(\g.we_clk [13048]));
Q_ASSIGN U3343 ( .B(clk), .A(\g.we_clk [13047]));
Q_ASSIGN U3344 ( .B(clk), .A(\g.we_clk [13046]));
Q_ASSIGN U3345 ( .B(clk), .A(\g.we_clk [13045]));
Q_ASSIGN U3346 ( .B(clk), .A(\g.we_clk [13044]));
Q_ASSIGN U3347 ( .B(clk), .A(\g.we_clk [13043]));
Q_ASSIGN U3348 ( .B(clk), .A(\g.we_clk [13042]));
Q_ASSIGN U3349 ( .B(clk), .A(\g.we_clk [13041]));
Q_ASSIGN U3350 ( .B(clk), .A(\g.we_clk [13040]));
Q_ASSIGN U3351 ( .B(clk), .A(\g.we_clk [13039]));
Q_ASSIGN U3352 ( .B(clk), .A(\g.we_clk [13038]));
Q_ASSIGN U3353 ( .B(clk), .A(\g.we_clk [13037]));
Q_ASSIGN U3354 ( .B(clk), .A(\g.we_clk [13036]));
Q_ASSIGN U3355 ( .B(clk), .A(\g.we_clk [13035]));
Q_ASSIGN U3356 ( .B(clk), .A(\g.we_clk [13034]));
Q_ASSIGN U3357 ( .B(clk), .A(\g.we_clk [13033]));
Q_ASSIGN U3358 ( .B(clk), .A(\g.we_clk [13032]));
Q_ASSIGN U3359 ( .B(clk), .A(\g.we_clk [13031]));
Q_ASSIGN U3360 ( .B(clk), .A(\g.we_clk [13030]));
Q_ASSIGN U3361 ( .B(clk), .A(\g.we_clk [13029]));
Q_ASSIGN U3362 ( .B(clk), .A(\g.we_clk [13028]));
Q_ASSIGN U3363 ( .B(clk), .A(\g.we_clk [13027]));
Q_ASSIGN U3364 ( .B(clk), .A(\g.we_clk [13026]));
Q_ASSIGN U3365 ( .B(clk), .A(\g.we_clk [13025]));
Q_ASSIGN U3366 ( .B(clk), .A(\g.we_clk [13024]));
Q_ASSIGN U3367 ( .B(clk), .A(\g.we_clk [13023]));
Q_ASSIGN U3368 ( .B(clk), .A(\g.we_clk [13022]));
Q_ASSIGN U3369 ( .B(clk), .A(\g.we_clk [13021]));
Q_ASSIGN U3370 ( .B(clk), .A(\g.we_clk [13020]));
Q_ASSIGN U3371 ( .B(clk), .A(\g.we_clk [13019]));
Q_ASSIGN U3372 ( .B(clk), .A(\g.we_clk [13018]));
Q_ASSIGN U3373 ( .B(clk), .A(\g.we_clk [13017]));
Q_ASSIGN U3374 ( .B(clk), .A(\g.we_clk [13016]));
Q_ASSIGN U3375 ( .B(clk), .A(\g.we_clk [13015]));
Q_ASSIGN U3376 ( .B(clk), .A(\g.we_clk [13014]));
Q_ASSIGN U3377 ( .B(clk), .A(\g.we_clk [13013]));
Q_ASSIGN U3378 ( .B(clk), .A(\g.we_clk [13012]));
Q_ASSIGN U3379 ( .B(clk), .A(\g.we_clk [13011]));
Q_ASSIGN U3380 ( .B(clk), .A(\g.we_clk [13010]));
Q_ASSIGN U3381 ( .B(clk), .A(\g.we_clk [13009]));
Q_ASSIGN U3382 ( .B(clk), .A(\g.we_clk [13008]));
Q_ASSIGN U3383 ( .B(clk), .A(\g.we_clk [13007]));
Q_ASSIGN U3384 ( .B(clk), .A(\g.we_clk [13006]));
Q_ASSIGN U3385 ( .B(clk), .A(\g.we_clk [13005]));
Q_ASSIGN U3386 ( .B(clk), .A(\g.we_clk [13004]));
Q_ASSIGN U3387 ( .B(clk), .A(\g.we_clk [13003]));
Q_ASSIGN U3388 ( .B(clk), .A(\g.we_clk [13002]));
Q_ASSIGN U3389 ( .B(clk), .A(\g.we_clk [13001]));
Q_ASSIGN U3390 ( .B(clk), .A(\g.we_clk [13000]));
Q_ASSIGN U3391 ( .B(clk), .A(\g.we_clk [12999]));
Q_ASSIGN U3392 ( .B(clk), .A(\g.we_clk [12998]));
Q_ASSIGN U3393 ( .B(clk), .A(\g.we_clk [12997]));
Q_ASSIGN U3394 ( .B(clk), .A(\g.we_clk [12996]));
Q_ASSIGN U3395 ( .B(clk), .A(\g.we_clk [12995]));
Q_ASSIGN U3396 ( .B(clk), .A(\g.we_clk [12994]));
Q_ASSIGN U3397 ( .B(clk), .A(\g.we_clk [12993]));
Q_ASSIGN U3398 ( .B(clk), .A(\g.we_clk [12992]));
Q_ASSIGN U3399 ( .B(clk), .A(\g.we_clk [12991]));
Q_ASSIGN U3400 ( .B(clk), .A(\g.we_clk [12990]));
Q_ASSIGN U3401 ( .B(clk), .A(\g.we_clk [12989]));
Q_ASSIGN U3402 ( .B(clk), .A(\g.we_clk [12988]));
Q_ASSIGN U3403 ( .B(clk), .A(\g.we_clk [12987]));
Q_ASSIGN U3404 ( .B(clk), .A(\g.we_clk [12986]));
Q_ASSIGN U3405 ( .B(clk), .A(\g.we_clk [12985]));
Q_ASSIGN U3406 ( .B(clk), .A(\g.we_clk [12984]));
Q_ASSIGN U3407 ( .B(clk), .A(\g.we_clk [12983]));
Q_ASSIGN U3408 ( .B(clk), .A(\g.we_clk [12982]));
Q_ASSIGN U3409 ( .B(clk), .A(\g.we_clk [12981]));
Q_ASSIGN U3410 ( .B(clk), .A(\g.we_clk [12980]));
Q_ASSIGN U3411 ( .B(clk), .A(\g.we_clk [12979]));
Q_ASSIGN U3412 ( .B(clk), .A(\g.we_clk [12978]));
Q_ASSIGN U3413 ( .B(clk), .A(\g.we_clk [12977]));
Q_ASSIGN U3414 ( .B(clk), .A(\g.we_clk [12976]));
Q_ASSIGN U3415 ( .B(clk), .A(\g.we_clk [12975]));
Q_ASSIGN U3416 ( .B(clk), .A(\g.we_clk [12974]));
Q_ASSIGN U3417 ( .B(clk), .A(\g.we_clk [12973]));
Q_ASSIGN U3418 ( .B(clk), .A(\g.we_clk [12972]));
Q_ASSIGN U3419 ( .B(clk), .A(\g.we_clk [12971]));
Q_ASSIGN U3420 ( .B(clk), .A(\g.we_clk [12970]));
Q_ASSIGN U3421 ( .B(clk), .A(\g.we_clk [12969]));
Q_ASSIGN U3422 ( .B(clk), .A(\g.we_clk [12968]));
Q_ASSIGN U3423 ( .B(clk), .A(\g.we_clk [12967]));
Q_ASSIGN U3424 ( .B(clk), .A(\g.we_clk [12966]));
Q_ASSIGN U3425 ( .B(clk), .A(\g.we_clk [12965]));
Q_ASSIGN U3426 ( .B(clk), .A(\g.we_clk [12964]));
Q_ASSIGN U3427 ( .B(clk), .A(\g.we_clk [12963]));
Q_ASSIGN U3428 ( .B(clk), .A(\g.we_clk [12962]));
Q_ASSIGN U3429 ( .B(clk), .A(\g.we_clk [12961]));
Q_ASSIGN U3430 ( .B(clk), .A(\g.we_clk [12960]));
Q_ASSIGN U3431 ( .B(clk), .A(\g.we_clk [12959]));
Q_ASSIGN U3432 ( .B(clk), .A(\g.we_clk [12958]));
Q_ASSIGN U3433 ( .B(clk), .A(\g.we_clk [12957]));
Q_ASSIGN U3434 ( .B(clk), .A(\g.we_clk [12956]));
Q_ASSIGN U3435 ( .B(clk), .A(\g.we_clk [12955]));
Q_ASSIGN U3436 ( .B(clk), .A(\g.we_clk [12954]));
Q_ASSIGN U3437 ( .B(clk), .A(\g.we_clk [12953]));
Q_ASSIGN U3438 ( .B(clk), .A(\g.we_clk [12952]));
Q_ASSIGN U3439 ( .B(clk), .A(\g.we_clk [12951]));
Q_ASSIGN U3440 ( .B(clk), .A(\g.we_clk [12950]));
Q_ASSIGN U3441 ( .B(clk), .A(\g.we_clk [12949]));
Q_ASSIGN U3442 ( .B(clk), .A(\g.we_clk [12948]));
Q_ASSIGN U3443 ( .B(clk), .A(\g.we_clk [12947]));
Q_ASSIGN U3444 ( .B(clk), .A(\g.we_clk [12946]));
Q_ASSIGN U3445 ( .B(clk), .A(\g.we_clk [12945]));
Q_ASSIGN U3446 ( .B(clk), .A(\g.we_clk [12944]));
Q_ASSIGN U3447 ( .B(clk), .A(\g.we_clk [12943]));
Q_ASSIGN U3448 ( .B(clk), .A(\g.we_clk [12942]));
Q_ASSIGN U3449 ( .B(clk), .A(\g.we_clk [12941]));
Q_ASSIGN U3450 ( .B(clk), .A(\g.we_clk [12940]));
Q_ASSIGN U3451 ( .B(clk), .A(\g.we_clk [12939]));
Q_ASSIGN U3452 ( .B(clk), .A(\g.we_clk [12938]));
Q_ASSIGN U3453 ( .B(clk), .A(\g.we_clk [12937]));
Q_ASSIGN U3454 ( .B(clk), .A(\g.we_clk [12936]));
Q_ASSIGN U3455 ( .B(clk), .A(\g.we_clk [12935]));
Q_ASSIGN U3456 ( .B(clk), .A(\g.we_clk [12934]));
Q_ASSIGN U3457 ( .B(clk), .A(\g.we_clk [12933]));
Q_ASSIGN U3458 ( .B(clk), .A(\g.we_clk [12932]));
Q_ASSIGN U3459 ( .B(clk), .A(\g.we_clk [12931]));
Q_ASSIGN U3460 ( .B(clk), .A(\g.we_clk [12930]));
Q_ASSIGN U3461 ( .B(clk), .A(\g.we_clk [12929]));
Q_ASSIGN U3462 ( .B(clk), .A(\g.we_clk [12928]));
Q_ASSIGN U3463 ( .B(clk), .A(\g.we_clk [12927]));
Q_ASSIGN U3464 ( .B(clk), .A(\g.we_clk [12926]));
Q_ASSIGN U3465 ( .B(clk), .A(\g.we_clk [12925]));
Q_ASSIGN U3466 ( .B(clk), .A(\g.we_clk [12924]));
Q_ASSIGN U3467 ( .B(clk), .A(\g.we_clk [12923]));
Q_ASSIGN U3468 ( .B(clk), .A(\g.we_clk [12922]));
Q_ASSIGN U3469 ( .B(clk), .A(\g.we_clk [12921]));
Q_ASSIGN U3470 ( .B(clk), .A(\g.we_clk [12920]));
Q_ASSIGN U3471 ( .B(clk), .A(\g.we_clk [12919]));
Q_ASSIGN U3472 ( .B(clk), .A(\g.we_clk [12918]));
Q_ASSIGN U3473 ( .B(clk), .A(\g.we_clk [12917]));
Q_ASSIGN U3474 ( .B(clk), .A(\g.we_clk [12916]));
Q_ASSIGN U3475 ( .B(clk), .A(\g.we_clk [12915]));
Q_ASSIGN U3476 ( .B(clk), .A(\g.we_clk [12914]));
Q_ASSIGN U3477 ( .B(clk), .A(\g.we_clk [12913]));
Q_ASSIGN U3478 ( .B(clk), .A(\g.we_clk [12912]));
Q_ASSIGN U3479 ( .B(clk), .A(\g.we_clk [12911]));
Q_ASSIGN U3480 ( .B(clk), .A(\g.we_clk [12910]));
Q_ASSIGN U3481 ( .B(clk), .A(\g.we_clk [12909]));
Q_ASSIGN U3482 ( .B(clk), .A(\g.we_clk [12908]));
Q_ASSIGN U3483 ( .B(clk), .A(\g.we_clk [12907]));
Q_ASSIGN U3484 ( .B(clk), .A(\g.we_clk [12906]));
Q_ASSIGN U3485 ( .B(clk), .A(\g.we_clk [12905]));
Q_ASSIGN U3486 ( .B(clk), .A(\g.we_clk [12904]));
Q_ASSIGN U3487 ( .B(clk), .A(\g.we_clk [12903]));
Q_ASSIGN U3488 ( .B(clk), .A(\g.we_clk [12902]));
Q_ASSIGN U3489 ( .B(clk), .A(\g.we_clk [12901]));
Q_ASSIGN U3490 ( .B(clk), .A(\g.we_clk [12900]));
Q_ASSIGN U3491 ( .B(clk), .A(\g.we_clk [12899]));
Q_ASSIGN U3492 ( .B(clk), .A(\g.we_clk [12898]));
Q_ASSIGN U3493 ( .B(clk), .A(\g.we_clk [12897]));
Q_ASSIGN U3494 ( .B(clk), .A(\g.we_clk [12896]));
Q_ASSIGN U3495 ( .B(clk), .A(\g.we_clk [12895]));
Q_ASSIGN U3496 ( .B(clk), .A(\g.we_clk [12894]));
Q_ASSIGN U3497 ( .B(clk), .A(\g.we_clk [12893]));
Q_ASSIGN U3498 ( .B(clk), .A(\g.we_clk [12892]));
Q_ASSIGN U3499 ( .B(clk), .A(\g.we_clk [12891]));
Q_ASSIGN U3500 ( .B(clk), .A(\g.we_clk [12890]));
Q_ASSIGN U3501 ( .B(clk), .A(\g.we_clk [12889]));
Q_ASSIGN U3502 ( .B(clk), .A(\g.we_clk [12888]));
Q_ASSIGN U3503 ( .B(clk), .A(\g.we_clk [12887]));
Q_ASSIGN U3504 ( .B(clk), .A(\g.we_clk [12886]));
Q_ASSIGN U3505 ( .B(clk), .A(\g.we_clk [12885]));
Q_ASSIGN U3506 ( .B(clk), .A(\g.we_clk [12884]));
Q_ASSIGN U3507 ( .B(clk), .A(\g.we_clk [12883]));
Q_ASSIGN U3508 ( .B(clk), .A(\g.we_clk [12882]));
Q_ASSIGN U3509 ( .B(clk), .A(\g.we_clk [12881]));
Q_ASSIGN U3510 ( .B(clk), .A(\g.we_clk [12880]));
Q_ASSIGN U3511 ( .B(clk), .A(\g.we_clk [12879]));
Q_ASSIGN U3512 ( .B(clk), .A(\g.we_clk [12878]));
Q_ASSIGN U3513 ( .B(clk), .A(\g.we_clk [12877]));
Q_ASSIGN U3514 ( .B(clk), .A(\g.we_clk [12876]));
Q_ASSIGN U3515 ( .B(clk), .A(\g.we_clk [12875]));
Q_ASSIGN U3516 ( .B(clk), .A(\g.we_clk [12874]));
Q_ASSIGN U3517 ( .B(clk), .A(\g.we_clk [12873]));
Q_ASSIGN U3518 ( .B(clk), .A(\g.we_clk [12872]));
Q_ASSIGN U3519 ( .B(clk), .A(\g.we_clk [12871]));
Q_ASSIGN U3520 ( .B(clk), .A(\g.we_clk [12870]));
Q_ASSIGN U3521 ( .B(clk), .A(\g.we_clk [12869]));
Q_ASSIGN U3522 ( .B(clk), .A(\g.we_clk [12868]));
Q_ASSIGN U3523 ( .B(clk), .A(\g.we_clk [12867]));
Q_ASSIGN U3524 ( .B(clk), .A(\g.we_clk [12866]));
Q_ASSIGN U3525 ( .B(clk), .A(\g.we_clk [12865]));
Q_ASSIGN U3526 ( .B(clk), .A(\g.we_clk [12864]));
Q_ASSIGN U3527 ( .B(clk), .A(\g.we_clk [12863]));
Q_ASSIGN U3528 ( .B(clk), .A(\g.we_clk [12862]));
Q_ASSIGN U3529 ( .B(clk), .A(\g.we_clk [12861]));
Q_ASSIGN U3530 ( .B(clk), .A(\g.we_clk [12860]));
Q_ASSIGN U3531 ( .B(clk), .A(\g.we_clk [12859]));
Q_ASSIGN U3532 ( .B(clk), .A(\g.we_clk [12858]));
Q_ASSIGN U3533 ( .B(clk), .A(\g.we_clk [12857]));
Q_ASSIGN U3534 ( .B(clk), .A(\g.we_clk [12856]));
Q_ASSIGN U3535 ( .B(clk), .A(\g.we_clk [12855]));
Q_ASSIGN U3536 ( .B(clk), .A(\g.we_clk [12854]));
Q_ASSIGN U3537 ( .B(clk), .A(\g.we_clk [12853]));
Q_ASSIGN U3538 ( .B(clk), .A(\g.we_clk [12852]));
Q_ASSIGN U3539 ( .B(clk), .A(\g.we_clk [12851]));
Q_ASSIGN U3540 ( .B(clk), .A(\g.we_clk [12850]));
Q_ASSIGN U3541 ( .B(clk), .A(\g.we_clk [12849]));
Q_ASSIGN U3542 ( .B(clk), .A(\g.we_clk [12848]));
Q_ASSIGN U3543 ( .B(clk), .A(\g.we_clk [12847]));
Q_ASSIGN U3544 ( .B(clk), .A(\g.we_clk [12846]));
Q_ASSIGN U3545 ( .B(clk), .A(\g.we_clk [12845]));
Q_ASSIGN U3546 ( .B(clk), .A(\g.we_clk [12844]));
Q_ASSIGN U3547 ( .B(clk), .A(\g.we_clk [12843]));
Q_ASSIGN U3548 ( .B(clk), .A(\g.we_clk [12842]));
Q_ASSIGN U3549 ( .B(clk), .A(\g.we_clk [12841]));
Q_ASSIGN U3550 ( .B(clk), .A(\g.we_clk [12840]));
Q_ASSIGN U3551 ( .B(clk), .A(\g.we_clk [12839]));
Q_ASSIGN U3552 ( .B(clk), .A(\g.we_clk [12838]));
Q_ASSIGN U3553 ( .B(clk), .A(\g.we_clk [12837]));
Q_ASSIGN U3554 ( .B(clk), .A(\g.we_clk [12836]));
Q_ASSIGN U3555 ( .B(clk), .A(\g.we_clk [12835]));
Q_ASSIGN U3556 ( .B(clk), .A(\g.we_clk [12834]));
Q_ASSIGN U3557 ( .B(clk), .A(\g.we_clk [12833]));
Q_ASSIGN U3558 ( .B(clk), .A(\g.we_clk [12832]));
Q_ASSIGN U3559 ( .B(clk), .A(\g.we_clk [12831]));
Q_ASSIGN U3560 ( .B(clk), .A(\g.we_clk [12830]));
Q_ASSIGN U3561 ( .B(clk), .A(\g.we_clk [12829]));
Q_ASSIGN U3562 ( .B(clk), .A(\g.we_clk [12828]));
Q_ASSIGN U3563 ( .B(clk), .A(\g.we_clk [12827]));
Q_ASSIGN U3564 ( .B(clk), .A(\g.we_clk [12826]));
Q_ASSIGN U3565 ( .B(clk), .A(\g.we_clk [12825]));
Q_ASSIGN U3566 ( .B(clk), .A(\g.we_clk [12824]));
Q_ASSIGN U3567 ( .B(clk), .A(\g.we_clk [12823]));
Q_ASSIGN U3568 ( .B(clk), .A(\g.we_clk [12822]));
Q_ASSIGN U3569 ( .B(clk), .A(\g.we_clk [12821]));
Q_ASSIGN U3570 ( .B(clk), .A(\g.we_clk [12820]));
Q_ASSIGN U3571 ( .B(clk), .A(\g.we_clk [12819]));
Q_ASSIGN U3572 ( .B(clk), .A(\g.we_clk [12818]));
Q_ASSIGN U3573 ( .B(clk), .A(\g.we_clk [12817]));
Q_ASSIGN U3574 ( .B(clk), .A(\g.we_clk [12816]));
Q_ASSIGN U3575 ( .B(clk), .A(\g.we_clk [12815]));
Q_ASSIGN U3576 ( .B(clk), .A(\g.we_clk [12814]));
Q_ASSIGN U3577 ( .B(clk), .A(\g.we_clk [12813]));
Q_ASSIGN U3578 ( .B(clk), .A(\g.we_clk [12812]));
Q_ASSIGN U3579 ( .B(clk), .A(\g.we_clk [12811]));
Q_ASSIGN U3580 ( .B(clk), .A(\g.we_clk [12810]));
Q_ASSIGN U3581 ( .B(clk), .A(\g.we_clk [12809]));
Q_ASSIGN U3582 ( .B(clk), .A(\g.we_clk [12808]));
Q_ASSIGN U3583 ( .B(clk), .A(\g.we_clk [12807]));
Q_ASSIGN U3584 ( .B(clk), .A(\g.we_clk [12806]));
Q_ASSIGN U3585 ( .B(clk), .A(\g.we_clk [12805]));
Q_ASSIGN U3586 ( .B(clk), .A(\g.we_clk [12804]));
Q_ASSIGN U3587 ( .B(clk), .A(\g.we_clk [12803]));
Q_ASSIGN U3588 ( .B(clk), .A(\g.we_clk [12802]));
Q_ASSIGN U3589 ( .B(clk), .A(\g.we_clk [12801]));
Q_ASSIGN U3590 ( .B(clk), .A(\g.we_clk [12800]));
Q_ASSIGN U3591 ( .B(clk), .A(\g.we_clk [12799]));
Q_ASSIGN U3592 ( .B(clk), .A(\g.we_clk [12798]));
Q_ASSIGN U3593 ( .B(clk), .A(\g.we_clk [12797]));
Q_ASSIGN U3594 ( .B(clk), .A(\g.we_clk [12796]));
Q_ASSIGN U3595 ( .B(clk), .A(\g.we_clk [12795]));
Q_ASSIGN U3596 ( .B(clk), .A(\g.we_clk [12794]));
Q_ASSIGN U3597 ( .B(clk), .A(\g.we_clk [12793]));
Q_ASSIGN U3598 ( .B(clk), .A(\g.we_clk [12792]));
Q_ASSIGN U3599 ( .B(clk), .A(\g.we_clk [12791]));
Q_ASSIGN U3600 ( .B(clk), .A(\g.we_clk [12790]));
Q_ASSIGN U3601 ( .B(clk), .A(\g.we_clk [12789]));
Q_ASSIGN U3602 ( .B(clk), .A(\g.we_clk [12788]));
Q_ASSIGN U3603 ( .B(clk), .A(\g.we_clk [12787]));
Q_ASSIGN U3604 ( .B(clk), .A(\g.we_clk [12786]));
Q_ASSIGN U3605 ( .B(clk), .A(\g.we_clk [12785]));
Q_ASSIGN U3606 ( .B(clk), .A(\g.we_clk [12784]));
Q_ASSIGN U3607 ( .B(clk), .A(\g.we_clk [12783]));
Q_ASSIGN U3608 ( .B(clk), .A(\g.we_clk [12782]));
Q_ASSIGN U3609 ( .B(clk), .A(\g.we_clk [12781]));
Q_ASSIGN U3610 ( .B(clk), .A(\g.we_clk [12780]));
Q_ASSIGN U3611 ( .B(clk), .A(\g.we_clk [12779]));
Q_ASSIGN U3612 ( .B(clk), .A(\g.we_clk [12778]));
Q_ASSIGN U3613 ( .B(clk), .A(\g.we_clk [12777]));
Q_ASSIGN U3614 ( .B(clk), .A(\g.we_clk [12776]));
Q_ASSIGN U3615 ( .B(clk), .A(\g.we_clk [12775]));
Q_ASSIGN U3616 ( .B(clk), .A(\g.we_clk [12774]));
Q_ASSIGN U3617 ( .B(clk), .A(\g.we_clk [12773]));
Q_ASSIGN U3618 ( .B(clk), .A(\g.we_clk [12772]));
Q_ASSIGN U3619 ( .B(clk), .A(\g.we_clk [12771]));
Q_ASSIGN U3620 ( .B(clk), .A(\g.we_clk [12770]));
Q_ASSIGN U3621 ( .B(clk), .A(\g.we_clk [12769]));
Q_ASSIGN U3622 ( .B(clk), .A(\g.we_clk [12768]));
Q_ASSIGN U3623 ( .B(clk), .A(\g.we_clk [12767]));
Q_ASSIGN U3624 ( .B(clk), .A(\g.we_clk [12766]));
Q_ASSIGN U3625 ( .B(clk), .A(\g.we_clk [12765]));
Q_ASSIGN U3626 ( .B(clk), .A(\g.we_clk [12764]));
Q_ASSIGN U3627 ( .B(clk), .A(\g.we_clk [12763]));
Q_ASSIGN U3628 ( .B(clk), .A(\g.we_clk [12762]));
Q_ASSIGN U3629 ( .B(clk), .A(\g.we_clk [12761]));
Q_ASSIGN U3630 ( .B(clk), .A(\g.we_clk [12760]));
Q_ASSIGN U3631 ( .B(clk), .A(\g.we_clk [12759]));
Q_ASSIGN U3632 ( .B(clk), .A(\g.we_clk [12758]));
Q_ASSIGN U3633 ( .B(clk), .A(\g.we_clk [12757]));
Q_ASSIGN U3634 ( .B(clk), .A(\g.we_clk [12756]));
Q_ASSIGN U3635 ( .B(clk), .A(\g.we_clk [12755]));
Q_ASSIGN U3636 ( .B(clk), .A(\g.we_clk [12754]));
Q_ASSIGN U3637 ( .B(clk), .A(\g.we_clk [12753]));
Q_ASSIGN U3638 ( .B(clk), .A(\g.we_clk [12752]));
Q_ASSIGN U3639 ( .B(clk), .A(\g.we_clk [12751]));
Q_ASSIGN U3640 ( .B(clk), .A(\g.we_clk [12750]));
Q_ASSIGN U3641 ( .B(clk), .A(\g.we_clk [12749]));
Q_ASSIGN U3642 ( .B(clk), .A(\g.we_clk [12748]));
Q_ASSIGN U3643 ( .B(clk), .A(\g.we_clk [12747]));
Q_ASSIGN U3644 ( .B(clk), .A(\g.we_clk [12746]));
Q_ASSIGN U3645 ( .B(clk), .A(\g.we_clk [12745]));
Q_ASSIGN U3646 ( .B(clk), .A(\g.we_clk [12744]));
Q_ASSIGN U3647 ( .B(clk), .A(\g.we_clk [12743]));
Q_ASSIGN U3648 ( .B(clk), .A(\g.we_clk [12742]));
Q_ASSIGN U3649 ( .B(clk), .A(\g.we_clk [12741]));
Q_ASSIGN U3650 ( .B(clk), .A(\g.we_clk [12740]));
Q_ASSIGN U3651 ( .B(clk), .A(\g.we_clk [12739]));
Q_ASSIGN U3652 ( .B(clk), .A(\g.we_clk [12738]));
Q_ASSIGN U3653 ( .B(clk), .A(\g.we_clk [12737]));
Q_ASSIGN U3654 ( .B(clk), .A(\g.we_clk [12736]));
Q_ASSIGN U3655 ( .B(clk), .A(\g.we_clk [12735]));
Q_ASSIGN U3656 ( .B(clk), .A(\g.we_clk [12734]));
Q_ASSIGN U3657 ( .B(clk), .A(\g.we_clk [12733]));
Q_ASSIGN U3658 ( .B(clk), .A(\g.we_clk [12732]));
Q_ASSIGN U3659 ( .B(clk), .A(\g.we_clk [12731]));
Q_ASSIGN U3660 ( .B(clk), .A(\g.we_clk [12730]));
Q_ASSIGN U3661 ( .B(clk), .A(\g.we_clk [12729]));
Q_ASSIGN U3662 ( .B(clk), .A(\g.we_clk [12728]));
Q_ASSIGN U3663 ( .B(clk), .A(\g.we_clk [12727]));
Q_ASSIGN U3664 ( .B(clk), .A(\g.we_clk [12726]));
Q_ASSIGN U3665 ( .B(clk), .A(\g.we_clk [12725]));
Q_ASSIGN U3666 ( .B(clk), .A(\g.we_clk [12724]));
Q_ASSIGN U3667 ( .B(clk), .A(\g.we_clk [12723]));
Q_ASSIGN U3668 ( .B(clk), .A(\g.we_clk [12722]));
Q_ASSIGN U3669 ( .B(clk), .A(\g.we_clk [12721]));
Q_ASSIGN U3670 ( .B(clk), .A(\g.we_clk [12720]));
Q_ASSIGN U3671 ( .B(clk), .A(\g.we_clk [12719]));
Q_ASSIGN U3672 ( .B(clk), .A(\g.we_clk [12718]));
Q_ASSIGN U3673 ( .B(clk), .A(\g.we_clk [12717]));
Q_ASSIGN U3674 ( .B(clk), .A(\g.we_clk [12716]));
Q_ASSIGN U3675 ( .B(clk), .A(\g.we_clk [12715]));
Q_ASSIGN U3676 ( .B(clk), .A(\g.we_clk [12714]));
Q_ASSIGN U3677 ( .B(clk), .A(\g.we_clk [12713]));
Q_ASSIGN U3678 ( .B(clk), .A(\g.we_clk [12712]));
Q_ASSIGN U3679 ( .B(clk), .A(\g.we_clk [12711]));
Q_ASSIGN U3680 ( .B(clk), .A(\g.we_clk [12710]));
Q_ASSIGN U3681 ( .B(clk), .A(\g.we_clk [12709]));
Q_ASSIGN U3682 ( .B(clk), .A(\g.we_clk [12708]));
Q_ASSIGN U3683 ( .B(clk), .A(\g.we_clk [12707]));
Q_ASSIGN U3684 ( .B(clk), .A(\g.we_clk [12706]));
Q_ASSIGN U3685 ( .B(clk), .A(\g.we_clk [12705]));
Q_ASSIGN U3686 ( .B(clk), .A(\g.we_clk [12704]));
Q_ASSIGN U3687 ( .B(clk), .A(\g.we_clk [12703]));
Q_ASSIGN U3688 ( .B(clk), .A(\g.we_clk [12702]));
Q_ASSIGN U3689 ( .B(clk), .A(\g.we_clk [12701]));
Q_ASSIGN U3690 ( .B(clk), .A(\g.we_clk [12700]));
Q_ASSIGN U3691 ( .B(clk), .A(\g.we_clk [12699]));
Q_ASSIGN U3692 ( .B(clk), .A(\g.we_clk [12698]));
Q_ASSIGN U3693 ( .B(clk), .A(\g.we_clk [12697]));
Q_ASSIGN U3694 ( .B(clk), .A(\g.we_clk [12696]));
Q_ASSIGN U3695 ( .B(clk), .A(\g.we_clk [12695]));
Q_ASSIGN U3696 ( .B(clk), .A(\g.we_clk [12694]));
Q_ASSIGN U3697 ( .B(clk), .A(\g.we_clk [12693]));
Q_ASSIGN U3698 ( .B(clk), .A(\g.we_clk [12692]));
Q_ASSIGN U3699 ( .B(clk), .A(\g.we_clk [12691]));
Q_ASSIGN U3700 ( .B(clk), .A(\g.we_clk [12690]));
Q_ASSIGN U3701 ( .B(clk), .A(\g.we_clk [12689]));
Q_ASSIGN U3702 ( .B(clk), .A(\g.we_clk [12688]));
Q_ASSIGN U3703 ( .B(clk), .A(\g.we_clk [12687]));
Q_ASSIGN U3704 ( .B(clk), .A(\g.we_clk [12686]));
Q_ASSIGN U3705 ( .B(clk), .A(\g.we_clk [12685]));
Q_ASSIGN U3706 ( .B(clk), .A(\g.we_clk [12684]));
Q_ASSIGN U3707 ( .B(clk), .A(\g.we_clk [12683]));
Q_ASSIGN U3708 ( .B(clk), .A(\g.we_clk [12682]));
Q_ASSIGN U3709 ( .B(clk), .A(\g.we_clk [12681]));
Q_ASSIGN U3710 ( .B(clk), .A(\g.we_clk [12680]));
Q_ASSIGN U3711 ( .B(clk), .A(\g.we_clk [12679]));
Q_ASSIGN U3712 ( .B(clk), .A(\g.we_clk [12678]));
Q_ASSIGN U3713 ( .B(clk), .A(\g.we_clk [12677]));
Q_ASSIGN U3714 ( .B(clk), .A(\g.we_clk [12676]));
Q_ASSIGN U3715 ( .B(clk), .A(\g.we_clk [12675]));
Q_ASSIGN U3716 ( .B(clk), .A(\g.we_clk [12674]));
Q_ASSIGN U3717 ( .B(clk), .A(\g.we_clk [12673]));
Q_ASSIGN U3718 ( .B(clk), .A(\g.we_clk [12672]));
Q_ASSIGN U3719 ( .B(clk), .A(\g.we_clk [12671]));
Q_ASSIGN U3720 ( .B(clk), .A(\g.we_clk [12670]));
Q_ASSIGN U3721 ( .B(clk), .A(\g.we_clk [12669]));
Q_ASSIGN U3722 ( .B(clk), .A(\g.we_clk [12668]));
Q_ASSIGN U3723 ( .B(clk), .A(\g.we_clk [12667]));
Q_ASSIGN U3724 ( .B(clk), .A(\g.we_clk [12666]));
Q_ASSIGN U3725 ( .B(clk), .A(\g.we_clk [12665]));
Q_ASSIGN U3726 ( .B(clk), .A(\g.we_clk [12664]));
Q_ASSIGN U3727 ( .B(clk), .A(\g.we_clk [12663]));
Q_ASSIGN U3728 ( .B(clk), .A(\g.we_clk [12662]));
Q_ASSIGN U3729 ( .B(clk), .A(\g.we_clk [12661]));
Q_ASSIGN U3730 ( .B(clk), .A(\g.we_clk [12660]));
Q_ASSIGN U3731 ( .B(clk), .A(\g.we_clk [12659]));
Q_ASSIGN U3732 ( .B(clk), .A(\g.we_clk [12658]));
Q_ASSIGN U3733 ( .B(clk), .A(\g.we_clk [12657]));
Q_ASSIGN U3734 ( .B(clk), .A(\g.we_clk [12656]));
Q_ASSIGN U3735 ( .B(clk), .A(\g.we_clk [12655]));
Q_ASSIGN U3736 ( .B(clk), .A(\g.we_clk [12654]));
Q_ASSIGN U3737 ( .B(clk), .A(\g.we_clk [12653]));
Q_ASSIGN U3738 ( .B(clk), .A(\g.we_clk [12652]));
Q_ASSIGN U3739 ( .B(clk), .A(\g.we_clk [12651]));
Q_ASSIGN U3740 ( .B(clk), .A(\g.we_clk [12650]));
Q_ASSIGN U3741 ( .B(clk), .A(\g.we_clk [12649]));
Q_ASSIGN U3742 ( .B(clk), .A(\g.we_clk [12648]));
Q_ASSIGN U3743 ( .B(clk), .A(\g.we_clk [12647]));
Q_ASSIGN U3744 ( .B(clk), .A(\g.we_clk [12646]));
Q_ASSIGN U3745 ( .B(clk), .A(\g.we_clk [12645]));
Q_ASSIGN U3746 ( .B(clk), .A(\g.we_clk [12644]));
Q_ASSIGN U3747 ( .B(clk), .A(\g.we_clk [12643]));
Q_ASSIGN U3748 ( .B(clk), .A(\g.we_clk [12642]));
Q_ASSIGN U3749 ( .B(clk), .A(\g.we_clk [12641]));
Q_ASSIGN U3750 ( .B(clk), .A(\g.we_clk [12640]));
Q_ASSIGN U3751 ( .B(clk), .A(\g.we_clk [12639]));
Q_ASSIGN U3752 ( .B(clk), .A(\g.we_clk [12638]));
Q_ASSIGN U3753 ( .B(clk), .A(\g.we_clk [12637]));
Q_ASSIGN U3754 ( .B(clk), .A(\g.we_clk [12636]));
Q_ASSIGN U3755 ( .B(clk), .A(\g.we_clk [12635]));
Q_ASSIGN U3756 ( .B(clk), .A(\g.we_clk [12634]));
Q_ASSIGN U3757 ( .B(clk), .A(\g.we_clk [12633]));
Q_ASSIGN U3758 ( .B(clk), .A(\g.we_clk [12632]));
Q_ASSIGN U3759 ( .B(clk), .A(\g.we_clk [12631]));
Q_ASSIGN U3760 ( .B(clk), .A(\g.we_clk [12630]));
Q_ASSIGN U3761 ( .B(clk), .A(\g.we_clk [12629]));
Q_ASSIGN U3762 ( .B(clk), .A(\g.we_clk [12628]));
Q_ASSIGN U3763 ( .B(clk), .A(\g.we_clk [12627]));
Q_ASSIGN U3764 ( .B(clk), .A(\g.we_clk [12626]));
Q_ASSIGN U3765 ( .B(clk), .A(\g.we_clk [12625]));
Q_ASSIGN U3766 ( .B(clk), .A(\g.we_clk [12624]));
Q_ASSIGN U3767 ( .B(clk), .A(\g.we_clk [12623]));
Q_ASSIGN U3768 ( .B(clk), .A(\g.we_clk [12622]));
Q_ASSIGN U3769 ( .B(clk), .A(\g.we_clk [12621]));
Q_ASSIGN U3770 ( .B(clk), .A(\g.we_clk [12620]));
Q_ASSIGN U3771 ( .B(clk), .A(\g.we_clk [12619]));
Q_ASSIGN U3772 ( .B(clk), .A(\g.we_clk [12618]));
Q_ASSIGN U3773 ( .B(clk), .A(\g.we_clk [12617]));
Q_ASSIGN U3774 ( .B(clk), .A(\g.we_clk [12616]));
Q_ASSIGN U3775 ( .B(clk), .A(\g.we_clk [12615]));
Q_ASSIGN U3776 ( .B(clk), .A(\g.we_clk [12614]));
Q_ASSIGN U3777 ( .B(clk), .A(\g.we_clk [12613]));
Q_ASSIGN U3778 ( .B(clk), .A(\g.we_clk [12612]));
Q_ASSIGN U3779 ( .B(clk), .A(\g.we_clk [12611]));
Q_ASSIGN U3780 ( .B(clk), .A(\g.we_clk [12610]));
Q_ASSIGN U3781 ( .B(clk), .A(\g.we_clk [12609]));
Q_ASSIGN U3782 ( .B(clk), .A(\g.we_clk [12608]));
Q_ASSIGN U3783 ( .B(clk), .A(\g.we_clk [12607]));
Q_ASSIGN U3784 ( .B(clk), .A(\g.we_clk [12606]));
Q_ASSIGN U3785 ( .B(clk), .A(\g.we_clk [12605]));
Q_ASSIGN U3786 ( .B(clk), .A(\g.we_clk [12604]));
Q_ASSIGN U3787 ( .B(clk), .A(\g.we_clk [12603]));
Q_ASSIGN U3788 ( .B(clk), .A(\g.we_clk [12602]));
Q_ASSIGN U3789 ( .B(clk), .A(\g.we_clk [12601]));
Q_ASSIGN U3790 ( .B(clk), .A(\g.we_clk [12600]));
Q_ASSIGN U3791 ( .B(clk), .A(\g.we_clk [12599]));
Q_ASSIGN U3792 ( .B(clk), .A(\g.we_clk [12598]));
Q_ASSIGN U3793 ( .B(clk), .A(\g.we_clk [12597]));
Q_ASSIGN U3794 ( .B(clk), .A(\g.we_clk [12596]));
Q_ASSIGN U3795 ( .B(clk), .A(\g.we_clk [12595]));
Q_ASSIGN U3796 ( .B(clk), .A(\g.we_clk [12594]));
Q_ASSIGN U3797 ( .B(clk), .A(\g.we_clk [12593]));
Q_ASSIGN U3798 ( .B(clk), .A(\g.we_clk [12592]));
Q_ASSIGN U3799 ( .B(clk), .A(\g.we_clk [12591]));
Q_ASSIGN U3800 ( .B(clk), .A(\g.we_clk [12590]));
Q_ASSIGN U3801 ( .B(clk), .A(\g.we_clk [12589]));
Q_ASSIGN U3802 ( .B(clk), .A(\g.we_clk [12588]));
Q_ASSIGN U3803 ( .B(clk), .A(\g.we_clk [12587]));
Q_ASSIGN U3804 ( .B(clk), .A(\g.we_clk [12586]));
Q_ASSIGN U3805 ( .B(clk), .A(\g.we_clk [12585]));
Q_ASSIGN U3806 ( .B(clk), .A(\g.we_clk [12584]));
Q_ASSIGN U3807 ( .B(clk), .A(\g.we_clk [12583]));
Q_ASSIGN U3808 ( .B(clk), .A(\g.we_clk [12582]));
Q_ASSIGN U3809 ( .B(clk), .A(\g.we_clk [12581]));
Q_ASSIGN U3810 ( .B(clk), .A(\g.we_clk [12580]));
Q_ASSIGN U3811 ( .B(clk), .A(\g.we_clk [12579]));
Q_ASSIGN U3812 ( .B(clk), .A(\g.we_clk [12578]));
Q_ASSIGN U3813 ( .B(clk), .A(\g.we_clk [12577]));
Q_ASSIGN U3814 ( .B(clk), .A(\g.we_clk [12576]));
Q_ASSIGN U3815 ( .B(clk), .A(\g.we_clk [12575]));
Q_ASSIGN U3816 ( .B(clk), .A(\g.we_clk [12574]));
Q_ASSIGN U3817 ( .B(clk), .A(\g.we_clk [12573]));
Q_ASSIGN U3818 ( .B(clk), .A(\g.we_clk [12572]));
Q_ASSIGN U3819 ( .B(clk), .A(\g.we_clk [12571]));
Q_ASSIGN U3820 ( .B(clk), .A(\g.we_clk [12570]));
Q_ASSIGN U3821 ( .B(clk), .A(\g.we_clk [12569]));
Q_ASSIGN U3822 ( .B(clk), .A(\g.we_clk [12568]));
Q_ASSIGN U3823 ( .B(clk), .A(\g.we_clk [12567]));
Q_ASSIGN U3824 ( .B(clk), .A(\g.we_clk [12566]));
Q_ASSIGN U3825 ( .B(clk), .A(\g.we_clk [12565]));
Q_ASSIGN U3826 ( .B(clk), .A(\g.we_clk [12564]));
Q_ASSIGN U3827 ( .B(clk), .A(\g.we_clk [12563]));
Q_ASSIGN U3828 ( .B(clk), .A(\g.we_clk [12562]));
Q_ASSIGN U3829 ( .B(clk), .A(\g.we_clk [12561]));
Q_ASSIGN U3830 ( .B(clk), .A(\g.we_clk [12560]));
Q_ASSIGN U3831 ( .B(clk), .A(\g.we_clk [12559]));
Q_ASSIGN U3832 ( .B(clk), .A(\g.we_clk [12558]));
Q_ASSIGN U3833 ( .B(clk), .A(\g.we_clk [12557]));
Q_ASSIGN U3834 ( .B(clk), .A(\g.we_clk [12556]));
Q_ASSIGN U3835 ( .B(clk), .A(\g.we_clk [12555]));
Q_ASSIGN U3836 ( .B(clk), .A(\g.we_clk [12554]));
Q_ASSIGN U3837 ( .B(clk), .A(\g.we_clk [12553]));
Q_ASSIGN U3838 ( .B(clk), .A(\g.we_clk [12552]));
Q_ASSIGN U3839 ( .B(clk), .A(\g.we_clk [12551]));
Q_ASSIGN U3840 ( .B(clk), .A(\g.we_clk [12550]));
Q_ASSIGN U3841 ( .B(clk), .A(\g.we_clk [12549]));
Q_ASSIGN U3842 ( .B(clk), .A(\g.we_clk [12548]));
Q_ASSIGN U3843 ( .B(clk), .A(\g.we_clk [12547]));
Q_ASSIGN U3844 ( .B(clk), .A(\g.we_clk [12546]));
Q_ASSIGN U3845 ( .B(clk), .A(\g.we_clk [12545]));
Q_ASSIGN U3846 ( .B(clk), .A(\g.we_clk [12544]));
Q_ASSIGN U3847 ( .B(clk), .A(\g.we_clk [12543]));
Q_ASSIGN U3848 ( .B(clk), .A(\g.we_clk [12542]));
Q_ASSIGN U3849 ( .B(clk), .A(\g.we_clk [12541]));
Q_ASSIGN U3850 ( .B(clk), .A(\g.we_clk [12540]));
Q_ASSIGN U3851 ( .B(clk), .A(\g.we_clk [12539]));
Q_ASSIGN U3852 ( .B(clk), .A(\g.we_clk [12538]));
Q_ASSIGN U3853 ( .B(clk), .A(\g.we_clk [12537]));
Q_ASSIGN U3854 ( .B(clk), .A(\g.we_clk [12536]));
Q_ASSIGN U3855 ( .B(clk), .A(\g.we_clk [12535]));
Q_ASSIGN U3856 ( .B(clk), .A(\g.we_clk [12534]));
Q_ASSIGN U3857 ( .B(clk), .A(\g.we_clk [12533]));
Q_ASSIGN U3858 ( .B(clk), .A(\g.we_clk [12532]));
Q_ASSIGN U3859 ( .B(clk), .A(\g.we_clk [12531]));
Q_ASSIGN U3860 ( .B(clk), .A(\g.we_clk [12530]));
Q_ASSIGN U3861 ( .B(clk), .A(\g.we_clk [12529]));
Q_ASSIGN U3862 ( .B(clk), .A(\g.we_clk [12528]));
Q_ASSIGN U3863 ( .B(clk), .A(\g.we_clk [12527]));
Q_ASSIGN U3864 ( .B(clk), .A(\g.we_clk [12526]));
Q_ASSIGN U3865 ( .B(clk), .A(\g.we_clk [12525]));
Q_ASSIGN U3866 ( .B(clk), .A(\g.we_clk [12524]));
Q_ASSIGN U3867 ( .B(clk), .A(\g.we_clk [12523]));
Q_ASSIGN U3868 ( .B(clk), .A(\g.we_clk [12522]));
Q_ASSIGN U3869 ( .B(clk), .A(\g.we_clk [12521]));
Q_ASSIGN U3870 ( .B(clk), .A(\g.we_clk [12520]));
Q_ASSIGN U3871 ( .B(clk), .A(\g.we_clk [12519]));
Q_ASSIGN U3872 ( .B(clk), .A(\g.we_clk [12518]));
Q_ASSIGN U3873 ( .B(clk), .A(\g.we_clk [12517]));
Q_ASSIGN U3874 ( .B(clk), .A(\g.we_clk [12516]));
Q_ASSIGN U3875 ( .B(clk), .A(\g.we_clk [12515]));
Q_ASSIGN U3876 ( .B(clk), .A(\g.we_clk [12514]));
Q_ASSIGN U3877 ( .B(clk), .A(\g.we_clk [12513]));
Q_ASSIGN U3878 ( .B(clk), .A(\g.we_clk [12512]));
Q_ASSIGN U3879 ( .B(clk), .A(\g.we_clk [12511]));
Q_ASSIGN U3880 ( .B(clk), .A(\g.we_clk [12510]));
Q_ASSIGN U3881 ( .B(clk), .A(\g.we_clk [12509]));
Q_ASSIGN U3882 ( .B(clk), .A(\g.we_clk [12508]));
Q_ASSIGN U3883 ( .B(clk), .A(\g.we_clk [12507]));
Q_ASSIGN U3884 ( .B(clk), .A(\g.we_clk [12506]));
Q_ASSIGN U3885 ( .B(clk), .A(\g.we_clk [12505]));
Q_ASSIGN U3886 ( .B(clk), .A(\g.we_clk [12504]));
Q_ASSIGN U3887 ( .B(clk), .A(\g.we_clk [12503]));
Q_ASSIGN U3888 ( .B(clk), .A(\g.we_clk [12502]));
Q_ASSIGN U3889 ( .B(clk), .A(\g.we_clk [12501]));
Q_ASSIGN U3890 ( .B(clk), .A(\g.we_clk [12500]));
Q_ASSIGN U3891 ( .B(clk), .A(\g.we_clk [12499]));
Q_ASSIGN U3892 ( .B(clk), .A(\g.we_clk [12498]));
Q_ASSIGN U3893 ( .B(clk), .A(\g.we_clk [12497]));
Q_ASSIGN U3894 ( .B(clk), .A(\g.we_clk [12496]));
Q_ASSIGN U3895 ( .B(clk), .A(\g.we_clk [12495]));
Q_ASSIGN U3896 ( .B(clk), .A(\g.we_clk [12494]));
Q_ASSIGN U3897 ( .B(clk), .A(\g.we_clk [12493]));
Q_ASSIGN U3898 ( .B(clk), .A(\g.we_clk [12492]));
Q_ASSIGN U3899 ( .B(clk), .A(\g.we_clk [12491]));
Q_ASSIGN U3900 ( .B(clk), .A(\g.we_clk [12490]));
Q_ASSIGN U3901 ( .B(clk), .A(\g.we_clk [12489]));
Q_ASSIGN U3902 ( .B(clk), .A(\g.we_clk [12488]));
Q_ASSIGN U3903 ( .B(clk), .A(\g.we_clk [12487]));
Q_ASSIGN U3904 ( .B(clk), .A(\g.we_clk [12486]));
Q_ASSIGN U3905 ( .B(clk), .A(\g.we_clk [12485]));
Q_ASSIGN U3906 ( .B(clk), .A(\g.we_clk [12484]));
Q_ASSIGN U3907 ( .B(clk), .A(\g.we_clk [12483]));
Q_ASSIGN U3908 ( .B(clk), .A(\g.we_clk [12482]));
Q_ASSIGN U3909 ( .B(clk), .A(\g.we_clk [12481]));
Q_ASSIGN U3910 ( .B(clk), .A(\g.we_clk [12480]));
Q_ASSIGN U3911 ( .B(clk), .A(\g.we_clk [12479]));
Q_ASSIGN U3912 ( .B(clk), .A(\g.we_clk [12478]));
Q_ASSIGN U3913 ( .B(clk), .A(\g.we_clk [12477]));
Q_ASSIGN U3914 ( .B(clk), .A(\g.we_clk [12476]));
Q_ASSIGN U3915 ( .B(clk), .A(\g.we_clk [12475]));
Q_ASSIGN U3916 ( .B(clk), .A(\g.we_clk [12474]));
Q_ASSIGN U3917 ( .B(clk), .A(\g.we_clk [12473]));
Q_ASSIGN U3918 ( .B(clk), .A(\g.we_clk [12472]));
Q_ASSIGN U3919 ( .B(clk), .A(\g.we_clk [12471]));
Q_ASSIGN U3920 ( .B(clk), .A(\g.we_clk [12470]));
Q_ASSIGN U3921 ( .B(clk), .A(\g.we_clk [12469]));
Q_ASSIGN U3922 ( .B(clk), .A(\g.we_clk [12468]));
Q_ASSIGN U3923 ( .B(clk), .A(\g.we_clk [12467]));
Q_ASSIGN U3924 ( .B(clk), .A(\g.we_clk [12466]));
Q_ASSIGN U3925 ( .B(clk), .A(\g.we_clk [12465]));
Q_ASSIGN U3926 ( .B(clk), .A(\g.we_clk [12464]));
Q_ASSIGN U3927 ( .B(clk), .A(\g.we_clk [12463]));
Q_ASSIGN U3928 ( .B(clk), .A(\g.we_clk [12462]));
Q_ASSIGN U3929 ( .B(clk), .A(\g.we_clk [12461]));
Q_ASSIGN U3930 ( .B(clk), .A(\g.we_clk [12460]));
Q_ASSIGN U3931 ( .B(clk), .A(\g.we_clk [12459]));
Q_ASSIGN U3932 ( .B(clk), .A(\g.we_clk [12458]));
Q_ASSIGN U3933 ( .B(clk), .A(\g.we_clk [12457]));
Q_ASSIGN U3934 ( .B(clk), .A(\g.we_clk [12456]));
Q_ASSIGN U3935 ( .B(clk), .A(\g.we_clk [12455]));
Q_ASSIGN U3936 ( .B(clk), .A(\g.we_clk [12454]));
Q_ASSIGN U3937 ( .B(clk), .A(\g.we_clk [12453]));
Q_ASSIGN U3938 ( .B(clk), .A(\g.we_clk [12452]));
Q_ASSIGN U3939 ( .B(clk), .A(\g.we_clk [12451]));
Q_ASSIGN U3940 ( .B(clk), .A(\g.we_clk [12450]));
Q_ASSIGN U3941 ( .B(clk), .A(\g.we_clk [12449]));
Q_ASSIGN U3942 ( .B(clk), .A(\g.we_clk [12448]));
Q_ASSIGN U3943 ( .B(clk), .A(\g.we_clk [12447]));
Q_ASSIGN U3944 ( .B(clk), .A(\g.we_clk [12446]));
Q_ASSIGN U3945 ( .B(clk), .A(\g.we_clk [12445]));
Q_ASSIGN U3946 ( .B(clk), .A(\g.we_clk [12444]));
Q_ASSIGN U3947 ( .B(clk), .A(\g.we_clk [12443]));
Q_ASSIGN U3948 ( .B(clk), .A(\g.we_clk [12442]));
Q_ASSIGN U3949 ( .B(clk), .A(\g.we_clk [12441]));
Q_ASSIGN U3950 ( .B(clk), .A(\g.we_clk [12440]));
Q_ASSIGN U3951 ( .B(clk), .A(\g.we_clk [12439]));
Q_ASSIGN U3952 ( .B(clk), .A(\g.we_clk [12438]));
Q_ASSIGN U3953 ( .B(clk), .A(\g.we_clk [12437]));
Q_ASSIGN U3954 ( .B(clk), .A(\g.we_clk [12436]));
Q_ASSIGN U3955 ( .B(clk), .A(\g.we_clk [12435]));
Q_ASSIGN U3956 ( .B(clk), .A(\g.we_clk [12434]));
Q_ASSIGN U3957 ( .B(clk), .A(\g.we_clk [12433]));
Q_ASSIGN U3958 ( .B(clk), .A(\g.we_clk [12432]));
Q_ASSIGN U3959 ( .B(clk), .A(\g.we_clk [12431]));
Q_ASSIGN U3960 ( .B(clk), .A(\g.we_clk [12430]));
Q_ASSIGN U3961 ( .B(clk), .A(\g.we_clk [12429]));
Q_ASSIGN U3962 ( .B(clk), .A(\g.we_clk [12428]));
Q_ASSIGN U3963 ( .B(clk), .A(\g.we_clk [12427]));
Q_ASSIGN U3964 ( .B(clk), .A(\g.we_clk [12426]));
Q_ASSIGN U3965 ( .B(clk), .A(\g.we_clk [12425]));
Q_ASSIGN U3966 ( .B(clk), .A(\g.we_clk [12424]));
Q_ASSIGN U3967 ( .B(clk), .A(\g.we_clk [12423]));
Q_ASSIGN U3968 ( .B(clk), .A(\g.we_clk [12422]));
Q_ASSIGN U3969 ( .B(clk), .A(\g.we_clk [12421]));
Q_ASSIGN U3970 ( .B(clk), .A(\g.we_clk [12420]));
Q_ASSIGN U3971 ( .B(clk), .A(\g.we_clk [12419]));
Q_ASSIGN U3972 ( .B(clk), .A(\g.we_clk [12418]));
Q_ASSIGN U3973 ( .B(clk), .A(\g.we_clk [12417]));
Q_ASSIGN U3974 ( .B(clk), .A(\g.we_clk [12416]));
Q_ASSIGN U3975 ( .B(clk), .A(\g.we_clk [12415]));
Q_ASSIGN U3976 ( .B(clk), .A(\g.we_clk [12414]));
Q_ASSIGN U3977 ( .B(clk), .A(\g.we_clk [12413]));
Q_ASSIGN U3978 ( .B(clk), .A(\g.we_clk [12412]));
Q_ASSIGN U3979 ( .B(clk), .A(\g.we_clk [12411]));
Q_ASSIGN U3980 ( .B(clk), .A(\g.we_clk [12410]));
Q_ASSIGN U3981 ( .B(clk), .A(\g.we_clk [12409]));
Q_ASSIGN U3982 ( .B(clk), .A(\g.we_clk [12408]));
Q_ASSIGN U3983 ( .B(clk), .A(\g.we_clk [12407]));
Q_ASSIGN U3984 ( .B(clk), .A(\g.we_clk [12406]));
Q_ASSIGN U3985 ( .B(clk), .A(\g.we_clk [12405]));
Q_ASSIGN U3986 ( .B(clk), .A(\g.we_clk [12404]));
Q_ASSIGN U3987 ( .B(clk), .A(\g.we_clk [12403]));
Q_ASSIGN U3988 ( .B(clk), .A(\g.we_clk [12402]));
Q_ASSIGN U3989 ( .B(clk), .A(\g.we_clk [12401]));
Q_ASSIGN U3990 ( .B(clk), .A(\g.we_clk [12400]));
Q_ASSIGN U3991 ( .B(clk), .A(\g.we_clk [12399]));
Q_ASSIGN U3992 ( .B(clk), .A(\g.we_clk [12398]));
Q_ASSIGN U3993 ( .B(clk), .A(\g.we_clk [12397]));
Q_ASSIGN U3994 ( .B(clk), .A(\g.we_clk [12396]));
Q_ASSIGN U3995 ( .B(clk), .A(\g.we_clk [12395]));
Q_ASSIGN U3996 ( .B(clk), .A(\g.we_clk [12394]));
Q_ASSIGN U3997 ( .B(clk), .A(\g.we_clk [12393]));
Q_ASSIGN U3998 ( .B(clk), .A(\g.we_clk [12392]));
Q_ASSIGN U3999 ( .B(clk), .A(\g.we_clk [12391]));
Q_ASSIGN U4000 ( .B(clk), .A(\g.we_clk [12390]));
Q_ASSIGN U4001 ( .B(clk), .A(\g.we_clk [12389]));
Q_ASSIGN U4002 ( .B(clk), .A(\g.we_clk [12388]));
Q_ASSIGN U4003 ( .B(clk), .A(\g.we_clk [12387]));
Q_ASSIGN U4004 ( .B(clk), .A(\g.we_clk [12386]));
Q_ASSIGN U4005 ( .B(clk), .A(\g.we_clk [12385]));
Q_ASSIGN U4006 ( .B(clk), .A(\g.we_clk [12384]));
Q_ASSIGN U4007 ( .B(clk), .A(\g.we_clk [12383]));
Q_ASSIGN U4008 ( .B(clk), .A(\g.we_clk [12382]));
Q_ASSIGN U4009 ( .B(clk), .A(\g.we_clk [12381]));
Q_ASSIGN U4010 ( .B(clk), .A(\g.we_clk [12380]));
Q_ASSIGN U4011 ( .B(clk), .A(\g.we_clk [12379]));
Q_ASSIGN U4012 ( .B(clk), .A(\g.we_clk [12378]));
Q_ASSIGN U4013 ( .B(clk), .A(\g.we_clk [12377]));
Q_ASSIGN U4014 ( .B(clk), .A(\g.we_clk [12376]));
Q_ASSIGN U4015 ( .B(clk), .A(\g.we_clk [12375]));
Q_ASSIGN U4016 ( .B(clk), .A(\g.we_clk [12374]));
Q_ASSIGN U4017 ( .B(clk), .A(\g.we_clk [12373]));
Q_ASSIGN U4018 ( .B(clk), .A(\g.we_clk [12372]));
Q_ASSIGN U4019 ( .B(clk), .A(\g.we_clk [12371]));
Q_ASSIGN U4020 ( .B(clk), .A(\g.we_clk [12370]));
Q_ASSIGN U4021 ( .B(clk), .A(\g.we_clk [12369]));
Q_ASSIGN U4022 ( .B(clk), .A(\g.we_clk [12368]));
Q_ASSIGN U4023 ( .B(clk), .A(\g.we_clk [12367]));
Q_ASSIGN U4024 ( .B(clk), .A(\g.we_clk [12366]));
Q_ASSIGN U4025 ( .B(clk), .A(\g.we_clk [12365]));
Q_ASSIGN U4026 ( .B(clk), .A(\g.we_clk [12364]));
Q_ASSIGN U4027 ( .B(clk), .A(\g.we_clk [12363]));
Q_ASSIGN U4028 ( .B(clk), .A(\g.we_clk [12362]));
Q_ASSIGN U4029 ( .B(clk), .A(\g.we_clk [12361]));
Q_ASSIGN U4030 ( .B(clk), .A(\g.we_clk [12360]));
Q_ASSIGN U4031 ( .B(clk), .A(\g.we_clk [12359]));
Q_ASSIGN U4032 ( .B(clk), .A(\g.we_clk [12358]));
Q_ASSIGN U4033 ( .B(clk), .A(\g.we_clk [12357]));
Q_ASSIGN U4034 ( .B(clk), .A(\g.we_clk [12356]));
Q_ASSIGN U4035 ( .B(clk), .A(\g.we_clk [12355]));
Q_ASSIGN U4036 ( .B(clk), .A(\g.we_clk [12354]));
Q_ASSIGN U4037 ( .B(clk), .A(\g.we_clk [12353]));
Q_ASSIGN U4038 ( .B(clk), .A(\g.we_clk [12352]));
Q_ASSIGN U4039 ( .B(clk), .A(\g.we_clk [12351]));
Q_ASSIGN U4040 ( .B(clk), .A(\g.we_clk [12350]));
Q_ASSIGN U4041 ( .B(clk), .A(\g.we_clk [12349]));
Q_ASSIGN U4042 ( .B(clk), .A(\g.we_clk [12348]));
Q_ASSIGN U4043 ( .B(clk), .A(\g.we_clk [12347]));
Q_ASSIGN U4044 ( .B(clk), .A(\g.we_clk [12346]));
Q_ASSIGN U4045 ( .B(clk), .A(\g.we_clk [12345]));
Q_ASSIGN U4046 ( .B(clk), .A(\g.we_clk [12344]));
Q_ASSIGN U4047 ( .B(clk), .A(\g.we_clk [12343]));
Q_ASSIGN U4048 ( .B(clk), .A(\g.we_clk [12342]));
Q_ASSIGN U4049 ( .B(clk), .A(\g.we_clk [12341]));
Q_ASSIGN U4050 ( .B(clk), .A(\g.we_clk [12340]));
Q_ASSIGN U4051 ( .B(clk), .A(\g.we_clk [12339]));
Q_ASSIGN U4052 ( .B(clk), .A(\g.we_clk [12338]));
Q_ASSIGN U4053 ( .B(clk), .A(\g.we_clk [12337]));
Q_ASSIGN U4054 ( .B(clk), .A(\g.we_clk [12336]));
Q_ASSIGN U4055 ( .B(clk), .A(\g.we_clk [12335]));
Q_ASSIGN U4056 ( .B(clk), .A(\g.we_clk [12334]));
Q_ASSIGN U4057 ( .B(clk), .A(\g.we_clk [12333]));
Q_ASSIGN U4058 ( .B(clk), .A(\g.we_clk [12332]));
Q_ASSIGN U4059 ( .B(clk), .A(\g.we_clk [12331]));
Q_ASSIGN U4060 ( .B(clk), .A(\g.we_clk [12330]));
Q_ASSIGN U4061 ( .B(clk), .A(\g.we_clk [12329]));
Q_ASSIGN U4062 ( .B(clk), .A(\g.we_clk [12328]));
Q_ASSIGN U4063 ( .B(clk), .A(\g.we_clk [12327]));
Q_ASSIGN U4064 ( .B(clk), .A(\g.we_clk [12326]));
Q_ASSIGN U4065 ( .B(clk), .A(\g.we_clk [12325]));
Q_ASSIGN U4066 ( .B(clk), .A(\g.we_clk [12324]));
Q_ASSIGN U4067 ( .B(clk), .A(\g.we_clk [12323]));
Q_ASSIGN U4068 ( .B(clk), .A(\g.we_clk [12322]));
Q_ASSIGN U4069 ( .B(clk), .A(\g.we_clk [12321]));
Q_ASSIGN U4070 ( .B(clk), .A(\g.we_clk [12320]));
Q_ASSIGN U4071 ( .B(clk), .A(\g.we_clk [12319]));
Q_ASSIGN U4072 ( .B(clk), .A(\g.we_clk [12318]));
Q_ASSIGN U4073 ( .B(clk), .A(\g.we_clk [12317]));
Q_ASSIGN U4074 ( .B(clk), .A(\g.we_clk [12316]));
Q_ASSIGN U4075 ( .B(clk), .A(\g.we_clk [12315]));
Q_ASSIGN U4076 ( .B(clk), .A(\g.we_clk [12314]));
Q_ASSIGN U4077 ( .B(clk), .A(\g.we_clk [12313]));
Q_ASSIGN U4078 ( .B(clk), .A(\g.we_clk [12312]));
Q_ASSIGN U4079 ( .B(clk), .A(\g.we_clk [12311]));
Q_ASSIGN U4080 ( .B(clk), .A(\g.we_clk [12310]));
Q_ASSIGN U4081 ( .B(clk), .A(\g.we_clk [12309]));
Q_ASSIGN U4082 ( .B(clk), .A(\g.we_clk [12308]));
Q_ASSIGN U4083 ( .B(clk), .A(\g.we_clk [12307]));
Q_ASSIGN U4084 ( .B(clk), .A(\g.we_clk [12306]));
Q_ASSIGN U4085 ( .B(clk), .A(\g.we_clk [12305]));
Q_ASSIGN U4086 ( .B(clk), .A(\g.we_clk [12304]));
Q_ASSIGN U4087 ( .B(clk), .A(\g.we_clk [12303]));
Q_ASSIGN U4088 ( .B(clk), .A(\g.we_clk [12302]));
Q_ASSIGN U4089 ( .B(clk), .A(\g.we_clk [12301]));
Q_ASSIGN U4090 ( .B(clk), .A(\g.we_clk [12300]));
Q_ASSIGN U4091 ( .B(clk), .A(\g.we_clk [12299]));
Q_ASSIGN U4092 ( .B(clk), .A(\g.we_clk [12298]));
Q_ASSIGN U4093 ( .B(clk), .A(\g.we_clk [12297]));
Q_ASSIGN U4094 ( .B(clk), .A(\g.we_clk [12296]));
Q_ASSIGN U4095 ( .B(clk), .A(\g.we_clk [12295]));
Q_ASSIGN U4096 ( .B(clk), .A(\g.we_clk [12294]));
Q_ASSIGN U4097 ( .B(clk), .A(\g.we_clk [12293]));
Q_ASSIGN U4098 ( .B(clk), .A(\g.we_clk [12292]));
Q_ASSIGN U4099 ( .B(clk), .A(\g.we_clk [12291]));
Q_ASSIGN U4100 ( .B(clk), .A(\g.we_clk [12290]));
Q_ASSIGN U4101 ( .B(clk), .A(\g.we_clk [12289]));
Q_ASSIGN U4102 ( .B(clk), .A(\g.we_clk [12288]));
Q_ASSIGN U4103 ( .B(clk), .A(\g.we_clk [12287]));
Q_ASSIGN U4104 ( .B(clk), .A(\g.we_clk [12286]));
Q_ASSIGN U4105 ( .B(clk), .A(\g.we_clk [12285]));
Q_ASSIGN U4106 ( .B(clk), .A(\g.we_clk [12284]));
Q_ASSIGN U4107 ( .B(clk), .A(\g.we_clk [12283]));
Q_ASSIGN U4108 ( .B(clk), .A(\g.we_clk [12282]));
Q_ASSIGN U4109 ( .B(clk), .A(\g.we_clk [12281]));
Q_ASSIGN U4110 ( .B(clk), .A(\g.we_clk [12280]));
Q_ASSIGN U4111 ( .B(clk), .A(\g.we_clk [12279]));
Q_ASSIGN U4112 ( .B(clk), .A(\g.we_clk [12278]));
Q_ASSIGN U4113 ( .B(clk), .A(\g.we_clk [12277]));
Q_ASSIGN U4114 ( .B(clk), .A(\g.we_clk [12276]));
Q_ASSIGN U4115 ( .B(clk), .A(\g.we_clk [12275]));
Q_ASSIGN U4116 ( .B(clk), .A(\g.we_clk [12274]));
Q_ASSIGN U4117 ( .B(clk), .A(\g.we_clk [12273]));
Q_ASSIGN U4118 ( .B(clk), .A(\g.we_clk [12272]));
Q_ASSIGN U4119 ( .B(clk), .A(\g.we_clk [12271]));
Q_ASSIGN U4120 ( .B(clk), .A(\g.we_clk [12270]));
Q_ASSIGN U4121 ( .B(clk), .A(\g.we_clk [12269]));
Q_ASSIGN U4122 ( .B(clk), .A(\g.we_clk [12268]));
Q_ASSIGN U4123 ( .B(clk), .A(\g.we_clk [12267]));
Q_ASSIGN U4124 ( .B(clk), .A(\g.we_clk [12266]));
Q_ASSIGN U4125 ( .B(clk), .A(\g.we_clk [12265]));
Q_ASSIGN U4126 ( .B(clk), .A(\g.we_clk [12264]));
Q_ASSIGN U4127 ( .B(clk), .A(\g.we_clk [12263]));
Q_ASSIGN U4128 ( .B(clk), .A(\g.we_clk [12262]));
Q_ASSIGN U4129 ( .B(clk), .A(\g.we_clk [12261]));
Q_ASSIGN U4130 ( .B(clk), .A(\g.we_clk [12260]));
Q_ASSIGN U4131 ( .B(clk), .A(\g.we_clk [12259]));
Q_ASSIGN U4132 ( .B(clk), .A(\g.we_clk [12258]));
Q_ASSIGN U4133 ( .B(clk), .A(\g.we_clk [12257]));
Q_ASSIGN U4134 ( .B(clk), .A(\g.we_clk [12256]));
Q_ASSIGN U4135 ( .B(clk), .A(\g.we_clk [12255]));
Q_ASSIGN U4136 ( .B(clk), .A(\g.we_clk [12254]));
Q_ASSIGN U4137 ( .B(clk), .A(\g.we_clk [12253]));
Q_ASSIGN U4138 ( .B(clk), .A(\g.we_clk [12252]));
Q_ASSIGN U4139 ( .B(clk), .A(\g.we_clk [12251]));
Q_ASSIGN U4140 ( .B(clk), .A(\g.we_clk [12250]));
Q_ASSIGN U4141 ( .B(clk), .A(\g.we_clk [12249]));
Q_ASSIGN U4142 ( .B(clk), .A(\g.we_clk [12248]));
Q_ASSIGN U4143 ( .B(clk), .A(\g.we_clk [12247]));
Q_ASSIGN U4144 ( .B(clk), .A(\g.we_clk [12246]));
Q_ASSIGN U4145 ( .B(clk), .A(\g.we_clk [12245]));
Q_ASSIGN U4146 ( .B(clk), .A(\g.we_clk [12244]));
Q_ASSIGN U4147 ( .B(clk), .A(\g.we_clk [12243]));
Q_ASSIGN U4148 ( .B(clk), .A(\g.we_clk [12242]));
Q_ASSIGN U4149 ( .B(clk), .A(\g.we_clk [12241]));
Q_ASSIGN U4150 ( .B(clk), .A(\g.we_clk [12240]));
Q_ASSIGN U4151 ( .B(clk), .A(\g.we_clk [12239]));
Q_ASSIGN U4152 ( .B(clk), .A(\g.we_clk [12238]));
Q_ASSIGN U4153 ( .B(clk), .A(\g.we_clk [12237]));
Q_ASSIGN U4154 ( .B(clk), .A(\g.we_clk [12236]));
Q_ASSIGN U4155 ( .B(clk), .A(\g.we_clk [12235]));
Q_ASSIGN U4156 ( .B(clk), .A(\g.we_clk [12234]));
Q_ASSIGN U4157 ( .B(clk), .A(\g.we_clk [12233]));
Q_ASSIGN U4158 ( .B(clk), .A(\g.we_clk [12232]));
Q_ASSIGN U4159 ( .B(clk), .A(\g.we_clk [12231]));
Q_ASSIGN U4160 ( .B(clk), .A(\g.we_clk [12230]));
Q_ASSIGN U4161 ( .B(clk), .A(\g.we_clk [12229]));
Q_ASSIGN U4162 ( .B(clk), .A(\g.we_clk [12228]));
Q_ASSIGN U4163 ( .B(clk), .A(\g.we_clk [12227]));
Q_ASSIGN U4164 ( .B(clk), .A(\g.we_clk [12226]));
Q_ASSIGN U4165 ( .B(clk), .A(\g.we_clk [12225]));
Q_ASSIGN U4166 ( .B(clk), .A(\g.we_clk [12224]));
Q_ASSIGN U4167 ( .B(clk), .A(\g.we_clk [12223]));
Q_ASSIGN U4168 ( .B(clk), .A(\g.we_clk [12222]));
Q_ASSIGN U4169 ( .B(clk), .A(\g.we_clk [12221]));
Q_ASSIGN U4170 ( .B(clk), .A(\g.we_clk [12220]));
Q_ASSIGN U4171 ( .B(clk), .A(\g.we_clk [12219]));
Q_ASSIGN U4172 ( .B(clk), .A(\g.we_clk [12218]));
Q_ASSIGN U4173 ( .B(clk), .A(\g.we_clk [12217]));
Q_ASSIGN U4174 ( .B(clk), .A(\g.we_clk [12216]));
Q_ASSIGN U4175 ( .B(clk), .A(\g.we_clk [12215]));
Q_ASSIGN U4176 ( .B(clk), .A(\g.we_clk [12214]));
Q_ASSIGN U4177 ( .B(clk), .A(\g.we_clk [12213]));
Q_ASSIGN U4178 ( .B(clk), .A(\g.we_clk [12212]));
Q_ASSIGN U4179 ( .B(clk), .A(\g.we_clk [12211]));
Q_ASSIGN U4180 ( .B(clk), .A(\g.we_clk [12210]));
Q_ASSIGN U4181 ( .B(clk), .A(\g.we_clk [12209]));
Q_ASSIGN U4182 ( .B(clk), .A(\g.we_clk [12208]));
Q_ASSIGN U4183 ( .B(clk), .A(\g.we_clk [12207]));
Q_ASSIGN U4184 ( .B(clk), .A(\g.we_clk [12206]));
Q_ASSIGN U4185 ( .B(clk), .A(\g.we_clk [12205]));
Q_ASSIGN U4186 ( .B(clk), .A(\g.we_clk [12204]));
Q_ASSIGN U4187 ( .B(clk), .A(\g.we_clk [12203]));
Q_ASSIGN U4188 ( .B(clk), .A(\g.we_clk [12202]));
Q_ASSIGN U4189 ( .B(clk), .A(\g.we_clk [12201]));
Q_ASSIGN U4190 ( .B(clk), .A(\g.we_clk [12200]));
Q_ASSIGN U4191 ( .B(clk), .A(\g.we_clk [12199]));
Q_ASSIGN U4192 ( .B(clk), .A(\g.we_clk [12198]));
Q_ASSIGN U4193 ( .B(clk), .A(\g.we_clk [12197]));
Q_ASSIGN U4194 ( .B(clk), .A(\g.we_clk [12196]));
Q_ASSIGN U4195 ( .B(clk), .A(\g.we_clk [12195]));
Q_ASSIGN U4196 ( .B(clk), .A(\g.we_clk [12194]));
Q_ASSIGN U4197 ( .B(clk), .A(\g.we_clk [12193]));
Q_ASSIGN U4198 ( .B(clk), .A(\g.we_clk [12192]));
Q_ASSIGN U4199 ( .B(clk), .A(\g.we_clk [12191]));
Q_ASSIGN U4200 ( .B(clk), .A(\g.we_clk [12190]));
Q_ASSIGN U4201 ( .B(clk), .A(\g.we_clk [12189]));
Q_ASSIGN U4202 ( .B(clk), .A(\g.we_clk [12188]));
Q_ASSIGN U4203 ( .B(clk), .A(\g.we_clk [12187]));
Q_ASSIGN U4204 ( .B(clk), .A(\g.we_clk [12186]));
Q_ASSIGN U4205 ( .B(clk), .A(\g.we_clk [12185]));
Q_ASSIGN U4206 ( .B(clk), .A(\g.we_clk [12184]));
Q_ASSIGN U4207 ( .B(clk), .A(\g.we_clk [12183]));
Q_ASSIGN U4208 ( .B(clk), .A(\g.we_clk [12182]));
Q_ASSIGN U4209 ( .B(clk), .A(\g.we_clk [12181]));
Q_ASSIGN U4210 ( .B(clk), .A(\g.we_clk [12180]));
Q_ASSIGN U4211 ( .B(clk), .A(\g.we_clk [12179]));
Q_ASSIGN U4212 ( .B(clk), .A(\g.we_clk [12178]));
Q_ASSIGN U4213 ( .B(clk), .A(\g.we_clk [12177]));
Q_ASSIGN U4214 ( .B(clk), .A(\g.we_clk [12176]));
Q_ASSIGN U4215 ( .B(clk), .A(\g.we_clk [12175]));
Q_ASSIGN U4216 ( .B(clk), .A(\g.we_clk [12174]));
Q_ASSIGN U4217 ( .B(clk), .A(\g.we_clk [12173]));
Q_ASSIGN U4218 ( .B(clk), .A(\g.we_clk [12172]));
Q_ASSIGN U4219 ( .B(clk), .A(\g.we_clk [12171]));
Q_ASSIGN U4220 ( .B(clk), .A(\g.we_clk [12170]));
Q_ASSIGN U4221 ( .B(clk), .A(\g.we_clk [12169]));
Q_ASSIGN U4222 ( .B(clk), .A(\g.we_clk [12168]));
Q_ASSIGN U4223 ( .B(clk), .A(\g.we_clk [12167]));
Q_ASSIGN U4224 ( .B(clk), .A(\g.we_clk [12166]));
Q_ASSIGN U4225 ( .B(clk), .A(\g.we_clk [12165]));
Q_ASSIGN U4226 ( .B(clk), .A(\g.we_clk [12164]));
Q_ASSIGN U4227 ( .B(clk), .A(\g.we_clk [12163]));
Q_ASSIGN U4228 ( .B(clk), .A(\g.we_clk [12162]));
Q_ASSIGN U4229 ( .B(clk), .A(\g.we_clk [12161]));
Q_ASSIGN U4230 ( .B(clk), .A(\g.we_clk [12160]));
Q_ASSIGN U4231 ( .B(clk), .A(\g.we_clk [12159]));
Q_ASSIGN U4232 ( .B(clk), .A(\g.we_clk [12158]));
Q_ASSIGN U4233 ( .B(clk), .A(\g.we_clk [12157]));
Q_ASSIGN U4234 ( .B(clk), .A(\g.we_clk [12156]));
Q_ASSIGN U4235 ( .B(clk), .A(\g.we_clk [12155]));
Q_ASSIGN U4236 ( .B(clk), .A(\g.we_clk [12154]));
Q_ASSIGN U4237 ( .B(clk), .A(\g.we_clk [12153]));
Q_ASSIGN U4238 ( .B(clk), .A(\g.we_clk [12152]));
Q_ASSIGN U4239 ( .B(clk), .A(\g.we_clk [12151]));
Q_ASSIGN U4240 ( .B(clk), .A(\g.we_clk [12150]));
Q_ASSIGN U4241 ( .B(clk), .A(\g.we_clk [12149]));
Q_ASSIGN U4242 ( .B(clk), .A(\g.we_clk [12148]));
Q_ASSIGN U4243 ( .B(clk), .A(\g.we_clk [12147]));
Q_ASSIGN U4244 ( .B(clk), .A(\g.we_clk [12146]));
Q_ASSIGN U4245 ( .B(clk), .A(\g.we_clk [12145]));
Q_ASSIGN U4246 ( .B(clk), .A(\g.we_clk [12144]));
Q_ASSIGN U4247 ( .B(clk), .A(\g.we_clk [12143]));
Q_ASSIGN U4248 ( .B(clk), .A(\g.we_clk [12142]));
Q_ASSIGN U4249 ( .B(clk), .A(\g.we_clk [12141]));
Q_ASSIGN U4250 ( .B(clk), .A(\g.we_clk [12140]));
Q_ASSIGN U4251 ( .B(clk), .A(\g.we_clk [12139]));
Q_ASSIGN U4252 ( .B(clk), .A(\g.we_clk [12138]));
Q_ASSIGN U4253 ( .B(clk), .A(\g.we_clk [12137]));
Q_ASSIGN U4254 ( .B(clk), .A(\g.we_clk [12136]));
Q_ASSIGN U4255 ( .B(clk), .A(\g.we_clk [12135]));
Q_ASSIGN U4256 ( .B(clk), .A(\g.we_clk [12134]));
Q_ASSIGN U4257 ( .B(clk), .A(\g.we_clk [12133]));
Q_ASSIGN U4258 ( .B(clk), .A(\g.we_clk [12132]));
Q_ASSIGN U4259 ( .B(clk), .A(\g.we_clk [12131]));
Q_ASSIGN U4260 ( .B(clk), .A(\g.we_clk [12130]));
Q_ASSIGN U4261 ( .B(clk), .A(\g.we_clk [12129]));
Q_ASSIGN U4262 ( .B(clk), .A(\g.we_clk [12128]));
Q_ASSIGN U4263 ( .B(clk), .A(\g.we_clk [12127]));
Q_ASSIGN U4264 ( .B(clk), .A(\g.we_clk [12126]));
Q_ASSIGN U4265 ( .B(clk), .A(\g.we_clk [12125]));
Q_ASSIGN U4266 ( .B(clk), .A(\g.we_clk [12124]));
Q_ASSIGN U4267 ( .B(clk), .A(\g.we_clk [12123]));
Q_ASSIGN U4268 ( .B(clk), .A(\g.we_clk [12122]));
Q_ASSIGN U4269 ( .B(clk), .A(\g.we_clk [12121]));
Q_ASSIGN U4270 ( .B(clk), .A(\g.we_clk [12120]));
Q_ASSIGN U4271 ( .B(clk), .A(\g.we_clk [12119]));
Q_ASSIGN U4272 ( .B(clk), .A(\g.we_clk [12118]));
Q_ASSIGN U4273 ( .B(clk), .A(\g.we_clk [12117]));
Q_ASSIGN U4274 ( .B(clk), .A(\g.we_clk [12116]));
Q_ASSIGN U4275 ( .B(clk), .A(\g.we_clk [12115]));
Q_ASSIGN U4276 ( .B(clk), .A(\g.we_clk [12114]));
Q_ASSIGN U4277 ( .B(clk), .A(\g.we_clk [12113]));
Q_ASSIGN U4278 ( .B(clk), .A(\g.we_clk [12112]));
Q_ASSIGN U4279 ( .B(clk), .A(\g.we_clk [12111]));
Q_ASSIGN U4280 ( .B(clk), .A(\g.we_clk [12110]));
Q_ASSIGN U4281 ( .B(clk), .A(\g.we_clk [12109]));
Q_ASSIGN U4282 ( .B(clk), .A(\g.we_clk [12108]));
Q_ASSIGN U4283 ( .B(clk), .A(\g.we_clk [12107]));
Q_ASSIGN U4284 ( .B(clk), .A(\g.we_clk [12106]));
Q_ASSIGN U4285 ( .B(clk), .A(\g.we_clk [12105]));
Q_ASSIGN U4286 ( .B(clk), .A(\g.we_clk [12104]));
Q_ASSIGN U4287 ( .B(clk), .A(\g.we_clk [12103]));
Q_ASSIGN U4288 ( .B(clk), .A(\g.we_clk [12102]));
Q_ASSIGN U4289 ( .B(clk), .A(\g.we_clk [12101]));
Q_ASSIGN U4290 ( .B(clk), .A(\g.we_clk [12100]));
Q_ASSIGN U4291 ( .B(clk), .A(\g.we_clk [12099]));
Q_ASSIGN U4292 ( .B(clk), .A(\g.we_clk [12098]));
Q_ASSIGN U4293 ( .B(clk), .A(\g.we_clk [12097]));
Q_ASSIGN U4294 ( .B(clk), .A(\g.we_clk [12096]));
Q_ASSIGN U4295 ( .B(clk), .A(\g.we_clk [12095]));
Q_ASSIGN U4296 ( .B(clk), .A(\g.we_clk [12094]));
Q_ASSIGN U4297 ( .B(clk), .A(\g.we_clk [12093]));
Q_ASSIGN U4298 ( .B(clk), .A(\g.we_clk [12092]));
Q_ASSIGN U4299 ( .B(clk), .A(\g.we_clk [12091]));
Q_ASSIGN U4300 ( .B(clk), .A(\g.we_clk [12090]));
Q_ASSIGN U4301 ( .B(clk), .A(\g.we_clk [12089]));
Q_ASSIGN U4302 ( .B(clk), .A(\g.we_clk [12088]));
Q_ASSIGN U4303 ( .B(clk), .A(\g.we_clk [12087]));
Q_ASSIGN U4304 ( .B(clk), .A(\g.we_clk [12086]));
Q_ASSIGN U4305 ( .B(clk), .A(\g.we_clk [12085]));
Q_ASSIGN U4306 ( .B(clk), .A(\g.we_clk [12084]));
Q_ASSIGN U4307 ( .B(clk), .A(\g.we_clk [12083]));
Q_ASSIGN U4308 ( .B(clk), .A(\g.we_clk [12082]));
Q_ASSIGN U4309 ( .B(clk), .A(\g.we_clk [12081]));
Q_ASSIGN U4310 ( .B(clk), .A(\g.we_clk [12080]));
Q_ASSIGN U4311 ( .B(clk), .A(\g.we_clk [12079]));
Q_ASSIGN U4312 ( .B(clk), .A(\g.we_clk [12078]));
Q_ASSIGN U4313 ( .B(clk), .A(\g.we_clk [12077]));
Q_ASSIGN U4314 ( .B(clk), .A(\g.we_clk [12076]));
Q_ASSIGN U4315 ( .B(clk), .A(\g.we_clk [12075]));
Q_ASSIGN U4316 ( .B(clk), .A(\g.we_clk [12074]));
Q_ASSIGN U4317 ( .B(clk), .A(\g.we_clk [12073]));
Q_ASSIGN U4318 ( .B(clk), .A(\g.we_clk [12072]));
Q_ASSIGN U4319 ( .B(clk), .A(\g.we_clk [12071]));
Q_ASSIGN U4320 ( .B(clk), .A(\g.we_clk [12070]));
Q_ASSIGN U4321 ( .B(clk), .A(\g.we_clk [12069]));
Q_ASSIGN U4322 ( .B(clk), .A(\g.we_clk [12068]));
Q_ASSIGN U4323 ( .B(clk), .A(\g.we_clk [12067]));
Q_ASSIGN U4324 ( .B(clk), .A(\g.we_clk [12066]));
Q_ASSIGN U4325 ( .B(clk), .A(\g.we_clk [12065]));
Q_ASSIGN U4326 ( .B(clk), .A(\g.we_clk [12064]));
Q_ASSIGN U4327 ( .B(clk), .A(\g.we_clk [12063]));
Q_ASSIGN U4328 ( .B(clk), .A(\g.we_clk [12062]));
Q_ASSIGN U4329 ( .B(clk), .A(\g.we_clk [12061]));
Q_ASSIGN U4330 ( .B(clk), .A(\g.we_clk [12060]));
Q_ASSIGN U4331 ( .B(clk), .A(\g.we_clk [12059]));
Q_ASSIGN U4332 ( .B(clk), .A(\g.we_clk [12058]));
Q_ASSIGN U4333 ( .B(clk), .A(\g.we_clk [12057]));
Q_ASSIGN U4334 ( .B(clk), .A(\g.we_clk [12056]));
Q_ASSIGN U4335 ( .B(clk), .A(\g.we_clk [12055]));
Q_ASSIGN U4336 ( .B(clk), .A(\g.we_clk [12054]));
Q_ASSIGN U4337 ( .B(clk), .A(\g.we_clk [12053]));
Q_ASSIGN U4338 ( .B(clk), .A(\g.we_clk [12052]));
Q_ASSIGN U4339 ( .B(clk), .A(\g.we_clk [12051]));
Q_ASSIGN U4340 ( .B(clk), .A(\g.we_clk [12050]));
Q_ASSIGN U4341 ( .B(clk), .A(\g.we_clk [12049]));
Q_ASSIGN U4342 ( .B(clk), .A(\g.we_clk [12048]));
Q_ASSIGN U4343 ( .B(clk), .A(\g.we_clk [12047]));
Q_ASSIGN U4344 ( .B(clk), .A(\g.we_clk [12046]));
Q_ASSIGN U4345 ( .B(clk), .A(\g.we_clk [12045]));
Q_ASSIGN U4346 ( .B(clk), .A(\g.we_clk [12044]));
Q_ASSIGN U4347 ( .B(clk), .A(\g.we_clk [12043]));
Q_ASSIGN U4348 ( .B(clk), .A(\g.we_clk [12042]));
Q_ASSIGN U4349 ( .B(clk), .A(\g.we_clk [12041]));
Q_ASSIGN U4350 ( .B(clk), .A(\g.we_clk [12040]));
Q_ASSIGN U4351 ( .B(clk), .A(\g.we_clk [12039]));
Q_ASSIGN U4352 ( .B(clk), .A(\g.we_clk [12038]));
Q_ASSIGN U4353 ( .B(clk), .A(\g.we_clk [12037]));
Q_ASSIGN U4354 ( .B(clk), .A(\g.we_clk [12036]));
Q_ASSIGN U4355 ( .B(clk), .A(\g.we_clk [12035]));
Q_ASSIGN U4356 ( .B(clk), .A(\g.we_clk [12034]));
Q_ASSIGN U4357 ( .B(clk), .A(\g.we_clk [12033]));
Q_ASSIGN U4358 ( .B(clk), .A(\g.we_clk [12032]));
Q_ASSIGN U4359 ( .B(clk), .A(\g.we_clk [12031]));
Q_ASSIGN U4360 ( .B(clk), .A(\g.we_clk [12030]));
Q_ASSIGN U4361 ( .B(clk), .A(\g.we_clk [12029]));
Q_ASSIGN U4362 ( .B(clk), .A(\g.we_clk [12028]));
Q_ASSIGN U4363 ( .B(clk), .A(\g.we_clk [12027]));
Q_ASSIGN U4364 ( .B(clk), .A(\g.we_clk [12026]));
Q_ASSIGN U4365 ( .B(clk), .A(\g.we_clk [12025]));
Q_ASSIGN U4366 ( .B(clk), .A(\g.we_clk [12024]));
Q_ASSIGN U4367 ( .B(clk), .A(\g.we_clk [12023]));
Q_ASSIGN U4368 ( .B(clk), .A(\g.we_clk [12022]));
Q_ASSIGN U4369 ( .B(clk), .A(\g.we_clk [12021]));
Q_ASSIGN U4370 ( .B(clk), .A(\g.we_clk [12020]));
Q_ASSIGN U4371 ( .B(clk), .A(\g.we_clk [12019]));
Q_ASSIGN U4372 ( .B(clk), .A(\g.we_clk [12018]));
Q_ASSIGN U4373 ( .B(clk), .A(\g.we_clk [12017]));
Q_ASSIGN U4374 ( .B(clk), .A(\g.we_clk [12016]));
Q_ASSIGN U4375 ( .B(clk), .A(\g.we_clk [12015]));
Q_ASSIGN U4376 ( .B(clk), .A(\g.we_clk [12014]));
Q_ASSIGN U4377 ( .B(clk), .A(\g.we_clk [12013]));
Q_ASSIGN U4378 ( .B(clk), .A(\g.we_clk [12012]));
Q_ASSIGN U4379 ( .B(clk), .A(\g.we_clk [12011]));
Q_ASSIGN U4380 ( .B(clk), .A(\g.we_clk [12010]));
Q_ASSIGN U4381 ( .B(clk), .A(\g.we_clk [12009]));
Q_ASSIGN U4382 ( .B(clk), .A(\g.we_clk [12008]));
Q_ASSIGN U4383 ( .B(clk), .A(\g.we_clk [12007]));
Q_ASSIGN U4384 ( .B(clk), .A(\g.we_clk [12006]));
Q_ASSIGN U4385 ( .B(clk), .A(\g.we_clk [12005]));
Q_ASSIGN U4386 ( .B(clk), .A(\g.we_clk [12004]));
Q_ASSIGN U4387 ( .B(clk), .A(\g.we_clk [12003]));
Q_ASSIGN U4388 ( .B(clk), .A(\g.we_clk [12002]));
Q_ASSIGN U4389 ( .B(clk), .A(\g.we_clk [12001]));
Q_ASSIGN U4390 ( .B(clk), .A(\g.we_clk [12000]));
Q_ASSIGN U4391 ( .B(clk), .A(\g.we_clk [11999]));
Q_ASSIGN U4392 ( .B(clk), .A(\g.we_clk [11998]));
Q_ASSIGN U4393 ( .B(clk), .A(\g.we_clk [11997]));
Q_ASSIGN U4394 ( .B(clk), .A(\g.we_clk [11996]));
Q_ASSIGN U4395 ( .B(clk), .A(\g.we_clk [11995]));
Q_ASSIGN U4396 ( .B(clk), .A(\g.we_clk [11994]));
Q_ASSIGN U4397 ( .B(clk), .A(\g.we_clk [11993]));
Q_ASSIGN U4398 ( .B(clk), .A(\g.we_clk [11992]));
Q_ASSIGN U4399 ( .B(clk), .A(\g.we_clk [11991]));
Q_ASSIGN U4400 ( .B(clk), .A(\g.we_clk [11990]));
Q_ASSIGN U4401 ( .B(clk), .A(\g.we_clk [11989]));
Q_ASSIGN U4402 ( .B(clk), .A(\g.we_clk [11988]));
Q_ASSIGN U4403 ( .B(clk), .A(\g.we_clk [11987]));
Q_ASSIGN U4404 ( .B(clk), .A(\g.we_clk [11986]));
Q_ASSIGN U4405 ( .B(clk), .A(\g.we_clk [11985]));
Q_ASSIGN U4406 ( .B(clk), .A(\g.we_clk [11984]));
Q_ASSIGN U4407 ( .B(clk), .A(\g.we_clk [11983]));
Q_ASSIGN U4408 ( .B(clk), .A(\g.we_clk [11982]));
Q_ASSIGN U4409 ( .B(clk), .A(\g.we_clk [11981]));
Q_ASSIGN U4410 ( .B(clk), .A(\g.we_clk [11980]));
Q_ASSIGN U4411 ( .B(clk), .A(\g.we_clk [11979]));
Q_ASSIGN U4412 ( .B(clk), .A(\g.we_clk [11978]));
Q_ASSIGN U4413 ( .B(clk), .A(\g.we_clk [11977]));
Q_ASSIGN U4414 ( .B(clk), .A(\g.we_clk [11976]));
Q_ASSIGN U4415 ( .B(clk), .A(\g.we_clk [11975]));
Q_ASSIGN U4416 ( .B(clk), .A(\g.we_clk [11974]));
Q_ASSIGN U4417 ( .B(clk), .A(\g.we_clk [11973]));
Q_ASSIGN U4418 ( .B(clk), .A(\g.we_clk [11972]));
Q_ASSIGN U4419 ( .B(clk), .A(\g.we_clk [11971]));
Q_ASSIGN U4420 ( .B(clk), .A(\g.we_clk [11970]));
Q_ASSIGN U4421 ( .B(clk), .A(\g.we_clk [11969]));
Q_ASSIGN U4422 ( .B(clk), .A(\g.we_clk [11968]));
Q_ASSIGN U4423 ( .B(clk), .A(\g.we_clk [11967]));
Q_ASSIGN U4424 ( .B(clk), .A(\g.we_clk [11966]));
Q_ASSIGN U4425 ( .B(clk), .A(\g.we_clk [11965]));
Q_ASSIGN U4426 ( .B(clk), .A(\g.we_clk [11964]));
Q_ASSIGN U4427 ( .B(clk), .A(\g.we_clk [11963]));
Q_ASSIGN U4428 ( .B(clk), .A(\g.we_clk [11962]));
Q_ASSIGN U4429 ( .B(clk), .A(\g.we_clk [11961]));
Q_ASSIGN U4430 ( .B(clk), .A(\g.we_clk [11960]));
Q_ASSIGN U4431 ( .B(clk), .A(\g.we_clk [11959]));
Q_ASSIGN U4432 ( .B(clk), .A(\g.we_clk [11958]));
Q_ASSIGN U4433 ( .B(clk), .A(\g.we_clk [11957]));
Q_ASSIGN U4434 ( .B(clk), .A(\g.we_clk [11956]));
Q_ASSIGN U4435 ( .B(clk), .A(\g.we_clk [11955]));
Q_ASSIGN U4436 ( .B(clk), .A(\g.we_clk [11954]));
Q_ASSIGN U4437 ( .B(clk), .A(\g.we_clk [11953]));
Q_ASSIGN U4438 ( .B(clk), .A(\g.we_clk [11952]));
Q_ASSIGN U4439 ( .B(clk), .A(\g.we_clk [11951]));
Q_ASSIGN U4440 ( .B(clk), .A(\g.we_clk [11950]));
Q_ASSIGN U4441 ( .B(clk), .A(\g.we_clk [11949]));
Q_ASSIGN U4442 ( .B(clk), .A(\g.we_clk [11948]));
Q_ASSIGN U4443 ( .B(clk), .A(\g.we_clk [11947]));
Q_ASSIGN U4444 ( .B(clk), .A(\g.we_clk [11946]));
Q_ASSIGN U4445 ( .B(clk), .A(\g.we_clk [11945]));
Q_ASSIGN U4446 ( .B(clk), .A(\g.we_clk [11944]));
Q_ASSIGN U4447 ( .B(clk), .A(\g.we_clk [11943]));
Q_ASSIGN U4448 ( .B(clk), .A(\g.we_clk [11942]));
Q_ASSIGN U4449 ( .B(clk), .A(\g.we_clk [11941]));
Q_ASSIGN U4450 ( .B(clk), .A(\g.we_clk [11940]));
Q_ASSIGN U4451 ( .B(clk), .A(\g.we_clk [11939]));
Q_ASSIGN U4452 ( .B(clk), .A(\g.we_clk [11938]));
Q_ASSIGN U4453 ( .B(clk), .A(\g.we_clk [11937]));
Q_ASSIGN U4454 ( .B(clk), .A(\g.we_clk [11936]));
Q_ASSIGN U4455 ( .B(clk), .A(\g.we_clk [11935]));
Q_ASSIGN U4456 ( .B(clk), .A(\g.we_clk [11934]));
Q_ASSIGN U4457 ( .B(clk), .A(\g.we_clk [11933]));
Q_ASSIGN U4458 ( .B(clk), .A(\g.we_clk [11932]));
Q_ASSIGN U4459 ( .B(clk), .A(\g.we_clk [11931]));
Q_ASSIGN U4460 ( .B(clk), .A(\g.we_clk [11930]));
Q_ASSIGN U4461 ( .B(clk), .A(\g.we_clk [11929]));
Q_ASSIGN U4462 ( .B(clk), .A(\g.we_clk [11928]));
Q_ASSIGN U4463 ( .B(clk), .A(\g.we_clk [11927]));
Q_ASSIGN U4464 ( .B(clk), .A(\g.we_clk [11926]));
Q_ASSIGN U4465 ( .B(clk), .A(\g.we_clk [11925]));
Q_ASSIGN U4466 ( .B(clk), .A(\g.we_clk [11924]));
Q_ASSIGN U4467 ( .B(clk), .A(\g.we_clk [11923]));
Q_ASSIGN U4468 ( .B(clk), .A(\g.we_clk [11922]));
Q_ASSIGN U4469 ( .B(clk), .A(\g.we_clk [11921]));
Q_ASSIGN U4470 ( .B(clk), .A(\g.we_clk [11920]));
Q_ASSIGN U4471 ( .B(clk), .A(\g.we_clk [11919]));
Q_ASSIGN U4472 ( .B(clk), .A(\g.we_clk [11918]));
Q_ASSIGN U4473 ( .B(clk), .A(\g.we_clk [11917]));
Q_ASSIGN U4474 ( .B(clk), .A(\g.we_clk [11916]));
Q_ASSIGN U4475 ( .B(clk), .A(\g.we_clk [11915]));
Q_ASSIGN U4476 ( .B(clk), .A(\g.we_clk [11914]));
Q_ASSIGN U4477 ( .B(clk), .A(\g.we_clk [11913]));
Q_ASSIGN U4478 ( .B(clk), .A(\g.we_clk [11912]));
Q_ASSIGN U4479 ( .B(clk), .A(\g.we_clk [11911]));
Q_ASSIGN U4480 ( .B(clk), .A(\g.we_clk [11910]));
Q_ASSIGN U4481 ( .B(clk), .A(\g.we_clk [11909]));
Q_ASSIGN U4482 ( .B(clk), .A(\g.we_clk [11908]));
Q_ASSIGN U4483 ( .B(clk), .A(\g.we_clk [11907]));
Q_ASSIGN U4484 ( .B(clk), .A(\g.we_clk [11906]));
Q_ASSIGN U4485 ( .B(clk), .A(\g.we_clk [11905]));
Q_ASSIGN U4486 ( .B(clk), .A(\g.we_clk [11904]));
Q_ASSIGN U4487 ( .B(clk), .A(\g.we_clk [11903]));
Q_ASSIGN U4488 ( .B(clk), .A(\g.we_clk [11902]));
Q_ASSIGN U4489 ( .B(clk), .A(\g.we_clk [11901]));
Q_ASSIGN U4490 ( .B(clk), .A(\g.we_clk [11900]));
Q_ASSIGN U4491 ( .B(clk), .A(\g.we_clk [11899]));
Q_ASSIGN U4492 ( .B(clk), .A(\g.we_clk [11898]));
Q_ASSIGN U4493 ( .B(clk), .A(\g.we_clk [11897]));
Q_ASSIGN U4494 ( .B(clk), .A(\g.we_clk [11896]));
Q_ASSIGN U4495 ( .B(clk), .A(\g.we_clk [11895]));
Q_ASSIGN U4496 ( .B(clk), .A(\g.we_clk [11894]));
Q_ASSIGN U4497 ( .B(clk), .A(\g.we_clk [11893]));
Q_ASSIGN U4498 ( .B(clk), .A(\g.we_clk [11892]));
Q_ASSIGN U4499 ( .B(clk), .A(\g.we_clk [11891]));
Q_ASSIGN U4500 ( .B(clk), .A(\g.we_clk [11890]));
Q_ASSIGN U4501 ( .B(clk), .A(\g.we_clk [11889]));
Q_ASSIGN U4502 ( .B(clk), .A(\g.we_clk [11888]));
Q_ASSIGN U4503 ( .B(clk), .A(\g.we_clk [11887]));
Q_ASSIGN U4504 ( .B(clk), .A(\g.we_clk [11886]));
Q_ASSIGN U4505 ( .B(clk), .A(\g.we_clk [11885]));
Q_ASSIGN U4506 ( .B(clk), .A(\g.we_clk [11884]));
Q_ASSIGN U4507 ( .B(clk), .A(\g.we_clk [11883]));
Q_ASSIGN U4508 ( .B(clk), .A(\g.we_clk [11882]));
Q_ASSIGN U4509 ( .B(clk), .A(\g.we_clk [11881]));
Q_ASSIGN U4510 ( .B(clk), .A(\g.we_clk [11880]));
Q_ASSIGN U4511 ( .B(clk), .A(\g.we_clk [11879]));
Q_ASSIGN U4512 ( .B(clk), .A(\g.we_clk [11878]));
Q_ASSIGN U4513 ( .B(clk), .A(\g.we_clk [11877]));
Q_ASSIGN U4514 ( .B(clk), .A(\g.we_clk [11876]));
Q_ASSIGN U4515 ( .B(clk), .A(\g.we_clk [11875]));
Q_ASSIGN U4516 ( .B(clk), .A(\g.we_clk [11874]));
Q_ASSIGN U4517 ( .B(clk), .A(\g.we_clk [11873]));
Q_ASSIGN U4518 ( .B(clk), .A(\g.we_clk [11872]));
Q_ASSIGN U4519 ( .B(clk), .A(\g.we_clk [11871]));
Q_ASSIGN U4520 ( .B(clk), .A(\g.we_clk [11870]));
Q_ASSIGN U4521 ( .B(clk), .A(\g.we_clk [11869]));
Q_ASSIGN U4522 ( .B(clk), .A(\g.we_clk [11868]));
Q_ASSIGN U4523 ( .B(clk), .A(\g.we_clk [11867]));
Q_ASSIGN U4524 ( .B(clk), .A(\g.we_clk [11866]));
Q_ASSIGN U4525 ( .B(clk), .A(\g.we_clk [11865]));
Q_ASSIGN U4526 ( .B(clk), .A(\g.we_clk [11864]));
Q_ASSIGN U4527 ( .B(clk), .A(\g.we_clk [11863]));
Q_ASSIGN U4528 ( .B(clk), .A(\g.we_clk [11862]));
Q_ASSIGN U4529 ( .B(clk), .A(\g.we_clk [11861]));
Q_ASSIGN U4530 ( .B(clk), .A(\g.we_clk [11860]));
Q_ASSIGN U4531 ( .B(clk), .A(\g.we_clk [11859]));
Q_ASSIGN U4532 ( .B(clk), .A(\g.we_clk [11858]));
Q_ASSIGN U4533 ( .B(clk), .A(\g.we_clk [11857]));
Q_ASSIGN U4534 ( .B(clk), .A(\g.we_clk [11856]));
Q_ASSIGN U4535 ( .B(clk), .A(\g.we_clk [11855]));
Q_ASSIGN U4536 ( .B(clk), .A(\g.we_clk [11854]));
Q_ASSIGN U4537 ( .B(clk), .A(\g.we_clk [11853]));
Q_ASSIGN U4538 ( .B(clk), .A(\g.we_clk [11852]));
Q_ASSIGN U4539 ( .B(clk), .A(\g.we_clk [11851]));
Q_ASSIGN U4540 ( .B(clk), .A(\g.we_clk [11850]));
Q_ASSIGN U4541 ( .B(clk), .A(\g.we_clk [11849]));
Q_ASSIGN U4542 ( .B(clk), .A(\g.we_clk [11848]));
Q_ASSIGN U4543 ( .B(clk), .A(\g.we_clk [11847]));
Q_ASSIGN U4544 ( .B(clk), .A(\g.we_clk [11846]));
Q_ASSIGN U4545 ( .B(clk), .A(\g.we_clk [11845]));
Q_ASSIGN U4546 ( .B(clk), .A(\g.we_clk [11844]));
Q_ASSIGN U4547 ( .B(clk), .A(\g.we_clk [11843]));
Q_ASSIGN U4548 ( .B(clk), .A(\g.we_clk [11842]));
Q_ASSIGN U4549 ( .B(clk), .A(\g.we_clk [11841]));
Q_ASSIGN U4550 ( .B(clk), .A(\g.we_clk [11840]));
Q_ASSIGN U4551 ( .B(clk), .A(\g.we_clk [11839]));
Q_ASSIGN U4552 ( .B(clk), .A(\g.we_clk [11838]));
Q_ASSIGN U4553 ( .B(clk), .A(\g.we_clk [11837]));
Q_ASSIGN U4554 ( .B(clk), .A(\g.we_clk [11836]));
Q_ASSIGN U4555 ( .B(clk), .A(\g.we_clk [11835]));
Q_ASSIGN U4556 ( .B(clk), .A(\g.we_clk [11834]));
Q_ASSIGN U4557 ( .B(clk), .A(\g.we_clk [11833]));
Q_ASSIGN U4558 ( .B(clk), .A(\g.we_clk [11832]));
Q_ASSIGN U4559 ( .B(clk), .A(\g.we_clk [11831]));
Q_ASSIGN U4560 ( .B(clk), .A(\g.we_clk [11830]));
Q_ASSIGN U4561 ( .B(clk), .A(\g.we_clk [11829]));
Q_ASSIGN U4562 ( .B(clk), .A(\g.we_clk [11828]));
Q_ASSIGN U4563 ( .B(clk), .A(\g.we_clk [11827]));
Q_ASSIGN U4564 ( .B(clk), .A(\g.we_clk [11826]));
Q_ASSIGN U4565 ( .B(clk), .A(\g.we_clk [11825]));
Q_ASSIGN U4566 ( .B(clk), .A(\g.we_clk [11824]));
Q_ASSIGN U4567 ( .B(clk), .A(\g.we_clk [11823]));
Q_ASSIGN U4568 ( .B(clk), .A(\g.we_clk [11822]));
Q_ASSIGN U4569 ( .B(clk), .A(\g.we_clk [11821]));
Q_ASSIGN U4570 ( .B(clk), .A(\g.we_clk [11820]));
Q_ASSIGN U4571 ( .B(clk), .A(\g.we_clk [11819]));
Q_ASSIGN U4572 ( .B(clk), .A(\g.we_clk [11818]));
Q_ASSIGN U4573 ( .B(clk), .A(\g.we_clk [11817]));
Q_ASSIGN U4574 ( .B(clk), .A(\g.we_clk [11816]));
Q_ASSIGN U4575 ( .B(clk), .A(\g.we_clk [11815]));
Q_ASSIGN U4576 ( .B(clk), .A(\g.we_clk [11814]));
Q_ASSIGN U4577 ( .B(clk), .A(\g.we_clk [11813]));
Q_ASSIGN U4578 ( .B(clk), .A(\g.we_clk [11812]));
Q_ASSIGN U4579 ( .B(clk), .A(\g.we_clk [11811]));
Q_ASSIGN U4580 ( .B(clk), .A(\g.we_clk [11810]));
Q_ASSIGN U4581 ( .B(clk), .A(\g.we_clk [11809]));
Q_ASSIGN U4582 ( .B(clk), .A(\g.we_clk [11808]));
Q_ASSIGN U4583 ( .B(clk), .A(\g.we_clk [11807]));
Q_ASSIGN U4584 ( .B(clk), .A(\g.we_clk [11806]));
Q_ASSIGN U4585 ( .B(clk), .A(\g.we_clk [11805]));
Q_ASSIGN U4586 ( .B(clk), .A(\g.we_clk [11804]));
Q_ASSIGN U4587 ( .B(clk), .A(\g.we_clk [11803]));
Q_ASSIGN U4588 ( .B(clk), .A(\g.we_clk [11802]));
Q_ASSIGN U4589 ( .B(clk), .A(\g.we_clk [11801]));
Q_ASSIGN U4590 ( .B(clk), .A(\g.we_clk [11800]));
Q_ASSIGN U4591 ( .B(clk), .A(\g.we_clk [11799]));
Q_ASSIGN U4592 ( .B(clk), .A(\g.we_clk [11798]));
Q_ASSIGN U4593 ( .B(clk), .A(\g.we_clk [11797]));
Q_ASSIGN U4594 ( .B(clk), .A(\g.we_clk [11796]));
Q_ASSIGN U4595 ( .B(clk), .A(\g.we_clk [11795]));
Q_ASSIGN U4596 ( .B(clk), .A(\g.we_clk [11794]));
Q_ASSIGN U4597 ( .B(clk), .A(\g.we_clk [11793]));
Q_ASSIGN U4598 ( .B(clk), .A(\g.we_clk [11792]));
Q_ASSIGN U4599 ( .B(clk), .A(\g.we_clk [11791]));
Q_ASSIGN U4600 ( .B(clk), .A(\g.we_clk [11790]));
Q_ASSIGN U4601 ( .B(clk), .A(\g.we_clk [11789]));
Q_ASSIGN U4602 ( .B(clk), .A(\g.we_clk [11788]));
Q_ASSIGN U4603 ( .B(clk), .A(\g.we_clk [11787]));
Q_ASSIGN U4604 ( .B(clk), .A(\g.we_clk [11786]));
Q_ASSIGN U4605 ( .B(clk), .A(\g.we_clk [11785]));
Q_ASSIGN U4606 ( .B(clk), .A(\g.we_clk [11784]));
Q_ASSIGN U4607 ( .B(clk), .A(\g.we_clk [11783]));
Q_ASSIGN U4608 ( .B(clk), .A(\g.we_clk [11782]));
Q_ASSIGN U4609 ( .B(clk), .A(\g.we_clk [11781]));
Q_ASSIGN U4610 ( .B(clk), .A(\g.we_clk [11780]));
Q_ASSIGN U4611 ( .B(clk), .A(\g.we_clk [11779]));
Q_ASSIGN U4612 ( .B(clk), .A(\g.we_clk [11778]));
Q_ASSIGN U4613 ( .B(clk), .A(\g.we_clk [11777]));
Q_ASSIGN U4614 ( .B(clk), .A(\g.we_clk [11776]));
Q_ASSIGN U4615 ( .B(clk), .A(\g.we_clk [11775]));
Q_ASSIGN U4616 ( .B(clk), .A(\g.we_clk [11774]));
Q_ASSIGN U4617 ( .B(clk), .A(\g.we_clk [11773]));
Q_ASSIGN U4618 ( .B(clk), .A(\g.we_clk [11772]));
Q_ASSIGN U4619 ( .B(clk), .A(\g.we_clk [11771]));
Q_ASSIGN U4620 ( .B(clk), .A(\g.we_clk [11770]));
Q_ASSIGN U4621 ( .B(clk), .A(\g.we_clk [11769]));
Q_ASSIGN U4622 ( .B(clk), .A(\g.we_clk [11768]));
Q_ASSIGN U4623 ( .B(clk), .A(\g.we_clk [11767]));
Q_ASSIGN U4624 ( .B(clk), .A(\g.we_clk [11766]));
Q_ASSIGN U4625 ( .B(clk), .A(\g.we_clk [11765]));
Q_ASSIGN U4626 ( .B(clk), .A(\g.we_clk [11764]));
Q_ASSIGN U4627 ( .B(clk), .A(\g.we_clk [11763]));
Q_ASSIGN U4628 ( .B(clk), .A(\g.we_clk [11762]));
Q_ASSIGN U4629 ( .B(clk), .A(\g.we_clk [11761]));
Q_ASSIGN U4630 ( .B(clk), .A(\g.we_clk [11760]));
Q_ASSIGN U4631 ( .B(clk), .A(\g.we_clk [11759]));
Q_ASSIGN U4632 ( .B(clk), .A(\g.we_clk [11758]));
Q_ASSIGN U4633 ( .B(clk), .A(\g.we_clk [11757]));
Q_ASSIGN U4634 ( .B(clk), .A(\g.we_clk [11756]));
Q_ASSIGN U4635 ( .B(clk), .A(\g.we_clk [11755]));
Q_ASSIGN U4636 ( .B(clk), .A(\g.we_clk [11754]));
Q_ASSIGN U4637 ( .B(clk), .A(\g.we_clk [11753]));
Q_ASSIGN U4638 ( .B(clk), .A(\g.we_clk [11752]));
Q_ASSIGN U4639 ( .B(clk), .A(\g.we_clk [11751]));
Q_ASSIGN U4640 ( .B(clk), .A(\g.we_clk [11750]));
Q_ASSIGN U4641 ( .B(clk), .A(\g.we_clk [11749]));
Q_ASSIGN U4642 ( .B(clk), .A(\g.we_clk [11748]));
Q_ASSIGN U4643 ( .B(clk), .A(\g.we_clk [11747]));
Q_ASSIGN U4644 ( .B(clk), .A(\g.we_clk [11746]));
Q_ASSIGN U4645 ( .B(clk), .A(\g.we_clk [11745]));
Q_ASSIGN U4646 ( .B(clk), .A(\g.we_clk [11744]));
Q_ASSIGN U4647 ( .B(clk), .A(\g.we_clk [11743]));
Q_ASSIGN U4648 ( .B(clk), .A(\g.we_clk [11742]));
Q_ASSIGN U4649 ( .B(clk), .A(\g.we_clk [11741]));
Q_ASSIGN U4650 ( .B(clk), .A(\g.we_clk [11740]));
Q_ASSIGN U4651 ( .B(clk), .A(\g.we_clk [11739]));
Q_ASSIGN U4652 ( .B(clk), .A(\g.we_clk [11738]));
Q_ASSIGN U4653 ( .B(clk), .A(\g.we_clk [11737]));
Q_ASSIGN U4654 ( .B(clk), .A(\g.we_clk [11736]));
Q_ASSIGN U4655 ( .B(clk), .A(\g.we_clk [11735]));
Q_ASSIGN U4656 ( .B(clk), .A(\g.we_clk [11734]));
Q_ASSIGN U4657 ( .B(clk), .A(\g.we_clk [11733]));
Q_ASSIGN U4658 ( .B(clk), .A(\g.we_clk [11732]));
Q_ASSIGN U4659 ( .B(clk), .A(\g.we_clk [11731]));
Q_ASSIGN U4660 ( .B(clk), .A(\g.we_clk [11730]));
Q_ASSIGN U4661 ( .B(clk), .A(\g.we_clk [11729]));
Q_ASSIGN U4662 ( .B(clk), .A(\g.we_clk [11728]));
Q_ASSIGN U4663 ( .B(clk), .A(\g.we_clk [11727]));
Q_ASSIGN U4664 ( .B(clk), .A(\g.we_clk [11726]));
Q_ASSIGN U4665 ( .B(clk), .A(\g.we_clk [11725]));
Q_ASSIGN U4666 ( .B(clk), .A(\g.we_clk [11724]));
Q_ASSIGN U4667 ( .B(clk), .A(\g.we_clk [11723]));
Q_ASSIGN U4668 ( .B(clk), .A(\g.we_clk [11722]));
Q_ASSIGN U4669 ( .B(clk), .A(\g.we_clk [11721]));
Q_ASSIGN U4670 ( .B(clk), .A(\g.we_clk [11720]));
Q_ASSIGN U4671 ( .B(clk), .A(\g.we_clk [11719]));
Q_ASSIGN U4672 ( .B(clk), .A(\g.we_clk [11718]));
Q_ASSIGN U4673 ( .B(clk), .A(\g.we_clk [11717]));
Q_ASSIGN U4674 ( .B(clk), .A(\g.we_clk [11716]));
Q_ASSIGN U4675 ( .B(clk), .A(\g.we_clk [11715]));
Q_ASSIGN U4676 ( .B(clk), .A(\g.we_clk [11714]));
Q_ASSIGN U4677 ( .B(clk), .A(\g.we_clk [11713]));
Q_ASSIGN U4678 ( .B(clk), .A(\g.we_clk [11712]));
Q_ASSIGN U4679 ( .B(clk), .A(\g.we_clk [11711]));
Q_ASSIGN U4680 ( .B(clk), .A(\g.we_clk [11710]));
Q_ASSIGN U4681 ( .B(clk), .A(\g.we_clk [11709]));
Q_ASSIGN U4682 ( .B(clk), .A(\g.we_clk [11708]));
Q_ASSIGN U4683 ( .B(clk), .A(\g.we_clk [11707]));
Q_ASSIGN U4684 ( .B(clk), .A(\g.we_clk [11706]));
Q_ASSIGN U4685 ( .B(clk), .A(\g.we_clk [11705]));
Q_ASSIGN U4686 ( .B(clk), .A(\g.we_clk [11704]));
Q_ASSIGN U4687 ( .B(clk), .A(\g.we_clk [11703]));
Q_ASSIGN U4688 ( .B(clk), .A(\g.we_clk [11702]));
Q_ASSIGN U4689 ( .B(clk), .A(\g.we_clk [11701]));
Q_ASSIGN U4690 ( .B(clk), .A(\g.we_clk [11700]));
Q_ASSIGN U4691 ( .B(clk), .A(\g.we_clk [11699]));
Q_ASSIGN U4692 ( .B(clk), .A(\g.we_clk [11698]));
Q_ASSIGN U4693 ( .B(clk), .A(\g.we_clk [11697]));
Q_ASSIGN U4694 ( .B(clk), .A(\g.we_clk [11696]));
Q_ASSIGN U4695 ( .B(clk), .A(\g.we_clk [11695]));
Q_ASSIGN U4696 ( .B(clk), .A(\g.we_clk [11694]));
Q_ASSIGN U4697 ( .B(clk), .A(\g.we_clk [11693]));
Q_ASSIGN U4698 ( .B(clk), .A(\g.we_clk [11692]));
Q_ASSIGN U4699 ( .B(clk), .A(\g.we_clk [11691]));
Q_ASSIGN U4700 ( .B(clk), .A(\g.we_clk [11690]));
Q_ASSIGN U4701 ( .B(clk), .A(\g.we_clk [11689]));
Q_ASSIGN U4702 ( .B(clk), .A(\g.we_clk [11688]));
Q_ASSIGN U4703 ( .B(clk), .A(\g.we_clk [11687]));
Q_ASSIGN U4704 ( .B(clk), .A(\g.we_clk [11686]));
Q_ASSIGN U4705 ( .B(clk), .A(\g.we_clk [11685]));
Q_ASSIGN U4706 ( .B(clk), .A(\g.we_clk [11684]));
Q_ASSIGN U4707 ( .B(clk), .A(\g.we_clk [11683]));
Q_ASSIGN U4708 ( .B(clk), .A(\g.we_clk [11682]));
Q_ASSIGN U4709 ( .B(clk), .A(\g.we_clk [11681]));
Q_ASSIGN U4710 ( .B(clk), .A(\g.we_clk [11680]));
Q_ASSIGN U4711 ( .B(clk), .A(\g.we_clk [11679]));
Q_ASSIGN U4712 ( .B(clk), .A(\g.we_clk [11678]));
Q_ASSIGN U4713 ( .B(clk), .A(\g.we_clk [11677]));
Q_ASSIGN U4714 ( .B(clk), .A(\g.we_clk [11676]));
Q_ASSIGN U4715 ( .B(clk), .A(\g.we_clk [11675]));
Q_ASSIGN U4716 ( .B(clk), .A(\g.we_clk [11674]));
Q_ASSIGN U4717 ( .B(clk), .A(\g.we_clk [11673]));
Q_ASSIGN U4718 ( .B(clk), .A(\g.we_clk [11672]));
Q_ASSIGN U4719 ( .B(clk), .A(\g.we_clk [11671]));
Q_ASSIGN U4720 ( .B(clk), .A(\g.we_clk [11670]));
Q_ASSIGN U4721 ( .B(clk), .A(\g.we_clk [11669]));
Q_ASSIGN U4722 ( .B(clk), .A(\g.we_clk [11668]));
Q_ASSIGN U4723 ( .B(clk), .A(\g.we_clk [11667]));
Q_ASSIGN U4724 ( .B(clk), .A(\g.we_clk [11666]));
Q_ASSIGN U4725 ( .B(clk), .A(\g.we_clk [11665]));
Q_ASSIGN U4726 ( .B(clk), .A(\g.we_clk [11664]));
Q_ASSIGN U4727 ( .B(clk), .A(\g.we_clk [11663]));
Q_ASSIGN U4728 ( .B(clk), .A(\g.we_clk [11662]));
Q_ASSIGN U4729 ( .B(clk), .A(\g.we_clk [11661]));
Q_ASSIGN U4730 ( .B(clk), .A(\g.we_clk [11660]));
Q_ASSIGN U4731 ( .B(clk), .A(\g.we_clk [11659]));
Q_ASSIGN U4732 ( .B(clk), .A(\g.we_clk [11658]));
Q_ASSIGN U4733 ( .B(clk), .A(\g.we_clk [11657]));
Q_ASSIGN U4734 ( .B(clk), .A(\g.we_clk [11656]));
Q_ASSIGN U4735 ( .B(clk), .A(\g.we_clk [11655]));
Q_ASSIGN U4736 ( .B(clk), .A(\g.we_clk [11654]));
Q_ASSIGN U4737 ( .B(clk), .A(\g.we_clk [11653]));
Q_ASSIGN U4738 ( .B(clk), .A(\g.we_clk [11652]));
Q_ASSIGN U4739 ( .B(clk), .A(\g.we_clk [11651]));
Q_ASSIGN U4740 ( .B(clk), .A(\g.we_clk [11650]));
Q_ASSIGN U4741 ( .B(clk), .A(\g.we_clk [11649]));
Q_ASSIGN U4742 ( .B(clk), .A(\g.we_clk [11648]));
Q_ASSIGN U4743 ( .B(clk), .A(\g.we_clk [11647]));
Q_ASSIGN U4744 ( .B(clk), .A(\g.we_clk [11646]));
Q_ASSIGN U4745 ( .B(clk), .A(\g.we_clk [11645]));
Q_ASSIGN U4746 ( .B(clk), .A(\g.we_clk [11644]));
Q_ASSIGN U4747 ( .B(clk), .A(\g.we_clk [11643]));
Q_ASSIGN U4748 ( .B(clk), .A(\g.we_clk [11642]));
Q_ASSIGN U4749 ( .B(clk), .A(\g.we_clk [11641]));
Q_ASSIGN U4750 ( .B(clk), .A(\g.we_clk [11640]));
Q_ASSIGN U4751 ( .B(clk), .A(\g.we_clk [11639]));
Q_ASSIGN U4752 ( .B(clk), .A(\g.we_clk [11638]));
Q_ASSIGN U4753 ( .B(clk), .A(\g.we_clk [11637]));
Q_ASSIGN U4754 ( .B(clk), .A(\g.we_clk [11636]));
Q_ASSIGN U4755 ( .B(clk), .A(\g.we_clk [11635]));
Q_ASSIGN U4756 ( .B(clk), .A(\g.we_clk [11634]));
Q_ASSIGN U4757 ( .B(clk), .A(\g.we_clk [11633]));
Q_ASSIGN U4758 ( .B(clk), .A(\g.we_clk [11632]));
Q_ASSIGN U4759 ( .B(clk), .A(\g.we_clk [11631]));
Q_ASSIGN U4760 ( .B(clk), .A(\g.we_clk [11630]));
Q_ASSIGN U4761 ( .B(clk), .A(\g.we_clk [11629]));
Q_ASSIGN U4762 ( .B(clk), .A(\g.we_clk [11628]));
Q_ASSIGN U4763 ( .B(clk), .A(\g.we_clk [11627]));
Q_ASSIGN U4764 ( .B(clk), .A(\g.we_clk [11626]));
Q_ASSIGN U4765 ( .B(clk), .A(\g.we_clk [11625]));
Q_ASSIGN U4766 ( .B(clk), .A(\g.we_clk [11624]));
Q_ASSIGN U4767 ( .B(clk), .A(\g.we_clk [11623]));
Q_ASSIGN U4768 ( .B(clk), .A(\g.we_clk [11622]));
Q_ASSIGN U4769 ( .B(clk), .A(\g.we_clk [11621]));
Q_ASSIGN U4770 ( .B(clk), .A(\g.we_clk [11620]));
Q_ASSIGN U4771 ( .B(clk), .A(\g.we_clk [11619]));
Q_ASSIGN U4772 ( .B(clk), .A(\g.we_clk [11618]));
Q_ASSIGN U4773 ( .B(clk), .A(\g.we_clk [11617]));
Q_ASSIGN U4774 ( .B(clk), .A(\g.we_clk [11616]));
Q_ASSIGN U4775 ( .B(clk), .A(\g.we_clk [11615]));
Q_ASSIGN U4776 ( .B(clk), .A(\g.we_clk [11614]));
Q_ASSIGN U4777 ( .B(clk), .A(\g.we_clk [11613]));
Q_ASSIGN U4778 ( .B(clk), .A(\g.we_clk [11612]));
Q_ASSIGN U4779 ( .B(clk), .A(\g.we_clk [11611]));
Q_ASSIGN U4780 ( .B(clk), .A(\g.we_clk [11610]));
Q_ASSIGN U4781 ( .B(clk), .A(\g.we_clk [11609]));
Q_ASSIGN U4782 ( .B(clk), .A(\g.we_clk [11608]));
Q_ASSIGN U4783 ( .B(clk), .A(\g.we_clk [11607]));
Q_ASSIGN U4784 ( .B(clk), .A(\g.we_clk [11606]));
Q_ASSIGN U4785 ( .B(clk), .A(\g.we_clk [11605]));
Q_ASSIGN U4786 ( .B(clk), .A(\g.we_clk [11604]));
Q_ASSIGN U4787 ( .B(clk), .A(\g.we_clk [11603]));
Q_ASSIGN U4788 ( .B(clk), .A(\g.we_clk [11602]));
Q_ASSIGN U4789 ( .B(clk), .A(\g.we_clk [11601]));
Q_ASSIGN U4790 ( .B(clk), .A(\g.we_clk [11600]));
Q_ASSIGN U4791 ( .B(clk), .A(\g.we_clk [11599]));
Q_ASSIGN U4792 ( .B(clk), .A(\g.we_clk [11598]));
Q_ASSIGN U4793 ( .B(clk), .A(\g.we_clk [11597]));
Q_ASSIGN U4794 ( .B(clk), .A(\g.we_clk [11596]));
Q_ASSIGN U4795 ( .B(clk), .A(\g.we_clk [11595]));
Q_ASSIGN U4796 ( .B(clk), .A(\g.we_clk [11594]));
Q_ASSIGN U4797 ( .B(clk), .A(\g.we_clk [11593]));
Q_ASSIGN U4798 ( .B(clk), .A(\g.we_clk [11592]));
Q_ASSIGN U4799 ( .B(clk), .A(\g.we_clk [11591]));
Q_ASSIGN U4800 ( .B(clk), .A(\g.we_clk [11590]));
Q_ASSIGN U4801 ( .B(clk), .A(\g.we_clk [11589]));
Q_ASSIGN U4802 ( .B(clk), .A(\g.we_clk [11588]));
Q_ASSIGN U4803 ( .B(clk), .A(\g.we_clk [11587]));
Q_ASSIGN U4804 ( .B(clk), .A(\g.we_clk [11586]));
Q_ASSIGN U4805 ( .B(clk), .A(\g.we_clk [11585]));
Q_ASSIGN U4806 ( .B(clk), .A(\g.we_clk [11584]));
Q_ASSIGN U4807 ( .B(clk), .A(\g.we_clk [11583]));
Q_ASSIGN U4808 ( .B(clk), .A(\g.we_clk [11582]));
Q_ASSIGN U4809 ( .B(clk), .A(\g.we_clk [11581]));
Q_ASSIGN U4810 ( .B(clk), .A(\g.we_clk [11580]));
Q_ASSIGN U4811 ( .B(clk), .A(\g.we_clk [11579]));
Q_ASSIGN U4812 ( .B(clk), .A(\g.we_clk [11578]));
Q_ASSIGN U4813 ( .B(clk), .A(\g.we_clk [11577]));
Q_ASSIGN U4814 ( .B(clk), .A(\g.we_clk [11576]));
Q_ASSIGN U4815 ( .B(clk), .A(\g.we_clk [11575]));
Q_ASSIGN U4816 ( .B(clk), .A(\g.we_clk [11574]));
Q_ASSIGN U4817 ( .B(clk), .A(\g.we_clk [11573]));
Q_ASSIGN U4818 ( .B(clk), .A(\g.we_clk [11572]));
Q_ASSIGN U4819 ( .B(clk), .A(\g.we_clk [11571]));
Q_ASSIGN U4820 ( .B(clk), .A(\g.we_clk [11570]));
Q_ASSIGN U4821 ( .B(clk), .A(\g.we_clk [11569]));
Q_ASSIGN U4822 ( .B(clk), .A(\g.we_clk [11568]));
Q_ASSIGN U4823 ( .B(clk), .A(\g.we_clk [11567]));
Q_ASSIGN U4824 ( .B(clk), .A(\g.we_clk [11566]));
Q_ASSIGN U4825 ( .B(clk), .A(\g.we_clk [11565]));
Q_ASSIGN U4826 ( .B(clk), .A(\g.we_clk [11564]));
Q_ASSIGN U4827 ( .B(clk), .A(\g.we_clk [11563]));
Q_ASSIGN U4828 ( .B(clk), .A(\g.we_clk [11562]));
Q_ASSIGN U4829 ( .B(clk), .A(\g.we_clk [11561]));
Q_ASSIGN U4830 ( .B(clk), .A(\g.we_clk [11560]));
Q_ASSIGN U4831 ( .B(clk), .A(\g.we_clk [11559]));
Q_ASSIGN U4832 ( .B(clk), .A(\g.we_clk [11558]));
Q_ASSIGN U4833 ( .B(clk), .A(\g.we_clk [11557]));
Q_ASSIGN U4834 ( .B(clk), .A(\g.we_clk [11556]));
Q_ASSIGN U4835 ( .B(clk), .A(\g.we_clk [11555]));
Q_ASSIGN U4836 ( .B(clk), .A(\g.we_clk [11554]));
Q_ASSIGN U4837 ( .B(clk), .A(\g.we_clk [11553]));
Q_ASSIGN U4838 ( .B(clk), .A(\g.we_clk [11552]));
Q_ASSIGN U4839 ( .B(clk), .A(\g.we_clk [11551]));
Q_ASSIGN U4840 ( .B(clk), .A(\g.we_clk [11550]));
Q_ASSIGN U4841 ( .B(clk), .A(\g.we_clk [11549]));
Q_ASSIGN U4842 ( .B(clk), .A(\g.we_clk [11548]));
Q_ASSIGN U4843 ( .B(clk), .A(\g.we_clk [11547]));
Q_ASSIGN U4844 ( .B(clk), .A(\g.we_clk [11546]));
Q_ASSIGN U4845 ( .B(clk), .A(\g.we_clk [11545]));
Q_ASSIGN U4846 ( .B(clk), .A(\g.we_clk [11544]));
Q_ASSIGN U4847 ( .B(clk), .A(\g.we_clk [11543]));
Q_ASSIGN U4848 ( .B(clk), .A(\g.we_clk [11542]));
Q_ASSIGN U4849 ( .B(clk), .A(\g.we_clk [11541]));
Q_ASSIGN U4850 ( .B(clk), .A(\g.we_clk [11540]));
Q_ASSIGN U4851 ( .B(clk), .A(\g.we_clk [11539]));
Q_ASSIGN U4852 ( .B(clk), .A(\g.we_clk [11538]));
Q_ASSIGN U4853 ( .B(clk), .A(\g.we_clk [11537]));
Q_ASSIGN U4854 ( .B(clk), .A(\g.we_clk [11536]));
Q_ASSIGN U4855 ( .B(clk), .A(\g.we_clk [11535]));
Q_ASSIGN U4856 ( .B(clk), .A(\g.we_clk [11534]));
Q_ASSIGN U4857 ( .B(clk), .A(\g.we_clk [11533]));
Q_ASSIGN U4858 ( .B(clk), .A(\g.we_clk [11532]));
Q_ASSIGN U4859 ( .B(clk), .A(\g.we_clk [11531]));
Q_ASSIGN U4860 ( .B(clk), .A(\g.we_clk [11530]));
Q_ASSIGN U4861 ( .B(clk), .A(\g.we_clk [11529]));
Q_ASSIGN U4862 ( .B(clk), .A(\g.we_clk [11528]));
Q_ASSIGN U4863 ( .B(clk), .A(\g.we_clk [11527]));
Q_ASSIGN U4864 ( .B(clk), .A(\g.we_clk [11526]));
Q_ASSIGN U4865 ( .B(clk), .A(\g.we_clk [11525]));
Q_ASSIGN U4866 ( .B(clk), .A(\g.we_clk [11524]));
Q_ASSIGN U4867 ( .B(clk), .A(\g.we_clk [11523]));
Q_ASSIGN U4868 ( .B(clk), .A(\g.we_clk [11522]));
Q_ASSIGN U4869 ( .B(clk), .A(\g.we_clk [11521]));
Q_ASSIGN U4870 ( .B(clk), .A(\g.we_clk [11520]));
Q_ASSIGN U4871 ( .B(clk), .A(\g.we_clk [11519]));
Q_ASSIGN U4872 ( .B(clk), .A(\g.we_clk [11518]));
Q_ASSIGN U4873 ( .B(clk), .A(\g.we_clk [11517]));
Q_ASSIGN U4874 ( .B(clk), .A(\g.we_clk [11516]));
Q_ASSIGN U4875 ( .B(clk), .A(\g.we_clk [11515]));
Q_ASSIGN U4876 ( .B(clk), .A(\g.we_clk [11514]));
Q_ASSIGN U4877 ( .B(clk), .A(\g.we_clk [11513]));
Q_ASSIGN U4878 ( .B(clk), .A(\g.we_clk [11512]));
Q_ASSIGN U4879 ( .B(clk), .A(\g.we_clk [11511]));
Q_ASSIGN U4880 ( .B(clk), .A(\g.we_clk [11510]));
Q_ASSIGN U4881 ( .B(clk), .A(\g.we_clk [11509]));
Q_ASSIGN U4882 ( .B(clk), .A(\g.we_clk [11508]));
Q_ASSIGN U4883 ( .B(clk), .A(\g.we_clk [11507]));
Q_ASSIGN U4884 ( .B(clk), .A(\g.we_clk [11506]));
Q_ASSIGN U4885 ( .B(clk), .A(\g.we_clk [11505]));
Q_ASSIGN U4886 ( .B(clk), .A(\g.we_clk [11504]));
Q_ASSIGN U4887 ( .B(clk), .A(\g.we_clk [11503]));
Q_ASSIGN U4888 ( .B(clk), .A(\g.we_clk [11502]));
Q_ASSIGN U4889 ( .B(clk), .A(\g.we_clk [11501]));
Q_ASSIGN U4890 ( .B(clk), .A(\g.we_clk [11500]));
Q_ASSIGN U4891 ( .B(clk), .A(\g.we_clk [11499]));
Q_ASSIGN U4892 ( .B(clk), .A(\g.we_clk [11498]));
Q_ASSIGN U4893 ( .B(clk), .A(\g.we_clk [11497]));
Q_ASSIGN U4894 ( .B(clk), .A(\g.we_clk [11496]));
Q_ASSIGN U4895 ( .B(clk), .A(\g.we_clk [11495]));
Q_ASSIGN U4896 ( .B(clk), .A(\g.we_clk [11494]));
Q_ASSIGN U4897 ( .B(clk), .A(\g.we_clk [11493]));
Q_ASSIGN U4898 ( .B(clk), .A(\g.we_clk [11492]));
Q_ASSIGN U4899 ( .B(clk), .A(\g.we_clk [11491]));
Q_ASSIGN U4900 ( .B(clk), .A(\g.we_clk [11490]));
Q_ASSIGN U4901 ( .B(clk), .A(\g.we_clk [11489]));
Q_ASSIGN U4902 ( .B(clk), .A(\g.we_clk [11488]));
Q_ASSIGN U4903 ( .B(clk), .A(\g.we_clk [11487]));
Q_ASSIGN U4904 ( .B(clk), .A(\g.we_clk [11486]));
Q_ASSIGN U4905 ( .B(clk), .A(\g.we_clk [11485]));
Q_ASSIGN U4906 ( .B(clk), .A(\g.we_clk [11484]));
Q_ASSIGN U4907 ( .B(clk), .A(\g.we_clk [11483]));
Q_ASSIGN U4908 ( .B(clk), .A(\g.we_clk [11482]));
Q_ASSIGN U4909 ( .B(clk), .A(\g.we_clk [11481]));
Q_ASSIGN U4910 ( .B(clk), .A(\g.we_clk [11480]));
Q_ASSIGN U4911 ( .B(clk), .A(\g.we_clk [11479]));
Q_ASSIGN U4912 ( .B(clk), .A(\g.we_clk [11478]));
Q_ASSIGN U4913 ( .B(clk), .A(\g.we_clk [11477]));
Q_ASSIGN U4914 ( .B(clk), .A(\g.we_clk [11476]));
Q_ASSIGN U4915 ( .B(clk), .A(\g.we_clk [11475]));
Q_ASSIGN U4916 ( .B(clk), .A(\g.we_clk [11474]));
Q_ASSIGN U4917 ( .B(clk), .A(\g.we_clk [11473]));
Q_ASSIGN U4918 ( .B(clk), .A(\g.we_clk [11472]));
Q_ASSIGN U4919 ( .B(clk), .A(\g.we_clk [11471]));
Q_ASSIGN U4920 ( .B(clk), .A(\g.we_clk [11470]));
Q_ASSIGN U4921 ( .B(clk), .A(\g.we_clk [11469]));
Q_ASSIGN U4922 ( .B(clk), .A(\g.we_clk [11468]));
Q_ASSIGN U4923 ( .B(clk), .A(\g.we_clk [11467]));
Q_ASSIGN U4924 ( .B(clk), .A(\g.we_clk [11466]));
Q_ASSIGN U4925 ( .B(clk), .A(\g.we_clk [11465]));
Q_ASSIGN U4926 ( .B(clk), .A(\g.we_clk [11464]));
Q_ASSIGN U4927 ( .B(clk), .A(\g.we_clk [11463]));
Q_ASSIGN U4928 ( .B(clk), .A(\g.we_clk [11462]));
Q_ASSIGN U4929 ( .B(clk), .A(\g.we_clk [11461]));
Q_ASSIGN U4930 ( .B(clk), .A(\g.we_clk [11460]));
Q_ASSIGN U4931 ( .B(clk), .A(\g.we_clk [11459]));
Q_ASSIGN U4932 ( .B(clk), .A(\g.we_clk [11458]));
Q_ASSIGN U4933 ( .B(clk), .A(\g.we_clk [11457]));
Q_ASSIGN U4934 ( .B(clk), .A(\g.we_clk [11456]));
Q_ASSIGN U4935 ( .B(clk), .A(\g.we_clk [11455]));
Q_ASSIGN U4936 ( .B(clk), .A(\g.we_clk [11454]));
Q_ASSIGN U4937 ( .B(clk), .A(\g.we_clk [11453]));
Q_ASSIGN U4938 ( .B(clk), .A(\g.we_clk [11452]));
Q_ASSIGN U4939 ( .B(clk), .A(\g.we_clk [11451]));
Q_ASSIGN U4940 ( .B(clk), .A(\g.we_clk [11450]));
Q_ASSIGN U4941 ( .B(clk), .A(\g.we_clk [11449]));
Q_ASSIGN U4942 ( .B(clk), .A(\g.we_clk [11448]));
Q_ASSIGN U4943 ( .B(clk), .A(\g.we_clk [11447]));
Q_ASSIGN U4944 ( .B(clk), .A(\g.we_clk [11446]));
Q_ASSIGN U4945 ( .B(clk), .A(\g.we_clk [11445]));
Q_ASSIGN U4946 ( .B(clk), .A(\g.we_clk [11444]));
Q_ASSIGN U4947 ( .B(clk), .A(\g.we_clk [11443]));
Q_ASSIGN U4948 ( .B(clk), .A(\g.we_clk [11442]));
Q_ASSIGN U4949 ( .B(clk), .A(\g.we_clk [11441]));
Q_ASSIGN U4950 ( .B(clk), .A(\g.we_clk [11440]));
Q_ASSIGN U4951 ( .B(clk), .A(\g.we_clk [11439]));
Q_ASSIGN U4952 ( .B(clk), .A(\g.we_clk [11438]));
Q_ASSIGN U4953 ( .B(clk), .A(\g.we_clk [11437]));
Q_ASSIGN U4954 ( .B(clk), .A(\g.we_clk [11436]));
Q_ASSIGN U4955 ( .B(clk), .A(\g.we_clk [11435]));
Q_ASSIGN U4956 ( .B(clk), .A(\g.we_clk [11434]));
Q_ASSIGN U4957 ( .B(clk), .A(\g.we_clk [11433]));
Q_ASSIGN U4958 ( .B(clk), .A(\g.we_clk [11432]));
Q_ASSIGN U4959 ( .B(clk), .A(\g.we_clk [11431]));
Q_ASSIGN U4960 ( .B(clk), .A(\g.we_clk [11430]));
Q_ASSIGN U4961 ( .B(clk), .A(\g.we_clk [11429]));
Q_ASSIGN U4962 ( .B(clk), .A(\g.we_clk [11428]));
Q_ASSIGN U4963 ( .B(clk), .A(\g.we_clk [11427]));
Q_ASSIGN U4964 ( .B(clk), .A(\g.we_clk [11426]));
Q_ASSIGN U4965 ( .B(clk), .A(\g.we_clk [11425]));
Q_ASSIGN U4966 ( .B(clk), .A(\g.we_clk [11424]));
Q_ASSIGN U4967 ( .B(clk), .A(\g.we_clk [11423]));
Q_ASSIGN U4968 ( .B(clk), .A(\g.we_clk [11422]));
Q_ASSIGN U4969 ( .B(clk), .A(\g.we_clk [11421]));
Q_ASSIGN U4970 ( .B(clk), .A(\g.we_clk [11420]));
Q_ASSIGN U4971 ( .B(clk), .A(\g.we_clk [11419]));
Q_ASSIGN U4972 ( .B(clk), .A(\g.we_clk [11418]));
Q_ASSIGN U4973 ( .B(clk), .A(\g.we_clk [11417]));
Q_ASSIGN U4974 ( .B(clk), .A(\g.we_clk [11416]));
Q_ASSIGN U4975 ( .B(clk), .A(\g.we_clk [11415]));
Q_ASSIGN U4976 ( .B(clk), .A(\g.we_clk [11414]));
Q_ASSIGN U4977 ( .B(clk), .A(\g.we_clk [11413]));
Q_ASSIGN U4978 ( .B(clk), .A(\g.we_clk [11412]));
Q_ASSIGN U4979 ( .B(clk), .A(\g.we_clk [11411]));
Q_ASSIGN U4980 ( .B(clk), .A(\g.we_clk [11410]));
Q_ASSIGN U4981 ( .B(clk), .A(\g.we_clk [11409]));
Q_ASSIGN U4982 ( .B(clk), .A(\g.we_clk [11408]));
Q_ASSIGN U4983 ( .B(clk), .A(\g.we_clk [11407]));
Q_ASSIGN U4984 ( .B(clk), .A(\g.we_clk [11406]));
Q_ASSIGN U4985 ( .B(clk), .A(\g.we_clk [11405]));
Q_ASSIGN U4986 ( .B(clk), .A(\g.we_clk [11404]));
Q_ASSIGN U4987 ( .B(clk), .A(\g.we_clk [11403]));
Q_ASSIGN U4988 ( .B(clk), .A(\g.we_clk [11402]));
Q_ASSIGN U4989 ( .B(clk), .A(\g.we_clk [11401]));
Q_ASSIGN U4990 ( .B(clk), .A(\g.we_clk [11400]));
Q_ASSIGN U4991 ( .B(clk), .A(\g.we_clk [11399]));
Q_ASSIGN U4992 ( .B(clk), .A(\g.we_clk [11398]));
Q_ASSIGN U4993 ( .B(clk), .A(\g.we_clk [11397]));
Q_ASSIGN U4994 ( .B(clk), .A(\g.we_clk [11396]));
Q_ASSIGN U4995 ( .B(clk), .A(\g.we_clk [11395]));
Q_ASSIGN U4996 ( .B(clk), .A(\g.we_clk [11394]));
Q_ASSIGN U4997 ( .B(clk), .A(\g.we_clk [11393]));
Q_ASSIGN U4998 ( .B(clk), .A(\g.we_clk [11392]));
Q_ASSIGN U4999 ( .B(clk), .A(\g.we_clk [11391]));
Q_ASSIGN U5000 ( .B(clk), .A(\g.we_clk [11390]));
Q_ASSIGN U5001 ( .B(clk), .A(\g.we_clk [11389]));
Q_ASSIGN U5002 ( .B(clk), .A(\g.we_clk [11388]));
Q_ASSIGN U5003 ( .B(clk), .A(\g.we_clk [11387]));
Q_ASSIGN U5004 ( .B(clk), .A(\g.we_clk [11386]));
Q_ASSIGN U5005 ( .B(clk), .A(\g.we_clk [11385]));
Q_ASSIGN U5006 ( .B(clk), .A(\g.we_clk [11384]));
Q_ASSIGN U5007 ( .B(clk), .A(\g.we_clk [11383]));
Q_ASSIGN U5008 ( .B(clk), .A(\g.we_clk [11382]));
Q_ASSIGN U5009 ( .B(clk), .A(\g.we_clk [11381]));
Q_ASSIGN U5010 ( .B(clk), .A(\g.we_clk [11380]));
Q_ASSIGN U5011 ( .B(clk), .A(\g.we_clk [11379]));
Q_ASSIGN U5012 ( .B(clk), .A(\g.we_clk [11378]));
Q_ASSIGN U5013 ( .B(clk), .A(\g.we_clk [11377]));
Q_ASSIGN U5014 ( .B(clk), .A(\g.we_clk [11376]));
Q_ASSIGN U5015 ( .B(clk), .A(\g.we_clk [11375]));
Q_ASSIGN U5016 ( .B(clk), .A(\g.we_clk [11374]));
Q_ASSIGN U5017 ( .B(clk), .A(\g.we_clk [11373]));
Q_ASSIGN U5018 ( .B(clk), .A(\g.we_clk [11372]));
Q_ASSIGN U5019 ( .B(clk), .A(\g.we_clk [11371]));
Q_ASSIGN U5020 ( .B(clk), .A(\g.we_clk [11370]));
Q_ASSIGN U5021 ( .B(clk), .A(\g.we_clk [11369]));
Q_ASSIGN U5022 ( .B(clk), .A(\g.we_clk [11368]));
Q_ASSIGN U5023 ( .B(clk), .A(\g.we_clk [11367]));
Q_ASSIGN U5024 ( .B(clk), .A(\g.we_clk [11366]));
Q_ASSIGN U5025 ( .B(clk), .A(\g.we_clk [11365]));
Q_ASSIGN U5026 ( .B(clk), .A(\g.we_clk [11364]));
Q_ASSIGN U5027 ( .B(clk), .A(\g.we_clk [11363]));
Q_ASSIGN U5028 ( .B(clk), .A(\g.we_clk [11362]));
Q_ASSIGN U5029 ( .B(clk), .A(\g.we_clk [11361]));
Q_ASSIGN U5030 ( .B(clk), .A(\g.we_clk [11360]));
Q_ASSIGN U5031 ( .B(clk), .A(\g.we_clk [11359]));
Q_ASSIGN U5032 ( .B(clk), .A(\g.we_clk [11358]));
Q_ASSIGN U5033 ( .B(clk), .A(\g.we_clk [11357]));
Q_ASSIGN U5034 ( .B(clk), .A(\g.we_clk [11356]));
Q_ASSIGN U5035 ( .B(clk), .A(\g.we_clk [11355]));
Q_ASSIGN U5036 ( .B(clk), .A(\g.we_clk [11354]));
Q_ASSIGN U5037 ( .B(clk), .A(\g.we_clk [11353]));
Q_ASSIGN U5038 ( .B(clk), .A(\g.we_clk [11352]));
Q_ASSIGN U5039 ( .B(clk), .A(\g.we_clk [11351]));
Q_ASSIGN U5040 ( .B(clk), .A(\g.we_clk [11350]));
Q_ASSIGN U5041 ( .B(clk), .A(\g.we_clk [11349]));
Q_ASSIGN U5042 ( .B(clk), .A(\g.we_clk [11348]));
Q_ASSIGN U5043 ( .B(clk), .A(\g.we_clk [11347]));
Q_ASSIGN U5044 ( .B(clk), .A(\g.we_clk [11346]));
Q_ASSIGN U5045 ( .B(clk), .A(\g.we_clk [11345]));
Q_ASSIGN U5046 ( .B(clk), .A(\g.we_clk [11344]));
Q_ASSIGN U5047 ( .B(clk), .A(\g.we_clk [11343]));
Q_ASSIGN U5048 ( .B(clk), .A(\g.we_clk [11342]));
Q_ASSIGN U5049 ( .B(clk), .A(\g.we_clk [11341]));
Q_ASSIGN U5050 ( .B(clk), .A(\g.we_clk [11340]));
Q_ASSIGN U5051 ( .B(clk), .A(\g.we_clk [11339]));
Q_ASSIGN U5052 ( .B(clk), .A(\g.we_clk [11338]));
Q_ASSIGN U5053 ( .B(clk), .A(\g.we_clk [11337]));
Q_ASSIGN U5054 ( .B(clk), .A(\g.we_clk [11336]));
Q_ASSIGN U5055 ( .B(clk), .A(\g.we_clk [11335]));
Q_ASSIGN U5056 ( .B(clk), .A(\g.we_clk [11334]));
Q_ASSIGN U5057 ( .B(clk), .A(\g.we_clk [11333]));
Q_ASSIGN U5058 ( .B(clk), .A(\g.we_clk [11332]));
Q_ASSIGN U5059 ( .B(clk), .A(\g.we_clk [11331]));
Q_ASSIGN U5060 ( .B(clk), .A(\g.we_clk [11330]));
Q_ASSIGN U5061 ( .B(clk), .A(\g.we_clk [11329]));
Q_ASSIGN U5062 ( .B(clk), .A(\g.we_clk [11328]));
Q_ASSIGN U5063 ( .B(clk), .A(\g.we_clk [11327]));
Q_ASSIGN U5064 ( .B(clk), .A(\g.we_clk [11326]));
Q_ASSIGN U5065 ( .B(clk), .A(\g.we_clk [11325]));
Q_ASSIGN U5066 ( .B(clk), .A(\g.we_clk [11324]));
Q_ASSIGN U5067 ( .B(clk), .A(\g.we_clk [11323]));
Q_ASSIGN U5068 ( .B(clk), .A(\g.we_clk [11322]));
Q_ASSIGN U5069 ( .B(clk), .A(\g.we_clk [11321]));
Q_ASSIGN U5070 ( .B(clk), .A(\g.we_clk [11320]));
Q_ASSIGN U5071 ( .B(clk), .A(\g.we_clk [11319]));
Q_ASSIGN U5072 ( .B(clk), .A(\g.we_clk [11318]));
Q_ASSIGN U5073 ( .B(clk), .A(\g.we_clk [11317]));
Q_ASSIGN U5074 ( .B(clk), .A(\g.we_clk [11316]));
Q_ASSIGN U5075 ( .B(clk), .A(\g.we_clk [11315]));
Q_ASSIGN U5076 ( .B(clk), .A(\g.we_clk [11314]));
Q_ASSIGN U5077 ( .B(clk), .A(\g.we_clk [11313]));
Q_ASSIGN U5078 ( .B(clk), .A(\g.we_clk [11312]));
Q_ASSIGN U5079 ( .B(clk), .A(\g.we_clk [11311]));
Q_ASSIGN U5080 ( .B(clk), .A(\g.we_clk [11310]));
Q_ASSIGN U5081 ( .B(clk), .A(\g.we_clk [11309]));
Q_ASSIGN U5082 ( .B(clk), .A(\g.we_clk [11308]));
Q_ASSIGN U5083 ( .B(clk), .A(\g.we_clk [11307]));
Q_ASSIGN U5084 ( .B(clk), .A(\g.we_clk [11306]));
Q_ASSIGN U5085 ( .B(clk), .A(\g.we_clk [11305]));
Q_ASSIGN U5086 ( .B(clk), .A(\g.we_clk [11304]));
Q_ASSIGN U5087 ( .B(clk), .A(\g.we_clk [11303]));
Q_ASSIGN U5088 ( .B(clk), .A(\g.we_clk [11302]));
Q_ASSIGN U5089 ( .B(clk), .A(\g.we_clk [11301]));
Q_ASSIGN U5090 ( .B(clk), .A(\g.we_clk [11300]));
Q_ASSIGN U5091 ( .B(clk), .A(\g.we_clk [11299]));
Q_ASSIGN U5092 ( .B(clk), .A(\g.we_clk [11298]));
Q_ASSIGN U5093 ( .B(clk), .A(\g.we_clk [11297]));
Q_ASSIGN U5094 ( .B(clk), .A(\g.we_clk [11296]));
Q_ASSIGN U5095 ( .B(clk), .A(\g.we_clk [11295]));
Q_ASSIGN U5096 ( .B(clk), .A(\g.we_clk [11294]));
Q_ASSIGN U5097 ( .B(clk), .A(\g.we_clk [11293]));
Q_ASSIGN U5098 ( .B(clk), .A(\g.we_clk [11292]));
Q_ASSIGN U5099 ( .B(clk), .A(\g.we_clk [11291]));
Q_ASSIGN U5100 ( .B(clk), .A(\g.we_clk [11290]));
Q_ASSIGN U5101 ( .B(clk), .A(\g.we_clk [11289]));
Q_ASSIGN U5102 ( .B(clk), .A(\g.we_clk [11288]));
Q_ASSIGN U5103 ( .B(clk), .A(\g.we_clk [11287]));
Q_ASSIGN U5104 ( .B(clk), .A(\g.we_clk [11286]));
Q_ASSIGN U5105 ( .B(clk), .A(\g.we_clk [11285]));
Q_ASSIGN U5106 ( .B(clk), .A(\g.we_clk [11284]));
Q_ASSIGN U5107 ( .B(clk), .A(\g.we_clk [11283]));
Q_ASSIGN U5108 ( .B(clk), .A(\g.we_clk [11282]));
Q_ASSIGN U5109 ( .B(clk), .A(\g.we_clk [11281]));
Q_ASSIGN U5110 ( .B(clk), .A(\g.we_clk [11280]));
Q_ASSIGN U5111 ( .B(clk), .A(\g.we_clk [11279]));
Q_ASSIGN U5112 ( .B(clk), .A(\g.we_clk [11278]));
Q_ASSIGN U5113 ( .B(clk), .A(\g.we_clk [11277]));
Q_ASSIGN U5114 ( .B(clk), .A(\g.we_clk [11276]));
Q_ASSIGN U5115 ( .B(clk), .A(\g.we_clk [11275]));
Q_ASSIGN U5116 ( .B(clk), .A(\g.we_clk [11274]));
Q_ASSIGN U5117 ( .B(clk), .A(\g.we_clk [11273]));
Q_ASSIGN U5118 ( .B(clk), .A(\g.we_clk [11272]));
Q_ASSIGN U5119 ( .B(clk), .A(\g.we_clk [11271]));
Q_ASSIGN U5120 ( .B(clk), .A(\g.we_clk [11270]));
Q_ASSIGN U5121 ( .B(clk), .A(\g.we_clk [11269]));
Q_ASSIGN U5122 ( .B(clk), .A(\g.we_clk [11268]));
Q_ASSIGN U5123 ( .B(clk), .A(\g.we_clk [11267]));
Q_ASSIGN U5124 ( .B(clk), .A(\g.we_clk [11266]));
Q_ASSIGN U5125 ( .B(clk), .A(\g.we_clk [11265]));
Q_ASSIGN U5126 ( .B(clk), .A(\g.we_clk [11264]));
Q_ASSIGN U5127 ( .B(clk), .A(\g.we_clk [11263]));
Q_ASSIGN U5128 ( .B(clk), .A(\g.we_clk [11262]));
Q_ASSIGN U5129 ( .B(clk), .A(\g.we_clk [11261]));
Q_ASSIGN U5130 ( .B(clk), .A(\g.we_clk [11260]));
Q_ASSIGN U5131 ( .B(clk), .A(\g.we_clk [11259]));
Q_ASSIGN U5132 ( .B(clk), .A(\g.we_clk [11258]));
Q_ASSIGN U5133 ( .B(clk), .A(\g.we_clk [11257]));
Q_ASSIGN U5134 ( .B(clk), .A(\g.we_clk [11256]));
Q_ASSIGN U5135 ( .B(clk), .A(\g.we_clk [11255]));
Q_ASSIGN U5136 ( .B(clk), .A(\g.we_clk [11254]));
Q_ASSIGN U5137 ( .B(clk), .A(\g.we_clk [11253]));
Q_ASSIGN U5138 ( .B(clk), .A(\g.we_clk [11252]));
Q_ASSIGN U5139 ( .B(clk), .A(\g.we_clk [11251]));
Q_ASSIGN U5140 ( .B(clk), .A(\g.we_clk [11250]));
Q_ASSIGN U5141 ( .B(clk), .A(\g.we_clk [11249]));
Q_ASSIGN U5142 ( .B(clk), .A(\g.we_clk [11248]));
Q_ASSIGN U5143 ( .B(clk), .A(\g.we_clk [11247]));
Q_ASSIGN U5144 ( .B(clk), .A(\g.we_clk [11246]));
Q_ASSIGN U5145 ( .B(clk), .A(\g.we_clk [11245]));
Q_ASSIGN U5146 ( .B(clk), .A(\g.we_clk [11244]));
Q_ASSIGN U5147 ( .B(clk), .A(\g.we_clk [11243]));
Q_ASSIGN U5148 ( .B(clk), .A(\g.we_clk [11242]));
Q_ASSIGN U5149 ( .B(clk), .A(\g.we_clk [11241]));
Q_ASSIGN U5150 ( .B(clk), .A(\g.we_clk [11240]));
Q_ASSIGN U5151 ( .B(clk), .A(\g.we_clk [11239]));
Q_ASSIGN U5152 ( .B(clk), .A(\g.we_clk [11238]));
Q_ASSIGN U5153 ( .B(clk), .A(\g.we_clk [11237]));
Q_ASSIGN U5154 ( .B(clk), .A(\g.we_clk [11236]));
Q_ASSIGN U5155 ( .B(clk), .A(\g.we_clk [11235]));
Q_ASSIGN U5156 ( .B(clk), .A(\g.we_clk [11234]));
Q_ASSIGN U5157 ( .B(clk), .A(\g.we_clk [11233]));
Q_ASSIGN U5158 ( .B(clk), .A(\g.we_clk [11232]));
Q_ASSIGN U5159 ( .B(clk), .A(\g.we_clk [11231]));
Q_ASSIGN U5160 ( .B(clk), .A(\g.we_clk [11230]));
Q_ASSIGN U5161 ( .B(clk), .A(\g.we_clk [11229]));
Q_ASSIGN U5162 ( .B(clk), .A(\g.we_clk [11228]));
Q_ASSIGN U5163 ( .B(clk), .A(\g.we_clk [11227]));
Q_ASSIGN U5164 ( .B(clk), .A(\g.we_clk [11226]));
Q_ASSIGN U5165 ( .B(clk), .A(\g.we_clk [11225]));
Q_ASSIGN U5166 ( .B(clk), .A(\g.we_clk [11224]));
Q_ASSIGN U5167 ( .B(clk), .A(\g.we_clk [11223]));
Q_ASSIGN U5168 ( .B(clk), .A(\g.we_clk [11222]));
Q_ASSIGN U5169 ( .B(clk), .A(\g.we_clk [11221]));
Q_ASSIGN U5170 ( .B(clk), .A(\g.we_clk [11220]));
Q_ASSIGN U5171 ( .B(clk), .A(\g.we_clk [11219]));
Q_ASSIGN U5172 ( .B(clk), .A(\g.we_clk [11218]));
Q_ASSIGN U5173 ( .B(clk), .A(\g.we_clk [11217]));
Q_ASSIGN U5174 ( .B(clk), .A(\g.we_clk [11216]));
Q_ASSIGN U5175 ( .B(clk), .A(\g.we_clk [11215]));
Q_ASSIGN U5176 ( .B(clk), .A(\g.we_clk [11214]));
Q_ASSIGN U5177 ( .B(clk), .A(\g.we_clk [11213]));
Q_ASSIGN U5178 ( .B(clk), .A(\g.we_clk [11212]));
Q_ASSIGN U5179 ( .B(clk), .A(\g.we_clk [11211]));
Q_ASSIGN U5180 ( .B(clk), .A(\g.we_clk [11210]));
Q_ASSIGN U5181 ( .B(clk), .A(\g.we_clk [11209]));
Q_ASSIGN U5182 ( .B(clk), .A(\g.we_clk [11208]));
Q_ASSIGN U5183 ( .B(clk), .A(\g.we_clk [11207]));
Q_ASSIGN U5184 ( .B(clk), .A(\g.we_clk [11206]));
Q_ASSIGN U5185 ( .B(clk), .A(\g.we_clk [11205]));
Q_ASSIGN U5186 ( .B(clk), .A(\g.we_clk [11204]));
Q_ASSIGN U5187 ( .B(clk), .A(\g.we_clk [11203]));
Q_ASSIGN U5188 ( .B(clk), .A(\g.we_clk [11202]));
Q_ASSIGN U5189 ( .B(clk), .A(\g.we_clk [11201]));
Q_ASSIGN U5190 ( .B(clk), .A(\g.we_clk [11200]));
Q_ASSIGN U5191 ( .B(clk), .A(\g.we_clk [11199]));
Q_ASSIGN U5192 ( .B(clk), .A(\g.we_clk [11198]));
Q_ASSIGN U5193 ( .B(clk), .A(\g.we_clk [11197]));
Q_ASSIGN U5194 ( .B(clk), .A(\g.we_clk [11196]));
Q_ASSIGN U5195 ( .B(clk), .A(\g.we_clk [11195]));
Q_ASSIGN U5196 ( .B(clk), .A(\g.we_clk [11194]));
Q_ASSIGN U5197 ( .B(clk), .A(\g.we_clk [11193]));
Q_ASSIGN U5198 ( .B(clk), .A(\g.we_clk [11192]));
Q_ASSIGN U5199 ( .B(clk), .A(\g.we_clk [11191]));
Q_ASSIGN U5200 ( .B(clk), .A(\g.we_clk [11190]));
Q_ASSIGN U5201 ( .B(clk), .A(\g.we_clk [11189]));
Q_ASSIGN U5202 ( .B(clk), .A(\g.we_clk [11188]));
Q_ASSIGN U5203 ( .B(clk), .A(\g.we_clk [11187]));
Q_ASSIGN U5204 ( .B(clk), .A(\g.we_clk [11186]));
Q_ASSIGN U5205 ( .B(clk), .A(\g.we_clk [11185]));
Q_ASSIGN U5206 ( .B(clk), .A(\g.we_clk [11184]));
Q_ASSIGN U5207 ( .B(clk), .A(\g.we_clk [11183]));
Q_ASSIGN U5208 ( .B(clk), .A(\g.we_clk [11182]));
Q_ASSIGN U5209 ( .B(clk), .A(\g.we_clk [11181]));
Q_ASSIGN U5210 ( .B(clk), .A(\g.we_clk [11180]));
Q_ASSIGN U5211 ( .B(clk), .A(\g.we_clk [11179]));
Q_ASSIGN U5212 ( .B(clk), .A(\g.we_clk [11178]));
Q_ASSIGN U5213 ( .B(clk), .A(\g.we_clk [11177]));
Q_ASSIGN U5214 ( .B(clk), .A(\g.we_clk [11176]));
Q_ASSIGN U5215 ( .B(clk), .A(\g.we_clk [11175]));
Q_ASSIGN U5216 ( .B(clk), .A(\g.we_clk [11174]));
Q_ASSIGN U5217 ( .B(clk), .A(\g.we_clk [11173]));
Q_ASSIGN U5218 ( .B(clk), .A(\g.we_clk [11172]));
Q_ASSIGN U5219 ( .B(clk), .A(\g.we_clk [11171]));
Q_ASSIGN U5220 ( .B(clk), .A(\g.we_clk [11170]));
Q_ASSIGN U5221 ( .B(clk), .A(\g.we_clk [11169]));
Q_ASSIGN U5222 ( .B(clk), .A(\g.we_clk [11168]));
Q_ASSIGN U5223 ( .B(clk), .A(\g.we_clk [11167]));
Q_ASSIGN U5224 ( .B(clk), .A(\g.we_clk [11166]));
Q_ASSIGN U5225 ( .B(clk), .A(\g.we_clk [11165]));
Q_ASSIGN U5226 ( .B(clk), .A(\g.we_clk [11164]));
Q_ASSIGN U5227 ( .B(clk), .A(\g.we_clk [11163]));
Q_ASSIGN U5228 ( .B(clk), .A(\g.we_clk [11162]));
Q_ASSIGN U5229 ( .B(clk), .A(\g.we_clk [11161]));
Q_ASSIGN U5230 ( .B(clk), .A(\g.we_clk [11160]));
Q_ASSIGN U5231 ( .B(clk), .A(\g.we_clk [11159]));
Q_ASSIGN U5232 ( .B(clk), .A(\g.we_clk [11158]));
Q_ASSIGN U5233 ( .B(clk), .A(\g.we_clk [11157]));
Q_ASSIGN U5234 ( .B(clk), .A(\g.we_clk [11156]));
Q_ASSIGN U5235 ( .B(clk), .A(\g.we_clk [11155]));
Q_ASSIGN U5236 ( .B(clk), .A(\g.we_clk [11154]));
Q_ASSIGN U5237 ( .B(clk), .A(\g.we_clk [11153]));
Q_ASSIGN U5238 ( .B(clk), .A(\g.we_clk [11152]));
Q_ASSIGN U5239 ( .B(clk), .A(\g.we_clk [11151]));
Q_ASSIGN U5240 ( .B(clk), .A(\g.we_clk [11150]));
Q_ASSIGN U5241 ( .B(clk), .A(\g.we_clk [11149]));
Q_ASSIGN U5242 ( .B(clk), .A(\g.we_clk [11148]));
Q_ASSIGN U5243 ( .B(clk), .A(\g.we_clk [11147]));
Q_ASSIGN U5244 ( .B(clk), .A(\g.we_clk [11146]));
Q_ASSIGN U5245 ( .B(clk), .A(\g.we_clk [11145]));
Q_ASSIGN U5246 ( .B(clk), .A(\g.we_clk [11144]));
Q_ASSIGN U5247 ( .B(clk), .A(\g.we_clk [11143]));
Q_ASSIGN U5248 ( .B(clk), .A(\g.we_clk [11142]));
Q_ASSIGN U5249 ( .B(clk), .A(\g.we_clk [11141]));
Q_ASSIGN U5250 ( .B(clk), .A(\g.we_clk [11140]));
Q_ASSIGN U5251 ( .B(clk), .A(\g.we_clk [11139]));
Q_ASSIGN U5252 ( .B(clk), .A(\g.we_clk [11138]));
Q_ASSIGN U5253 ( .B(clk), .A(\g.we_clk [11137]));
Q_ASSIGN U5254 ( .B(clk), .A(\g.we_clk [11136]));
Q_ASSIGN U5255 ( .B(clk), .A(\g.we_clk [11135]));
Q_ASSIGN U5256 ( .B(clk), .A(\g.we_clk [11134]));
Q_ASSIGN U5257 ( .B(clk), .A(\g.we_clk [11133]));
Q_ASSIGN U5258 ( .B(clk), .A(\g.we_clk [11132]));
Q_ASSIGN U5259 ( .B(clk), .A(\g.we_clk [11131]));
Q_ASSIGN U5260 ( .B(clk), .A(\g.we_clk [11130]));
Q_ASSIGN U5261 ( .B(clk), .A(\g.we_clk [11129]));
Q_ASSIGN U5262 ( .B(clk), .A(\g.we_clk [11128]));
Q_ASSIGN U5263 ( .B(clk), .A(\g.we_clk [11127]));
Q_ASSIGN U5264 ( .B(clk), .A(\g.we_clk [11126]));
Q_ASSIGN U5265 ( .B(clk), .A(\g.we_clk [11125]));
Q_ASSIGN U5266 ( .B(clk), .A(\g.we_clk [11124]));
Q_ASSIGN U5267 ( .B(clk), .A(\g.we_clk [11123]));
Q_ASSIGN U5268 ( .B(clk), .A(\g.we_clk [11122]));
Q_ASSIGN U5269 ( .B(clk), .A(\g.we_clk [11121]));
Q_ASSIGN U5270 ( .B(clk), .A(\g.we_clk [11120]));
Q_ASSIGN U5271 ( .B(clk), .A(\g.we_clk [11119]));
Q_ASSIGN U5272 ( .B(clk), .A(\g.we_clk [11118]));
Q_ASSIGN U5273 ( .B(clk), .A(\g.we_clk [11117]));
Q_ASSIGN U5274 ( .B(clk), .A(\g.we_clk [11116]));
Q_ASSIGN U5275 ( .B(clk), .A(\g.we_clk [11115]));
Q_ASSIGN U5276 ( .B(clk), .A(\g.we_clk [11114]));
Q_ASSIGN U5277 ( .B(clk), .A(\g.we_clk [11113]));
Q_ASSIGN U5278 ( .B(clk), .A(\g.we_clk [11112]));
Q_ASSIGN U5279 ( .B(clk), .A(\g.we_clk [11111]));
Q_ASSIGN U5280 ( .B(clk), .A(\g.we_clk [11110]));
Q_ASSIGN U5281 ( .B(clk), .A(\g.we_clk [11109]));
Q_ASSIGN U5282 ( .B(clk), .A(\g.we_clk [11108]));
Q_ASSIGN U5283 ( .B(clk), .A(\g.we_clk [11107]));
Q_ASSIGN U5284 ( .B(clk), .A(\g.we_clk [11106]));
Q_ASSIGN U5285 ( .B(clk), .A(\g.we_clk [11105]));
Q_ASSIGN U5286 ( .B(clk), .A(\g.we_clk [11104]));
Q_ASSIGN U5287 ( .B(clk), .A(\g.we_clk [11103]));
Q_ASSIGN U5288 ( .B(clk), .A(\g.we_clk [11102]));
Q_ASSIGN U5289 ( .B(clk), .A(\g.we_clk [11101]));
Q_ASSIGN U5290 ( .B(clk), .A(\g.we_clk [11100]));
Q_ASSIGN U5291 ( .B(clk), .A(\g.we_clk [11099]));
Q_ASSIGN U5292 ( .B(clk), .A(\g.we_clk [11098]));
Q_ASSIGN U5293 ( .B(clk), .A(\g.we_clk [11097]));
Q_ASSIGN U5294 ( .B(clk), .A(\g.we_clk [11096]));
Q_ASSIGN U5295 ( .B(clk), .A(\g.we_clk [11095]));
Q_ASSIGN U5296 ( .B(clk), .A(\g.we_clk [11094]));
Q_ASSIGN U5297 ( .B(clk), .A(\g.we_clk [11093]));
Q_ASSIGN U5298 ( .B(clk), .A(\g.we_clk [11092]));
Q_ASSIGN U5299 ( .B(clk), .A(\g.we_clk [11091]));
Q_ASSIGN U5300 ( .B(clk), .A(\g.we_clk [11090]));
Q_ASSIGN U5301 ( .B(clk), .A(\g.we_clk [11089]));
Q_ASSIGN U5302 ( .B(clk), .A(\g.we_clk [11088]));
Q_ASSIGN U5303 ( .B(clk), .A(\g.we_clk [11087]));
Q_ASSIGN U5304 ( .B(clk), .A(\g.we_clk [11086]));
Q_ASSIGN U5305 ( .B(clk), .A(\g.we_clk [11085]));
Q_ASSIGN U5306 ( .B(clk), .A(\g.we_clk [11084]));
Q_ASSIGN U5307 ( .B(clk), .A(\g.we_clk [11083]));
Q_ASSIGN U5308 ( .B(clk), .A(\g.we_clk [11082]));
Q_ASSIGN U5309 ( .B(clk), .A(\g.we_clk [11081]));
Q_ASSIGN U5310 ( .B(clk), .A(\g.we_clk [11080]));
Q_ASSIGN U5311 ( .B(clk), .A(\g.we_clk [11079]));
Q_ASSIGN U5312 ( .B(clk), .A(\g.we_clk [11078]));
Q_ASSIGN U5313 ( .B(clk), .A(\g.we_clk [11077]));
Q_ASSIGN U5314 ( .B(clk), .A(\g.we_clk [11076]));
Q_ASSIGN U5315 ( .B(clk), .A(\g.we_clk [11075]));
Q_ASSIGN U5316 ( .B(clk), .A(\g.we_clk [11074]));
Q_ASSIGN U5317 ( .B(clk), .A(\g.we_clk [11073]));
Q_ASSIGN U5318 ( .B(clk), .A(\g.we_clk [11072]));
Q_ASSIGN U5319 ( .B(clk), .A(\g.we_clk [11071]));
Q_ASSIGN U5320 ( .B(clk), .A(\g.we_clk [11070]));
Q_ASSIGN U5321 ( .B(clk), .A(\g.we_clk [11069]));
Q_ASSIGN U5322 ( .B(clk), .A(\g.we_clk [11068]));
Q_ASSIGN U5323 ( .B(clk), .A(\g.we_clk [11067]));
Q_ASSIGN U5324 ( .B(clk), .A(\g.we_clk [11066]));
Q_ASSIGN U5325 ( .B(clk), .A(\g.we_clk [11065]));
Q_ASSIGN U5326 ( .B(clk), .A(\g.we_clk [11064]));
Q_ASSIGN U5327 ( .B(clk), .A(\g.we_clk [11063]));
Q_ASSIGN U5328 ( .B(clk), .A(\g.we_clk [11062]));
Q_ASSIGN U5329 ( .B(clk), .A(\g.we_clk [11061]));
Q_ASSIGN U5330 ( .B(clk), .A(\g.we_clk [11060]));
Q_ASSIGN U5331 ( .B(clk), .A(\g.we_clk [11059]));
Q_ASSIGN U5332 ( .B(clk), .A(\g.we_clk [11058]));
Q_ASSIGN U5333 ( .B(clk), .A(\g.we_clk [11057]));
Q_ASSIGN U5334 ( .B(clk), .A(\g.we_clk [11056]));
Q_ASSIGN U5335 ( .B(clk), .A(\g.we_clk [11055]));
Q_ASSIGN U5336 ( .B(clk), .A(\g.we_clk [11054]));
Q_ASSIGN U5337 ( .B(clk), .A(\g.we_clk [11053]));
Q_ASSIGN U5338 ( .B(clk), .A(\g.we_clk [11052]));
Q_ASSIGN U5339 ( .B(clk), .A(\g.we_clk [11051]));
Q_ASSIGN U5340 ( .B(clk), .A(\g.we_clk [11050]));
Q_ASSIGN U5341 ( .B(clk), .A(\g.we_clk [11049]));
Q_ASSIGN U5342 ( .B(clk), .A(\g.we_clk [11048]));
Q_ASSIGN U5343 ( .B(clk), .A(\g.we_clk [11047]));
Q_ASSIGN U5344 ( .B(clk), .A(\g.we_clk [11046]));
Q_ASSIGN U5345 ( .B(clk), .A(\g.we_clk [11045]));
Q_ASSIGN U5346 ( .B(clk), .A(\g.we_clk [11044]));
Q_ASSIGN U5347 ( .B(clk), .A(\g.we_clk [11043]));
Q_ASSIGN U5348 ( .B(clk), .A(\g.we_clk [11042]));
Q_ASSIGN U5349 ( .B(clk), .A(\g.we_clk [11041]));
Q_ASSIGN U5350 ( .B(clk), .A(\g.we_clk [11040]));
Q_ASSIGN U5351 ( .B(clk), .A(\g.we_clk [11039]));
Q_ASSIGN U5352 ( .B(clk), .A(\g.we_clk [11038]));
Q_ASSIGN U5353 ( .B(clk), .A(\g.we_clk [11037]));
Q_ASSIGN U5354 ( .B(clk), .A(\g.we_clk [11036]));
Q_ASSIGN U5355 ( .B(clk), .A(\g.we_clk [11035]));
Q_ASSIGN U5356 ( .B(clk), .A(\g.we_clk [11034]));
Q_ASSIGN U5357 ( .B(clk), .A(\g.we_clk [11033]));
Q_ASSIGN U5358 ( .B(clk), .A(\g.we_clk [11032]));
Q_ASSIGN U5359 ( .B(clk), .A(\g.we_clk [11031]));
Q_ASSIGN U5360 ( .B(clk), .A(\g.we_clk [11030]));
Q_ASSIGN U5361 ( .B(clk), .A(\g.we_clk [11029]));
Q_ASSIGN U5362 ( .B(clk), .A(\g.we_clk [11028]));
Q_ASSIGN U5363 ( .B(clk), .A(\g.we_clk [11027]));
Q_ASSIGN U5364 ( .B(clk), .A(\g.we_clk [11026]));
Q_ASSIGN U5365 ( .B(clk), .A(\g.we_clk [11025]));
Q_ASSIGN U5366 ( .B(clk), .A(\g.we_clk [11024]));
Q_ASSIGN U5367 ( .B(clk), .A(\g.we_clk [11023]));
Q_ASSIGN U5368 ( .B(clk), .A(\g.we_clk [11022]));
Q_ASSIGN U5369 ( .B(clk), .A(\g.we_clk [11021]));
Q_ASSIGN U5370 ( .B(clk), .A(\g.we_clk [11020]));
Q_ASSIGN U5371 ( .B(clk), .A(\g.we_clk [11019]));
Q_ASSIGN U5372 ( .B(clk), .A(\g.we_clk [11018]));
Q_ASSIGN U5373 ( .B(clk), .A(\g.we_clk [11017]));
Q_ASSIGN U5374 ( .B(clk), .A(\g.we_clk [11016]));
Q_ASSIGN U5375 ( .B(clk), .A(\g.we_clk [11015]));
Q_ASSIGN U5376 ( .B(clk), .A(\g.we_clk [11014]));
Q_ASSIGN U5377 ( .B(clk), .A(\g.we_clk [11013]));
Q_ASSIGN U5378 ( .B(clk), .A(\g.we_clk [11012]));
Q_ASSIGN U5379 ( .B(clk), .A(\g.we_clk [11011]));
Q_ASSIGN U5380 ( .B(clk), .A(\g.we_clk [11010]));
Q_ASSIGN U5381 ( .B(clk), .A(\g.we_clk [11009]));
Q_ASSIGN U5382 ( .B(clk), .A(\g.we_clk [11008]));
Q_ASSIGN U5383 ( .B(clk), .A(\g.we_clk [11007]));
Q_ASSIGN U5384 ( .B(clk), .A(\g.we_clk [11006]));
Q_ASSIGN U5385 ( .B(clk), .A(\g.we_clk [11005]));
Q_ASSIGN U5386 ( .B(clk), .A(\g.we_clk [11004]));
Q_ASSIGN U5387 ( .B(clk), .A(\g.we_clk [11003]));
Q_ASSIGN U5388 ( .B(clk), .A(\g.we_clk [11002]));
Q_ASSIGN U5389 ( .B(clk), .A(\g.we_clk [11001]));
Q_ASSIGN U5390 ( .B(clk), .A(\g.we_clk [11000]));
Q_ASSIGN U5391 ( .B(clk), .A(\g.we_clk [10999]));
Q_ASSIGN U5392 ( .B(clk), .A(\g.we_clk [10998]));
Q_ASSIGN U5393 ( .B(clk), .A(\g.we_clk [10997]));
Q_ASSIGN U5394 ( .B(clk), .A(\g.we_clk [10996]));
Q_ASSIGN U5395 ( .B(clk), .A(\g.we_clk [10995]));
Q_ASSIGN U5396 ( .B(clk), .A(\g.we_clk [10994]));
Q_ASSIGN U5397 ( .B(clk), .A(\g.we_clk [10993]));
Q_ASSIGN U5398 ( .B(clk), .A(\g.we_clk [10992]));
Q_ASSIGN U5399 ( .B(clk), .A(\g.we_clk [10991]));
Q_ASSIGN U5400 ( .B(clk), .A(\g.we_clk [10990]));
Q_ASSIGN U5401 ( .B(clk), .A(\g.we_clk [10989]));
Q_ASSIGN U5402 ( .B(clk), .A(\g.we_clk [10988]));
Q_ASSIGN U5403 ( .B(clk), .A(\g.we_clk [10987]));
Q_ASSIGN U5404 ( .B(clk), .A(\g.we_clk [10986]));
Q_ASSIGN U5405 ( .B(clk), .A(\g.we_clk [10985]));
Q_ASSIGN U5406 ( .B(clk), .A(\g.we_clk [10984]));
Q_ASSIGN U5407 ( .B(clk), .A(\g.we_clk [10983]));
Q_ASSIGN U5408 ( .B(clk), .A(\g.we_clk [10982]));
Q_ASSIGN U5409 ( .B(clk), .A(\g.we_clk [10981]));
Q_ASSIGN U5410 ( .B(clk), .A(\g.we_clk [10980]));
Q_ASSIGN U5411 ( .B(clk), .A(\g.we_clk [10979]));
Q_ASSIGN U5412 ( .B(clk), .A(\g.we_clk [10978]));
Q_ASSIGN U5413 ( .B(clk), .A(\g.we_clk [10977]));
Q_ASSIGN U5414 ( .B(clk), .A(\g.we_clk [10976]));
Q_ASSIGN U5415 ( .B(clk), .A(\g.we_clk [10975]));
Q_ASSIGN U5416 ( .B(clk), .A(\g.we_clk [10974]));
Q_ASSIGN U5417 ( .B(clk), .A(\g.we_clk [10973]));
Q_ASSIGN U5418 ( .B(clk), .A(\g.we_clk [10972]));
Q_ASSIGN U5419 ( .B(clk), .A(\g.we_clk [10971]));
Q_ASSIGN U5420 ( .B(clk), .A(\g.we_clk [10970]));
Q_ASSIGN U5421 ( .B(clk), .A(\g.we_clk [10969]));
Q_ASSIGN U5422 ( .B(clk), .A(\g.we_clk [10968]));
Q_ASSIGN U5423 ( .B(clk), .A(\g.we_clk [10967]));
Q_ASSIGN U5424 ( .B(clk), .A(\g.we_clk [10966]));
Q_ASSIGN U5425 ( .B(clk), .A(\g.we_clk [10965]));
Q_ASSIGN U5426 ( .B(clk), .A(\g.we_clk [10964]));
Q_ASSIGN U5427 ( .B(clk), .A(\g.we_clk [10963]));
Q_ASSIGN U5428 ( .B(clk), .A(\g.we_clk [10962]));
Q_ASSIGN U5429 ( .B(clk), .A(\g.we_clk [10961]));
Q_ASSIGN U5430 ( .B(clk), .A(\g.we_clk [10960]));
Q_ASSIGN U5431 ( .B(clk), .A(\g.we_clk [10959]));
Q_ASSIGN U5432 ( .B(clk), .A(\g.we_clk [10958]));
Q_ASSIGN U5433 ( .B(clk), .A(\g.we_clk [10957]));
Q_ASSIGN U5434 ( .B(clk), .A(\g.we_clk [10956]));
Q_ASSIGN U5435 ( .B(clk), .A(\g.we_clk [10955]));
Q_ASSIGN U5436 ( .B(clk), .A(\g.we_clk [10954]));
Q_ASSIGN U5437 ( .B(clk), .A(\g.we_clk [10953]));
Q_ASSIGN U5438 ( .B(clk), .A(\g.we_clk [10952]));
Q_ASSIGN U5439 ( .B(clk), .A(\g.we_clk [10951]));
Q_ASSIGN U5440 ( .B(clk), .A(\g.we_clk [10950]));
Q_ASSIGN U5441 ( .B(clk), .A(\g.we_clk [10949]));
Q_ASSIGN U5442 ( .B(clk), .A(\g.we_clk [10948]));
Q_ASSIGN U5443 ( .B(clk), .A(\g.we_clk [10947]));
Q_ASSIGN U5444 ( .B(clk), .A(\g.we_clk [10946]));
Q_ASSIGN U5445 ( .B(clk), .A(\g.we_clk [10945]));
Q_ASSIGN U5446 ( .B(clk), .A(\g.we_clk [10944]));
Q_ASSIGN U5447 ( .B(clk), .A(\g.we_clk [10943]));
Q_ASSIGN U5448 ( .B(clk), .A(\g.we_clk [10942]));
Q_ASSIGN U5449 ( .B(clk), .A(\g.we_clk [10941]));
Q_ASSIGN U5450 ( .B(clk), .A(\g.we_clk [10940]));
Q_ASSIGN U5451 ( .B(clk), .A(\g.we_clk [10939]));
Q_ASSIGN U5452 ( .B(clk), .A(\g.we_clk [10938]));
Q_ASSIGN U5453 ( .B(clk), .A(\g.we_clk [10937]));
Q_ASSIGN U5454 ( .B(clk), .A(\g.we_clk [10936]));
Q_ASSIGN U5455 ( .B(clk), .A(\g.we_clk [10935]));
Q_ASSIGN U5456 ( .B(clk), .A(\g.we_clk [10934]));
Q_ASSIGN U5457 ( .B(clk), .A(\g.we_clk [10933]));
Q_ASSIGN U5458 ( .B(clk), .A(\g.we_clk [10932]));
Q_ASSIGN U5459 ( .B(clk), .A(\g.we_clk [10931]));
Q_ASSIGN U5460 ( .B(clk), .A(\g.we_clk [10930]));
Q_ASSIGN U5461 ( .B(clk), .A(\g.we_clk [10929]));
Q_ASSIGN U5462 ( .B(clk), .A(\g.we_clk [10928]));
Q_ASSIGN U5463 ( .B(clk), .A(\g.we_clk [10927]));
Q_ASSIGN U5464 ( .B(clk), .A(\g.we_clk [10926]));
Q_ASSIGN U5465 ( .B(clk), .A(\g.we_clk [10925]));
Q_ASSIGN U5466 ( .B(clk), .A(\g.we_clk [10924]));
Q_ASSIGN U5467 ( .B(clk), .A(\g.we_clk [10923]));
Q_ASSIGN U5468 ( .B(clk), .A(\g.we_clk [10922]));
Q_ASSIGN U5469 ( .B(clk), .A(\g.we_clk [10921]));
Q_ASSIGN U5470 ( .B(clk), .A(\g.we_clk [10920]));
Q_ASSIGN U5471 ( .B(clk), .A(\g.we_clk [10919]));
Q_ASSIGN U5472 ( .B(clk), .A(\g.we_clk [10918]));
Q_ASSIGN U5473 ( .B(clk), .A(\g.we_clk [10917]));
Q_ASSIGN U5474 ( .B(clk), .A(\g.we_clk [10916]));
Q_ASSIGN U5475 ( .B(clk), .A(\g.we_clk [10915]));
Q_ASSIGN U5476 ( .B(clk), .A(\g.we_clk [10914]));
Q_ASSIGN U5477 ( .B(clk), .A(\g.we_clk [10913]));
Q_ASSIGN U5478 ( .B(clk), .A(\g.we_clk [10912]));
Q_ASSIGN U5479 ( .B(clk), .A(\g.we_clk [10911]));
Q_ASSIGN U5480 ( .B(clk), .A(\g.we_clk [10910]));
Q_ASSIGN U5481 ( .B(clk), .A(\g.we_clk [10909]));
Q_ASSIGN U5482 ( .B(clk), .A(\g.we_clk [10908]));
Q_ASSIGN U5483 ( .B(clk), .A(\g.we_clk [10907]));
Q_ASSIGN U5484 ( .B(clk), .A(\g.we_clk [10906]));
Q_ASSIGN U5485 ( .B(clk), .A(\g.we_clk [10905]));
Q_ASSIGN U5486 ( .B(clk), .A(\g.we_clk [10904]));
Q_ASSIGN U5487 ( .B(clk), .A(\g.we_clk [10903]));
Q_ASSIGN U5488 ( .B(clk), .A(\g.we_clk [10902]));
Q_ASSIGN U5489 ( .B(clk), .A(\g.we_clk [10901]));
Q_ASSIGN U5490 ( .B(clk), .A(\g.we_clk [10900]));
Q_ASSIGN U5491 ( .B(clk), .A(\g.we_clk [10899]));
Q_ASSIGN U5492 ( .B(clk), .A(\g.we_clk [10898]));
Q_ASSIGN U5493 ( .B(clk), .A(\g.we_clk [10897]));
Q_ASSIGN U5494 ( .B(clk), .A(\g.we_clk [10896]));
Q_ASSIGN U5495 ( .B(clk), .A(\g.we_clk [10895]));
Q_ASSIGN U5496 ( .B(clk), .A(\g.we_clk [10894]));
Q_ASSIGN U5497 ( .B(clk), .A(\g.we_clk [10893]));
Q_ASSIGN U5498 ( .B(clk), .A(\g.we_clk [10892]));
Q_ASSIGN U5499 ( .B(clk), .A(\g.we_clk [10891]));
Q_ASSIGN U5500 ( .B(clk), .A(\g.we_clk [10890]));
Q_ASSIGN U5501 ( .B(clk), .A(\g.we_clk [10889]));
Q_ASSIGN U5502 ( .B(clk), .A(\g.we_clk [10888]));
Q_ASSIGN U5503 ( .B(clk), .A(\g.we_clk [10887]));
Q_ASSIGN U5504 ( .B(clk), .A(\g.we_clk [10886]));
Q_ASSIGN U5505 ( .B(clk), .A(\g.we_clk [10885]));
Q_ASSIGN U5506 ( .B(clk), .A(\g.we_clk [10884]));
Q_ASSIGN U5507 ( .B(clk), .A(\g.we_clk [10883]));
Q_ASSIGN U5508 ( .B(clk), .A(\g.we_clk [10882]));
Q_ASSIGN U5509 ( .B(clk), .A(\g.we_clk [10881]));
Q_ASSIGN U5510 ( .B(clk), .A(\g.we_clk [10880]));
Q_ASSIGN U5511 ( .B(clk), .A(\g.we_clk [10879]));
Q_ASSIGN U5512 ( .B(clk), .A(\g.we_clk [10878]));
Q_ASSIGN U5513 ( .B(clk), .A(\g.we_clk [10877]));
Q_ASSIGN U5514 ( .B(clk), .A(\g.we_clk [10876]));
Q_ASSIGN U5515 ( .B(clk), .A(\g.we_clk [10875]));
Q_ASSIGN U5516 ( .B(clk), .A(\g.we_clk [10874]));
Q_ASSIGN U5517 ( .B(clk), .A(\g.we_clk [10873]));
Q_ASSIGN U5518 ( .B(clk), .A(\g.we_clk [10872]));
Q_ASSIGN U5519 ( .B(clk), .A(\g.we_clk [10871]));
Q_ASSIGN U5520 ( .B(clk), .A(\g.we_clk [10870]));
Q_ASSIGN U5521 ( .B(clk), .A(\g.we_clk [10869]));
Q_ASSIGN U5522 ( .B(clk), .A(\g.we_clk [10868]));
Q_ASSIGN U5523 ( .B(clk), .A(\g.we_clk [10867]));
Q_ASSIGN U5524 ( .B(clk), .A(\g.we_clk [10866]));
Q_ASSIGN U5525 ( .B(clk), .A(\g.we_clk [10865]));
Q_ASSIGN U5526 ( .B(clk), .A(\g.we_clk [10864]));
Q_ASSIGN U5527 ( .B(clk), .A(\g.we_clk [10863]));
Q_ASSIGN U5528 ( .B(clk), .A(\g.we_clk [10862]));
Q_ASSIGN U5529 ( .B(clk), .A(\g.we_clk [10861]));
Q_ASSIGN U5530 ( .B(clk), .A(\g.we_clk [10860]));
Q_ASSIGN U5531 ( .B(clk), .A(\g.we_clk [10859]));
Q_ASSIGN U5532 ( .B(clk), .A(\g.we_clk [10858]));
Q_ASSIGN U5533 ( .B(clk), .A(\g.we_clk [10857]));
Q_ASSIGN U5534 ( .B(clk), .A(\g.we_clk [10856]));
Q_ASSIGN U5535 ( .B(clk), .A(\g.we_clk [10855]));
Q_ASSIGN U5536 ( .B(clk), .A(\g.we_clk [10854]));
Q_ASSIGN U5537 ( .B(clk), .A(\g.we_clk [10853]));
Q_ASSIGN U5538 ( .B(clk), .A(\g.we_clk [10852]));
Q_ASSIGN U5539 ( .B(clk), .A(\g.we_clk [10851]));
Q_ASSIGN U5540 ( .B(clk), .A(\g.we_clk [10850]));
Q_ASSIGN U5541 ( .B(clk), .A(\g.we_clk [10849]));
Q_ASSIGN U5542 ( .B(clk), .A(\g.we_clk [10848]));
Q_ASSIGN U5543 ( .B(clk), .A(\g.we_clk [10847]));
Q_ASSIGN U5544 ( .B(clk), .A(\g.we_clk [10846]));
Q_ASSIGN U5545 ( .B(clk), .A(\g.we_clk [10845]));
Q_ASSIGN U5546 ( .B(clk), .A(\g.we_clk [10844]));
Q_ASSIGN U5547 ( .B(clk), .A(\g.we_clk [10843]));
Q_ASSIGN U5548 ( .B(clk), .A(\g.we_clk [10842]));
Q_ASSIGN U5549 ( .B(clk), .A(\g.we_clk [10841]));
Q_ASSIGN U5550 ( .B(clk), .A(\g.we_clk [10840]));
Q_ASSIGN U5551 ( .B(clk), .A(\g.we_clk [10839]));
Q_ASSIGN U5552 ( .B(clk), .A(\g.we_clk [10838]));
Q_ASSIGN U5553 ( .B(clk), .A(\g.we_clk [10837]));
Q_ASSIGN U5554 ( .B(clk), .A(\g.we_clk [10836]));
Q_ASSIGN U5555 ( .B(clk), .A(\g.we_clk [10835]));
Q_ASSIGN U5556 ( .B(clk), .A(\g.we_clk [10834]));
Q_ASSIGN U5557 ( .B(clk), .A(\g.we_clk [10833]));
Q_ASSIGN U5558 ( .B(clk), .A(\g.we_clk [10832]));
Q_ASSIGN U5559 ( .B(clk), .A(\g.we_clk [10831]));
Q_ASSIGN U5560 ( .B(clk), .A(\g.we_clk [10830]));
Q_ASSIGN U5561 ( .B(clk), .A(\g.we_clk [10829]));
Q_ASSIGN U5562 ( .B(clk), .A(\g.we_clk [10828]));
Q_ASSIGN U5563 ( .B(clk), .A(\g.we_clk [10827]));
Q_ASSIGN U5564 ( .B(clk), .A(\g.we_clk [10826]));
Q_ASSIGN U5565 ( .B(clk), .A(\g.we_clk [10825]));
Q_ASSIGN U5566 ( .B(clk), .A(\g.we_clk [10824]));
Q_ASSIGN U5567 ( .B(clk), .A(\g.we_clk [10823]));
Q_ASSIGN U5568 ( .B(clk), .A(\g.we_clk [10822]));
Q_ASSIGN U5569 ( .B(clk), .A(\g.we_clk [10821]));
Q_ASSIGN U5570 ( .B(clk), .A(\g.we_clk [10820]));
Q_ASSIGN U5571 ( .B(clk), .A(\g.we_clk [10819]));
Q_ASSIGN U5572 ( .B(clk), .A(\g.we_clk [10818]));
Q_ASSIGN U5573 ( .B(clk), .A(\g.we_clk [10817]));
Q_ASSIGN U5574 ( .B(clk), .A(\g.we_clk [10816]));
Q_ASSIGN U5575 ( .B(clk), .A(\g.we_clk [10815]));
Q_ASSIGN U5576 ( .B(clk), .A(\g.we_clk [10814]));
Q_ASSIGN U5577 ( .B(clk), .A(\g.we_clk [10813]));
Q_ASSIGN U5578 ( .B(clk), .A(\g.we_clk [10812]));
Q_ASSIGN U5579 ( .B(clk), .A(\g.we_clk [10811]));
Q_ASSIGN U5580 ( .B(clk), .A(\g.we_clk [10810]));
Q_ASSIGN U5581 ( .B(clk), .A(\g.we_clk [10809]));
Q_ASSIGN U5582 ( .B(clk), .A(\g.we_clk [10808]));
Q_ASSIGN U5583 ( .B(clk), .A(\g.we_clk [10807]));
Q_ASSIGN U5584 ( .B(clk), .A(\g.we_clk [10806]));
Q_ASSIGN U5585 ( .B(clk), .A(\g.we_clk [10805]));
Q_ASSIGN U5586 ( .B(clk), .A(\g.we_clk [10804]));
Q_ASSIGN U5587 ( .B(clk), .A(\g.we_clk [10803]));
Q_ASSIGN U5588 ( .B(clk), .A(\g.we_clk [10802]));
Q_ASSIGN U5589 ( .B(clk), .A(\g.we_clk [10801]));
Q_ASSIGN U5590 ( .B(clk), .A(\g.we_clk [10800]));
Q_ASSIGN U5591 ( .B(clk), .A(\g.we_clk [10799]));
Q_ASSIGN U5592 ( .B(clk), .A(\g.we_clk [10798]));
Q_ASSIGN U5593 ( .B(clk), .A(\g.we_clk [10797]));
Q_ASSIGN U5594 ( .B(clk), .A(\g.we_clk [10796]));
Q_ASSIGN U5595 ( .B(clk), .A(\g.we_clk [10795]));
Q_ASSIGN U5596 ( .B(clk), .A(\g.we_clk [10794]));
Q_ASSIGN U5597 ( .B(clk), .A(\g.we_clk [10793]));
Q_ASSIGN U5598 ( .B(clk), .A(\g.we_clk [10792]));
Q_ASSIGN U5599 ( .B(clk), .A(\g.we_clk [10791]));
Q_ASSIGN U5600 ( .B(clk), .A(\g.we_clk [10790]));
Q_ASSIGN U5601 ( .B(clk), .A(\g.we_clk [10789]));
Q_ASSIGN U5602 ( .B(clk), .A(\g.we_clk [10788]));
Q_ASSIGN U5603 ( .B(clk), .A(\g.we_clk [10787]));
Q_ASSIGN U5604 ( .B(clk), .A(\g.we_clk [10786]));
Q_ASSIGN U5605 ( .B(clk), .A(\g.we_clk [10785]));
Q_ASSIGN U5606 ( .B(clk), .A(\g.we_clk [10784]));
Q_ASSIGN U5607 ( .B(clk), .A(\g.we_clk [10783]));
Q_ASSIGN U5608 ( .B(clk), .A(\g.we_clk [10782]));
Q_ASSIGN U5609 ( .B(clk), .A(\g.we_clk [10781]));
Q_ASSIGN U5610 ( .B(clk), .A(\g.we_clk [10780]));
Q_ASSIGN U5611 ( .B(clk), .A(\g.we_clk [10779]));
Q_ASSIGN U5612 ( .B(clk), .A(\g.we_clk [10778]));
Q_ASSIGN U5613 ( .B(clk), .A(\g.we_clk [10777]));
Q_ASSIGN U5614 ( .B(clk), .A(\g.we_clk [10776]));
Q_ASSIGN U5615 ( .B(clk), .A(\g.we_clk [10775]));
Q_ASSIGN U5616 ( .B(clk), .A(\g.we_clk [10774]));
Q_ASSIGN U5617 ( .B(clk), .A(\g.we_clk [10773]));
Q_ASSIGN U5618 ( .B(clk), .A(\g.we_clk [10772]));
Q_ASSIGN U5619 ( .B(clk), .A(\g.we_clk [10771]));
Q_ASSIGN U5620 ( .B(clk), .A(\g.we_clk [10770]));
Q_ASSIGN U5621 ( .B(clk), .A(\g.we_clk [10769]));
Q_ASSIGN U5622 ( .B(clk), .A(\g.we_clk [10768]));
Q_ASSIGN U5623 ( .B(clk), .A(\g.we_clk [10767]));
Q_ASSIGN U5624 ( .B(clk), .A(\g.we_clk [10766]));
Q_ASSIGN U5625 ( .B(clk), .A(\g.we_clk [10765]));
Q_ASSIGN U5626 ( .B(clk), .A(\g.we_clk [10764]));
Q_ASSIGN U5627 ( .B(clk), .A(\g.we_clk [10763]));
Q_ASSIGN U5628 ( .B(clk), .A(\g.we_clk [10762]));
Q_ASSIGN U5629 ( .B(clk), .A(\g.we_clk [10761]));
Q_ASSIGN U5630 ( .B(clk), .A(\g.we_clk [10760]));
Q_ASSIGN U5631 ( .B(clk), .A(\g.we_clk [10759]));
Q_ASSIGN U5632 ( .B(clk), .A(\g.we_clk [10758]));
Q_ASSIGN U5633 ( .B(clk), .A(\g.we_clk [10757]));
Q_ASSIGN U5634 ( .B(clk), .A(\g.we_clk [10756]));
Q_ASSIGN U5635 ( .B(clk), .A(\g.we_clk [10755]));
Q_ASSIGN U5636 ( .B(clk), .A(\g.we_clk [10754]));
Q_ASSIGN U5637 ( .B(clk), .A(\g.we_clk [10753]));
Q_ASSIGN U5638 ( .B(clk), .A(\g.we_clk [10752]));
Q_ASSIGN U5639 ( .B(clk), .A(\g.we_clk [10751]));
Q_ASSIGN U5640 ( .B(clk), .A(\g.we_clk [10750]));
Q_ASSIGN U5641 ( .B(clk), .A(\g.we_clk [10749]));
Q_ASSIGN U5642 ( .B(clk), .A(\g.we_clk [10748]));
Q_ASSIGN U5643 ( .B(clk), .A(\g.we_clk [10747]));
Q_ASSIGN U5644 ( .B(clk), .A(\g.we_clk [10746]));
Q_ASSIGN U5645 ( .B(clk), .A(\g.we_clk [10745]));
Q_ASSIGN U5646 ( .B(clk), .A(\g.we_clk [10744]));
Q_ASSIGN U5647 ( .B(clk), .A(\g.we_clk [10743]));
Q_ASSIGN U5648 ( .B(clk), .A(\g.we_clk [10742]));
Q_ASSIGN U5649 ( .B(clk), .A(\g.we_clk [10741]));
Q_ASSIGN U5650 ( .B(clk), .A(\g.we_clk [10740]));
Q_ASSIGN U5651 ( .B(clk), .A(\g.we_clk [10739]));
Q_ASSIGN U5652 ( .B(clk), .A(\g.we_clk [10738]));
Q_ASSIGN U5653 ( .B(clk), .A(\g.we_clk [10737]));
Q_ASSIGN U5654 ( .B(clk), .A(\g.we_clk [10736]));
Q_ASSIGN U5655 ( .B(clk), .A(\g.we_clk [10735]));
Q_ASSIGN U5656 ( .B(clk), .A(\g.we_clk [10734]));
Q_ASSIGN U5657 ( .B(clk), .A(\g.we_clk [10733]));
Q_ASSIGN U5658 ( .B(clk), .A(\g.we_clk [10732]));
Q_ASSIGN U5659 ( .B(clk), .A(\g.we_clk [10731]));
Q_ASSIGN U5660 ( .B(clk), .A(\g.we_clk [10730]));
Q_ASSIGN U5661 ( .B(clk), .A(\g.we_clk [10729]));
Q_ASSIGN U5662 ( .B(clk), .A(\g.we_clk [10728]));
Q_ASSIGN U5663 ( .B(clk), .A(\g.we_clk [10727]));
Q_ASSIGN U5664 ( .B(clk), .A(\g.we_clk [10726]));
Q_ASSIGN U5665 ( .B(clk), .A(\g.we_clk [10725]));
Q_ASSIGN U5666 ( .B(clk), .A(\g.we_clk [10724]));
Q_ASSIGN U5667 ( .B(clk), .A(\g.we_clk [10723]));
Q_ASSIGN U5668 ( .B(clk), .A(\g.we_clk [10722]));
Q_ASSIGN U5669 ( .B(clk), .A(\g.we_clk [10721]));
Q_ASSIGN U5670 ( .B(clk), .A(\g.we_clk [10720]));
Q_ASSIGN U5671 ( .B(clk), .A(\g.we_clk [10719]));
Q_ASSIGN U5672 ( .B(clk), .A(\g.we_clk [10718]));
Q_ASSIGN U5673 ( .B(clk), .A(\g.we_clk [10717]));
Q_ASSIGN U5674 ( .B(clk), .A(\g.we_clk [10716]));
Q_ASSIGN U5675 ( .B(clk), .A(\g.we_clk [10715]));
Q_ASSIGN U5676 ( .B(clk), .A(\g.we_clk [10714]));
Q_ASSIGN U5677 ( .B(clk), .A(\g.we_clk [10713]));
Q_ASSIGN U5678 ( .B(clk), .A(\g.we_clk [10712]));
Q_ASSIGN U5679 ( .B(clk), .A(\g.we_clk [10711]));
Q_ASSIGN U5680 ( .B(clk), .A(\g.we_clk [10710]));
Q_ASSIGN U5681 ( .B(clk), .A(\g.we_clk [10709]));
Q_ASSIGN U5682 ( .B(clk), .A(\g.we_clk [10708]));
Q_ASSIGN U5683 ( .B(clk), .A(\g.we_clk [10707]));
Q_ASSIGN U5684 ( .B(clk), .A(\g.we_clk [10706]));
Q_ASSIGN U5685 ( .B(clk), .A(\g.we_clk [10705]));
Q_ASSIGN U5686 ( .B(clk), .A(\g.we_clk [10704]));
Q_ASSIGN U5687 ( .B(clk), .A(\g.we_clk [10703]));
Q_ASSIGN U5688 ( .B(clk), .A(\g.we_clk [10702]));
Q_ASSIGN U5689 ( .B(clk), .A(\g.we_clk [10701]));
Q_ASSIGN U5690 ( .B(clk), .A(\g.we_clk [10700]));
Q_ASSIGN U5691 ( .B(clk), .A(\g.we_clk [10699]));
Q_ASSIGN U5692 ( .B(clk), .A(\g.we_clk [10698]));
Q_ASSIGN U5693 ( .B(clk), .A(\g.we_clk [10697]));
Q_ASSIGN U5694 ( .B(clk), .A(\g.we_clk [10696]));
Q_ASSIGN U5695 ( .B(clk), .A(\g.we_clk [10695]));
Q_ASSIGN U5696 ( .B(clk), .A(\g.we_clk [10694]));
Q_ASSIGN U5697 ( .B(clk), .A(\g.we_clk [10693]));
Q_ASSIGN U5698 ( .B(clk), .A(\g.we_clk [10692]));
Q_ASSIGN U5699 ( .B(clk), .A(\g.we_clk [10691]));
Q_ASSIGN U5700 ( .B(clk), .A(\g.we_clk [10690]));
Q_ASSIGN U5701 ( .B(clk), .A(\g.we_clk [10689]));
Q_ASSIGN U5702 ( .B(clk), .A(\g.we_clk [10688]));
Q_ASSIGN U5703 ( .B(clk), .A(\g.we_clk [10687]));
Q_ASSIGN U5704 ( .B(clk), .A(\g.we_clk [10686]));
Q_ASSIGN U5705 ( .B(clk), .A(\g.we_clk [10685]));
Q_ASSIGN U5706 ( .B(clk), .A(\g.we_clk [10684]));
Q_ASSIGN U5707 ( .B(clk), .A(\g.we_clk [10683]));
Q_ASSIGN U5708 ( .B(clk), .A(\g.we_clk [10682]));
Q_ASSIGN U5709 ( .B(clk), .A(\g.we_clk [10681]));
Q_ASSIGN U5710 ( .B(clk), .A(\g.we_clk [10680]));
Q_ASSIGN U5711 ( .B(clk), .A(\g.we_clk [10679]));
Q_ASSIGN U5712 ( .B(clk), .A(\g.we_clk [10678]));
Q_ASSIGN U5713 ( .B(clk), .A(\g.we_clk [10677]));
Q_ASSIGN U5714 ( .B(clk), .A(\g.we_clk [10676]));
Q_ASSIGN U5715 ( .B(clk), .A(\g.we_clk [10675]));
Q_ASSIGN U5716 ( .B(clk), .A(\g.we_clk [10674]));
Q_ASSIGN U5717 ( .B(clk), .A(\g.we_clk [10673]));
Q_ASSIGN U5718 ( .B(clk), .A(\g.we_clk [10672]));
Q_ASSIGN U5719 ( .B(clk), .A(\g.we_clk [10671]));
Q_ASSIGN U5720 ( .B(clk), .A(\g.we_clk [10670]));
Q_ASSIGN U5721 ( .B(clk), .A(\g.we_clk [10669]));
Q_ASSIGN U5722 ( .B(clk), .A(\g.we_clk [10668]));
Q_ASSIGN U5723 ( .B(clk), .A(\g.we_clk [10667]));
Q_ASSIGN U5724 ( .B(clk), .A(\g.we_clk [10666]));
Q_ASSIGN U5725 ( .B(clk), .A(\g.we_clk [10665]));
Q_ASSIGN U5726 ( .B(clk), .A(\g.we_clk [10664]));
Q_ASSIGN U5727 ( .B(clk), .A(\g.we_clk [10663]));
Q_ASSIGN U5728 ( .B(clk), .A(\g.we_clk [10662]));
Q_ASSIGN U5729 ( .B(clk), .A(\g.we_clk [10661]));
Q_ASSIGN U5730 ( .B(clk), .A(\g.we_clk [10660]));
Q_ASSIGN U5731 ( .B(clk), .A(\g.we_clk [10659]));
Q_ASSIGN U5732 ( .B(clk), .A(\g.we_clk [10658]));
Q_ASSIGN U5733 ( .B(clk), .A(\g.we_clk [10657]));
Q_ASSIGN U5734 ( .B(clk), .A(\g.we_clk [10656]));
Q_ASSIGN U5735 ( .B(clk), .A(\g.we_clk [10655]));
Q_ASSIGN U5736 ( .B(clk), .A(\g.we_clk [10654]));
Q_ASSIGN U5737 ( .B(clk), .A(\g.we_clk [10653]));
Q_ASSIGN U5738 ( .B(clk), .A(\g.we_clk [10652]));
Q_ASSIGN U5739 ( .B(clk), .A(\g.we_clk [10651]));
Q_ASSIGN U5740 ( .B(clk), .A(\g.we_clk [10650]));
Q_ASSIGN U5741 ( .B(clk), .A(\g.we_clk [10649]));
Q_ASSIGN U5742 ( .B(clk), .A(\g.we_clk [10648]));
Q_ASSIGN U5743 ( .B(clk), .A(\g.we_clk [10647]));
Q_ASSIGN U5744 ( .B(clk), .A(\g.we_clk [10646]));
Q_ASSIGN U5745 ( .B(clk), .A(\g.we_clk [10645]));
Q_ASSIGN U5746 ( .B(clk), .A(\g.we_clk [10644]));
Q_ASSIGN U5747 ( .B(clk), .A(\g.we_clk [10643]));
Q_ASSIGN U5748 ( .B(clk), .A(\g.we_clk [10642]));
Q_ASSIGN U5749 ( .B(clk), .A(\g.we_clk [10641]));
Q_ASSIGN U5750 ( .B(clk), .A(\g.we_clk [10640]));
Q_ASSIGN U5751 ( .B(clk), .A(\g.we_clk [10639]));
Q_ASSIGN U5752 ( .B(clk), .A(\g.we_clk [10638]));
Q_ASSIGN U5753 ( .B(clk), .A(\g.we_clk [10637]));
Q_ASSIGN U5754 ( .B(clk), .A(\g.we_clk [10636]));
Q_ASSIGN U5755 ( .B(clk), .A(\g.we_clk [10635]));
Q_ASSIGN U5756 ( .B(clk), .A(\g.we_clk [10634]));
Q_ASSIGN U5757 ( .B(clk), .A(\g.we_clk [10633]));
Q_ASSIGN U5758 ( .B(clk), .A(\g.we_clk [10632]));
Q_ASSIGN U5759 ( .B(clk), .A(\g.we_clk [10631]));
Q_ASSIGN U5760 ( .B(clk), .A(\g.we_clk [10630]));
Q_ASSIGN U5761 ( .B(clk), .A(\g.we_clk [10629]));
Q_ASSIGN U5762 ( .B(clk), .A(\g.we_clk [10628]));
Q_ASSIGN U5763 ( .B(clk), .A(\g.we_clk [10627]));
Q_ASSIGN U5764 ( .B(clk), .A(\g.we_clk [10626]));
Q_ASSIGN U5765 ( .B(clk), .A(\g.we_clk [10625]));
Q_ASSIGN U5766 ( .B(clk), .A(\g.we_clk [10624]));
Q_ASSIGN U5767 ( .B(clk), .A(\g.we_clk [10623]));
Q_ASSIGN U5768 ( .B(clk), .A(\g.we_clk [10622]));
Q_ASSIGN U5769 ( .B(clk), .A(\g.we_clk [10621]));
Q_ASSIGN U5770 ( .B(clk), .A(\g.we_clk [10620]));
Q_ASSIGN U5771 ( .B(clk), .A(\g.we_clk [10619]));
Q_ASSIGN U5772 ( .B(clk), .A(\g.we_clk [10618]));
Q_ASSIGN U5773 ( .B(clk), .A(\g.we_clk [10617]));
Q_ASSIGN U5774 ( .B(clk), .A(\g.we_clk [10616]));
Q_ASSIGN U5775 ( .B(clk), .A(\g.we_clk [10615]));
Q_ASSIGN U5776 ( .B(clk), .A(\g.we_clk [10614]));
Q_ASSIGN U5777 ( .B(clk), .A(\g.we_clk [10613]));
Q_ASSIGN U5778 ( .B(clk), .A(\g.we_clk [10612]));
Q_ASSIGN U5779 ( .B(clk), .A(\g.we_clk [10611]));
Q_ASSIGN U5780 ( .B(clk), .A(\g.we_clk [10610]));
Q_ASSIGN U5781 ( .B(clk), .A(\g.we_clk [10609]));
Q_ASSIGN U5782 ( .B(clk), .A(\g.we_clk [10608]));
Q_ASSIGN U5783 ( .B(clk), .A(\g.we_clk [10607]));
Q_ASSIGN U5784 ( .B(clk), .A(\g.we_clk [10606]));
Q_ASSIGN U5785 ( .B(clk), .A(\g.we_clk [10605]));
Q_ASSIGN U5786 ( .B(clk), .A(\g.we_clk [10604]));
Q_ASSIGN U5787 ( .B(clk), .A(\g.we_clk [10603]));
Q_ASSIGN U5788 ( .B(clk), .A(\g.we_clk [10602]));
Q_ASSIGN U5789 ( .B(clk), .A(\g.we_clk [10601]));
Q_ASSIGN U5790 ( .B(clk), .A(\g.we_clk [10600]));
Q_ASSIGN U5791 ( .B(clk), .A(\g.we_clk [10599]));
Q_ASSIGN U5792 ( .B(clk), .A(\g.we_clk [10598]));
Q_ASSIGN U5793 ( .B(clk), .A(\g.we_clk [10597]));
Q_ASSIGN U5794 ( .B(clk), .A(\g.we_clk [10596]));
Q_ASSIGN U5795 ( .B(clk), .A(\g.we_clk [10595]));
Q_ASSIGN U5796 ( .B(clk), .A(\g.we_clk [10594]));
Q_ASSIGN U5797 ( .B(clk), .A(\g.we_clk [10593]));
Q_ASSIGN U5798 ( .B(clk), .A(\g.we_clk [10592]));
Q_ASSIGN U5799 ( .B(clk), .A(\g.we_clk [10591]));
Q_ASSIGN U5800 ( .B(clk), .A(\g.we_clk [10590]));
Q_ASSIGN U5801 ( .B(clk), .A(\g.we_clk [10589]));
Q_ASSIGN U5802 ( .B(clk), .A(\g.we_clk [10588]));
Q_ASSIGN U5803 ( .B(clk), .A(\g.we_clk [10587]));
Q_ASSIGN U5804 ( .B(clk), .A(\g.we_clk [10586]));
Q_ASSIGN U5805 ( .B(clk), .A(\g.we_clk [10585]));
Q_ASSIGN U5806 ( .B(clk), .A(\g.we_clk [10584]));
Q_ASSIGN U5807 ( .B(clk), .A(\g.we_clk [10583]));
Q_ASSIGN U5808 ( .B(clk), .A(\g.we_clk [10582]));
Q_ASSIGN U5809 ( .B(clk), .A(\g.we_clk [10581]));
Q_ASSIGN U5810 ( .B(clk), .A(\g.we_clk [10580]));
Q_ASSIGN U5811 ( .B(clk), .A(\g.we_clk [10579]));
Q_ASSIGN U5812 ( .B(clk), .A(\g.we_clk [10578]));
Q_ASSIGN U5813 ( .B(clk), .A(\g.we_clk [10577]));
Q_ASSIGN U5814 ( .B(clk), .A(\g.we_clk [10576]));
Q_ASSIGN U5815 ( .B(clk), .A(\g.we_clk [10575]));
Q_ASSIGN U5816 ( .B(clk), .A(\g.we_clk [10574]));
Q_ASSIGN U5817 ( .B(clk), .A(\g.we_clk [10573]));
Q_ASSIGN U5818 ( .B(clk), .A(\g.we_clk [10572]));
Q_ASSIGN U5819 ( .B(clk), .A(\g.we_clk [10571]));
Q_ASSIGN U5820 ( .B(clk), .A(\g.we_clk [10570]));
Q_ASSIGN U5821 ( .B(clk), .A(\g.we_clk [10569]));
Q_ASSIGN U5822 ( .B(clk), .A(\g.we_clk [10568]));
Q_ASSIGN U5823 ( .B(clk), .A(\g.we_clk [10567]));
Q_ASSIGN U5824 ( .B(clk), .A(\g.we_clk [10566]));
Q_ASSIGN U5825 ( .B(clk), .A(\g.we_clk [10565]));
Q_ASSIGN U5826 ( .B(clk), .A(\g.we_clk [10564]));
Q_ASSIGN U5827 ( .B(clk), .A(\g.we_clk [10563]));
Q_ASSIGN U5828 ( .B(clk), .A(\g.we_clk [10562]));
Q_ASSIGN U5829 ( .B(clk), .A(\g.we_clk [10561]));
Q_ASSIGN U5830 ( .B(clk), .A(\g.we_clk [10560]));
Q_ASSIGN U5831 ( .B(clk), .A(\g.we_clk [10559]));
Q_ASSIGN U5832 ( .B(clk), .A(\g.we_clk [10558]));
Q_ASSIGN U5833 ( .B(clk), .A(\g.we_clk [10557]));
Q_ASSIGN U5834 ( .B(clk), .A(\g.we_clk [10556]));
Q_ASSIGN U5835 ( .B(clk), .A(\g.we_clk [10555]));
Q_ASSIGN U5836 ( .B(clk), .A(\g.we_clk [10554]));
Q_ASSIGN U5837 ( .B(clk), .A(\g.we_clk [10553]));
Q_ASSIGN U5838 ( .B(clk), .A(\g.we_clk [10552]));
Q_ASSIGN U5839 ( .B(clk), .A(\g.we_clk [10551]));
Q_ASSIGN U5840 ( .B(clk), .A(\g.we_clk [10550]));
Q_ASSIGN U5841 ( .B(clk), .A(\g.we_clk [10549]));
Q_ASSIGN U5842 ( .B(clk), .A(\g.we_clk [10548]));
Q_ASSIGN U5843 ( .B(clk), .A(\g.we_clk [10547]));
Q_ASSIGN U5844 ( .B(clk), .A(\g.we_clk [10546]));
Q_ASSIGN U5845 ( .B(clk), .A(\g.we_clk [10545]));
Q_ASSIGN U5846 ( .B(clk), .A(\g.we_clk [10544]));
Q_ASSIGN U5847 ( .B(clk), .A(\g.we_clk [10543]));
Q_ASSIGN U5848 ( .B(clk), .A(\g.we_clk [10542]));
Q_ASSIGN U5849 ( .B(clk), .A(\g.we_clk [10541]));
Q_ASSIGN U5850 ( .B(clk), .A(\g.we_clk [10540]));
Q_ASSIGN U5851 ( .B(clk), .A(\g.we_clk [10539]));
Q_ASSIGN U5852 ( .B(clk), .A(\g.we_clk [10538]));
Q_ASSIGN U5853 ( .B(clk), .A(\g.we_clk [10537]));
Q_ASSIGN U5854 ( .B(clk), .A(\g.we_clk [10536]));
Q_ASSIGN U5855 ( .B(clk), .A(\g.we_clk [10535]));
Q_ASSIGN U5856 ( .B(clk), .A(\g.we_clk [10534]));
Q_ASSIGN U5857 ( .B(clk), .A(\g.we_clk [10533]));
Q_ASSIGN U5858 ( .B(clk), .A(\g.we_clk [10532]));
Q_ASSIGN U5859 ( .B(clk), .A(\g.we_clk [10531]));
Q_ASSIGN U5860 ( .B(clk), .A(\g.we_clk [10530]));
Q_ASSIGN U5861 ( .B(clk), .A(\g.we_clk [10529]));
Q_ASSIGN U5862 ( .B(clk), .A(\g.we_clk [10528]));
Q_ASSIGN U5863 ( .B(clk), .A(\g.we_clk [10527]));
Q_ASSIGN U5864 ( .B(clk), .A(\g.we_clk [10526]));
Q_ASSIGN U5865 ( .B(clk), .A(\g.we_clk [10525]));
Q_ASSIGN U5866 ( .B(clk), .A(\g.we_clk [10524]));
Q_ASSIGN U5867 ( .B(clk), .A(\g.we_clk [10523]));
Q_ASSIGN U5868 ( .B(clk), .A(\g.we_clk [10522]));
Q_ASSIGN U5869 ( .B(clk), .A(\g.we_clk [10521]));
Q_ASSIGN U5870 ( .B(clk), .A(\g.we_clk [10520]));
Q_ASSIGN U5871 ( .B(clk), .A(\g.we_clk [10519]));
Q_ASSIGN U5872 ( .B(clk), .A(\g.we_clk [10518]));
Q_ASSIGN U5873 ( .B(clk), .A(\g.we_clk [10517]));
Q_ASSIGN U5874 ( .B(clk), .A(\g.we_clk [10516]));
Q_ASSIGN U5875 ( .B(clk), .A(\g.we_clk [10515]));
Q_ASSIGN U5876 ( .B(clk), .A(\g.we_clk [10514]));
Q_ASSIGN U5877 ( .B(clk), .A(\g.we_clk [10513]));
Q_ASSIGN U5878 ( .B(clk), .A(\g.we_clk [10512]));
Q_ASSIGN U5879 ( .B(clk), .A(\g.we_clk [10511]));
Q_ASSIGN U5880 ( .B(clk), .A(\g.we_clk [10510]));
Q_ASSIGN U5881 ( .B(clk), .A(\g.we_clk [10509]));
Q_ASSIGN U5882 ( .B(clk), .A(\g.we_clk [10508]));
Q_ASSIGN U5883 ( .B(clk), .A(\g.we_clk [10507]));
Q_ASSIGN U5884 ( .B(clk), .A(\g.we_clk [10506]));
Q_ASSIGN U5885 ( .B(clk), .A(\g.we_clk [10505]));
Q_ASSIGN U5886 ( .B(clk), .A(\g.we_clk [10504]));
Q_ASSIGN U5887 ( .B(clk), .A(\g.we_clk [10503]));
Q_ASSIGN U5888 ( .B(clk), .A(\g.we_clk [10502]));
Q_ASSIGN U5889 ( .B(clk), .A(\g.we_clk [10501]));
Q_ASSIGN U5890 ( .B(clk), .A(\g.we_clk [10500]));
Q_ASSIGN U5891 ( .B(clk), .A(\g.we_clk [10499]));
Q_ASSIGN U5892 ( .B(clk), .A(\g.we_clk [10498]));
Q_ASSIGN U5893 ( .B(clk), .A(\g.we_clk [10497]));
Q_ASSIGN U5894 ( .B(clk), .A(\g.we_clk [10496]));
Q_ASSIGN U5895 ( .B(clk), .A(\g.we_clk [10495]));
Q_ASSIGN U5896 ( .B(clk), .A(\g.we_clk [10494]));
Q_ASSIGN U5897 ( .B(clk), .A(\g.we_clk [10493]));
Q_ASSIGN U5898 ( .B(clk), .A(\g.we_clk [10492]));
Q_ASSIGN U5899 ( .B(clk), .A(\g.we_clk [10491]));
Q_ASSIGN U5900 ( .B(clk), .A(\g.we_clk [10490]));
Q_ASSIGN U5901 ( .B(clk), .A(\g.we_clk [10489]));
Q_ASSIGN U5902 ( .B(clk), .A(\g.we_clk [10488]));
Q_ASSIGN U5903 ( .B(clk), .A(\g.we_clk [10487]));
Q_ASSIGN U5904 ( .B(clk), .A(\g.we_clk [10486]));
Q_ASSIGN U5905 ( .B(clk), .A(\g.we_clk [10485]));
Q_ASSIGN U5906 ( .B(clk), .A(\g.we_clk [10484]));
Q_ASSIGN U5907 ( .B(clk), .A(\g.we_clk [10483]));
Q_ASSIGN U5908 ( .B(clk), .A(\g.we_clk [10482]));
Q_ASSIGN U5909 ( .B(clk), .A(\g.we_clk [10481]));
Q_ASSIGN U5910 ( .B(clk), .A(\g.we_clk [10480]));
Q_ASSIGN U5911 ( .B(clk), .A(\g.we_clk [10479]));
Q_ASSIGN U5912 ( .B(clk), .A(\g.we_clk [10478]));
Q_ASSIGN U5913 ( .B(clk), .A(\g.we_clk [10477]));
Q_ASSIGN U5914 ( .B(clk), .A(\g.we_clk [10476]));
Q_ASSIGN U5915 ( .B(clk), .A(\g.we_clk [10475]));
Q_ASSIGN U5916 ( .B(clk), .A(\g.we_clk [10474]));
Q_ASSIGN U5917 ( .B(clk), .A(\g.we_clk [10473]));
Q_ASSIGN U5918 ( .B(clk), .A(\g.we_clk [10472]));
Q_ASSIGN U5919 ( .B(clk), .A(\g.we_clk [10471]));
Q_ASSIGN U5920 ( .B(clk), .A(\g.we_clk [10470]));
Q_ASSIGN U5921 ( .B(clk), .A(\g.we_clk [10469]));
Q_ASSIGN U5922 ( .B(clk), .A(\g.we_clk [10468]));
Q_ASSIGN U5923 ( .B(clk), .A(\g.we_clk [10467]));
Q_ASSIGN U5924 ( .B(clk), .A(\g.we_clk [10466]));
Q_ASSIGN U5925 ( .B(clk), .A(\g.we_clk [10465]));
Q_ASSIGN U5926 ( .B(clk), .A(\g.we_clk [10464]));
Q_ASSIGN U5927 ( .B(clk), .A(\g.we_clk [10463]));
Q_ASSIGN U5928 ( .B(clk), .A(\g.we_clk [10462]));
Q_ASSIGN U5929 ( .B(clk), .A(\g.we_clk [10461]));
Q_ASSIGN U5930 ( .B(clk), .A(\g.we_clk [10460]));
Q_ASSIGN U5931 ( .B(clk), .A(\g.we_clk [10459]));
Q_ASSIGN U5932 ( .B(clk), .A(\g.we_clk [10458]));
Q_ASSIGN U5933 ( .B(clk), .A(\g.we_clk [10457]));
Q_ASSIGN U5934 ( .B(clk), .A(\g.we_clk [10456]));
Q_ASSIGN U5935 ( .B(clk), .A(\g.we_clk [10455]));
Q_ASSIGN U5936 ( .B(clk), .A(\g.we_clk [10454]));
Q_ASSIGN U5937 ( .B(clk), .A(\g.we_clk [10453]));
Q_ASSIGN U5938 ( .B(clk), .A(\g.we_clk [10452]));
Q_ASSIGN U5939 ( .B(clk), .A(\g.we_clk [10451]));
Q_ASSIGN U5940 ( .B(clk), .A(\g.we_clk [10450]));
Q_ASSIGN U5941 ( .B(clk), .A(\g.we_clk [10449]));
Q_ASSIGN U5942 ( .B(clk), .A(\g.we_clk [10448]));
Q_ASSIGN U5943 ( .B(clk), .A(\g.we_clk [10447]));
Q_ASSIGN U5944 ( .B(clk), .A(\g.we_clk [10446]));
Q_ASSIGN U5945 ( .B(clk), .A(\g.we_clk [10445]));
Q_ASSIGN U5946 ( .B(clk), .A(\g.we_clk [10444]));
Q_ASSIGN U5947 ( .B(clk), .A(\g.we_clk [10443]));
Q_ASSIGN U5948 ( .B(clk), .A(\g.we_clk [10442]));
Q_ASSIGN U5949 ( .B(clk), .A(\g.we_clk [10441]));
Q_ASSIGN U5950 ( .B(clk), .A(\g.we_clk [10440]));
Q_ASSIGN U5951 ( .B(clk), .A(\g.we_clk [10439]));
Q_ASSIGN U5952 ( .B(clk), .A(\g.we_clk [10438]));
Q_ASSIGN U5953 ( .B(clk), .A(\g.we_clk [10437]));
Q_ASSIGN U5954 ( .B(clk), .A(\g.we_clk [10436]));
Q_ASSIGN U5955 ( .B(clk), .A(\g.we_clk [10435]));
Q_ASSIGN U5956 ( .B(clk), .A(\g.we_clk [10434]));
Q_ASSIGN U5957 ( .B(clk), .A(\g.we_clk [10433]));
Q_ASSIGN U5958 ( .B(clk), .A(\g.we_clk [10432]));
Q_ASSIGN U5959 ( .B(clk), .A(\g.we_clk [10431]));
Q_ASSIGN U5960 ( .B(clk), .A(\g.we_clk [10430]));
Q_ASSIGN U5961 ( .B(clk), .A(\g.we_clk [10429]));
Q_ASSIGN U5962 ( .B(clk), .A(\g.we_clk [10428]));
Q_ASSIGN U5963 ( .B(clk), .A(\g.we_clk [10427]));
Q_ASSIGN U5964 ( .B(clk), .A(\g.we_clk [10426]));
Q_ASSIGN U5965 ( .B(clk), .A(\g.we_clk [10425]));
Q_ASSIGN U5966 ( .B(clk), .A(\g.we_clk [10424]));
Q_ASSIGN U5967 ( .B(clk), .A(\g.we_clk [10423]));
Q_ASSIGN U5968 ( .B(clk), .A(\g.we_clk [10422]));
Q_ASSIGN U5969 ( .B(clk), .A(\g.we_clk [10421]));
Q_ASSIGN U5970 ( .B(clk), .A(\g.we_clk [10420]));
Q_ASSIGN U5971 ( .B(clk), .A(\g.we_clk [10419]));
Q_ASSIGN U5972 ( .B(clk), .A(\g.we_clk [10418]));
Q_ASSIGN U5973 ( .B(clk), .A(\g.we_clk [10417]));
Q_ASSIGN U5974 ( .B(clk), .A(\g.we_clk [10416]));
Q_ASSIGN U5975 ( .B(clk), .A(\g.we_clk [10415]));
Q_ASSIGN U5976 ( .B(clk), .A(\g.we_clk [10414]));
Q_ASSIGN U5977 ( .B(clk), .A(\g.we_clk [10413]));
Q_ASSIGN U5978 ( .B(clk), .A(\g.we_clk [10412]));
Q_ASSIGN U5979 ( .B(clk), .A(\g.we_clk [10411]));
Q_ASSIGN U5980 ( .B(clk), .A(\g.we_clk [10410]));
Q_ASSIGN U5981 ( .B(clk), .A(\g.we_clk [10409]));
Q_ASSIGN U5982 ( .B(clk), .A(\g.we_clk [10408]));
Q_ASSIGN U5983 ( .B(clk), .A(\g.we_clk [10407]));
Q_ASSIGN U5984 ( .B(clk), .A(\g.we_clk [10406]));
Q_ASSIGN U5985 ( .B(clk), .A(\g.we_clk [10405]));
Q_ASSIGN U5986 ( .B(clk), .A(\g.we_clk [10404]));
Q_ASSIGN U5987 ( .B(clk), .A(\g.we_clk [10403]));
Q_ASSIGN U5988 ( .B(clk), .A(\g.we_clk [10402]));
Q_ASSIGN U5989 ( .B(clk), .A(\g.we_clk [10401]));
Q_ASSIGN U5990 ( .B(clk), .A(\g.we_clk [10400]));
Q_ASSIGN U5991 ( .B(clk), .A(\g.we_clk [10399]));
Q_ASSIGN U5992 ( .B(clk), .A(\g.we_clk [10398]));
Q_ASSIGN U5993 ( .B(clk), .A(\g.we_clk [10397]));
Q_ASSIGN U5994 ( .B(clk), .A(\g.we_clk [10396]));
Q_ASSIGN U5995 ( .B(clk), .A(\g.we_clk [10395]));
Q_ASSIGN U5996 ( .B(clk), .A(\g.we_clk [10394]));
Q_ASSIGN U5997 ( .B(clk), .A(\g.we_clk [10393]));
Q_ASSIGN U5998 ( .B(clk), .A(\g.we_clk [10392]));
Q_ASSIGN U5999 ( .B(clk), .A(\g.we_clk [10391]));
Q_ASSIGN U6000 ( .B(clk), .A(\g.we_clk [10390]));
Q_ASSIGN U6001 ( .B(clk), .A(\g.we_clk [10389]));
Q_ASSIGN U6002 ( .B(clk), .A(\g.we_clk [10388]));
Q_ASSIGN U6003 ( .B(clk), .A(\g.we_clk [10387]));
Q_ASSIGN U6004 ( .B(clk), .A(\g.we_clk [10386]));
Q_ASSIGN U6005 ( .B(clk), .A(\g.we_clk [10385]));
Q_ASSIGN U6006 ( .B(clk), .A(\g.we_clk [10384]));
Q_ASSIGN U6007 ( .B(clk), .A(\g.we_clk [10383]));
Q_ASSIGN U6008 ( .B(clk), .A(\g.we_clk [10382]));
Q_ASSIGN U6009 ( .B(clk), .A(\g.we_clk [10381]));
Q_ASSIGN U6010 ( .B(clk), .A(\g.we_clk [10380]));
Q_ASSIGN U6011 ( .B(clk), .A(\g.we_clk [10379]));
Q_ASSIGN U6012 ( .B(clk), .A(\g.we_clk [10378]));
Q_ASSIGN U6013 ( .B(clk), .A(\g.we_clk [10377]));
Q_ASSIGN U6014 ( .B(clk), .A(\g.we_clk [10376]));
Q_ASSIGN U6015 ( .B(clk), .A(\g.we_clk [10375]));
Q_ASSIGN U6016 ( .B(clk), .A(\g.we_clk [10374]));
Q_ASSIGN U6017 ( .B(clk), .A(\g.we_clk [10373]));
Q_ASSIGN U6018 ( .B(clk), .A(\g.we_clk [10372]));
Q_ASSIGN U6019 ( .B(clk), .A(\g.we_clk [10371]));
Q_ASSIGN U6020 ( .B(clk), .A(\g.we_clk [10370]));
Q_ASSIGN U6021 ( .B(clk), .A(\g.we_clk [10369]));
Q_ASSIGN U6022 ( .B(clk), .A(\g.we_clk [10368]));
Q_ASSIGN U6023 ( .B(clk), .A(\g.we_clk [10367]));
Q_ASSIGN U6024 ( .B(clk), .A(\g.we_clk [10366]));
Q_ASSIGN U6025 ( .B(clk), .A(\g.we_clk [10365]));
Q_ASSIGN U6026 ( .B(clk), .A(\g.we_clk [10364]));
Q_ASSIGN U6027 ( .B(clk), .A(\g.we_clk [10363]));
Q_ASSIGN U6028 ( .B(clk), .A(\g.we_clk [10362]));
Q_ASSIGN U6029 ( .B(clk), .A(\g.we_clk [10361]));
Q_ASSIGN U6030 ( .B(clk), .A(\g.we_clk [10360]));
Q_ASSIGN U6031 ( .B(clk), .A(\g.we_clk [10359]));
Q_ASSIGN U6032 ( .B(clk), .A(\g.we_clk [10358]));
Q_ASSIGN U6033 ( .B(clk), .A(\g.we_clk [10357]));
Q_ASSIGN U6034 ( .B(clk), .A(\g.we_clk [10356]));
Q_ASSIGN U6035 ( .B(clk), .A(\g.we_clk [10355]));
Q_ASSIGN U6036 ( .B(clk), .A(\g.we_clk [10354]));
Q_ASSIGN U6037 ( .B(clk), .A(\g.we_clk [10353]));
Q_ASSIGN U6038 ( .B(clk), .A(\g.we_clk [10352]));
Q_ASSIGN U6039 ( .B(clk), .A(\g.we_clk [10351]));
Q_ASSIGN U6040 ( .B(clk), .A(\g.we_clk [10350]));
Q_ASSIGN U6041 ( .B(clk), .A(\g.we_clk [10349]));
Q_ASSIGN U6042 ( .B(clk), .A(\g.we_clk [10348]));
Q_ASSIGN U6043 ( .B(clk), .A(\g.we_clk [10347]));
Q_ASSIGN U6044 ( .B(clk), .A(\g.we_clk [10346]));
Q_ASSIGN U6045 ( .B(clk), .A(\g.we_clk [10345]));
Q_ASSIGN U6046 ( .B(clk), .A(\g.we_clk [10344]));
Q_ASSIGN U6047 ( .B(clk), .A(\g.we_clk [10343]));
Q_ASSIGN U6048 ( .B(clk), .A(\g.we_clk [10342]));
Q_ASSIGN U6049 ( .B(clk), .A(\g.we_clk [10341]));
Q_ASSIGN U6050 ( .B(clk), .A(\g.we_clk [10340]));
Q_ASSIGN U6051 ( .B(clk), .A(\g.we_clk [10339]));
Q_ASSIGN U6052 ( .B(clk), .A(\g.we_clk [10338]));
Q_ASSIGN U6053 ( .B(clk), .A(\g.we_clk [10337]));
Q_ASSIGN U6054 ( .B(clk), .A(\g.we_clk [10336]));
Q_ASSIGN U6055 ( .B(clk), .A(\g.we_clk [10335]));
Q_ASSIGN U6056 ( .B(clk), .A(\g.we_clk [10334]));
Q_ASSIGN U6057 ( .B(clk), .A(\g.we_clk [10333]));
Q_ASSIGN U6058 ( .B(clk), .A(\g.we_clk [10332]));
Q_ASSIGN U6059 ( .B(clk), .A(\g.we_clk [10331]));
Q_ASSIGN U6060 ( .B(clk), .A(\g.we_clk [10330]));
Q_ASSIGN U6061 ( .B(clk), .A(\g.we_clk [10329]));
Q_ASSIGN U6062 ( .B(clk), .A(\g.we_clk [10328]));
Q_ASSIGN U6063 ( .B(clk), .A(\g.we_clk [10327]));
Q_ASSIGN U6064 ( .B(clk), .A(\g.we_clk [10326]));
Q_ASSIGN U6065 ( .B(clk), .A(\g.we_clk [10325]));
Q_ASSIGN U6066 ( .B(clk), .A(\g.we_clk [10324]));
Q_ASSIGN U6067 ( .B(clk), .A(\g.we_clk [10323]));
Q_ASSIGN U6068 ( .B(clk), .A(\g.we_clk [10322]));
Q_ASSIGN U6069 ( .B(clk), .A(\g.we_clk [10321]));
Q_ASSIGN U6070 ( .B(clk), .A(\g.we_clk [10320]));
Q_ASSIGN U6071 ( .B(clk), .A(\g.we_clk [10319]));
Q_ASSIGN U6072 ( .B(clk), .A(\g.we_clk [10318]));
Q_ASSIGN U6073 ( .B(clk), .A(\g.we_clk [10317]));
Q_ASSIGN U6074 ( .B(clk), .A(\g.we_clk [10316]));
Q_ASSIGN U6075 ( .B(clk), .A(\g.we_clk [10315]));
Q_ASSIGN U6076 ( .B(clk), .A(\g.we_clk [10314]));
Q_ASSIGN U6077 ( .B(clk), .A(\g.we_clk [10313]));
Q_ASSIGN U6078 ( .B(clk), .A(\g.we_clk [10312]));
Q_ASSIGN U6079 ( .B(clk), .A(\g.we_clk [10311]));
Q_ASSIGN U6080 ( .B(clk), .A(\g.we_clk [10310]));
Q_ASSIGN U6081 ( .B(clk), .A(\g.we_clk [10309]));
Q_ASSIGN U6082 ( .B(clk), .A(\g.we_clk [10308]));
Q_ASSIGN U6083 ( .B(clk), .A(\g.we_clk [10307]));
Q_ASSIGN U6084 ( .B(clk), .A(\g.we_clk [10306]));
Q_ASSIGN U6085 ( .B(clk), .A(\g.we_clk [10305]));
Q_ASSIGN U6086 ( .B(clk), .A(\g.we_clk [10304]));
Q_ASSIGN U6087 ( .B(clk), .A(\g.we_clk [10303]));
Q_ASSIGN U6088 ( .B(clk), .A(\g.we_clk [10302]));
Q_ASSIGN U6089 ( .B(clk), .A(\g.we_clk [10301]));
Q_ASSIGN U6090 ( .B(clk), .A(\g.we_clk [10300]));
Q_ASSIGN U6091 ( .B(clk), .A(\g.we_clk [10299]));
Q_ASSIGN U6092 ( .B(clk), .A(\g.we_clk [10298]));
Q_ASSIGN U6093 ( .B(clk), .A(\g.we_clk [10297]));
Q_ASSIGN U6094 ( .B(clk), .A(\g.we_clk [10296]));
Q_ASSIGN U6095 ( .B(clk), .A(\g.we_clk [10295]));
Q_ASSIGN U6096 ( .B(clk), .A(\g.we_clk [10294]));
Q_ASSIGN U6097 ( .B(clk), .A(\g.we_clk [10293]));
Q_ASSIGN U6098 ( .B(clk), .A(\g.we_clk [10292]));
Q_ASSIGN U6099 ( .B(clk), .A(\g.we_clk [10291]));
Q_ASSIGN U6100 ( .B(clk), .A(\g.we_clk [10290]));
Q_ASSIGN U6101 ( .B(clk), .A(\g.we_clk [10289]));
Q_ASSIGN U6102 ( .B(clk), .A(\g.we_clk [10288]));
Q_ASSIGN U6103 ( .B(clk), .A(\g.we_clk [10287]));
Q_ASSIGN U6104 ( .B(clk), .A(\g.we_clk [10286]));
Q_ASSIGN U6105 ( .B(clk), .A(\g.we_clk [10285]));
Q_ASSIGN U6106 ( .B(clk), .A(\g.we_clk [10284]));
Q_ASSIGN U6107 ( .B(clk), .A(\g.we_clk [10283]));
Q_ASSIGN U6108 ( .B(clk), .A(\g.we_clk [10282]));
Q_ASSIGN U6109 ( .B(clk), .A(\g.we_clk [10281]));
Q_ASSIGN U6110 ( .B(clk), .A(\g.we_clk [10280]));
Q_ASSIGN U6111 ( .B(clk), .A(\g.we_clk [10279]));
Q_ASSIGN U6112 ( .B(clk), .A(\g.we_clk [10278]));
Q_ASSIGN U6113 ( .B(clk), .A(\g.we_clk [10277]));
Q_ASSIGN U6114 ( .B(clk), .A(\g.we_clk [10276]));
Q_ASSIGN U6115 ( .B(clk), .A(\g.we_clk [10275]));
Q_ASSIGN U6116 ( .B(clk), .A(\g.we_clk [10274]));
Q_ASSIGN U6117 ( .B(clk), .A(\g.we_clk [10273]));
Q_ASSIGN U6118 ( .B(clk), .A(\g.we_clk [10272]));
Q_ASSIGN U6119 ( .B(clk), .A(\g.we_clk [10271]));
Q_ASSIGN U6120 ( .B(clk), .A(\g.we_clk [10270]));
Q_ASSIGN U6121 ( .B(clk), .A(\g.we_clk [10269]));
Q_ASSIGN U6122 ( .B(clk), .A(\g.we_clk [10268]));
Q_ASSIGN U6123 ( .B(clk), .A(\g.we_clk [10267]));
Q_ASSIGN U6124 ( .B(clk), .A(\g.we_clk [10266]));
Q_ASSIGN U6125 ( .B(clk), .A(\g.we_clk [10265]));
Q_ASSIGN U6126 ( .B(clk), .A(\g.we_clk [10264]));
Q_ASSIGN U6127 ( .B(clk), .A(\g.we_clk [10263]));
Q_ASSIGN U6128 ( .B(clk), .A(\g.we_clk [10262]));
Q_ASSIGN U6129 ( .B(clk), .A(\g.we_clk [10261]));
Q_ASSIGN U6130 ( .B(clk), .A(\g.we_clk [10260]));
Q_ASSIGN U6131 ( .B(clk), .A(\g.we_clk [10259]));
Q_ASSIGN U6132 ( .B(clk), .A(\g.we_clk [10258]));
Q_ASSIGN U6133 ( .B(clk), .A(\g.we_clk [10257]));
Q_ASSIGN U6134 ( .B(clk), .A(\g.we_clk [10256]));
Q_ASSIGN U6135 ( .B(clk), .A(\g.we_clk [10255]));
Q_ASSIGN U6136 ( .B(clk), .A(\g.we_clk [10254]));
Q_ASSIGN U6137 ( .B(clk), .A(\g.we_clk [10253]));
Q_ASSIGN U6138 ( .B(clk), .A(\g.we_clk [10252]));
Q_ASSIGN U6139 ( .B(clk), .A(\g.we_clk [10251]));
Q_ASSIGN U6140 ( .B(clk), .A(\g.we_clk [10250]));
Q_ASSIGN U6141 ( .B(clk), .A(\g.we_clk [10249]));
Q_ASSIGN U6142 ( .B(clk), .A(\g.we_clk [10248]));
Q_ASSIGN U6143 ( .B(clk), .A(\g.we_clk [10247]));
Q_ASSIGN U6144 ( .B(clk), .A(\g.we_clk [10246]));
Q_ASSIGN U6145 ( .B(clk), .A(\g.we_clk [10245]));
Q_ASSIGN U6146 ( .B(clk), .A(\g.we_clk [10244]));
Q_ASSIGN U6147 ( .B(clk), .A(\g.we_clk [10243]));
Q_ASSIGN U6148 ( .B(clk), .A(\g.we_clk [10242]));
Q_ASSIGN U6149 ( .B(clk), .A(\g.we_clk [10241]));
Q_ASSIGN U6150 ( .B(clk), .A(\g.we_clk [10240]));
Q_ASSIGN U6151 ( .B(clk), .A(\g.we_clk [10239]));
Q_ASSIGN U6152 ( .B(clk), .A(\g.we_clk [10238]));
Q_ASSIGN U6153 ( .B(clk), .A(\g.we_clk [10237]));
Q_ASSIGN U6154 ( .B(clk), .A(\g.we_clk [10236]));
Q_ASSIGN U6155 ( .B(clk), .A(\g.we_clk [10235]));
Q_ASSIGN U6156 ( .B(clk), .A(\g.we_clk [10234]));
Q_ASSIGN U6157 ( .B(clk), .A(\g.we_clk [10233]));
Q_ASSIGN U6158 ( .B(clk), .A(\g.we_clk [10232]));
Q_ASSIGN U6159 ( .B(clk), .A(\g.we_clk [10231]));
Q_ASSIGN U6160 ( .B(clk), .A(\g.we_clk [10230]));
Q_ASSIGN U6161 ( .B(clk), .A(\g.we_clk [10229]));
Q_ASSIGN U6162 ( .B(clk), .A(\g.we_clk [10228]));
Q_ASSIGN U6163 ( .B(clk), .A(\g.we_clk [10227]));
Q_ASSIGN U6164 ( .B(clk), .A(\g.we_clk [10226]));
Q_ASSIGN U6165 ( .B(clk), .A(\g.we_clk [10225]));
Q_ASSIGN U6166 ( .B(clk), .A(\g.we_clk [10224]));
Q_ASSIGN U6167 ( .B(clk), .A(\g.we_clk [10223]));
Q_ASSIGN U6168 ( .B(clk), .A(\g.we_clk [10222]));
Q_ASSIGN U6169 ( .B(clk), .A(\g.we_clk [10221]));
Q_ASSIGN U6170 ( .B(clk), .A(\g.we_clk [10220]));
Q_ASSIGN U6171 ( .B(clk), .A(\g.we_clk [10219]));
Q_ASSIGN U6172 ( .B(clk), .A(\g.we_clk [10218]));
Q_ASSIGN U6173 ( .B(clk), .A(\g.we_clk [10217]));
Q_ASSIGN U6174 ( .B(clk), .A(\g.we_clk [10216]));
Q_ASSIGN U6175 ( .B(clk), .A(\g.we_clk [10215]));
Q_ASSIGN U6176 ( .B(clk), .A(\g.we_clk [10214]));
Q_ASSIGN U6177 ( .B(clk), .A(\g.we_clk [10213]));
Q_ASSIGN U6178 ( .B(clk), .A(\g.we_clk [10212]));
Q_ASSIGN U6179 ( .B(clk), .A(\g.we_clk [10211]));
Q_ASSIGN U6180 ( .B(clk), .A(\g.we_clk [10210]));
Q_ASSIGN U6181 ( .B(clk), .A(\g.we_clk [10209]));
Q_ASSIGN U6182 ( .B(clk), .A(\g.we_clk [10208]));
Q_ASSIGN U6183 ( .B(clk), .A(\g.we_clk [10207]));
Q_ASSIGN U6184 ( .B(clk), .A(\g.we_clk [10206]));
Q_ASSIGN U6185 ( .B(clk), .A(\g.we_clk [10205]));
Q_ASSIGN U6186 ( .B(clk), .A(\g.we_clk [10204]));
Q_ASSIGN U6187 ( .B(clk), .A(\g.we_clk [10203]));
Q_ASSIGN U6188 ( .B(clk), .A(\g.we_clk [10202]));
Q_ASSIGN U6189 ( .B(clk), .A(\g.we_clk [10201]));
Q_ASSIGN U6190 ( .B(clk), .A(\g.we_clk [10200]));
Q_ASSIGN U6191 ( .B(clk), .A(\g.we_clk [10199]));
Q_ASSIGN U6192 ( .B(clk), .A(\g.we_clk [10198]));
Q_ASSIGN U6193 ( .B(clk), .A(\g.we_clk [10197]));
Q_ASSIGN U6194 ( .B(clk), .A(\g.we_clk [10196]));
Q_ASSIGN U6195 ( .B(clk), .A(\g.we_clk [10195]));
Q_ASSIGN U6196 ( .B(clk), .A(\g.we_clk [10194]));
Q_ASSIGN U6197 ( .B(clk), .A(\g.we_clk [10193]));
Q_ASSIGN U6198 ( .B(clk), .A(\g.we_clk [10192]));
Q_ASSIGN U6199 ( .B(clk), .A(\g.we_clk [10191]));
Q_ASSIGN U6200 ( .B(clk), .A(\g.we_clk [10190]));
Q_ASSIGN U6201 ( .B(clk), .A(\g.we_clk [10189]));
Q_ASSIGN U6202 ( .B(clk), .A(\g.we_clk [10188]));
Q_ASSIGN U6203 ( .B(clk), .A(\g.we_clk [10187]));
Q_ASSIGN U6204 ( .B(clk), .A(\g.we_clk [10186]));
Q_ASSIGN U6205 ( .B(clk), .A(\g.we_clk [10185]));
Q_ASSIGN U6206 ( .B(clk), .A(\g.we_clk [10184]));
Q_ASSIGN U6207 ( .B(clk), .A(\g.we_clk [10183]));
Q_ASSIGN U6208 ( .B(clk), .A(\g.we_clk [10182]));
Q_ASSIGN U6209 ( .B(clk), .A(\g.we_clk [10181]));
Q_ASSIGN U6210 ( .B(clk), .A(\g.we_clk [10180]));
Q_ASSIGN U6211 ( .B(clk), .A(\g.we_clk [10179]));
Q_ASSIGN U6212 ( .B(clk), .A(\g.we_clk [10178]));
Q_ASSIGN U6213 ( .B(clk), .A(\g.we_clk [10177]));
Q_ASSIGN U6214 ( .B(clk), .A(\g.we_clk [10176]));
Q_ASSIGN U6215 ( .B(clk), .A(\g.we_clk [10175]));
Q_ASSIGN U6216 ( .B(clk), .A(\g.we_clk [10174]));
Q_ASSIGN U6217 ( .B(clk), .A(\g.we_clk [10173]));
Q_ASSIGN U6218 ( .B(clk), .A(\g.we_clk [10172]));
Q_ASSIGN U6219 ( .B(clk), .A(\g.we_clk [10171]));
Q_ASSIGN U6220 ( .B(clk), .A(\g.we_clk [10170]));
Q_ASSIGN U6221 ( .B(clk), .A(\g.we_clk [10169]));
Q_ASSIGN U6222 ( .B(clk), .A(\g.we_clk [10168]));
Q_ASSIGN U6223 ( .B(clk), .A(\g.we_clk [10167]));
Q_ASSIGN U6224 ( .B(clk), .A(\g.we_clk [10166]));
Q_ASSIGN U6225 ( .B(clk), .A(\g.we_clk [10165]));
Q_ASSIGN U6226 ( .B(clk), .A(\g.we_clk [10164]));
Q_ASSIGN U6227 ( .B(clk), .A(\g.we_clk [10163]));
Q_ASSIGN U6228 ( .B(clk), .A(\g.we_clk [10162]));
Q_ASSIGN U6229 ( .B(clk), .A(\g.we_clk [10161]));
Q_ASSIGN U6230 ( .B(clk), .A(\g.we_clk [10160]));
Q_ASSIGN U6231 ( .B(clk), .A(\g.we_clk [10159]));
Q_ASSIGN U6232 ( .B(clk), .A(\g.we_clk [10158]));
Q_ASSIGN U6233 ( .B(clk), .A(\g.we_clk [10157]));
Q_ASSIGN U6234 ( .B(clk), .A(\g.we_clk [10156]));
Q_ASSIGN U6235 ( .B(clk), .A(\g.we_clk [10155]));
Q_ASSIGN U6236 ( .B(clk), .A(\g.we_clk [10154]));
Q_ASSIGN U6237 ( .B(clk), .A(\g.we_clk [10153]));
Q_ASSIGN U6238 ( .B(clk), .A(\g.we_clk [10152]));
Q_ASSIGN U6239 ( .B(clk), .A(\g.we_clk [10151]));
Q_ASSIGN U6240 ( .B(clk), .A(\g.we_clk [10150]));
Q_ASSIGN U6241 ( .B(clk), .A(\g.we_clk [10149]));
Q_ASSIGN U6242 ( .B(clk), .A(\g.we_clk [10148]));
Q_ASSIGN U6243 ( .B(clk), .A(\g.we_clk [10147]));
Q_ASSIGN U6244 ( .B(clk), .A(\g.we_clk [10146]));
Q_ASSIGN U6245 ( .B(clk), .A(\g.we_clk [10145]));
Q_ASSIGN U6246 ( .B(clk), .A(\g.we_clk [10144]));
Q_ASSIGN U6247 ( .B(clk), .A(\g.we_clk [10143]));
Q_ASSIGN U6248 ( .B(clk), .A(\g.we_clk [10142]));
Q_ASSIGN U6249 ( .B(clk), .A(\g.we_clk [10141]));
Q_ASSIGN U6250 ( .B(clk), .A(\g.we_clk [10140]));
Q_ASSIGN U6251 ( .B(clk), .A(\g.we_clk [10139]));
Q_ASSIGN U6252 ( .B(clk), .A(\g.we_clk [10138]));
Q_ASSIGN U6253 ( .B(clk), .A(\g.we_clk [10137]));
Q_ASSIGN U6254 ( .B(clk), .A(\g.we_clk [10136]));
Q_ASSIGN U6255 ( .B(clk), .A(\g.we_clk [10135]));
Q_ASSIGN U6256 ( .B(clk), .A(\g.we_clk [10134]));
Q_ASSIGN U6257 ( .B(clk), .A(\g.we_clk [10133]));
Q_ASSIGN U6258 ( .B(clk), .A(\g.we_clk [10132]));
Q_ASSIGN U6259 ( .B(clk), .A(\g.we_clk [10131]));
Q_ASSIGN U6260 ( .B(clk), .A(\g.we_clk [10130]));
Q_ASSIGN U6261 ( .B(clk), .A(\g.we_clk [10129]));
Q_ASSIGN U6262 ( .B(clk), .A(\g.we_clk [10128]));
Q_ASSIGN U6263 ( .B(clk), .A(\g.we_clk [10127]));
Q_ASSIGN U6264 ( .B(clk), .A(\g.we_clk [10126]));
Q_ASSIGN U6265 ( .B(clk), .A(\g.we_clk [10125]));
Q_ASSIGN U6266 ( .B(clk), .A(\g.we_clk [10124]));
Q_ASSIGN U6267 ( .B(clk), .A(\g.we_clk [10123]));
Q_ASSIGN U6268 ( .B(clk), .A(\g.we_clk [10122]));
Q_ASSIGN U6269 ( .B(clk), .A(\g.we_clk [10121]));
Q_ASSIGN U6270 ( .B(clk), .A(\g.we_clk [10120]));
Q_ASSIGN U6271 ( .B(clk), .A(\g.we_clk [10119]));
Q_ASSIGN U6272 ( .B(clk), .A(\g.we_clk [10118]));
Q_ASSIGN U6273 ( .B(clk), .A(\g.we_clk [10117]));
Q_ASSIGN U6274 ( .B(clk), .A(\g.we_clk [10116]));
Q_ASSIGN U6275 ( .B(clk), .A(\g.we_clk [10115]));
Q_ASSIGN U6276 ( .B(clk), .A(\g.we_clk [10114]));
Q_ASSIGN U6277 ( .B(clk), .A(\g.we_clk [10113]));
Q_ASSIGN U6278 ( .B(clk), .A(\g.we_clk [10112]));
Q_ASSIGN U6279 ( .B(clk), .A(\g.we_clk [10111]));
Q_ASSIGN U6280 ( .B(clk), .A(\g.we_clk [10110]));
Q_ASSIGN U6281 ( .B(clk), .A(\g.we_clk [10109]));
Q_ASSIGN U6282 ( .B(clk), .A(\g.we_clk [10108]));
Q_ASSIGN U6283 ( .B(clk), .A(\g.we_clk [10107]));
Q_ASSIGN U6284 ( .B(clk), .A(\g.we_clk [10106]));
Q_ASSIGN U6285 ( .B(clk), .A(\g.we_clk [10105]));
Q_ASSIGN U6286 ( .B(clk), .A(\g.we_clk [10104]));
Q_ASSIGN U6287 ( .B(clk), .A(\g.we_clk [10103]));
Q_ASSIGN U6288 ( .B(clk), .A(\g.we_clk [10102]));
Q_ASSIGN U6289 ( .B(clk), .A(\g.we_clk [10101]));
Q_ASSIGN U6290 ( .B(clk), .A(\g.we_clk [10100]));
Q_ASSIGN U6291 ( .B(clk), .A(\g.we_clk [10099]));
Q_ASSIGN U6292 ( .B(clk), .A(\g.we_clk [10098]));
Q_ASSIGN U6293 ( .B(clk), .A(\g.we_clk [10097]));
Q_ASSIGN U6294 ( .B(clk), .A(\g.we_clk [10096]));
Q_ASSIGN U6295 ( .B(clk), .A(\g.we_clk [10095]));
Q_ASSIGN U6296 ( .B(clk), .A(\g.we_clk [10094]));
Q_ASSIGN U6297 ( .B(clk), .A(\g.we_clk [10093]));
Q_ASSIGN U6298 ( .B(clk), .A(\g.we_clk [10092]));
Q_ASSIGN U6299 ( .B(clk), .A(\g.we_clk [10091]));
Q_ASSIGN U6300 ( .B(clk), .A(\g.we_clk [10090]));
Q_ASSIGN U6301 ( .B(clk), .A(\g.we_clk [10089]));
Q_ASSIGN U6302 ( .B(clk), .A(\g.we_clk [10088]));
Q_ASSIGN U6303 ( .B(clk), .A(\g.we_clk [10087]));
Q_ASSIGN U6304 ( .B(clk), .A(\g.we_clk [10086]));
Q_ASSIGN U6305 ( .B(clk), .A(\g.we_clk [10085]));
Q_ASSIGN U6306 ( .B(clk), .A(\g.we_clk [10084]));
Q_ASSIGN U6307 ( .B(clk), .A(\g.we_clk [10083]));
Q_ASSIGN U6308 ( .B(clk), .A(\g.we_clk [10082]));
Q_ASSIGN U6309 ( .B(clk), .A(\g.we_clk [10081]));
Q_ASSIGN U6310 ( .B(clk), .A(\g.we_clk [10080]));
Q_ASSIGN U6311 ( .B(clk), .A(\g.we_clk [10079]));
Q_ASSIGN U6312 ( .B(clk), .A(\g.we_clk [10078]));
Q_ASSIGN U6313 ( .B(clk), .A(\g.we_clk [10077]));
Q_ASSIGN U6314 ( .B(clk), .A(\g.we_clk [10076]));
Q_ASSIGN U6315 ( .B(clk), .A(\g.we_clk [10075]));
Q_ASSIGN U6316 ( .B(clk), .A(\g.we_clk [10074]));
Q_ASSIGN U6317 ( .B(clk), .A(\g.we_clk [10073]));
Q_ASSIGN U6318 ( .B(clk), .A(\g.we_clk [10072]));
Q_ASSIGN U6319 ( .B(clk), .A(\g.we_clk [10071]));
Q_ASSIGN U6320 ( .B(clk), .A(\g.we_clk [10070]));
Q_ASSIGN U6321 ( .B(clk), .A(\g.we_clk [10069]));
Q_ASSIGN U6322 ( .B(clk), .A(\g.we_clk [10068]));
Q_ASSIGN U6323 ( .B(clk), .A(\g.we_clk [10067]));
Q_ASSIGN U6324 ( .B(clk), .A(\g.we_clk [10066]));
Q_ASSIGN U6325 ( .B(clk), .A(\g.we_clk [10065]));
Q_ASSIGN U6326 ( .B(clk), .A(\g.we_clk [10064]));
Q_ASSIGN U6327 ( .B(clk), .A(\g.we_clk [10063]));
Q_ASSIGN U6328 ( .B(clk), .A(\g.we_clk [10062]));
Q_ASSIGN U6329 ( .B(clk), .A(\g.we_clk [10061]));
Q_ASSIGN U6330 ( .B(clk), .A(\g.we_clk [10060]));
Q_ASSIGN U6331 ( .B(clk), .A(\g.we_clk [10059]));
Q_ASSIGN U6332 ( .B(clk), .A(\g.we_clk [10058]));
Q_ASSIGN U6333 ( .B(clk), .A(\g.we_clk [10057]));
Q_ASSIGN U6334 ( .B(clk), .A(\g.we_clk [10056]));
Q_ASSIGN U6335 ( .B(clk), .A(\g.we_clk [10055]));
Q_ASSIGN U6336 ( .B(clk), .A(\g.we_clk [10054]));
Q_ASSIGN U6337 ( .B(clk), .A(\g.we_clk [10053]));
Q_ASSIGN U6338 ( .B(clk), .A(\g.we_clk [10052]));
Q_ASSIGN U6339 ( .B(clk), .A(\g.we_clk [10051]));
Q_ASSIGN U6340 ( .B(clk), .A(\g.we_clk [10050]));
Q_ASSIGN U6341 ( .B(clk), .A(\g.we_clk [10049]));
Q_ASSIGN U6342 ( .B(clk), .A(\g.we_clk [10048]));
Q_ASSIGN U6343 ( .B(clk), .A(\g.we_clk [10047]));
Q_ASSIGN U6344 ( .B(clk), .A(\g.we_clk [10046]));
Q_ASSIGN U6345 ( .B(clk), .A(\g.we_clk [10045]));
Q_ASSIGN U6346 ( .B(clk), .A(\g.we_clk [10044]));
Q_ASSIGN U6347 ( .B(clk), .A(\g.we_clk [10043]));
Q_ASSIGN U6348 ( .B(clk), .A(\g.we_clk [10042]));
Q_ASSIGN U6349 ( .B(clk), .A(\g.we_clk [10041]));
Q_ASSIGN U6350 ( .B(clk), .A(\g.we_clk [10040]));
Q_ASSIGN U6351 ( .B(clk), .A(\g.we_clk [10039]));
Q_ASSIGN U6352 ( .B(clk), .A(\g.we_clk [10038]));
Q_ASSIGN U6353 ( .B(clk), .A(\g.we_clk [10037]));
Q_ASSIGN U6354 ( .B(clk), .A(\g.we_clk [10036]));
Q_ASSIGN U6355 ( .B(clk), .A(\g.we_clk [10035]));
Q_ASSIGN U6356 ( .B(clk), .A(\g.we_clk [10034]));
Q_ASSIGN U6357 ( .B(clk), .A(\g.we_clk [10033]));
Q_ASSIGN U6358 ( .B(clk), .A(\g.we_clk [10032]));
Q_ASSIGN U6359 ( .B(clk), .A(\g.we_clk [10031]));
Q_ASSIGN U6360 ( .B(clk), .A(\g.we_clk [10030]));
Q_ASSIGN U6361 ( .B(clk), .A(\g.we_clk [10029]));
Q_ASSIGN U6362 ( .B(clk), .A(\g.we_clk [10028]));
Q_ASSIGN U6363 ( .B(clk), .A(\g.we_clk [10027]));
Q_ASSIGN U6364 ( .B(clk), .A(\g.we_clk [10026]));
Q_ASSIGN U6365 ( .B(clk), .A(\g.we_clk [10025]));
Q_ASSIGN U6366 ( .B(clk), .A(\g.we_clk [10024]));
Q_ASSIGN U6367 ( .B(clk), .A(\g.we_clk [10023]));
Q_ASSIGN U6368 ( .B(clk), .A(\g.we_clk [10022]));
Q_ASSIGN U6369 ( .B(clk), .A(\g.we_clk [10021]));
Q_ASSIGN U6370 ( .B(clk), .A(\g.we_clk [10020]));
Q_ASSIGN U6371 ( .B(clk), .A(\g.we_clk [10019]));
Q_ASSIGN U6372 ( .B(clk), .A(\g.we_clk [10018]));
Q_ASSIGN U6373 ( .B(clk), .A(\g.we_clk [10017]));
Q_ASSIGN U6374 ( .B(clk), .A(\g.we_clk [10016]));
Q_ASSIGN U6375 ( .B(clk), .A(\g.we_clk [10015]));
Q_ASSIGN U6376 ( .B(clk), .A(\g.we_clk [10014]));
Q_ASSIGN U6377 ( .B(clk), .A(\g.we_clk [10013]));
Q_ASSIGN U6378 ( .B(clk), .A(\g.we_clk [10012]));
Q_ASSIGN U6379 ( .B(clk), .A(\g.we_clk [10011]));
Q_ASSIGN U6380 ( .B(clk), .A(\g.we_clk [10010]));
Q_ASSIGN U6381 ( .B(clk), .A(\g.we_clk [10009]));
Q_ASSIGN U6382 ( .B(clk), .A(\g.we_clk [10008]));
Q_ASSIGN U6383 ( .B(clk), .A(\g.we_clk [10007]));
Q_ASSIGN U6384 ( .B(clk), .A(\g.we_clk [10006]));
Q_ASSIGN U6385 ( .B(clk), .A(\g.we_clk [10005]));
Q_ASSIGN U6386 ( .B(clk), .A(\g.we_clk [10004]));
Q_ASSIGN U6387 ( .B(clk), .A(\g.we_clk [10003]));
Q_ASSIGN U6388 ( .B(clk), .A(\g.we_clk [10002]));
Q_ASSIGN U6389 ( .B(clk), .A(\g.we_clk [10001]));
Q_ASSIGN U6390 ( .B(clk), .A(\g.we_clk [10000]));
Q_ASSIGN U6391 ( .B(clk), .A(\g.we_clk [9999]));
Q_ASSIGN U6392 ( .B(clk), .A(\g.we_clk [9998]));
Q_ASSIGN U6393 ( .B(clk), .A(\g.we_clk [9997]));
Q_ASSIGN U6394 ( .B(clk), .A(\g.we_clk [9996]));
Q_ASSIGN U6395 ( .B(clk), .A(\g.we_clk [9995]));
Q_ASSIGN U6396 ( .B(clk), .A(\g.we_clk [9994]));
Q_ASSIGN U6397 ( .B(clk), .A(\g.we_clk [9993]));
Q_ASSIGN U6398 ( .B(clk), .A(\g.we_clk [9992]));
Q_ASSIGN U6399 ( .B(clk), .A(\g.we_clk [9991]));
Q_ASSIGN U6400 ( .B(clk), .A(\g.we_clk [9990]));
Q_ASSIGN U6401 ( .B(clk), .A(\g.we_clk [9989]));
Q_ASSIGN U6402 ( .B(clk), .A(\g.we_clk [9988]));
Q_ASSIGN U6403 ( .B(clk), .A(\g.we_clk [9987]));
Q_ASSIGN U6404 ( .B(clk), .A(\g.we_clk [9986]));
Q_ASSIGN U6405 ( .B(clk), .A(\g.we_clk [9985]));
Q_ASSIGN U6406 ( .B(clk), .A(\g.we_clk [9984]));
Q_ASSIGN U6407 ( .B(clk), .A(\g.we_clk [9983]));
Q_ASSIGN U6408 ( .B(clk), .A(\g.we_clk [9982]));
Q_ASSIGN U6409 ( .B(clk), .A(\g.we_clk [9981]));
Q_ASSIGN U6410 ( .B(clk), .A(\g.we_clk [9980]));
Q_ASSIGN U6411 ( .B(clk), .A(\g.we_clk [9979]));
Q_ASSIGN U6412 ( .B(clk), .A(\g.we_clk [9978]));
Q_ASSIGN U6413 ( .B(clk), .A(\g.we_clk [9977]));
Q_ASSIGN U6414 ( .B(clk), .A(\g.we_clk [9976]));
Q_ASSIGN U6415 ( .B(clk), .A(\g.we_clk [9975]));
Q_ASSIGN U6416 ( .B(clk), .A(\g.we_clk [9974]));
Q_ASSIGN U6417 ( .B(clk), .A(\g.we_clk [9973]));
Q_ASSIGN U6418 ( .B(clk), .A(\g.we_clk [9972]));
Q_ASSIGN U6419 ( .B(clk), .A(\g.we_clk [9971]));
Q_ASSIGN U6420 ( .B(clk), .A(\g.we_clk [9970]));
Q_ASSIGN U6421 ( .B(clk), .A(\g.we_clk [9969]));
Q_ASSIGN U6422 ( .B(clk), .A(\g.we_clk [9968]));
Q_ASSIGN U6423 ( .B(clk), .A(\g.we_clk [9967]));
Q_ASSIGN U6424 ( .B(clk), .A(\g.we_clk [9966]));
Q_ASSIGN U6425 ( .B(clk), .A(\g.we_clk [9965]));
Q_ASSIGN U6426 ( .B(clk), .A(\g.we_clk [9964]));
Q_ASSIGN U6427 ( .B(clk), .A(\g.we_clk [9963]));
Q_ASSIGN U6428 ( .B(clk), .A(\g.we_clk [9962]));
Q_ASSIGN U6429 ( .B(clk), .A(\g.we_clk [9961]));
Q_ASSIGN U6430 ( .B(clk), .A(\g.we_clk [9960]));
Q_ASSIGN U6431 ( .B(clk), .A(\g.we_clk [9959]));
Q_ASSIGN U6432 ( .B(clk), .A(\g.we_clk [9958]));
Q_ASSIGN U6433 ( .B(clk), .A(\g.we_clk [9957]));
Q_ASSIGN U6434 ( .B(clk), .A(\g.we_clk [9956]));
Q_ASSIGN U6435 ( .B(clk), .A(\g.we_clk [9955]));
Q_ASSIGN U6436 ( .B(clk), .A(\g.we_clk [9954]));
Q_ASSIGN U6437 ( .B(clk), .A(\g.we_clk [9953]));
Q_ASSIGN U6438 ( .B(clk), .A(\g.we_clk [9952]));
Q_ASSIGN U6439 ( .B(clk), .A(\g.we_clk [9951]));
Q_ASSIGN U6440 ( .B(clk), .A(\g.we_clk [9950]));
Q_ASSIGN U6441 ( .B(clk), .A(\g.we_clk [9949]));
Q_ASSIGN U6442 ( .B(clk), .A(\g.we_clk [9948]));
Q_ASSIGN U6443 ( .B(clk), .A(\g.we_clk [9947]));
Q_ASSIGN U6444 ( .B(clk), .A(\g.we_clk [9946]));
Q_ASSIGN U6445 ( .B(clk), .A(\g.we_clk [9945]));
Q_ASSIGN U6446 ( .B(clk), .A(\g.we_clk [9944]));
Q_ASSIGN U6447 ( .B(clk), .A(\g.we_clk [9943]));
Q_ASSIGN U6448 ( .B(clk), .A(\g.we_clk [9942]));
Q_ASSIGN U6449 ( .B(clk), .A(\g.we_clk [9941]));
Q_ASSIGN U6450 ( .B(clk), .A(\g.we_clk [9940]));
Q_ASSIGN U6451 ( .B(clk), .A(\g.we_clk [9939]));
Q_ASSIGN U6452 ( .B(clk), .A(\g.we_clk [9938]));
Q_ASSIGN U6453 ( .B(clk), .A(\g.we_clk [9937]));
Q_ASSIGN U6454 ( .B(clk), .A(\g.we_clk [9936]));
Q_ASSIGN U6455 ( .B(clk), .A(\g.we_clk [9935]));
Q_ASSIGN U6456 ( .B(clk), .A(\g.we_clk [9934]));
Q_ASSIGN U6457 ( .B(clk), .A(\g.we_clk [9933]));
Q_ASSIGN U6458 ( .B(clk), .A(\g.we_clk [9932]));
Q_ASSIGN U6459 ( .B(clk), .A(\g.we_clk [9931]));
Q_ASSIGN U6460 ( .B(clk), .A(\g.we_clk [9930]));
Q_ASSIGN U6461 ( .B(clk), .A(\g.we_clk [9929]));
Q_ASSIGN U6462 ( .B(clk), .A(\g.we_clk [9928]));
Q_ASSIGN U6463 ( .B(clk), .A(\g.we_clk [9927]));
Q_ASSIGN U6464 ( .B(clk), .A(\g.we_clk [9926]));
Q_ASSIGN U6465 ( .B(clk), .A(\g.we_clk [9925]));
Q_ASSIGN U6466 ( .B(clk), .A(\g.we_clk [9924]));
Q_ASSIGN U6467 ( .B(clk), .A(\g.we_clk [9923]));
Q_ASSIGN U6468 ( .B(clk), .A(\g.we_clk [9922]));
Q_ASSIGN U6469 ( .B(clk), .A(\g.we_clk [9921]));
Q_ASSIGN U6470 ( .B(clk), .A(\g.we_clk [9920]));
Q_ASSIGN U6471 ( .B(clk), .A(\g.we_clk [9919]));
Q_ASSIGN U6472 ( .B(clk), .A(\g.we_clk [9918]));
Q_ASSIGN U6473 ( .B(clk), .A(\g.we_clk [9917]));
Q_ASSIGN U6474 ( .B(clk), .A(\g.we_clk [9916]));
Q_ASSIGN U6475 ( .B(clk), .A(\g.we_clk [9915]));
Q_ASSIGN U6476 ( .B(clk), .A(\g.we_clk [9914]));
Q_ASSIGN U6477 ( .B(clk), .A(\g.we_clk [9913]));
Q_ASSIGN U6478 ( .B(clk), .A(\g.we_clk [9912]));
Q_ASSIGN U6479 ( .B(clk), .A(\g.we_clk [9911]));
Q_ASSIGN U6480 ( .B(clk), .A(\g.we_clk [9910]));
Q_ASSIGN U6481 ( .B(clk), .A(\g.we_clk [9909]));
Q_ASSIGN U6482 ( .B(clk), .A(\g.we_clk [9908]));
Q_ASSIGN U6483 ( .B(clk), .A(\g.we_clk [9907]));
Q_ASSIGN U6484 ( .B(clk), .A(\g.we_clk [9906]));
Q_ASSIGN U6485 ( .B(clk), .A(\g.we_clk [9905]));
Q_ASSIGN U6486 ( .B(clk), .A(\g.we_clk [9904]));
Q_ASSIGN U6487 ( .B(clk), .A(\g.we_clk [9903]));
Q_ASSIGN U6488 ( .B(clk), .A(\g.we_clk [9902]));
Q_ASSIGN U6489 ( .B(clk), .A(\g.we_clk [9901]));
Q_ASSIGN U6490 ( .B(clk), .A(\g.we_clk [9900]));
Q_ASSIGN U6491 ( .B(clk), .A(\g.we_clk [9899]));
Q_ASSIGN U6492 ( .B(clk), .A(\g.we_clk [9898]));
Q_ASSIGN U6493 ( .B(clk), .A(\g.we_clk [9897]));
Q_ASSIGN U6494 ( .B(clk), .A(\g.we_clk [9896]));
Q_ASSIGN U6495 ( .B(clk), .A(\g.we_clk [9895]));
Q_ASSIGN U6496 ( .B(clk), .A(\g.we_clk [9894]));
Q_ASSIGN U6497 ( .B(clk), .A(\g.we_clk [9893]));
Q_ASSIGN U6498 ( .B(clk), .A(\g.we_clk [9892]));
Q_ASSIGN U6499 ( .B(clk), .A(\g.we_clk [9891]));
Q_ASSIGN U6500 ( .B(clk), .A(\g.we_clk [9890]));
Q_ASSIGN U6501 ( .B(clk), .A(\g.we_clk [9889]));
Q_ASSIGN U6502 ( .B(clk), .A(\g.we_clk [9888]));
Q_ASSIGN U6503 ( .B(clk), .A(\g.we_clk [9887]));
Q_ASSIGN U6504 ( .B(clk), .A(\g.we_clk [9886]));
Q_ASSIGN U6505 ( .B(clk), .A(\g.we_clk [9885]));
Q_ASSIGN U6506 ( .B(clk), .A(\g.we_clk [9884]));
Q_ASSIGN U6507 ( .B(clk), .A(\g.we_clk [9883]));
Q_ASSIGN U6508 ( .B(clk), .A(\g.we_clk [9882]));
Q_ASSIGN U6509 ( .B(clk), .A(\g.we_clk [9881]));
Q_ASSIGN U6510 ( .B(clk), .A(\g.we_clk [9880]));
Q_ASSIGN U6511 ( .B(clk), .A(\g.we_clk [9879]));
Q_ASSIGN U6512 ( .B(clk), .A(\g.we_clk [9878]));
Q_ASSIGN U6513 ( .B(clk), .A(\g.we_clk [9877]));
Q_ASSIGN U6514 ( .B(clk), .A(\g.we_clk [9876]));
Q_ASSIGN U6515 ( .B(clk), .A(\g.we_clk [9875]));
Q_ASSIGN U6516 ( .B(clk), .A(\g.we_clk [9874]));
Q_ASSIGN U6517 ( .B(clk), .A(\g.we_clk [9873]));
Q_ASSIGN U6518 ( .B(clk), .A(\g.we_clk [9872]));
Q_ASSIGN U6519 ( .B(clk), .A(\g.we_clk [9871]));
Q_ASSIGN U6520 ( .B(clk), .A(\g.we_clk [9870]));
Q_ASSIGN U6521 ( .B(clk), .A(\g.we_clk [9869]));
Q_ASSIGN U6522 ( .B(clk), .A(\g.we_clk [9868]));
Q_ASSIGN U6523 ( .B(clk), .A(\g.we_clk [9867]));
Q_ASSIGN U6524 ( .B(clk), .A(\g.we_clk [9866]));
Q_ASSIGN U6525 ( .B(clk), .A(\g.we_clk [9865]));
Q_ASSIGN U6526 ( .B(clk), .A(\g.we_clk [9864]));
Q_ASSIGN U6527 ( .B(clk), .A(\g.we_clk [9863]));
Q_ASSIGN U6528 ( .B(clk), .A(\g.we_clk [9862]));
Q_ASSIGN U6529 ( .B(clk), .A(\g.we_clk [9861]));
Q_ASSIGN U6530 ( .B(clk), .A(\g.we_clk [9860]));
Q_ASSIGN U6531 ( .B(clk), .A(\g.we_clk [9859]));
Q_ASSIGN U6532 ( .B(clk), .A(\g.we_clk [9858]));
Q_ASSIGN U6533 ( .B(clk), .A(\g.we_clk [9857]));
Q_ASSIGN U6534 ( .B(clk), .A(\g.we_clk [9856]));
Q_ASSIGN U6535 ( .B(clk), .A(\g.we_clk [9855]));
Q_ASSIGN U6536 ( .B(clk), .A(\g.we_clk [9854]));
Q_ASSIGN U6537 ( .B(clk), .A(\g.we_clk [9853]));
Q_ASSIGN U6538 ( .B(clk), .A(\g.we_clk [9852]));
Q_ASSIGN U6539 ( .B(clk), .A(\g.we_clk [9851]));
Q_ASSIGN U6540 ( .B(clk), .A(\g.we_clk [9850]));
Q_ASSIGN U6541 ( .B(clk), .A(\g.we_clk [9849]));
Q_ASSIGN U6542 ( .B(clk), .A(\g.we_clk [9848]));
Q_ASSIGN U6543 ( .B(clk), .A(\g.we_clk [9847]));
Q_ASSIGN U6544 ( .B(clk), .A(\g.we_clk [9846]));
Q_ASSIGN U6545 ( .B(clk), .A(\g.we_clk [9845]));
Q_ASSIGN U6546 ( .B(clk), .A(\g.we_clk [9844]));
Q_ASSIGN U6547 ( .B(clk), .A(\g.we_clk [9843]));
Q_ASSIGN U6548 ( .B(clk), .A(\g.we_clk [9842]));
Q_ASSIGN U6549 ( .B(clk), .A(\g.we_clk [9841]));
Q_ASSIGN U6550 ( .B(clk), .A(\g.we_clk [9840]));
Q_ASSIGN U6551 ( .B(clk), .A(\g.we_clk [9839]));
Q_ASSIGN U6552 ( .B(clk), .A(\g.we_clk [9838]));
Q_ASSIGN U6553 ( .B(clk), .A(\g.we_clk [9837]));
Q_ASSIGN U6554 ( .B(clk), .A(\g.we_clk [9836]));
Q_ASSIGN U6555 ( .B(clk), .A(\g.we_clk [9835]));
Q_ASSIGN U6556 ( .B(clk), .A(\g.we_clk [9834]));
Q_ASSIGN U6557 ( .B(clk), .A(\g.we_clk [9833]));
Q_ASSIGN U6558 ( .B(clk), .A(\g.we_clk [9832]));
Q_ASSIGN U6559 ( .B(clk), .A(\g.we_clk [9831]));
Q_ASSIGN U6560 ( .B(clk), .A(\g.we_clk [9830]));
Q_ASSIGN U6561 ( .B(clk), .A(\g.we_clk [9829]));
Q_ASSIGN U6562 ( .B(clk), .A(\g.we_clk [9828]));
Q_ASSIGN U6563 ( .B(clk), .A(\g.we_clk [9827]));
Q_ASSIGN U6564 ( .B(clk), .A(\g.we_clk [9826]));
Q_ASSIGN U6565 ( .B(clk), .A(\g.we_clk [9825]));
Q_ASSIGN U6566 ( .B(clk), .A(\g.we_clk [9824]));
Q_ASSIGN U6567 ( .B(clk), .A(\g.we_clk [9823]));
Q_ASSIGN U6568 ( .B(clk), .A(\g.we_clk [9822]));
Q_ASSIGN U6569 ( .B(clk), .A(\g.we_clk [9821]));
Q_ASSIGN U6570 ( .B(clk), .A(\g.we_clk [9820]));
Q_ASSIGN U6571 ( .B(clk), .A(\g.we_clk [9819]));
Q_ASSIGN U6572 ( .B(clk), .A(\g.we_clk [9818]));
Q_ASSIGN U6573 ( .B(clk), .A(\g.we_clk [9817]));
Q_ASSIGN U6574 ( .B(clk), .A(\g.we_clk [9816]));
Q_ASSIGN U6575 ( .B(clk), .A(\g.we_clk [9815]));
Q_ASSIGN U6576 ( .B(clk), .A(\g.we_clk [9814]));
Q_ASSIGN U6577 ( .B(clk), .A(\g.we_clk [9813]));
Q_ASSIGN U6578 ( .B(clk), .A(\g.we_clk [9812]));
Q_ASSIGN U6579 ( .B(clk), .A(\g.we_clk [9811]));
Q_ASSIGN U6580 ( .B(clk), .A(\g.we_clk [9810]));
Q_ASSIGN U6581 ( .B(clk), .A(\g.we_clk [9809]));
Q_ASSIGN U6582 ( .B(clk), .A(\g.we_clk [9808]));
Q_ASSIGN U6583 ( .B(clk), .A(\g.we_clk [9807]));
Q_ASSIGN U6584 ( .B(clk), .A(\g.we_clk [9806]));
Q_ASSIGN U6585 ( .B(clk), .A(\g.we_clk [9805]));
Q_ASSIGN U6586 ( .B(clk), .A(\g.we_clk [9804]));
Q_ASSIGN U6587 ( .B(clk), .A(\g.we_clk [9803]));
Q_ASSIGN U6588 ( .B(clk), .A(\g.we_clk [9802]));
Q_ASSIGN U6589 ( .B(clk), .A(\g.we_clk [9801]));
Q_ASSIGN U6590 ( .B(clk), .A(\g.we_clk [9800]));
Q_ASSIGN U6591 ( .B(clk), .A(\g.we_clk [9799]));
Q_ASSIGN U6592 ( .B(clk), .A(\g.we_clk [9798]));
Q_ASSIGN U6593 ( .B(clk), .A(\g.we_clk [9797]));
Q_ASSIGN U6594 ( .B(clk), .A(\g.we_clk [9796]));
Q_ASSIGN U6595 ( .B(clk), .A(\g.we_clk [9795]));
Q_ASSIGN U6596 ( .B(clk), .A(\g.we_clk [9794]));
Q_ASSIGN U6597 ( .B(clk), .A(\g.we_clk [9793]));
Q_ASSIGN U6598 ( .B(clk), .A(\g.we_clk [9792]));
Q_ASSIGN U6599 ( .B(clk), .A(\g.we_clk [9791]));
Q_ASSIGN U6600 ( .B(clk), .A(\g.we_clk [9790]));
Q_ASSIGN U6601 ( .B(clk), .A(\g.we_clk [9789]));
Q_ASSIGN U6602 ( .B(clk), .A(\g.we_clk [9788]));
Q_ASSIGN U6603 ( .B(clk), .A(\g.we_clk [9787]));
Q_ASSIGN U6604 ( .B(clk), .A(\g.we_clk [9786]));
Q_ASSIGN U6605 ( .B(clk), .A(\g.we_clk [9785]));
Q_ASSIGN U6606 ( .B(clk), .A(\g.we_clk [9784]));
Q_ASSIGN U6607 ( .B(clk), .A(\g.we_clk [9783]));
Q_ASSIGN U6608 ( .B(clk), .A(\g.we_clk [9782]));
Q_ASSIGN U6609 ( .B(clk), .A(\g.we_clk [9781]));
Q_ASSIGN U6610 ( .B(clk), .A(\g.we_clk [9780]));
Q_ASSIGN U6611 ( .B(clk), .A(\g.we_clk [9779]));
Q_ASSIGN U6612 ( .B(clk), .A(\g.we_clk [9778]));
Q_ASSIGN U6613 ( .B(clk), .A(\g.we_clk [9777]));
Q_ASSIGN U6614 ( .B(clk), .A(\g.we_clk [9776]));
Q_ASSIGN U6615 ( .B(clk), .A(\g.we_clk [9775]));
Q_ASSIGN U6616 ( .B(clk), .A(\g.we_clk [9774]));
Q_ASSIGN U6617 ( .B(clk), .A(\g.we_clk [9773]));
Q_ASSIGN U6618 ( .B(clk), .A(\g.we_clk [9772]));
Q_ASSIGN U6619 ( .B(clk), .A(\g.we_clk [9771]));
Q_ASSIGN U6620 ( .B(clk), .A(\g.we_clk [9770]));
Q_ASSIGN U6621 ( .B(clk), .A(\g.we_clk [9769]));
Q_ASSIGN U6622 ( .B(clk), .A(\g.we_clk [9768]));
Q_ASSIGN U6623 ( .B(clk), .A(\g.we_clk [9767]));
Q_ASSIGN U6624 ( .B(clk), .A(\g.we_clk [9766]));
Q_ASSIGN U6625 ( .B(clk), .A(\g.we_clk [9765]));
Q_ASSIGN U6626 ( .B(clk), .A(\g.we_clk [9764]));
Q_ASSIGN U6627 ( .B(clk), .A(\g.we_clk [9763]));
Q_ASSIGN U6628 ( .B(clk), .A(\g.we_clk [9762]));
Q_ASSIGN U6629 ( .B(clk), .A(\g.we_clk [9761]));
Q_ASSIGN U6630 ( .B(clk), .A(\g.we_clk [9760]));
Q_ASSIGN U6631 ( .B(clk), .A(\g.we_clk [9759]));
Q_ASSIGN U6632 ( .B(clk), .A(\g.we_clk [9758]));
Q_ASSIGN U6633 ( .B(clk), .A(\g.we_clk [9757]));
Q_ASSIGN U6634 ( .B(clk), .A(\g.we_clk [9756]));
Q_ASSIGN U6635 ( .B(clk), .A(\g.we_clk [9755]));
Q_ASSIGN U6636 ( .B(clk), .A(\g.we_clk [9754]));
Q_ASSIGN U6637 ( .B(clk), .A(\g.we_clk [9753]));
Q_ASSIGN U6638 ( .B(clk), .A(\g.we_clk [9752]));
Q_ASSIGN U6639 ( .B(clk), .A(\g.we_clk [9751]));
Q_ASSIGN U6640 ( .B(clk), .A(\g.we_clk [9750]));
Q_ASSIGN U6641 ( .B(clk), .A(\g.we_clk [9749]));
Q_ASSIGN U6642 ( .B(clk), .A(\g.we_clk [9748]));
Q_ASSIGN U6643 ( .B(clk), .A(\g.we_clk [9747]));
Q_ASSIGN U6644 ( .B(clk), .A(\g.we_clk [9746]));
Q_ASSIGN U6645 ( .B(clk), .A(\g.we_clk [9745]));
Q_ASSIGN U6646 ( .B(clk), .A(\g.we_clk [9744]));
Q_ASSIGN U6647 ( .B(clk), .A(\g.we_clk [9743]));
Q_ASSIGN U6648 ( .B(clk), .A(\g.we_clk [9742]));
Q_ASSIGN U6649 ( .B(clk), .A(\g.we_clk [9741]));
Q_ASSIGN U6650 ( .B(clk), .A(\g.we_clk [9740]));
Q_ASSIGN U6651 ( .B(clk), .A(\g.we_clk [9739]));
Q_ASSIGN U6652 ( .B(clk), .A(\g.we_clk [9738]));
Q_ASSIGN U6653 ( .B(clk), .A(\g.we_clk [9737]));
Q_ASSIGN U6654 ( .B(clk), .A(\g.we_clk [9736]));
Q_ASSIGN U6655 ( .B(clk), .A(\g.we_clk [9735]));
Q_ASSIGN U6656 ( .B(clk), .A(\g.we_clk [9734]));
Q_ASSIGN U6657 ( .B(clk), .A(\g.we_clk [9733]));
Q_ASSIGN U6658 ( .B(clk), .A(\g.we_clk [9732]));
Q_ASSIGN U6659 ( .B(clk), .A(\g.we_clk [9731]));
Q_ASSIGN U6660 ( .B(clk), .A(\g.we_clk [9730]));
Q_ASSIGN U6661 ( .B(clk), .A(\g.we_clk [9729]));
Q_ASSIGN U6662 ( .B(clk), .A(\g.we_clk [9728]));
Q_ASSIGN U6663 ( .B(clk), .A(\g.we_clk [9727]));
Q_ASSIGN U6664 ( .B(clk), .A(\g.we_clk [9726]));
Q_ASSIGN U6665 ( .B(clk), .A(\g.we_clk [9725]));
Q_ASSIGN U6666 ( .B(clk), .A(\g.we_clk [9724]));
Q_ASSIGN U6667 ( .B(clk), .A(\g.we_clk [9723]));
Q_ASSIGN U6668 ( .B(clk), .A(\g.we_clk [9722]));
Q_ASSIGN U6669 ( .B(clk), .A(\g.we_clk [9721]));
Q_ASSIGN U6670 ( .B(clk), .A(\g.we_clk [9720]));
Q_ASSIGN U6671 ( .B(clk), .A(\g.we_clk [9719]));
Q_ASSIGN U6672 ( .B(clk), .A(\g.we_clk [9718]));
Q_ASSIGN U6673 ( .B(clk), .A(\g.we_clk [9717]));
Q_ASSIGN U6674 ( .B(clk), .A(\g.we_clk [9716]));
Q_ASSIGN U6675 ( .B(clk), .A(\g.we_clk [9715]));
Q_ASSIGN U6676 ( .B(clk), .A(\g.we_clk [9714]));
Q_ASSIGN U6677 ( .B(clk), .A(\g.we_clk [9713]));
Q_ASSIGN U6678 ( .B(clk), .A(\g.we_clk [9712]));
Q_ASSIGN U6679 ( .B(clk), .A(\g.we_clk [9711]));
Q_ASSIGN U6680 ( .B(clk), .A(\g.we_clk [9710]));
Q_ASSIGN U6681 ( .B(clk), .A(\g.we_clk [9709]));
Q_ASSIGN U6682 ( .B(clk), .A(\g.we_clk [9708]));
Q_ASSIGN U6683 ( .B(clk), .A(\g.we_clk [9707]));
Q_ASSIGN U6684 ( .B(clk), .A(\g.we_clk [9706]));
Q_ASSIGN U6685 ( .B(clk), .A(\g.we_clk [9705]));
Q_ASSIGN U6686 ( .B(clk), .A(\g.we_clk [9704]));
Q_ASSIGN U6687 ( .B(clk), .A(\g.we_clk [9703]));
Q_ASSIGN U6688 ( .B(clk), .A(\g.we_clk [9702]));
Q_ASSIGN U6689 ( .B(clk), .A(\g.we_clk [9701]));
Q_ASSIGN U6690 ( .B(clk), .A(\g.we_clk [9700]));
Q_ASSIGN U6691 ( .B(clk), .A(\g.we_clk [9699]));
Q_ASSIGN U6692 ( .B(clk), .A(\g.we_clk [9698]));
Q_ASSIGN U6693 ( .B(clk), .A(\g.we_clk [9697]));
Q_ASSIGN U6694 ( .B(clk), .A(\g.we_clk [9696]));
Q_ASSIGN U6695 ( .B(clk), .A(\g.we_clk [9695]));
Q_ASSIGN U6696 ( .B(clk), .A(\g.we_clk [9694]));
Q_ASSIGN U6697 ( .B(clk), .A(\g.we_clk [9693]));
Q_ASSIGN U6698 ( .B(clk), .A(\g.we_clk [9692]));
Q_ASSIGN U6699 ( .B(clk), .A(\g.we_clk [9691]));
Q_ASSIGN U6700 ( .B(clk), .A(\g.we_clk [9690]));
Q_ASSIGN U6701 ( .B(clk), .A(\g.we_clk [9689]));
Q_ASSIGN U6702 ( .B(clk), .A(\g.we_clk [9688]));
Q_ASSIGN U6703 ( .B(clk), .A(\g.we_clk [9687]));
Q_ASSIGN U6704 ( .B(clk), .A(\g.we_clk [9686]));
Q_ASSIGN U6705 ( .B(clk), .A(\g.we_clk [9685]));
Q_ASSIGN U6706 ( .B(clk), .A(\g.we_clk [9684]));
Q_ASSIGN U6707 ( .B(clk), .A(\g.we_clk [9683]));
Q_ASSIGN U6708 ( .B(clk), .A(\g.we_clk [9682]));
Q_ASSIGN U6709 ( .B(clk), .A(\g.we_clk [9681]));
Q_ASSIGN U6710 ( .B(clk), .A(\g.we_clk [9680]));
Q_ASSIGN U6711 ( .B(clk), .A(\g.we_clk [9679]));
Q_ASSIGN U6712 ( .B(clk), .A(\g.we_clk [9678]));
Q_ASSIGN U6713 ( .B(clk), .A(\g.we_clk [9677]));
Q_ASSIGN U6714 ( .B(clk), .A(\g.we_clk [9676]));
Q_ASSIGN U6715 ( .B(clk), .A(\g.we_clk [9675]));
Q_ASSIGN U6716 ( .B(clk), .A(\g.we_clk [9674]));
Q_ASSIGN U6717 ( .B(clk), .A(\g.we_clk [9673]));
Q_ASSIGN U6718 ( .B(clk), .A(\g.we_clk [9672]));
Q_ASSIGN U6719 ( .B(clk), .A(\g.we_clk [9671]));
Q_ASSIGN U6720 ( .B(clk), .A(\g.we_clk [9670]));
Q_ASSIGN U6721 ( .B(clk), .A(\g.we_clk [9669]));
Q_ASSIGN U6722 ( .B(clk), .A(\g.we_clk [9668]));
Q_ASSIGN U6723 ( .B(clk), .A(\g.we_clk [9667]));
Q_ASSIGN U6724 ( .B(clk), .A(\g.we_clk [9666]));
Q_ASSIGN U6725 ( .B(clk), .A(\g.we_clk [9665]));
Q_ASSIGN U6726 ( .B(clk), .A(\g.we_clk [9664]));
Q_ASSIGN U6727 ( .B(clk), .A(\g.we_clk [9663]));
Q_ASSIGN U6728 ( .B(clk), .A(\g.we_clk [9662]));
Q_ASSIGN U6729 ( .B(clk), .A(\g.we_clk [9661]));
Q_ASSIGN U6730 ( .B(clk), .A(\g.we_clk [9660]));
Q_ASSIGN U6731 ( .B(clk), .A(\g.we_clk [9659]));
Q_ASSIGN U6732 ( .B(clk), .A(\g.we_clk [9658]));
Q_ASSIGN U6733 ( .B(clk), .A(\g.we_clk [9657]));
Q_ASSIGN U6734 ( .B(clk), .A(\g.we_clk [9656]));
Q_ASSIGN U6735 ( .B(clk), .A(\g.we_clk [9655]));
Q_ASSIGN U6736 ( .B(clk), .A(\g.we_clk [9654]));
Q_ASSIGN U6737 ( .B(clk), .A(\g.we_clk [9653]));
Q_ASSIGN U6738 ( .B(clk), .A(\g.we_clk [9652]));
Q_ASSIGN U6739 ( .B(clk), .A(\g.we_clk [9651]));
Q_ASSIGN U6740 ( .B(clk), .A(\g.we_clk [9650]));
Q_ASSIGN U6741 ( .B(clk), .A(\g.we_clk [9649]));
Q_ASSIGN U6742 ( .B(clk), .A(\g.we_clk [9648]));
Q_ASSIGN U6743 ( .B(clk), .A(\g.we_clk [9647]));
Q_ASSIGN U6744 ( .B(clk), .A(\g.we_clk [9646]));
Q_ASSIGN U6745 ( .B(clk), .A(\g.we_clk [9645]));
Q_ASSIGN U6746 ( .B(clk), .A(\g.we_clk [9644]));
Q_ASSIGN U6747 ( .B(clk), .A(\g.we_clk [9643]));
Q_ASSIGN U6748 ( .B(clk), .A(\g.we_clk [9642]));
Q_ASSIGN U6749 ( .B(clk), .A(\g.we_clk [9641]));
Q_ASSIGN U6750 ( .B(clk), .A(\g.we_clk [9640]));
Q_ASSIGN U6751 ( .B(clk), .A(\g.we_clk [9639]));
Q_ASSIGN U6752 ( .B(clk), .A(\g.we_clk [9638]));
Q_ASSIGN U6753 ( .B(clk), .A(\g.we_clk [9637]));
Q_ASSIGN U6754 ( .B(clk), .A(\g.we_clk [9636]));
Q_ASSIGN U6755 ( .B(clk), .A(\g.we_clk [9635]));
Q_ASSIGN U6756 ( .B(clk), .A(\g.we_clk [9634]));
Q_ASSIGN U6757 ( .B(clk), .A(\g.we_clk [9633]));
Q_ASSIGN U6758 ( .B(clk), .A(\g.we_clk [9632]));
Q_ASSIGN U6759 ( .B(clk), .A(\g.we_clk [9631]));
Q_ASSIGN U6760 ( .B(clk), .A(\g.we_clk [9630]));
Q_ASSIGN U6761 ( .B(clk), .A(\g.we_clk [9629]));
Q_ASSIGN U6762 ( .B(clk), .A(\g.we_clk [9628]));
Q_ASSIGN U6763 ( .B(clk), .A(\g.we_clk [9627]));
Q_ASSIGN U6764 ( .B(clk), .A(\g.we_clk [9626]));
Q_ASSIGN U6765 ( .B(clk), .A(\g.we_clk [9625]));
Q_ASSIGN U6766 ( .B(clk), .A(\g.we_clk [9624]));
Q_ASSIGN U6767 ( .B(clk), .A(\g.we_clk [9623]));
Q_ASSIGN U6768 ( .B(clk), .A(\g.we_clk [9622]));
Q_ASSIGN U6769 ( .B(clk), .A(\g.we_clk [9621]));
Q_ASSIGN U6770 ( .B(clk), .A(\g.we_clk [9620]));
Q_ASSIGN U6771 ( .B(clk), .A(\g.we_clk [9619]));
Q_ASSIGN U6772 ( .B(clk), .A(\g.we_clk [9618]));
Q_ASSIGN U6773 ( .B(clk), .A(\g.we_clk [9617]));
Q_ASSIGN U6774 ( .B(clk), .A(\g.we_clk [9616]));
Q_ASSIGN U6775 ( .B(clk), .A(\g.we_clk [9615]));
Q_ASSIGN U6776 ( .B(clk), .A(\g.we_clk [9614]));
Q_ASSIGN U6777 ( .B(clk), .A(\g.we_clk [9613]));
Q_ASSIGN U6778 ( .B(clk), .A(\g.we_clk [9612]));
Q_ASSIGN U6779 ( .B(clk), .A(\g.we_clk [9611]));
Q_ASSIGN U6780 ( .B(clk), .A(\g.we_clk [9610]));
Q_ASSIGN U6781 ( .B(clk), .A(\g.we_clk [9609]));
Q_ASSIGN U6782 ( .B(clk), .A(\g.we_clk [9608]));
Q_ASSIGN U6783 ( .B(clk), .A(\g.we_clk [9607]));
Q_ASSIGN U6784 ( .B(clk), .A(\g.we_clk [9606]));
Q_ASSIGN U6785 ( .B(clk), .A(\g.we_clk [9605]));
Q_ASSIGN U6786 ( .B(clk), .A(\g.we_clk [9604]));
Q_ASSIGN U6787 ( .B(clk), .A(\g.we_clk [9603]));
Q_ASSIGN U6788 ( .B(clk), .A(\g.we_clk [9602]));
Q_ASSIGN U6789 ( .B(clk), .A(\g.we_clk [9601]));
Q_ASSIGN U6790 ( .B(clk), .A(\g.we_clk [9600]));
Q_ASSIGN U6791 ( .B(clk), .A(\g.we_clk [9599]));
Q_ASSIGN U6792 ( .B(clk), .A(\g.we_clk [9598]));
Q_ASSIGN U6793 ( .B(clk), .A(\g.we_clk [9597]));
Q_ASSIGN U6794 ( .B(clk), .A(\g.we_clk [9596]));
Q_ASSIGN U6795 ( .B(clk), .A(\g.we_clk [9595]));
Q_ASSIGN U6796 ( .B(clk), .A(\g.we_clk [9594]));
Q_ASSIGN U6797 ( .B(clk), .A(\g.we_clk [9593]));
Q_ASSIGN U6798 ( .B(clk), .A(\g.we_clk [9592]));
Q_ASSIGN U6799 ( .B(clk), .A(\g.we_clk [9591]));
Q_ASSIGN U6800 ( .B(clk), .A(\g.we_clk [9590]));
Q_ASSIGN U6801 ( .B(clk), .A(\g.we_clk [9589]));
Q_ASSIGN U6802 ( .B(clk), .A(\g.we_clk [9588]));
Q_ASSIGN U6803 ( .B(clk), .A(\g.we_clk [9587]));
Q_ASSIGN U6804 ( .B(clk), .A(\g.we_clk [9586]));
Q_ASSIGN U6805 ( .B(clk), .A(\g.we_clk [9585]));
Q_ASSIGN U6806 ( .B(clk), .A(\g.we_clk [9584]));
Q_ASSIGN U6807 ( .B(clk), .A(\g.we_clk [9583]));
Q_ASSIGN U6808 ( .B(clk), .A(\g.we_clk [9582]));
Q_ASSIGN U6809 ( .B(clk), .A(\g.we_clk [9581]));
Q_ASSIGN U6810 ( .B(clk), .A(\g.we_clk [9580]));
Q_ASSIGN U6811 ( .B(clk), .A(\g.we_clk [9579]));
Q_ASSIGN U6812 ( .B(clk), .A(\g.we_clk [9578]));
Q_ASSIGN U6813 ( .B(clk), .A(\g.we_clk [9577]));
Q_ASSIGN U6814 ( .B(clk), .A(\g.we_clk [9576]));
Q_ASSIGN U6815 ( .B(clk), .A(\g.we_clk [9575]));
Q_ASSIGN U6816 ( .B(clk), .A(\g.we_clk [9574]));
Q_ASSIGN U6817 ( .B(clk), .A(\g.we_clk [9573]));
Q_ASSIGN U6818 ( .B(clk), .A(\g.we_clk [9572]));
Q_ASSIGN U6819 ( .B(clk), .A(\g.we_clk [9571]));
Q_ASSIGN U6820 ( .B(clk), .A(\g.we_clk [9570]));
Q_ASSIGN U6821 ( .B(clk), .A(\g.we_clk [9569]));
Q_ASSIGN U6822 ( .B(clk), .A(\g.we_clk [9568]));
Q_ASSIGN U6823 ( .B(clk), .A(\g.we_clk [9567]));
Q_ASSIGN U6824 ( .B(clk), .A(\g.we_clk [9566]));
Q_ASSIGN U6825 ( .B(clk), .A(\g.we_clk [9565]));
Q_ASSIGN U6826 ( .B(clk), .A(\g.we_clk [9564]));
Q_ASSIGN U6827 ( .B(clk), .A(\g.we_clk [9563]));
Q_ASSIGN U6828 ( .B(clk), .A(\g.we_clk [9562]));
Q_ASSIGN U6829 ( .B(clk), .A(\g.we_clk [9561]));
Q_ASSIGN U6830 ( .B(clk), .A(\g.we_clk [9560]));
Q_ASSIGN U6831 ( .B(clk), .A(\g.we_clk [9559]));
Q_ASSIGN U6832 ( .B(clk), .A(\g.we_clk [9558]));
Q_ASSIGN U6833 ( .B(clk), .A(\g.we_clk [9557]));
Q_ASSIGN U6834 ( .B(clk), .A(\g.we_clk [9556]));
Q_ASSIGN U6835 ( .B(clk), .A(\g.we_clk [9555]));
Q_ASSIGN U6836 ( .B(clk), .A(\g.we_clk [9554]));
Q_ASSIGN U6837 ( .B(clk), .A(\g.we_clk [9553]));
Q_ASSIGN U6838 ( .B(clk), .A(\g.we_clk [9552]));
Q_ASSIGN U6839 ( .B(clk), .A(\g.we_clk [9551]));
Q_ASSIGN U6840 ( .B(clk), .A(\g.we_clk [9550]));
Q_ASSIGN U6841 ( .B(clk), .A(\g.we_clk [9549]));
Q_ASSIGN U6842 ( .B(clk), .A(\g.we_clk [9548]));
Q_ASSIGN U6843 ( .B(clk), .A(\g.we_clk [9547]));
Q_ASSIGN U6844 ( .B(clk), .A(\g.we_clk [9546]));
Q_ASSIGN U6845 ( .B(clk), .A(\g.we_clk [9545]));
Q_ASSIGN U6846 ( .B(clk), .A(\g.we_clk [9544]));
Q_ASSIGN U6847 ( .B(clk), .A(\g.we_clk [9543]));
Q_ASSIGN U6848 ( .B(clk), .A(\g.we_clk [9542]));
Q_ASSIGN U6849 ( .B(clk), .A(\g.we_clk [9541]));
Q_ASSIGN U6850 ( .B(clk), .A(\g.we_clk [9540]));
Q_ASSIGN U6851 ( .B(clk), .A(\g.we_clk [9539]));
Q_ASSIGN U6852 ( .B(clk), .A(\g.we_clk [9538]));
Q_ASSIGN U6853 ( .B(clk), .A(\g.we_clk [9537]));
Q_ASSIGN U6854 ( .B(clk), .A(\g.we_clk [9536]));
Q_ASSIGN U6855 ( .B(clk), .A(\g.we_clk [9535]));
Q_ASSIGN U6856 ( .B(clk), .A(\g.we_clk [9534]));
Q_ASSIGN U6857 ( .B(clk), .A(\g.we_clk [9533]));
Q_ASSIGN U6858 ( .B(clk), .A(\g.we_clk [9532]));
Q_ASSIGN U6859 ( .B(clk), .A(\g.we_clk [9531]));
Q_ASSIGN U6860 ( .B(clk), .A(\g.we_clk [9530]));
Q_ASSIGN U6861 ( .B(clk), .A(\g.we_clk [9529]));
Q_ASSIGN U6862 ( .B(clk), .A(\g.we_clk [9528]));
Q_ASSIGN U6863 ( .B(clk), .A(\g.we_clk [9527]));
Q_ASSIGN U6864 ( .B(clk), .A(\g.we_clk [9526]));
Q_ASSIGN U6865 ( .B(clk), .A(\g.we_clk [9525]));
Q_ASSIGN U6866 ( .B(clk), .A(\g.we_clk [9524]));
Q_ASSIGN U6867 ( .B(clk), .A(\g.we_clk [9523]));
Q_ASSIGN U6868 ( .B(clk), .A(\g.we_clk [9522]));
Q_ASSIGN U6869 ( .B(clk), .A(\g.we_clk [9521]));
Q_ASSIGN U6870 ( .B(clk), .A(\g.we_clk [9520]));
Q_ASSIGN U6871 ( .B(clk), .A(\g.we_clk [9519]));
Q_ASSIGN U6872 ( .B(clk), .A(\g.we_clk [9518]));
Q_ASSIGN U6873 ( .B(clk), .A(\g.we_clk [9517]));
Q_ASSIGN U6874 ( .B(clk), .A(\g.we_clk [9516]));
Q_ASSIGN U6875 ( .B(clk), .A(\g.we_clk [9515]));
Q_ASSIGN U6876 ( .B(clk), .A(\g.we_clk [9514]));
Q_ASSIGN U6877 ( .B(clk), .A(\g.we_clk [9513]));
Q_ASSIGN U6878 ( .B(clk), .A(\g.we_clk [9512]));
Q_ASSIGN U6879 ( .B(clk), .A(\g.we_clk [9511]));
Q_ASSIGN U6880 ( .B(clk), .A(\g.we_clk [9510]));
Q_ASSIGN U6881 ( .B(clk), .A(\g.we_clk [9509]));
Q_ASSIGN U6882 ( .B(clk), .A(\g.we_clk [9508]));
Q_ASSIGN U6883 ( .B(clk), .A(\g.we_clk [9507]));
Q_ASSIGN U6884 ( .B(clk), .A(\g.we_clk [9506]));
Q_ASSIGN U6885 ( .B(clk), .A(\g.we_clk [9505]));
Q_ASSIGN U6886 ( .B(clk), .A(\g.we_clk [9504]));
Q_ASSIGN U6887 ( .B(clk), .A(\g.we_clk [9503]));
Q_ASSIGN U6888 ( .B(clk), .A(\g.we_clk [9502]));
Q_ASSIGN U6889 ( .B(clk), .A(\g.we_clk [9501]));
Q_ASSIGN U6890 ( .B(clk), .A(\g.we_clk [9500]));
Q_ASSIGN U6891 ( .B(clk), .A(\g.we_clk [9499]));
Q_ASSIGN U6892 ( .B(clk), .A(\g.we_clk [9498]));
Q_ASSIGN U6893 ( .B(clk), .A(\g.we_clk [9497]));
Q_ASSIGN U6894 ( .B(clk), .A(\g.we_clk [9496]));
Q_ASSIGN U6895 ( .B(clk), .A(\g.we_clk [9495]));
Q_ASSIGN U6896 ( .B(clk), .A(\g.we_clk [9494]));
Q_ASSIGN U6897 ( .B(clk), .A(\g.we_clk [9493]));
Q_ASSIGN U6898 ( .B(clk), .A(\g.we_clk [9492]));
Q_ASSIGN U6899 ( .B(clk), .A(\g.we_clk [9491]));
Q_ASSIGN U6900 ( .B(clk), .A(\g.we_clk [9490]));
Q_ASSIGN U6901 ( .B(clk), .A(\g.we_clk [9489]));
Q_ASSIGN U6902 ( .B(clk), .A(\g.we_clk [9488]));
Q_ASSIGN U6903 ( .B(clk), .A(\g.we_clk [9487]));
Q_ASSIGN U6904 ( .B(clk), .A(\g.we_clk [9486]));
Q_ASSIGN U6905 ( .B(clk), .A(\g.we_clk [9485]));
Q_ASSIGN U6906 ( .B(clk), .A(\g.we_clk [9484]));
Q_ASSIGN U6907 ( .B(clk), .A(\g.we_clk [9483]));
Q_ASSIGN U6908 ( .B(clk), .A(\g.we_clk [9482]));
Q_ASSIGN U6909 ( .B(clk), .A(\g.we_clk [9481]));
Q_ASSIGN U6910 ( .B(clk), .A(\g.we_clk [9480]));
Q_ASSIGN U6911 ( .B(clk), .A(\g.we_clk [9479]));
Q_ASSIGN U6912 ( .B(clk), .A(\g.we_clk [9478]));
Q_ASSIGN U6913 ( .B(clk), .A(\g.we_clk [9477]));
Q_ASSIGN U6914 ( .B(clk), .A(\g.we_clk [9476]));
Q_ASSIGN U6915 ( .B(clk), .A(\g.we_clk [9475]));
Q_ASSIGN U6916 ( .B(clk), .A(\g.we_clk [9474]));
Q_ASSIGN U6917 ( .B(clk), .A(\g.we_clk [9473]));
Q_ASSIGN U6918 ( .B(clk), .A(\g.we_clk [9472]));
Q_ASSIGN U6919 ( .B(clk), .A(\g.we_clk [9471]));
Q_ASSIGN U6920 ( .B(clk), .A(\g.we_clk [9470]));
Q_ASSIGN U6921 ( .B(clk), .A(\g.we_clk [9469]));
Q_ASSIGN U6922 ( .B(clk), .A(\g.we_clk [9468]));
Q_ASSIGN U6923 ( .B(clk), .A(\g.we_clk [9467]));
Q_ASSIGN U6924 ( .B(clk), .A(\g.we_clk [9466]));
Q_ASSIGN U6925 ( .B(clk), .A(\g.we_clk [9465]));
Q_ASSIGN U6926 ( .B(clk), .A(\g.we_clk [9464]));
Q_ASSIGN U6927 ( .B(clk), .A(\g.we_clk [9463]));
Q_ASSIGN U6928 ( .B(clk), .A(\g.we_clk [9462]));
Q_ASSIGN U6929 ( .B(clk), .A(\g.we_clk [9461]));
Q_ASSIGN U6930 ( .B(clk), .A(\g.we_clk [9460]));
Q_ASSIGN U6931 ( .B(clk), .A(\g.we_clk [9459]));
Q_ASSIGN U6932 ( .B(clk), .A(\g.we_clk [9458]));
Q_ASSIGN U6933 ( .B(clk), .A(\g.we_clk [9457]));
Q_ASSIGN U6934 ( .B(clk), .A(\g.we_clk [9456]));
Q_ASSIGN U6935 ( .B(clk), .A(\g.we_clk [9455]));
Q_ASSIGN U6936 ( .B(clk), .A(\g.we_clk [9454]));
Q_ASSIGN U6937 ( .B(clk), .A(\g.we_clk [9453]));
Q_ASSIGN U6938 ( .B(clk), .A(\g.we_clk [9452]));
Q_ASSIGN U6939 ( .B(clk), .A(\g.we_clk [9451]));
Q_ASSIGN U6940 ( .B(clk), .A(\g.we_clk [9450]));
Q_ASSIGN U6941 ( .B(clk), .A(\g.we_clk [9449]));
Q_ASSIGN U6942 ( .B(clk), .A(\g.we_clk [9448]));
Q_ASSIGN U6943 ( .B(clk), .A(\g.we_clk [9447]));
Q_ASSIGN U6944 ( .B(clk), .A(\g.we_clk [9446]));
Q_ASSIGN U6945 ( .B(clk), .A(\g.we_clk [9445]));
Q_ASSIGN U6946 ( .B(clk), .A(\g.we_clk [9444]));
Q_ASSIGN U6947 ( .B(clk), .A(\g.we_clk [9443]));
Q_ASSIGN U6948 ( .B(clk), .A(\g.we_clk [9442]));
Q_ASSIGN U6949 ( .B(clk), .A(\g.we_clk [9441]));
Q_ASSIGN U6950 ( .B(clk), .A(\g.we_clk [9440]));
Q_ASSIGN U6951 ( .B(clk), .A(\g.we_clk [9439]));
Q_ASSIGN U6952 ( .B(clk), .A(\g.we_clk [9438]));
Q_ASSIGN U6953 ( .B(clk), .A(\g.we_clk [9437]));
Q_ASSIGN U6954 ( .B(clk), .A(\g.we_clk [9436]));
Q_ASSIGN U6955 ( .B(clk), .A(\g.we_clk [9435]));
Q_ASSIGN U6956 ( .B(clk), .A(\g.we_clk [9434]));
Q_ASSIGN U6957 ( .B(clk), .A(\g.we_clk [9433]));
Q_ASSIGN U6958 ( .B(clk), .A(\g.we_clk [9432]));
Q_ASSIGN U6959 ( .B(clk), .A(\g.we_clk [9431]));
Q_ASSIGN U6960 ( .B(clk), .A(\g.we_clk [9430]));
Q_ASSIGN U6961 ( .B(clk), .A(\g.we_clk [9429]));
Q_ASSIGN U6962 ( .B(clk), .A(\g.we_clk [9428]));
Q_ASSIGN U6963 ( .B(clk), .A(\g.we_clk [9427]));
Q_ASSIGN U6964 ( .B(clk), .A(\g.we_clk [9426]));
Q_ASSIGN U6965 ( .B(clk), .A(\g.we_clk [9425]));
Q_ASSIGN U6966 ( .B(clk), .A(\g.we_clk [9424]));
Q_ASSIGN U6967 ( .B(clk), .A(\g.we_clk [9423]));
Q_ASSIGN U6968 ( .B(clk), .A(\g.we_clk [9422]));
Q_ASSIGN U6969 ( .B(clk), .A(\g.we_clk [9421]));
Q_ASSIGN U6970 ( .B(clk), .A(\g.we_clk [9420]));
Q_ASSIGN U6971 ( .B(clk), .A(\g.we_clk [9419]));
Q_ASSIGN U6972 ( .B(clk), .A(\g.we_clk [9418]));
Q_ASSIGN U6973 ( .B(clk), .A(\g.we_clk [9417]));
Q_ASSIGN U6974 ( .B(clk), .A(\g.we_clk [9416]));
Q_ASSIGN U6975 ( .B(clk), .A(\g.we_clk [9415]));
Q_ASSIGN U6976 ( .B(clk), .A(\g.we_clk [9414]));
Q_ASSIGN U6977 ( .B(clk), .A(\g.we_clk [9413]));
Q_ASSIGN U6978 ( .B(clk), .A(\g.we_clk [9412]));
Q_ASSIGN U6979 ( .B(clk), .A(\g.we_clk [9411]));
Q_ASSIGN U6980 ( .B(clk), .A(\g.we_clk [9410]));
Q_ASSIGN U6981 ( .B(clk), .A(\g.we_clk [9409]));
Q_ASSIGN U6982 ( .B(clk), .A(\g.we_clk [9408]));
Q_ASSIGN U6983 ( .B(clk), .A(\g.we_clk [9407]));
Q_ASSIGN U6984 ( .B(clk), .A(\g.we_clk [9406]));
Q_ASSIGN U6985 ( .B(clk), .A(\g.we_clk [9405]));
Q_ASSIGN U6986 ( .B(clk), .A(\g.we_clk [9404]));
Q_ASSIGN U6987 ( .B(clk), .A(\g.we_clk [9403]));
Q_ASSIGN U6988 ( .B(clk), .A(\g.we_clk [9402]));
Q_ASSIGN U6989 ( .B(clk), .A(\g.we_clk [9401]));
Q_ASSIGN U6990 ( .B(clk), .A(\g.we_clk [9400]));
Q_ASSIGN U6991 ( .B(clk), .A(\g.we_clk [9399]));
Q_ASSIGN U6992 ( .B(clk), .A(\g.we_clk [9398]));
Q_ASSIGN U6993 ( .B(clk), .A(\g.we_clk [9397]));
Q_ASSIGN U6994 ( .B(clk), .A(\g.we_clk [9396]));
Q_ASSIGN U6995 ( .B(clk), .A(\g.we_clk [9395]));
Q_ASSIGN U6996 ( .B(clk), .A(\g.we_clk [9394]));
Q_ASSIGN U6997 ( .B(clk), .A(\g.we_clk [9393]));
Q_ASSIGN U6998 ( .B(clk), .A(\g.we_clk [9392]));
Q_ASSIGN U6999 ( .B(clk), .A(\g.we_clk [9391]));
Q_ASSIGN U7000 ( .B(clk), .A(\g.we_clk [9390]));
Q_ASSIGN U7001 ( .B(clk), .A(\g.we_clk [9389]));
Q_ASSIGN U7002 ( .B(clk), .A(\g.we_clk [9388]));
Q_ASSIGN U7003 ( .B(clk), .A(\g.we_clk [9387]));
Q_ASSIGN U7004 ( .B(clk), .A(\g.we_clk [9386]));
Q_ASSIGN U7005 ( .B(clk), .A(\g.we_clk [9385]));
Q_ASSIGN U7006 ( .B(clk), .A(\g.we_clk [9384]));
Q_ASSIGN U7007 ( .B(clk), .A(\g.we_clk [9383]));
Q_ASSIGN U7008 ( .B(clk), .A(\g.we_clk [9382]));
Q_ASSIGN U7009 ( .B(clk), .A(\g.we_clk [9381]));
Q_ASSIGN U7010 ( .B(clk), .A(\g.we_clk [9380]));
Q_ASSIGN U7011 ( .B(clk), .A(\g.we_clk [9379]));
Q_ASSIGN U7012 ( .B(clk), .A(\g.we_clk [9378]));
Q_ASSIGN U7013 ( .B(clk), .A(\g.we_clk [9377]));
Q_ASSIGN U7014 ( .B(clk), .A(\g.we_clk [9376]));
Q_ASSIGN U7015 ( .B(clk), .A(\g.we_clk [9375]));
Q_ASSIGN U7016 ( .B(clk), .A(\g.we_clk [9374]));
Q_ASSIGN U7017 ( .B(clk), .A(\g.we_clk [9373]));
Q_ASSIGN U7018 ( .B(clk), .A(\g.we_clk [9372]));
Q_ASSIGN U7019 ( .B(clk), .A(\g.we_clk [9371]));
Q_ASSIGN U7020 ( .B(clk), .A(\g.we_clk [9370]));
Q_ASSIGN U7021 ( .B(clk), .A(\g.we_clk [9369]));
Q_ASSIGN U7022 ( .B(clk), .A(\g.we_clk [9368]));
Q_ASSIGN U7023 ( .B(clk), .A(\g.we_clk [9367]));
Q_ASSIGN U7024 ( .B(clk), .A(\g.we_clk [9366]));
Q_ASSIGN U7025 ( .B(clk), .A(\g.we_clk [9365]));
Q_ASSIGN U7026 ( .B(clk), .A(\g.we_clk [9364]));
Q_ASSIGN U7027 ( .B(clk), .A(\g.we_clk [9363]));
Q_ASSIGN U7028 ( .B(clk), .A(\g.we_clk [9362]));
Q_ASSIGN U7029 ( .B(clk), .A(\g.we_clk [9361]));
Q_ASSIGN U7030 ( .B(clk), .A(\g.we_clk [9360]));
Q_ASSIGN U7031 ( .B(clk), .A(\g.we_clk [9359]));
Q_ASSIGN U7032 ( .B(clk), .A(\g.we_clk [9358]));
Q_ASSIGN U7033 ( .B(clk), .A(\g.we_clk [9357]));
Q_ASSIGN U7034 ( .B(clk), .A(\g.we_clk [9356]));
Q_ASSIGN U7035 ( .B(clk), .A(\g.we_clk [9355]));
Q_ASSIGN U7036 ( .B(clk), .A(\g.we_clk [9354]));
Q_ASSIGN U7037 ( .B(clk), .A(\g.we_clk [9353]));
Q_ASSIGN U7038 ( .B(clk), .A(\g.we_clk [9352]));
Q_ASSIGN U7039 ( .B(clk), .A(\g.we_clk [9351]));
Q_ASSIGN U7040 ( .B(clk), .A(\g.we_clk [9350]));
Q_ASSIGN U7041 ( .B(clk), .A(\g.we_clk [9349]));
Q_ASSIGN U7042 ( .B(clk), .A(\g.we_clk [9348]));
Q_ASSIGN U7043 ( .B(clk), .A(\g.we_clk [9347]));
Q_ASSIGN U7044 ( .B(clk), .A(\g.we_clk [9346]));
Q_ASSIGN U7045 ( .B(clk), .A(\g.we_clk [9345]));
Q_ASSIGN U7046 ( .B(clk), .A(\g.we_clk [9344]));
Q_ASSIGN U7047 ( .B(clk), .A(\g.we_clk [9343]));
Q_ASSIGN U7048 ( .B(clk), .A(\g.we_clk [9342]));
Q_ASSIGN U7049 ( .B(clk), .A(\g.we_clk [9341]));
Q_ASSIGN U7050 ( .B(clk), .A(\g.we_clk [9340]));
Q_ASSIGN U7051 ( .B(clk), .A(\g.we_clk [9339]));
Q_ASSIGN U7052 ( .B(clk), .A(\g.we_clk [9338]));
Q_ASSIGN U7053 ( .B(clk), .A(\g.we_clk [9337]));
Q_ASSIGN U7054 ( .B(clk), .A(\g.we_clk [9336]));
Q_ASSIGN U7055 ( .B(clk), .A(\g.we_clk [9335]));
Q_ASSIGN U7056 ( .B(clk), .A(\g.we_clk [9334]));
Q_ASSIGN U7057 ( .B(clk), .A(\g.we_clk [9333]));
Q_ASSIGN U7058 ( .B(clk), .A(\g.we_clk [9332]));
Q_ASSIGN U7059 ( .B(clk), .A(\g.we_clk [9331]));
Q_ASSIGN U7060 ( .B(clk), .A(\g.we_clk [9330]));
Q_ASSIGN U7061 ( .B(clk), .A(\g.we_clk [9329]));
Q_ASSIGN U7062 ( .B(clk), .A(\g.we_clk [9328]));
Q_ASSIGN U7063 ( .B(clk), .A(\g.we_clk [9327]));
Q_ASSIGN U7064 ( .B(clk), .A(\g.we_clk [9326]));
Q_ASSIGN U7065 ( .B(clk), .A(\g.we_clk [9325]));
Q_ASSIGN U7066 ( .B(clk), .A(\g.we_clk [9324]));
Q_ASSIGN U7067 ( .B(clk), .A(\g.we_clk [9323]));
Q_ASSIGN U7068 ( .B(clk), .A(\g.we_clk [9322]));
Q_ASSIGN U7069 ( .B(clk), .A(\g.we_clk [9321]));
Q_ASSIGN U7070 ( .B(clk), .A(\g.we_clk [9320]));
Q_ASSIGN U7071 ( .B(clk), .A(\g.we_clk [9319]));
Q_ASSIGN U7072 ( .B(clk), .A(\g.we_clk [9318]));
Q_ASSIGN U7073 ( .B(clk), .A(\g.we_clk [9317]));
Q_ASSIGN U7074 ( .B(clk), .A(\g.we_clk [9316]));
Q_ASSIGN U7075 ( .B(clk), .A(\g.we_clk [9315]));
Q_ASSIGN U7076 ( .B(clk), .A(\g.we_clk [9314]));
Q_ASSIGN U7077 ( .B(clk), .A(\g.we_clk [9313]));
Q_ASSIGN U7078 ( .B(clk), .A(\g.we_clk [9312]));
Q_ASSIGN U7079 ( .B(clk), .A(\g.we_clk [9311]));
Q_ASSIGN U7080 ( .B(clk), .A(\g.we_clk [9310]));
Q_ASSIGN U7081 ( .B(clk), .A(\g.we_clk [9309]));
Q_ASSIGN U7082 ( .B(clk), .A(\g.we_clk [9308]));
Q_ASSIGN U7083 ( .B(clk), .A(\g.we_clk [9307]));
Q_ASSIGN U7084 ( .B(clk), .A(\g.we_clk [9306]));
Q_ASSIGN U7085 ( .B(clk), .A(\g.we_clk [9305]));
Q_ASSIGN U7086 ( .B(clk), .A(\g.we_clk [9304]));
Q_ASSIGN U7087 ( .B(clk), .A(\g.we_clk [9303]));
Q_ASSIGN U7088 ( .B(clk), .A(\g.we_clk [9302]));
Q_ASSIGN U7089 ( .B(clk), .A(\g.we_clk [9301]));
Q_ASSIGN U7090 ( .B(clk), .A(\g.we_clk [9300]));
Q_ASSIGN U7091 ( .B(clk), .A(\g.we_clk [9299]));
Q_ASSIGN U7092 ( .B(clk), .A(\g.we_clk [9298]));
Q_ASSIGN U7093 ( .B(clk), .A(\g.we_clk [9297]));
Q_ASSIGN U7094 ( .B(clk), .A(\g.we_clk [9296]));
Q_ASSIGN U7095 ( .B(clk), .A(\g.we_clk [9295]));
Q_ASSIGN U7096 ( .B(clk), .A(\g.we_clk [9294]));
Q_ASSIGN U7097 ( .B(clk), .A(\g.we_clk [9293]));
Q_ASSIGN U7098 ( .B(clk), .A(\g.we_clk [9292]));
Q_ASSIGN U7099 ( .B(clk), .A(\g.we_clk [9291]));
Q_ASSIGN U7100 ( .B(clk), .A(\g.we_clk [9290]));
Q_ASSIGN U7101 ( .B(clk), .A(\g.we_clk [9289]));
Q_ASSIGN U7102 ( .B(clk), .A(\g.we_clk [9288]));
Q_ASSIGN U7103 ( .B(clk), .A(\g.we_clk [9287]));
Q_ASSIGN U7104 ( .B(clk), .A(\g.we_clk [9286]));
Q_ASSIGN U7105 ( .B(clk), .A(\g.we_clk [9285]));
Q_ASSIGN U7106 ( .B(clk), .A(\g.we_clk [9284]));
Q_ASSIGN U7107 ( .B(clk), .A(\g.we_clk [9283]));
Q_ASSIGN U7108 ( .B(clk), .A(\g.we_clk [9282]));
Q_ASSIGN U7109 ( .B(clk), .A(\g.we_clk [9281]));
Q_ASSIGN U7110 ( .B(clk), .A(\g.we_clk [9280]));
Q_ASSIGN U7111 ( .B(clk), .A(\g.we_clk [9279]));
Q_ASSIGN U7112 ( .B(clk), .A(\g.we_clk [9278]));
Q_ASSIGN U7113 ( .B(clk), .A(\g.we_clk [9277]));
Q_ASSIGN U7114 ( .B(clk), .A(\g.we_clk [9276]));
Q_ASSIGN U7115 ( .B(clk), .A(\g.we_clk [9275]));
Q_ASSIGN U7116 ( .B(clk), .A(\g.we_clk [9274]));
Q_ASSIGN U7117 ( .B(clk), .A(\g.we_clk [9273]));
Q_ASSIGN U7118 ( .B(clk), .A(\g.we_clk [9272]));
Q_ASSIGN U7119 ( .B(clk), .A(\g.we_clk [9271]));
Q_ASSIGN U7120 ( .B(clk), .A(\g.we_clk [9270]));
Q_ASSIGN U7121 ( .B(clk), .A(\g.we_clk [9269]));
Q_ASSIGN U7122 ( .B(clk), .A(\g.we_clk [9268]));
Q_ASSIGN U7123 ( .B(clk), .A(\g.we_clk [9267]));
Q_ASSIGN U7124 ( .B(clk), .A(\g.we_clk [9266]));
Q_ASSIGN U7125 ( .B(clk), .A(\g.we_clk [9265]));
Q_ASSIGN U7126 ( .B(clk), .A(\g.we_clk [9264]));
Q_ASSIGN U7127 ( .B(clk), .A(\g.we_clk [9263]));
Q_ASSIGN U7128 ( .B(clk), .A(\g.we_clk [9262]));
Q_ASSIGN U7129 ( .B(clk), .A(\g.we_clk [9261]));
Q_ASSIGN U7130 ( .B(clk), .A(\g.we_clk [9260]));
Q_ASSIGN U7131 ( .B(clk), .A(\g.we_clk [9259]));
Q_ASSIGN U7132 ( .B(clk), .A(\g.we_clk [9258]));
Q_ASSIGN U7133 ( .B(clk), .A(\g.we_clk [9257]));
Q_ASSIGN U7134 ( .B(clk), .A(\g.we_clk [9256]));
Q_ASSIGN U7135 ( .B(clk), .A(\g.we_clk [9255]));
Q_ASSIGN U7136 ( .B(clk), .A(\g.we_clk [9254]));
Q_ASSIGN U7137 ( .B(clk), .A(\g.we_clk [9253]));
Q_ASSIGN U7138 ( .B(clk), .A(\g.we_clk [9252]));
Q_ASSIGN U7139 ( .B(clk), .A(\g.we_clk [9251]));
Q_ASSIGN U7140 ( .B(clk), .A(\g.we_clk [9250]));
Q_ASSIGN U7141 ( .B(clk), .A(\g.we_clk [9249]));
Q_ASSIGN U7142 ( .B(clk), .A(\g.we_clk [9248]));
Q_ASSIGN U7143 ( .B(clk), .A(\g.we_clk [9247]));
Q_ASSIGN U7144 ( .B(clk), .A(\g.we_clk [9246]));
Q_ASSIGN U7145 ( .B(clk), .A(\g.we_clk [9245]));
Q_ASSIGN U7146 ( .B(clk), .A(\g.we_clk [9244]));
Q_ASSIGN U7147 ( .B(clk), .A(\g.we_clk [9243]));
Q_ASSIGN U7148 ( .B(clk), .A(\g.we_clk [9242]));
Q_ASSIGN U7149 ( .B(clk), .A(\g.we_clk [9241]));
Q_ASSIGN U7150 ( .B(clk), .A(\g.we_clk [9240]));
Q_ASSIGN U7151 ( .B(clk), .A(\g.we_clk [9239]));
Q_ASSIGN U7152 ( .B(clk), .A(\g.we_clk [9238]));
Q_ASSIGN U7153 ( .B(clk), .A(\g.we_clk [9237]));
Q_ASSIGN U7154 ( .B(clk), .A(\g.we_clk [9236]));
Q_ASSIGN U7155 ( .B(clk), .A(\g.we_clk [9235]));
Q_ASSIGN U7156 ( .B(clk), .A(\g.we_clk [9234]));
Q_ASSIGN U7157 ( .B(clk), .A(\g.we_clk [9233]));
Q_ASSIGN U7158 ( .B(clk), .A(\g.we_clk [9232]));
Q_ASSIGN U7159 ( .B(clk), .A(\g.we_clk [9231]));
Q_ASSIGN U7160 ( .B(clk), .A(\g.we_clk [9230]));
Q_ASSIGN U7161 ( .B(clk), .A(\g.we_clk [9229]));
Q_ASSIGN U7162 ( .B(clk), .A(\g.we_clk [9228]));
Q_ASSIGN U7163 ( .B(clk), .A(\g.we_clk [9227]));
Q_ASSIGN U7164 ( .B(clk), .A(\g.we_clk [9226]));
Q_ASSIGN U7165 ( .B(clk), .A(\g.we_clk [9225]));
Q_ASSIGN U7166 ( .B(clk), .A(\g.we_clk [9224]));
Q_ASSIGN U7167 ( .B(clk), .A(\g.we_clk [9223]));
Q_ASSIGN U7168 ( .B(clk), .A(\g.we_clk [9222]));
Q_ASSIGN U7169 ( .B(clk), .A(\g.we_clk [9221]));
Q_ASSIGN U7170 ( .B(clk), .A(\g.we_clk [9220]));
Q_ASSIGN U7171 ( .B(clk), .A(\g.we_clk [9219]));
Q_ASSIGN U7172 ( .B(clk), .A(\g.we_clk [9218]));
Q_ASSIGN U7173 ( .B(clk), .A(\g.we_clk [9217]));
Q_ASSIGN U7174 ( .B(clk), .A(\g.we_clk [9216]));
Q_ASSIGN U7175 ( .B(clk), .A(\g.we_clk [9215]));
Q_ASSIGN U7176 ( .B(clk), .A(\g.we_clk [9214]));
Q_ASSIGN U7177 ( .B(clk), .A(\g.we_clk [9213]));
Q_ASSIGN U7178 ( .B(clk), .A(\g.we_clk [9212]));
Q_ASSIGN U7179 ( .B(clk), .A(\g.we_clk [9211]));
Q_ASSIGN U7180 ( .B(clk), .A(\g.we_clk [9210]));
Q_ASSIGN U7181 ( .B(clk), .A(\g.we_clk [9209]));
Q_ASSIGN U7182 ( .B(clk), .A(\g.we_clk [9208]));
Q_ASSIGN U7183 ( .B(clk), .A(\g.we_clk [9207]));
Q_ASSIGN U7184 ( .B(clk), .A(\g.we_clk [9206]));
Q_ASSIGN U7185 ( .B(clk), .A(\g.we_clk [9205]));
Q_ASSIGN U7186 ( .B(clk), .A(\g.we_clk [9204]));
Q_ASSIGN U7187 ( .B(clk), .A(\g.we_clk [9203]));
Q_ASSIGN U7188 ( .B(clk), .A(\g.we_clk [9202]));
Q_ASSIGN U7189 ( .B(clk), .A(\g.we_clk [9201]));
Q_ASSIGN U7190 ( .B(clk), .A(\g.we_clk [9200]));
Q_ASSIGN U7191 ( .B(clk), .A(\g.we_clk [9199]));
Q_ASSIGN U7192 ( .B(clk), .A(\g.we_clk [9198]));
Q_ASSIGN U7193 ( .B(clk), .A(\g.we_clk [9197]));
Q_ASSIGN U7194 ( .B(clk), .A(\g.we_clk [9196]));
Q_ASSIGN U7195 ( .B(clk), .A(\g.we_clk [9195]));
Q_ASSIGN U7196 ( .B(clk), .A(\g.we_clk [9194]));
Q_ASSIGN U7197 ( .B(clk), .A(\g.we_clk [9193]));
Q_ASSIGN U7198 ( .B(clk), .A(\g.we_clk [9192]));
Q_ASSIGN U7199 ( .B(clk), .A(\g.we_clk [9191]));
Q_ASSIGN U7200 ( .B(clk), .A(\g.we_clk [9190]));
Q_ASSIGN U7201 ( .B(clk), .A(\g.we_clk [9189]));
Q_ASSIGN U7202 ( .B(clk), .A(\g.we_clk [9188]));
Q_ASSIGN U7203 ( .B(clk), .A(\g.we_clk [9187]));
Q_ASSIGN U7204 ( .B(clk), .A(\g.we_clk [9186]));
Q_ASSIGN U7205 ( .B(clk), .A(\g.we_clk [9185]));
Q_ASSIGN U7206 ( .B(clk), .A(\g.we_clk [9184]));
Q_ASSIGN U7207 ( .B(clk), .A(\g.we_clk [9183]));
Q_ASSIGN U7208 ( .B(clk), .A(\g.we_clk [9182]));
Q_ASSIGN U7209 ( .B(clk), .A(\g.we_clk [9181]));
Q_ASSIGN U7210 ( .B(clk), .A(\g.we_clk [9180]));
Q_ASSIGN U7211 ( .B(clk), .A(\g.we_clk [9179]));
Q_ASSIGN U7212 ( .B(clk), .A(\g.we_clk [9178]));
Q_ASSIGN U7213 ( .B(clk), .A(\g.we_clk [9177]));
Q_ASSIGN U7214 ( .B(clk), .A(\g.we_clk [9176]));
Q_ASSIGN U7215 ( .B(clk), .A(\g.we_clk [9175]));
Q_ASSIGN U7216 ( .B(clk), .A(\g.we_clk [9174]));
Q_ASSIGN U7217 ( .B(clk), .A(\g.we_clk [9173]));
Q_ASSIGN U7218 ( .B(clk), .A(\g.we_clk [9172]));
Q_ASSIGN U7219 ( .B(clk), .A(\g.we_clk [9171]));
Q_ASSIGN U7220 ( .B(clk), .A(\g.we_clk [9170]));
Q_ASSIGN U7221 ( .B(clk), .A(\g.we_clk [9169]));
Q_ASSIGN U7222 ( .B(clk), .A(\g.we_clk [9168]));
Q_ASSIGN U7223 ( .B(clk), .A(\g.we_clk [9167]));
Q_ASSIGN U7224 ( .B(clk), .A(\g.we_clk [9166]));
Q_ASSIGN U7225 ( .B(clk), .A(\g.we_clk [9165]));
Q_ASSIGN U7226 ( .B(clk), .A(\g.we_clk [9164]));
Q_ASSIGN U7227 ( .B(clk), .A(\g.we_clk [9163]));
Q_ASSIGN U7228 ( .B(clk), .A(\g.we_clk [9162]));
Q_ASSIGN U7229 ( .B(clk), .A(\g.we_clk [9161]));
Q_ASSIGN U7230 ( .B(clk), .A(\g.we_clk [9160]));
Q_ASSIGN U7231 ( .B(clk), .A(\g.we_clk [9159]));
Q_ASSIGN U7232 ( .B(clk), .A(\g.we_clk [9158]));
Q_ASSIGN U7233 ( .B(clk), .A(\g.we_clk [9157]));
Q_ASSIGN U7234 ( .B(clk), .A(\g.we_clk [9156]));
Q_ASSIGN U7235 ( .B(clk), .A(\g.we_clk [9155]));
Q_ASSIGN U7236 ( .B(clk), .A(\g.we_clk [9154]));
Q_ASSIGN U7237 ( .B(clk), .A(\g.we_clk [9153]));
Q_ASSIGN U7238 ( .B(clk), .A(\g.we_clk [9152]));
Q_ASSIGN U7239 ( .B(clk), .A(\g.we_clk [9151]));
Q_ASSIGN U7240 ( .B(clk), .A(\g.we_clk [9150]));
Q_ASSIGN U7241 ( .B(clk), .A(\g.we_clk [9149]));
Q_ASSIGN U7242 ( .B(clk), .A(\g.we_clk [9148]));
Q_ASSIGN U7243 ( .B(clk), .A(\g.we_clk [9147]));
Q_ASSIGN U7244 ( .B(clk), .A(\g.we_clk [9146]));
Q_ASSIGN U7245 ( .B(clk), .A(\g.we_clk [9145]));
Q_ASSIGN U7246 ( .B(clk), .A(\g.we_clk [9144]));
Q_ASSIGN U7247 ( .B(clk), .A(\g.we_clk [9143]));
Q_ASSIGN U7248 ( .B(clk), .A(\g.we_clk [9142]));
Q_ASSIGN U7249 ( .B(clk), .A(\g.we_clk [9141]));
Q_ASSIGN U7250 ( .B(clk), .A(\g.we_clk [9140]));
Q_ASSIGN U7251 ( .B(clk), .A(\g.we_clk [9139]));
Q_ASSIGN U7252 ( .B(clk), .A(\g.we_clk [9138]));
Q_ASSIGN U7253 ( .B(clk), .A(\g.we_clk [9137]));
Q_ASSIGN U7254 ( .B(clk), .A(\g.we_clk [9136]));
Q_ASSIGN U7255 ( .B(clk), .A(\g.we_clk [9135]));
Q_ASSIGN U7256 ( .B(clk), .A(\g.we_clk [9134]));
Q_ASSIGN U7257 ( .B(clk), .A(\g.we_clk [9133]));
Q_ASSIGN U7258 ( .B(clk), .A(\g.we_clk [9132]));
Q_ASSIGN U7259 ( .B(clk), .A(\g.we_clk [9131]));
Q_ASSIGN U7260 ( .B(clk), .A(\g.we_clk [9130]));
Q_ASSIGN U7261 ( .B(clk), .A(\g.we_clk [9129]));
Q_ASSIGN U7262 ( .B(clk), .A(\g.we_clk [9128]));
Q_ASSIGN U7263 ( .B(clk), .A(\g.we_clk [9127]));
Q_ASSIGN U7264 ( .B(clk), .A(\g.we_clk [9126]));
Q_ASSIGN U7265 ( .B(clk), .A(\g.we_clk [9125]));
Q_ASSIGN U7266 ( .B(clk), .A(\g.we_clk [9124]));
Q_ASSIGN U7267 ( .B(clk), .A(\g.we_clk [9123]));
Q_ASSIGN U7268 ( .B(clk), .A(\g.we_clk [9122]));
Q_ASSIGN U7269 ( .B(clk), .A(\g.we_clk [9121]));
Q_ASSIGN U7270 ( .B(clk), .A(\g.we_clk [9120]));
Q_ASSIGN U7271 ( .B(clk), .A(\g.we_clk [9119]));
Q_ASSIGN U7272 ( .B(clk), .A(\g.we_clk [9118]));
Q_ASSIGN U7273 ( .B(clk), .A(\g.we_clk [9117]));
Q_ASSIGN U7274 ( .B(clk), .A(\g.we_clk [9116]));
Q_ASSIGN U7275 ( .B(clk), .A(\g.we_clk [9115]));
Q_ASSIGN U7276 ( .B(clk), .A(\g.we_clk [9114]));
Q_ASSIGN U7277 ( .B(clk), .A(\g.we_clk [9113]));
Q_ASSIGN U7278 ( .B(clk), .A(\g.we_clk [9112]));
Q_ASSIGN U7279 ( .B(clk), .A(\g.we_clk [9111]));
Q_ASSIGN U7280 ( .B(clk), .A(\g.we_clk [9110]));
Q_ASSIGN U7281 ( .B(clk), .A(\g.we_clk [9109]));
Q_ASSIGN U7282 ( .B(clk), .A(\g.we_clk [9108]));
Q_ASSIGN U7283 ( .B(clk), .A(\g.we_clk [9107]));
Q_ASSIGN U7284 ( .B(clk), .A(\g.we_clk [9106]));
Q_ASSIGN U7285 ( .B(clk), .A(\g.we_clk [9105]));
Q_ASSIGN U7286 ( .B(clk), .A(\g.we_clk [9104]));
Q_ASSIGN U7287 ( .B(clk), .A(\g.we_clk [9103]));
Q_ASSIGN U7288 ( .B(clk), .A(\g.we_clk [9102]));
Q_ASSIGN U7289 ( .B(clk), .A(\g.we_clk [9101]));
Q_ASSIGN U7290 ( .B(clk), .A(\g.we_clk [9100]));
Q_ASSIGN U7291 ( .B(clk), .A(\g.we_clk [9099]));
Q_ASSIGN U7292 ( .B(clk), .A(\g.we_clk [9098]));
Q_ASSIGN U7293 ( .B(clk), .A(\g.we_clk [9097]));
Q_ASSIGN U7294 ( .B(clk), .A(\g.we_clk [9096]));
Q_ASSIGN U7295 ( .B(clk), .A(\g.we_clk [9095]));
Q_ASSIGN U7296 ( .B(clk), .A(\g.we_clk [9094]));
Q_ASSIGN U7297 ( .B(clk), .A(\g.we_clk [9093]));
Q_ASSIGN U7298 ( .B(clk), .A(\g.we_clk [9092]));
Q_ASSIGN U7299 ( .B(clk), .A(\g.we_clk [9091]));
Q_ASSIGN U7300 ( .B(clk), .A(\g.we_clk [9090]));
Q_ASSIGN U7301 ( .B(clk), .A(\g.we_clk [9089]));
Q_ASSIGN U7302 ( .B(clk), .A(\g.we_clk [9088]));
Q_ASSIGN U7303 ( .B(clk), .A(\g.we_clk [9087]));
Q_ASSIGN U7304 ( .B(clk), .A(\g.we_clk [9086]));
Q_ASSIGN U7305 ( .B(clk), .A(\g.we_clk [9085]));
Q_ASSIGN U7306 ( .B(clk), .A(\g.we_clk [9084]));
Q_ASSIGN U7307 ( .B(clk), .A(\g.we_clk [9083]));
Q_ASSIGN U7308 ( .B(clk), .A(\g.we_clk [9082]));
Q_ASSIGN U7309 ( .B(clk), .A(\g.we_clk [9081]));
Q_ASSIGN U7310 ( .B(clk), .A(\g.we_clk [9080]));
Q_ASSIGN U7311 ( .B(clk), .A(\g.we_clk [9079]));
Q_ASSIGN U7312 ( .B(clk), .A(\g.we_clk [9078]));
Q_ASSIGN U7313 ( .B(clk), .A(\g.we_clk [9077]));
Q_ASSIGN U7314 ( .B(clk), .A(\g.we_clk [9076]));
Q_ASSIGN U7315 ( .B(clk), .A(\g.we_clk [9075]));
Q_ASSIGN U7316 ( .B(clk), .A(\g.we_clk [9074]));
Q_ASSIGN U7317 ( .B(clk), .A(\g.we_clk [9073]));
Q_ASSIGN U7318 ( .B(clk), .A(\g.we_clk [9072]));
Q_ASSIGN U7319 ( .B(clk), .A(\g.we_clk [9071]));
Q_ASSIGN U7320 ( .B(clk), .A(\g.we_clk [9070]));
Q_ASSIGN U7321 ( .B(clk), .A(\g.we_clk [9069]));
Q_ASSIGN U7322 ( .B(clk), .A(\g.we_clk [9068]));
Q_ASSIGN U7323 ( .B(clk), .A(\g.we_clk [9067]));
Q_ASSIGN U7324 ( .B(clk), .A(\g.we_clk [9066]));
Q_ASSIGN U7325 ( .B(clk), .A(\g.we_clk [9065]));
Q_ASSIGN U7326 ( .B(clk), .A(\g.we_clk [9064]));
Q_ASSIGN U7327 ( .B(clk), .A(\g.we_clk [9063]));
Q_ASSIGN U7328 ( .B(clk), .A(\g.we_clk [9062]));
Q_ASSIGN U7329 ( .B(clk), .A(\g.we_clk [9061]));
Q_ASSIGN U7330 ( .B(clk), .A(\g.we_clk [9060]));
Q_ASSIGN U7331 ( .B(clk), .A(\g.we_clk [9059]));
Q_ASSIGN U7332 ( .B(clk), .A(\g.we_clk [9058]));
Q_ASSIGN U7333 ( .B(clk), .A(\g.we_clk [9057]));
Q_ASSIGN U7334 ( .B(clk), .A(\g.we_clk [9056]));
Q_ASSIGN U7335 ( .B(clk), .A(\g.we_clk [9055]));
Q_ASSIGN U7336 ( .B(clk), .A(\g.we_clk [9054]));
Q_ASSIGN U7337 ( .B(clk), .A(\g.we_clk [9053]));
Q_ASSIGN U7338 ( .B(clk), .A(\g.we_clk [9052]));
Q_ASSIGN U7339 ( .B(clk), .A(\g.we_clk [9051]));
Q_ASSIGN U7340 ( .B(clk), .A(\g.we_clk [9050]));
Q_ASSIGN U7341 ( .B(clk), .A(\g.we_clk [9049]));
Q_ASSIGN U7342 ( .B(clk), .A(\g.we_clk [9048]));
Q_ASSIGN U7343 ( .B(clk), .A(\g.we_clk [9047]));
Q_ASSIGN U7344 ( .B(clk), .A(\g.we_clk [9046]));
Q_ASSIGN U7345 ( .B(clk), .A(\g.we_clk [9045]));
Q_ASSIGN U7346 ( .B(clk), .A(\g.we_clk [9044]));
Q_ASSIGN U7347 ( .B(clk), .A(\g.we_clk [9043]));
Q_ASSIGN U7348 ( .B(clk), .A(\g.we_clk [9042]));
Q_ASSIGN U7349 ( .B(clk), .A(\g.we_clk [9041]));
Q_ASSIGN U7350 ( .B(clk), .A(\g.we_clk [9040]));
Q_ASSIGN U7351 ( .B(clk), .A(\g.we_clk [9039]));
Q_ASSIGN U7352 ( .B(clk), .A(\g.we_clk [9038]));
Q_ASSIGN U7353 ( .B(clk), .A(\g.we_clk [9037]));
Q_ASSIGN U7354 ( .B(clk), .A(\g.we_clk [9036]));
Q_ASSIGN U7355 ( .B(clk), .A(\g.we_clk [9035]));
Q_ASSIGN U7356 ( .B(clk), .A(\g.we_clk [9034]));
Q_ASSIGN U7357 ( .B(clk), .A(\g.we_clk [9033]));
Q_ASSIGN U7358 ( .B(clk), .A(\g.we_clk [9032]));
Q_ASSIGN U7359 ( .B(clk), .A(\g.we_clk [9031]));
Q_ASSIGN U7360 ( .B(clk), .A(\g.we_clk [9030]));
Q_ASSIGN U7361 ( .B(clk), .A(\g.we_clk [9029]));
Q_ASSIGN U7362 ( .B(clk), .A(\g.we_clk [9028]));
Q_ASSIGN U7363 ( .B(clk), .A(\g.we_clk [9027]));
Q_ASSIGN U7364 ( .B(clk), .A(\g.we_clk [9026]));
Q_ASSIGN U7365 ( .B(clk), .A(\g.we_clk [9025]));
Q_ASSIGN U7366 ( .B(clk), .A(\g.we_clk [9024]));
Q_ASSIGN U7367 ( .B(clk), .A(\g.we_clk [9023]));
Q_ASSIGN U7368 ( .B(clk), .A(\g.we_clk [9022]));
Q_ASSIGN U7369 ( .B(clk), .A(\g.we_clk [9021]));
Q_ASSIGN U7370 ( .B(clk), .A(\g.we_clk [9020]));
Q_ASSIGN U7371 ( .B(clk), .A(\g.we_clk [9019]));
Q_ASSIGN U7372 ( .B(clk), .A(\g.we_clk [9018]));
Q_ASSIGN U7373 ( .B(clk), .A(\g.we_clk [9017]));
Q_ASSIGN U7374 ( .B(clk), .A(\g.we_clk [9016]));
Q_ASSIGN U7375 ( .B(clk), .A(\g.we_clk [9015]));
Q_ASSIGN U7376 ( .B(clk), .A(\g.we_clk [9014]));
Q_ASSIGN U7377 ( .B(clk), .A(\g.we_clk [9013]));
Q_ASSIGN U7378 ( .B(clk), .A(\g.we_clk [9012]));
Q_ASSIGN U7379 ( .B(clk), .A(\g.we_clk [9011]));
Q_ASSIGN U7380 ( .B(clk), .A(\g.we_clk [9010]));
Q_ASSIGN U7381 ( .B(clk), .A(\g.we_clk [9009]));
Q_ASSIGN U7382 ( .B(clk), .A(\g.we_clk [9008]));
Q_ASSIGN U7383 ( .B(clk), .A(\g.we_clk [9007]));
Q_ASSIGN U7384 ( .B(clk), .A(\g.we_clk [9006]));
Q_ASSIGN U7385 ( .B(clk), .A(\g.we_clk [9005]));
Q_ASSIGN U7386 ( .B(clk), .A(\g.we_clk [9004]));
Q_ASSIGN U7387 ( .B(clk), .A(\g.we_clk [9003]));
Q_ASSIGN U7388 ( .B(clk), .A(\g.we_clk [9002]));
Q_ASSIGN U7389 ( .B(clk), .A(\g.we_clk [9001]));
Q_ASSIGN U7390 ( .B(clk), .A(\g.we_clk [9000]));
Q_ASSIGN U7391 ( .B(clk), .A(\g.we_clk [8999]));
Q_ASSIGN U7392 ( .B(clk), .A(\g.we_clk [8998]));
Q_ASSIGN U7393 ( .B(clk), .A(\g.we_clk [8997]));
Q_ASSIGN U7394 ( .B(clk), .A(\g.we_clk [8996]));
Q_ASSIGN U7395 ( .B(clk), .A(\g.we_clk [8995]));
Q_ASSIGN U7396 ( .B(clk), .A(\g.we_clk [8994]));
Q_ASSIGN U7397 ( .B(clk), .A(\g.we_clk [8993]));
Q_ASSIGN U7398 ( .B(clk), .A(\g.we_clk [8992]));
Q_ASSIGN U7399 ( .B(clk), .A(\g.we_clk [8991]));
Q_ASSIGN U7400 ( .B(clk), .A(\g.we_clk [8990]));
Q_ASSIGN U7401 ( .B(clk), .A(\g.we_clk [8989]));
Q_ASSIGN U7402 ( .B(clk), .A(\g.we_clk [8988]));
Q_ASSIGN U7403 ( .B(clk), .A(\g.we_clk [8987]));
Q_ASSIGN U7404 ( .B(clk), .A(\g.we_clk [8986]));
Q_ASSIGN U7405 ( .B(clk), .A(\g.we_clk [8985]));
Q_ASSIGN U7406 ( .B(clk), .A(\g.we_clk [8984]));
Q_ASSIGN U7407 ( .B(clk), .A(\g.we_clk [8983]));
Q_ASSIGN U7408 ( .B(clk), .A(\g.we_clk [8982]));
Q_ASSIGN U7409 ( .B(clk), .A(\g.we_clk [8981]));
Q_ASSIGN U7410 ( .B(clk), .A(\g.we_clk [8980]));
Q_ASSIGN U7411 ( .B(clk), .A(\g.we_clk [8979]));
Q_ASSIGN U7412 ( .B(clk), .A(\g.we_clk [8978]));
Q_ASSIGN U7413 ( .B(clk), .A(\g.we_clk [8977]));
Q_ASSIGN U7414 ( .B(clk), .A(\g.we_clk [8976]));
Q_ASSIGN U7415 ( .B(clk), .A(\g.we_clk [8975]));
Q_ASSIGN U7416 ( .B(clk), .A(\g.we_clk [8974]));
Q_ASSIGN U7417 ( .B(clk), .A(\g.we_clk [8973]));
Q_ASSIGN U7418 ( .B(clk), .A(\g.we_clk [8972]));
Q_ASSIGN U7419 ( .B(clk), .A(\g.we_clk [8971]));
Q_ASSIGN U7420 ( .B(clk), .A(\g.we_clk [8970]));
Q_ASSIGN U7421 ( .B(clk), .A(\g.we_clk [8969]));
Q_ASSIGN U7422 ( .B(clk), .A(\g.we_clk [8968]));
Q_ASSIGN U7423 ( .B(clk), .A(\g.we_clk [8967]));
Q_ASSIGN U7424 ( .B(clk), .A(\g.we_clk [8966]));
Q_ASSIGN U7425 ( .B(clk), .A(\g.we_clk [8965]));
Q_ASSIGN U7426 ( .B(clk), .A(\g.we_clk [8964]));
Q_ASSIGN U7427 ( .B(clk), .A(\g.we_clk [8963]));
Q_ASSIGN U7428 ( .B(clk), .A(\g.we_clk [8962]));
Q_ASSIGN U7429 ( .B(clk), .A(\g.we_clk [8961]));
Q_ASSIGN U7430 ( .B(clk), .A(\g.we_clk [8960]));
Q_ASSIGN U7431 ( .B(clk), .A(\g.we_clk [8959]));
Q_ASSIGN U7432 ( .B(clk), .A(\g.we_clk [8958]));
Q_ASSIGN U7433 ( .B(clk), .A(\g.we_clk [8957]));
Q_ASSIGN U7434 ( .B(clk), .A(\g.we_clk [8956]));
Q_ASSIGN U7435 ( .B(clk), .A(\g.we_clk [8955]));
Q_ASSIGN U7436 ( .B(clk), .A(\g.we_clk [8954]));
Q_ASSIGN U7437 ( .B(clk), .A(\g.we_clk [8953]));
Q_ASSIGN U7438 ( .B(clk), .A(\g.we_clk [8952]));
Q_ASSIGN U7439 ( .B(clk), .A(\g.we_clk [8951]));
Q_ASSIGN U7440 ( .B(clk), .A(\g.we_clk [8950]));
Q_ASSIGN U7441 ( .B(clk), .A(\g.we_clk [8949]));
Q_ASSIGN U7442 ( .B(clk), .A(\g.we_clk [8948]));
Q_ASSIGN U7443 ( .B(clk), .A(\g.we_clk [8947]));
Q_ASSIGN U7444 ( .B(clk), .A(\g.we_clk [8946]));
Q_ASSIGN U7445 ( .B(clk), .A(\g.we_clk [8945]));
Q_ASSIGN U7446 ( .B(clk), .A(\g.we_clk [8944]));
Q_ASSIGN U7447 ( .B(clk), .A(\g.we_clk [8943]));
Q_ASSIGN U7448 ( .B(clk), .A(\g.we_clk [8942]));
Q_ASSIGN U7449 ( .B(clk), .A(\g.we_clk [8941]));
Q_ASSIGN U7450 ( .B(clk), .A(\g.we_clk [8940]));
Q_ASSIGN U7451 ( .B(clk), .A(\g.we_clk [8939]));
Q_ASSIGN U7452 ( .B(clk), .A(\g.we_clk [8938]));
Q_ASSIGN U7453 ( .B(clk), .A(\g.we_clk [8937]));
Q_ASSIGN U7454 ( .B(clk), .A(\g.we_clk [8936]));
Q_ASSIGN U7455 ( .B(clk), .A(\g.we_clk [8935]));
Q_ASSIGN U7456 ( .B(clk), .A(\g.we_clk [8934]));
Q_ASSIGN U7457 ( .B(clk), .A(\g.we_clk [8933]));
Q_ASSIGN U7458 ( .B(clk), .A(\g.we_clk [8932]));
Q_ASSIGN U7459 ( .B(clk), .A(\g.we_clk [8931]));
Q_ASSIGN U7460 ( .B(clk), .A(\g.we_clk [8930]));
Q_ASSIGN U7461 ( .B(clk), .A(\g.we_clk [8929]));
Q_ASSIGN U7462 ( .B(clk), .A(\g.we_clk [8928]));
Q_ASSIGN U7463 ( .B(clk), .A(\g.we_clk [8927]));
Q_ASSIGN U7464 ( .B(clk), .A(\g.we_clk [8926]));
Q_ASSIGN U7465 ( .B(clk), .A(\g.we_clk [8925]));
Q_ASSIGN U7466 ( .B(clk), .A(\g.we_clk [8924]));
Q_ASSIGN U7467 ( .B(clk), .A(\g.we_clk [8923]));
Q_ASSIGN U7468 ( .B(clk), .A(\g.we_clk [8922]));
Q_ASSIGN U7469 ( .B(clk), .A(\g.we_clk [8921]));
Q_ASSIGN U7470 ( .B(clk), .A(\g.we_clk [8920]));
Q_ASSIGN U7471 ( .B(clk), .A(\g.we_clk [8919]));
Q_ASSIGN U7472 ( .B(clk), .A(\g.we_clk [8918]));
Q_ASSIGN U7473 ( .B(clk), .A(\g.we_clk [8917]));
Q_ASSIGN U7474 ( .B(clk), .A(\g.we_clk [8916]));
Q_ASSIGN U7475 ( .B(clk), .A(\g.we_clk [8915]));
Q_ASSIGN U7476 ( .B(clk), .A(\g.we_clk [8914]));
Q_ASSIGN U7477 ( .B(clk), .A(\g.we_clk [8913]));
Q_ASSIGN U7478 ( .B(clk), .A(\g.we_clk [8912]));
Q_ASSIGN U7479 ( .B(clk), .A(\g.we_clk [8911]));
Q_ASSIGN U7480 ( .B(clk), .A(\g.we_clk [8910]));
Q_ASSIGN U7481 ( .B(clk), .A(\g.we_clk [8909]));
Q_ASSIGN U7482 ( .B(clk), .A(\g.we_clk [8908]));
Q_ASSIGN U7483 ( .B(clk), .A(\g.we_clk [8907]));
Q_ASSIGN U7484 ( .B(clk), .A(\g.we_clk [8906]));
Q_ASSIGN U7485 ( .B(clk), .A(\g.we_clk [8905]));
Q_ASSIGN U7486 ( .B(clk), .A(\g.we_clk [8904]));
Q_ASSIGN U7487 ( .B(clk), .A(\g.we_clk [8903]));
Q_ASSIGN U7488 ( .B(clk), .A(\g.we_clk [8902]));
Q_ASSIGN U7489 ( .B(clk), .A(\g.we_clk [8901]));
Q_ASSIGN U7490 ( .B(clk), .A(\g.we_clk [8900]));
Q_ASSIGN U7491 ( .B(clk), .A(\g.we_clk [8899]));
Q_ASSIGN U7492 ( .B(clk), .A(\g.we_clk [8898]));
Q_ASSIGN U7493 ( .B(clk), .A(\g.we_clk [8897]));
Q_ASSIGN U7494 ( .B(clk), .A(\g.we_clk [8896]));
Q_ASSIGN U7495 ( .B(clk), .A(\g.we_clk [8895]));
Q_ASSIGN U7496 ( .B(clk), .A(\g.we_clk [8894]));
Q_ASSIGN U7497 ( .B(clk), .A(\g.we_clk [8893]));
Q_ASSIGN U7498 ( .B(clk), .A(\g.we_clk [8892]));
Q_ASSIGN U7499 ( .B(clk), .A(\g.we_clk [8891]));
Q_ASSIGN U7500 ( .B(clk), .A(\g.we_clk [8890]));
Q_ASSIGN U7501 ( .B(clk), .A(\g.we_clk [8889]));
Q_ASSIGN U7502 ( .B(clk), .A(\g.we_clk [8888]));
Q_ASSIGN U7503 ( .B(clk), .A(\g.we_clk [8887]));
Q_ASSIGN U7504 ( .B(clk), .A(\g.we_clk [8886]));
Q_ASSIGN U7505 ( .B(clk), .A(\g.we_clk [8885]));
Q_ASSIGN U7506 ( .B(clk), .A(\g.we_clk [8884]));
Q_ASSIGN U7507 ( .B(clk), .A(\g.we_clk [8883]));
Q_ASSIGN U7508 ( .B(clk), .A(\g.we_clk [8882]));
Q_ASSIGN U7509 ( .B(clk), .A(\g.we_clk [8881]));
Q_ASSIGN U7510 ( .B(clk), .A(\g.we_clk [8880]));
Q_ASSIGN U7511 ( .B(clk), .A(\g.we_clk [8879]));
Q_ASSIGN U7512 ( .B(clk), .A(\g.we_clk [8878]));
Q_ASSIGN U7513 ( .B(clk), .A(\g.we_clk [8877]));
Q_ASSIGN U7514 ( .B(clk), .A(\g.we_clk [8876]));
Q_ASSIGN U7515 ( .B(clk), .A(\g.we_clk [8875]));
Q_ASSIGN U7516 ( .B(clk), .A(\g.we_clk [8874]));
Q_ASSIGN U7517 ( .B(clk), .A(\g.we_clk [8873]));
Q_ASSIGN U7518 ( .B(clk), .A(\g.we_clk [8872]));
Q_ASSIGN U7519 ( .B(clk), .A(\g.we_clk [8871]));
Q_ASSIGN U7520 ( .B(clk), .A(\g.we_clk [8870]));
Q_ASSIGN U7521 ( .B(clk), .A(\g.we_clk [8869]));
Q_ASSIGN U7522 ( .B(clk), .A(\g.we_clk [8868]));
Q_ASSIGN U7523 ( .B(clk), .A(\g.we_clk [8867]));
Q_ASSIGN U7524 ( .B(clk), .A(\g.we_clk [8866]));
Q_ASSIGN U7525 ( .B(clk), .A(\g.we_clk [8865]));
Q_ASSIGN U7526 ( .B(clk), .A(\g.we_clk [8864]));
Q_ASSIGN U7527 ( .B(clk), .A(\g.we_clk [8863]));
Q_ASSIGN U7528 ( .B(clk), .A(\g.we_clk [8862]));
Q_ASSIGN U7529 ( .B(clk), .A(\g.we_clk [8861]));
Q_ASSIGN U7530 ( .B(clk), .A(\g.we_clk [8860]));
Q_ASSIGN U7531 ( .B(clk), .A(\g.we_clk [8859]));
Q_ASSIGN U7532 ( .B(clk), .A(\g.we_clk [8858]));
Q_ASSIGN U7533 ( .B(clk), .A(\g.we_clk [8857]));
Q_ASSIGN U7534 ( .B(clk), .A(\g.we_clk [8856]));
Q_ASSIGN U7535 ( .B(clk), .A(\g.we_clk [8855]));
Q_ASSIGN U7536 ( .B(clk), .A(\g.we_clk [8854]));
Q_ASSIGN U7537 ( .B(clk), .A(\g.we_clk [8853]));
Q_ASSIGN U7538 ( .B(clk), .A(\g.we_clk [8852]));
Q_ASSIGN U7539 ( .B(clk), .A(\g.we_clk [8851]));
Q_ASSIGN U7540 ( .B(clk), .A(\g.we_clk [8850]));
Q_ASSIGN U7541 ( .B(clk), .A(\g.we_clk [8849]));
Q_ASSIGN U7542 ( .B(clk), .A(\g.we_clk [8848]));
Q_ASSIGN U7543 ( .B(clk), .A(\g.we_clk [8847]));
Q_ASSIGN U7544 ( .B(clk), .A(\g.we_clk [8846]));
Q_ASSIGN U7545 ( .B(clk), .A(\g.we_clk [8845]));
Q_ASSIGN U7546 ( .B(clk), .A(\g.we_clk [8844]));
Q_ASSIGN U7547 ( .B(clk), .A(\g.we_clk [8843]));
Q_ASSIGN U7548 ( .B(clk), .A(\g.we_clk [8842]));
Q_ASSIGN U7549 ( .B(clk), .A(\g.we_clk [8841]));
Q_ASSIGN U7550 ( .B(clk), .A(\g.we_clk [8840]));
Q_ASSIGN U7551 ( .B(clk), .A(\g.we_clk [8839]));
Q_ASSIGN U7552 ( .B(clk), .A(\g.we_clk [8838]));
Q_ASSIGN U7553 ( .B(clk), .A(\g.we_clk [8837]));
Q_ASSIGN U7554 ( .B(clk), .A(\g.we_clk [8836]));
Q_ASSIGN U7555 ( .B(clk), .A(\g.we_clk [8835]));
Q_ASSIGN U7556 ( .B(clk), .A(\g.we_clk [8834]));
Q_ASSIGN U7557 ( .B(clk), .A(\g.we_clk [8833]));
Q_ASSIGN U7558 ( .B(clk), .A(\g.we_clk [8832]));
Q_ASSIGN U7559 ( .B(clk), .A(\g.we_clk [8831]));
Q_ASSIGN U7560 ( .B(clk), .A(\g.we_clk [8830]));
Q_ASSIGN U7561 ( .B(clk), .A(\g.we_clk [8829]));
Q_ASSIGN U7562 ( .B(clk), .A(\g.we_clk [8828]));
Q_ASSIGN U7563 ( .B(clk), .A(\g.we_clk [8827]));
Q_ASSIGN U7564 ( .B(clk), .A(\g.we_clk [8826]));
Q_ASSIGN U7565 ( .B(clk), .A(\g.we_clk [8825]));
Q_ASSIGN U7566 ( .B(clk), .A(\g.we_clk [8824]));
Q_ASSIGN U7567 ( .B(clk), .A(\g.we_clk [8823]));
Q_ASSIGN U7568 ( .B(clk), .A(\g.we_clk [8822]));
Q_ASSIGN U7569 ( .B(clk), .A(\g.we_clk [8821]));
Q_ASSIGN U7570 ( .B(clk), .A(\g.we_clk [8820]));
Q_ASSIGN U7571 ( .B(clk), .A(\g.we_clk [8819]));
Q_ASSIGN U7572 ( .B(clk), .A(\g.we_clk [8818]));
Q_ASSIGN U7573 ( .B(clk), .A(\g.we_clk [8817]));
Q_ASSIGN U7574 ( .B(clk), .A(\g.we_clk [8816]));
Q_ASSIGN U7575 ( .B(clk), .A(\g.we_clk [8815]));
Q_ASSIGN U7576 ( .B(clk), .A(\g.we_clk [8814]));
Q_ASSIGN U7577 ( .B(clk), .A(\g.we_clk [8813]));
Q_ASSIGN U7578 ( .B(clk), .A(\g.we_clk [8812]));
Q_ASSIGN U7579 ( .B(clk), .A(\g.we_clk [8811]));
Q_ASSIGN U7580 ( .B(clk), .A(\g.we_clk [8810]));
Q_ASSIGN U7581 ( .B(clk), .A(\g.we_clk [8809]));
Q_ASSIGN U7582 ( .B(clk), .A(\g.we_clk [8808]));
Q_ASSIGN U7583 ( .B(clk), .A(\g.we_clk [8807]));
Q_ASSIGN U7584 ( .B(clk), .A(\g.we_clk [8806]));
Q_ASSIGN U7585 ( .B(clk), .A(\g.we_clk [8805]));
Q_ASSIGN U7586 ( .B(clk), .A(\g.we_clk [8804]));
Q_ASSIGN U7587 ( .B(clk), .A(\g.we_clk [8803]));
Q_ASSIGN U7588 ( .B(clk), .A(\g.we_clk [8802]));
Q_ASSIGN U7589 ( .B(clk), .A(\g.we_clk [8801]));
Q_ASSIGN U7590 ( .B(clk), .A(\g.we_clk [8800]));
Q_ASSIGN U7591 ( .B(clk), .A(\g.we_clk [8799]));
Q_ASSIGN U7592 ( .B(clk), .A(\g.we_clk [8798]));
Q_ASSIGN U7593 ( .B(clk), .A(\g.we_clk [8797]));
Q_ASSIGN U7594 ( .B(clk), .A(\g.we_clk [8796]));
Q_ASSIGN U7595 ( .B(clk), .A(\g.we_clk [8795]));
Q_ASSIGN U7596 ( .B(clk), .A(\g.we_clk [8794]));
Q_ASSIGN U7597 ( .B(clk), .A(\g.we_clk [8793]));
Q_ASSIGN U7598 ( .B(clk), .A(\g.we_clk [8792]));
Q_ASSIGN U7599 ( .B(clk), .A(\g.we_clk [8791]));
Q_ASSIGN U7600 ( .B(clk), .A(\g.we_clk [8790]));
Q_ASSIGN U7601 ( .B(clk), .A(\g.we_clk [8789]));
Q_ASSIGN U7602 ( .B(clk), .A(\g.we_clk [8788]));
Q_ASSIGN U7603 ( .B(clk), .A(\g.we_clk [8787]));
Q_ASSIGN U7604 ( .B(clk), .A(\g.we_clk [8786]));
Q_ASSIGN U7605 ( .B(clk), .A(\g.we_clk [8785]));
Q_ASSIGN U7606 ( .B(clk), .A(\g.we_clk [8784]));
Q_ASSIGN U7607 ( .B(clk), .A(\g.we_clk [8783]));
Q_ASSIGN U7608 ( .B(clk), .A(\g.we_clk [8782]));
Q_ASSIGN U7609 ( .B(clk), .A(\g.we_clk [8781]));
Q_ASSIGN U7610 ( .B(clk), .A(\g.we_clk [8780]));
Q_ASSIGN U7611 ( .B(clk), .A(\g.we_clk [8779]));
Q_ASSIGN U7612 ( .B(clk), .A(\g.we_clk [8778]));
Q_ASSIGN U7613 ( .B(clk), .A(\g.we_clk [8777]));
Q_ASSIGN U7614 ( .B(clk), .A(\g.we_clk [8776]));
Q_ASSIGN U7615 ( .B(clk), .A(\g.we_clk [8775]));
Q_ASSIGN U7616 ( .B(clk), .A(\g.we_clk [8774]));
Q_ASSIGN U7617 ( .B(clk), .A(\g.we_clk [8773]));
Q_ASSIGN U7618 ( .B(clk), .A(\g.we_clk [8772]));
Q_ASSIGN U7619 ( .B(clk), .A(\g.we_clk [8771]));
Q_ASSIGN U7620 ( .B(clk), .A(\g.we_clk [8770]));
Q_ASSIGN U7621 ( .B(clk), .A(\g.we_clk [8769]));
Q_ASSIGN U7622 ( .B(clk), .A(\g.we_clk [8768]));
Q_ASSIGN U7623 ( .B(clk), .A(\g.we_clk [8767]));
Q_ASSIGN U7624 ( .B(clk), .A(\g.we_clk [8766]));
Q_ASSIGN U7625 ( .B(clk), .A(\g.we_clk [8765]));
Q_ASSIGN U7626 ( .B(clk), .A(\g.we_clk [8764]));
Q_ASSIGN U7627 ( .B(clk), .A(\g.we_clk [8763]));
Q_ASSIGN U7628 ( .B(clk), .A(\g.we_clk [8762]));
Q_ASSIGN U7629 ( .B(clk), .A(\g.we_clk [8761]));
Q_ASSIGN U7630 ( .B(clk), .A(\g.we_clk [8760]));
Q_ASSIGN U7631 ( .B(clk), .A(\g.we_clk [8759]));
Q_ASSIGN U7632 ( .B(clk), .A(\g.we_clk [8758]));
Q_ASSIGN U7633 ( .B(clk), .A(\g.we_clk [8757]));
Q_ASSIGN U7634 ( .B(clk), .A(\g.we_clk [8756]));
Q_ASSIGN U7635 ( .B(clk), .A(\g.we_clk [8755]));
Q_ASSIGN U7636 ( .B(clk), .A(\g.we_clk [8754]));
Q_ASSIGN U7637 ( .B(clk), .A(\g.we_clk [8753]));
Q_ASSIGN U7638 ( .B(clk), .A(\g.we_clk [8752]));
Q_ASSIGN U7639 ( .B(clk), .A(\g.we_clk [8751]));
Q_ASSIGN U7640 ( .B(clk), .A(\g.we_clk [8750]));
Q_ASSIGN U7641 ( .B(clk), .A(\g.we_clk [8749]));
Q_ASSIGN U7642 ( .B(clk), .A(\g.we_clk [8748]));
Q_ASSIGN U7643 ( .B(clk), .A(\g.we_clk [8747]));
Q_ASSIGN U7644 ( .B(clk), .A(\g.we_clk [8746]));
Q_ASSIGN U7645 ( .B(clk), .A(\g.we_clk [8745]));
Q_ASSIGN U7646 ( .B(clk), .A(\g.we_clk [8744]));
Q_ASSIGN U7647 ( .B(clk), .A(\g.we_clk [8743]));
Q_ASSIGN U7648 ( .B(clk), .A(\g.we_clk [8742]));
Q_ASSIGN U7649 ( .B(clk), .A(\g.we_clk [8741]));
Q_ASSIGN U7650 ( .B(clk), .A(\g.we_clk [8740]));
Q_ASSIGN U7651 ( .B(clk), .A(\g.we_clk [8739]));
Q_ASSIGN U7652 ( .B(clk), .A(\g.we_clk [8738]));
Q_ASSIGN U7653 ( .B(clk), .A(\g.we_clk [8737]));
Q_ASSIGN U7654 ( .B(clk), .A(\g.we_clk [8736]));
Q_ASSIGN U7655 ( .B(clk), .A(\g.we_clk [8735]));
Q_ASSIGN U7656 ( .B(clk), .A(\g.we_clk [8734]));
Q_ASSIGN U7657 ( .B(clk), .A(\g.we_clk [8733]));
Q_ASSIGN U7658 ( .B(clk), .A(\g.we_clk [8732]));
Q_ASSIGN U7659 ( .B(clk), .A(\g.we_clk [8731]));
Q_ASSIGN U7660 ( .B(clk), .A(\g.we_clk [8730]));
Q_ASSIGN U7661 ( .B(clk), .A(\g.we_clk [8729]));
Q_ASSIGN U7662 ( .B(clk), .A(\g.we_clk [8728]));
Q_ASSIGN U7663 ( .B(clk), .A(\g.we_clk [8727]));
Q_ASSIGN U7664 ( .B(clk), .A(\g.we_clk [8726]));
Q_ASSIGN U7665 ( .B(clk), .A(\g.we_clk [8725]));
Q_ASSIGN U7666 ( .B(clk), .A(\g.we_clk [8724]));
Q_ASSIGN U7667 ( .B(clk), .A(\g.we_clk [8723]));
Q_ASSIGN U7668 ( .B(clk), .A(\g.we_clk [8722]));
Q_ASSIGN U7669 ( .B(clk), .A(\g.we_clk [8721]));
Q_ASSIGN U7670 ( .B(clk), .A(\g.we_clk [8720]));
Q_ASSIGN U7671 ( .B(clk), .A(\g.we_clk [8719]));
Q_ASSIGN U7672 ( .B(clk), .A(\g.we_clk [8718]));
Q_ASSIGN U7673 ( .B(clk), .A(\g.we_clk [8717]));
Q_ASSIGN U7674 ( .B(clk), .A(\g.we_clk [8716]));
Q_ASSIGN U7675 ( .B(clk), .A(\g.we_clk [8715]));
Q_ASSIGN U7676 ( .B(clk), .A(\g.we_clk [8714]));
Q_ASSIGN U7677 ( .B(clk), .A(\g.we_clk [8713]));
Q_ASSIGN U7678 ( .B(clk), .A(\g.we_clk [8712]));
Q_ASSIGN U7679 ( .B(clk), .A(\g.we_clk [8711]));
Q_ASSIGN U7680 ( .B(clk), .A(\g.we_clk [8710]));
Q_ASSIGN U7681 ( .B(clk), .A(\g.we_clk [8709]));
Q_ASSIGN U7682 ( .B(clk), .A(\g.we_clk [8708]));
Q_ASSIGN U7683 ( .B(clk), .A(\g.we_clk [8707]));
Q_ASSIGN U7684 ( .B(clk), .A(\g.we_clk [8706]));
Q_ASSIGN U7685 ( .B(clk), .A(\g.we_clk [8705]));
Q_ASSIGN U7686 ( .B(clk), .A(\g.we_clk [8704]));
Q_ASSIGN U7687 ( .B(clk), .A(\g.we_clk [8703]));
Q_ASSIGN U7688 ( .B(clk), .A(\g.we_clk [8702]));
Q_ASSIGN U7689 ( .B(clk), .A(\g.we_clk [8701]));
Q_ASSIGN U7690 ( .B(clk), .A(\g.we_clk [8700]));
Q_ASSIGN U7691 ( .B(clk), .A(\g.we_clk [8699]));
Q_ASSIGN U7692 ( .B(clk), .A(\g.we_clk [8698]));
Q_ASSIGN U7693 ( .B(clk), .A(\g.we_clk [8697]));
Q_ASSIGN U7694 ( .B(clk), .A(\g.we_clk [8696]));
Q_ASSIGN U7695 ( .B(clk), .A(\g.we_clk [8695]));
Q_ASSIGN U7696 ( .B(clk), .A(\g.we_clk [8694]));
Q_ASSIGN U7697 ( .B(clk), .A(\g.we_clk [8693]));
Q_ASSIGN U7698 ( .B(clk), .A(\g.we_clk [8692]));
Q_ASSIGN U7699 ( .B(clk), .A(\g.we_clk [8691]));
Q_ASSIGN U7700 ( .B(clk), .A(\g.we_clk [8690]));
Q_ASSIGN U7701 ( .B(clk), .A(\g.we_clk [8689]));
Q_ASSIGN U7702 ( .B(clk), .A(\g.we_clk [8688]));
Q_ASSIGN U7703 ( .B(clk), .A(\g.we_clk [8687]));
Q_ASSIGN U7704 ( .B(clk), .A(\g.we_clk [8686]));
Q_ASSIGN U7705 ( .B(clk), .A(\g.we_clk [8685]));
Q_ASSIGN U7706 ( .B(clk), .A(\g.we_clk [8684]));
Q_ASSIGN U7707 ( .B(clk), .A(\g.we_clk [8683]));
Q_ASSIGN U7708 ( .B(clk), .A(\g.we_clk [8682]));
Q_ASSIGN U7709 ( .B(clk), .A(\g.we_clk [8681]));
Q_ASSIGN U7710 ( .B(clk), .A(\g.we_clk [8680]));
Q_ASSIGN U7711 ( .B(clk), .A(\g.we_clk [8679]));
Q_ASSIGN U7712 ( .B(clk), .A(\g.we_clk [8678]));
Q_ASSIGN U7713 ( .B(clk), .A(\g.we_clk [8677]));
Q_ASSIGN U7714 ( .B(clk), .A(\g.we_clk [8676]));
Q_ASSIGN U7715 ( .B(clk), .A(\g.we_clk [8675]));
Q_ASSIGN U7716 ( .B(clk), .A(\g.we_clk [8674]));
Q_ASSIGN U7717 ( .B(clk), .A(\g.we_clk [8673]));
Q_ASSIGN U7718 ( .B(clk), .A(\g.we_clk [8672]));
Q_ASSIGN U7719 ( .B(clk), .A(\g.we_clk [8671]));
Q_ASSIGN U7720 ( .B(clk), .A(\g.we_clk [8670]));
Q_ASSIGN U7721 ( .B(clk), .A(\g.we_clk [8669]));
Q_ASSIGN U7722 ( .B(clk), .A(\g.we_clk [8668]));
Q_ASSIGN U7723 ( .B(clk), .A(\g.we_clk [8667]));
Q_ASSIGN U7724 ( .B(clk), .A(\g.we_clk [8666]));
Q_ASSIGN U7725 ( .B(clk), .A(\g.we_clk [8665]));
Q_ASSIGN U7726 ( .B(clk), .A(\g.we_clk [8664]));
Q_ASSIGN U7727 ( .B(clk), .A(\g.we_clk [8663]));
Q_ASSIGN U7728 ( .B(clk), .A(\g.we_clk [8662]));
Q_ASSIGN U7729 ( .B(clk), .A(\g.we_clk [8661]));
Q_ASSIGN U7730 ( .B(clk), .A(\g.we_clk [8660]));
Q_ASSIGN U7731 ( .B(clk), .A(\g.we_clk [8659]));
Q_ASSIGN U7732 ( .B(clk), .A(\g.we_clk [8658]));
Q_ASSIGN U7733 ( .B(clk), .A(\g.we_clk [8657]));
Q_ASSIGN U7734 ( .B(clk), .A(\g.we_clk [8656]));
Q_ASSIGN U7735 ( .B(clk), .A(\g.we_clk [8655]));
Q_ASSIGN U7736 ( .B(clk), .A(\g.we_clk [8654]));
Q_ASSIGN U7737 ( .B(clk), .A(\g.we_clk [8653]));
Q_ASSIGN U7738 ( .B(clk), .A(\g.we_clk [8652]));
Q_ASSIGN U7739 ( .B(clk), .A(\g.we_clk [8651]));
Q_ASSIGN U7740 ( .B(clk), .A(\g.we_clk [8650]));
Q_ASSIGN U7741 ( .B(clk), .A(\g.we_clk [8649]));
Q_ASSIGN U7742 ( .B(clk), .A(\g.we_clk [8648]));
Q_ASSIGN U7743 ( .B(clk), .A(\g.we_clk [8647]));
Q_ASSIGN U7744 ( .B(clk), .A(\g.we_clk [8646]));
Q_ASSIGN U7745 ( .B(clk), .A(\g.we_clk [8645]));
Q_ASSIGN U7746 ( .B(clk), .A(\g.we_clk [8644]));
Q_ASSIGN U7747 ( .B(clk), .A(\g.we_clk [8643]));
Q_ASSIGN U7748 ( .B(clk), .A(\g.we_clk [8642]));
Q_ASSIGN U7749 ( .B(clk), .A(\g.we_clk [8641]));
Q_ASSIGN U7750 ( .B(clk), .A(\g.we_clk [8640]));
Q_ASSIGN U7751 ( .B(clk), .A(\g.we_clk [8639]));
Q_ASSIGN U7752 ( .B(clk), .A(\g.we_clk [8638]));
Q_ASSIGN U7753 ( .B(clk), .A(\g.we_clk [8637]));
Q_ASSIGN U7754 ( .B(clk), .A(\g.we_clk [8636]));
Q_ASSIGN U7755 ( .B(clk), .A(\g.we_clk [8635]));
Q_ASSIGN U7756 ( .B(clk), .A(\g.we_clk [8634]));
Q_ASSIGN U7757 ( .B(clk), .A(\g.we_clk [8633]));
Q_ASSIGN U7758 ( .B(clk), .A(\g.we_clk [8632]));
Q_ASSIGN U7759 ( .B(clk), .A(\g.we_clk [8631]));
Q_ASSIGN U7760 ( .B(clk), .A(\g.we_clk [8630]));
Q_ASSIGN U7761 ( .B(clk), .A(\g.we_clk [8629]));
Q_ASSIGN U7762 ( .B(clk), .A(\g.we_clk [8628]));
Q_ASSIGN U7763 ( .B(clk), .A(\g.we_clk [8627]));
Q_ASSIGN U7764 ( .B(clk), .A(\g.we_clk [8626]));
Q_ASSIGN U7765 ( .B(clk), .A(\g.we_clk [8625]));
Q_ASSIGN U7766 ( .B(clk), .A(\g.we_clk [8624]));
Q_ASSIGN U7767 ( .B(clk), .A(\g.we_clk [8623]));
Q_ASSIGN U7768 ( .B(clk), .A(\g.we_clk [8622]));
Q_ASSIGN U7769 ( .B(clk), .A(\g.we_clk [8621]));
Q_ASSIGN U7770 ( .B(clk), .A(\g.we_clk [8620]));
Q_ASSIGN U7771 ( .B(clk), .A(\g.we_clk [8619]));
Q_ASSIGN U7772 ( .B(clk), .A(\g.we_clk [8618]));
Q_ASSIGN U7773 ( .B(clk), .A(\g.we_clk [8617]));
Q_ASSIGN U7774 ( .B(clk), .A(\g.we_clk [8616]));
Q_ASSIGN U7775 ( .B(clk), .A(\g.we_clk [8615]));
Q_ASSIGN U7776 ( .B(clk), .A(\g.we_clk [8614]));
Q_ASSIGN U7777 ( .B(clk), .A(\g.we_clk [8613]));
Q_ASSIGN U7778 ( .B(clk), .A(\g.we_clk [8612]));
Q_ASSIGN U7779 ( .B(clk), .A(\g.we_clk [8611]));
Q_ASSIGN U7780 ( .B(clk), .A(\g.we_clk [8610]));
Q_ASSIGN U7781 ( .B(clk), .A(\g.we_clk [8609]));
Q_ASSIGN U7782 ( .B(clk), .A(\g.we_clk [8608]));
Q_ASSIGN U7783 ( .B(clk), .A(\g.we_clk [8607]));
Q_ASSIGN U7784 ( .B(clk), .A(\g.we_clk [8606]));
Q_ASSIGN U7785 ( .B(clk), .A(\g.we_clk [8605]));
Q_ASSIGN U7786 ( .B(clk), .A(\g.we_clk [8604]));
Q_ASSIGN U7787 ( .B(clk), .A(\g.we_clk [8603]));
Q_ASSIGN U7788 ( .B(clk), .A(\g.we_clk [8602]));
Q_ASSIGN U7789 ( .B(clk), .A(\g.we_clk [8601]));
Q_ASSIGN U7790 ( .B(clk), .A(\g.we_clk [8600]));
Q_ASSIGN U7791 ( .B(clk), .A(\g.we_clk [8599]));
Q_ASSIGN U7792 ( .B(clk), .A(\g.we_clk [8598]));
Q_ASSIGN U7793 ( .B(clk), .A(\g.we_clk [8597]));
Q_ASSIGN U7794 ( .B(clk), .A(\g.we_clk [8596]));
Q_ASSIGN U7795 ( .B(clk), .A(\g.we_clk [8595]));
Q_ASSIGN U7796 ( .B(clk), .A(\g.we_clk [8594]));
Q_ASSIGN U7797 ( .B(clk), .A(\g.we_clk [8593]));
Q_ASSIGN U7798 ( .B(clk), .A(\g.we_clk [8592]));
Q_ASSIGN U7799 ( .B(clk), .A(\g.we_clk [8591]));
Q_ASSIGN U7800 ( .B(clk), .A(\g.we_clk [8590]));
Q_ASSIGN U7801 ( .B(clk), .A(\g.we_clk [8589]));
Q_ASSIGN U7802 ( .B(clk), .A(\g.we_clk [8588]));
Q_ASSIGN U7803 ( .B(clk), .A(\g.we_clk [8587]));
Q_ASSIGN U7804 ( .B(clk), .A(\g.we_clk [8586]));
Q_ASSIGN U7805 ( .B(clk), .A(\g.we_clk [8585]));
Q_ASSIGN U7806 ( .B(clk), .A(\g.we_clk [8584]));
Q_ASSIGN U7807 ( .B(clk), .A(\g.we_clk [8583]));
Q_ASSIGN U7808 ( .B(clk), .A(\g.we_clk [8582]));
Q_ASSIGN U7809 ( .B(clk), .A(\g.we_clk [8581]));
Q_ASSIGN U7810 ( .B(clk), .A(\g.we_clk [8580]));
Q_ASSIGN U7811 ( .B(clk), .A(\g.we_clk [8579]));
Q_ASSIGN U7812 ( .B(clk), .A(\g.we_clk [8578]));
Q_ASSIGN U7813 ( .B(clk), .A(\g.we_clk [8577]));
Q_ASSIGN U7814 ( .B(clk), .A(\g.we_clk [8576]));
Q_ASSIGN U7815 ( .B(clk), .A(\g.we_clk [8575]));
Q_ASSIGN U7816 ( .B(clk), .A(\g.we_clk [8574]));
Q_ASSIGN U7817 ( .B(clk), .A(\g.we_clk [8573]));
Q_ASSIGN U7818 ( .B(clk), .A(\g.we_clk [8572]));
Q_ASSIGN U7819 ( .B(clk), .A(\g.we_clk [8571]));
Q_ASSIGN U7820 ( .B(clk), .A(\g.we_clk [8570]));
Q_ASSIGN U7821 ( .B(clk), .A(\g.we_clk [8569]));
Q_ASSIGN U7822 ( .B(clk), .A(\g.we_clk [8568]));
Q_ASSIGN U7823 ( .B(clk), .A(\g.we_clk [8567]));
Q_ASSIGN U7824 ( .B(clk), .A(\g.we_clk [8566]));
Q_ASSIGN U7825 ( .B(clk), .A(\g.we_clk [8565]));
Q_ASSIGN U7826 ( .B(clk), .A(\g.we_clk [8564]));
Q_ASSIGN U7827 ( .B(clk), .A(\g.we_clk [8563]));
Q_ASSIGN U7828 ( .B(clk), .A(\g.we_clk [8562]));
Q_ASSIGN U7829 ( .B(clk), .A(\g.we_clk [8561]));
Q_ASSIGN U7830 ( .B(clk), .A(\g.we_clk [8560]));
Q_ASSIGN U7831 ( .B(clk), .A(\g.we_clk [8559]));
Q_ASSIGN U7832 ( .B(clk), .A(\g.we_clk [8558]));
Q_ASSIGN U7833 ( .B(clk), .A(\g.we_clk [8557]));
Q_ASSIGN U7834 ( .B(clk), .A(\g.we_clk [8556]));
Q_ASSIGN U7835 ( .B(clk), .A(\g.we_clk [8555]));
Q_ASSIGN U7836 ( .B(clk), .A(\g.we_clk [8554]));
Q_ASSIGN U7837 ( .B(clk), .A(\g.we_clk [8553]));
Q_ASSIGN U7838 ( .B(clk), .A(\g.we_clk [8552]));
Q_ASSIGN U7839 ( .B(clk), .A(\g.we_clk [8551]));
Q_ASSIGN U7840 ( .B(clk), .A(\g.we_clk [8550]));
Q_ASSIGN U7841 ( .B(clk), .A(\g.we_clk [8549]));
Q_ASSIGN U7842 ( .B(clk), .A(\g.we_clk [8548]));
Q_ASSIGN U7843 ( .B(clk), .A(\g.we_clk [8547]));
Q_ASSIGN U7844 ( .B(clk), .A(\g.we_clk [8546]));
Q_ASSIGN U7845 ( .B(clk), .A(\g.we_clk [8545]));
Q_ASSIGN U7846 ( .B(clk), .A(\g.we_clk [8544]));
Q_ASSIGN U7847 ( .B(clk), .A(\g.we_clk [8543]));
Q_ASSIGN U7848 ( .B(clk), .A(\g.we_clk [8542]));
Q_ASSIGN U7849 ( .B(clk), .A(\g.we_clk [8541]));
Q_ASSIGN U7850 ( .B(clk), .A(\g.we_clk [8540]));
Q_ASSIGN U7851 ( .B(clk), .A(\g.we_clk [8539]));
Q_ASSIGN U7852 ( .B(clk), .A(\g.we_clk [8538]));
Q_ASSIGN U7853 ( .B(clk), .A(\g.we_clk [8537]));
Q_ASSIGN U7854 ( .B(clk), .A(\g.we_clk [8536]));
Q_ASSIGN U7855 ( .B(clk), .A(\g.we_clk [8535]));
Q_ASSIGN U7856 ( .B(clk), .A(\g.we_clk [8534]));
Q_ASSIGN U7857 ( .B(clk), .A(\g.we_clk [8533]));
Q_ASSIGN U7858 ( .B(clk), .A(\g.we_clk [8532]));
Q_ASSIGN U7859 ( .B(clk), .A(\g.we_clk [8531]));
Q_ASSIGN U7860 ( .B(clk), .A(\g.we_clk [8530]));
Q_ASSIGN U7861 ( .B(clk), .A(\g.we_clk [8529]));
Q_ASSIGN U7862 ( .B(clk), .A(\g.we_clk [8528]));
Q_ASSIGN U7863 ( .B(clk), .A(\g.we_clk [8527]));
Q_ASSIGN U7864 ( .B(clk), .A(\g.we_clk [8526]));
Q_ASSIGN U7865 ( .B(clk), .A(\g.we_clk [8525]));
Q_ASSIGN U7866 ( .B(clk), .A(\g.we_clk [8524]));
Q_ASSIGN U7867 ( .B(clk), .A(\g.we_clk [8523]));
Q_ASSIGN U7868 ( .B(clk), .A(\g.we_clk [8522]));
Q_ASSIGN U7869 ( .B(clk), .A(\g.we_clk [8521]));
Q_ASSIGN U7870 ( .B(clk), .A(\g.we_clk [8520]));
Q_ASSIGN U7871 ( .B(clk), .A(\g.we_clk [8519]));
Q_ASSIGN U7872 ( .B(clk), .A(\g.we_clk [8518]));
Q_ASSIGN U7873 ( .B(clk), .A(\g.we_clk [8517]));
Q_ASSIGN U7874 ( .B(clk), .A(\g.we_clk [8516]));
Q_ASSIGN U7875 ( .B(clk), .A(\g.we_clk [8515]));
Q_ASSIGN U7876 ( .B(clk), .A(\g.we_clk [8514]));
Q_ASSIGN U7877 ( .B(clk), .A(\g.we_clk [8513]));
Q_ASSIGN U7878 ( .B(clk), .A(\g.we_clk [8512]));
Q_ASSIGN U7879 ( .B(clk), .A(\g.we_clk [8511]));
Q_ASSIGN U7880 ( .B(clk), .A(\g.we_clk [8510]));
Q_ASSIGN U7881 ( .B(clk), .A(\g.we_clk [8509]));
Q_ASSIGN U7882 ( .B(clk), .A(\g.we_clk [8508]));
Q_ASSIGN U7883 ( .B(clk), .A(\g.we_clk [8507]));
Q_ASSIGN U7884 ( .B(clk), .A(\g.we_clk [8506]));
Q_ASSIGN U7885 ( .B(clk), .A(\g.we_clk [8505]));
Q_ASSIGN U7886 ( .B(clk), .A(\g.we_clk [8504]));
Q_ASSIGN U7887 ( .B(clk), .A(\g.we_clk [8503]));
Q_ASSIGN U7888 ( .B(clk), .A(\g.we_clk [8502]));
Q_ASSIGN U7889 ( .B(clk), .A(\g.we_clk [8501]));
Q_ASSIGN U7890 ( .B(clk), .A(\g.we_clk [8500]));
Q_ASSIGN U7891 ( .B(clk), .A(\g.we_clk [8499]));
Q_ASSIGN U7892 ( .B(clk), .A(\g.we_clk [8498]));
Q_ASSIGN U7893 ( .B(clk), .A(\g.we_clk [8497]));
Q_ASSIGN U7894 ( .B(clk), .A(\g.we_clk [8496]));
Q_ASSIGN U7895 ( .B(clk), .A(\g.we_clk [8495]));
Q_ASSIGN U7896 ( .B(clk), .A(\g.we_clk [8494]));
Q_ASSIGN U7897 ( .B(clk), .A(\g.we_clk [8493]));
Q_ASSIGN U7898 ( .B(clk), .A(\g.we_clk [8492]));
Q_ASSIGN U7899 ( .B(clk), .A(\g.we_clk [8491]));
Q_ASSIGN U7900 ( .B(clk), .A(\g.we_clk [8490]));
Q_ASSIGN U7901 ( .B(clk), .A(\g.we_clk [8489]));
Q_ASSIGN U7902 ( .B(clk), .A(\g.we_clk [8488]));
Q_ASSIGN U7903 ( .B(clk), .A(\g.we_clk [8487]));
Q_ASSIGN U7904 ( .B(clk), .A(\g.we_clk [8486]));
Q_ASSIGN U7905 ( .B(clk), .A(\g.we_clk [8485]));
Q_ASSIGN U7906 ( .B(clk), .A(\g.we_clk [8484]));
Q_ASSIGN U7907 ( .B(clk), .A(\g.we_clk [8483]));
Q_ASSIGN U7908 ( .B(clk), .A(\g.we_clk [8482]));
Q_ASSIGN U7909 ( .B(clk), .A(\g.we_clk [8481]));
Q_ASSIGN U7910 ( .B(clk), .A(\g.we_clk [8480]));
Q_ASSIGN U7911 ( .B(clk), .A(\g.we_clk [8479]));
Q_ASSIGN U7912 ( .B(clk), .A(\g.we_clk [8478]));
Q_ASSIGN U7913 ( .B(clk), .A(\g.we_clk [8477]));
Q_ASSIGN U7914 ( .B(clk), .A(\g.we_clk [8476]));
Q_ASSIGN U7915 ( .B(clk), .A(\g.we_clk [8475]));
Q_ASSIGN U7916 ( .B(clk), .A(\g.we_clk [8474]));
Q_ASSIGN U7917 ( .B(clk), .A(\g.we_clk [8473]));
Q_ASSIGN U7918 ( .B(clk), .A(\g.we_clk [8472]));
Q_ASSIGN U7919 ( .B(clk), .A(\g.we_clk [8471]));
Q_ASSIGN U7920 ( .B(clk), .A(\g.we_clk [8470]));
Q_ASSIGN U7921 ( .B(clk), .A(\g.we_clk [8469]));
Q_ASSIGN U7922 ( .B(clk), .A(\g.we_clk [8468]));
Q_ASSIGN U7923 ( .B(clk), .A(\g.we_clk [8467]));
Q_ASSIGN U7924 ( .B(clk), .A(\g.we_clk [8466]));
Q_ASSIGN U7925 ( .B(clk), .A(\g.we_clk [8465]));
Q_ASSIGN U7926 ( .B(clk), .A(\g.we_clk [8464]));
Q_ASSIGN U7927 ( .B(clk), .A(\g.we_clk [8463]));
Q_ASSIGN U7928 ( .B(clk), .A(\g.we_clk [8462]));
Q_ASSIGN U7929 ( .B(clk), .A(\g.we_clk [8461]));
Q_ASSIGN U7930 ( .B(clk), .A(\g.we_clk [8460]));
Q_ASSIGN U7931 ( .B(clk), .A(\g.we_clk [8459]));
Q_ASSIGN U7932 ( .B(clk), .A(\g.we_clk [8458]));
Q_ASSIGN U7933 ( .B(clk), .A(\g.we_clk [8457]));
Q_ASSIGN U7934 ( .B(clk), .A(\g.we_clk [8456]));
Q_ASSIGN U7935 ( .B(clk), .A(\g.we_clk [8455]));
Q_ASSIGN U7936 ( .B(clk), .A(\g.we_clk [8454]));
Q_ASSIGN U7937 ( .B(clk), .A(\g.we_clk [8453]));
Q_ASSIGN U7938 ( .B(clk), .A(\g.we_clk [8452]));
Q_ASSIGN U7939 ( .B(clk), .A(\g.we_clk [8451]));
Q_ASSIGN U7940 ( .B(clk), .A(\g.we_clk [8450]));
Q_ASSIGN U7941 ( .B(clk), .A(\g.we_clk [8449]));
Q_ASSIGN U7942 ( .B(clk), .A(\g.we_clk [8448]));
Q_ASSIGN U7943 ( .B(clk), .A(\g.we_clk [8447]));
Q_ASSIGN U7944 ( .B(clk), .A(\g.we_clk [8446]));
Q_ASSIGN U7945 ( .B(clk), .A(\g.we_clk [8445]));
Q_ASSIGN U7946 ( .B(clk), .A(\g.we_clk [8444]));
Q_ASSIGN U7947 ( .B(clk), .A(\g.we_clk [8443]));
Q_ASSIGN U7948 ( .B(clk), .A(\g.we_clk [8442]));
Q_ASSIGN U7949 ( .B(clk), .A(\g.we_clk [8441]));
Q_ASSIGN U7950 ( .B(clk), .A(\g.we_clk [8440]));
Q_ASSIGN U7951 ( .B(clk), .A(\g.we_clk [8439]));
Q_ASSIGN U7952 ( .B(clk), .A(\g.we_clk [8438]));
Q_ASSIGN U7953 ( .B(clk), .A(\g.we_clk [8437]));
Q_ASSIGN U7954 ( .B(clk), .A(\g.we_clk [8436]));
Q_ASSIGN U7955 ( .B(clk), .A(\g.we_clk [8435]));
Q_ASSIGN U7956 ( .B(clk), .A(\g.we_clk [8434]));
Q_ASSIGN U7957 ( .B(clk), .A(\g.we_clk [8433]));
Q_ASSIGN U7958 ( .B(clk), .A(\g.we_clk [8432]));
Q_ASSIGN U7959 ( .B(clk), .A(\g.we_clk [8431]));
Q_ASSIGN U7960 ( .B(clk), .A(\g.we_clk [8430]));
Q_ASSIGN U7961 ( .B(clk), .A(\g.we_clk [8429]));
Q_ASSIGN U7962 ( .B(clk), .A(\g.we_clk [8428]));
Q_ASSIGN U7963 ( .B(clk), .A(\g.we_clk [8427]));
Q_ASSIGN U7964 ( .B(clk), .A(\g.we_clk [8426]));
Q_ASSIGN U7965 ( .B(clk), .A(\g.we_clk [8425]));
Q_ASSIGN U7966 ( .B(clk), .A(\g.we_clk [8424]));
Q_ASSIGN U7967 ( .B(clk), .A(\g.we_clk [8423]));
Q_ASSIGN U7968 ( .B(clk), .A(\g.we_clk [8422]));
Q_ASSIGN U7969 ( .B(clk), .A(\g.we_clk [8421]));
Q_ASSIGN U7970 ( .B(clk), .A(\g.we_clk [8420]));
Q_ASSIGN U7971 ( .B(clk), .A(\g.we_clk [8419]));
Q_ASSIGN U7972 ( .B(clk), .A(\g.we_clk [8418]));
Q_ASSIGN U7973 ( .B(clk), .A(\g.we_clk [8417]));
Q_ASSIGN U7974 ( .B(clk), .A(\g.we_clk [8416]));
Q_ASSIGN U7975 ( .B(clk), .A(\g.we_clk [8415]));
Q_ASSIGN U7976 ( .B(clk), .A(\g.we_clk [8414]));
Q_ASSIGN U7977 ( .B(clk), .A(\g.we_clk [8413]));
Q_ASSIGN U7978 ( .B(clk), .A(\g.we_clk [8412]));
Q_ASSIGN U7979 ( .B(clk), .A(\g.we_clk [8411]));
Q_ASSIGN U7980 ( .B(clk), .A(\g.we_clk [8410]));
Q_ASSIGN U7981 ( .B(clk), .A(\g.we_clk [8409]));
Q_ASSIGN U7982 ( .B(clk), .A(\g.we_clk [8408]));
Q_ASSIGN U7983 ( .B(clk), .A(\g.we_clk [8407]));
Q_ASSIGN U7984 ( .B(clk), .A(\g.we_clk [8406]));
Q_ASSIGN U7985 ( .B(clk), .A(\g.we_clk [8405]));
Q_ASSIGN U7986 ( .B(clk), .A(\g.we_clk [8404]));
Q_ASSIGN U7987 ( .B(clk), .A(\g.we_clk [8403]));
Q_ASSIGN U7988 ( .B(clk), .A(\g.we_clk [8402]));
Q_ASSIGN U7989 ( .B(clk), .A(\g.we_clk [8401]));
Q_ASSIGN U7990 ( .B(clk), .A(\g.we_clk [8400]));
Q_ASSIGN U7991 ( .B(clk), .A(\g.we_clk [8399]));
Q_ASSIGN U7992 ( .B(clk), .A(\g.we_clk [8398]));
Q_ASSIGN U7993 ( .B(clk), .A(\g.we_clk [8397]));
Q_ASSIGN U7994 ( .B(clk), .A(\g.we_clk [8396]));
Q_ASSIGN U7995 ( .B(clk), .A(\g.we_clk [8395]));
Q_ASSIGN U7996 ( .B(clk), .A(\g.we_clk [8394]));
Q_ASSIGN U7997 ( .B(clk), .A(\g.we_clk [8393]));
Q_ASSIGN U7998 ( .B(clk), .A(\g.we_clk [8392]));
Q_ASSIGN U7999 ( .B(clk), .A(\g.we_clk [8391]));
Q_ASSIGN U8000 ( .B(clk), .A(\g.we_clk [8390]));
Q_ASSIGN U8001 ( .B(clk), .A(\g.we_clk [8389]));
Q_ASSIGN U8002 ( .B(clk), .A(\g.we_clk [8388]));
Q_ASSIGN U8003 ( .B(clk), .A(\g.we_clk [8387]));
Q_ASSIGN U8004 ( .B(clk), .A(\g.we_clk [8386]));
Q_ASSIGN U8005 ( .B(clk), .A(\g.we_clk [8385]));
Q_ASSIGN U8006 ( .B(clk), .A(\g.we_clk [8384]));
Q_ASSIGN U8007 ( .B(clk), .A(\g.we_clk [8383]));
Q_ASSIGN U8008 ( .B(clk), .A(\g.we_clk [8382]));
Q_ASSIGN U8009 ( .B(clk), .A(\g.we_clk [8381]));
Q_ASSIGN U8010 ( .B(clk), .A(\g.we_clk [8380]));
Q_ASSIGN U8011 ( .B(clk), .A(\g.we_clk [8379]));
Q_ASSIGN U8012 ( .B(clk), .A(\g.we_clk [8378]));
Q_ASSIGN U8013 ( .B(clk), .A(\g.we_clk [8377]));
Q_ASSIGN U8014 ( .B(clk), .A(\g.we_clk [8376]));
Q_ASSIGN U8015 ( .B(clk), .A(\g.we_clk [8375]));
Q_ASSIGN U8016 ( .B(clk), .A(\g.we_clk [8374]));
Q_ASSIGN U8017 ( .B(clk), .A(\g.we_clk [8373]));
Q_ASSIGN U8018 ( .B(clk), .A(\g.we_clk [8372]));
Q_ASSIGN U8019 ( .B(clk), .A(\g.we_clk [8371]));
Q_ASSIGN U8020 ( .B(clk), .A(\g.we_clk [8370]));
Q_ASSIGN U8021 ( .B(clk), .A(\g.we_clk [8369]));
Q_ASSIGN U8022 ( .B(clk), .A(\g.we_clk [8368]));
Q_ASSIGN U8023 ( .B(clk), .A(\g.we_clk [8367]));
Q_ASSIGN U8024 ( .B(clk), .A(\g.we_clk [8366]));
Q_ASSIGN U8025 ( .B(clk), .A(\g.we_clk [8365]));
Q_ASSIGN U8026 ( .B(clk), .A(\g.we_clk [8364]));
Q_ASSIGN U8027 ( .B(clk), .A(\g.we_clk [8363]));
Q_ASSIGN U8028 ( .B(clk), .A(\g.we_clk [8362]));
Q_ASSIGN U8029 ( .B(clk), .A(\g.we_clk [8361]));
Q_ASSIGN U8030 ( .B(clk), .A(\g.we_clk [8360]));
Q_ASSIGN U8031 ( .B(clk), .A(\g.we_clk [8359]));
Q_ASSIGN U8032 ( .B(clk), .A(\g.we_clk [8358]));
Q_ASSIGN U8033 ( .B(clk), .A(\g.we_clk [8357]));
Q_ASSIGN U8034 ( .B(clk), .A(\g.we_clk [8356]));
Q_ASSIGN U8035 ( .B(clk), .A(\g.we_clk [8355]));
Q_ASSIGN U8036 ( .B(clk), .A(\g.we_clk [8354]));
Q_ASSIGN U8037 ( .B(clk), .A(\g.we_clk [8353]));
Q_ASSIGN U8038 ( .B(clk), .A(\g.we_clk [8352]));
Q_ASSIGN U8039 ( .B(clk), .A(\g.we_clk [8351]));
Q_ASSIGN U8040 ( .B(clk), .A(\g.we_clk [8350]));
Q_ASSIGN U8041 ( .B(clk), .A(\g.we_clk [8349]));
Q_ASSIGN U8042 ( .B(clk), .A(\g.we_clk [8348]));
Q_ASSIGN U8043 ( .B(clk), .A(\g.we_clk [8347]));
Q_ASSIGN U8044 ( .B(clk), .A(\g.we_clk [8346]));
Q_ASSIGN U8045 ( .B(clk), .A(\g.we_clk [8345]));
Q_ASSIGN U8046 ( .B(clk), .A(\g.we_clk [8344]));
Q_ASSIGN U8047 ( .B(clk), .A(\g.we_clk [8343]));
Q_ASSIGN U8048 ( .B(clk), .A(\g.we_clk [8342]));
Q_ASSIGN U8049 ( .B(clk), .A(\g.we_clk [8341]));
Q_ASSIGN U8050 ( .B(clk), .A(\g.we_clk [8340]));
Q_ASSIGN U8051 ( .B(clk), .A(\g.we_clk [8339]));
Q_ASSIGN U8052 ( .B(clk), .A(\g.we_clk [8338]));
Q_ASSIGN U8053 ( .B(clk), .A(\g.we_clk [8337]));
Q_ASSIGN U8054 ( .B(clk), .A(\g.we_clk [8336]));
Q_ASSIGN U8055 ( .B(clk), .A(\g.we_clk [8335]));
Q_ASSIGN U8056 ( .B(clk), .A(\g.we_clk [8334]));
Q_ASSIGN U8057 ( .B(clk), .A(\g.we_clk [8333]));
Q_ASSIGN U8058 ( .B(clk), .A(\g.we_clk [8332]));
Q_ASSIGN U8059 ( .B(clk), .A(\g.we_clk [8331]));
Q_ASSIGN U8060 ( .B(clk), .A(\g.we_clk [8330]));
Q_ASSIGN U8061 ( .B(clk), .A(\g.we_clk [8329]));
Q_ASSIGN U8062 ( .B(clk), .A(\g.we_clk [8328]));
Q_ASSIGN U8063 ( .B(clk), .A(\g.we_clk [8327]));
Q_ASSIGN U8064 ( .B(clk), .A(\g.we_clk [8326]));
Q_ASSIGN U8065 ( .B(clk), .A(\g.we_clk [8325]));
Q_ASSIGN U8066 ( .B(clk), .A(\g.we_clk [8324]));
Q_ASSIGN U8067 ( .B(clk), .A(\g.we_clk [8323]));
Q_ASSIGN U8068 ( .B(clk), .A(\g.we_clk [8322]));
Q_ASSIGN U8069 ( .B(clk), .A(\g.we_clk [8321]));
Q_ASSIGN U8070 ( .B(clk), .A(\g.we_clk [8320]));
Q_ASSIGN U8071 ( .B(clk), .A(\g.we_clk [8319]));
Q_ASSIGN U8072 ( .B(clk), .A(\g.we_clk [8318]));
Q_ASSIGN U8073 ( .B(clk), .A(\g.we_clk [8317]));
Q_ASSIGN U8074 ( .B(clk), .A(\g.we_clk [8316]));
Q_ASSIGN U8075 ( .B(clk), .A(\g.we_clk [8315]));
Q_ASSIGN U8076 ( .B(clk), .A(\g.we_clk [8314]));
Q_ASSIGN U8077 ( .B(clk), .A(\g.we_clk [8313]));
Q_ASSIGN U8078 ( .B(clk), .A(\g.we_clk [8312]));
Q_ASSIGN U8079 ( .B(clk), .A(\g.we_clk [8311]));
Q_ASSIGN U8080 ( .B(clk), .A(\g.we_clk [8310]));
Q_ASSIGN U8081 ( .B(clk), .A(\g.we_clk [8309]));
Q_ASSIGN U8082 ( .B(clk), .A(\g.we_clk [8308]));
Q_ASSIGN U8083 ( .B(clk), .A(\g.we_clk [8307]));
Q_ASSIGN U8084 ( .B(clk), .A(\g.we_clk [8306]));
Q_ASSIGN U8085 ( .B(clk), .A(\g.we_clk [8305]));
Q_ASSIGN U8086 ( .B(clk), .A(\g.we_clk [8304]));
Q_ASSIGN U8087 ( .B(clk), .A(\g.we_clk [8303]));
Q_ASSIGN U8088 ( .B(clk), .A(\g.we_clk [8302]));
Q_ASSIGN U8089 ( .B(clk), .A(\g.we_clk [8301]));
Q_ASSIGN U8090 ( .B(clk), .A(\g.we_clk [8300]));
Q_ASSIGN U8091 ( .B(clk), .A(\g.we_clk [8299]));
Q_ASSIGN U8092 ( .B(clk), .A(\g.we_clk [8298]));
Q_ASSIGN U8093 ( .B(clk), .A(\g.we_clk [8297]));
Q_ASSIGN U8094 ( .B(clk), .A(\g.we_clk [8296]));
Q_ASSIGN U8095 ( .B(clk), .A(\g.we_clk [8295]));
Q_ASSIGN U8096 ( .B(clk), .A(\g.we_clk [8294]));
Q_ASSIGN U8097 ( .B(clk), .A(\g.we_clk [8293]));
Q_ASSIGN U8098 ( .B(clk), .A(\g.we_clk [8292]));
Q_ASSIGN U8099 ( .B(clk), .A(\g.we_clk [8291]));
Q_ASSIGN U8100 ( .B(clk), .A(\g.we_clk [8290]));
Q_ASSIGN U8101 ( .B(clk), .A(\g.we_clk [8289]));
Q_ASSIGN U8102 ( .B(clk), .A(\g.we_clk [8288]));
Q_ASSIGN U8103 ( .B(clk), .A(\g.we_clk [8287]));
Q_ASSIGN U8104 ( .B(clk), .A(\g.we_clk [8286]));
Q_ASSIGN U8105 ( .B(clk), .A(\g.we_clk [8285]));
Q_ASSIGN U8106 ( .B(clk), .A(\g.we_clk [8284]));
Q_ASSIGN U8107 ( .B(clk), .A(\g.we_clk [8283]));
Q_ASSIGN U8108 ( .B(clk), .A(\g.we_clk [8282]));
Q_ASSIGN U8109 ( .B(clk), .A(\g.we_clk [8281]));
Q_ASSIGN U8110 ( .B(clk), .A(\g.we_clk [8280]));
Q_ASSIGN U8111 ( .B(clk), .A(\g.we_clk [8279]));
Q_ASSIGN U8112 ( .B(clk), .A(\g.we_clk [8278]));
Q_ASSIGN U8113 ( .B(clk), .A(\g.we_clk [8277]));
Q_ASSIGN U8114 ( .B(clk), .A(\g.we_clk [8276]));
Q_ASSIGN U8115 ( .B(clk), .A(\g.we_clk [8275]));
Q_ASSIGN U8116 ( .B(clk), .A(\g.we_clk [8274]));
Q_ASSIGN U8117 ( .B(clk), .A(\g.we_clk [8273]));
Q_ASSIGN U8118 ( .B(clk), .A(\g.we_clk [8272]));
Q_ASSIGN U8119 ( .B(clk), .A(\g.we_clk [8271]));
Q_ASSIGN U8120 ( .B(clk), .A(\g.we_clk [8270]));
Q_ASSIGN U8121 ( .B(clk), .A(\g.we_clk [8269]));
Q_ASSIGN U8122 ( .B(clk), .A(\g.we_clk [8268]));
Q_ASSIGN U8123 ( .B(clk), .A(\g.we_clk [8267]));
Q_ASSIGN U8124 ( .B(clk), .A(\g.we_clk [8266]));
Q_ASSIGN U8125 ( .B(clk), .A(\g.we_clk [8265]));
Q_ASSIGN U8126 ( .B(clk), .A(\g.we_clk [8264]));
Q_ASSIGN U8127 ( .B(clk), .A(\g.we_clk [8263]));
Q_ASSIGN U8128 ( .B(clk), .A(\g.we_clk [8262]));
Q_ASSIGN U8129 ( .B(clk), .A(\g.we_clk [8261]));
Q_ASSIGN U8130 ( .B(clk), .A(\g.we_clk [8260]));
Q_ASSIGN U8131 ( .B(clk), .A(\g.we_clk [8259]));
Q_ASSIGN U8132 ( .B(clk), .A(\g.we_clk [8258]));
Q_ASSIGN U8133 ( .B(clk), .A(\g.we_clk [8257]));
Q_ASSIGN U8134 ( .B(clk), .A(\g.we_clk [8256]));
Q_ASSIGN U8135 ( .B(clk), .A(\g.we_clk [8255]));
Q_ASSIGN U8136 ( .B(clk), .A(\g.we_clk [8254]));
Q_ASSIGN U8137 ( .B(clk), .A(\g.we_clk [8253]));
Q_ASSIGN U8138 ( .B(clk), .A(\g.we_clk [8252]));
Q_ASSIGN U8139 ( .B(clk), .A(\g.we_clk [8251]));
Q_ASSIGN U8140 ( .B(clk), .A(\g.we_clk [8250]));
Q_ASSIGN U8141 ( .B(clk), .A(\g.we_clk [8249]));
Q_ASSIGN U8142 ( .B(clk), .A(\g.we_clk [8248]));
Q_ASSIGN U8143 ( .B(clk), .A(\g.we_clk [8247]));
Q_ASSIGN U8144 ( .B(clk), .A(\g.we_clk [8246]));
Q_ASSIGN U8145 ( .B(clk), .A(\g.we_clk [8245]));
Q_ASSIGN U8146 ( .B(clk), .A(\g.we_clk [8244]));
Q_ASSIGN U8147 ( .B(clk), .A(\g.we_clk [8243]));
Q_ASSIGN U8148 ( .B(clk), .A(\g.we_clk [8242]));
Q_ASSIGN U8149 ( .B(clk), .A(\g.we_clk [8241]));
Q_ASSIGN U8150 ( .B(clk), .A(\g.we_clk [8240]));
Q_ASSIGN U8151 ( .B(clk), .A(\g.we_clk [8239]));
Q_ASSIGN U8152 ( .B(clk), .A(\g.we_clk [8238]));
Q_ASSIGN U8153 ( .B(clk), .A(\g.we_clk [8237]));
Q_ASSIGN U8154 ( .B(clk), .A(\g.we_clk [8236]));
Q_ASSIGN U8155 ( .B(clk), .A(\g.we_clk [8235]));
Q_ASSIGN U8156 ( .B(clk), .A(\g.we_clk [8234]));
Q_ASSIGN U8157 ( .B(clk), .A(\g.we_clk [8233]));
Q_ASSIGN U8158 ( .B(clk), .A(\g.we_clk [8232]));
Q_ASSIGN U8159 ( .B(clk), .A(\g.we_clk [8231]));
Q_ASSIGN U8160 ( .B(clk), .A(\g.we_clk [8230]));
Q_ASSIGN U8161 ( .B(clk), .A(\g.we_clk [8229]));
Q_ASSIGN U8162 ( .B(clk), .A(\g.we_clk [8228]));
Q_ASSIGN U8163 ( .B(clk), .A(\g.we_clk [8227]));
Q_ASSIGN U8164 ( .B(clk), .A(\g.we_clk [8226]));
Q_ASSIGN U8165 ( .B(clk), .A(\g.we_clk [8225]));
Q_ASSIGN U8166 ( .B(clk), .A(\g.we_clk [8224]));
Q_ASSIGN U8167 ( .B(clk), .A(\g.we_clk [8223]));
Q_ASSIGN U8168 ( .B(clk), .A(\g.we_clk [8222]));
Q_ASSIGN U8169 ( .B(clk), .A(\g.we_clk [8221]));
Q_ASSIGN U8170 ( .B(clk), .A(\g.we_clk [8220]));
Q_ASSIGN U8171 ( .B(clk), .A(\g.we_clk [8219]));
Q_ASSIGN U8172 ( .B(clk), .A(\g.we_clk [8218]));
Q_ASSIGN U8173 ( .B(clk), .A(\g.we_clk [8217]));
Q_ASSIGN U8174 ( .B(clk), .A(\g.we_clk [8216]));
Q_ASSIGN U8175 ( .B(clk), .A(\g.we_clk [8215]));
Q_ASSIGN U8176 ( .B(clk), .A(\g.we_clk [8214]));
Q_ASSIGN U8177 ( .B(clk), .A(\g.we_clk [8213]));
Q_ASSIGN U8178 ( .B(clk), .A(\g.we_clk [8212]));
Q_ASSIGN U8179 ( .B(clk), .A(\g.we_clk [8211]));
Q_ASSIGN U8180 ( .B(clk), .A(\g.we_clk [8210]));
Q_ASSIGN U8181 ( .B(clk), .A(\g.we_clk [8209]));
Q_ASSIGN U8182 ( .B(clk), .A(\g.we_clk [8208]));
Q_ASSIGN U8183 ( .B(clk), .A(\g.we_clk [8207]));
Q_ASSIGN U8184 ( .B(clk), .A(\g.we_clk [8206]));
Q_ASSIGN U8185 ( .B(clk), .A(\g.we_clk [8205]));
Q_ASSIGN U8186 ( .B(clk), .A(\g.we_clk [8204]));
Q_ASSIGN U8187 ( .B(clk), .A(\g.we_clk [8203]));
Q_ASSIGN U8188 ( .B(clk), .A(\g.we_clk [8202]));
Q_ASSIGN U8189 ( .B(clk), .A(\g.we_clk [8201]));
Q_ASSIGN U8190 ( .B(clk), .A(\g.we_clk [8200]));
Q_ASSIGN U8191 ( .B(clk), .A(\g.we_clk [8199]));
Q_ASSIGN U8192 ( .B(clk), .A(\g.we_clk [8198]));
Q_ASSIGN U8193 ( .B(clk), .A(\g.we_clk [8197]));
Q_ASSIGN U8194 ( .B(clk), .A(\g.we_clk [8196]));
Q_ASSIGN U8195 ( .B(clk), .A(\g.we_clk [8195]));
Q_ASSIGN U8196 ( .B(clk), .A(\g.we_clk [8194]));
Q_ASSIGN U8197 ( .B(clk), .A(\g.we_clk [8193]));
Q_ASSIGN U8198 ( .B(clk), .A(\g.we_clk [8192]));
Q_ASSIGN U8199 ( .B(clk), .A(\g.we_clk [8191]));
Q_ASSIGN U8200 ( .B(clk), .A(\g.we_clk [8190]));
Q_ASSIGN U8201 ( .B(clk), .A(\g.we_clk [8189]));
Q_ASSIGN U8202 ( .B(clk), .A(\g.we_clk [8188]));
Q_ASSIGN U8203 ( .B(clk), .A(\g.we_clk [8187]));
Q_ASSIGN U8204 ( .B(clk), .A(\g.we_clk [8186]));
Q_ASSIGN U8205 ( .B(clk), .A(\g.we_clk [8185]));
Q_ASSIGN U8206 ( .B(clk), .A(\g.we_clk [8184]));
Q_ASSIGN U8207 ( .B(clk), .A(\g.we_clk [8183]));
Q_ASSIGN U8208 ( .B(clk), .A(\g.we_clk [8182]));
Q_ASSIGN U8209 ( .B(clk), .A(\g.we_clk [8181]));
Q_ASSIGN U8210 ( .B(clk), .A(\g.we_clk [8180]));
Q_ASSIGN U8211 ( .B(clk), .A(\g.we_clk [8179]));
Q_ASSIGN U8212 ( .B(clk), .A(\g.we_clk [8178]));
Q_ASSIGN U8213 ( .B(clk), .A(\g.we_clk [8177]));
Q_ASSIGN U8214 ( .B(clk), .A(\g.we_clk [8176]));
Q_ASSIGN U8215 ( .B(clk), .A(\g.we_clk [8175]));
Q_ASSIGN U8216 ( .B(clk), .A(\g.we_clk [8174]));
Q_ASSIGN U8217 ( .B(clk), .A(\g.we_clk [8173]));
Q_ASSIGN U8218 ( .B(clk), .A(\g.we_clk [8172]));
Q_ASSIGN U8219 ( .B(clk), .A(\g.we_clk [8171]));
Q_ASSIGN U8220 ( .B(clk), .A(\g.we_clk [8170]));
Q_ASSIGN U8221 ( .B(clk), .A(\g.we_clk [8169]));
Q_ASSIGN U8222 ( .B(clk), .A(\g.we_clk [8168]));
Q_ASSIGN U8223 ( .B(clk), .A(\g.we_clk [8167]));
Q_ASSIGN U8224 ( .B(clk), .A(\g.we_clk [8166]));
Q_ASSIGN U8225 ( .B(clk), .A(\g.we_clk [8165]));
Q_ASSIGN U8226 ( .B(clk), .A(\g.we_clk [8164]));
Q_ASSIGN U8227 ( .B(clk), .A(\g.we_clk [8163]));
Q_ASSIGN U8228 ( .B(clk), .A(\g.we_clk [8162]));
Q_ASSIGN U8229 ( .B(clk), .A(\g.we_clk [8161]));
Q_ASSIGN U8230 ( .B(clk), .A(\g.we_clk [8160]));
Q_ASSIGN U8231 ( .B(clk), .A(\g.we_clk [8159]));
Q_ASSIGN U8232 ( .B(clk), .A(\g.we_clk [8158]));
Q_ASSIGN U8233 ( .B(clk), .A(\g.we_clk [8157]));
Q_ASSIGN U8234 ( .B(clk), .A(\g.we_clk [8156]));
Q_ASSIGN U8235 ( .B(clk), .A(\g.we_clk [8155]));
Q_ASSIGN U8236 ( .B(clk), .A(\g.we_clk [8154]));
Q_ASSIGN U8237 ( .B(clk), .A(\g.we_clk [8153]));
Q_ASSIGN U8238 ( .B(clk), .A(\g.we_clk [8152]));
Q_ASSIGN U8239 ( .B(clk), .A(\g.we_clk [8151]));
Q_ASSIGN U8240 ( .B(clk), .A(\g.we_clk [8150]));
Q_ASSIGN U8241 ( .B(clk), .A(\g.we_clk [8149]));
Q_ASSIGN U8242 ( .B(clk), .A(\g.we_clk [8148]));
Q_ASSIGN U8243 ( .B(clk), .A(\g.we_clk [8147]));
Q_ASSIGN U8244 ( .B(clk), .A(\g.we_clk [8146]));
Q_ASSIGN U8245 ( .B(clk), .A(\g.we_clk [8145]));
Q_ASSIGN U8246 ( .B(clk), .A(\g.we_clk [8144]));
Q_ASSIGN U8247 ( .B(clk), .A(\g.we_clk [8143]));
Q_ASSIGN U8248 ( .B(clk), .A(\g.we_clk [8142]));
Q_ASSIGN U8249 ( .B(clk), .A(\g.we_clk [8141]));
Q_ASSIGN U8250 ( .B(clk), .A(\g.we_clk [8140]));
Q_ASSIGN U8251 ( .B(clk), .A(\g.we_clk [8139]));
Q_ASSIGN U8252 ( .B(clk), .A(\g.we_clk [8138]));
Q_ASSIGN U8253 ( .B(clk), .A(\g.we_clk [8137]));
Q_ASSIGN U8254 ( .B(clk), .A(\g.we_clk [8136]));
Q_ASSIGN U8255 ( .B(clk), .A(\g.we_clk [8135]));
Q_ASSIGN U8256 ( .B(clk), .A(\g.we_clk [8134]));
Q_ASSIGN U8257 ( .B(clk), .A(\g.we_clk [8133]));
Q_ASSIGN U8258 ( .B(clk), .A(\g.we_clk [8132]));
Q_ASSIGN U8259 ( .B(clk), .A(\g.we_clk [8131]));
Q_ASSIGN U8260 ( .B(clk), .A(\g.we_clk [8130]));
Q_ASSIGN U8261 ( .B(clk), .A(\g.we_clk [8129]));
Q_ASSIGN U8262 ( .B(clk), .A(\g.we_clk [8128]));
Q_ASSIGN U8263 ( .B(clk), .A(\g.we_clk [8127]));
Q_ASSIGN U8264 ( .B(clk), .A(\g.we_clk [8126]));
Q_ASSIGN U8265 ( .B(clk), .A(\g.we_clk [8125]));
Q_ASSIGN U8266 ( .B(clk), .A(\g.we_clk [8124]));
Q_ASSIGN U8267 ( .B(clk), .A(\g.we_clk [8123]));
Q_ASSIGN U8268 ( .B(clk), .A(\g.we_clk [8122]));
Q_ASSIGN U8269 ( .B(clk), .A(\g.we_clk [8121]));
Q_ASSIGN U8270 ( .B(clk), .A(\g.we_clk [8120]));
Q_ASSIGN U8271 ( .B(clk), .A(\g.we_clk [8119]));
Q_ASSIGN U8272 ( .B(clk), .A(\g.we_clk [8118]));
Q_ASSIGN U8273 ( .B(clk), .A(\g.we_clk [8117]));
Q_ASSIGN U8274 ( .B(clk), .A(\g.we_clk [8116]));
Q_ASSIGN U8275 ( .B(clk), .A(\g.we_clk [8115]));
Q_ASSIGN U8276 ( .B(clk), .A(\g.we_clk [8114]));
Q_ASSIGN U8277 ( .B(clk), .A(\g.we_clk [8113]));
Q_ASSIGN U8278 ( .B(clk), .A(\g.we_clk [8112]));
Q_ASSIGN U8279 ( .B(clk), .A(\g.we_clk [8111]));
Q_ASSIGN U8280 ( .B(clk), .A(\g.we_clk [8110]));
Q_ASSIGN U8281 ( .B(clk), .A(\g.we_clk [8109]));
Q_ASSIGN U8282 ( .B(clk), .A(\g.we_clk [8108]));
Q_ASSIGN U8283 ( .B(clk), .A(\g.we_clk [8107]));
Q_ASSIGN U8284 ( .B(clk), .A(\g.we_clk [8106]));
Q_ASSIGN U8285 ( .B(clk), .A(\g.we_clk [8105]));
Q_ASSIGN U8286 ( .B(clk), .A(\g.we_clk [8104]));
Q_ASSIGN U8287 ( .B(clk), .A(\g.we_clk [8103]));
Q_ASSIGN U8288 ( .B(clk), .A(\g.we_clk [8102]));
Q_ASSIGN U8289 ( .B(clk), .A(\g.we_clk [8101]));
Q_ASSIGN U8290 ( .B(clk), .A(\g.we_clk [8100]));
Q_ASSIGN U8291 ( .B(clk), .A(\g.we_clk [8099]));
Q_ASSIGN U8292 ( .B(clk), .A(\g.we_clk [8098]));
Q_ASSIGN U8293 ( .B(clk), .A(\g.we_clk [8097]));
Q_ASSIGN U8294 ( .B(clk), .A(\g.we_clk [8096]));
Q_ASSIGN U8295 ( .B(clk), .A(\g.we_clk [8095]));
Q_ASSIGN U8296 ( .B(clk), .A(\g.we_clk [8094]));
Q_ASSIGN U8297 ( .B(clk), .A(\g.we_clk [8093]));
Q_ASSIGN U8298 ( .B(clk), .A(\g.we_clk [8092]));
Q_ASSIGN U8299 ( .B(clk), .A(\g.we_clk [8091]));
Q_ASSIGN U8300 ( .B(clk), .A(\g.we_clk [8090]));
Q_ASSIGN U8301 ( .B(clk), .A(\g.we_clk [8089]));
Q_ASSIGN U8302 ( .B(clk), .A(\g.we_clk [8088]));
Q_ASSIGN U8303 ( .B(clk), .A(\g.we_clk [8087]));
Q_ASSIGN U8304 ( .B(clk), .A(\g.we_clk [8086]));
Q_ASSIGN U8305 ( .B(clk), .A(\g.we_clk [8085]));
Q_ASSIGN U8306 ( .B(clk), .A(\g.we_clk [8084]));
Q_ASSIGN U8307 ( .B(clk), .A(\g.we_clk [8083]));
Q_ASSIGN U8308 ( .B(clk), .A(\g.we_clk [8082]));
Q_ASSIGN U8309 ( .B(clk), .A(\g.we_clk [8081]));
Q_ASSIGN U8310 ( .B(clk), .A(\g.we_clk [8080]));
Q_ASSIGN U8311 ( .B(clk), .A(\g.we_clk [8079]));
Q_ASSIGN U8312 ( .B(clk), .A(\g.we_clk [8078]));
Q_ASSIGN U8313 ( .B(clk), .A(\g.we_clk [8077]));
Q_ASSIGN U8314 ( .B(clk), .A(\g.we_clk [8076]));
Q_ASSIGN U8315 ( .B(clk), .A(\g.we_clk [8075]));
Q_ASSIGN U8316 ( .B(clk), .A(\g.we_clk [8074]));
Q_ASSIGN U8317 ( .B(clk), .A(\g.we_clk [8073]));
Q_ASSIGN U8318 ( .B(clk), .A(\g.we_clk [8072]));
Q_ASSIGN U8319 ( .B(clk), .A(\g.we_clk [8071]));
Q_ASSIGN U8320 ( .B(clk), .A(\g.we_clk [8070]));
Q_ASSIGN U8321 ( .B(clk), .A(\g.we_clk [8069]));
Q_ASSIGN U8322 ( .B(clk), .A(\g.we_clk [8068]));
Q_ASSIGN U8323 ( .B(clk), .A(\g.we_clk [8067]));
Q_ASSIGN U8324 ( .B(clk), .A(\g.we_clk [8066]));
Q_ASSIGN U8325 ( .B(clk), .A(\g.we_clk [8065]));
Q_ASSIGN U8326 ( .B(clk), .A(\g.we_clk [8064]));
Q_ASSIGN U8327 ( .B(clk), .A(\g.we_clk [8063]));
Q_ASSIGN U8328 ( .B(clk), .A(\g.we_clk [8062]));
Q_ASSIGN U8329 ( .B(clk), .A(\g.we_clk [8061]));
Q_ASSIGN U8330 ( .B(clk), .A(\g.we_clk [8060]));
Q_ASSIGN U8331 ( .B(clk), .A(\g.we_clk [8059]));
Q_ASSIGN U8332 ( .B(clk), .A(\g.we_clk [8058]));
Q_ASSIGN U8333 ( .B(clk), .A(\g.we_clk [8057]));
Q_ASSIGN U8334 ( .B(clk), .A(\g.we_clk [8056]));
Q_ASSIGN U8335 ( .B(clk), .A(\g.we_clk [8055]));
Q_ASSIGN U8336 ( .B(clk), .A(\g.we_clk [8054]));
Q_ASSIGN U8337 ( .B(clk), .A(\g.we_clk [8053]));
Q_ASSIGN U8338 ( .B(clk), .A(\g.we_clk [8052]));
Q_ASSIGN U8339 ( .B(clk), .A(\g.we_clk [8051]));
Q_ASSIGN U8340 ( .B(clk), .A(\g.we_clk [8050]));
Q_ASSIGN U8341 ( .B(clk), .A(\g.we_clk [8049]));
Q_ASSIGN U8342 ( .B(clk), .A(\g.we_clk [8048]));
Q_ASSIGN U8343 ( .B(clk), .A(\g.we_clk [8047]));
Q_ASSIGN U8344 ( .B(clk), .A(\g.we_clk [8046]));
Q_ASSIGN U8345 ( .B(clk), .A(\g.we_clk [8045]));
Q_ASSIGN U8346 ( .B(clk), .A(\g.we_clk [8044]));
Q_ASSIGN U8347 ( .B(clk), .A(\g.we_clk [8043]));
Q_ASSIGN U8348 ( .B(clk), .A(\g.we_clk [8042]));
Q_ASSIGN U8349 ( .B(clk), .A(\g.we_clk [8041]));
Q_ASSIGN U8350 ( .B(clk), .A(\g.we_clk [8040]));
Q_ASSIGN U8351 ( .B(clk), .A(\g.we_clk [8039]));
Q_ASSIGN U8352 ( .B(clk), .A(\g.we_clk [8038]));
Q_ASSIGN U8353 ( .B(clk), .A(\g.we_clk [8037]));
Q_ASSIGN U8354 ( .B(clk), .A(\g.we_clk [8036]));
Q_ASSIGN U8355 ( .B(clk), .A(\g.we_clk [8035]));
Q_ASSIGN U8356 ( .B(clk), .A(\g.we_clk [8034]));
Q_ASSIGN U8357 ( .B(clk), .A(\g.we_clk [8033]));
Q_ASSIGN U8358 ( .B(clk), .A(\g.we_clk [8032]));
Q_ASSIGN U8359 ( .B(clk), .A(\g.we_clk [8031]));
Q_ASSIGN U8360 ( .B(clk), .A(\g.we_clk [8030]));
Q_ASSIGN U8361 ( .B(clk), .A(\g.we_clk [8029]));
Q_ASSIGN U8362 ( .B(clk), .A(\g.we_clk [8028]));
Q_ASSIGN U8363 ( .B(clk), .A(\g.we_clk [8027]));
Q_ASSIGN U8364 ( .B(clk), .A(\g.we_clk [8026]));
Q_ASSIGN U8365 ( .B(clk), .A(\g.we_clk [8025]));
Q_ASSIGN U8366 ( .B(clk), .A(\g.we_clk [8024]));
Q_ASSIGN U8367 ( .B(clk), .A(\g.we_clk [8023]));
Q_ASSIGN U8368 ( .B(clk), .A(\g.we_clk [8022]));
Q_ASSIGN U8369 ( .B(clk), .A(\g.we_clk [8021]));
Q_ASSIGN U8370 ( .B(clk), .A(\g.we_clk [8020]));
Q_ASSIGN U8371 ( .B(clk), .A(\g.we_clk [8019]));
Q_ASSIGN U8372 ( .B(clk), .A(\g.we_clk [8018]));
Q_ASSIGN U8373 ( .B(clk), .A(\g.we_clk [8017]));
Q_ASSIGN U8374 ( .B(clk), .A(\g.we_clk [8016]));
Q_ASSIGN U8375 ( .B(clk), .A(\g.we_clk [8015]));
Q_ASSIGN U8376 ( .B(clk), .A(\g.we_clk [8014]));
Q_ASSIGN U8377 ( .B(clk), .A(\g.we_clk [8013]));
Q_ASSIGN U8378 ( .B(clk), .A(\g.we_clk [8012]));
Q_ASSIGN U8379 ( .B(clk), .A(\g.we_clk [8011]));
Q_ASSIGN U8380 ( .B(clk), .A(\g.we_clk [8010]));
Q_ASSIGN U8381 ( .B(clk), .A(\g.we_clk [8009]));
Q_ASSIGN U8382 ( .B(clk), .A(\g.we_clk [8008]));
Q_ASSIGN U8383 ( .B(clk), .A(\g.we_clk [8007]));
Q_ASSIGN U8384 ( .B(clk), .A(\g.we_clk [8006]));
Q_ASSIGN U8385 ( .B(clk), .A(\g.we_clk [8005]));
Q_ASSIGN U8386 ( .B(clk), .A(\g.we_clk [8004]));
Q_ASSIGN U8387 ( .B(clk), .A(\g.we_clk [8003]));
Q_ASSIGN U8388 ( .B(clk), .A(\g.we_clk [8002]));
Q_ASSIGN U8389 ( .B(clk), .A(\g.we_clk [8001]));
Q_ASSIGN U8390 ( .B(clk), .A(\g.we_clk [8000]));
Q_ASSIGN U8391 ( .B(clk), .A(\g.we_clk [7999]));
Q_ASSIGN U8392 ( .B(clk), .A(\g.we_clk [7998]));
Q_ASSIGN U8393 ( .B(clk), .A(\g.we_clk [7997]));
Q_ASSIGN U8394 ( .B(clk), .A(\g.we_clk [7996]));
Q_ASSIGN U8395 ( .B(clk), .A(\g.we_clk [7995]));
Q_ASSIGN U8396 ( .B(clk), .A(\g.we_clk [7994]));
Q_ASSIGN U8397 ( .B(clk), .A(\g.we_clk [7993]));
Q_ASSIGN U8398 ( .B(clk), .A(\g.we_clk [7992]));
Q_ASSIGN U8399 ( .B(clk), .A(\g.we_clk [7991]));
Q_ASSIGN U8400 ( .B(clk), .A(\g.we_clk [7990]));
Q_ASSIGN U8401 ( .B(clk), .A(\g.we_clk [7989]));
Q_ASSIGN U8402 ( .B(clk), .A(\g.we_clk [7988]));
Q_ASSIGN U8403 ( .B(clk), .A(\g.we_clk [7987]));
Q_ASSIGN U8404 ( .B(clk), .A(\g.we_clk [7986]));
Q_ASSIGN U8405 ( .B(clk), .A(\g.we_clk [7985]));
Q_ASSIGN U8406 ( .B(clk), .A(\g.we_clk [7984]));
Q_ASSIGN U8407 ( .B(clk), .A(\g.we_clk [7983]));
Q_ASSIGN U8408 ( .B(clk), .A(\g.we_clk [7982]));
Q_ASSIGN U8409 ( .B(clk), .A(\g.we_clk [7981]));
Q_ASSIGN U8410 ( .B(clk), .A(\g.we_clk [7980]));
Q_ASSIGN U8411 ( .B(clk), .A(\g.we_clk [7979]));
Q_ASSIGN U8412 ( .B(clk), .A(\g.we_clk [7978]));
Q_ASSIGN U8413 ( .B(clk), .A(\g.we_clk [7977]));
Q_ASSIGN U8414 ( .B(clk), .A(\g.we_clk [7976]));
Q_ASSIGN U8415 ( .B(clk), .A(\g.we_clk [7975]));
Q_ASSIGN U8416 ( .B(clk), .A(\g.we_clk [7974]));
Q_ASSIGN U8417 ( .B(clk), .A(\g.we_clk [7973]));
Q_ASSIGN U8418 ( .B(clk), .A(\g.we_clk [7972]));
Q_ASSIGN U8419 ( .B(clk), .A(\g.we_clk [7971]));
Q_ASSIGN U8420 ( .B(clk), .A(\g.we_clk [7970]));
Q_ASSIGN U8421 ( .B(clk), .A(\g.we_clk [7969]));
Q_ASSIGN U8422 ( .B(clk), .A(\g.we_clk [7968]));
Q_ASSIGN U8423 ( .B(clk), .A(\g.we_clk [7967]));
Q_ASSIGN U8424 ( .B(clk), .A(\g.we_clk [7966]));
Q_ASSIGN U8425 ( .B(clk), .A(\g.we_clk [7965]));
Q_ASSIGN U8426 ( .B(clk), .A(\g.we_clk [7964]));
Q_ASSIGN U8427 ( .B(clk), .A(\g.we_clk [7963]));
Q_ASSIGN U8428 ( .B(clk), .A(\g.we_clk [7962]));
Q_ASSIGN U8429 ( .B(clk), .A(\g.we_clk [7961]));
Q_ASSIGN U8430 ( .B(clk), .A(\g.we_clk [7960]));
Q_ASSIGN U8431 ( .B(clk), .A(\g.we_clk [7959]));
Q_ASSIGN U8432 ( .B(clk), .A(\g.we_clk [7958]));
Q_ASSIGN U8433 ( .B(clk), .A(\g.we_clk [7957]));
Q_ASSIGN U8434 ( .B(clk), .A(\g.we_clk [7956]));
Q_ASSIGN U8435 ( .B(clk), .A(\g.we_clk [7955]));
Q_ASSIGN U8436 ( .B(clk), .A(\g.we_clk [7954]));
Q_ASSIGN U8437 ( .B(clk), .A(\g.we_clk [7953]));
Q_ASSIGN U8438 ( .B(clk), .A(\g.we_clk [7952]));
Q_ASSIGN U8439 ( .B(clk), .A(\g.we_clk [7951]));
Q_ASSIGN U8440 ( .B(clk), .A(\g.we_clk [7950]));
Q_ASSIGN U8441 ( .B(clk), .A(\g.we_clk [7949]));
Q_ASSIGN U8442 ( .B(clk), .A(\g.we_clk [7948]));
Q_ASSIGN U8443 ( .B(clk), .A(\g.we_clk [7947]));
Q_ASSIGN U8444 ( .B(clk), .A(\g.we_clk [7946]));
Q_ASSIGN U8445 ( .B(clk), .A(\g.we_clk [7945]));
Q_ASSIGN U8446 ( .B(clk), .A(\g.we_clk [7944]));
Q_ASSIGN U8447 ( .B(clk), .A(\g.we_clk [7943]));
Q_ASSIGN U8448 ( .B(clk), .A(\g.we_clk [7942]));
Q_ASSIGN U8449 ( .B(clk), .A(\g.we_clk [7941]));
Q_ASSIGN U8450 ( .B(clk), .A(\g.we_clk [7940]));
Q_ASSIGN U8451 ( .B(clk), .A(\g.we_clk [7939]));
Q_ASSIGN U8452 ( .B(clk), .A(\g.we_clk [7938]));
Q_ASSIGN U8453 ( .B(clk), .A(\g.we_clk [7937]));
Q_ASSIGN U8454 ( .B(clk), .A(\g.we_clk [7936]));
Q_ASSIGN U8455 ( .B(clk), .A(\g.we_clk [7935]));
Q_ASSIGN U8456 ( .B(clk), .A(\g.we_clk [7934]));
Q_ASSIGN U8457 ( .B(clk), .A(\g.we_clk [7933]));
Q_ASSIGN U8458 ( .B(clk), .A(\g.we_clk [7932]));
Q_ASSIGN U8459 ( .B(clk), .A(\g.we_clk [7931]));
Q_ASSIGN U8460 ( .B(clk), .A(\g.we_clk [7930]));
Q_ASSIGN U8461 ( .B(clk), .A(\g.we_clk [7929]));
Q_ASSIGN U8462 ( .B(clk), .A(\g.we_clk [7928]));
Q_ASSIGN U8463 ( .B(clk), .A(\g.we_clk [7927]));
Q_ASSIGN U8464 ( .B(clk), .A(\g.we_clk [7926]));
Q_ASSIGN U8465 ( .B(clk), .A(\g.we_clk [7925]));
Q_ASSIGN U8466 ( .B(clk), .A(\g.we_clk [7924]));
Q_ASSIGN U8467 ( .B(clk), .A(\g.we_clk [7923]));
Q_ASSIGN U8468 ( .B(clk), .A(\g.we_clk [7922]));
Q_ASSIGN U8469 ( .B(clk), .A(\g.we_clk [7921]));
Q_ASSIGN U8470 ( .B(clk), .A(\g.we_clk [7920]));
Q_ASSIGN U8471 ( .B(clk), .A(\g.we_clk [7919]));
Q_ASSIGN U8472 ( .B(clk), .A(\g.we_clk [7918]));
Q_ASSIGN U8473 ( .B(clk), .A(\g.we_clk [7917]));
Q_ASSIGN U8474 ( .B(clk), .A(\g.we_clk [7916]));
Q_ASSIGN U8475 ( .B(clk), .A(\g.we_clk [7915]));
Q_ASSIGN U8476 ( .B(clk), .A(\g.we_clk [7914]));
Q_ASSIGN U8477 ( .B(clk), .A(\g.we_clk [7913]));
Q_ASSIGN U8478 ( .B(clk), .A(\g.we_clk [7912]));
Q_ASSIGN U8479 ( .B(clk), .A(\g.we_clk [7911]));
Q_ASSIGN U8480 ( .B(clk), .A(\g.we_clk [7910]));
Q_ASSIGN U8481 ( .B(clk), .A(\g.we_clk [7909]));
Q_ASSIGN U8482 ( .B(clk), .A(\g.we_clk [7908]));
Q_ASSIGN U8483 ( .B(clk), .A(\g.we_clk [7907]));
Q_ASSIGN U8484 ( .B(clk), .A(\g.we_clk [7906]));
Q_ASSIGN U8485 ( .B(clk), .A(\g.we_clk [7905]));
Q_ASSIGN U8486 ( .B(clk), .A(\g.we_clk [7904]));
Q_ASSIGN U8487 ( .B(clk), .A(\g.we_clk [7903]));
Q_ASSIGN U8488 ( .B(clk), .A(\g.we_clk [7902]));
Q_ASSIGN U8489 ( .B(clk), .A(\g.we_clk [7901]));
Q_ASSIGN U8490 ( .B(clk), .A(\g.we_clk [7900]));
Q_ASSIGN U8491 ( .B(clk), .A(\g.we_clk [7899]));
Q_ASSIGN U8492 ( .B(clk), .A(\g.we_clk [7898]));
Q_ASSIGN U8493 ( .B(clk), .A(\g.we_clk [7897]));
Q_ASSIGN U8494 ( .B(clk), .A(\g.we_clk [7896]));
Q_ASSIGN U8495 ( .B(clk), .A(\g.we_clk [7895]));
Q_ASSIGN U8496 ( .B(clk), .A(\g.we_clk [7894]));
Q_ASSIGN U8497 ( .B(clk), .A(\g.we_clk [7893]));
Q_ASSIGN U8498 ( .B(clk), .A(\g.we_clk [7892]));
Q_ASSIGN U8499 ( .B(clk), .A(\g.we_clk [7891]));
Q_ASSIGN U8500 ( .B(clk), .A(\g.we_clk [7890]));
Q_ASSIGN U8501 ( .B(clk), .A(\g.we_clk [7889]));
Q_ASSIGN U8502 ( .B(clk), .A(\g.we_clk [7888]));
Q_ASSIGN U8503 ( .B(clk), .A(\g.we_clk [7887]));
Q_ASSIGN U8504 ( .B(clk), .A(\g.we_clk [7886]));
Q_ASSIGN U8505 ( .B(clk), .A(\g.we_clk [7885]));
Q_ASSIGN U8506 ( .B(clk), .A(\g.we_clk [7884]));
Q_ASSIGN U8507 ( .B(clk), .A(\g.we_clk [7883]));
Q_ASSIGN U8508 ( .B(clk), .A(\g.we_clk [7882]));
Q_ASSIGN U8509 ( .B(clk), .A(\g.we_clk [7881]));
Q_ASSIGN U8510 ( .B(clk), .A(\g.we_clk [7880]));
Q_ASSIGN U8511 ( .B(clk), .A(\g.we_clk [7879]));
Q_ASSIGN U8512 ( .B(clk), .A(\g.we_clk [7878]));
Q_ASSIGN U8513 ( .B(clk), .A(\g.we_clk [7877]));
Q_ASSIGN U8514 ( .B(clk), .A(\g.we_clk [7876]));
Q_ASSIGN U8515 ( .B(clk), .A(\g.we_clk [7875]));
Q_ASSIGN U8516 ( .B(clk), .A(\g.we_clk [7874]));
Q_ASSIGN U8517 ( .B(clk), .A(\g.we_clk [7873]));
Q_ASSIGN U8518 ( .B(clk), .A(\g.we_clk [7872]));
Q_ASSIGN U8519 ( .B(clk), .A(\g.we_clk [7871]));
Q_ASSIGN U8520 ( .B(clk), .A(\g.we_clk [7870]));
Q_ASSIGN U8521 ( .B(clk), .A(\g.we_clk [7869]));
Q_ASSIGN U8522 ( .B(clk), .A(\g.we_clk [7868]));
Q_ASSIGN U8523 ( .B(clk), .A(\g.we_clk [7867]));
Q_ASSIGN U8524 ( .B(clk), .A(\g.we_clk [7866]));
Q_ASSIGN U8525 ( .B(clk), .A(\g.we_clk [7865]));
Q_ASSIGN U8526 ( .B(clk), .A(\g.we_clk [7864]));
Q_ASSIGN U8527 ( .B(clk), .A(\g.we_clk [7863]));
Q_ASSIGN U8528 ( .B(clk), .A(\g.we_clk [7862]));
Q_ASSIGN U8529 ( .B(clk), .A(\g.we_clk [7861]));
Q_ASSIGN U8530 ( .B(clk), .A(\g.we_clk [7860]));
Q_ASSIGN U8531 ( .B(clk), .A(\g.we_clk [7859]));
Q_ASSIGN U8532 ( .B(clk), .A(\g.we_clk [7858]));
Q_ASSIGN U8533 ( .B(clk), .A(\g.we_clk [7857]));
Q_ASSIGN U8534 ( .B(clk), .A(\g.we_clk [7856]));
Q_ASSIGN U8535 ( .B(clk), .A(\g.we_clk [7855]));
Q_ASSIGN U8536 ( .B(clk), .A(\g.we_clk [7854]));
Q_ASSIGN U8537 ( .B(clk), .A(\g.we_clk [7853]));
Q_ASSIGN U8538 ( .B(clk), .A(\g.we_clk [7852]));
Q_ASSIGN U8539 ( .B(clk), .A(\g.we_clk [7851]));
Q_ASSIGN U8540 ( .B(clk), .A(\g.we_clk [7850]));
Q_ASSIGN U8541 ( .B(clk), .A(\g.we_clk [7849]));
Q_ASSIGN U8542 ( .B(clk), .A(\g.we_clk [7848]));
Q_ASSIGN U8543 ( .B(clk), .A(\g.we_clk [7847]));
Q_ASSIGN U8544 ( .B(clk), .A(\g.we_clk [7846]));
Q_ASSIGN U8545 ( .B(clk), .A(\g.we_clk [7845]));
Q_ASSIGN U8546 ( .B(clk), .A(\g.we_clk [7844]));
Q_ASSIGN U8547 ( .B(clk), .A(\g.we_clk [7843]));
Q_ASSIGN U8548 ( .B(clk), .A(\g.we_clk [7842]));
Q_ASSIGN U8549 ( .B(clk), .A(\g.we_clk [7841]));
Q_ASSIGN U8550 ( .B(clk), .A(\g.we_clk [7840]));
Q_ASSIGN U8551 ( .B(clk), .A(\g.we_clk [7839]));
Q_ASSIGN U8552 ( .B(clk), .A(\g.we_clk [7838]));
Q_ASSIGN U8553 ( .B(clk), .A(\g.we_clk [7837]));
Q_ASSIGN U8554 ( .B(clk), .A(\g.we_clk [7836]));
Q_ASSIGN U8555 ( .B(clk), .A(\g.we_clk [7835]));
Q_ASSIGN U8556 ( .B(clk), .A(\g.we_clk [7834]));
Q_ASSIGN U8557 ( .B(clk), .A(\g.we_clk [7833]));
Q_ASSIGN U8558 ( .B(clk), .A(\g.we_clk [7832]));
Q_ASSIGN U8559 ( .B(clk), .A(\g.we_clk [7831]));
Q_ASSIGN U8560 ( .B(clk), .A(\g.we_clk [7830]));
Q_ASSIGN U8561 ( .B(clk), .A(\g.we_clk [7829]));
Q_ASSIGN U8562 ( .B(clk), .A(\g.we_clk [7828]));
Q_ASSIGN U8563 ( .B(clk), .A(\g.we_clk [7827]));
Q_ASSIGN U8564 ( .B(clk), .A(\g.we_clk [7826]));
Q_ASSIGN U8565 ( .B(clk), .A(\g.we_clk [7825]));
Q_ASSIGN U8566 ( .B(clk), .A(\g.we_clk [7824]));
Q_ASSIGN U8567 ( .B(clk), .A(\g.we_clk [7823]));
Q_ASSIGN U8568 ( .B(clk), .A(\g.we_clk [7822]));
Q_ASSIGN U8569 ( .B(clk), .A(\g.we_clk [7821]));
Q_ASSIGN U8570 ( .B(clk), .A(\g.we_clk [7820]));
Q_ASSIGN U8571 ( .B(clk), .A(\g.we_clk [7819]));
Q_ASSIGN U8572 ( .B(clk), .A(\g.we_clk [7818]));
Q_ASSIGN U8573 ( .B(clk), .A(\g.we_clk [7817]));
Q_ASSIGN U8574 ( .B(clk), .A(\g.we_clk [7816]));
Q_ASSIGN U8575 ( .B(clk), .A(\g.we_clk [7815]));
Q_ASSIGN U8576 ( .B(clk), .A(\g.we_clk [7814]));
Q_ASSIGN U8577 ( .B(clk), .A(\g.we_clk [7813]));
Q_ASSIGN U8578 ( .B(clk), .A(\g.we_clk [7812]));
Q_ASSIGN U8579 ( .B(clk), .A(\g.we_clk [7811]));
Q_ASSIGN U8580 ( .B(clk), .A(\g.we_clk [7810]));
Q_ASSIGN U8581 ( .B(clk), .A(\g.we_clk [7809]));
Q_ASSIGN U8582 ( .B(clk), .A(\g.we_clk [7808]));
Q_ASSIGN U8583 ( .B(clk), .A(\g.we_clk [7807]));
Q_ASSIGN U8584 ( .B(clk), .A(\g.we_clk [7806]));
Q_ASSIGN U8585 ( .B(clk), .A(\g.we_clk [7805]));
Q_ASSIGN U8586 ( .B(clk), .A(\g.we_clk [7804]));
Q_ASSIGN U8587 ( .B(clk), .A(\g.we_clk [7803]));
Q_ASSIGN U8588 ( .B(clk), .A(\g.we_clk [7802]));
Q_ASSIGN U8589 ( .B(clk), .A(\g.we_clk [7801]));
Q_ASSIGN U8590 ( .B(clk), .A(\g.we_clk [7800]));
Q_ASSIGN U8591 ( .B(clk), .A(\g.we_clk [7799]));
Q_ASSIGN U8592 ( .B(clk), .A(\g.we_clk [7798]));
Q_ASSIGN U8593 ( .B(clk), .A(\g.we_clk [7797]));
Q_ASSIGN U8594 ( .B(clk), .A(\g.we_clk [7796]));
Q_ASSIGN U8595 ( .B(clk), .A(\g.we_clk [7795]));
Q_ASSIGN U8596 ( .B(clk), .A(\g.we_clk [7794]));
Q_ASSIGN U8597 ( .B(clk), .A(\g.we_clk [7793]));
Q_ASSIGN U8598 ( .B(clk), .A(\g.we_clk [7792]));
Q_ASSIGN U8599 ( .B(clk), .A(\g.we_clk [7791]));
Q_ASSIGN U8600 ( .B(clk), .A(\g.we_clk [7790]));
Q_ASSIGN U8601 ( .B(clk), .A(\g.we_clk [7789]));
Q_ASSIGN U8602 ( .B(clk), .A(\g.we_clk [7788]));
Q_ASSIGN U8603 ( .B(clk), .A(\g.we_clk [7787]));
Q_ASSIGN U8604 ( .B(clk), .A(\g.we_clk [7786]));
Q_ASSIGN U8605 ( .B(clk), .A(\g.we_clk [7785]));
Q_ASSIGN U8606 ( .B(clk), .A(\g.we_clk [7784]));
Q_ASSIGN U8607 ( .B(clk), .A(\g.we_clk [7783]));
Q_ASSIGN U8608 ( .B(clk), .A(\g.we_clk [7782]));
Q_ASSIGN U8609 ( .B(clk), .A(\g.we_clk [7781]));
Q_ASSIGN U8610 ( .B(clk), .A(\g.we_clk [7780]));
Q_ASSIGN U8611 ( .B(clk), .A(\g.we_clk [7779]));
Q_ASSIGN U8612 ( .B(clk), .A(\g.we_clk [7778]));
Q_ASSIGN U8613 ( .B(clk), .A(\g.we_clk [7777]));
Q_ASSIGN U8614 ( .B(clk), .A(\g.we_clk [7776]));
Q_ASSIGN U8615 ( .B(clk), .A(\g.we_clk [7775]));
Q_ASSIGN U8616 ( .B(clk), .A(\g.we_clk [7774]));
Q_ASSIGN U8617 ( .B(clk), .A(\g.we_clk [7773]));
Q_ASSIGN U8618 ( .B(clk), .A(\g.we_clk [7772]));
Q_ASSIGN U8619 ( .B(clk), .A(\g.we_clk [7771]));
Q_ASSIGN U8620 ( .B(clk), .A(\g.we_clk [7770]));
Q_ASSIGN U8621 ( .B(clk), .A(\g.we_clk [7769]));
Q_ASSIGN U8622 ( .B(clk), .A(\g.we_clk [7768]));
Q_ASSIGN U8623 ( .B(clk), .A(\g.we_clk [7767]));
Q_ASSIGN U8624 ( .B(clk), .A(\g.we_clk [7766]));
Q_ASSIGN U8625 ( .B(clk), .A(\g.we_clk [7765]));
Q_ASSIGN U8626 ( .B(clk), .A(\g.we_clk [7764]));
Q_ASSIGN U8627 ( .B(clk), .A(\g.we_clk [7763]));
Q_ASSIGN U8628 ( .B(clk), .A(\g.we_clk [7762]));
Q_ASSIGN U8629 ( .B(clk), .A(\g.we_clk [7761]));
Q_ASSIGN U8630 ( .B(clk), .A(\g.we_clk [7760]));
Q_ASSIGN U8631 ( .B(clk), .A(\g.we_clk [7759]));
Q_ASSIGN U8632 ( .B(clk), .A(\g.we_clk [7758]));
Q_ASSIGN U8633 ( .B(clk), .A(\g.we_clk [7757]));
Q_ASSIGN U8634 ( .B(clk), .A(\g.we_clk [7756]));
Q_ASSIGN U8635 ( .B(clk), .A(\g.we_clk [7755]));
Q_ASSIGN U8636 ( .B(clk), .A(\g.we_clk [7754]));
Q_ASSIGN U8637 ( .B(clk), .A(\g.we_clk [7753]));
Q_ASSIGN U8638 ( .B(clk), .A(\g.we_clk [7752]));
Q_ASSIGN U8639 ( .B(clk), .A(\g.we_clk [7751]));
Q_ASSIGN U8640 ( .B(clk), .A(\g.we_clk [7750]));
Q_ASSIGN U8641 ( .B(clk), .A(\g.we_clk [7749]));
Q_ASSIGN U8642 ( .B(clk), .A(\g.we_clk [7748]));
Q_ASSIGN U8643 ( .B(clk), .A(\g.we_clk [7747]));
Q_ASSIGN U8644 ( .B(clk), .A(\g.we_clk [7746]));
Q_ASSIGN U8645 ( .B(clk), .A(\g.we_clk [7745]));
Q_ASSIGN U8646 ( .B(clk), .A(\g.we_clk [7744]));
Q_ASSIGN U8647 ( .B(clk), .A(\g.we_clk [7743]));
Q_ASSIGN U8648 ( .B(clk), .A(\g.we_clk [7742]));
Q_ASSIGN U8649 ( .B(clk), .A(\g.we_clk [7741]));
Q_ASSIGN U8650 ( .B(clk), .A(\g.we_clk [7740]));
Q_ASSIGN U8651 ( .B(clk), .A(\g.we_clk [7739]));
Q_ASSIGN U8652 ( .B(clk), .A(\g.we_clk [7738]));
Q_ASSIGN U8653 ( .B(clk), .A(\g.we_clk [7737]));
Q_ASSIGN U8654 ( .B(clk), .A(\g.we_clk [7736]));
Q_ASSIGN U8655 ( .B(clk), .A(\g.we_clk [7735]));
Q_ASSIGN U8656 ( .B(clk), .A(\g.we_clk [7734]));
Q_ASSIGN U8657 ( .B(clk), .A(\g.we_clk [7733]));
Q_ASSIGN U8658 ( .B(clk), .A(\g.we_clk [7732]));
Q_ASSIGN U8659 ( .B(clk), .A(\g.we_clk [7731]));
Q_ASSIGN U8660 ( .B(clk), .A(\g.we_clk [7730]));
Q_ASSIGN U8661 ( .B(clk), .A(\g.we_clk [7729]));
Q_ASSIGN U8662 ( .B(clk), .A(\g.we_clk [7728]));
Q_ASSIGN U8663 ( .B(clk), .A(\g.we_clk [7727]));
Q_ASSIGN U8664 ( .B(clk), .A(\g.we_clk [7726]));
Q_ASSIGN U8665 ( .B(clk), .A(\g.we_clk [7725]));
Q_ASSIGN U8666 ( .B(clk), .A(\g.we_clk [7724]));
Q_ASSIGN U8667 ( .B(clk), .A(\g.we_clk [7723]));
Q_ASSIGN U8668 ( .B(clk), .A(\g.we_clk [7722]));
Q_ASSIGN U8669 ( .B(clk), .A(\g.we_clk [7721]));
Q_ASSIGN U8670 ( .B(clk), .A(\g.we_clk [7720]));
Q_ASSIGN U8671 ( .B(clk), .A(\g.we_clk [7719]));
Q_ASSIGN U8672 ( .B(clk), .A(\g.we_clk [7718]));
Q_ASSIGN U8673 ( .B(clk), .A(\g.we_clk [7717]));
Q_ASSIGN U8674 ( .B(clk), .A(\g.we_clk [7716]));
Q_ASSIGN U8675 ( .B(clk), .A(\g.we_clk [7715]));
Q_ASSIGN U8676 ( .B(clk), .A(\g.we_clk [7714]));
Q_ASSIGN U8677 ( .B(clk), .A(\g.we_clk [7713]));
Q_ASSIGN U8678 ( .B(clk), .A(\g.we_clk [7712]));
Q_ASSIGN U8679 ( .B(clk), .A(\g.we_clk [7711]));
Q_ASSIGN U8680 ( .B(clk), .A(\g.we_clk [7710]));
Q_ASSIGN U8681 ( .B(clk), .A(\g.we_clk [7709]));
Q_ASSIGN U8682 ( .B(clk), .A(\g.we_clk [7708]));
Q_ASSIGN U8683 ( .B(clk), .A(\g.we_clk [7707]));
Q_ASSIGN U8684 ( .B(clk), .A(\g.we_clk [7706]));
Q_ASSIGN U8685 ( .B(clk), .A(\g.we_clk [7705]));
Q_ASSIGN U8686 ( .B(clk), .A(\g.we_clk [7704]));
Q_ASSIGN U8687 ( .B(clk), .A(\g.we_clk [7703]));
Q_ASSIGN U8688 ( .B(clk), .A(\g.we_clk [7702]));
Q_ASSIGN U8689 ( .B(clk), .A(\g.we_clk [7701]));
Q_ASSIGN U8690 ( .B(clk), .A(\g.we_clk [7700]));
Q_ASSIGN U8691 ( .B(clk), .A(\g.we_clk [7699]));
Q_ASSIGN U8692 ( .B(clk), .A(\g.we_clk [7698]));
Q_ASSIGN U8693 ( .B(clk), .A(\g.we_clk [7697]));
Q_ASSIGN U8694 ( .B(clk), .A(\g.we_clk [7696]));
Q_ASSIGN U8695 ( .B(clk), .A(\g.we_clk [7695]));
Q_ASSIGN U8696 ( .B(clk), .A(\g.we_clk [7694]));
Q_ASSIGN U8697 ( .B(clk), .A(\g.we_clk [7693]));
Q_ASSIGN U8698 ( .B(clk), .A(\g.we_clk [7692]));
Q_ASSIGN U8699 ( .B(clk), .A(\g.we_clk [7691]));
Q_ASSIGN U8700 ( .B(clk), .A(\g.we_clk [7690]));
Q_ASSIGN U8701 ( .B(clk), .A(\g.we_clk [7689]));
Q_ASSIGN U8702 ( .B(clk), .A(\g.we_clk [7688]));
Q_ASSIGN U8703 ( .B(clk), .A(\g.we_clk [7687]));
Q_ASSIGN U8704 ( .B(clk), .A(\g.we_clk [7686]));
Q_ASSIGN U8705 ( .B(clk), .A(\g.we_clk [7685]));
Q_ASSIGN U8706 ( .B(clk), .A(\g.we_clk [7684]));
Q_ASSIGN U8707 ( .B(clk), .A(\g.we_clk [7683]));
Q_ASSIGN U8708 ( .B(clk), .A(\g.we_clk [7682]));
Q_ASSIGN U8709 ( .B(clk), .A(\g.we_clk [7681]));
Q_ASSIGN U8710 ( .B(clk), .A(\g.we_clk [7680]));
Q_ASSIGN U8711 ( .B(clk), .A(\g.we_clk [7679]));
Q_ASSIGN U8712 ( .B(clk), .A(\g.we_clk [7678]));
Q_ASSIGN U8713 ( .B(clk), .A(\g.we_clk [7677]));
Q_ASSIGN U8714 ( .B(clk), .A(\g.we_clk [7676]));
Q_ASSIGN U8715 ( .B(clk), .A(\g.we_clk [7675]));
Q_ASSIGN U8716 ( .B(clk), .A(\g.we_clk [7674]));
Q_ASSIGN U8717 ( .B(clk), .A(\g.we_clk [7673]));
Q_ASSIGN U8718 ( .B(clk), .A(\g.we_clk [7672]));
Q_ASSIGN U8719 ( .B(clk), .A(\g.we_clk [7671]));
Q_ASSIGN U8720 ( .B(clk), .A(\g.we_clk [7670]));
Q_ASSIGN U8721 ( .B(clk), .A(\g.we_clk [7669]));
Q_ASSIGN U8722 ( .B(clk), .A(\g.we_clk [7668]));
Q_ASSIGN U8723 ( .B(clk), .A(\g.we_clk [7667]));
Q_ASSIGN U8724 ( .B(clk), .A(\g.we_clk [7666]));
Q_ASSIGN U8725 ( .B(clk), .A(\g.we_clk [7665]));
Q_ASSIGN U8726 ( .B(clk), .A(\g.we_clk [7664]));
Q_ASSIGN U8727 ( .B(clk), .A(\g.we_clk [7663]));
Q_ASSIGN U8728 ( .B(clk), .A(\g.we_clk [7662]));
Q_ASSIGN U8729 ( .B(clk), .A(\g.we_clk [7661]));
Q_ASSIGN U8730 ( .B(clk), .A(\g.we_clk [7660]));
Q_ASSIGN U8731 ( .B(clk), .A(\g.we_clk [7659]));
Q_ASSIGN U8732 ( .B(clk), .A(\g.we_clk [7658]));
Q_ASSIGN U8733 ( .B(clk), .A(\g.we_clk [7657]));
Q_ASSIGN U8734 ( .B(clk), .A(\g.we_clk [7656]));
Q_ASSIGN U8735 ( .B(clk), .A(\g.we_clk [7655]));
Q_ASSIGN U8736 ( .B(clk), .A(\g.we_clk [7654]));
Q_ASSIGN U8737 ( .B(clk), .A(\g.we_clk [7653]));
Q_ASSIGN U8738 ( .B(clk), .A(\g.we_clk [7652]));
Q_ASSIGN U8739 ( .B(clk), .A(\g.we_clk [7651]));
Q_ASSIGN U8740 ( .B(clk), .A(\g.we_clk [7650]));
Q_ASSIGN U8741 ( .B(clk), .A(\g.we_clk [7649]));
Q_ASSIGN U8742 ( .B(clk), .A(\g.we_clk [7648]));
Q_ASSIGN U8743 ( .B(clk), .A(\g.we_clk [7647]));
Q_ASSIGN U8744 ( .B(clk), .A(\g.we_clk [7646]));
Q_ASSIGN U8745 ( .B(clk), .A(\g.we_clk [7645]));
Q_ASSIGN U8746 ( .B(clk), .A(\g.we_clk [7644]));
Q_ASSIGN U8747 ( .B(clk), .A(\g.we_clk [7643]));
Q_ASSIGN U8748 ( .B(clk), .A(\g.we_clk [7642]));
Q_ASSIGN U8749 ( .B(clk), .A(\g.we_clk [7641]));
Q_ASSIGN U8750 ( .B(clk), .A(\g.we_clk [7640]));
Q_ASSIGN U8751 ( .B(clk), .A(\g.we_clk [7639]));
Q_ASSIGN U8752 ( .B(clk), .A(\g.we_clk [7638]));
Q_ASSIGN U8753 ( .B(clk), .A(\g.we_clk [7637]));
Q_ASSIGN U8754 ( .B(clk), .A(\g.we_clk [7636]));
Q_ASSIGN U8755 ( .B(clk), .A(\g.we_clk [7635]));
Q_ASSIGN U8756 ( .B(clk), .A(\g.we_clk [7634]));
Q_ASSIGN U8757 ( .B(clk), .A(\g.we_clk [7633]));
Q_ASSIGN U8758 ( .B(clk), .A(\g.we_clk [7632]));
Q_ASSIGN U8759 ( .B(clk), .A(\g.we_clk [7631]));
Q_ASSIGN U8760 ( .B(clk), .A(\g.we_clk [7630]));
Q_ASSIGN U8761 ( .B(clk), .A(\g.we_clk [7629]));
Q_ASSIGN U8762 ( .B(clk), .A(\g.we_clk [7628]));
Q_ASSIGN U8763 ( .B(clk), .A(\g.we_clk [7627]));
Q_ASSIGN U8764 ( .B(clk), .A(\g.we_clk [7626]));
Q_ASSIGN U8765 ( .B(clk), .A(\g.we_clk [7625]));
Q_ASSIGN U8766 ( .B(clk), .A(\g.we_clk [7624]));
Q_ASSIGN U8767 ( .B(clk), .A(\g.we_clk [7623]));
Q_ASSIGN U8768 ( .B(clk), .A(\g.we_clk [7622]));
Q_ASSIGN U8769 ( .B(clk), .A(\g.we_clk [7621]));
Q_ASSIGN U8770 ( .B(clk), .A(\g.we_clk [7620]));
Q_ASSIGN U8771 ( .B(clk), .A(\g.we_clk [7619]));
Q_ASSIGN U8772 ( .B(clk), .A(\g.we_clk [7618]));
Q_ASSIGN U8773 ( .B(clk), .A(\g.we_clk [7617]));
Q_ASSIGN U8774 ( .B(clk), .A(\g.we_clk [7616]));
Q_ASSIGN U8775 ( .B(clk), .A(\g.we_clk [7615]));
Q_ASSIGN U8776 ( .B(clk), .A(\g.we_clk [7614]));
Q_ASSIGN U8777 ( .B(clk), .A(\g.we_clk [7613]));
Q_ASSIGN U8778 ( .B(clk), .A(\g.we_clk [7612]));
Q_ASSIGN U8779 ( .B(clk), .A(\g.we_clk [7611]));
Q_ASSIGN U8780 ( .B(clk), .A(\g.we_clk [7610]));
Q_ASSIGN U8781 ( .B(clk), .A(\g.we_clk [7609]));
Q_ASSIGN U8782 ( .B(clk), .A(\g.we_clk [7608]));
Q_ASSIGN U8783 ( .B(clk), .A(\g.we_clk [7607]));
Q_ASSIGN U8784 ( .B(clk), .A(\g.we_clk [7606]));
Q_ASSIGN U8785 ( .B(clk), .A(\g.we_clk [7605]));
Q_ASSIGN U8786 ( .B(clk), .A(\g.we_clk [7604]));
Q_ASSIGN U8787 ( .B(clk), .A(\g.we_clk [7603]));
Q_ASSIGN U8788 ( .B(clk), .A(\g.we_clk [7602]));
Q_ASSIGN U8789 ( .B(clk), .A(\g.we_clk [7601]));
Q_ASSIGN U8790 ( .B(clk), .A(\g.we_clk [7600]));
Q_ASSIGN U8791 ( .B(clk), .A(\g.we_clk [7599]));
Q_ASSIGN U8792 ( .B(clk), .A(\g.we_clk [7598]));
Q_ASSIGN U8793 ( .B(clk), .A(\g.we_clk [7597]));
Q_ASSIGN U8794 ( .B(clk), .A(\g.we_clk [7596]));
Q_ASSIGN U8795 ( .B(clk), .A(\g.we_clk [7595]));
Q_ASSIGN U8796 ( .B(clk), .A(\g.we_clk [7594]));
Q_ASSIGN U8797 ( .B(clk), .A(\g.we_clk [7593]));
Q_ASSIGN U8798 ( .B(clk), .A(\g.we_clk [7592]));
Q_ASSIGN U8799 ( .B(clk), .A(\g.we_clk [7591]));
Q_ASSIGN U8800 ( .B(clk), .A(\g.we_clk [7590]));
Q_ASSIGN U8801 ( .B(clk), .A(\g.we_clk [7589]));
Q_ASSIGN U8802 ( .B(clk), .A(\g.we_clk [7588]));
Q_ASSIGN U8803 ( .B(clk), .A(\g.we_clk [7587]));
Q_ASSIGN U8804 ( .B(clk), .A(\g.we_clk [7586]));
Q_ASSIGN U8805 ( .B(clk), .A(\g.we_clk [7585]));
Q_ASSIGN U8806 ( .B(clk), .A(\g.we_clk [7584]));
Q_ASSIGN U8807 ( .B(clk), .A(\g.we_clk [7583]));
Q_ASSIGN U8808 ( .B(clk), .A(\g.we_clk [7582]));
Q_ASSIGN U8809 ( .B(clk), .A(\g.we_clk [7581]));
Q_ASSIGN U8810 ( .B(clk), .A(\g.we_clk [7580]));
Q_ASSIGN U8811 ( .B(clk), .A(\g.we_clk [7579]));
Q_ASSIGN U8812 ( .B(clk), .A(\g.we_clk [7578]));
Q_ASSIGN U8813 ( .B(clk), .A(\g.we_clk [7577]));
Q_ASSIGN U8814 ( .B(clk), .A(\g.we_clk [7576]));
Q_ASSIGN U8815 ( .B(clk), .A(\g.we_clk [7575]));
Q_ASSIGN U8816 ( .B(clk), .A(\g.we_clk [7574]));
Q_ASSIGN U8817 ( .B(clk), .A(\g.we_clk [7573]));
Q_ASSIGN U8818 ( .B(clk), .A(\g.we_clk [7572]));
Q_ASSIGN U8819 ( .B(clk), .A(\g.we_clk [7571]));
Q_ASSIGN U8820 ( .B(clk), .A(\g.we_clk [7570]));
Q_ASSIGN U8821 ( .B(clk), .A(\g.we_clk [7569]));
Q_ASSIGN U8822 ( .B(clk), .A(\g.we_clk [7568]));
Q_ASSIGN U8823 ( .B(clk), .A(\g.we_clk [7567]));
Q_ASSIGN U8824 ( .B(clk), .A(\g.we_clk [7566]));
Q_ASSIGN U8825 ( .B(clk), .A(\g.we_clk [7565]));
Q_ASSIGN U8826 ( .B(clk), .A(\g.we_clk [7564]));
Q_ASSIGN U8827 ( .B(clk), .A(\g.we_clk [7563]));
Q_ASSIGN U8828 ( .B(clk), .A(\g.we_clk [7562]));
Q_ASSIGN U8829 ( .B(clk), .A(\g.we_clk [7561]));
Q_ASSIGN U8830 ( .B(clk), .A(\g.we_clk [7560]));
Q_ASSIGN U8831 ( .B(clk), .A(\g.we_clk [7559]));
Q_ASSIGN U8832 ( .B(clk), .A(\g.we_clk [7558]));
Q_ASSIGN U8833 ( .B(clk), .A(\g.we_clk [7557]));
Q_ASSIGN U8834 ( .B(clk), .A(\g.we_clk [7556]));
Q_ASSIGN U8835 ( .B(clk), .A(\g.we_clk [7555]));
Q_ASSIGN U8836 ( .B(clk), .A(\g.we_clk [7554]));
Q_ASSIGN U8837 ( .B(clk), .A(\g.we_clk [7553]));
Q_ASSIGN U8838 ( .B(clk), .A(\g.we_clk [7552]));
Q_ASSIGN U8839 ( .B(clk), .A(\g.we_clk [7551]));
Q_ASSIGN U8840 ( .B(clk), .A(\g.we_clk [7550]));
Q_ASSIGN U8841 ( .B(clk), .A(\g.we_clk [7549]));
Q_ASSIGN U8842 ( .B(clk), .A(\g.we_clk [7548]));
Q_ASSIGN U8843 ( .B(clk), .A(\g.we_clk [7547]));
Q_ASSIGN U8844 ( .B(clk), .A(\g.we_clk [7546]));
Q_ASSIGN U8845 ( .B(clk), .A(\g.we_clk [7545]));
Q_ASSIGN U8846 ( .B(clk), .A(\g.we_clk [7544]));
Q_ASSIGN U8847 ( .B(clk), .A(\g.we_clk [7543]));
Q_ASSIGN U8848 ( .B(clk), .A(\g.we_clk [7542]));
Q_ASSIGN U8849 ( .B(clk), .A(\g.we_clk [7541]));
Q_ASSIGN U8850 ( .B(clk), .A(\g.we_clk [7540]));
Q_ASSIGN U8851 ( .B(clk), .A(\g.we_clk [7539]));
Q_ASSIGN U8852 ( .B(clk), .A(\g.we_clk [7538]));
Q_ASSIGN U8853 ( .B(clk), .A(\g.we_clk [7537]));
Q_ASSIGN U8854 ( .B(clk), .A(\g.we_clk [7536]));
Q_ASSIGN U8855 ( .B(clk), .A(\g.we_clk [7535]));
Q_ASSIGN U8856 ( .B(clk), .A(\g.we_clk [7534]));
Q_ASSIGN U8857 ( .B(clk), .A(\g.we_clk [7533]));
Q_ASSIGN U8858 ( .B(clk), .A(\g.we_clk [7532]));
Q_ASSIGN U8859 ( .B(clk), .A(\g.we_clk [7531]));
Q_ASSIGN U8860 ( .B(clk), .A(\g.we_clk [7530]));
Q_ASSIGN U8861 ( .B(clk), .A(\g.we_clk [7529]));
Q_ASSIGN U8862 ( .B(clk), .A(\g.we_clk [7528]));
Q_ASSIGN U8863 ( .B(clk), .A(\g.we_clk [7527]));
Q_ASSIGN U8864 ( .B(clk), .A(\g.we_clk [7526]));
Q_ASSIGN U8865 ( .B(clk), .A(\g.we_clk [7525]));
Q_ASSIGN U8866 ( .B(clk), .A(\g.we_clk [7524]));
Q_ASSIGN U8867 ( .B(clk), .A(\g.we_clk [7523]));
Q_ASSIGN U8868 ( .B(clk), .A(\g.we_clk [7522]));
Q_ASSIGN U8869 ( .B(clk), .A(\g.we_clk [7521]));
Q_ASSIGN U8870 ( .B(clk), .A(\g.we_clk [7520]));
Q_ASSIGN U8871 ( .B(clk), .A(\g.we_clk [7519]));
Q_ASSIGN U8872 ( .B(clk), .A(\g.we_clk [7518]));
Q_ASSIGN U8873 ( .B(clk), .A(\g.we_clk [7517]));
Q_ASSIGN U8874 ( .B(clk), .A(\g.we_clk [7516]));
Q_ASSIGN U8875 ( .B(clk), .A(\g.we_clk [7515]));
Q_ASSIGN U8876 ( .B(clk), .A(\g.we_clk [7514]));
Q_ASSIGN U8877 ( .B(clk), .A(\g.we_clk [7513]));
Q_ASSIGN U8878 ( .B(clk), .A(\g.we_clk [7512]));
Q_ASSIGN U8879 ( .B(clk), .A(\g.we_clk [7511]));
Q_ASSIGN U8880 ( .B(clk), .A(\g.we_clk [7510]));
Q_ASSIGN U8881 ( .B(clk), .A(\g.we_clk [7509]));
Q_ASSIGN U8882 ( .B(clk), .A(\g.we_clk [7508]));
Q_ASSIGN U8883 ( .B(clk), .A(\g.we_clk [7507]));
Q_ASSIGN U8884 ( .B(clk), .A(\g.we_clk [7506]));
Q_ASSIGN U8885 ( .B(clk), .A(\g.we_clk [7505]));
Q_ASSIGN U8886 ( .B(clk), .A(\g.we_clk [7504]));
Q_ASSIGN U8887 ( .B(clk), .A(\g.we_clk [7503]));
Q_ASSIGN U8888 ( .B(clk), .A(\g.we_clk [7502]));
Q_ASSIGN U8889 ( .B(clk), .A(\g.we_clk [7501]));
Q_ASSIGN U8890 ( .B(clk), .A(\g.we_clk [7500]));
Q_ASSIGN U8891 ( .B(clk), .A(\g.we_clk [7499]));
Q_ASSIGN U8892 ( .B(clk), .A(\g.we_clk [7498]));
Q_ASSIGN U8893 ( .B(clk), .A(\g.we_clk [7497]));
Q_ASSIGN U8894 ( .B(clk), .A(\g.we_clk [7496]));
Q_ASSIGN U8895 ( .B(clk), .A(\g.we_clk [7495]));
Q_ASSIGN U8896 ( .B(clk), .A(\g.we_clk [7494]));
Q_ASSIGN U8897 ( .B(clk), .A(\g.we_clk [7493]));
Q_ASSIGN U8898 ( .B(clk), .A(\g.we_clk [7492]));
Q_ASSIGN U8899 ( .B(clk), .A(\g.we_clk [7491]));
Q_ASSIGN U8900 ( .B(clk), .A(\g.we_clk [7490]));
Q_ASSIGN U8901 ( .B(clk), .A(\g.we_clk [7489]));
Q_ASSIGN U8902 ( .B(clk), .A(\g.we_clk [7488]));
Q_ASSIGN U8903 ( .B(clk), .A(\g.we_clk [7487]));
Q_ASSIGN U8904 ( .B(clk), .A(\g.we_clk [7486]));
Q_ASSIGN U8905 ( .B(clk), .A(\g.we_clk [7485]));
Q_ASSIGN U8906 ( .B(clk), .A(\g.we_clk [7484]));
Q_ASSIGN U8907 ( .B(clk), .A(\g.we_clk [7483]));
Q_ASSIGN U8908 ( .B(clk), .A(\g.we_clk [7482]));
Q_ASSIGN U8909 ( .B(clk), .A(\g.we_clk [7481]));
Q_ASSIGN U8910 ( .B(clk), .A(\g.we_clk [7480]));
Q_ASSIGN U8911 ( .B(clk), .A(\g.we_clk [7479]));
Q_ASSIGN U8912 ( .B(clk), .A(\g.we_clk [7478]));
Q_ASSIGN U8913 ( .B(clk), .A(\g.we_clk [7477]));
Q_ASSIGN U8914 ( .B(clk), .A(\g.we_clk [7476]));
Q_ASSIGN U8915 ( .B(clk), .A(\g.we_clk [7475]));
Q_ASSIGN U8916 ( .B(clk), .A(\g.we_clk [7474]));
Q_ASSIGN U8917 ( .B(clk), .A(\g.we_clk [7473]));
Q_ASSIGN U8918 ( .B(clk), .A(\g.we_clk [7472]));
Q_ASSIGN U8919 ( .B(clk), .A(\g.we_clk [7471]));
Q_ASSIGN U8920 ( .B(clk), .A(\g.we_clk [7470]));
Q_ASSIGN U8921 ( .B(clk), .A(\g.we_clk [7469]));
Q_ASSIGN U8922 ( .B(clk), .A(\g.we_clk [7468]));
Q_ASSIGN U8923 ( .B(clk), .A(\g.we_clk [7467]));
Q_ASSIGN U8924 ( .B(clk), .A(\g.we_clk [7466]));
Q_ASSIGN U8925 ( .B(clk), .A(\g.we_clk [7465]));
Q_ASSIGN U8926 ( .B(clk), .A(\g.we_clk [7464]));
Q_ASSIGN U8927 ( .B(clk), .A(\g.we_clk [7463]));
Q_ASSIGN U8928 ( .B(clk), .A(\g.we_clk [7462]));
Q_ASSIGN U8929 ( .B(clk), .A(\g.we_clk [7461]));
Q_ASSIGN U8930 ( .B(clk), .A(\g.we_clk [7460]));
Q_ASSIGN U8931 ( .B(clk), .A(\g.we_clk [7459]));
Q_ASSIGN U8932 ( .B(clk), .A(\g.we_clk [7458]));
Q_ASSIGN U8933 ( .B(clk), .A(\g.we_clk [7457]));
Q_ASSIGN U8934 ( .B(clk), .A(\g.we_clk [7456]));
Q_ASSIGN U8935 ( .B(clk), .A(\g.we_clk [7455]));
Q_ASSIGN U8936 ( .B(clk), .A(\g.we_clk [7454]));
Q_ASSIGN U8937 ( .B(clk), .A(\g.we_clk [7453]));
Q_ASSIGN U8938 ( .B(clk), .A(\g.we_clk [7452]));
Q_ASSIGN U8939 ( .B(clk), .A(\g.we_clk [7451]));
Q_ASSIGN U8940 ( .B(clk), .A(\g.we_clk [7450]));
Q_ASSIGN U8941 ( .B(clk), .A(\g.we_clk [7449]));
Q_ASSIGN U8942 ( .B(clk), .A(\g.we_clk [7448]));
Q_ASSIGN U8943 ( .B(clk), .A(\g.we_clk [7447]));
Q_ASSIGN U8944 ( .B(clk), .A(\g.we_clk [7446]));
Q_ASSIGN U8945 ( .B(clk), .A(\g.we_clk [7445]));
Q_ASSIGN U8946 ( .B(clk), .A(\g.we_clk [7444]));
Q_ASSIGN U8947 ( .B(clk), .A(\g.we_clk [7443]));
Q_ASSIGN U8948 ( .B(clk), .A(\g.we_clk [7442]));
Q_ASSIGN U8949 ( .B(clk), .A(\g.we_clk [7441]));
Q_ASSIGN U8950 ( .B(clk), .A(\g.we_clk [7440]));
Q_ASSIGN U8951 ( .B(clk), .A(\g.we_clk [7439]));
Q_ASSIGN U8952 ( .B(clk), .A(\g.we_clk [7438]));
Q_ASSIGN U8953 ( .B(clk), .A(\g.we_clk [7437]));
Q_ASSIGN U8954 ( .B(clk), .A(\g.we_clk [7436]));
Q_ASSIGN U8955 ( .B(clk), .A(\g.we_clk [7435]));
Q_ASSIGN U8956 ( .B(clk), .A(\g.we_clk [7434]));
Q_ASSIGN U8957 ( .B(clk), .A(\g.we_clk [7433]));
Q_ASSIGN U8958 ( .B(clk), .A(\g.we_clk [7432]));
Q_ASSIGN U8959 ( .B(clk), .A(\g.we_clk [7431]));
Q_ASSIGN U8960 ( .B(clk), .A(\g.we_clk [7430]));
Q_ASSIGN U8961 ( .B(clk), .A(\g.we_clk [7429]));
Q_ASSIGN U8962 ( .B(clk), .A(\g.we_clk [7428]));
Q_ASSIGN U8963 ( .B(clk), .A(\g.we_clk [7427]));
Q_ASSIGN U8964 ( .B(clk), .A(\g.we_clk [7426]));
Q_ASSIGN U8965 ( .B(clk), .A(\g.we_clk [7425]));
Q_ASSIGN U8966 ( .B(clk), .A(\g.we_clk [7424]));
Q_ASSIGN U8967 ( .B(clk), .A(\g.we_clk [7423]));
Q_ASSIGN U8968 ( .B(clk), .A(\g.we_clk [7422]));
Q_ASSIGN U8969 ( .B(clk), .A(\g.we_clk [7421]));
Q_ASSIGN U8970 ( .B(clk), .A(\g.we_clk [7420]));
Q_ASSIGN U8971 ( .B(clk), .A(\g.we_clk [7419]));
Q_ASSIGN U8972 ( .B(clk), .A(\g.we_clk [7418]));
Q_ASSIGN U8973 ( .B(clk), .A(\g.we_clk [7417]));
Q_ASSIGN U8974 ( .B(clk), .A(\g.we_clk [7416]));
Q_ASSIGN U8975 ( .B(clk), .A(\g.we_clk [7415]));
Q_ASSIGN U8976 ( .B(clk), .A(\g.we_clk [7414]));
Q_ASSIGN U8977 ( .B(clk), .A(\g.we_clk [7413]));
Q_ASSIGN U8978 ( .B(clk), .A(\g.we_clk [7412]));
Q_ASSIGN U8979 ( .B(clk), .A(\g.we_clk [7411]));
Q_ASSIGN U8980 ( .B(clk), .A(\g.we_clk [7410]));
Q_ASSIGN U8981 ( .B(clk), .A(\g.we_clk [7409]));
Q_ASSIGN U8982 ( .B(clk), .A(\g.we_clk [7408]));
Q_ASSIGN U8983 ( .B(clk), .A(\g.we_clk [7407]));
Q_ASSIGN U8984 ( .B(clk), .A(\g.we_clk [7406]));
Q_ASSIGN U8985 ( .B(clk), .A(\g.we_clk [7405]));
Q_ASSIGN U8986 ( .B(clk), .A(\g.we_clk [7404]));
Q_ASSIGN U8987 ( .B(clk), .A(\g.we_clk [7403]));
Q_ASSIGN U8988 ( .B(clk), .A(\g.we_clk [7402]));
Q_ASSIGN U8989 ( .B(clk), .A(\g.we_clk [7401]));
Q_ASSIGN U8990 ( .B(clk), .A(\g.we_clk [7400]));
Q_ASSIGN U8991 ( .B(clk), .A(\g.we_clk [7399]));
Q_ASSIGN U8992 ( .B(clk), .A(\g.we_clk [7398]));
Q_ASSIGN U8993 ( .B(clk), .A(\g.we_clk [7397]));
Q_ASSIGN U8994 ( .B(clk), .A(\g.we_clk [7396]));
Q_ASSIGN U8995 ( .B(clk), .A(\g.we_clk [7395]));
Q_ASSIGN U8996 ( .B(clk), .A(\g.we_clk [7394]));
Q_ASSIGN U8997 ( .B(clk), .A(\g.we_clk [7393]));
Q_ASSIGN U8998 ( .B(clk), .A(\g.we_clk [7392]));
Q_ASSIGN U8999 ( .B(clk), .A(\g.we_clk [7391]));
Q_ASSIGN U9000 ( .B(clk), .A(\g.we_clk [7390]));
Q_ASSIGN U9001 ( .B(clk), .A(\g.we_clk [7389]));
Q_ASSIGN U9002 ( .B(clk), .A(\g.we_clk [7388]));
Q_ASSIGN U9003 ( .B(clk), .A(\g.we_clk [7387]));
Q_ASSIGN U9004 ( .B(clk), .A(\g.we_clk [7386]));
Q_ASSIGN U9005 ( .B(clk), .A(\g.we_clk [7385]));
Q_ASSIGN U9006 ( .B(clk), .A(\g.we_clk [7384]));
Q_ASSIGN U9007 ( .B(clk), .A(\g.we_clk [7383]));
Q_ASSIGN U9008 ( .B(clk), .A(\g.we_clk [7382]));
Q_ASSIGN U9009 ( .B(clk), .A(\g.we_clk [7381]));
Q_ASSIGN U9010 ( .B(clk), .A(\g.we_clk [7380]));
Q_ASSIGN U9011 ( .B(clk), .A(\g.we_clk [7379]));
Q_ASSIGN U9012 ( .B(clk), .A(\g.we_clk [7378]));
Q_ASSIGN U9013 ( .B(clk), .A(\g.we_clk [7377]));
Q_ASSIGN U9014 ( .B(clk), .A(\g.we_clk [7376]));
Q_ASSIGN U9015 ( .B(clk), .A(\g.we_clk [7375]));
Q_ASSIGN U9016 ( .B(clk), .A(\g.we_clk [7374]));
Q_ASSIGN U9017 ( .B(clk), .A(\g.we_clk [7373]));
Q_ASSIGN U9018 ( .B(clk), .A(\g.we_clk [7372]));
Q_ASSIGN U9019 ( .B(clk), .A(\g.we_clk [7371]));
Q_ASSIGN U9020 ( .B(clk), .A(\g.we_clk [7370]));
Q_ASSIGN U9021 ( .B(clk), .A(\g.we_clk [7369]));
Q_ASSIGN U9022 ( .B(clk), .A(\g.we_clk [7368]));
Q_ASSIGN U9023 ( .B(clk), .A(\g.we_clk [7367]));
Q_ASSIGN U9024 ( .B(clk), .A(\g.we_clk [7366]));
Q_ASSIGN U9025 ( .B(clk), .A(\g.we_clk [7365]));
Q_ASSIGN U9026 ( .B(clk), .A(\g.we_clk [7364]));
Q_ASSIGN U9027 ( .B(clk), .A(\g.we_clk [7363]));
Q_ASSIGN U9028 ( .B(clk), .A(\g.we_clk [7362]));
Q_ASSIGN U9029 ( .B(clk), .A(\g.we_clk [7361]));
Q_ASSIGN U9030 ( .B(clk), .A(\g.we_clk [7360]));
Q_ASSIGN U9031 ( .B(clk), .A(\g.we_clk [7359]));
Q_ASSIGN U9032 ( .B(clk), .A(\g.we_clk [7358]));
Q_ASSIGN U9033 ( .B(clk), .A(\g.we_clk [7357]));
Q_ASSIGN U9034 ( .B(clk), .A(\g.we_clk [7356]));
Q_ASSIGN U9035 ( .B(clk), .A(\g.we_clk [7355]));
Q_ASSIGN U9036 ( .B(clk), .A(\g.we_clk [7354]));
Q_ASSIGN U9037 ( .B(clk), .A(\g.we_clk [7353]));
Q_ASSIGN U9038 ( .B(clk), .A(\g.we_clk [7352]));
Q_ASSIGN U9039 ( .B(clk), .A(\g.we_clk [7351]));
Q_ASSIGN U9040 ( .B(clk), .A(\g.we_clk [7350]));
Q_ASSIGN U9041 ( .B(clk), .A(\g.we_clk [7349]));
Q_ASSIGN U9042 ( .B(clk), .A(\g.we_clk [7348]));
Q_ASSIGN U9043 ( .B(clk), .A(\g.we_clk [7347]));
Q_ASSIGN U9044 ( .B(clk), .A(\g.we_clk [7346]));
Q_ASSIGN U9045 ( .B(clk), .A(\g.we_clk [7345]));
Q_ASSIGN U9046 ( .B(clk), .A(\g.we_clk [7344]));
Q_ASSIGN U9047 ( .B(clk), .A(\g.we_clk [7343]));
Q_ASSIGN U9048 ( .B(clk), .A(\g.we_clk [7342]));
Q_ASSIGN U9049 ( .B(clk), .A(\g.we_clk [7341]));
Q_ASSIGN U9050 ( .B(clk), .A(\g.we_clk [7340]));
Q_ASSIGN U9051 ( .B(clk), .A(\g.we_clk [7339]));
Q_ASSIGN U9052 ( .B(clk), .A(\g.we_clk [7338]));
Q_ASSIGN U9053 ( .B(clk), .A(\g.we_clk [7337]));
Q_ASSIGN U9054 ( .B(clk), .A(\g.we_clk [7336]));
Q_ASSIGN U9055 ( .B(clk), .A(\g.we_clk [7335]));
Q_ASSIGN U9056 ( .B(clk), .A(\g.we_clk [7334]));
Q_ASSIGN U9057 ( .B(clk), .A(\g.we_clk [7333]));
Q_ASSIGN U9058 ( .B(clk), .A(\g.we_clk [7332]));
Q_ASSIGN U9059 ( .B(clk), .A(\g.we_clk [7331]));
Q_ASSIGN U9060 ( .B(clk), .A(\g.we_clk [7330]));
Q_ASSIGN U9061 ( .B(clk), .A(\g.we_clk [7329]));
Q_ASSIGN U9062 ( .B(clk), .A(\g.we_clk [7328]));
Q_ASSIGN U9063 ( .B(clk), .A(\g.we_clk [7327]));
Q_ASSIGN U9064 ( .B(clk), .A(\g.we_clk [7326]));
Q_ASSIGN U9065 ( .B(clk), .A(\g.we_clk [7325]));
Q_ASSIGN U9066 ( .B(clk), .A(\g.we_clk [7324]));
Q_ASSIGN U9067 ( .B(clk), .A(\g.we_clk [7323]));
Q_ASSIGN U9068 ( .B(clk), .A(\g.we_clk [7322]));
Q_ASSIGN U9069 ( .B(clk), .A(\g.we_clk [7321]));
Q_ASSIGN U9070 ( .B(clk), .A(\g.we_clk [7320]));
Q_ASSIGN U9071 ( .B(clk), .A(\g.we_clk [7319]));
Q_ASSIGN U9072 ( .B(clk), .A(\g.we_clk [7318]));
Q_ASSIGN U9073 ( .B(clk), .A(\g.we_clk [7317]));
Q_ASSIGN U9074 ( .B(clk), .A(\g.we_clk [7316]));
Q_ASSIGN U9075 ( .B(clk), .A(\g.we_clk [7315]));
Q_ASSIGN U9076 ( .B(clk), .A(\g.we_clk [7314]));
Q_ASSIGN U9077 ( .B(clk), .A(\g.we_clk [7313]));
Q_ASSIGN U9078 ( .B(clk), .A(\g.we_clk [7312]));
Q_ASSIGN U9079 ( .B(clk), .A(\g.we_clk [7311]));
Q_ASSIGN U9080 ( .B(clk), .A(\g.we_clk [7310]));
Q_ASSIGN U9081 ( .B(clk), .A(\g.we_clk [7309]));
Q_ASSIGN U9082 ( .B(clk), .A(\g.we_clk [7308]));
Q_ASSIGN U9083 ( .B(clk), .A(\g.we_clk [7307]));
Q_ASSIGN U9084 ( .B(clk), .A(\g.we_clk [7306]));
Q_ASSIGN U9085 ( .B(clk), .A(\g.we_clk [7305]));
Q_ASSIGN U9086 ( .B(clk), .A(\g.we_clk [7304]));
Q_ASSIGN U9087 ( .B(clk), .A(\g.we_clk [7303]));
Q_ASSIGN U9088 ( .B(clk), .A(\g.we_clk [7302]));
Q_ASSIGN U9089 ( .B(clk), .A(\g.we_clk [7301]));
Q_ASSIGN U9090 ( .B(clk), .A(\g.we_clk [7300]));
Q_ASSIGN U9091 ( .B(clk), .A(\g.we_clk [7299]));
Q_ASSIGN U9092 ( .B(clk), .A(\g.we_clk [7298]));
Q_ASSIGN U9093 ( .B(clk), .A(\g.we_clk [7297]));
Q_ASSIGN U9094 ( .B(clk), .A(\g.we_clk [7296]));
Q_ASSIGN U9095 ( .B(clk), .A(\g.we_clk [7295]));
Q_ASSIGN U9096 ( .B(clk), .A(\g.we_clk [7294]));
Q_ASSIGN U9097 ( .B(clk), .A(\g.we_clk [7293]));
Q_ASSIGN U9098 ( .B(clk), .A(\g.we_clk [7292]));
Q_ASSIGN U9099 ( .B(clk), .A(\g.we_clk [7291]));
Q_ASSIGN U9100 ( .B(clk), .A(\g.we_clk [7290]));
Q_ASSIGN U9101 ( .B(clk), .A(\g.we_clk [7289]));
Q_ASSIGN U9102 ( .B(clk), .A(\g.we_clk [7288]));
Q_ASSIGN U9103 ( .B(clk), .A(\g.we_clk [7287]));
Q_ASSIGN U9104 ( .B(clk), .A(\g.we_clk [7286]));
Q_ASSIGN U9105 ( .B(clk), .A(\g.we_clk [7285]));
Q_ASSIGN U9106 ( .B(clk), .A(\g.we_clk [7284]));
Q_ASSIGN U9107 ( .B(clk), .A(\g.we_clk [7283]));
Q_ASSIGN U9108 ( .B(clk), .A(\g.we_clk [7282]));
Q_ASSIGN U9109 ( .B(clk), .A(\g.we_clk [7281]));
Q_ASSIGN U9110 ( .B(clk), .A(\g.we_clk [7280]));
Q_ASSIGN U9111 ( .B(clk), .A(\g.we_clk [7279]));
Q_ASSIGN U9112 ( .B(clk), .A(\g.we_clk [7278]));
Q_ASSIGN U9113 ( .B(clk), .A(\g.we_clk [7277]));
Q_ASSIGN U9114 ( .B(clk), .A(\g.we_clk [7276]));
Q_ASSIGN U9115 ( .B(clk), .A(\g.we_clk [7275]));
Q_ASSIGN U9116 ( .B(clk), .A(\g.we_clk [7274]));
Q_ASSIGN U9117 ( .B(clk), .A(\g.we_clk [7273]));
Q_ASSIGN U9118 ( .B(clk), .A(\g.we_clk [7272]));
Q_ASSIGN U9119 ( .B(clk), .A(\g.we_clk [7271]));
Q_ASSIGN U9120 ( .B(clk), .A(\g.we_clk [7270]));
Q_ASSIGN U9121 ( .B(clk), .A(\g.we_clk [7269]));
Q_ASSIGN U9122 ( .B(clk), .A(\g.we_clk [7268]));
Q_ASSIGN U9123 ( .B(clk), .A(\g.we_clk [7267]));
Q_ASSIGN U9124 ( .B(clk), .A(\g.we_clk [7266]));
Q_ASSIGN U9125 ( .B(clk), .A(\g.we_clk [7265]));
Q_ASSIGN U9126 ( .B(clk), .A(\g.we_clk [7264]));
Q_ASSIGN U9127 ( .B(clk), .A(\g.we_clk [7263]));
Q_ASSIGN U9128 ( .B(clk), .A(\g.we_clk [7262]));
Q_ASSIGN U9129 ( .B(clk), .A(\g.we_clk [7261]));
Q_ASSIGN U9130 ( .B(clk), .A(\g.we_clk [7260]));
Q_ASSIGN U9131 ( .B(clk), .A(\g.we_clk [7259]));
Q_ASSIGN U9132 ( .B(clk), .A(\g.we_clk [7258]));
Q_ASSIGN U9133 ( .B(clk), .A(\g.we_clk [7257]));
Q_ASSIGN U9134 ( .B(clk), .A(\g.we_clk [7256]));
Q_ASSIGN U9135 ( .B(clk), .A(\g.we_clk [7255]));
Q_ASSIGN U9136 ( .B(clk), .A(\g.we_clk [7254]));
Q_ASSIGN U9137 ( .B(clk), .A(\g.we_clk [7253]));
Q_ASSIGN U9138 ( .B(clk), .A(\g.we_clk [7252]));
Q_ASSIGN U9139 ( .B(clk), .A(\g.we_clk [7251]));
Q_ASSIGN U9140 ( .B(clk), .A(\g.we_clk [7250]));
Q_ASSIGN U9141 ( .B(clk), .A(\g.we_clk [7249]));
Q_ASSIGN U9142 ( .B(clk), .A(\g.we_clk [7248]));
Q_ASSIGN U9143 ( .B(clk), .A(\g.we_clk [7247]));
Q_ASSIGN U9144 ( .B(clk), .A(\g.we_clk [7246]));
Q_ASSIGN U9145 ( .B(clk), .A(\g.we_clk [7245]));
Q_ASSIGN U9146 ( .B(clk), .A(\g.we_clk [7244]));
Q_ASSIGN U9147 ( .B(clk), .A(\g.we_clk [7243]));
Q_ASSIGN U9148 ( .B(clk), .A(\g.we_clk [7242]));
Q_ASSIGN U9149 ( .B(clk), .A(\g.we_clk [7241]));
Q_ASSIGN U9150 ( .B(clk), .A(\g.we_clk [7240]));
Q_ASSIGN U9151 ( .B(clk), .A(\g.we_clk [7239]));
Q_ASSIGN U9152 ( .B(clk), .A(\g.we_clk [7238]));
Q_ASSIGN U9153 ( .B(clk), .A(\g.we_clk [7237]));
Q_ASSIGN U9154 ( .B(clk), .A(\g.we_clk [7236]));
Q_ASSIGN U9155 ( .B(clk), .A(\g.we_clk [7235]));
Q_ASSIGN U9156 ( .B(clk), .A(\g.we_clk [7234]));
Q_ASSIGN U9157 ( .B(clk), .A(\g.we_clk [7233]));
Q_ASSIGN U9158 ( .B(clk), .A(\g.we_clk [7232]));
Q_ASSIGN U9159 ( .B(clk), .A(\g.we_clk [7231]));
Q_ASSIGN U9160 ( .B(clk), .A(\g.we_clk [7230]));
Q_ASSIGN U9161 ( .B(clk), .A(\g.we_clk [7229]));
Q_ASSIGN U9162 ( .B(clk), .A(\g.we_clk [7228]));
Q_ASSIGN U9163 ( .B(clk), .A(\g.we_clk [7227]));
Q_ASSIGN U9164 ( .B(clk), .A(\g.we_clk [7226]));
Q_ASSIGN U9165 ( .B(clk), .A(\g.we_clk [7225]));
Q_ASSIGN U9166 ( .B(clk), .A(\g.we_clk [7224]));
Q_ASSIGN U9167 ( .B(clk), .A(\g.we_clk [7223]));
Q_ASSIGN U9168 ( .B(clk), .A(\g.we_clk [7222]));
Q_ASSIGN U9169 ( .B(clk), .A(\g.we_clk [7221]));
Q_ASSIGN U9170 ( .B(clk), .A(\g.we_clk [7220]));
Q_ASSIGN U9171 ( .B(clk), .A(\g.we_clk [7219]));
Q_ASSIGN U9172 ( .B(clk), .A(\g.we_clk [7218]));
Q_ASSIGN U9173 ( .B(clk), .A(\g.we_clk [7217]));
Q_ASSIGN U9174 ( .B(clk), .A(\g.we_clk [7216]));
Q_ASSIGN U9175 ( .B(clk), .A(\g.we_clk [7215]));
Q_ASSIGN U9176 ( .B(clk), .A(\g.we_clk [7214]));
Q_ASSIGN U9177 ( .B(clk), .A(\g.we_clk [7213]));
Q_ASSIGN U9178 ( .B(clk), .A(\g.we_clk [7212]));
Q_ASSIGN U9179 ( .B(clk), .A(\g.we_clk [7211]));
Q_ASSIGN U9180 ( .B(clk), .A(\g.we_clk [7210]));
Q_ASSIGN U9181 ( .B(clk), .A(\g.we_clk [7209]));
Q_ASSIGN U9182 ( .B(clk), .A(\g.we_clk [7208]));
Q_ASSIGN U9183 ( .B(clk), .A(\g.we_clk [7207]));
Q_ASSIGN U9184 ( .B(clk), .A(\g.we_clk [7206]));
Q_ASSIGN U9185 ( .B(clk), .A(\g.we_clk [7205]));
Q_ASSIGN U9186 ( .B(clk), .A(\g.we_clk [7204]));
Q_ASSIGN U9187 ( .B(clk), .A(\g.we_clk [7203]));
Q_ASSIGN U9188 ( .B(clk), .A(\g.we_clk [7202]));
Q_ASSIGN U9189 ( .B(clk), .A(\g.we_clk [7201]));
Q_ASSIGN U9190 ( .B(clk), .A(\g.we_clk [7200]));
Q_ASSIGN U9191 ( .B(clk), .A(\g.we_clk [7199]));
Q_ASSIGN U9192 ( .B(clk), .A(\g.we_clk [7198]));
Q_ASSIGN U9193 ( .B(clk), .A(\g.we_clk [7197]));
Q_ASSIGN U9194 ( .B(clk), .A(\g.we_clk [7196]));
Q_ASSIGN U9195 ( .B(clk), .A(\g.we_clk [7195]));
Q_ASSIGN U9196 ( .B(clk), .A(\g.we_clk [7194]));
Q_ASSIGN U9197 ( .B(clk), .A(\g.we_clk [7193]));
Q_ASSIGN U9198 ( .B(clk), .A(\g.we_clk [7192]));
Q_ASSIGN U9199 ( .B(clk), .A(\g.we_clk [7191]));
Q_ASSIGN U9200 ( .B(clk), .A(\g.we_clk [7190]));
Q_ASSIGN U9201 ( .B(clk), .A(\g.we_clk [7189]));
Q_ASSIGN U9202 ( .B(clk), .A(\g.we_clk [7188]));
Q_ASSIGN U9203 ( .B(clk), .A(\g.we_clk [7187]));
Q_ASSIGN U9204 ( .B(clk), .A(\g.we_clk [7186]));
Q_ASSIGN U9205 ( .B(clk), .A(\g.we_clk [7185]));
Q_ASSIGN U9206 ( .B(clk), .A(\g.we_clk [7184]));
Q_ASSIGN U9207 ( .B(clk), .A(\g.we_clk [7183]));
Q_ASSIGN U9208 ( .B(clk), .A(\g.we_clk [7182]));
Q_ASSIGN U9209 ( .B(clk), .A(\g.we_clk [7181]));
Q_ASSIGN U9210 ( .B(clk), .A(\g.we_clk [7180]));
Q_ASSIGN U9211 ( .B(clk), .A(\g.we_clk [7179]));
Q_ASSIGN U9212 ( .B(clk), .A(\g.we_clk [7178]));
Q_ASSIGN U9213 ( .B(clk), .A(\g.we_clk [7177]));
Q_ASSIGN U9214 ( .B(clk), .A(\g.we_clk [7176]));
Q_ASSIGN U9215 ( .B(clk), .A(\g.we_clk [7175]));
Q_ASSIGN U9216 ( .B(clk), .A(\g.we_clk [7174]));
Q_ASSIGN U9217 ( .B(clk), .A(\g.we_clk [7173]));
Q_ASSIGN U9218 ( .B(clk), .A(\g.we_clk [7172]));
Q_ASSIGN U9219 ( .B(clk), .A(\g.we_clk [7171]));
Q_ASSIGN U9220 ( .B(clk), .A(\g.we_clk [7170]));
Q_ASSIGN U9221 ( .B(clk), .A(\g.we_clk [7169]));
Q_ASSIGN U9222 ( .B(clk), .A(\g.we_clk [7168]));
Q_ASSIGN U9223 ( .B(clk), .A(\g.we_clk [7167]));
Q_ASSIGN U9224 ( .B(clk), .A(\g.we_clk [7166]));
Q_ASSIGN U9225 ( .B(clk), .A(\g.we_clk [7165]));
Q_ASSIGN U9226 ( .B(clk), .A(\g.we_clk [7164]));
Q_ASSIGN U9227 ( .B(clk), .A(\g.we_clk [7163]));
Q_ASSIGN U9228 ( .B(clk), .A(\g.we_clk [7162]));
Q_ASSIGN U9229 ( .B(clk), .A(\g.we_clk [7161]));
Q_ASSIGN U9230 ( .B(clk), .A(\g.we_clk [7160]));
Q_ASSIGN U9231 ( .B(clk), .A(\g.we_clk [7159]));
Q_ASSIGN U9232 ( .B(clk), .A(\g.we_clk [7158]));
Q_ASSIGN U9233 ( .B(clk), .A(\g.we_clk [7157]));
Q_ASSIGN U9234 ( .B(clk), .A(\g.we_clk [7156]));
Q_ASSIGN U9235 ( .B(clk), .A(\g.we_clk [7155]));
Q_ASSIGN U9236 ( .B(clk), .A(\g.we_clk [7154]));
Q_ASSIGN U9237 ( .B(clk), .A(\g.we_clk [7153]));
Q_ASSIGN U9238 ( .B(clk), .A(\g.we_clk [7152]));
Q_ASSIGN U9239 ( .B(clk), .A(\g.we_clk [7151]));
Q_ASSIGN U9240 ( .B(clk), .A(\g.we_clk [7150]));
Q_ASSIGN U9241 ( .B(clk), .A(\g.we_clk [7149]));
Q_ASSIGN U9242 ( .B(clk), .A(\g.we_clk [7148]));
Q_ASSIGN U9243 ( .B(clk), .A(\g.we_clk [7147]));
Q_ASSIGN U9244 ( .B(clk), .A(\g.we_clk [7146]));
Q_ASSIGN U9245 ( .B(clk), .A(\g.we_clk [7145]));
Q_ASSIGN U9246 ( .B(clk), .A(\g.we_clk [7144]));
Q_ASSIGN U9247 ( .B(clk), .A(\g.we_clk [7143]));
Q_ASSIGN U9248 ( .B(clk), .A(\g.we_clk [7142]));
Q_ASSIGN U9249 ( .B(clk), .A(\g.we_clk [7141]));
Q_ASSIGN U9250 ( .B(clk), .A(\g.we_clk [7140]));
Q_ASSIGN U9251 ( .B(clk), .A(\g.we_clk [7139]));
Q_ASSIGN U9252 ( .B(clk), .A(\g.we_clk [7138]));
Q_ASSIGN U9253 ( .B(clk), .A(\g.we_clk [7137]));
Q_ASSIGN U9254 ( .B(clk), .A(\g.we_clk [7136]));
Q_ASSIGN U9255 ( .B(clk), .A(\g.we_clk [7135]));
Q_ASSIGN U9256 ( .B(clk), .A(\g.we_clk [7134]));
Q_ASSIGN U9257 ( .B(clk), .A(\g.we_clk [7133]));
Q_ASSIGN U9258 ( .B(clk), .A(\g.we_clk [7132]));
Q_ASSIGN U9259 ( .B(clk), .A(\g.we_clk [7131]));
Q_ASSIGN U9260 ( .B(clk), .A(\g.we_clk [7130]));
Q_ASSIGN U9261 ( .B(clk), .A(\g.we_clk [7129]));
Q_ASSIGN U9262 ( .B(clk), .A(\g.we_clk [7128]));
Q_ASSIGN U9263 ( .B(clk), .A(\g.we_clk [7127]));
Q_ASSIGN U9264 ( .B(clk), .A(\g.we_clk [7126]));
Q_ASSIGN U9265 ( .B(clk), .A(\g.we_clk [7125]));
Q_ASSIGN U9266 ( .B(clk), .A(\g.we_clk [7124]));
Q_ASSIGN U9267 ( .B(clk), .A(\g.we_clk [7123]));
Q_ASSIGN U9268 ( .B(clk), .A(\g.we_clk [7122]));
Q_ASSIGN U9269 ( .B(clk), .A(\g.we_clk [7121]));
Q_ASSIGN U9270 ( .B(clk), .A(\g.we_clk [7120]));
Q_ASSIGN U9271 ( .B(clk), .A(\g.we_clk [7119]));
Q_ASSIGN U9272 ( .B(clk), .A(\g.we_clk [7118]));
Q_ASSIGN U9273 ( .B(clk), .A(\g.we_clk [7117]));
Q_ASSIGN U9274 ( .B(clk), .A(\g.we_clk [7116]));
Q_ASSIGN U9275 ( .B(clk), .A(\g.we_clk [7115]));
Q_ASSIGN U9276 ( .B(clk), .A(\g.we_clk [7114]));
Q_ASSIGN U9277 ( .B(clk), .A(\g.we_clk [7113]));
Q_ASSIGN U9278 ( .B(clk), .A(\g.we_clk [7112]));
Q_ASSIGN U9279 ( .B(clk), .A(\g.we_clk [7111]));
Q_ASSIGN U9280 ( .B(clk), .A(\g.we_clk [7110]));
Q_ASSIGN U9281 ( .B(clk), .A(\g.we_clk [7109]));
Q_ASSIGN U9282 ( .B(clk), .A(\g.we_clk [7108]));
Q_ASSIGN U9283 ( .B(clk), .A(\g.we_clk [7107]));
Q_ASSIGN U9284 ( .B(clk), .A(\g.we_clk [7106]));
Q_ASSIGN U9285 ( .B(clk), .A(\g.we_clk [7105]));
Q_ASSIGN U9286 ( .B(clk), .A(\g.we_clk [7104]));
Q_ASSIGN U9287 ( .B(clk), .A(\g.we_clk [7103]));
Q_ASSIGN U9288 ( .B(clk), .A(\g.we_clk [7102]));
Q_ASSIGN U9289 ( .B(clk), .A(\g.we_clk [7101]));
Q_ASSIGN U9290 ( .B(clk), .A(\g.we_clk [7100]));
Q_ASSIGN U9291 ( .B(clk), .A(\g.we_clk [7099]));
Q_ASSIGN U9292 ( .B(clk), .A(\g.we_clk [7098]));
Q_ASSIGN U9293 ( .B(clk), .A(\g.we_clk [7097]));
Q_ASSIGN U9294 ( .B(clk), .A(\g.we_clk [7096]));
Q_ASSIGN U9295 ( .B(clk), .A(\g.we_clk [7095]));
Q_ASSIGN U9296 ( .B(clk), .A(\g.we_clk [7094]));
Q_ASSIGN U9297 ( .B(clk), .A(\g.we_clk [7093]));
Q_ASSIGN U9298 ( .B(clk), .A(\g.we_clk [7092]));
Q_ASSIGN U9299 ( .B(clk), .A(\g.we_clk [7091]));
Q_ASSIGN U9300 ( .B(clk), .A(\g.we_clk [7090]));
Q_ASSIGN U9301 ( .B(clk), .A(\g.we_clk [7089]));
Q_ASSIGN U9302 ( .B(clk), .A(\g.we_clk [7088]));
Q_ASSIGN U9303 ( .B(clk), .A(\g.we_clk [7087]));
Q_ASSIGN U9304 ( .B(clk), .A(\g.we_clk [7086]));
Q_ASSIGN U9305 ( .B(clk), .A(\g.we_clk [7085]));
Q_ASSIGN U9306 ( .B(clk), .A(\g.we_clk [7084]));
Q_ASSIGN U9307 ( .B(clk), .A(\g.we_clk [7083]));
Q_ASSIGN U9308 ( .B(clk), .A(\g.we_clk [7082]));
Q_ASSIGN U9309 ( .B(clk), .A(\g.we_clk [7081]));
Q_ASSIGN U9310 ( .B(clk), .A(\g.we_clk [7080]));
Q_ASSIGN U9311 ( .B(clk), .A(\g.we_clk [7079]));
Q_ASSIGN U9312 ( .B(clk), .A(\g.we_clk [7078]));
Q_ASSIGN U9313 ( .B(clk), .A(\g.we_clk [7077]));
Q_ASSIGN U9314 ( .B(clk), .A(\g.we_clk [7076]));
Q_ASSIGN U9315 ( .B(clk), .A(\g.we_clk [7075]));
Q_ASSIGN U9316 ( .B(clk), .A(\g.we_clk [7074]));
Q_ASSIGN U9317 ( .B(clk), .A(\g.we_clk [7073]));
Q_ASSIGN U9318 ( .B(clk), .A(\g.we_clk [7072]));
Q_ASSIGN U9319 ( .B(clk), .A(\g.we_clk [7071]));
Q_ASSIGN U9320 ( .B(clk), .A(\g.we_clk [7070]));
Q_ASSIGN U9321 ( .B(clk), .A(\g.we_clk [7069]));
Q_ASSIGN U9322 ( .B(clk), .A(\g.we_clk [7068]));
Q_ASSIGN U9323 ( .B(clk), .A(\g.we_clk [7067]));
Q_ASSIGN U9324 ( .B(clk), .A(\g.we_clk [7066]));
Q_ASSIGN U9325 ( .B(clk), .A(\g.we_clk [7065]));
Q_ASSIGN U9326 ( .B(clk), .A(\g.we_clk [7064]));
Q_ASSIGN U9327 ( .B(clk), .A(\g.we_clk [7063]));
Q_ASSIGN U9328 ( .B(clk), .A(\g.we_clk [7062]));
Q_ASSIGN U9329 ( .B(clk), .A(\g.we_clk [7061]));
Q_ASSIGN U9330 ( .B(clk), .A(\g.we_clk [7060]));
Q_ASSIGN U9331 ( .B(clk), .A(\g.we_clk [7059]));
Q_ASSIGN U9332 ( .B(clk), .A(\g.we_clk [7058]));
Q_ASSIGN U9333 ( .B(clk), .A(\g.we_clk [7057]));
Q_ASSIGN U9334 ( .B(clk), .A(\g.we_clk [7056]));
Q_ASSIGN U9335 ( .B(clk), .A(\g.we_clk [7055]));
Q_ASSIGN U9336 ( .B(clk), .A(\g.we_clk [7054]));
Q_ASSIGN U9337 ( .B(clk), .A(\g.we_clk [7053]));
Q_ASSIGN U9338 ( .B(clk), .A(\g.we_clk [7052]));
Q_ASSIGN U9339 ( .B(clk), .A(\g.we_clk [7051]));
Q_ASSIGN U9340 ( .B(clk), .A(\g.we_clk [7050]));
Q_ASSIGN U9341 ( .B(clk), .A(\g.we_clk [7049]));
Q_ASSIGN U9342 ( .B(clk), .A(\g.we_clk [7048]));
Q_ASSIGN U9343 ( .B(clk), .A(\g.we_clk [7047]));
Q_ASSIGN U9344 ( .B(clk), .A(\g.we_clk [7046]));
Q_ASSIGN U9345 ( .B(clk), .A(\g.we_clk [7045]));
Q_ASSIGN U9346 ( .B(clk), .A(\g.we_clk [7044]));
Q_ASSIGN U9347 ( .B(clk), .A(\g.we_clk [7043]));
Q_ASSIGN U9348 ( .B(clk), .A(\g.we_clk [7042]));
Q_ASSIGN U9349 ( .B(clk), .A(\g.we_clk [7041]));
Q_ASSIGN U9350 ( .B(clk), .A(\g.we_clk [7040]));
Q_ASSIGN U9351 ( .B(clk), .A(\g.we_clk [7039]));
Q_ASSIGN U9352 ( .B(clk), .A(\g.we_clk [7038]));
Q_ASSIGN U9353 ( .B(clk), .A(\g.we_clk [7037]));
Q_ASSIGN U9354 ( .B(clk), .A(\g.we_clk [7036]));
Q_ASSIGN U9355 ( .B(clk), .A(\g.we_clk [7035]));
Q_ASSIGN U9356 ( .B(clk), .A(\g.we_clk [7034]));
Q_ASSIGN U9357 ( .B(clk), .A(\g.we_clk [7033]));
Q_ASSIGN U9358 ( .B(clk), .A(\g.we_clk [7032]));
Q_ASSIGN U9359 ( .B(clk), .A(\g.we_clk [7031]));
Q_ASSIGN U9360 ( .B(clk), .A(\g.we_clk [7030]));
Q_ASSIGN U9361 ( .B(clk), .A(\g.we_clk [7029]));
Q_ASSIGN U9362 ( .B(clk), .A(\g.we_clk [7028]));
Q_ASSIGN U9363 ( .B(clk), .A(\g.we_clk [7027]));
Q_ASSIGN U9364 ( .B(clk), .A(\g.we_clk [7026]));
Q_ASSIGN U9365 ( .B(clk), .A(\g.we_clk [7025]));
Q_ASSIGN U9366 ( .B(clk), .A(\g.we_clk [7024]));
Q_ASSIGN U9367 ( .B(clk), .A(\g.we_clk [7023]));
Q_ASSIGN U9368 ( .B(clk), .A(\g.we_clk [7022]));
Q_ASSIGN U9369 ( .B(clk), .A(\g.we_clk [7021]));
Q_ASSIGN U9370 ( .B(clk), .A(\g.we_clk [7020]));
Q_ASSIGN U9371 ( .B(clk), .A(\g.we_clk [7019]));
Q_ASSIGN U9372 ( .B(clk), .A(\g.we_clk [7018]));
Q_ASSIGN U9373 ( .B(clk), .A(\g.we_clk [7017]));
Q_ASSIGN U9374 ( .B(clk), .A(\g.we_clk [7016]));
Q_ASSIGN U9375 ( .B(clk), .A(\g.we_clk [7015]));
Q_ASSIGN U9376 ( .B(clk), .A(\g.we_clk [7014]));
Q_ASSIGN U9377 ( .B(clk), .A(\g.we_clk [7013]));
Q_ASSIGN U9378 ( .B(clk), .A(\g.we_clk [7012]));
Q_ASSIGN U9379 ( .B(clk), .A(\g.we_clk [7011]));
Q_ASSIGN U9380 ( .B(clk), .A(\g.we_clk [7010]));
Q_ASSIGN U9381 ( .B(clk), .A(\g.we_clk [7009]));
Q_ASSIGN U9382 ( .B(clk), .A(\g.we_clk [7008]));
Q_ASSIGN U9383 ( .B(clk), .A(\g.we_clk [7007]));
Q_ASSIGN U9384 ( .B(clk), .A(\g.we_clk [7006]));
Q_ASSIGN U9385 ( .B(clk), .A(\g.we_clk [7005]));
Q_ASSIGN U9386 ( .B(clk), .A(\g.we_clk [7004]));
Q_ASSIGN U9387 ( .B(clk), .A(\g.we_clk [7003]));
Q_ASSIGN U9388 ( .B(clk), .A(\g.we_clk [7002]));
Q_ASSIGN U9389 ( .B(clk), .A(\g.we_clk [7001]));
Q_ASSIGN U9390 ( .B(clk), .A(\g.we_clk [7000]));
Q_ASSIGN U9391 ( .B(clk), .A(\g.we_clk [6999]));
Q_ASSIGN U9392 ( .B(clk), .A(\g.we_clk [6998]));
Q_ASSIGN U9393 ( .B(clk), .A(\g.we_clk [6997]));
Q_ASSIGN U9394 ( .B(clk), .A(\g.we_clk [6996]));
Q_ASSIGN U9395 ( .B(clk), .A(\g.we_clk [6995]));
Q_ASSIGN U9396 ( .B(clk), .A(\g.we_clk [6994]));
Q_ASSIGN U9397 ( .B(clk), .A(\g.we_clk [6993]));
Q_ASSIGN U9398 ( .B(clk), .A(\g.we_clk [6992]));
Q_ASSIGN U9399 ( .B(clk), .A(\g.we_clk [6991]));
Q_ASSIGN U9400 ( .B(clk), .A(\g.we_clk [6990]));
Q_ASSIGN U9401 ( .B(clk), .A(\g.we_clk [6989]));
Q_ASSIGN U9402 ( .B(clk), .A(\g.we_clk [6988]));
Q_ASSIGN U9403 ( .B(clk), .A(\g.we_clk [6987]));
Q_ASSIGN U9404 ( .B(clk), .A(\g.we_clk [6986]));
Q_ASSIGN U9405 ( .B(clk), .A(\g.we_clk [6985]));
Q_ASSIGN U9406 ( .B(clk), .A(\g.we_clk [6984]));
Q_ASSIGN U9407 ( .B(clk), .A(\g.we_clk [6983]));
Q_ASSIGN U9408 ( .B(clk), .A(\g.we_clk [6982]));
Q_ASSIGN U9409 ( .B(clk), .A(\g.we_clk [6981]));
Q_ASSIGN U9410 ( .B(clk), .A(\g.we_clk [6980]));
Q_ASSIGN U9411 ( .B(clk), .A(\g.we_clk [6979]));
Q_ASSIGN U9412 ( .B(clk), .A(\g.we_clk [6978]));
Q_ASSIGN U9413 ( .B(clk), .A(\g.we_clk [6977]));
Q_ASSIGN U9414 ( .B(clk), .A(\g.we_clk [6976]));
Q_ASSIGN U9415 ( .B(clk), .A(\g.we_clk [6975]));
Q_ASSIGN U9416 ( .B(clk), .A(\g.we_clk [6974]));
Q_ASSIGN U9417 ( .B(clk), .A(\g.we_clk [6973]));
Q_ASSIGN U9418 ( .B(clk), .A(\g.we_clk [6972]));
Q_ASSIGN U9419 ( .B(clk), .A(\g.we_clk [6971]));
Q_ASSIGN U9420 ( .B(clk), .A(\g.we_clk [6970]));
Q_ASSIGN U9421 ( .B(clk), .A(\g.we_clk [6969]));
Q_ASSIGN U9422 ( .B(clk), .A(\g.we_clk [6968]));
Q_ASSIGN U9423 ( .B(clk), .A(\g.we_clk [6967]));
Q_ASSIGN U9424 ( .B(clk), .A(\g.we_clk [6966]));
Q_ASSIGN U9425 ( .B(clk), .A(\g.we_clk [6965]));
Q_ASSIGN U9426 ( .B(clk), .A(\g.we_clk [6964]));
Q_ASSIGN U9427 ( .B(clk), .A(\g.we_clk [6963]));
Q_ASSIGN U9428 ( .B(clk), .A(\g.we_clk [6962]));
Q_ASSIGN U9429 ( .B(clk), .A(\g.we_clk [6961]));
Q_ASSIGN U9430 ( .B(clk), .A(\g.we_clk [6960]));
Q_ASSIGN U9431 ( .B(clk), .A(\g.we_clk [6959]));
Q_ASSIGN U9432 ( .B(clk), .A(\g.we_clk [6958]));
Q_ASSIGN U9433 ( .B(clk), .A(\g.we_clk [6957]));
Q_ASSIGN U9434 ( .B(clk), .A(\g.we_clk [6956]));
Q_ASSIGN U9435 ( .B(clk), .A(\g.we_clk [6955]));
Q_ASSIGN U9436 ( .B(clk), .A(\g.we_clk [6954]));
Q_ASSIGN U9437 ( .B(clk), .A(\g.we_clk [6953]));
Q_ASSIGN U9438 ( .B(clk), .A(\g.we_clk [6952]));
Q_ASSIGN U9439 ( .B(clk), .A(\g.we_clk [6951]));
Q_ASSIGN U9440 ( .B(clk), .A(\g.we_clk [6950]));
Q_ASSIGN U9441 ( .B(clk), .A(\g.we_clk [6949]));
Q_ASSIGN U9442 ( .B(clk), .A(\g.we_clk [6948]));
Q_ASSIGN U9443 ( .B(clk), .A(\g.we_clk [6947]));
Q_ASSIGN U9444 ( .B(clk), .A(\g.we_clk [6946]));
Q_ASSIGN U9445 ( .B(clk), .A(\g.we_clk [6945]));
Q_ASSIGN U9446 ( .B(clk), .A(\g.we_clk [6944]));
Q_ASSIGN U9447 ( .B(clk), .A(\g.we_clk [6943]));
Q_ASSIGN U9448 ( .B(clk), .A(\g.we_clk [6942]));
Q_ASSIGN U9449 ( .B(clk), .A(\g.we_clk [6941]));
Q_ASSIGN U9450 ( .B(clk), .A(\g.we_clk [6940]));
Q_ASSIGN U9451 ( .B(clk), .A(\g.we_clk [6939]));
Q_ASSIGN U9452 ( .B(clk), .A(\g.we_clk [6938]));
Q_ASSIGN U9453 ( .B(clk), .A(\g.we_clk [6937]));
Q_ASSIGN U9454 ( .B(clk), .A(\g.we_clk [6936]));
Q_ASSIGN U9455 ( .B(clk), .A(\g.we_clk [6935]));
Q_ASSIGN U9456 ( .B(clk), .A(\g.we_clk [6934]));
Q_ASSIGN U9457 ( .B(clk), .A(\g.we_clk [6933]));
Q_ASSIGN U9458 ( .B(clk), .A(\g.we_clk [6932]));
Q_ASSIGN U9459 ( .B(clk), .A(\g.we_clk [6931]));
Q_ASSIGN U9460 ( .B(clk), .A(\g.we_clk [6930]));
Q_ASSIGN U9461 ( .B(clk), .A(\g.we_clk [6929]));
Q_ASSIGN U9462 ( .B(clk), .A(\g.we_clk [6928]));
Q_ASSIGN U9463 ( .B(clk), .A(\g.we_clk [6927]));
Q_ASSIGN U9464 ( .B(clk), .A(\g.we_clk [6926]));
Q_ASSIGN U9465 ( .B(clk), .A(\g.we_clk [6925]));
Q_ASSIGN U9466 ( .B(clk), .A(\g.we_clk [6924]));
Q_ASSIGN U9467 ( .B(clk), .A(\g.we_clk [6923]));
Q_ASSIGN U9468 ( .B(clk), .A(\g.we_clk [6922]));
Q_ASSIGN U9469 ( .B(clk), .A(\g.we_clk [6921]));
Q_ASSIGN U9470 ( .B(clk), .A(\g.we_clk [6920]));
Q_ASSIGN U9471 ( .B(clk), .A(\g.we_clk [6919]));
Q_ASSIGN U9472 ( .B(clk), .A(\g.we_clk [6918]));
Q_ASSIGN U9473 ( .B(clk), .A(\g.we_clk [6917]));
Q_ASSIGN U9474 ( .B(clk), .A(\g.we_clk [6916]));
Q_ASSIGN U9475 ( .B(clk), .A(\g.we_clk [6915]));
Q_ASSIGN U9476 ( .B(clk), .A(\g.we_clk [6914]));
Q_ASSIGN U9477 ( .B(clk), .A(\g.we_clk [6913]));
Q_ASSIGN U9478 ( .B(clk), .A(\g.we_clk [6912]));
Q_ASSIGN U9479 ( .B(clk), .A(\g.we_clk [6911]));
Q_ASSIGN U9480 ( .B(clk), .A(\g.we_clk [6910]));
Q_ASSIGN U9481 ( .B(clk), .A(\g.we_clk [6909]));
Q_ASSIGN U9482 ( .B(clk), .A(\g.we_clk [6908]));
Q_ASSIGN U9483 ( .B(clk), .A(\g.we_clk [6907]));
Q_ASSIGN U9484 ( .B(clk), .A(\g.we_clk [6906]));
Q_ASSIGN U9485 ( .B(clk), .A(\g.we_clk [6905]));
Q_ASSIGN U9486 ( .B(clk), .A(\g.we_clk [6904]));
Q_ASSIGN U9487 ( .B(clk), .A(\g.we_clk [6903]));
Q_ASSIGN U9488 ( .B(clk), .A(\g.we_clk [6902]));
Q_ASSIGN U9489 ( .B(clk), .A(\g.we_clk [6901]));
Q_ASSIGN U9490 ( .B(clk), .A(\g.we_clk [6900]));
Q_ASSIGN U9491 ( .B(clk), .A(\g.we_clk [6899]));
Q_ASSIGN U9492 ( .B(clk), .A(\g.we_clk [6898]));
Q_ASSIGN U9493 ( .B(clk), .A(\g.we_clk [6897]));
Q_ASSIGN U9494 ( .B(clk), .A(\g.we_clk [6896]));
Q_ASSIGN U9495 ( .B(clk), .A(\g.we_clk [6895]));
Q_ASSIGN U9496 ( .B(clk), .A(\g.we_clk [6894]));
Q_ASSIGN U9497 ( .B(clk), .A(\g.we_clk [6893]));
Q_ASSIGN U9498 ( .B(clk), .A(\g.we_clk [6892]));
Q_ASSIGN U9499 ( .B(clk), .A(\g.we_clk [6891]));
Q_ASSIGN U9500 ( .B(clk), .A(\g.we_clk [6890]));
Q_ASSIGN U9501 ( .B(clk), .A(\g.we_clk [6889]));
Q_ASSIGN U9502 ( .B(clk), .A(\g.we_clk [6888]));
Q_ASSIGN U9503 ( .B(clk), .A(\g.we_clk [6887]));
Q_ASSIGN U9504 ( .B(clk), .A(\g.we_clk [6886]));
Q_ASSIGN U9505 ( .B(clk), .A(\g.we_clk [6885]));
Q_ASSIGN U9506 ( .B(clk), .A(\g.we_clk [6884]));
Q_ASSIGN U9507 ( .B(clk), .A(\g.we_clk [6883]));
Q_ASSIGN U9508 ( .B(clk), .A(\g.we_clk [6882]));
Q_ASSIGN U9509 ( .B(clk), .A(\g.we_clk [6881]));
Q_ASSIGN U9510 ( .B(clk), .A(\g.we_clk [6880]));
Q_ASSIGN U9511 ( .B(clk), .A(\g.we_clk [6879]));
Q_ASSIGN U9512 ( .B(clk), .A(\g.we_clk [6878]));
Q_ASSIGN U9513 ( .B(clk), .A(\g.we_clk [6877]));
Q_ASSIGN U9514 ( .B(clk), .A(\g.we_clk [6876]));
Q_ASSIGN U9515 ( .B(clk), .A(\g.we_clk [6875]));
Q_ASSIGN U9516 ( .B(clk), .A(\g.we_clk [6874]));
Q_ASSIGN U9517 ( .B(clk), .A(\g.we_clk [6873]));
Q_ASSIGN U9518 ( .B(clk), .A(\g.we_clk [6872]));
Q_ASSIGN U9519 ( .B(clk), .A(\g.we_clk [6871]));
Q_ASSIGN U9520 ( .B(clk), .A(\g.we_clk [6870]));
Q_ASSIGN U9521 ( .B(clk), .A(\g.we_clk [6869]));
Q_ASSIGN U9522 ( .B(clk), .A(\g.we_clk [6868]));
Q_ASSIGN U9523 ( .B(clk), .A(\g.we_clk [6867]));
Q_ASSIGN U9524 ( .B(clk), .A(\g.we_clk [6866]));
Q_ASSIGN U9525 ( .B(clk), .A(\g.we_clk [6865]));
Q_ASSIGN U9526 ( .B(clk), .A(\g.we_clk [6864]));
Q_ASSIGN U9527 ( .B(clk), .A(\g.we_clk [6863]));
Q_ASSIGN U9528 ( .B(clk), .A(\g.we_clk [6862]));
Q_ASSIGN U9529 ( .B(clk), .A(\g.we_clk [6861]));
Q_ASSIGN U9530 ( .B(clk), .A(\g.we_clk [6860]));
Q_ASSIGN U9531 ( .B(clk), .A(\g.we_clk [6859]));
Q_ASSIGN U9532 ( .B(clk), .A(\g.we_clk [6858]));
Q_ASSIGN U9533 ( .B(clk), .A(\g.we_clk [6857]));
Q_ASSIGN U9534 ( .B(clk), .A(\g.we_clk [6856]));
Q_ASSIGN U9535 ( .B(clk), .A(\g.we_clk [6855]));
Q_ASSIGN U9536 ( .B(clk), .A(\g.we_clk [6854]));
Q_ASSIGN U9537 ( .B(clk), .A(\g.we_clk [6853]));
Q_ASSIGN U9538 ( .B(clk), .A(\g.we_clk [6852]));
Q_ASSIGN U9539 ( .B(clk), .A(\g.we_clk [6851]));
Q_ASSIGN U9540 ( .B(clk), .A(\g.we_clk [6850]));
Q_ASSIGN U9541 ( .B(clk), .A(\g.we_clk [6849]));
Q_ASSIGN U9542 ( .B(clk), .A(\g.we_clk [6848]));
Q_ASSIGN U9543 ( .B(clk), .A(\g.we_clk [6847]));
Q_ASSIGN U9544 ( .B(clk), .A(\g.we_clk [6846]));
Q_ASSIGN U9545 ( .B(clk), .A(\g.we_clk [6845]));
Q_ASSIGN U9546 ( .B(clk), .A(\g.we_clk [6844]));
Q_ASSIGN U9547 ( .B(clk), .A(\g.we_clk [6843]));
Q_ASSIGN U9548 ( .B(clk), .A(\g.we_clk [6842]));
Q_ASSIGN U9549 ( .B(clk), .A(\g.we_clk [6841]));
Q_ASSIGN U9550 ( .B(clk), .A(\g.we_clk [6840]));
Q_ASSIGN U9551 ( .B(clk), .A(\g.we_clk [6839]));
Q_ASSIGN U9552 ( .B(clk), .A(\g.we_clk [6838]));
Q_ASSIGN U9553 ( .B(clk), .A(\g.we_clk [6837]));
Q_ASSIGN U9554 ( .B(clk), .A(\g.we_clk [6836]));
Q_ASSIGN U9555 ( .B(clk), .A(\g.we_clk [6835]));
Q_ASSIGN U9556 ( .B(clk), .A(\g.we_clk [6834]));
Q_ASSIGN U9557 ( .B(clk), .A(\g.we_clk [6833]));
Q_ASSIGN U9558 ( .B(clk), .A(\g.we_clk [6832]));
Q_ASSIGN U9559 ( .B(clk), .A(\g.we_clk [6831]));
Q_ASSIGN U9560 ( .B(clk), .A(\g.we_clk [6830]));
Q_ASSIGN U9561 ( .B(clk), .A(\g.we_clk [6829]));
Q_ASSIGN U9562 ( .B(clk), .A(\g.we_clk [6828]));
Q_ASSIGN U9563 ( .B(clk), .A(\g.we_clk [6827]));
Q_ASSIGN U9564 ( .B(clk), .A(\g.we_clk [6826]));
Q_ASSIGN U9565 ( .B(clk), .A(\g.we_clk [6825]));
Q_ASSIGN U9566 ( .B(clk), .A(\g.we_clk [6824]));
Q_ASSIGN U9567 ( .B(clk), .A(\g.we_clk [6823]));
Q_ASSIGN U9568 ( .B(clk), .A(\g.we_clk [6822]));
Q_ASSIGN U9569 ( .B(clk), .A(\g.we_clk [6821]));
Q_ASSIGN U9570 ( .B(clk), .A(\g.we_clk [6820]));
Q_ASSIGN U9571 ( .B(clk), .A(\g.we_clk [6819]));
Q_ASSIGN U9572 ( .B(clk), .A(\g.we_clk [6818]));
Q_ASSIGN U9573 ( .B(clk), .A(\g.we_clk [6817]));
Q_ASSIGN U9574 ( .B(clk), .A(\g.we_clk [6816]));
Q_ASSIGN U9575 ( .B(clk), .A(\g.we_clk [6815]));
Q_ASSIGN U9576 ( .B(clk), .A(\g.we_clk [6814]));
Q_ASSIGN U9577 ( .B(clk), .A(\g.we_clk [6813]));
Q_ASSIGN U9578 ( .B(clk), .A(\g.we_clk [6812]));
Q_ASSIGN U9579 ( .B(clk), .A(\g.we_clk [6811]));
Q_ASSIGN U9580 ( .B(clk), .A(\g.we_clk [6810]));
Q_ASSIGN U9581 ( .B(clk), .A(\g.we_clk [6809]));
Q_ASSIGN U9582 ( .B(clk), .A(\g.we_clk [6808]));
Q_ASSIGN U9583 ( .B(clk), .A(\g.we_clk [6807]));
Q_ASSIGN U9584 ( .B(clk), .A(\g.we_clk [6806]));
Q_ASSIGN U9585 ( .B(clk), .A(\g.we_clk [6805]));
Q_ASSIGN U9586 ( .B(clk), .A(\g.we_clk [6804]));
Q_ASSIGN U9587 ( .B(clk), .A(\g.we_clk [6803]));
Q_ASSIGN U9588 ( .B(clk), .A(\g.we_clk [6802]));
Q_ASSIGN U9589 ( .B(clk), .A(\g.we_clk [6801]));
Q_ASSIGN U9590 ( .B(clk), .A(\g.we_clk [6800]));
Q_ASSIGN U9591 ( .B(clk), .A(\g.we_clk [6799]));
Q_ASSIGN U9592 ( .B(clk), .A(\g.we_clk [6798]));
Q_ASSIGN U9593 ( .B(clk), .A(\g.we_clk [6797]));
Q_ASSIGN U9594 ( .B(clk), .A(\g.we_clk [6796]));
Q_ASSIGN U9595 ( .B(clk), .A(\g.we_clk [6795]));
Q_ASSIGN U9596 ( .B(clk), .A(\g.we_clk [6794]));
Q_ASSIGN U9597 ( .B(clk), .A(\g.we_clk [6793]));
Q_ASSIGN U9598 ( .B(clk), .A(\g.we_clk [6792]));
Q_ASSIGN U9599 ( .B(clk), .A(\g.we_clk [6791]));
Q_ASSIGN U9600 ( .B(clk), .A(\g.we_clk [6790]));
Q_ASSIGN U9601 ( .B(clk), .A(\g.we_clk [6789]));
Q_ASSIGN U9602 ( .B(clk), .A(\g.we_clk [6788]));
Q_ASSIGN U9603 ( .B(clk), .A(\g.we_clk [6787]));
Q_ASSIGN U9604 ( .B(clk), .A(\g.we_clk [6786]));
Q_ASSIGN U9605 ( .B(clk), .A(\g.we_clk [6785]));
Q_ASSIGN U9606 ( .B(clk), .A(\g.we_clk [6784]));
Q_ASSIGN U9607 ( .B(clk), .A(\g.we_clk [6783]));
Q_ASSIGN U9608 ( .B(clk), .A(\g.we_clk [6782]));
Q_ASSIGN U9609 ( .B(clk), .A(\g.we_clk [6781]));
Q_ASSIGN U9610 ( .B(clk), .A(\g.we_clk [6780]));
Q_ASSIGN U9611 ( .B(clk), .A(\g.we_clk [6779]));
Q_ASSIGN U9612 ( .B(clk), .A(\g.we_clk [6778]));
Q_ASSIGN U9613 ( .B(clk), .A(\g.we_clk [6777]));
Q_ASSIGN U9614 ( .B(clk), .A(\g.we_clk [6776]));
Q_ASSIGN U9615 ( .B(clk), .A(\g.we_clk [6775]));
Q_ASSIGN U9616 ( .B(clk), .A(\g.we_clk [6774]));
Q_ASSIGN U9617 ( .B(clk), .A(\g.we_clk [6773]));
Q_ASSIGN U9618 ( .B(clk), .A(\g.we_clk [6772]));
Q_ASSIGN U9619 ( .B(clk), .A(\g.we_clk [6771]));
Q_ASSIGN U9620 ( .B(clk), .A(\g.we_clk [6770]));
Q_ASSIGN U9621 ( .B(clk), .A(\g.we_clk [6769]));
Q_ASSIGN U9622 ( .B(clk), .A(\g.we_clk [6768]));
Q_ASSIGN U9623 ( .B(clk), .A(\g.we_clk [6767]));
Q_ASSIGN U9624 ( .B(clk), .A(\g.we_clk [6766]));
Q_ASSIGN U9625 ( .B(clk), .A(\g.we_clk [6765]));
Q_ASSIGN U9626 ( .B(clk), .A(\g.we_clk [6764]));
Q_ASSIGN U9627 ( .B(clk), .A(\g.we_clk [6763]));
Q_ASSIGN U9628 ( .B(clk), .A(\g.we_clk [6762]));
Q_ASSIGN U9629 ( .B(clk), .A(\g.we_clk [6761]));
Q_ASSIGN U9630 ( .B(clk), .A(\g.we_clk [6760]));
Q_ASSIGN U9631 ( .B(clk), .A(\g.we_clk [6759]));
Q_ASSIGN U9632 ( .B(clk), .A(\g.we_clk [6758]));
Q_ASSIGN U9633 ( .B(clk), .A(\g.we_clk [6757]));
Q_ASSIGN U9634 ( .B(clk), .A(\g.we_clk [6756]));
Q_ASSIGN U9635 ( .B(clk), .A(\g.we_clk [6755]));
Q_ASSIGN U9636 ( .B(clk), .A(\g.we_clk [6754]));
Q_ASSIGN U9637 ( .B(clk), .A(\g.we_clk [6753]));
Q_ASSIGN U9638 ( .B(clk), .A(\g.we_clk [6752]));
Q_ASSIGN U9639 ( .B(clk), .A(\g.we_clk [6751]));
Q_ASSIGN U9640 ( .B(clk), .A(\g.we_clk [6750]));
Q_ASSIGN U9641 ( .B(clk), .A(\g.we_clk [6749]));
Q_ASSIGN U9642 ( .B(clk), .A(\g.we_clk [6748]));
Q_ASSIGN U9643 ( .B(clk), .A(\g.we_clk [6747]));
Q_ASSIGN U9644 ( .B(clk), .A(\g.we_clk [6746]));
Q_ASSIGN U9645 ( .B(clk), .A(\g.we_clk [6745]));
Q_ASSIGN U9646 ( .B(clk), .A(\g.we_clk [6744]));
Q_ASSIGN U9647 ( .B(clk), .A(\g.we_clk [6743]));
Q_ASSIGN U9648 ( .B(clk), .A(\g.we_clk [6742]));
Q_ASSIGN U9649 ( .B(clk), .A(\g.we_clk [6741]));
Q_ASSIGN U9650 ( .B(clk), .A(\g.we_clk [6740]));
Q_ASSIGN U9651 ( .B(clk), .A(\g.we_clk [6739]));
Q_ASSIGN U9652 ( .B(clk), .A(\g.we_clk [6738]));
Q_ASSIGN U9653 ( .B(clk), .A(\g.we_clk [6737]));
Q_ASSIGN U9654 ( .B(clk), .A(\g.we_clk [6736]));
Q_ASSIGN U9655 ( .B(clk), .A(\g.we_clk [6735]));
Q_ASSIGN U9656 ( .B(clk), .A(\g.we_clk [6734]));
Q_ASSIGN U9657 ( .B(clk), .A(\g.we_clk [6733]));
Q_ASSIGN U9658 ( .B(clk), .A(\g.we_clk [6732]));
Q_ASSIGN U9659 ( .B(clk), .A(\g.we_clk [6731]));
Q_ASSIGN U9660 ( .B(clk), .A(\g.we_clk [6730]));
Q_ASSIGN U9661 ( .B(clk), .A(\g.we_clk [6729]));
Q_ASSIGN U9662 ( .B(clk), .A(\g.we_clk [6728]));
Q_ASSIGN U9663 ( .B(clk), .A(\g.we_clk [6727]));
Q_ASSIGN U9664 ( .B(clk), .A(\g.we_clk [6726]));
Q_ASSIGN U9665 ( .B(clk), .A(\g.we_clk [6725]));
Q_ASSIGN U9666 ( .B(clk), .A(\g.we_clk [6724]));
Q_ASSIGN U9667 ( .B(clk), .A(\g.we_clk [6723]));
Q_ASSIGN U9668 ( .B(clk), .A(\g.we_clk [6722]));
Q_ASSIGN U9669 ( .B(clk), .A(\g.we_clk [6721]));
Q_ASSIGN U9670 ( .B(clk), .A(\g.we_clk [6720]));
Q_ASSIGN U9671 ( .B(clk), .A(\g.we_clk [6719]));
Q_ASSIGN U9672 ( .B(clk), .A(\g.we_clk [6718]));
Q_ASSIGN U9673 ( .B(clk), .A(\g.we_clk [6717]));
Q_ASSIGN U9674 ( .B(clk), .A(\g.we_clk [6716]));
Q_ASSIGN U9675 ( .B(clk), .A(\g.we_clk [6715]));
Q_ASSIGN U9676 ( .B(clk), .A(\g.we_clk [6714]));
Q_ASSIGN U9677 ( .B(clk), .A(\g.we_clk [6713]));
Q_ASSIGN U9678 ( .B(clk), .A(\g.we_clk [6712]));
Q_ASSIGN U9679 ( .B(clk), .A(\g.we_clk [6711]));
Q_ASSIGN U9680 ( .B(clk), .A(\g.we_clk [6710]));
Q_ASSIGN U9681 ( .B(clk), .A(\g.we_clk [6709]));
Q_ASSIGN U9682 ( .B(clk), .A(\g.we_clk [6708]));
Q_ASSIGN U9683 ( .B(clk), .A(\g.we_clk [6707]));
Q_ASSIGN U9684 ( .B(clk), .A(\g.we_clk [6706]));
Q_ASSIGN U9685 ( .B(clk), .A(\g.we_clk [6705]));
Q_ASSIGN U9686 ( .B(clk), .A(\g.we_clk [6704]));
Q_ASSIGN U9687 ( .B(clk), .A(\g.we_clk [6703]));
Q_ASSIGN U9688 ( .B(clk), .A(\g.we_clk [6702]));
Q_ASSIGN U9689 ( .B(clk), .A(\g.we_clk [6701]));
Q_ASSIGN U9690 ( .B(clk), .A(\g.we_clk [6700]));
Q_ASSIGN U9691 ( .B(clk), .A(\g.we_clk [6699]));
Q_ASSIGN U9692 ( .B(clk), .A(\g.we_clk [6698]));
Q_ASSIGN U9693 ( .B(clk), .A(\g.we_clk [6697]));
Q_ASSIGN U9694 ( .B(clk), .A(\g.we_clk [6696]));
Q_ASSIGN U9695 ( .B(clk), .A(\g.we_clk [6695]));
Q_ASSIGN U9696 ( .B(clk), .A(\g.we_clk [6694]));
Q_ASSIGN U9697 ( .B(clk), .A(\g.we_clk [6693]));
Q_ASSIGN U9698 ( .B(clk), .A(\g.we_clk [6692]));
Q_ASSIGN U9699 ( .B(clk), .A(\g.we_clk [6691]));
Q_ASSIGN U9700 ( .B(clk), .A(\g.we_clk [6690]));
Q_ASSIGN U9701 ( .B(clk), .A(\g.we_clk [6689]));
Q_ASSIGN U9702 ( .B(clk), .A(\g.we_clk [6688]));
Q_ASSIGN U9703 ( .B(clk), .A(\g.we_clk [6687]));
Q_ASSIGN U9704 ( .B(clk), .A(\g.we_clk [6686]));
Q_ASSIGN U9705 ( .B(clk), .A(\g.we_clk [6685]));
Q_ASSIGN U9706 ( .B(clk), .A(\g.we_clk [6684]));
Q_ASSIGN U9707 ( .B(clk), .A(\g.we_clk [6683]));
Q_ASSIGN U9708 ( .B(clk), .A(\g.we_clk [6682]));
Q_ASSIGN U9709 ( .B(clk), .A(\g.we_clk [6681]));
Q_ASSIGN U9710 ( .B(clk), .A(\g.we_clk [6680]));
Q_ASSIGN U9711 ( .B(clk), .A(\g.we_clk [6679]));
Q_ASSIGN U9712 ( .B(clk), .A(\g.we_clk [6678]));
Q_ASSIGN U9713 ( .B(clk), .A(\g.we_clk [6677]));
Q_ASSIGN U9714 ( .B(clk), .A(\g.we_clk [6676]));
Q_ASSIGN U9715 ( .B(clk), .A(\g.we_clk [6675]));
Q_ASSIGN U9716 ( .B(clk), .A(\g.we_clk [6674]));
Q_ASSIGN U9717 ( .B(clk), .A(\g.we_clk [6673]));
Q_ASSIGN U9718 ( .B(clk), .A(\g.we_clk [6672]));
Q_ASSIGN U9719 ( .B(clk), .A(\g.we_clk [6671]));
Q_ASSIGN U9720 ( .B(clk), .A(\g.we_clk [6670]));
Q_ASSIGN U9721 ( .B(clk), .A(\g.we_clk [6669]));
Q_ASSIGN U9722 ( .B(clk), .A(\g.we_clk [6668]));
Q_ASSIGN U9723 ( .B(clk), .A(\g.we_clk [6667]));
Q_ASSIGN U9724 ( .B(clk), .A(\g.we_clk [6666]));
Q_ASSIGN U9725 ( .B(clk), .A(\g.we_clk [6665]));
Q_ASSIGN U9726 ( .B(clk), .A(\g.we_clk [6664]));
Q_ASSIGN U9727 ( .B(clk), .A(\g.we_clk [6663]));
Q_ASSIGN U9728 ( .B(clk), .A(\g.we_clk [6662]));
Q_ASSIGN U9729 ( .B(clk), .A(\g.we_clk [6661]));
Q_ASSIGN U9730 ( .B(clk), .A(\g.we_clk [6660]));
Q_ASSIGN U9731 ( .B(clk), .A(\g.we_clk [6659]));
Q_ASSIGN U9732 ( .B(clk), .A(\g.we_clk [6658]));
Q_ASSIGN U9733 ( .B(clk), .A(\g.we_clk [6657]));
Q_ASSIGN U9734 ( .B(clk), .A(\g.we_clk [6656]));
Q_ASSIGN U9735 ( .B(clk), .A(\g.we_clk [6655]));
Q_ASSIGN U9736 ( .B(clk), .A(\g.we_clk [6654]));
Q_ASSIGN U9737 ( .B(clk), .A(\g.we_clk [6653]));
Q_ASSIGN U9738 ( .B(clk), .A(\g.we_clk [6652]));
Q_ASSIGN U9739 ( .B(clk), .A(\g.we_clk [6651]));
Q_ASSIGN U9740 ( .B(clk), .A(\g.we_clk [6650]));
Q_ASSIGN U9741 ( .B(clk), .A(\g.we_clk [6649]));
Q_ASSIGN U9742 ( .B(clk), .A(\g.we_clk [6648]));
Q_ASSIGN U9743 ( .B(clk), .A(\g.we_clk [6647]));
Q_ASSIGN U9744 ( .B(clk), .A(\g.we_clk [6646]));
Q_ASSIGN U9745 ( .B(clk), .A(\g.we_clk [6645]));
Q_ASSIGN U9746 ( .B(clk), .A(\g.we_clk [6644]));
Q_ASSIGN U9747 ( .B(clk), .A(\g.we_clk [6643]));
Q_ASSIGN U9748 ( .B(clk), .A(\g.we_clk [6642]));
Q_ASSIGN U9749 ( .B(clk), .A(\g.we_clk [6641]));
Q_ASSIGN U9750 ( .B(clk), .A(\g.we_clk [6640]));
Q_ASSIGN U9751 ( .B(clk), .A(\g.we_clk [6639]));
Q_ASSIGN U9752 ( .B(clk), .A(\g.we_clk [6638]));
Q_ASSIGN U9753 ( .B(clk), .A(\g.we_clk [6637]));
Q_ASSIGN U9754 ( .B(clk), .A(\g.we_clk [6636]));
Q_ASSIGN U9755 ( .B(clk), .A(\g.we_clk [6635]));
Q_ASSIGN U9756 ( .B(clk), .A(\g.we_clk [6634]));
Q_ASSIGN U9757 ( .B(clk), .A(\g.we_clk [6633]));
Q_ASSIGN U9758 ( .B(clk), .A(\g.we_clk [6632]));
Q_ASSIGN U9759 ( .B(clk), .A(\g.we_clk [6631]));
Q_ASSIGN U9760 ( .B(clk), .A(\g.we_clk [6630]));
Q_ASSIGN U9761 ( .B(clk), .A(\g.we_clk [6629]));
Q_ASSIGN U9762 ( .B(clk), .A(\g.we_clk [6628]));
Q_ASSIGN U9763 ( .B(clk), .A(\g.we_clk [6627]));
Q_ASSIGN U9764 ( .B(clk), .A(\g.we_clk [6626]));
Q_ASSIGN U9765 ( .B(clk), .A(\g.we_clk [6625]));
Q_ASSIGN U9766 ( .B(clk), .A(\g.we_clk [6624]));
Q_ASSIGN U9767 ( .B(clk), .A(\g.we_clk [6623]));
Q_ASSIGN U9768 ( .B(clk), .A(\g.we_clk [6622]));
Q_ASSIGN U9769 ( .B(clk), .A(\g.we_clk [6621]));
Q_ASSIGN U9770 ( .B(clk), .A(\g.we_clk [6620]));
Q_ASSIGN U9771 ( .B(clk), .A(\g.we_clk [6619]));
Q_ASSIGN U9772 ( .B(clk), .A(\g.we_clk [6618]));
Q_ASSIGN U9773 ( .B(clk), .A(\g.we_clk [6617]));
Q_ASSIGN U9774 ( .B(clk), .A(\g.we_clk [6616]));
Q_ASSIGN U9775 ( .B(clk), .A(\g.we_clk [6615]));
Q_ASSIGN U9776 ( .B(clk), .A(\g.we_clk [6614]));
Q_ASSIGN U9777 ( .B(clk), .A(\g.we_clk [6613]));
Q_ASSIGN U9778 ( .B(clk), .A(\g.we_clk [6612]));
Q_ASSIGN U9779 ( .B(clk), .A(\g.we_clk [6611]));
Q_ASSIGN U9780 ( .B(clk), .A(\g.we_clk [6610]));
Q_ASSIGN U9781 ( .B(clk), .A(\g.we_clk [6609]));
Q_ASSIGN U9782 ( .B(clk), .A(\g.we_clk [6608]));
Q_ASSIGN U9783 ( .B(clk), .A(\g.we_clk [6607]));
Q_ASSIGN U9784 ( .B(clk), .A(\g.we_clk [6606]));
Q_ASSIGN U9785 ( .B(clk), .A(\g.we_clk [6605]));
Q_ASSIGN U9786 ( .B(clk), .A(\g.we_clk [6604]));
Q_ASSIGN U9787 ( .B(clk), .A(\g.we_clk [6603]));
Q_ASSIGN U9788 ( .B(clk), .A(\g.we_clk [6602]));
Q_ASSIGN U9789 ( .B(clk), .A(\g.we_clk [6601]));
Q_ASSIGN U9790 ( .B(clk), .A(\g.we_clk [6600]));
Q_ASSIGN U9791 ( .B(clk), .A(\g.we_clk [6599]));
Q_ASSIGN U9792 ( .B(clk), .A(\g.we_clk [6598]));
Q_ASSIGN U9793 ( .B(clk), .A(\g.we_clk [6597]));
Q_ASSIGN U9794 ( .B(clk), .A(\g.we_clk [6596]));
Q_ASSIGN U9795 ( .B(clk), .A(\g.we_clk [6595]));
Q_ASSIGN U9796 ( .B(clk), .A(\g.we_clk [6594]));
Q_ASSIGN U9797 ( .B(clk), .A(\g.we_clk [6593]));
Q_ASSIGN U9798 ( .B(clk), .A(\g.we_clk [6592]));
Q_ASSIGN U9799 ( .B(clk), .A(\g.we_clk [6591]));
Q_ASSIGN U9800 ( .B(clk), .A(\g.we_clk [6590]));
Q_ASSIGN U9801 ( .B(clk), .A(\g.we_clk [6589]));
Q_ASSIGN U9802 ( .B(clk), .A(\g.we_clk [6588]));
Q_ASSIGN U9803 ( .B(clk), .A(\g.we_clk [6587]));
Q_ASSIGN U9804 ( .B(clk), .A(\g.we_clk [6586]));
Q_ASSIGN U9805 ( .B(clk), .A(\g.we_clk [6585]));
Q_ASSIGN U9806 ( .B(clk), .A(\g.we_clk [6584]));
Q_ASSIGN U9807 ( .B(clk), .A(\g.we_clk [6583]));
Q_ASSIGN U9808 ( .B(clk), .A(\g.we_clk [6582]));
Q_ASSIGN U9809 ( .B(clk), .A(\g.we_clk [6581]));
Q_ASSIGN U9810 ( .B(clk), .A(\g.we_clk [6580]));
Q_ASSIGN U9811 ( .B(clk), .A(\g.we_clk [6579]));
Q_ASSIGN U9812 ( .B(clk), .A(\g.we_clk [6578]));
Q_ASSIGN U9813 ( .B(clk), .A(\g.we_clk [6577]));
Q_ASSIGN U9814 ( .B(clk), .A(\g.we_clk [6576]));
Q_ASSIGN U9815 ( .B(clk), .A(\g.we_clk [6575]));
Q_ASSIGN U9816 ( .B(clk), .A(\g.we_clk [6574]));
Q_ASSIGN U9817 ( .B(clk), .A(\g.we_clk [6573]));
Q_ASSIGN U9818 ( .B(clk), .A(\g.we_clk [6572]));
Q_ASSIGN U9819 ( .B(clk), .A(\g.we_clk [6571]));
Q_ASSIGN U9820 ( .B(clk), .A(\g.we_clk [6570]));
Q_ASSIGN U9821 ( .B(clk), .A(\g.we_clk [6569]));
Q_ASSIGN U9822 ( .B(clk), .A(\g.we_clk [6568]));
Q_ASSIGN U9823 ( .B(clk), .A(\g.we_clk [6567]));
Q_ASSIGN U9824 ( .B(clk), .A(\g.we_clk [6566]));
Q_ASSIGN U9825 ( .B(clk), .A(\g.we_clk [6565]));
Q_ASSIGN U9826 ( .B(clk), .A(\g.we_clk [6564]));
Q_ASSIGN U9827 ( .B(clk), .A(\g.we_clk [6563]));
Q_ASSIGN U9828 ( .B(clk), .A(\g.we_clk [6562]));
Q_ASSIGN U9829 ( .B(clk), .A(\g.we_clk [6561]));
Q_ASSIGN U9830 ( .B(clk), .A(\g.we_clk [6560]));
Q_ASSIGN U9831 ( .B(clk), .A(\g.we_clk [6559]));
Q_ASSIGN U9832 ( .B(clk), .A(\g.we_clk [6558]));
Q_ASSIGN U9833 ( .B(clk), .A(\g.we_clk [6557]));
Q_ASSIGN U9834 ( .B(clk), .A(\g.we_clk [6556]));
Q_ASSIGN U9835 ( .B(clk), .A(\g.we_clk [6555]));
Q_ASSIGN U9836 ( .B(clk), .A(\g.we_clk [6554]));
Q_ASSIGN U9837 ( .B(clk), .A(\g.we_clk [6553]));
Q_ASSIGN U9838 ( .B(clk), .A(\g.we_clk [6552]));
Q_ASSIGN U9839 ( .B(clk), .A(\g.we_clk [6551]));
Q_ASSIGN U9840 ( .B(clk), .A(\g.we_clk [6550]));
Q_ASSIGN U9841 ( .B(clk), .A(\g.we_clk [6549]));
Q_ASSIGN U9842 ( .B(clk), .A(\g.we_clk [6548]));
Q_ASSIGN U9843 ( .B(clk), .A(\g.we_clk [6547]));
Q_ASSIGN U9844 ( .B(clk), .A(\g.we_clk [6546]));
Q_ASSIGN U9845 ( .B(clk), .A(\g.we_clk [6545]));
Q_ASSIGN U9846 ( .B(clk), .A(\g.we_clk [6544]));
Q_ASSIGN U9847 ( .B(clk), .A(\g.we_clk [6543]));
Q_ASSIGN U9848 ( .B(clk), .A(\g.we_clk [6542]));
Q_ASSIGN U9849 ( .B(clk), .A(\g.we_clk [6541]));
Q_ASSIGN U9850 ( .B(clk), .A(\g.we_clk [6540]));
Q_ASSIGN U9851 ( .B(clk), .A(\g.we_clk [6539]));
Q_ASSIGN U9852 ( .B(clk), .A(\g.we_clk [6538]));
Q_ASSIGN U9853 ( .B(clk), .A(\g.we_clk [6537]));
Q_ASSIGN U9854 ( .B(clk), .A(\g.we_clk [6536]));
Q_ASSIGN U9855 ( .B(clk), .A(\g.we_clk [6535]));
Q_ASSIGN U9856 ( .B(clk), .A(\g.we_clk [6534]));
Q_ASSIGN U9857 ( .B(clk), .A(\g.we_clk [6533]));
Q_ASSIGN U9858 ( .B(clk), .A(\g.we_clk [6532]));
Q_ASSIGN U9859 ( .B(clk), .A(\g.we_clk [6531]));
Q_ASSIGN U9860 ( .B(clk), .A(\g.we_clk [6530]));
Q_ASSIGN U9861 ( .B(clk), .A(\g.we_clk [6529]));
Q_ASSIGN U9862 ( .B(clk), .A(\g.we_clk [6528]));
Q_ASSIGN U9863 ( .B(clk), .A(\g.we_clk [6527]));
Q_ASSIGN U9864 ( .B(clk), .A(\g.we_clk [6526]));
Q_ASSIGN U9865 ( .B(clk), .A(\g.we_clk [6525]));
Q_ASSIGN U9866 ( .B(clk), .A(\g.we_clk [6524]));
Q_ASSIGN U9867 ( .B(clk), .A(\g.we_clk [6523]));
Q_ASSIGN U9868 ( .B(clk), .A(\g.we_clk [6522]));
Q_ASSIGN U9869 ( .B(clk), .A(\g.we_clk [6521]));
Q_ASSIGN U9870 ( .B(clk), .A(\g.we_clk [6520]));
Q_ASSIGN U9871 ( .B(clk), .A(\g.we_clk [6519]));
Q_ASSIGN U9872 ( .B(clk), .A(\g.we_clk [6518]));
Q_ASSIGN U9873 ( .B(clk), .A(\g.we_clk [6517]));
Q_ASSIGN U9874 ( .B(clk), .A(\g.we_clk [6516]));
Q_ASSIGN U9875 ( .B(clk), .A(\g.we_clk [6515]));
Q_ASSIGN U9876 ( .B(clk), .A(\g.we_clk [6514]));
Q_ASSIGN U9877 ( .B(clk), .A(\g.we_clk [6513]));
Q_ASSIGN U9878 ( .B(clk), .A(\g.we_clk [6512]));
Q_ASSIGN U9879 ( .B(clk), .A(\g.we_clk [6511]));
Q_ASSIGN U9880 ( .B(clk), .A(\g.we_clk [6510]));
Q_ASSIGN U9881 ( .B(clk), .A(\g.we_clk [6509]));
Q_ASSIGN U9882 ( .B(clk), .A(\g.we_clk [6508]));
Q_ASSIGN U9883 ( .B(clk), .A(\g.we_clk [6507]));
Q_ASSIGN U9884 ( .B(clk), .A(\g.we_clk [6506]));
Q_ASSIGN U9885 ( .B(clk), .A(\g.we_clk [6505]));
Q_ASSIGN U9886 ( .B(clk), .A(\g.we_clk [6504]));
Q_ASSIGN U9887 ( .B(clk), .A(\g.we_clk [6503]));
Q_ASSIGN U9888 ( .B(clk), .A(\g.we_clk [6502]));
Q_ASSIGN U9889 ( .B(clk), .A(\g.we_clk [6501]));
Q_ASSIGN U9890 ( .B(clk), .A(\g.we_clk [6500]));
Q_ASSIGN U9891 ( .B(clk), .A(\g.we_clk [6499]));
Q_ASSIGN U9892 ( .B(clk), .A(\g.we_clk [6498]));
Q_ASSIGN U9893 ( .B(clk), .A(\g.we_clk [6497]));
Q_ASSIGN U9894 ( .B(clk), .A(\g.we_clk [6496]));
Q_ASSIGN U9895 ( .B(clk), .A(\g.we_clk [6495]));
Q_ASSIGN U9896 ( .B(clk), .A(\g.we_clk [6494]));
Q_ASSIGN U9897 ( .B(clk), .A(\g.we_clk [6493]));
Q_ASSIGN U9898 ( .B(clk), .A(\g.we_clk [6492]));
Q_ASSIGN U9899 ( .B(clk), .A(\g.we_clk [6491]));
Q_ASSIGN U9900 ( .B(clk), .A(\g.we_clk [6490]));
Q_ASSIGN U9901 ( .B(clk), .A(\g.we_clk [6489]));
Q_ASSIGN U9902 ( .B(clk), .A(\g.we_clk [6488]));
Q_ASSIGN U9903 ( .B(clk), .A(\g.we_clk [6487]));
Q_ASSIGN U9904 ( .B(clk), .A(\g.we_clk [6486]));
Q_ASSIGN U9905 ( .B(clk), .A(\g.we_clk [6485]));
Q_ASSIGN U9906 ( .B(clk), .A(\g.we_clk [6484]));
Q_ASSIGN U9907 ( .B(clk), .A(\g.we_clk [6483]));
Q_ASSIGN U9908 ( .B(clk), .A(\g.we_clk [6482]));
Q_ASSIGN U9909 ( .B(clk), .A(\g.we_clk [6481]));
Q_ASSIGN U9910 ( .B(clk), .A(\g.we_clk [6480]));
Q_ASSIGN U9911 ( .B(clk), .A(\g.we_clk [6479]));
Q_ASSIGN U9912 ( .B(clk), .A(\g.we_clk [6478]));
Q_ASSIGN U9913 ( .B(clk), .A(\g.we_clk [6477]));
Q_ASSIGN U9914 ( .B(clk), .A(\g.we_clk [6476]));
Q_ASSIGN U9915 ( .B(clk), .A(\g.we_clk [6475]));
Q_ASSIGN U9916 ( .B(clk), .A(\g.we_clk [6474]));
Q_ASSIGN U9917 ( .B(clk), .A(\g.we_clk [6473]));
Q_ASSIGN U9918 ( .B(clk), .A(\g.we_clk [6472]));
Q_ASSIGN U9919 ( .B(clk), .A(\g.we_clk [6471]));
Q_ASSIGN U9920 ( .B(clk), .A(\g.we_clk [6470]));
Q_ASSIGN U9921 ( .B(clk), .A(\g.we_clk [6469]));
Q_ASSIGN U9922 ( .B(clk), .A(\g.we_clk [6468]));
Q_ASSIGN U9923 ( .B(clk), .A(\g.we_clk [6467]));
Q_ASSIGN U9924 ( .B(clk), .A(\g.we_clk [6466]));
Q_ASSIGN U9925 ( .B(clk), .A(\g.we_clk [6465]));
Q_ASSIGN U9926 ( .B(clk), .A(\g.we_clk [6464]));
Q_ASSIGN U9927 ( .B(clk), .A(\g.we_clk [6463]));
Q_ASSIGN U9928 ( .B(clk), .A(\g.we_clk [6462]));
Q_ASSIGN U9929 ( .B(clk), .A(\g.we_clk [6461]));
Q_ASSIGN U9930 ( .B(clk), .A(\g.we_clk [6460]));
Q_ASSIGN U9931 ( .B(clk), .A(\g.we_clk [6459]));
Q_ASSIGN U9932 ( .B(clk), .A(\g.we_clk [6458]));
Q_ASSIGN U9933 ( .B(clk), .A(\g.we_clk [6457]));
Q_ASSIGN U9934 ( .B(clk), .A(\g.we_clk [6456]));
Q_ASSIGN U9935 ( .B(clk), .A(\g.we_clk [6455]));
Q_ASSIGN U9936 ( .B(clk), .A(\g.we_clk [6454]));
Q_ASSIGN U9937 ( .B(clk), .A(\g.we_clk [6453]));
Q_ASSIGN U9938 ( .B(clk), .A(\g.we_clk [6452]));
Q_ASSIGN U9939 ( .B(clk), .A(\g.we_clk [6451]));
Q_ASSIGN U9940 ( .B(clk), .A(\g.we_clk [6450]));
Q_ASSIGN U9941 ( .B(clk), .A(\g.we_clk [6449]));
Q_ASSIGN U9942 ( .B(clk), .A(\g.we_clk [6448]));
Q_ASSIGN U9943 ( .B(clk), .A(\g.we_clk [6447]));
Q_ASSIGN U9944 ( .B(clk), .A(\g.we_clk [6446]));
Q_ASSIGN U9945 ( .B(clk), .A(\g.we_clk [6445]));
Q_ASSIGN U9946 ( .B(clk), .A(\g.we_clk [6444]));
Q_ASSIGN U9947 ( .B(clk), .A(\g.we_clk [6443]));
Q_ASSIGN U9948 ( .B(clk), .A(\g.we_clk [6442]));
Q_ASSIGN U9949 ( .B(clk), .A(\g.we_clk [6441]));
Q_ASSIGN U9950 ( .B(clk), .A(\g.we_clk [6440]));
Q_ASSIGN U9951 ( .B(clk), .A(\g.we_clk [6439]));
Q_ASSIGN U9952 ( .B(clk), .A(\g.we_clk [6438]));
Q_ASSIGN U9953 ( .B(clk), .A(\g.we_clk [6437]));
Q_ASSIGN U9954 ( .B(clk), .A(\g.we_clk [6436]));
Q_ASSIGN U9955 ( .B(clk), .A(\g.we_clk [6435]));
Q_ASSIGN U9956 ( .B(clk), .A(\g.we_clk [6434]));
Q_ASSIGN U9957 ( .B(clk), .A(\g.we_clk [6433]));
Q_ASSIGN U9958 ( .B(clk), .A(\g.we_clk [6432]));
Q_ASSIGN U9959 ( .B(clk), .A(\g.we_clk [6431]));
Q_ASSIGN U9960 ( .B(clk), .A(\g.we_clk [6430]));
Q_ASSIGN U9961 ( .B(clk), .A(\g.we_clk [6429]));
Q_ASSIGN U9962 ( .B(clk), .A(\g.we_clk [6428]));
Q_ASSIGN U9963 ( .B(clk), .A(\g.we_clk [6427]));
Q_ASSIGN U9964 ( .B(clk), .A(\g.we_clk [6426]));
Q_ASSIGN U9965 ( .B(clk), .A(\g.we_clk [6425]));
Q_ASSIGN U9966 ( .B(clk), .A(\g.we_clk [6424]));
Q_ASSIGN U9967 ( .B(clk), .A(\g.we_clk [6423]));
Q_ASSIGN U9968 ( .B(clk), .A(\g.we_clk [6422]));
Q_ASSIGN U9969 ( .B(clk), .A(\g.we_clk [6421]));
Q_ASSIGN U9970 ( .B(clk), .A(\g.we_clk [6420]));
Q_ASSIGN U9971 ( .B(clk), .A(\g.we_clk [6419]));
Q_ASSIGN U9972 ( .B(clk), .A(\g.we_clk [6418]));
Q_ASSIGN U9973 ( .B(clk), .A(\g.we_clk [6417]));
Q_ASSIGN U9974 ( .B(clk), .A(\g.we_clk [6416]));
Q_ASSIGN U9975 ( .B(clk), .A(\g.we_clk [6415]));
Q_ASSIGN U9976 ( .B(clk), .A(\g.we_clk [6414]));
Q_ASSIGN U9977 ( .B(clk), .A(\g.we_clk [6413]));
Q_ASSIGN U9978 ( .B(clk), .A(\g.we_clk [6412]));
Q_ASSIGN U9979 ( .B(clk), .A(\g.we_clk [6411]));
Q_ASSIGN U9980 ( .B(clk), .A(\g.we_clk [6410]));
Q_ASSIGN U9981 ( .B(clk), .A(\g.we_clk [6409]));
Q_ASSIGN U9982 ( .B(clk), .A(\g.we_clk [6408]));
Q_ASSIGN U9983 ( .B(clk), .A(\g.we_clk [6407]));
Q_ASSIGN U9984 ( .B(clk), .A(\g.we_clk [6406]));
Q_ASSIGN U9985 ( .B(clk), .A(\g.we_clk [6405]));
Q_ASSIGN U9986 ( .B(clk), .A(\g.we_clk [6404]));
Q_ASSIGN U9987 ( .B(clk), .A(\g.we_clk [6403]));
Q_ASSIGN U9988 ( .B(clk), .A(\g.we_clk [6402]));
Q_ASSIGN U9989 ( .B(clk), .A(\g.we_clk [6401]));
Q_ASSIGN U9990 ( .B(clk), .A(\g.we_clk [6400]));
Q_ASSIGN U9991 ( .B(clk), .A(\g.we_clk [6399]));
Q_ASSIGN U9992 ( .B(clk), .A(\g.we_clk [6398]));
Q_ASSIGN U9993 ( .B(clk), .A(\g.we_clk [6397]));
Q_ASSIGN U9994 ( .B(clk), .A(\g.we_clk [6396]));
Q_ASSIGN U9995 ( .B(clk), .A(\g.we_clk [6395]));
Q_ASSIGN U9996 ( .B(clk), .A(\g.we_clk [6394]));
Q_ASSIGN U9997 ( .B(clk), .A(\g.we_clk [6393]));
Q_ASSIGN U9998 ( .B(clk), .A(\g.we_clk [6392]));
Q_ASSIGN U9999 ( .B(clk), .A(\g.we_clk [6391]));
Q_ASSIGN U10000 ( .B(clk), .A(\g.we_clk [6390]));
Q_ASSIGN U10001 ( .B(clk), .A(\g.we_clk [6389]));
Q_ASSIGN U10002 ( .B(clk), .A(\g.we_clk [6388]));
Q_ASSIGN U10003 ( .B(clk), .A(\g.we_clk [6387]));
Q_ASSIGN U10004 ( .B(clk), .A(\g.we_clk [6386]));
Q_ASSIGN U10005 ( .B(clk), .A(\g.we_clk [6385]));
Q_ASSIGN U10006 ( .B(clk), .A(\g.we_clk [6384]));
Q_ASSIGN U10007 ( .B(clk), .A(\g.we_clk [6383]));
Q_ASSIGN U10008 ( .B(clk), .A(\g.we_clk [6382]));
Q_ASSIGN U10009 ( .B(clk), .A(\g.we_clk [6381]));
Q_ASSIGN U10010 ( .B(clk), .A(\g.we_clk [6380]));
Q_ASSIGN U10011 ( .B(clk), .A(\g.we_clk [6379]));
Q_ASSIGN U10012 ( .B(clk), .A(\g.we_clk [6378]));
Q_ASSIGN U10013 ( .B(clk), .A(\g.we_clk [6377]));
Q_ASSIGN U10014 ( .B(clk), .A(\g.we_clk [6376]));
Q_ASSIGN U10015 ( .B(clk), .A(\g.we_clk [6375]));
Q_ASSIGN U10016 ( .B(clk), .A(\g.we_clk [6374]));
Q_ASSIGN U10017 ( .B(clk), .A(\g.we_clk [6373]));
Q_ASSIGN U10018 ( .B(clk), .A(\g.we_clk [6372]));
Q_ASSIGN U10019 ( .B(clk), .A(\g.we_clk [6371]));
Q_ASSIGN U10020 ( .B(clk), .A(\g.we_clk [6370]));
Q_ASSIGN U10021 ( .B(clk), .A(\g.we_clk [6369]));
Q_ASSIGN U10022 ( .B(clk), .A(\g.we_clk [6368]));
Q_ASSIGN U10023 ( .B(clk), .A(\g.we_clk [6367]));
Q_ASSIGN U10024 ( .B(clk), .A(\g.we_clk [6366]));
Q_ASSIGN U10025 ( .B(clk), .A(\g.we_clk [6365]));
Q_ASSIGN U10026 ( .B(clk), .A(\g.we_clk [6364]));
Q_ASSIGN U10027 ( .B(clk), .A(\g.we_clk [6363]));
Q_ASSIGN U10028 ( .B(clk), .A(\g.we_clk [6362]));
Q_ASSIGN U10029 ( .B(clk), .A(\g.we_clk [6361]));
Q_ASSIGN U10030 ( .B(clk), .A(\g.we_clk [6360]));
Q_ASSIGN U10031 ( .B(clk), .A(\g.we_clk [6359]));
Q_ASSIGN U10032 ( .B(clk), .A(\g.we_clk [6358]));
Q_ASSIGN U10033 ( .B(clk), .A(\g.we_clk [6357]));
Q_ASSIGN U10034 ( .B(clk), .A(\g.we_clk [6356]));
Q_ASSIGN U10035 ( .B(clk), .A(\g.we_clk [6355]));
Q_ASSIGN U10036 ( .B(clk), .A(\g.we_clk [6354]));
Q_ASSIGN U10037 ( .B(clk), .A(\g.we_clk [6353]));
Q_ASSIGN U10038 ( .B(clk), .A(\g.we_clk [6352]));
Q_ASSIGN U10039 ( .B(clk), .A(\g.we_clk [6351]));
Q_ASSIGN U10040 ( .B(clk), .A(\g.we_clk [6350]));
Q_ASSIGN U10041 ( .B(clk), .A(\g.we_clk [6349]));
Q_ASSIGN U10042 ( .B(clk), .A(\g.we_clk [6348]));
Q_ASSIGN U10043 ( .B(clk), .A(\g.we_clk [6347]));
Q_ASSIGN U10044 ( .B(clk), .A(\g.we_clk [6346]));
Q_ASSIGN U10045 ( .B(clk), .A(\g.we_clk [6345]));
Q_ASSIGN U10046 ( .B(clk), .A(\g.we_clk [6344]));
Q_ASSIGN U10047 ( .B(clk), .A(\g.we_clk [6343]));
Q_ASSIGN U10048 ( .B(clk), .A(\g.we_clk [6342]));
Q_ASSIGN U10049 ( .B(clk), .A(\g.we_clk [6341]));
Q_ASSIGN U10050 ( .B(clk), .A(\g.we_clk [6340]));
Q_ASSIGN U10051 ( .B(clk), .A(\g.we_clk [6339]));
Q_ASSIGN U10052 ( .B(clk), .A(\g.we_clk [6338]));
Q_ASSIGN U10053 ( .B(clk), .A(\g.we_clk [6337]));
Q_ASSIGN U10054 ( .B(clk), .A(\g.we_clk [6336]));
Q_ASSIGN U10055 ( .B(clk), .A(\g.we_clk [6335]));
Q_ASSIGN U10056 ( .B(clk), .A(\g.we_clk [6334]));
Q_ASSIGN U10057 ( .B(clk), .A(\g.we_clk [6333]));
Q_ASSIGN U10058 ( .B(clk), .A(\g.we_clk [6332]));
Q_ASSIGN U10059 ( .B(clk), .A(\g.we_clk [6331]));
Q_ASSIGN U10060 ( .B(clk), .A(\g.we_clk [6330]));
Q_ASSIGN U10061 ( .B(clk), .A(\g.we_clk [6329]));
Q_ASSIGN U10062 ( .B(clk), .A(\g.we_clk [6328]));
Q_ASSIGN U10063 ( .B(clk), .A(\g.we_clk [6327]));
Q_ASSIGN U10064 ( .B(clk), .A(\g.we_clk [6326]));
Q_ASSIGN U10065 ( .B(clk), .A(\g.we_clk [6325]));
Q_ASSIGN U10066 ( .B(clk), .A(\g.we_clk [6324]));
Q_ASSIGN U10067 ( .B(clk), .A(\g.we_clk [6323]));
Q_ASSIGN U10068 ( .B(clk), .A(\g.we_clk [6322]));
Q_ASSIGN U10069 ( .B(clk), .A(\g.we_clk [6321]));
Q_ASSIGN U10070 ( .B(clk), .A(\g.we_clk [6320]));
Q_ASSIGN U10071 ( .B(clk), .A(\g.we_clk [6319]));
Q_ASSIGN U10072 ( .B(clk), .A(\g.we_clk [6318]));
Q_ASSIGN U10073 ( .B(clk), .A(\g.we_clk [6317]));
Q_ASSIGN U10074 ( .B(clk), .A(\g.we_clk [6316]));
Q_ASSIGN U10075 ( .B(clk), .A(\g.we_clk [6315]));
Q_ASSIGN U10076 ( .B(clk), .A(\g.we_clk [6314]));
Q_ASSIGN U10077 ( .B(clk), .A(\g.we_clk [6313]));
Q_ASSIGN U10078 ( .B(clk), .A(\g.we_clk [6312]));
Q_ASSIGN U10079 ( .B(clk), .A(\g.we_clk [6311]));
Q_ASSIGN U10080 ( .B(clk), .A(\g.we_clk [6310]));
Q_ASSIGN U10081 ( .B(clk), .A(\g.we_clk [6309]));
Q_ASSIGN U10082 ( .B(clk), .A(\g.we_clk [6308]));
Q_ASSIGN U10083 ( .B(clk), .A(\g.we_clk [6307]));
Q_ASSIGN U10084 ( .B(clk), .A(\g.we_clk [6306]));
Q_ASSIGN U10085 ( .B(clk), .A(\g.we_clk [6305]));
Q_ASSIGN U10086 ( .B(clk), .A(\g.we_clk [6304]));
Q_ASSIGN U10087 ( .B(clk), .A(\g.we_clk [6303]));
Q_ASSIGN U10088 ( .B(clk), .A(\g.we_clk [6302]));
Q_ASSIGN U10089 ( .B(clk), .A(\g.we_clk [6301]));
Q_ASSIGN U10090 ( .B(clk), .A(\g.we_clk [6300]));
Q_ASSIGN U10091 ( .B(clk), .A(\g.we_clk [6299]));
Q_ASSIGN U10092 ( .B(clk), .A(\g.we_clk [6298]));
Q_ASSIGN U10093 ( .B(clk), .A(\g.we_clk [6297]));
Q_ASSIGN U10094 ( .B(clk), .A(\g.we_clk [6296]));
Q_ASSIGN U10095 ( .B(clk), .A(\g.we_clk [6295]));
Q_ASSIGN U10096 ( .B(clk), .A(\g.we_clk [6294]));
Q_ASSIGN U10097 ( .B(clk), .A(\g.we_clk [6293]));
Q_ASSIGN U10098 ( .B(clk), .A(\g.we_clk [6292]));
Q_ASSIGN U10099 ( .B(clk), .A(\g.we_clk [6291]));
Q_ASSIGN U10100 ( .B(clk), .A(\g.we_clk [6290]));
Q_ASSIGN U10101 ( .B(clk), .A(\g.we_clk [6289]));
Q_ASSIGN U10102 ( .B(clk), .A(\g.we_clk [6288]));
Q_ASSIGN U10103 ( .B(clk), .A(\g.we_clk [6287]));
Q_ASSIGN U10104 ( .B(clk), .A(\g.we_clk [6286]));
Q_ASSIGN U10105 ( .B(clk), .A(\g.we_clk [6285]));
Q_ASSIGN U10106 ( .B(clk), .A(\g.we_clk [6284]));
Q_ASSIGN U10107 ( .B(clk), .A(\g.we_clk [6283]));
Q_ASSIGN U10108 ( .B(clk), .A(\g.we_clk [6282]));
Q_ASSIGN U10109 ( .B(clk), .A(\g.we_clk [6281]));
Q_ASSIGN U10110 ( .B(clk), .A(\g.we_clk [6280]));
Q_ASSIGN U10111 ( .B(clk), .A(\g.we_clk [6279]));
Q_ASSIGN U10112 ( .B(clk), .A(\g.we_clk [6278]));
Q_ASSIGN U10113 ( .B(clk), .A(\g.we_clk [6277]));
Q_ASSIGN U10114 ( .B(clk), .A(\g.we_clk [6276]));
Q_ASSIGN U10115 ( .B(clk), .A(\g.we_clk [6275]));
Q_ASSIGN U10116 ( .B(clk), .A(\g.we_clk [6274]));
Q_ASSIGN U10117 ( .B(clk), .A(\g.we_clk [6273]));
Q_ASSIGN U10118 ( .B(clk), .A(\g.we_clk [6272]));
Q_ASSIGN U10119 ( .B(clk), .A(\g.we_clk [6271]));
Q_ASSIGN U10120 ( .B(clk), .A(\g.we_clk [6270]));
Q_ASSIGN U10121 ( .B(clk), .A(\g.we_clk [6269]));
Q_ASSIGN U10122 ( .B(clk), .A(\g.we_clk [6268]));
Q_ASSIGN U10123 ( .B(clk), .A(\g.we_clk [6267]));
Q_ASSIGN U10124 ( .B(clk), .A(\g.we_clk [6266]));
Q_ASSIGN U10125 ( .B(clk), .A(\g.we_clk [6265]));
Q_ASSIGN U10126 ( .B(clk), .A(\g.we_clk [6264]));
Q_ASSIGN U10127 ( .B(clk), .A(\g.we_clk [6263]));
Q_ASSIGN U10128 ( .B(clk), .A(\g.we_clk [6262]));
Q_ASSIGN U10129 ( .B(clk), .A(\g.we_clk [6261]));
Q_ASSIGN U10130 ( .B(clk), .A(\g.we_clk [6260]));
Q_ASSIGN U10131 ( .B(clk), .A(\g.we_clk [6259]));
Q_ASSIGN U10132 ( .B(clk), .A(\g.we_clk [6258]));
Q_ASSIGN U10133 ( .B(clk), .A(\g.we_clk [6257]));
Q_ASSIGN U10134 ( .B(clk), .A(\g.we_clk [6256]));
Q_ASSIGN U10135 ( .B(clk), .A(\g.we_clk [6255]));
Q_ASSIGN U10136 ( .B(clk), .A(\g.we_clk [6254]));
Q_ASSIGN U10137 ( .B(clk), .A(\g.we_clk [6253]));
Q_ASSIGN U10138 ( .B(clk), .A(\g.we_clk [6252]));
Q_ASSIGN U10139 ( .B(clk), .A(\g.we_clk [6251]));
Q_ASSIGN U10140 ( .B(clk), .A(\g.we_clk [6250]));
Q_ASSIGN U10141 ( .B(clk), .A(\g.we_clk [6249]));
Q_ASSIGN U10142 ( .B(clk), .A(\g.we_clk [6248]));
Q_ASSIGN U10143 ( .B(clk), .A(\g.we_clk [6247]));
Q_ASSIGN U10144 ( .B(clk), .A(\g.we_clk [6246]));
Q_ASSIGN U10145 ( .B(clk), .A(\g.we_clk [6245]));
Q_ASSIGN U10146 ( .B(clk), .A(\g.we_clk [6244]));
Q_ASSIGN U10147 ( .B(clk), .A(\g.we_clk [6243]));
Q_ASSIGN U10148 ( .B(clk), .A(\g.we_clk [6242]));
Q_ASSIGN U10149 ( .B(clk), .A(\g.we_clk [6241]));
Q_ASSIGN U10150 ( .B(clk), .A(\g.we_clk [6240]));
Q_ASSIGN U10151 ( .B(clk), .A(\g.we_clk [6239]));
Q_ASSIGN U10152 ( .B(clk), .A(\g.we_clk [6238]));
Q_ASSIGN U10153 ( .B(clk), .A(\g.we_clk [6237]));
Q_ASSIGN U10154 ( .B(clk), .A(\g.we_clk [6236]));
Q_ASSIGN U10155 ( .B(clk), .A(\g.we_clk [6235]));
Q_ASSIGN U10156 ( .B(clk), .A(\g.we_clk [6234]));
Q_ASSIGN U10157 ( .B(clk), .A(\g.we_clk [6233]));
Q_ASSIGN U10158 ( .B(clk), .A(\g.we_clk [6232]));
Q_ASSIGN U10159 ( .B(clk), .A(\g.we_clk [6231]));
Q_ASSIGN U10160 ( .B(clk), .A(\g.we_clk [6230]));
Q_ASSIGN U10161 ( .B(clk), .A(\g.we_clk [6229]));
Q_ASSIGN U10162 ( .B(clk), .A(\g.we_clk [6228]));
Q_ASSIGN U10163 ( .B(clk), .A(\g.we_clk [6227]));
Q_ASSIGN U10164 ( .B(clk), .A(\g.we_clk [6226]));
Q_ASSIGN U10165 ( .B(clk), .A(\g.we_clk [6225]));
Q_ASSIGN U10166 ( .B(clk), .A(\g.we_clk [6224]));
Q_ASSIGN U10167 ( .B(clk), .A(\g.we_clk [6223]));
Q_ASSIGN U10168 ( .B(clk), .A(\g.we_clk [6222]));
Q_ASSIGN U10169 ( .B(clk), .A(\g.we_clk [6221]));
Q_ASSIGN U10170 ( .B(clk), .A(\g.we_clk [6220]));
Q_ASSIGN U10171 ( .B(clk), .A(\g.we_clk [6219]));
Q_ASSIGN U10172 ( .B(clk), .A(\g.we_clk [6218]));
Q_ASSIGN U10173 ( .B(clk), .A(\g.we_clk [6217]));
Q_ASSIGN U10174 ( .B(clk), .A(\g.we_clk [6216]));
Q_ASSIGN U10175 ( .B(clk), .A(\g.we_clk [6215]));
Q_ASSIGN U10176 ( .B(clk), .A(\g.we_clk [6214]));
Q_ASSIGN U10177 ( .B(clk), .A(\g.we_clk [6213]));
Q_ASSIGN U10178 ( .B(clk), .A(\g.we_clk [6212]));
Q_ASSIGN U10179 ( .B(clk), .A(\g.we_clk [6211]));
Q_ASSIGN U10180 ( .B(clk), .A(\g.we_clk [6210]));
Q_ASSIGN U10181 ( .B(clk), .A(\g.we_clk [6209]));
Q_ASSIGN U10182 ( .B(clk), .A(\g.we_clk [6208]));
Q_ASSIGN U10183 ( .B(clk), .A(\g.we_clk [6207]));
Q_ASSIGN U10184 ( .B(clk), .A(\g.we_clk [6206]));
Q_ASSIGN U10185 ( .B(clk), .A(\g.we_clk [6205]));
Q_ASSIGN U10186 ( .B(clk), .A(\g.we_clk [6204]));
Q_ASSIGN U10187 ( .B(clk), .A(\g.we_clk [6203]));
Q_ASSIGN U10188 ( .B(clk), .A(\g.we_clk [6202]));
Q_ASSIGN U10189 ( .B(clk), .A(\g.we_clk [6201]));
Q_ASSIGN U10190 ( .B(clk), .A(\g.we_clk [6200]));
Q_ASSIGN U10191 ( .B(clk), .A(\g.we_clk [6199]));
Q_ASSIGN U10192 ( .B(clk), .A(\g.we_clk [6198]));
Q_ASSIGN U10193 ( .B(clk), .A(\g.we_clk [6197]));
Q_ASSIGN U10194 ( .B(clk), .A(\g.we_clk [6196]));
Q_ASSIGN U10195 ( .B(clk), .A(\g.we_clk [6195]));
Q_ASSIGN U10196 ( .B(clk), .A(\g.we_clk [6194]));
Q_ASSIGN U10197 ( .B(clk), .A(\g.we_clk [6193]));
Q_ASSIGN U10198 ( .B(clk), .A(\g.we_clk [6192]));
Q_ASSIGN U10199 ( .B(clk), .A(\g.we_clk [6191]));
Q_ASSIGN U10200 ( .B(clk), .A(\g.we_clk [6190]));
Q_ASSIGN U10201 ( .B(clk), .A(\g.we_clk [6189]));
Q_ASSIGN U10202 ( .B(clk), .A(\g.we_clk [6188]));
Q_ASSIGN U10203 ( .B(clk), .A(\g.we_clk [6187]));
Q_ASSIGN U10204 ( .B(clk), .A(\g.we_clk [6186]));
Q_ASSIGN U10205 ( .B(clk), .A(\g.we_clk [6185]));
Q_ASSIGN U10206 ( .B(clk), .A(\g.we_clk [6184]));
Q_ASSIGN U10207 ( .B(clk), .A(\g.we_clk [6183]));
Q_ASSIGN U10208 ( .B(clk), .A(\g.we_clk [6182]));
Q_ASSIGN U10209 ( .B(clk), .A(\g.we_clk [6181]));
Q_ASSIGN U10210 ( .B(clk), .A(\g.we_clk [6180]));
Q_ASSIGN U10211 ( .B(clk), .A(\g.we_clk [6179]));
Q_ASSIGN U10212 ( .B(clk), .A(\g.we_clk [6178]));
Q_ASSIGN U10213 ( .B(clk), .A(\g.we_clk [6177]));
Q_ASSIGN U10214 ( .B(clk), .A(\g.we_clk [6176]));
Q_ASSIGN U10215 ( .B(clk), .A(\g.we_clk [6175]));
Q_ASSIGN U10216 ( .B(clk), .A(\g.we_clk [6174]));
Q_ASSIGN U10217 ( .B(clk), .A(\g.we_clk [6173]));
Q_ASSIGN U10218 ( .B(clk), .A(\g.we_clk [6172]));
Q_ASSIGN U10219 ( .B(clk), .A(\g.we_clk [6171]));
Q_ASSIGN U10220 ( .B(clk), .A(\g.we_clk [6170]));
Q_ASSIGN U10221 ( .B(clk), .A(\g.we_clk [6169]));
Q_ASSIGN U10222 ( .B(clk), .A(\g.we_clk [6168]));
Q_ASSIGN U10223 ( .B(clk), .A(\g.we_clk [6167]));
Q_ASSIGN U10224 ( .B(clk), .A(\g.we_clk [6166]));
Q_ASSIGN U10225 ( .B(clk), .A(\g.we_clk [6165]));
Q_ASSIGN U10226 ( .B(clk), .A(\g.we_clk [6164]));
Q_ASSIGN U10227 ( .B(clk), .A(\g.we_clk [6163]));
Q_ASSIGN U10228 ( .B(clk), .A(\g.we_clk [6162]));
Q_ASSIGN U10229 ( .B(clk), .A(\g.we_clk [6161]));
Q_ASSIGN U10230 ( .B(clk), .A(\g.we_clk [6160]));
Q_ASSIGN U10231 ( .B(clk), .A(\g.we_clk [6159]));
Q_ASSIGN U10232 ( .B(clk), .A(\g.we_clk [6158]));
Q_ASSIGN U10233 ( .B(clk), .A(\g.we_clk [6157]));
Q_ASSIGN U10234 ( .B(clk), .A(\g.we_clk [6156]));
Q_ASSIGN U10235 ( .B(clk), .A(\g.we_clk [6155]));
Q_ASSIGN U10236 ( .B(clk), .A(\g.we_clk [6154]));
Q_ASSIGN U10237 ( .B(clk), .A(\g.we_clk [6153]));
Q_ASSIGN U10238 ( .B(clk), .A(\g.we_clk [6152]));
Q_ASSIGN U10239 ( .B(clk), .A(\g.we_clk [6151]));
Q_ASSIGN U10240 ( .B(clk), .A(\g.we_clk [6150]));
Q_ASSIGN U10241 ( .B(clk), .A(\g.we_clk [6149]));
Q_ASSIGN U10242 ( .B(clk), .A(\g.we_clk [6148]));
Q_ASSIGN U10243 ( .B(clk), .A(\g.we_clk [6147]));
Q_ASSIGN U10244 ( .B(clk), .A(\g.we_clk [6146]));
Q_ASSIGN U10245 ( .B(clk), .A(\g.we_clk [6145]));
Q_ASSIGN U10246 ( .B(clk), .A(\g.we_clk [6144]));
Q_ASSIGN U10247 ( .B(clk), .A(\g.we_clk [6143]));
Q_ASSIGN U10248 ( .B(clk), .A(\g.we_clk [6142]));
Q_ASSIGN U10249 ( .B(clk), .A(\g.we_clk [6141]));
Q_ASSIGN U10250 ( .B(clk), .A(\g.we_clk [6140]));
Q_ASSIGN U10251 ( .B(clk), .A(\g.we_clk [6139]));
Q_ASSIGN U10252 ( .B(clk), .A(\g.we_clk [6138]));
Q_ASSIGN U10253 ( .B(clk), .A(\g.we_clk [6137]));
Q_ASSIGN U10254 ( .B(clk), .A(\g.we_clk [6136]));
Q_ASSIGN U10255 ( .B(clk), .A(\g.we_clk [6135]));
Q_ASSIGN U10256 ( .B(clk), .A(\g.we_clk [6134]));
Q_ASSIGN U10257 ( .B(clk), .A(\g.we_clk [6133]));
Q_ASSIGN U10258 ( .B(clk), .A(\g.we_clk [6132]));
Q_ASSIGN U10259 ( .B(clk), .A(\g.we_clk [6131]));
Q_ASSIGN U10260 ( .B(clk), .A(\g.we_clk [6130]));
Q_ASSIGN U10261 ( .B(clk), .A(\g.we_clk [6129]));
Q_ASSIGN U10262 ( .B(clk), .A(\g.we_clk [6128]));
Q_ASSIGN U10263 ( .B(clk), .A(\g.we_clk [6127]));
Q_ASSIGN U10264 ( .B(clk), .A(\g.we_clk [6126]));
Q_ASSIGN U10265 ( .B(clk), .A(\g.we_clk [6125]));
Q_ASSIGN U10266 ( .B(clk), .A(\g.we_clk [6124]));
Q_ASSIGN U10267 ( .B(clk), .A(\g.we_clk [6123]));
Q_ASSIGN U10268 ( .B(clk), .A(\g.we_clk [6122]));
Q_ASSIGN U10269 ( .B(clk), .A(\g.we_clk [6121]));
Q_ASSIGN U10270 ( .B(clk), .A(\g.we_clk [6120]));
Q_ASSIGN U10271 ( .B(clk), .A(\g.we_clk [6119]));
Q_ASSIGN U10272 ( .B(clk), .A(\g.we_clk [6118]));
Q_ASSIGN U10273 ( .B(clk), .A(\g.we_clk [6117]));
Q_ASSIGN U10274 ( .B(clk), .A(\g.we_clk [6116]));
Q_ASSIGN U10275 ( .B(clk), .A(\g.we_clk [6115]));
Q_ASSIGN U10276 ( .B(clk), .A(\g.we_clk [6114]));
Q_ASSIGN U10277 ( .B(clk), .A(\g.we_clk [6113]));
Q_ASSIGN U10278 ( .B(clk), .A(\g.we_clk [6112]));
Q_ASSIGN U10279 ( .B(clk), .A(\g.we_clk [6111]));
Q_ASSIGN U10280 ( .B(clk), .A(\g.we_clk [6110]));
Q_ASSIGN U10281 ( .B(clk), .A(\g.we_clk [6109]));
Q_ASSIGN U10282 ( .B(clk), .A(\g.we_clk [6108]));
Q_ASSIGN U10283 ( .B(clk), .A(\g.we_clk [6107]));
Q_ASSIGN U10284 ( .B(clk), .A(\g.we_clk [6106]));
Q_ASSIGN U10285 ( .B(clk), .A(\g.we_clk [6105]));
Q_ASSIGN U10286 ( .B(clk), .A(\g.we_clk [6104]));
Q_ASSIGN U10287 ( .B(clk), .A(\g.we_clk [6103]));
Q_ASSIGN U10288 ( .B(clk), .A(\g.we_clk [6102]));
Q_ASSIGN U10289 ( .B(clk), .A(\g.we_clk [6101]));
Q_ASSIGN U10290 ( .B(clk), .A(\g.we_clk [6100]));
Q_ASSIGN U10291 ( .B(clk), .A(\g.we_clk [6099]));
Q_ASSIGN U10292 ( .B(clk), .A(\g.we_clk [6098]));
Q_ASSIGN U10293 ( .B(clk), .A(\g.we_clk [6097]));
Q_ASSIGN U10294 ( .B(clk), .A(\g.we_clk [6096]));
Q_ASSIGN U10295 ( .B(clk), .A(\g.we_clk [6095]));
Q_ASSIGN U10296 ( .B(clk), .A(\g.we_clk [6094]));
Q_ASSIGN U10297 ( .B(clk), .A(\g.we_clk [6093]));
Q_ASSIGN U10298 ( .B(clk), .A(\g.we_clk [6092]));
Q_ASSIGN U10299 ( .B(clk), .A(\g.we_clk [6091]));
Q_ASSIGN U10300 ( .B(clk), .A(\g.we_clk [6090]));
Q_ASSIGN U10301 ( .B(clk), .A(\g.we_clk [6089]));
Q_ASSIGN U10302 ( .B(clk), .A(\g.we_clk [6088]));
Q_ASSIGN U10303 ( .B(clk), .A(\g.we_clk [6087]));
Q_ASSIGN U10304 ( .B(clk), .A(\g.we_clk [6086]));
Q_ASSIGN U10305 ( .B(clk), .A(\g.we_clk [6085]));
Q_ASSIGN U10306 ( .B(clk), .A(\g.we_clk [6084]));
Q_ASSIGN U10307 ( .B(clk), .A(\g.we_clk [6083]));
Q_ASSIGN U10308 ( .B(clk), .A(\g.we_clk [6082]));
Q_ASSIGN U10309 ( .B(clk), .A(\g.we_clk [6081]));
Q_ASSIGN U10310 ( .B(clk), .A(\g.we_clk [6080]));
Q_ASSIGN U10311 ( .B(clk), .A(\g.we_clk [6079]));
Q_ASSIGN U10312 ( .B(clk), .A(\g.we_clk [6078]));
Q_ASSIGN U10313 ( .B(clk), .A(\g.we_clk [6077]));
Q_ASSIGN U10314 ( .B(clk), .A(\g.we_clk [6076]));
Q_ASSIGN U10315 ( .B(clk), .A(\g.we_clk [6075]));
Q_ASSIGN U10316 ( .B(clk), .A(\g.we_clk [6074]));
Q_ASSIGN U10317 ( .B(clk), .A(\g.we_clk [6073]));
Q_ASSIGN U10318 ( .B(clk), .A(\g.we_clk [6072]));
Q_ASSIGN U10319 ( .B(clk), .A(\g.we_clk [6071]));
Q_ASSIGN U10320 ( .B(clk), .A(\g.we_clk [6070]));
Q_ASSIGN U10321 ( .B(clk), .A(\g.we_clk [6069]));
Q_ASSIGN U10322 ( .B(clk), .A(\g.we_clk [6068]));
Q_ASSIGN U10323 ( .B(clk), .A(\g.we_clk [6067]));
Q_ASSIGN U10324 ( .B(clk), .A(\g.we_clk [6066]));
Q_ASSIGN U10325 ( .B(clk), .A(\g.we_clk [6065]));
Q_ASSIGN U10326 ( .B(clk), .A(\g.we_clk [6064]));
Q_ASSIGN U10327 ( .B(clk), .A(\g.we_clk [6063]));
Q_ASSIGN U10328 ( .B(clk), .A(\g.we_clk [6062]));
Q_ASSIGN U10329 ( .B(clk), .A(\g.we_clk [6061]));
Q_ASSIGN U10330 ( .B(clk), .A(\g.we_clk [6060]));
Q_ASSIGN U10331 ( .B(clk), .A(\g.we_clk [6059]));
Q_ASSIGN U10332 ( .B(clk), .A(\g.we_clk [6058]));
Q_ASSIGN U10333 ( .B(clk), .A(\g.we_clk [6057]));
Q_ASSIGN U10334 ( .B(clk), .A(\g.we_clk [6056]));
Q_ASSIGN U10335 ( .B(clk), .A(\g.we_clk [6055]));
Q_ASSIGN U10336 ( .B(clk), .A(\g.we_clk [6054]));
Q_ASSIGN U10337 ( .B(clk), .A(\g.we_clk [6053]));
Q_ASSIGN U10338 ( .B(clk), .A(\g.we_clk [6052]));
Q_ASSIGN U10339 ( .B(clk), .A(\g.we_clk [6051]));
Q_ASSIGN U10340 ( .B(clk), .A(\g.we_clk [6050]));
Q_ASSIGN U10341 ( .B(clk), .A(\g.we_clk [6049]));
Q_ASSIGN U10342 ( .B(clk), .A(\g.we_clk [6048]));
Q_ASSIGN U10343 ( .B(clk), .A(\g.we_clk [6047]));
Q_ASSIGN U10344 ( .B(clk), .A(\g.we_clk [6046]));
Q_ASSIGN U10345 ( .B(clk), .A(\g.we_clk [6045]));
Q_ASSIGN U10346 ( .B(clk), .A(\g.we_clk [6044]));
Q_ASSIGN U10347 ( .B(clk), .A(\g.we_clk [6043]));
Q_ASSIGN U10348 ( .B(clk), .A(\g.we_clk [6042]));
Q_ASSIGN U10349 ( .B(clk), .A(\g.we_clk [6041]));
Q_ASSIGN U10350 ( .B(clk), .A(\g.we_clk [6040]));
Q_ASSIGN U10351 ( .B(clk), .A(\g.we_clk [6039]));
Q_ASSIGN U10352 ( .B(clk), .A(\g.we_clk [6038]));
Q_ASSIGN U10353 ( .B(clk), .A(\g.we_clk [6037]));
Q_ASSIGN U10354 ( .B(clk), .A(\g.we_clk [6036]));
Q_ASSIGN U10355 ( .B(clk), .A(\g.we_clk [6035]));
Q_ASSIGN U10356 ( .B(clk), .A(\g.we_clk [6034]));
Q_ASSIGN U10357 ( .B(clk), .A(\g.we_clk [6033]));
Q_ASSIGN U10358 ( .B(clk), .A(\g.we_clk [6032]));
Q_ASSIGN U10359 ( .B(clk), .A(\g.we_clk [6031]));
Q_ASSIGN U10360 ( .B(clk), .A(\g.we_clk [6030]));
Q_ASSIGN U10361 ( .B(clk), .A(\g.we_clk [6029]));
Q_ASSIGN U10362 ( .B(clk), .A(\g.we_clk [6028]));
Q_ASSIGN U10363 ( .B(clk), .A(\g.we_clk [6027]));
Q_ASSIGN U10364 ( .B(clk), .A(\g.we_clk [6026]));
Q_ASSIGN U10365 ( .B(clk), .A(\g.we_clk [6025]));
Q_ASSIGN U10366 ( .B(clk), .A(\g.we_clk [6024]));
Q_ASSIGN U10367 ( .B(clk), .A(\g.we_clk [6023]));
Q_ASSIGN U10368 ( .B(clk), .A(\g.we_clk [6022]));
Q_ASSIGN U10369 ( .B(clk), .A(\g.we_clk [6021]));
Q_ASSIGN U10370 ( .B(clk), .A(\g.we_clk [6020]));
Q_ASSIGN U10371 ( .B(clk), .A(\g.we_clk [6019]));
Q_ASSIGN U10372 ( .B(clk), .A(\g.we_clk [6018]));
Q_ASSIGN U10373 ( .B(clk), .A(\g.we_clk [6017]));
Q_ASSIGN U10374 ( .B(clk), .A(\g.we_clk [6016]));
Q_ASSIGN U10375 ( .B(clk), .A(\g.we_clk [6015]));
Q_ASSIGN U10376 ( .B(clk), .A(\g.we_clk [6014]));
Q_ASSIGN U10377 ( .B(clk), .A(\g.we_clk [6013]));
Q_ASSIGN U10378 ( .B(clk), .A(\g.we_clk [6012]));
Q_ASSIGN U10379 ( .B(clk), .A(\g.we_clk [6011]));
Q_ASSIGN U10380 ( .B(clk), .A(\g.we_clk [6010]));
Q_ASSIGN U10381 ( .B(clk), .A(\g.we_clk [6009]));
Q_ASSIGN U10382 ( .B(clk), .A(\g.we_clk [6008]));
Q_ASSIGN U10383 ( .B(clk), .A(\g.we_clk [6007]));
Q_ASSIGN U10384 ( .B(clk), .A(\g.we_clk [6006]));
Q_ASSIGN U10385 ( .B(clk), .A(\g.we_clk [6005]));
Q_ASSIGN U10386 ( .B(clk), .A(\g.we_clk [6004]));
Q_ASSIGN U10387 ( .B(clk), .A(\g.we_clk [6003]));
Q_ASSIGN U10388 ( .B(clk), .A(\g.we_clk [6002]));
Q_ASSIGN U10389 ( .B(clk), .A(\g.we_clk [6001]));
Q_ASSIGN U10390 ( .B(clk), .A(\g.we_clk [6000]));
Q_ASSIGN U10391 ( .B(clk), .A(\g.we_clk [5999]));
Q_ASSIGN U10392 ( .B(clk), .A(\g.we_clk [5998]));
Q_ASSIGN U10393 ( .B(clk), .A(\g.we_clk [5997]));
Q_ASSIGN U10394 ( .B(clk), .A(\g.we_clk [5996]));
Q_ASSIGN U10395 ( .B(clk), .A(\g.we_clk [5995]));
Q_ASSIGN U10396 ( .B(clk), .A(\g.we_clk [5994]));
Q_ASSIGN U10397 ( .B(clk), .A(\g.we_clk [5993]));
Q_ASSIGN U10398 ( .B(clk), .A(\g.we_clk [5992]));
Q_ASSIGN U10399 ( .B(clk), .A(\g.we_clk [5991]));
Q_ASSIGN U10400 ( .B(clk), .A(\g.we_clk [5990]));
Q_ASSIGN U10401 ( .B(clk), .A(\g.we_clk [5989]));
Q_ASSIGN U10402 ( .B(clk), .A(\g.we_clk [5988]));
Q_ASSIGN U10403 ( .B(clk), .A(\g.we_clk [5987]));
Q_ASSIGN U10404 ( .B(clk), .A(\g.we_clk [5986]));
Q_ASSIGN U10405 ( .B(clk), .A(\g.we_clk [5985]));
Q_ASSIGN U10406 ( .B(clk), .A(\g.we_clk [5984]));
Q_ASSIGN U10407 ( .B(clk), .A(\g.we_clk [5983]));
Q_ASSIGN U10408 ( .B(clk), .A(\g.we_clk [5982]));
Q_ASSIGN U10409 ( .B(clk), .A(\g.we_clk [5981]));
Q_ASSIGN U10410 ( .B(clk), .A(\g.we_clk [5980]));
Q_ASSIGN U10411 ( .B(clk), .A(\g.we_clk [5979]));
Q_ASSIGN U10412 ( .B(clk), .A(\g.we_clk [5978]));
Q_ASSIGN U10413 ( .B(clk), .A(\g.we_clk [5977]));
Q_ASSIGN U10414 ( .B(clk), .A(\g.we_clk [5976]));
Q_ASSIGN U10415 ( .B(clk), .A(\g.we_clk [5975]));
Q_ASSIGN U10416 ( .B(clk), .A(\g.we_clk [5974]));
Q_ASSIGN U10417 ( .B(clk), .A(\g.we_clk [5973]));
Q_ASSIGN U10418 ( .B(clk), .A(\g.we_clk [5972]));
Q_ASSIGN U10419 ( .B(clk), .A(\g.we_clk [5971]));
Q_ASSIGN U10420 ( .B(clk), .A(\g.we_clk [5970]));
Q_ASSIGN U10421 ( .B(clk), .A(\g.we_clk [5969]));
Q_ASSIGN U10422 ( .B(clk), .A(\g.we_clk [5968]));
Q_ASSIGN U10423 ( .B(clk), .A(\g.we_clk [5967]));
Q_ASSIGN U10424 ( .B(clk), .A(\g.we_clk [5966]));
Q_ASSIGN U10425 ( .B(clk), .A(\g.we_clk [5965]));
Q_ASSIGN U10426 ( .B(clk), .A(\g.we_clk [5964]));
Q_ASSIGN U10427 ( .B(clk), .A(\g.we_clk [5963]));
Q_ASSIGN U10428 ( .B(clk), .A(\g.we_clk [5962]));
Q_ASSIGN U10429 ( .B(clk), .A(\g.we_clk [5961]));
Q_ASSIGN U10430 ( .B(clk), .A(\g.we_clk [5960]));
Q_ASSIGN U10431 ( .B(clk), .A(\g.we_clk [5959]));
Q_ASSIGN U10432 ( .B(clk), .A(\g.we_clk [5958]));
Q_ASSIGN U10433 ( .B(clk), .A(\g.we_clk [5957]));
Q_ASSIGN U10434 ( .B(clk), .A(\g.we_clk [5956]));
Q_ASSIGN U10435 ( .B(clk), .A(\g.we_clk [5955]));
Q_ASSIGN U10436 ( .B(clk), .A(\g.we_clk [5954]));
Q_ASSIGN U10437 ( .B(clk), .A(\g.we_clk [5953]));
Q_ASSIGN U10438 ( .B(clk), .A(\g.we_clk [5952]));
Q_ASSIGN U10439 ( .B(clk), .A(\g.we_clk [5951]));
Q_ASSIGN U10440 ( .B(clk), .A(\g.we_clk [5950]));
Q_ASSIGN U10441 ( .B(clk), .A(\g.we_clk [5949]));
Q_ASSIGN U10442 ( .B(clk), .A(\g.we_clk [5948]));
Q_ASSIGN U10443 ( .B(clk), .A(\g.we_clk [5947]));
Q_ASSIGN U10444 ( .B(clk), .A(\g.we_clk [5946]));
Q_ASSIGN U10445 ( .B(clk), .A(\g.we_clk [5945]));
Q_ASSIGN U10446 ( .B(clk), .A(\g.we_clk [5944]));
Q_ASSIGN U10447 ( .B(clk), .A(\g.we_clk [5943]));
Q_ASSIGN U10448 ( .B(clk), .A(\g.we_clk [5942]));
Q_ASSIGN U10449 ( .B(clk), .A(\g.we_clk [5941]));
Q_ASSIGN U10450 ( .B(clk), .A(\g.we_clk [5940]));
Q_ASSIGN U10451 ( .B(clk), .A(\g.we_clk [5939]));
Q_ASSIGN U10452 ( .B(clk), .A(\g.we_clk [5938]));
Q_ASSIGN U10453 ( .B(clk), .A(\g.we_clk [5937]));
Q_ASSIGN U10454 ( .B(clk), .A(\g.we_clk [5936]));
Q_ASSIGN U10455 ( .B(clk), .A(\g.we_clk [5935]));
Q_ASSIGN U10456 ( .B(clk), .A(\g.we_clk [5934]));
Q_ASSIGN U10457 ( .B(clk), .A(\g.we_clk [5933]));
Q_ASSIGN U10458 ( .B(clk), .A(\g.we_clk [5932]));
Q_ASSIGN U10459 ( .B(clk), .A(\g.we_clk [5931]));
Q_ASSIGN U10460 ( .B(clk), .A(\g.we_clk [5930]));
Q_ASSIGN U10461 ( .B(clk), .A(\g.we_clk [5929]));
Q_ASSIGN U10462 ( .B(clk), .A(\g.we_clk [5928]));
Q_ASSIGN U10463 ( .B(clk), .A(\g.we_clk [5927]));
Q_ASSIGN U10464 ( .B(clk), .A(\g.we_clk [5926]));
Q_ASSIGN U10465 ( .B(clk), .A(\g.we_clk [5925]));
Q_ASSIGN U10466 ( .B(clk), .A(\g.we_clk [5924]));
Q_ASSIGN U10467 ( .B(clk), .A(\g.we_clk [5923]));
Q_ASSIGN U10468 ( .B(clk), .A(\g.we_clk [5922]));
Q_ASSIGN U10469 ( .B(clk), .A(\g.we_clk [5921]));
Q_ASSIGN U10470 ( .B(clk), .A(\g.we_clk [5920]));
Q_ASSIGN U10471 ( .B(clk), .A(\g.we_clk [5919]));
Q_ASSIGN U10472 ( .B(clk), .A(\g.we_clk [5918]));
Q_ASSIGN U10473 ( .B(clk), .A(\g.we_clk [5917]));
Q_ASSIGN U10474 ( .B(clk), .A(\g.we_clk [5916]));
Q_ASSIGN U10475 ( .B(clk), .A(\g.we_clk [5915]));
Q_ASSIGN U10476 ( .B(clk), .A(\g.we_clk [5914]));
Q_ASSIGN U10477 ( .B(clk), .A(\g.we_clk [5913]));
Q_ASSIGN U10478 ( .B(clk), .A(\g.we_clk [5912]));
Q_ASSIGN U10479 ( .B(clk), .A(\g.we_clk [5911]));
Q_ASSIGN U10480 ( .B(clk), .A(\g.we_clk [5910]));
Q_ASSIGN U10481 ( .B(clk), .A(\g.we_clk [5909]));
Q_ASSIGN U10482 ( .B(clk), .A(\g.we_clk [5908]));
Q_ASSIGN U10483 ( .B(clk), .A(\g.we_clk [5907]));
Q_ASSIGN U10484 ( .B(clk), .A(\g.we_clk [5906]));
Q_ASSIGN U10485 ( .B(clk), .A(\g.we_clk [5905]));
Q_ASSIGN U10486 ( .B(clk), .A(\g.we_clk [5904]));
Q_ASSIGN U10487 ( .B(clk), .A(\g.we_clk [5903]));
Q_ASSIGN U10488 ( .B(clk), .A(\g.we_clk [5902]));
Q_ASSIGN U10489 ( .B(clk), .A(\g.we_clk [5901]));
Q_ASSIGN U10490 ( .B(clk), .A(\g.we_clk [5900]));
Q_ASSIGN U10491 ( .B(clk), .A(\g.we_clk [5899]));
Q_ASSIGN U10492 ( .B(clk), .A(\g.we_clk [5898]));
Q_ASSIGN U10493 ( .B(clk), .A(\g.we_clk [5897]));
Q_ASSIGN U10494 ( .B(clk), .A(\g.we_clk [5896]));
Q_ASSIGN U10495 ( .B(clk), .A(\g.we_clk [5895]));
Q_ASSIGN U10496 ( .B(clk), .A(\g.we_clk [5894]));
Q_ASSIGN U10497 ( .B(clk), .A(\g.we_clk [5893]));
Q_ASSIGN U10498 ( .B(clk), .A(\g.we_clk [5892]));
Q_ASSIGN U10499 ( .B(clk), .A(\g.we_clk [5891]));
Q_ASSIGN U10500 ( .B(clk), .A(\g.we_clk [5890]));
Q_ASSIGN U10501 ( .B(clk), .A(\g.we_clk [5889]));
Q_ASSIGN U10502 ( .B(clk), .A(\g.we_clk [5888]));
Q_ASSIGN U10503 ( .B(clk), .A(\g.we_clk [5887]));
Q_ASSIGN U10504 ( .B(clk), .A(\g.we_clk [5886]));
Q_ASSIGN U10505 ( .B(clk), .A(\g.we_clk [5885]));
Q_ASSIGN U10506 ( .B(clk), .A(\g.we_clk [5884]));
Q_ASSIGN U10507 ( .B(clk), .A(\g.we_clk [5883]));
Q_ASSIGN U10508 ( .B(clk), .A(\g.we_clk [5882]));
Q_ASSIGN U10509 ( .B(clk), .A(\g.we_clk [5881]));
Q_ASSIGN U10510 ( .B(clk), .A(\g.we_clk [5880]));
Q_ASSIGN U10511 ( .B(clk), .A(\g.we_clk [5879]));
Q_ASSIGN U10512 ( .B(clk), .A(\g.we_clk [5878]));
Q_ASSIGN U10513 ( .B(clk), .A(\g.we_clk [5877]));
Q_ASSIGN U10514 ( .B(clk), .A(\g.we_clk [5876]));
Q_ASSIGN U10515 ( .B(clk), .A(\g.we_clk [5875]));
Q_ASSIGN U10516 ( .B(clk), .A(\g.we_clk [5874]));
Q_ASSIGN U10517 ( .B(clk), .A(\g.we_clk [5873]));
Q_ASSIGN U10518 ( .B(clk), .A(\g.we_clk [5872]));
Q_ASSIGN U10519 ( .B(clk), .A(\g.we_clk [5871]));
Q_ASSIGN U10520 ( .B(clk), .A(\g.we_clk [5870]));
Q_ASSIGN U10521 ( .B(clk), .A(\g.we_clk [5869]));
Q_ASSIGN U10522 ( .B(clk), .A(\g.we_clk [5868]));
Q_ASSIGN U10523 ( .B(clk), .A(\g.we_clk [5867]));
Q_ASSIGN U10524 ( .B(clk), .A(\g.we_clk [5866]));
Q_ASSIGN U10525 ( .B(clk), .A(\g.we_clk [5865]));
Q_ASSIGN U10526 ( .B(clk), .A(\g.we_clk [5864]));
Q_ASSIGN U10527 ( .B(clk), .A(\g.we_clk [5863]));
Q_ASSIGN U10528 ( .B(clk), .A(\g.we_clk [5862]));
Q_ASSIGN U10529 ( .B(clk), .A(\g.we_clk [5861]));
Q_ASSIGN U10530 ( .B(clk), .A(\g.we_clk [5860]));
Q_ASSIGN U10531 ( .B(clk), .A(\g.we_clk [5859]));
Q_ASSIGN U10532 ( .B(clk), .A(\g.we_clk [5858]));
Q_ASSIGN U10533 ( .B(clk), .A(\g.we_clk [5857]));
Q_ASSIGN U10534 ( .B(clk), .A(\g.we_clk [5856]));
Q_ASSIGN U10535 ( .B(clk), .A(\g.we_clk [5855]));
Q_ASSIGN U10536 ( .B(clk), .A(\g.we_clk [5854]));
Q_ASSIGN U10537 ( .B(clk), .A(\g.we_clk [5853]));
Q_ASSIGN U10538 ( .B(clk), .A(\g.we_clk [5852]));
Q_ASSIGN U10539 ( .B(clk), .A(\g.we_clk [5851]));
Q_ASSIGN U10540 ( .B(clk), .A(\g.we_clk [5850]));
Q_ASSIGN U10541 ( .B(clk), .A(\g.we_clk [5849]));
Q_ASSIGN U10542 ( .B(clk), .A(\g.we_clk [5848]));
Q_ASSIGN U10543 ( .B(clk), .A(\g.we_clk [5847]));
Q_ASSIGN U10544 ( .B(clk), .A(\g.we_clk [5846]));
Q_ASSIGN U10545 ( .B(clk), .A(\g.we_clk [5845]));
Q_ASSIGN U10546 ( .B(clk), .A(\g.we_clk [5844]));
Q_ASSIGN U10547 ( .B(clk), .A(\g.we_clk [5843]));
Q_ASSIGN U10548 ( .B(clk), .A(\g.we_clk [5842]));
Q_ASSIGN U10549 ( .B(clk), .A(\g.we_clk [5841]));
Q_ASSIGN U10550 ( .B(clk), .A(\g.we_clk [5840]));
Q_ASSIGN U10551 ( .B(clk), .A(\g.we_clk [5839]));
Q_ASSIGN U10552 ( .B(clk), .A(\g.we_clk [5838]));
Q_ASSIGN U10553 ( .B(clk), .A(\g.we_clk [5837]));
Q_ASSIGN U10554 ( .B(clk), .A(\g.we_clk [5836]));
Q_ASSIGN U10555 ( .B(clk), .A(\g.we_clk [5835]));
Q_ASSIGN U10556 ( .B(clk), .A(\g.we_clk [5834]));
Q_ASSIGN U10557 ( .B(clk), .A(\g.we_clk [5833]));
Q_ASSIGN U10558 ( .B(clk), .A(\g.we_clk [5832]));
Q_ASSIGN U10559 ( .B(clk), .A(\g.we_clk [5831]));
Q_ASSIGN U10560 ( .B(clk), .A(\g.we_clk [5830]));
Q_ASSIGN U10561 ( .B(clk), .A(\g.we_clk [5829]));
Q_ASSIGN U10562 ( .B(clk), .A(\g.we_clk [5828]));
Q_ASSIGN U10563 ( .B(clk), .A(\g.we_clk [5827]));
Q_ASSIGN U10564 ( .B(clk), .A(\g.we_clk [5826]));
Q_ASSIGN U10565 ( .B(clk), .A(\g.we_clk [5825]));
Q_ASSIGN U10566 ( .B(clk), .A(\g.we_clk [5824]));
Q_ASSIGN U10567 ( .B(clk), .A(\g.we_clk [5823]));
Q_ASSIGN U10568 ( .B(clk), .A(\g.we_clk [5822]));
Q_ASSIGN U10569 ( .B(clk), .A(\g.we_clk [5821]));
Q_ASSIGN U10570 ( .B(clk), .A(\g.we_clk [5820]));
Q_ASSIGN U10571 ( .B(clk), .A(\g.we_clk [5819]));
Q_ASSIGN U10572 ( .B(clk), .A(\g.we_clk [5818]));
Q_ASSIGN U10573 ( .B(clk), .A(\g.we_clk [5817]));
Q_ASSIGN U10574 ( .B(clk), .A(\g.we_clk [5816]));
Q_ASSIGN U10575 ( .B(clk), .A(\g.we_clk [5815]));
Q_ASSIGN U10576 ( .B(clk), .A(\g.we_clk [5814]));
Q_ASSIGN U10577 ( .B(clk), .A(\g.we_clk [5813]));
Q_ASSIGN U10578 ( .B(clk), .A(\g.we_clk [5812]));
Q_ASSIGN U10579 ( .B(clk), .A(\g.we_clk [5811]));
Q_ASSIGN U10580 ( .B(clk), .A(\g.we_clk [5810]));
Q_ASSIGN U10581 ( .B(clk), .A(\g.we_clk [5809]));
Q_ASSIGN U10582 ( .B(clk), .A(\g.we_clk [5808]));
Q_ASSIGN U10583 ( .B(clk), .A(\g.we_clk [5807]));
Q_ASSIGN U10584 ( .B(clk), .A(\g.we_clk [5806]));
Q_ASSIGN U10585 ( .B(clk), .A(\g.we_clk [5805]));
Q_ASSIGN U10586 ( .B(clk), .A(\g.we_clk [5804]));
Q_ASSIGN U10587 ( .B(clk), .A(\g.we_clk [5803]));
Q_ASSIGN U10588 ( .B(clk), .A(\g.we_clk [5802]));
Q_ASSIGN U10589 ( .B(clk), .A(\g.we_clk [5801]));
Q_ASSIGN U10590 ( .B(clk), .A(\g.we_clk [5800]));
Q_ASSIGN U10591 ( .B(clk), .A(\g.we_clk [5799]));
Q_ASSIGN U10592 ( .B(clk), .A(\g.we_clk [5798]));
Q_ASSIGN U10593 ( .B(clk), .A(\g.we_clk [5797]));
Q_ASSIGN U10594 ( .B(clk), .A(\g.we_clk [5796]));
Q_ASSIGN U10595 ( .B(clk), .A(\g.we_clk [5795]));
Q_ASSIGN U10596 ( .B(clk), .A(\g.we_clk [5794]));
Q_ASSIGN U10597 ( .B(clk), .A(\g.we_clk [5793]));
Q_ASSIGN U10598 ( .B(clk), .A(\g.we_clk [5792]));
Q_ASSIGN U10599 ( .B(clk), .A(\g.we_clk [5791]));
Q_ASSIGN U10600 ( .B(clk), .A(\g.we_clk [5790]));
Q_ASSIGN U10601 ( .B(clk), .A(\g.we_clk [5789]));
Q_ASSIGN U10602 ( .B(clk), .A(\g.we_clk [5788]));
Q_ASSIGN U10603 ( .B(clk), .A(\g.we_clk [5787]));
Q_ASSIGN U10604 ( .B(clk), .A(\g.we_clk [5786]));
Q_ASSIGN U10605 ( .B(clk), .A(\g.we_clk [5785]));
Q_ASSIGN U10606 ( .B(clk), .A(\g.we_clk [5784]));
Q_ASSIGN U10607 ( .B(clk), .A(\g.we_clk [5783]));
Q_ASSIGN U10608 ( .B(clk), .A(\g.we_clk [5782]));
Q_ASSIGN U10609 ( .B(clk), .A(\g.we_clk [5781]));
Q_ASSIGN U10610 ( .B(clk), .A(\g.we_clk [5780]));
Q_ASSIGN U10611 ( .B(clk), .A(\g.we_clk [5779]));
Q_ASSIGN U10612 ( .B(clk), .A(\g.we_clk [5778]));
Q_ASSIGN U10613 ( .B(clk), .A(\g.we_clk [5777]));
Q_ASSIGN U10614 ( .B(clk), .A(\g.we_clk [5776]));
Q_ASSIGN U10615 ( .B(clk), .A(\g.we_clk [5775]));
Q_ASSIGN U10616 ( .B(clk), .A(\g.we_clk [5774]));
Q_ASSIGN U10617 ( .B(clk), .A(\g.we_clk [5773]));
Q_ASSIGN U10618 ( .B(clk), .A(\g.we_clk [5772]));
Q_ASSIGN U10619 ( .B(clk), .A(\g.we_clk [5771]));
Q_ASSIGN U10620 ( .B(clk), .A(\g.we_clk [5770]));
Q_ASSIGN U10621 ( .B(clk), .A(\g.we_clk [5769]));
Q_ASSIGN U10622 ( .B(clk), .A(\g.we_clk [5768]));
Q_ASSIGN U10623 ( .B(clk), .A(\g.we_clk [5767]));
Q_ASSIGN U10624 ( .B(clk), .A(\g.we_clk [5766]));
Q_ASSIGN U10625 ( .B(clk), .A(\g.we_clk [5765]));
Q_ASSIGN U10626 ( .B(clk), .A(\g.we_clk [5764]));
Q_ASSIGN U10627 ( .B(clk), .A(\g.we_clk [5763]));
Q_ASSIGN U10628 ( .B(clk), .A(\g.we_clk [5762]));
Q_ASSIGN U10629 ( .B(clk), .A(\g.we_clk [5761]));
Q_ASSIGN U10630 ( .B(clk), .A(\g.we_clk [5760]));
Q_ASSIGN U10631 ( .B(clk), .A(\g.we_clk [5759]));
Q_ASSIGN U10632 ( .B(clk), .A(\g.we_clk [5758]));
Q_ASSIGN U10633 ( .B(clk), .A(\g.we_clk [5757]));
Q_ASSIGN U10634 ( .B(clk), .A(\g.we_clk [5756]));
Q_ASSIGN U10635 ( .B(clk), .A(\g.we_clk [5755]));
Q_ASSIGN U10636 ( .B(clk), .A(\g.we_clk [5754]));
Q_ASSIGN U10637 ( .B(clk), .A(\g.we_clk [5753]));
Q_ASSIGN U10638 ( .B(clk), .A(\g.we_clk [5752]));
Q_ASSIGN U10639 ( .B(clk), .A(\g.we_clk [5751]));
Q_ASSIGN U10640 ( .B(clk), .A(\g.we_clk [5750]));
Q_ASSIGN U10641 ( .B(clk), .A(\g.we_clk [5749]));
Q_ASSIGN U10642 ( .B(clk), .A(\g.we_clk [5748]));
Q_ASSIGN U10643 ( .B(clk), .A(\g.we_clk [5747]));
Q_ASSIGN U10644 ( .B(clk), .A(\g.we_clk [5746]));
Q_ASSIGN U10645 ( .B(clk), .A(\g.we_clk [5745]));
Q_ASSIGN U10646 ( .B(clk), .A(\g.we_clk [5744]));
Q_ASSIGN U10647 ( .B(clk), .A(\g.we_clk [5743]));
Q_ASSIGN U10648 ( .B(clk), .A(\g.we_clk [5742]));
Q_ASSIGN U10649 ( .B(clk), .A(\g.we_clk [5741]));
Q_ASSIGN U10650 ( .B(clk), .A(\g.we_clk [5740]));
Q_ASSIGN U10651 ( .B(clk), .A(\g.we_clk [5739]));
Q_ASSIGN U10652 ( .B(clk), .A(\g.we_clk [5738]));
Q_ASSIGN U10653 ( .B(clk), .A(\g.we_clk [5737]));
Q_ASSIGN U10654 ( .B(clk), .A(\g.we_clk [5736]));
Q_ASSIGN U10655 ( .B(clk), .A(\g.we_clk [5735]));
Q_ASSIGN U10656 ( .B(clk), .A(\g.we_clk [5734]));
Q_ASSIGN U10657 ( .B(clk), .A(\g.we_clk [5733]));
Q_ASSIGN U10658 ( .B(clk), .A(\g.we_clk [5732]));
Q_ASSIGN U10659 ( .B(clk), .A(\g.we_clk [5731]));
Q_ASSIGN U10660 ( .B(clk), .A(\g.we_clk [5730]));
Q_ASSIGN U10661 ( .B(clk), .A(\g.we_clk [5729]));
Q_ASSIGN U10662 ( .B(clk), .A(\g.we_clk [5728]));
Q_ASSIGN U10663 ( .B(clk), .A(\g.we_clk [5727]));
Q_ASSIGN U10664 ( .B(clk), .A(\g.we_clk [5726]));
Q_ASSIGN U10665 ( .B(clk), .A(\g.we_clk [5725]));
Q_ASSIGN U10666 ( .B(clk), .A(\g.we_clk [5724]));
Q_ASSIGN U10667 ( .B(clk), .A(\g.we_clk [5723]));
Q_ASSIGN U10668 ( .B(clk), .A(\g.we_clk [5722]));
Q_ASSIGN U10669 ( .B(clk), .A(\g.we_clk [5721]));
Q_ASSIGN U10670 ( .B(clk), .A(\g.we_clk [5720]));
Q_ASSIGN U10671 ( .B(clk), .A(\g.we_clk [5719]));
Q_ASSIGN U10672 ( .B(clk), .A(\g.we_clk [5718]));
Q_ASSIGN U10673 ( .B(clk), .A(\g.we_clk [5717]));
Q_ASSIGN U10674 ( .B(clk), .A(\g.we_clk [5716]));
Q_ASSIGN U10675 ( .B(clk), .A(\g.we_clk [5715]));
Q_ASSIGN U10676 ( .B(clk), .A(\g.we_clk [5714]));
Q_ASSIGN U10677 ( .B(clk), .A(\g.we_clk [5713]));
Q_ASSIGN U10678 ( .B(clk), .A(\g.we_clk [5712]));
Q_ASSIGN U10679 ( .B(clk), .A(\g.we_clk [5711]));
Q_ASSIGN U10680 ( .B(clk), .A(\g.we_clk [5710]));
Q_ASSIGN U10681 ( .B(clk), .A(\g.we_clk [5709]));
Q_ASSIGN U10682 ( .B(clk), .A(\g.we_clk [5708]));
Q_ASSIGN U10683 ( .B(clk), .A(\g.we_clk [5707]));
Q_ASSIGN U10684 ( .B(clk), .A(\g.we_clk [5706]));
Q_ASSIGN U10685 ( .B(clk), .A(\g.we_clk [5705]));
Q_ASSIGN U10686 ( .B(clk), .A(\g.we_clk [5704]));
Q_ASSIGN U10687 ( .B(clk), .A(\g.we_clk [5703]));
Q_ASSIGN U10688 ( .B(clk), .A(\g.we_clk [5702]));
Q_ASSIGN U10689 ( .B(clk), .A(\g.we_clk [5701]));
Q_ASSIGN U10690 ( .B(clk), .A(\g.we_clk [5700]));
Q_ASSIGN U10691 ( .B(clk), .A(\g.we_clk [5699]));
Q_ASSIGN U10692 ( .B(clk), .A(\g.we_clk [5698]));
Q_ASSIGN U10693 ( .B(clk), .A(\g.we_clk [5697]));
Q_ASSIGN U10694 ( .B(clk), .A(\g.we_clk [5696]));
Q_ASSIGN U10695 ( .B(clk), .A(\g.we_clk [5695]));
Q_ASSIGN U10696 ( .B(clk), .A(\g.we_clk [5694]));
Q_ASSIGN U10697 ( .B(clk), .A(\g.we_clk [5693]));
Q_ASSIGN U10698 ( .B(clk), .A(\g.we_clk [5692]));
Q_ASSIGN U10699 ( .B(clk), .A(\g.we_clk [5691]));
Q_ASSIGN U10700 ( .B(clk), .A(\g.we_clk [5690]));
Q_ASSIGN U10701 ( .B(clk), .A(\g.we_clk [5689]));
Q_ASSIGN U10702 ( .B(clk), .A(\g.we_clk [5688]));
Q_ASSIGN U10703 ( .B(clk), .A(\g.we_clk [5687]));
Q_ASSIGN U10704 ( .B(clk), .A(\g.we_clk [5686]));
Q_ASSIGN U10705 ( .B(clk), .A(\g.we_clk [5685]));
Q_ASSIGN U10706 ( .B(clk), .A(\g.we_clk [5684]));
Q_ASSIGN U10707 ( .B(clk), .A(\g.we_clk [5683]));
Q_ASSIGN U10708 ( .B(clk), .A(\g.we_clk [5682]));
Q_ASSIGN U10709 ( .B(clk), .A(\g.we_clk [5681]));
Q_ASSIGN U10710 ( .B(clk), .A(\g.we_clk [5680]));
Q_ASSIGN U10711 ( .B(clk), .A(\g.we_clk [5679]));
Q_ASSIGN U10712 ( .B(clk), .A(\g.we_clk [5678]));
Q_ASSIGN U10713 ( .B(clk), .A(\g.we_clk [5677]));
Q_ASSIGN U10714 ( .B(clk), .A(\g.we_clk [5676]));
Q_ASSIGN U10715 ( .B(clk), .A(\g.we_clk [5675]));
Q_ASSIGN U10716 ( .B(clk), .A(\g.we_clk [5674]));
Q_ASSIGN U10717 ( .B(clk), .A(\g.we_clk [5673]));
Q_ASSIGN U10718 ( .B(clk), .A(\g.we_clk [5672]));
Q_ASSIGN U10719 ( .B(clk), .A(\g.we_clk [5671]));
Q_ASSIGN U10720 ( .B(clk), .A(\g.we_clk [5670]));
Q_ASSIGN U10721 ( .B(clk), .A(\g.we_clk [5669]));
Q_ASSIGN U10722 ( .B(clk), .A(\g.we_clk [5668]));
Q_ASSIGN U10723 ( .B(clk), .A(\g.we_clk [5667]));
Q_ASSIGN U10724 ( .B(clk), .A(\g.we_clk [5666]));
Q_ASSIGN U10725 ( .B(clk), .A(\g.we_clk [5665]));
Q_ASSIGN U10726 ( .B(clk), .A(\g.we_clk [5664]));
Q_ASSIGN U10727 ( .B(clk), .A(\g.we_clk [5663]));
Q_ASSIGN U10728 ( .B(clk), .A(\g.we_clk [5662]));
Q_ASSIGN U10729 ( .B(clk), .A(\g.we_clk [5661]));
Q_ASSIGN U10730 ( .B(clk), .A(\g.we_clk [5660]));
Q_ASSIGN U10731 ( .B(clk), .A(\g.we_clk [5659]));
Q_ASSIGN U10732 ( .B(clk), .A(\g.we_clk [5658]));
Q_ASSIGN U10733 ( .B(clk), .A(\g.we_clk [5657]));
Q_ASSIGN U10734 ( .B(clk), .A(\g.we_clk [5656]));
Q_ASSIGN U10735 ( .B(clk), .A(\g.we_clk [5655]));
Q_ASSIGN U10736 ( .B(clk), .A(\g.we_clk [5654]));
Q_ASSIGN U10737 ( .B(clk), .A(\g.we_clk [5653]));
Q_ASSIGN U10738 ( .B(clk), .A(\g.we_clk [5652]));
Q_ASSIGN U10739 ( .B(clk), .A(\g.we_clk [5651]));
Q_ASSIGN U10740 ( .B(clk), .A(\g.we_clk [5650]));
Q_ASSIGN U10741 ( .B(clk), .A(\g.we_clk [5649]));
Q_ASSIGN U10742 ( .B(clk), .A(\g.we_clk [5648]));
Q_ASSIGN U10743 ( .B(clk), .A(\g.we_clk [5647]));
Q_ASSIGN U10744 ( .B(clk), .A(\g.we_clk [5646]));
Q_ASSIGN U10745 ( .B(clk), .A(\g.we_clk [5645]));
Q_ASSIGN U10746 ( .B(clk), .A(\g.we_clk [5644]));
Q_ASSIGN U10747 ( .B(clk), .A(\g.we_clk [5643]));
Q_ASSIGN U10748 ( .B(clk), .A(\g.we_clk [5642]));
Q_ASSIGN U10749 ( .B(clk), .A(\g.we_clk [5641]));
Q_ASSIGN U10750 ( .B(clk), .A(\g.we_clk [5640]));
Q_ASSIGN U10751 ( .B(clk), .A(\g.we_clk [5639]));
Q_ASSIGN U10752 ( .B(clk), .A(\g.we_clk [5638]));
Q_ASSIGN U10753 ( .B(clk), .A(\g.we_clk [5637]));
Q_ASSIGN U10754 ( .B(clk), .A(\g.we_clk [5636]));
Q_ASSIGN U10755 ( .B(clk), .A(\g.we_clk [5635]));
Q_ASSIGN U10756 ( .B(clk), .A(\g.we_clk [5634]));
Q_ASSIGN U10757 ( .B(clk), .A(\g.we_clk [5633]));
Q_ASSIGN U10758 ( .B(clk), .A(\g.we_clk [5632]));
Q_ASSIGN U10759 ( .B(clk), .A(\g.we_clk [5631]));
Q_ASSIGN U10760 ( .B(clk), .A(\g.we_clk [5630]));
Q_ASSIGN U10761 ( .B(clk), .A(\g.we_clk [5629]));
Q_ASSIGN U10762 ( .B(clk), .A(\g.we_clk [5628]));
Q_ASSIGN U10763 ( .B(clk), .A(\g.we_clk [5627]));
Q_ASSIGN U10764 ( .B(clk), .A(\g.we_clk [5626]));
Q_ASSIGN U10765 ( .B(clk), .A(\g.we_clk [5625]));
Q_ASSIGN U10766 ( .B(clk), .A(\g.we_clk [5624]));
Q_ASSIGN U10767 ( .B(clk), .A(\g.we_clk [5623]));
Q_ASSIGN U10768 ( .B(clk), .A(\g.we_clk [5622]));
Q_ASSIGN U10769 ( .B(clk), .A(\g.we_clk [5621]));
Q_ASSIGN U10770 ( .B(clk), .A(\g.we_clk [5620]));
Q_ASSIGN U10771 ( .B(clk), .A(\g.we_clk [5619]));
Q_ASSIGN U10772 ( .B(clk), .A(\g.we_clk [5618]));
Q_ASSIGN U10773 ( .B(clk), .A(\g.we_clk [5617]));
Q_ASSIGN U10774 ( .B(clk), .A(\g.we_clk [5616]));
Q_ASSIGN U10775 ( .B(clk), .A(\g.we_clk [5615]));
Q_ASSIGN U10776 ( .B(clk), .A(\g.we_clk [5614]));
Q_ASSIGN U10777 ( .B(clk), .A(\g.we_clk [5613]));
Q_ASSIGN U10778 ( .B(clk), .A(\g.we_clk [5612]));
Q_ASSIGN U10779 ( .B(clk), .A(\g.we_clk [5611]));
Q_ASSIGN U10780 ( .B(clk), .A(\g.we_clk [5610]));
Q_ASSIGN U10781 ( .B(clk), .A(\g.we_clk [5609]));
Q_ASSIGN U10782 ( .B(clk), .A(\g.we_clk [5608]));
Q_ASSIGN U10783 ( .B(clk), .A(\g.we_clk [5607]));
Q_ASSIGN U10784 ( .B(clk), .A(\g.we_clk [5606]));
Q_ASSIGN U10785 ( .B(clk), .A(\g.we_clk [5605]));
Q_ASSIGN U10786 ( .B(clk), .A(\g.we_clk [5604]));
Q_ASSIGN U10787 ( .B(clk), .A(\g.we_clk [5603]));
Q_ASSIGN U10788 ( .B(clk), .A(\g.we_clk [5602]));
Q_ASSIGN U10789 ( .B(clk), .A(\g.we_clk [5601]));
Q_ASSIGN U10790 ( .B(clk), .A(\g.we_clk [5600]));
Q_ASSIGN U10791 ( .B(clk), .A(\g.we_clk [5599]));
Q_ASSIGN U10792 ( .B(clk), .A(\g.we_clk [5598]));
Q_ASSIGN U10793 ( .B(clk), .A(\g.we_clk [5597]));
Q_ASSIGN U10794 ( .B(clk), .A(\g.we_clk [5596]));
Q_ASSIGN U10795 ( .B(clk), .A(\g.we_clk [5595]));
Q_ASSIGN U10796 ( .B(clk), .A(\g.we_clk [5594]));
Q_ASSIGN U10797 ( .B(clk), .A(\g.we_clk [5593]));
Q_ASSIGN U10798 ( .B(clk), .A(\g.we_clk [5592]));
Q_ASSIGN U10799 ( .B(clk), .A(\g.we_clk [5591]));
Q_ASSIGN U10800 ( .B(clk), .A(\g.we_clk [5590]));
Q_ASSIGN U10801 ( .B(clk), .A(\g.we_clk [5589]));
Q_ASSIGN U10802 ( .B(clk), .A(\g.we_clk [5588]));
Q_ASSIGN U10803 ( .B(clk), .A(\g.we_clk [5587]));
Q_ASSIGN U10804 ( .B(clk), .A(\g.we_clk [5586]));
Q_ASSIGN U10805 ( .B(clk), .A(\g.we_clk [5585]));
Q_ASSIGN U10806 ( .B(clk), .A(\g.we_clk [5584]));
Q_ASSIGN U10807 ( .B(clk), .A(\g.we_clk [5583]));
Q_ASSIGN U10808 ( .B(clk), .A(\g.we_clk [5582]));
Q_ASSIGN U10809 ( .B(clk), .A(\g.we_clk [5581]));
Q_ASSIGN U10810 ( .B(clk), .A(\g.we_clk [5580]));
Q_ASSIGN U10811 ( .B(clk), .A(\g.we_clk [5579]));
Q_ASSIGN U10812 ( .B(clk), .A(\g.we_clk [5578]));
Q_ASSIGN U10813 ( .B(clk), .A(\g.we_clk [5577]));
Q_ASSIGN U10814 ( .B(clk), .A(\g.we_clk [5576]));
Q_ASSIGN U10815 ( .B(clk), .A(\g.we_clk [5575]));
Q_ASSIGN U10816 ( .B(clk), .A(\g.we_clk [5574]));
Q_ASSIGN U10817 ( .B(clk), .A(\g.we_clk [5573]));
Q_ASSIGN U10818 ( .B(clk), .A(\g.we_clk [5572]));
Q_ASSIGN U10819 ( .B(clk), .A(\g.we_clk [5571]));
Q_ASSIGN U10820 ( .B(clk), .A(\g.we_clk [5570]));
Q_ASSIGN U10821 ( .B(clk), .A(\g.we_clk [5569]));
Q_ASSIGN U10822 ( .B(clk), .A(\g.we_clk [5568]));
Q_ASSIGN U10823 ( .B(clk), .A(\g.we_clk [5567]));
Q_ASSIGN U10824 ( .B(clk), .A(\g.we_clk [5566]));
Q_ASSIGN U10825 ( .B(clk), .A(\g.we_clk [5565]));
Q_ASSIGN U10826 ( .B(clk), .A(\g.we_clk [5564]));
Q_ASSIGN U10827 ( .B(clk), .A(\g.we_clk [5563]));
Q_ASSIGN U10828 ( .B(clk), .A(\g.we_clk [5562]));
Q_ASSIGN U10829 ( .B(clk), .A(\g.we_clk [5561]));
Q_ASSIGN U10830 ( .B(clk), .A(\g.we_clk [5560]));
Q_ASSIGN U10831 ( .B(clk), .A(\g.we_clk [5559]));
Q_ASSIGN U10832 ( .B(clk), .A(\g.we_clk [5558]));
Q_ASSIGN U10833 ( .B(clk), .A(\g.we_clk [5557]));
Q_ASSIGN U10834 ( .B(clk), .A(\g.we_clk [5556]));
Q_ASSIGN U10835 ( .B(clk), .A(\g.we_clk [5555]));
Q_ASSIGN U10836 ( .B(clk), .A(\g.we_clk [5554]));
Q_ASSIGN U10837 ( .B(clk), .A(\g.we_clk [5553]));
Q_ASSIGN U10838 ( .B(clk), .A(\g.we_clk [5552]));
Q_ASSIGN U10839 ( .B(clk), .A(\g.we_clk [5551]));
Q_ASSIGN U10840 ( .B(clk), .A(\g.we_clk [5550]));
Q_ASSIGN U10841 ( .B(clk), .A(\g.we_clk [5549]));
Q_ASSIGN U10842 ( .B(clk), .A(\g.we_clk [5548]));
Q_ASSIGN U10843 ( .B(clk), .A(\g.we_clk [5547]));
Q_ASSIGN U10844 ( .B(clk), .A(\g.we_clk [5546]));
Q_ASSIGN U10845 ( .B(clk), .A(\g.we_clk [5545]));
Q_ASSIGN U10846 ( .B(clk), .A(\g.we_clk [5544]));
Q_ASSIGN U10847 ( .B(clk), .A(\g.we_clk [5543]));
Q_ASSIGN U10848 ( .B(clk), .A(\g.we_clk [5542]));
Q_ASSIGN U10849 ( .B(clk), .A(\g.we_clk [5541]));
Q_ASSIGN U10850 ( .B(clk), .A(\g.we_clk [5540]));
Q_ASSIGN U10851 ( .B(clk), .A(\g.we_clk [5539]));
Q_ASSIGN U10852 ( .B(clk), .A(\g.we_clk [5538]));
Q_ASSIGN U10853 ( .B(clk), .A(\g.we_clk [5537]));
Q_ASSIGN U10854 ( .B(clk), .A(\g.we_clk [5536]));
Q_ASSIGN U10855 ( .B(clk), .A(\g.we_clk [5535]));
Q_ASSIGN U10856 ( .B(clk), .A(\g.we_clk [5534]));
Q_ASSIGN U10857 ( .B(clk), .A(\g.we_clk [5533]));
Q_ASSIGN U10858 ( .B(clk), .A(\g.we_clk [5532]));
Q_ASSIGN U10859 ( .B(clk), .A(\g.we_clk [5531]));
Q_ASSIGN U10860 ( .B(clk), .A(\g.we_clk [5530]));
Q_ASSIGN U10861 ( .B(clk), .A(\g.we_clk [5529]));
Q_ASSIGN U10862 ( .B(clk), .A(\g.we_clk [5528]));
Q_ASSIGN U10863 ( .B(clk), .A(\g.we_clk [5527]));
Q_ASSIGN U10864 ( .B(clk), .A(\g.we_clk [5526]));
Q_ASSIGN U10865 ( .B(clk), .A(\g.we_clk [5525]));
Q_ASSIGN U10866 ( .B(clk), .A(\g.we_clk [5524]));
Q_ASSIGN U10867 ( .B(clk), .A(\g.we_clk [5523]));
Q_ASSIGN U10868 ( .B(clk), .A(\g.we_clk [5522]));
Q_ASSIGN U10869 ( .B(clk), .A(\g.we_clk [5521]));
Q_ASSIGN U10870 ( .B(clk), .A(\g.we_clk [5520]));
Q_ASSIGN U10871 ( .B(clk), .A(\g.we_clk [5519]));
Q_ASSIGN U10872 ( .B(clk), .A(\g.we_clk [5518]));
Q_ASSIGN U10873 ( .B(clk), .A(\g.we_clk [5517]));
Q_ASSIGN U10874 ( .B(clk), .A(\g.we_clk [5516]));
Q_ASSIGN U10875 ( .B(clk), .A(\g.we_clk [5515]));
Q_ASSIGN U10876 ( .B(clk), .A(\g.we_clk [5514]));
Q_ASSIGN U10877 ( .B(clk), .A(\g.we_clk [5513]));
Q_ASSIGN U10878 ( .B(clk), .A(\g.we_clk [5512]));
Q_ASSIGN U10879 ( .B(clk), .A(\g.we_clk [5511]));
Q_ASSIGN U10880 ( .B(clk), .A(\g.we_clk [5510]));
Q_ASSIGN U10881 ( .B(clk), .A(\g.we_clk [5509]));
Q_ASSIGN U10882 ( .B(clk), .A(\g.we_clk [5508]));
Q_ASSIGN U10883 ( .B(clk), .A(\g.we_clk [5507]));
Q_ASSIGN U10884 ( .B(clk), .A(\g.we_clk [5506]));
Q_ASSIGN U10885 ( .B(clk), .A(\g.we_clk [5505]));
Q_ASSIGN U10886 ( .B(clk), .A(\g.we_clk [5504]));
Q_ASSIGN U10887 ( .B(clk), .A(\g.we_clk [5503]));
Q_ASSIGN U10888 ( .B(clk), .A(\g.we_clk [5502]));
Q_ASSIGN U10889 ( .B(clk), .A(\g.we_clk [5501]));
Q_ASSIGN U10890 ( .B(clk), .A(\g.we_clk [5500]));
Q_ASSIGN U10891 ( .B(clk), .A(\g.we_clk [5499]));
Q_ASSIGN U10892 ( .B(clk), .A(\g.we_clk [5498]));
Q_ASSIGN U10893 ( .B(clk), .A(\g.we_clk [5497]));
Q_ASSIGN U10894 ( .B(clk), .A(\g.we_clk [5496]));
Q_ASSIGN U10895 ( .B(clk), .A(\g.we_clk [5495]));
Q_ASSIGN U10896 ( .B(clk), .A(\g.we_clk [5494]));
Q_ASSIGN U10897 ( .B(clk), .A(\g.we_clk [5493]));
Q_ASSIGN U10898 ( .B(clk), .A(\g.we_clk [5492]));
Q_ASSIGN U10899 ( .B(clk), .A(\g.we_clk [5491]));
Q_ASSIGN U10900 ( .B(clk), .A(\g.we_clk [5490]));
Q_ASSIGN U10901 ( .B(clk), .A(\g.we_clk [5489]));
Q_ASSIGN U10902 ( .B(clk), .A(\g.we_clk [5488]));
Q_ASSIGN U10903 ( .B(clk), .A(\g.we_clk [5487]));
Q_ASSIGN U10904 ( .B(clk), .A(\g.we_clk [5486]));
Q_ASSIGN U10905 ( .B(clk), .A(\g.we_clk [5485]));
Q_ASSIGN U10906 ( .B(clk), .A(\g.we_clk [5484]));
Q_ASSIGN U10907 ( .B(clk), .A(\g.we_clk [5483]));
Q_ASSIGN U10908 ( .B(clk), .A(\g.we_clk [5482]));
Q_ASSIGN U10909 ( .B(clk), .A(\g.we_clk [5481]));
Q_ASSIGN U10910 ( .B(clk), .A(\g.we_clk [5480]));
Q_ASSIGN U10911 ( .B(clk), .A(\g.we_clk [5479]));
Q_ASSIGN U10912 ( .B(clk), .A(\g.we_clk [5478]));
Q_ASSIGN U10913 ( .B(clk), .A(\g.we_clk [5477]));
Q_ASSIGN U10914 ( .B(clk), .A(\g.we_clk [5476]));
Q_ASSIGN U10915 ( .B(clk), .A(\g.we_clk [5475]));
Q_ASSIGN U10916 ( .B(clk), .A(\g.we_clk [5474]));
Q_ASSIGN U10917 ( .B(clk), .A(\g.we_clk [5473]));
Q_ASSIGN U10918 ( .B(clk), .A(\g.we_clk [5472]));
Q_ASSIGN U10919 ( .B(clk), .A(\g.we_clk [5471]));
Q_ASSIGN U10920 ( .B(clk), .A(\g.we_clk [5470]));
Q_ASSIGN U10921 ( .B(clk), .A(\g.we_clk [5469]));
Q_ASSIGN U10922 ( .B(clk), .A(\g.we_clk [5468]));
Q_ASSIGN U10923 ( .B(clk), .A(\g.we_clk [5467]));
Q_ASSIGN U10924 ( .B(clk), .A(\g.we_clk [5466]));
Q_ASSIGN U10925 ( .B(clk), .A(\g.we_clk [5465]));
Q_ASSIGN U10926 ( .B(clk), .A(\g.we_clk [5464]));
Q_ASSIGN U10927 ( .B(clk), .A(\g.we_clk [5463]));
Q_ASSIGN U10928 ( .B(clk), .A(\g.we_clk [5462]));
Q_ASSIGN U10929 ( .B(clk), .A(\g.we_clk [5461]));
Q_ASSIGN U10930 ( .B(clk), .A(\g.we_clk [5460]));
Q_ASSIGN U10931 ( .B(clk), .A(\g.we_clk [5459]));
Q_ASSIGN U10932 ( .B(clk), .A(\g.we_clk [5458]));
Q_ASSIGN U10933 ( .B(clk), .A(\g.we_clk [5457]));
Q_ASSIGN U10934 ( .B(clk), .A(\g.we_clk [5456]));
Q_ASSIGN U10935 ( .B(clk), .A(\g.we_clk [5455]));
Q_ASSIGN U10936 ( .B(clk), .A(\g.we_clk [5454]));
Q_ASSIGN U10937 ( .B(clk), .A(\g.we_clk [5453]));
Q_ASSIGN U10938 ( .B(clk), .A(\g.we_clk [5452]));
Q_ASSIGN U10939 ( .B(clk), .A(\g.we_clk [5451]));
Q_ASSIGN U10940 ( .B(clk), .A(\g.we_clk [5450]));
Q_ASSIGN U10941 ( .B(clk), .A(\g.we_clk [5449]));
Q_ASSIGN U10942 ( .B(clk), .A(\g.we_clk [5448]));
Q_ASSIGN U10943 ( .B(clk), .A(\g.we_clk [5447]));
Q_ASSIGN U10944 ( .B(clk), .A(\g.we_clk [5446]));
Q_ASSIGN U10945 ( .B(clk), .A(\g.we_clk [5445]));
Q_ASSIGN U10946 ( .B(clk), .A(\g.we_clk [5444]));
Q_ASSIGN U10947 ( .B(clk), .A(\g.we_clk [5443]));
Q_ASSIGN U10948 ( .B(clk), .A(\g.we_clk [5442]));
Q_ASSIGN U10949 ( .B(clk), .A(\g.we_clk [5441]));
Q_ASSIGN U10950 ( .B(clk), .A(\g.we_clk [5440]));
Q_ASSIGN U10951 ( .B(clk), .A(\g.we_clk [5439]));
Q_ASSIGN U10952 ( .B(clk), .A(\g.we_clk [5438]));
Q_ASSIGN U10953 ( .B(clk), .A(\g.we_clk [5437]));
Q_ASSIGN U10954 ( .B(clk), .A(\g.we_clk [5436]));
Q_ASSIGN U10955 ( .B(clk), .A(\g.we_clk [5435]));
Q_ASSIGN U10956 ( .B(clk), .A(\g.we_clk [5434]));
Q_ASSIGN U10957 ( .B(clk), .A(\g.we_clk [5433]));
Q_ASSIGN U10958 ( .B(clk), .A(\g.we_clk [5432]));
Q_ASSIGN U10959 ( .B(clk), .A(\g.we_clk [5431]));
Q_ASSIGN U10960 ( .B(clk), .A(\g.we_clk [5430]));
Q_ASSIGN U10961 ( .B(clk), .A(\g.we_clk [5429]));
Q_ASSIGN U10962 ( .B(clk), .A(\g.we_clk [5428]));
Q_ASSIGN U10963 ( .B(clk), .A(\g.we_clk [5427]));
Q_ASSIGN U10964 ( .B(clk), .A(\g.we_clk [5426]));
Q_ASSIGN U10965 ( .B(clk), .A(\g.we_clk [5425]));
Q_ASSIGN U10966 ( .B(clk), .A(\g.we_clk [5424]));
Q_ASSIGN U10967 ( .B(clk), .A(\g.we_clk [5423]));
Q_ASSIGN U10968 ( .B(clk), .A(\g.we_clk [5422]));
Q_ASSIGN U10969 ( .B(clk), .A(\g.we_clk [5421]));
Q_ASSIGN U10970 ( .B(clk), .A(\g.we_clk [5420]));
Q_ASSIGN U10971 ( .B(clk), .A(\g.we_clk [5419]));
Q_ASSIGN U10972 ( .B(clk), .A(\g.we_clk [5418]));
Q_ASSIGN U10973 ( .B(clk), .A(\g.we_clk [5417]));
Q_ASSIGN U10974 ( .B(clk), .A(\g.we_clk [5416]));
Q_ASSIGN U10975 ( .B(clk), .A(\g.we_clk [5415]));
Q_ASSIGN U10976 ( .B(clk), .A(\g.we_clk [5414]));
Q_ASSIGN U10977 ( .B(clk), .A(\g.we_clk [5413]));
Q_ASSIGN U10978 ( .B(clk), .A(\g.we_clk [5412]));
Q_ASSIGN U10979 ( .B(clk), .A(\g.we_clk [5411]));
Q_ASSIGN U10980 ( .B(clk), .A(\g.we_clk [5410]));
Q_ASSIGN U10981 ( .B(clk), .A(\g.we_clk [5409]));
Q_ASSIGN U10982 ( .B(clk), .A(\g.we_clk [5408]));
Q_ASSIGN U10983 ( .B(clk), .A(\g.we_clk [5407]));
Q_ASSIGN U10984 ( .B(clk), .A(\g.we_clk [5406]));
Q_ASSIGN U10985 ( .B(clk), .A(\g.we_clk [5405]));
Q_ASSIGN U10986 ( .B(clk), .A(\g.we_clk [5404]));
Q_ASSIGN U10987 ( .B(clk), .A(\g.we_clk [5403]));
Q_ASSIGN U10988 ( .B(clk), .A(\g.we_clk [5402]));
Q_ASSIGN U10989 ( .B(clk), .A(\g.we_clk [5401]));
Q_ASSIGN U10990 ( .B(clk), .A(\g.we_clk [5400]));
Q_ASSIGN U10991 ( .B(clk), .A(\g.we_clk [5399]));
Q_ASSIGN U10992 ( .B(clk), .A(\g.we_clk [5398]));
Q_ASSIGN U10993 ( .B(clk), .A(\g.we_clk [5397]));
Q_ASSIGN U10994 ( .B(clk), .A(\g.we_clk [5396]));
Q_ASSIGN U10995 ( .B(clk), .A(\g.we_clk [5395]));
Q_ASSIGN U10996 ( .B(clk), .A(\g.we_clk [5394]));
Q_ASSIGN U10997 ( .B(clk), .A(\g.we_clk [5393]));
Q_ASSIGN U10998 ( .B(clk), .A(\g.we_clk [5392]));
Q_ASSIGN U10999 ( .B(clk), .A(\g.we_clk [5391]));
Q_ASSIGN U11000 ( .B(clk), .A(\g.we_clk [5390]));
Q_ASSIGN U11001 ( .B(clk), .A(\g.we_clk [5389]));
Q_ASSIGN U11002 ( .B(clk), .A(\g.we_clk [5388]));
Q_ASSIGN U11003 ( .B(clk), .A(\g.we_clk [5387]));
Q_ASSIGN U11004 ( .B(clk), .A(\g.we_clk [5386]));
Q_ASSIGN U11005 ( .B(clk), .A(\g.we_clk [5385]));
Q_ASSIGN U11006 ( .B(clk), .A(\g.we_clk [5384]));
Q_ASSIGN U11007 ( .B(clk), .A(\g.we_clk [5383]));
Q_ASSIGN U11008 ( .B(clk), .A(\g.we_clk [5382]));
Q_ASSIGN U11009 ( .B(clk), .A(\g.we_clk [5381]));
Q_ASSIGN U11010 ( .B(clk), .A(\g.we_clk [5380]));
Q_ASSIGN U11011 ( .B(clk), .A(\g.we_clk [5379]));
Q_ASSIGN U11012 ( .B(clk), .A(\g.we_clk [5378]));
Q_ASSIGN U11013 ( .B(clk), .A(\g.we_clk [5377]));
Q_ASSIGN U11014 ( .B(clk), .A(\g.we_clk [5376]));
Q_ASSIGN U11015 ( .B(clk), .A(\g.we_clk [5375]));
Q_ASSIGN U11016 ( .B(clk), .A(\g.we_clk [5374]));
Q_ASSIGN U11017 ( .B(clk), .A(\g.we_clk [5373]));
Q_ASSIGN U11018 ( .B(clk), .A(\g.we_clk [5372]));
Q_ASSIGN U11019 ( .B(clk), .A(\g.we_clk [5371]));
Q_ASSIGN U11020 ( .B(clk), .A(\g.we_clk [5370]));
Q_ASSIGN U11021 ( .B(clk), .A(\g.we_clk [5369]));
Q_ASSIGN U11022 ( .B(clk), .A(\g.we_clk [5368]));
Q_ASSIGN U11023 ( .B(clk), .A(\g.we_clk [5367]));
Q_ASSIGN U11024 ( .B(clk), .A(\g.we_clk [5366]));
Q_ASSIGN U11025 ( .B(clk), .A(\g.we_clk [5365]));
Q_ASSIGN U11026 ( .B(clk), .A(\g.we_clk [5364]));
Q_ASSIGN U11027 ( .B(clk), .A(\g.we_clk [5363]));
Q_ASSIGN U11028 ( .B(clk), .A(\g.we_clk [5362]));
Q_ASSIGN U11029 ( .B(clk), .A(\g.we_clk [5361]));
Q_ASSIGN U11030 ( .B(clk), .A(\g.we_clk [5360]));
Q_ASSIGN U11031 ( .B(clk), .A(\g.we_clk [5359]));
Q_ASSIGN U11032 ( .B(clk), .A(\g.we_clk [5358]));
Q_ASSIGN U11033 ( .B(clk), .A(\g.we_clk [5357]));
Q_ASSIGN U11034 ( .B(clk), .A(\g.we_clk [5356]));
Q_ASSIGN U11035 ( .B(clk), .A(\g.we_clk [5355]));
Q_ASSIGN U11036 ( .B(clk), .A(\g.we_clk [5354]));
Q_ASSIGN U11037 ( .B(clk), .A(\g.we_clk [5353]));
Q_ASSIGN U11038 ( .B(clk), .A(\g.we_clk [5352]));
Q_ASSIGN U11039 ( .B(clk), .A(\g.we_clk [5351]));
Q_ASSIGN U11040 ( .B(clk), .A(\g.we_clk [5350]));
Q_ASSIGN U11041 ( .B(clk), .A(\g.we_clk [5349]));
Q_ASSIGN U11042 ( .B(clk), .A(\g.we_clk [5348]));
Q_ASSIGN U11043 ( .B(clk), .A(\g.we_clk [5347]));
Q_ASSIGN U11044 ( .B(clk), .A(\g.we_clk [5346]));
Q_ASSIGN U11045 ( .B(clk), .A(\g.we_clk [5345]));
Q_ASSIGN U11046 ( .B(clk), .A(\g.we_clk [5344]));
Q_ASSIGN U11047 ( .B(clk), .A(\g.we_clk [5343]));
Q_ASSIGN U11048 ( .B(clk), .A(\g.we_clk [5342]));
Q_ASSIGN U11049 ( .B(clk), .A(\g.we_clk [5341]));
Q_ASSIGN U11050 ( .B(clk), .A(\g.we_clk [5340]));
Q_ASSIGN U11051 ( .B(clk), .A(\g.we_clk [5339]));
Q_ASSIGN U11052 ( .B(clk), .A(\g.we_clk [5338]));
Q_ASSIGN U11053 ( .B(clk), .A(\g.we_clk [5337]));
Q_ASSIGN U11054 ( .B(clk), .A(\g.we_clk [5336]));
Q_ASSIGN U11055 ( .B(clk), .A(\g.we_clk [5335]));
Q_ASSIGN U11056 ( .B(clk), .A(\g.we_clk [5334]));
Q_ASSIGN U11057 ( .B(clk), .A(\g.we_clk [5333]));
Q_ASSIGN U11058 ( .B(clk), .A(\g.we_clk [5332]));
Q_ASSIGN U11059 ( .B(clk), .A(\g.we_clk [5331]));
Q_ASSIGN U11060 ( .B(clk), .A(\g.we_clk [5330]));
Q_ASSIGN U11061 ( .B(clk), .A(\g.we_clk [5329]));
Q_ASSIGN U11062 ( .B(clk), .A(\g.we_clk [5328]));
Q_ASSIGN U11063 ( .B(clk), .A(\g.we_clk [5327]));
Q_ASSIGN U11064 ( .B(clk), .A(\g.we_clk [5326]));
Q_ASSIGN U11065 ( .B(clk), .A(\g.we_clk [5325]));
Q_ASSIGN U11066 ( .B(clk), .A(\g.we_clk [5324]));
Q_ASSIGN U11067 ( .B(clk), .A(\g.we_clk [5323]));
Q_ASSIGN U11068 ( .B(clk), .A(\g.we_clk [5322]));
Q_ASSIGN U11069 ( .B(clk), .A(\g.we_clk [5321]));
Q_ASSIGN U11070 ( .B(clk), .A(\g.we_clk [5320]));
Q_ASSIGN U11071 ( .B(clk), .A(\g.we_clk [5319]));
Q_ASSIGN U11072 ( .B(clk), .A(\g.we_clk [5318]));
Q_ASSIGN U11073 ( .B(clk), .A(\g.we_clk [5317]));
Q_ASSIGN U11074 ( .B(clk), .A(\g.we_clk [5316]));
Q_ASSIGN U11075 ( .B(clk), .A(\g.we_clk [5315]));
Q_ASSIGN U11076 ( .B(clk), .A(\g.we_clk [5314]));
Q_ASSIGN U11077 ( .B(clk), .A(\g.we_clk [5313]));
Q_ASSIGN U11078 ( .B(clk), .A(\g.we_clk [5312]));
Q_ASSIGN U11079 ( .B(clk), .A(\g.we_clk [5311]));
Q_ASSIGN U11080 ( .B(clk), .A(\g.we_clk [5310]));
Q_ASSIGN U11081 ( .B(clk), .A(\g.we_clk [5309]));
Q_ASSIGN U11082 ( .B(clk), .A(\g.we_clk [5308]));
Q_ASSIGN U11083 ( .B(clk), .A(\g.we_clk [5307]));
Q_ASSIGN U11084 ( .B(clk), .A(\g.we_clk [5306]));
Q_ASSIGN U11085 ( .B(clk), .A(\g.we_clk [5305]));
Q_ASSIGN U11086 ( .B(clk), .A(\g.we_clk [5304]));
Q_ASSIGN U11087 ( .B(clk), .A(\g.we_clk [5303]));
Q_ASSIGN U11088 ( .B(clk), .A(\g.we_clk [5302]));
Q_ASSIGN U11089 ( .B(clk), .A(\g.we_clk [5301]));
Q_ASSIGN U11090 ( .B(clk), .A(\g.we_clk [5300]));
Q_ASSIGN U11091 ( .B(clk), .A(\g.we_clk [5299]));
Q_ASSIGN U11092 ( .B(clk), .A(\g.we_clk [5298]));
Q_ASSIGN U11093 ( .B(clk), .A(\g.we_clk [5297]));
Q_ASSIGN U11094 ( .B(clk), .A(\g.we_clk [5296]));
Q_ASSIGN U11095 ( .B(clk), .A(\g.we_clk [5295]));
Q_ASSIGN U11096 ( .B(clk), .A(\g.we_clk [5294]));
Q_ASSIGN U11097 ( .B(clk), .A(\g.we_clk [5293]));
Q_ASSIGN U11098 ( .B(clk), .A(\g.we_clk [5292]));
Q_ASSIGN U11099 ( .B(clk), .A(\g.we_clk [5291]));
Q_ASSIGN U11100 ( .B(clk), .A(\g.we_clk [5290]));
Q_ASSIGN U11101 ( .B(clk), .A(\g.we_clk [5289]));
Q_ASSIGN U11102 ( .B(clk), .A(\g.we_clk [5288]));
Q_ASSIGN U11103 ( .B(clk), .A(\g.we_clk [5287]));
Q_ASSIGN U11104 ( .B(clk), .A(\g.we_clk [5286]));
Q_ASSIGN U11105 ( .B(clk), .A(\g.we_clk [5285]));
Q_ASSIGN U11106 ( .B(clk), .A(\g.we_clk [5284]));
Q_ASSIGN U11107 ( .B(clk), .A(\g.we_clk [5283]));
Q_ASSIGN U11108 ( .B(clk), .A(\g.we_clk [5282]));
Q_ASSIGN U11109 ( .B(clk), .A(\g.we_clk [5281]));
Q_ASSIGN U11110 ( .B(clk), .A(\g.we_clk [5280]));
Q_ASSIGN U11111 ( .B(clk), .A(\g.we_clk [5279]));
Q_ASSIGN U11112 ( .B(clk), .A(\g.we_clk [5278]));
Q_ASSIGN U11113 ( .B(clk), .A(\g.we_clk [5277]));
Q_ASSIGN U11114 ( .B(clk), .A(\g.we_clk [5276]));
Q_ASSIGN U11115 ( .B(clk), .A(\g.we_clk [5275]));
Q_ASSIGN U11116 ( .B(clk), .A(\g.we_clk [5274]));
Q_ASSIGN U11117 ( .B(clk), .A(\g.we_clk [5273]));
Q_ASSIGN U11118 ( .B(clk), .A(\g.we_clk [5272]));
Q_ASSIGN U11119 ( .B(clk), .A(\g.we_clk [5271]));
Q_ASSIGN U11120 ( .B(clk), .A(\g.we_clk [5270]));
Q_ASSIGN U11121 ( .B(clk), .A(\g.we_clk [5269]));
Q_ASSIGN U11122 ( .B(clk), .A(\g.we_clk [5268]));
Q_ASSIGN U11123 ( .B(clk), .A(\g.we_clk [5267]));
Q_ASSIGN U11124 ( .B(clk), .A(\g.we_clk [5266]));
Q_ASSIGN U11125 ( .B(clk), .A(\g.we_clk [5265]));
Q_ASSIGN U11126 ( .B(clk), .A(\g.we_clk [5264]));
Q_ASSIGN U11127 ( .B(clk), .A(\g.we_clk [5263]));
Q_ASSIGN U11128 ( .B(clk), .A(\g.we_clk [5262]));
Q_ASSIGN U11129 ( .B(clk), .A(\g.we_clk [5261]));
Q_ASSIGN U11130 ( .B(clk), .A(\g.we_clk [5260]));
Q_ASSIGN U11131 ( .B(clk), .A(\g.we_clk [5259]));
Q_ASSIGN U11132 ( .B(clk), .A(\g.we_clk [5258]));
Q_ASSIGN U11133 ( .B(clk), .A(\g.we_clk [5257]));
Q_ASSIGN U11134 ( .B(clk), .A(\g.we_clk [5256]));
Q_ASSIGN U11135 ( .B(clk), .A(\g.we_clk [5255]));
Q_ASSIGN U11136 ( .B(clk), .A(\g.we_clk [5254]));
Q_ASSIGN U11137 ( .B(clk), .A(\g.we_clk [5253]));
Q_ASSIGN U11138 ( .B(clk), .A(\g.we_clk [5252]));
Q_ASSIGN U11139 ( .B(clk), .A(\g.we_clk [5251]));
Q_ASSIGN U11140 ( .B(clk), .A(\g.we_clk [5250]));
Q_ASSIGN U11141 ( .B(clk), .A(\g.we_clk [5249]));
Q_ASSIGN U11142 ( .B(clk), .A(\g.we_clk [5248]));
Q_ASSIGN U11143 ( .B(clk), .A(\g.we_clk [5247]));
Q_ASSIGN U11144 ( .B(clk), .A(\g.we_clk [5246]));
Q_ASSIGN U11145 ( .B(clk), .A(\g.we_clk [5245]));
Q_ASSIGN U11146 ( .B(clk), .A(\g.we_clk [5244]));
Q_ASSIGN U11147 ( .B(clk), .A(\g.we_clk [5243]));
Q_ASSIGN U11148 ( .B(clk), .A(\g.we_clk [5242]));
Q_ASSIGN U11149 ( .B(clk), .A(\g.we_clk [5241]));
Q_ASSIGN U11150 ( .B(clk), .A(\g.we_clk [5240]));
Q_ASSIGN U11151 ( .B(clk), .A(\g.we_clk [5239]));
Q_ASSIGN U11152 ( .B(clk), .A(\g.we_clk [5238]));
Q_ASSIGN U11153 ( .B(clk), .A(\g.we_clk [5237]));
Q_ASSIGN U11154 ( .B(clk), .A(\g.we_clk [5236]));
Q_ASSIGN U11155 ( .B(clk), .A(\g.we_clk [5235]));
Q_ASSIGN U11156 ( .B(clk), .A(\g.we_clk [5234]));
Q_ASSIGN U11157 ( .B(clk), .A(\g.we_clk [5233]));
Q_ASSIGN U11158 ( .B(clk), .A(\g.we_clk [5232]));
Q_ASSIGN U11159 ( .B(clk), .A(\g.we_clk [5231]));
Q_ASSIGN U11160 ( .B(clk), .A(\g.we_clk [5230]));
Q_ASSIGN U11161 ( .B(clk), .A(\g.we_clk [5229]));
Q_ASSIGN U11162 ( .B(clk), .A(\g.we_clk [5228]));
Q_ASSIGN U11163 ( .B(clk), .A(\g.we_clk [5227]));
Q_ASSIGN U11164 ( .B(clk), .A(\g.we_clk [5226]));
Q_ASSIGN U11165 ( .B(clk), .A(\g.we_clk [5225]));
Q_ASSIGN U11166 ( .B(clk), .A(\g.we_clk [5224]));
Q_ASSIGN U11167 ( .B(clk), .A(\g.we_clk [5223]));
Q_ASSIGN U11168 ( .B(clk), .A(\g.we_clk [5222]));
Q_ASSIGN U11169 ( .B(clk), .A(\g.we_clk [5221]));
Q_ASSIGN U11170 ( .B(clk), .A(\g.we_clk [5220]));
Q_ASSIGN U11171 ( .B(clk), .A(\g.we_clk [5219]));
Q_ASSIGN U11172 ( .B(clk), .A(\g.we_clk [5218]));
Q_ASSIGN U11173 ( .B(clk), .A(\g.we_clk [5217]));
Q_ASSIGN U11174 ( .B(clk), .A(\g.we_clk [5216]));
Q_ASSIGN U11175 ( .B(clk), .A(\g.we_clk [5215]));
Q_ASSIGN U11176 ( .B(clk), .A(\g.we_clk [5214]));
Q_ASSIGN U11177 ( .B(clk), .A(\g.we_clk [5213]));
Q_ASSIGN U11178 ( .B(clk), .A(\g.we_clk [5212]));
Q_ASSIGN U11179 ( .B(clk), .A(\g.we_clk [5211]));
Q_ASSIGN U11180 ( .B(clk), .A(\g.we_clk [5210]));
Q_ASSIGN U11181 ( .B(clk), .A(\g.we_clk [5209]));
Q_ASSIGN U11182 ( .B(clk), .A(\g.we_clk [5208]));
Q_ASSIGN U11183 ( .B(clk), .A(\g.we_clk [5207]));
Q_ASSIGN U11184 ( .B(clk), .A(\g.we_clk [5206]));
Q_ASSIGN U11185 ( .B(clk), .A(\g.we_clk [5205]));
Q_ASSIGN U11186 ( .B(clk), .A(\g.we_clk [5204]));
Q_ASSIGN U11187 ( .B(clk), .A(\g.we_clk [5203]));
Q_ASSIGN U11188 ( .B(clk), .A(\g.we_clk [5202]));
Q_ASSIGN U11189 ( .B(clk), .A(\g.we_clk [5201]));
Q_ASSIGN U11190 ( .B(clk), .A(\g.we_clk [5200]));
Q_ASSIGN U11191 ( .B(clk), .A(\g.we_clk [5199]));
Q_ASSIGN U11192 ( .B(clk), .A(\g.we_clk [5198]));
Q_ASSIGN U11193 ( .B(clk), .A(\g.we_clk [5197]));
Q_ASSIGN U11194 ( .B(clk), .A(\g.we_clk [5196]));
Q_ASSIGN U11195 ( .B(clk), .A(\g.we_clk [5195]));
Q_ASSIGN U11196 ( .B(clk), .A(\g.we_clk [5194]));
Q_ASSIGN U11197 ( .B(clk), .A(\g.we_clk [5193]));
Q_ASSIGN U11198 ( .B(clk), .A(\g.we_clk [5192]));
Q_ASSIGN U11199 ( .B(clk), .A(\g.we_clk [5191]));
Q_ASSIGN U11200 ( .B(clk), .A(\g.we_clk [5190]));
Q_ASSIGN U11201 ( .B(clk), .A(\g.we_clk [5189]));
Q_ASSIGN U11202 ( .B(clk), .A(\g.we_clk [5188]));
Q_ASSIGN U11203 ( .B(clk), .A(\g.we_clk [5187]));
Q_ASSIGN U11204 ( .B(clk), .A(\g.we_clk [5186]));
Q_ASSIGN U11205 ( .B(clk), .A(\g.we_clk [5185]));
Q_ASSIGN U11206 ( .B(clk), .A(\g.we_clk [5184]));
Q_ASSIGN U11207 ( .B(clk), .A(\g.we_clk [5183]));
Q_ASSIGN U11208 ( .B(clk), .A(\g.we_clk [5182]));
Q_ASSIGN U11209 ( .B(clk), .A(\g.we_clk [5181]));
Q_ASSIGN U11210 ( .B(clk), .A(\g.we_clk [5180]));
Q_ASSIGN U11211 ( .B(clk), .A(\g.we_clk [5179]));
Q_ASSIGN U11212 ( .B(clk), .A(\g.we_clk [5178]));
Q_ASSIGN U11213 ( .B(clk), .A(\g.we_clk [5177]));
Q_ASSIGN U11214 ( .B(clk), .A(\g.we_clk [5176]));
Q_ASSIGN U11215 ( .B(clk), .A(\g.we_clk [5175]));
Q_ASSIGN U11216 ( .B(clk), .A(\g.we_clk [5174]));
Q_ASSIGN U11217 ( .B(clk), .A(\g.we_clk [5173]));
Q_ASSIGN U11218 ( .B(clk), .A(\g.we_clk [5172]));
Q_ASSIGN U11219 ( .B(clk), .A(\g.we_clk [5171]));
Q_ASSIGN U11220 ( .B(clk), .A(\g.we_clk [5170]));
Q_ASSIGN U11221 ( .B(clk), .A(\g.we_clk [5169]));
Q_ASSIGN U11222 ( .B(clk), .A(\g.we_clk [5168]));
Q_ASSIGN U11223 ( .B(clk), .A(\g.we_clk [5167]));
Q_ASSIGN U11224 ( .B(clk), .A(\g.we_clk [5166]));
Q_ASSIGN U11225 ( .B(clk), .A(\g.we_clk [5165]));
Q_ASSIGN U11226 ( .B(clk), .A(\g.we_clk [5164]));
Q_ASSIGN U11227 ( .B(clk), .A(\g.we_clk [5163]));
Q_ASSIGN U11228 ( .B(clk), .A(\g.we_clk [5162]));
Q_ASSIGN U11229 ( .B(clk), .A(\g.we_clk [5161]));
Q_ASSIGN U11230 ( .B(clk), .A(\g.we_clk [5160]));
Q_ASSIGN U11231 ( .B(clk), .A(\g.we_clk [5159]));
Q_ASSIGN U11232 ( .B(clk), .A(\g.we_clk [5158]));
Q_ASSIGN U11233 ( .B(clk), .A(\g.we_clk [5157]));
Q_ASSIGN U11234 ( .B(clk), .A(\g.we_clk [5156]));
Q_ASSIGN U11235 ( .B(clk), .A(\g.we_clk [5155]));
Q_ASSIGN U11236 ( .B(clk), .A(\g.we_clk [5154]));
Q_ASSIGN U11237 ( .B(clk), .A(\g.we_clk [5153]));
Q_ASSIGN U11238 ( .B(clk), .A(\g.we_clk [5152]));
Q_ASSIGN U11239 ( .B(clk), .A(\g.we_clk [5151]));
Q_ASSIGN U11240 ( .B(clk), .A(\g.we_clk [5150]));
Q_ASSIGN U11241 ( .B(clk), .A(\g.we_clk [5149]));
Q_ASSIGN U11242 ( .B(clk), .A(\g.we_clk [5148]));
Q_ASSIGN U11243 ( .B(clk), .A(\g.we_clk [5147]));
Q_ASSIGN U11244 ( .B(clk), .A(\g.we_clk [5146]));
Q_ASSIGN U11245 ( .B(clk), .A(\g.we_clk [5145]));
Q_ASSIGN U11246 ( .B(clk), .A(\g.we_clk [5144]));
Q_ASSIGN U11247 ( .B(clk), .A(\g.we_clk [5143]));
Q_ASSIGN U11248 ( .B(clk), .A(\g.we_clk [5142]));
Q_ASSIGN U11249 ( .B(clk), .A(\g.we_clk [5141]));
Q_ASSIGN U11250 ( .B(clk), .A(\g.we_clk [5140]));
Q_ASSIGN U11251 ( .B(clk), .A(\g.we_clk [5139]));
Q_ASSIGN U11252 ( .B(clk), .A(\g.we_clk [5138]));
Q_ASSIGN U11253 ( .B(clk), .A(\g.we_clk [5137]));
Q_ASSIGN U11254 ( .B(clk), .A(\g.we_clk [5136]));
Q_ASSIGN U11255 ( .B(clk), .A(\g.we_clk [5135]));
Q_ASSIGN U11256 ( .B(clk), .A(\g.we_clk [5134]));
Q_ASSIGN U11257 ( .B(clk), .A(\g.we_clk [5133]));
Q_ASSIGN U11258 ( .B(clk), .A(\g.we_clk [5132]));
Q_ASSIGN U11259 ( .B(clk), .A(\g.we_clk [5131]));
Q_ASSIGN U11260 ( .B(clk), .A(\g.we_clk [5130]));
Q_ASSIGN U11261 ( .B(clk), .A(\g.we_clk [5129]));
Q_ASSIGN U11262 ( .B(clk), .A(\g.we_clk [5128]));
Q_ASSIGN U11263 ( .B(clk), .A(\g.we_clk [5127]));
Q_ASSIGN U11264 ( .B(clk), .A(\g.we_clk [5126]));
Q_ASSIGN U11265 ( .B(clk), .A(\g.we_clk [5125]));
Q_ASSIGN U11266 ( .B(clk), .A(\g.we_clk [5124]));
Q_ASSIGN U11267 ( .B(clk), .A(\g.we_clk [5123]));
Q_ASSIGN U11268 ( .B(clk), .A(\g.we_clk [5122]));
Q_ASSIGN U11269 ( .B(clk), .A(\g.we_clk [5121]));
Q_ASSIGN U11270 ( .B(clk), .A(\g.we_clk [5120]));
Q_ASSIGN U11271 ( .B(clk), .A(\g.we_clk [5119]));
Q_ASSIGN U11272 ( .B(clk), .A(\g.we_clk [5118]));
Q_ASSIGN U11273 ( .B(clk), .A(\g.we_clk [5117]));
Q_ASSIGN U11274 ( .B(clk), .A(\g.we_clk [5116]));
Q_ASSIGN U11275 ( .B(clk), .A(\g.we_clk [5115]));
Q_ASSIGN U11276 ( .B(clk), .A(\g.we_clk [5114]));
Q_ASSIGN U11277 ( .B(clk), .A(\g.we_clk [5113]));
Q_ASSIGN U11278 ( .B(clk), .A(\g.we_clk [5112]));
Q_ASSIGN U11279 ( .B(clk), .A(\g.we_clk [5111]));
Q_ASSIGN U11280 ( .B(clk), .A(\g.we_clk [5110]));
Q_ASSIGN U11281 ( .B(clk), .A(\g.we_clk [5109]));
Q_ASSIGN U11282 ( .B(clk), .A(\g.we_clk [5108]));
Q_ASSIGN U11283 ( .B(clk), .A(\g.we_clk [5107]));
Q_ASSIGN U11284 ( .B(clk), .A(\g.we_clk [5106]));
Q_ASSIGN U11285 ( .B(clk), .A(\g.we_clk [5105]));
Q_ASSIGN U11286 ( .B(clk), .A(\g.we_clk [5104]));
Q_ASSIGN U11287 ( .B(clk), .A(\g.we_clk [5103]));
Q_ASSIGN U11288 ( .B(clk), .A(\g.we_clk [5102]));
Q_ASSIGN U11289 ( .B(clk), .A(\g.we_clk [5101]));
Q_ASSIGN U11290 ( .B(clk), .A(\g.we_clk [5100]));
Q_ASSIGN U11291 ( .B(clk), .A(\g.we_clk [5099]));
Q_ASSIGN U11292 ( .B(clk), .A(\g.we_clk [5098]));
Q_ASSIGN U11293 ( .B(clk), .A(\g.we_clk [5097]));
Q_ASSIGN U11294 ( .B(clk), .A(\g.we_clk [5096]));
Q_ASSIGN U11295 ( .B(clk), .A(\g.we_clk [5095]));
Q_ASSIGN U11296 ( .B(clk), .A(\g.we_clk [5094]));
Q_ASSIGN U11297 ( .B(clk), .A(\g.we_clk [5093]));
Q_ASSIGN U11298 ( .B(clk), .A(\g.we_clk [5092]));
Q_ASSIGN U11299 ( .B(clk), .A(\g.we_clk [5091]));
Q_ASSIGN U11300 ( .B(clk), .A(\g.we_clk [5090]));
Q_ASSIGN U11301 ( .B(clk), .A(\g.we_clk [5089]));
Q_ASSIGN U11302 ( .B(clk), .A(\g.we_clk [5088]));
Q_ASSIGN U11303 ( .B(clk), .A(\g.we_clk [5087]));
Q_ASSIGN U11304 ( .B(clk), .A(\g.we_clk [5086]));
Q_ASSIGN U11305 ( .B(clk), .A(\g.we_clk [5085]));
Q_ASSIGN U11306 ( .B(clk), .A(\g.we_clk [5084]));
Q_ASSIGN U11307 ( .B(clk), .A(\g.we_clk [5083]));
Q_ASSIGN U11308 ( .B(clk), .A(\g.we_clk [5082]));
Q_ASSIGN U11309 ( .B(clk), .A(\g.we_clk [5081]));
Q_ASSIGN U11310 ( .B(clk), .A(\g.we_clk [5080]));
Q_ASSIGN U11311 ( .B(clk), .A(\g.we_clk [5079]));
Q_ASSIGN U11312 ( .B(clk), .A(\g.we_clk [5078]));
Q_ASSIGN U11313 ( .B(clk), .A(\g.we_clk [5077]));
Q_ASSIGN U11314 ( .B(clk), .A(\g.we_clk [5076]));
Q_ASSIGN U11315 ( .B(clk), .A(\g.we_clk [5075]));
Q_ASSIGN U11316 ( .B(clk), .A(\g.we_clk [5074]));
Q_ASSIGN U11317 ( .B(clk), .A(\g.we_clk [5073]));
Q_ASSIGN U11318 ( .B(clk), .A(\g.we_clk [5072]));
Q_ASSIGN U11319 ( .B(clk), .A(\g.we_clk [5071]));
Q_ASSIGN U11320 ( .B(clk), .A(\g.we_clk [5070]));
Q_ASSIGN U11321 ( .B(clk), .A(\g.we_clk [5069]));
Q_ASSIGN U11322 ( .B(clk), .A(\g.we_clk [5068]));
Q_ASSIGN U11323 ( .B(clk), .A(\g.we_clk [5067]));
Q_ASSIGN U11324 ( .B(clk), .A(\g.we_clk [5066]));
Q_ASSIGN U11325 ( .B(clk), .A(\g.we_clk [5065]));
Q_ASSIGN U11326 ( .B(clk), .A(\g.we_clk [5064]));
Q_ASSIGN U11327 ( .B(clk), .A(\g.we_clk [5063]));
Q_ASSIGN U11328 ( .B(clk), .A(\g.we_clk [5062]));
Q_ASSIGN U11329 ( .B(clk), .A(\g.we_clk [5061]));
Q_ASSIGN U11330 ( .B(clk), .A(\g.we_clk [5060]));
Q_ASSIGN U11331 ( .B(clk), .A(\g.we_clk [5059]));
Q_ASSIGN U11332 ( .B(clk), .A(\g.we_clk [5058]));
Q_ASSIGN U11333 ( .B(clk), .A(\g.we_clk [5057]));
Q_ASSIGN U11334 ( .B(clk), .A(\g.we_clk [5056]));
Q_ASSIGN U11335 ( .B(clk), .A(\g.we_clk [5055]));
Q_ASSIGN U11336 ( .B(clk), .A(\g.we_clk [5054]));
Q_ASSIGN U11337 ( .B(clk), .A(\g.we_clk [5053]));
Q_ASSIGN U11338 ( .B(clk), .A(\g.we_clk [5052]));
Q_ASSIGN U11339 ( .B(clk), .A(\g.we_clk [5051]));
Q_ASSIGN U11340 ( .B(clk), .A(\g.we_clk [5050]));
Q_ASSIGN U11341 ( .B(clk), .A(\g.we_clk [5049]));
Q_ASSIGN U11342 ( .B(clk), .A(\g.we_clk [5048]));
Q_ASSIGN U11343 ( .B(clk), .A(\g.we_clk [5047]));
Q_ASSIGN U11344 ( .B(clk), .A(\g.we_clk [5046]));
Q_ASSIGN U11345 ( .B(clk), .A(\g.we_clk [5045]));
Q_ASSIGN U11346 ( .B(clk), .A(\g.we_clk [5044]));
Q_ASSIGN U11347 ( .B(clk), .A(\g.we_clk [5043]));
Q_ASSIGN U11348 ( .B(clk), .A(\g.we_clk [5042]));
Q_ASSIGN U11349 ( .B(clk), .A(\g.we_clk [5041]));
Q_ASSIGN U11350 ( .B(clk), .A(\g.we_clk [5040]));
Q_ASSIGN U11351 ( .B(clk), .A(\g.we_clk [5039]));
Q_ASSIGN U11352 ( .B(clk), .A(\g.we_clk [5038]));
Q_ASSIGN U11353 ( .B(clk), .A(\g.we_clk [5037]));
Q_ASSIGN U11354 ( .B(clk), .A(\g.we_clk [5036]));
Q_ASSIGN U11355 ( .B(clk), .A(\g.we_clk [5035]));
Q_ASSIGN U11356 ( .B(clk), .A(\g.we_clk [5034]));
Q_ASSIGN U11357 ( .B(clk), .A(\g.we_clk [5033]));
Q_ASSIGN U11358 ( .B(clk), .A(\g.we_clk [5032]));
Q_ASSIGN U11359 ( .B(clk), .A(\g.we_clk [5031]));
Q_ASSIGN U11360 ( .B(clk), .A(\g.we_clk [5030]));
Q_ASSIGN U11361 ( .B(clk), .A(\g.we_clk [5029]));
Q_ASSIGN U11362 ( .B(clk), .A(\g.we_clk [5028]));
Q_ASSIGN U11363 ( .B(clk), .A(\g.we_clk [5027]));
Q_ASSIGN U11364 ( .B(clk), .A(\g.we_clk [5026]));
Q_ASSIGN U11365 ( .B(clk), .A(\g.we_clk [5025]));
Q_ASSIGN U11366 ( .B(clk), .A(\g.we_clk [5024]));
Q_ASSIGN U11367 ( .B(clk), .A(\g.we_clk [5023]));
Q_ASSIGN U11368 ( .B(clk), .A(\g.we_clk [5022]));
Q_ASSIGN U11369 ( .B(clk), .A(\g.we_clk [5021]));
Q_ASSIGN U11370 ( .B(clk), .A(\g.we_clk [5020]));
Q_ASSIGN U11371 ( .B(clk), .A(\g.we_clk [5019]));
Q_ASSIGN U11372 ( .B(clk), .A(\g.we_clk [5018]));
Q_ASSIGN U11373 ( .B(clk), .A(\g.we_clk [5017]));
Q_ASSIGN U11374 ( .B(clk), .A(\g.we_clk [5016]));
Q_ASSIGN U11375 ( .B(clk), .A(\g.we_clk [5015]));
Q_ASSIGN U11376 ( .B(clk), .A(\g.we_clk [5014]));
Q_ASSIGN U11377 ( .B(clk), .A(\g.we_clk [5013]));
Q_ASSIGN U11378 ( .B(clk), .A(\g.we_clk [5012]));
Q_ASSIGN U11379 ( .B(clk), .A(\g.we_clk [5011]));
Q_ASSIGN U11380 ( .B(clk), .A(\g.we_clk [5010]));
Q_ASSIGN U11381 ( .B(clk), .A(\g.we_clk [5009]));
Q_ASSIGN U11382 ( .B(clk), .A(\g.we_clk [5008]));
Q_ASSIGN U11383 ( .B(clk), .A(\g.we_clk [5007]));
Q_ASSIGN U11384 ( .B(clk), .A(\g.we_clk [5006]));
Q_ASSIGN U11385 ( .B(clk), .A(\g.we_clk [5005]));
Q_ASSIGN U11386 ( .B(clk), .A(\g.we_clk [5004]));
Q_ASSIGN U11387 ( .B(clk), .A(\g.we_clk [5003]));
Q_ASSIGN U11388 ( .B(clk), .A(\g.we_clk [5002]));
Q_ASSIGN U11389 ( .B(clk), .A(\g.we_clk [5001]));
Q_ASSIGN U11390 ( .B(clk), .A(\g.we_clk [5000]));
Q_ASSIGN U11391 ( .B(clk), .A(\g.we_clk [4999]));
Q_ASSIGN U11392 ( .B(clk), .A(\g.we_clk [4998]));
Q_ASSIGN U11393 ( .B(clk), .A(\g.we_clk [4997]));
Q_ASSIGN U11394 ( .B(clk), .A(\g.we_clk [4996]));
Q_ASSIGN U11395 ( .B(clk), .A(\g.we_clk [4995]));
Q_ASSIGN U11396 ( .B(clk), .A(\g.we_clk [4994]));
Q_ASSIGN U11397 ( .B(clk), .A(\g.we_clk [4993]));
Q_ASSIGN U11398 ( .B(clk), .A(\g.we_clk [4992]));
Q_ASSIGN U11399 ( .B(clk), .A(\g.we_clk [4991]));
Q_ASSIGN U11400 ( .B(clk), .A(\g.we_clk [4990]));
Q_ASSIGN U11401 ( .B(clk), .A(\g.we_clk [4989]));
Q_ASSIGN U11402 ( .B(clk), .A(\g.we_clk [4988]));
Q_ASSIGN U11403 ( .B(clk), .A(\g.we_clk [4987]));
Q_ASSIGN U11404 ( .B(clk), .A(\g.we_clk [4986]));
Q_ASSIGN U11405 ( .B(clk), .A(\g.we_clk [4985]));
Q_ASSIGN U11406 ( .B(clk), .A(\g.we_clk [4984]));
Q_ASSIGN U11407 ( .B(clk), .A(\g.we_clk [4983]));
Q_ASSIGN U11408 ( .B(clk), .A(\g.we_clk [4982]));
Q_ASSIGN U11409 ( .B(clk), .A(\g.we_clk [4981]));
Q_ASSIGN U11410 ( .B(clk), .A(\g.we_clk [4980]));
Q_ASSIGN U11411 ( .B(clk), .A(\g.we_clk [4979]));
Q_ASSIGN U11412 ( .B(clk), .A(\g.we_clk [4978]));
Q_ASSIGN U11413 ( .B(clk), .A(\g.we_clk [4977]));
Q_ASSIGN U11414 ( .B(clk), .A(\g.we_clk [4976]));
Q_ASSIGN U11415 ( .B(clk), .A(\g.we_clk [4975]));
Q_ASSIGN U11416 ( .B(clk), .A(\g.we_clk [4974]));
Q_ASSIGN U11417 ( .B(clk), .A(\g.we_clk [4973]));
Q_ASSIGN U11418 ( .B(clk), .A(\g.we_clk [4972]));
Q_ASSIGN U11419 ( .B(clk), .A(\g.we_clk [4971]));
Q_ASSIGN U11420 ( .B(clk), .A(\g.we_clk [4970]));
Q_ASSIGN U11421 ( .B(clk), .A(\g.we_clk [4969]));
Q_ASSIGN U11422 ( .B(clk), .A(\g.we_clk [4968]));
Q_ASSIGN U11423 ( .B(clk), .A(\g.we_clk [4967]));
Q_ASSIGN U11424 ( .B(clk), .A(\g.we_clk [4966]));
Q_ASSIGN U11425 ( .B(clk), .A(\g.we_clk [4965]));
Q_ASSIGN U11426 ( .B(clk), .A(\g.we_clk [4964]));
Q_ASSIGN U11427 ( .B(clk), .A(\g.we_clk [4963]));
Q_ASSIGN U11428 ( .B(clk), .A(\g.we_clk [4962]));
Q_ASSIGN U11429 ( .B(clk), .A(\g.we_clk [4961]));
Q_ASSIGN U11430 ( .B(clk), .A(\g.we_clk [4960]));
Q_ASSIGN U11431 ( .B(clk), .A(\g.we_clk [4959]));
Q_ASSIGN U11432 ( .B(clk), .A(\g.we_clk [4958]));
Q_ASSIGN U11433 ( .B(clk), .A(\g.we_clk [4957]));
Q_ASSIGN U11434 ( .B(clk), .A(\g.we_clk [4956]));
Q_ASSIGN U11435 ( .B(clk), .A(\g.we_clk [4955]));
Q_ASSIGN U11436 ( .B(clk), .A(\g.we_clk [4954]));
Q_ASSIGN U11437 ( .B(clk), .A(\g.we_clk [4953]));
Q_ASSIGN U11438 ( .B(clk), .A(\g.we_clk [4952]));
Q_ASSIGN U11439 ( .B(clk), .A(\g.we_clk [4951]));
Q_ASSIGN U11440 ( .B(clk), .A(\g.we_clk [4950]));
Q_ASSIGN U11441 ( .B(clk), .A(\g.we_clk [4949]));
Q_ASSIGN U11442 ( .B(clk), .A(\g.we_clk [4948]));
Q_ASSIGN U11443 ( .B(clk), .A(\g.we_clk [4947]));
Q_ASSIGN U11444 ( .B(clk), .A(\g.we_clk [4946]));
Q_ASSIGN U11445 ( .B(clk), .A(\g.we_clk [4945]));
Q_ASSIGN U11446 ( .B(clk), .A(\g.we_clk [4944]));
Q_ASSIGN U11447 ( .B(clk), .A(\g.we_clk [4943]));
Q_ASSIGN U11448 ( .B(clk), .A(\g.we_clk [4942]));
Q_ASSIGN U11449 ( .B(clk), .A(\g.we_clk [4941]));
Q_ASSIGN U11450 ( .B(clk), .A(\g.we_clk [4940]));
Q_ASSIGN U11451 ( .B(clk), .A(\g.we_clk [4939]));
Q_ASSIGN U11452 ( .B(clk), .A(\g.we_clk [4938]));
Q_ASSIGN U11453 ( .B(clk), .A(\g.we_clk [4937]));
Q_ASSIGN U11454 ( .B(clk), .A(\g.we_clk [4936]));
Q_ASSIGN U11455 ( .B(clk), .A(\g.we_clk [4935]));
Q_ASSIGN U11456 ( .B(clk), .A(\g.we_clk [4934]));
Q_ASSIGN U11457 ( .B(clk), .A(\g.we_clk [4933]));
Q_ASSIGN U11458 ( .B(clk), .A(\g.we_clk [4932]));
Q_ASSIGN U11459 ( .B(clk), .A(\g.we_clk [4931]));
Q_ASSIGN U11460 ( .B(clk), .A(\g.we_clk [4930]));
Q_ASSIGN U11461 ( .B(clk), .A(\g.we_clk [4929]));
Q_ASSIGN U11462 ( .B(clk), .A(\g.we_clk [4928]));
Q_ASSIGN U11463 ( .B(clk), .A(\g.we_clk [4927]));
Q_ASSIGN U11464 ( .B(clk), .A(\g.we_clk [4926]));
Q_ASSIGN U11465 ( .B(clk), .A(\g.we_clk [4925]));
Q_ASSIGN U11466 ( .B(clk), .A(\g.we_clk [4924]));
Q_ASSIGN U11467 ( .B(clk), .A(\g.we_clk [4923]));
Q_ASSIGN U11468 ( .B(clk), .A(\g.we_clk [4922]));
Q_ASSIGN U11469 ( .B(clk), .A(\g.we_clk [4921]));
Q_ASSIGN U11470 ( .B(clk), .A(\g.we_clk [4920]));
Q_ASSIGN U11471 ( .B(clk), .A(\g.we_clk [4919]));
Q_ASSIGN U11472 ( .B(clk), .A(\g.we_clk [4918]));
Q_ASSIGN U11473 ( .B(clk), .A(\g.we_clk [4917]));
Q_ASSIGN U11474 ( .B(clk), .A(\g.we_clk [4916]));
Q_ASSIGN U11475 ( .B(clk), .A(\g.we_clk [4915]));
Q_ASSIGN U11476 ( .B(clk), .A(\g.we_clk [4914]));
Q_ASSIGN U11477 ( .B(clk), .A(\g.we_clk [4913]));
Q_ASSIGN U11478 ( .B(clk), .A(\g.we_clk [4912]));
Q_ASSIGN U11479 ( .B(clk), .A(\g.we_clk [4911]));
Q_ASSIGN U11480 ( .B(clk), .A(\g.we_clk [4910]));
Q_ASSIGN U11481 ( .B(clk), .A(\g.we_clk [4909]));
Q_ASSIGN U11482 ( .B(clk), .A(\g.we_clk [4908]));
Q_ASSIGN U11483 ( .B(clk), .A(\g.we_clk [4907]));
Q_ASSIGN U11484 ( .B(clk), .A(\g.we_clk [4906]));
Q_ASSIGN U11485 ( .B(clk), .A(\g.we_clk [4905]));
Q_ASSIGN U11486 ( .B(clk), .A(\g.we_clk [4904]));
Q_ASSIGN U11487 ( .B(clk), .A(\g.we_clk [4903]));
Q_ASSIGN U11488 ( .B(clk), .A(\g.we_clk [4902]));
Q_ASSIGN U11489 ( .B(clk), .A(\g.we_clk [4901]));
Q_ASSIGN U11490 ( .B(clk), .A(\g.we_clk [4900]));
Q_ASSIGN U11491 ( .B(clk), .A(\g.we_clk [4899]));
Q_ASSIGN U11492 ( .B(clk), .A(\g.we_clk [4898]));
Q_ASSIGN U11493 ( .B(clk), .A(\g.we_clk [4897]));
Q_ASSIGN U11494 ( .B(clk), .A(\g.we_clk [4896]));
Q_ASSIGN U11495 ( .B(clk), .A(\g.we_clk [4895]));
Q_ASSIGN U11496 ( .B(clk), .A(\g.we_clk [4894]));
Q_ASSIGN U11497 ( .B(clk), .A(\g.we_clk [4893]));
Q_ASSIGN U11498 ( .B(clk), .A(\g.we_clk [4892]));
Q_ASSIGN U11499 ( .B(clk), .A(\g.we_clk [4891]));
Q_ASSIGN U11500 ( .B(clk), .A(\g.we_clk [4890]));
Q_ASSIGN U11501 ( .B(clk), .A(\g.we_clk [4889]));
Q_ASSIGN U11502 ( .B(clk), .A(\g.we_clk [4888]));
Q_ASSIGN U11503 ( .B(clk), .A(\g.we_clk [4887]));
Q_ASSIGN U11504 ( .B(clk), .A(\g.we_clk [4886]));
Q_ASSIGN U11505 ( .B(clk), .A(\g.we_clk [4885]));
Q_ASSIGN U11506 ( .B(clk), .A(\g.we_clk [4884]));
Q_ASSIGN U11507 ( .B(clk), .A(\g.we_clk [4883]));
Q_ASSIGN U11508 ( .B(clk), .A(\g.we_clk [4882]));
Q_ASSIGN U11509 ( .B(clk), .A(\g.we_clk [4881]));
Q_ASSIGN U11510 ( .B(clk), .A(\g.we_clk [4880]));
Q_ASSIGN U11511 ( .B(clk), .A(\g.we_clk [4879]));
Q_ASSIGN U11512 ( .B(clk), .A(\g.we_clk [4878]));
Q_ASSIGN U11513 ( .B(clk), .A(\g.we_clk [4877]));
Q_ASSIGN U11514 ( .B(clk), .A(\g.we_clk [4876]));
Q_ASSIGN U11515 ( .B(clk), .A(\g.we_clk [4875]));
Q_ASSIGN U11516 ( .B(clk), .A(\g.we_clk [4874]));
Q_ASSIGN U11517 ( .B(clk), .A(\g.we_clk [4873]));
Q_ASSIGN U11518 ( .B(clk), .A(\g.we_clk [4872]));
Q_ASSIGN U11519 ( .B(clk), .A(\g.we_clk [4871]));
Q_ASSIGN U11520 ( .B(clk), .A(\g.we_clk [4870]));
Q_ASSIGN U11521 ( .B(clk), .A(\g.we_clk [4869]));
Q_ASSIGN U11522 ( .B(clk), .A(\g.we_clk [4868]));
Q_ASSIGN U11523 ( .B(clk), .A(\g.we_clk [4867]));
Q_ASSIGN U11524 ( .B(clk), .A(\g.we_clk [4866]));
Q_ASSIGN U11525 ( .B(clk), .A(\g.we_clk [4865]));
Q_ASSIGN U11526 ( .B(clk), .A(\g.we_clk [4864]));
Q_ASSIGN U11527 ( .B(clk), .A(\g.we_clk [4863]));
Q_ASSIGN U11528 ( .B(clk), .A(\g.we_clk [4862]));
Q_ASSIGN U11529 ( .B(clk), .A(\g.we_clk [4861]));
Q_ASSIGN U11530 ( .B(clk), .A(\g.we_clk [4860]));
Q_ASSIGN U11531 ( .B(clk), .A(\g.we_clk [4859]));
Q_ASSIGN U11532 ( .B(clk), .A(\g.we_clk [4858]));
Q_ASSIGN U11533 ( .B(clk), .A(\g.we_clk [4857]));
Q_ASSIGN U11534 ( .B(clk), .A(\g.we_clk [4856]));
Q_ASSIGN U11535 ( .B(clk), .A(\g.we_clk [4855]));
Q_ASSIGN U11536 ( .B(clk), .A(\g.we_clk [4854]));
Q_ASSIGN U11537 ( .B(clk), .A(\g.we_clk [4853]));
Q_ASSIGN U11538 ( .B(clk), .A(\g.we_clk [4852]));
Q_ASSIGN U11539 ( .B(clk), .A(\g.we_clk [4851]));
Q_ASSIGN U11540 ( .B(clk), .A(\g.we_clk [4850]));
Q_ASSIGN U11541 ( .B(clk), .A(\g.we_clk [4849]));
Q_ASSIGN U11542 ( .B(clk), .A(\g.we_clk [4848]));
Q_ASSIGN U11543 ( .B(clk), .A(\g.we_clk [4847]));
Q_ASSIGN U11544 ( .B(clk), .A(\g.we_clk [4846]));
Q_ASSIGN U11545 ( .B(clk), .A(\g.we_clk [4845]));
Q_ASSIGN U11546 ( .B(clk), .A(\g.we_clk [4844]));
Q_ASSIGN U11547 ( .B(clk), .A(\g.we_clk [4843]));
Q_ASSIGN U11548 ( .B(clk), .A(\g.we_clk [4842]));
Q_ASSIGN U11549 ( .B(clk), .A(\g.we_clk [4841]));
Q_ASSIGN U11550 ( .B(clk), .A(\g.we_clk [4840]));
Q_ASSIGN U11551 ( .B(clk), .A(\g.we_clk [4839]));
Q_ASSIGN U11552 ( .B(clk), .A(\g.we_clk [4838]));
Q_ASSIGN U11553 ( .B(clk), .A(\g.we_clk [4837]));
Q_ASSIGN U11554 ( .B(clk), .A(\g.we_clk [4836]));
Q_ASSIGN U11555 ( .B(clk), .A(\g.we_clk [4835]));
Q_ASSIGN U11556 ( .B(clk), .A(\g.we_clk [4834]));
Q_ASSIGN U11557 ( .B(clk), .A(\g.we_clk [4833]));
Q_ASSIGN U11558 ( .B(clk), .A(\g.we_clk [4832]));
Q_ASSIGN U11559 ( .B(clk), .A(\g.we_clk [4831]));
Q_ASSIGN U11560 ( .B(clk), .A(\g.we_clk [4830]));
Q_ASSIGN U11561 ( .B(clk), .A(\g.we_clk [4829]));
Q_ASSIGN U11562 ( .B(clk), .A(\g.we_clk [4828]));
Q_ASSIGN U11563 ( .B(clk), .A(\g.we_clk [4827]));
Q_ASSIGN U11564 ( .B(clk), .A(\g.we_clk [4826]));
Q_ASSIGN U11565 ( .B(clk), .A(\g.we_clk [4825]));
Q_ASSIGN U11566 ( .B(clk), .A(\g.we_clk [4824]));
Q_ASSIGN U11567 ( .B(clk), .A(\g.we_clk [4823]));
Q_ASSIGN U11568 ( .B(clk), .A(\g.we_clk [4822]));
Q_ASSIGN U11569 ( .B(clk), .A(\g.we_clk [4821]));
Q_ASSIGN U11570 ( .B(clk), .A(\g.we_clk [4820]));
Q_ASSIGN U11571 ( .B(clk), .A(\g.we_clk [4819]));
Q_ASSIGN U11572 ( .B(clk), .A(\g.we_clk [4818]));
Q_ASSIGN U11573 ( .B(clk), .A(\g.we_clk [4817]));
Q_ASSIGN U11574 ( .B(clk), .A(\g.we_clk [4816]));
Q_ASSIGN U11575 ( .B(clk), .A(\g.we_clk [4815]));
Q_ASSIGN U11576 ( .B(clk), .A(\g.we_clk [4814]));
Q_ASSIGN U11577 ( .B(clk), .A(\g.we_clk [4813]));
Q_ASSIGN U11578 ( .B(clk), .A(\g.we_clk [4812]));
Q_ASSIGN U11579 ( .B(clk), .A(\g.we_clk [4811]));
Q_ASSIGN U11580 ( .B(clk), .A(\g.we_clk [4810]));
Q_ASSIGN U11581 ( .B(clk), .A(\g.we_clk [4809]));
Q_ASSIGN U11582 ( .B(clk), .A(\g.we_clk [4808]));
Q_ASSIGN U11583 ( .B(clk), .A(\g.we_clk [4807]));
Q_ASSIGN U11584 ( .B(clk), .A(\g.we_clk [4806]));
Q_ASSIGN U11585 ( .B(clk), .A(\g.we_clk [4805]));
Q_ASSIGN U11586 ( .B(clk), .A(\g.we_clk [4804]));
Q_ASSIGN U11587 ( .B(clk), .A(\g.we_clk [4803]));
Q_ASSIGN U11588 ( .B(clk), .A(\g.we_clk [4802]));
Q_ASSIGN U11589 ( .B(clk), .A(\g.we_clk [4801]));
Q_ASSIGN U11590 ( .B(clk), .A(\g.we_clk [4800]));
Q_ASSIGN U11591 ( .B(clk), .A(\g.we_clk [4799]));
Q_ASSIGN U11592 ( .B(clk), .A(\g.we_clk [4798]));
Q_ASSIGN U11593 ( .B(clk), .A(\g.we_clk [4797]));
Q_ASSIGN U11594 ( .B(clk), .A(\g.we_clk [4796]));
Q_ASSIGN U11595 ( .B(clk), .A(\g.we_clk [4795]));
Q_ASSIGN U11596 ( .B(clk), .A(\g.we_clk [4794]));
Q_ASSIGN U11597 ( .B(clk), .A(\g.we_clk [4793]));
Q_ASSIGN U11598 ( .B(clk), .A(\g.we_clk [4792]));
Q_ASSIGN U11599 ( .B(clk), .A(\g.we_clk [4791]));
Q_ASSIGN U11600 ( .B(clk), .A(\g.we_clk [4790]));
Q_ASSIGN U11601 ( .B(clk), .A(\g.we_clk [4789]));
Q_ASSIGN U11602 ( .B(clk), .A(\g.we_clk [4788]));
Q_ASSIGN U11603 ( .B(clk), .A(\g.we_clk [4787]));
Q_ASSIGN U11604 ( .B(clk), .A(\g.we_clk [4786]));
Q_ASSIGN U11605 ( .B(clk), .A(\g.we_clk [4785]));
Q_ASSIGN U11606 ( .B(clk), .A(\g.we_clk [4784]));
Q_ASSIGN U11607 ( .B(clk), .A(\g.we_clk [4783]));
Q_ASSIGN U11608 ( .B(clk), .A(\g.we_clk [4782]));
Q_ASSIGN U11609 ( .B(clk), .A(\g.we_clk [4781]));
Q_ASSIGN U11610 ( .B(clk), .A(\g.we_clk [4780]));
Q_ASSIGN U11611 ( .B(clk), .A(\g.we_clk [4779]));
Q_ASSIGN U11612 ( .B(clk), .A(\g.we_clk [4778]));
Q_ASSIGN U11613 ( .B(clk), .A(\g.we_clk [4777]));
Q_ASSIGN U11614 ( .B(clk), .A(\g.we_clk [4776]));
Q_ASSIGN U11615 ( .B(clk), .A(\g.we_clk [4775]));
Q_ASSIGN U11616 ( .B(clk), .A(\g.we_clk [4774]));
Q_ASSIGN U11617 ( .B(clk), .A(\g.we_clk [4773]));
Q_ASSIGN U11618 ( .B(clk), .A(\g.we_clk [4772]));
Q_ASSIGN U11619 ( .B(clk), .A(\g.we_clk [4771]));
Q_ASSIGN U11620 ( .B(clk), .A(\g.we_clk [4770]));
Q_ASSIGN U11621 ( .B(clk), .A(\g.we_clk [4769]));
Q_ASSIGN U11622 ( .B(clk), .A(\g.we_clk [4768]));
Q_ASSIGN U11623 ( .B(clk), .A(\g.we_clk [4767]));
Q_ASSIGN U11624 ( .B(clk), .A(\g.we_clk [4766]));
Q_ASSIGN U11625 ( .B(clk), .A(\g.we_clk [4765]));
Q_ASSIGN U11626 ( .B(clk), .A(\g.we_clk [4764]));
Q_ASSIGN U11627 ( .B(clk), .A(\g.we_clk [4763]));
Q_ASSIGN U11628 ( .B(clk), .A(\g.we_clk [4762]));
Q_ASSIGN U11629 ( .B(clk), .A(\g.we_clk [4761]));
Q_ASSIGN U11630 ( .B(clk), .A(\g.we_clk [4760]));
Q_ASSIGN U11631 ( .B(clk), .A(\g.we_clk [4759]));
Q_ASSIGN U11632 ( .B(clk), .A(\g.we_clk [4758]));
Q_ASSIGN U11633 ( .B(clk), .A(\g.we_clk [4757]));
Q_ASSIGN U11634 ( .B(clk), .A(\g.we_clk [4756]));
Q_ASSIGN U11635 ( .B(clk), .A(\g.we_clk [4755]));
Q_ASSIGN U11636 ( .B(clk), .A(\g.we_clk [4754]));
Q_ASSIGN U11637 ( .B(clk), .A(\g.we_clk [4753]));
Q_ASSIGN U11638 ( .B(clk), .A(\g.we_clk [4752]));
Q_ASSIGN U11639 ( .B(clk), .A(\g.we_clk [4751]));
Q_ASSIGN U11640 ( .B(clk), .A(\g.we_clk [4750]));
Q_ASSIGN U11641 ( .B(clk), .A(\g.we_clk [4749]));
Q_ASSIGN U11642 ( .B(clk), .A(\g.we_clk [4748]));
Q_ASSIGN U11643 ( .B(clk), .A(\g.we_clk [4747]));
Q_ASSIGN U11644 ( .B(clk), .A(\g.we_clk [4746]));
Q_ASSIGN U11645 ( .B(clk), .A(\g.we_clk [4745]));
Q_ASSIGN U11646 ( .B(clk), .A(\g.we_clk [4744]));
Q_ASSIGN U11647 ( .B(clk), .A(\g.we_clk [4743]));
Q_ASSIGN U11648 ( .B(clk), .A(\g.we_clk [4742]));
Q_ASSIGN U11649 ( .B(clk), .A(\g.we_clk [4741]));
Q_ASSIGN U11650 ( .B(clk), .A(\g.we_clk [4740]));
Q_ASSIGN U11651 ( .B(clk), .A(\g.we_clk [4739]));
Q_ASSIGN U11652 ( .B(clk), .A(\g.we_clk [4738]));
Q_ASSIGN U11653 ( .B(clk), .A(\g.we_clk [4737]));
Q_ASSIGN U11654 ( .B(clk), .A(\g.we_clk [4736]));
Q_ASSIGN U11655 ( .B(clk), .A(\g.we_clk [4735]));
Q_ASSIGN U11656 ( .B(clk), .A(\g.we_clk [4734]));
Q_ASSIGN U11657 ( .B(clk), .A(\g.we_clk [4733]));
Q_ASSIGN U11658 ( .B(clk), .A(\g.we_clk [4732]));
Q_ASSIGN U11659 ( .B(clk), .A(\g.we_clk [4731]));
Q_ASSIGN U11660 ( .B(clk), .A(\g.we_clk [4730]));
Q_ASSIGN U11661 ( .B(clk), .A(\g.we_clk [4729]));
Q_ASSIGN U11662 ( .B(clk), .A(\g.we_clk [4728]));
Q_ASSIGN U11663 ( .B(clk), .A(\g.we_clk [4727]));
Q_ASSIGN U11664 ( .B(clk), .A(\g.we_clk [4726]));
Q_ASSIGN U11665 ( .B(clk), .A(\g.we_clk [4725]));
Q_ASSIGN U11666 ( .B(clk), .A(\g.we_clk [4724]));
Q_ASSIGN U11667 ( .B(clk), .A(\g.we_clk [4723]));
Q_ASSIGN U11668 ( .B(clk), .A(\g.we_clk [4722]));
Q_ASSIGN U11669 ( .B(clk), .A(\g.we_clk [4721]));
Q_ASSIGN U11670 ( .B(clk), .A(\g.we_clk [4720]));
Q_ASSIGN U11671 ( .B(clk), .A(\g.we_clk [4719]));
Q_ASSIGN U11672 ( .B(clk), .A(\g.we_clk [4718]));
Q_ASSIGN U11673 ( .B(clk), .A(\g.we_clk [4717]));
Q_ASSIGN U11674 ( .B(clk), .A(\g.we_clk [4716]));
Q_ASSIGN U11675 ( .B(clk), .A(\g.we_clk [4715]));
Q_ASSIGN U11676 ( .B(clk), .A(\g.we_clk [4714]));
Q_ASSIGN U11677 ( .B(clk), .A(\g.we_clk [4713]));
Q_ASSIGN U11678 ( .B(clk), .A(\g.we_clk [4712]));
Q_ASSIGN U11679 ( .B(clk), .A(\g.we_clk [4711]));
Q_ASSIGN U11680 ( .B(clk), .A(\g.we_clk [4710]));
Q_ASSIGN U11681 ( .B(clk), .A(\g.we_clk [4709]));
Q_ASSIGN U11682 ( .B(clk), .A(\g.we_clk [4708]));
Q_ASSIGN U11683 ( .B(clk), .A(\g.we_clk [4707]));
Q_ASSIGN U11684 ( .B(clk), .A(\g.we_clk [4706]));
Q_ASSIGN U11685 ( .B(clk), .A(\g.we_clk [4705]));
Q_ASSIGN U11686 ( .B(clk), .A(\g.we_clk [4704]));
Q_ASSIGN U11687 ( .B(clk), .A(\g.we_clk [4703]));
Q_ASSIGN U11688 ( .B(clk), .A(\g.we_clk [4702]));
Q_ASSIGN U11689 ( .B(clk), .A(\g.we_clk [4701]));
Q_ASSIGN U11690 ( .B(clk), .A(\g.we_clk [4700]));
Q_ASSIGN U11691 ( .B(clk), .A(\g.we_clk [4699]));
Q_ASSIGN U11692 ( .B(clk), .A(\g.we_clk [4698]));
Q_ASSIGN U11693 ( .B(clk), .A(\g.we_clk [4697]));
Q_ASSIGN U11694 ( .B(clk), .A(\g.we_clk [4696]));
Q_ASSIGN U11695 ( .B(clk), .A(\g.we_clk [4695]));
Q_ASSIGN U11696 ( .B(clk), .A(\g.we_clk [4694]));
Q_ASSIGN U11697 ( .B(clk), .A(\g.we_clk [4693]));
Q_ASSIGN U11698 ( .B(clk), .A(\g.we_clk [4692]));
Q_ASSIGN U11699 ( .B(clk), .A(\g.we_clk [4691]));
Q_ASSIGN U11700 ( .B(clk), .A(\g.we_clk [4690]));
Q_ASSIGN U11701 ( .B(clk), .A(\g.we_clk [4689]));
Q_ASSIGN U11702 ( .B(clk), .A(\g.we_clk [4688]));
Q_ASSIGN U11703 ( .B(clk), .A(\g.we_clk [4687]));
Q_ASSIGN U11704 ( .B(clk), .A(\g.we_clk [4686]));
Q_ASSIGN U11705 ( .B(clk), .A(\g.we_clk [4685]));
Q_ASSIGN U11706 ( .B(clk), .A(\g.we_clk [4684]));
Q_ASSIGN U11707 ( .B(clk), .A(\g.we_clk [4683]));
Q_ASSIGN U11708 ( .B(clk), .A(\g.we_clk [4682]));
Q_ASSIGN U11709 ( .B(clk), .A(\g.we_clk [4681]));
Q_ASSIGN U11710 ( .B(clk), .A(\g.we_clk [4680]));
Q_ASSIGN U11711 ( .B(clk), .A(\g.we_clk [4679]));
Q_ASSIGN U11712 ( .B(clk), .A(\g.we_clk [4678]));
Q_ASSIGN U11713 ( .B(clk), .A(\g.we_clk [4677]));
Q_ASSIGN U11714 ( .B(clk), .A(\g.we_clk [4676]));
Q_ASSIGN U11715 ( .B(clk), .A(\g.we_clk [4675]));
Q_ASSIGN U11716 ( .B(clk), .A(\g.we_clk [4674]));
Q_ASSIGN U11717 ( .B(clk), .A(\g.we_clk [4673]));
Q_ASSIGN U11718 ( .B(clk), .A(\g.we_clk [4672]));
Q_ASSIGN U11719 ( .B(clk), .A(\g.we_clk [4671]));
Q_ASSIGN U11720 ( .B(clk), .A(\g.we_clk [4670]));
Q_ASSIGN U11721 ( .B(clk), .A(\g.we_clk [4669]));
Q_ASSIGN U11722 ( .B(clk), .A(\g.we_clk [4668]));
Q_ASSIGN U11723 ( .B(clk), .A(\g.we_clk [4667]));
Q_ASSIGN U11724 ( .B(clk), .A(\g.we_clk [4666]));
Q_ASSIGN U11725 ( .B(clk), .A(\g.we_clk [4665]));
Q_ASSIGN U11726 ( .B(clk), .A(\g.we_clk [4664]));
Q_ASSIGN U11727 ( .B(clk), .A(\g.we_clk [4663]));
Q_ASSIGN U11728 ( .B(clk), .A(\g.we_clk [4662]));
Q_ASSIGN U11729 ( .B(clk), .A(\g.we_clk [4661]));
Q_ASSIGN U11730 ( .B(clk), .A(\g.we_clk [4660]));
Q_ASSIGN U11731 ( .B(clk), .A(\g.we_clk [4659]));
Q_ASSIGN U11732 ( .B(clk), .A(\g.we_clk [4658]));
Q_ASSIGN U11733 ( .B(clk), .A(\g.we_clk [4657]));
Q_ASSIGN U11734 ( .B(clk), .A(\g.we_clk [4656]));
Q_ASSIGN U11735 ( .B(clk), .A(\g.we_clk [4655]));
Q_ASSIGN U11736 ( .B(clk), .A(\g.we_clk [4654]));
Q_ASSIGN U11737 ( .B(clk), .A(\g.we_clk [4653]));
Q_ASSIGN U11738 ( .B(clk), .A(\g.we_clk [4652]));
Q_ASSIGN U11739 ( .B(clk), .A(\g.we_clk [4651]));
Q_ASSIGN U11740 ( .B(clk), .A(\g.we_clk [4650]));
Q_ASSIGN U11741 ( .B(clk), .A(\g.we_clk [4649]));
Q_ASSIGN U11742 ( .B(clk), .A(\g.we_clk [4648]));
Q_ASSIGN U11743 ( .B(clk), .A(\g.we_clk [4647]));
Q_ASSIGN U11744 ( .B(clk), .A(\g.we_clk [4646]));
Q_ASSIGN U11745 ( .B(clk), .A(\g.we_clk [4645]));
Q_ASSIGN U11746 ( .B(clk), .A(\g.we_clk [4644]));
Q_ASSIGN U11747 ( .B(clk), .A(\g.we_clk [4643]));
Q_ASSIGN U11748 ( .B(clk), .A(\g.we_clk [4642]));
Q_ASSIGN U11749 ( .B(clk), .A(\g.we_clk [4641]));
Q_ASSIGN U11750 ( .B(clk), .A(\g.we_clk [4640]));
Q_ASSIGN U11751 ( .B(clk), .A(\g.we_clk [4639]));
Q_ASSIGN U11752 ( .B(clk), .A(\g.we_clk [4638]));
Q_ASSIGN U11753 ( .B(clk), .A(\g.we_clk [4637]));
Q_ASSIGN U11754 ( .B(clk), .A(\g.we_clk [4636]));
Q_ASSIGN U11755 ( .B(clk), .A(\g.we_clk [4635]));
Q_ASSIGN U11756 ( .B(clk), .A(\g.we_clk [4634]));
Q_ASSIGN U11757 ( .B(clk), .A(\g.we_clk [4633]));
Q_ASSIGN U11758 ( .B(clk), .A(\g.we_clk [4632]));
Q_ASSIGN U11759 ( .B(clk), .A(\g.we_clk [4631]));
Q_ASSIGN U11760 ( .B(clk), .A(\g.we_clk [4630]));
Q_ASSIGN U11761 ( .B(clk), .A(\g.we_clk [4629]));
Q_ASSIGN U11762 ( .B(clk), .A(\g.we_clk [4628]));
Q_ASSIGN U11763 ( .B(clk), .A(\g.we_clk [4627]));
Q_ASSIGN U11764 ( .B(clk), .A(\g.we_clk [4626]));
Q_ASSIGN U11765 ( .B(clk), .A(\g.we_clk [4625]));
Q_ASSIGN U11766 ( .B(clk), .A(\g.we_clk [4624]));
Q_ASSIGN U11767 ( .B(clk), .A(\g.we_clk [4623]));
Q_ASSIGN U11768 ( .B(clk), .A(\g.we_clk [4622]));
Q_ASSIGN U11769 ( .B(clk), .A(\g.we_clk [4621]));
Q_ASSIGN U11770 ( .B(clk), .A(\g.we_clk [4620]));
Q_ASSIGN U11771 ( .B(clk), .A(\g.we_clk [4619]));
Q_ASSIGN U11772 ( .B(clk), .A(\g.we_clk [4618]));
Q_ASSIGN U11773 ( .B(clk), .A(\g.we_clk [4617]));
Q_ASSIGN U11774 ( .B(clk), .A(\g.we_clk [4616]));
Q_ASSIGN U11775 ( .B(clk), .A(\g.we_clk [4615]));
Q_ASSIGN U11776 ( .B(clk), .A(\g.we_clk [4614]));
Q_ASSIGN U11777 ( .B(clk), .A(\g.we_clk [4613]));
Q_ASSIGN U11778 ( .B(clk), .A(\g.we_clk [4612]));
Q_ASSIGN U11779 ( .B(clk), .A(\g.we_clk [4611]));
Q_ASSIGN U11780 ( .B(clk), .A(\g.we_clk [4610]));
Q_ASSIGN U11781 ( .B(clk), .A(\g.we_clk [4609]));
Q_ASSIGN U11782 ( .B(clk), .A(\g.we_clk [4608]));
Q_ASSIGN U11783 ( .B(clk), .A(\g.we_clk [4607]));
Q_ASSIGN U11784 ( .B(clk), .A(\g.we_clk [4606]));
Q_ASSIGN U11785 ( .B(clk), .A(\g.we_clk [4605]));
Q_ASSIGN U11786 ( .B(clk), .A(\g.we_clk [4604]));
Q_ASSIGN U11787 ( .B(clk), .A(\g.we_clk [4603]));
Q_ASSIGN U11788 ( .B(clk), .A(\g.we_clk [4602]));
Q_ASSIGN U11789 ( .B(clk), .A(\g.we_clk [4601]));
Q_ASSIGN U11790 ( .B(clk), .A(\g.we_clk [4600]));
Q_ASSIGN U11791 ( .B(clk), .A(\g.we_clk [4599]));
Q_ASSIGN U11792 ( .B(clk), .A(\g.we_clk [4598]));
Q_ASSIGN U11793 ( .B(clk), .A(\g.we_clk [4597]));
Q_ASSIGN U11794 ( .B(clk), .A(\g.we_clk [4596]));
Q_ASSIGN U11795 ( .B(clk), .A(\g.we_clk [4595]));
Q_ASSIGN U11796 ( .B(clk), .A(\g.we_clk [4594]));
Q_ASSIGN U11797 ( .B(clk), .A(\g.we_clk [4593]));
Q_ASSIGN U11798 ( .B(clk), .A(\g.we_clk [4592]));
Q_ASSIGN U11799 ( .B(clk), .A(\g.we_clk [4591]));
Q_ASSIGN U11800 ( .B(clk), .A(\g.we_clk [4590]));
Q_ASSIGN U11801 ( .B(clk), .A(\g.we_clk [4589]));
Q_ASSIGN U11802 ( .B(clk), .A(\g.we_clk [4588]));
Q_ASSIGN U11803 ( .B(clk), .A(\g.we_clk [4587]));
Q_ASSIGN U11804 ( .B(clk), .A(\g.we_clk [4586]));
Q_ASSIGN U11805 ( .B(clk), .A(\g.we_clk [4585]));
Q_ASSIGN U11806 ( .B(clk), .A(\g.we_clk [4584]));
Q_ASSIGN U11807 ( .B(clk), .A(\g.we_clk [4583]));
Q_ASSIGN U11808 ( .B(clk), .A(\g.we_clk [4582]));
Q_ASSIGN U11809 ( .B(clk), .A(\g.we_clk [4581]));
Q_ASSIGN U11810 ( .B(clk), .A(\g.we_clk [4580]));
Q_ASSIGN U11811 ( .B(clk), .A(\g.we_clk [4579]));
Q_ASSIGN U11812 ( .B(clk), .A(\g.we_clk [4578]));
Q_ASSIGN U11813 ( .B(clk), .A(\g.we_clk [4577]));
Q_ASSIGN U11814 ( .B(clk), .A(\g.we_clk [4576]));
Q_ASSIGN U11815 ( .B(clk), .A(\g.we_clk [4575]));
Q_ASSIGN U11816 ( .B(clk), .A(\g.we_clk [4574]));
Q_ASSIGN U11817 ( .B(clk), .A(\g.we_clk [4573]));
Q_ASSIGN U11818 ( .B(clk), .A(\g.we_clk [4572]));
Q_ASSIGN U11819 ( .B(clk), .A(\g.we_clk [4571]));
Q_ASSIGN U11820 ( .B(clk), .A(\g.we_clk [4570]));
Q_ASSIGN U11821 ( .B(clk), .A(\g.we_clk [4569]));
Q_ASSIGN U11822 ( .B(clk), .A(\g.we_clk [4568]));
Q_ASSIGN U11823 ( .B(clk), .A(\g.we_clk [4567]));
Q_ASSIGN U11824 ( .B(clk), .A(\g.we_clk [4566]));
Q_ASSIGN U11825 ( .B(clk), .A(\g.we_clk [4565]));
Q_ASSIGN U11826 ( .B(clk), .A(\g.we_clk [4564]));
Q_ASSIGN U11827 ( .B(clk), .A(\g.we_clk [4563]));
Q_ASSIGN U11828 ( .B(clk), .A(\g.we_clk [4562]));
Q_ASSIGN U11829 ( .B(clk), .A(\g.we_clk [4561]));
Q_ASSIGN U11830 ( .B(clk), .A(\g.we_clk [4560]));
Q_ASSIGN U11831 ( .B(clk), .A(\g.we_clk [4559]));
Q_ASSIGN U11832 ( .B(clk), .A(\g.we_clk [4558]));
Q_ASSIGN U11833 ( .B(clk), .A(\g.we_clk [4557]));
Q_ASSIGN U11834 ( .B(clk), .A(\g.we_clk [4556]));
Q_ASSIGN U11835 ( .B(clk), .A(\g.we_clk [4555]));
Q_ASSIGN U11836 ( .B(clk), .A(\g.we_clk [4554]));
Q_ASSIGN U11837 ( .B(clk), .A(\g.we_clk [4553]));
Q_ASSIGN U11838 ( .B(clk), .A(\g.we_clk [4552]));
Q_ASSIGN U11839 ( .B(clk), .A(\g.we_clk [4551]));
Q_ASSIGN U11840 ( .B(clk), .A(\g.we_clk [4550]));
Q_ASSIGN U11841 ( .B(clk), .A(\g.we_clk [4549]));
Q_ASSIGN U11842 ( .B(clk), .A(\g.we_clk [4548]));
Q_ASSIGN U11843 ( .B(clk), .A(\g.we_clk [4547]));
Q_ASSIGN U11844 ( .B(clk), .A(\g.we_clk [4546]));
Q_ASSIGN U11845 ( .B(clk), .A(\g.we_clk [4545]));
Q_ASSIGN U11846 ( .B(clk), .A(\g.we_clk [4544]));
Q_ASSIGN U11847 ( .B(clk), .A(\g.we_clk [4543]));
Q_ASSIGN U11848 ( .B(clk), .A(\g.we_clk [4542]));
Q_ASSIGN U11849 ( .B(clk), .A(\g.we_clk [4541]));
Q_ASSIGN U11850 ( .B(clk), .A(\g.we_clk [4540]));
Q_ASSIGN U11851 ( .B(clk), .A(\g.we_clk [4539]));
Q_ASSIGN U11852 ( .B(clk), .A(\g.we_clk [4538]));
Q_ASSIGN U11853 ( .B(clk), .A(\g.we_clk [4537]));
Q_ASSIGN U11854 ( .B(clk), .A(\g.we_clk [4536]));
Q_ASSIGN U11855 ( .B(clk), .A(\g.we_clk [4535]));
Q_ASSIGN U11856 ( .B(clk), .A(\g.we_clk [4534]));
Q_ASSIGN U11857 ( .B(clk), .A(\g.we_clk [4533]));
Q_ASSIGN U11858 ( .B(clk), .A(\g.we_clk [4532]));
Q_ASSIGN U11859 ( .B(clk), .A(\g.we_clk [4531]));
Q_ASSIGN U11860 ( .B(clk), .A(\g.we_clk [4530]));
Q_ASSIGN U11861 ( .B(clk), .A(\g.we_clk [4529]));
Q_ASSIGN U11862 ( .B(clk), .A(\g.we_clk [4528]));
Q_ASSIGN U11863 ( .B(clk), .A(\g.we_clk [4527]));
Q_ASSIGN U11864 ( .B(clk), .A(\g.we_clk [4526]));
Q_ASSIGN U11865 ( .B(clk), .A(\g.we_clk [4525]));
Q_ASSIGN U11866 ( .B(clk), .A(\g.we_clk [4524]));
Q_ASSIGN U11867 ( .B(clk), .A(\g.we_clk [4523]));
Q_ASSIGN U11868 ( .B(clk), .A(\g.we_clk [4522]));
Q_ASSIGN U11869 ( .B(clk), .A(\g.we_clk [4521]));
Q_ASSIGN U11870 ( .B(clk), .A(\g.we_clk [4520]));
Q_ASSIGN U11871 ( .B(clk), .A(\g.we_clk [4519]));
Q_ASSIGN U11872 ( .B(clk), .A(\g.we_clk [4518]));
Q_ASSIGN U11873 ( .B(clk), .A(\g.we_clk [4517]));
Q_ASSIGN U11874 ( .B(clk), .A(\g.we_clk [4516]));
Q_ASSIGN U11875 ( .B(clk), .A(\g.we_clk [4515]));
Q_ASSIGN U11876 ( .B(clk), .A(\g.we_clk [4514]));
Q_ASSIGN U11877 ( .B(clk), .A(\g.we_clk [4513]));
Q_ASSIGN U11878 ( .B(clk), .A(\g.we_clk [4512]));
Q_ASSIGN U11879 ( .B(clk), .A(\g.we_clk [4511]));
Q_ASSIGN U11880 ( .B(clk), .A(\g.we_clk [4510]));
Q_ASSIGN U11881 ( .B(clk), .A(\g.we_clk [4509]));
Q_ASSIGN U11882 ( .B(clk), .A(\g.we_clk [4508]));
Q_ASSIGN U11883 ( .B(clk), .A(\g.we_clk [4507]));
Q_ASSIGN U11884 ( .B(clk), .A(\g.we_clk [4506]));
Q_ASSIGN U11885 ( .B(clk), .A(\g.we_clk [4505]));
Q_ASSIGN U11886 ( .B(clk), .A(\g.we_clk [4504]));
Q_ASSIGN U11887 ( .B(clk), .A(\g.we_clk [4503]));
Q_ASSIGN U11888 ( .B(clk), .A(\g.we_clk [4502]));
Q_ASSIGN U11889 ( .B(clk), .A(\g.we_clk [4501]));
Q_ASSIGN U11890 ( .B(clk), .A(\g.we_clk [4500]));
Q_ASSIGN U11891 ( .B(clk), .A(\g.we_clk [4499]));
Q_ASSIGN U11892 ( .B(clk), .A(\g.we_clk [4498]));
Q_ASSIGN U11893 ( .B(clk), .A(\g.we_clk [4497]));
Q_ASSIGN U11894 ( .B(clk), .A(\g.we_clk [4496]));
Q_ASSIGN U11895 ( .B(clk), .A(\g.we_clk [4495]));
Q_ASSIGN U11896 ( .B(clk), .A(\g.we_clk [4494]));
Q_ASSIGN U11897 ( .B(clk), .A(\g.we_clk [4493]));
Q_ASSIGN U11898 ( .B(clk), .A(\g.we_clk [4492]));
Q_ASSIGN U11899 ( .B(clk), .A(\g.we_clk [4491]));
Q_ASSIGN U11900 ( .B(clk), .A(\g.we_clk [4490]));
Q_ASSIGN U11901 ( .B(clk), .A(\g.we_clk [4489]));
Q_ASSIGN U11902 ( .B(clk), .A(\g.we_clk [4488]));
Q_ASSIGN U11903 ( .B(clk), .A(\g.we_clk [4487]));
Q_ASSIGN U11904 ( .B(clk), .A(\g.we_clk [4486]));
Q_ASSIGN U11905 ( .B(clk), .A(\g.we_clk [4485]));
Q_ASSIGN U11906 ( .B(clk), .A(\g.we_clk [4484]));
Q_ASSIGN U11907 ( .B(clk), .A(\g.we_clk [4483]));
Q_ASSIGN U11908 ( .B(clk), .A(\g.we_clk [4482]));
Q_ASSIGN U11909 ( .B(clk), .A(\g.we_clk [4481]));
Q_ASSIGN U11910 ( .B(clk), .A(\g.we_clk [4480]));
Q_ASSIGN U11911 ( .B(clk), .A(\g.we_clk [4479]));
Q_ASSIGN U11912 ( .B(clk), .A(\g.we_clk [4478]));
Q_ASSIGN U11913 ( .B(clk), .A(\g.we_clk [4477]));
Q_ASSIGN U11914 ( .B(clk), .A(\g.we_clk [4476]));
Q_ASSIGN U11915 ( .B(clk), .A(\g.we_clk [4475]));
Q_ASSIGN U11916 ( .B(clk), .A(\g.we_clk [4474]));
Q_ASSIGN U11917 ( .B(clk), .A(\g.we_clk [4473]));
Q_ASSIGN U11918 ( .B(clk), .A(\g.we_clk [4472]));
Q_ASSIGN U11919 ( .B(clk), .A(\g.we_clk [4471]));
Q_ASSIGN U11920 ( .B(clk), .A(\g.we_clk [4470]));
Q_ASSIGN U11921 ( .B(clk), .A(\g.we_clk [4469]));
Q_ASSIGN U11922 ( .B(clk), .A(\g.we_clk [4468]));
Q_ASSIGN U11923 ( .B(clk), .A(\g.we_clk [4467]));
Q_ASSIGN U11924 ( .B(clk), .A(\g.we_clk [4466]));
Q_ASSIGN U11925 ( .B(clk), .A(\g.we_clk [4465]));
Q_ASSIGN U11926 ( .B(clk), .A(\g.we_clk [4464]));
Q_ASSIGN U11927 ( .B(clk), .A(\g.we_clk [4463]));
Q_ASSIGN U11928 ( .B(clk), .A(\g.we_clk [4462]));
Q_ASSIGN U11929 ( .B(clk), .A(\g.we_clk [4461]));
Q_ASSIGN U11930 ( .B(clk), .A(\g.we_clk [4460]));
Q_ASSIGN U11931 ( .B(clk), .A(\g.we_clk [4459]));
Q_ASSIGN U11932 ( .B(clk), .A(\g.we_clk [4458]));
Q_ASSIGN U11933 ( .B(clk), .A(\g.we_clk [4457]));
Q_ASSIGN U11934 ( .B(clk), .A(\g.we_clk [4456]));
Q_ASSIGN U11935 ( .B(clk), .A(\g.we_clk [4455]));
Q_ASSIGN U11936 ( .B(clk), .A(\g.we_clk [4454]));
Q_ASSIGN U11937 ( .B(clk), .A(\g.we_clk [4453]));
Q_ASSIGN U11938 ( .B(clk), .A(\g.we_clk [4452]));
Q_ASSIGN U11939 ( .B(clk), .A(\g.we_clk [4451]));
Q_ASSIGN U11940 ( .B(clk), .A(\g.we_clk [4450]));
Q_ASSIGN U11941 ( .B(clk), .A(\g.we_clk [4449]));
Q_ASSIGN U11942 ( .B(clk), .A(\g.we_clk [4448]));
Q_ASSIGN U11943 ( .B(clk), .A(\g.we_clk [4447]));
Q_ASSIGN U11944 ( .B(clk), .A(\g.we_clk [4446]));
Q_ASSIGN U11945 ( .B(clk), .A(\g.we_clk [4445]));
Q_ASSIGN U11946 ( .B(clk), .A(\g.we_clk [4444]));
Q_ASSIGN U11947 ( .B(clk), .A(\g.we_clk [4443]));
Q_ASSIGN U11948 ( .B(clk), .A(\g.we_clk [4442]));
Q_ASSIGN U11949 ( .B(clk), .A(\g.we_clk [4441]));
Q_ASSIGN U11950 ( .B(clk), .A(\g.we_clk [4440]));
Q_ASSIGN U11951 ( .B(clk), .A(\g.we_clk [4439]));
Q_ASSIGN U11952 ( .B(clk), .A(\g.we_clk [4438]));
Q_ASSIGN U11953 ( .B(clk), .A(\g.we_clk [4437]));
Q_ASSIGN U11954 ( .B(clk), .A(\g.we_clk [4436]));
Q_ASSIGN U11955 ( .B(clk), .A(\g.we_clk [4435]));
Q_ASSIGN U11956 ( .B(clk), .A(\g.we_clk [4434]));
Q_ASSIGN U11957 ( .B(clk), .A(\g.we_clk [4433]));
Q_ASSIGN U11958 ( .B(clk), .A(\g.we_clk [4432]));
Q_ASSIGN U11959 ( .B(clk), .A(\g.we_clk [4431]));
Q_ASSIGN U11960 ( .B(clk), .A(\g.we_clk [4430]));
Q_ASSIGN U11961 ( .B(clk), .A(\g.we_clk [4429]));
Q_ASSIGN U11962 ( .B(clk), .A(\g.we_clk [4428]));
Q_ASSIGN U11963 ( .B(clk), .A(\g.we_clk [4427]));
Q_ASSIGN U11964 ( .B(clk), .A(\g.we_clk [4426]));
Q_ASSIGN U11965 ( .B(clk), .A(\g.we_clk [4425]));
Q_ASSIGN U11966 ( .B(clk), .A(\g.we_clk [4424]));
Q_ASSIGN U11967 ( .B(clk), .A(\g.we_clk [4423]));
Q_ASSIGN U11968 ( .B(clk), .A(\g.we_clk [4422]));
Q_ASSIGN U11969 ( .B(clk), .A(\g.we_clk [4421]));
Q_ASSIGN U11970 ( .B(clk), .A(\g.we_clk [4420]));
Q_ASSIGN U11971 ( .B(clk), .A(\g.we_clk [4419]));
Q_ASSIGN U11972 ( .B(clk), .A(\g.we_clk [4418]));
Q_ASSIGN U11973 ( .B(clk), .A(\g.we_clk [4417]));
Q_ASSIGN U11974 ( .B(clk), .A(\g.we_clk [4416]));
Q_ASSIGN U11975 ( .B(clk), .A(\g.we_clk [4415]));
Q_ASSIGN U11976 ( .B(clk), .A(\g.we_clk [4414]));
Q_ASSIGN U11977 ( .B(clk), .A(\g.we_clk [4413]));
Q_ASSIGN U11978 ( .B(clk), .A(\g.we_clk [4412]));
Q_ASSIGN U11979 ( .B(clk), .A(\g.we_clk [4411]));
Q_ASSIGN U11980 ( .B(clk), .A(\g.we_clk [4410]));
Q_ASSIGN U11981 ( .B(clk), .A(\g.we_clk [4409]));
Q_ASSIGN U11982 ( .B(clk), .A(\g.we_clk [4408]));
Q_ASSIGN U11983 ( .B(clk), .A(\g.we_clk [4407]));
Q_ASSIGN U11984 ( .B(clk), .A(\g.we_clk [4406]));
Q_ASSIGN U11985 ( .B(clk), .A(\g.we_clk [4405]));
Q_ASSIGN U11986 ( .B(clk), .A(\g.we_clk [4404]));
Q_ASSIGN U11987 ( .B(clk), .A(\g.we_clk [4403]));
Q_ASSIGN U11988 ( .B(clk), .A(\g.we_clk [4402]));
Q_ASSIGN U11989 ( .B(clk), .A(\g.we_clk [4401]));
Q_ASSIGN U11990 ( .B(clk), .A(\g.we_clk [4400]));
Q_ASSIGN U11991 ( .B(clk), .A(\g.we_clk [4399]));
Q_ASSIGN U11992 ( .B(clk), .A(\g.we_clk [4398]));
Q_ASSIGN U11993 ( .B(clk), .A(\g.we_clk [4397]));
Q_ASSIGN U11994 ( .B(clk), .A(\g.we_clk [4396]));
Q_ASSIGN U11995 ( .B(clk), .A(\g.we_clk [4395]));
Q_ASSIGN U11996 ( .B(clk), .A(\g.we_clk [4394]));
Q_ASSIGN U11997 ( .B(clk), .A(\g.we_clk [4393]));
Q_ASSIGN U11998 ( .B(clk), .A(\g.we_clk [4392]));
Q_ASSIGN U11999 ( .B(clk), .A(\g.we_clk [4391]));
Q_ASSIGN U12000 ( .B(clk), .A(\g.we_clk [4390]));
Q_ASSIGN U12001 ( .B(clk), .A(\g.we_clk [4389]));
Q_ASSIGN U12002 ( .B(clk), .A(\g.we_clk [4388]));
Q_ASSIGN U12003 ( .B(clk), .A(\g.we_clk [4387]));
Q_ASSIGN U12004 ( .B(clk), .A(\g.we_clk [4386]));
Q_ASSIGN U12005 ( .B(clk), .A(\g.we_clk [4385]));
Q_ASSIGN U12006 ( .B(clk), .A(\g.we_clk [4384]));
Q_ASSIGN U12007 ( .B(clk), .A(\g.we_clk [4383]));
Q_ASSIGN U12008 ( .B(clk), .A(\g.we_clk [4382]));
Q_ASSIGN U12009 ( .B(clk), .A(\g.we_clk [4381]));
Q_ASSIGN U12010 ( .B(clk), .A(\g.we_clk [4380]));
Q_ASSIGN U12011 ( .B(clk), .A(\g.we_clk [4379]));
Q_ASSIGN U12012 ( .B(clk), .A(\g.we_clk [4378]));
Q_ASSIGN U12013 ( .B(clk), .A(\g.we_clk [4377]));
Q_ASSIGN U12014 ( .B(clk), .A(\g.we_clk [4376]));
Q_ASSIGN U12015 ( .B(clk), .A(\g.we_clk [4375]));
Q_ASSIGN U12016 ( .B(clk), .A(\g.we_clk [4374]));
Q_ASSIGN U12017 ( .B(clk), .A(\g.we_clk [4373]));
Q_ASSIGN U12018 ( .B(clk), .A(\g.we_clk [4372]));
Q_ASSIGN U12019 ( .B(clk), .A(\g.we_clk [4371]));
Q_ASSIGN U12020 ( .B(clk), .A(\g.we_clk [4370]));
Q_ASSIGN U12021 ( .B(clk), .A(\g.we_clk [4369]));
Q_ASSIGN U12022 ( .B(clk), .A(\g.we_clk [4368]));
Q_ASSIGN U12023 ( .B(clk), .A(\g.we_clk [4367]));
Q_ASSIGN U12024 ( .B(clk), .A(\g.we_clk [4366]));
Q_ASSIGN U12025 ( .B(clk), .A(\g.we_clk [4365]));
Q_ASSIGN U12026 ( .B(clk), .A(\g.we_clk [4364]));
Q_ASSIGN U12027 ( .B(clk), .A(\g.we_clk [4363]));
Q_ASSIGN U12028 ( .B(clk), .A(\g.we_clk [4362]));
Q_ASSIGN U12029 ( .B(clk), .A(\g.we_clk [4361]));
Q_ASSIGN U12030 ( .B(clk), .A(\g.we_clk [4360]));
Q_ASSIGN U12031 ( .B(clk), .A(\g.we_clk [4359]));
Q_ASSIGN U12032 ( .B(clk), .A(\g.we_clk [4358]));
Q_ASSIGN U12033 ( .B(clk), .A(\g.we_clk [4357]));
Q_ASSIGN U12034 ( .B(clk), .A(\g.we_clk [4356]));
Q_ASSIGN U12035 ( .B(clk), .A(\g.we_clk [4355]));
Q_ASSIGN U12036 ( .B(clk), .A(\g.we_clk [4354]));
Q_ASSIGN U12037 ( .B(clk), .A(\g.we_clk [4353]));
Q_ASSIGN U12038 ( .B(clk), .A(\g.we_clk [4352]));
Q_ASSIGN U12039 ( .B(clk), .A(\g.we_clk [4351]));
Q_ASSIGN U12040 ( .B(clk), .A(\g.we_clk [4350]));
Q_ASSIGN U12041 ( .B(clk), .A(\g.we_clk [4349]));
Q_ASSIGN U12042 ( .B(clk), .A(\g.we_clk [4348]));
Q_ASSIGN U12043 ( .B(clk), .A(\g.we_clk [4347]));
Q_ASSIGN U12044 ( .B(clk), .A(\g.we_clk [4346]));
Q_ASSIGN U12045 ( .B(clk), .A(\g.we_clk [4345]));
Q_ASSIGN U12046 ( .B(clk), .A(\g.we_clk [4344]));
Q_ASSIGN U12047 ( .B(clk), .A(\g.we_clk [4343]));
Q_ASSIGN U12048 ( .B(clk), .A(\g.we_clk [4342]));
Q_ASSIGN U12049 ( .B(clk), .A(\g.we_clk [4341]));
Q_ASSIGN U12050 ( .B(clk), .A(\g.we_clk [4340]));
Q_ASSIGN U12051 ( .B(clk), .A(\g.we_clk [4339]));
Q_ASSIGN U12052 ( .B(clk), .A(\g.we_clk [4338]));
Q_ASSIGN U12053 ( .B(clk), .A(\g.we_clk [4337]));
Q_ASSIGN U12054 ( .B(clk), .A(\g.we_clk [4336]));
Q_ASSIGN U12055 ( .B(clk), .A(\g.we_clk [4335]));
Q_ASSIGN U12056 ( .B(clk), .A(\g.we_clk [4334]));
Q_ASSIGN U12057 ( .B(clk), .A(\g.we_clk [4333]));
Q_ASSIGN U12058 ( .B(clk), .A(\g.we_clk [4332]));
Q_ASSIGN U12059 ( .B(clk), .A(\g.we_clk [4331]));
Q_ASSIGN U12060 ( .B(clk), .A(\g.we_clk [4330]));
Q_ASSIGN U12061 ( .B(clk), .A(\g.we_clk [4329]));
Q_ASSIGN U12062 ( .B(clk), .A(\g.we_clk [4328]));
Q_ASSIGN U12063 ( .B(clk), .A(\g.we_clk [4327]));
Q_ASSIGN U12064 ( .B(clk), .A(\g.we_clk [4326]));
Q_ASSIGN U12065 ( .B(clk), .A(\g.we_clk [4325]));
Q_ASSIGN U12066 ( .B(clk), .A(\g.we_clk [4324]));
Q_ASSIGN U12067 ( .B(clk), .A(\g.we_clk [4323]));
Q_ASSIGN U12068 ( .B(clk), .A(\g.we_clk [4322]));
Q_ASSIGN U12069 ( .B(clk), .A(\g.we_clk [4321]));
Q_ASSIGN U12070 ( .B(clk), .A(\g.we_clk [4320]));
Q_ASSIGN U12071 ( .B(clk), .A(\g.we_clk [4319]));
Q_ASSIGN U12072 ( .B(clk), .A(\g.we_clk [4318]));
Q_ASSIGN U12073 ( .B(clk), .A(\g.we_clk [4317]));
Q_ASSIGN U12074 ( .B(clk), .A(\g.we_clk [4316]));
Q_ASSIGN U12075 ( .B(clk), .A(\g.we_clk [4315]));
Q_ASSIGN U12076 ( .B(clk), .A(\g.we_clk [4314]));
Q_ASSIGN U12077 ( .B(clk), .A(\g.we_clk [4313]));
Q_ASSIGN U12078 ( .B(clk), .A(\g.we_clk [4312]));
Q_ASSIGN U12079 ( .B(clk), .A(\g.we_clk [4311]));
Q_ASSIGN U12080 ( .B(clk), .A(\g.we_clk [4310]));
Q_ASSIGN U12081 ( .B(clk), .A(\g.we_clk [4309]));
Q_ASSIGN U12082 ( .B(clk), .A(\g.we_clk [4308]));
Q_ASSIGN U12083 ( .B(clk), .A(\g.we_clk [4307]));
Q_ASSIGN U12084 ( .B(clk), .A(\g.we_clk [4306]));
Q_ASSIGN U12085 ( .B(clk), .A(\g.we_clk [4305]));
Q_ASSIGN U12086 ( .B(clk), .A(\g.we_clk [4304]));
Q_ASSIGN U12087 ( .B(clk), .A(\g.we_clk [4303]));
Q_ASSIGN U12088 ( .B(clk), .A(\g.we_clk [4302]));
Q_ASSIGN U12089 ( .B(clk), .A(\g.we_clk [4301]));
Q_ASSIGN U12090 ( .B(clk), .A(\g.we_clk [4300]));
Q_ASSIGN U12091 ( .B(clk), .A(\g.we_clk [4299]));
Q_ASSIGN U12092 ( .B(clk), .A(\g.we_clk [4298]));
Q_ASSIGN U12093 ( .B(clk), .A(\g.we_clk [4297]));
Q_ASSIGN U12094 ( .B(clk), .A(\g.we_clk [4296]));
Q_ASSIGN U12095 ( .B(clk), .A(\g.we_clk [4295]));
Q_ASSIGN U12096 ( .B(clk), .A(\g.we_clk [4294]));
Q_ASSIGN U12097 ( .B(clk), .A(\g.we_clk [4293]));
Q_ASSIGN U12098 ( .B(clk), .A(\g.we_clk [4292]));
Q_ASSIGN U12099 ( .B(clk), .A(\g.we_clk [4291]));
Q_ASSIGN U12100 ( .B(clk), .A(\g.we_clk [4290]));
Q_ASSIGN U12101 ( .B(clk), .A(\g.we_clk [4289]));
Q_ASSIGN U12102 ( .B(clk), .A(\g.we_clk [4288]));
Q_ASSIGN U12103 ( .B(clk), .A(\g.we_clk [4287]));
Q_ASSIGN U12104 ( .B(clk), .A(\g.we_clk [4286]));
Q_ASSIGN U12105 ( .B(clk), .A(\g.we_clk [4285]));
Q_ASSIGN U12106 ( .B(clk), .A(\g.we_clk [4284]));
Q_ASSIGN U12107 ( .B(clk), .A(\g.we_clk [4283]));
Q_ASSIGN U12108 ( .B(clk), .A(\g.we_clk [4282]));
Q_ASSIGN U12109 ( .B(clk), .A(\g.we_clk [4281]));
Q_ASSIGN U12110 ( .B(clk), .A(\g.we_clk [4280]));
Q_ASSIGN U12111 ( .B(clk), .A(\g.we_clk [4279]));
Q_ASSIGN U12112 ( .B(clk), .A(\g.we_clk [4278]));
Q_ASSIGN U12113 ( .B(clk), .A(\g.we_clk [4277]));
Q_ASSIGN U12114 ( .B(clk), .A(\g.we_clk [4276]));
Q_ASSIGN U12115 ( .B(clk), .A(\g.we_clk [4275]));
Q_ASSIGN U12116 ( .B(clk), .A(\g.we_clk [4274]));
Q_ASSIGN U12117 ( .B(clk), .A(\g.we_clk [4273]));
Q_ASSIGN U12118 ( .B(clk), .A(\g.we_clk [4272]));
Q_ASSIGN U12119 ( .B(clk), .A(\g.we_clk [4271]));
Q_ASSIGN U12120 ( .B(clk), .A(\g.we_clk [4270]));
Q_ASSIGN U12121 ( .B(clk), .A(\g.we_clk [4269]));
Q_ASSIGN U12122 ( .B(clk), .A(\g.we_clk [4268]));
Q_ASSIGN U12123 ( .B(clk), .A(\g.we_clk [4267]));
Q_ASSIGN U12124 ( .B(clk), .A(\g.we_clk [4266]));
Q_ASSIGN U12125 ( .B(clk), .A(\g.we_clk [4265]));
Q_ASSIGN U12126 ( .B(clk), .A(\g.we_clk [4264]));
Q_ASSIGN U12127 ( .B(clk), .A(\g.we_clk [4263]));
Q_ASSIGN U12128 ( .B(clk), .A(\g.we_clk [4262]));
Q_ASSIGN U12129 ( .B(clk), .A(\g.we_clk [4261]));
Q_ASSIGN U12130 ( .B(clk), .A(\g.we_clk [4260]));
Q_ASSIGN U12131 ( .B(clk), .A(\g.we_clk [4259]));
Q_ASSIGN U12132 ( .B(clk), .A(\g.we_clk [4258]));
Q_ASSIGN U12133 ( .B(clk), .A(\g.we_clk [4257]));
Q_ASSIGN U12134 ( .B(clk), .A(\g.we_clk [4256]));
Q_ASSIGN U12135 ( .B(clk), .A(\g.we_clk [4255]));
Q_ASSIGN U12136 ( .B(clk), .A(\g.we_clk [4254]));
Q_ASSIGN U12137 ( .B(clk), .A(\g.we_clk [4253]));
Q_ASSIGN U12138 ( .B(clk), .A(\g.we_clk [4252]));
Q_ASSIGN U12139 ( .B(clk), .A(\g.we_clk [4251]));
Q_ASSIGN U12140 ( .B(clk), .A(\g.we_clk [4250]));
Q_ASSIGN U12141 ( .B(clk), .A(\g.we_clk [4249]));
Q_ASSIGN U12142 ( .B(clk), .A(\g.we_clk [4248]));
Q_ASSIGN U12143 ( .B(clk), .A(\g.we_clk [4247]));
Q_ASSIGN U12144 ( .B(clk), .A(\g.we_clk [4246]));
Q_ASSIGN U12145 ( .B(clk), .A(\g.we_clk [4245]));
Q_ASSIGN U12146 ( .B(clk), .A(\g.we_clk [4244]));
Q_ASSIGN U12147 ( .B(clk), .A(\g.we_clk [4243]));
Q_ASSIGN U12148 ( .B(clk), .A(\g.we_clk [4242]));
Q_ASSIGN U12149 ( .B(clk), .A(\g.we_clk [4241]));
Q_ASSIGN U12150 ( .B(clk), .A(\g.we_clk [4240]));
Q_ASSIGN U12151 ( .B(clk), .A(\g.we_clk [4239]));
Q_ASSIGN U12152 ( .B(clk), .A(\g.we_clk [4238]));
Q_ASSIGN U12153 ( .B(clk), .A(\g.we_clk [4237]));
Q_ASSIGN U12154 ( .B(clk), .A(\g.we_clk [4236]));
Q_ASSIGN U12155 ( .B(clk), .A(\g.we_clk [4235]));
Q_ASSIGN U12156 ( .B(clk), .A(\g.we_clk [4234]));
Q_ASSIGN U12157 ( .B(clk), .A(\g.we_clk [4233]));
Q_ASSIGN U12158 ( .B(clk), .A(\g.we_clk [4232]));
Q_ASSIGN U12159 ( .B(clk), .A(\g.we_clk [4231]));
Q_ASSIGN U12160 ( .B(clk), .A(\g.we_clk [4230]));
Q_ASSIGN U12161 ( .B(clk), .A(\g.we_clk [4229]));
Q_ASSIGN U12162 ( .B(clk), .A(\g.we_clk [4228]));
Q_ASSIGN U12163 ( .B(clk), .A(\g.we_clk [4227]));
Q_ASSIGN U12164 ( .B(clk), .A(\g.we_clk [4226]));
Q_ASSIGN U12165 ( .B(clk), .A(\g.we_clk [4225]));
Q_ASSIGN U12166 ( .B(clk), .A(\g.we_clk [4224]));
Q_ASSIGN U12167 ( .B(clk), .A(\g.we_clk [4223]));
Q_ASSIGN U12168 ( .B(clk), .A(\g.we_clk [4222]));
Q_ASSIGN U12169 ( .B(clk), .A(\g.we_clk [4221]));
Q_ASSIGN U12170 ( .B(clk), .A(\g.we_clk [4220]));
Q_ASSIGN U12171 ( .B(clk), .A(\g.we_clk [4219]));
Q_ASSIGN U12172 ( .B(clk), .A(\g.we_clk [4218]));
Q_ASSIGN U12173 ( .B(clk), .A(\g.we_clk [4217]));
Q_ASSIGN U12174 ( .B(clk), .A(\g.we_clk [4216]));
Q_ASSIGN U12175 ( .B(clk), .A(\g.we_clk [4215]));
Q_ASSIGN U12176 ( .B(clk), .A(\g.we_clk [4214]));
Q_ASSIGN U12177 ( .B(clk), .A(\g.we_clk [4213]));
Q_ASSIGN U12178 ( .B(clk), .A(\g.we_clk [4212]));
Q_ASSIGN U12179 ( .B(clk), .A(\g.we_clk [4211]));
Q_ASSIGN U12180 ( .B(clk), .A(\g.we_clk [4210]));
Q_ASSIGN U12181 ( .B(clk), .A(\g.we_clk [4209]));
Q_ASSIGN U12182 ( .B(clk), .A(\g.we_clk [4208]));
Q_ASSIGN U12183 ( .B(clk), .A(\g.we_clk [4207]));
Q_ASSIGN U12184 ( .B(clk), .A(\g.we_clk [4206]));
Q_ASSIGN U12185 ( .B(clk), .A(\g.we_clk [4205]));
Q_ASSIGN U12186 ( .B(clk), .A(\g.we_clk [4204]));
Q_ASSIGN U12187 ( .B(clk), .A(\g.we_clk [4203]));
Q_ASSIGN U12188 ( .B(clk), .A(\g.we_clk [4202]));
Q_ASSIGN U12189 ( .B(clk), .A(\g.we_clk [4201]));
Q_ASSIGN U12190 ( .B(clk), .A(\g.we_clk [4200]));
Q_ASSIGN U12191 ( .B(clk), .A(\g.we_clk [4199]));
Q_ASSIGN U12192 ( .B(clk), .A(\g.we_clk [4198]));
Q_ASSIGN U12193 ( .B(clk), .A(\g.we_clk [4197]));
Q_ASSIGN U12194 ( .B(clk), .A(\g.we_clk [4196]));
Q_ASSIGN U12195 ( .B(clk), .A(\g.we_clk [4195]));
Q_ASSIGN U12196 ( .B(clk), .A(\g.we_clk [4194]));
Q_ASSIGN U12197 ( .B(clk), .A(\g.we_clk [4193]));
Q_ASSIGN U12198 ( .B(clk), .A(\g.we_clk [4192]));
Q_ASSIGN U12199 ( .B(clk), .A(\g.we_clk [4191]));
Q_ASSIGN U12200 ( .B(clk), .A(\g.we_clk [4190]));
Q_ASSIGN U12201 ( .B(clk), .A(\g.we_clk [4189]));
Q_ASSIGN U12202 ( .B(clk), .A(\g.we_clk [4188]));
Q_ASSIGN U12203 ( .B(clk), .A(\g.we_clk [4187]));
Q_ASSIGN U12204 ( .B(clk), .A(\g.we_clk [4186]));
Q_ASSIGN U12205 ( .B(clk), .A(\g.we_clk [4185]));
Q_ASSIGN U12206 ( .B(clk), .A(\g.we_clk [4184]));
Q_ASSIGN U12207 ( .B(clk), .A(\g.we_clk [4183]));
Q_ASSIGN U12208 ( .B(clk), .A(\g.we_clk [4182]));
Q_ASSIGN U12209 ( .B(clk), .A(\g.we_clk [4181]));
Q_ASSIGN U12210 ( .B(clk), .A(\g.we_clk [4180]));
Q_ASSIGN U12211 ( .B(clk), .A(\g.we_clk [4179]));
Q_ASSIGN U12212 ( .B(clk), .A(\g.we_clk [4178]));
Q_ASSIGN U12213 ( .B(clk), .A(\g.we_clk [4177]));
Q_ASSIGN U12214 ( .B(clk), .A(\g.we_clk [4176]));
Q_ASSIGN U12215 ( .B(clk), .A(\g.we_clk [4175]));
Q_ASSIGN U12216 ( .B(clk), .A(\g.we_clk [4174]));
Q_ASSIGN U12217 ( .B(clk), .A(\g.we_clk [4173]));
Q_ASSIGN U12218 ( .B(clk), .A(\g.we_clk [4172]));
Q_ASSIGN U12219 ( .B(clk), .A(\g.we_clk [4171]));
Q_ASSIGN U12220 ( .B(clk), .A(\g.we_clk [4170]));
Q_ASSIGN U12221 ( .B(clk), .A(\g.we_clk [4169]));
Q_ASSIGN U12222 ( .B(clk), .A(\g.we_clk [4168]));
Q_ASSIGN U12223 ( .B(clk), .A(\g.we_clk [4167]));
Q_ASSIGN U12224 ( .B(clk), .A(\g.we_clk [4166]));
Q_ASSIGN U12225 ( .B(clk), .A(\g.we_clk [4165]));
Q_ASSIGN U12226 ( .B(clk), .A(\g.we_clk [4164]));
Q_ASSIGN U12227 ( .B(clk), .A(\g.we_clk [4163]));
Q_ASSIGN U12228 ( .B(clk), .A(\g.we_clk [4162]));
Q_ASSIGN U12229 ( .B(clk), .A(\g.we_clk [4161]));
Q_ASSIGN U12230 ( .B(clk), .A(\g.we_clk [4160]));
Q_ASSIGN U12231 ( .B(clk), .A(\g.we_clk [4159]));
Q_ASSIGN U12232 ( .B(clk), .A(\g.we_clk [4158]));
Q_ASSIGN U12233 ( .B(clk), .A(\g.we_clk [4157]));
Q_ASSIGN U12234 ( .B(clk), .A(\g.we_clk [4156]));
Q_ASSIGN U12235 ( .B(clk), .A(\g.we_clk [4155]));
Q_ASSIGN U12236 ( .B(clk), .A(\g.we_clk [4154]));
Q_ASSIGN U12237 ( .B(clk), .A(\g.we_clk [4153]));
Q_ASSIGN U12238 ( .B(clk), .A(\g.we_clk [4152]));
Q_ASSIGN U12239 ( .B(clk), .A(\g.we_clk [4151]));
Q_ASSIGN U12240 ( .B(clk), .A(\g.we_clk [4150]));
Q_ASSIGN U12241 ( .B(clk), .A(\g.we_clk [4149]));
Q_ASSIGN U12242 ( .B(clk), .A(\g.we_clk [4148]));
Q_ASSIGN U12243 ( .B(clk), .A(\g.we_clk [4147]));
Q_ASSIGN U12244 ( .B(clk), .A(\g.we_clk [4146]));
Q_ASSIGN U12245 ( .B(clk), .A(\g.we_clk [4145]));
Q_ASSIGN U12246 ( .B(clk), .A(\g.we_clk [4144]));
Q_ASSIGN U12247 ( .B(clk), .A(\g.we_clk [4143]));
Q_ASSIGN U12248 ( .B(clk), .A(\g.we_clk [4142]));
Q_ASSIGN U12249 ( .B(clk), .A(\g.we_clk [4141]));
Q_ASSIGN U12250 ( .B(clk), .A(\g.we_clk [4140]));
Q_ASSIGN U12251 ( .B(clk), .A(\g.we_clk [4139]));
Q_ASSIGN U12252 ( .B(clk), .A(\g.we_clk [4138]));
Q_ASSIGN U12253 ( .B(clk), .A(\g.we_clk [4137]));
Q_ASSIGN U12254 ( .B(clk), .A(\g.we_clk [4136]));
Q_ASSIGN U12255 ( .B(clk), .A(\g.we_clk [4135]));
Q_ASSIGN U12256 ( .B(clk), .A(\g.we_clk [4134]));
Q_ASSIGN U12257 ( .B(clk), .A(\g.we_clk [4133]));
Q_ASSIGN U12258 ( .B(clk), .A(\g.we_clk [4132]));
Q_ASSIGN U12259 ( .B(clk), .A(\g.we_clk [4131]));
Q_ASSIGN U12260 ( .B(clk), .A(\g.we_clk [4130]));
Q_ASSIGN U12261 ( .B(clk), .A(\g.we_clk [4129]));
Q_ASSIGN U12262 ( .B(clk), .A(\g.we_clk [4128]));
Q_ASSIGN U12263 ( .B(clk), .A(\g.we_clk [4127]));
Q_ASSIGN U12264 ( .B(clk), .A(\g.we_clk [4126]));
Q_ASSIGN U12265 ( .B(clk), .A(\g.we_clk [4125]));
Q_ASSIGN U12266 ( .B(clk), .A(\g.we_clk [4124]));
Q_ASSIGN U12267 ( .B(clk), .A(\g.we_clk [4123]));
Q_ASSIGN U12268 ( .B(clk), .A(\g.we_clk [4122]));
Q_ASSIGN U12269 ( .B(clk), .A(\g.we_clk [4121]));
Q_ASSIGN U12270 ( .B(clk), .A(\g.we_clk [4120]));
Q_ASSIGN U12271 ( .B(clk), .A(\g.we_clk [4119]));
Q_ASSIGN U12272 ( .B(clk), .A(\g.we_clk [4118]));
Q_ASSIGN U12273 ( .B(clk), .A(\g.we_clk [4117]));
Q_ASSIGN U12274 ( .B(clk), .A(\g.we_clk [4116]));
Q_ASSIGN U12275 ( .B(clk), .A(\g.we_clk [4115]));
Q_ASSIGN U12276 ( .B(clk), .A(\g.we_clk [4114]));
Q_ASSIGN U12277 ( .B(clk), .A(\g.we_clk [4113]));
Q_ASSIGN U12278 ( .B(clk), .A(\g.we_clk [4112]));
Q_ASSIGN U12279 ( .B(clk), .A(\g.we_clk [4111]));
Q_ASSIGN U12280 ( .B(clk), .A(\g.we_clk [4110]));
Q_ASSIGN U12281 ( .B(clk), .A(\g.we_clk [4109]));
Q_ASSIGN U12282 ( .B(clk), .A(\g.we_clk [4108]));
Q_ASSIGN U12283 ( .B(clk), .A(\g.we_clk [4107]));
Q_ASSIGN U12284 ( .B(clk), .A(\g.we_clk [4106]));
Q_ASSIGN U12285 ( .B(clk), .A(\g.we_clk [4105]));
Q_ASSIGN U12286 ( .B(clk), .A(\g.we_clk [4104]));
Q_ASSIGN U12287 ( .B(clk), .A(\g.we_clk [4103]));
Q_ASSIGN U12288 ( .B(clk), .A(\g.we_clk [4102]));
Q_ASSIGN U12289 ( .B(clk), .A(\g.we_clk [4101]));
Q_ASSIGN U12290 ( .B(clk), .A(\g.we_clk [4100]));
Q_ASSIGN U12291 ( .B(clk), .A(\g.we_clk [4099]));
Q_ASSIGN U12292 ( .B(clk), .A(\g.we_clk [4098]));
Q_ASSIGN U12293 ( .B(clk), .A(\g.we_clk [4097]));
Q_ASSIGN U12294 ( .B(clk), .A(\g.we_clk [4096]));
Q_ASSIGN U12295 ( .B(clk), .A(\g.we_clk [4095]));
Q_ASSIGN U12296 ( .B(clk), .A(\g.we_clk [4094]));
Q_ASSIGN U12297 ( .B(clk), .A(\g.we_clk [4093]));
Q_ASSIGN U12298 ( .B(clk), .A(\g.we_clk [4092]));
Q_ASSIGN U12299 ( .B(clk), .A(\g.we_clk [4091]));
Q_ASSIGN U12300 ( .B(clk), .A(\g.we_clk [4090]));
Q_ASSIGN U12301 ( .B(clk), .A(\g.we_clk [4089]));
Q_ASSIGN U12302 ( .B(clk), .A(\g.we_clk [4088]));
Q_ASSIGN U12303 ( .B(clk), .A(\g.we_clk [4087]));
Q_ASSIGN U12304 ( .B(clk), .A(\g.we_clk [4086]));
Q_ASSIGN U12305 ( .B(clk), .A(\g.we_clk [4085]));
Q_ASSIGN U12306 ( .B(clk), .A(\g.we_clk [4084]));
Q_ASSIGN U12307 ( .B(clk), .A(\g.we_clk [4083]));
Q_ASSIGN U12308 ( .B(clk), .A(\g.we_clk [4082]));
Q_ASSIGN U12309 ( .B(clk), .A(\g.we_clk [4081]));
Q_ASSIGN U12310 ( .B(clk), .A(\g.we_clk [4080]));
Q_ASSIGN U12311 ( .B(clk), .A(\g.we_clk [4079]));
Q_ASSIGN U12312 ( .B(clk), .A(\g.we_clk [4078]));
Q_ASSIGN U12313 ( .B(clk), .A(\g.we_clk [4077]));
Q_ASSIGN U12314 ( .B(clk), .A(\g.we_clk [4076]));
Q_ASSIGN U12315 ( .B(clk), .A(\g.we_clk [4075]));
Q_ASSIGN U12316 ( .B(clk), .A(\g.we_clk [4074]));
Q_ASSIGN U12317 ( .B(clk), .A(\g.we_clk [4073]));
Q_ASSIGN U12318 ( .B(clk), .A(\g.we_clk [4072]));
Q_ASSIGN U12319 ( .B(clk), .A(\g.we_clk [4071]));
Q_ASSIGN U12320 ( .B(clk), .A(\g.we_clk [4070]));
Q_ASSIGN U12321 ( .B(clk), .A(\g.we_clk [4069]));
Q_ASSIGN U12322 ( .B(clk), .A(\g.we_clk [4068]));
Q_ASSIGN U12323 ( .B(clk), .A(\g.we_clk [4067]));
Q_ASSIGN U12324 ( .B(clk), .A(\g.we_clk [4066]));
Q_ASSIGN U12325 ( .B(clk), .A(\g.we_clk [4065]));
Q_ASSIGN U12326 ( .B(clk), .A(\g.we_clk [4064]));
Q_ASSIGN U12327 ( .B(clk), .A(\g.we_clk [4063]));
Q_ASSIGN U12328 ( .B(clk), .A(\g.we_clk [4062]));
Q_ASSIGN U12329 ( .B(clk), .A(\g.we_clk [4061]));
Q_ASSIGN U12330 ( .B(clk), .A(\g.we_clk [4060]));
Q_ASSIGN U12331 ( .B(clk), .A(\g.we_clk [4059]));
Q_ASSIGN U12332 ( .B(clk), .A(\g.we_clk [4058]));
Q_ASSIGN U12333 ( .B(clk), .A(\g.we_clk [4057]));
Q_ASSIGN U12334 ( .B(clk), .A(\g.we_clk [4056]));
Q_ASSIGN U12335 ( .B(clk), .A(\g.we_clk [4055]));
Q_ASSIGN U12336 ( .B(clk), .A(\g.we_clk [4054]));
Q_ASSIGN U12337 ( .B(clk), .A(\g.we_clk [4053]));
Q_ASSIGN U12338 ( .B(clk), .A(\g.we_clk [4052]));
Q_ASSIGN U12339 ( .B(clk), .A(\g.we_clk [4051]));
Q_ASSIGN U12340 ( .B(clk), .A(\g.we_clk [4050]));
Q_ASSIGN U12341 ( .B(clk), .A(\g.we_clk [4049]));
Q_ASSIGN U12342 ( .B(clk), .A(\g.we_clk [4048]));
Q_ASSIGN U12343 ( .B(clk), .A(\g.we_clk [4047]));
Q_ASSIGN U12344 ( .B(clk), .A(\g.we_clk [4046]));
Q_ASSIGN U12345 ( .B(clk), .A(\g.we_clk [4045]));
Q_ASSIGN U12346 ( .B(clk), .A(\g.we_clk [4044]));
Q_ASSIGN U12347 ( .B(clk), .A(\g.we_clk [4043]));
Q_ASSIGN U12348 ( .B(clk), .A(\g.we_clk [4042]));
Q_ASSIGN U12349 ( .B(clk), .A(\g.we_clk [4041]));
Q_ASSIGN U12350 ( .B(clk), .A(\g.we_clk [4040]));
Q_ASSIGN U12351 ( .B(clk), .A(\g.we_clk [4039]));
Q_ASSIGN U12352 ( .B(clk), .A(\g.we_clk [4038]));
Q_ASSIGN U12353 ( .B(clk), .A(\g.we_clk [4037]));
Q_ASSIGN U12354 ( .B(clk), .A(\g.we_clk [4036]));
Q_ASSIGN U12355 ( .B(clk), .A(\g.we_clk [4035]));
Q_ASSIGN U12356 ( .B(clk), .A(\g.we_clk [4034]));
Q_ASSIGN U12357 ( .B(clk), .A(\g.we_clk [4033]));
Q_ASSIGN U12358 ( .B(clk), .A(\g.we_clk [4032]));
Q_ASSIGN U12359 ( .B(clk), .A(\g.we_clk [4031]));
Q_ASSIGN U12360 ( .B(clk), .A(\g.we_clk [4030]));
Q_ASSIGN U12361 ( .B(clk), .A(\g.we_clk [4029]));
Q_ASSIGN U12362 ( .B(clk), .A(\g.we_clk [4028]));
Q_ASSIGN U12363 ( .B(clk), .A(\g.we_clk [4027]));
Q_ASSIGN U12364 ( .B(clk), .A(\g.we_clk [4026]));
Q_ASSIGN U12365 ( .B(clk), .A(\g.we_clk [4025]));
Q_ASSIGN U12366 ( .B(clk), .A(\g.we_clk [4024]));
Q_ASSIGN U12367 ( .B(clk), .A(\g.we_clk [4023]));
Q_ASSIGN U12368 ( .B(clk), .A(\g.we_clk [4022]));
Q_ASSIGN U12369 ( .B(clk), .A(\g.we_clk [4021]));
Q_ASSIGN U12370 ( .B(clk), .A(\g.we_clk [4020]));
Q_ASSIGN U12371 ( .B(clk), .A(\g.we_clk [4019]));
Q_ASSIGN U12372 ( .B(clk), .A(\g.we_clk [4018]));
Q_ASSIGN U12373 ( .B(clk), .A(\g.we_clk [4017]));
Q_ASSIGN U12374 ( .B(clk), .A(\g.we_clk [4016]));
Q_ASSIGN U12375 ( .B(clk), .A(\g.we_clk [4015]));
Q_ASSIGN U12376 ( .B(clk), .A(\g.we_clk [4014]));
Q_ASSIGN U12377 ( .B(clk), .A(\g.we_clk [4013]));
Q_ASSIGN U12378 ( .B(clk), .A(\g.we_clk [4012]));
Q_ASSIGN U12379 ( .B(clk), .A(\g.we_clk [4011]));
Q_ASSIGN U12380 ( .B(clk), .A(\g.we_clk [4010]));
Q_ASSIGN U12381 ( .B(clk), .A(\g.we_clk [4009]));
Q_ASSIGN U12382 ( .B(clk), .A(\g.we_clk [4008]));
Q_ASSIGN U12383 ( .B(clk), .A(\g.we_clk [4007]));
Q_ASSIGN U12384 ( .B(clk), .A(\g.we_clk [4006]));
Q_ASSIGN U12385 ( .B(clk), .A(\g.we_clk [4005]));
Q_ASSIGN U12386 ( .B(clk), .A(\g.we_clk [4004]));
Q_ASSIGN U12387 ( .B(clk), .A(\g.we_clk [4003]));
Q_ASSIGN U12388 ( .B(clk), .A(\g.we_clk [4002]));
Q_ASSIGN U12389 ( .B(clk), .A(\g.we_clk [4001]));
Q_ASSIGN U12390 ( .B(clk), .A(\g.we_clk [4000]));
Q_ASSIGN U12391 ( .B(clk), .A(\g.we_clk [3999]));
Q_ASSIGN U12392 ( .B(clk), .A(\g.we_clk [3998]));
Q_ASSIGN U12393 ( .B(clk), .A(\g.we_clk [3997]));
Q_ASSIGN U12394 ( .B(clk), .A(\g.we_clk [3996]));
Q_ASSIGN U12395 ( .B(clk), .A(\g.we_clk [3995]));
Q_ASSIGN U12396 ( .B(clk), .A(\g.we_clk [3994]));
Q_ASSIGN U12397 ( .B(clk), .A(\g.we_clk [3993]));
Q_ASSIGN U12398 ( .B(clk), .A(\g.we_clk [3992]));
Q_ASSIGN U12399 ( .B(clk), .A(\g.we_clk [3991]));
Q_ASSIGN U12400 ( .B(clk), .A(\g.we_clk [3990]));
Q_ASSIGN U12401 ( .B(clk), .A(\g.we_clk [3989]));
Q_ASSIGN U12402 ( .B(clk), .A(\g.we_clk [3988]));
Q_ASSIGN U12403 ( .B(clk), .A(\g.we_clk [3987]));
Q_ASSIGN U12404 ( .B(clk), .A(\g.we_clk [3986]));
Q_ASSIGN U12405 ( .B(clk), .A(\g.we_clk [3985]));
Q_ASSIGN U12406 ( .B(clk), .A(\g.we_clk [3984]));
Q_ASSIGN U12407 ( .B(clk), .A(\g.we_clk [3983]));
Q_ASSIGN U12408 ( .B(clk), .A(\g.we_clk [3982]));
Q_ASSIGN U12409 ( .B(clk), .A(\g.we_clk [3981]));
Q_ASSIGN U12410 ( .B(clk), .A(\g.we_clk [3980]));
Q_ASSIGN U12411 ( .B(clk), .A(\g.we_clk [3979]));
Q_ASSIGN U12412 ( .B(clk), .A(\g.we_clk [3978]));
Q_ASSIGN U12413 ( .B(clk), .A(\g.we_clk [3977]));
Q_ASSIGN U12414 ( .B(clk), .A(\g.we_clk [3976]));
Q_ASSIGN U12415 ( .B(clk), .A(\g.we_clk [3975]));
Q_ASSIGN U12416 ( .B(clk), .A(\g.we_clk [3974]));
Q_ASSIGN U12417 ( .B(clk), .A(\g.we_clk [3973]));
Q_ASSIGN U12418 ( .B(clk), .A(\g.we_clk [3972]));
Q_ASSIGN U12419 ( .B(clk), .A(\g.we_clk [3971]));
Q_ASSIGN U12420 ( .B(clk), .A(\g.we_clk [3970]));
Q_ASSIGN U12421 ( .B(clk), .A(\g.we_clk [3969]));
Q_ASSIGN U12422 ( .B(clk), .A(\g.we_clk [3968]));
Q_ASSIGN U12423 ( .B(clk), .A(\g.we_clk [3967]));
Q_ASSIGN U12424 ( .B(clk), .A(\g.we_clk [3966]));
Q_ASSIGN U12425 ( .B(clk), .A(\g.we_clk [3965]));
Q_ASSIGN U12426 ( .B(clk), .A(\g.we_clk [3964]));
Q_ASSIGN U12427 ( .B(clk), .A(\g.we_clk [3963]));
Q_ASSIGN U12428 ( .B(clk), .A(\g.we_clk [3962]));
Q_ASSIGN U12429 ( .B(clk), .A(\g.we_clk [3961]));
Q_ASSIGN U12430 ( .B(clk), .A(\g.we_clk [3960]));
Q_ASSIGN U12431 ( .B(clk), .A(\g.we_clk [3959]));
Q_ASSIGN U12432 ( .B(clk), .A(\g.we_clk [3958]));
Q_ASSIGN U12433 ( .B(clk), .A(\g.we_clk [3957]));
Q_ASSIGN U12434 ( .B(clk), .A(\g.we_clk [3956]));
Q_ASSIGN U12435 ( .B(clk), .A(\g.we_clk [3955]));
Q_ASSIGN U12436 ( .B(clk), .A(\g.we_clk [3954]));
Q_ASSIGN U12437 ( .B(clk), .A(\g.we_clk [3953]));
Q_ASSIGN U12438 ( .B(clk), .A(\g.we_clk [3952]));
Q_ASSIGN U12439 ( .B(clk), .A(\g.we_clk [3951]));
Q_ASSIGN U12440 ( .B(clk), .A(\g.we_clk [3950]));
Q_ASSIGN U12441 ( .B(clk), .A(\g.we_clk [3949]));
Q_ASSIGN U12442 ( .B(clk), .A(\g.we_clk [3948]));
Q_ASSIGN U12443 ( .B(clk), .A(\g.we_clk [3947]));
Q_ASSIGN U12444 ( .B(clk), .A(\g.we_clk [3946]));
Q_ASSIGN U12445 ( .B(clk), .A(\g.we_clk [3945]));
Q_ASSIGN U12446 ( .B(clk), .A(\g.we_clk [3944]));
Q_ASSIGN U12447 ( .B(clk), .A(\g.we_clk [3943]));
Q_ASSIGN U12448 ( .B(clk), .A(\g.we_clk [3942]));
Q_ASSIGN U12449 ( .B(clk), .A(\g.we_clk [3941]));
Q_ASSIGN U12450 ( .B(clk), .A(\g.we_clk [3940]));
Q_ASSIGN U12451 ( .B(clk), .A(\g.we_clk [3939]));
Q_ASSIGN U12452 ( .B(clk), .A(\g.we_clk [3938]));
Q_ASSIGN U12453 ( .B(clk), .A(\g.we_clk [3937]));
Q_ASSIGN U12454 ( .B(clk), .A(\g.we_clk [3936]));
Q_ASSIGN U12455 ( .B(clk), .A(\g.we_clk [3935]));
Q_ASSIGN U12456 ( .B(clk), .A(\g.we_clk [3934]));
Q_ASSIGN U12457 ( .B(clk), .A(\g.we_clk [3933]));
Q_ASSIGN U12458 ( .B(clk), .A(\g.we_clk [3932]));
Q_ASSIGN U12459 ( .B(clk), .A(\g.we_clk [3931]));
Q_ASSIGN U12460 ( .B(clk), .A(\g.we_clk [3930]));
Q_ASSIGN U12461 ( .B(clk), .A(\g.we_clk [3929]));
Q_ASSIGN U12462 ( .B(clk), .A(\g.we_clk [3928]));
Q_ASSIGN U12463 ( .B(clk), .A(\g.we_clk [3927]));
Q_ASSIGN U12464 ( .B(clk), .A(\g.we_clk [3926]));
Q_ASSIGN U12465 ( .B(clk), .A(\g.we_clk [3925]));
Q_ASSIGN U12466 ( .B(clk), .A(\g.we_clk [3924]));
Q_ASSIGN U12467 ( .B(clk), .A(\g.we_clk [3923]));
Q_ASSIGN U12468 ( .B(clk), .A(\g.we_clk [3922]));
Q_ASSIGN U12469 ( .B(clk), .A(\g.we_clk [3921]));
Q_ASSIGN U12470 ( .B(clk), .A(\g.we_clk [3920]));
Q_ASSIGN U12471 ( .B(clk), .A(\g.we_clk [3919]));
Q_ASSIGN U12472 ( .B(clk), .A(\g.we_clk [3918]));
Q_ASSIGN U12473 ( .B(clk), .A(\g.we_clk [3917]));
Q_ASSIGN U12474 ( .B(clk), .A(\g.we_clk [3916]));
Q_ASSIGN U12475 ( .B(clk), .A(\g.we_clk [3915]));
Q_ASSIGN U12476 ( .B(clk), .A(\g.we_clk [3914]));
Q_ASSIGN U12477 ( .B(clk), .A(\g.we_clk [3913]));
Q_ASSIGN U12478 ( .B(clk), .A(\g.we_clk [3912]));
Q_ASSIGN U12479 ( .B(clk), .A(\g.we_clk [3911]));
Q_ASSIGN U12480 ( .B(clk), .A(\g.we_clk [3910]));
Q_ASSIGN U12481 ( .B(clk), .A(\g.we_clk [3909]));
Q_ASSIGN U12482 ( .B(clk), .A(\g.we_clk [3908]));
Q_ASSIGN U12483 ( .B(clk), .A(\g.we_clk [3907]));
Q_ASSIGN U12484 ( .B(clk), .A(\g.we_clk [3906]));
Q_ASSIGN U12485 ( .B(clk), .A(\g.we_clk [3905]));
Q_ASSIGN U12486 ( .B(clk), .A(\g.we_clk [3904]));
Q_ASSIGN U12487 ( .B(clk), .A(\g.we_clk [3903]));
Q_ASSIGN U12488 ( .B(clk), .A(\g.we_clk [3902]));
Q_ASSIGN U12489 ( .B(clk), .A(\g.we_clk [3901]));
Q_ASSIGN U12490 ( .B(clk), .A(\g.we_clk [3900]));
Q_ASSIGN U12491 ( .B(clk), .A(\g.we_clk [3899]));
Q_ASSIGN U12492 ( .B(clk), .A(\g.we_clk [3898]));
Q_ASSIGN U12493 ( .B(clk), .A(\g.we_clk [3897]));
Q_ASSIGN U12494 ( .B(clk), .A(\g.we_clk [3896]));
Q_ASSIGN U12495 ( .B(clk), .A(\g.we_clk [3895]));
Q_ASSIGN U12496 ( .B(clk), .A(\g.we_clk [3894]));
Q_ASSIGN U12497 ( .B(clk), .A(\g.we_clk [3893]));
Q_ASSIGN U12498 ( .B(clk), .A(\g.we_clk [3892]));
Q_ASSIGN U12499 ( .B(clk), .A(\g.we_clk [3891]));
Q_ASSIGN U12500 ( .B(clk), .A(\g.we_clk [3890]));
Q_ASSIGN U12501 ( .B(clk), .A(\g.we_clk [3889]));
Q_ASSIGN U12502 ( .B(clk), .A(\g.we_clk [3888]));
Q_ASSIGN U12503 ( .B(clk), .A(\g.we_clk [3887]));
Q_ASSIGN U12504 ( .B(clk), .A(\g.we_clk [3886]));
Q_ASSIGN U12505 ( .B(clk), .A(\g.we_clk [3885]));
Q_ASSIGN U12506 ( .B(clk), .A(\g.we_clk [3884]));
Q_ASSIGN U12507 ( .B(clk), .A(\g.we_clk [3883]));
Q_ASSIGN U12508 ( .B(clk), .A(\g.we_clk [3882]));
Q_ASSIGN U12509 ( .B(clk), .A(\g.we_clk [3881]));
Q_ASSIGN U12510 ( .B(clk), .A(\g.we_clk [3880]));
Q_ASSIGN U12511 ( .B(clk), .A(\g.we_clk [3879]));
Q_ASSIGN U12512 ( .B(clk), .A(\g.we_clk [3878]));
Q_ASSIGN U12513 ( .B(clk), .A(\g.we_clk [3877]));
Q_ASSIGN U12514 ( .B(clk), .A(\g.we_clk [3876]));
Q_ASSIGN U12515 ( .B(clk), .A(\g.we_clk [3875]));
Q_ASSIGN U12516 ( .B(clk), .A(\g.we_clk [3874]));
Q_ASSIGN U12517 ( .B(clk), .A(\g.we_clk [3873]));
Q_ASSIGN U12518 ( .B(clk), .A(\g.we_clk [3872]));
Q_ASSIGN U12519 ( .B(clk), .A(\g.we_clk [3871]));
Q_ASSIGN U12520 ( .B(clk), .A(\g.we_clk [3870]));
Q_ASSIGN U12521 ( .B(clk), .A(\g.we_clk [3869]));
Q_ASSIGN U12522 ( .B(clk), .A(\g.we_clk [3868]));
Q_ASSIGN U12523 ( .B(clk), .A(\g.we_clk [3867]));
Q_ASSIGN U12524 ( .B(clk), .A(\g.we_clk [3866]));
Q_ASSIGN U12525 ( .B(clk), .A(\g.we_clk [3865]));
Q_ASSIGN U12526 ( .B(clk), .A(\g.we_clk [3864]));
Q_ASSIGN U12527 ( .B(clk), .A(\g.we_clk [3863]));
Q_ASSIGN U12528 ( .B(clk), .A(\g.we_clk [3862]));
Q_ASSIGN U12529 ( .B(clk), .A(\g.we_clk [3861]));
Q_ASSIGN U12530 ( .B(clk), .A(\g.we_clk [3860]));
Q_ASSIGN U12531 ( .B(clk), .A(\g.we_clk [3859]));
Q_ASSIGN U12532 ( .B(clk), .A(\g.we_clk [3858]));
Q_ASSIGN U12533 ( .B(clk), .A(\g.we_clk [3857]));
Q_ASSIGN U12534 ( .B(clk), .A(\g.we_clk [3856]));
Q_ASSIGN U12535 ( .B(clk), .A(\g.we_clk [3855]));
Q_ASSIGN U12536 ( .B(clk), .A(\g.we_clk [3854]));
Q_ASSIGN U12537 ( .B(clk), .A(\g.we_clk [3853]));
Q_ASSIGN U12538 ( .B(clk), .A(\g.we_clk [3852]));
Q_ASSIGN U12539 ( .B(clk), .A(\g.we_clk [3851]));
Q_ASSIGN U12540 ( .B(clk), .A(\g.we_clk [3850]));
Q_ASSIGN U12541 ( .B(clk), .A(\g.we_clk [3849]));
Q_ASSIGN U12542 ( .B(clk), .A(\g.we_clk [3848]));
Q_ASSIGN U12543 ( .B(clk), .A(\g.we_clk [3847]));
Q_ASSIGN U12544 ( .B(clk), .A(\g.we_clk [3846]));
Q_ASSIGN U12545 ( .B(clk), .A(\g.we_clk [3845]));
Q_ASSIGN U12546 ( .B(clk), .A(\g.we_clk [3844]));
Q_ASSIGN U12547 ( .B(clk), .A(\g.we_clk [3843]));
Q_ASSIGN U12548 ( .B(clk), .A(\g.we_clk [3842]));
Q_ASSIGN U12549 ( .B(clk), .A(\g.we_clk [3841]));
Q_ASSIGN U12550 ( .B(clk), .A(\g.we_clk [3840]));
Q_ASSIGN U12551 ( .B(clk), .A(\g.we_clk [3839]));
Q_ASSIGN U12552 ( .B(clk), .A(\g.we_clk [3838]));
Q_ASSIGN U12553 ( .B(clk), .A(\g.we_clk [3837]));
Q_ASSIGN U12554 ( .B(clk), .A(\g.we_clk [3836]));
Q_ASSIGN U12555 ( .B(clk), .A(\g.we_clk [3835]));
Q_ASSIGN U12556 ( .B(clk), .A(\g.we_clk [3834]));
Q_ASSIGN U12557 ( .B(clk), .A(\g.we_clk [3833]));
Q_ASSIGN U12558 ( .B(clk), .A(\g.we_clk [3832]));
Q_ASSIGN U12559 ( .B(clk), .A(\g.we_clk [3831]));
Q_ASSIGN U12560 ( .B(clk), .A(\g.we_clk [3830]));
Q_ASSIGN U12561 ( .B(clk), .A(\g.we_clk [3829]));
Q_ASSIGN U12562 ( .B(clk), .A(\g.we_clk [3828]));
Q_ASSIGN U12563 ( .B(clk), .A(\g.we_clk [3827]));
Q_ASSIGN U12564 ( .B(clk), .A(\g.we_clk [3826]));
Q_ASSIGN U12565 ( .B(clk), .A(\g.we_clk [3825]));
Q_ASSIGN U12566 ( .B(clk), .A(\g.we_clk [3824]));
Q_ASSIGN U12567 ( .B(clk), .A(\g.we_clk [3823]));
Q_ASSIGN U12568 ( .B(clk), .A(\g.we_clk [3822]));
Q_ASSIGN U12569 ( .B(clk), .A(\g.we_clk [3821]));
Q_ASSIGN U12570 ( .B(clk), .A(\g.we_clk [3820]));
Q_ASSIGN U12571 ( .B(clk), .A(\g.we_clk [3819]));
Q_ASSIGN U12572 ( .B(clk), .A(\g.we_clk [3818]));
Q_ASSIGN U12573 ( .B(clk), .A(\g.we_clk [3817]));
Q_ASSIGN U12574 ( .B(clk), .A(\g.we_clk [3816]));
Q_ASSIGN U12575 ( .B(clk), .A(\g.we_clk [3815]));
Q_ASSIGN U12576 ( .B(clk), .A(\g.we_clk [3814]));
Q_ASSIGN U12577 ( .B(clk), .A(\g.we_clk [3813]));
Q_ASSIGN U12578 ( .B(clk), .A(\g.we_clk [3812]));
Q_ASSIGN U12579 ( .B(clk), .A(\g.we_clk [3811]));
Q_ASSIGN U12580 ( .B(clk), .A(\g.we_clk [3810]));
Q_ASSIGN U12581 ( .B(clk), .A(\g.we_clk [3809]));
Q_ASSIGN U12582 ( .B(clk), .A(\g.we_clk [3808]));
Q_ASSIGN U12583 ( .B(clk), .A(\g.we_clk [3807]));
Q_ASSIGN U12584 ( .B(clk), .A(\g.we_clk [3806]));
Q_ASSIGN U12585 ( .B(clk), .A(\g.we_clk [3805]));
Q_ASSIGN U12586 ( .B(clk), .A(\g.we_clk [3804]));
Q_ASSIGN U12587 ( .B(clk), .A(\g.we_clk [3803]));
Q_ASSIGN U12588 ( .B(clk), .A(\g.we_clk [3802]));
Q_ASSIGN U12589 ( .B(clk), .A(\g.we_clk [3801]));
Q_ASSIGN U12590 ( .B(clk), .A(\g.we_clk [3800]));
Q_ASSIGN U12591 ( .B(clk), .A(\g.we_clk [3799]));
Q_ASSIGN U12592 ( .B(clk), .A(\g.we_clk [3798]));
Q_ASSIGN U12593 ( .B(clk), .A(\g.we_clk [3797]));
Q_ASSIGN U12594 ( .B(clk), .A(\g.we_clk [3796]));
Q_ASSIGN U12595 ( .B(clk), .A(\g.we_clk [3795]));
Q_ASSIGN U12596 ( .B(clk), .A(\g.we_clk [3794]));
Q_ASSIGN U12597 ( .B(clk), .A(\g.we_clk [3793]));
Q_ASSIGN U12598 ( .B(clk), .A(\g.we_clk [3792]));
Q_ASSIGN U12599 ( .B(clk), .A(\g.we_clk [3791]));
Q_ASSIGN U12600 ( .B(clk), .A(\g.we_clk [3790]));
Q_ASSIGN U12601 ( .B(clk), .A(\g.we_clk [3789]));
Q_ASSIGN U12602 ( .B(clk), .A(\g.we_clk [3788]));
Q_ASSIGN U12603 ( .B(clk), .A(\g.we_clk [3787]));
Q_ASSIGN U12604 ( .B(clk), .A(\g.we_clk [3786]));
Q_ASSIGN U12605 ( .B(clk), .A(\g.we_clk [3785]));
Q_ASSIGN U12606 ( .B(clk), .A(\g.we_clk [3784]));
Q_ASSIGN U12607 ( .B(clk), .A(\g.we_clk [3783]));
Q_ASSIGN U12608 ( .B(clk), .A(\g.we_clk [3782]));
Q_ASSIGN U12609 ( .B(clk), .A(\g.we_clk [3781]));
Q_ASSIGN U12610 ( .B(clk), .A(\g.we_clk [3780]));
Q_ASSIGN U12611 ( .B(clk), .A(\g.we_clk [3779]));
Q_ASSIGN U12612 ( .B(clk), .A(\g.we_clk [3778]));
Q_ASSIGN U12613 ( .B(clk), .A(\g.we_clk [3777]));
Q_ASSIGN U12614 ( .B(clk), .A(\g.we_clk [3776]));
Q_ASSIGN U12615 ( .B(clk), .A(\g.we_clk [3775]));
Q_ASSIGN U12616 ( .B(clk), .A(\g.we_clk [3774]));
Q_ASSIGN U12617 ( .B(clk), .A(\g.we_clk [3773]));
Q_ASSIGN U12618 ( .B(clk), .A(\g.we_clk [3772]));
Q_ASSIGN U12619 ( .B(clk), .A(\g.we_clk [3771]));
Q_ASSIGN U12620 ( .B(clk), .A(\g.we_clk [3770]));
Q_ASSIGN U12621 ( .B(clk), .A(\g.we_clk [3769]));
Q_ASSIGN U12622 ( .B(clk), .A(\g.we_clk [3768]));
Q_ASSIGN U12623 ( .B(clk), .A(\g.we_clk [3767]));
Q_ASSIGN U12624 ( .B(clk), .A(\g.we_clk [3766]));
Q_ASSIGN U12625 ( .B(clk), .A(\g.we_clk [3765]));
Q_ASSIGN U12626 ( .B(clk), .A(\g.we_clk [3764]));
Q_ASSIGN U12627 ( .B(clk), .A(\g.we_clk [3763]));
Q_ASSIGN U12628 ( .B(clk), .A(\g.we_clk [3762]));
Q_ASSIGN U12629 ( .B(clk), .A(\g.we_clk [3761]));
Q_ASSIGN U12630 ( .B(clk), .A(\g.we_clk [3760]));
Q_ASSIGN U12631 ( .B(clk), .A(\g.we_clk [3759]));
Q_ASSIGN U12632 ( .B(clk), .A(\g.we_clk [3758]));
Q_ASSIGN U12633 ( .B(clk), .A(\g.we_clk [3757]));
Q_ASSIGN U12634 ( .B(clk), .A(\g.we_clk [3756]));
Q_ASSIGN U12635 ( .B(clk), .A(\g.we_clk [3755]));
Q_ASSIGN U12636 ( .B(clk), .A(\g.we_clk [3754]));
Q_ASSIGN U12637 ( .B(clk), .A(\g.we_clk [3753]));
Q_ASSIGN U12638 ( .B(clk), .A(\g.we_clk [3752]));
Q_ASSIGN U12639 ( .B(clk), .A(\g.we_clk [3751]));
Q_ASSIGN U12640 ( .B(clk), .A(\g.we_clk [3750]));
Q_ASSIGN U12641 ( .B(clk), .A(\g.we_clk [3749]));
Q_ASSIGN U12642 ( .B(clk), .A(\g.we_clk [3748]));
Q_ASSIGN U12643 ( .B(clk), .A(\g.we_clk [3747]));
Q_ASSIGN U12644 ( .B(clk), .A(\g.we_clk [3746]));
Q_ASSIGN U12645 ( .B(clk), .A(\g.we_clk [3745]));
Q_ASSIGN U12646 ( .B(clk), .A(\g.we_clk [3744]));
Q_ASSIGN U12647 ( .B(clk), .A(\g.we_clk [3743]));
Q_ASSIGN U12648 ( .B(clk), .A(\g.we_clk [3742]));
Q_ASSIGN U12649 ( .B(clk), .A(\g.we_clk [3741]));
Q_ASSIGN U12650 ( .B(clk), .A(\g.we_clk [3740]));
Q_ASSIGN U12651 ( .B(clk), .A(\g.we_clk [3739]));
Q_ASSIGN U12652 ( .B(clk), .A(\g.we_clk [3738]));
Q_ASSIGN U12653 ( .B(clk), .A(\g.we_clk [3737]));
Q_ASSIGN U12654 ( .B(clk), .A(\g.we_clk [3736]));
Q_ASSIGN U12655 ( .B(clk), .A(\g.we_clk [3735]));
Q_ASSIGN U12656 ( .B(clk), .A(\g.we_clk [3734]));
Q_ASSIGN U12657 ( .B(clk), .A(\g.we_clk [3733]));
Q_ASSIGN U12658 ( .B(clk), .A(\g.we_clk [3732]));
Q_ASSIGN U12659 ( .B(clk), .A(\g.we_clk [3731]));
Q_ASSIGN U12660 ( .B(clk), .A(\g.we_clk [3730]));
Q_ASSIGN U12661 ( .B(clk), .A(\g.we_clk [3729]));
Q_ASSIGN U12662 ( .B(clk), .A(\g.we_clk [3728]));
Q_ASSIGN U12663 ( .B(clk), .A(\g.we_clk [3727]));
Q_ASSIGN U12664 ( .B(clk), .A(\g.we_clk [3726]));
Q_ASSIGN U12665 ( .B(clk), .A(\g.we_clk [3725]));
Q_ASSIGN U12666 ( .B(clk), .A(\g.we_clk [3724]));
Q_ASSIGN U12667 ( .B(clk), .A(\g.we_clk [3723]));
Q_ASSIGN U12668 ( .B(clk), .A(\g.we_clk [3722]));
Q_ASSIGN U12669 ( .B(clk), .A(\g.we_clk [3721]));
Q_ASSIGN U12670 ( .B(clk), .A(\g.we_clk [3720]));
Q_ASSIGN U12671 ( .B(clk), .A(\g.we_clk [3719]));
Q_ASSIGN U12672 ( .B(clk), .A(\g.we_clk [3718]));
Q_ASSIGN U12673 ( .B(clk), .A(\g.we_clk [3717]));
Q_ASSIGN U12674 ( .B(clk), .A(\g.we_clk [3716]));
Q_ASSIGN U12675 ( .B(clk), .A(\g.we_clk [3715]));
Q_ASSIGN U12676 ( .B(clk), .A(\g.we_clk [3714]));
Q_ASSIGN U12677 ( .B(clk), .A(\g.we_clk [3713]));
Q_ASSIGN U12678 ( .B(clk), .A(\g.we_clk [3712]));
Q_ASSIGN U12679 ( .B(clk), .A(\g.we_clk [3711]));
Q_ASSIGN U12680 ( .B(clk), .A(\g.we_clk [3710]));
Q_ASSIGN U12681 ( .B(clk), .A(\g.we_clk [3709]));
Q_ASSIGN U12682 ( .B(clk), .A(\g.we_clk [3708]));
Q_ASSIGN U12683 ( .B(clk), .A(\g.we_clk [3707]));
Q_ASSIGN U12684 ( .B(clk), .A(\g.we_clk [3706]));
Q_ASSIGN U12685 ( .B(clk), .A(\g.we_clk [3705]));
Q_ASSIGN U12686 ( .B(clk), .A(\g.we_clk [3704]));
Q_ASSIGN U12687 ( .B(clk), .A(\g.we_clk [3703]));
Q_ASSIGN U12688 ( .B(clk), .A(\g.we_clk [3702]));
Q_ASSIGN U12689 ( .B(clk), .A(\g.we_clk [3701]));
Q_ASSIGN U12690 ( .B(clk), .A(\g.we_clk [3700]));
Q_ASSIGN U12691 ( .B(clk), .A(\g.we_clk [3699]));
Q_ASSIGN U12692 ( .B(clk), .A(\g.we_clk [3698]));
Q_ASSIGN U12693 ( .B(clk), .A(\g.we_clk [3697]));
Q_ASSIGN U12694 ( .B(clk), .A(\g.we_clk [3696]));
Q_ASSIGN U12695 ( .B(clk), .A(\g.we_clk [3695]));
Q_ASSIGN U12696 ( .B(clk), .A(\g.we_clk [3694]));
Q_ASSIGN U12697 ( .B(clk), .A(\g.we_clk [3693]));
Q_ASSIGN U12698 ( .B(clk), .A(\g.we_clk [3692]));
Q_ASSIGN U12699 ( .B(clk), .A(\g.we_clk [3691]));
Q_ASSIGN U12700 ( .B(clk), .A(\g.we_clk [3690]));
Q_ASSIGN U12701 ( .B(clk), .A(\g.we_clk [3689]));
Q_ASSIGN U12702 ( .B(clk), .A(\g.we_clk [3688]));
Q_ASSIGN U12703 ( .B(clk), .A(\g.we_clk [3687]));
Q_ASSIGN U12704 ( .B(clk), .A(\g.we_clk [3686]));
Q_ASSIGN U12705 ( .B(clk), .A(\g.we_clk [3685]));
Q_ASSIGN U12706 ( .B(clk), .A(\g.we_clk [3684]));
Q_ASSIGN U12707 ( .B(clk), .A(\g.we_clk [3683]));
Q_ASSIGN U12708 ( .B(clk), .A(\g.we_clk [3682]));
Q_ASSIGN U12709 ( .B(clk), .A(\g.we_clk [3681]));
Q_ASSIGN U12710 ( .B(clk), .A(\g.we_clk [3680]));
Q_ASSIGN U12711 ( .B(clk), .A(\g.we_clk [3679]));
Q_ASSIGN U12712 ( .B(clk), .A(\g.we_clk [3678]));
Q_ASSIGN U12713 ( .B(clk), .A(\g.we_clk [3677]));
Q_ASSIGN U12714 ( .B(clk), .A(\g.we_clk [3676]));
Q_ASSIGN U12715 ( .B(clk), .A(\g.we_clk [3675]));
Q_ASSIGN U12716 ( .B(clk), .A(\g.we_clk [3674]));
Q_ASSIGN U12717 ( .B(clk), .A(\g.we_clk [3673]));
Q_ASSIGN U12718 ( .B(clk), .A(\g.we_clk [3672]));
Q_ASSIGN U12719 ( .B(clk), .A(\g.we_clk [3671]));
Q_ASSIGN U12720 ( .B(clk), .A(\g.we_clk [3670]));
Q_ASSIGN U12721 ( .B(clk), .A(\g.we_clk [3669]));
Q_ASSIGN U12722 ( .B(clk), .A(\g.we_clk [3668]));
Q_ASSIGN U12723 ( .B(clk), .A(\g.we_clk [3667]));
Q_ASSIGN U12724 ( .B(clk), .A(\g.we_clk [3666]));
Q_ASSIGN U12725 ( .B(clk), .A(\g.we_clk [3665]));
Q_ASSIGN U12726 ( .B(clk), .A(\g.we_clk [3664]));
Q_ASSIGN U12727 ( .B(clk), .A(\g.we_clk [3663]));
Q_ASSIGN U12728 ( .B(clk), .A(\g.we_clk [3662]));
Q_ASSIGN U12729 ( .B(clk), .A(\g.we_clk [3661]));
Q_ASSIGN U12730 ( .B(clk), .A(\g.we_clk [3660]));
Q_ASSIGN U12731 ( .B(clk), .A(\g.we_clk [3659]));
Q_ASSIGN U12732 ( .B(clk), .A(\g.we_clk [3658]));
Q_ASSIGN U12733 ( .B(clk), .A(\g.we_clk [3657]));
Q_ASSIGN U12734 ( .B(clk), .A(\g.we_clk [3656]));
Q_ASSIGN U12735 ( .B(clk), .A(\g.we_clk [3655]));
Q_ASSIGN U12736 ( .B(clk), .A(\g.we_clk [3654]));
Q_ASSIGN U12737 ( .B(clk), .A(\g.we_clk [3653]));
Q_ASSIGN U12738 ( .B(clk), .A(\g.we_clk [3652]));
Q_ASSIGN U12739 ( .B(clk), .A(\g.we_clk [3651]));
Q_ASSIGN U12740 ( .B(clk), .A(\g.we_clk [3650]));
Q_ASSIGN U12741 ( .B(clk), .A(\g.we_clk [3649]));
Q_ASSIGN U12742 ( .B(clk), .A(\g.we_clk [3648]));
Q_ASSIGN U12743 ( .B(clk), .A(\g.we_clk [3647]));
Q_ASSIGN U12744 ( .B(clk), .A(\g.we_clk [3646]));
Q_ASSIGN U12745 ( .B(clk), .A(\g.we_clk [3645]));
Q_ASSIGN U12746 ( .B(clk), .A(\g.we_clk [3644]));
Q_ASSIGN U12747 ( .B(clk), .A(\g.we_clk [3643]));
Q_ASSIGN U12748 ( .B(clk), .A(\g.we_clk [3642]));
Q_ASSIGN U12749 ( .B(clk), .A(\g.we_clk [3641]));
Q_ASSIGN U12750 ( .B(clk), .A(\g.we_clk [3640]));
Q_ASSIGN U12751 ( .B(clk), .A(\g.we_clk [3639]));
Q_ASSIGN U12752 ( .B(clk), .A(\g.we_clk [3638]));
Q_ASSIGN U12753 ( .B(clk), .A(\g.we_clk [3637]));
Q_ASSIGN U12754 ( .B(clk), .A(\g.we_clk [3636]));
Q_ASSIGN U12755 ( .B(clk), .A(\g.we_clk [3635]));
Q_ASSIGN U12756 ( .B(clk), .A(\g.we_clk [3634]));
Q_ASSIGN U12757 ( .B(clk), .A(\g.we_clk [3633]));
Q_ASSIGN U12758 ( .B(clk), .A(\g.we_clk [3632]));
Q_ASSIGN U12759 ( .B(clk), .A(\g.we_clk [3631]));
Q_ASSIGN U12760 ( .B(clk), .A(\g.we_clk [3630]));
Q_ASSIGN U12761 ( .B(clk), .A(\g.we_clk [3629]));
Q_ASSIGN U12762 ( .B(clk), .A(\g.we_clk [3628]));
Q_ASSIGN U12763 ( .B(clk), .A(\g.we_clk [3627]));
Q_ASSIGN U12764 ( .B(clk), .A(\g.we_clk [3626]));
Q_ASSIGN U12765 ( .B(clk), .A(\g.we_clk [3625]));
Q_ASSIGN U12766 ( .B(clk), .A(\g.we_clk [3624]));
Q_ASSIGN U12767 ( .B(clk), .A(\g.we_clk [3623]));
Q_ASSIGN U12768 ( .B(clk), .A(\g.we_clk [3622]));
Q_ASSIGN U12769 ( .B(clk), .A(\g.we_clk [3621]));
Q_ASSIGN U12770 ( .B(clk), .A(\g.we_clk [3620]));
Q_ASSIGN U12771 ( .B(clk), .A(\g.we_clk [3619]));
Q_ASSIGN U12772 ( .B(clk), .A(\g.we_clk [3618]));
Q_ASSIGN U12773 ( .B(clk), .A(\g.we_clk [3617]));
Q_ASSIGN U12774 ( .B(clk), .A(\g.we_clk [3616]));
Q_ASSIGN U12775 ( .B(clk), .A(\g.we_clk [3615]));
Q_ASSIGN U12776 ( .B(clk), .A(\g.we_clk [3614]));
Q_ASSIGN U12777 ( .B(clk), .A(\g.we_clk [3613]));
Q_ASSIGN U12778 ( .B(clk), .A(\g.we_clk [3612]));
Q_ASSIGN U12779 ( .B(clk), .A(\g.we_clk [3611]));
Q_ASSIGN U12780 ( .B(clk), .A(\g.we_clk [3610]));
Q_ASSIGN U12781 ( .B(clk), .A(\g.we_clk [3609]));
Q_ASSIGN U12782 ( .B(clk), .A(\g.we_clk [3608]));
Q_ASSIGN U12783 ( .B(clk), .A(\g.we_clk [3607]));
Q_ASSIGN U12784 ( .B(clk), .A(\g.we_clk [3606]));
Q_ASSIGN U12785 ( .B(clk), .A(\g.we_clk [3605]));
Q_ASSIGN U12786 ( .B(clk), .A(\g.we_clk [3604]));
Q_ASSIGN U12787 ( .B(clk), .A(\g.we_clk [3603]));
Q_ASSIGN U12788 ( .B(clk), .A(\g.we_clk [3602]));
Q_ASSIGN U12789 ( .B(clk), .A(\g.we_clk [3601]));
Q_ASSIGN U12790 ( .B(clk), .A(\g.we_clk [3600]));
Q_ASSIGN U12791 ( .B(clk), .A(\g.we_clk [3599]));
Q_ASSIGN U12792 ( .B(clk), .A(\g.we_clk [3598]));
Q_ASSIGN U12793 ( .B(clk), .A(\g.we_clk [3597]));
Q_ASSIGN U12794 ( .B(clk), .A(\g.we_clk [3596]));
Q_ASSIGN U12795 ( .B(clk), .A(\g.we_clk [3595]));
Q_ASSIGN U12796 ( .B(clk), .A(\g.we_clk [3594]));
Q_ASSIGN U12797 ( .B(clk), .A(\g.we_clk [3593]));
Q_ASSIGN U12798 ( .B(clk), .A(\g.we_clk [3592]));
Q_ASSIGN U12799 ( .B(clk), .A(\g.we_clk [3591]));
Q_ASSIGN U12800 ( .B(clk), .A(\g.we_clk [3590]));
Q_ASSIGN U12801 ( .B(clk), .A(\g.we_clk [3589]));
Q_ASSIGN U12802 ( .B(clk), .A(\g.we_clk [3588]));
Q_ASSIGN U12803 ( .B(clk), .A(\g.we_clk [3587]));
Q_ASSIGN U12804 ( .B(clk), .A(\g.we_clk [3586]));
Q_ASSIGN U12805 ( .B(clk), .A(\g.we_clk [3585]));
Q_ASSIGN U12806 ( .B(clk), .A(\g.we_clk [3584]));
Q_ASSIGN U12807 ( .B(clk), .A(\g.we_clk [3583]));
Q_ASSIGN U12808 ( .B(clk), .A(\g.we_clk [3582]));
Q_ASSIGN U12809 ( .B(clk), .A(\g.we_clk [3581]));
Q_ASSIGN U12810 ( .B(clk), .A(\g.we_clk [3580]));
Q_ASSIGN U12811 ( .B(clk), .A(\g.we_clk [3579]));
Q_ASSIGN U12812 ( .B(clk), .A(\g.we_clk [3578]));
Q_ASSIGN U12813 ( .B(clk), .A(\g.we_clk [3577]));
Q_ASSIGN U12814 ( .B(clk), .A(\g.we_clk [3576]));
Q_ASSIGN U12815 ( .B(clk), .A(\g.we_clk [3575]));
Q_ASSIGN U12816 ( .B(clk), .A(\g.we_clk [3574]));
Q_ASSIGN U12817 ( .B(clk), .A(\g.we_clk [3573]));
Q_ASSIGN U12818 ( .B(clk), .A(\g.we_clk [3572]));
Q_ASSIGN U12819 ( .B(clk), .A(\g.we_clk [3571]));
Q_ASSIGN U12820 ( .B(clk), .A(\g.we_clk [3570]));
Q_ASSIGN U12821 ( .B(clk), .A(\g.we_clk [3569]));
Q_ASSIGN U12822 ( .B(clk), .A(\g.we_clk [3568]));
Q_ASSIGN U12823 ( .B(clk), .A(\g.we_clk [3567]));
Q_ASSIGN U12824 ( .B(clk), .A(\g.we_clk [3566]));
Q_ASSIGN U12825 ( .B(clk), .A(\g.we_clk [3565]));
Q_ASSIGN U12826 ( .B(clk), .A(\g.we_clk [3564]));
Q_ASSIGN U12827 ( .B(clk), .A(\g.we_clk [3563]));
Q_ASSIGN U12828 ( .B(clk), .A(\g.we_clk [3562]));
Q_ASSIGN U12829 ( .B(clk), .A(\g.we_clk [3561]));
Q_ASSIGN U12830 ( .B(clk), .A(\g.we_clk [3560]));
Q_ASSIGN U12831 ( .B(clk), .A(\g.we_clk [3559]));
Q_ASSIGN U12832 ( .B(clk), .A(\g.we_clk [3558]));
Q_ASSIGN U12833 ( .B(clk), .A(\g.we_clk [3557]));
Q_ASSIGN U12834 ( .B(clk), .A(\g.we_clk [3556]));
Q_ASSIGN U12835 ( .B(clk), .A(\g.we_clk [3555]));
Q_ASSIGN U12836 ( .B(clk), .A(\g.we_clk [3554]));
Q_ASSIGN U12837 ( .B(clk), .A(\g.we_clk [3553]));
Q_ASSIGN U12838 ( .B(clk), .A(\g.we_clk [3552]));
Q_ASSIGN U12839 ( .B(clk), .A(\g.we_clk [3551]));
Q_ASSIGN U12840 ( .B(clk), .A(\g.we_clk [3550]));
Q_ASSIGN U12841 ( .B(clk), .A(\g.we_clk [3549]));
Q_ASSIGN U12842 ( .B(clk), .A(\g.we_clk [3548]));
Q_ASSIGN U12843 ( .B(clk), .A(\g.we_clk [3547]));
Q_ASSIGN U12844 ( .B(clk), .A(\g.we_clk [3546]));
Q_ASSIGN U12845 ( .B(clk), .A(\g.we_clk [3545]));
Q_ASSIGN U12846 ( .B(clk), .A(\g.we_clk [3544]));
Q_ASSIGN U12847 ( .B(clk), .A(\g.we_clk [3543]));
Q_ASSIGN U12848 ( .B(clk), .A(\g.we_clk [3542]));
Q_ASSIGN U12849 ( .B(clk), .A(\g.we_clk [3541]));
Q_ASSIGN U12850 ( .B(clk), .A(\g.we_clk [3540]));
Q_ASSIGN U12851 ( .B(clk), .A(\g.we_clk [3539]));
Q_ASSIGN U12852 ( .B(clk), .A(\g.we_clk [3538]));
Q_ASSIGN U12853 ( .B(clk), .A(\g.we_clk [3537]));
Q_ASSIGN U12854 ( .B(clk), .A(\g.we_clk [3536]));
Q_ASSIGN U12855 ( .B(clk), .A(\g.we_clk [3535]));
Q_ASSIGN U12856 ( .B(clk), .A(\g.we_clk [3534]));
Q_ASSIGN U12857 ( .B(clk), .A(\g.we_clk [3533]));
Q_ASSIGN U12858 ( .B(clk), .A(\g.we_clk [3532]));
Q_ASSIGN U12859 ( .B(clk), .A(\g.we_clk [3531]));
Q_ASSIGN U12860 ( .B(clk), .A(\g.we_clk [3530]));
Q_ASSIGN U12861 ( .B(clk), .A(\g.we_clk [3529]));
Q_ASSIGN U12862 ( .B(clk), .A(\g.we_clk [3528]));
Q_ASSIGN U12863 ( .B(clk), .A(\g.we_clk [3527]));
Q_ASSIGN U12864 ( .B(clk), .A(\g.we_clk [3526]));
Q_ASSIGN U12865 ( .B(clk), .A(\g.we_clk [3525]));
Q_ASSIGN U12866 ( .B(clk), .A(\g.we_clk [3524]));
Q_ASSIGN U12867 ( .B(clk), .A(\g.we_clk [3523]));
Q_ASSIGN U12868 ( .B(clk), .A(\g.we_clk [3522]));
Q_ASSIGN U12869 ( .B(clk), .A(\g.we_clk [3521]));
Q_ASSIGN U12870 ( .B(clk), .A(\g.we_clk [3520]));
Q_ASSIGN U12871 ( .B(clk), .A(\g.we_clk [3519]));
Q_ASSIGN U12872 ( .B(clk), .A(\g.we_clk [3518]));
Q_ASSIGN U12873 ( .B(clk), .A(\g.we_clk [3517]));
Q_ASSIGN U12874 ( .B(clk), .A(\g.we_clk [3516]));
Q_ASSIGN U12875 ( .B(clk), .A(\g.we_clk [3515]));
Q_ASSIGN U12876 ( .B(clk), .A(\g.we_clk [3514]));
Q_ASSIGN U12877 ( .B(clk), .A(\g.we_clk [3513]));
Q_ASSIGN U12878 ( .B(clk), .A(\g.we_clk [3512]));
Q_ASSIGN U12879 ( .B(clk), .A(\g.we_clk [3511]));
Q_ASSIGN U12880 ( .B(clk), .A(\g.we_clk [3510]));
Q_ASSIGN U12881 ( .B(clk), .A(\g.we_clk [3509]));
Q_ASSIGN U12882 ( .B(clk), .A(\g.we_clk [3508]));
Q_ASSIGN U12883 ( .B(clk), .A(\g.we_clk [3507]));
Q_ASSIGN U12884 ( .B(clk), .A(\g.we_clk [3506]));
Q_ASSIGN U12885 ( .B(clk), .A(\g.we_clk [3505]));
Q_ASSIGN U12886 ( .B(clk), .A(\g.we_clk [3504]));
Q_ASSIGN U12887 ( .B(clk), .A(\g.we_clk [3503]));
Q_ASSIGN U12888 ( .B(clk), .A(\g.we_clk [3502]));
Q_ASSIGN U12889 ( .B(clk), .A(\g.we_clk [3501]));
Q_ASSIGN U12890 ( .B(clk), .A(\g.we_clk [3500]));
Q_ASSIGN U12891 ( .B(clk), .A(\g.we_clk [3499]));
Q_ASSIGN U12892 ( .B(clk), .A(\g.we_clk [3498]));
Q_ASSIGN U12893 ( .B(clk), .A(\g.we_clk [3497]));
Q_ASSIGN U12894 ( .B(clk), .A(\g.we_clk [3496]));
Q_ASSIGN U12895 ( .B(clk), .A(\g.we_clk [3495]));
Q_ASSIGN U12896 ( .B(clk), .A(\g.we_clk [3494]));
Q_ASSIGN U12897 ( .B(clk), .A(\g.we_clk [3493]));
Q_ASSIGN U12898 ( .B(clk), .A(\g.we_clk [3492]));
Q_ASSIGN U12899 ( .B(clk), .A(\g.we_clk [3491]));
Q_ASSIGN U12900 ( .B(clk), .A(\g.we_clk [3490]));
Q_ASSIGN U12901 ( .B(clk), .A(\g.we_clk [3489]));
Q_ASSIGN U12902 ( .B(clk), .A(\g.we_clk [3488]));
Q_ASSIGN U12903 ( .B(clk), .A(\g.we_clk [3487]));
Q_ASSIGN U12904 ( .B(clk), .A(\g.we_clk [3486]));
Q_ASSIGN U12905 ( .B(clk), .A(\g.we_clk [3485]));
Q_ASSIGN U12906 ( .B(clk), .A(\g.we_clk [3484]));
Q_ASSIGN U12907 ( .B(clk), .A(\g.we_clk [3483]));
Q_ASSIGN U12908 ( .B(clk), .A(\g.we_clk [3482]));
Q_ASSIGN U12909 ( .B(clk), .A(\g.we_clk [3481]));
Q_ASSIGN U12910 ( .B(clk), .A(\g.we_clk [3480]));
Q_ASSIGN U12911 ( .B(clk), .A(\g.we_clk [3479]));
Q_ASSIGN U12912 ( .B(clk), .A(\g.we_clk [3478]));
Q_ASSIGN U12913 ( .B(clk), .A(\g.we_clk [3477]));
Q_ASSIGN U12914 ( .B(clk), .A(\g.we_clk [3476]));
Q_ASSIGN U12915 ( .B(clk), .A(\g.we_clk [3475]));
Q_ASSIGN U12916 ( .B(clk), .A(\g.we_clk [3474]));
Q_ASSIGN U12917 ( .B(clk), .A(\g.we_clk [3473]));
Q_ASSIGN U12918 ( .B(clk), .A(\g.we_clk [3472]));
Q_ASSIGN U12919 ( .B(clk), .A(\g.we_clk [3471]));
Q_ASSIGN U12920 ( .B(clk), .A(\g.we_clk [3470]));
Q_ASSIGN U12921 ( .B(clk), .A(\g.we_clk [3469]));
Q_ASSIGN U12922 ( .B(clk), .A(\g.we_clk [3468]));
Q_ASSIGN U12923 ( .B(clk), .A(\g.we_clk [3467]));
Q_ASSIGN U12924 ( .B(clk), .A(\g.we_clk [3466]));
Q_ASSIGN U12925 ( .B(clk), .A(\g.we_clk [3465]));
Q_ASSIGN U12926 ( .B(clk), .A(\g.we_clk [3464]));
Q_ASSIGN U12927 ( .B(clk), .A(\g.we_clk [3463]));
Q_ASSIGN U12928 ( .B(clk), .A(\g.we_clk [3462]));
Q_ASSIGN U12929 ( .B(clk), .A(\g.we_clk [3461]));
Q_ASSIGN U12930 ( .B(clk), .A(\g.we_clk [3460]));
Q_ASSIGN U12931 ( .B(clk), .A(\g.we_clk [3459]));
Q_ASSIGN U12932 ( .B(clk), .A(\g.we_clk [3458]));
Q_ASSIGN U12933 ( .B(clk), .A(\g.we_clk [3457]));
Q_ASSIGN U12934 ( .B(clk), .A(\g.we_clk [3456]));
Q_ASSIGN U12935 ( .B(clk), .A(\g.we_clk [3455]));
Q_ASSIGN U12936 ( .B(clk), .A(\g.we_clk [3454]));
Q_ASSIGN U12937 ( .B(clk), .A(\g.we_clk [3453]));
Q_ASSIGN U12938 ( .B(clk), .A(\g.we_clk [3452]));
Q_ASSIGN U12939 ( .B(clk), .A(\g.we_clk [3451]));
Q_ASSIGN U12940 ( .B(clk), .A(\g.we_clk [3450]));
Q_ASSIGN U12941 ( .B(clk), .A(\g.we_clk [3449]));
Q_ASSIGN U12942 ( .B(clk), .A(\g.we_clk [3448]));
Q_ASSIGN U12943 ( .B(clk), .A(\g.we_clk [3447]));
Q_ASSIGN U12944 ( .B(clk), .A(\g.we_clk [3446]));
Q_ASSIGN U12945 ( .B(clk), .A(\g.we_clk [3445]));
Q_ASSIGN U12946 ( .B(clk), .A(\g.we_clk [3444]));
Q_ASSIGN U12947 ( .B(clk), .A(\g.we_clk [3443]));
Q_ASSIGN U12948 ( .B(clk), .A(\g.we_clk [3442]));
Q_ASSIGN U12949 ( .B(clk), .A(\g.we_clk [3441]));
Q_ASSIGN U12950 ( .B(clk), .A(\g.we_clk [3440]));
Q_ASSIGN U12951 ( .B(clk), .A(\g.we_clk [3439]));
Q_ASSIGN U12952 ( .B(clk), .A(\g.we_clk [3438]));
Q_ASSIGN U12953 ( .B(clk), .A(\g.we_clk [3437]));
Q_ASSIGN U12954 ( .B(clk), .A(\g.we_clk [3436]));
Q_ASSIGN U12955 ( .B(clk), .A(\g.we_clk [3435]));
Q_ASSIGN U12956 ( .B(clk), .A(\g.we_clk [3434]));
Q_ASSIGN U12957 ( .B(clk), .A(\g.we_clk [3433]));
Q_ASSIGN U12958 ( .B(clk), .A(\g.we_clk [3432]));
Q_ASSIGN U12959 ( .B(clk), .A(\g.we_clk [3431]));
Q_ASSIGN U12960 ( .B(clk), .A(\g.we_clk [3430]));
Q_ASSIGN U12961 ( .B(clk), .A(\g.we_clk [3429]));
Q_ASSIGN U12962 ( .B(clk), .A(\g.we_clk [3428]));
Q_ASSIGN U12963 ( .B(clk), .A(\g.we_clk [3427]));
Q_ASSIGN U12964 ( .B(clk), .A(\g.we_clk [3426]));
Q_ASSIGN U12965 ( .B(clk), .A(\g.we_clk [3425]));
Q_ASSIGN U12966 ( .B(clk), .A(\g.we_clk [3424]));
Q_ASSIGN U12967 ( .B(clk), .A(\g.we_clk [3423]));
Q_ASSIGN U12968 ( .B(clk), .A(\g.we_clk [3422]));
Q_ASSIGN U12969 ( .B(clk), .A(\g.we_clk [3421]));
Q_ASSIGN U12970 ( .B(clk), .A(\g.we_clk [3420]));
Q_ASSIGN U12971 ( .B(clk), .A(\g.we_clk [3419]));
Q_ASSIGN U12972 ( .B(clk), .A(\g.we_clk [3418]));
Q_ASSIGN U12973 ( .B(clk), .A(\g.we_clk [3417]));
Q_ASSIGN U12974 ( .B(clk), .A(\g.we_clk [3416]));
Q_ASSIGN U12975 ( .B(clk), .A(\g.we_clk [3415]));
Q_ASSIGN U12976 ( .B(clk), .A(\g.we_clk [3414]));
Q_ASSIGN U12977 ( .B(clk), .A(\g.we_clk [3413]));
Q_ASSIGN U12978 ( .B(clk), .A(\g.we_clk [3412]));
Q_ASSIGN U12979 ( .B(clk), .A(\g.we_clk [3411]));
Q_ASSIGN U12980 ( .B(clk), .A(\g.we_clk [3410]));
Q_ASSIGN U12981 ( .B(clk), .A(\g.we_clk [3409]));
Q_ASSIGN U12982 ( .B(clk), .A(\g.we_clk [3408]));
Q_ASSIGN U12983 ( .B(clk), .A(\g.we_clk [3407]));
Q_ASSIGN U12984 ( .B(clk), .A(\g.we_clk [3406]));
Q_ASSIGN U12985 ( .B(clk), .A(\g.we_clk [3405]));
Q_ASSIGN U12986 ( .B(clk), .A(\g.we_clk [3404]));
Q_ASSIGN U12987 ( .B(clk), .A(\g.we_clk [3403]));
Q_ASSIGN U12988 ( .B(clk), .A(\g.we_clk [3402]));
Q_ASSIGN U12989 ( .B(clk), .A(\g.we_clk [3401]));
Q_ASSIGN U12990 ( .B(clk), .A(\g.we_clk [3400]));
Q_ASSIGN U12991 ( .B(clk), .A(\g.we_clk [3399]));
Q_ASSIGN U12992 ( .B(clk), .A(\g.we_clk [3398]));
Q_ASSIGN U12993 ( .B(clk), .A(\g.we_clk [3397]));
Q_ASSIGN U12994 ( .B(clk), .A(\g.we_clk [3396]));
Q_ASSIGN U12995 ( .B(clk), .A(\g.we_clk [3395]));
Q_ASSIGN U12996 ( .B(clk), .A(\g.we_clk [3394]));
Q_ASSIGN U12997 ( .B(clk), .A(\g.we_clk [3393]));
Q_ASSIGN U12998 ( .B(clk), .A(\g.we_clk [3392]));
Q_ASSIGN U12999 ( .B(clk), .A(\g.we_clk [3391]));
Q_ASSIGN U13000 ( .B(clk), .A(\g.we_clk [3390]));
Q_ASSIGN U13001 ( .B(clk), .A(\g.we_clk [3389]));
Q_ASSIGN U13002 ( .B(clk), .A(\g.we_clk [3388]));
Q_ASSIGN U13003 ( .B(clk), .A(\g.we_clk [3387]));
Q_ASSIGN U13004 ( .B(clk), .A(\g.we_clk [3386]));
Q_ASSIGN U13005 ( .B(clk), .A(\g.we_clk [3385]));
Q_ASSIGN U13006 ( .B(clk), .A(\g.we_clk [3384]));
Q_ASSIGN U13007 ( .B(clk), .A(\g.we_clk [3383]));
Q_ASSIGN U13008 ( .B(clk), .A(\g.we_clk [3382]));
Q_ASSIGN U13009 ( .B(clk), .A(\g.we_clk [3381]));
Q_ASSIGN U13010 ( .B(clk), .A(\g.we_clk [3380]));
Q_ASSIGN U13011 ( .B(clk), .A(\g.we_clk [3379]));
Q_ASSIGN U13012 ( .B(clk), .A(\g.we_clk [3378]));
Q_ASSIGN U13013 ( .B(clk), .A(\g.we_clk [3377]));
Q_ASSIGN U13014 ( .B(clk), .A(\g.we_clk [3376]));
Q_ASSIGN U13015 ( .B(clk), .A(\g.we_clk [3375]));
Q_ASSIGN U13016 ( .B(clk), .A(\g.we_clk [3374]));
Q_ASSIGN U13017 ( .B(clk), .A(\g.we_clk [3373]));
Q_ASSIGN U13018 ( .B(clk), .A(\g.we_clk [3372]));
Q_ASSIGN U13019 ( .B(clk), .A(\g.we_clk [3371]));
Q_ASSIGN U13020 ( .B(clk), .A(\g.we_clk [3370]));
Q_ASSIGN U13021 ( .B(clk), .A(\g.we_clk [3369]));
Q_ASSIGN U13022 ( .B(clk), .A(\g.we_clk [3368]));
Q_ASSIGN U13023 ( .B(clk), .A(\g.we_clk [3367]));
Q_ASSIGN U13024 ( .B(clk), .A(\g.we_clk [3366]));
Q_ASSIGN U13025 ( .B(clk), .A(\g.we_clk [3365]));
Q_ASSIGN U13026 ( .B(clk), .A(\g.we_clk [3364]));
Q_ASSIGN U13027 ( .B(clk), .A(\g.we_clk [3363]));
Q_ASSIGN U13028 ( .B(clk), .A(\g.we_clk [3362]));
Q_ASSIGN U13029 ( .B(clk), .A(\g.we_clk [3361]));
Q_ASSIGN U13030 ( .B(clk), .A(\g.we_clk [3360]));
Q_ASSIGN U13031 ( .B(clk), .A(\g.we_clk [3359]));
Q_ASSIGN U13032 ( .B(clk), .A(\g.we_clk [3358]));
Q_ASSIGN U13033 ( .B(clk), .A(\g.we_clk [3357]));
Q_ASSIGN U13034 ( .B(clk), .A(\g.we_clk [3356]));
Q_ASSIGN U13035 ( .B(clk), .A(\g.we_clk [3355]));
Q_ASSIGN U13036 ( .B(clk), .A(\g.we_clk [3354]));
Q_ASSIGN U13037 ( .B(clk), .A(\g.we_clk [3353]));
Q_ASSIGN U13038 ( .B(clk), .A(\g.we_clk [3352]));
Q_ASSIGN U13039 ( .B(clk), .A(\g.we_clk [3351]));
Q_ASSIGN U13040 ( .B(clk), .A(\g.we_clk [3350]));
Q_ASSIGN U13041 ( .B(clk), .A(\g.we_clk [3349]));
Q_ASSIGN U13042 ( .B(clk), .A(\g.we_clk [3348]));
Q_ASSIGN U13043 ( .B(clk), .A(\g.we_clk [3347]));
Q_ASSIGN U13044 ( .B(clk), .A(\g.we_clk [3346]));
Q_ASSIGN U13045 ( .B(clk), .A(\g.we_clk [3345]));
Q_ASSIGN U13046 ( .B(clk), .A(\g.we_clk [3344]));
Q_ASSIGN U13047 ( .B(clk), .A(\g.we_clk [3343]));
Q_ASSIGN U13048 ( .B(clk), .A(\g.we_clk [3342]));
Q_ASSIGN U13049 ( .B(clk), .A(\g.we_clk [3341]));
Q_ASSIGN U13050 ( .B(clk), .A(\g.we_clk [3340]));
Q_ASSIGN U13051 ( .B(clk), .A(\g.we_clk [3339]));
Q_ASSIGN U13052 ( .B(clk), .A(\g.we_clk [3338]));
Q_ASSIGN U13053 ( .B(clk), .A(\g.we_clk [3337]));
Q_ASSIGN U13054 ( .B(clk), .A(\g.we_clk [3336]));
Q_ASSIGN U13055 ( .B(clk), .A(\g.we_clk [3335]));
Q_ASSIGN U13056 ( .B(clk), .A(\g.we_clk [3334]));
Q_ASSIGN U13057 ( .B(clk), .A(\g.we_clk [3333]));
Q_ASSIGN U13058 ( .B(clk), .A(\g.we_clk [3332]));
Q_ASSIGN U13059 ( .B(clk), .A(\g.we_clk [3331]));
Q_ASSIGN U13060 ( .B(clk), .A(\g.we_clk [3330]));
Q_ASSIGN U13061 ( .B(clk), .A(\g.we_clk [3329]));
Q_ASSIGN U13062 ( .B(clk), .A(\g.we_clk [3328]));
Q_ASSIGN U13063 ( .B(clk), .A(\g.we_clk [3327]));
Q_ASSIGN U13064 ( .B(clk), .A(\g.we_clk [3326]));
Q_ASSIGN U13065 ( .B(clk), .A(\g.we_clk [3325]));
Q_ASSIGN U13066 ( .B(clk), .A(\g.we_clk [3324]));
Q_ASSIGN U13067 ( .B(clk), .A(\g.we_clk [3323]));
Q_ASSIGN U13068 ( .B(clk), .A(\g.we_clk [3322]));
Q_ASSIGN U13069 ( .B(clk), .A(\g.we_clk [3321]));
Q_ASSIGN U13070 ( .B(clk), .A(\g.we_clk [3320]));
Q_ASSIGN U13071 ( .B(clk), .A(\g.we_clk [3319]));
Q_ASSIGN U13072 ( .B(clk), .A(\g.we_clk [3318]));
Q_ASSIGN U13073 ( .B(clk), .A(\g.we_clk [3317]));
Q_ASSIGN U13074 ( .B(clk), .A(\g.we_clk [3316]));
Q_ASSIGN U13075 ( .B(clk), .A(\g.we_clk [3315]));
Q_ASSIGN U13076 ( .B(clk), .A(\g.we_clk [3314]));
Q_ASSIGN U13077 ( .B(clk), .A(\g.we_clk [3313]));
Q_ASSIGN U13078 ( .B(clk), .A(\g.we_clk [3312]));
Q_ASSIGN U13079 ( .B(clk), .A(\g.we_clk [3311]));
Q_ASSIGN U13080 ( .B(clk), .A(\g.we_clk [3310]));
Q_ASSIGN U13081 ( .B(clk), .A(\g.we_clk [3309]));
Q_ASSIGN U13082 ( .B(clk), .A(\g.we_clk [3308]));
Q_ASSIGN U13083 ( .B(clk), .A(\g.we_clk [3307]));
Q_ASSIGN U13084 ( .B(clk), .A(\g.we_clk [3306]));
Q_ASSIGN U13085 ( .B(clk), .A(\g.we_clk [3305]));
Q_ASSIGN U13086 ( .B(clk), .A(\g.we_clk [3304]));
Q_ASSIGN U13087 ( .B(clk), .A(\g.we_clk [3303]));
Q_ASSIGN U13088 ( .B(clk), .A(\g.we_clk [3302]));
Q_ASSIGN U13089 ( .B(clk), .A(\g.we_clk [3301]));
Q_ASSIGN U13090 ( .B(clk), .A(\g.we_clk [3300]));
Q_ASSIGN U13091 ( .B(clk), .A(\g.we_clk [3299]));
Q_ASSIGN U13092 ( .B(clk), .A(\g.we_clk [3298]));
Q_ASSIGN U13093 ( .B(clk), .A(\g.we_clk [3297]));
Q_ASSIGN U13094 ( .B(clk), .A(\g.we_clk [3296]));
Q_ASSIGN U13095 ( .B(clk), .A(\g.we_clk [3295]));
Q_ASSIGN U13096 ( .B(clk), .A(\g.we_clk [3294]));
Q_ASSIGN U13097 ( .B(clk), .A(\g.we_clk [3293]));
Q_ASSIGN U13098 ( .B(clk), .A(\g.we_clk [3292]));
Q_ASSIGN U13099 ( .B(clk), .A(\g.we_clk [3291]));
Q_ASSIGN U13100 ( .B(clk), .A(\g.we_clk [3290]));
Q_ASSIGN U13101 ( .B(clk), .A(\g.we_clk [3289]));
Q_ASSIGN U13102 ( .B(clk), .A(\g.we_clk [3288]));
Q_ASSIGN U13103 ( .B(clk), .A(\g.we_clk [3287]));
Q_ASSIGN U13104 ( .B(clk), .A(\g.we_clk [3286]));
Q_ASSIGN U13105 ( .B(clk), .A(\g.we_clk [3285]));
Q_ASSIGN U13106 ( .B(clk), .A(\g.we_clk [3284]));
Q_ASSIGN U13107 ( .B(clk), .A(\g.we_clk [3283]));
Q_ASSIGN U13108 ( .B(clk), .A(\g.we_clk [3282]));
Q_ASSIGN U13109 ( .B(clk), .A(\g.we_clk [3281]));
Q_ASSIGN U13110 ( .B(clk), .A(\g.we_clk [3280]));
Q_ASSIGN U13111 ( .B(clk), .A(\g.we_clk [3279]));
Q_ASSIGN U13112 ( .B(clk), .A(\g.we_clk [3278]));
Q_ASSIGN U13113 ( .B(clk), .A(\g.we_clk [3277]));
Q_ASSIGN U13114 ( .B(clk), .A(\g.we_clk [3276]));
Q_ASSIGN U13115 ( .B(clk), .A(\g.we_clk [3275]));
Q_ASSIGN U13116 ( .B(clk), .A(\g.we_clk [3274]));
Q_ASSIGN U13117 ( .B(clk), .A(\g.we_clk [3273]));
Q_ASSIGN U13118 ( .B(clk), .A(\g.we_clk [3272]));
Q_ASSIGN U13119 ( .B(clk), .A(\g.we_clk [3271]));
Q_ASSIGN U13120 ( .B(clk), .A(\g.we_clk [3270]));
Q_ASSIGN U13121 ( .B(clk), .A(\g.we_clk [3269]));
Q_ASSIGN U13122 ( .B(clk), .A(\g.we_clk [3268]));
Q_ASSIGN U13123 ( .B(clk), .A(\g.we_clk [3267]));
Q_ASSIGN U13124 ( .B(clk), .A(\g.we_clk [3266]));
Q_ASSIGN U13125 ( .B(clk), .A(\g.we_clk [3265]));
Q_ASSIGN U13126 ( .B(clk), .A(\g.we_clk [3264]));
Q_ASSIGN U13127 ( .B(clk), .A(\g.we_clk [3263]));
Q_ASSIGN U13128 ( .B(clk), .A(\g.we_clk [3262]));
Q_ASSIGN U13129 ( .B(clk), .A(\g.we_clk [3261]));
Q_ASSIGN U13130 ( .B(clk), .A(\g.we_clk [3260]));
Q_ASSIGN U13131 ( .B(clk), .A(\g.we_clk [3259]));
Q_ASSIGN U13132 ( .B(clk), .A(\g.we_clk [3258]));
Q_ASSIGN U13133 ( .B(clk), .A(\g.we_clk [3257]));
Q_ASSIGN U13134 ( .B(clk), .A(\g.we_clk [3256]));
Q_ASSIGN U13135 ( .B(clk), .A(\g.we_clk [3255]));
Q_ASSIGN U13136 ( .B(clk), .A(\g.we_clk [3254]));
Q_ASSIGN U13137 ( .B(clk), .A(\g.we_clk [3253]));
Q_ASSIGN U13138 ( .B(clk), .A(\g.we_clk [3252]));
Q_ASSIGN U13139 ( .B(clk), .A(\g.we_clk [3251]));
Q_ASSIGN U13140 ( .B(clk), .A(\g.we_clk [3250]));
Q_ASSIGN U13141 ( .B(clk), .A(\g.we_clk [3249]));
Q_ASSIGN U13142 ( .B(clk), .A(\g.we_clk [3248]));
Q_ASSIGN U13143 ( .B(clk), .A(\g.we_clk [3247]));
Q_ASSIGN U13144 ( .B(clk), .A(\g.we_clk [3246]));
Q_ASSIGN U13145 ( .B(clk), .A(\g.we_clk [3245]));
Q_ASSIGN U13146 ( .B(clk), .A(\g.we_clk [3244]));
Q_ASSIGN U13147 ( .B(clk), .A(\g.we_clk [3243]));
Q_ASSIGN U13148 ( .B(clk), .A(\g.we_clk [3242]));
Q_ASSIGN U13149 ( .B(clk), .A(\g.we_clk [3241]));
Q_ASSIGN U13150 ( .B(clk), .A(\g.we_clk [3240]));
Q_ASSIGN U13151 ( .B(clk), .A(\g.we_clk [3239]));
Q_ASSIGN U13152 ( .B(clk), .A(\g.we_clk [3238]));
Q_ASSIGN U13153 ( .B(clk), .A(\g.we_clk [3237]));
Q_ASSIGN U13154 ( .B(clk), .A(\g.we_clk [3236]));
Q_ASSIGN U13155 ( .B(clk), .A(\g.we_clk [3235]));
Q_ASSIGN U13156 ( .B(clk), .A(\g.we_clk [3234]));
Q_ASSIGN U13157 ( .B(clk), .A(\g.we_clk [3233]));
Q_ASSIGN U13158 ( .B(clk), .A(\g.we_clk [3232]));
Q_ASSIGN U13159 ( .B(clk), .A(\g.we_clk [3231]));
Q_ASSIGN U13160 ( .B(clk), .A(\g.we_clk [3230]));
Q_ASSIGN U13161 ( .B(clk), .A(\g.we_clk [3229]));
Q_ASSIGN U13162 ( .B(clk), .A(\g.we_clk [3228]));
Q_ASSIGN U13163 ( .B(clk), .A(\g.we_clk [3227]));
Q_ASSIGN U13164 ( .B(clk), .A(\g.we_clk [3226]));
Q_ASSIGN U13165 ( .B(clk), .A(\g.we_clk [3225]));
Q_ASSIGN U13166 ( .B(clk), .A(\g.we_clk [3224]));
Q_ASSIGN U13167 ( .B(clk), .A(\g.we_clk [3223]));
Q_ASSIGN U13168 ( .B(clk), .A(\g.we_clk [3222]));
Q_ASSIGN U13169 ( .B(clk), .A(\g.we_clk [3221]));
Q_ASSIGN U13170 ( .B(clk), .A(\g.we_clk [3220]));
Q_ASSIGN U13171 ( .B(clk), .A(\g.we_clk [3219]));
Q_ASSIGN U13172 ( .B(clk), .A(\g.we_clk [3218]));
Q_ASSIGN U13173 ( .B(clk), .A(\g.we_clk [3217]));
Q_ASSIGN U13174 ( .B(clk), .A(\g.we_clk [3216]));
Q_ASSIGN U13175 ( .B(clk), .A(\g.we_clk [3215]));
Q_ASSIGN U13176 ( .B(clk), .A(\g.we_clk [3214]));
Q_ASSIGN U13177 ( .B(clk), .A(\g.we_clk [3213]));
Q_ASSIGN U13178 ( .B(clk), .A(\g.we_clk [3212]));
Q_ASSIGN U13179 ( .B(clk), .A(\g.we_clk [3211]));
Q_ASSIGN U13180 ( .B(clk), .A(\g.we_clk [3210]));
Q_ASSIGN U13181 ( .B(clk), .A(\g.we_clk [3209]));
Q_ASSIGN U13182 ( .B(clk), .A(\g.we_clk [3208]));
Q_ASSIGN U13183 ( .B(clk), .A(\g.we_clk [3207]));
Q_ASSIGN U13184 ( .B(clk), .A(\g.we_clk [3206]));
Q_ASSIGN U13185 ( .B(clk), .A(\g.we_clk [3205]));
Q_ASSIGN U13186 ( .B(clk), .A(\g.we_clk [3204]));
Q_ASSIGN U13187 ( .B(clk), .A(\g.we_clk [3203]));
Q_ASSIGN U13188 ( .B(clk), .A(\g.we_clk [3202]));
Q_ASSIGN U13189 ( .B(clk), .A(\g.we_clk [3201]));
Q_ASSIGN U13190 ( .B(clk), .A(\g.we_clk [3200]));
Q_ASSIGN U13191 ( .B(clk), .A(\g.we_clk [3199]));
Q_ASSIGN U13192 ( .B(clk), .A(\g.we_clk [3198]));
Q_ASSIGN U13193 ( .B(clk), .A(\g.we_clk [3197]));
Q_ASSIGN U13194 ( .B(clk), .A(\g.we_clk [3196]));
Q_ASSIGN U13195 ( .B(clk), .A(\g.we_clk [3195]));
Q_ASSIGN U13196 ( .B(clk), .A(\g.we_clk [3194]));
Q_ASSIGN U13197 ( .B(clk), .A(\g.we_clk [3193]));
Q_ASSIGN U13198 ( .B(clk), .A(\g.we_clk [3192]));
Q_ASSIGN U13199 ( .B(clk), .A(\g.we_clk [3191]));
Q_ASSIGN U13200 ( .B(clk), .A(\g.we_clk [3190]));
Q_ASSIGN U13201 ( .B(clk), .A(\g.we_clk [3189]));
Q_ASSIGN U13202 ( .B(clk), .A(\g.we_clk [3188]));
Q_ASSIGN U13203 ( .B(clk), .A(\g.we_clk [3187]));
Q_ASSIGN U13204 ( .B(clk), .A(\g.we_clk [3186]));
Q_ASSIGN U13205 ( .B(clk), .A(\g.we_clk [3185]));
Q_ASSIGN U13206 ( .B(clk), .A(\g.we_clk [3184]));
Q_ASSIGN U13207 ( .B(clk), .A(\g.we_clk [3183]));
Q_ASSIGN U13208 ( .B(clk), .A(\g.we_clk [3182]));
Q_ASSIGN U13209 ( .B(clk), .A(\g.we_clk [3181]));
Q_ASSIGN U13210 ( .B(clk), .A(\g.we_clk [3180]));
Q_ASSIGN U13211 ( .B(clk), .A(\g.we_clk [3179]));
Q_ASSIGN U13212 ( .B(clk), .A(\g.we_clk [3178]));
Q_ASSIGN U13213 ( .B(clk), .A(\g.we_clk [3177]));
Q_ASSIGN U13214 ( .B(clk), .A(\g.we_clk [3176]));
Q_ASSIGN U13215 ( .B(clk), .A(\g.we_clk [3175]));
Q_ASSIGN U13216 ( .B(clk), .A(\g.we_clk [3174]));
Q_ASSIGN U13217 ( .B(clk), .A(\g.we_clk [3173]));
Q_ASSIGN U13218 ( .B(clk), .A(\g.we_clk [3172]));
Q_ASSIGN U13219 ( .B(clk), .A(\g.we_clk [3171]));
Q_ASSIGN U13220 ( .B(clk), .A(\g.we_clk [3170]));
Q_ASSIGN U13221 ( .B(clk), .A(\g.we_clk [3169]));
Q_ASSIGN U13222 ( .B(clk), .A(\g.we_clk [3168]));
Q_ASSIGN U13223 ( .B(clk), .A(\g.we_clk [3167]));
Q_ASSIGN U13224 ( .B(clk), .A(\g.we_clk [3166]));
Q_ASSIGN U13225 ( .B(clk), .A(\g.we_clk [3165]));
Q_ASSIGN U13226 ( .B(clk), .A(\g.we_clk [3164]));
Q_ASSIGN U13227 ( .B(clk), .A(\g.we_clk [3163]));
Q_ASSIGN U13228 ( .B(clk), .A(\g.we_clk [3162]));
Q_ASSIGN U13229 ( .B(clk), .A(\g.we_clk [3161]));
Q_ASSIGN U13230 ( .B(clk), .A(\g.we_clk [3160]));
Q_ASSIGN U13231 ( .B(clk), .A(\g.we_clk [3159]));
Q_ASSIGN U13232 ( .B(clk), .A(\g.we_clk [3158]));
Q_ASSIGN U13233 ( .B(clk), .A(\g.we_clk [3157]));
Q_ASSIGN U13234 ( .B(clk), .A(\g.we_clk [3156]));
Q_ASSIGN U13235 ( .B(clk), .A(\g.we_clk [3155]));
Q_ASSIGN U13236 ( .B(clk), .A(\g.we_clk [3154]));
Q_ASSIGN U13237 ( .B(clk), .A(\g.we_clk [3153]));
Q_ASSIGN U13238 ( .B(clk), .A(\g.we_clk [3152]));
Q_ASSIGN U13239 ( .B(clk), .A(\g.we_clk [3151]));
Q_ASSIGN U13240 ( .B(clk), .A(\g.we_clk [3150]));
Q_ASSIGN U13241 ( .B(clk), .A(\g.we_clk [3149]));
Q_ASSIGN U13242 ( .B(clk), .A(\g.we_clk [3148]));
Q_ASSIGN U13243 ( .B(clk), .A(\g.we_clk [3147]));
Q_ASSIGN U13244 ( .B(clk), .A(\g.we_clk [3146]));
Q_ASSIGN U13245 ( .B(clk), .A(\g.we_clk [3145]));
Q_ASSIGN U13246 ( .B(clk), .A(\g.we_clk [3144]));
Q_ASSIGN U13247 ( .B(clk), .A(\g.we_clk [3143]));
Q_ASSIGN U13248 ( .B(clk), .A(\g.we_clk [3142]));
Q_ASSIGN U13249 ( .B(clk), .A(\g.we_clk [3141]));
Q_ASSIGN U13250 ( .B(clk), .A(\g.we_clk [3140]));
Q_ASSIGN U13251 ( .B(clk), .A(\g.we_clk [3139]));
Q_ASSIGN U13252 ( .B(clk), .A(\g.we_clk [3138]));
Q_ASSIGN U13253 ( .B(clk), .A(\g.we_clk [3137]));
Q_ASSIGN U13254 ( .B(clk), .A(\g.we_clk [3136]));
Q_ASSIGN U13255 ( .B(clk), .A(\g.we_clk [3135]));
Q_ASSIGN U13256 ( .B(clk), .A(\g.we_clk [3134]));
Q_ASSIGN U13257 ( .B(clk), .A(\g.we_clk [3133]));
Q_ASSIGN U13258 ( .B(clk), .A(\g.we_clk [3132]));
Q_ASSIGN U13259 ( .B(clk), .A(\g.we_clk [3131]));
Q_ASSIGN U13260 ( .B(clk), .A(\g.we_clk [3130]));
Q_ASSIGN U13261 ( .B(clk), .A(\g.we_clk [3129]));
Q_ASSIGN U13262 ( .B(clk), .A(\g.we_clk [3128]));
Q_ASSIGN U13263 ( .B(clk), .A(\g.we_clk [3127]));
Q_ASSIGN U13264 ( .B(clk), .A(\g.we_clk [3126]));
Q_ASSIGN U13265 ( .B(clk), .A(\g.we_clk [3125]));
Q_ASSIGN U13266 ( .B(clk), .A(\g.we_clk [3124]));
Q_ASSIGN U13267 ( .B(clk), .A(\g.we_clk [3123]));
Q_ASSIGN U13268 ( .B(clk), .A(\g.we_clk [3122]));
Q_ASSIGN U13269 ( .B(clk), .A(\g.we_clk [3121]));
Q_ASSIGN U13270 ( .B(clk), .A(\g.we_clk [3120]));
Q_ASSIGN U13271 ( .B(clk), .A(\g.we_clk [3119]));
Q_ASSIGN U13272 ( .B(clk), .A(\g.we_clk [3118]));
Q_ASSIGN U13273 ( .B(clk), .A(\g.we_clk [3117]));
Q_ASSIGN U13274 ( .B(clk), .A(\g.we_clk [3116]));
Q_ASSIGN U13275 ( .B(clk), .A(\g.we_clk [3115]));
Q_ASSIGN U13276 ( .B(clk), .A(\g.we_clk [3114]));
Q_ASSIGN U13277 ( .B(clk), .A(\g.we_clk [3113]));
Q_ASSIGN U13278 ( .B(clk), .A(\g.we_clk [3112]));
Q_ASSIGN U13279 ( .B(clk), .A(\g.we_clk [3111]));
Q_ASSIGN U13280 ( .B(clk), .A(\g.we_clk [3110]));
Q_ASSIGN U13281 ( .B(clk), .A(\g.we_clk [3109]));
Q_ASSIGN U13282 ( .B(clk), .A(\g.we_clk [3108]));
Q_ASSIGN U13283 ( .B(clk), .A(\g.we_clk [3107]));
Q_ASSIGN U13284 ( .B(clk), .A(\g.we_clk [3106]));
Q_ASSIGN U13285 ( .B(clk), .A(\g.we_clk [3105]));
Q_ASSIGN U13286 ( .B(clk), .A(\g.we_clk [3104]));
Q_ASSIGN U13287 ( .B(clk), .A(\g.we_clk [3103]));
Q_ASSIGN U13288 ( .B(clk), .A(\g.we_clk [3102]));
Q_ASSIGN U13289 ( .B(clk), .A(\g.we_clk [3101]));
Q_ASSIGN U13290 ( .B(clk), .A(\g.we_clk [3100]));
Q_ASSIGN U13291 ( .B(clk), .A(\g.we_clk [3099]));
Q_ASSIGN U13292 ( .B(clk), .A(\g.we_clk [3098]));
Q_ASSIGN U13293 ( .B(clk), .A(\g.we_clk [3097]));
Q_ASSIGN U13294 ( .B(clk), .A(\g.we_clk [3096]));
Q_ASSIGN U13295 ( .B(clk), .A(\g.we_clk [3095]));
Q_ASSIGN U13296 ( .B(clk), .A(\g.we_clk [3094]));
Q_ASSIGN U13297 ( .B(clk), .A(\g.we_clk [3093]));
Q_ASSIGN U13298 ( .B(clk), .A(\g.we_clk [3092]));
Q_ASSIGN U13299 ( .B(clk), .A(\g.we_clk [3091]));
Q_ASSIGN U13300 ( .B(clk), .A(\g.we_clk [3090]));
Q_ASSIGN U13301 ( .B(clk), .A(\g.we_clk [3089]));
Q_ASSIGN U13302 ( .B(clk), .A(\g.we_clk [3088]));
Q_ASSIGN U13303 ( .B(clk), .A(\g.we_clk [3087]));
Q_ASSIGN U13304 ( .B(clk), .A(\g.we_clk [3086]));
Q_ASSIGN U13305 ( .B(clk), .A(\g.we_clk [3085]));
Q_ASSIGN U13306 ( .B(clk), .A(\g.we_clk [3084]));
Q_ASSIGN U13307 ( .B(clk), .A(\g.we_clk [3083]));
Q_ASSIGN U13308 ( .B(clk), .A(\g.we_clk [3082]));
Q_ASSIGN U13309 ( .B(clk), .A(\g.we_clk [3081]));
Q_ASSIGN U13310 ( .B(clk), .A(\g.we_clk [3080]));
Q_ASSIGN U13311 ( .B(clk), .A(\g.we_clk [3079]));
Q_ASSIGN U13312 ( .B(clk), .A(\g.we_clk [3078]));
Q_ASSIGN U13313 ( .B(clk), .A(\g.we_clk [3077]));
Q_ASSIGN U13314 ( .B(clk), .A(\g.we_clk [3076]));
Q_ASSIGN U13315 ( .B(clk), .A(\g.we_clk [3075]));
Q_ASSIGN U13316 ( .B(clk), .A(\g.we_clk [3074]));
Q_ASSIGN U13317 ( .B(clk), .A(\g.we_clk [3073]));
Q_ASSIGN U13318 ( .B(clk), .A(\g.we_clk [3072]));
Q_ASSIGN U13319 ( .B(clk), .A(\g.we_clk [3071]));
Q_ASSIGN U13320 ( .B(clk), .A(\g.we_clk [3070]));
Q_ASSIGN U13321 ( .B(clk), .A(\g.we_clk [3069]));
Q_ASSIGN U13322 ( .B(clk), .A(\g.we_clk [3068]));
Q_ASSIGN U13323 ( .B(clk), .A(\g.we_clk [3067]));
Q_ASSIGN U13324 ( .B(clk), .A(\g.we_clk [3066]));
Q_ASSIGN U13325 ( .B(clk), .A(\g.we_clk [3065]));
Q_ASSIGN U13326 ( .B(clk), .A(\g.we_clk [3064]));
Q_ASSIGN U13327 ( .B(clk), .A(\g.we_clk [3063]));
Q_ASSIGN U13328 ( .B(clk), .A(\g.we_clk [3062]));
Q_ASSIGN U13329 ( .B(clk), .A(\g.we_clk [3061]));
Q_ASSIGN U13330 ( .B(clk), .A(\g.we_clk [3060]));
Q_ASSIGN U13331 ( .B(clk), .A(\g.we_clk [3059]));
Q_ASSIGN U13332 ( .B(clk), .A(\g.we_clk [3058]));
Q_ASSIGN U13333 ( .B(clk), .A(\g.we_clk [3057]));
Q_ASSIGN U13334 ( .B(clk), .A(\g.we_clk [3056]));
Q_ASSIGN U13335 ( .B(clk), .A(\g.we_clk [3055]));
Q_ASSIGN U13336 ( .B(clk), .A(\g.we_clk [3054]));
Q_ASSIGN U13337 ( .B(clk), .A(\g.we_clk [3053]));
Q_ASSIGN U13338 ( .B(clk), .A(\g.we_clk [3052]));
Q_ASSIGN U13339 ( .B(clk), .A(\g.we_clk [3051]));
Q_ASSIGN U13340 ( .B(clk), .A(\g.we_clk [3050]));
Q_ASSIGN U13341 ( .B(clk), .A(\g.we_clk [3049]));
Q_ASSIGN U13342 ( .B(clk), .A(\g.we_clk [3048]));
Q_ASSIGN U13343 ( .B(clk), .A(\g.we_clk [3047]));
Q_ASSIGN U13344 ( .B(clk), .A(\g.we_clk [3046]));
Q_ASSIGN U13345 ( .B(clk), .A(\g.we_clk [3045]));
Q_ASSIGN U13346 ( .B(clk), .A(\g.we_clk [3044]));
Q_ASSIGN U13347 ( .B(clk), .A(\g.we_clk [3043]));
Q_ASSIGN U13348 ( .B(clk), .A(\g.we_clk [3042]));
Q_ASSIGN U13349 ( .B(clk), .A(\g.we_clk [3041]));
Q_ASSIGN U13350 ( .B(clk), .A(\g.we_clk [3040]));
Q_ASSIGN U13351 ( .B(clk), .A(\g.we_clk [3039]));
Q_ASSIGN U13352 ( .B(clk), .A(\g.we_clk [3038]));
Q_ASSIGN U13353 ( .B(clk), .A(\g.we_clk [3037]));
Q_ASSIGN U13354 ( .B(clk), .A(\g.we_clk [3036]));
Q_ASSIGN U13355 ( .B(clk), .A(\g.we_clk [3035]));
Q_ASSIGN U13356 ( .B(clk), .A(\g.we_clk [3034]));
Q_ASSIGN U13357 ( .B(clk), .A(\g.we_clk [3033]));
Q_ASSIGN U13358 ( .B(clk), .A(\g.we_clk [3032]));
Q_ASSIGN U13359 ( .B(clk), .A(\g.we_clk [3031]));
Q_ASSIGN U13360 ( .B(clk), .A(\g.we_clk [3030]));
Q_ASSIGN U13361 ( .B(clk), .A(\g.we_clk [3029]));
Q_ASSIGN U13362 ( .B(clk), .A(\g.we_clk [3028]));
Q_ASSIGN U13363 ( .B(clk), .A(\g.we_clk [3027]));
Q_ASSIGN U13364 ( .B(clk), .A(\g.we_clk [3026]));
Q_ASSIGN U13365 ( .B(clk), .A(\g.we_clk [3025]));
Q_ASSIGN U13366 ( .B(clk), .A(\g.we_clk [3024]));
Q_ASSIGN U13367 ( .B(clk), .A(\g.we_clk [3023]));
Q_ASSIGN U13368 ( .B(clk), .A(\g.we_clk [3022]));
Q_ASSIGN U13369 ( .B(clk), .A(\g.we_clk [3021]));
Q_ASSIGN U13370 ( .B(clk), .A(\g.we_clk [3020]));
Q_ASSIGN U13371 ( .B(clk), .A(\g.we_clk [3019]));
Q_ASSIGN U13372 ( .B(clk), .A(\g.we_clk [3018]));
Q_ASSIGN U13373 ( .B(clk), .A(\g.we_clk [3017]));
Q_ASSIGN U13374 ( .B(clk), .A(\g.we_clk [3016]));
Q_ASSIGN U13375 ( .B(clk), .A(\g.we_clk [3015]));
Q_ASSIGN U13376 ( .B(clk), .A(\g.we_clk [3014]));
Q_ASSIGN U13377 ( .B(clk), .A(\g.we_clk [3013]));
Q_ASSIGN U13378 ( .B(clk), .A(\g.we_clk [3012]));
Q_ASSIGN U13379 ( .B(clk), .A(\g.we_clk [3011]));
Q_ASSIGN U13380 ( .B(clk), .A(\g.we_clk [3010]));
Q_ASSIGN U13381 ( .B(clk), .A(\g.we_clk [3009]));
Q_ASSIGN U13382 ( .B(clk), .A(\g.we_clk [3008]));
Q_ASSIGN U13383 ( .B(clk), .A(\g.we_clk [3007]));
Q_ASSIGN U13384 ( .B(clk), .A(\g.we_clk [3006]));
Q_ASSIGN U13385 ( .B(clk), .A(\g.we_clk [3005]));
Q_ASSIGN U13386 ( .B(clk), .A(\g.we_clk [3004]));
Q_ASSIGN U13387 ( .B(clk), .A(\g.we_clk [3003]));
Q_ASSIGN U13388 ( .B(clk), .A(\g.we_clk [3002]));
Q_ASSIGN U13389 ( .B(clk), .A(\g.we_clk [3001]));
Q_ASSIGN U13390 ( .B(clk), .A(\g.we_clk [3000]));
Q_ASSIGN U13391 ( .B(clk), .A(\g.we_clk [2999]));
Q_ASSIGN U13392 ( .B(clk), .A(\g.we_clk [2998]));
Q_ASSIGN U13393 ( .B(clk), .A(\g.we_clk [2997]));
Q_ASSIGN U13394 ( .B(clk), .A(\g.we_clk [2996]));
Q_ASSIGN U13395 ( .B(clk), .A(\g.we_clk [2995]));
Q_ASSIGN U13396 ( .B(clk), .A(\g.we_clk [2994]));
Q_ASSIGN U13397 ( .B(clk), .A(\g.we_clk [2993]));
Q_ASSIGN U13398 ( .B(clk), .A(\g.we_clk [2992]));
Q_ASSIGN U13399 ( .B(clk), .A(\g.we_clk [2991]));
Q_ASSIGN U13400 ( .B(clk), .A(\g.we_clk [2990]));
Q_ASSIGN U13401 ( .B(clk), .A(\g.we_clk [2989]));
Q_ASSIGN U13402 ( .B(clk), .A(\g.we_clk [2988]));
Q_ASSIGN U13403 ( .B(clk), .A(\g.we_clk [2987]));
Q_ASSIGN U13404 ( .B(clk), .A(\g.we_clk [2986]));
Q_ASSIGN U13405 ( .B(clk), .A(\g.we_clk [2985]));
Q_ASSIGN U13406 ( .B(clk), .A(\g.we_clk [2984]));
Q_ASSIGN U13407 ( .B(clk), .A(\g.we_clk [2983]));
Q_ASSIGN U13408 ( .B(clk), .A(\g.we_clk [2982]));
Q_ASSIGN U13409 ( .B(clk), .A(\g.we_clk [2981]));
Q_ASSIGN U13410 ( .B(clk), .A(\g.we_clk [2980]));
Q_ASSIGN U13411 ( .B(clk), .A(\g.we_clk [2979]));
Q_ASSIGN U13412 ( .B(clk), .A(\g.we_clk [2978]));
Q_ASSIGN U13413 ( .B(clk), .A(\g.we_clk [2977]));
Q_ASSIGN U13414 ( .B(clk), .A(\g.we_clk [2976]));
Q_ASSIGN U13415 ( .B(clk), .A(\g.we_clk [2975]));
Q_ASSIGN U13416 ( .B(clk), .A(\g.we_clk [2974]));
Q_ASSIGN U13417 ( .B(clk), .A(\g.we_clk [2973]));
Q_ASSIGN U13418 ( .B(clk), .A(\g.we_clk [2972]));
Q_ASSIGN U13419 ( .B(clk), .A(\g.we_clk [2971]));
Q_ASSIGN U13420 ( .B(clk), .A(\g.we_clk [2970]));
Q_ASSIGN U13421 ( .B(clk), .A(\g.we_clk [2969]));
Q_ASSIGN U13422 ( .B(clk), .A(\g.we_clk [2968]));
Q_ASSIGN U13423 ( .B(clk), .A(\g.we_clk [2967]));
Q_ASSIGN U13424 ( .B(clk), .A(\g.we_clk [2966]));
Q_ASSIGN U13425 ( .B(clk), .A(\g.we_clk [2965]));
Q_ASSIGN U13426 ( .B(clk), .A(\g.we_clk [2964]));
Q_ASSIGN U13427 ( .B(clk), .A(\g.we_clk [2963]));
Q_ASSIGN U13428 ( .B(clk), .A(\g.we_clk [2962]));
Q_ASSIGN U13429 ( .B(clk), .A(\g.we_clk [2961]));
Q_ASSIGN U13430 ( .B(clk), .A(\g.we_clk [2960]));
Q_ASSIGN U13431 ( .B(clk), .A(\g.we_clk [2959]));
Q_ASSIGN U13432 ( .B(clk), .A(\g.we_clk [2958]));
Q_ASSIGN U13433 ( .B(clk), .A(\g.we_clk [2957]));
Q_ASSIGN U13434 ( .B(clk), .A(\g.we_clk [2956]));
Q_ASSIGN U13435 ( .B(clk), .A(\g.we_clk [2955]));
Q_ASSIGN U13436 ( .B(clk), .A(\g.we_clk [2954]));
Q_ASSIGN U13437 ( .B(clk), .A(\g.we_clk [2953]));
Q_ASSIGN U13438 ( .B(clk), .A(\g.we_clk [2952]));
Q_ASSIGN U13439 ( .B(clk), .A(\g.we_clk [2951]));
Q_ASSIGN U13440 ( .B(clk), .A(\g.we_clk [2950]));
Q_ASSIGN U13441 ( .B(clk), .A(\g.we_clk [2949]));
Q_ASSIGN U13442 ( .B(clk), .A(\g.we_clk [2948]));
Q_ASSIGN U13443 ( .B(clk), .A(\g.we_clk [2947]));
Q_ASSIGN U13444 ( .B(clk), .A(\g.we_clk [2946]));
Q_ASSIGN U13445 ( .B(clk), .A(\g.we_clk [2945]));
Q_ASSIGN U13446 ( .B(clk), .A(\g.we_clk [2944]));
Q_ASSIGN U13447 ( .B(clk), .A(\g.we_clk [2943]));
Q_ASSIGN U13448 ( .B(clk), .A(\g.we_clk [2942]));
Q_ASSIGN U13449 ( .B(clk), .A(\g.we_clk [2941]));
Q_ASSIGN U13450 ( .B(clk), .A(\g.we_clk [2940]));
Q_ASSIGN U13451 ( .B(clk), .A(\g.we_clk [2939]));
Q_ASSIGN U13452 ( .B(clk), .A(\g.we_clk [2938]));
Q_ASSIGN U13453 ( .B(clk), .A(\g.we_clk [2937]));
Q_ASSIGN U13454 ( .B(clk), .A(\g.we_clk [2936]));
Q_ASSIGN U13455 ( .B(clk), .A(\g.we_clk [2935]));
Q_ASSIGN U13456 ( .B(clk), .A(\g.we_clk [2934]));
Q_ASSIGN U13457 ( .B(clk), .A(\g.we_clk [2933]));
Q_ASSIGN U13458 ( .B(clk), .A(\g.we_clk [2932]));
Q_ASSIGN U13459 ( .B(clk), .A(\g.we_clk [2931]));
Q_ASSIGN U13460 ( .B(clk), .A(\g.we_clk [2930]));
Q_ASSIGN U13461 ( .B(clk), .A(\g.we_clk [2929]));
Q_ASSIGN U13462 ( .B(clk), .A(\g.we_clk [2928]));
Q_ASSIGN U13463 ( .B(clk), .A(\g.we_clk [2927]));
Q_ASSIGN U13464 ( .B(clk), .A(\g.we_clk [2926]));
Q_ASSIGN U13465 ( .B(clk), .A(\g.we_clk [2925]));
Q_ASSIGN U13466 ( .B(clk), .A(\g.we_clk [2924]));
Q_ASSIGN U13467 ( .B(clk), .A(\g.we_clk [2923]));
Q_ASSIGN U13468 ( .B(clk), .A(\g.we_clk [2922]));
Q_ASSIGN U13469 ( .B(clk), .A(\g.we_clk [2921]));
Q_ASSIGN U13470 ( .B(clk), .A(\g.we_clk [2920]));
Q_ASSIGN U13471 ( .B(clk), .A(\g.we_clk [2919]));
Q_ASSIGN U13472 ( .B(clk), .A(\g.we_clk [2918]));
Q_ASSIGN U13473 ( .B(clk), .A(\g.we_clk [2917]));
Q_ASSIGN U13474 ( .B(clk), .A(\g.we_clk [2916]));
Q_ASSIGN U13475 ( .B(clk), .A(\g.we_clk [2915]));
Q_ASSIGN U13476 ( .B(clk), .A(\g.we_clk [2914]));
Q_ASSIGN U13477 ( .B(clk), .A(\g.we_clk [2913]));
Q_ASSIGN U13478 ( .B(clk), .A(\g.we_clk [2912]));
Q_ASSIGN U13479 ( .B(clk), .A(\g.we_clk [2911]));
Q_ASSIGN U13480 ( .B(clk), .A(\g.we_clk [2910]));
Q_ASSIGN U13481 ( .B(clk), .A(\g.we_clk [2909]));
Q_ASSIGN U13482 ( .B(clk), .A(\g.we_clk [2908]));
Q_ASSIGN U13483 ( .B(clk), .A(\g.we_clk [2907]));
Q_ASSIGN U13484 ( .B(clk), .A(\g.we_clk [2906]));
Q_ASSIGN U13485 ( .B(clk), .A(\g.we_clk [2905]));
Q_ASSIGN U13486 ( .B(clk), .A(\g.we_clk [2904]));
Q_ASSIGN U13487 ( .B(clk), .A(\g.we_clk [2903]));
Q_ASSIGN U13488 ( .B(clk), .A(\g.we_clk [2902]));
Q_ASSIGN U13489 ( .B(clk), .A(\g.we_clk [2901]));
Q_ASSIGN U13490 ( .B(clk), .A(\g.we_clk [2900]));
Q_ASSIGN U13491 ( .B(clk), .A(\g.we_clk [2899]));
Q_ASSIGN U13492 ( .B(clk), .A(\g.we_clk [2898]));
Q_ASSIGN U13493 ( .B(clk), .A(\g.we_clk [2897]));
Q_ASSIGN U13494 ( .B(clk), .A(\g.we_clk [2896]));
Q_ASSIGN U13495 ( .B(clk), .A(\g.we_clk [2895]));
Q_ASSIGN U13496 ( .B(clk), .A(\g.we_clk [2894]));
Q_ASSIGN U13497 ( .B(clk), .A(\g.we_clk [2893]));
Q_ASSIGN U13498 ( .B(clk), .A(\g.we_clk [2892]));
Q_ASSIGN U13499 ( .B(clk), .A(\g.we_clk [2891]));
Q_ASSIGN U13500 ( .B(clk), .A(\g.we_clk [2890]));
Q_ASSIGN U13501 ( .B(clk), .A(\g.we_clk [2889]));
Q_ASSIGN U13502 ( .B(clk), .A(\g.we_clk [2888]));
Q_ASSIGN U13503 ( .B(clk), .A(\g.we_clk [2887]));
Q_ASSIGN U13504 ( .B(clk), .A(\g.we_clk [2886]));
Q_ASSIGN U13505 ( .B(clk), .A(\g.we_clk [2885]));
Q_ASSIGN U13506 ( .B(clk), .A(\g.we_clk [2884]));
Q_ASSIGN U13507 ( .B(clk), .A(\g.we_clk [2883]));
Q_ASSIGN U13508 ( .B(clk), .A(\g.we_clk [2882]));
Q_ASSIGN U13509 ( .B(clk), .A(\g.we_clk [2881]));
Q_ASSIGN U13510 ( .B(clk), .A(\g.we_clk [2880]));
Q_ASSIGN U13511 ( .B(clk), .A(\g.we_clk [2879]));
Q_ASSIGN U13512 ( .B(clk), .A(\g.we_clk [2878]));
Q_ASSIGN U13513 ( .B(clk), .A(\g.we_clk [2877]));
Q_ASSIGN U13514 ( .B(clk), .A(\g.we_clk [2876]));
Q_ASSIGN U13515 ( .B(clk), .A(\g.we_clk [2875]));
Q_ASSIGN U13516 ( .B(clk), .A(\g.we_clk [2874]));
Q_ASSIGN U13517 ( .B(clk), .A(\g.we_clk [2873]));
Q_ASSIGN U13518 ( .B(clk), .A(\g.we_clk [2872]));
Q_ASSIGN U13519 ( .B(clk), .A(\g.we_clk [2871]));
Q_ASSIGN U13520 ( .B(clk), .A(\g.we_clk [2870]));
Q_ASSIGN U13521 ( .B(clk), .A(\g.we_clk [2869]));
Q_ASSIGN U13522 ( .B(clk), .A(\g.we_clk [2868]));
Q_ASSIGN U13523 ( .B(clk), .A(\g.we_clk [2867]));
Q_ASSIGN U13524 ( .B(clk), .A(\g.we_clk [2866]));
Q_ASSIGN U13525 ( .B(clk), .A(\g.we_clk [2865]));
Q_ASSIGN U13526 ( .B(clk), .A(\g.we_clk [2864]));
Q_ASSIGN U13527 ( .B(clk), .A(\g.we_clk [2863]));
Q_ASSIGN U13528 ( .B(clk), .A(\g.we_clk [2862]));
Q_ASSIGN U13529 ( .B(clk), .A(\g.we_clk [2861]));
Q_ASSIGN U13530 ( .B(clk), .A(\g.we_clk [2860]));
Q_ASSIGN U13531 ( .B(clk), .A(\g.we_clk [2859]));
Q_ASSIGN U13532 ( .B(clk), .A(\g.we_clk [2858]));
Q_ASSIGN U13533 ( .B(clk), .A(\g.we_clk [2857]));
Q_ASSIGN U13534 ( .B(clk), .A(\g.we_clk [2856]));
Q_ASSIGN U13535 ( .B(clk), .A(\g.we_clk [2855]));
Q_ASSIGN U13536 ( .B(clk), .A(\g.we_clk [2854]));
Q_ASSIGN U13537 ( .B(clk), .A(\g.we_clk [2853]));
Q_ASSIGN U13538 ( .B(clk), .A(\g.we_clk [2852]));
Q_ASSIGN U13539 ( .B(clk), .A(\g.we_clk [2851]));
Q_ASSIGN U13540 ( .B(clk), .A(\g.we_clk [2850]));
Q_ASSIGN U13541 ( .B(clk), .A(\g.we_clk [2849]));
Q_ASSIGN U13542 ( .B(clk), .A(\g.we_clk [2848]));
Q_ASSIGN U13543 ( .B(clk), .A(\g.we_clk [2847]));
Q_ASSIGN U13544 ( .B(clk), .A(\g.we_clk [2846]));
Q_ASSIGN U13545 ( .B(clk), .A(\g.we_clk [2845]));
Q_ASSIGN U13546 ( .B(clk), .A(\g.we_clk [2844]));
Q_ASSIGN U13547 ( .B(clk), .A(\g.we_clk [2843]));
Q_ASSIGN U13548 ( .B(clk), .A(\g.we_clk [2842]));
Q_ASSIGN U13549 ( .B(clk), .A(\g.we_clk [2841]));
Q_ASSIGN U13550 ( .B(clk), .A(\g.we_clk [2840]));
Q_ASSIGN U13551 ( .B(clk), .A(\g.we_clk [2839]));
Q_ASSIGN U13552 ( .B(clk), .A(\g.we_clk [2838]));
Q_ASSIGN U13553 ( .B(clk), .A(\g.we_clk [2837]));
Q_ASSIGN U13554 ( .B(clk), .A(\g.we_clk [2836]));
Q_ASSIGN U13555 ( .B(clk), .A(\g.we_clk [2835]));
Q_ASSIGN U13556 ( .B(clk), .A(\g.we_clk [2834]));
Q_ASSIGN U13557 ( .B(clk), .A(\g.we_clk [2833]));
Q_ASSIGN U13558 ( .B(clk), .A(\g.we_clk [2832]));
Q_ASSIGN U13559 ( .B(clk), .A(\g.we_clk [2831]));
Q_ASSIGN U13560 ( .B(clk), .A(\g.we_clk [2830]));
Q_ASSIGN U13561 ( .B(clk), .A(\g.we_clk [2829]));
Q_ASSIGN U13562 ( .B(clk), .A(\g.we_clk [2828]));
Q_ASSIGN U13563 ( .B(clk), .A(\g.we_clk [2827]));
Q_ASSIGN U13564 ( .B(clk), .A(\g.we_clk [2826]));
Q_ASSIGN U13565 ( .B(clk), .A(\g.we_clk [2825]));
Q_ASSIGN U13566 ( .B(clk), .A(\g.we_clk [2824]));
Q_ASSIGN U13567 ( .B(clk), .A(\g.we_clk [2823]));
Q_ASSIGN U13568 ( .B(clk), .A(\g.we_clk [2822]));
Q_ASSIGN U13569 ( .B(clk), .A(\g.we_clk [2821]));
Q_ASSIGN U13570 ( .B(clk), .A(\g.we_clk [2820]));
Q_ASSIGN U13571 ( .B(clk), .A(\g.we_clk [2819]));
Q_ASSIGN U13572 ( .B(clk), .A(\g.we_clk [2818]));
Q_ASSIGN U13573 ( .B(clk), .A(\g.we_clk [2817]));
Q_ASSIGN U13574 ( .B(clk), .A(\g.we_clk [2816]));
Q_ASSIGN U13575 ( .B(clk), .A(\g.we_clk [2815]));
Q_ASSIGN U13576 ( .B(clk), .A(\g.we_clk [2814]));
Q_ASSIGN U13577 ( .B(clk), .A(\g.we_clk [2813]));
Q_ASSIGN U13578 ( .B(clk), .A(\g.we_clk [2812]));
Q_ASSIGN U13579 ( .B(clk), .A(\g.we_clk [2811]));
Q_ASSIGN U13580 ( .B(clk), .A(\g.we_clk [2810]));
Q_ASSIGN U13581 ( .B(clk), .A(\g.we_clk [2809]));
Q_ASSIGN U13582 ( .B(clk), .A(\g.we_clk [2808]));
Q_ASSIGN U13583 ( .B(clk), .A(\g.we_clk [2807]));
Q_ASSIGN U13584 ( .B(clk), .A(\g.we_clk [2806]));
Q_ASSIGN U13585 ( .B(clk), .A(\g.we_clk [2805]));
Q_ASSIGN U13586 ( .B(clk), .A(\g.we_clk [2804]));
Q_ASSIGN U13587 ( .B(clk), .A(\g.we_clk [2803]));
Q_ASSIGN U13588 ( .B(clk), .A(\g.we_clk [2802]));
Q_ASSIGN U13589 ( .B(clk), .A(\g.we_clk [2801]));
Q_ASSIGN U13590 ( .B(clk), .A(\g.we_clk [2800]));
Q_ASSIGN U13591 ( .B(clk), .A(\g.we_clk [2799]));
Q_ASSIGN U13592 ( .B(clk), .A(\g.we_clk [2798]));
Q_ASSIGN U13593 ( .B(clk), .A(\g.we_clk [2797]));
Q_ASSIGN U13594 ( .B(clk), .A(\g.we_clk [2796]));
Q_ASSIGN U13595 ( .B(clk), .A(\g.we_clk [2795]));
Q_ASSIGN U13596 ( .B(clk), .A(\g.we_clk [2794]));
Q_ASSIGN U13597 ( .B(clk), .A(\g.we_clk [2793]));
Q_ASSIGN U13598 ( .B(clk), .A(\g.we_clk [2792]));
Q_ASSIGN U13599 ( .B(clk), .A(\g.we_clk [2791]));
Q_ASSIGN U13600 ( .B(clk), .A(\g.we_clk [2790]));
Q_ASSIGN U13601 ( .B(clk), .A(\g.we_clk [2789]));
Q_ASSIGN U13602 ( .B(clk), .A(\g.we_clk [2788]));
Q_ASSIGN U13603 ( .B(clk), .A(\g.we_clk [2787]));
Q_ASSIGN U13604 ( .B(clk), .A(\g.we_clk [2786]));
Q_ASSIGN U13605 ( .B(clk), .A(\g.we_clk [2785]));
Q_ASSIGN U13606 ( .B(clk), .A(\g.we_clk [2784]));
Q_ASSIGN U13607 ( .B(clk), .A(\g.we_clk [2783]));
Q_ASSIGN U13608 ( .B(clk), .A(\g.we_clk [2782]));
Q_ASSIGN U13609 ( .B(clk), .A(\g.we_clk [2781]));
Q_ASSIGN U13610 ( .B(clk), .A(\g.we_clk [2780]));
Q_ASSIGN U13611 ( .B(clk), .A(\g.we_clk [2779]));
Q_ASSIGN U13612 ( .B(clk), .A(\g.we_clk [2778]));
Q_ASSIGN U13613 ( .B(clk), .A(\g.we_clk [2777]));
Q_ASSIGN U13614 ( .B(clk), .A(\g.we_clk [2776]));
Q_ASSIGN U13615 ( .B(clk), .A(\g.we_clk [2775]));
Q_ASSIGN U13616 ( .B(clk), .A(\g.we_clk [2774]));
Q_ASSIGN U13617 ( .B(clk), .A(\g.we_clk [2773]));
Q_ASSIGN U13618 ( .B(clk), .A(\g.we_clk [2772]));
Q_ASSIGN U13619 ( .B(clk), .A(\g.we_clk [2771]));
Q_ASSIGN U13620 ( .B(clk), .A(\g.we_clk [2770]));
Q_ASSIGN U13621 ( .B(clk), .A(\g.we_clk [2769]));
Q_ASSIGN U13622 ( .B(clk), .A(\g.we_clk [2768]));
Q_ASSIGN U13623 ( .B(clk), .A(\g.we_clk [2767]));
Q_ASSIGN U13624 ( .B(clk), .A(\g.we_clk [2766]));
Q_ASSIGN U13625 ( .B(clk), .A(\g.we_clk [2765]));
Q_ASSIGN U13626 ( .B(clk), .A(\g.we_clk [2764]));
Q_ASSIGN U13627 ( .B(clk), .A(\g.we_clk [2763]));
Q_ASSIGN U13628 ( .B(clk), .A(\g.we_clk [2762]));
Q_ASSIGN U13629 ( .B(clk), .A(\g.we_clk [2761]));
Q_ASSIGN U13630 ( .B(clk), .A(\g.we_clk [2760]));
Q_ASSIGN U13631 ( .B(clk), .A(\g.we_clk [2759]));
Q_ASSIGN U13632 ( .B(clk), .A(\g.we_clk [2758]));
Q_ASSIGN U13633 ( .B(clk), .A(\g.we_clk [2757]));
Q_ASSIGN U13634 ( .B(clk), .A(\g.we_clk [2756]));
Q_ASSIGN U13635 ( .B(clk), .A(\g.we_clk [2755]));
Q_ASSIGN U13636 ( .B(clk), .A(\g.we_clk [2754]));
Q_ASSIGN U13637 ( .B(clk), .A(\g.we_clk [2753]));
Q_ASSIGN U13638 ( .B(clk), .A(\g.we_clk [2752]));
Q_ASSIGN U13639 ( .B(clk), .A(\g.we_clk [2751]));
Q_ASSIGN U13640 ( .B(clk), .A(\g.we_clk [2750]));
Q_ASSIGN U13641 ( .B(clk), .A(\g.we_clk [2749]));
Q_ASSIGN U13642 ( .B(clk), .A(\g.we_clk [2748]));
Q_ASSIGN U13643 ( .B(clk), .A(\g.we_clk [2747]));
Q_ASSIGN U13644 ( .B(clk), .A(\g.we_clk [2746]));
Q_ASSIGN U13645 ( .B(clk), .A(\g.we_clk [2745]));
Q_ASSIGN U13646 ( .B(clk), .A(\g.we_clk [2744]));
Q_ASSIGN U13647 ( .B(clk), .A(\g.we_clk [2743]));
Q_ASSIGN U13648 ( .B(clk), .A(\g.we_clk [2742]));
Q_ASSIGN U13649 ( .B(clk), .A(\g.we_clk [2741]));
Q_ASSIGN U13650 ( .B(clk), .A(\g.we_clk [2740]));
Q_ASSIGN U13651 ( .B(clk), .A(\g.we_clk [2739]));
Q_ASSIGN U13652 ( .B(clk), .A(\g.we_clk [2738]));
Q_ASSIGN U13653 ( .B(clk), .A(\g.we_clk [2737]));
Q_ASSIGN U13654 ( .B(clk), .A(\g.we_clk [2736]));
Q_ASSIGN U13655 ( .B(clk), .A(\g.we_clk [2735]));
Q_ASSIGN U13656 ( .B(clk), .A(\g.we_clk [2734]));
Q_ASSIGN U13657 ( .B(clk), .A(\g.we_clk [2733]));
Q_ASSIGN U13658 ( .B(clk), .A(\g.we_clk [2732]));
Q_ASSIGN U13659 ( .B(clk), .A(\g.we_clk [2731]));
Q_ASSIGN U13660 ( .B(clk), .A(\g.we_clk [2730]));
Q_ASSIGN U13661 ( .B(clk), .A(\g.we_clk [2729]));
Q_ASSIGN U13662 ( .B(clk), .A(\g.we_clk [2728]));
Q_ASSIGN U13663 ( .B(clk), .A(\g.we_clk [2727]));
Q_ASSIGN U13664 ( .B(clk), .A(\g.we_clk [2726]));
Q_ASSIGN U13665 ( .B(clk), .A(\g.we_clk [2725]));
Q_ASSIGN U13666 ( .B(clk), .A(\g.we_clk [2724]));
Q_ASSIGN U13667 ( .B(clk), .A(\g.we_clk [2723]));
Q_ASSIGN U13668 ( .B(clk), .A(\g.we_clk [2722]));
Q_ASSIGN U13669 ( .B(clk), .A(\g.we_clk [2721]));
Q_ASSIGN U13670 ( .B(clk), .A(\g.we_clk [2720]));
Q_ASSIGN U13671 ( .B(clk), .A(\g.we_clk [2719]));
Q_ASSIGN U13672 ( .B(clk), .A(\g.we_clk [2718]));
Q_ASSIGN U13673 ( .B(clk), .A(\g.we_clk [2717]));
Q_ASSIGN U13674 ( .B(clk), .A(\g.we_clk [2716]));
Q_ASSIGN U13675 ( .B(clk), .A(\g.we_clk [2715]));
Q_ASSIGN U13676 ( .B(clk), .A(\g.we_clk [2714]));
Q_ASSIGN U13677 ( .B(clk), .A(\g.we_clk [2713]));
Q_ASSIGN U13678 ( .B(clk), .A(\g.we_clk [2712]));
Q_ASSIGN U13679 ( .B(clk), .A(\g.we_clk [2711]));
Q_ASSIGN U13680 ( .B(clk), .A(\g.we_clk [2710]));
Q_ASSIGN U13681 ( .B(clk), .A(\g.we_clk [2709]));
Q_ASSIGN U13682 ( .B(clk), .A(\g.we_clk [2708]));
Q_ASSIGN U13683 ( .B(clk), .A(\g.we_clk [2707]));
Q_ASSIGN U13684 ( .B(clk), .A(\g.we_clk [2706]));
Q_ASSIGN U13685 ( .B(clk), .A(\g.we_clk [2705]));
Q_ASSIGN U13686 ( .B(clk), .A(\g.we_clk [2704]));
Q_ASSIGN U13687 ( .B(clk), .A(\g.we_clk [2703]));
Q_ASSIGN U13688 ( .B(clk), .A(\g.we_clk [2702]));
Q_ASSIGN U13689 ( .B(clk), .A(\g.we_clk [2701]));
Q_ASSIGN U13690 ( .B(clk), .A(\g.we_clk [2700]));
Q_ASSIGN U13691 ( .B(clk), .A(\g.we_clk [2699]));
Q_ASSIGN U13692 ( .B(clk), .A(\g.we_clk [2698]));
Q_ASSIGN U13693 ( .B(clk), .A(\g.we_clk [2697]));
Q_ASSIGN U13694 ( .B(clk), .A(\g.we_clk [2696]));
Q_ASSIGN U13695 ( .B(clk), .A(\g.we_clk [2695]));
Q_ASSIGN U13696 ( .B(clk), .A(\g.we_clk [2694]));
Q_ASSIGN U13697 ( .B(clk), .A(\g.we_clk [2693]));
Q_ASSIGN U13698 ( .B(clk), .A(\g.we_clk [2692]));
Q_ASSIGN U13699 ( .B(clk), .A(\g.we_clk [2691]));
Q_ASSIGN U13700 ( .B(clk), .A(\g.we_clk [2690]));
Q_ASSIGN U13701 ( .B(clk), .A(\g.we_clk [2689]));
Q_ASSIGN U13702 ( .B(clk), .A(\g.we_clk [2688]));
Q_ASSIGN U13703 ( .B(clk), .A(\g.we_clk [2687]));
Q_ASSIGN U13704 ( .B(clk), .A(\g.we_clk [2686]));
Q_ASSIGN U13705 ( .B(clk), .A(\g.we_clk [2685]));
Q_ASSIGN U13706 ( .B(clk), .A(\g.we_clk [2684]));
Q_ASSIGN U13707 ( .B(clk), .A(\g.we_clk [2683]));
Q_ASSIGN U13708 ( .B(clk), .A(\g.we_clk [2682]));
Q_ASSIGN U13709 ( .B(clk), .A(\g.we_clk [2681]));
Q_ASSIGN U13710 ( .B(clk), .A(\g.we_clk [2680]));
Q_ASSIGN U13711 ( .B(clk), .A(\g.we_clk [2679]));
Q_ASSIGN U13712 ( .B(clk), .A(\g.we_clk [2678]));
Q_ASSIGN U13713 ( .B(clk), .A(\g.we_clk [2677]));
Q_ASSIGN U13714 ( .B(clk), .A(\g.we_clk [2676]));
Q_ASSIGN U13715 ( .B(clk), .A(\g.we_clk [2675]));
Q_ASSIGN U13716 ( .B(clk), .A(\g.we_clk [2674]));
Q_ASSIGN U13717 ( .B(clk), .A(\g.we_clk [2673]));
Q_ASSIGN U13718 ( .B(clk), .A(\g.we_clk [2672]));
Q_ASSIGN U13719 ( .B(clk), .A(\g.we_clk [2671]));
Q_ASSIGN U13720 ( .B(clk), .A(\g.we_clk [2670]));
Q_ASSIGN U13721 ( .B(clk), .A(\g.we_clk [2669]));
Q_ASSIGN U13722 ( .B(clk), .A(\g.we_clk [2668]));
Q_ASSIGN U13723 ( .B(clk), .A(\g.we_clk [2667]));
Q_ASSIGN U13724 ( .B(clk), .A(\g.we_clk [2666]));
Q_ASSIGN U13725 ( .B(clk), .A(\g.we_clk [2665]));
Q_ASSIGN U13726 ( .B(clk), .A(\g.we_clk [2664]));
Q_ASSIGN U13727 ( .B(clk), .A(\g.we_clk [2663]));
Q_ASSIGN U13728 ( .B(clk), .A(\g.we_clk [2662]));
Q_ASSIGN U13729 ( .B(clk), .A(\g.we_clk [2661]));
Q_ASSIGN U13730 ( .B(clk), .A(\g.we_clk [2660]));
Q_ASSIGN U13731 ( .B(clk), .A(\g.we_clk [2659]));
Q_ASSIGN U13732 ( .B(clk), .A(\g.we_clk [2658]));
Q_ASSIGN U13733 ( .B(clk), .A(\g.we_clk [2657]));
Q_ASSIGN U13734 ( .B(clk), .A(\g.we_clk [2656]));
Q_ASSIGN U13735 ( .B(clk), .A(\g.we_clk [2655]));
Q_ASSIGN U13736 ( .B(clk), .A(\g.we_clk [2654]));
Q_ASSIGN U13737 ( .B(clk), .A(\g.we_clk [2653]));
Q_ASSIGN U13738 ( .B(clk), .A(\g.we_clk [2652]));
Q_ASSIGN U13739 ( .B(clk), .A(\g.we_clk [2651]));
Q_ASSIGN U13740 ( .B(clk), .A(\g.we_clk [2650]));
Q_ASSIGN U13741 ( .B(clk), .A(\g.we_clk [2649]));
Q_ASSIGN U13742 ( .B(clk), .A(\g.we_clk [2648]));
Q_ASSIGN U13743 ( .B(clk), .A(\g.we_clk [2647]));
Q_ASSIGN U13744 ( .B(clk), .A(\g.we_clk [2646]));
Q_ASSIGN U13745 ( .B(clk), .A(\g.we_clk [2645]));
Q_ASSIGN U13746 ( .B(clk), .A(\g.we_clk [2644]));
Q_ASSIGN U13747 ( .B(clk), .A(\g.we_clk [2643]));
Q_ASSIGN U13748 ( .B(clk), .A(\g.we_clk [2642]));
Q_ASSIGN U13749 ( .B(clk), .A(\g.we_clk [2641]));
Q_ASSIGN U13750 ( .B(clk), .A(\g.we_clk [2640]));
Q_ASSIGN U13751 ( .B(clk), .A(\g.we_clk [2639]));
Q_ASSIGN U13752 ( .B(clk), .A(\g.we_clk [2638]));
Q_ASSIGN U13753 ( .B(clk), .A(\g.we_clk [2637]));
Q_ASSIGN U13754 ( .B(clk), .A(\g.we_clk [2636]));
Q_ASSIGN U13755 ( .B(clk), .A(\g.we_clk [2635]));
Q_ASSIGN U13756 ( .B(clk), .A(\g.we_clk [2634]));
Q_ASSIGN U13757 ( .B(clk), .A(\g.we_clk [2633]));
Q_ASSIGN U13758 ( .B(clk), .A(\g.we_clk [2632]));
Q_ASSIGN U13759 ( .B(clk), .A(\g.we_clk [2631]));
Q_ASSIGN U13760 ( .B(clk), .A(\g.we_clk [2630]));
Q_ASSIGN U13761 ( .B(clk), .A(\g.we_clk [2629]));
Q_ASSIGN U13762 ( .B(clk), .A(\g.we_clk [2628]));
Q_ASSIGN U13763 ( .B(clk), .A(\g.we_clk [2627]));
Q_ASSIGN U13764 ( .B(clk), .A(\g.we_clk [2626]));
Q_ASSIGN U13765 ( .B(clk), .A(\g.we_clk [2625]));
Q_ASSIGN U13766 ( .B(clk), .A(\g.we_clk [2624]));
Q_ASSIGN U13767 ( .B(clk), .A(\g.we_clk [2623]));
Q_ASSIGN U13768 ( .B(clk), .A(\g.we_clk [2622]));
Q_ASSIGN U13769 ( .B(clk), .A(\g.we_clk [2621]));
Q_ASSIGN U13770 ( .B(clk), .A(\g.we_clk [2620]));
Q_ASSIGN U13771 ( .B(clk), .A(\g.we_clk [2619]));
Q_ASSIGN U13772 ( .B(clk), .A(\g.we_clk [2618]));
Q_ASSIGN U13773 ( .B(clk), .A(\g.we_clk [2617]));
Q_ASSIGN U13774 ( .B(clk), .A(\g.we_clk [2616]));
Q_ASSIGN U13775 ( .B(clk), .A(\g.we_clk [2615]));
Q_ASSIGN U13776 ( .B(clk), .A(\g.we_clk [2614]));
Q_ASSIGN U13777 ( .B(clk), .A(\g.we_clk [2613]));
Q_ASSIGN U13778 ( .B(clk), .A(\g.we_clk [2612]));
Q_ASSIGN U13779 ( .B(clk), .A(\g.we_clk [2611]));
Q_ASSIGN U13780 ( .B(clk), .A(\g.we_clk [2610]));
Q_ASSIGN U13781 ( .B(clk), .A(\g.we_clk [2609]));
Q_ASSIGN U13782 ( .B(clk), .A(\g.we_clk [2608]));
Q_ASSIGN U13783 ( .B(clk), .A(\g.we_clk [2607]));
Q_ASSIGN U13784 ( .B(clk), .A(\g.we_clk [2606]));
Q_ASSIGN U13785 ( .B(clk), .A(\g.we_clk [2605]));
Q_ASSIGN U13786 ( .B(clk), .A(\g.we_clk [2604]));
Q_ASSIGN U13787 ( .B(clk), .A(\g.we_clk [2603]));
Q_ASSIGN U13788 ( .B(clk), .A(\g.we_clk [2602]));
Q_ASSIGN U13789 ( .B(clk), .A(\g.we_clk [2601]));
Q_ASSIGN U13790 ( .B(clk), .A(\g.we_clk [2600]));
Q_ASSIGN U13791 ( .B(clk), .A(\g.we_clk [2599]));
Q_ASSIGN U13792 ( .B(clk), .A(\g.we_clk [2598]));
Q_ASSIGN U13793 ( .B(clk), .A(\g.we_clk [2597]));
Q_ASSIGN U13794 ( .B(clk), .A(\g.we_clk [2596]));
Q_ASSIGN U13795 ( .B(clk), .A(\g.we_clk [2595]));
Q_ASSIGN U13796 ( .B(clk), .A(\g.we_clk [2594]));
Q_ASSIGN U13797 ( .B(clk), .A(\g.we_clk [2593]));
Q_ASSIGN U13798 ( .B(clk), .A(\g.we_clk [2592]));
Q_ASSIGN U13799 ( .B(clk), .A(\g.we_clk [2591]));
Q_ASSIGN U13800 ( .B(clk), .A(\g.we_clk [2590]));
Q_ASSIGN U13801 ( .B(clk), .A(\g.we_clk [2589]));
Q_ASSIGN U13802 ( .B(clk), .A(\g.we_clk [2588]));
Q_ASSIGN U13803 ( .B(clk), .A(\g.we_clk [2587]));
Q_ASSIGN U13804 ( .B(clk), .A(\g.we_clk [2586]));
Q_ASSIGN U13805 ( .B(clk), .A(\g.we_clk [2585]));
Q_ASSIGN U13806 ( .B(clk), .A(\g.we_clk [2584]));
Q_ASSIGN U13807 ( .B(clk), .A(\g.we_clk [2583]));
Q_ASSIGN U13808 ( .B(clk), .A(\g.we_clk [2582]));
Q_ASSIGN U13809 ( .B(clk), .A(\g.we_clk [2581]));
Q_ASSIGN U13810 ( .B(clk), .A(\g.we_clk [2580]));
Q_ASSIGN U13811 ( .B(clk), .A(\g.we_clk [2579]));
Q_ASSIGN U13812 ( .B(clk), .A(\g.we_clk [2578]));
Q_ASSIGN U13813 ( .B(clk), .A(\g.we_clk [2577]));
Q_ASSIGN U13814 ( .B(clk), .A(\g.we_clk [2576]));
Q_ASSIGN U13815 ( .B(clk), .A(\g.we_clk [2575]));
Q_ASSIGN U13816 ( .B(clk), .A(\g.we_clk [2574]));
Q_ASSIGN U13817 ( .B(clk), .A(\g.we_clk [2573]));
Q_ASSIGN U13818 ( .B(clk), .A(\g.we_clk [2572]));
Q_ASSIGN U13819 ( .B(clk), .A(\g.we_clk [2571]));
Q_ASSIGN U13820 ( .B(clk), .A(\g.we_clk [2570]));
Q_ASSIGN U13821 ( .B(clk), .A(\g.we_clk [2569]));
Q_ASSIGN U13822 ( .B(clk), .A(\g.we_clk [2568]));
Q_ASSIGN U13823 ( .B(clk), .A(\g.we_clk [2567]));
Q_ASSIGN U13824 ( .B(clk), .A(\g.we_clk [2566]));
Q_ASSIGN U13825 ( .B(clk), .A(\g.we_clk [2565]));
Q_ASSIGN U13826 ( .B(clk), .A(\g.we_clk [2564]));
Q_ASSIGN U13827 ( .B(clk), .A(\g.we_clk [2563]));
Q_ASSIGN U13828 ( .B(clk), .A(\g.we_clk [2562]));
Q_ASSIGN U13829 ( .B(clk), .A(\g.we_clk [2561]));
Q_ASSIGN U13830 ( .B(clk), .A(\g.we_clk [2560]));
Q_ASSIGN U13831 ( .B(clk), .A(\g.we_clk [2559]));
Q_ASSIGN U13832 ( .B(clk), .A(\g.we_clk [2558]));
Q_ASSIGN U13833 ( .B(clk), .A(\g.we_clk [2557]));
Q_ASSIGN U13834 ( .B(clk), .A(\g.we_clk [2556]));
Q_ASSIGN U13835 ( .B(clk), .A(\g.we_clk [2555]));
Q_ASSIGN U13836 ( .B(clk), .A(\g.we_clk [2554]));
Q_ASSIGN U13837 ( .B(clk), .A(\g.we_clk [2553]));
Q_ASSIGN U13838 ( .B(clk), .A(\g.we_clk [2552]));
Q_ASSIGN U13839 ( .B(clk), .A(\g.we_clk [2551]));
Q_ASSIGN U13840 ( .B(clk), .A(\g.we_clk [2550]));
Q_ASSIGN U13841 ( .B(clk), .A(\g.we_clk [2549]));
Q_ASSIGN U13842 ( .B(clk), .A(\g.we_clk [2548]));
Q_ASSIGN U13843 ( .B(clk), .A(\g.we_clk [2547]));
Q_ASSIGN U13844 ( .B(clk), .A(\g.we_clk [2546]));
Q_ASSIGN U13845 ( .B(clk), .A(\g.we_clk [2545]));
Q_ASSIGN U13846 ( .B(clk), .A(\g.we_clk [2544]));
Q_ASSIGN U13847 ( .B(clk), .A(\g.we_clk [2543]));
Q_ASSIGN U13848 ( .B(clk), .A(\g.we_clk [2542]));
Q_ASSIGN U13849 ( .B(clk), .A(\g.we_clk [2541]));
Q_ASSIGN U13850 ( .B(clk), .A(\g.we_clk [2540]));
Q_ASSIGN U13851 ( .B(clk), .A(\g.we_clk [2539]));
Q_ASSIGN U13852 ( .B(clk), .A(\g.we_clk [2538]));
Q_ASSIGN U13853 ( .B(clk), .A(\g.we_clk [2537]));
Q_ASSIGN U13854 ( .B(clk), .A(\g.we_clk [2536]));
Q_ASSIGN U13855 ( .B(clk), .A(\g.we_clk [2535]));
Q_ASSIGN U13856 ( .B(clk), .A(\g.we_clk [2534]));
Q_ASSIGN U13857 ( .B(clk), .A(\g.we_clk [2533]));
Q_ASSIGN U13858 ( .B(clk), .A(\g.we_clk [2532]));
Q_ASSIGN U13859 ( .B(clk), .A(\g.we_clk [2531]));
Q_ASSIGN U13860 ( .B(clk), .A(\g.we_clk [2530]));
Q_ASSIGN U13861 ( .B(clk), .A(\g.we_clk [2529]));
Q_ASSIGN U13862 ( .B(clk), .A(\g.we_clk [2528]));
Q_ASSIGN U13863 ( .B(clk), .A(\g.we_clk [2527]));
Q_ASSIGN U13864 ( .B(clk), .A(\g.we_clk [2526]));
Q_ASSIGN U13865 ( .B(clk), .A(\g.we_clk [2525]));
Q_ASSIGN U13866 ( .B(clk), .A(\g.we_clk [2524]));
Q_ASSIGN U13867 ( .B(clk), .A(\g.we_clk [2523]));
Q_ASSIGN U13868 ( .B(clk), .A(\g.we_clk [2522]));
Q_ASSIGN U13869 ( .B(clk), .A(\g.we_clk [2521]));
Q_ASSIGN U13870 ( .B(clk), .A(\g.we_clk [2520]));
Q_ASSIGN U13871 ( .B(clk), .A(\g.we_clk [2519]));
Q_ASSIGN U13872 ( .B(clk), .A(\g.we_clk [2518]));
Q_ASSIGN U13873 ( .B(clk), .A(\g.we_clk [2517]));
Q_ASSIGN U13874 ( .B(clk), .A(\g.we_clk [2516]));
Q_ASSIGN U13875 ( .B(clk), .A(\g.we_clk [2515]));
Q_ASSIGN U13876 ( .B(clk), .A(\g.we_clk [2514]));
Q_ASSIGN U13877 ( .B(clk), .A(\g.we_clk [2513]));
Q_ASSIGN U13878 ( .B(clk), .A(\g.we_clk [2512]));
Q_ASSIGN U13879 ( .B(clk), .A(\g.we_clk [2511]));
Q_ASSIGN U13880 ( .B(clk), .A(\g.we_clk [2510]));
Q_ASSIGN U13881 ( .B(clk), .A(\g.we_clk [2509]));
Q_ASSIGN U13882 ( .B(clk), .A(\g.we_clk [2508]));
Q_ASSIGN U13883 ( .B(clk), .A(\g.we_clk [2507]));
Q_ASSIGN U13884 ( .B(clk), .A(\g.we_clk [2506]));
Q_ASSIGN U13885 ( .B(clk), .A(\g.we_clk [2505]));
Q_ASSIGN U13886 ( .B(clk), .A(\g.we_clk [2504]));
Q_ASSIGN U13887 ( .B(clk), .A(\g.we_clk [2503]));
Q_ASSIGN U13888 ( .B(clk), .A(\g.we_clk [2502]));
Q_ASSIGN U13889 ( .B(clk), .A(\g.we_clk [2501]));
Q_ASSIGN U13890 ( .B(clk), .A(\g.we_clk [2500]));
Q_ASSIGN U13891 ( .B(clk), .A(\g.we_clk [2499]));
Q_ASSIGN U13892 ( .B(clk), .A(\g.we_clk [2498]));
Q_ASSIGN U13893 ( .B(clk), .A(\g.we_clk [2497]));
Q_ASSIGN U13894 ( .B(clk), .A(\g.we_clk [2496]));
Q_ASSIGN U13895 ( .B(clk), .A(\g.we_clk [2495]));
Q_ASSIGN U13896 ( .B(clk), .A(\g.we_clk [2494]));
Q_ASSIGN U13897 ( .B(clk), .A(\g.we_clk [2493]));
Q_ASSIGN U13898 ( .B(clk), .A(\g.we_clk [2492]));
Q_ASSIGN U13899 ( .B(clk), .A(\g.we_clk [2491]));
Q_ASSIGN U13900 ( .B(clk), .A(\g.we_clk [2490]));
Q_ASSIGN U13901 ( .B(clk), .A(\g.we_clk [2489]));
Q_ASSIGN U13902 ( .B(clk), .A(\g.we_clk [2488]));
Q_ASSIGN U13903 ( .B(clk), .A(\g.we_clk [2487]));
Q_ASSIGN U13904 ( .B(clk), .A(\g.we_clk [2486]));
Q_ASSIGN U13905 ( .B(clk), .A(\g.we_clk [2485]));
Q_ASSIGN U13906 ( .B(clk), .A(\g.we_clk [2484]));
Q_ASSIGN U13907 ( .B(clk), .A(\g.we_clk [2483]));
Q_ASSIGN U13908 ( .B(clk), .A(\g.we_clk [2482]));
Q_ASSIGN U13909 ( .B(clk), .A(\g.we_clk [2481]));
Q_ASSIGN U13910 ( .B(clk), .A(\g.we_clk [2480]));
Q_ASSIGN U13911 ( .B(clk), .A(\g.we_clk [2479]));
Q_ASSIGN U13912 ( .B(clk), .A(\g.we_clk [2478]));
Q_ASSIGN U13913 ( .B(clk), .A(\g.we_clk [2477]));
Q_ASSIGN U13914 ( .B(clk), .A(\g.we_clk [2476]));
Q_ASSIGN U13915 ( .B(clk), .A(\g.we_clk [2475]));
Q_ASSIGN U13916 ( .B(clk), .A(\g.we_clk [2474]));
Q_ASSIGN U13917 ( .B(clk), .A(\g.we_clk [2473]));
Q_ASSIGN U13918 ( .B(clk), .A(\g.we_clk [2472]));
Q_ASSIGN U13919 ( .B(clk), .A(\g.we_clk [2471]));
Q_ASSIGN U13920 ( .B(clk), .A(\g.we_clk [2470]));
Q_ASSIGN U13921 ( .B(clk), .A(\g.we_clk [2469]));
Q_ASSIGN U13922 ( .B(clk), .A(\g.we_clk [2468]));
Q_ASSIGN U13923 ( .B(clk), .A(\g.we_clk [2467]));
Q_ASSIGN U13924 ( .B(clk), .A(\g.we_clk [2466]));
Q_ASSIGN U13925 ( .B(clk), .A(\g.we_clk [2465]));
Q_ASSIGN U13926 ( .B(clk), .A(\g.we_clk [2464]));
Q_ASSIGN U13927 ( .B(clk), .A(\g.we_clk [2463]));
Q_ASSIGN U13928 ( .B(clk), .A(\g.we_clk [2462]));
Q_ASSIGN U13929 ( .B(clk), .A(\g.we_clk [2461]));
Q_ASSIGN U13930 ( .B(clk), .A(\g.we_clk [2460]));
Q_ASSIGN U13931 ( .B(clk), .A(\g.we_clk [2459]));
Q_ASSIGN U13932 ( .B(clk), .A(\g.we_clk [2458]));
Q_ASSIGN U13933 ( .B(clk), .A(\g.we_clk [2457]));
Q_ASSIGN U13934 ( .B(clk), .A(\g.we_clk [2456]));
Q_ASSIGN U13935 ( .B(clk), .A(\g.we_clk [2455]));
Q_ASSIGN U13936 ( .B(clk), .A(\g.we_clk [2454]));
Q_ASSIGN U13937 ( .B(clk), .A(\g.we_clk [2453]));
Q_ASSIGN U13938 ( .B(clk), .A(\g.we_clk [2452]));
Q_ASSIGN U13939 ( .B(clk), .A(\g.we_clk [2451]));
Q_ASSIGN U13940 ( .B(clk), .A(\g.we_clk [2450]));
Q_ASSIGN U13941 ( .B(clk), .A(\g.we_clk [2449]));
Q_ASSIGN U13942 ( .B(clk), .A(\g.we_clk [2448]));
Q_ASSIGN U13943 ( .B(clk), .A(\g.we_clk [2447]));
Q_ASSIGN U13944 ( .B(clk), .A(\g.we_clk [2446]));
Q_ASSIGN U13945 ( .B(clk), .A(\g.we_clk [2445]));
Q_ASSIGN U13946 ( .B(clk), .A(\g.we_clk [2444]));
Q_ASSIGN U13947 ( .B(clk), .A(\g.we_clk [2443]));
Q_ASSIGN U13948 ( .B(clk), .A(\g.we_clk [2442]));
Q_ASSIGN U13949 ( .B(clk), .A(\g.we_clk [2441]));
Q_ASSIGN U13950 ( .B(clk), .A(\g.we_clk [2440]));
Q_ASSIGN U13951 ( .B(clk), .A(\g.we_clk [2439]));
Q_ASSIGN U13952 ( .B(clk), .A(\g.we_clk [2438]));
Q_ASSIGN U13953 ( .B(clk), .A(\g.we_clk [2437]));
Q_ASSIGN U13954 ( .B(clk), .A(\g.we_clk [2436]));
Q_ASSIGN U13955 ( .B(clk), .A(\g.we_clk [2435]));
Q_ASSIGN U13956 ( .B(clk), .A(\g.we_clk [2434]));
Q_ASSIGN U13957 ( .B(clk), .A(\g.we_clk [2433]));
Q_ASSIGN U13958 ( .B(clk), .A(\g.we_clk [2432]));
Q_ASSIGN U13959 ( .B(clk), .A(\g.we_clk [2431]));
Q_ASSIGN U13960 ( .B(clk), .A(\g.we_clk [2430]));
Q_ASSIGN U13961 ( .B(clk), .A(\g.we_clk [2429]));
Q_ASSIGN U13962 ( .B(clk), .A(\g.we_clk [2428]));
Q_ASSIGN U13963 ( .B(clk), .A(\g.we_clk [2427]));
Q_ASSIGN U13964 ( .B(clk), .A(\g.we_clk [2426]));
Q_ASSIGN U13965 ( .B(clk), .A(\g.we_clk [2425]));
Q_ASSIGN U13966 ( .B(clk), .A(\g.we_clk [2424]));
Q_ASSIGN U13967 ( .B(clk), .A(\g.we_clk [2423]));
Q_ASSIGN U13968 ( .B(clk), .A(\g.we_clk [2422]));
Q_ASSIGN U13969 ( .B(clk), .A(\g.we_clk [2421]));
Q_ASSIGN U13970 ( .B(clk), .A(\g.we_clk [2420]));
Q_ASSIGN U13971 ( .B(clk), .A(\g.we_clk [2419]));
Q_ASSIGN U13972 ( .B(clk), .A(\g.we_clk [2418]));
Q_ASSIGN U13973 ( .B(clk), .A(\g.we_clk [2417]));
Q_ASSIGN U13974 ( .B(clk), .A(\g.we_clk [2416]));
Q_ASSIGN U13975 ( .B(clk), .A(\g.we_clk [2415]));
Q_ASSIGN U13976 ( .B(clk), .A(\g.we_clk [2414]));
Q_ASSIGN U13977 ( .B(clk), .A(\g.we_clk [2413]));
Q_ASSIGN U13978 ( .B(clk), .A(\g.we_clk [2412]));
Q_ASSIGN U13979 ( .B(clk), .A(\g.we_clk [2411]));
Q_ASSIGN U13980 ( .B(clk), .A(\g.we_clk [2410]));
Q_ASSIGN U13981 ( .B(clk), .A(\g.we_clk [2409]));
Q_ASSIGN U13982 ( .B(clk), .A(\g.we_clk [2408]));
Q_ASSIGN U13983 ( .B(clk), .A(\g.we_clk [2407]));
Q_ASSIGN U13984 ( .B(clk), .A(\g.we_clk [2406]));
Q_ASSIGN U13985 ( .B(clk), .A(\g.we_clk [2405]));
Q_ASSIGN U13986 ( .B(clk), .A(\g.we_clk [2404]));
Q_ASSIGN U13987 ( .B(clk), .A(\g.we_clk [2403]));
Q_ASSIGN U13988 ( .B(clk), .A(\g.we_clk [2402]));
Q_ASSIGN U13989 ( .B(clk), .A(\g.we_clk [2401]));
Q_ASSIGN U13990 ( .B(clk), .A(\g.we_clk [2400]));
Q_ASSIGN U13991 ( .B(clk), .A(\g.we_clk [2399]));
Q_ASSIGN U13992 ( .B(clk), .A(\g.we_clk [2398]));
Q_ASSIGN U13993 ( .B(clk), .A(\g.we_clk [2397]));
Q_ASSIGN U13994 ( .B(clk), .A(\g.we_clk [2396]));
Q_ASSIGN U13995 ( .B(clk), .A(\g.we_clk [2395]));
Q_ASSIGN U13996 ( .B(clk), .A(\g.we_clk [2394]));
Q_ASSIGN U13997 ( .B(clk), .A(\g.we_clk [2393]));
Q_ASSIGN U13998 ( .B(clk), .A(\g.we_clk [2392]));
Q_ASSIGN U13999 ( .B(clk), .A(\g.we_clk [2391]));
Q_ASSIGN U14000 ( .B(clk), .A(\g.we_clk [2390]));
Q_ASSIGN U14001 ( .B(clk), .A(\g.we_clk [2389]));
Q_ASSIGN U14002 ( .B(clk), .A(\g.we_clk [2388]));
Q_ASSIGN U14003 ( .B(clk), .A(\g.we_clk [2387]));
Q_ASSIGN U14004 ( .B(clk), .A(\g.we_clk [2386]));
Q_ASSIGN U14005 ( .B(clk), .A(\g.we_clk [2385]));
Q_ASSIGN U14006 ( .B(clk), .A(\g.we_clk [2384]));
Q_ASSIGN U14007 ( .B(clk), .A(\g.we_clk [2383]));
Q_ASSIGN U14008 ( .B(clk), .A(\g.we_clk [2382]));
Q_ASSIGN U14009 ( .B(clk), .A(\g.we_clk [2381]));
Q_ASSIGN U14010 ( .B(clk), .A(\g.we_clk [2380]));
Q_ASSIGN U14011 ( .B(clk), .A(\g.we_clk [2379]));
Q_ASSIGN U14012 ( .B(clk), .A(\g.we_clk [2378]));
Q_ASSIGN U14013 ( .B(clk), .A(\g.we_clk [2377]));
Q_ASSIGN U14014 ( .B(clk), .A(\g.we_clk [2376]));
Q_ASSIGN U14015 ( .B(clk), .A(\g.we_clk [2375]));
Q_ASSIGN U14016 ( .B(clk), .A(\g.we_clk [2374]));
Q_ASSIGN U14017 ( .B(clk), .A(\g.we_clk [2373]));
Q_ASSIGN U14018 ( .B(clk), .A(\g.we_clk [2372]));
Q_ASSIGN U14019 ( .B(clk), .A(\g.we_clk [2371]));
Q_ASSIGN U14020 ( .B(clk), .A(\g.we_clk [2370]));
Q_ASSIGN U14021 ( .B(clk), .A(\g.we_clk [2369]));
Q_ASSIGN U14022 ( .B(clk), .A(\g.we_clk [2368]));
Q_ASSIGN U14023 ( .B(clk), .A(\g.we_clk [2367]));
Q_ASSIGN U14024 ( .B(clk), .A(\g.we_clk [2366]));
Q_ASSIGN U14025 ( .B(clk), .A(\g.we_clk [2365]));
Q_ASSIGN U14026 ( .B(clk), .A(\g.we_clk [2364]));
Q_ASSIGN U14027 ( .B(clk), .A(\g.we_clk [2363]));
Q_ASSIGN U14028 ( .B(clk), .A(\g.we_clk [2362]));
Q_ASSIGN U14029 ( .B(clk), .A(\g.we_clk [2361]));
Q_ASSIGN U14030 ( .B(clk), .A(\g.we_clk [2360]));
Q_ASSIGN U14031 ( .B(clk), .A(\g.we_clk [2359]));
Q_ASSIGN U14032 ( .B(clk), .A(\g.we_clk [2358]));
Q_ASSIGN U14033 ( .B(clk), .A(\g.we_clk [2357]));
Q_ASSIGN U14034 ( .B(clk), .A(\g.we_clk [2356]));
Q_ASSIGN U14035 ( .B(clk), .A(\g.we_clk [2355]));
Q_ASSIGN U14036 ( .B(clk), .A(\g.we_clk [2354]));
Q_ASSIGN U14037 ( .B(clk), .A(\g.we_clk [2353]));
Q_ASSIGN U14038 ( .B(clk), .A(\g.we_clk [2352]));
Q_ASSIGN U14039 ( .B(clk), .A(\g.we_clk [2351]));
Q_ASSIGN U14040 ( .B(clk), .A(\g.we_clk [2350]));
Q_ASSIGN U14041 ( .B(clk), .A(\g.we_clk [2349]));
Q_ASSIGN U14042 ( .B(clk), .A(\g.we_clk [2348]));
Q_ASSIGN U14043 ( .B(clk), .A(\g.we_clk [2347]));
Q_ASSIGN U14044 ( .B(clk), .A(\g.we_clk [2346]));
Q_ASSIGN U14045 ( .B(clk), .A(\g.we_clk [2345]));
Q_ASSIGN U14046 ( .B(clk), .A(\g.we_clk [2344]));
Q_ASSIGN U14047 ( .B(clk), .A(\g.we_clk [2343]));
Q_ASSIGN U14048 ( .B(clk), .A(\g.we_clk [2342]));
Q_ASSIGN U14049 ( .B(clk), .A(\g.we_clk [2341]));
Q_ASSIGN U14050 ( .B(clk), .A(\g.we_clk [2340]));
Q_ASSIGN U14051 ( .B(clk), .A(\g.we_clk [2339]));
Q_ASSIGN U14052 ( .B(clk), .A(\g.we_clk [2338]));
Q_ASSIGN U14053 ( .B(clk), .A(\g.we_clk [2337]));
Q_ASSIGN U14054 ( .B(clk), .A(\g.we_clk [2336]));
Q_ASSIGN U14055 ( .B(clk), .A(\g.we_clk [2335]));
Q_ASSIGN U14056 ( .B(clk), .A(\g.we_clk [2334]));
Q_ASSIGN U14057 ( .B(clk), .A(\g.we_clk [2333]));
Q_ASSIGN U14058 ( .B(clk), .A(\g.we_clk [2332]));
Q_ASSIGN U14059 ( .B(clk), .A(\g.we_clk [2331]));
Q_ASSIGN U14060 ( .B(clk), .A(\g.we_clk [2330]));
Q_ASSIGN U14061 ( .B(clk), .A(\g.we_clk [2329]));
Q_ASSIGN U14062 ( .B(clk), .A(\g.we_clk [2328]));
Q_ASSIGN U14063 ( .B(clk), .A(\g.we_clk [2327]));
Q_ASSIGN U14064 ( .B(clk), .A(\g.we_clk [2326]));
Q_ASSIGN U14065 ( .B(clk), .A(\g.we_clk [2325]));
Q_ASSIGN U14066 ( .B(clk), .A(\g.we_clk [2324]));
Q_ASSIGN U14067 ( .B(clk), .A(\g.we_clk [2323]));
Q_ASSIGN U14068 ( .B(clk), .A(\g.we_clk [2322]));
Q_ASSIGN U14069 ( .B(clk), .A(\g.we_clk [2321]));
Q_ASSIGN U14070 ( .B(clk), .A(\g.we_clk [2320]));
Q_ASSIGN U14071 ( .B(clk), .A(\g.we_clk [2319]));
Q_ASSIGN U14072 ( .B(clk), .A(\g.we_clk [2318]));
Q_ASSIGN U14073 ( .B(clk), .A(\g.we_clk [2317]));
Q_ASSIGN U14074 ( .B(clk), .A(\g.we_clk [2316]));
Q_ASSIGN U14075 ( .B(clk), .A(\g.we_clk [2315]));
Q_ASSIGN U14076 ( .B(clk), .A(\g.we_clk [2314]));
Q_ASSIGN U14077 ( .B(clk), .A(\g.we_clk [2313]));
Q_ASSIGN U14078 ( .B(clk), .A(\g.we_clk [2312]));
Q_ASSIGN U14079 ( .B(clk), .A(\g.we_clk [2311]));
Q_ASSIGN U14080 ( .B(clk), .A(\g.we_clk [2310]));
Q_ASSIGN U14081 ( .B(clk), .A(\g.we_clk [2309]));
Q_ASSIGN U14082 ( .B(clk), .A(\g.we_clk [2308]));
Q_ASSIGN U14083 ( .B(clk), .A(\g.we_clk [2307]));
Q_ASSIGN U14084 ( .B(clk), .A(\g.we_clk [2306]));
Q_ASSIGN U14085 ( .B(clk), .A(\g.we_clk [2305]));
Q_ASSIGN U14086 ( .B(clk), .A(\g.we_clk [2304]));
Q_ASSIGN U14087 ( .B(clk), .A(\g.we_clk [2303]));
Q_ASSIGN U14088 ( .B(clk), .A(\g.we_clk [2302]));
Q_ASSIGN U14089 ( .B(clk), .A(\g.we_clk [2301]));
Q_ASSIGN U14090 ( .B(clk), .A(\g.we_clk [2300]));
Q_ASSIGN U14091 ( .B(clk), .A(\g.we_clk [2299]));
Q_ASSIGN U14092 ( .B(clk), .A(\g.we_clk [2298]));
Q_ASSIGN U14093 ( .B(clk), .A(\g.we_clk [2297]));
Q_ASSIGN U14094 ( .B(clk), .A(\g.we_clk [2296]));
Q_ASSIGN U14095 ( .B(clk), .A(\g.we_clk [2295]));
Q_ASSIGN U14096 ( .B(clk), .A(\g.we_clk [2294]));
Q_ASSIGN U14097 ( .B(clk), .A(\g.we_clk [2293]));
Q_ASSIGN U14098 ( .B(clk), .A(\g.we_clk [2292]));
Q_ASSIGN U14099 ( .B(clk), .A(\g.we_clk [2291]));
Q_ASSIGN U14100 ( .B(clk), .A(\g.we_clk [2290]));
Q_ASSIGN U14101 ( .B(clk), .A(\g.we_clk [2289]));
Q_ASSIGN U14102 ( .B(clk), .A(\g.we_clk [2288]));
Q_ASSIGN U14103 ( .B(clk), .A(\g.we_clk [2287]));
Q_ASSIGN U14104 ( .B(clk), .A(\g.we_clk [2286]));
Q_ASSIGN U14105 ( .B(clk), .A(\g.we_clk [2285]));
Q_ASSIGN U14106 ( .B(clk), .A(\g.we_clk [2284]));
Q_ASSIGN U14107 ( .B(clk), .A(\g.we_clk [2283]));
Q_ASSIGN U14108 ( .B(clk), .A(\g.we_clk [2282]));
Q_ASSIGN U14109 ( .B(clk), .A(\g.we_clk [2281]));
Q_ASSIGN U14110 ( .B(clk), .A(\g.we_clk [2280]));
Q_ASSIGN U14111 ( .B(clk), .A(\g.we_clk [2279]));
Q_ASSIGN U14112 ( .B(clk), .A(\g.we_clk [2278]));
Q_ASSIGN U14113 ( .B(clk), .A(\g.we_clk [2277]));
Q_ASSIGN U14114 ( .B(clk), .A(\g.we_clk [2276]));
Q_ASSIGN U14115 ( .B(clk), .A(\g.we_clk [2275]));
Q_ASSIGN U14116 ( .B(clk), .A(\g.we_clk [2274]));
Q_ASSIGN U14117 ( .B(clk), .A(\g.we_clk [2273]));
Q_ASSIGN U14118 ( .B(clk), .A(\g.we_clk [2272]));
Q_ASSIGN U14119 ( .B(clk), .A(\g.we_clk [2271]));
Q_ASSIGN U14120 ( .B(clk), .A(\g.we_clk [2270]));
Q_ASSIGN U14121 ( .B(clk), .A(\g.we_clk [2269]));
Q_ASSIGN U14122 ( .B(clk), .A(\g.we_clk [2268]));
Q_ASSIGN U14123 ( .B(clk), .A(\g.we_clk [2267]));
Q_ASSIGN U14124 ( .B(clk), .A(\g.we_clk [2266]));
Q_ASSIGN U14125 ( .B(clk), .A(\g.we_clk [2265]));
Q_ASSIGN U14126 ( .B(clk), .A(\g.we_clk [2264]));
Q_ASSIGN U14127 ( .B(clk), .A(\g.we_clk [2263]));
Q_ASSIGN U14128 ( .B(clk), .A(\g.we_clk [2262]));
Q_ASSIGN U14129 ( .B(clk), .A(\g.we_clk [2261]));
Q_ASSIGN U14130 ( .B(clk), .A(\g.we_clk [2260]));
Q_ASSIGN U14131 ( .B(clk), .A(\g.we_clk [2259]));
Q_ASSIGN U14132 ( .B(clk), .A(\g.we_clk [2258]));
Q_ASSIGN U14133 ( .B(clk), .A(\g.we_clk [2257]));
Q_ASSIGN U14134 ( .B(clk), .A(\g.we_clk [2256]));
Q_ASSIGN U14135 ( .B(clk), .A(\g.we_clk [2255]));
Q_ASSIGN U14136 ( .B(clk), .A(\g.we_clk [2254]));
Q_ASSIGN U14137 ( .B(clk), .A(\g.we_clk [2253]));
Q_ASSIGN U14138 ( .B(clk), .A(\g.we_clk [2252]));
Q_ASSIGN U14139 ( .B(clk), .A(\g.we_clk [2251]));
Q_ASSIGN U14140 ( .B(clk), .A(\g.we_clk [2250]));
Q_ASSIGN U14141 ( .B(clk), .A(\g.we_clk [2249]));
Q_ASSIGN U14142 ( .B(clk), .A(\g.we_clk [2248]));
Q_ASSIGN U14143 ( .B(clk), .A(\g.we_clk [2247]));
Q_ASSIGN U14144 ( .B(clk), .A(\g.we_clk [2246]));
Q_ASSIGN U14145 ( .B(clk), .A(\g.we_clk [2245]));
Q_ASSIGN U14146 ( .B(clk), .A(\g.we_clk [2244]));
Q_ASSIGN U14147 ( .B(clk), .A(\g.we_clk [2243]));
Q_ASSIGN U14148 ( .B(clk), .A(\g.we_clk [2242]));
Q_ASSIGN U14149 ( .B(clk), .A(\g.we_clk [2241]));
Q_ASSIGN U14150 ( .B(clk), .A(\g.we_clk [2240]));
Q_ASSIGN U14151 ( .B(clk), .A(\g.we_clk [2239]));
Q_ASSIGN U14152 ( .B(clk), .A(\g.we_clk [2238]));
Q_ASSIGN U14153 ( .B(clk), .A(\g.we_clk [2237]));
Q_ASSIGN U14154 ( .B(clk), .A(\g.we_clk [2236]));
Q_ASSIGN U14155 ( .B(clk), .A(\g.we_clk [2235]));
Q_ASSIGN U14156 ( .B(clk), .A(\g.we_clk [2234]));
Q_ASSIGN U14157 ( .B(clk), .A(\g.we_clk [2233]));
Q_ASSIGN U14158 ( .B(clk), .A(\g.we_clk [2232]));
Q_ASSIGN U14159 ( .B(clk), .A(\g.we_clk [2231]));
Q_ASSIGN U14160 ( .B(clk), .A(\g.we_clk [2230]));
Q_ASSIGN U14161 ( .B(clk), .A(\g.we_clk [2229]));
Q_ASSIGN U14162 ( .B(clk), .A(\g.we_clk [2228]));
Q_ASSIGN U14163 ( .B(clk), .A(\g.we_clk [2227]));
Q_ASSIGN U14164 ( .B(clk), .A(\g.we_clk [2226]));
Q_ASSIGN U14165 ( .B(clk), .A(\g.we_clk [2225]));
Q_ASSIGN U14166 ( .B(clk), .A(\g.we_clk [2224]));
Q_ASSIGN U14167 ( .B(clk), .A(\g.we_clk [2223]));
Q_ASSIGN U14168 ( .B(clk), .A(\g.we_clk [2222]));
Q_ASSIGN U14169 ( .B(clk), .A(\g.we_clk [2221]));
Q_ASSIGN U14170 ( .B(clk), .A(\g.we_clk [2220]));
Q_ASSIGN U14171 ( .B(clk), .A(\g.we_clk [2219]));
Q_ASSIGN U14172 ( .B(clk), .A(\g.we_clk [2218]));
Q_ASSIGN U14173 ( .B(clk), .A(\g.we_clk [2217]));
Q_ASSIGN U14174 ( .B(clk), .A(\g.we_clk [2216]));
Q_ASSIGN U14175 ( .B(clk), .A(\g.we_clk [2215]));
Q_ASSIGN U14176 ( .B(clk), .A(\g.we_clk [2214]));
Q_ASSIGN U14177 ( .B(clk), .A(\g.we_clk [2213]));
Q_ASSIGN U14178 ( .B(clk), .A(\g.we_clk [2212]));
Q_ASSIGN U14179 ( .B(clk), .A(\g.we_clk [2211]));
Q_ASSIGN U14180 ( .B(clk), .A(\g.we_clk [2210]));
Q_ASSIGN U14181 ( .B(clk), .A(\g.we_clk [2209]));
Q_ASSIGN U14182 ( .B(clk), .A(\g.we_clk [2208]));
Q_ASSIGN U14183 ( .B(clk), .A(\g.we_clk [2207]));
Q_ASSIGN U14184 ( .B(clk), .A(\g.we_clk [2206]));
Q_ASSIGN U14185 ( .B(clk), .A(\g.we_clk [2205]));
Q_ASSIGN U14186 ( .B(clk), .A(\g.we_clk [2204]));
Q_ASSIGN U14187 ( .B(clk), .A(\g.we_clk [2203]));
Q_ASSIGN U14188 ( .B(clk), .A(\g.we_clk [2202]));
Q_ASSIGN U14189 ( .B(clk), .A(\g.we_clk [2201]));
Q_ASSIGN U14190 ( .B(clk), .A(\g.we_clk [2200]));
Q_ASSIGN U14191 ( .B(clk), .A(\g.we_clk [2199]));
Q_ASSIGN U14192 ( .B(clk), .A(\g.we_clk [2198]));
Q_ASSIGN U14193 ( .B(clk), .A(\g.we_clk [2197]));
Q_ASSIGN U14194 ( .B(clk), .A(\g.we_clk [2196]));
Q_ASSIGN U14195 ( .B(clk), .A(\g.we_clk [2195]));
Q_ASSIGN U14196 ( .B(clk), .A(\g.we_clk [2194]));
Q_ASSIGN U14197 ( .B(clk), .A(\g.we_clk [2193]));
Q_ASSIGN U14198 ( .B(clk), .A(\g.we_clk [2192]));
Q_ASSIGN U14199 ( .B(clk), .A(\g.we_clk [2191]));
Q_ASSIGN U14200 ( .B(clk), .A(\g.we_clk [2190]));
Q_ASSIGN U14201 ( .B(clk), .A(\g.we_clk [2189]));
Q_ASSIGN U14202 ( .B(clk), .A(\g.we_clk [2188]));
Q_ASSIGN U14203 ( .B(clk), .A(\g.we_clk [2187]));
Q_ASSIGN U14204 ( .B(clk), .A(\g.we_clk [2186]));
Q_ASSIGN U14205 ( .B(clk), .A(\g.we_clk [2185]));
Q_ASSIGN U14206 ( .B(clk), .A(\g.we_clk [2184]));
Q_ASSIGN U14207 ( .B(clk), .A(\g.we_clk [2183]));
Q_ASSIGN U14208 ( .B(clk), .A(\g.we_clk [2182]));
Q_ASSIGN U14209 ( .B(clk), .A(\g.we_clk [2181]));
Q_ASSIGN U14210 ( .B(clk), .A(\g.we_clk [2180]));
Q_ASSIGN U14211 ( .B(clk), .A(\g.we_clk [2179]));
Q_ASSIGN U14212 ( .B(clk), .A(\g.we_clk [2178]));
Q_ASSIGN U14213 ( .B(clk), .A(\g.we_clk [2177]));
Q_ASSIGN U14214 ( .B(clk), .A(\g.we_clk [2176]));
Q_ASSIGN U14215 ( .B(clk), .A(\g.we_clk [2175]));
Q_ASSIGN U14216 ( .B(clk), .A(\g.we_clk [2174]));
Q_ASSIGN U14217 ( .B(clk), .A(\g.we_clk [2173]));
Q_ASSIGN U14218 ( .B(clk), .A(\g.we_clk [2172]));
Q_ASSIGN U14219 ( .B(clk), .A(\g.we_clk [2171]));
Q_ASSIGN U14220 ( .B(clk), .A(\g.we_clk [2170]));
Q_ASSIGN U14221 ( .B(clk), .A(\g.we_clk [2169]));
Q_ASSIGN U14222 ( .B(clk), .A(\g.we_clk [2168]));
Q_ASSIGN U14223 ( .B(clk), .A(\g.we_clk [2167]));
Q_ASSIGN U14224 ( .B(clk), .A(\g.we_clk [2166]));
Q_ASSIGN U14225 ( .B(clk), .A(\g.we_clk [2165]));
Q_ASSIGN U14226 ( .B(clk), .A(\g.we_clk [2164]));
Q_ASSIGN U14227 ( .B(clk), .A(\g.we_clk [2163]));
Q_ASSIGN U14228 ( .B(clk), .A(\g.we_clk [2162]));
Q_ASSIGN U14229 ( .B(clk), .A(\g.we_clk [2161]));
Q_ASSIGN U14230 ( .B(clk), .A(\g.we_clk [2160]));
Q_ASSIGN U14231 ( .B(clk), .A(\g.we_clk [2159]));
Q_ASSIGN U14232 ( .B(clk), .A(\g.we_clk [2158]));
Q_ASSIGN U14233 ( .B(clk), .A(\g.we_clk [2157]));
Q_ASSIGN U14234 ( .B(clk), .A(\g.we_clk [2156]));
Q_ASSIGN U14235 ( .B(clk), .A(\g.we_clk [2155]));
Q_ASSIGN U14236 ( .B(clk), .A(\g.we_clk [2154]));
Q_ASSIGN U14237 ( .B(clk), .A(\g.we_clk [2153]));
Q_ASSIGN U14238 ( .B(clk), .A(\g.we_clk [2152]));
Q_ASSIGN U14239 ( .B(clk), .A(\g.we_clk [2151]));
Q_ASSIGN U14240 ( .B(clk), .A(\g.we_clk [2150]));
Q_ASSIGN U14241 ( .B(clk), .A(\g.we_clk [2149]));
Q_ASSIGN U14242 ( .B(clk), .A(\g.we_clk [2148]));
Q_ASSIGN U14243 ( .B(clk), .A(\g.we_clk [2147]));
Q_ASSIGN U14244 ( .B(clk), .A(\g.we_clk [2146]));
Q_ASSIGN U14245 ( .B(clk), .A(\g.we_clk [2145]));
Q_ASSIGN U14246 ( .B(clk), .A(\g.we_clk [2144]));
Q_ASSIGN U14247 ( .B(clk), .A(\g.we_clk [2143]));
Q_ASSIGN U14248 ( .B(clk), .A(\g.we_clk [2142]));
Q_ASSIGN U14249 ( .B(clk), .A(\g.we_clk [2141]));
Q_ASSIGN U14250 ( .B(clk), .A(\g.we_clk [2140]));
Q_ASSIGN U14251 ( .B(clk), .A(\g.we_clk [2139]));
Q_ASSIGN U14252 ( .B(clk), .A(\g.we_clk [2138]));
Q_ASSIGN U14253 ( .B(clk), .A(\g.we_clk [2137]));
Q_ASSIGN U14254 ( .B(clk), .A(\g.we_clk [2136]));
Q_ASSIGN U14255 ( .B(clk), .A(\g.we_clk [2135]));
Q_ASSIGN U14256 ( .B(clk), .A(\g.we_clk [2134]));
Q_ASSIGN U14257 ( .B(clk), .A(\g.we_clk [2133]));
Q_ASSIGN U14258 ( .B(clk), .A(\g.we_clk [2132]));
Q_ASSIGN U14259 ( .B(clk), .A(\g.we_clk [2131]));
Q_ASSIGN U14260 ( .B(clk), .A(\g.we_clk [2130]));
Q_ASSIGN U14261 ( .B(clk), .A(\g.we_clk [2129]));
Q_ASSIGN U14262 ( .B(clk), .A(\g.we_clk [2128]));
Q_ASSIGN U14263 ( .B(clk), .A(\g.we_clk [2127]));
Q_ASSIGN U14264 ( .B(clk), .A(\g.we_clk [2126]));
Q_ASSIGN U14265 ( .B(clk), .A(\g.we_clk [2125]));
Q_ASSIGN U14266 ( .B(clk), .A(\g.we_clk [2124]));
Q_ASSIGN U14267 ( .B(clk), .A(\g.we_clk [2123]));
Q_ASSIGN U14268 ( .B(clk), .A(\g.we_clk [2122]));
Q_ASSIGN U14269 ( .B(clk), .A(\g.we_clk [2121]));
Q_ASSIGN U14270 ( .B(clk), .A(\g.we_clk [2120]));
Q_ASSIGN U14271 ( .B(clk), .A(\g.we_clk [2119]));
Q_ASSIGN U14272 ( .B(clk), .A(\g.we_clk [2118]));
Q_ASSIGN U14273 ( .B(clk), .A(\g.we_clk [2117]));
Q_ASSIGN U14274 ( .B(clk), .A(\g.we_clk [2116]));
Q_ASSIGN U14275 ( .B(clk), .A(\g.we_clk [2115]));
Q_ASSIGN U14276 ( .B(clk), .A(\g.we_clk [2114]));
Q_ASSIGN U14277 ( .B(clk), .A(\g.we_clk [2113]));
Q_ASSIGN U14278 ( .B(clk), .A(\g.we_clk [2112]));
Q_ASSIGN U14279 ( .B(clk), .A(\g.we_clk [2111]));
Q_ASSIGN U14280 ( .B(clk), .A(\g.we_clk [2110]));
Q_ASSIGN U14281 ( .B(clk), .A(\g.we_clk [2109]));
Q_ASSIGN U14282 ( .B(clk), .A(\g.we_clk [2108]));
Q_ASSIGN U14283 ( .B(clk), .A(\g.we_clk [2107]));
Q_ASSIGN U14284 ( .B(clk), .A(\g.we_clk [2106]));
Q_ASSIGN U14285 ( .B(clk), .A(\g.we_clk [2105]));
Q_ASSIGN U14286 ( .B(clk), .A(\g.we_clk [2104]));
Q_ASSIGN U14287 ( .B(clk), .A(\g.we_clk [2103]));
Q_ASSIGN U14288 ( .B(clk), .A(\g.we_clk [2102]));
Q_ASSIGN U14289 ( .B(clk), .A(\g.we_clk [2101]));
Q_ASSIGN U14290 ( .B(clk), .A(\g.we_clk [2100]));
Q_ASSIGN U14291 ( .B(clk), .A(\g.we_clk [2099]));
Q_ASSIGN U14292 ( .B(clk), .A(\g.we_clk [2098]));
Q_ASSIGN U14293 ( .B(clk), .A(\g.we_clk [2097]));
Q_ASSIGN U14294 ( .B(clk), .A(\g.we_clk [2096]));
Q_ASSIGN U14295 ( .B(clk), .A(\g.we_clk [2095]));
Q_ASSIGN U14296 ( .B(clk), .A(\g.we_clk [2094]));
Q_ASSIGN U14297 ( .B(clk), .A(\g.we_clk [2093]));
Q_ASSIGN U14298 ( .B(clk), .A(\g.we_clk [2092]));
Q_ASSIGN U14299 ( .B(clk), .A(\g.we_clk [2091]));
Q_ASSIGN U14300 ( .B(clk), .A(\g.we_clk [2090]));
Q_ASSIGN U14301 ( .B(clk), .A(\g.we_clk [2089]));
Q_ASSIGN U14302 ( .B(clk), .A(\g.we_clk [2088]));
Q_ASSIGN U14303 ( .B(clk), .A(\g.we_clk [2087]));
Q_ASSIGN U14304 ( .B(clk), .A(\g.we_clk [2086]));
Q_ASSIGN U14305 ( .B(clk), .A(\g.we_clk [2085]));
Q_ASSIGN U14306 ( .B(clk), .A(\g.we_clk [2084]));
Q_ASSIGN U14307 ( .B(clk), .A(\g.we_clk [2083]));
Q_ASSIGN U14308 ( .B(clk), .A(\g.we_clk [2082]));
Q_ASSIGN U14309 ( .B(clk), .A(\g.we_clk [2081]));
Q_ASSIGN U14310 ( .B(clk), .A(\g.we_clk [2080]));
Q_ASSIGN U14311 ( .B(clk), .A(\g.we_clk [2079]));
Q_ASSIGN U14312 ( .B(clk), .A(\g.we_clk [2078]));
Q_ASSIGN U14313 ( .B(clk), .A(\g.we_clk [2077]));
Q_ASSIGN U14314 ( .B(clk), .A(\g.we_clk [2076]));
Q_ASSIGN U14315 ( .B(clk), .A(\g.we_clk [2075]));
Q_ASSIGN U14316 ( .B(clk), .A(\g.we_clk [2074]));
Q_ASSIGN U14317 ( .B(clk), .A(\g.we_clk [2073]));
Q_ASSIGN U14318 ( .B(clk), .A(\g.we_clk [2072]));
Q_ASSIGN U14319 ( .B(clk), .A(\g.we_clk [2071]));
Q_ASSIGN U14320 ( .B(clk), .A(\g.we_clk [2070]));
Q_ASSIGN U14321 ( .B(clk), .A(\g.we_clk [2069]));
Q_ASSIGN U14322 ( .B(clk), .A(\g.we_clk [2068]));
Q_ASSIGN U14323 ( .B(clk), .A(\g.we_clk [2067]));
Q_ASSIGN U14324 ( .B(clk), .A(\g.we_clk [2066]));
Q_ASSIGN U14325 ( .B(clk), .A(\g.we_clk [2065]));
Q_ASSIGN U14326 ( .B(clk), .A(\g.we_clk [2064]));
Q_ASSIGN U14327 ( .B(clk), .A(\g.we_clk [2063]));
Q_ASSIGN U14328 ( .B(clk), .A(\g.we_clk [2062]));
Q_ASSIGN U14329 ( .B(clk), .A(\g.we_clk [2061]));
Q_ASSIGN U14330 ( .B(clk), .A(\g.we_clk [2060]));
Q_ASSIGN U14331 ( .B(clk), .A(\g.we_clk [2059]));
Q_ASSIGN U14332 ( .B(clk), .A(\g.we_clk [2058]));
Q_ASSIGN U14333 ( .B(clk), .A(\g.we_clk [2057]));
Q_ASSIGN U14334 ( .B(clk), .A(\g.we_clk [2056]));
Q_ASSIGN U14335 ( .B(clk), .A(\g.we_clk [2055]));
Q_ASSIGN U14336 ( .B(clk), .A(\g.we_clk [2054]));
Q_ASSIGN U14337 ( .B(clk), .A(\g.we_clk [2053]));
Q_ASSIGN U14338 ( .B(clk), .A(\g.we_clk [2052]));
Q_ASSIGN U14339 ( .B(clk), .A(\g.we_clk [2051]));
Q_ASSIGN U14340 ( .B(clk), .A(\g.we_clk [2050]));
Q_ASSIGN U14341 ( .B(clk), .A(\g.we_clk [2049]));
Q_ASSIGN U14342 ( .B(clk), .A(\g.we_clk [2048]));
Q_ASSIGN U14343 ( .B(clk), .A(\g.we_clk [2047]));
Q_ASSIGN U14344 ( .B(clk), .A(\g.we_clk [2046]));
Q_ASSIGN U14345 ( .B(clk), .A(\g.we_clk [2045]));
Q_ASSIGN U14346 ( .B(clk), .A(\g.we_clk [2044]));
Q_ASSIGN U14347 ( .B(clk), .A(\g.we_clk [2043]));
Q_ASSIGN U14348 ( .B(clk), .A(\g.we_clk [2042]));
Q_ASSIGN U14349 ( .B(clk), .A(\g.we_clk [2041]));
Q_ASSIGN U14350 ( .B(clk), .A(\g.we_clk [2040]));
Q_ASSIGN U14351 ( .B(clk), .A(\g.we_clk [2039]));
Q_ASSIGN U14352 ( .B(clk), .A(\g.we_clk [2038]));
Q_ASSIGN U14353 ( .B(clk), .A(\g.we_clk [2037]));
Q_ASSIGN U14354 ( .B(clk), .A(\g.we_clk [2036]));
Q_ASSIGN U14355 ( .B(clk), .A(\g.we_clk [2035]));
Q_ASSIGN U14356 ( .B(clk), .A(\g.we_clk [2034]));
Q_ASSIGN U14357 ( .B(clk), .A(\g.we_clk [2033]));
Q_ASSIGN U14358 ( .B(clk), .A(\g.we_clk [2032]));
Q_ASSIGN U14359 ( .B(clk), .A(\g.we_clk [2031]));
Q_ASSIGN U14360 ( .B(clk), .A(\g.we_clk [2030]));
Q_ASSIGN U14361 ( .B(clk), .A(\g.we_clk [2029]));
Q_ASSIGN U14362 ( .B(clk), .A(\g.we_clk [2028]));
Q_ASSIGN U14363 ( .B(clk), .A(\g.we_clk [2027]));
Q_ASSIGN U14364 ( .B(clk), .A(\g.we_clk [2026]));
Q_ASSIGN U14365 ( .B(clk), .A(\g.we_clk [2025]));
Q_ASSIGN U14366 ( .B(clk), .A(\g.we_clk [2024]));
Q_ASSIGN U14367 ( .B(clk), .A(\g.we_clk [2023]));
Q_ASSIGN U14368 ( .B(clk), .A(\g.we_clk [2022]));
Q_ASSIGN U14369 ( .B(clk), .A(\g.we_clk [2021]));
Q_ASSIGN U14370 ( .B(clk), .A(\g.we_clk [2020]));
Q_ASSIGN U14371 ( .B(clk), .A(\g.we_clk [2019]));
Q_ASSIGN U14372 ( .B(clk), .A(\g.we_clk [2018]));
Q_ASSIGN U14373 ( .B(clk), .A(\g.we_clk [2017]));
Q_ASSIGN U14374 ( .B(clk), .A(\g.we_clk [2016]));
Q_ASSIGN U14375 ( .B(clk), .A(\g.we_clk [2015]));
Q_ASSIGN U14376 ( .B(clk), .A(\g.we_clk [2014]));
Q_ASSIGN U14377 ( .B(clk), .A(\g.we_clk [2013]));
Q_ASSIGN U14378 ( .B(clk), .A(\g.we_clk [2012]));
Q_ASSIGN U14379 ( .B(clk), .A(\g.we_clk [2011]));
Q_ASSIGN U14380 ( .B(clk), .A(\g.we_clk [2010]));
Q_ASSIGN U14381 ( .B(clk), .A(\g.we_clk [2009]));
Q_ASSIGN U14382 ( .B(clk), .A(\g.we_clk [2008]));
Q_ASSIGN U14383 ( .B(clk), .A(\g.we_clk [2007]));
Q_ASSIGN U14384 ( .B(clk), .A(\g.we_clk [2006]));
Q_ASSIGN U14385 ( .B(clk), .A(\g.we_clk [2005]));
Q_ASSIGN U14386 ( .B(clk), .A(\g.we_clk [2004]));
Q_ASSIGN U14387 ( .B(clk), .A(\g.we_clk [2003]));
Q_ASSIGN U14388 ( .B(clk), .A(\g.we_clk [2002]));
Q_ASSIGN U14389 ( .B(clk), .A(\g.we_clk [2001]));
Q_ASSIGN U14390 ( .B(clk), .A(\g.we_clk [2000]));
Q_ASSIGN U14391 ( .B(clk), .A(\g.we_clk [1999]));
Q_ASSIGN U14392 ( .B(clk), .A(\g.we_clk [1998]));
Q_ASSIGN U14393 ( .B(clk), .A(\g.we_clk [1997]));
Q_ASSIGN U14394 ( .B(clk), .A(\g.we_clk [1996]));
Q_ASSIGN U14395 ( .B(clk), .A(\g.we_clk [1995]));
Q_ASSIGN U14396 ( .B(clk), .A(\g.we_clk [1994]));
Q_ASSIGN U14397 ( .B(clk), .A(\g.we_clk [1993]));
Q_ASSIGN U14398 ( .B(clk), .A(\g.we_clk [1992]));
Q_ASSIGN U14399 ( .B(clk), .A(\g.we_clk [1991]));
Q_ASSIGN U14400 ( .B(clk), .A(\g.we_clk [1990]));
Q_ASSIGN U14401 ( .B(clk), .A(\g.we_clk [1989]));
Q_ASSIGN U14402 ( .B(clk), .A(\g.we_clk [1988]));
Q_ASSIGN U14403 ( .B(clk), .A(\g.we_clk [1987]));
Q_ASSIGN U14404 ( .B(clk), .A(\g.we_clk [1986]));
Q_ASSIGN U14405 ( .B(clk), .A(\g.we_clk [1985]));
Q_ASSIGN U14406 ( .B(clk), .A(\g.we_clk [1984]));
Q_ASSIGN U14407 ( .B(clk), .A(\g.we_clk [1983]));
Q_ASSIGN U14408 ( .B(clk), .A(\g.we_clk [1982]));
Q_ASSIGN U14409 ( .B(clk), .A(\g.we_clk [1981]));
Q_ASSIGN U14410 ( .B(clk), .A(\g.we_clk [1980]));
Q_ASSIGN U14411 ( .B(clk), .A(\g.we_clk [1979]));
Q_ASSIGN U14412 ( .B(clk), .A(\g.we_clk [1978]));
Q_ASSIGN U14413 ( .B(clk), .A(\g.we_clk [1977]));
Q_ASSIGN U14414 ( .B(clk), .A(\g.we_clk [1976]));
Q_ASSIGN U14415 ( .B(clk), .A(\g.we_clk [1975]));
Q_ASSIGN U14416 ( .B(clk), .A(\g.we_clk [1974]));
Q_ASSIGN U14417 ( .B(clk), .A(\g.we_clk [1973]));
Q_ASSIGN U14418 ( .B(clk), .A(\g.we_clk [1972]));
Q_ASSIGN U14419 ( .B(clk), .A(\g.we_clk [1971]));
Q_ASSIGN U14420 ( .B(clk), .A(\g.we_clk [1970]));
Q_ASSIGN U14421 ( .B(clk), .A(\g.we_clk [1969]));
Q_ASSIGN U14422 ( .B(clk), .A(\g.we_clk [1968]));
Q_ASSIGN U14423 ( .B(clk), .A(\g.we_clk [1967]));
Q_ASSIGN U14424 ( .B(clk), .A(\g.we_clk [1966]));
Q_ASSIGN U14425 ( .B(clk), .A(\g.we_clk [1965]));
Q_ASSIGN U14426 ( .B(clk), .A(\g.we_clk [1964]));
Q_ASSIGN U14427 ( .B(clk), .A(\g.we_clk [1963]));
Q_ASSIGN U14428 ( .B(clk), .A(\g.we_clk [1962]));
Q_ASSIGN U14429 ( .B(clk), .A(\g.we_clk [1961]));
Q_ASSIGN U14430 ( .B(clk), .A(\g.we_clk [1960]));
Q_ASSIGN U14431 ( .B(clk), .A(\g.we_clk [1959]));
Q_ASSIGN U14432 ( .B(clk), .A(\g.we_clk [1958]));
Q_ASSIGN U14433 ( .B(clk), .A(\g.we_clk [1957]));
Q_ASSIGN U14434 ( .B(clk), .A(\g.we_clk [1956]));
Q_ASSIGN U14435 ( .B(clk), .A(\g.we_clk [1955]));
Q_ASSIGN U14436 ( .B(clk), .A(\g.we_clk [1954]));
Q_ASSIGN U14437 ( .B(clk), .A(\g.we_clk [1953]));
Q_ASSIGN U14438 ( .B(clk), .A(\g.we_clk [1952]));
Q_ASSIGN U14439 ( .B(clk), .A(\g.we_clk [1951]));
Q_ASSIGN U14440 ( .B(clk), .A(\g.we_clk [1950]));
Q_ASSIGN U14441 ( .B(clk), .A(\g.we_clk [1949]));
Q_ASSIGN U14442 ( .B(clk), .A(\g.we_clk [1948]));
Q_ASSIGN U14443 ( .B(clk), .A(\g.we_clk [1947]));
Q_ASSIGN U14444 ( .B(clk), .A(\g.we_clk [1946]));
Q_ASSIGN U14445 ( .B(clk), .A(\g.we_clk [1945]));
Q_ASSIGN U14446 ( .B(clk), .A(\g.we_clk [1944]));
Q_ASSIGN U14447 ( .B(clk), .A(\g.we_clk [1943]));
Q_ASSIGN U14448 ( .B(clk), .A(\g.we_clk [1942]));
Q_ASSIGN U14449 ( .B(clk), .A(\g.we_clk [1941]));
Q_ASSIGN U14450 ( .B(clk), .A(\g.we_clk [1940]));
Q_ASSIGN U14451 ( .B(clk), .A(\g.we_clk [1939]));
Q_ASSIGN U14452 ( .B(clk), .A(\g.we_clk [1938]));
Q_ASSIGN U14453 ( .B(clk), .A(\g.we_clk [1937]));
Q_ASSIGN U14454 ( .B(clk), .A(\g.we_clk [1936]));
Q_ASSIGN U14455 ( .B(clk), .A(\g.we_clk [1935]));
Q_ASSIGN U14456 ( .B(clk), .A(\g.we_clk [1934]));
Q_ASSIGN U14457 ( .B(clk), .A(\g.we_clk [1933]));
Q_ASSIGN U14458 ( .B(clk), .A(\g.we_clk [1932]));
Q_ASSIGN U14459 ( .B(clk), .A(\g.we_clk [1931]));
Q_ASSIGN U14460 ( .B(clk), .A(\g.we_clk [1930]));
Q_ASSIGN U14461 ( .B(clk), .A(\g.we_clk [1929]));
Q_ASSIGN U14462 ( .B(clk), .A(\g.we_clk [1928]));
Q_ASSIGN U14463 ( .B(clk), .A(\g.we_clk [1927]));
Q_ASSIGN U14464 ( .B(clk), .A(\g.we_clk [1926]));
Q_ASSIGN U14465 ( .B(clk), .A(\g.we_clk [1925]));
Q_ASSIGN U14466 ( .B(clk), .A(\g.we_clk [1924]));
Q_ASSIGN U14467 ( .B(clk), .A(\g.we_clk [1923]));
Q_ASSIGN U14468 ( .B(clk), .A(\g.we_clk [1922]));
Q_ASSIGN U14469 ( .B(clk), .A(\g.we_clk [1921]));
Q_ASSIGN U14470 ( .B(clk), .A(\g.we_clk [1920]));
Q_ASSIGN U14471 ( .B(clk), .A(\g.we_clk [1919]));
Q_ASSIGN U14472 ( .B(clk), .A(\g.we_clk [1918]));
Q_ASSIGN U14473 ( .B(clk), .A(\g.we_clk [1917]));
Q_ASSIGN U14474 ( .B(clk), .A(\g.we_clk [1916]));
Q_ASSIGN U14475 ( .B(clk), .A(\g.we_clk [1915]));
Q_ASSIGN U14476 ( .B(clk), .A(\g.we_clk [1914]));
Q_ASSIGN U14477 ( .B(clk), .A(\g.we_clk [1913]));
Q_ASSIGN U14478 ( .B(clk), .A(\g.we_clk [1912]));
Q_ASSIGN U14479 ( .B(clk), .A(\g.we_clk [1911]));
Q_ASSIGN U14480 ( .B(clk), .A(\g.we_clk [1910]));
Q_ASSIGN U14481 ( .B(clk), .A(\g.we_clk [1909]));
Q_ASSIGN U14482 ( .B(clk), .A(\g.we_clk [1908]));
Q_ASSIGN U14483 ( .B(clk), .A(\g.we_clk [1907]));
Q_ASSIGN U14484 ( .B(clk), .A(\g.we_clk [1906]));
Q_ASSIGN U14485 ( .B(clk), .A(\g.we_clk [1905]));
Q_ASSIGN U14486 ( .B(clk), .A(\g.we_clk [1904]));
Q_ASSIGN U14487 ( .B(clk), .A(\g.we_clk [1903]));
Q_ASSIGN U14488 ( .B(clk), .A(\g.we_clk [1902]));
Q_ASSIGN U14489 ( .B(clk), .A(\g.we_clk [1901]));
Q_ASSIGN U14490 ( .B(clk), .A(\g.we_clk [1900]));
Q_ASSIGN U14491 ( .B(clk), .A(\g.we_clk [1899]));
Q_ASSIGN U14492 ( .B(clk), .A(\g.we_clk [1898]));
Q_ASSIGN U14493 ( .B(clk), .A(\g.we_clk [1897]));
Q_ASSIGN U14494 ( .B(clk), .A(\g.we_clk [1896]));
Q_ASSIGN U14495 ( .B(clk), .A(\g.we_clk [1895]));
Q_ASSIGN U14496 ( .B(clk), .A(\g.we_clk [1894]));
Q_ASSIGN U14497 ( .B(clk), .A(\g.we_clk [1893]));
Q_ASSIGN U14498 ( .B(clk), .A(\g.we_clk [1892]));
Q_ASSIGN U14499 ( .B(clk), .A(\g.we_clk [1891]));
Q_ASSIGN U14500 ( .B(clk), .A(\g.we_clk [1890]));
Q_ASSIGN U14501 ( .B(clk), .A(\g.we_clk [1889]));
Q_ASSIGN U14502 ( .B(clk), .A(\g.we_clk [1888]));
Q_ASSIGN U14503 ( .B(clk), .A(\g.we_clk [1887]));
Q_ASSIGN U14504 ( .B(clk), .A(\g.we_clk [1886]));
Q_ASSIGN U14505 ( .B(clk), .A(\g.we_clk [1885]));
Q_ASSIGN U14506 ( .B(clk), .A(\g.we_clk [1884]));
Q_ASSIGN U14507 ( .B(clk), .A(\g.we_clk [1883]));
Q_ASSIGN U14508 ( .B(clk), .A(\g.we_clk [1882]));
Q_ASSIGN U14509 ( .B(clk), .A(\g.we_clk [1881]));
Q_ASSIGN U14510 ( .B(clk), .A(\g.we_clk [1880]));
Q_ASSIGN U14511 ( .B(clk), .A(\g.we_clk [1879]));
Q_ASSIGN U14512 ( .B(clk), .A(\g.we_clk [1878]));
Q_ASSIGN U14513 ( .B(clk), .A(\g.we_clk [1877]));
Q_ASSIGN U14514 ( .B(clk), .A(\g.we_clk [1876]));
Q_ASSIGN U14515 ( .B(clk), .A(\g.we_clk [1875]));
Q_ASSIGN U14516 ( .B(clk), .A(\g.we_clk [1874]));
Q_ASSIGN U14517 ( .B(clk), .A(\g.we_clk [1873]));
Q_ASSIGN U14518 ( .B(clk), .A(\g.we_clk [1872]));
Q_ASSIGN U14519 ( .B(clk), .A(\g.we_clk [1871]));
Q_ASSIGN U14520 ( .B(clk), .A(\g.we_clk [1870]));
Q_ASSIGN U14521 ( .B(clk), .A(\g.we_clk [1869]));
Q_ASSIGN U14522 ( .B(clk), .A(\g.we_clk [1868]));
Q_ASSIGN U14523 ( .B(clk), .A(\g.we_clk [1867]));
Q_ASSIGN U14524 ( .B(clk), .A(\g.we_clk [1866]));
Q_ASSIGN U14525 ( .B(clk), .A(\g.we_clk [1865]));
Q_ASSIGN U14526 ( .B(clk), .A(\g.we_clk [1864]));
Q_ASSIGN U14527 ( .B(clk), .A(\g.we_clk [1863]));
Q_ASSIGN U14528 ( .B(clk), .A(\g.we_clk [1862]));
Q_ASSIGN U14529 ( .B(clk), .A(\g.we_clk [1861]));
Q_ASSIGN U14530 ( .B(clk), .A(\g.we_clk [1860]));
Q_ASSIGN U14531 ( .B(clk), .A(\g.we_clk [1859]));
Q_ASSIGN U14532 ( .B(clk), .A(\g.we_clk [1858]));
Q_ASSIGN U14533 ( .B(clk), .A(\g.we_clk [1857]));
Q_ASSIGN U14534 ( .B(clk), .A(\g.we_clk [1856]));
Q_ASSIGN U14535 ( .B(clk), .A(\g.we_clk [1855]));
Q_ASSIGN U14536 ( .B(clk), .A(\g.we_clk [1854]));
Q_ASSIGN U14537 ( .B(clk), .A(\g.we_clk [1853]));
Q_ASSIGN U14538 ( .B(clk), .A(\g.we_clk [1852]));
Q_ASSIGN U14539 ( .B(clk), .A(\g.we_clk [1851]));
Q_ASSIGN U14540 ( .B(clk), .A(\g.we_clk [1850]));
Q_ASSIGN U14541 ( .B(clk), .A(\g.we_clk [1849]));
Q_ASSIGN U14542 ( .B(clk), .A(\g.we_clk [1848]));
Q_ASSIGN U14543 ( .B(clk), .A(\g.we_clk [1847]));
Q_ASSIGN U14544 ( .B(clk), .A(\g.we_clk [1846]));
Q_ASSIGN U14545 ( .B(clk), .A(\g.we_clk [1845]));
Q_ASSIGN U14546 ( .B(clk), .A(\g.we_clk [1844]));
Q_ASSIGN U14547 ( .B(clk), .A(\g.we_clk [1843]));
Q_ASSIGN U14548 ( .B(clk), .A(\g.we_clk [1842]));
Q_ASSIGN U14549 ( .B(clk), .A(\g.we_clk [1841]));
Q_ASSIGN U14550 ( .B(clk), .A(\g.we_clk [1840]));
Q_ASSIGN U14551 ( .B(clk), .A(\g.we_clk [1839]));
Q_ASSIGN U14552 ( .B(clk), .A(\g.we_clk [1838]));
Q_ASSIGN U14553 ( .B(clk), .A(\g.we_clk [1837]));
Q_ASSIGN U14554 ( .B(clk), .A(\g.we_clk [1836]));
Q_ASSIGN U14555 ( .B(clk), .A(\g.we_clk [1835]));
Q_ASSIGN U14556 ( .B(clk), .A(\g.we_clk [1834]));
Q_ASSIGN U14557 ( .B(clk), .A(\g.we_clk [1833]));
Q_ASSIGN U14558 ( .B(clk), .A(\g.we_clk [1832]));
Q_ASSIGN U14559 ( .B(clk), .A(\g.we_clk [1831]));
Q_ASSIGN U14560 ( .B(clk), .A(\g.we_clk [1830]));
Q_ASSIGN U14561 ( .B(clk), .A(\g.we_clk [1829]));
Q_ASSIGN U14562 ( .B(clk), .A(\g.we_clk [1828]));
Q_ASSIGN U14563 ( .B(clk), .A(\g.we_clk [1827]));
Q_ASSIGN U14564 ( .B(clk), .A(\g.we_clk [1826]));
Q_ASSIGN U14565 ( .B(clk), .A(\g.we_clk [1825]));
Q_ASSIGN U14566 ( .B(clk), .A(\g.we_clk [1824]));
Q_ASSIGN U14567 ( .B(clk), .A(\g.we_clk [1823]));
Q_ASSIGN U14568 ( .B(clk), .A(\g.we_clk [1822]));
Q_ASSIGN U14569 ( .B(clk), .A(\g.we_clk [1821]));
Q_ASSIGN U14570 ( .B(clk), .A(\g.we_clk [1820]));
Q_ASSIGN U14571 ( .B(clk), .A(\g.we_clk [1819]));
Q_ASSIGN U14572 ( .B(clk), .A(\g.we_clk [1818]));
Q_ASSIGN U14573 ( .B(clk), .A(\g.we_clk [1817]));
Q_ASSIGN U14574 ( .B(clk), .A(\g.we_clk [1816]));
Q_ASSIGN U14575 ( .B(clk), .A(\g.we_clk [1815]));
Q_ASSIGN U14576 ( .B(clk), .A(\g.we_clk [1814]));
Q_ASSIGN U14577 ( .B(clk), .A(\g.we_clk [1813]));
Q_ASSIGN U14578 ( .B(clk), .A(\g.we_clk [1812]));
Q_ASSIGN U14579 ( .B(clk), .A(\g.we_clk [1811]));
Q_ASSIGN U14580 ( .B(clk), .A(\g.we_clk [1810]));
Q_ASSIGN U14581 ( .B(clk), .A(\g.we_clk [1809]));
Q_ASSIGN U14582 ( .B(clk), .A(\g.we_clk [1808]));
Q_ASSIGN U14583 ( .B(clk), .A(\g.we_clk [1807]));
Q_ASSIGN U14584 ( .B(clk), .A(\g.we_clk [1806]));
Q_ASSIGN U14585 ( .B(clk), .A(\g.we_clk [1805]));
Q_ASSIGN U14586 ( .B(clk), .A(\g.we_clk [1804]));
Q_ASSIGN U14587 ( .B(clk), .A(\g.we_clk [1803]));
Q_ASSIGN U14588 ( .B(clk), .A(\g.we_clk [1802]));
Q_ASSIGN U14589 ( .B(clk), .A(\g.we_clk [1801]));
Q_ASSIGN U14590 ( .B(clk), .A(\g.we_clk [1800]));
Q_ASSIGN U14591 ( .B(clk), .A(\g.we_clk [1799]));
Q_ASSIGN U14592 ( .B(clk), .A(\g.we_clk [1798]));
Q_ASSIGN U14593 ( .B(clk), .A(\g.we_clk [1797]));
Q_ASSIGN U14594 ( .B(clk), .A(\g.we_clk [1796]));
Q_ASSIGN U14595 ( .B(clk), .A(\g.we_clk [1795]));
Q_ASSIGN U14596 ( .B(clk), .A(\g.we_clk [1794]));
Q_ASSIGN U14597 ( .B(clk), .A(\g.we_clk [1793]));
Q_ASSIGN U14598 ( .B(clk), .A(\g.we_clk [1792]));
Q_ASSIGN U14599 ( .B(clk), .A(\g.we_clk [1791]));
Q_ASSIGN U14600 ( .B(clk), .A(\g.we_clk [1790]));
Q_ASSIGN U14601 ( .B(clk), .A(\g.we_clk [1789]));
Q_ASSIGN U14602 ( .B(clk), .A(\g.we_clk [1788]));
Q_ASSIGN U14603 ( .B(clk), .A(\g.we_clk [1787]));
Q_ASSIGN U14604 ( .B(clk), .A(\g.we_clk [1786]));
Q_ASSIGN U14605 ( .B(clk), .A(\g.we_clk [1785]));
Q_ASSIGN U14606 ( .B(clk), .A(\g.we_clk [1784]));
Q_ASSIGN U14607 ( .B(clk), .A(\g.we_clk [1783]));
Q_ASSIGN U14608 ( .B(clk), .A(\g.we_clk [1782]));
Q_ASSIGN U14609 ( .B(clk), .A(\g.we_clk [1781]));
Q_ASSIGN U14610 ( .B(clk), .A(\g.we_clk [1780]));
Q_ASSIGN U14611 ( .B(clk), .A(\g.we_clk [1779]));
Q_ASSIGN U14612 ( .B(clk), .A(\g.we_clk [1778]));
Q_ASSIGN U14613 ( .B(clk), .A(\g.we_clk [1777]));
Q_ASSIGN U14614 ( .B(clk), .A(\g.we_clk [1776]));
Q_ASSIGN U14615 ( .B(clk), .A(\g.we_clk [1775]));
Q_ASSIGN U14616 ( .B(clk), .A(\g.we_clk [1774]));
Q_ASSIGN U14617 ( .B(clk), .A(\g.we_clk [1773]));
Q_ASSIGN U14618 ( .B(clk), .A(\g.we_clk [1772]));
Q_ASSIGN U14619 ( .B(clk), .A(\g.we_clk [1771]));
Q_ASSIGN U14620 ( .B(clk), .A(\g.we_clk [1770]));
Q_ASSIGN U14621 ( .B(clk), .A(\g.we_clk [1769]));
Q_ASSIGN U14622 ( .B(clk), .A(\g.we_clk [1768]));
Q_ASSIGN U14623 ( .B(clk), .A(\g.we_clk [1767]));
Q_ASSIGN U14624 ( .B(clk), .A(\g.we_clk [1766]));
Q_ASSIGN U14625 ( .B(clk), .A(\g.we_clk [1765]));
Q_ASSIGN U14626 ( .B(clk), .A(\g.we_clk [1764]));
Q_ASSIGN U14627 ( .B(clk), .A(\g.we_clk [1763]));
Q_ASSIGN U14628 ( .B(clk), .A(\g.we_clk [1762]));
Q_ASSIGN U14629 ( .B(clk), .A(\g.we_clk [1761]));
Q_ASSIGN U14630 ( .B(clk), .A(\g.we_clk [1760]));
Q_ASSIGN U14631 ( .B(clk), .A(\g.we_clk [1759]));
Q_ASSIGN U14632 ( .B(clk), .A(\g.we_clk [1758]));
Q_ASSIGN U14633 ( .B(clk), .A(\g.we_clk [1757]));
Q_ASSIGN U14634 ( .B(clk), .A(\g.we_clk [1756]));
Q_ASSIGN U14635 ( .B(clk), .A(\g.we_clk [1755]));
Q_ASSIGN U14636 ( .B(clk), .A(\g.we_clk [1754]));
Q_ASSIGN U14637 ( .B(clk), .A(\g.we_clk [1753]));
Q_ASSIGN U14638 ( .B(clk), .A(\g.we_clk [1752]));
Q_ASSIGN U14639 ( .B(clk), .A(\g.we_clk [1751]));
Q_ASSIGN U14640 ( .B(clk), .A(\g.we_clk [1750]));
Q_ASSIGN U14641 ( .B(clk), .A(\g.we_clk [1749]));
Q_ASSIGN U14642 ( .B(clk), .A(\g.we_clk [1748]));
Q_ASSIGN U14643 ( .B(clk), .A(\g.we_clk [1747]));
Q_ASSIGN U14644 ( .B(clk), .A(\g.we_clk [1746]));
Q_ASSIGN U14645 ( .B(clk), .A(\g.we_clk [1745]));
Q_ASSIGN U14646 ( .B(clk), .A(\g.we_clk [1744]));
Q_ASSIGN U14647 ( .B(clk), .A(\g.we_clk [1743]));
Q_ASSIGN U14648 ( .B(clk), .A(\g.we_clk [1742]));
Q_ASSIGN U14649 ( .B(clk), .A(\g.we_clk [1741]));
Q_ASSIGN U14650 ( .B(clk), .A(\g.we_clk [1740]));
Q_ASSIGN U14651 ( .B(clk), .A(\g.we_clk [1739]));
Q_ASSIGN U14652 ( .B(clk), .A(\g.we_clk [1738]));
Q_ASSIGN U14653 ( .B(clk), .A(\g.we_clk [1737]));
Q_ASSIGN U14654 ( .B(clk), .A(\g.we_clk [1736]));
Q_ASSIGN U14655 ( .B(clk), .A(\g.we_clk [1735]));
Q_ASSIGN U14656 ( .B(clk), .A(\g.we_clk [1734]));
Q_ASSIGN U14657 ( .B(clk), .A(\g.we_clk [1733]));
Q_ASSIGN U14658 ( .B(clk), .A(\g.we_clk [1732]));
Q_ASSIGN U14659 ( .B(clk), .A(\g.we_clk [1731]));
Q_ASSIGN U14660 ( .B(clk), .A(\g.we_clk [1730]));
Q_ASSIGN U14661 ( .B(clk), .A(\g.we_clk [1729]));
Q_ASSIGN U14662 ( .B(clk), .A(\g.we_clk [1728]));
Q_ASSIGN U14663 ( .B(clk), .A(\g.we_clk [1727]));
Q_ASSIGN U14664 ( .B(clk), .A(\g.we_clk [1726]));
Q_ASSIGN U14665 ( .B(clk), .A(\g.we_clk [1725]));
Q_ASSIGN U14666 ( .B(clk), .A(\g.we_clk [1724]));
Q_ASSIGN U14667 ( .B(clk), .A(\g.we_clk [1723]));
Q_ASSIGN U14668 ( .B(clk), .A(\g.we_clk [1722]));
Q_ASSIGN U14669 ( .B(clk), .A(\g.we_clk [1721]));
Q_ASSIGN U14670 ( .B(clk), .A(\g.we_clk [1720]));
Q_ASSIGN U14671 ( .B(clk), .A(\g.we_clk [1719]));
Q_ASSIGN U14672 ( .B(clk), .A(\g.we_clk [1718]));
Q_ASSIGN U14673 ( .B(clk), .A(\g.we_clk [1717]));
Q_ASSIGN U14674 ( .B(clk), .A(\g.we_clk [1716]));
Q_ASSIGN U14675 ( .B(clk), .A(\g.we_clk [1715]));
Q_ASSIGN U14676 ( .B(clk), .A(\g.we_clk [1714]));
Q_ASSIGN U14677 ( .B(clk), .A(\g.we_clk [1713]));
Q_ASSIGN U14678 ( .B(clk), .A(\g.we_clk [1712]));
Q_ASSIGN U14679 ( .B(clk), .A(\g.we_clk [1711]));
Q_ASSIGN U14680 ( .B(clk), .A(\g.we_clk [1710]));
Q_ASSIGN U14681 ( .B(clk), .A(\g.we_clk [1709]));
Q_ASSIGN U14682 ( .B(clk), .A(\g.we_clk [1708]));
Q_ASSIGN U14683 ( .B(clk), .A(\g.we_clk [1707]));
Q_ASSIGN U14684 ( .B(clk), .A(\g.we_clk [1706]));
Q_ASSIGN U14685 ( .B(clk), .A(\g.we_clk [1705]));
Q_ASSIGN U14686 ( .B(clk), .A(\g.we_clk [1704]));
Q_ASSIGN U14687 ( .B(clk), .A(\g.we_clk [1703]));
Q_ASSIGN U14688 ( .B(clk), .A(\g.we_clk [1702]));
Q_ASSIGN U14689 ( .B(clk), .A(\g.we_clk [1701]));
Q_ASSIGN U14690 ( .B(clk), .A(\g.we_clk [1700]));
Q_ASSIGN U14691 ( .B(clk), .A(\g.we_clk [1699]));
Q_ASSIGN U14692 ( .B(clk), .A(\g.we_clk [1698]));
Q_ASSIGN U14693 ( .B(clk), .A(\g.we_clk [1697]));
Q_ASSIGN U14694 ( .B(clk), .A(\g.we_clk [1696]));
Q_ASSIGN U14695 ( .B(clk), .A(\g.we_clk [1695]));
Q_ASSIGN U14696 ( .B(clk), .A(\g.we_clk [1694]));
Q_ASSIGN U14697 ( .B(clk), .A(\g.we_clk [1693]));
Q_ASSIGN U14698 ( .B(clk), .A(\g.we_clk [1692]));
Q_ASSIGN U14699 ( .B(clk), .A(\g.we_clk [1691]));
Q_ASSIGN U14700 ( .B(clk), .A(\g.we_clk [1690]));
Q_ASSIGN U14701 ( .B(clk), .A(\g.we_clk [1689]));
Q_ASSIGN U14702 ( .B(clk), .A(\g.we_clk [1688]));
Q_ASSIGN U14703 ( .B(clk), .A(\g.we_clk [1687]));
Q_ASSIGN U14704 ( .B(clk), .A(\g.we_clk [1686]));
Q_ASSIGN U14705 ( .B(clk), .A(\g.we_clk [1685]));
Q_ASSIGN U14706 ( .B(clk), .A(\g.we_clk [1684]));
Q_ASSIGN U14707 ( .B(clk), .A(\g.we_clk [1683]));
Q_ASSIGN U14708 ( .B(clk), .A(\g.we_clk [1682]));
Q_ASSIGN U14709 ( .B(clk), .A(\g.we_clk [1681]));
Q_ASSIGN U14710 ( .B(clk), .A(\g.we_clk [1680]));
Q_ASSIGN U14711 ( .B(clk), .A(\g.we_clk [1679]));
Q_ASSIGN U14712 ( .B(clk), .A(\g.we_clk [1678]));
Q_ASSIGN U14713 ( .B(clk), .A(\g.we_clk [1677]));
Q_ASSIGN U14714 ( .B(clk), .A(\g.we_clk [1676]));
Q_ASSIGN U14715 ( .B(clk), .A(\g.we_clk [1675]));
Q_ASSIGN U14716 ( .B(clk), .A(\g.we_clk [1674]));
Q_ASSIGN U14717 ( .B(clk), .A(\g.we_clk [1673]));
Q_ASSIGN U14718 ( .B(clk), .A(\g.we_clk [1672]));
Q_ASSIGN U14719 ( .B(clk), .A(\g.we_clk [1671]));
Q_ASSIGN U14720 ( .B(clk), .A(\g.we_clk [1670]));
Q_ASSIGN U14721 ( .B(clk), .A(\g.we_clk [1669]));
Q_ASSIGN U14722 ( .B(clk), .A(\g.we_clk [1668]));
Q_ASSIGN U14723 ( .B(clk), .A(\g.we_clk [1667]));
Q_ASSIGN U14724 ( .B(clk), .A(\g.we_clk [1666]));
Q_ASSIGN U14725 ( .B(clk), .A(\g.we_clk [1665]));
Q_ASSIGN U14726 ( .B(clk), .A(\g.we_clk [1664]));
Q_ASSIGN U14727 ( .B(clk), .A(\g.we_clk [1663]));
Q_ASSIGN U14728 ( .B(clk), .A(\g.we_clk [1662]));
Q_ASSIGN U14729 ( .B(clk), .A(\g.we_clk [1661]));
Q_ASSIGN U14730 ( .B(clk), .A(\g.we_clk [1660]));
Q_ASSIGN U14731 ( .B(clk), .A(\g.we_clk [1659]));
Q_ASSIGN U14732 ( .B(clk), .A(\g.we_clk [1658]));
Q_ASSIGN U14733 ( .B(clk), .A(\g.we_clk [1657]));
Q_ASSIGN U14734 ( .B(clk), .A(\g.we_clk [1656]));
Q_ASSIGN U14735 ( .B(clk), .A(\g.we_clk [1655]));
Q_ASSIGN U14736 ( .B(clk), .A(\g.we_clk [1654]));
Q_ASSIGN U14737 ( .B(clk), .A(\g.we_clk [1653]));
Q_ASSIGN U14738 ( .B(clk), .A(\g.we_clk [1652]));
Q_ASSIGN U14739 ( .B(clk), .A(\g.we_clk [1651]));
Q_ASSIGN U14740 ( .B(clk), .A(\g.we_clk [1650]));
Q_ASSIGN U14741 ( .B(clk), .A(\g.we_clk [1649]));
Q_ASSIGN U14742 ( .B(clk), .A(\g.we_clk [1648]));
Q_ASSIGN U14743 ( .B(clk), .A(\g.we_clk [1647]));
Q_ASSIGN U14744 ( .B(clk), .A(\g.we_clk [1646]));
Q_ASSIGN U14745 ( .B(clk), .A(\g.we_clk [1645]));
Q_ASSIGN U14746 ( .B(clk), .A(\g.we_clk [1644]));
Q_ASSIGN U14747 ( .B(clk), .A(\g.we_clk [1643]));
Q_ASSIGN U14748 ( .B(clk), .A(\g.we_clk [1642]));
Q_ASSIGN U14749 ( .B(clk), .A(\g.we_clk [1641]));
Q_ASSIGN U14750 ( .B(clk), .A(\g.we_clk [1640]));
Q_ASSIGN U14751 ( .B(clk), .A(\g.we_clk [1639]));
Q_ASSIGN U14752 ( .B(clk), .A(\g.we_clk [1638]));
Q_ASSIGN U14753 ( .B(clk), .A(\g.we_clk [1637]));
Q_ASSIGN U14754 ( .B(clk), .A(\g.we_clk [1636]));
Q_ASSIGN U14755 ( .B(clk), .A(\g.we_clk [1635]));
Q_ASSIGN U14756 ( .B(clk), .A(\g.we_clk [1634]));
Q_ASSIGN U14757 ( .B(clk), .A(\g.we_clk [1633]));
Q_ASSIGN U14758 ( .B(clk), .A(\g.we_clk [1632]));
Q_ASSIGN U14759 ( .B(clk), .A(\g.we_clk [1631]));
Q_ASSIGN U14760 ( .B(clk), .A(\g.we_clk [1630]));
Q_ASSIGN U14761 ( .B(clk), .A(\g.we_clk [1629]));
Q_ASSIGN U14762 ( .B(clk), .A(\g.we_clk [1628]));
Q_ASSIGN U14763 ( .B(clk), .A(\g.we_clk [1627]));
Q_ASSIGN U14764 ( .B(clk), .A(\g.we_clk [1626]));
Q_ASSIGN U14765 ( .B(clk), .A(\g.we_clk [1625]));
Q_ASSIGN U14766 ( .B(clk), .A(\g.we_clk [1624]));
Q_ASSIGN U14767 ( .B(clk), .A(\g.we_clk [1623]));
Q_ASSIGN U14768 ( .B(clk), .A(\g.we_clk [1622]));
Q_ASSIGN U14769 ( .B(clk), .A(\g.we_clk [1621]));
Q_ASSIGN U14770 ( .B(clk), .A(\g.we_clk [1620]));
Q_ASSIGN U14771 ( .B(clk), .A(\g.we_clk [1619]));
Q_ASSIGN U14772 ( .B(clk), .A(\g.we_clk [1618]));
Q_ASSIGN U14773 ( .B(clk), .A(\g.we_clk [1617]));
Q_ASSIGN U14774 ( .B(clk), .A(\g.we_clk [1616]));
Q_ASSIGN U14775 ( .B(clk), .A(\g.we_clk [1615]));
Q_ASSIGN U14776 ( .B(clk), .A(\g.we_clk [1614]));
Q_ASSIGN U14777 ( .B(clk), .A(\g.we_clk [1613]));
Q_ASSIGN U14778 ( .B(clk), .A(\g.we_clk [1612]));
Q_ASSIGN U14779 ( .B(clk), .A(\g.we_clk [1611]));
Q_ASSIGN U14780 ( .B(clk), .A(\g.we_clk [1610]));
Q_ASSIGN U14781 ( .B(clk), .A(\g.we_clk [1609]));
Q_ASSIGN U14782 ( .B(clk), .A(\g.we_clk [1608]));
Q_ASSIGN U14783 ( .B(clk), .A(\g.we_clk [1607]));
Q_ASSIGN U14784 ( .B(clk), .A(\g.we_clk [1606]));
Q_ASSIGN U14785 ( .B(clk), .A(\g.we_clk [1605]));
Q_ASSIGN U14786 ( .B(clk), .A(\g.we_clk [1604]));
Q_ASSIGN U14787 ( .B(clk), .A(\g.we_clk [1603]));
Q_ASSIGN U14788 ( .B(clk), .A(\g.we_clk [1602]));
Q_ASSIGN U14789 ( .B(clk), .A(\g.we_clk [1601]));
Q_ASSIGN U14790 ( .B(clk), .A(\g.we_clk [1600]));
Q_ASSIGN U14791 ( .B(clk), .A(\g.we_clk [1599]));
Q_ASSIGN U14792 ( .B(clk), .A(\g.we_clk [1598]));
Q_ASSIGN U14793 ( .B(clk), .A(\g.we_clk [1597]));
Q_ASSIGN U14794 ( .B(clk), .A(\g.we_clk [1596]));
Q_ASSIGN U14795 ( .B(clk), .A(\g.we_clk [1595]));
Q_ASSIGN U14796 ( .B(clk), .A(\g.we_clk [1594]));
Q_ASSIGN U14797 ( .B(clk), .A(\g.we_clk [1593]));
Q_ASSIGN U14798 ( .B(clk), .A(\g.we_clk [1592]));
Q_ASSIGN U14799 ( .B(clk), .A(\g.we_clk [1591]));
Q_ASSIGN U14800 ( .B(clk), .A(\g.we_clk [1590]));
Q_ASSIGN U14801 ( .B(clk), .A(\g.we_clk [1589]));
Q_ASSIGN U14802 ( .B(clk), .A(\g.we_clk [1588]));
Q_ASSIGN U14803 ( .B(clk), .A(\g.we_clk [1587]));
Q_ASSIGN U14804 ( .B(clk), .A(\g.we_clk [1586]));
Q_ASSIGN U14805 ( .B(clk), .A(\g.we_clk [1585]));
Q_ASSIGN U14806 ( .B(clk), .A(\g.we_clk [1584]));
Q_ASSIGN U14807 ( .B(clk), .A(\g.we_clk [1583]));
Q_ASSIGN U14808 ( .B(clk), .A(\g.we_clk [1582]));
Q_ASSIGN U14809 ( .B(clk), .A(\g.we_clk [1581]));
Q_ASSIGN U14810 ( .B(clk), .A(\g.we_clk [1580]));
Q_ASSIGN U14811 ( .B(clk), .A(\g.we_clk [1579]));
Q_ASSIGN U14812 ( .B(clk), .A(\g.we_clk [1578]));
Q_ASSIGN U14813 ( .B(clk), .A(\g.we_clk [1577]));
Q_ASSIGN U14814 ( .B(clk), .A(\g.we_clk [1576]));
Q_ASSIGN U14815 ( .B(clk), .A(\g.we_clk [1575]));
Q_ASSIGN U14816 ( .B(clk), .A(\g.we_clk [1574]));
Q_ASSIGN U14817 ( .B(clk), .A(\g.we_clk [1573]));
Q_ASSIGN U14818 ( .B(clk), .A(\g.we_clk [1572]));
Q_ASSIGN U14819 ( .B(clk), .A(\g.we_clk [1571]));
Q_ASSIGN U14820 ( .B(clk), .A(\g.we_clk [1570]));
Q_ASSIGN U14821 ( .B(clk), .A(\g.we_clk [1569]));
Q_ASSIGN U14822 ( .B(clk), .A(\g.we_clk [1568]));
Q_ASSIGN U14823 ( .B(clk), .A(\g.we_clk [1567]));
Q_ASSIGN U14824 ( .B(clk), .A(\g.we_clk [1566]));
Q_ASSIGN U14825 ( .B(clk), .A(\g.we_clk [1565]));
Q_ASSIGN U14826 ( .B(clk), .A(\g.we_clk [1564]));
Q_ASSIGN U14827 ( .B(clk), .A(\g.we_clk [1563]));
Q_ASSIGN U14828 ( .B(clk), .A(\g.we_clk [1562]));
Q_ASSIGN U14829 ( .B(clk), .A(\g.we_clk [1561]));
Q_ASSIGN U14830 ( .B(clk), .A(\g.we_clk [1560]));
Q_ASSIGN U14831 ( .B(clk), .A(\g.we_clk [1559]));
Q_ASSIGN U14832 ( .B(clk), .A(\g.we_clk [1558]));
Q_ASSIGN U14833 ( .B(clk), .A(\g.we_clk [1557]));
Q_ASSIGN U14834 ( .B(clk), .A(\g.we_clk [1556]));
Q_ASSIGN U14835 ( .B(clk), .A(\g.we_clk [1555]));
Q_ASSIGN U14836 ( .B(clk), .A(\g.we_clk [1554]));
Q_ASSIGN U14837 ( .B(clk), .A(\g.we_clk [1553]));
Q_ASSIGN U14838 ( .B(clk), .A(\g.we_clk [1552]));
Q_ASSIGN U14839 ( .B(clk), .A(\g.we_clk [1551]));
Q_ASSIGN U14840 ( .B(clk), .A(\g.we_clk [1550]));
Q_ASSIGN U14841 ( .B(clk), .A(\g.we_clk [1549]));
Q_ASSIGN U14842 ( .B(clk), .A(\g.we_clk [1548]));
Q_ASSIGN U14843 ( .B(clk), .A(\g.we_clk [1547]));
Q_ASSIGN U14844 ( .B(clk), .A(\g.we_clk [1546]));
Q_ASSIGN U14845 ( .B(clk), .A(\g.we_clk [1545]));
Q_ASSIGN U14846 ( .B(clk), .A(\g.we_clk [1544]));
Q_ASSIGN U14847 ( .B(clk), .A(\g.we_clk [1543]));
Q_ASSIGN U14848 ( .B(clk), .A(\g.we_clk [1542]));
Q_ASSIGN U14849 ( .B(clk), .A(\g.we_clk [1541]));
Q_ASSIGN U14850 ( .B(clk), .A(\g.we_clk [1540]));
Q_ASSIGN U14851 ( .B(clk), .A(\g.we_clk [1539]));
Q_ASSIGN U14852 ( .B(clk), .A(\g.we_clk [1538]));
Q_ASSIGN U14853 ( .B(clk), .A(\g.we_clk [1537]));
Q_ASSIGN U14854 ( .B(clk), .A(\g.we_clk [1536]));
Q_ASSIGN U14855 ( .B(clk), .A(\g.we_clk [1535]));
Q_ASSIGN U14856 ( .B(clk), .A(\g.we_clk [1534]));
Q_ASSIGN U14857 ( .B(clk), .A(\g.we_clk [1533]));
Q_ASSIGN U14858 ( .B(clk), .A(\g.we_clk [1532]));
Q_ASSIGN U14859 ( .B(clk), .A(\g.we_clk [1531]));
Q_ASSIGN U14860 ( .B(clk), .A(\g.we_clk [1530]));
Q_ASSIGN U14861 ( .B(clk), .A(\g.we_clk [1529]));
Q_ASSIGN U14862 ( .B(clk), .A(\g.we_clk [1528]));
Q_ASSIGN U14863 ( .B(clk), .A(\g.we_clk [1527]));
Q_ASSIGN U14864 ( .B(clk), .A(\g.we_clk [1526]));
Q_ASSIGN U14865 ( .B(clk), .A(\g.we_clk [1525]));
Q_ASSIGN U14866 ( .B(clk), .A(\g.we_clk [1524]));
Q_ASSIGN U14867 ( .B(clk), .A(\g.we_clk [1523]));
Q_ASSIGN U14868 ( .B(clk), .A(\g.we_clk [1522]));
Q_ASSIGN U14869 ( .B(clk), .A(\g.we_clk [1521]));
Q_ASSIGN U14870 ( .B(clk), .A(\g.we_clk [1520]));
Q_ASSIGN U14871 ( .B(clk), .A(\g.we_clk [1519]));
Q_ASSIGN U14872 ( .B(clk), .A(\g.we_clk [1518]));
Q_ASSIGN U14873 ( .B(clk), .A(\g.we_clk [1517]));
Q_ASSIGN U14874 ( .B(clk), .A(\g.we_clk [1516]));
Q_ASSIGN U14875 ( .B(clk), .A(\g.we_clk [1515]));
Q_ASSIGN U14876 ( .B(clk), .A(\g.we_clk [1514]));
Q_ASSIGN U14877 ( .B(clk), .A(\g.we_clk [1513]));
Q_ASSIGN U14878 ( .B(clk), .A(\g.we_clk [1512]));
Q_ASSIGN U14879 ( .B(clk), .A(\g.we_clk [1511]));
Q_ASSIGN U14880 ( .B(clk), .A(\g.we_clk [1510]));
Q_ASSIGN U14881 ( .B(clk), .A(\g.we_clk [1509]));
Q_ASSIGN U14882 ( .B(clk), .A(\g.we_clk [1508]));
Q_ASSIGN U14883 ( .B(clk), .A(\g.we_clk [1507]));
Q_ASSIGN U14884 ( .B(clk), .A(\g.we_clk [1506]));
Q_ASSIGN U14885 ( .B(clk), .A(\g.we_clk [1505]));
Q_ASSIGN U14886 ( .B(clk), .A(\g.we_clk [1504]));
Q_ASSIGN U14887 ( .B(clk), .A(\g.we_clk [1503]));
Q_ASSIGN U14888 ( .B(clk), .A(\g.we_clk [1502]));
Q_ASSIGN U14889 ( .B(clk), .A(\g.we_clk [1501]));
Q_ASSIGN U14890 ( .B(clk), .A(\g.we_clk [1500]));
Q_ASSIGN U14891 ( .B(clk), .A(\g.we_clk [1499]));
Q_ASSIGN U14892 ( .B(clk), .A(\g.we_clk [1498]));
Q_ASSIGN U14893 ( .B(clk), .A(\g.we_clk [1497]));
Q_ASSIGN U14894 ( .B(clk), .A(\g.we_clk [1496]));
Q_ASSIGN U14895 ( .B(clk), .A(\g.we_clk [1495]));
Q_ASSIGN U14896 ( .B(clk), .A(\g.we_clk [1494]));
Q_ASSIGN U14897 ( .B(clk), .A(\g.we_clk [1493]));
Q_ASSIGN U14898 ( .B(clk), .A(\g.we_clk [1492]));
Q_ASSIGN U14899 ( .B(clk), .A(\g.we_clk [1491]));
Q_ASSIGN U14900 ( .B(clk), .A(\g.we_clk [1490]));
Q_ASSIGN U14901 ( .B(clk), .A(\g.we_clk [1489]));
Q_ASSIGN U14902 ( .B(clk), .A(\g.we_clk [1488]));
Q_ASSIGN U14903 ( .B(clk), .A(\g.we_clk [1487]));
Q_ASSIGN U14904 ( .B(clk), .A(\g.we_clk [1486]));
Q_ASSIGN U14905 ( .B(clk), .A(\g.we_clk [1485]));
Q_ASSIGN U14906 ( .B(clk), .A(\g.we_clk [1484]));
Q_ASSIGN U14907 ( .B(clk), .A(\g.we_clk [1483]));
Q_ASSIGN U14908 ( .B(clk), .A(\g.we_clk [1482]));
Q_ASSIGN U14909 ( .B(clk), .A(\g.we_clk [1481]));
Q_ASSIGN U14910 ( .B(clk), .A(\g.we_clk [1480]));
Q_ASSIGN U14911 ( .B(clk), .A(\g.we_clk [1479]));
Q_ASSIGN U14912 ( .B(clk), .A(\g.we_clk [1478]));
Q_ASSIGN U14913 ( .B(clk), .A(\g.we_clk [1477]));
Q_ASSIGN U14914 ( .B(clk), .A(\g.we_clk [1476]));
Q_ASSIGN U14915 ( .B(clk), .A(\g.we_clk [1475]));
Q_ASSIGN U14916 ( .B(clk), .A(\g.we_clk [1474]));
Q_ASSIGN U14917 ( .B(clk), .A(\g.we_clk [1473]));
Q_ASSIGN U14918 ( .B(clk), .A(\g.we_clk [1472]));
Q_ASSIGN U14919 ( .B(clk), .A(\g.we_clk [1471]));
Q_ASSIGN U14920 ( .B(clk), .A(\g.we_clk [1470]));
Q_ASSIGN U14921 ( .B(clk), .A(\g.we_clk [1469]));
Q_ASSIGN U14922 ( .B(clk), .A(\g.we_clk [1468]));
Q_ASSIGN U14923 ( .B(clk), .A(\g.we_clk [1467]));
Q_ASSIGN U14924 ( .B(clk), .A(\g.we_clk [1466]));
Q_ASSIGN U14925 ( .B(clk), .A(\g.we_clk [1465]));
Q_ASSIGN U14926 ( .B(clk), .A(\g.we_clk [1464]));
Q_ASSIGN U14927 ( .B(clk), .A(\g.we_clk [1463]));
Q_ASSIGN U14928 ( .B(clk), .A(\g.we_clk [1462]));
Q_ASSIGN U14929 ( .B(clk), .A(\g.we_clk [1461]));
Q_ASSIGN U14930 ( .B(clk), .A(\g.we_clk [1460]));
Q_ASSIGN U14931 ( .B(clk), .A(\g.we_clk [1459]));
Q_ASSIGN U14932 ( .B(clk), .A(\g.we_clk [1458]));
Q_ASSIGN U14933 ( .B(clk), .A(\g.we_clk [1457]));
Q_ASSIGN U14934 ( .B(clk), .A(\g.we_clk [1456]));
Q_ASSIGN U14935 ( .B(clk), .A(\g.we_clk [1455]));
Q_ASSIGN U14936 ( .B(clk), .A(\g.we_clk [1454]));
Q_ASSIGN U14937 ( .B(clk), .A(\g.we_clk [1453]));
Q_ASSIGN U14938 ( .B(clk), .A(\g.we_clk [1452]));
Q_ASSIGN U14939 ( .B(clk), .A(\g.we_clk [1451]));
Q_ASSIGN U14940 ( .B(clk), .A(\g.we_clk [1450]));
Q_ASSIGN U14941 ( .B(clk), .A(\g.we_clk [1449]));
Q_ASSIGN U14942 ( .B(clk), .A(\g.we_clk [1448]));
Q_ASSIGN U14943 ( .B(clk), .A(\g.we_clk [1447]));
Q_ASSIGN U14944 ( .B(clk), .A(\g.we_clk [1446]));
Q_ASSIGN U14945 ( .B(clk), .A(\g.we_clk [1445]));
Q_ASSIGN U14946 ( .B(clk), .A(\g.we_clk [1444]));
Q_ASSIGN U14947 ( .B(clk), .A(\g.we_clk [1443]));
Q_ASSIGN U14948 ( .B(clk), .A(\g.we_clk [1442]));
Q_ASSIGN U14949 ( .B(clk), .A(\g.we_clk [1441]));
Q_ASSIGN U14950 ( .B(clk), .A(\g.we_clk [1440]));
Q_ASSIGN U14951 ( .B(clk), .A(\g.we_clk [1439]));
Q_ASSIGN U14952 ( .B(clk), .A(\g.we_clk [1438]));
Q_ASSIGN U14953 ( .B(clk), .A(\g.we_clk [1437]));
Q_ASSIGN U14954 ( .B(clk), .A(\g.we_clk [1436]));
Q_ASSIGN U14955 ( .B(clk), .A(\g.we_clk [1435]));
Q_ASSIGN U14956 ( .B(clk), .A(\g.we_clk [1434]));
Q_ASSIGN U14957 ( .B(clk), .A(\g.we_clk [1433]));
Q_ASSIGN U14958 ( .B(clk), .A(\g.we_clk [1432]));
Q_ASSIGN U14959 ( .B(clk), .A(\g.we_clk [1431]));
Q_ASSIGN U14960 ( .B(clk), .A(\g.we_clk [1430]));
Q_ASSIGN U14961 ( .B(clk), .A(\g.we_clk [1429]));
Q_ASSIGN U14962 ( .B(clk), .A(\g.we_clk [1428]));
Q_ASSIGN U14963 ( .B(clk), .A(\g.we_clk [1427]));
Q_ASSIGN U14964 ( .B(clk), .A(\g.we_clk [1426]));
Q_ASSIGN U14965 ( .B(clk), .A(\g.we_clk [1425]));
Q_ASSIGN U14966 ( .B(clk), .A(\g.we_clk [1424]));
Q_ASSIGN U14967 ( .B(clk), .A(\g.we_clk [1423]));
Q_ASSIGN U14968 ( .B(clk), .A(\g.we_clk [1422]));
Q_ASSIGN U14969 ( .B(clk), .A(\g.we_clk [1421]));
Q_ASSIGN U14970 ( .B(clk), .A(\g.we_clk [1420]));
Q_ASSIGN U14971 ( .B(clk), .A(\g.we_clk [1419]));
Q_ASSIGN U14972 ( .B(clk), .A(\g.we_clk [1418]));
Q_ASSIGN U14973 ( .B(clk), .A(\g.we_clk [1417]));
Q_ASSIGN U14974 ( .B(clk), .A(\g.we_clk [1416]));
Q_ASSIGN U14975 ( .B(clk), .A(\g.we_clk [1415]));
Q_ASSIGN U14976 ( .B(clk), .A(\g.we_clk [1414]));
Q_ASSIGN U14977 ( .B(clk), .A(\g.we_clk [1413]));
Q_ASSIGN U14978 ( .B(clk), .A(\g.we_clk [1412]));
Q_ASSIGN U14979 ( .B(clk), .A(\g.we_clk [1411]));
Q_ASSIGN U14980 ( .B(clk), .A(\g.we_clk [1410]));
Q_ASSIGN U14981 ( .B(clk), .A(\g.we_clk [1409]));
Q_ASSIGN U14982 ( .B(clk), .A(\g.we_clk [1408]));
Q_ASSIGN U14983 ( .B(clk), .A(\g.we_clk [1407]));
Q_ASSIGN U14984 ( .B(clk), .A(\g.we_clk [1406]));
Q_ASSIGN U14985 ( .B(clk), .A(\g.we_clk [1405]));
Q_ASSIGN U14986 ( .B(clk), .A(\g.we_clk [1404]));
Q_ASSIGN U14987 ( .B(clk), .A(\g.we_clk [1403]));
Q_ASSIGN U14988 ( .B(clk), .A(\g.we_clk [1402]));
Q_ASSIGN U14989 ( .B(clk), .A(\g.we_clk [1401]));
Q_ASSIGN U14990 ( .B(clk), .A(\g.we_clk [1400]));
Q_ASSIGN U14991 ( .B(clk), .A(\g.we_clk [1399]));
Q_ASSIGN U14992 ( .B(clk), .A(\g.we_clk [1398]));
Q_ASSIGN U14993 ( .B(clk), .A(\g.we_clk [1397]));
Q_ASSIGN U14994 ( .B(clk), .A(\g.we_clk [1396]));
Q_ASSIGN U14995 ( .B(clk), .A(\g.we_clk [1395]));
Q_ASSIGN U14996 ( .B(clk), .A(\g.we_clk [1394]));
Q_ASSIGN U14997 ( .B(clk), .A(\g.we_clk [1393]));
Q_ASSIGN U14998 ( .B(clk), .A(\g.we_clk [1392]));
Q_ASSIGN U14999 ( .B(clk), .A(\g.we_clk [1391]));
Q_ASSIGN U15000 ( .B(clk), .A(\g.we_clk [1390]));
Q_ASSIGN U15001 ( .B(clk), .A(\g.we_clk [1389]));
Q_ASSIGN U15002 ( .B(clk), .A(\g.we_clk [1388]));
Q_ASSIGN U15003 ( .B(clk), .A(\g.we_clk [1387]));
Q_ASSIGN U15004 ( .B(clk), .A(\g.we_clk [1386]));
Q_ASSIGN U15005 ( .B(clk), .A(\g.we_clk [1385]));
Q_ASSIGN U15006 ( .B(clk), .A(\g.we_clk [1384]));
Q_ASSIGN U15007 ( .B(clk), .A(\g.we_clk [1383]));
Q_ASSIGN U15008 ( .B(clk), .A(\g.we_clk [1382]));
Q_ASSIGN U15009 ( .B(clk), .A(\g.we_clk [1381]));
Q_ASSIGN U15010 ( .B(clk), .A(\g.we_clk [1380]));
Q_ASSIGN U15011 ( .B(clk), .A(\g.we_clk [1379]));
Q_ASSIGN U15012 ( .B(clk), .A(\g.we_clk [1378]));
Q_ASSIGN U15013 ( .B(clk), .A(\g.we_clk [1377]));
Q_ASSIGN U15014 ( .B(clk), .A(\g.we_clk [1376]));
Q_ASSIGN U15015 ( .B(clk), .A(\g.we_clk [1375]));
Q_ASSIGN U15016 ( .B(clk), .A(\g.we_clk [1374]));
Q_ASSIGN U15017 ( .B(clk), .A(\g.we_clk [1373]));
Q_ASSIGN U15018 ( .B(clk), .A(\g.we_clk [1372]));
Q_ASSIGN U15019 ( .B(clk), .A(\g.we_clk [1371]));
Q_ASSIGN U15020 ( .B(clk), .A(\g.we_clk [1370]));
Q_ASSIGN U15021 ( .B(clk), .A(\g.we_clk [1369]));
Q_ASSIGN U15022 ( .B(clk), .A(\g.we_clk [1368]));
Q_ASSIGN U15023 ( .B(clk), .A(\g.we_clk [1367]));
Q_ASSIGN U15024 ( .B(clk), .A(\g.we_clk [1366]));
Q_ASSIGN U15025 ( .B(clk), .A(\g.we_clk [1365]));
Q_ASSIGN U15026 ( .B(clk), .A(\g.we_clk [1364]));
Q_ASSIGN U15027 ( .B(clk), .A(\g.we_clk [1363]));
Q_ASSIGN U15028 ( .B(clk), .A(\g.we_clk [1362]));
Q_ASSIGN U15029 ( .B(clk), .A(\g.we_clk [1361]));
Q_ASSIGN U15030 ( .B(clk), .A(\g.we_clk [1360]));
Q_ASSIGN U15031 ( .B(clk), .A(\g.we_clk [1359]));
Q_ASSIGN U15032 ( .B(clk), .A(\g.we_clk [1358]));
Q_ASSIGN U15033 ( .B(clk), .A(\g.we_clk [1357]));
Q_ASSIGN U15034 ( .B(clk), .A(\g.we_clk [1356]));
Q_ASSIGN U15035 ( .B(clk), .A(\g.we_clk [1355]));
Q_ASSIGN U15036 ( .B(clk), .A(\g.we_clk [1354]));
Q_ASSIGN U15037 ( .B(clk), .A(\g.we_clk [1353]));
Q_ASSIGN U15038 ( .B(clk), .A(\g.we_clk [1352]));
Q_ASSIGN U15039 ( .B(clk), .A(\g.we_clk [1351]));
Q_ASSIGN U15040 ( .B(clk), .A(\g.we_clk [1350]));
Q_ASSIGN U15041 ( .B(clk), .A(\g.we_clk [1349]));
Q_ASSIGN U15042 ( .B(clk), .A(\g.we_clk [1348]));
Q_ASSIGN U15043 ( .B(clk), .A(\g.we_clk [1347]));
Q_ASSIGN U15044 ( .B(clk), .A(\g.we_clk [1346]));
Q_ASSIGN U15045 ( .B(clk), .A(\g.we_clk [1345]));
Q_ASSIGN U15046 ( .B(clk), .A(\g.we_clk [1344]));
Q_ASSIGN U15047 ( .B(clk), .A(\g.we_clk [1343]));
Q_ASSIGN U15048 ( .B(clk), .A(\g.we_clk [1342]));
Q_ASSIGN U15049 ( .B(clk), .A(\g.we_clk [1341]));
Q_ASSIGN U15050 ( .B(clk), .A(\g.we_clk [1340]));
Q_ASSIGN U15051 ( .B(clk), .A(\g.we_clk [1339]));
Q_ASSIGN U15052 ( .B(clk), .A(\g.we_clk [1338]));
Q_ASSIGN U15053 ( .B(clk), .A(\g.we_clk [1337]));
Q_ASSIGN U15054 ( .B(clk), .A(\g.we_clk [1336]));
Q_ASSIGN U15055 ( .B(clk), .A(\g.we_clk [1335]));
Q_ASSIGN U15056 ( .B(clk), .A(\g.we_clk [1334]));
Q_ASSIGN U15057 ( .B(clk), .A(\g.we_clk [1333]));
Q_ASSIGN U15058 ( .B(clk), .A(\g.we_clk [1332]));
Q_ASSIGN U15059 ( .B(clk), .A(\g.we_clk [1331]));
Q_ASSIGN U15060 ( .B(clk), .A(\g.we_clk [1330]));
Q_ASSIGN U15061 ( .B(clk), .A(\g.we_clk [1329]));
Q_ASSIGN U15062 ( .B(clk), .A(\g.we_clk [1328]));
Q_ASSIGN U15063 ( .B(clk), .A(\g.we_clk [1327]));
Q_ASSIGN U15064 ( .B(clk), .A(\g.we_clk [1326]));
Q_ASSIGN U15065 ( .B(clk), .A(\g.we_clk [1325]));
Q_ASSIGN U15066 ( .B(clk), .A(\g.we_clk [1324]));
Q_ASSIGN U15067 ( .B(clk), .A(\g.we_clk [1323]));
Q_ASSIGN U15068 ( .B(clk), .A(\g.we_clk [1322]));
Q_ASSIGN U15069 ( .B(clk), .A(\g.we_clk [1321]));
Q_ASSIGN U15070 ( .B(clk), .A(\g.we_clk [1320]));
Q_ASSIGN U15071 ( .B(clk), .A(\g.we_clk [1319]));
Q_ASSIGN U15072 ( .B(clk), .A(\g.we_clk [1318]));
Q_ASSIGN U15073 ( .B(clk), .A(\g.we_clk [1317]));
Q_ASSIGN U15074 ( .B(clk), .A(\g.we_clk [1316]));
Q_ASSIGN U15075 ( .B(clk), .A(\g.we_clk [1315]));
Q_ASSIGN U15076 ( .B(clk), .A(\g.we_clk [1314]));
Q_ASSIGN U15077 ( .B(clk), .A(\g.we_clk [1313]));
Q_ASSIGN U15078 ( .B(clk), .A(\g.we_clk [1312]));
Q_ASSIGN U15079 ( .B(clk), .A(\g.we_clk [1311]));
Q_ASSIGN U15080 ( .B(clk), .A(\g.we_clk [1310]));
Q_ASSIGN U15081 ( .B(clk), .A(\g.we_clk [1309]));
Q_ASSIGN U15082 ( .B(clk), .A(\g.we_clk [1308]));
Q_ASSIGN U15083 ( .B(clk), .A(\g.we_clk [1307]));
Q_ASSIGN U15084 ( .B(clk), .A(\g.we_clk [1306]));
Q_ASSIGN U15085 ( .B(clk), .A(\g.we_clk [1305]));
Q_ASSIGN U15086 ( .B(clk), .A(\g.we_clk [1304]));
Q_ASSIGN U15087 ( .B(clk), .A(\g.we_clk [1303]));
Q_ASSIGN U15088 ( .B(clk), .A(\g.we_clk [1302]));
Q_ASSIGN U15089 ( .B(clk), .A(\g.we_clk [1301]));
Q_ASSIGN U15090 ( .B(clk), .A(\g.we_clk [1300]));
Q_ASSIGN U15091 ( .B(clk), .A(\g.we_clk [1299]));
Q_ASSIGN U15092 ( .B(clk), .A(\g.we_clk [1298]));
Q_ASSIGN U15093 ( .B(clk), .A(\g.we_clk [1297]));
Q_ASSIGN U15094 ( .B(clk), .A(\g.we_clk [1296]));
Q_ASSIGN U15095 ( .B(clk), .A(\g.we_clk [1295]));
Q_ASSIGN U15096 ( .B(clk), .A(\g.we_clk [1294]));
Q_ASSIGN U15097 ( .B(clk), .A(\g.we_clk [1293]));
Q_ASSIGN U15098 ( .B(clk), .A(\g.we_clk [1292]));
Q_ASSIGN U15099 ( .B(clk), .A(\g.we_clk [1291]));
Q_ASSIGN U15100 ( .B(clk), .A(\g.we_clk [1290]));
Q_ASSIGN U15101 ( .B(clk), .A(\g.we_clk [1289]));
Q_ASSIGN U15102 ( .B(clk), .A(\g.we_clk [1288]));
Q_ASSIGN U15103 ( .B(clk), .A(\g.we_clk [1287]));
Q_ASSIGN U15104 ( .B(clk), .A(\g.we_clk [1286]));
Q_ASSIGN U15105 ( .B(clk), .A(\g.we_clk [1285]));
Q_ASSIGN U15106 ( .B(clk), .A(\g.we_clk [1284]));
Q_ASSIGN U15107 ( .B(clk), .A(\g.we_clk [1283]));
Q_ASSIGN U15108 ( .B(clk), .A(\g.we_clk [1282]));
Q_ASSIGN U15109 ( .B(clk), .A(\g.we_clk [1281]));
Q_ASSIGN U15110 ( .B(clk), .A(\g.we_clk [1280]));
Q_ASSIGN U15111 ( .B(clk), .A(\g.we_clk [1279]));
Q_ASSIGN U15112 ( .B(clk), .A(\g.we_clk [1278]));
Q_ASSIGN U15113 ( .B(clk), .A(\g.we_clk [1277]));
Q_ASSIGN U15114 ( .B(clk), .A(\g.we_clk [1276]));
Q_ASSIGN U15115 ( .B(clk), .A(\g.we_clk [1275]));
Q_ASSIGN U15116 ( .B(clk), .A(\g.we_clk [1274]));
Q_ASSIGN U15117 ( .B(clk), .A(\g.we_clk [1273]));
Q_ASSIGN U15118 ( .B(clk), .A(\g.we_clk [1272]));
Q_ASSIGN U15119 ( .B(clk), .A(\g.we_clk [1271]));
Q_ASSIGN U15120 ( .B(clk), .A(\g.we_clk [1270]));
Q_ASSIGN U15121 ( .B(clk), .A(\g.we_clk [1269]));
Q_ASSIGN U15122 ( .B(clk), .A(\g.we_clk [1268]));
Q_ASSIGN U15123 ( .B(clk), .A(\g.we_clk [1267]));
Q_ASSIGN U15124 ( .B(clk), .A(\g.we_clk [1266]));
Q_ASSIGN U15125 ( .B(clk), .A(\g.we_clk [1265]));
Q_ASSIGN U15126 ( .B(clk), .A(\g.we_clk [1264]));
Q_ASSIGN U15127 ( .B(clk), .A(\g.we_clk [1263]));
Q_ASSIGN U15128 ( .B(clk), .A(\g.we_clk [1262]));
Q_ASSIGN U15129 ( .B(clk), .A(\g.we_clk [1261]));
Q_ASSIGN U15130 ( .B(clk), .A(\g.we_clk [1260]));
Q_ASSIGN U15131 ( .B(clk), .A(\g.we_clk [1259]));
Q_ASSIGN U15132 ( .B(clk), .A(\g.we_clk [1258]));
Q_ASSIGN U15133 ( .B(clk), .A(\g.we_clk [1257]));
Q_ASSIGN U15134 ( .B(clk), .A(\g.we_clk [1256]));
Q_ASSIGN U15135 ( .B(clk), .A(\g.we_clk [1255]));
Q_ASSIGN U15136 ( .B(clk), .A(\g.we_clk [1254]));
Q_ASSIGN U15137 ( .B(clk), .A(\g.we_clk [1253]));
Q_ASSIGN U15138 ( .B(clk), .A(\g.we_clk [1252]));
Q_ASSIGN U15139 ( .B(clk), .A(\g.we_clk [1251]));
Q_ASSIGN U15140 ( .B(clk), .A(\g.we_clk [1250]));
Q_ASSIGN U15141 ( .B(clk), .A(\g.we_clk [1249]));
Q_ASSIGN U15142 ( .B(clk), .A(\g.we_clk [1248]));
Q_ASSIGN U15143 ( .B(clk), .A(\g.we_clk [1247]));
Q_ASSIGN U15144 ( .B(clk), .A(\g.we_clk [1246]));
Q_ASSIGN U15145 ( .B(clk), .A(\g.we_clk [1245]));
Q_ASSIGN U15146 ( .B(clk), .A(\g.we_clk [1244]));
Q_ASSIGN U15147 ( .B(clk), .A(\g.we_clk [1243]));
Q_ASSIGN U15148 ( .B(clk), .A(\g.we_clk [1242]));
Q_ASSIGN U15149 ( .B(clk), .A(\g.we_clk [1241]));
Q_ASSIGN U15150 ( .B(clk), .A(\g.we_clk [1240]));
Q_ASSIGN U15151 ( .B(clk), .A(\g.we_clk [1239]));
Q_ASSIGN U15152 ( .B(clk), .A(\g.we_clk [1238]));
Q_ASSIGN U15153 ( .B(clk), .A(\g.we_clk [1237]));
Q_ASSIGN U15154 ( .B(clk), .A(\g.we_clk [1236]));
Q_ASSIGN U15155 ( .B(clk), .A(\g.we_clk [1235]));
Q_ASSIGN U15156 ( .B(clk), .A(\g.we_clk [1234]));
Q_ASSIGN U15157 ( .B(clk), .A(\g.we_clk [1233]));
Q_ASSIGN U15158 ( .B(clk), .A(\g.we_clk [1232]));
Q_ASSIGN U15159 ( .B(clk), .A(\g.we_clk [1231]));
Q_ASSIGN U15160 ( .B(clk), .A(\g.we_clk [1230]));
Q_ASSIGN U15161 ( .B(clk), .A(\g.we_clk [1229]));
Q_ASSIGN U15162 ( .B(clk), .A(\g.we_clk [1228]));
Q_ASSIGN U15163 ( .B(clk), .A(\g.we_clk [1227]));
Q_ASSIGN U15164 ( .B(clk), .A(\g.we_clk [1226]));
Q_ASSIGN U15165 ( .B(clk), .A(\g.we_clk [1225]));
Q_ASSIGN U15166 ( .B(clk), .A(\g.we_clk [1224]));
Q_ASSIGN U15167 ( .B(clk), .A(\g.we_clk [1223]));
Q_ASSIGN U15168 ( .B(clk), .A(\g.we_clk [1222]));
Q_ASSIGN U15169 ( .B(clk), .A(\g.we_clk [1221]));
Q_ASSIGN U15170 ( .B(clk), .A(\g.we_clk [1220]));
Q_ASSIGN U15171 ( .B(clk), .A(\g.we_clk [1219]));
Q_ASSIGN U15172 ( .B(clk), .A(\g.we_clk [1218]));
Q_ASSIGN U15173 ( .B(clk), .A(\g.we_clk [1217]));
Q_ASSIGN U15174 ( .B(clk), .A(\g.we_clk [1216]));
Q_ASSIGN U15175 ( .B(clk), .A(\g.we_clk [1215]));
Q_ASSIGN U15176 ( .B(clk), .A(\g.we_clk [1214]));
Q_ASSIGN U15177 ( .B(clk), .A(\g.we_clk [1213]));
Q_ASSIGN U15178 ( .B(clk), .A(\g.we_clk [1212]));
Q_ASSIGN U15179 ( .B(clk), .A(\g.we_clk [1211]));
Q_ASSIGN U15180 ( .B(clk), .A(\g.we_clk [1210]));
Q_ASSIGN U15181 ( .B(clk), .A(\g.we_clk [1209]));
Q_ASSIGN U15182 ( .B(clk), .A(\g.we_clk [1208]));
Q_ASSIGN U15183 ( .B(clk), .A(\g.we_clk [1207]));
Q_ASSIGN U15184 ( .B(clk), .A(\g.we_clk [1206]));
Q_ASSIGN U15185 ( .B(clk), .A(\g.we_clk [1205]));
Q_ASSIGN U15186 ( .B(clk), .A(\g.we_clk [1204]));
Q_ASSIGN U15187 ( .B(clk), .A(\g.we_clk [1203]));
Q_ASSIGN U15188 ( .B(clk), .A(\g.we_clk [1202]));
Q_ASSIGN U15189 ( .B(clk), .A(\g.we_clk [1201]));
Q_ASSIGN U15190 ( .B(clk), .A(\g.we_clk [1200]));
Q_ASSIGN U15191 ( .B(clk), .A(\g.we_clk [1199]));
Q_ASSIGN U15192 ( .B(clk), .A(\g.we_clk [1198]));
Q_ASSIGN U15193 ( .B(clk), .A(\g.we_clk [1197]));
Q_ASSIGN U15194 ( .B(clk), .A(\g.we_clk [1196]));
Q_ASSIGN U15195 ( .B(clk), .A(\g.we_clk [1195]));
Q_ASSIGN U15196 ( .B(clk), .A(\g.we_clk [1194]));
Q_ASSIGN U15197 ( .B(clk), .A(\g.we_clk [1193]));
Q_ASSIGN U15198 ( .B(clk), .A(\g.we_clk [1192]));
Q_ASSIGN U15199 ( .B(clk), .A(\g.we_clk [1191]));
Q_ASSIGN U15200 ( .B(clk), .A(\g.we_clk [1190]));
Q_ASSIGN U15201 ( .B(clk), .A(\g.we_clk [1189]));
Q_ASSIGN U15202 ( .B(clk), .A(\g.we_clk [1188]));
Q_ASSIGN U15203 ( .B(clk), .A(\g.we_clk [1187]));
Q_ASSIGN U15204 ( .B(clk), .A(\g.we_clk [1186]));
Q_ASSIGN U15205 ( .B(clk), .A(\g.we_clk [1185]));
Q_ASSIGN U15206 ( .B(clk), .A(\g.we_clk [1184]));
Q_ASSIGN U15207 ( .B(clk), .A(\g.we_clk [1183]));
Q_ASSIGN U15208 ( .B(clk), .A(\g.we_clk [1182]));
Q_ASSIGN U15209 ( .B(clk), .A(\g.we_clk [1181]));
Q_ASSIGN U15210 ( .B(clk), .A(\g.we_clk [1180]));
Q_ASSIGN U15211 ( .B(clk), .A(\g.we_clk [1179]));
Q_ASSIGN U15212 ( .B(clk), .A(\g.we_clk [1178]));
Q_ASSIGN U15213 ( .B(clk), .A(\g.we_clk [1177]));
Q_ASSIGN U15214 ( .B(clk), .A(\g.we_clk [1176]));
Q_ASSIGN U15215 ( .B(clk), .A(\g.we_clk [1175]));
Q_ASSIGN U15216 ( .B(clk), .A(\g.we_clk [1174]));
Q_ASSIGN U15217 ( .B(clk), .A(\g.we_clk [1173]));
Q_ASSIGN U15218 ( .B(clk), .A(\g.we_clk [1172]));
Q_ASSIGN U15219 ( .B(clk), .A(\g.we_clk [1171]));
Q_ASSIGN U15220 ( .B(clk), .A(\g.we_clk [1170]));
Q_ASSIGN U15221 ( .B(clk), .A(\g.we_clk [1169]));
Q_ASSIGN U15222 ( .B(clk), .A(\g.we_clk [1168]));
Q_ASSIGN U15223 ( .B(clk), .A(\g.we_clk [1167]));
Q_ASSIGN U15224 ( .B(clk), .A(\g.we_clk [1166]));
Q_ASSIGN U15225 ( .B(clk), .A(\g.we_clk [1165]));
Q_ASSIGN U15226 ( .B(clk), .A(\g.we_clk [1164]));
Q_ASSIGN U15227 ( .B(clk), .A(\g.we_clk [1163]));
Q_ASSIGN U15228 ( .B(clk), .A(\g.we_clk [1162]));
Q_ASSIGN U15229 ( .B(clk), .A(\g.we_clk [1161]));
Q_ASSIGN U15230 ( .B(clk), .A(\g.we_clk [1160]));
Q_ASSIGN U15231 ( .B(clk), .A(\g.we_clk [1159]));
Q_ASSIGN U15232 ( .B(clk), .A(\g.we_clk [1158]));
Q_ASSIGN U15233 ( .B(clk), .A(\g.we_clk [1157]));
Q_ASSIGN U15234 ( .B(clk), .A(\g.we_clk [1156]));
Q_ASSIGN U15235 ( .B(clk), .A(\g.we_clk [1155]));
Q_ASSIGN U15236 ( .B(clk), .A(\g.we_clk [1154]));
Q_ASSIGN U15237 ( .B(clk), .A(\g.we_clk [1153]));
Q_ASSIGN U15238 ( .B(clk), .A(\g.we_clk [1152]));
Q_ASSIGN U15239 ( .B(clk), .A(\g.we_clk [1151]));
Q_ASSIGN U15240 ( .B(clk), .A(\g.we_clk [1150]));
Q_ASSIGN U15241 ( .B(clk), .A(\g.we_clk [1149]));
Q_ASSIGN U15242 ( .B(clk), .A(\g.we_clk [1148]));
Q_ASSIGN U15243 ( .B(clk), .A(\g.we_clk [1147]));
Q_ASSIGN U15244 ( .B(clk), .A(\g.we_clk [1146]));
Q_ASSIGN U15245 ( .B(clk), .A(\g.we_clk [1145]));
Q_ASSIGN U15246 ( .B(clk), .A(\g.we_clk [1144]));
Q_ASSIGN U15247 ( .B(clk), .A(\g.we_clk [1143]));
Q_ASSIGN U15248 ( .B(clk), .A(\g.we_clk [1142]));
Q_ASSIGN U15249 ( .B(clk), .A(\g.we_clk [1141]));
Q_ASSIGN U15250 ( .B(clk), .A(\g.we_clk [1140]));
Q_ASSIGN U15251 ( .B(clk), .A(\g.we_clk [1139]));
Q_ASSIGN U15252 ( .B(clk), .A(\g.we_clk [1138]));
Q_ASSIGN U15253 ( .B(clk), .A(\g.we_clk [1137]));
Q_ASSIGN U15254 ( .B(clk), .A(\g.we_clk [1136]));
Q_ASSIGN U15255 ( .B(clk), .A(\g.we_clk [1135]));
Q_ASSIGN U15256 ( .B(clk), .A(\g.we_clk [1134]));
Q_ASSIGN U15257 ( .B(clk), .A(\g.we_clk [1133]));
Q_ASSIGN U15258 ( .B(clk), .A(\g.we_clk [1132]));
Q_ASSIGN U15259 ( .B(clk), .A(\g.we_clk [1131]));
Q_ASSIGN U15260 ( .B(clk), .A(\g.we_clk [1130]));
Q_ASSIGN U15261 ( .B(clk), .A(\g.we_clk [1129]));
Q_ASSIGN U15262 ( .B(clk), .A(\g.we_clk [1128]));
Q_ASSIGN U15263 ( .B(clk), .A(\g.we_clk [1127]));
Q_ASSIGN U15264 ( .B(clk), .A(\g.we_clk [1126]));
Q_ASSIGN U15265 ( .B(clk), .A(\g.we_clk [1125]));
Q_ASSIGN U15266 ( .B(clk), .A(\g.we_clk [1124]));
Q_ASSIGN U15267 ( .B(clk), .A(\g.we_clk [1123]));
Q_ASSIGN U15268 ( .B(clk), .A(\g.we_clk [1122]));
Q_ASSIGN U15269 ( .B(clk), .A(\g.we_clk [1121]));
Q_ASSIGN U15270 ( .B(clk), .A(\g.we_clk [1120]));
Q_ASSIGN U15271 ( .B(clk), .A(\g.we_clk [1119]));
Q_ASSIGN U15272 ( .B(clk), .A(\g.we_clk [1118]));
Q_ASSIGN U15273 ( .B(clk), .A(\g.we_clk [1117]));
Q_ASSIGN U15274 ( .B(clk), .A(\g.we_clk [1116]));
Q_ASSIGN U15275 ( .B(clk), .A(\g.we_clk [1115]));
Q_ASSIGN U15276 ( .B(clk), .A(\g.we_clk [1114]));
Q_ASSIGN U15277 ( .B(clk), .A(\g.we_clk [1113]));
Q_ASSIGN U15278 ( .B(clk), .A(\g.we_clk [1112]));
Q_ASSIGN U15279 ( .B(clk), .A(\g.we_clk [1111]));
Q_ASSIGN U15280 ( .B(clk), .A(\g.we_clk [1110]));
Q_ASSIGN U15281 ( .B(clk), .A(\g.we_clk [1109]));
Q_ASSIGN U15282 ( .B(clk), .A(\g.we_clk [1108]));
Q_ASSIGN U15283 ( .B(clk), .A(\g.we_clk [1107]));
Q_ASSIGN U15284 ( .B(clk), .A(\g.we_clk [1106]));
Q_ASSIGN U15285 ( .B(clk), .A(\g.we_clk [1105]));
Q_ASSIGN U15286 ( .B(clk), .A(\g.we_clk [1104]));
Q_ASSIGN U15287 ( .B(clk), .A(\g.we_clk [1103]));
Q_ASSIGN U15288 ( .B(clk), .A(\g.we_clk [1102]));
Q_ASSIGN U15289 ( .B(clk), .A(\g.we_clk [1101]));
Q_ASSIGN U15290 ( .B(clk), .A(\g.we_clk [1100]));
Q_ASSIGN U15291 ( .B(clk), .A(\g.we_clk [1099]));
Q_ASSIGN U15292 ( .B(clk), .A(\g.we_clk [1098]));
Q_ASSIGN U15293 ( .B(clk), .A(\g.we_clk [1097]));
Q_ASSIGN U15294 ( .B(clk), .A(\g.we_clk [1096]));
Q_ASSIGN U15295 ( .B(clk), .A(\g.we_clk [1095]));
Q_ASSIGN U15296 ( .B(clk), .A(\g.we_clk [1094]));
Q_ASSIGN U15297 ( .B(clk), .A(\g.we_clk [1093]));
Q_ASSIGN U15298 ( .B(clk), .A(\g.we_clk [1092]));
Q_ASSIGN U15299 ( .B(clk), .A(\g.we_clk [1091]));
Q_ASSIGN U15300 ( .B(clk), .A(\g.we_clk [1090]));
Q_ASSIGN U15301 ( .B(clk), .A(\g.we_clk [1089]));
Q_ASSIGN U15302 ( .B(clk), .A(\g.we_clk [1088]));
Q_ASSIGN U15303 ( .B(clk), .A(\g.we_clk [1087]));
Q_ASSIGN U15304 ( .B(clk), .A(\g.we_clk [1086]));
Q_ASSIGN U15305 ( .B(clk), .A(\g.we_clk [1085]));
Q_ASSIGN U15306 ( .B(clk), .A(\g.we_clk [1084]));
Q_ASSIGN U15307 ( .B(clk), .A(\g.we_clk [1083]));
Q_ASSIGN U15308 ( .B(clk), .A(\g.we_clk [1082]));
Q_ASSIGN U15309 ( .B(clk), .A(\g.we_clk [1081]));
Q_ASSIGN U15310 ( .B(clk), .A(\g.we_clk [1080]));
Q_ASSIGN U15311 ( .B(clk), .A(\g.we_clk [1079]));
Q_ASSIGN U15312 ( .B(clk), .A(\g.we_clk [1078]));
Q_ASSIGN U15313 ( .B(clk), .A(\g.we_clk [1077]));
Q_ASSIGN U15314 ( .B(clk), .A(\g.we_clk [1076]));
Q_ASSIGN U15315 ( .B(clk), .A(\g.we_clk [1075]));
Q_ASSIGN U15316 ( .B(clk), .A(\g.we_clk [1074]));
Q_ASSIGN U15317 ( .B(clk), .A(\g.we_clk [1073]));
Q_ASSIGN U15318 ( .B(clk), .A(\g.we_clk [1072]));
Q_ASSIGN U15319 ( .B(clk), .A(\g.we_clk [1071]));
Q_ASSIGN U15320 ( .B(clk), .A(\g.we_clk [1070]));
Q_ASSIGN U15321 ( .B(clk), .A(\g.we_clk [1069]));
Q_ASSIGN U15322 ( .B(clk), .A(\g.we_clk [1068]));
Q_ASSIGN U15323 ( .B(clk), .A(\g.we_clk [1067]));
Q_ASSIGN U15324 ( .B(clk), .A(\g.we_clk [1066]));
Q_ASSIGN U15325 ( .B(clk), .A(\g.we_clk [1065]));
Q_ASSIGN U15326 ( .B(clk), .A(\g.we_clk [1064]));
Q_ASSIGN U15327 ( .B(clk), .A(\g.we_clk [1063]));
Q_ASSIGN U15328 ( .B(clk), .A(\g.we_clk [1062]));
Q_ASSIGN U15329 ( .B(clk), .A(\g.we_clk [1061]));
Q_ASSIGN U15330 ( .B(clk), .A(\g.we_clk [1060]));
Q_ASSIGN U15331 ( .B(clk), .A(\g.we_clk [1059]));
Q_ASSIGN U15332 ( .B(clk), .A(\g.we_clk [1058]));
Q_ASSIGN U15333 ( .B(clk), .A(\g.we_clk [1057]));
Q_ASSIGN U15334 ( .B(clk), .A(\g.we_clk [1056]));
Q_ASSIGN U15335 ( .B(clk), .A(\g.we_clk [1055]));
Q_ASSIGN U15336 ( .B(clk), .A(\g.we_clk [1054]));
Q_ASSIGN U15337 ( .B(clk), .A(\g.we_clk [1053]));
Q_ASSIGN U15338 ( .B(clk), .A(\g.we_clk [1052]));
Q_ASSIGN U15339 ( .B(clk), .A(\g.we_clk [1051]));
Q_ASSIGN U15340 ( .B(clk), .A(\g.we_clk [1050]));
Q_ASSIGN U15341 ( .B(clk), .A(\g.we_clk [1049]));
Q_ASSIGN U15342 ( .B(clk), .A(\g.we_clk [1048]));
Q_ASSIGN U15343 ( .B(clk), .A(\g.we_clk [1047]));
Q_ASSIGN U15344 ( .B(clk), .A(\g.we_clk [1046]));
Q_ASSIGN U15345 ( .B(clk), .A(\g.we_clk [1045]));
Q_ASSIGN U15346 ( .B(clk), .A(\g.we_clk [1044]));
Q_ASSIGN U15347 ( .B(clk), .A(\g.we_clk [1043]));
Q_ASSIGN U15348 ( .B(clk), .A(\g.we_clk [1042]));
Q_ASSIGN U15349 ( .B(clk), .A(\g.we_clk [1041]));
Q_ASSIGN U15350 ( .B(clk), .A(\g.we_clk [1040]));
Q_ASSIGN U15351 ( .B(clk), .A(\g.we_clk [1039]));
Q_ASSIGN U15352 ( .B(clk), .A(\g.we_clk [1038]));
Q_ASSIGN U15353 ( .B(clk), .A(\g.we_clk [1037]));
Q_ASSIGN U15354 ( .B(clk), .A(\g.we_clk [1036]));
Q_ASSIGN U15355 ( .B(clk), .A(\g.we_clk [1035]));
Q_ASSIGN U15356 ( .B(clk), .A(\g.we_clk [1034]));
Q_ASSIGN U15357 ( .B(clk), .A(\g.we_clk [1033]));
Q_ASSIGN U15358 ( .B(clk), .A(\g.we_clk [1032]));
Q_ASSIGN U15359 ( .B(clk), .A(\g.we_clk [1031]));
Q_ASSIGN U15360 ( .B(clk), .A(\g.we_clk [1030]));
Q_ASSIGN U15361 ( .B(clk), .A(\g.we_clk [1029]));
Q_ASSIGN U15362 ( .B(clk), .A(\g.we_clk [1028]));
Q_ASSIGN U15363 ( .B(clk), .A(\g.we_clk [1027]));
Q_ASSIGN U15364 ( .B(clk), .A(\g.we_clk [1026]));
Q_ASSIGN U15365 ( .B(clk), .A(\g.we_clk [1025]));
Q_ASSIGN U15366 ( .B(clk), .A(\g.we_clk [1024]));
Q_ASSIGN U15367 ( .B(clk), .A(\g.we_clk [1023]));
Q_ASSIGN U15368 ( .B(clk), .A(\g.we_clk [1022]));
Q_ASSIGN U15369 ( .B(clk), .A(\g.we_clk [1021]));
Q_ASSIGN U15370 ( .B(clk), .A(\g.we_clk [1020]));
Q_ASSIGN U15371 ( .B(clk), .A(\g.we_clk [1019]));
Q_ASSIGN U15372 ( .B(clk), .A(\g.we_clk [1018]));
Q_ASSIGN U15373 ( .B(clk), .A(\g.we_clk [1017]));
Q_ASSIGN U15374 ( .B(clk), .A(\g.we_clk [1016]));
Q_ASSIGN U15375 ( .B(clk), .A(\g.we_clk [1015]));
Q_ASSIGN U15376 ( .B(clk), .A(\g.we_clk [1014]));
Q_ASSIGN U15377 ( .B(clk), .A(\g.we_clk [1013]));
Q_ASSIGN U15378 ( .B(clk), .A(\g.we_clk [1012]));
Q_ASSIGN U15379 ( .B(clk), .A(\g.we_clk [1011]));
Q_ASSIGN U15380 ( .B(clk), .A(\g.we_clk [1010]));
Q_ASSIGN U15381 ( .B(clk), .A(\g.we_clk [1009]));
Q_ASSIGN U15382 ( .B(clk), .A(\g.we_clk [1008]));
Q_ASSIGN U15383 ( .B(clk), .A(\g.we_clk [1007]));
Q_ASSIGN U15384 ( .B(clk), .A(\g.we_clk [1006]));
Q_ASSIGN U15385 ( .B(clk), .A(\g.we_clk [1005]));
Q_ASSIGN U15386 ( .B(clk), .A(\g.we_clk [1004]));
Q_ASSIGN U15387 ( .B(clk), .A(\g.we_clk [1003]));
Q_ASSIGN U15388 ( .B(clk), .A(\g.we_clk [1002]));
Q_ASSIGN U15389 ( .B(clk), .A(\g.we_clk [1001]));
Q_ASSIGN U15390 ( .B(clk), .A(\g.we_clk [1000]));
Q_ASSIGN U15391 ( .B(clk), .A(\g.we_clk [999]));
Q_ASSIGN U15392 ( .B(clk), .A(\g.we_clk [998]));
Q_ASSIGN U15393 ( .B(clk), .A(\g.we_clk [997]));
Q_ASSIGN U15394 ( .B(clk), .A(\g.we_clk [996]));
Q_ASSIGN U15395 ( .B(clk), .A(\g.we_clk [995]));
Q_ASSIGN U15396 ( .B(clk), .A(\g.we_clk [994]));
Q_ASSIGN U15397 ( .B(clk), .A(\g.we_clk [993]));
Q_ASSIGN U15398 ( .B(clk), .A(\g.we_clk [992]));
Q_ASSIGN U15399 ( .B(clk), .A(\g.we_clk [991]));
Q_ASSIGN U15400 ( .B(clk), .A(\g.we_clk [990]));
Q_ASSIGN U15401 ( .B(clk), .A(\g.we_clk [989]));
Q_ASSIGN U15402 ( .B(clk), .A(\g.we_clk [988]));
Q_ASSIGN U15403 ( .B(clk), .A(\g.we_clk [987]));
Q_ASSIGN U15404 ( .B(clk), .A(\g.we_clk [986]));
Q_ASSIGN U15405 ( .B(clk), .A(\g.we_clk [985]));
Q_ASSIGN U15406 ( .B(clk), .A(\g.we_clk [984]));
Q_ASSIGN U15407 ( .B(clk), .A(\g.we_clk [983]));
Q_ASSIGN U15408 ( .B(clk), .A(\g.we_clk [982]));
Q_ASSIGN U15409 ( .B(clk), .A(\g.we_clk [981]));
Q_ASSIGN U15410 ( .B(clk), .A(\g.we_clk [980]));
Q_ASSIGN U15411 ( .B(clk), .A(\g.we_clk [979]));
Q_ASSIGN U15412 ( .B(clk), .A(\g.we_clk [978]));
Q_ASSIGN U15413 ( .B(clk), .A(\g.we_clk [977]));
Q_ASSIGN U15414 ( .B(clk), .A(\g.we_clk [976]));
Q_ASSIGN U15415 ( .B(clk), .A(\g.we_clk [975]));
Q_ASSIGN U15416 ( .B(clk), .A(\g.we_clk [974]));
Q_ASSIGN U15417 ( .B(clk), .A(\g.we_clk [973]));
Q_ASSIGN U15418 ( .B(clk), .A(\g.we_clk [972]));
Q_ASSIGN U15419 ( .B(clk), .A(\g.we_clk [971]));
Q_ASSIGN U15420 ( .B(clk), .A(\g.we_clk [970]));
Q_ASSIGN U15421 ( .B(clk), .A(\g.we_clk [969]));
Q_ASSIGN U15422 ( .B(clk), .A(\g.we_clk [968]));
Q_ASSIGN U15423 ( .B(clk), .A(\g.we_clk [967]));
Q_ASSIGN U15424 ( .B(clk), .A(\g.we_clk [966]));
Q_ASSIGN U15425 ( .B(clk), .A(\g.we_clk [965]));
Q_ASSIGN U15426 ( .B(clk), .A(\g.we_clk [964]));
Q_ASSIGN U15427 ( .B(clk), .A(\g.we_clk [963]));
Q_ASSIGN U15428 ( .B(clk), .A(\g.we_clk [962]));
Q_ASSIGN U15429 ( .B(clk), .A(\g.we_clk [961]));
Q_ASSIGN U15430 ( .B(clk), .A(\g.we_clk [960]));
Q_ASSIGN U15431 ( .B(clk), .A(\g.we_clk [959]));
Q_ASSIGN U15432 ( .B(clk), .A(\g.we_clk [958]));
Q_ASSIGN U15433 ( .B(clk), .A(\g.we_clk [957]));
Q_ASSIGN U15434 ( .B(clk), .A(\g.we_clk [956]));
Q_ASSIGN U15435 ( .B(clk), .A(\g.we_clk [955]));
Q_ASSIGN U15436 ( .B(clk), .A(\g.we_clk [954]));
Q_ASSIGN U15437 ( .B(clk), .A(\g.we_clk [953]));
Q_ASSIGN U15438 ( .B(clk), .A(\g.we_clk [952]));
Q_ASSIGN U15439 ( .B(clk), .A(\g.we_clk [951]));
Q_ASSIGN U15440 ( .B(clk), .A(\g.we_clk [950]));
Q_ASSIGN U15441 ( .B(clk), .A(\g.we_clk [949]));
Q_ASSIGN U15442 ( .B(clk), .A(\g.we_clk [948]));
Q_ASSIGN U15443 ( .B(clk), .A(\g.we_clk [947]));
Q_ASSIGN U15444 ( .B(clk), .A(\g.we_clk [946]));
Q_ASSIGN U15445 ( .B(clk), .A(\g.we_clk [945]));
Q_ASSIGN U15446 ( .B(clk), .A(\g.we_clk [944]));
Q_ASSIGN U15447 ( .B(clk), .A(\g.we_clk [943]));
Q_ASSIGN U15448 ( .B(clk), .A(\g.we_clk [942]));
Q_ASSIGN U15449 ( .B(clk), .A(\g.we_clk [941]));
Q_ASSIGN U15450 ( .B(clk), .A(\g.we_clk [940]));
Q_ASSIGN U15451 ( .B(clk), .A(\g.we_clk [939]));
Q_ASSIGN U15452 ( .B(clk), .A(\g.we_clk [938]));
Q_ASSIGN U15453 ( .B(clk), .A(\g.we_clk [937]));
Q_ASSIGN U15454 ( .B(clk), .A(\g.we_clk [936]));
Q_ASSIGN U15455 ( .B(clk), .A(\g.we_clk [935]));
Q_ASSIGN U15456 ( .B(clk), .A(\g.we_clk [934]));
Q_ASSIGN U15457 ( .B(clk), .A(\g.we_clk [933]));
Q_ASSIGN U15458 ( .B(clk), .A(\g.we_clk [932]));
Q_ASSIGN U15459 ( .B(clk), .A(\g.we_clk [931]));
Q_ASSIGN U15460 ( .B(clk), .A(\g.we_clk [930]));
Q_ASSIGN U15461 ( .B(clk), .A(\g.we_clk [929]));
Q_ASSIGN U15462 ( .B(clk), .A(\g.we_clk [928]));
Q_ASSIGN U15463 ( .B(clk), .A(\g.we_clk [927]));
Q_ASSIGN U15464 ( .B(clk), .A(\g.we_clk [926]));
Q_ASSIGN U15465 ( .B(clk), .A(\g.we_clk [925]));
Q_ASSIGN U15466 ( .B(clk), .A(\g.we_clk [924]));
Q_ASSIGN U15467 ( .B(clk), .A(\g.we_clk [923]));
Q_ASSIGN U15468 ( .B(clk), .A(\g.we_clk [922]));
Q_ASSIGN U15469 ( .B(clk), .A(\g.we_clk [921]));
Q_ASSIGN U15470 ( .B(clk), .A(\g.we_clk [920]));
Q_ASSIGN U15471 ( .B(clk), .A(\g.we_clk [919]));
Q_ASSIGN U15472 ( .B(clk), .A(\g.we_clk [918]));
Q_ASSIGN U15473 ( .B(clk), .A(\g.we_clk [917]));
Q_ASSIGN U15474 ( .B(clk), .A(\g.we_clk [916]));
Q_ASSIGN U15475 ( .B(clk), .A(\g.we_clk [915]));
Q_ASSIGN U15476 ( .B(clk), .A(\g.we_clk [914]));
Q_ASSIGN U15477 ( .B(clk), .A(\g.we_clk [913]));
Q_ASSIGN U15478 ( .B(clk), .A(\g.we_clk [912]));
Q_ASSIGN U15479 ( .B(clk), .A(\g.we_clk [911]));
Q_ASSIGN U15480 ( .B(clk), .A(\g.we_clk [910]));
Q_ASSIGN U15481 ( .B(clk), .A(\g.we_clk [909]));
Q_ASSIGN U15482 ( .B(clk), .A(\g.we_clk [908]));
Q_ASSIGN U15483 ( .B(clk), .A(\g.we_clk [907]));
Q_ASSIGN U15484 ( .B(clk), .A(\g.we_clk [906]));
Q_ASSIGN U15485 ( .B(clk), .A(\g.we_clk [905]));
Q_ASSIGN U15486 ( .B(clk), .A(\g.we_clk [904]));
Q_ASSIGN U15487 ( .B(clk), .A(\g.we_clk [903]));
Q_ASSIGN U15488 ( .B(clk), .A(\g.we_clk [902]));
Q_ASSIGN U15489 ( .B(clk), .A(\g.we_clk [901]));
Q_ASSIGN U15490 ( .B(clk), .A(\g.we_clk [900]));
Q_ASSIGN U15491 ( .B(clk), .A(\g.we_clk [899]));
Q_ASSIGN U15492 ( .B(clk), .A(\g.we_clk [898]));
Q_ASSIGN U15493 ( .B(clk), .A(\g.we_clk [897]));
Q_ASSIGN U15494 ( .B(clk), .A(\g.we_clk [896]));
Q_ASSIGN U15495 ( .B(clk), .A(\g.we_clk [895]));
Q_ASSIGN U15496 ( .B(clk), .A(\g.we_clk [894]));
Q_ASSIGN U15497 ( .B(clk), .A(\g.we_clk [893]));
Q_ASSIGN U15498 ( .B(clk), .A(\g.we_clk [892]));
Q_ASSIGN U15499 ( .B(clk), .A(\g.we_clk [891]));
Q_ASSIGN U15500 ( .B(clk), .A(\g.we_clk [890]));
Q_ASSIGN U15501 ( .B(clk), .A(\g.we_clk [889]));
Q_ASSIGN U15502 ( .B(clk), .A(\g.we_clk [888]));
Q_ASSIGN U15503 ( .B(clk), .A(\g.we_clk [887]));
Q_ASSIGN U15504 ( .B(clk), .A(\g.we_clk [886]));
Q_ASSIGN U15505 ( .B(clk), .A(\g.we_clk [885]));
Q_ASSIGN U15506 ( .B(clk), .A(\g.we_clk [884]));
Q_ASSIGN U15507 ( .B(clk), .A(\g.we_clk [883]));
Q_ASSIGN U15508 ( .B(clk), .A(\g.we_clk [882]));
Q_ASSIGN U15509 ( .B(clk), .A(\g.we_clk [881]));
Q_ASSIGN U15510 ( .B(clk), .A(\g.we_clk [880]));
Q_ASSIGN U15511 ( .B(clk), .A(\g.we_clk [879]));
Q_ASSIGN U15512 ( .B(clk), .A(\g.we_clk [878]));
Q_ASSIGN U15513 ( .B(clk), .A(\g.we_clk [877]));
Q_ASSIGN U15514 ( .B(clk), .A(\g.we_clk [876]));
Q_ASSIGN U15515 ( .B(clk), .A(\g.we_clk [875]));
Q_ASSIGN U15516 ( .B(clk), .A(\g.we_clk [874]));
Q_ASSIGN U15517 ( .B(clk), .A(\g.we_clk [873]));
Q_ASSIGN U15518 ( .B(clk), .A(\g.we_clk [872]));
Q_ASSIGN U15519 ( .B(clk), .A(\g.we_clk [871]));
Q_ASSIGN U15520 ( .B(clk), .A(\g.we_clk [870]));
Q_ASSIGN U15521 ( .B(clk), .A(\g.we_clk [869]));
Q_ASSIGN U15522 ( .B(clk), .A(\g.we_clk [868]));
Q_ASSIGN U15523 ( .B(clk), .A(\g.we_clk [867]));
Q_ASSIGN U15524 ( .B(clk), .A(\g.we_clk [866]));
Q_ASSIGN U15525 ( .B(clk), .A(\g.we_clk [865]));
Q_ASSIGN U15526 ( .B(clk), .A(\g.we_clk [864]));
Q_ASSIGN U15527 ( .B(clk), .A(\g.we_clk [863]));
Q_ASSIGN U15528 ( .B(clk), .A(\g.we_clk [862]));
Q_ASSIGN U15529 ( .B(clk), .A(\g.we_clk [861]));
Q_ASSIGN U15530 ( .B(clk), .A(\g.we_clk [860]));
Q_ASSIGN U15531 ( .B(clk), .A(\g.we_clk [859]));
Q_ASSIGN U15532 ( .B(clk), .A(\g.we_clk [858]));
Q_ASSIGN U15533 ( .B(clk), .A(\g.we_clk [857]));
Q_ASSIGN U15534 ( .B(clk), .A(\g.we_clk [856]));
Q_ASSIGN U15535 ( .B(clk), .A(\g.we_clk [855]));
Q_ASSIGN U15536 ( .B(clk), .A(\g.we_clk [854]));
Q_ASSIGN U15537 ( .B(clk), .A(\g.we_clk [853]));
Q_ASSIGN U15538 ( .B(clk), .A(\g.we_clk [852]));
Q_ASSIGN U15539 ( .B(clk), .A(\g.we_clk [851]));
Q_ASSIGN U15540 ( .B(clk), .A(\g.we_clk [850]));
Q_ASSIGN U15541 ( .B(clk), .A(\g.we_clk [849]));
Q_ASSIGN U15542 ( .B(clk), .A(\g.we_clk [848]));
Q_ASSIGN U15543 ( .B(clk), .A(\g.we_clk [847]));
Q_ASSIGN U15544 ( .B(clk), .A(\g.we_clk [846]));
Q_ASSIGN U15545 ( .B(clk), .A(\g.we_clk [845]));
Q_ASSIGN U15546 ( .B(clk), .A(\g.we_clk [844]));
Q_ASSIGN U15547 ( .B(clk), .A(\g.we_clk [843]));
Q_ASSIGN U15548 ( .B(clk), .A(\g.we_clk [842]));
Q_ASSIGN U15549 ( .B(clk), .A(\g.we_clk [841]));
Q_ASSIGN U15550 ( .B(clk), .A(\g.we_clk [840]));
Q_ASSIGN U15551 ( .B(clk), .A(\g.we_clk [839]));
Q_ASSIGN U15552 ( .B(clk), .A(\g.we_clk [838]));
Q_ASSIGN U15553 ( .B(clk), .A(\g.we_clk [837]));
Q_ASSIGN U15554 ( .B(clk), .A(\g.we_clk [836]));
Q_ASSIGN U15555 ( .B(clk), .A(\g.we_clk [835]));
Q_ASSIGN U15556 ( .B(clk), .A(\g.we_clk [834]));
Q_ASSIGN U15557 ( .B(clk), .A(\g.we_clk [833]));
Q_ASSIGN U15558 ( .B(clk), .A(\g.we_clk [832]));
Q_ASSIGN U15559 ( .B(clk), .A(\g.we_clk [831]));
Q_ASSIGN U15560 ( .B(clk), .A(\g.we_clk [830]));
Q_ASSIGN U15561 ( .B(clk), .A(\g.we_clk [829]));
Q_ASSIGN U15562 ( .B(clk), .A(\g.we_clk [828]));
Q_ASSIGN U15563 ( .B(clk), .A(\g.we_clk [827]));
Q_ASSIGN U15564 ( .B(clk), .A(\g.we_clk [826]));
Q_ASSIGN U15565 ( .B(clk), .A(\g.we_clk [825]));
Q_ASSIGN U15566 ( .B(clk), .A(\g.we_clk [824]));
Q_ASSIGN U15567 ( .B(clk), .A(\g.we_clk [823]));
Q_ASSIGN U15568 ( .B(clk), .A(\g.we_clk [822]));
Q_ASSIGN U15569 ( .B(clk), .A(\g.we_clk [821]));
Q_ASSIGN U15570 ( .B(clk), .A(\g.we_clk [820]));
Q_ASSIGN U15571 ( .B(clk), .A(\g.we_clk [819]));
Q_ASSIGN U15572 ( .B(clk), .A(\g.we_clk [818]));
Q_ASSIGN U15573 ( .B(clk), .A(\g.we_clk [817]));
Q_ASSIGN U15574 ( .B(clk), .A(\g.we_clk [816]));
Q_ASSIGN U15575 ( .B(clk), .A(\g.we_clk [815]));
Q_ASSIGN U15576 ( .B(clk), .A(\g.we_clk [814]));
Q_ASSIGN U15577 ( .B(clk), .A(\g.we_clk [813]));
Q_ASSIGN U15578 ( .B(clk), .A(\g.we_clk [812]));
Q_ASSIGN U15579 ( .B(clk), .A(\g.we_clk [811]));
Q_ASSIGN U15580 ( .B(clk), .A(\g.we_clk [810]));
Q_ASSIGN U15581 ( .B(clk), .A(\g.we_clk [809]));
Q_ASSIGN U15582 ( .B(clk), .A(\g.we_clk [808]));
Q_ASSIGN U15583 ( .B(clk), .A(\g.we_clk [807]));
Q_ASSIGN U15584 ( .B(clk), .A(\g.we_clk [806]));
Q_ASSIGN U15585 ( .B(clk), .A(\g.we_clk [805]));
Q_ASSIGN U15586 ( .B(clk), .A(\g.we_clk [804]));
Q_ASSIGN U15587 ( .B(clk), .A(\g.we_clk [803]));
Q_ASSIGN U15588 ( .B(clk), .A(\g.we_clk [802]));
Q_ASSIGN U15589 ( .B(clk), .A(\g.we_clk [801]));
Q_ASSIGN U15590 ( .B(clk), .A(\g.we_clk [800]));
Q_ASSIGN U15591 ( .B(clk), .A(\g.we_clk [799]));
Q_ASSIGN U15592 ( .B(clk), .A(\g.we_clk [798]));
Q_ASSIGN U15593 ( .B(clk), .A(\g.we_clk [797]));
Q_ASSIGN U15594 ( .B(clk), .A(\g.we_clk [796]));
Q_ASSIGN U15595 ( .B(clk), .A(\g.we_clk [795]));
Q_ASSIGN U15596 ( .B(clk), .A(\g.we_clk [794]));
Q_ASSIGN U15597 ( .B(clk), .A(\g.we_clk [793]));
Q_ASSIGN U15598 ( .B(clk), .A(\g.we_clk [792]));
Q_ASSIGN U15599 ( .B(clk), .A(\g.we_clk [791]));
Q_ASSIGN U15600 ( .B(clk), .A(\g.we_clk [790]));
Q_ASSIGN U15601 ( .B(clk), .A(\g.we_clk [789]));
Q_ASSIGN U15602 ( .B(clk), .A(\g.we_clk [788]));
Q_ASSIGN U15603 ( .B(clk), .A(\g.we_clk [787]));
Q_ASSIGN U15604 ( .B(clk), .A(\g.we_clk [786]));
Q_ASSIGN U15605 ( .B(clk), .A(\g.we_clk [785]));
Q_ASSIGN U15606 ( .B(clk), .A(\g.we_clk [784]));
Q_ASSIGN U15607 ( .B(clk), .A(\g.we_clk [783]));
Q_ASSIGN U15608 ( .B(clk), .A(\g.we_clk [782]));
Q_ASSIGN U15609 ( .B(clk), .A(\g.we_clk [781]));
Q_ASSIGN U15610 ( .B(clk), .A(\g.we_clk [780]));
Q_ASSIGN U15611 ( .B(clk), .A(\g.we_clk [779]));
Q_ASSIGN U15612 ( .B(clk), .A(\g.we_clk [778]));
Q_ASSIGN U15613 ( .B(clk), .A(\g.we_clk [777]));
Q_ASSIGN U15614 ( .B(clk), .A(\g.we_clk [776]));
Q_ASSIGN U15615 ( .B(clk), .A(\g.we_clk [775]));
Q_ASSIGN U15616 ( .B(clk), .A(\g.we_clk [774]));
Q_ASSIGN U15617 ( .B(clk), .A(\g.we_clk [773]));
Q_ASSIGN U15618 ( .B(clk), .A(\g.we_clk [772]));
Q_ASSIGN U15619 ( .B(clk), .A(\g.we_clk [771]));
Q_ASSIGN U15620 ( .B(clk), .A(\g.we_clk [770]));
Q_ASSIGN U15621 ( .B(clk), .A(\g.we_clk [769]));
Q_ASSIGN U15622 ( .B(clk), .A(\g.we_clk [768]));
Q_ASSIGN U15623 ( .B(clk), .A(\g.we_clk [767]));
Q_ASSIGN U15624 ( .B(clk), .A(\g.we_clk [766]));
Q_ASSIGN U15625 ( .B(clk), .A(\g.we_clk [765]));
Q_ASSIGN U15626 ( .B(clk), .A(\g.we_clk [764]));
Q_ASSIGN U15627 ( .B(clk), .A(\g.we_clk [763]));
Q_ASSIGN U15628 ( .B(clk), .A(\g.we_clk [762]));
Q_ASSIGN U15629 ( .B(clk), .A(\g.we_clk [761]));
Q_ASSIGN U15630 ( .B(clk), .A(\g.we_clk [760]));
Q_ASSIGN U15631 ( .B(clk), .A(\g.we_clk [759]));
Q_ASSIGN U15632 ( .B(clk), .A(\g.we_clk [758]));
Q_ASSIGN U15633 ( .B(clk), .A(\g.we_clk [757]));
Q_ASSIGN U15634 ( .B(clk), .A(\g.we_clk [756]));
Q_ASSIGN U15635 ( .B(clk), .A(\g.we_clk [755]));
Q_ASSIGN U15636 ( .B(clk), .A(\g.we_clk [754]));
Q_ASSIGN U15637 ( .B(clk), .A(\g.we_clk [753]));
Q_ASSIGN U15638 ( .B(clk), .A(\g.we_clk [752]));
Q_ASSIGN U15639 ( .B(clk), .A(\g.we_clk [751]));
Q_ASSIGN U15640 ( .B(clk), .A(\g.we_clk [750]));
Q_ASSIGN U15641 ( .B(clk), .A(\g.we_clk [749]));
Q_ASSIGN U15642 ( .B(clk), .A(\g.we_clk [748]));
Q_ASSIGN U15643 ( .B(clk), .A(\g.we_clk [747]));
Q_ASSIGN U15644 ( .B(clk), .A(\g.we_clk [746]));
Q_ASSIGN U15645 ( .B(clk), .A(\g.we_clk [745]));
Q_ASSIGN U15646 ( .B(clk), .A(\g.we_clk [744]));
Q_ASSIGN U15647 ( .B(clk), .A(\g.we_clk [743]));
Q_ASSIGN U15648 ( .B(clk), .A(\g.we_clk [742]));
Q_ASSIGN U15649 ( .B(clk), .A(\g.we_clk [741]));
Q_ASSIGN U15650 ( .B(clk), .A(\g.we_clk [740]));
Q_ASSIGN U15651 ( .B(clk), .A(\g.we_clk [739]));
Q_ASSIGN U15652 ( .B(clk), .A(\g.we_clk [738]));
Q_ASSIGN U15653 ( .B(clk), .A(\g.we_clk [737]));
Q_ASSIGN U15654 ( .B(clk), .A(\g.we_clk [736]));
Q_ASSIGN U15655 ( .B(clk), .A(\g.we_clk [735]));
Q_ASSIGN U15656 ( .B(clk), .A(\g.we_clk [734]));
Q_ASSIGN U15657 ( .B(clk), .A(\g.we_clk [733]));
Q_ASSIGN U15658 ( .B(clk), .A(\g.we_clk [732]));
Q_ASSIGN U15659 ( .B(clk), .A(\g.we_clk [731]));
Q_ASSIGN U15660 ( .B(clk), .A(\g.we_clk [730]));
Q_ASSIGN U15661 ( .B(clk), .A(\g.we_clk [729]));
Q_ASSIGN U15662 ( .B(clk), .A(\g.we_clk [728]));
Q_ASSIGN U15663 ( .B(clk), .A(\g.we_clk [727]));
Q_ASSIGN U15664 ( .B(clk), .A(\g.we_clk [726]));
Q_ASSIGN U15665 ( .B(clk), .A(\g.we_clk [725]));
Q_ASSIGN U15666 ( .B(clk), .A(\g.we_clk [724]));
Q_ASSIGN U15667 ( .B(clk), .A(\g.we_clk [723]));
Q_ASSIGN U15668 ( .B(clk), .A(\g.we_clk [722]));
Q_ASSIGN U15669 ( .B(clk), .A(\g.we_clk [721]));
Q_ASSIGN U15670 ( .B(clk), .A(\g.we_clk [720]));
Q_ASSIGN U15671 ( .B(clk), .A(\g.we_clk [719]));
Q_ASSIGN U15672 ( .B(clk), .A(\g.we_clk [718]));
Q_ASSIGN U15673 ( .B(clk), .A(\g.we_clk [717]));
Q_ASSIGN U15674 ( .B(clk), .A(\g.we_clk [716]));
Q_ASSIGN U15675 ( .B(clk), .A(\g.we_clk [715]));
Q_ASSIGN U15676 ( .B(clk), .A(\g.we_clk [714]));
Q_ASSIGN U15677 ( .B(clk), .A(\g.we_clk [713]));
Q_ASSIGN U15678 ( .B(clk), .A(\g.we_clk [712]));
Q_ASSIGN U15679 ( .B(clk), .A(\g.we_clk [711]));
Q_ASSIGN U15680 ( .B(clk), .A(\g.we_clk [710]));
Q_ASSIGN U15681 ( .B(clk), .A(\g.we_clk [709]));
Q_ASSIGN U15682 ( .B(clk), .A(\g.we_clk [708]));
Q_ASSIGN U15683 ( .B(clk), .A(\g.we_clk [707]));
Q_ASSIGN U15684 ( .B(clk), .A(\g.we_clk [706]));
Q_ASSIGN U15685 ( .B(clk), .A(\g.we_clk [705]));
Q_ASSIGN U15686 ( .B(clk), .A(\g.we_clk [704]));
Q_ASSIGN U15687 ( .B(clk), .A(\g.we_clk [703]));
Q_ASSIGN U15688 ( .B(clk), .A(\g.we_clk [702]));
Q_ASSIGN U15689 ( .B(clk), .A(\g.we_clk [701]));
Q_ASSIGN U15690 ( .B(clk), .A(\g.we_clk [700]));
Q_ASSIGN U15691 ( .B(clk), .A(\g.we_clk [699]));
Q_ASSIGN U15692 ( .B(clk), .A(\g.we_clk [698]));
Q_ASSIGN U15693 ( .B(clk), .A(\g.we_clk [697]));
Q_ASSIGN U15694 ( .B(clk), .A(\g.we_clk [696]));
Q_ASSIGN U15695 ( .B(clk), .A(\g.we_clk [695]));
Q_ASSIGN U15696 ( .B(clk), .A(\g.we_clk [694]));
Q_ASSIGN U15697 ( .B(clk), .A(\g.we_clk [693]));
Q_ASSIGN U15698 ( .B(clk), .A(\g.we_clk [692]));
Q_ASSIGN U15699 ( .B(clk), .A(\g.we_clk [691]));
Q_ASSIGN U15700 ( .B(clk), .A(\g.we_clk [690]));
Q_ASSIGN U15701 ( .B(clk), .A(\g.we_clk [689]));
Q_ASSIGN U15702 ( .B(clk), .A(\g.we_clk [688]));
Q_ASSIGN U15703 ( .B(clk), .A(\g.we_clk [687]));
Q_ASSIGN U15704 ( .B(clk), .A(\g.we_clk [686]));
Q_ASSIGN U15705 ( .B(clk), .A(\g.we_clk [685]));
Q_ASSIGN U15706 ( .B(clk), .A(\g.we_clk [684]));
Q_ASSIGN U15707 ( .B(clk), .A(\g.we_clk [683]));
Q_ASSIGN U15708 ( .B(clk), .A(\g.we_clk [682]));
Q_ASSIGN U15709 ( .B(clk), .A(\g.we_clk [681]));
Q_ASSIGN U15710 ( .B(clk), .A(\g.we_clk [680]));
Q_ASSIGN U15711 ( .B(clk), .A(\g.we_clk [679]));
Q_ASSIGN U15712 ( .B(clk), .A(\g.we_clk [678]));
Q_ASSIGN U15713 ( .B(clk), .A(\g.we_clk [677]));
Q_ASSIGN U15714 ( .B(clk), .A(\g.we_clk [676]));
Q_ASSIGN U15715 ( .B(clk), .A(\g.we_clk [675]));
Q_ASSIGN U15716 ( .B(clk), .A(\g.we_clk [674]));
Q_ASSIGN U15717 ( .B(clk), .A(\g.we_clk [673]));
Q_ASSIGN U15718 ( .B(clk), .A(\g.we_clk [672]));
Q_ASSIGN U15719 ( .B(clk), .A(\g.we_clk [671]));
Q_ASSIGN U15720 ( .B(clk), .A(\g.we_clk [670]));
Q_ASSIGN U15721 ( .B(clk), .A(\g.we_clk [669]));
Q_ASSIGN U15722 ( .B(clk), .A(\g.we_clk [668]));
Q_ASSIGN U15723 ( .B(clk), .A(\g.we_clk [667]));
Q_ASSIGN U15724 ( .B(clk), .A(\g.we_clk [666]));
Q_ASSIGN U15725 ( .B(clk), .A(\g.we_clk [665]));
Q_ASSIGN U15726 ( .B(clk), .A(\g.we_clk [664]));
Q_ASSIGN U15727 ( .B(clk), .A(\g.we_clk [663]));
Q_ASSIGN U15728 ( .B(clk), .A(\g.we_clk [662]));
Q_ASSIGN U15729 ( .B(clk), .A(\g.we_clk [661]));
Q_ASSIGN U15730 ( .B(clk), .A(\g.we_clk [660]));
Q_ASSIGN U15731 ( .B(clk), .A(\g.we_clk [659]));
Q_ASSIGN U15732 ( .B(clk), .A(\g.we_clk [658]));
Q_ASSIGN U15733 ( .B(clk), .A(\g.we_clk [657]));
Q_ASSIGN U15734 ( .B(clk), .A(\g.we_clk [656]));
Q_ASSIGN U15735 ( .B(clk), .A(\g.we_clk [655]));
Q_ASSIGN U15736 ( .B(clk), .A(\g.we_clk [654]));
Q_ASSIGN U15737 ( .B(clk), .A(\g.we_clk [653]));
Q_ASSIGN U15738 ( .B(clk), .A(\g.we_clk [652]));
Q_ASSIGN U15739 ( .B(clk), .A(\g.we_clk [651]));
Q_ASSIGN U15740 ( .B(clk), .A(\g.we_clk [650]));
Q_ASSIGN U15741 ( .B(clk), .A(\g.we_clk [649]));
Q_ASSIGN U15742 ( .B(clk), .A(\g.we_clk [648]));
Q_ASSIGN U15743 ( .B(clk), .A(\g.we_clk [647]));
Q_ASSIGN U15744 ( .B(clk), .A(\g.we_clk [646]));
Q_ASSIGN U15745 ( .B(clk), .A(\g.we_clk [645]));
Q_ASSIGN U15746 ( .B(clk), .A(\g.we_clk [644]));
Q_ASSIGN U15747 ( .B(clk), .A(\g.we_clk [643]));
Q_ASSIGN U15748 ( .B(clk), .A(\g.we_clk [642]));
Q_ASSIGN U15749 ( .B(clk), .A(\g.we_clk [641]));
Q_ASSIGN U15750 ( .B(clk), .A(\g.we_clk [640]));
Q_ASSIGN U15751 ( .B(clk), .A(\g.we_clk [639]));
Q_ASSIGN U15752 ( .B(clk), .A(\g.we_clk [638]));
Q_ASSIGN U15753 ( .B(clk), .A(\g.we_clk [637]));
Q_ASSIGN U15754 ( .B(clk), .A(\g.we_clk [636]));
Q_ASSIGN U15755 ( .B(clk), .A(\g.we_clk [635]));
Q_ASSIGN U15756 ( .B(clk), .A(\g.we_clk [634]));
Q_ASSIGN U15757 ( .B(clk), .A(\g.we_clk [633]));
Q_ASSIGN U15758 ( .B(clk), .A(\g.we_clk [632]));
Q_ASSIGN U15759 ( .B(clk), .A(\g.we_clk [631]));
Q_ASSIGN U15760 ( .B(clk), .A(\g.we_clk [630]));
Q_ASSIGN U15761 ( .B(clk), .A(\g.we_clk [629]));
Q_ASSIGN U15762 ( .B(clk), .A(\g.we_clk [628]));
Q_ASSIGN U15763 ( .B(clk), .A(\g.we_clk [627]));
Q_ASSIGN U15764 ( .B(clk), .A(\g.we_clk [626]));
Q_ASSIGN U15765 ( .B(clk), .A(\g.we_clk [625]));
Q_ASSIGN U15766 ( .B(clk), .A(\g.we_clk [624]));
Q_ASSIGN U15767 ( .B(clk), .A(\g.we_clk [623]));
Q_ASSIGN U15768 ( .B(clk), .A(\g.we_clk [622]));
Q_ASSIGN U15769 ( .B(clk), .A(\g.we_clk [621]));
Q_ASSIGN U15770 ( .B(clk), .A(\g.we_clk [620]));
Q_ASSIGN U15771 ( .B(clk), .A(\g.we_clk [619]));
Q_ASSIGN U15772 ( .B(clk), .A(\g.we_clk [618]));
Q_ASSIGN U15773 ( .B(clk), .A(\g.we_clk [617]));
Q_ASSIGN U15774 ( .B(clk), .A(\g.we_clk [616]));
Q_ASSIGN U15775 ( .B(clk), .A(\g.we_clk [615]));
Q_ASSIGN U15776 ( .B(clk), .A(\g.we_clk [614]));
Q_ASSIGN U15777 ( .B(clk), .A(\g.we_clk [613]));
Q_ASSIGN U15778 ( .B(clk), .A(\g.we_clk [612]));
Q_ASSIGN U15779 ( .B(clk), .A(\g.we_clk [611]));
Q_ASSIGN U15780 ( .B(clk), .A(\g.we_clk [610]));
Q_ASSIGN U15781 ( .B(clk), .A(\g.we_clk [609]));
Q_ASSIGN U15782 ( .B(clk), .A(\g.we_clk [608]));
Q_ASSIGN U15783 ( .B(clk), .A(\g.we_clk [607]));
Q_ASSIGN U15784 ( .B(clk), .A(\g.we_clk [606]));
Q_ASSIGN U15785 ( .B(clk), .A(\g.we_clk [605]));
Q_ASSIGN U15786 ( .B(clk), .A(\g.we_clk [604]));
Q_ASSIGN U15787 ( .B(clk), .A(\g.we_clk [603]));
Q_ASSIGN U15788 ( .B(clk), .A(\g.we_clk [602]));
Q_ASSIGN U15789 ( .B(clk), .A(\g.we_clk [601]));
Q_ASSIGN U15790 ( .B(clk), .A(\g.we_clk [600]));
Q_ASSIGN U15791 ( .B(clk), .A(\g.we_clk [599]));
Q_ASSIGN U15792 ( .B(clk), .A(\g.we_clk [598]));
Q_ASSIGN U15793 ( .B(clk), .A(\g.we_clk [597]));
Q_ASSIGN U15794 ( .B(clk), .A(\g.we_clk [596]));
Q_ASSIGN U15795 ( .B(clk), .A(\g.we_clk [595]));
Q_ASSIGN U15796 ( .B(clk), .A(\g.we_clk [594]));
Q_ASSIGN U15797 ( .B(clk), .A(\g.we_clk [593]));
Q_ASSIGN U15798 ( .B(clk), .A(\g.we_clk [592]));
Q_ASSIGN U15799 ( .B(clk), .A(\g.we_clk [591]));
Q_ASSIGN U15800 ( .B(clk), .A(\g.we_clk [590]));
Q_ASSIGN U15801 ( .B(clk), .A(\g.we_clk [589]));
Q_ASSIGN U15802 ( .B(clk), .A(\g.we_clk [588]));
Q_ASSIGN U15803 ( .B(clk), .A(\g.we_clk [587]));
Q_ASSIGN U15804 ( .B(clk), .A(\g.we_clk [586]));
Q_ASSIGN U15805 ( .B(clk), .A(\g.we_clk [585]));
Q_ASSIGN U15806 ( .B(clk), .A(\g.we_clk [584]));
Q_ASSIGN U15807 ( .B(clk), .A(\g.we_clk [583]));
Q_ASSIGN U15808 ( .B(clk), .A(\g.we_clk [582]));
Q_ASSIGN U15809 ( .B(clk), .A(\g.we_clk [581]));
Q_ASSIGN U15810 ( .B(clk), .A(\g.we_clk [580]));
Q_ASSIGN U15811 ( .B(clk), .A(\g.we_clk [579]));
Q_ASSIGN U15812 ( .B(clk), .A(\g.we_clk [578]));
Q_ASSIGN U15813 ( .B(clk), .A(\g.we_clk [577]));
Q_ASSIGN U15814 ( .B(clk), .A(\g.we_clk [576]));
Q_ASSIGN U15815 ( .B(clk), .A(\g.we_clk [575]));
Q_ASSIGN U15816 ( .B(clk), .A(\g.we_clk [574]));
Q_ASSIGN U15817 ( .B(clk), .A(\g.we_clk [573]));
Q_ASSIGN U15818 ( .B(clk), .A(\g.we_clk [572]));
Q_ASSIGN U15819 ( .B(clk), .A(\g.we_clk [571]));
Q_ASSIGN U15820 ( .B(clk), .A(\g.we_clk [570]));
Q_ASSIGN U15821 ( .B(clk), .A(\g.we_clk [569]));
Q_ASSIGN U15822 ( .B(clk), .A(\g.we_clk [568]));
Q_ASSIGN U15823 ( .B(clk), .A(\g.we_clk [567]));
Q_ASSIGN U15824 ( .B(clk), .A(\g.we_clk [566]));
Q_ASSIGN U15825 ( .B(clk), .A(\g.we_clk [565]));
Q_ASSIGN U15826 ( .B(clk), .A(\g.we_clk [564]));
Q_ASSIGN U15827 ( .B(clk), .A(\g.we_clk [563]));
Q_ASSIGN U15828 ( .B(clk), .A(\g.we_clk [562]));
Q_ASSIGN U15829 ( .B(clk), .A(\g.we_clk [561]));
Q_ASSIGN U15830 ( .B(clk), .A(\g.we_clk [560]));
Q_ASSIGN U15831 ( .B(clk), .A(\g.we_clk [559]));
Q_ASSIGN U15832 ( .B(clk), .A(\g.we_clk [558]));
Q_ASSIGN U15833 ( .B(clk), .A(\g.we_clk [557]));
Q_ASSIGN U15834 ( .B(clk), .A(\g.we_clk [556]));
Q_ASSIGN U15835 ( .B(clk), .A(\g.we_clk [555]));
Q_ASSIGN U15836 ( .B(clk), .A(\g.we_clk [554]));
Q_ASSIGN U15837 ( .B(clk), .A(\g.we_clk [553]));
Q_ASSIGN U15838 ( .B(clk), .A(\g.we_clk [552]));
Q_ASSIGN U15839 ( .B(clk), .A(\g.we_clk [551]));
Q_ASSIGN U15840 ( .B(clk), .A(\g.we_clk [550]));
Q_ASSIGN U15841 ( .B(clk), .A(\g.we_clk [549]));
Q_ASSIGN U15842 ( .B(clk), .A(\g.we_clk [548]));
Q_ASSIGN U15843 ( .B(clk), .A(\g.we_clk [547]));
Q_ASSIGN U15844 ( .B(clk), .A(\g.we_clk [546]));
Q_ASSIGN U15845 ( .B(clk), .A(\g.we_clk [545]));
Q_ASSIGN U15846 ( .B(clk), .A(\g.we_clk [544]));
Q_ASSIGN U15847 ( .B(clk), .A(\g.we_clk [543]));
Q_ASSIGN U15848 ( .B(clk), .A(\g.we_clk [542]));
Q_ASSIGN U15849 ( .B(clk), .A(\g.we_clk [541]));
Q_ASSIGN U15850 ( .B(clk), .A(\g.we_clk [540]));
Q_ASSIGN U15851 ( .B(clk), .A(\g.we_clk [539]));
Q_ASSIGN U15852 ( .B(clk), .A(\g.we_clk [538]));
Q_ASSIGN U15853 ( .B(clk), .A(\g.we_clk [537]));
Q_ASSIGN U15854 ( .B(clk), .A(\g.we_clk [536]));
Q_ASSIGN U15855 ( .B(clk), .A(\g.we_clk [535]));
Q_ASSIGN U15856 ( .B(clk), .A(\g.we_clk [534]));
Q_ASSIGN U15857 ( .B(clk), .A(\g.we_clk [533]));
Q_ASSIGN U15858 ( .B(clk), .A(\g.we_clk [532]));
Q_ASSIGN U15859 ( .B(clk), .A(\g.we_clk [531]));
Q_ASSIGN U15860 ( .B(clk), .A(\g.we_clk [530]));
Q_ASSIGN U15861 ( .B(clk), .A(\g.we_clk [529]));
Q_ASSIGN U15862 ( .B(clk), .A(\g.we_clk [528]));
Q_ASSIGN U15863 ( .B(clk), .A(\g.we_clk [527]));
Q_ASSIGN U15864 ( .B(clk), .A(\g.we_clk [526]));
Q_ASSIGN U15865 ( .B(clk), .A(\g.we_clk [525]));
Q_ASSIGN U15866 ( .B(clk), .A(\g.we_clk [524]));
Q_ASSIGN U15867 ( .B(clk), .A(\g.we_clk [523]));
Q_ASSIGN U15868 ( .B(clk), .A(\g.we_clk [522]));
Q_ASSIGN U15869 ( .B(clk), .A(\g.we_clk [521]));
Q_ASSIGN U15870 ( .B(clk), .A(\g.we_clk [520]));
Q_ASSIGN U15871 ( .B(clk), .A(\g.we_clk [519]));
Q_ASSIGN U15872 ( .B(clk), .A(\g.we_clk [518]));
Q_ASSIGN U15873 ( .B(clk), .A(\g.we_clk [517]));
Q_ASSIGN U15874 ( .B(clk), .A(\g.we_clk [516]));
Q_ASSIGN U15875 ( .B(clk), .A(\g.we_clk [515]));
Q_ASSIGN U15876 ( .B(clk), .A(\g.we_clk [514]));
Q_ASSIGN U15877 ( .B(clk), .A(\g.we_clk [513]));
Q_ASSIGN U15878 ( .B(clk), .A(\g.we_clk [512]));
Q_ASSIGN U15879 ( .B(clk), .A(\g.we_clk [511]));
Q_ASSIGN U15880 ( .B(clk), .A(\g.we_clk [510]));
Q_ASSIGN U15881 ( .B(clk), .A(\g.we_clk [509]));
Q_ASSIGN U15882 ( .B(clk), .A(\g.we_clk [508]));
Q_ASSIGN U15883 ( .B(clk), .A(\g.we_clk [507]));
Q_ASSIGN U15884 ( .B(clk), .A(\g.we_clk [506]));
Q_ASSIGN U15885 ( .B(clk), .A(\g.we_clk [505]));
Q_ASSIGN U15886 ( .B(clk), .A(\g.we_clk [504]));
Q_ASSIGN U15887 ( .B(clk), .A(\g.we_clk [503]));
Q_ASSIGN U15888 ( .B(clk), .A(\g.we_clk [502]));
Q_ASSIGN U15889 ( .B(clk), .A(\g.we_clk [501]));
Q_ASSIGN U15890 ( .B(clk), .A(\g.we_clk [500]));
Q_ASSIGN U15891 ( .B(clk), .A(\g.we_clk [499]));
Q_ASSIGN U15892 ( .B(clk), .A(\g.we_clk [498]));
Q_ASSIGN U15893 ( .B(clk), .A(\g.we_clk [497]));
Q_ASSIGN U15894 ( .B(clk), .A(\g.we_clk [496]));
Q_ASSIGN U15895 ( .B(clk), .A(\g.we_clk [495]));
Q_ASSIGN U15896 ( .B(clk), .A(\g.we_clk [494]));
Q_ASSIGN U15897 ( .B(clk), .A(\g.we_clk [493]));
Q_ASSIGN U15898 ( .B(clk), .A(\g.we_clk [492]));
Q_ASSIGN U15899 ( .B(clk), .A(\g.we_clk [491]));
Q_ASSIGN U15900 ( .B(clk), .A(\g.we_clk [490]));
Q_ASSIGN U15901 ( .B(clk), .A(\g.we_clk [489]));
Q_ASSIGN U15902 ( .B(clk), .A(\g.we_clk [488]));
Q_ASSIGN U15903 ( .B(clk), .A(\g.we_clk [487]));
Q_ASSIGN U15904 ( .B(clk), .A(\g.we_clk [486]));
Q_ASSIGN U15905 ( .B(clk), .A(\g.we_clk [485]));
Q_ASSIGN U15906 ( .B(clk), .A(\g.we_clk [484]));
Q_ASSIGN U15907 ( .B(clk), .A(\g.we_clk [483]));
Q_ASSIGN U15908 ( .B(clk), .A(\g.we_clk [482]));
Q_ASSIGN U15909 ( .B(clk), .A(\g.we_clk [481]));
Q_ASSIGN U15910 ( .B(clk), .A(\g.we_clk [480]));
Q_ASSIGN U15911 ( .B(clk), .A(\g.we_clk [479]));
Q_ASSIGN U15912 ( .B(clk), .A(\g.we_clk [478]));
Q_ASSIGN U15913 ( .B(clk), .A(\g.we_clk [477]));
Q_ASSIGN U15914 ( .B(clk), .A(\g.we_clk [476]));
Q_ASSIGN U15915 ( .B(clk), .A(\g.we_clk [475]));
Q_ASSIGN U15916 ( .B(clk), .A(\g.we_clk [474]));
Q_ASSIGN U15917 ( .B(clk), .A(\g.we_clk [473]));
Q_ASSIGN U15918 ( .B(clk), .A(\g.we_clk [472]));
Q_ASSIGN U15919 ( .B(clk), .A(\g.we_clk [471]));
Q_ASSIGN U15920 ( .B(clk), .A(\g.we_clk [470]));
Q_ASSIGN U15921 ( .B(clk), .A(\g.we_clk [469]));
Q_ASSIGN U15922 ( .B(clk), .A(\g.we_clk [468]));
Q_ASSIGN U15923 ( .B(clk), .A(\g.we_clk [467]));
Q_ASSIGN U15924 ( .B(clk), .A(\g.we_clk [466]));
Q_ASSIGN U15925 ( .B(clk), .A(\g.we_clk [465]));
Q_ASSIGN U15926 ( .B(clk), .A(\g.we_clk [464]));
Q_ASSIGN U15927 ( .B(clk), .A(\g.we_clk [463]));
Q_ASSIGN U15928 ( .B(clk), .A(\g.we_clk [462]));
Q_ASSIGN U15929 ( .B(clk), .A(\g.we_clk [461]));
Q_ASSIGN U15930 ( .B(clk), .A(\g.we_clk [460]));
Q_ASSIGN U15931 ( .B(clk), .A(\g.we_clk [459]));
Q_ASSIGN U15932 ( .B(clk), .A(\g.we_clk [458]));
Q_ASSIGN U15933 ( .B(clk), .A(\g.we_clk [457]));
Q_ASSIGN U15934 ( .B(clk), .A(\g.we_clk [456]));
Q_ASSIGN U15935 ( .B(clk), .A(\g.we_clk [455]));
Q_ASSIGN U15936 ( .B(clk), .A(\g.we_clk [454]));
Q_ASSIGN U15937 ( .B(clk), .A(\g.we_clk [453]));
Q_ASSIGN U15938 ( .B(clk), .A(\g.we_clk [452]));
Q_ASSIGN U15939 ( .B(clk), .A(\g.we_clk [451]));
Q_ASSIGN U15940 ( .B(clk), .A(\g.we_clk [450]));
Q_ASSIGN U15941 ( .B(clk), .A(\g.we_clk [449]));
Q_ASSIGN U15942 ( .B(clk), .A(\g.we_clk [448]));
Q_ASSIGN U15943 ( .B(clk), .A(\g.we_clk [447]));
Q_ASSIGN U15944 ( .B(clk), .A(\g.we_clk [446]));
Q_ASSIGN U15945 ( .B(clk), .A(\g.we_clk [445]));
Q_ASSIGN U15946 ( .B(clk), .A(\g.we_clk [444]));
Q_ASSIGN U15947 ( .B(clk), .A(\g.we_clk [443]));
Q_ASSIGN U15948 ( .B(clk), .A(\g.we_clk [442]));
Q_ASSIGN U15949 ( .B(clk), .A(\g.we_clk [441]));
Q_ASSIGN U15950 ( .B(clk), .A(\g.we_clk [440]));
Q_ASSIGN U15951 ( .B(clk), .A(\g.we_clk [439]));
Q_ASSIGN U15952 ( .B(clk), .A(\g.we_clk [438]));
Q_ASSIGN U15953 ( .B(clk), .A(\g.we_clk [437]));
Q_ASSIGN U15954 ( .B(clk), .A(\g.we_clk [436]));
Q_ASSIGN U15955 ( .B(clk), .A(\g.we_clk [435]));
Q_ASSIGN U15956 ( .B(clk), .A(\g.we_clk [434]));
Q_ASSIGN U15957 ( .B(clk), .A(\g.we_clk [433]));
Q_ASSIGN U15958 ( .B(clk), .A(\g.we_clk [432]));
Q_ASSIGN U15959 ( .B(clk), .A(\g.we_clk [431]));
Q_ASSIGN U15960 ( .B(clk), .A(\g.we_clk [430]));
Q_ASSIGN U15961 ( .B(clk), .A(\g.we_clk [429]));
Q_ASSIGN U15962 ( .B(clk), .A(\g.we_clk [428]));
Q_ASSIGN U15963 ( .B(clk), .A(\g.we_clk [427]));
Q_ASSIGN U15964 ( .B(clk), .A(\g.we_clk [426]));
Q_ASSIGN U15965 ( .B(clk), .A(\g.we_clk [425]));
Q_ASSIGN U15966 ( .B(clk), .A(\g.we_clk [424]));
Q_ASSIGN U15967 ( .B(clk), .A(\g.we_clk [423]));
Q_ASSIGN U15968 ( .B(clk), .A(\g.we_clk [422]));
Q_ASSIGN U15969 ( .B(clk), .A(\g.we_clk [421]));
Q_ASSIGN U15970 ( .B(clk), .A(\g.we_clk [420]));
Q_ASSIGN U15971 ( .B(clk), .A(\g.we_clk [419]));
Q_ASSIGN U15972 ( .B(clk), .A(\g.we_clk [418]));
Q_ASSIGN U15973 ( .B(clk), .A(\g.we_clk [417]));
Q_ASSIGN U15974 ( .B(clk), .A(\g.we_clk [416]));
Q_ASSIGN U15975 ( .B(clk), .A(\g.we_clk [415]));
Q_ASSIGN U15976 ( .B(clk), .A(\g.we_clk [414]));
Q_ASSIGN U15977 ( .B(clk), .A(\g.we_clk [413]));
Q_ASSIGN U15978 ( .B(clk), .A(\g.we_clk [412]));
Q_ASSIGN U15979 ( .B(clk), .A(\g.we_clk [411]));
Q_ASSIGN U15980 ( .B(clk), .A(\g.we_clk [410]));
Q_ASSIGN U15981 ( .B(clk), .A(\g.we_clk [409]));
Q_ASSIGN U15982 ( .B(clk), .A(\g.we_clk [408]));
Q_ASSIGN U15983 ( .B(clk), .A(\g.we_clk [407]));
Q_ASSIGN U15984 ( .B(clk), .A(\g.we_clk [406]));
Q_ASSIGN U15985 ( .B(clk), .A(\g.we_clk [405]));
Q_ASSIGN U15986 ( .B(clk), .A(\g.we_clk [404]));
Q_ASSIGN U15987 ( .B(clk), .A(\g.we_clk [403]));
Q_ASSIGN U15988 ( .B(clk), .A(\g.we_clk [402]));
Q_ASSIGN U15989 ( .B(clk), .A(\g.we_clk [401]));
Q_ASSIGN U15990 ( .B(clk), .A(\g.we_clk [400]));
Q_ASSIGN U15991 ( .B(clk), .A(\g.we_clk [399]));
Q_ASSIGN U15992 ( .B(clk), .A(\g.we_clk [398]));
Q_ASSIGN U15993 ( .B(clk), .A(\g.we_clk [397]));
Q_ASSIGN U15994 ( .B(clk), .A(\g.we_clk [396]));
Q_ASSIGN U15995 ( .B(clk), .A(\g.we_clk [395]));
Q_ASSIGN U15996 ( .B(clk), .A(\g.we_clk [394]));
Q_ASSIGN U15997 ( .B(clk), .A(\g.we_clk [393]));
Q_ASSIGN U15998 ( .B(clk), .A(\g.we_clk [392]));
Q_ASSIGN U15999 ( .B(clk), .A(\g.we_clk [391]));
Q_ASSIGN U16000 ( .B(clk), .A(\g.we_clk [390]));
Q_ASSIGN U16001 ( .B(clk), .A(\g.we_clk [389]));
Q_ASSIGN U16002 ( .B(clk), .A(\g.we_clk [388]));
Q_ASSIGN U16003 ( .B(clk), .A(\g.we_clk [387]));
Q_ASSIGN U16004 ( .B(clk), .A(\g.we_clk [386]));
Q_ASSIGN U16005 ( .B(clk), .A(\g.we_clk [385]));
Q_ASSIGN U16006 ( .B(clk), .A(\g.we_clk [384]));
Q_ASSIGN U16007 ( .B(clk), .A(\g.we_clk [383]));
Q_ASSIGN U16008 ( .B(clk), .A(\g.we_clk [382]));
Q_ASSIGN U16009 ( .B(clk), .A(\g.we_clk [381]));
Q_ASSIGN U16010 ( .B(clk), .A(\g.we_clk [380]));
Q_ASSIGN U16011 ( .B(clk), .A(\g.we_clk [379]));
Q_ASSIGN U16012 ( .B(clk), .A(\g.we_clk [378]));
Q_ASSIGN U16013 ( .B(clk), .A(\g.we_clk [377]));
Q_ASSIGN U16014 ( .B(clk), .A(\g.we_clk [376]));
Q_ASSIGN U16015 ( .B(clk), .A(\g.we_clk [375]));
Q_ASSIGN U16016 ( .B(clk), .A(\g.we_clk [374]));
Q_ASSIGN U16017 ( .B(clk), .A(\g.we_clk [373]));
Q_ASSIGN U16018 ( .B(clk), .A(\g.we_clk [372]));
Q_ASSIGN U16019 ( .B(clk), .A(\g.we_clk [371]));
Q_ASSIGN U16020 ( .B(clk), .A(\g.we_clk [370]));
Q_ASSIGN U16021 ( .B(clk), .A(\g.we_clk [369]));
Q_ASSIGN U16022 ( .B(clk), .A(\g.we_clk [368]));
Q_ASSIGN U16023 ( .B(clk), .A(\g.we_clk [367]));
Q_ASSIGN U16024 ( .B(clk), .A(\g.we_clk [366]));
Q_ASSIGN U16025 ( .B(clk), .A(\g.we_clk [365]));
Q_ASSIGN U16026 ( .B(clk), .A(\g.we_clk [364]));
Q_ASSIGN U16027 ( .B(clk), .A(\g.we_clk [363]));
Q_ASSIGN U16028 ( .B(clk), .A(\g.we_clk [362]));
Q_ASSIGN U16029 ( .B(clk), .A(\g.we_clk [361]));
Q_ASSIGN U16030 ( .B(clk), .A(\g.we_clk [360]));
Q_ASSIGN U16031 ( .B(clk), .A(\g.we_clk [359]));
Q_ASSIGN U16032 ( .B(clk), .A(\g.we_clk [358]));
Q_ASSIGN U16033 ( .B(clk), .A(\g.we_clk [357]));
Q_ASSIGN U16034 ( .B(clk), .A(\g.we_clk [356]));
Q_ASSIGN U16035 ( .B(clk), .A(\g.we_clk [355]));
Q_ASSIGN U16036 ( .B(clk), .A(\g.we_clk [354]));
Q_ASSIGN U16037 ( .B(clk), .A(\g.we_clk [353]));
Q_ASSIGN U16038 ( .B(clk), .A(\g.we_clk [352]));
Q_ASSIGN U16039 ( .B(clk), .A(\g.we_clk [351]));
Q_ASSIGN U16040 ( .B(clk), .A(\g.we_clk [350]));
Q_ASSIGN U16041 ( .B(clk), .A(\g.we_clk [349]));
Q_ASSIGN U16042 ( .B(clk), .A(\g.we_clk [348]));
Q_ASSIGN U16043 ( .B(clk), .A(\g.we_clk [347]));
Q_ASSIGN U16044 ( .B(clk), .A(\g.we_clk [346]));
Q_ASSIGN U16045 ( .B(clk), .A(\g.we_clk [345]));
Q_ASSIGN U16046 ( .B(clk), .A(\g.we_clk [344]));
Q_ASSIGN U16047 ( .B(clk), .A(\g.we_clk [343]));
Q_ASSIGN U16048 ( .B(clk), .A(\g.we_clk [342]));
Q_ASSIGN U16049 ( .B(clk), .A(\g.we_clk [341]));
Q_ASSIGN U16050 ( .B(clk), .A(\g.we_clk [340]));
Q_ASSIGN U16051 ( .B(clk), .A(\g.we_clk [339]));
Q_ASSIGN U16052 ( .B(clk), .A(\g.we_clk [338]));
Q_ASSIGN U16053 ( .B(clk), .A(\g.we_clk [337]));
Q_ASSIGN U16054 ( .B(clk), .A(\g.we_clk [336]));
Q_ASSIGN U16055 ( .B(clk), .A(\g.we_clk [335]));
Q_ASSIGN U16056 ( .B(clk), .A(\g.we_clk [334]));
Q_ASSIGN U16057 ( .B(clk), .A(\g.we_clk [333]));
Q_ASSIGN U16058 ( .B(clk), .A(\g.we_clk [332]));
Q_ASSIGN U16059 ( .B(clk), .A(\g.we_clk [331]));
Q_ASSIGN U16060 ( .B(clk), .A(\g.we_clk [330]));
Q_ASSIGN U16061 ( .B(clk), .A(\g.we_clk [329]));
Q_ASSIGN U16062 ( .B(clk), .A(\g.we_clk [328]));
Q_ASSIGN U16063 ( .B(clk), .A(\g.we_clk [327]));
Q_ASSIGN U16064 ( .B(clk), .A(\g.we_clk [326]));
Q_ASSIGN U16065 ( .B(clk), .A(\g.we_clk [325]));
Q_ASSIGN U16066 ( .B(clk), .A(\g.we_clk [324]));
Q_ASSIGN U16067 ( .B(clk), .A(\g.we_clk [323]));
Q_ASSIGN U16068 ( .B(clk), .A(\g.we_clk [322]));
Q_ASSIGN U16069 ( .B(clk), .A(\g.we_clk [321]));
Q_ASSIGN U16070 ( .B(clk), .A(\g.we_clk [320]));
Q_ASSIGN U16071 ( .B(clk), .A(\g.we_clk [319]));
Q_ASSIGN U16072 ( .B(clk), .A(\g.we_clk [318]));
Q_ASSIGN U16073 ( .B(clk), .A(\g.we_clk [317]));
Q_ASSIGN U16074 ( .B(clk), .A(\g.we_clk [316]));
Q_ASSIGN U16075 ( .B(clk), .A(\g.we_clk [315]));
Q_ASSIGN U16076 ( .B(clk), .A(\g.we_clk [314]));
Q_ASSIGN U16077 ( .B(clk), .A(\g.we_clk [313]));
Q_ASSIGN U16078 ( .B(clk), .A(\g.we_clk [312]));
Q_ASSIGN U16079 ( .B(clk), .A(\g.we_clk [311]));
Q_ASSIGN U16080 ( .B(clk), .A(\g.we_clk [310]));
Q_ASSIGN U16081 ( .B(clk), .A(\g.we_clk [309]));
Q_ASSIGN U16082 ( .B(clk), .A(\g.we_clk [308]));
Q_ASSIGN U16083 ( .B(clk), .A(\g.we_clk [307]));
Q_ASSIGN U16084 ( .B(clk), .A(\g.we_clk [306]));
Q_ASSIGN U16085 ( .B(clk), .A(\g.we_clk [305]));
Q_ASSIGN U16086 ( .B(clk), .A(\g.we_clk [304]));
Q_ASSIGN U16087 ( .B(clk), .A(\g.we_clk [303]));
Q_ASSIGN U16088 ( .B(clk), .A(\g.we_clk [302]));
Q_ASSIGN U16089 ( .B(clk), .A(\g.we_clk [301]));
Q_ASSIGN U16090 ( .B(clk), .A(\g.we_clk [300]));
Q_ASSIGN U16091 ( .B(clk), .A(\g.we_clk [299]));
Q_ASSIGN U16092 ( .B(clk), .A(\g.we_clk [298]));
Q_ASSIGN U16093 ( .B(clk), .A(\g.we_clk [297]));
Q_ASSIGN U16094 ( .B(clk), .A(\g.we_clk [296]));
Q_ASSIGN U16095 ( .B(clk), .A(\g.we_clk [295]));
Q_ASSIGN U16096 ( .B(clk), .A(\g.we_clk [294]));
Q_ASSIGN U16097 ( .B(clk), .A(\g.we_clk [293]));
Q_ASSIGN U16098 ( .B(clk), .A(\g.we_clk [292]));
Q_ASSIGN U16099 ( .B(clk), .A(\g.we_clk [291]));
Q_ASSIGN U16100 ( .B(clk), .A(\g.we_clk [290]));
Q_ASSIGN U16101 ( .B(clk), .A(\g.we_clk [289]));
Q_ASSIGN U16102 ( .B(clk), .A(\g.we_clk [288]));
Q_ASSIGN U16103 ( .B(clk), .A(\g.we_clk [287]));
Q_ASSIGN U16104 ( .B(clk), .A(\g.we_clk [286]));
Q_ASSIGN U16105 ( .B(clk), .A(\g.we_clk [285]));
Q_ASSIGN U16106 ( .B(clk), .A(\g.we_clk [284]));
Q_ASSIGN U16107 ( .B(clk), .A(\g.we_clk [283]));
Q_ASSIGN U16108 ( .B(clk), .A(\g.we_clk [282]));
Q_ASSIGN U16109 ( .B(clk), .A(\g.we_clk [281]));
Q_ASSIGN U16110 ( .B(clk), .A(\g.we_clk [280]));
Q_ASSIGN U16111 ( .B(clk), .A(\g.we_clk [279]));
Q_ASSIGN U16112 ( .B(clk), .A(\g.we_clk [278]));
Q_ASSIGN U16113 ( .B(clk), .A(\g.we_clk [277]));
Q_ASSIGN U16114 ( .B(clk), .A(\g.we_clk [276]));
Q_ASSIGN U16115 ( .B(clk), .A(\g.we_clk [275]));
Q_ASSIGN U16116 ( .B(clk), .A(\g.we_clk [274]));
Q_ASSIGN U16117 ( .B(clk), .A(\g.we_clk [273]));
Q_ASSIGN U16118 ( .B(clk), .A(\g.we_clk [272]));
Q_ASSIGN U16119 ( .B(clk), .A(\g.we_clk [271]));
Q_ASSIGN U16120 ( .B(clk), .A(\g.we_clk [270]));
Q_ASSIGN U16121 ( .B(clk), .A(\g.we_clk [269]));
Q_ASSIGN U16122 ( .B(clk), .A(\g.we_clk [268]));
Q_ASSIGN U16123 ( .B(clk), .A(\g.we_clk [267]));
Q_ASSIGN U16124 ( .B(clk), .A(\g.we_clk [266]));
Q_ASSIGN U16125 ( .B(clk), .A(\g.we_clk [265]));
Q_ASSIGN U16126 ( .B(clk), .A(\g.we_clk [264]));
Q_ASSIGN U16127 ( .B(clk), .A(\g.we_clk [263]));
Q_ASSIGN U16128 ( .B(clk), .A(\g.we_clk [262]));
Q_ASSIGN U16129 ( .B(clk), .A(\g.we_clk [261]));
Q_ASSIGN U16130 ( .B(clk), .A(\g.we_clk [260]));
Q_ASSIGN U16131 ( .B(clk), .A(\g.we_clk [259]));
Q_ASSIGN U16132 ( .B(clk), .A(\g.we_clk [258]));
Q_ASSIGN U16133 ( .B(clk), .A(\g.we_clk [257]));
Q_ASSIGN U16134 ( .B(clk), .A(\g.we_clk [256]));
Q_ASSIGN U16135 ( .B(clk), .A(\g.we_clk [255]));
Q_ASSIGN U16136 ( .B(clk), .A(\g.we_clk [254]));
Q_ASSIGN U16137 ( .B(clk), .A(\g.we_clk [253]));
Q_ASSIGN U16138 ( .B(clk), .A(\g.we_clk [252]));
Q_ASSIGN U16139 ( .B(clk), .A(\g.we_clk [251]));
Q_ASSIGN U16140 ( .B(clk), .A(\g.we_clk [250]));
Q_ASSIGN U16141 ( .B(clk), .A(\g.we_clk [249]));
Q_ASSIGN U16142 ( .B(clk), .A(\g.we_clk [248]));
Q_ASSIGN U16143 ( .B(clk), .A(\g.we_clk [247]));
Q_ASSIGN U16144 ( .B(clk), .A(\g.we_clk [246]));
Q_ASSIGN U16145 ( .B(clk), .A(\g.we_clk [245]));
Q_ASSIGN U16146 ( .B(clk), .A(\g.we_clk [244]));
Q_ASSIGN U16147 ( .B(clk), .A(\g.we_clk [243]));
Q_ASSIGN U16148 ( .B(clk), .A(\g.we_clk [242]));
Q_ASSIGN U16149 ( .B(clk), .A(\g.we_clk [241]));
Q_ASSIGN U16150 ( .B(clk), .A(\g.we_clk [240]));
Q_ASSIGN U16151 ( .B(clk), .A(\g.we_clk [239]));
Q_ASSIGN U16152 ( .B(clk), .A(\g.we_clk [238]));
Q_ASSIGN U16153 ( .B(clk), .A(\g.we_clk [237]));
Q_ASSIGN U16154 ( .B(clk), .A(\g.we_clk [236]));
Q_ASSIGN U16155 ( .B(clk), .A(\g.we_clk [235]));
Q_ASSIGN U16156 ( .B(clk), .A(\g.we_clk [234]));
Q_ASSIGN U16157 ( .B(clk), .A(\g.we_clk [233]));
Q_ASSIGN U16158 ( .B(clk), .A(\g.we_clk [232]));
Q_ASSIGN U16159 ( .B(clk), .A(\g.we_clk [231]));
Q_ASSIGN U16160 ( .B(clk), .A(\g.we_clk [230]));
Q_ASSIGN U16161 ( .B(clk), .A(\g.we_clk [229]));
Q_ASSIGN U16162 ( .B(clk), .A(\g.we_clk [228]));
Q_ASSIGN U16163 ( .B(clk), .A(\g.we_clk [227]));
Q_ASSIGN U16164 ( .B(clk), .A(\g.we_clk [226]));
Q_ASSIGN U16165 ( .B(clk), .A(\g.we_clk [225]));
Q_ASSIGN U16166 ( .B(clk), .A(\g.we_clk [224]));
Q_ASSIGN U16167 ( .B(clk), .A(\g.we_clk [223]));
Q_ASSIGN U16168 ( .B(clk), .A(\g.we_clk [222]));
Q_ASSIGN U16169 ( .B(clk), .A(\g.we_clk [221]));
Q_ASSIGN U16170 ( .B(clk), .A(\g.we_clk [220]));
Q_ASSIGN U16171 ( .B(clk), .A(\g.we_clk [219]));
Q_ASSIGN U16172 ( .B(clk), .A(\g.we_clk [218]));
Q_ASSIGN U16173 ( .B(clk), .A(\g.we_clk [217]));
Q_ASSIGN U16174 ( .B(clk), .A(\g.we_clk [216]));
Q_ASSIGN U16175 ( .B(clk), .A(\g.we_clk [215]));
Q_ASSIGN U16176 ( .B(clk), .A(\g.we_clk [214]));
Q_ASSIGN U16177 ( .B(clk), .A(\g.we_clk [213]));
Q_ASSIGN U16178 ( .B(clk), .A(\g.we_clk [212]));
Q_ASSIGN U16179 ( .B(clk), .A(\g.we_clk [211]));
Q_ASSIGN U16180 ( .B(clk), .A(\g.we_clk [210]));
Q_ASSIGN U16181 ( .B(clk), .A(\g.we_clk [209]));
Q_ASSIGN U16182 ( .B(clk), .A(\g.we_clk [208]));
Q_ASSIGN U16183 ( .B(clk), .A(\g.we_clk [207]));
Q_ASSIGN U16184 ( .B(clk), .A(\g.we_clk [206]));
Q_ASSIGN U16185 ( .B(clk), .A(\g.we_clk [205]));
Q_ASSIGN U16186 ( .B(clk), .A(\g.we_clk [204]));
Q_ASSIGN U16187 ( .B(clk), .A(\g.we_clk [203]));
Q_ASSIGN U16188 ( .B(clk), .A(\g.we_clk [202]));
Q_ASSIGN U16189 ( .B(clk), .A(\g.we_clk [201]));
Q_ASSIGN U16190 ( .B(clk), .A(\g.we_clk [200]));
Q_ASSIGN U16191 ( .B(clk), .A(\g.we_clk [199]));
Q_ASSIGN U16192 ( .B(clk), .A(\g.we_clk [198]));
Q_ASSIGN U16193 ( .B(clk), .A(\g.we_clk [197]));
Q_ASSIGN U16194 ( .B(clk), .A(\g.we_clk [196]));
Q_ASSIGN U16195 ( .B(clk), .A(\g.we_clk [195]));
Q_ASSIGN U16196 ( .B(clk), .A(\g.we_clk [194]));
Q_ASSIGN U16197 ( .B(clk), .A(\g.we_clk [193]));
Q_ASSIGN U16198 ( .B(clk), .A(\g.we_clk [192]));
Q_ASSIGN U16199 ( .B(clk), .A(\g.we_clk [191]));
Q_ASSIGN U16200 ( .B(clk), .A(\g.we_clk [190]));
Q_ASSIGN U16201 ( .B(clk), .A(\g.we_clk [189]));
Q_ASSIGN U16202 ( .B(clk), .A(\g.we_clk [188]));
Q_ASSIGN U16203 ( .B(clk), .A(\g.we_clk [187]));
Q_ASSIGN U16204 ( .B(clk), .A(\g.we_clk [186]));
Q_ASSIGN U16205 ( .B(clk), .A(\g.we_clk [185]));
Q_ASSIGN U16206 ( .B(clk), .A(\g.we_clk [184]));
Q_ASSIGN U16207 ( .B(clk), .A(\g.we_clk [183]));
Q_ASSIGN U16208 ( .B(clk), .A(\g.we_clk [182]));
Q_ASSIGN U16209 ( .B(clk), .A(\g.we_clk [181]));
Q_ASSIGN U16210 ( .B(clk), .A(\g.we_clk [180]));
Q_ASSIGN U16211 ( .B(clk), .A(\g.we_clk [179]));
Q_ASSIGN U16212 ( .B(clk), .A(\g.we_clk [178]));
Q_ASSIGN U16213 ( .B(clk), .A(\g.we_clk [177]));
Q_ASSIGN U16214 ( .B(clk), .A(\g.we_clk [176]));
Q_ASSIGN U16215 ( .B(clk), .A(\g.we_clk [175]));
Q_ASSIGN U16216 ( .B(clk), .A(\g.we_clk [174]));
Q_ASSIGN U16217 ( .B(clk), .A(\g.we_clk [173]));
Q_ASSIGN U16218 ( .B(clk), .A(\g.we_clk [172]));
Q_ASSIGN U16219 ( .B(clk), .A(\g.we_clk [171]));
Q_ASSIGN U16220 ( .B(clk), .A(\g.we_clk [170]));
Q_ASSIGN U16221 ( .B(clk), .A(\g.we_clk [169]));
Q_ASSIGN U16222 ( .B(clk), .A(\g.we_clk [168]));
Q_ASSIGN U16223 ( .B(clk), .A(\g.we_clk [167]));
Q_ASSIGN U16224 ( .B(clk), .A(\g.we_clk [166]));
Q_ASSIGN U16225 ( .B(clk), .A(\g.we_clk [165]));
Q_ASSIGN U16226 ( .B(clk), .A(\g.we_clk [164]));
Q_ASSIGN U16227 ( .B(clk), .A(\g.we_clk [163]));
Q_ASSIGN U16228 ( .B(clk), .A(\g.we_clk [162]));
Q_ASSIGN U16229 ( .B(clk), .A(\g.we_clk [161]));
Q_ASSIGN U16230 ( .B(clk), .A(\g.we_clk [160]));
Q_ASSIGN U16231 ( .B(clk), .A(\g.we_clk [159]));
Q_ASSIGN U16232 ( .B(clk), .A(\g.we_clk [158]));
Q_ASSIGN U16233 ( .B(clk), .A(\g.we_clk [157]));
Q_ASSIGN U16234 ( .B(clk), .A(\g.we_clk [156]));
Q_ASSIGN U16235 ( .B(clk), .A(\g.we_clk [155]));
Q_ASSIGN U16236 ( .B(clk), .A(\g.we_clk [154]));
Q_ASSIGN U16237 ( .B(clk), .A(\g.we_clk [153]));
Q_ASSIGN U16238 ( .B(clk), .A(\g.we_clk [152]));
Q_ASSIGN U16239 ( .B(clk), .A(\g.we_clk [151]));
Q_ASSIGN U16240 ( .B(clk), .A(\g.we_clk [150]));
Q_ASSIGN U16241 ( .B(clk), .A(\g.we_clk [149]));
Q_ASSIGN U16242 ( .B(clk), .A(\g.we_clk [148]));
Q_ASSIGN U16243 ( .B(clk), .A(\g.we_clk [147]));
Q_ASSIGN U16244 ( .B(clk), .A(\g.we_clk [146]));
Q_ASSIGN U16245 ( .B(clk), .A(\g.we_clk [145]));
Q_ASSIGN U16246 ( .B(clk), .A(\g.we_clk [144]));
Q_ASSIGN U16247 ( .B(clk), .A(\g.we_clk [143]));
Q_ASSIGN U16248 ( .B(clk), .A(\g.we_clk [142]));
Q_ASSIGN U16249 ( .B(clk), .A(\g.we_clk [141]));
Q_ASSIGN U16250 ( .B(clk), .A(\g.we_clk [140]));
Q_ASSIGN U16251 ( .B(clk), .A(\g.we_clk [139]));
Q_ASSIGN U16252 ( .B(clk), .A(\g.we_clk [138]));
Q_ASSIGN U16253 ( .B(clk), .A(\g.we_clk [137]));
Q_ASSIGN U16254 ( .B(clk), .A(\g.we_clk [136]));
Q_ASSIGN U16255 ( .B(clk), .A(\g.we_clk [135]));
Q_ASSIGN U16256 ( .B(clk), .A(\g.we_clk [134]));
Q_ASSIGN U16257 ( .B(clk), .A(\g.we_clk [133]));
Q_ASSIGN U16258 ( .B(clk), .A(\g.we_clk [132]));
Q_ASSIGN U16259 ( .B(clk), .A(\g.we_clk [131]));
Q_ASSIGN U16260 ( .B(clk), .A(\g.we_clk [130]));
Q_ASSIGN U16261 ( .B(clk), .A(\g.we_clk [129]));
Q_ASSIGN U16262 ( .B(clk), .A(\g.we_clk [128]));
Q_ASSIGN U16263 ( .B(clk), .A(\g.we_clk [127]));
Q_ASSIGN U16264 ( .B(clk), .A(\g.we_clk [126]));
Q_ASSIGN U16265 ( .B(clk), .A(\g.we_clk [125]));
Q_ASSIGN U16266 ( .B(clk), .A(\g.we_clk [124]));
Q_ASSIGN U16267 ( .B(clk), .A(\g.we_clk [123]));
Q_ASSIGN U16268 ( .B(clk), .A(\g.we_clk [122]));
Q_ASSIGN U16269 ( .B(clk), .A(\g.we_clk [121]));
Q_ASSIGN U16270 ( .B(clk), .A(\g.we_clk [120]));
Q_ASSIGN U16271 ( .B(clk), .A(\g.we_clk [119]));
Q_ASSIGN U16272 ( .B(clk), .A(\g.we_clk [118]));
Q_ASSIGN U16273 ( .B(clk), .A(\g.we_clk [117]));
Q_ASSIGN U16274 ( .B(clk), .A(\g.we_clk [116]));
Q_ASSIGN U16275 ( .B(clk), .A(\g.we_clk [115]));
Q_ASSIGN U16276 ( .B(clk), .A(\g.we_clk [114]));
Q_ASSIGN U16277 ( .B(clk), .A(\g.we_clk [113]));
Q_ASSIGN U16278 ( .B(clk), .A(\g.we_clk [112]));
Q_ASSIGN U16279 ( .B(clk), .A(\g.we_clk [111]));
Q_ASSIGN U16280 ( .B(clk), .A(\g.we_clk [110]));
Q_ASSIGN U16281 ( .B(clk), .A(\g.we_clk [109]));
Q_ASSIGN U16282 ( .B(clk), .A(\g.we_clk [108]));
Q_ASSIGN U16283 ( .B(clk), .A(\g.we_clk [107]));
Q_ASSIGN U16284 ( .B(clk), .A(\g.we_clk [106]));
Q_ASSIGN U16285 ( .B(clk), .A(\g.we_clk [105]));
Q_ASSIGN U16286 ( .B(clk), .A(\g.we_clk [104]));
Q_ASSIGN U16287 ( .B(clk), .A(\g.we_clk [103]));
Q_ASSIGN U16288 ( .B(clk), .A(\g.we_clk [102]));
Q_ASSIGN U16289 ( .B(clk), .A(\g.we_clk [101]));
Q_ASSIGN U16290 ( .B(clk), .A(\g.we_clk [100]));
Q_ASSIGN U16291 ( .B(clk), .A(\g.we_clk [99]));
Q_ASSIGN U16292 ( .B(clk), .A(\g.we_clk [98]));
Q_ASSIGN U16293 ( .B(clk), .A(\g.we_clk [97]));
Q_ASSIGN U16294 ( .B(clk), .A(\g.we_clk [96]));
Q_ASSIGN U16295 ( .B(clk), .A(\g.we_clk [95]));
Q_ASSIGN U16296 ( .B(clk), .A(\g.we_clk [94]));
Q_ASSIGN U16297 ( .B(clk), .A(\g.we_clk [93]));
Q_ASSIGN U16298 ( .B(clk), .A(\g.we_clk [92]));
Q_ASSIGN U16299 ( .B(clk), .A(\g.we_clk [91]));
Q_ASSIGN U16300 ( .B(clk), .A(\g.we_clk [90]));
Q_ASSIGN U16301 ( .B(clk), .A(\g.we_clk [89]));
Q_ASSIGN U16302 ( .B(clk), .A(\g.we_clk [88]));
Q_ASSIGN U16303 ( .B(clk), .A(\g.we_clk [87]));
Q_ASSIGN U16304 ( .B(clk), .A(\g.we_clk [86]));
Q_ASSIGN U16305 ( .B(clk), .A(\g.we_clk [85]));
Q_ASSIGN U16306 ( .B(clk), .A(\g.we_clk [84]));
Q_ASSIGN U16307 ( .B(clk), .A(\g.we_clk [83]));
Q_ASSIGN U16308 ( .B(clk), .A(\g.we_clk [82]));
Q_ASSIGN U16309 ( .B(clk), .A(\g.we_clk [81]));
Q_ASSIGN U16310 ( .B(clk), .A(\g.we_clk [80]));
Q_ASSIGN U16311 ( .B(clk), .A(\g.we_clk [79]));
Q_ASSIGN U16312 ( .B(clk), .A(\g.we_clk [78]));
Q_ASSIGN U16313 ( .B(clk), .A(\g.we_clk [77]));
Q_ASSIGN U16314 ( .B(clk), .A(\g.we_clk [76]));
Q_ASSIGN U16315 ( .B(clk), .A(\g.we_clk [75]));
Q_ASSIGN U16316 ( .B(clk), .A(\g.we_clk [74]));
Q_ASSIGN U16317 ( .B(clk), .A(\g.we_clk [73]));
Q_ASSIGN U16318 ( .B(clk), .A(\g.we_clk [72]));
Q_ASSIGN U16319 ( .B(clk), .A(\g.we_clk [71]));
Q_ASSIGN U16320 ( .B(clk), .A(\g.we_clk [70]));
Q_ASSIGN U16321 ( .B(clk), .A(\g.we_clk [69]));
Q_ASSIGN U16322 ( .B(clk), .A(\g.we_clk [68]));
Q_ASSIGN U16323 ( .B(clk), .A(\g.we_clk [67]));
Q_ASSIGN U16324 ( .B(clk), .A(\g.we_clk [66]));
Q_ASSIGN U16325 ( .B(clk), .A(\g.we_clk [65]));
Q_ASSIGN U16326 ( .B(clk), .A(\g.we_clk [64]));
Q_ASSIGN U16327 ( .B(clk), .A(\g.we_clk [63]));
Q_ASSIGN U16328 ( .B(clk), .A(\g.we_clk [62]));
Q_ASSIGN U16329 ( .B(clk), .A(\g.we_clk [61]));
Q_ASSIGN U16330 ( .B(clk), .A(\g.we_clk [60]));
Q_ASSIGN U16331 ( .B(clk), .A(\g.we_clk [59]));
Q_ASSIGN U16332 ( .B(clk), .A(\g.we_clk [58]));
Q_ASSIGN U16333 ( .B(clk), .A(\g.we_clk [57]));
Q_ASSIGN U16334 ( .B(clk), .A(\g.we_clk [56]));
Q_ASSIGN U16335 ( .B(clk), .A(\g.we_clk [55]));
Q_ASSIGN U16336 ( .B(clk), .A(\g.we_clk [54]));
Q_ASSIGN U16337 ( .B(clk), .A(\g.we_clk [53]));
Q_ASSIGN U16338 ( .B(clk), .A(\g.we_clk [52]));
Q_ASSIGN U16339 ( .B(clk), .A(\g.we_clk [51]));
Q_ASSIGN U16340 ( .B(clk), .A(\g.we_clk [50]));
Q_ASSIGN U16341 ( .B(clk), .A(\g.we_clk [49]));
Q_ASSIGN U16342 ( .B(clk), .A(\g.we_clk [48]));
Q_ASSIGN U16343 ( .B(clk), .A(\g.we_clk [47]));
Q_ASSIGN U16344 ( .B(clk), .A(\g.we_clk [46]));
Q_ASSIGN U16345 ( .B(clk), .A(\g.we_clk [45]));
Q_ASSIGN U16346 ( .B(clk), .A(\g.we_clk [44]));
Q_ASSIGN U16347 ( .B(clk), .A(\g.we_clk [43]));
Q_ASSIGN U16348 ( .B(clk), .A(\g.we_clk [42]));
Q_ASSIGN U16349 ( .B(clk), .A(\g.we_clk [41]));
Q_ASSIGN U16350 ( .B(clk), .A(\g.we_clk [40]));
Q_ASSIGN U16351 ( .B(clk), .A(\g.we_clk [39]));
Q_ASSIGN U16352 ( .B(clk), .A(\g.we_clk [38]));
Q_ASSIGN U16353 ( .B(clk), .A(\g.we_clk [37]));
Q_ASSIGN U16354 ( .B(clk), .A(\g.we_clk [36]));
Q_ASSIGN U16355 ( .B(clk), .A(\g.we_clk [35]));
Q_ASSIGN U16356 ( .B(clk), .A(\g.we_clk [34]));
Q_ASSIGN U16357 ( .B(clk), .A(\g.we_clk [33]));
Q_ASSIGN U16358 ( .B(clk), .A(\g.we_clk [32]));
Q_ASSIGN U16359 ( .B(clk), .A(\g.we_clk [31]));
Q_ASSIGN U16360 ( .B(clk), .A(\g.we_clk [30]));
Q_ASSIGN U16361 ( .B(clk), .A(\g.we_clk [29]));
Q_ASSIGN U16362 ( .B(clk), .A(\g.we_clk [28]));
Q_ASSIGN U16363 ( .B(clk), .A(\g.we_clk [27]));
Q_ASSIGN U16364 ( .B(clk), .A(\g.we_clk [26]));
Q_ASSIGN U16365 ( .B(clk), .A(\g.we_clk [25]));
Q_ASSIGN U16366 ( .B(clk), .A(\g.we_clk [24]));
Q_ASSIGN U16367 ( .B(clk), .A(\g.we_clk [23]));
Q_ASSIGN U16368 ( .B(clk), .A(\g.we_clk [22]));
Q_ASSIGN U16369 ( .B(clk), .A(\g.we_clk [21]));
Q_ASSIGN U16370 ( .B(clk), .A(\g.we_clk [20]));
Q_ASSIGN U16371 ( .B(clk), .A(\g.we_clk [19]));
Q_ASSIGN U16372 ( .B(clk), .A(\g.we_clk [18]));
Q_ASSIGN U16373 ( .B(clk), .A(\g.we_clk [17]));
Q_ASSIGN U16374 ( .B(clk), .A(\g.we_clk [16]));
Q_ASSIGN U16375 ( .B(clk), .A(\g.we_clk [15]));
Q_ASSIGN U16376 ( .B(clk), .A(\g.we_clk [14]));
Q_ASSIGN U16377 ( .B(clk), .A(\g.we_clk [13]));
Q_ASSIGN U16378 ( .B(clk), .A(\g.we_clk [12]));
Q_ASSIGN U16379 ( .B(clk), .A(\g.we_clk [11]));
Q_ASSIGN U16380 ( .B(clk), .A(\g.we_clk [10]));
Q_ASSIGN U16381 ( .B(clk), .A(\g.we_clk [9]));
Q_ASSIGN U16382 ( .B(clk), .A(\g.we_clk [8]));
Q_ASSIGN U16383 ( .B(clk), .A(\g.we_clk [7]));
Q_ASSIGN U16384 ( .B(clk), .A(\g.we_clk [6]));
Q_ASSIGN U16385 ( .B(clk), .A(\g.we_clk [5]));
Q_ASSIGN U16386 ( .B(clk), .A(\g.we_clk [4]));
Q_ASSIGN U16387 ( .B(clk), .A(\g.we_clk [3]));
Q_ASSIGN U16388 ( .B(clk), .A(\g.we_clk [2]));
Q_ASSIGN U16389 ( .B(clk), .A(\g.we_clk [1]));
Q_ASSIGN U16390 ( .B(clk), .A(\g.we_clk [0]));
Q_BUF U16391 ( .A(n138), .Z(ro_uncorrectable_ecc_error));
ixc_assign _zz_strnp_10 ( _zy_simnet_ro_uncorrectable_ecc_error_2_w$, n138);
ixc_assign _zz_strnp_9 ( _zy_simnet_bimc_osync_1_w$, bimc_osync);
ixc_assign _zz_strnp_8 ( _zy_simnet_bimc_odat_0_w$, bimc_odat);
Q_INV U16395 ( .A(n137), .Z(web));
Q_AN02 U16396 ( .A0(cs), .A1(we), .Z(n137));
ixc_assign _zz_strnp_7 ( rst_rclk_n, rst_n);
ixc_assign _zz_strnp_6 ( rst_clk_n, rst_n);
ixc_assign _zz_strnp_5 ( bimc_irstn, bimc_rst_n);
ixc_assign _zz_strnp_4 ( bimc_iclk, clk);
Q_FDP0 U16401 ( .CK(clk), .D(\g.din_i [37]), .Q(n136), .QN( ));
Q_FDP0 U16402 ( .CK(clk), .D(\g.din_i [36]), .Q(n135), .QN( ));
Q_FDP0 U16403 ( .CK(clk), .D(\g.din_i [35]), .Q(n134), .QN( ));
Q_FDP0 U16404 ( .CK(clk), .D(\g.din_i [34]), .Q(n133), .QN( ));
Q_FDP0 U16405 ( .CK(clk), .D(\g.din_i [33]), .Q(n132), .QN( ));
Q_FDP0 U16406 ( .CK(clk), .D(\g.din_i [32]), .Q(n131), .QN( ));
Q_FDP0 U16407 ( .CK(clk), .D(\g.din_i [31]), .Q(n130), .QN( ));
Q_FDP0 U16408 ( .CK(clk), .D(\g.din_i [30]), .Q(n129), .QN( ));
Q_FDP0 U16409 ( .CK(clk), .D(\g.din_i [29]), .Q(n128), .QN( ));
Q_FDP0 U16410 ( .CK(clk), .D(\g.din_i [28]), .Q(n127), .QN( ));
Q_FDP0 U16411 ( .CK(clk), .D(\g.din_i [27]), .Q(n126), .QN( ));
Q_FDP0 U16412 ( .CK(clk), .D(\g.din_i [26]), .Q(n125), .QN( ));
Q_FDP0 U16413 ( .CK(clk), .D(\g.din_i [25]), .Q(n124), .QN( ));
Q_FDP0 U16414 ( .CK(clk), .D(\g.din_i [24]), .Q(n123), .QN( ));
Q_FDP0 U16415 ( .CK(clk), .D(\g.din_i [23]), .Q(n122), .QN( ));
Q_FDP0 U16416 ( .CK(clk), .D(\g.din_i [22]), .Q(n121), .QN( ));
Q_FDP0 U16417 ( .CK(clk), .D(\g.din_i [21]), .Q(n120), .QN( ));
Q_FDP0 U16418 ( .CK(clk), .D(\g.din_i [20]), .Q(n119), .QN( ));
Q_FDP0 U16419 ( .CK(clk), .D(\g.din_i [19]), .Q(n118), .QN( ));
Q_FDP0 U16420 ( .CK(clk), .D(\g.din_i [18]), .Q(n117), .QN( ));
Q_FDP0 U16421 ( .CK(clk), .D(\g.din_i [17]), .Q(n116), .QN( ));
Q_FDP0 U16422 ( .CK(clk), .D(\g.din_i [16]), .Q(n115), .QN( ));
Q_FDP0 U16423 ( .CK(clk), .D(\g.din_i [15]), .Q(n114), .QN( ));
Q_FDP0 U16424 ( .CK(clk), .D(\g.din_i [14]), .Q(n113), .QN( ));
Q_FDP0 U16425 ( .CK(clk), .D(\g.din_i [13]), .Q(n112), .QN( ));
Q_FDP0 U16426 ( .CK(clk), .D(\g.din_i [12]), .Q(n111), .QN( ));
Q_FDP0 U16427 ( .CK(clk), .D(\g.din_i [11]), .Q(n110), .QN( ));
Q_FDP0 U16428 ( .CK(clk), .D(\g.din_i [10]), .Q(n109), .QN( ));
Q_FDP0 U16429 ( .CK(clk), .D(\g.din_i [9]), .Q(n108), .QN( ));
Q_FDP0 U16430 ( .CK(clk), .D(\g.din_i [8]), .Q(n107), .QN( ));
Q_FDP0 U16431 ( .CK(clk), .D(\g.din_i [7]), .Q(n106), .QN( ));
Q_FDP0 U16432 ( .CK(clk), .D(\g.din_i [6]), .Q(n105), .QN( ));
Q_FDP0 U16433 ( .CK(clk), .D(\g.din_i [5]), .Q(n104), .QN( ));
Q_FDP0 U16434 ( .CK(clk), .D(\g.din_i [4]), .Q(n103), .QN( ));
Q_FDP0 U16435 ( .CK(clk), .D(\g.din_i [3]), .Q(n102), .QN( ));
Q_FDP0 U16436 ( .CK(clk), .D(\g.din_i [2]), .Q(n101), .QN( ));
Q_FDP0 U16437 ( .CK(clk), .D(\g.din_i [1]), .Q(n100), .QN( ));
Q_FDP0 U16438 ( .CK(clk), .D(\g.din_i [0]), .Q(n99), .QN( ));
Q_FDP0 U16439 ( .CK(clk), .D(add[13]), .Q(n98), .QN( ));
Q_FDP0 U16440 ( .CK(clk), .D(add[12]), .Q(n97), .QN( ));
Q_FDP0 U16441 ( .CK(clk), .D(add[11]), .Q(n96), .QN( ));
Q_FDP0 U16442 ( .CK(clk), .D(add[10]), .Q(n95), .QN( ));
Q_FDP0 U16443 ( .CK(clk), .D(add[9]), .Q(n94), .QN( ));
Q_FDP0 U16444 ( .CK(clk), .D(add[8]), .Q(n93), .QN( ));
Q_FDP0 U16445 ( .CK(clk), .D(add[7]), .Q(n92), .QN( ));
Q_FDP0 U16446 ( .CK(clk), .D(add[6]), .Q(n91), .QN( ));
Q_FDP0 U16447 ( .CK(clk), .D(add[5]), .Q(n90), .QN( ));
Q_FDP0 U16448 ( .CK(clk), .D(add[4]), .Q(n89), .QN( ));
Q_FDP0 U16449 ( .CK(clk), .D(add[3]), .Q(n88), .QN( ));
Q_FDP0 U16450 ( .CK(clk), .D(add[2]), .Q(n87), .QN( ));
Q_FDP0 U16451 ( .CK(clk), .D(add[1]), .Q(n86), .QN( ));
Q_FDP0 U16452 ( .CK(clk), .D(add[0]), .Q(n85), .QN( ));
Q_AN02 U16453 ( .A0(n80), .A1(n83), .Z(n84));
Q_XOR2 U16454 ( .A0(n79), .A1(n82), .Z(n83));
// pragma CVAINTPROP NET n79 _2_state_ 1
// pragma CVAINTPROP INSTANCE U16454 NOBREAKS 1
Q_FDP0B U16455 ( .D(n79), .QTFCLK( ), .Q(n82));
Q_FDP0 U16456 ( .CK(clk), .D(n137), .Q(n80), .QN( ));
Q_FDP0 U16457 ( .CK(clk), .D(n81), .Q(n79), .QN(n81));
Q_MX02 U16458 ( .S(we), .A0(\g.dout_i [37]), .A1(\g.din_i [37]), .Z(n78));
Q_MX02 U16459 ( .S(we), .A0(\g.dout_i [36]), .A1(\g.din_i [36]), .Z(n77));
Q_MX02 U16460 ( .S(we), .A0(\g.dout_i [35]), .A1(\g.din_i [35]), .Z(n76));
Q_MX02 U16461 ( .S(we), .A0(\g.dout_i [34]), .A1(\g.din_i [34]), .Z(n75));
Q_MX02 U16462 ( .S(we), .A0(\g.dout_i [33]), .A1(\g.din_i [33]), .Z(n74));
Q_MX02 U16463 ( .S(we), .A0(\g.dout_i [32]), .A1(\g.din_i [32]), .Z(n73));
Q_MX02 U16464 ( .S(we), .A0(\g.dout_i [31]), .A1(\g.din_i [31]), .Z(n72));
Q_MX02 U16465 ( .S(we), .A0(\g.dout_i [30]), .A1(\g.din_i [30]), .Z(n71));
Q_MX02 U16466 ( .S(we), .A0(\g.dout_i [29]), .A1(\g.din_i [29]), .Z(n70));
Q_MX02 U16467 ( .S(we), .A0(\g.dout_i [28]), .A1(\g.din_i [28]), .Z(n69));
Q_MX02 U16468 ( .S(we), .A0(\g.dout_i [27]), .A1(\g.din_i [27]), .Z(n68));
Q_MX02 U16469 ( .S(we), .A0(\g.dout_i [26]), .A1(\g.din_i [26]), .Z(n67));
Q_MX02 U16470 ( .S(we), .A0(\g.dout_i [25]), .A1(\g.din_i [25]), .Z(n66));
Q_MX02 U16471 ( .S(we), .A0(\g.dout_i [24]), .A1(\g.din_i [24]), .Z(n65));
Q_MX02 U16472 ( .S(we), .A0(\g.dout_i [23]), .A1(\g.din_i [23]), .Z(n64));
Q_MX02 U16473 ( .S(we), .A0(\g.dout_i [22]), .A1(\g.din_i [22]), .Z(n63));
Q_MX02 U16474 ( .S(we), .A0(\g.dout_i [21]), .A1(\g.din_i [21]), .Z(n62));
Q_MX02 U16475 ( .S(we), .A0(\g.dout_i [20]), .A1(\g.din_i [20]), .Z(n61));
Q_MX02 U16476 ( .S(we), .A0(\g.dout_i [19]), .A1(\g.din_i [19]), .Z(n60));
Q_MX02 U16477 ( .S(we), .A0(\g.dout_i [18]), .A1(\g.din_i [18]), .Z(n59));
Q_MX02 U16478 ( .S(we), .A0(\g.dout_i [17]), .A1(\g.din_i [17]), .Z(n58));
Q_MX02 U16479 ( .S(we), .A0(\g.dout_i [16]), .A1(\g.din_i [16]), .Z(n57));
Q_MX02 U16480 ( .S(we), .A0(\g.dout_i [15]), .A1(\g.din_i [15]), .Z(n56));
Q_MX02 U16481 ( .S(we), .A0(\g.dout_i [14]), .A1(\g.din_i [14]), .Z(n55));
Q_MX02 U16482 ( .S(we), .A0(\g.dout_i [13]), .A1(\g.din_i [13]), .Z(n54));
Q_MX02 U16483 ( .S(we), .A0(\g.dout_i [12]), .A1(\g.din_i [12]), .Z(n53));
Q_MX02 U16484 ( .S(we), .A0(\g.dout_i [11]), .A1(\g.din_i [11]), .Z(n52));
Q_MX02 U16485 ( .S(we), .A0(\g.dout_i [10]), .A1(\g.din_i [10]), .Z(n51));
Q_MX02 U16486 ( .S(we), .A0(\g.dout_i [9]), .A1(\g.din_i [9]), .Z(n50));
Q_MX02 U16487 ( .S(we), .A0(\g.dout_i [8]), .A1(\g.din_i [8]), .Z(n49));
Q_MX02 U16488 ( .S(we), .A0(\g.dout_i [7]), .A1(\g.din_i [7]), .Z(n48));
Q_MX02 U16489 ( .S(we), .A0(\g.dout_i [6]), .A1(\g.din_i [6]), .Z(n47));
Q_MX02 U16490 ( .S(we), .A0(\g.dout_i [5]), .A1(\g.din_i [5]), .Z(n46));
Q_MX02 U16491 ( .S(we), .A0(\g.dout_i [4]), .A1(\g.din_i [4]), .Z(n45));
Q_MX02 U16492 ( .S(we), .A0(\g.dout_i [3]), .A1(\g.din_i [3]), .Z(n44));
Q_MX02 U16493 ( .S(we), .A0(\g.dout_i [2]), .A1(\g.din_i [2]), .Z(n43));
Q_MX02 U16494 ( .S(we), .A0(\g.dout_i [1]), .A1(\g.din_i [1]), .Z(n42));
Q_MX02 U16495 ( .S(we), .A0(\g.dout_i [0]), .A1(\g.din_i [0]), .Z(n41));
ixc_assign_38 \g._zz_strnp_0 ( \g.dout_i [37:0], { n40, n39, n38, n37, n36, 
	n35, n34, n33, n32, n31, n30, n29, n28, n27, n26, n25, n24, n23, n22, 
	n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10, n9, n8, 
	n7, n6, n5, n4, n3});
ixc_assign \g._zz_strnp_3 ( bimc_osync, bimc_isync);
ixc_assign \g._zz_strnp_2 ( bimc_odat, bimc_idat);
ixc_assign_38 \g._zz_strnp_1 ( dout[37:0], \g.dat_r [37:0]);
Q_MX02 U16500 ( .S(bwe[37]), .A0(\g.dout_i [37]), .A1(din[37]), .Z(\g.din_i [37]));
Q_MX02 U16501 ( .S(bwe[36]), .A0(\g.dout_i [36]), .A1(din[36]), .Z(\g.din_i [36]));
Q_MX02 U16502 ( .S(bwe[35]), .A0(\g.dout_i [35]), .A1(din[35]), .Z(\g.din_i [35]));
Q_MX02 U16503 ( .S(bwe[34]), .A0(\g.dout_i [34]), .A1(din[34]), .Z(\g.din_i [34]));
Q_MX02 U16504 ( .S(bwe[33]), .A0(\g.dout_i [33]), .A1(din[33]), .Z(\g.din_i [33]));
Q_MX02 U16505 ( .S(bwe[32]), .A0(\g.dout_i [32]), .A1(din[32]), .Z(\g.din_i [32]));
Q_MX02 U16506 ( .S(bwe[31]), .A0(\g.dout_i [31]), .A1(din[31]), .Z(\g.din_i [31]));
Q_MX02 U16507 ( .S(bwe[30]), .A0(\g.dout_i [30]), .A1(din[30]), .Z(\g.din_i [30]));
Q_MX02 U16508 ( .S(bwe[29]), .A0(\g.dout_i [29]), .A1(din[29]), .Z(\g.din_i [29]));
Q_MX02 U16509 ( .S(bwe[28]), .A0(\g.dout_i [28]), .A1(din[28]), .Z(\g.din_i [28]));
Q_MX02 U16510 ( .S(bwe[27]), .A0(\g.dout_i [27]), .A1(din[27]), .Z(\g.din_i [27]));
Q_MX02 U16511 ( .S(bwe[26]), .A0(\g.dout_i [26]), .A1(din[26]), .Z(\g.din_i [26]));
Q_MX02 U16512 ( .S(bwe[25]), .A0(\g.dout_i [25]), .A1(din[25]), .Z(\g.din_i [25]));
Q_MX02 U16513 ( .S(bwe[24]), .A0(\g.dout_i [24]), .A1(din[24]), .Z(\g.din_i [24]));
Q_MX02 U16514 ( .S(bwe[23]), .A0(\g.dout_i [23]), .A1(din[23]), .Z(\g.din_i [23]));
Q_MX02 U16515 ( .S(bwe[22]), .A0(\g.dout_i [22]), .A1(din[22]), .Z(\g.din_i [22]));
Q_MX02 U16516 ( .S(bwe[21]), .A0(\g.dout_i [21]), .A1(din[21]), .Z(\g.din_i [21]));
Q_MX02 U16517 ( .S(bwe[20]), .A0(\g.dout_i [20]), .A1(din[20]), .Z(\g.din_i [20]));
Q_MX02 U16518 ( .S(bwe[19]), .A0(\g.dout_i [19]), .A1(din[19]), .Z(\g.din_i [19]));
Q_MX02 U16519 ( .S(bwe[18]), .A0(\g.dout_i [18]), .A1(din[18]), .Z(\g.din_i [18]));
Q_MX02 U16520 ( .S(bwe[17]), .A0(\g.dout_i [17]), .A1(din[17]), .Z(\g.din_i [17]));
Q_MX02 U16521 ( .S(bwe[16]), .A0(\g.dout_i [16]), .A1(din[16]), .Z(\g.din_i [16]));
Q_MX02 U16522 ( .S(bwe[15]), .A0(\g.dout_i [15]), .A1(din[15]), .Z(\g.din_i [15]));
Q_MX02 U16523 ( .S(bwe[14]), .A0(\g.dout_i [14]), .A1(din[14]), .Z(\g.din_i [14]));
Q_MX02 U16524 ( .S(bwe[13]), .A0(\g.dout_i [13]), .A1(din[13]), .Z(\g.din_i [13]));
Q_MX02 U16525 ( .S(bwe[12]), .A0(\g.dout_i [12]), .A1(din[12]), .Z(\g.din_i [12]));
Q_MX02 U16526 ( .S(bwe[11]), .A0(\g.dout_i [11]), .A1(din[11]), .Z(\g.din_i [11]));
Q_MX02 U16527 ( .S(bwe[10]), .A0(\g.dout_i [10]), .A1(din[10]), .Z(\g.din_i [10]));
Q_MX02 U16528 ( .S(bwe[9]), .A0(\g.dout_i [9]), .A1(din[9]), .Z(\g.din_i [9]));
Q_MX02 U16529 ( .S(bwe[8]), .A0(\g.dout_i [8]), .A1(din[8]), .Z(\g.din_i [8]));
Q_MX02 U16530 ( .S(bwe[7]), .A0(\g.dout_i [7]), .A1(din[7]), .Z(\g.din_i [7]));
Q_MX02 U16531 ( .S(bwe[6]), .A0(\g.dout_i [6]), .A1(din[6]), .Z(\g.din_i [6]));
Q_MX02 U16532 ( .S(bwe[5]), .A0(\g.dout_i [5]), .A1(din[5]), .Z(\g.din_i [5]));
Q_MX02 U16533 ( .S(bwe[4]), .A0(\g.dout_i [4]), .A1(din[4]), .Z(\g.din_i [4]));
Q_MX02 U16534 ( .S(bwe[3]), .A0(\g.dout_i [3]), .A1(din[3]), .Z(\g.din_i [3]));
Q_MX02 U16535 ( .S(bwe[2]), .A0(\g.dout_i [2]), .A1(din[2]), .Z(\g.din_i [2]));
Q_MX02 U16536 ( .S(bwe[1]), .A0(\g.dout_i [1]), .A1(din[1]), .Z(\g.din_i [1]));
Q_MX02 U16537 ( .S(bwe[0]), .A0(\g.dout_i [0]), .A1(din[0]), .Z(\g.din_i [0]));
Q_FDP4EP \g.dat_r_REG[37] ( .CK(clk), .CE(cs), .R(n1), .D(n78), .Q(\g.dat_r [37]));
Q_INV U16539 ( .A(rst_n), .Z(n1));
Q_FDP4EP \g.dat_r_REG[36] ( .CK(clk), .CE(cs), .R(n1), .D(n77), .Q(\g.dat_r [36]));
Q_FDP4EP \g.dat_r_REG[35] ( .CK(clk), .CE(cs), .R(n1), .D(n76), .Q(\g.dat_r [35]));
Q_FDP4EP \g.dat_r_REG[34] ( .CK(clk), .CE(cs), .R(n1), .D(n75), .Q(\g.dat_r [34]));
Q_FDP4EP \g.dat_r_REG[33] ( .CK(clk), .CE(cs), .R(n1), .D(n74), .Q(\g.dat_r [33]));
Q_FDP4EP \g.dat_r_REG[32] ( .CK(clk), .CE(cs), .R(n1), .D(n73), .Q(\g.dat_r [32]));
Q_FDP4EP \g.dat_r_REG[31] ( .CK(clk), .CE(cs), .R(n1), .D(n72), .Q(\g.dat_r [31]));
Q_FDP4EP \g.dat_r_REG[30] ( .CK(clk), .CE(cs), .R(n1), .D(n71), .Q(\g.dat_r [30]));
Q_FDP4EP \g.dat_r_REG[29] ( .CK(clk), .CE(cs), .R(n1), .D(n70), .Q(\g.dat_r [29]));
Q_FDP4EP \g.dat_r_REG[28] ( .CK(clk), .CE(cs), .R(n1), .D(n69), .Q(\g.dat_r [28]));
Q_FDP4EP \g.dat_r_REG[27] ( .CK(clk), .CE(cs), .R(n1), .D(n68), .Q(\g.dat_r [27]));
Q_FDP4EP \g.dat_r_REG[26] ( .CK(clk), .CE(cs), .R(n1), .D(n67), .Q(\g.dat_r [26]));
Q_FDP4EP \g.dat_r_REG[25] ( .CK(clk), .CE(cs), .R(n1), .D(n66), .Q(\g.dat_r [25]));
Q_FDP4EP \g.dat_r_REG[24] ( .CK(clk), .CE(cs), .R(n1), .D(n65), .Q(\g.dat_r [24]));
Q_FDP4EP \g.dat_r_REG[23] ( .CK(clk), .CE(cs), .R(n1), .D(n64), .Q(\g.dat_r [23]));
Q_FDP4EP \g.dat_r_REG[22] ( .CK(clk), .CE(cs), .R(n1), .D(n63), .Q(\g.dat_r [22]));
Q_FDP4EP \g.dat_r_REG[21] ( .CK(clk), .CE(cs), .R(n1), .D(n62), .Q(\g.dat_r [21]));
Q_FDP4EP \g.dat_r_REG[20] ( .CK(clk), .CE(cs), .R(n1), .D(n61), .Q(\g.dat_r [20]));
Q_FDP4EP \g.dat_r_REG[19] ( .CK(clk), .CE(cs), .R(n1), .D(n60), .Q(\g.dat_r [19]));
Q_FDP4EP \g.dat_r_REG[18] ( .CK(clk), .CE(cs), .R(n1), .D(n59), .Q(\g.dat_r [18]));
Q_FDP4EP \g.dat_r_REG[17] ( .CK(clk), .CE(cs), .R(n1), .D(n58), .Q(\g.dat_r [17]));
Q_FDP4EP \g.dat_r_REG[16] ( .CK(clk), .CE(cs), .R(n1), .D(n57), .Q(\g.dat_r [16]));
Q_FDP4EP \g.dat_r_REG[15] ( .CK(clk), .CE(cs), .R(n1), .D(n56), .Q(\g.dat_r [15]));
Q_FDP4EP \g.dat_r_REG[14] ( .CK(clk), .CE(cs), .R(n1), .D(n55), .Q(\g.dat_r [14]));
Q_FDP4EP \g.dat_r_REG[13] ( .CK(clk), .CE(cs), .R(n1), .D(n54), .Q(\g.dat_r [13]));
Q_FDP4EP \g.dat_r_REG[12] ( .CK(clk), .CE(cs), .R(n1), .D(n53), .Q(\g.dat_r [12]));
Q_FDP4EP \g.dat_r_REG[11] ( .CK(clk), .CE(cs), .R(n1), .D(n52), .Q(\g.dat_r [11]));
Q_FDP4EP \g.dat_r_REG[10] ( .CK(clk), .CE(cs), .R(n1), .D(n51), .Q(\g.dat_r [10]));
Q_FDP4EP \g.dat_r_REG[9] ( .CK(clk), .CE(cs), .R(n1), .D(n50), .Q(\g.dat_r [9]));
Q_FDP4EP \g.dat_r_REG[8] ( .CK(clk), .CE(cs), .R(n1), .D(n49), .Q(\g.dat_r [8]));
Q_FDP4EP \g.dat_r_REG[7] ( .CK(clk), .CE(cs), .R(n1), .D(n48), .Q(\g.dat_r [7]));
Q_FDP4EP \g.dat_r_REG[6] ( .CK(clk), .CE(cs), .R(n1), .D(n47), .Q(\g.dat_r [6]));
Q_FDP4EP \g.dat_r_REG[5] ( .CK(clk), .CE(cs), .R(n1), .D(n46), .Q(\g.dat_r [5]));
Q_FDP4EP \g.dat_r_REG[4] ( .CK(clk), .CE(cs), .R(n1), .D(n45), .Q(\g.dat_r [4]));
Q_FDP4EP \g.dat_r_REG[3] ( .CK(clk), .CE(cs), .R(n1), .D(n44), .Q(\g.dat_r [3]));
Q_FDP4EP \g.dat_r_REG[2] ( .CK(clk), .CE(cs), .R(n1), .D(n43), .Q(\g.dat_r [2]));
Q_FDP4EP \g.dat_r_REG[1] ( .CK(clk), .CE(cs), .R(n1), .D(n42), .Q(\g.dat_r [1]));
Q_FDP4EP \g.dat_r_REG[0] ( .CK(clk), .CE(cs), .R(n1), .D(n41), .Q(\g.dat_r [0]));
`ifdef CBV

reg [37:0] \g.mem  [0:16383];
initial begin: U16577
  integer i;
  for (i=0; i<=16383; i=i+1) \g.mem [i] =
`ifdef CBV_MEM_INIT1
  {38{1'b1}};
`else
  38'b0;
`endif
end
reg [37:0] n139;
assign {n40, n39, n38, n37, n36, n35, n34,
n33, n32, n31, n30, n29, n28, n27, n26,
n25, n24, n23, n22, n21, n20, n19, n18,
n17, n16, n15, n14, n13, n12, n11, n10,
n9, n8, n7, n6, n5, n4, n3} = n139; 
always @(n98 or n97 or n96 or n95 or n94
 or n93 or n92 or n91 or n90 or n89 or n88 or n87 or n86
 or n85 or n136 or n135 or n134 or n133 or n132 or n131 or n130
 or n129 or n128 or n127 or n126 or n125 or n124 or n123 or n122
 or n121 or n120 or n119 or n118 or n117 or n116 or n115 or n114
 or n113 or n112 or n111 or n110 or n109 or n108 or n107 or n106
 or n105 or n104 or n103 or n102 or n101 or n100 or n99 or n84
 or add[13] or add[12] or add[11] or add[10] or add[9] or add[8] or add[7] or add[6]
 or add[5] or add[4] or add[3] or add[2] or add[1] or add[0])
#0 begin
if (n84)
\g.mem [{n98, n97, n96, n95, n94,
 n93, n92, n91, n90, n89, n88, n87, n86,
 n85}] =
{n136, n135, n134, n133, n132,
 n131, n130, n129, n128, n127, n126, n125, n124,
 n123, n122, n121, n120, n119, n118, n117, n116,
 n115, n114, n113, n112, n111, n110, n109, n108,
 n107, n106, n105, n104, n103, n102, n101, n100,
 n99};
n139 = \g.mem [{add[13], add[12], add[11], add[10], add[9],
 add[8], add[7], add[6], add[5], add[4], add[3], add[2], add[1],
 add[0]}];
end
`else

MPW16KX38 \g.mem  ( .A13(n98), .A12(n97), .A11(n96), .A10(n95), .A9(n94), .A8(n93),
 .A7(n92), .A6(n91), .A5(n90), .A4(n89), .A3(n88), .A2(n87), .A1(n86), .A0(n85),
 .DI37(n136), .DI36(n135), .DI35(n134), .DI34(n133), .DI33(n132), .DI32(n131), .DI31(n130), .DI30(n129),
 .DI29(n128), .DI28(n127), .DI27(n126), .DI26(n125), .DI25(n124), .DI24(n123), .DI23(n122), .DI22(n121),
 .DI21(n120), .DI20(n119), .DI19(n118), .DI18(n117), .DI17(n116), .DI16(n115), .DI15(n114), .DI14(n113),
 .DI13(n112), .DI12(n111), .DI11(n110), .DI10(n109), .DI9(n108), .DI8(n107), .DI7(n106), .DI6(n105),
 .DI5(n104), .DI4(n103), .DI3(n102), .DI2(n101), .DI1(n100), .DI0(n99), .WE(n84), .SYNC_IN(n138),
 .SYNC_OUT(n139));
// pragma CVASTRPROP INSTANCE "\g.mem " HDL_MEMORY_DECL "1 37 0 0 16383"
MPR16KX38 U16578 ( .A13(add[13]), .A12(add[12]), .A11(add[11]), .A10(add[10]), .A9(add[9]), .A8(add[8]),
 .A7(add[7]), .A6(add[6]), .A5(add[5]), .A4(add[4]), .A3(add[3]), .A2(add[2]), .A1(add[1]), .A0(add[0]),
 .SYNC_IN(n139), .DO37(n40), .DO36(n39), .DO35(n38), .DO34(n37), .DO33(n36), .DO32(n35), .DO31(n34),
 .DO30(n33), .DO29(n32), .DO28(n31), .DO27(n30), .DO26(n29), .DO25(n28), .DO24(n27), .DO23(n26),
 .DO22(n25), .DO21(n24), .DO20(n23), .DO19(n22), .DO18(n21), .DO17(n20), .DO16(n19), .DO15(n18),
 .DO14(n17), .DO13(n16), .DO12(n15), .DO11(n14), .DO10(n13), .DO9(n12), .DO8(n11), .DO7(n10),
 .DO6(n9), .DO5(n8), .DO4(n7), .DO3(n6), .DO2(n5), .DO1(n4), .DO0(n3), .SYNC_OUT( ));
`endif
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_1 "0 u_ram  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate_0 "-1 g  "
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "g.u_ram"
// pragma CVASTRPROP MODULE HDLICE cva_for_generate "g"
endmodule
`ifdef CBV
`else
`ifdef MPW16KX38_MPR16KX38
`else
module MPW16KX38( A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, DI37,
 DI36, DI35, DI34, DI33, DI32, DI31, DI30, DI29,
 DI28, DI27, DI26, DI25, DI24, DI23, DI22, DI21,
 DI20, DI19, DI18, DI17, DI16, DI15, DI14, DI13,
 DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5,
 DI4, DI3, DI2, DI1, DI0, WE, SYNC_IN, SYNC_OUT);
input  A13, A12, A11, A10, A9, A8, A7, A6,
 A5, A4, A3, A2, A1, A0, DI37, DI36, DI35, DI34,
 DI33, DI32, DI31, DI30, DI29, DI28, DI27, DI26, DI25, DI24,
 DI23, DI22, DI21, DI20, DI19, DI18, DI17, DI16, DI15, DI14,
 DI13, DI12, DI11, DI10, DI9, DI8, DI7, DI6, DI5, DI4,
 DI3, DI2, DI1, DI0, WE, SYNC_IN;
output  SYNC_OUT;
endmodule
`ifdef _MPR16KX38_
`else
module MPR16KX38( A13, A12, A11, A10, A9, A8, A7,
 A6, A5, A4, A3, A2, A1, A0, SYNC_IN,
 DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30,
 DO29, DO28, DO27, DO26, DO25, DO24, DO23, DO22,
 DO21, DO20, DO19, DO18, DO17, DO16, DO15, DO14,
 DO13, DO12, DO11, DO10, DO9, DO8, DO7, DO6,
 DO5, DO4, DO3, DO2, DO1, DO0, SYNC_OUT);
input  A13, A12, A11, A10, A9, A8, A7, A6,
 A5, A4, A3, A2, A1, A0, SYNC_IN;
output  DO37, DO36, DO35, DO34, DO33, DO32, DO31, DO30,
 DO29, DO28, DO27, DO26, DO25, DO24, DO23, DO22, DO21, DO20,
 DO19, DO18, DO17, DO16, DO15, DO14, DO13, DO12, DO11, DO10,
 DO9, DO8, DO7, DO6, DO5, DO4, DO3, DO2, DO1, DO0,
 SYNC_OUT;
endmodule
`define _MPR16KX38_
`endif
`define MPW16KX38_MPR16KX38
`endif
`endif
